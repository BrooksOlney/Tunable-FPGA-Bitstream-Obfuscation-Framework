module sqrt_qmap_map (ax126x, ax127x, ax124x, ax125x, ax122x, ax123x, ax120x, ax121x, ax118x, ax119x, ax116x, ax117x, ax114x, ax115x, ax112x, ax113x, ax110x, ax111x, ax108x, ax109x, ax106x, ax107x, ax104x, ax105x, ax102x, ax103x, ax100x, ax101x, ax98x, ax99x, ax96x, ax97x, ax94x, ax95x, ax92x, ax93x, ax90x, ax91x, ax88x, ax89x, ax86x, ax87x, ax84x, ax85x, ax82x, ax83x, ax80x, ax81x, ax78x, ax79x, ax76x, ax77x, ax74x, ax75x, ax72x, ax73x, ax70x, ax71x, ax68x, ax69x, ax66x, ax67x, ax64x, ax65x, ax62x, ax63x, ax60x, ax61x, ax58x, ax59x, ax56x, ax57x, ax54x, ax55x, ax52x, ax53x, ax50x, ax51x, ax48x, ax49x, ax46x, ax47x, ax44x, ax45x, ax42x, ax43x, ax40x, ax41x, ax38x, ax39x, ax36x, ax37x, ax34x, ax35x, ax32x, ax33x, ax30x, ax31x, ax28x, ax29x, ax26x, ax27x, ax24x, ax25x, ax22x, ax23x, ax20x, ax21x, ax18x, ax19x, ax16x, ax17x, ax14x, ax15x, ax12x, ax13x, ax10x, ax11x, ax8x, ax9x, ax6x, ax7x, ax4x, ax5x, ax2x, ax3x, ax0x, ax1x, asqrtx0x, asqrtx1x, asqrtx2x, asqrtx3x, asqrtx4x, asqrtx5x, asqrtx6x, asqrtx7x, asqrtx8x, asqrtx9x, asqrtx10x, asqrtx11x, asqrtx12x, asqrtx13x, asqrtx14x, asqrtx15x, asqrtx16x, asqrtx17x, asqrtx18x, asqrtx19x, asqrtx20x, asqrtx21x, asqrtx22x, asqrtx23x, asqrtx24x, asqrtx25x, asqrtx26x, asqrtx27x, asqrtx28x, asqrtx29x, asqrtx30x, asqrtx31x, asqrtx32x, asqrtx33x, asqrtx34x, asqrtx35x, asqrtx36x, asqrtx37x, asqrtx38x, asqrtx39x, asqrtx40x, asqrtx41x, asqrtx42x, asqrtx43x, asqrtx44x, asqrtx45x, asqrtx46x, asqrtx47x, asqrtx48x, asqrtx49x, asqrtx50x, asqrtx51x, asqrtx52x, asqrtx53x, asqrtx54x, asqrtx55x, asqrtx56x, asqrtx57x, asqrtx58x, asqrtx59x, asqrtx60x, asqrtx61x, asqrtx62x, asqrtx63x);

	input ax126x;
	input ax127x;
	input ax124x;
	input ax125x;
	input ax122x;
	input ax123x;
	input ax120x;
	input ax121x;
	input ax118x;
	input ax119x;
	input ax116x;
	input ax117x;
	input ax114x;
	input ax115x;
	input ax112x;
	input ax113x;
	input ax110x;
	input ax111x;
	input ax108x;
	input ax109x;
	input ax106x;
	input ax107x;
	input ax104x;
	input ax105x;
	input ax102x;
	input ax103x;
	input ax100x;
	input ax101x;
	input ax98x;
	input ax99x;
	input ax96x;
	input ax97x;
	input ax94x;
	input ax95x;
	input ax92x;
	input ax93x;
	input ax90x;
	input ax91x;
	input ax88x;
	input ax89x;
	input ax86x;
	input ax87x;
	input ax84x;
	input ax85x;
	input ax82x;
	input ax83x;
	input ax80x;
	input ax81x;
	input ax78x;
	input ax79x;
	input ax76x;
	input ax77x;
	input ax74x;
	input ax75x;
	input ax72x;
	input ax73x;
	input ax70x;
	input ax71x;
	input ax68x;
	input ax69x;
	input ax66x;
	input ax67x;
	input ax64x;
	input ax65x;
	input ax62x;
	input ax63x;
	input ax60x;
	input ax61x;
	input ax58x;
	input ax59x;
	input ax56x;
	input ax57x;
	input ax54x;
	input ax55x;
	input ax52x;
	input ax53x;
	input ax50x;
	input ax51x;
	input ax48x;
	input ax49x;
	input ax46x;
	input ax47x;
	input ax44x;
	input ax45x;
	input ax42x;
	input ax43x;
	input ax40x;
	input ax41x;
	input ax38x;
	input ax39x;
	input ax36x;
	input ax37x;
	input ax34x;
	input ax35x;
	input ax32x;
	input ax33x;
	input ax30x;
	input ax31x;
	input ax28x;
	input ax29x;
	input ax26x;
	input ax27x;
	input ax24x;
	input ax25x;
	input ax22x;
	input ax23x;
	input ax20x;
	input ax21x;
	input ax18x;
	input ax19x;
	input ax16x;
	input ax17x;
	input ax14x;
	input ax15x;
	input ax12x;
	input ax13x;
	input ax10x;
	input ax11x;
	input ax8x;
	input ax9x;
	input ax6x;
	input ax7x;
	input ax4x;
	input ax5x;
	input ax2x;
	input ax3x;
	input ax0x;
	input ax1x;
	output asqrtx0x;
	output asqrtx1x;
	output asqrtx2x;
	output asqrtx3x;
	output asqrtx4x;
	output asqrtx5x;
	output asqrtx6x;
	output asqrtx7x;
	output asqrtx8x;
	output asqrtx9x;
	output asqrtx10x;
	output asqrtx11x;
	output asqrtx12x;
	output asqrtx13x;
	output asqrtx14x;
	output asqrtx15x;
	output asqrtx16x;
	output asqrtx17x;
	output asqrtx18x;
	output asqrtx19x;
	output asqrtx20x;
	output asqrtx21x;
	output asqrtx22x;
	output asqrtx23x;
	output asqrtx24x;
	output asqrtx25x;
	output asqrtx26x;
	output asqrtx27x;
	output asqrtx28x;
	output asqrtx29x;
	output asqrtx30x;
	output asqrtx31x;
	output asqrtx32x;
	output asqrtx33x;
	output asqrtx34x;
	output asqrtx35x;
	output asqrtx36x;
	output asqrtx37x;
	output asqrtx38x;
	output asqrtx39x;
	output asqrtx40x;
	output asqrtx41x;
	output asqrtx42x;
	output asqrtx43x;
	output asqrtx44x;
	output asqrtx45x;
	output asqrtx46x;
	output asqrtx47x;
	output asqrtx48x;
	output asqrtx49x;
	output asqrtx50x;
	output asqrtx51x;
	output asqrtx52x;
	output asqrtx53x;
	output asqrtx54x;
	output asqrtx55x;
	output asqrtx56x;
	output asqrtx57x;
	output asqrtx58x;
	output asqrtx59x;
	output asqrtx60x;
	output asqrtx61x;
	output asqrtx62x;
	output asqrtx63x;



	wire g3496, g3400, g3395, g3187, g3178, g2980, g3030, g2779, g2825, g2585, g2627;
	wire g2398, g2436, g2218, g2252, g2045, g2075, g1879, g1905, g1720, g1742, g1568;
	wire g1586, g1423, g1437, g1285, g1295, g1154, g1160, g1030, g1032, g914, g851;
	wire g803, g744, g700, g645, g604, g553, g515, g468, g433, g390, g358;
	wire g319, g290, g255, g229, g198, g174, g147, g127, g104, g87, g68;
	wire g54, g39, g27, g18, g8, g2, g4, g1, g3, g5, g6;
	wire g7, g9, g10, g11, g12, g13, g14, g15, g16, g17, g19;
	wire g20, g21, g22, g23, g24, g25, g26, g28, g29, g30, g31;
	wire g32, g33, g34, g35, g36, g37, g38, g40, g41, g42, g43;
	wire g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g55;
	wire g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66;
	wire g67, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78;
	wire g79, g80, g81, g82, g83, g84, g85, g86, g88, g89, g90;
	wire g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101;
	wire g102, g103, g105, g106, g107, g108, g109, g110, g111, g112, g113;
	wire g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124;
	wire g125, g126, g128, g129, g130, g131, g132, g133, g134, g135, g136;
	wire g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g148;
	wire g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159;
	wire g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g170;
	wire g171, g172, g173, g175, g176, g177, g178, g179, g180, g181, g182;
	wire g183, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193;
	wire g194, g195, g196, g197, g199, g200, g201, g202, g203, g204, g205;
	wire g206, g207, g208, g209, g210, g211, g212, g213, g214, g215, g216;
	wire g217, g218, g219, g220, g221, g222, g223, g224, g225, g226, g227;
	wire g228, g230, g231, g232, g233, g234, g235, g236, g237, g238, g239;
	wire g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250;
	wire g251, g252, g253, g254, g256, g257, g258, g259, g260, g261, g262;
	wire g263, g264, g265, g266, g267, g268, g269, g270, g271, g272, g273;
	wire g274, g275, g276, g277, g278, g279, g280, g281, g282, g283, g284;
	wire g285, g286, g287, g288, g289, g291, g292, g293, g294, g295, g296;
	wire g297, g298, g299, g300, g301, g302, g303, g304, g305, g306, g307;
	wire g308, g309, g310, g311, g312, g313, g314, g315, g316, g317, g318;
	wire g320, g321, g322, g323, g324, g325, g326, g327, g328, g329, g330;
	wire g331, g332, g333, g334, g335, g336, g337, g338, g339, g340, g341;
	wire g342, g343, g344, g345, g346, g347, g348, g349, g350, g351, g352;
	wire g353, g354, g355, g356, g357, g359, g360, g361, g362, g363, g364;
	wire g365, g366, g367, g368, g369, g370, g371, g372, g373, g374, g375;
	wire g376, g377, g378, g379, g380, g381, g382, g383, g384, g385, g386;
	wire g387, g388, g389, g391, g392, g393, g394, g395, g396, g397, g398;
	wire g399, g400, g401, g402, g403, g404, g405, g406, g407, g408, g409;
	wire g410, g411, g412, g413, g414, g415, g416, g417, g418, g419, g420;
	wire g421, g422, g423, g424, g425, g426, g427, g428, g429, g430, g431;
	wire g432, g434, g435, g436, g437, g438, g439, g440, g441, g442, g443;
	wire g444, g445, g446, g447, g448, g449, g450, g451, g452, g453, g454;
	wire g455, g456, g457, g458, g459, g460, g461, g462, g463, g464, g465;
	wire g466, g467, g469, g470, g471, g472, g473, g474, g475, g476, g477;
	wire g478, g479, g480, g481, g482, g483, g484, g485, g486, g487, g488;
	wire g489, g490, g491, g492, g493, g494, g495, g496, g497, g498, g499;
	wire g500, g501, g502, g503, g504, g505, g506, g507, g508, g509, g510;
	wire g511, g512, g513, g514, g516, g517, g518, g519, g520, g521, g522;
	wire g523, g524, g525, g526, g527, g528, g529, g530, g531, g532, g533;
	wire g534, g535, g536, g537, g538, g539, g540, g541, g542, g543, g544;
	wire g545, g546, g547, g548, g549, g550, g551, g552, g554, g555, g556;
	wire g557, g558, g559, g560, g561, g562, g563, g564, g565, g566, g567;
	wire g568, g569, g570, g571, g572, g573, g574, g575, g576, g577, g578;
	wire g579, g580, g581, g582, g583, g584, g585, g586, g587, g588, g589;
	wire g590, g591, g592, g593, g594, g595, g596, g597, g598, g599, g600;
	wire g601, g602, g603, g605, g606, g607, g608, g609, g610, g611, g612;
	wire g613, g614, g615, g616, g617, g618, g619, g620, g621, g622, g623;
	wire g624, g625, g626, g627, g628, g629, g630, g631, g632, g633, g634;
	wire g635, g636, g637, g638, g639, g640, g641, g642, g643, g644, g646;
	wire g647, g648, g649, g650, g651, g652, g653, g654, g655, g656, g657;
	wire g658, g659, g660, g661, g662, g663, g664, g665, g666, g667, g668;
	wire g669, g670, g671, g672, g673, g674, g675, g676, g677, g678, g679;
	wire g680, g681, g682, g683, g684, g685, g686, g687, g688, g689, g690;
	wire g691, g692, g693, g694, g695, g696, g697, g698, g699, g701, g702;
	wire g703, g704, g705, g706, g707, g708, g709, g710, g711, g712, g713;
	wire g714, g715, g716, g717, g718, g719, g720, g721, g722, g723, g724;
	wire g725, g726, g727, g728, g729, g730, g731, g732, g733, g734, g735;
	wire g736, g737, g738, g739, g740, g741, g742, g743, g745, g746, g747;
	wire g748, g749, g750, g751, g752, g753, g754, g755, g756, g757, g758;
	wire g759, g760, g761, g762, g763, g764, g765, g766, g767, g768, g769;
	wire g770, g771, g772, g773, g774, g775, g776, g777, g778, g779, g780;
	wire g781, g782, g783, g784, g785, g786, g787, g788, g789, g790, g791;
	wire g792, g793, g794, g795, g796, g797, g798, g799, g800, g801, g802;
	wire g804, g805, g806, g807, g808, g809, g810, g811, g812, g813, g814;
	wire g815, g816, g817, g818, g819, g820, g821, g822, g823, g824, g825;
	wire g826, g827, g828, g829, g830, g831, g832, g833, g834, g835, g836;
	wire g837, g838, g839, g840, g841, g842, g843, g844, g845, g846, g847;
	wire g848, g849, g850, g852, g853, g854, g855, g856, g857, g858, g859;
	wire g860, g861, g862, g863, g864, g865, g866, g867, g868, g869, g870;
	wire g871, g872, g873, g874, g875, g876, g877, g878, g879, g880, g881;
	wire g882, g883, g884, g885, g886, g887, g888, g889, g890, g891, g892;
	wire g893, g894, g895, g896, g897, g898, g899, g900, g901, g902, g903;
	wire g904, g905, g906, g907, g908, g909, g910, g911, g912, g913, g915;
	wire g916, g917, g918, g919, g920, g921, g922, g923, g924, g925, g926;
	wire g927, g928, g929, g930, g931, g932, g933, g934, g935, g936, g937;
	wire g938, g939, g940, g941, g942, g943, g944, g945, g946, g947, g948;
	wire g949, g950, g951, g952, g953, g954, g955, g956, g957, g958, g959;
	wire g960, g961, g962, g963, g964, g965, g966, g967, g968, g969, g970;
	wire g971, g972, g973, g974, g975, g976, g977, g978, g979, g980, g981;
	wire g982, g983, g984, g985, g986, g987, g988, g989, g990, g991, g992;
	wire g993, g994, g995, g996, g997, g998, g999, g1000, g1001, g1002, g1003;
	wire g1004, g1005, g1006, g1007, g1008, g1009, g1010, g1011, g1012, g1013, g1014;
	wire g1015, g1016, g1017, g1018, g1019, g1020, g1021, g1022, g1023, g1024, g1025;
	wire g1026, g1027, g1028, g1029, g1031, g1033, g1034, g1035, g1036, g1037, g1038;
	wire g1039, g1040, g1041, g1042, g1043, g1044, g1045, g1046, g1047, g1048, g1049;
	wire g1050, g1051, g1052, g1053, g1054, g1055, g1056, g1057, g1058, g1059, g1060;
	wire g1061, g1062, g1063, g1064, g1065, g1066, g1067, g1068, g1069, g1070, g1071;
	wire g1072, g1073, g1074, g1075, g1076, g1077, g1078, g1079, g1080, g1081, g1082;
	wire g1083, g1084, g1085, g1086, g1087, g1088, g1089, g1090, g1091, g1092, g1093;
	wire g1094, g1095, g1096, g1097, g1098, g1099, g1100, g1101, g1102, g1103, g1104;
	wire g1105, g1106, g1107, g1108, g1109, g1110, g1111, g1112, g1113, g1114, g1115;
	wire g1116, g1117, g1118, g1119, g1120, g1121, g1122, g1123, g1124, g1125, g1126;
	wire g1127, g1128, g1129, g1130, g1131, g1132, g1133, g1134, g1135, g1136, g1137;
	wire g1138, g1139, g1140, g1141, g1142, g1143, g1144, g1145, g1146, g1147, g1148;
	wire g1149, g1150, g1151, g1152, g1153, g1155, g1156, g1157, g1158, g1159, g1161;
	wire g1162, g1163, g1164, g1165, g1166, g1167, g1168, g1169, g1170, g1171, g1172;
	wire g1173, g1174, g1175, g1176, g1177, g1178, g1179, g1180, g1181, g1182, g1183;
	wire g1184, g1185, g1186, g1187, g1188, g1189, g1190, g1191, g1192, g1193, g1194;
	wire g1195, g1196, g1197, g1198, g1199, g1200, g1201, g1202, g1203, g1204, g1205;
	wire g1206, g1207, g1208, g1209, g1210, g1211, g1212, g1213, g1214, g1215, g1216;
	wire g1217, g1218, g1219, g1220, g1221, g1222, g1223, g1224, g1225, g1226, g1227;
	wire g1228, g1229, g1230, g1231, g1232, g1233, g1234, g1235, g1236, g1237, g1238;
	wire g1239, g1240, g1241, g1242, g1243, g1244, g1245, g1246, g1247, g1248, g1249;
	wire g1250, g1251, g1252, g1253, g1254, g1255, g1256, g1257, g1258, g1259, g1260;
	wire g1261, g1262, g1263, g1264, g1265, g1266, g1267, g1268, g1269, g1270, g1271;
	wire g1272, g1273, g1274, g1275, g1276, g1277, g1278, g1279, g1280, g1281, g1282;
	wire g1283, g1284, g1286, g1287, g1288, g1289, g1290, g1291, g1292, g1293, g1294;
	wire g1296, g1297, g1298, g1299, g1300, g1301, g1302, g1303, g1304, g1305, g1306;
	wire g1307, g1308, g1309, g1310, g1311, g1312, g1313, g1314, g1315, g1316, g1317;
	wire g1318, g1319, g1320, g1321, g1322, g1323, g1324, g1325, g1326, g1327, g1328;
	wire g1329, g1330, g1331, g1332, g1333, g1334, g1335, g1336, g1337, g1338, g1339;
	wire g1340, g1341, g1342, g1343, g1344, g1345, g1346, g1347, g1348, g1349, g1350;
	wire g1351, g1352, g1353, g1354, g1355, g1356, g1357, g1358, g1359, g1360, g1361;
	wire g1362, g1363, g1364, g1365, g1366, g1367, g1368, g1369, g1370, g1371, g1372;
	wire g1373, g1374, g1375, g1376, g1377, g1378, g1379, g1380, g1381, g1382, g1383;
	wire g1384, g1385, g1386, g1387, g1388, g1389, g1390, g1391, g1392, g1393, g1394;
	wire g1395, g1396, g1397, g1398, g1399, g1400, g1401, g1402, g1403, g1404, g1405;
	wire g1406, g1407, g1408, g1409, g1410, g1411, g1412, g1413, g1414, g1415, g1416;
	wire g1417, g1418, g1419, g1420, g1421, g1422, g1424, g1425, g1426, g1427, g1428;
	wire g1429, g1430, g1431, g1432, g1433, g1434, g1435, g1436, g1438, g1439, g1440;
	wire g1441, g1442, g1443, g1444, g1445, g1446, g1447, g1448, g1449, g1450, g1451;
	wire g1452, g1453, g1454, g1455, g1456, g1457, g1458, g1459, g1460, g1461, g1462;
	wire g1463, g1464, g1465, g1466, g1467, g1468, g1469, g1470, g1471, g1472, g1473;
	wire g1474, g1475, g1476, g1477, g1478, g1479, g1480, g1481, g1482, g1483, g1484;
	wire g1485, g1486, g1487, g1488, g1489, g1490, g1491, g1492, g1493, g1494, g1495;
	wire g1496, g1497, g1498, g1499, g1500, g1501, g1502, g1503, g1504, g1505, g1506;
	wire g1507, g1508, g1509, g1510, g1511, g1512, g1513, g1514, g1515, g1516, g1517;
	wire g1518, g1519, g1520, g1521, g1522, g1523, g1524, g1525, g1526, g1527, g1528;
	wire g1529, g1530, g1531, g1532, g1533, g1534, g1535, g1536, g1537, g1538, g1539;
	wire g1540, g1541, g1542, g1543, g1544, g1545, g1546, g1547, g1548, g1549, g1550;
	wire g1551, g1552, g1553, g1554, g1555, g1556, g1557, g1558, g1559, g1560, g1561;
	wire g1562, g1563, g1564, g1565, g1566, g1567, g1569, g1570, g1571, g1572, g1573;
	wire g1574, g1575, g1576, g1577, g1578, g1579, g1580, g1581, g1582, g1583, g1584;
	wire g1585, g1587, g1588, g1589, g1590, g1591, g1592, g1593, g1594, g1595, g1596;
	wire g1597, g1598, g1599, g1600, g1601, g1602, g1603, g1604, g1605, g1606, g1607;
	wire g1608, g1609, g1610, g1611, g1612, g1613, g1614, g1615, g1616, g1617, g1618;
	wire g1619, g1620, g1621, g1622, g1623, g1624, g1625, g1626, g1627, g1628, g1629;
	wire g1630, g1631, g1632, g1633, g1634, g1635, g1636, g1637, g1638, g1639, g1640;
	wire g1641, g1642, g1643, g1644, g1645, g1646, g1647, g1648, g1649, g1650, g1651;
	wire g1652, g1653, g1654, g1655, g1656, g1657, g1658, g1659, g1660, g1661, g1662;
	wire g1663, g1664, g1665, g1666, g1667, g1668, g1669, g1670, g1671, g1672, g1673;
	wire g1674, g1675, g1676, g1677, g1678, g1679, g1680, g1681, g1682, g1683, g1684;
	wire g1685, g1686, g1687, g1688, g1689, g1690, g1691, g1692, g1693, g1694, g1695;
	wire g1696, g1697, g1698, g1699, g1700, g1701, g1702, g1703, g1704, g1705, g1706;
	wire g1707, g1708, g1709, g1710, g1711, g1712, g1713, g1714, g1715, g1716, g1717;
	wire g1718, g1719, g1721, g1722, g1723, g1724, g1725, g1726, g1727, g1728, g1729;
	wire g1730, g1731, g1732, g1733, g1734, g1735, g1736, g1737, g1738, g1739, g1740;
	wire g1741, g1743, g1744, g1745, g1746, g1747, g1748, g1749, g1750, g1751, g1752;
	wire g1753, g1754, g1755, g1756, g1757, g1758, g1759, g1760, g1761, g1762, g1763;
	wire g1764, g1765, g1766, g1767, g1768, g1769, g1770, g1771, g1772, g1773, g1774;
	wire g1775, g1776, g1777, g1778, g1779, g1780, g1781, g1782, g1783, g1784, g1785;
	wire g1786, g1787, g1788, g1789, g1790, g1791, g1792, g1793, g1794, g1795, g1796;
	wire g1797, g1798, g1799, g1800, g1801, g1802, g1803, g1804, g1805, g1806, g1807;
	wire g1808, g1809, g1810, g1811, g1812, g1813, g1814, g1815, g1816, g1817, g1818;
	wire g1819, g1820, g1821, g1822, g1823, g1824, g1825, g1826, g1827, g1828, g1829;
	wire g1830, g1831, g1832, g1833, g1834, g1835, g1836, g1837, g1838, g1839, g1840;
	wire g1841, g1842, g1843, g1844, g1845, g1846, g1847, g1848, g1849, g1850, g1851;
	wire g1852, g1853, g1854, g1855, g1856, g1857, g1858, g1859, g1860, g1861, g1862;
	wire g1863, g1864, g1865, g1866, g1867, g1868, g1869, g1870, g1871, g1872, g1873;
	wire g1874, g1875, g1876, g1877, g1878, g1880, g1881, g1882, g1883, g1884, g1885;
	wire g1886, g1887, g1888, g1889, g1890, g1891, g1892, g1893, g1894, g1895, g1896;
	wire g1897, g1898, g1899, g1900, g1901, g1902, g1903, g1904, g1906, g1907, g1908;
	wire g1909, g1910, g1911, g1912, g1913, g1914, g1915, g1916, g1917, g1918, g1919;
	wire g1920, g1921, g1922, g1923, g1924, g1925, g1926, g1927, g1928, g1929, g1930;
	wire g1931, g1932, g1933, g1934, g1935, g1936, g1937, g1938, g1939, g1940, g1941;
	wire g1942, g1943, g1944, g1945, g1946, g1947, g1948, g1949, g1950, g1951, g1952;
	wire g1953, g1954, g1955, g1956, g1957, g1958, g1959, g1960, g1961, g1962, g1963;
	wire g1964, g1965, g1966, g1967, g1968, g1969, g1970, g1971, g1972, g1973, g1974;
	wire g1975, g1976, g1977, g1978, g1979, g1980, g1981, g1982, g1983, g1984, g1985;
	wire g1986, g1987, g1988, g1989, g1990, g1991, g1992, g1993, g1994, g1995, g1996;
	wire g1997, g1998, g1999, g2000, g2001, g2002, g2003, g2004, g2005, g2006, g2007;
	wire g2008, g2009, g2010, g2011, g2012, g2013, g2014, g2015, g2016, g2017, g2018;
	wire g2019, g2020, g2021, g2022, g2023, g2024, g2025, g2026, g2027, g2028, g2029;
	wire g2030, g2031, g2032, g2033, g2034, g2035, g2036, g2037, g2038, g2039, g2040;
	wire g2041, g2042, g2043, g2044, g2046, g2047, g2048, g2049, g2050, g2051, g2052;
	wire g2053, g2054, g2055, g2056, g2057, g2058, g2059, g2060, g2061, g2062, g2063;
	wire g2064, g2065, g2066, g2067, g2068, g2069, g2070, g2071, g2072, g2073, g2074;
	wire g2076, g2077, g2078, g2079, g2080, g2081, g2082, g2083, g2084, g2085, g2086;
	wire g2087, g2088, g2089, g2090, g2091, g2092, g2093, g2094, g2095, g2096, g2097;
	wire g2098, g2099, g2100, g2101, g2102, g2103, g2104, g2105, g2106, g2107, g2108;
	wire g2109, g2110, g2111, g2112, g2113, g2114, g2115, g2116, g2117, g2118, g2119;
	wire g2120, g2121, g2122, g2123, g2124, g2125, g2126, g2127, g2128, g2129, g2130;
	wire g2131, g2132, g2133, g2134, g2135, g2136, g2137, g2138, g2139, g2140, g2141;
	wire g2142, g2143, g2144, g2145, g2146, g2147, g2148, g2149, g2150, g2151, g2152;
	wire g2153, g2154, g2155, g2156, g2157, g2158, g2159, g2160, g2161, g2162, g2163;
	wire g2164, g2165, g2166, g2167, g2168, g2169, g2170, g2171, g2172, g2173, g2174;
	wire g2175, g2176, g2177, g2178, g2179, g2180, g2181, g2182, g2183, g2184, g2185;
	wire g2186, g2187, g2188, g2189, g2190, g2191, g2192, g2193, g2194, g2195, g2196;
	wire g2197, g2198, g2199, g2200, g2201, g2202, g2203, g2204, g2205, g2206, g2207;
	wire g2208, g2209, g2210, g2211, g2212, g2213, g2214, g2215, g2216, g2217, g2219;
	wire g2220, g2221, g2222, g2223, g2224, g2225, g2226, g2227, g2228, g2229, g2230;
	wire g2231, g2232, g2233, g2234, g2235, g2236, g2237, g2238, g2239, g2240, g2241;
	wire g2242, g2243, g2244, g2245, g2246, g2247, g2248, g2249, g2250, g2251, g2253;
	wire g2254, g2255, g2256, g2257, g2258, g2259, g2260, g2261, g2262, g2263, g2264;
	wire g2265, g2266, g2267, g2268, g2269, g2270, g2271, g2272, g2273, g2274, g2275;
	wire g2276, g2277, g2278, g2279, g2280, g2281, g2282, g2283, g2284, g2285, g2286;
	wire g2287, g2288, g2289, g2290, g2291, g2292, g2293, g2294, g2295, g2296, g2297;
	wire g2298, g2299, g2300, g2301, g2302, g2303, g2304, g2305, g2306, g2307, g2308;
	wire g2309, g2310, g2311, g2312, g2313, g2314, g2315, g2316, g2317, g2318, g2319;
	wire g2320, g2321, g2322, g2323, g2324, g2325, g2326, g2327, g2328, g2329, g2330;
	wire g2331, g2332, g2333, g2334, g2335, g2336, g2337, g2338, g2339, g2340, g2341;
	wire g2342, g2343, g2344, g2345, g2346, g2347, g2348, g2349, g2350, g2351, g2352;
	wire g2353, g2354, g2355, g2356, g2357, g2358, g2359, g2360, g2361, g2362, g2363;
	wire g2364, g2365, g2366, g2367, g2368, g2369, g2370, g2371, g2372, g2373, g2374;
	wire g2375, g2376, g2377, g2378, g2379, g2380, g2381, g2382, g2383, g2384, g2385;
	wire g2386, g2387, g2388, g2389, g2390, g2391, g2392, g2393, g2394, g2395, g2396;
	wire g2397, g2399, g2400, g2401, g2402, g2403, g2404, g2405, g2406, g2407, g2408;
	wire g2409, g2410, g2411, g2412, g2413, g2414, g2415, g2416, g2417, g2418, g2419;
	wire g2420, g2421, g2422, g2423, g2424, g2425, g2426, g2427, g2428, g2429, g2430;
	wire g2431, g2432, g2433, g2434, g2435, g2437, g2438, g2439, g2440, g2441, g2442;
	wire g2443, g2444, g2445, g2446, g2447, g2448, g2449, g2450, g2451, g2452, g2453;
	wire g2454, g2455, g2456, g2457, g2458, g2459, g2460, g2461, g2462, g2463, g2464;
	wire g2465, g2466, g2467, g2468, g2469, g2470, g2471, g2472, g2473, g2474, g2475;
	wire g2476, g2477, g2478, g2479, g2480, g2481, g2482, g2483, g2484, g2485, g2486;
	wire g2487, g2488, g2489, g2490, g2491, g2492, g2493, g2494, g2495, g2496, g2497;
	wire g2498, g2499, g2500, g2501, g2502, g2503, g2504, g2505, g2506, g2507, g2508;
	wire g2509, g2510, g2511, g2512, g2513, g2514, g2515, g2516, g2517, g2518, g2519;
	wire g2520, g2521, g2522, g2523, g2524, g2525, g2526, g2527, g2528, g2529, g2530;
	wire g2531, g2532, g2533, g2534, g2535, g2536, g2537, g2538, g2539, g2540, g2541;
	wire g2542, g2543, g2544, g2545, g2546, g2547, g2548, g2549, g2550, g2551, g2552;
	wire g2553, g2554, g2555, g2556, g2557, g2558, g2559, g2560, g2561, g2562, g2563;
	wire g2564, g2565, g2566, g2567, g2568, g2569, g2570, g2571, g2572, g2573, g2574;
	wire g2575, g2576, g2577, g2578, g2579, g2580, g2581, g2582, g2583, g2584, g2586;
	wire g2587, g2588, g2589, g2590, g2591, g2592, g2593, g2594, g2595, g2596, g2597;
	wire g2598, g2599, g2600, g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608;
	wire g2609, g2610, g2611, g2612, g2613, g2614, g2615, g2616, g2617, g2618, g2619;
	wire g2620, g2621, g2622, g2623, g2624, g2625, g2626, g2628, g2629, g2630, g2631;
	wire g2632, g2633, g2634, g2635, g2636, g2637, g2638, g2639, g2640, g2641, g2642;
	wire g2643, g2644, g2645, g2646, g2647, g2648, g2649, g2650, g2651, g2652, g2653;
	wire g2654, g2655, g2656, g2657, g2658, g2659, g2660, g2661, g2662, g2663, g2664;
	wire g2665, g2666, g2667, g2668, g2669, g2670, g2671, g2672, g2673, g2674, g2675;
	wire g2676, g2677, g2678, g2679, g2680, g2681, g2682, g2683, g2684, g2685, g2686;
	wire g2687, g2688, g2689, g2690, g2691, g2692, g2693, g2694, g2695, g2696, g2697;
	wire g2698, g2699, g2700, g2701, g2702, g2703, g2704, g2705, g2706, g2707, g2708;
	wire g2709, g2710, g2711, g2712, g2713, g2714, g2715, g2716, g2717, g2718, g2719;
	wire g2720, g2721, g2722, g2723, g2724, g2725, g2726, g2727, g2728, g2729, g2730;
	wire g2731, g2732, g2733, g2734, g2735, g2736, g2737, g2738, g2739, g2740, g2741;
	wire g2742, g2743, g2744, g2745, g2746, g2747, g2748, g2749, g2750, g2751, g2752;
	wire g2753, g2754, g2755, g2756, g2757, g2758, g2759, g2760, g2761, g2762, g2763;
	wire g2764, g2765, g2766, g2767, g2768, g2769, g2770, g2771, g2772, g2773, g2774;
	wire g2775, g2776, g2777, g2778, g2780, g2781, g2782, g2783, g2784, g2785, g2786;
	wire g2787, g2788, g2789, g2790, g2791, g2792, g2793, g2794, g2795, g2796, g2797;
	wire g2798, g2799, g2800, g2801, g2802, g2803, g2804, g2805, g2806, g2807, g2808;
	wire g2809, g2810, g2811, g2812, g2813, g2814, g2815, g2816, g2817, g2818, g2819;
	wire g2820, g2821, g2822, g2823, g2824, g2826, g2827, g2828, g2829, g2830, g2831;
	wire g2832, g2833, g2834, g2835, g2836, g2837, g2838, g2839, g2840, g2841, g2842;
	wire g2843, g2844, g2845, g2846, g2847, g2848, g2849, g2850, g2851, g2852, g2853;
	wire g2854, g2855, g2856, g2857, g2858, g2859, g2860, g2861, g2862, g2863, g2864;
	wire g2865, g2866, g2867, g2868, g2869, g2870, g2871, g2872, g2873, g2874, g2875;
	wire g2876, g2877, g2878, g2879, g2880, g2881, g2882, g2883, g2884, g2885, g2886;
	wire g2887, g2888, g2889, g2890, g2891, g2892, g2893, g2894, g2895, g2896, g2897;
	wire g2898, g2899, g2900, g2901, g2902, g2903, g2904, g2905, g2906, g2907, g2908;
	wire g2909, g2910, g2911, g2912, g2913, g2914, g2915, g2916, g2917, g2918, g2919;
	wire g2920, g2921, g2922, g2923, g2924, g2925, g2926, g2927, g2928, g2929, g2930;
	wire g2931, g2932, g2933, g2934, g2935, g2936, g2937, g2938, g2939, g2940, g2941;
	wire g2942, g2943, g2944, g2945, g2946, g2947, g2948, g2949, g2950, g2951, g2952;
	wire g2953, g2954, g2955, g2956, g2957, g2958, g2959, g2960, g2961, g2962, g2963;
	wire g2964, g2965, g2966, g2967, g2968, g2969, g2970, g2971, g2972, g2973, g2974;
	wire g2975, g2976, g2977, g2978, g2979, g2981, g2982, g2983, g2984, g2985, g2986;
	wire g2987, g2988, g2989, g2990, g2991, g2992, g2993, g2994, g2995, g2996, g2997;
	wire g2998, g2999, g3000, g3001, g3002, g3003, g3004, g3005, g3006, g3007, g3008;
	wire g3009, g3010, g3011, g3012, g3013, g3014, g3015, g3016, g3017, g3018, g3019;
	wire g3020, g3021, g3022, g3023, g3024, g3025, g3026, g3027, g3028, g3029, g3031;
	wire g3032, g3033, g3034, g3035, g3036, g3037, g3038, g3039, g3040, g3041, g3042;
	wire g3043, g3044, g3045, g3046, g3047, g3048, g3049, g3050, g3051, g3052, g3053;
	wire g3054, g3055, g3056, g3057, g3058, g3059, g3060, g3061, g3062, g3063, g3064;
	wire g3065, g3066, g3067, g3068, g3069, g3070, g3071, g3072, g3073, g3074, g3075;
	wire g3076, g3077, g3078, g3079, g3080, g3081, g3082, g3083, g3084, g3085, g3086;
	wire g3087, g3088, g3089, g3090, g3091, g3092, g3093, g3094, g3095, g3096, g3097;
	wire g3098, g3099, g3100, g3101, g3102, g3103, g3104, g3105, g3106, g3107, g3108;
	wire g3109, g3110, g3111, g3112, g3113, g3114, g3115, g3116, g3117, g3118, g3119;
	wire g3120, g3121, g3122, g3123, g3124, g3125, g3126, g3127, g3128, g3129, g3130;
	wire g3131, g3132, g3133, g3134, g3135, g3136, g3137, g3138, g3139, g3140, g3141;
	wire g3142, g3143, g3144, g3145, g3146, g3147, g3148, g3149, g3150, g3151, g3152;
	wire g3153, g3154, g3155, g3156, g3157, g3158, g3159, g3160, g3161, g3162, g3163;
	wire g3164, g3165, g3166, g3167, g3168, g3169, g3170, g3171, g3172, g3173, g3174;
	wire g3175, g3176, g3177, g3179, g3180, g3181, g3182, g3183, g3184, g3185, g3186;
	wire g3188, g3189, g3190, g3191, g3192, g3193, g3194, g3195, g3196, g3197, g3198;
	wire g3199, g3200, g3201, g3202, g3203, g3204, g3205, g3206, g3207, g3208, g3209;
	wire g3210, g3211, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220;
	wire g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231;
	wire g3232, g3233, g3234, g3235, g3236, g3237, g3238, g3239, g3240, g3241, g3242;
	wire g3243, g3244, g3245, g3246, g3247, g3248, g3249, g3250, g3251, g3252, g3253;
	wire g3254, g3255, g3256, g3257, g3258, g3259, g3260, g3261, g3262, g3263, g3264;
	wire g3265, g3266, g3267, g3268, g3269, g3270, g3271, g3272, g3273, g3274, g3275;
	wire g3276, g3277, g3278, g3279, g3280, g3281, g3282, g3283, g3284, g3285, g3286;
	wire g3287, g3288, g3289, g3290, g3291, g3292, g3293, g3294, g3295, g3296, g3297;
	wire g3298, g3299, g3300, g3301, g3302, g3303, g3304, g3305, g3306, g3307, g3308;
	wire g3309, g3310, g3311, g3312, g3313, g3314, g3315, g3316, g3317, g3318, g3319;
	wire g3320, g3321, g3322, g3323, g3324, g3325, g3326, g3327, g3328, g3329, g3330;
	wire g3331, g3332, g3333, g3334, g3335, g3336, g3337, g3338, g3339, g3340, g3341;
	wire g3342, g3343, g3344, g3345, g3346, g3347, g3348, g3349, g3350, g3351, g3352;
	wire g3353, g3354, g3355, g3356, g3357, g3358, g3359, g3360, g3361, g3362, g3363;
	wire g3364, g3365, g3366, g3367, g3368, g3369, g3370, g3371, g3372, g3373, g3374;
	wire g3375, g3376, g3377, g3378, g3379, g3380, g3381, g3382, g3383, g3384, g3385;
	wire g3386, g3387, g3388, g3389, g3390, g3391, g3392, g3393, g3394, g3396, g3397;
	wire g3398, g3399, g3401, g3402, g3403, g3404, g3405, g3406, g3407, g3408, g3409;
	wire g3410, g3411, g3412, g3413, g3414, g3415, g3416, g3417, g3418, g3419, g3420;
	wire g3421, g3422, g3423, g3424, g3425, g3426, g3427, g3428, g3429, g3430, g3431;
	wire g3432, g3433, g3434, g3435, g3436, g3437, g3438, g3439, g3440, g3441, g3442;
	wire g3443, g3444, g3445, g3446, g3447, g3448, g3449, g3450, g3451, g3452, g3453;
	wire g3454, g3455, g3456, g3457, g3458, g3459, g3460, g3461, g3462, g3463, g3464;
	wire g3465, g3466, g3467, g3468, g3469, g3470, g3471, g3472, g3473, g3474, g3475;
	wire g3476, g3477, g3478, g3479, g3480, g3481, g3482, g3483, g3484, g3485, g3486;
	wire g3487, g3488, g3489, g3490, g3491, g3492, g3493, g3494, g3495, g3497, g3498;
	wire g3499, g3500, g3501, g3502, g3503, g3504, g3505, g3506, g3507, g3508, g3509;
	wire g3510, g3511, g3512, g3513, g3514, g3515, g3516, g3517, g3518, g3519, g3520;
	wire g3521, g3522, g3523, g3524, g3525, g3526, g3527, g3528, g3529, g3530, g3531;
	wire g3532, g3533, g3534, g3535, g3536, g3537, g3538, g3539, g3540, g3541, g3542;
	wire g3543, g3544, g3545, g3546, g3547, g3548, g3549, g3550, g3551, g3552, g3553;
	wire g3554, g3555, g3556, g3557, g3558, g3559, g3560, g3561, g3562, g3563, g3564;
	wire g3565, g3566, g3567, g3568, g3569, g3570, g3571, g3572, g3573, g3574, g3575;
	wire g3576, g3577, g3578, g3579, g3580, g3581, g3582, g3583, g3584, g3585, g3586;
	wire g3587, g3588, g3589, g3590, g3591, g3592, g3593, g3594, g3595, g3596, g3597;
	wire g3598, g3599, g3600, g3601, g3602, g3603, g3604, g3605, g3606, g3607, g3608;
	wire g3609, g3610, g3611, g3612, g3613, g3614, g3615, g3616, g3617, g3618, g3619;
	wire g3620, g3621, g3622, g3623;



	assign asqrtx1x = (((!g3496)));
	assign asqrtx2x = (((!g3400)));
	assign asqrtx3x = (((!g3395)));
	assign asqrtx4x = (((!g3187)));
	assign asqrtx5x = (((!g3178)));
	assign asqrtx6x = (((!g2980)));
	assign asqrtx7x = (((!g3030)));
	assign asqrtx8x = (((!g2779)));
	assign asqrtx9x = (((!g2825)));
	assign asqrtx10x = (((!g2585)));
	assign asqrtx11x = (((!g2627)));
	assign asqrtx12x = (((!g2398)));
	assign asqrtx13x = (((!g2436)));
	assign asqrtx14x = (((!g2218)));
	assign asqrtx15x = (((!g2252)));
	assign asqrtx16x = (((!g2045)));
	assign asqrtx17x = (((!g2075)));
	assign asqrtx18x = (((!g1879)));
	assign asqrtx19x = (((!g1905)));
	assign asqrtx20x = (((!g1720)));
	assign asqrtx21x = (((!g1742)));
	assign asqrtx22x = (((!g1568)));
	assign asqrtx23x = (((!g1586)));
	assign asqrtx24x = (((!g1423)));
	assign asqrtx25x = (((!g1437)));
	assign asqrtx26x = (((!g1285)));
	assign asqrtx27x = (((!g1295)));
	assign asqrtx28x = (((!g1154)));
	assign asqrtx29x = (((!g1160)));
	assign asqrtx30x = (((!g1030)));
	assign asqrtx31x = (((!g1032)));
	assign asqrtx32x = (((!g914)));
	assign asqrtx33x = (((!g851)));
	assign asqrtx34x = (((!g803)));
	assign asqrtx35x = (((!g744)));
	assign asqrtx36x = (((!g700)));
	assign asqrtx37x = (((!g645)));
	assign asqrtx38x = (((!g604)));
	assign asqrtx39x = (((!g553)));
	assign asqrtx40x = (((!g515)));
	assign asqrtx41x = (((!g468)));
	assign asqrtx42x = (((!g433)));
	assign asqrtx43x = (((!g390)));
	assign asqrtx44x = (((!g358)));
	assign asqrtx45x = (((!g319)));
	assign asqrtx46x = (((!g290)));
	assign asqrtx47x = (((!g255)));
	assign asqrtx48x = (((!g229)));
	assign asqrtx49x = (((!g198)));
	assign asqrtx50x = (((!g174)));
	assign asqrtx51x = (((!g147)));
	assign asqrtx52x = (((!g127)));
	assign asqrtx53x = (((!g104)));
	assign asqrtx54x = (((!g87)));
	assign asqrtx55x = (((!g68)));
	assign asqrtx56x = (((!g54)));
	assign asqrtx57x = (((!g39)));
	assign asqrtx58x = (((!g27)));
	assign asqrtx59x = (((!g18)));
	assign asqrtx60x = (((!g8)));
	assign asqrtx61x = (((!g2)));
	assign asqrtx62x = (((g4)));
	assign asqrtx63x = (((g1)));
	assign g1 = (((!ax126x) & (ax127x)) + ((ax126x) & (!ax127x)) + ((ax126x) & (ax127x)));
	assign g2 = (((!ax124x) & (!ax126x) & (!ax127x) & (!ax125x) & (!ax122x) & (!ax123x)) + ((!ax124x) & (!ax126x) & (!ax127x) & (ax125x) & (!ax122x) & (!ax123x)) + ((!ax124x) & (!ax126x) & (ax127x) & (ax125x) & (!ax122x) & (!ax123x)) + ((!ax124x) & (!ax126x) & (ax127x) & (ax125x) & (!ax122x) & (ax123x)) + ((!ax124x) & (!ax126x) & (ax127x) & (ax125x) & (ax122x) & (!ax123x)) + ((!ax124x) & (!ax126x) & (ax127x) & (ax125x) & (ax122x) & (ax123x)) + ((!ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (!ax122x) & (!ax123x)) + ((!ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (!ax122x) & (ax123x)) + ((!ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (ax122x) & (!ax123x)) + ((!ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (ax122x) & (ax123x)) + ((!ax124x) & (ax126x) & (!ax127x) & (ax125x) & (!ax122x) & (!ax123x)) + ((!ax124x) & (ax126x) & (ax127x) & (!ax125x) & (!ax122x) & (!ax123x)) + ((ax124x) & (!ax126x) & (!ax127x) & (!ax125x) & (!ax122x) & (!ax123x)) + ((ax124x) & (!ax126x) & (!ax127x) & (!ax125x) & (!ax122x) & (ax123x)) + ((ax124x) & (!ax126x) & (!ax127x) & (!ax125x) & (ax122x) & (!ax123x)) + ((ax124x) & (!ax126x) & (!ax127x) & (!ax125x) & (ax122x) & (ax123x)) + ((ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (!ax122x) & (!ax123x)) + ((ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (!ax122x) & (ax123x)) + ((ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (ax122x) & (!ax123x)) + ((ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (ax122x) & (ax123x)) + ((ax124x) & (!ax126x) & (ax127x) & (ax125x) & (!ax122x) & (!ax123x)) + ((ax124x) & (!ax126x) & (ax127x) & (ax125x) & (!ax122x) & (ax123x)) + ((ax124x) & (!ax126x) & (ax127x) & (ax125x) & (ax122x) & (!ax123x)) + ((ax124x) & (!ax126x) & (ax127x) & (ax125x) & (ax122x) & (ax123x)) + ((ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (!ax122x) & (!ax123x)) + ((ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (!ax122x) & (ax123x)) + ((ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (ax122x) & (!ax123x)) + ((ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (ax122x) & (ax123x)));
	assign g3 = (((!ax122x) & (!ax123x)));
	assign g4 = (((!ax124x) & (!ax126x) & (!ax127x) & (ax125x)) + ((!ax124x) & (!ax126x) & (ax127x) & (ax125x)) + ((!ax124x) & (ax126x) & (ax127x) & (!ax125x)) + ((!ax124x) & (ax126x) & (ax127x) & (ax125x)) + ((ax124x) & (!ax126x) & (!ax127x) & (!ax125x)) + ((ax124x) & (!ax126x) & (!ax127x) & (ax125x)) + ((ax124x) & (!ax126x) & (ax127x) & (!ax125x)) + ((ax124x) & (!ax126x) & (ax127x) & (ax125x)) + ((ax124x) & (ax126x) & (ax127x) & (!ax125x)) + ((ax124x) & (ax126x) & (ax127x) & (ax125x)));
	assign g5 = (((!ax120x) & (!ax121x)));
	assign g6 = (((!ax124x) & (!ax126x) & (!ax127x) & (!ax125x)) + ((!ax124x) & (!ax126x) & (ax127x) & (!ax125x)) + ((!ax124x) & (ax126x) & (!ax127x) & (!ax125x)) + ((!ax124x) & (ax126x) & (!ax127x) & (ax125x)) + ((ax124x) & (ax126x) & (!ax127x) & (!ax125x)) + ((ax124x) & (ax126x) & (!ax127x) & (ax125x)));
	assign g7 = (((!g4) & (!ax122x) & (!ax123x) & (!g2) & (!g5) & (!g6)) + ((!g4) & (!ax122x) & (!ax123x) & (!g2) & (!g5) & (g6)) + ((!g4) & (!ax122x) & (!ax123x) & (!g2) & (g5) & (!g6)) + ((!g4) & (!ax122x) & (!ax123x) & (!g2) & (g5) & (g6)) + ((!g4) & (!ax122x) & (!ax123x) & (g2) & (!g5) & (g6)) + ((!g4) & (!ax122x) & (ax123x) & (!g2) & (!g5) & (g6)) + ((!g4) & (!ax122x) & (ax123x) & (g2) & (!g5) & (!g6)) + ((!g4) & (!ax122x) & (ax123x) & (g2) & (!g5) & (g6)) + ((!g4) & (!ax122x) & (ax123x) & (g2) & (g5) & (!g6)) + ((!g4) & (!ax122x) & (ax123x) & (g2) & (g5) & (g6)) + ((!g4) & (ax122x) & (!ax123x) & (g2) & (!g5) & (g6)) + ((!g4) & (ax122x) & (!ax123x) & (g2) & (g5) & (g6)) + ((!g4) & (ax122x) & (ax123x) & (!g2) & (!g5) & (!g6)) + ((!g4) & (ax122x) & (ax123x) & (!g2) & (!g5) & (g6)) + ((!g4) & (ax122x) & (ax123x) & (!g2) & (g5) & (!g6)) + ((!g4) & (ax122x) & (ax123x) & (!g2) & (g5) & (g6)) + ((!g4) & (ax122x) & (ax123x) & (g2) & (!g5) & (!g6)) + ((!g4) & (ax122x) & (ax123x) & (g2) & (!g5) & (g6)) + ((!g4) & (ax122x) & (ax123x) & (g2) & (g5) & (!g6)) + ((!g4) & (ax122x) & (ax123x) & (g2) & (g5) & (g6)) + ((g4) & (!ax122x) & (!ax123x) & (!g2) & (!g5) & (!g6)) + ((g4) & (!ax122x) & (!ax123x) & (!g2) & (!g5) & (g6)) + ((g4) & (!ax122x) & (!ax123x) & (g2) & (!g5) & (g6)) + ((g4) & (!ax122x) & (ax123x) & (!g2) & (!g5) & (g6)) + ((g4) & (!ax122x) & (ax123x) & (g2) & (!g5) & (!g6)) + ((g4) & (!ax122x) & (ax123x) & (g2) & (!g5) & (g6)) + ((g4) & (ax122x) & (!ax123x) & (g2) & (!g5) & (g6)) + ((g4) & (ax122x) & (!ax123x) & (g2) & (g5) & (g6)) + ((g4) & (ax122x) & (ax123x) & (g2) & (!g5) & (!g6)) + ((g4) & (ax122x) & (ax123x) & (g2) & (!g5) & (g6)) + ((g4) & (ax122x) & (ax123x) & (g2) & (g5) & (!g6)) + ((g4) & (ax122x) & (ax123x) & (g2) & (g5) & (g6)));
	assign g8 = (((!ax124x) & (!ax126x) & (!ax127x) & (!ax125x) & (!g3) & (!g7)) + ((!ax124x) & (!ax126x) & (!ax127x) & (!ax125x) & (g3) & (!g7)) + ((!ax124x) & (!ax126x) & (!ax127x) & (ax125x) & (!g3) & (!g7)) + ((!ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (g3) & (!g7)) + ((!ax124x) & (!ax126x) & (ax127x) & (ax125x) & (!g3) & (!g7)) + ((!ax124x) & (!ax126x) & (ax127x) & (ax125x) & (g3) & (!g7)) + ((!ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (!g3) & (!g7)) + ((!ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (!g3) & (g7)) + ((!ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (g3) & (!g7)) + ((!ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (g3) & (g7)) + ((!ax124x) & (ax126x) & (!ax127x) & (ax125x) & (!g3) & (!g7)) + ((!ax124x) & (ax126x) & (!ax127x) & (ax125x) & (!g3) & (g7)) + ((!ax124x) & (ax126x) & (ax127x) & (!ax125x) & (!g3) & (!g7)) + ((!ax124x) & (ax126x) & (ax127x) & (!ax125x) & (!g3) & (g7)) + ((!ax124x) & (ax126x) & (ax127x) & (ax125x) & (g3) & (!g7)) + ((ax124x) & (!ax126x) & (!ax127x) & (!ax125x) & (!g3) & (!g7)) + ((ax124x) & (!ax126x) & (!ax127x) & (!ax125x) & (g3) & (!g7)) + ((ax124x) & (!ax126x) & (!ax127x) & (ax125x) & (g3) & (!g7)) + ((ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (!g3) & (!g7)) + ((ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (!g3) & (g7)) + ((ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (g3) & (!g7)) + ((ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (g3) & (g7)) + ((ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (!g3) & (!g7)) + ((ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (g3) & (!g7)) + ((ax124x) & (ax126x) & (!ax127x) & (ax125x) & (!g3) & (!g7)) + ((ax124x) & (ax126x) & (!ax127x) & (ax125x) & (g3) & (!g7)) + ((ax124x) & (ax126x) & (!ax127x) & (ax125x) & (g3) & (g7)) + ((ax124x) & (ax126x) & (ax127x) & (!ax125x) & (!g3) & (!g7)) + ((ax124x) & (ax126x) & (ax127x) & (!ax125x) & (g3) & (!g7)) + ((ax124x) & (ax126x) & (ax127x) & (!ax125x) & (g3) & (g7)));
	assign g9 = (((!g4) & (!ax122x) & (!g2) & (!g5) & (!g6)) + ((!g4) & (!ax122x) & (!g2) & (g5) & (!g6)) + ((!g4) & (!ax122x) & (!g2) & (g5) & (g6)) + ((!g4) & (!ax122x) & (g2) & (!g5) & (!g6)) + ((!g4) & (!ax122x) & (g2) & (g5) & (!g6)) + ((!g4) & (!ax122x) & (g2) & (g5) & (g6)) + ((!g4) & (ax122x) & (!g2) & (!g5) & (!g6)) + ((!g4) & (ax122x) & (!g2) & (!g5) & (g6)) + ((!g4) & (ax122x) & (!g2) & (g5) & (!g6)) + ((!g4) & (ax122x) & (!g2) & (g5) & (g6)) + ((!g4) & (ax122x) & (g2) & (!g5) & (!g6)) + ((!g4) & (ax122x) & (g2) & (g5) & (!g6)) + ((g4) & (!ax122x) & (!g2) & (!g5) & (!g6)) + ((g4) & (!ax122x) & (g2) & (!g5) & (!g6)) + ((g4) & (ax122x) & (g2) & (!g5) & (!g6)) + ((g4) & (ax122x) & (g2) & (g5) & (!g6)));
	assign g10 = (((!ax122x) & (!ax123x) & (!g2) & (!g8) & (!g9)) + ((!ax122x) & (!ax123x) & (!g2) & (g8) & (!g9)) + ((!ax122x) & (!ax123x) & (!g2) & (g8) & (g9)) + ((!ax122x) & (!ax123x) & (g2) & (!g8) & (g9)) + ((!ax122x) & (ax123x) & (!g2) & (!g8) & (g9)) + ((!ax122x) & (ax123x) & (g2) & (!g8) & (!g9)) + ((!ax122x) & (ax123x) & (g2) & (g8) & (!g9)) + ((!ax122x) & (ax123x) & (g2) & (g8) & (g9)) + ((ax122x) & (!ax123x) & (!g2) & (!g8) & (g9)) + ((ax122x) & (!ax123x) & (g2) & (!g8) & (g9)) + ((ax122x) & (ax123x) & (!g2) & (!g8) & (!g9)) + ((ax122x) & (ax123x) & (!g2) & (g8) & (!g9)) + ((ax122x) & (ax123x) & (!g2) & (g8) & (g9)) + ((ax122x) & (ax123x) & (g2) & (!g8) & (!g9)) + ((ax122x) & (ax123x) & (g2) & (g8) & (!g9)) + ((ax122x) & (ax123x) & (g2) & (g8) & (g9)));
	assign g11 = (((!ax118x) & (!ax119x)));
	assign g12 = (((!ax120x) & (!ax121x) & (!g2) & (!g8) & (!g11)) + ((!ax120x) & (!ax121x) & (g2) & (!g8) & (!g11)) + ((!ax120x) & (!ax121x) & (g2) & (!g8) & (g11)) + ((!ax120x) & (!ax121x) & (g2) & (g8) & (!g11)) + ((!ax120x) & (ax121x) & (!g2) & (g8) & (!g11)) + ((!ax120x) & (ax121x) & (g2) & (!g8) & (!g11)) + ((!ax120x) & (ax121x) & (g2) & (g8) & (!g11)) + ((!ax120x) & (ax121x) & (g2) & (g8) & (g11)) + ((ax120x) & (!ax121x) & (g2) & (g8) & (!g11)) + ((ax120x) & (!ax121x) & (g2) & (g8) & (g11)) + ((ax120x) & (ax121x) & (!g2) & (g8) & (!g11)) + ((ax120x) & (ax121x) & (!g2) & (g8) & (g11)) + ((ax120x) & (ax121x) & (g2) & (!g8) & (!g11)) + ((ax120x) & (ax121x) & (g2) & (!g8) & (g11)) + ((ax120x) & (ax121x) & (g2) & (g8) & (!g11)) + ((ax120x) & (ax121x) & (g2) & (g8) & (g11)));
	assign g13 = (((!ax122x) & (!g2) & (!g5) & (g8)) + ((!ax122x) & (!g2) & (g5) & (!g8)) + ((!ax122x) & (!g2) & (g5) & (g8)) + ((!ax122x) & (g2) & (g5) & (!g8)) + ((ax122x) & (!g2) & (!g5) & (!g8)) + ((ax122x) & (g2) & (!g5) & (!g8)) + ((ax122x) & (g2) & (!g5) & (g8)) + ((ax122x) & (g2) & (g5) & (g8)));
	assign g14 = (((!ax124x) & (!ax126x) & (!ax127x) & (ax125x) & (g3) & (g7)) + ((!ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (!g3) & (!g7)) + ((!ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (g3) & (g7)) + ((!ax124x) & (!ax126x) & (ax127x) & (ax125x) & (!g3) & (g7)) + ((!ax124x) & (!ax126x) & (ax127x) & (ax125x) & (g3) & (g7)) + ((!ax124x) & (ax126x) & (!ax127x) & (ax125x) & (g3) & (!g7)) + ((!ax124x) & (ax126x) & (ax127x) & (!ax125x) & (g3) & (g7)) + ((!ax124x) & (ax126x) & (ax127x) & (ax125x) & (!g3) & (!g7)) + ((!ax124x) & (ax126x) & (ax127x) & (ax125x) & (g3) & (g7)) + ((ax124x) & (!ax126x) & (!ax127x) & (ax125x) & (!g3) & (g7)) + ((ax124x) & (!ax126x) & (ax127x) & (ax125x) & (!g3) & (!g7)) + ((ax124x) & (!ax126x) & (ax127x) & (ax125x) & (g3) & (!g7)) + ((ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (!g3) & (g7)) + ((ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (g3) & (g7)) + ((ax124x) & (ax126x) & (!ax127x) & (ax125x) & (!g3) & (g7)) + ((ax124x) & (ax126x) & (ax127x) & (!ax125x) & (!g3) & (g7)) + ((ax124x) & (ax126x) & (ax127x) & (ax125x) & (!g3) & (g7)) + ((ax124x) & (ax126x) & (ax127x) & (ax125x) & (g3) & (!g7)));
	assign g15 = (((!g4) & (!g1) & (!g10) & (!g12) & (!g13) & (g14)) + ((!g4) & (!g1) & (!g10) & (!g12) & (g13) & (!g14)) + ((!g4) & (!g1) & (!g10) & (!g12) & (g13) & (g14)) + ((!g4) & (!g1) & (!g10) & (g12) & (!g13) & (!g14)) + ((!g4) & (!g1) & (!g10) & (g12) & (!g13) & (g14)) + ((!g4) & (!g1) & (!g10) & (g12) & (g13) & (!g14)) + ((!g4) & (!g1) & (!g10) & (g12) & (g13) & (g14)) + ((!g4) & (!g1) & (g10) & (!g12) & (!g13) & (!g14)) + ((!g4) & (!g1) & (g10) & (!g12) & (!g13) & (g14)) + ((!g4) & (!g1) & (g10) & (!g12) & (g13) & (!g14)) + ((!g4) & (!g1) & (g10) & (!g12) & (g13) & (g14)) + ((!g4) & (!g1) & (g10) & (g12) & (!g13) & (!g14)) + ((!g4) & (!g1) & (g10) & (g12) & (!g13) & (g14)) + ((!g4) & (!g1) & (g10) & (g12) & (g13) & (!g14)) + ((!g4) & (!g1) & (g10) & (g12) & (g13) & (g14)) + ((g4) & (!g1) & (!g10) & (!g12) & (!g13) & (g14)) + ((g4) & (!g1) & (!g10) & (!g12) & (g13) & (g14)) + ((g4) & (!g1) & (!g10) & (g12) & (!g13) & (g14)) + ((g4) & (!g1) & (!g10) & (g12) & (g13) & (!g14)) + ((g4) & (!g1) & (!g10) & (g12) & (g13) & (g14)) + ((g4) & (!g1) & (g10) & (!g12) & (!g13) & (!g14)) + ((g4) & (!g1) & (g10) & (!g12) & (!g13) & (g14)) + ((g4) & (!g1) & (g10) & (!g12) & (g13) & (!g14)) + ((g4) & (!g1) & (g10) & (!g12) & (g13) & (g14)) + ((g4) & (!g1) & (g10) & (g12) & (!g13) & (!g14)) + ((g4) & (!g1) & (g10) & (g12) & (!g13) & (g14)) + ((g4) & (!g1) & (g10) & (g12) & (g13) & (!g14)) + ((g4) & (!g1) & (g10) & (g12) & (g13) & (g14)));
	assign g16 = (((!ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (!g3) & (g7)) + ((!ax124x) & (!ax126x) & (ax127x) & (!ax125x) & (g3) & (!g7)) + ((!ax124x) & (!ax126x) & (ax127x) & (ax125x) & (!g3) & (!g7)) + ((!ax124x) & (!ax126x) & (ax127x) & (ax125x) & (g3) & (!g7)) + ((!ax124x) & (ax126x) & (!ax127x) & (ax125x) & (g3) & (g7)) + ((!ax124x) & (ax126x) & (ax127x) & (!ax125x) & (g3) & (!g7)) + ((!ax124x) & (ax126x) & (ax127x) & (ax125x) & (!g3) & (g7)) + ((!ax124x) & (ax126x) & (ax127x) & (ax125x) & (g3) & (!g7)) + ((ax124x) & (!ax126x) & (ax127x) & (ax125x) & (!g3) & (g7)) + ((ax124x) & (!ax126x) & (ax127x) & (ax125x) & (g3) & (g7)) + ((ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (!g3) & (!g7)) + ((ax124x) & (ax126x) & (!ax127x) & (!ax125x) & (g3) & (!g7)) + ((ax124x) & (ax126x) & (!ax127x) & (ax125x) & (!g3) & (!g7)) + ((ax124x) & (ax126x) & (ax127x) & (!ax125x) & (!g3) & (!g7)) + ((ax124x) & (ax126x) & (ax127x) & (ax125x) & (!g3) & (!g7)) + ((ax124x) & (ax126x) & (ax127x) & (ax125x) & (g3) & (g7)));
	assign g17 = (((!g4) & (!g10) & (!g12) & (!g13) & (!g16)) + ((!g4) & (!g10) & (!g12) & (g13) & (!g16)) + ((!g4) & (!g10) & (g12) & (!g13) & (!g16)) + ((!g4) & (!g10) & (g12) & (g13) & (!g16)) + ((!g4) & (g10) & (!g12) & (!g13) & (!g16)) + ((g4) & (!g10) & (!g12) & (!g13) & (!g16)) + ((g4) & (!g10) & (!g12) & (g13) & (!g16)) + ((g4) & (!g10) & (g12) & (!g13) & (!g16)) + ((g4) & (!g10) & (g12) & (g13) & (!g16)) + ((g4) & (g10) & (!g12) & (!g13) & (!g16)) + ((g4) & (g10) & (!g12) & (g13) & (!g16)) + ((g4) & (g10) & (g12) & (!g13) & (!g16)));
	assign g18 = (((!g15) & (g17)));
	assign g19 = (((!g4) & (!g12) & (g13)) + ((!g4) & (g12) & (!g13)) + ((!g4) & (g12) & (g13)) + ((g4) & (g12) & (g13)));
	assign g20 = (((!g4) & (!g12) & (!g13) & (!g15) & (!g17)) + ((!g4) & (!g12) & (!g13) & (g15) & (!g17)) + ((!g4) & (!g12) & (!g13) & (g15) & (g17)) + ((!g4) & (!g12) & (g13) & (!g15) & (g17)) + ((!g4) & (g12) & (g13) & (!g15) & (!g17)) + ((!g4) & (g12) & (g13) & (!g15) & (g17)) + ((!g4) & (g12) & (g13) & (g15) & (!g17)) + ((!g4) & (g12) & (g13) & (g15) & (g17)) + ((g4) & (!g12) & (g13) & (!g15) & (!g17)) + ((g4) & (!g12) & (g13) & (!g15) & (g17)) + ((g4) & (!g12) & (g13) & (g15) & (!g17)) + ((g4) & (!g12) & (g13) & (g15) & (g17)) + ((g4) & (g12) & (!g13) & (!g15) & (!g17)) + ((g4) & (g12) & (!g13) & (g15) & (!g17)) + ((g4) & (g12) & (!g13) & (g15) & (g17)) + ((g4) & (g12) & (g13) & (!g15) & (g17)));
	assign g21 = (((!ax120x) & (!g2) & (!g8) & (!g11)) + ((!ax120x) & (!g2) & (g8) & (!g11)) + ((!ax120x) & (g2) & (!g8) & (g11)) + ((!ax120x) & (g2) & (g8) & (g11)) + ((ax120x) & (!g2) & (g8) & (!g11)) + ((ax120x) & (!g2) & (g8) & (g11)) + ((ax120x) & (g2) & (!g8) & (!g11)) + ((ax120x) & (g2) & (!g8) & (g11)));
	assign g22 = (((!ax120x) & (!ax121x) & (!g8) & (!g15) & (!g17) & (!g21)) + ((!ax120x) & (!ax121x) & (!g8) & (!g15) & (g17) & (!g21)) + ((!ax120x) & (!ax121x) & (!g8) & (!g15) & (g17) & (g21)) + ((!ax120x) & (!ax121x) & (!g8) & (g15) & (!g17) & (!g21)) + ((!ax120x) & (!ax121x) & (!g8) & (g15) & (g17) & (!g21)) + ((!ax120x) & (!ax121x) & (g8) & (!g15) & (!g17) & (g21)) + ((!ax120x) & (!ax121x) & (g8) & (g15) & (!g17) & (g21)) + ((!ax120x) & (!ax121x) & (g8) & (g15) & (g17) & (g21)) + ((!ax120x) & (ax121x) & (!g8) & (!g15) & (!g17) & (g21)) + ((!ax120x) & (ax121x) & (!g8) & (g15) & (!g17) & (g21)) + ((!ax120x) & (ax121x) & (!g8) & (g15) & (g17) & (g21)) + ((!ax120x) & (ax121x) & (g8) & (!g15) & (!g17) & (!g21)) + ((!ax120x) & (ax121x) & (g8) & (!g15) & (g17) & (!g21)) + ((!ax120x) & (ax121x) & (g8) & (!g15) & (g17) & (g21)) + ((!ax120x) & (ax121x) & (g8) & (g15) & (!g17) & (!g21)) + ((!ax120x) & (ax121x) & (g8) & (g15) & (g17) & (!g21)) + ((ax120x) & (!ax121x) & (!g8) & (!g15) & (!g17) & (g21)) + ((ax120x) & (!ax121x) & (!g8) & (g15) & (!g17) & (g21)) + ((ax120x) & (!ax121x) & (!g8) & (g15) & (g17) & (g21)) + ((ax120x) & (!ax121x) & (g8) & (!g15) & (!g17) & (g21)) + ((ax120x) & (!ax121x) & (g8) & (g15) & (!g17) & (g21)) + ((ax120x) & (!ax121x) & (g8) & (g15) & (g17) & (g21)) + ((ax120x) & (ax121x) & (!g8) & (!g15) & (!g17) & (!g21)) + ((ax120x) & (ax121x) & (!g8) & (!g15) & (g17) & (!g21)) + ((ax120x) & (ax121x) & (!g8) & (!g15) & (g17) & (g21)) + ((ax120x) & (ax121x) & (!g8) & (g15) & (!g17) & (!g21)) + ((ax120x) & (ax121x) & (!g8) & (g15) & (g17) & (!g21)) + ((ax120x) & (ax121x) & (g8) & (!g15) & (!g17) & (!g21)) + ((ax120x) & (ax121x) & (g8) & (!g15) & (g17) & (!g21)) + ((ax120x) & (ax121x) & (g8) & (!g15) & (g17) & (g21)) + ((ax120x) & (ax121x) & (g8) & (g15) & (!g17) & (!g21)) + ((ax120x) & (ax121x) & (g8) & (g15) & (g17) & (!g21)));
	assign g23 = (((!ax120x) & (!g8) & (!g11) & (!g15) & (g17)) + ((!ax120x) & (!g8) & (g11) & (!g15) & (!g17)) + ((!ax120x) & (!g8) & (g11) & (!g15) & (g17)) + ((!ax120x) & (!g8) & (g11) & (g15) & (!g17)) + ((!ax120x) & (!g8) & (g11) & (g15) & (g17)) + ((!ax120x) & (g8) & (g11) & (!g15) & (!g17)) + ((!ax120x) & (g8) & (g11) & (g15) & (!g17)) + ((!ax120x) & (g8) & (g11) & (g15) & (g17)) + ((ax120x) & (!g8) & (!g11) & (!g15) & (!g17)) + ((ax120x) & (!g8) & (!g11) & (g15) & (!g17)) + ((ax120x) & (!g8) & (!g11) & (g15) & (g17)) + ((ax120x) & (g8) & (!g11) & (!g15) & (!g17)) + ((ax120x) & (g8) & (!g11) & (!g15) & (g17)) + ((ax120x) & (g8) & (!g11) & (g15) & (!g17)) + ((ax120x) & (g8) & (!g11) & (g15) & (g17)) + ((ax120x) & (g8) & (g11) & (!g15) & (g17)));
	assign g24 = (((!ax116x) & (!ax117x)));
	assign g25 = (((!g8) & (!ax118x) & (!ax119x) & (!g15) & (!g17) & (!g24)) + ((!g8) & (!ax118x) & (!ax119x) & (g15) & (!g17) & (!g24)) + ((!g8) & (!ax118x) & (!ax119x) & (g15) & (g17) & (!g24)) + ((!g8) & (!ax118x) & (ax119x) & (!g15) & (g17) & (!g24)) + ((!g8) & (ax118x) & (ax119x) & (!g15) & (g17) & (!g24)) + ((!g8) & (ax118x) & (ax119x) & (!g15) & (g17) & (g24)) + ((g8) & (!ax118x) & (!ax119x) & (!g15) & (!g17) & (!g24)) + ((g8) & (!ax118x) & (!ax119x) & (!g15) & (!g17) & (g24)) + ((g8) & (!ax118x) & (!ax119x) & (!g15) & (g17) & (!g24)) + ((g8) & (!ax118x) & (!ax119x) & (g15) & (!g17) & (!g24)) + ((g8) & (!ax118x) & (!ax119x) & (g15) & (!g17) & (g24)) + ((g8) & (!ax118x) & (!ax119x) & (g15) & (g17) & (!g24)) + ((g8) & (!ax118x) & (!ax119x) & (g15) & (g17) & (g24)) + ((g8) & (!ax118x) & (ax119x) & (!g15) & (!g17) & (!g24)) + ((g8) & (!ax118x) & (ax119x) & (!g15) & (g17) & (!g24)) + ((g8) & (!ax118x) & (ax119x) & (!g15) & (g17) & (g24)) + ((g8) & (!ax118x) & (ax119x) & (g15) & (!g17) & (!g24)) + ((g8) & (!ax118x) & (ax119x) & (g15) & (g17) & (!g24)) + ((g8) & (ax118x) & (!ax119x) & (!g15) & (g17) & (!g24)) + ((g8) & (ax118x) & (!ax119x) & (!g15) & (g17) & (g24)) + ((g8) & (ax118x) & (ax119x) & (!g15) & (!g17) & (!g24)) + ((g8) & (ax118x) & (ax119x) & (!g15) & (!g17) & (g24)) + ((g8) & (ax118x) & (ax119x) & (!g15) & (g17) & (!g24)) + ((g8) & (ax118x) & (ax119x) & (!g15) & (g17) & (g24)) + ((g8) & (ax118x) & (ax119x) & (g15) & (!g17) & (!g24)) + ((g8) & (ax118x) & (ax119x) & (g15) & (!g17) & (g24)) + ((g8) & (ax118x) & (ax119x) & (g15) & (g17) & (!g24)) + ((g8) & (ax118x) & (ax119x) & (g15) & (g17) & (g24)));
	assign g26 = (((!g4) & (!g2) & (!g22) & (g23) & (g25)) + ((!g4) & (!g2) & (g22) & (!g23) & (!g25)) + ((!g4) & (!g2) & (g22) & (!g23) & (g25)) + ((!g4) & (!g2) & (g22) & (g23) & (!g25)) + ((!g4) & (!g2) & (g22) & (g23) & (g25)) + ((!g4) & (g2) & (!g22) & (!g23) & (g25)) + ((!g4) & (g2) & (!g22) & (g23) & (!g25)) + ((!g4) & (g2) & (!g22) & (g23) & (g25)) + ((!g4) & (g2) & (g22) & (!g23) & (!g25)) + ((!g4) & (g2) & (g22) & (!g23) & (g25)) + ((!g4) & (g2) & (g22) & (g23) & (!g25)) + ((!g4) & (g2) & (g22) & (g23) & (g25)) + ((g4) & (!g2) & (g22) & (g23) & (g25)) + ((g4) & (g2) & (g22) & (!g23) & (g25)) + ((g4) & (g2) & (g22) & (g23) & (!g25)) + ((g4) & (g2) & (g22) & (g23) & (g25)));
	assign g27 = (((!g1) & (!g10) & (!g19) & (g18) & (!g20) & (!g26)) + ((!g1) & (!g10) & (g19) & (!g18) & (!g20) & (!g26)) + ((!g1) & (!g10) & (g19) & (g18) & (!g20) & (!g26)) + ((!g1) & (g10) & (!g19) & (!g18) & (!g20) & (!g26)) + ((g1) & (!g10) & (!g19) & (!g18) & (!g20) & (!g26)) + ((g1) & (!g10) & (!g19) & (!g18) & (!g20) & (g26)) + ((g1) & (!g10) & (!g19) & (!g18) & (g20) & (!g26)) + ((g1) & (!g10) & (!g19) & (g18) & (!g20) & (!g26)) + ((g1) & (!g10) & (!g19) & (g18) & (!g20) & (g26)) + ((g1) & (!g10) & (!g19) & (g18) & (g20) & (!g26)) + ((g1) & (!g10) & (g19) & (g18) & (!g20) & (!g26)) + ((g1) & (!g10) & (g19) & (g18) & (!g20) & (g26)) + ((g1) & (!g10) & (g19) & (g18) & (g20) & (!g26)) + ((g1) & (g10) & (g19) & (!g18) & (!g20) & (!g26)) + ((g1) & (g10) & (g19) & (!g18) & (!g20) & (g26)) + ((g1) & (g10) & (g19) & (!g18) & (g20) & (!g26)));
	assign g28 = (((!g4) & (!g2) & (!g22) & (!g23) & (!g25) & (!g27)) + ((!g4) & (!g2) & (!g22) & (!g23) & (g25) & (!g27)) + ((!g4) & (!g2) & (!g22) & (g23) & (!g25) & (!g27)) + ((!g4) & (!g2) & (g22) & (!g23) & (!g25) & (g27)) + ((!g4) & (!g2) & (g22) & (!g23) & (g25) & (g27)) + ((!g4) & (!g2) & (g22) & (g23) & (!g25) & (g27)) + ((!g4) & (!g2) & (g22) & (g23) & (g25) & (!g27)) + ((!g4) & (!g2) & (g22) & (g23) & (g25) & (g27)) + ((!g4) & (g2) & (!g22) & (!g23) & (!g25) & (!g27)) + ((!g4) & (g2) & (g22) & (!g23) & (!g25) & (g27)) + ((!g4) & (g2) & (g22) & (!g23) & (g25) & (!g27)) + ((!g4) & (g2) & (g22) & (!g23) & (g25) & (g27)) + ((!g4) & (g2) & (g22) & (g23) & (!g25) & (!g27)) + ((!g4) & (g2) & (g22) & (g23) & (!g25) & (g27)) + ((!g4) & (g2) & (g22) & (g23) & (g25) & (!g27)) + ((!g4) & (g2) & (g22) & (g23) & (g25) & (g27)) + ((g4) & (!g2) & (!g22) & (g23) & (g25) & (!g27)) + ((g4) & (!g2) & (g22) & (!g23) & (!g25) & (!g27)) + ((g4) & (!g2) & (g22) & (!g23) & (!g25) & (g27)) + ((g4) & (!g2) & (g22) & (!g23) & (g25) & (!g27)) + ((g4) & (!g2) & (g22) & (!g23) & (g25) & (g27)) + ((g4) & (!g2) & (g22) & (g23) & (!g25) & (!g27)) + ((g4) & (!g2) & (g22) & (g23) & (!g25) & (g27)) + ((g4) & (!g2) & (g22) & (g23) & (g25) & (g27)) + ((g4) & (g2) & (!g22) & (!g23) & (g25) & (!g27)) + ((g4) & (g2) & (!g22) & (g23) & (!g25) & (!g27)) + ((g4) & (g2) & (!g22) & (g23) & (g25) & (!g27)) + ((g4) & (g2) & (g22) & (!g23) & (!g25) & (!g27)) + ((g4) & (g2) & (g22) & (!g23) & (!g25) & (g27)) + ((g4) & (g2) & (g22) & (!g23) & (g25) & (g27)) + ((g4) & (g2) & (g22) & (g23) & (!g25) & (g27)) + ((g4) & (g2) & (g22) & (g23) & (g25) & (g27)));
	assign g29 = (((!g8) & (!ax118x) & (!ax119x) & (!g18) & (!g24) & (g27)) + ((!g8) & (!ax118x) & (!ax119x) & (!g18) & (g24) & (!g27)) + ((!g8) & (!ax118x) & (!ax119x) & (!g18) & (g24) & (g27)) + ((!g8) & (!ax118x) & (!ax119x) & (g18) & (!g24) & (!g27)) + ((!g8) & (!ax118x) & (ax119x) & (!g18) & (!g24) & (!g27)) + ((!g8) & (!ax118x) & (ax119x) & (g18) & (!g24) & (g27)) + ((!g8) & (!ax118x) & (ax119x) & (g18) & (g24) & (!g27)) + ((!g8) & (!ax118x) & (ax119x) & (g18) & (g24) & (g27)) + ((!g8) & (ax118x) & (!ax119x) & (g18) & (!g24) & (!g27)) + ((!g8) & (ax118x) & (!ax119x) & (g18) & (g24) & (!g27)) + ((!g8) & (ax118x) & (ax119x) & (!g18) & (!g24) & (!g27)) + ((!g8) & (ax118x) & (ax119x) & (!g18) & (!g24) & (g27)) + ((!g8) & (ax118x) & (ax119x) & (!g18) & (g24) & (!g27)) + ((!g8) & (ax118x) & (ax119x) & (!g18) & (g24) & (g27)) + ((!g8) & (ax118x) & (ax119x) & (g18) & (!g24) & (g27)) + ((!g8) & (ax118x) & (ax119x) & (g18) & (g24) & (g27)) + ((g8) & (!ax118x) & (!ax119x) & (!g18) & (!g24) & (!g27)) + ((g8) & (!ax118x) & (!ax119x) & (!g18) & (!g24) & (g27)) + ((g8) & (!ax118x) & (!ax119x) & (!g18) & (g24) & (g27)) + ((g8) & (!ax118x) & (!ax119x) & (g18) & (g24) & (!g27)) + ((g8) & (!ax118x) & (ax119x) & (!g18) & (g24) & (!g27)) + ((g8) & (!ax118x) & (ax119x) & (g18) & (!g24) & (!g27)) + ((g8) & (!ax118x) & (ax119x) & (g18) & (!g24) & (g27)) + ((g8) & (!ax118x) & (ax119x) & (g18) & (g24) & (g27)) + ((g8) & (ax118x) & (!ax119x) & (!g18) & (!g24) & (!g27)) + ((g8) & (ax118x) & (!ax119x) & (!g18) & (g24) & (!g27)) + ((g8) & (ax118x) & (ax119x) & (!g18) & (!g24) & (g27)) + ((g8) & (ax118x) & (ax119x) & (!g18) & (g24) & (g27)) + ((g8) & (ax118x) & (ax119x) & (g18) & (!g24) & (!g27)) + ((g8) & (ax118x) & (ax119x) & (g18) & (!g24) & (g27)) + ((g8) & (ax118x) & (ax119x) & (g18) & (g24) & (!g27)) + ((g8) & (ax118x) & (ax119x) & (g18) & (g24) & (g27)));
	assign g30 = (((!ax118x) & (!g18) & (!g24) & (g27)) + ((!ax118x) & (!g18) & (g24) & (!g27)) + ((!ax118x) & (!g18) & (g24) & (g27)) + ((!ax118x) & (g18) & (g24) & (!g27)) + ((ax118x) & (!g18) & (!g24) & (!g27)) + ((ax118x) & (g18) & (!g24) & (!g27)) + ((ax118x) & (g18) & (!g24) & (g27)) + ((ax118x) & (g18) & (g24) & (g27)));
	assign g31 = (((!ax114x) & (!ax115x)));
	assign g32 = (((!g18) & (!ax116x) & (!ax117x) & (!g27) & (!g31)) + ((!g18) & (!ax116x) & (ax117x) & (g27) & (!g31)) + ((!g18) & (ax116x) & (ax117x) & (g27) & (!g31)) + ((!g18) & (ax116x) & (ax117x) & (g27) & (g31)) + ((g18) & (!ax116x) & (!ax117x) & (!g27) & (!g31)) + ((g18) & (!ax116x) & (!ax117x) & (!g27) & (g31)) + ((g18) & (!ax116x) & (!ax117x) & (g27) & (!g31)) + ((g18) & (!ax116x) & (ax117x) & (!g27) & (!g31)) + ((g18) & (!ax116x) & (ax117x) & (g27) & (!g31)) + ((g18) & (!ax116x) & (ax117x) & (g27) & (g31)) + ((g18) & (ax116x) & (!ax117x) & (g27) & (!g31)) + ((g18) & (ax116x) & (!ax117x) & (g27) & (g31)) + ((g18) & (ax116x) & (ax117x) & (!g27) & (!g31)) + ((g18) & (ax116x) & (ax117x) & (!g27) & (g31)) + ((g18) & (ax116x) & (ax117x) & (g27) & (!g31)) + ((g18) & (ax116x) & (ax117x) & (g27) & (g31)));
	assign g33 = (((!g2) & (!g8) & (g29) & (g30) & (g32)) + ((!g2) & (g8) & (g29) & (!g30) & (g32)) + ((!g2) & (g8) & (g29) & (g30) & (!g32)) + ((!g2) & (g8) & (g29) & (g30) & (g32)) + ((g2) & (!g8) & (!g29) & (g30) & (g32)) + ((g2) & (!g8) & (g29) & (!g30) & (!g32)) + ((g2) & (!g8) & (g29) & (!g30) & (g32)) + ((g2) & (!g8) & (g29) & (g30) & (!g32)) + ((g2) & (!g8) & (g29) & (g30) & (g32)) + ((g2) & (g8) & (!g29) & (!g30) & (g32)) + ((g2) & (g8) & (!g29) & (g30) & (!g32)) + ((g2) & (g8) & (!g29) & (g30) & (g32)) + ((g2) & (g8) & (g29) & (!g30) & (!g32)) + ((g2) & (g8) & (g29) & (!g30) & (g32)) + ((g2) & (g8) & (g29) & (g30) & (!g32)) + ((g2) & (g8) & (g29) & (g30) & (g32)));
	assign g34 = (((!g2) & (!g23) & (g25) & (!g27)) + ((!g2) & (g23) & (!g25) & (!g27)) + ((!g2) & (g23) & (!g25) & (g27)) + ((!g2) & (g23) & (g25) & (g27)) + ((g2) & (!g23) & (!g25) & (!g27)) + ((g2) & (g23) & (!g25) & (g27)) + ((g2) & (g23) & (g25) & (!g27)) + ((g2) & (g23) & (g25) & (g27)));
	assign g35 = (((!g1) & (!g10) & (!g19) & (!g18) & (!g20) & (!g26)) + ((!g1) & (!g10) & (!g19) & (!g18) & (g20) & (g26)) + ((!g1) & (!g10) & (!g19) & (g18) & (g20) & (g26)) + ((!g1) & (!g10) & (g19) & (!g18) & (g20) & (g26)) + ((!g1) & (!g10) & (g19) & (g18) & (g20) & (g26)) + ((!g1) & (g10) & (!g19) & (!g18) & (g20) & (g26)) + ((!g1) & (g10) & (!g19) & (g18) & (!g20) & (!g26)) + ((!g1) & (g10) & (!g19) & (g18) & (g20) & (g26)) + ((!g1) & (g10) & (g19) & (!g18) & (!g20) & (!g26)) + ((!g1) & (g10) & (g19) & (!g18) & (g20) & (g26)) + ((!g1) & (g10) & (g19) & (g18) & (!g20) & (!g26)) + ((!g1) & (g10) & (g19) & (g18) & (g20) & (g26)) + ((g1) & (!g10) & (!g19) & (!g18) & (g20) & (g26)) + ((g1) & (!g10) & (!g19) & (g18) & (g20) & (g26)) + ((g1) & (!g10) & (g19) & (!g18) & (!g20) & (!g26)) + ((g1) & (!g10) & (g19) & (!g18) & (g20) & (g26)) + ((g1) & (!g10) & (g19) & (g18) & (g20) & (g26)) + ((g1) & (g10) & (!g19) & (!g18) & (!g20) & (!g26)) + ((g1) & (g10) & (!g19) & (!g18) & (g20) & (g26)) + ((g1) & (g10) & (!g19) & (g18) & (!g20) & (!g26)) + ((g1) & (g10) & (!g19) & (g18) & (g20) & (g26)) + ((g1) & (g10) & (g19) & (!g18) & (g20) & (g26)) + ((g1) & (g10) & (g19) & (g18) & (!g20) & (!g26)) + ((g1) & (g10) & (g19) & (g18) & (g20) & (g26)));
	assign g36 = (((!g4) & (!g1) & (!g28) & (!g33) & (!g34) & (g35)) + ((!g4) & (!g1) & (!g28) & (!g33) & (g34) & (!g35)) + ((!g4) & (!g1) & (!g28) & (!g33) & (g34) & (g35)) + ((!g4) & (!g1) & (!g28) & (g33) & (!g34) & (!g35)) + ((!g4) & (!g1) & (!g28) & (g33) & (!g34) & (g35)) + ((!g4) & (!g1) & (!g28) & (g33) & (g34) & (!g35)) + ((!g4) & (!g1) & (!g28) & (g33) & (g34) & (g35)) + ((!g4) & (!g1) & (g28) & (!g33) & (!g34) & (!g35)) + ((!g4) & (!g1) & (g28) & (!g33) & (!g34) & (g35)) + ((!g4) & (!g1) & (g28) & (!g33) & (g34) & (!g35)) + ((!g4) & (!g1) & (g28) & (!g33) & (g34) & (g35)) + ((!g4) & (!g1) & (g28) & (g33) & (!g34) & (!g35)) + ((!g4) & (!g1) & (g28) & (g33) & (!g34) & (g35)) + ((!g4) & (!g1) & (g28) & (g33) & (g34) & (!g35)) + ((!g4) & (!g1) & (g28) & (g33) & (g34) & (g35)) + ((g4) & (!g1) & (!g28) & (!g33) & (!g34) & (g35)) + ((g4) & (!g1) & (!g28) & (!g33) & (g34) & (g35)) + ((g4) & (!g1) & (!g28) & (g33) & (!g34) & (g35)) + ((g4) & (!g1) & (!g28) & (g33) & (g34) & (!g35)) + ((g4) & (!g1) & (!g28) & (g33) & (g34) & (g35)) + ((g4) & (!g1) & (g28) & (!g33) & (!g34) & (!g35)) + ((g4) & (!g1) & (g28) & (!g33) & (!g34) & (g35)) + ((g4) & (!g1) & (g28) & (!g33) & (g34) & (!g35)) + ((g4) & (!g1) & (g28) & (!g33) & (g34) & (g35)) + ((g4) & (!g1) & (g28) & (g33) & (!g34) & (!g35)) + ((g4) & (!g1) & (g28) & (g33) & (!g34) & (g35)) + ((g4) & (!g1) & (g28) & (g33) & (g34) & (!g35)) + ((g4) & (!g1) & (g28) & (g33) & (g34) & (g35)));
	assign g37 = (((g1) & (!g10) & (!g19) & (!g18) & (g20) & (!g26)) + ((g1) & (!g10) & (!g19) & (g18) & (g20) & (!g26)) + ((g1) & (!g10) & (g19) & (!g18) & (!g20) & (g26)) + ((g1) & (!g10) & (g19) & (!g18) & (g20) & (!g26)) + ((g1) & (!g10) & (g19) & (g18) & (g20) & (!g26)) + ((g1) & (g10) & (!g19) & (!g18) & (!g20) & (g26)) + ((g1) & (g10) & (!g19) & (!g18) & (g20) & (!g26)) + ((g1) & (g10) & (!g19) & (g18) & (!g20) & (g26)) + ((g1) & (g10) & (!g19) & (g18) & (g20) & (!g26)) + ((g1) & (g10) & (g19) & (!g18) & (g20) & (!g26)) + ((g1) & (g10) & (g19) & (g18) & (!g20) & (g26)) + ((g1) & (g10) & (g19) & (g18) & (g20) & (!g26)));
	assign g38 = (((!g4) & (!g28) & (!g33) & (!g34) & (!g37)) + ((!g4) & (!g28) & (!g33) & (g34) & (!g37)) + ((!g4) & (!g28) & (g33) & (!g34) & (!g37)) + ((!g4) & (!g28) & (g33) & (g34) & (!g37)) + ((!g4) & (g28) & (!g33) & (!g34) & (!g37)) + ((g4) & (!g28) & (!g33) & (!g34) & (!g37)) + ((g4) & (!g28) & (!g33) & (g34) & (!g37)) + ((g4) & (!g28) & (g33) & (!g34) & (!g37)) + ((g4) & (!g28) & (g33) & (g34) & (!g37)) + ((g4) & (g28) & (!g33) & (!g34) & (!g37)) + ((g4) & (g28) & (!g33) & (g34) & (!g37)) + ((g4) & (g28) & (g33) & (!g34) & (!g37)));
	assign g39 = (((!g36) & (g38)));
	assign g40 = (((!g4) & (!g33) & (!g34) & (!g36) & (!g38)) + ((!g4) & (!g33) & (!g34) & (g36) & (!g38)) + ((!g4) & (!g33) & (!g34) & (g36) & (g38)) + ((!g4) & (!g33) & (g34) & (!g36) & (g38)) + ((!g4) & (g33) & (g34) & (!g36) & (!g38)) + ((!g4) & (g33) & (g34) & (!g36) & (g38)) + ((!g4) & (g33) & (g34) & (g36) & (!g38)) + ((!g4) & (g33) & (g34) & (g36) & (g38)) + ((g4) & (!g33) & (g34) & (!g36) & (!g38)) + ((g4) & (!g33) & (g34) & (!g36) & (g38)) + ((g4) & (!g33) & (g34) & (g36) & (!g38)) + ((g4) & (!g33) & (g34) & (g36) & (g38)) + ((g4) & (g33) & (!g34) & (!g36) & (!g38)) + ((g4) & (g33) & (!g34) & (g36) & (!g38)) + ((g4) & (g33) & (!g34) & (g36) & (g38)) + ((g4) & (g33) & (g34) & (!g36) & (g38)));
	assign g41 = (((!g8) & (!g30) & (g32) & (!g36) & (!g38)) + ((!g8) & (!g30) & (g32) & (g36) & (!g38)) + ((!g8) & (!g30) & (g32) & (g36) & (g38)) + ((!g8) & (g30) & (!g32) & (!g36) & (!g38)) + ((!g8) & (g30) & (!g32) & (!g36) & (g38)) + ((!g8) & (g30) & (!g32) & (g36) & (!g38)) + ((!g8) & (g30) & (!g32) & (g36) & (g38)) + ((!g8) & (g30) & (g32) & (!g36) & (g38)) + ((g8) & (!g30) & (!g32) & (!g36) & (!g38)) + ((g8) & (!g30) & (!g32) & (g36) & (!g38)) + ((g8) & (!g30) & (!g32) & (g36) & (g38)) + ((g8) & (g30) & (!g32) & (!g36) & (g38)) + ((g8) & (g30) & (g32) & (!g36) & (!g38)) + ((g8) & (g30) & (g32) & (!g36) & (g38)) + ((g8) & (g30) & (g32) & (g36) & (!g38)) + ((g8) & (g30) & (g32) & (g36) & (g38)));
	assign g42 = (((!g18) & (!ax116x) & (!g27) & (g31)) + ((!g18) & (!ax116x) & (g27) & (g31)) + ((!g18) & (ax116x) & (!g27) & (!g31)) + ((!g18) & (ax116x) & (!g27) & (g31)) + ((g18) & (!ax116x) & (!g27) & (!g31)) + ((g18) & (!ax116x) & (g27) & (!g31)) + ((g18) & (ax116x) & (g27) & (!g31)) + ((g18) & (ax116x) & (g27) & (g31)));
	assign g43 = (((!ax116x) & (!ax117x) & (!g27) & (!g36) & (!g38) & (g42)) + ((!ax116x) & (!ax117x) & (!g27) & (!g36) & (g38) & (!g42)) + ((!ax116x) & (!ax117x) & (!g27) & (!g36) & (g38) & (g42)) + ((!ax116x) & (!ax117x) & (!g27) & (g36) & (!g38) & (g42)) + ((!ax116x) & (!ax117x) & (!g27) & (g36) & (g38) & (g42)) + ((!ax116x) & (!ax117x) & (g27) & (!g36) & (!g38) & (!g42)) + ((!ax116x) & (!ax117x) & (g27) & (g36) & (!g38) & (!g42)) + ((!ax116x) & (!ax117x) & (g27) & (g36) & (g38) & (!g42)) + ((!ax116x) & (ax117x) & (!g27) & (!g36) & (!g38) & (!g42)) + ((!ax116x) & (ax117x) & (!g27) & (g36) & (!g38) & (!g42)) + ((!ax116x) & (ax117x) & (!g27) & (g36) & (g38) & (!g42)) + ((!ax116x) & (ax117x) & (g27) & (!g36) & (!g38) & (g42)) + ((!ax116x) & (ax117x) & (g27) & (!g36) & (g38) & (!g42)) + ((!ax116x) & (ax117x) & (g27) & (!g36) & (g38) & (g42)) + ((!ax116x) & (ax117x) & (g27) & (g36) & (!g38) & (g42)) + ((!ax116x) & (ax117x) & (g27) & (g36) & (g38) & (g42)) + ((ax116x) & (!ax117x) & (!g27) & (!g36) & (!g38) & (!g42)) + ((ax116x) & (!ax117x) & (!g27) & (g36) & (!g38) & (!g42)) + ((ax116x) & (!ax117x) & (!g27) & (g36) & (g38) & (!g42)) + ((ax116x) & (!ax117x) & (g27) & (!g36) & (!g38) & (!g42)) + ((ax116x) & (!ax117x) & (g27) & (g36) & (!g38) & (!g42)) + ((ax116x) & (!ax117x) & (g27) & (g36) & (g38) & (!g42)) + ((ax116x) & (ax117x) & (!g27) & (!g36) & (!g38) & (g42)) + ((ax116x) & (ax117x) & (!g27) & (!g36) & (g38) & (!g42)) + ((ax116x) & (ax117x) & (!g27) & (!g36) & (g38) & (g42)) + ((ax116x) & (ax117x) & (!g27) & (g36) & (!g38) & (g42)) + ((ax116x) & (ax117x) & (!g27) & (g36) & (g38) & (g42)) + ((ax116x) & (ax117x) & (g27) & (!g36) & (!g38) & (g42)) + ((ax116x) & (ax117x) & (g27) & (!g36) & (g38) & (!g42)) + ((ax116x) & (ax117x) & (g27) & (!g36) & (g38) & (g42)) + ((ax116x) & (ax117x) & (g27) & (g36) & (!g38) & (g42)) + ((ax116x) & (ax117x) & (g27) & (g36) & (g38) & (g42)));
	assign g44 = (((!ax116x) & (!g27) & (!g31) & (!g36) & (g38)) + ((!ax116x) & (!g27) & (g31) & (!g36) & (!g38)) + ((!ax116x) & (!g27) & (g31) & (!g36) & (g38)) + ((!ax116x) & (!g27) & (g31) & (g36) & (!g38)) + ((!ax116x) & (!g27) & (g31) & (g36) & (g38)) + ((!ax116x) & (g27) & (g31) & (!g36) & (!g38)) + ((!ax116x) & (g27) & (g31) & (g36) & (!g38)) + ((!ax116x) & (g27) & (g31) & (g36) & (g38)) + ((ax116x) & (!g27) & (!g31) & (!g36) & (!g38)) + ((ax116x) & (!g27) & (!g31) & (g36) & (!g38)) + ((ax116x) & (!g27) & (!g31) & (g36) & (g38)) + ((ax116x) & (g27) & (!g31) & (!g36) & (!g38)) + ((ax116x) & (g27) & (!g31) & (!g36) & (g38)) + ((ax116x) & (g27) & (!g31) & (g36) & (!g38)) + ((ax116x) & (g27) & (!g31) & (g36) & (g38)) + ((ax116x) & (g27) & (g31) & (!g36) & (g38)));
	assign g45 = (((!ax112x) & (!ax113x)));
	assign g46 = (((!g27) & (!ax114x) & (!ax115x) & (!g36) & (!g38) & (!g45)) + ((!g27) & (!ax114x) & (!ax115x) & (g36) & (!g38) & (!g45)) + ((!g27) & (!ax114x) & (!ax115x) & (g36) & (g38) & (!g45)) + ((!g27) & (!ax114x) & (ax115x) & (!g36) & (g38) & (!g45)) + ((!g27) & (ax114x) & (ax115x) & (!g36) & (g38) & (!g45)) + ((!g27) & (ax114x) & (ax115x) & (!g36) & (g38) & (g45)) + ((g27) & (!ax114x) & (!ax115x) & (!g36) & (!g38) & (!g45)) + ((g27) & (!ax114x) & (!ax115x) & (!g36) & (!g38) & (g45)) + ((g27) & (!ax114x) & (!ax115x) & (!g36) & (g38) & (!g45)) + ((g27) & (!ax114x) & (!ax115x) & (g36) & (!g38) & (!g45)) + ((g27) & (!ax114x) & (!ax115x) & (g36) & (!g38) & (g45)) + ((g27) & (!ax114x) & (!ax115x) & (g36) & (g38) & (!g45)) + ((g27) & (!ax114x) & (!ax115x) & (g36) & (g38) & (g45)) + ((g27) & (!ax114x) & (ax115x) & (!g36) & (!g38) & (!g45)) + ((g27) & (!ax114x) & (ax115x) & (!g36) & (g38) & (!g45)) + ((g27) & (!ax114x) & (ax115x) & (!g36) & (g38) & (g45)) + ((g27) & (!ax114x) & (ax115x) & (g36) & (!g38) & (!g45)) + ((g27) & (!ax114x) & (ax115x) & (g36) & (g38) & (!g45)) + ((g27) & (ax114x) & (!ax115x) & (!g36) & (g38) & (!g45)) + ((g27) & (ax114x) & (!ax115x) & (!g36) & (g38) & (g45)) + ((g27) & (ax114x) & (ax115x) & (!g36) & (!g38) & (!g45)) + ((g27) & (ax114x) & (ax115x) & (!g36) & (!g38) & (g45)) + ((g27) & (ax114x) & (ax115x) & (!g36) & (g38) & (!g45)) + ((g27) & (ax114x) & (ax115x) & (!g36) & (g38) & (g45)) + ((g27) & (ax114x) & (ax115x) & (g36) & (!g38) & (!g45)) + ((g27) & (ax114x) & (ax115x) & (g36) & (!g38) & (g45)) + ((g27) & (ax114x) & (ax115x) & (g36) & (g38) & (!g45)) + ((g27) & (ax114x) & (ax115x) & (g36) & (g38) & (g45)));
	assign g47 = (((!g8) & (!g18) & (g43) & (g44) & (g46)) + ((!g8) & (g18) & (g43) & (!g44) & (g46)) + ((!g8) & (g18) & (g43) & (g44) & (!g46)) + ((!g8) & (g18) & (g43) & (g44) & (g46)) + ((g8) & (!g18) & (!g43) & (g44) & (g46)) + ((g8) & (!g18) & (g43) & (!g44) & (!g46)) + ((g8) & (!g18) & (g43) & (!g44) & (g46)) + ((g8) & (!g18) & (g43) & (g44) & (!g46)) + ((g8) & (!g18) & (g43) & (g44) & (g46)) + ((g8) & (g18) & (!g43) & (!g44) & (g46)) + ((g8) & (g18) & (!g43) & (g44) & (!g46)) + ((g8) & (g18) & (!g43) & (g44) & (g46)) + ((g8) & (g18) & (g43) & (!g44) & (!g46)) + ((g8) & (g18) & (g43) & (!g44) & (g46)) + ((g8) & (g18) & (g43) & (g44) & (!g46)) + ((g8) & (g18) & (g43) & (g44) & (g46)));
	assign g48 = (((!g2) & (!g8) & (g30) & (g32)) + ((!g2) & (g8) & (!g30) & (g32)) + ((!g2) & (g8) & (g30) & (!g32)) + ((!g2) & (g8) & (g30) & (g32)) + ((g2) & (!g8) & (!g30) & (!g32)) + ((g2) & (!g8) & (!g30) & (g32)) + ((g2) & (!g8) & (g30) & (!g32)) + ((g2) & (g8) & (!g30) & (!g32)));
	assign g49 = (((!g29) & (!g36) & (!g38) & (g48)) + ((!g29) & (g36) & (!g38) & (g48)) + ((!g29) & (g36) & (g38) & (g48)) + ((g29) & (!g36) & (!g38) & (!g48)) + ((g29) & (!g36) & (g38) & (!g48)) + ((g29) & (!g36) & (g38) & (g48)) + ((g29) & (g36) & (!g38) & (!g48)) + ((g29) & (g36) & (g38) & (!g48)));
	assign g50 = (((!g4) & (!g2) & (!g41) & (!g47) & (g49)) + ((!g4) & (!g2) & (!g41) & (g47) & (g49)) + ((!g4) & (!g2) & (g41) & (!g47) & (g49)) + ((!g4) & (!g2) & (g41) & (g47) & (!g49)) + ((!g4) & (!g2) & (g41) & (g47) & (g49)) + ((!g4) & (g2) & (!g41) & (!g47) & (g49)) + ((!g4) & (g2) & (!g41) & (g47) & (!g49)) + ((!g4) & (g2) & (!g41) & (g47) & (g49)) + ((!g4) & (g2) & (g41) & (!g47) & (!g49)) + ((!g4) & (g2) & (g41) & (!g47) & (g49)) + ((!g4) & (g2) & (g41) & (g47) & (!g49)) + ((!g4) & (g2) & (g41) & (g47) & (g49)) + ((g4) & (!g2) & (g41) & (g47) & (g49)) + ((g4) & (g2) & (!g41) & (g47) & (g49)) + ((g4) & (g2) & (g41) & (!g47) & (g49)) + ((g4) & (g2) & (g41) & (g47) & (g49)));
	assign g51 = (((!g4) & (!g33) & (g34)) + ((!g4) & (g33) & (!g34)) + ((!g4) & (g33) & (g34)) + ((g4) & (g33) & (g34)));
	assign g52 = (((!g28) & (!g51) & (!g36) & (!g38)) + ((!g28) & (!g51) & (g36) & (!g38)) + ((!g28) & (!g51) & (g36) & (g38)) + ((g28) & (g51) & (!g36) & (!g38)) + ((g28) & (g51) & (!g36) & (g38)) + ((g28) & (g51) & (g36) & (!g38)) + ((g28) & (g51) & (g36) & (g38)));
	assign g53 = (((!g1) & (g28) & (!g51) & (!g36) & (!g37)) + ((g1) & (!g28) & (g51) & (!g36) & (g37)) + ((g1) & (!g28) & (g51) & (g36) & (g37)) + ((g1) & (g28) & (!g51) & (!g36) & (!g37)) + ((g1) & (g28) & (!g51) & (!g36) & (g37)) + ((g1) & (g28) & (!g51) & (g36) & (!g37)) + ((g1) & (g28) & (!g51) & (g36) & (g37)));
	assign g54 = (((!g1) & (!g40) & (!g50) & (!g52) & (!g53)) + ((g1) & (!g40) & (!g50) & (!g52) & (!g53)) + ((g1) & (!g40) & (!g50) & (g52) & (!g53)) + ((g1) & (!g40) & (g50) & (!g52) & (!g53)) + ((g1) & (!g40) & (g50) & (g52) & (!g53)) + ((g1) & (g40) & (!g50) & (!g52) & (!g53)) + ((g1) & (g40) & (!g50) & (g52) & (!g53)));
	assign g55 = (((g1) & (!g40) & (g50) & (g53)) + ((g1) & (g40) & (!g50) & (!g53)) + ((g1) & (g40) & (!g50) & (g53)));
	assign g56 = (((!g4) & (!g2) & (!g41) & (!g47) & (!g49) & (!g54)) + ((!g4) & (!g2) & (!g41) & (!g47) & (g49) & (g54)) + ((!g4) & (!g2) & (!g41) & (g47) & (!g49) & (!g54)) + ((!g4) & (!g2) & (!g41) & (g47) & (g49) & (g54)) + ((!g4) & (!g2) & (g41) & (!g47) & (!g49) & (!g54)) + ((!g4) & (!g2) & (g41) & (!g47) & (g49) & (g54)) + ((!g4) & (!g2) & (g41) & (g47) & (g49) & (!g54)) + ((!g4) & (!g2) & (g41) & (g47) & (g49) & (g54)) + ((!g4) & (g2) & (!g41) & (!g47) & (!g49) & (!g54)) + ((!g4) & (g2) & (!g41) & (!g47) & (g49) & (g54)) + ((!g4) & (g2) & (!g41) & (g47) & (g49) & (!g54)) + ((!g4) & (g2) & (!g41) & (g47) & (g49) & (g54)) + ((!g4) & (g2) & (g41) & (!g47) & (g49) & (!g54)) + ((!g4) & (g2) & (g41) & (!g47) & (g49) & (g54)) + ((!g4) & (g2) & (g41) & (g47) & (g49) & (!g54)) + ((!g4) & (g2) & (g41) & (g47) & (g49) & (g54)) + ((g4) & (!g2) & (!g41) & (!g47) & (g49) & (!g54)) + ((g4) & (!g2) & (!g41) & (!g47) & (g49) & (g54)) + ((g4) & (!g2) & (!g41) & (g47) & (g49) & (!g54)) + ((g4) & (!g2) & (!g41) & (g47) & (g49) & (g54)) + ((g4) & (!g2) & (g41) & (!g47) & (g49) & (!g54)) + ((g4) & (!g2) & (g41) & (!g47) & (g49) & (g54)) + ((g4) & (!g2) & (g41) & (g47) & (!g49) & (!g54)) + ((g4) & (!g2) & (g41) & (g47) & (g49) & (g54)) + ((g4) & (g2) & (!g41) & (!g47) & (g49) & (!g54)) + ((g4) & (g2) & (!g41) & (!g47) & (g49) & (g54)) + ((g4) & (g2) & (!g41) & (g47) & (!g49) & (!g54)) + ((g4) & (g2) & (!g41) & (g47) & (g49) & (g54)) + ((g4) & (g2) & (g41) & (!g47) & (!g49) & (!g54)) + ((g4) & (g2) & (g41) & (!g47) & (g49) & (g54)) + ((g4) & (g2) & (g41) & (g47) & (!g49) & (!g54)) + ((g4) & (g2) & (g41) & (g47) & (g49) & (g54)));
	assign g57 = (((!g8) & (!g18) & (!g43) & (g44) & (g46) & (!g54)) + ((!g8) & (!g18) & (g43) & (!g44) & (!g46) & (!g54)) + ((!g8) & (!g18) & (g43) & (!g44) & (!g46) & (g54)) + ((!g8) & (!g18) & (g43) & (!g44) & (g46) & (!g54)) + ((!g8) & (!g18) & (g43) & (!g44) & (g46) & (g54)) + ((!g8) & (!g18) & (g43) & (g44) & (!g46) & (!g54)) + ((!g8) & (!g18) & (g43) & (g44) & (!g46) & (g54)) + ((!g8) & (!g18) & (g43) & (g44) & (g46) & (g54)) + ((!g8) & (g18) & (!g43) & (!g44) & (g46) & (!g54)) + ((!g8) & (g18) & (!g43) & (g44) & (!g46) & (!g54)) + ((!g8) & (g18) & (!g43) & (g44) & (g46) & (!g54)) + ((!g8) & (g18) & (g43) & (!g44) & (!g46) & (!g54)) + ((!g8) & (g18) & (g43) & (!g44) & (!g46) & (g54)) + ((!g8) & (g18) & (g43) & (!g44) & (g46) & (g54)) + ((!g8) & (g18) & (g43) & (g44) & (!g46) & (g54)) + ((!g8) & (g18) & (g43) & (g44) & (g46) & (g54)) + ((g8) & (!g18) & (!g43) & (!g44) & (!g46) & (!g54)) + ((g8) & (!g18) & (!g43) & (!g44) & (g46) & (!g54)) + ((g8) & (!g18) & (!g43) & (g44) & (!g46) & (!g54)) + ((g8) & (!g18) & (g43) & (!g44) & (!g46) & (g54)) + ((g8) & (!g18) & (g43) & (!g44) & (g46) & (g54)) + ((g8) & (!g18) & (g43) & (g44) & (!g46) & (g54)) + ((g8) & (!g18) & (g43) & (g44) & (g46) & (!g54)) + ((g8) & (!g18) & (g43) & (g44) & (g46) & (g54)) + ((g8) & (g18) & (!g43) & (!g44) & (!g46) & (!g54)) + ((g8) & (g18) & (g43) & (!g44) & (!g46) & (g54)) + ((g8) & (g18) & (g43) & (!g44) & (g46) & (!g54)) + ((g8) & (g18) & (g43) & (!g44) & (g46) & (g54)) + ((g8) & (g18) & (g43) & (g44) & (!g46) & (!g54)) + ((g8) & (g18) & (g43) & (g44) & (!g46) & (g54)) + ((g8) & (g18) & (g43) & (g44) & (g46) & (!g54)) + ((g8) & (g18) & (g43) & (g44) & (g46) & (g54)));
	assign g58 = (((!g18) & (!g44) & (g46) & (!g54)) + ((!g18) & (g44) & (!g46) & (!g54)) + ((!g18) & (g44) & (!g46) & (g54)) + ((!g18) & (g44) & (g46) & (g54)) + ((g18) & (!g44) & (!g46) & (!g54)) + ((g18) & (g44) & (!g46) & (g54)) + ((g18) & (g44) & (g46) & (!g54)) + ((g18) & (g44) & (g46) & (g54)));
	assign g59 = (((!g27) & (!ax114x) & (!ax115x) & (!g39) & (!g45) & (g54)) + ((!g27) & (!ax114x) & (!ax115x) & (!g39) & (g45) & (!g54)) + ((!g27) & (!ax114x) & (!ax115x) & (!g39) & (g45) & (g54)) + ((!g27) & (!ax114x) & (!ax115x) & (g39) & (!g45) & (!g54)) + ((!g27) & (!ax114x) & (ax115x) & (!g39) & (!g45) & (!g54)) + ((!g27) & (!ax114x) & (ax115x) & (g39) & (!g45) & (g54)) + ((!g27) & (!ax114x) & (ax115x) & (g39) & (g45) & (!g54)) + ((!g27) & (!ax114x) & (ax115x) & (g39) & (g45) & (g54)) + ((!g27) & (ax114x) & (!ax115x) & (g39) & (!g45) & (!g54)) + ((!g27) & (ax114x) & (!ax115x) & (g39) & (g45) & (!g54)) + ((!g27) & (ax114x) & (ax115x) & (!g39) & (!g45) & (!g54)) + ((!g27) & (ax114x) & (ax115x) & (!g39) & (!g45) & (g54)) + ((!g27) & (ax114x) & (ax115x) & (!g39) & (g45) & (!g54)) + ((!g27) & (ax114x) & (ax115x) & (!g39) & (g45) & (g54)) + ((!g27) & (ax114x) & (ax115x) & (g39) & (!g45) & (g54)) + ((!g27) & (ax114x) & (ax115x) & (g39) & (g45) & (g54)) + ((g27) & (!ax114x) & (!ax115x) & (!g39) & (!g45) & (!g54)) + ((g27) & (!ax114x) & (!ax115x) & (!g39) & (!g45) & (g54)) + ((g27) & (!ax114x) & (!ax115x) & (!g39) & (g45) & (g54)) + ((g27) & (!ax114x) & (!ax115x) & (g39) & (g45) & (!g54)) + ((g27) & (!ax114x) & (ax115x) & (!g39) & (g45) & (!g54)) + ((g27) & (!ax114x) & (ax115x) & (g39) & (!g45) & (!g54)) + ((g27) & (!ax114x) & (ax115x) & (g39) & (!g45) & (g54)) + ((g27) & (!ax114x) & (ax115x) & (g39) & (g45) & (g54)) + ((g27) & (ax114x) & (!ax115x) & (!g39) & (!g45) & (!g54)) + ((g27) & (ax114x) & (!ax115x) & (!g39) & (g45) & (!g54)) + ((g27) & (ax114x) & (ax115x) & (!g39) & (!g45) & (g54)) + ((g27) & (ax114x) & (ax115x) & (!g39) & (g45) & (g54)) + ((g27) & (ax114x) & (ax115x) & (g39) & (!g45) & (!g54)) + ((g27) & (ax114x) & (ax115x) & (g39) & (!g45) & (g54)) + ((g27) & (ax114x) & (ax115x) & (g39) & (g45) & (!g54)) + ((g27) & (ax114x) & (ax115x) & (g39) & (g45) & (g54)));
	assign g60 = (((!ax114x) & (!g39) & (!g45) & (g54)) + ((!ax114x) & (!g39) & (g45) & (!g54)) + ((!ax114x) & (!g39) & (g45) & (g54)) + ((!ax114x) & (g39) & (g45) & (!g54)) + ((ax114x) & (!g39) & (!g45) & (!g54)) + ((ax114x) & (g39) & (!g45) & (!g54)) + ((ax114x) & (g39) & (!g45) & (g54)) + ((ax114x) & (g39) & (g45) & (g54)));
	assign g61 = (((!ax110x) & (!ax111x)));
	assign g62 = (((!ax112x) & (!ax113x) & (!g39) & (!g54) & (!g61)) + ((!ax112x) & (!ax113x) & (g39) & (!g54) & (!g61)) + ((!ax112x) & (!ax113x) & (g39) & (!g54) & (g61)) + ((!ax112x) & (!ax113x) & (g39) & (g54) & (!g61)) + ((!ax112x) & (ax113x) & (!g39) & (g54) & (!g61)) + ((!ax112x) & (ax113x) & (g39) & (!g54) & (!g61)) + ((!ax112x) & (ax113x) & (g39) & (g54) & (!g61)) + ((!ax112x) & (ax113x) & (g39) & (g54) & (g61)) + ((ax112x) & (!ax113x) & (g39) & (g54) & (!g61)) + ((ax112x) & (!ax113x) & (g39) & (g54) & (g61)) + ((ax112x) & (ax113x) & (!g39) & (g54) & (!g61)) + ((ax112x) & (ax113x) & (!g39) & (g54) & (g61)) + ((ax112x) & (ax113x) & (g39) & (!g54) & (!g61)) + ((ax112x) & (ax113x) & (g39) & (!g54) & (g61)) + ((ax112x) & (ax113x) & (g39) & (g54) & (!g61)) + ((ax112x) & (ax113x) & (g39) & (g54) & (g61)));
	assign g63 = (((!g18) & (!g27) & (g59) & (g60) & (g62)) + ((!g18) & (g27) & (g59) & (!g60) & (g62)) + ((!g18) & (g27) & (g59) & (g60) & (!g62)) + ((!g18) & (g27) & (g59) & (g60) & (g62)) + ((g18) & (!g27) & (!g59) & (g60) & (g62)) + ((g18) & (!g27) & (g59) & (!g60) & (!g62)) + ((g18) & (!g27) & (g59) & (!g60) & (g62)) + ((g18) & (!g27) & (g59) & (g60) & (!g62)) + ((g18) & (!g27) & (g59) & (g60) & (g62)) + ((g18) & (g27) & (!g59) & (!g60) & (g62)) + ((g18) & (g27) & (!g59) & (g60) & (!g62)) + ((g18) & (g27) & (!g59) & (g60) & (g62)) + ((g18) & (g27) & (g59) & (!g60) & (!g62)) + ((g18) & (g27) & (g59) & (!g60) & (g62)) + ((g18) & (g27) & (g59) & (g60) & (!g62)) + ((g18) & (g27) & (g59) & (g60) & (g62)));
	assign g64 = (((!g2) & (!g8) & (g57) & (g58) & (g63)) + ((!g2) & (g8) & (g57) & (!g58) & (g63)) + ((!g2) & (g8) & (g57) & (g58) & (!g63)) + ((!g2) & (g8) & (g57) & (g58) & (g63)) + ((g2) & (!g8) & (!g57) & (g58) & (g63)) + ((g2) & (!g8) & (g57) & (!g58) & (!g63)) + ((g2) & (!g8) & (g57) & (!g58) & (g63)) + ((g2) & (!g8) & (g57) & (g58) & (!g63)) + ((g2) & (!g8) & (g57) & (g58) & (g63)) + ((g2) & (g8) & (!g57) & (!g58) & (g63)) + ((g2) & (g8) & (!g57) & (g58) & (!g63)) + ((g2) & (g8) & (!g57) & (g58) & (g63)) + ((g2) & (g8) & (g57) & (!g58) & (!g63)) + ((g2) & (g8) & (g57) & (!g58) & (g63)) + ((g2) & (g8) & (g57) & (g58) & (!g63)) + ((g2) & (g8) & (g57) & (g58) & (g63)));
	assign g65 = (((!g2) & (!g41) & (g47) & (!g54)) + ((!g2) & (g41) & (!g47) & (!g54)) + ((!g2) & (g41) & (!g47) & (g54)) + ((!g2) & (g41) & (g47) & (g54)) + ((g2) & (!g41) & (!g47) & (!g54)) + ((g2) & (g41) & (!g47) & (g54)) + ((g2) & (g41) & (g47) & (!g54)) + ((g2) & (g41) & (g47) & (g54)));
	assign g66 = (((!g1) & (!g40) & (!g50) & (!g52) & (g53)) + ((!g1) & (!g40) & (!g50) & (g52) & (!g53)) + ((!g1) & (!g40) & (!g50) & (g52) & (g53)) + ((!g1) & (g40) & (g50) & (!g52) & (!g53)) + ((!g1) & (g40) & (g50) & (!g52) & (g53)) + ((!g1) & (g40) & (g50) & (g52) & (!g53)) + ((!g1) & (g40) & (g50) & (g52) & (g53)) + ((g1) & (!g40) & (!g50) & (!g52) & (g53)) + ((g1) & (!g40) & (!g50) & (g52) & (g53)) + ((g1) & (g40) & (g50) & (!g52) & (!g53)) + ((g1) & (g40) & (g50) & (!g52) & (g53)) + ((g1) & (g40) & (g50) & (g52) & (!g53)) + ((g1) & (g40) & (g50) & (g52) & (g53)));
	assign g67 = (((!g4) & (!g1) & (!g56) & (!g64) & (!g65) & (!g66)) + ((!g4) & (g1) & (!g56) & (!g64) & (!g65) & (!g66)) + ((!g4) & (g1) & (!g56) & (!g64) & (!g65) & (g66)) + ((!g4) & (g1) & (!g56) & (!g64) & (g65) & (!g66)) + ((!g4) & (g1) & (!g56) & (!g64) & (g65) & (g66)) + ((!g4) & (g1) & (!g56) & (g64) & (!g65) & (!g66)) + ((!g4) & (g1) & (!g56) & (g64) & (!g65) & (g66)) + ((!g4) & (g1) & (!g56) & (g64) & (g65) & (!g66)) + ((!g4) & (g1) & (!g56) & (g64) & (g65) & (g66)) + ((!g4) & (g1) & (g56) & (!g64) & (!g65) & (!g66)) + ((!g4) & (g1) & (g56) & (!g64) & (!g65) & (g66)) + ((g4) & (!g1) & (!g56) & (!g64) & (!g65) & (!g66)) + ((g4) & (!g1) & (!g56) & (!g64) & (g65) & (!g66)) + ((g4) & (!g1) & (!g56) & (g64) & (!g65) & (!g66)) + ((g4) & (g1) & (!g56) & (!g64) & (!g65) & (!g66)) + ((g4) & (g1) & (!g56) & (!g64) & (!g65) & (g66)) + ((g4) & (g1) & (!g56) & (!g64) & (g65) & (!g66)) + ((g4) & (g1) & (!g56) & (!g64) & (g65) & (g66)) + ((g4) & (g1) & (!g56) & (g64) & (!g65) & (!g66)) + ((g4) & (g1) & (!g56) & (g64) & (!g65) & (g66)) + ((g4) & (g1) & (!g56) & (g64) & (g65) & (!g66)) + ((g4) & (g1) & (!g56) & (g64) & (g65) & (g66)) + ((g4) & (g1) & (g56) & (!g64) & (!g65) & (!g66)) + ((g4) & (g1) & (g56) & (!g64) & (!g65) & (g66)) + ((g4) & (g1) & (g56) & (!g64) & (g65) & (!g66)) + ((g4) & (g1) & (g56) & (!g64) & (g65) & (g66)) + ((g4) & (g1) & (g56) & (g64) & (!g65) & (!g66)) + ((g4) & (g1) & (g56) & (g64) & (!g65) & (g66)));
	assign g68 = (((!g55) & (g67)));
	assign g69 = (((!g4) & (!g64) & (!g65) & (!g55) & (!g67)) + ((!g4) & (!g64) & (!g65) & (g55) & (!g67)) + ((!g4) & (!g64) & (!g65) & (g55) & (g67)) + ((!g4) & (!g64) & (g65) & (!g55) & (g67)) + ((!g4) & (g64) & (g65) & (!g55) & (!g67)) + ((!g4) & (g64) & (g65) & (!g55) & (g67)) + ((!g4) & (g64) & (g65) & (g55) & (!g67)) + ((!g4) & (g64) & (g65) & (g55) & (g67)) + ((g4) & (!g64) & (g65) & (!g55) & (!g67)) + ((g4) & (!g64) & (g65) & (!g55) & (g67)) + ((g4) & (!g64) & (g65) & (g55) & (!g67)) + ((g4) & (!g64) & (g65) & (g55) & (g67)) + ((g4) & (g64) & (!g65) & (!g55) & (!g67)) + ((g4) & (g64) & (!g65) & (g55) & (!g67)) + ((g4) & (g64) & (!g65) & (g55) & (g67)) + ((g4) & (g64) & (g65) & (!g55) & (g67)));
	assign g70 = (((!g8) & (!g58) & (g63) & (!g55) & (!g67)) + ((!g8) & (!g58) & (g63) & (g55) & (!g67)) + ((!g8) & (!g58) & (g63) & (g55) & (g67)) + ((!g8) & (g58) & (!g63) & (!g55) & (!g67)) + ((!g8) & (g58) & (!g63) & (!g55) & (g67)) + ((!g8) & (g58) & (!g63) & (g55) & (!g67)) + ((!g8) & (g58) & (!g63) & (g55) & (g67)) + ((!g8) & (g58) & (g63) & (!g55) & (g67)) + ((g8) & (!g58) & (!g63) & (!g55) & (!g67)) + ((g8) & (!g58) & (!g63) & (g55) & (!g67)) + ((g8) & (!g58) & (!g63) & (g55) & (g67)) + ((g8) & (g58) & (!g63) & (!g55) & (g67)) + ((g8) & (g58) & (g63) & (!g55) & (!g67)) + ((g8) & (g58) & (g63) & (!g55) & (g67)) + ((g8) & (g58) & (g63) & (g55) & (!g67)) + ((g8) & (g58) & (g63) & (g55) & (g67)));
	assign g71 = (((!g18) & (!g27) & (g60) & (g62)) + ((!g18) & (g27) & (!g60) & (g62)) + ((!g18) & (g27) & (g60) & (!g62)) + ((!g18) & (g27) & (g60) & (g62)) + ((g18) & (!g27) & (!g60) & (!g62)) + ((g18) & (!g27) & (!g60) & (g62)) + ((g18) & (!g27) & (g60) & (!g62)) + ((g18) & (g27) & (!g60) & (!g62)));
	assign g72 = (((!g59) & (!g55) & (!g67) & (g71)) + ((!g59) & (g55) & (!g67) & (g71)) + ((!g59) & (g55) & (g67) & (g71)) + ((g59) & (!g55) & (!g67) & (!g71)) + ((g59) & (!g55) & (g67) & (!g71)) + ((g59) & (!g55) & (g67) & (g71)) + ((g59) & (g55) & (!g67) & (!g71)) + ((g59) & (g55) & (g67) & (!g71)));
	assign g73 = (((!g27) & (!g60) & (g62) & (!g55) & (!g67)) + ((!g27) & (!g60) & (g62) & (g55) & (!g67)) + ((!g27) & (!g60) & (g62) & (g55) & (g67)) + ((!g27) & (g60) & (!g62) & (!g55) & (!g67)) + ((!g27) & (g60) & (!g62) & (!g55) & (g67)) + ((!g27) & (g60) & (!g62) & (g55) & (!g67)) + ((!g27) & (g60) & (!g62) & (g55) & (g67)) + ((!g27) & (g60) & (g62) & (!g55) & (g67)) + ((g27) & (!g60) & (!g62) & (!g55) & (!g67)) + ((g27) & (!g60) & (!g62) & (g55) & (!g67)) + ((g27) & (!g60) & (!g62) & (g55) & (g67)) + ((g27) & (g60) & (!g62) & (!g55) & (g67)) + ((g27) & (g60) & (g62) & (!g55) & (!g67)) + ((g27) & (g60) & (g62) & (!g55) & (g67)) + ((g27) & (g60) & (g62) & (g55) & (!g67)) + ((g27) & (g60) & (g62) & (g55) & (g67)));
	assign g74 = (((!ax112x) & (!g39) & (!g54) & (!g61)) + ((!ax112x) & (!g39) & (g54) & (!g61)) + ((!ax112x) & (g39) & (!g54) & (g61)) + ((!ax112x) & (g39) & (g54) & (g61)) + ((ax112x) & (!g39) & (g54) & (!g61)) + ((ax112x) & (!g39) & (g54) & (g61)) + ((ax112x) & (g39) & (!g54) & (!g61)) + ((ax112x) & (g39) & (!g54) & (g61)));
	assign g75 = (((!ax112x) & (!ax113x) & (!g54) & (!g55) & (!g67) & (!g74)) + ((!ax112x) & (!ax113x) & (!g54) & (!g55) & (g67) & (!g74)) + ((!ax112x) & (!ax113x) & (!g54) & (!g55) & (g67) & (g74)) + ((!ax112x) & (!ax113x) & (!g54) & (g55) & (!g67) & (!g74)) + ((!ax112x) & (!ax113x) & (!g54) & (g55) & (g67) & (!g74)) + ((!ax112x) & (!ax113x) & (g54) & (!g55) & (!g67) & (g74)) + ((!ax112x) & (!ax113x) & (g54) & (g55) & (!g67) & (g74)) + ((!ax112x) & (!ax113x) & (g54) & (g55) & (g67) & (g74)) + ((!ax112x) & (ax113x) & (!g54) & (!g55) & (!g67) & (g74)) + ((!ax112x) & (ax113x) & (!g54) & (g55) & (!g67) & (g74)) + ((!ax112x) & (ax113x) & (!g54) & (g55) & (g67) & (g74)) + ((!ax112x) & (ax113x) & (g54) & (!g55) & (!g67) & (!g74)) + ((!ax112x) & (ax113x) & (g54) & (!g55) & (g67) & (!g74)) + ((!ax112x) & (ax113x) & (g54) & (!g55) & (g67) & (g74)) + ((!ax112x) & (ax113x) & (g54) & (g55) & (!g67) & (!g74)) + ((!ax112x) & (ax113x) & (g54) & (g55) & (g67) & (!g74)) + ((ax112x) & (!ax113x) & (!g54) & (!g55) & (!g67) & (g74)) + ((ax112x) & (!ax113x) & (!g54) & (g55) & (!g67) & (g74)) + ((ax112x) & (!ax113x) & (!g54) & (g55) & (g67) & (g74)) + ((ax112x) & (!ax113x) & (g54) & (!g55) & (!g67) & (g74)) + ((ax112x) & (!ax113x) & (g54) & (g55) & (!g67) & (g74)) + ((ax112x) & (!ax113x) & (g54) & (g55) & (g67) & (g74)) + ((ax112x) & (ax113x) & (!g54) & (!g55) & (!g67) & (!g74)) + ((ax112x) & (ax113x) & (!g54) & (!g55) & (g67) & (!g74)) + ((ax112x) & (ax113x) & (!g54) & (!g55) & (g67) & (g74)) + ((ax112x) & (ax113x) & (!g54) & (g55) & (!g67) & (!g74)) + ((ax112x) & (ax113x) & (!g54) & (g55) & (g67) & (!g74)) + ((ax112x) & (ax113x) & (g54) & (!g55) & (!g67) & (!g74)) + ((ax112x) & (ax113x) & (g54) & (!g55) & (g67) & (!g74)) + ((ax112x) & (ax113x) & (g54) & (!g55) & (g67) & (g74)) + ((ax112x) & (ax113x) & (g54) & (g55) & (!g67) & (!g74)) + ((ax112x) & (ax113x) & (g54) & (g55) & (g67) & (!g74)));
	assign g76 = (((!ax112x) & (!g54) & (!g61) & (!g55) & (g67)) + ((!ax112x) & (!g54) & (g61) & (!g55) & (!g67)) + ((!ax112x) & (!g54) & (g61) & (!g55) & (g67)) + ((!ax112x) & (!g54) & (g61) & (g55) & (!g67)) + ((!ax112x) & (!g54) & (g61) & (g55) & (g67)) + ((!ax112x) & (g54) & (g61) & (!g55) & (!g67)) + ((!ax112x) & (g54) & (g61) & (g55) & (!g67)) + ((!ax112x) & (g54) & (g61) & (g55) & (g67)) + ((ax112x) & (!g54) & (!g61) & (!g55) & (!g67)) + ((ax112x) & (!g54) & (!g61) & (g55) & (!g67)) + ((ax112x) & (!g54) & (!g61) & (g55) & (g67)) + ((ax112x) & (g54) & (!g61) & (!g55) & (!g67)) + ((ax112x) & (g54) & (!g61) & (!g55) & (g67)) + ((ax112x) & (g54) & (!g61) & (g55) & (!g67)) + ((ax112x) & (g54) & (!g61) & (g55) & (g67)) + ((ax112x) & (g54) & (g61) & (!g55) & (g67)));
	assign g77 = (((!ax108x) & (!ax109x)));
	assign g78 = (((!g54) & (!ax110x) & (!ax111x) & (!g55) & (!g67) & (!g77)) + ((!g54) & (!ax110x) & (!ax111x) & (g55) & (!g67) & (!g77)) + ((!g54) & (!ax110x) & (!ax111x) & (g55) & (g67) & (!g77)) + ((!g54) & (!ax110x) & (ax111x) & (!g55) & (g67) & (!g77)) + ((!g54) & (ax110x) & (ax111x) & (!g55) & (g67) & (!g77)) + ((!g54) & (ax110x) & (ax111x) & (!g55) & (g67) & (g77)) + ((g54) & (!ax110x) & (!ax111x) & (!g55) & (!g67) & (!g77)) + ((g54) & (!ax110x) & (!ax111x) & (!g55) & (!g67) & (g77)) + ((g54) & (!ax110x) & (!ax111x) & (!g55) & (g67) & (!g77)) + ((g54) & (!ax110x) & (!ax111x) & (g55) & (!g67) & (!g77)) + ((g54) & (!ax110x) & (!ax111x) & (g55) & (!g67) & (g77)) + ((g54) & (!ax110x) & (!ax111x) & (g55) & (g67) & (!g77)) + ((g54) & (!ax110x) & (!ax111x) & (g55) & (g67) & (g77)) + ((g54) & (!ax110x) & (ax111x) & (!g55) & (!g67) & (!g77)) + ((g54) & (!ax110x) & (ax111x) & (!g55) & (g67) & (!g77)) + ((g54) & (!ax110x) & (ax111x) & (!g55) & (g67) & (g77)) + ((g54) & (!ax110x) & (ax111x) & (g55) & (!g67) & (!g77)) + ((g54) & (!ax110x) & (ax111x) & (g55) & (g67) & (!g77)) + ((g54) & (ax110x) & (!ax111x) & (!g55) & (g67) & (!g77)) + ((g54) & (ax110x) & (!ax111x) & (!g55) & (g67) & (g77)) + ((g54) & (ax110x) & (ax111x) & (!g55) & (!g67) & (!g77)) + ((g54) & (ax110x) & (ax111x) & (!g55) & (!g67) & (g77)) + ((g54) & (ax110x) & (ax111x) & (!g55) & (g67) & (!g77)) + ((g54) & (ax110x) & (ax111x) & (!g55) & (g67) & (g77)) + ((g54) & (ax110x) & (ax111x) & (g55) & (!g67) & (!g77)) + ((g54) & (ax110x) & (ax111x) & (g55) & (!g67) & (g77)) + ((g54) & (ax110x) & (ax111x) & (g55) & (g67) & (!g77)) + ((g54) & (ax110x) & (ax111x) & (g55) & (g67) & (g77)));
	assign g79 = (((!g27) & (!g39) & (g75) & (g76) & (g78)) + ((!g27) & (g39) & (g75) & (!g76) & (g78)) + ((!g27) & (g39) & (g75) & (g76) & (!g78)) + ((!g27) & (g39) & (g75) & (g76) & (g78)) + ((g27) & (!g39) & (!g75) & (g76) & (g78)) + ((g27) & (!g39) & (g75) & (!g76) & (!g78)) + ((g27) & (!g39) & (g75) & (!g76) & (g78)) + ((g27) & (!g39) & (g75) & (g76) & (!g78)) + ((g27) & (!g39) & (g75) & (g76) & (g78)) + ((g27) & (g39) & (!g75) & (!g76) & (g78)) + ((g27) & (g39) & (!g75) & (g76) & (!g78)) + ((g27) & (g39) & (!g75) & (g76) & (g78)) + ((g27) & (g39) & (g75) & (!g76) & (!g78)) + ((g27) & (g39) & (g75) & (!g76) & (g78)) + ((g27) & (g39) & (g75) & (g76) & (!g78)) + ((g27) & (g39) & (g75) & (g76) & (g78)));
	assign g80 = (((!g8) & (!g18) & (g72) & (g73) & (g79)) + ((!g8) & (g18) & (g72) & (!g73) & (g79)) + ((!g8) & (g18) & (g72) & (g73) & (!g79)) + ((!g8) & (g18) & (g72) & (g73) & (g79)) + ((g8) & (!g18) & (!g72) & (g73) & (g79)) + ((g8) & (!g18) & (g72) & (!g73) & (!g79)) + ((g8) & (!g18) & (g72) & (!g73) & (g79)) + ((g8) & (!g18) & (g72) & (g73) & (!g79)) + ((g8) & (!g18) & (g72) & (g73) & (g79)) + ((g8) & (g18) & (!g72) & (!g73) & (g79)) + ((g8) & (g18) & (!g72) & (g73) & (!g79)) + ((g8) & (g18) & (!g72) & (g73) & (g79)) + ((g8) & (g18) & (g72) & (!g73) & (!g79)) + ((g8) & (g18) & (g72) & (!g73) & (g79)) + ((g8) & (g18) & (g72) & (g73) & (!g79)) + ((g8) & (g18) & (g72) & (g73) & (g79)));
	assign g81 = (((!g2) & (!g8) & (g58) & (g63)) + ((!g2) & (g8) & (!g58) & (g63)) + ((!g2) & (g8) & (g58) & (!g63)) + ((!g2) & (g8) & (g58) & (g63)) + ((g2) & (!g8) & (!g58) & (!g63)) + ((g2) & (!g8) & (!g58) & (g63)) + ((g2) & (!g8) & (g58) & (!g63)) + ((g2) & (g8) & (!g58) & (!g63)));
	assign g82 = (((!g57) & (!g55) & (!g67) & (g81)) + ((!g57) & (g55) & (!g67) & (g81)) + ((!g57) & (g55) & (g67) & (g81)) + ((g57) & (!g55) & (!g67) & (!g81)) + ((g57) & (!g55) & (g67) & (!g81)) + ((g57) & (!g55) & (g67) & (g81)) + ((g57) & (g55) & (!g67) & (!g81)) + ((g57) & (g55) & (g67) & (!g81)));
	assign g83 = (((!g4) & (!g2) & (!g70) & (!g80) & (g82)) + ((!g4) & (!g2) & (!g70) & (g80) & (g82)) + ((!g4) & (!g2) & (g70) & (!g80) & (g82)) + ((!g4) & (!g2) & (g70) & (g80) & (!g82)) + ((!g4) & (!g2) & (g70) & (g80) & (g82)) + ((!g4) & (g2) & (!g70) & (!g80) & (g82)) + ((!g4) & (g2) & (!g70) & (g80) & (!g82)) + ((!g4) & (g2) & (!g70) & (g80) & (g82)) + ((!g4) & (g2) & (g70) & (!g80) & (!g82)) + ((!g4) & (g2) & (g70) & (!g80) & (g82)) + ((!g4) & (g2) & (g70) & (g80) & (!g82)) + ((!g4) & (g2) & (g70) & (g80) & (g82)) + ((g4) & (!g2) & (g70) & (g80) & (g82)) + ((g4) & (g2) & (!g70) & (g80) & (g82)) + ((g4) & (g2) & (g70) & (!g80) & (g82)) + ((g4) & (g2) & (g70) & (g80) & (g82)));
	assign g84 = (((!g4) & (!g64) & (g65)) + ((!g4) & (g64) & (!g65)) + ((!g4) & (g64) & (g65)) + ((g4) & (g64) & (g65)));
	assign g85 = (((!g56) & (!g84) & (!g55) & (!g67)) + ((!g56) & (!g84) & (g55) & (!g67)) + ((!g56) & (!g84) & (g55) & (g67)) + ((g56) & (g84) & (!g55) & (!g67)) + ((g56) & (g84) & (!g55) & (g67)) + ((g56) & (g84) & (g55) & (!g67)) + ((g56) & (g84) & (g55) & (g67)));
	assign g86 = (((!g1) & (g56) & (!g84) & (!g55) & (g67)) + ((!g1) & (g56) & (g84) & (!g55) & (g67)) + ((g1) & (!g56) & (g84) & (g55) & (!g67)) + ((g1) & (!g56) & (g84) & (g55) & (g67)) + ((g1) & (g56) & (!g84) & (!g55) & (!g67)) + ((g1) & (g56) & (!g84) & (!g55) & (g67)) + ((g1) & (g56) & (!g84) & (g55) & (!g67)) + ((g1) & (g56) & (!g84) & (g55) & (g67)) + ((g1) & (g56) & (g84) & (!g55) & (g67)));
	assign g87 = (((!g1) & (!g69) & (!g83) & (!g85) & (!g86)) + ((g1) & (!g69) & (!g83) & (!g85) & (!g86)) + ((g1) & (!g69) & (!g83) & (g85) & (!g86)) + ((g1) & (!g69) & (g83) & (!g85) & (!g86)) + ((g1) & (!g69) & (g83) & (g85) & (!g86)) + ((g1) & (g69) & (!g83) & (!g85) & (!g86)) + ((g1) & (g69) & (!g83) & (g85) & (!g86)));
	assign g88 = (((g1) & (!g69) & (g83) & (g86)) + ((g1) & (g69) & (!g83) & (!g86)) + ((g1) & (g69) & (!g83) & (g86)));
	assign g89 = (((!g4) & (!g2) & (!g70) & (!g80) & (!g82) & (!g87)) + ((!g4) & (!g2) & (!g70) & (!g80) & (g82) & (g87)) + ((!g4) & (!g2) & (!g70) & (g80) & (!g82) & (!g87)) + ((!g4) & (!g2) & (!g70) & (g80) & (g82) & (g87)) + ((!g4) & (!g2) & (g70) & (!g80) & (!g82) & (!g87)) + ((!g4) & (!g2) & (g70) & (!g80) & (g82) & (g87)) + ((!g4) & (!g2) & (g70) & (g80) & (g82) & (!g87)) + ((!g4) & (!g2) & (g70) & (g80) & (g82) & (g87)) + ((!g4) & (g2) & (!g70) & (!g80) & (!g82) & (!g87)) + ((!g4) & (g2) & (!g70) & (!g80) & (g82) & (g87)) + ((!g4) & (g2) & (!g70) & (g80) & (g82) & (!g87)) + ((!g4) & (g2) & (!g70) & (g80) & (g82) & (g87)) + ((!g4) & (g2) & (g70) & (!g80) & (g82) & (!g87)) + ((!g4) & (g2) & (g70) & (!g80) & (g82) & (g87)) + ((!g4) & (g2) & (g70) & (g80) & (g82) & (!g87)) + ((!g4) & (g2) & (g70) & (g80) & (g82) & (g87)) + ((g4) & (!g2) & (!g70) & (!g80) & (g82) & (!g87)) + ((g4) & (!g2) & (!g70) & (!g80) & (g82) & (g87)) + ((g4) & (!g2) & (!g70) & (g80) & (g82) & (!g87)) + ((g4) & (!g2) & (!g70) & (g80) & (g82) & (g87)) + ((g4) & (!g2) & (g70) & (!g80) & (g82) & (!g87)) + ((g4) & (!g2) & (g70) & (!g80) & (g82) & (g87)) + ((g4) & (!g2) & (g70) & (g80) & (!g82) & (!g87)) + ((g4) & (!g2) & (g70) & (g80) & (g82) & (g87)) + ((g4) & (g2) & (!g70) & (!g80) & (g82) & (!g87)) + ((g4) & (g2) & (!g70) & (!g80) & (g82) & (g87)) + ((g4) & (g2) & (!g70) & (g80) & (!g82) & (!g87)) + ((g4) & (g2) & (!g70) & (g80) & (g82) & (g87)) + ((g4) & (g2) & (g70) & (!g80) & (!g82) & (!g87)) + ((g4) & (g2) & (g70) & (!g80) & (g82) & (g87)) + ((g4) & (g2) & (g70) & (g80) & (!g82) & (!g87)) + ((g4) & (g2) & (g70) & (g80) & (g82) & (g87)));
	assign g90 = (((!g8) & (!g18) & (!g72) & (g73) & (g79) & (!g87)) + ((!g8) & (!g18) & (g72) & (!g73) & (!g79) & (!g87)) + ((!g8) & (!g18) & (g72) & (!g73) & (!g79) & (g87)) + ((!g8) & (!g18) & (g72) & (!g73) & (g79) & (!g87)) + ((!g8) & (!g18) & (g72) & (!g73) & (g79) & (g87)) + ((!g8) & (!g18) & (g72) & (g73) & (!g79) & (!g87)) + ((!g8) & (!g18) & (g72) & (g73) & (!g79) & (g87)) + ((!g8) & (!g18) & (g72) & (g73) & (g79) & (g87)) + ((!g8) & (g18) & (!g72) & (!g73) & (g79) & (!g87)) + ((!g8) & (g18) & (!g72) & (g73) & (!g79) & (!g87)) + ((!g8) & (g18) & (!g72) & (g73) & (g79) & (!g87)) + ((!g8) & (g18) & (g72) & (!g73) & (!g79) & (!g87)) + ((!g8) & (g18) & (g72) & (!g73) & (!g79) & (g87)) + ((!g8) & (g18) & (g72) & (!g73) & (g79) & (g87)) + ((!g8) & (g18) & (g72) & (g73) & (!g79) & (g87)) + ((!g8) & (g18) & (g72) & (g73) & (g79) & (g87)) + ((g8) & (!g18) & (!g72) & (!g73) & (!g79) & (!g87)) + ((g8) & (!g18) & (!g72) & (!g73) & (g79) & (!g87)) + ((g8) & (!g18) & (!g72) & (g73) & (!g79) & (!g87)) + ((g8) & (!g18) & (g72) & (!g73) & (!g79) & (g87)) + ((g8) & (!g18) & (g72) & (!g73) & (g79) & (g87)) + ((g8) & (!g18) & (g72) & (g73) & (!g79) & (g87)) + ((g8) & (!g18) & (g72) & (g73) & (g79) & (!g87)) + ((g8) & (!g18) & (g72) & (g73) & (g79) & (g87)) + ((g8) & (g18) & (!g72) & (!g73) & (!g79) & (!g87)) + ((g8) & (g18) & (g72) & (!g73) & (!g79) & (g87)) + ((g8) & (g18) & (g72) & (!g73) & (g79) & (!g87)) + ((g8) & (g18) & (g72) & (!g73) & (g79) & (g87)) + ((g8) & (g18) & (g72) & (g73) & (!g79) & (!g87)) + ((g8) & (g18) & (g72) & (g73) & (!g79) & (g87)) + ((g8) & (g18) & (g72) & (g73) & (g79) & (!g87)) + ((g8) & (g18) & (g72) & (g73) & (g79) & (g87)));
	assign g91 = (((!g18) & (!g73) & (g79) & (!g87)) + ((!g18) & (g73) & (!g79) & (!g87)) + ((!g18) & (g73) & (!g79) & (g87)) + ((!g18) & (g73) & (g79) & (g87)) + ((g18) & (!g73) & (!g79) & (!g87)) + ((g18) & (g73) & (!g79) & (g87)) + ((g18) & (g73) & (g79) & (!g87)) + ((g18) & (g73) & (g79) & (g87)));
	assign g92 = (((!g27) & (!g39) & (!g75) & (g76) & (g78) & (!g87)) + ((!g27) & (!g39) & (g75) & (!g76) & (!g78) & (!g87)) + ((!g27) & (!g39) & (g75) & (!g76) & (!g78) & (g87)) + ((!g27) & (!g39) & (g75) & (!g76) & (g78) & (!g87)) + ((!g27) & (!g39) & (g75) & (!g76) & (g78) & (g87)) + ((!g27) & (!g39) & (g75) & (g76) & (!g78) & (!g87)) + ((!g27) & (!g39) & (g75) & (g76) & (!g78) & (g87)) + ((!g27) & (!g39) & (g75) & (g76) & (g78) & (g87)) + ((!g27) & (g39) & (!g75) & (!g76) & (g78) & (!g87)) + ((!g27) & (g39) & (!g75) & (g76) & (!g78) & (!g87)) + ((!g27) & (g39) & (!g75) & (g76) & (g78) & (!g87)) + ((!g27) & (g39) & (g75) & (!g76) & (!g78) & (!g87)) + ((!g27) & (g39) & (g75) & (!g76) & (!g78) & (g87)) + ((!g27) & (g39) & (g75) & (!g76) & (g78) & (g87)) + ((!g27) & (g39) & (g75) & (g76) & (!g78) & (g87)) + ((!g27) & (g39) & (g75) & (g76) & (g78) & (g87)) + ((g27) & (!g39) & (!g75) & (!g76) & (!g78) & (!g87)) + ((g27) & (!g39) & (!g75) & (!g76) & (g78) & (!g87)) + ((g27) & (!g39) & (!g75) & (g76) & (!g78) & (!g87)) + ((g27) & (!g39) & (g75) & (!g76) & (!g78) & (g87)) + ((g27) & (!g39) & (g75) & (!g76) & (g78) & (g87)) + ((g27) & (!g39) & (g75) & (g76) & (!g78) & (g87)) + ((g27) & (!g39) & (g75) & (g76) & (g78) & (!g87)) + ((g27) & (!g39) & (g75) & (g76) & (g78) & (g87)) + ((g27) & (g39) & (!g75) & (!g76) & (!g78) & (!g87)) + ((g27) & (g39) & (g75) & (!g76) & (!g78) & (g87)) + ((g27) & (g39) & (g75) & (!g76) & (g78) & (!g87)) + ((g27) & (g39) & (g75) & (!g76) & (g78) & (g87)) + ((g27) & (g39) & (g75) & (g76) & (!g78) & (!g87)) + ((g27) & (g39) & (g75) & (g76) & (!g78) & (g87)) + ((g27) & (g39) & (g75) & (g76) & (g78) & (!g87)) + ((g27) & (g39) & (g75) & (g76) & (g78) & (g87)));
	assign g93 = (((!g39) & (!g76) & (g78) & (!g87)) + ((!g39) & (g76) & (!g78) & (!g87)) + ((!g39) & (g76) & (!g78) & (g87)) + ((!g39) & (g76) & (g78) & (g87)) + ((g39) & (!g76) & (!g78) & (!g87)) + ((g39) & (g76) & (!g78) & (g87)) + ((g39) & (g76) & (g78) & (!g87)) + ((g39) & (g76) & (g78) & (g87)));
	assign g94 = (((!g54) & (!ax110x) & (!ax111x) & (!g68) & (!g77) & (g87)) + ((!g54) & (!ax110x) & (!ax111x) & (!g68) & (g77) & (!g87)) + ((!g54) & (!ax110x) & (!ax111x) & (!g68) & (g77) & (g87)) + ((!g54) & (!ax110x) & (!ax111x) & (g68) & (!g77) & (!g87)) + ((!g54) & (!ax110x) & (ax111x) & (!g68) & (!g77) & (!g87)) + ((!g54) & (!ax110x) & (ax111x) & (g68) & (!g77) & (g87)) + ((!g54) & (!ax110x) & (ax111x) & (g68) & (g77) & (!g87)) + ((!g54) & (!ax110x) & (ax111x) & (g68) & (g77) & (g87)) + ((!g54) & (ax110x) & (!ax111x) & (g68) & (!g77) & (!g87)) + ((!g54) & (ax110x) & (!ax111x) & (g68) & (g77) & (!g87)) + ((!g54) & (ax110x) & (ax111x) & (!g68) & (!g77) & (!g87)) + ((!g54) & (ax110x) & (ax111x) & (!g68) & (!g77) & (g87)) + ((!g54) & (ax110x) & (ax111x) & (!g68) & (g77) & (!g87)) + ((!g54) & (ax110x) & (ax111x) & (!g68) & (g77) & (g87)) + ((!g54) & (ax110x) & (ax111x) & (g68) & (!g77) & (g87)) + ((!g54) & (ax110x) & (ax111x) & (g68) & (g77) & (g87)) + ((g54) & (!ax110x) & (!ax111x) & (!g68) & (!g77) & (!g87)) + ((g54) & (!ax110x) & (!ax111x) & (!g68) & (!g77) & (g87)) + ((g54) & (!ax110x) & (!ax111x) & (!g68) & (g77) & (g87)) + ((g54) & (!ax110x) & (!ax111x) & (g68) & (g77) & (!g87)) + ((g54) & (!ax110x) & (ax111x) & (!g68) & (g77) & (!g87)) + ((g54) & (!ax110x) & (ax111x) & (g68) & (!g77) & (!g87)) + ((g54) & (!ax110x) & (ax111x) & (g68) & (!g77) & (g87)) + ((g54) & (!ax110x) & (ax111x) & (g68) & (g77) & (g87)) + ((g54) & (ax110x) & (!ax111x) & (!g68) & (!g77) & (!g87)) + ((g54) & (ax110x) & (!ax111x) & (!g68) & (g77) & (!g87)) + ((g54) & (ax110x) & (ax111x) & (!g68) & (!g77) & (g87)) + ((g54) & (ax110x) & (ax111x) & (!g68) & (g77) & (g87)) + ((g54) & (ax110x) & (ax111x) & (g68) & (!g77) & (!g87)) + ((g54) & (ax110x) & (ax111x) & (g68) & (!g77) & (g87)) + ((g54) & (ax110x) & (ax111x) & (g68) & (g77) & (!g87)) + ((g54) & (ax110x) & (ax111x) & (g68) & (g77) & (g87)));
	assign g95 = (((!ax110x) & (!g68) & (!g77) & (g87)) + ((!ax110x) & (!g68) & (g77) & (!g87)) + ((!ax110x) & (!g68) & (g77) & (g87)) + ((!ax110x) & (g68) & (g77) & (!g87)) + ((ax110x) & (!g68) & (!g77) & (!g87)) + ((ax110x) & (g68) & (!g77) & (!g87)) + ((ax110x) & (g68) & (!g77) & (g87)) + ((ax110x) & (g68) & (g77) & (g87)));
	assign g96 = (((!ax106x) & (!ax107x)));
	assign g97 = (((!g68) & (!ax108x) & (!ax109x) & (!g87) & (!g96)) + ((!g68) & (!ax108x) & (ax109x) & (g87) & (!g96)) + ((!g68) & (ax108x) & (ax109x) & (g87) & (!g96)) + ((!g68) & (ax108x) & (ax109x) & (g87) & (g96)) + ((g68) & (!ax108x) & (!ax109x) & (!g87) & (!g96)) + ((g68) & (!ax108x) & (!ax109x) & (!g87) & (g96)) + ((g68) & (!ax108x) & (!ax109x) & (g87) & (!g96)) + ((g68) & (!ax108x) & (ax109x) & (!g87) & (!g96)) + ((g68) & (!ax108x) & (ax109x) & (g87) & (!g96)) + ((g68) & (!ax108x) & (ax109x) & (g87) & (g96)) + ((g68) & (ax108x) & (!ax109x) & (g87) & (!g96)) + ((g68) & (ax108x) & (!ax109x) & (g87) & (g96)) + ((g68) & (ax108x) & (ax109x) & (!g87) & (!g96)) + ((g68) & (ax108x) & (ax109x) & (!g87) & (g96)) + ((g68) & (ax108x) & (ax109x) & (g87) & (!g96)) + ((g68) & (ax108x) & (ax109x) & (g87) & (g96)));
	assign g98 = (((!g39) & (!g54) & (g94) & (g95) & (g97)) + ((!g39) & (g54) & (g94) & (!g95) & (g97)) + ((!g39) & (g54) & (g94) & (g95) & (!g97)) + ((!g39) & (g54) & (g94) & (g95) & (g97)) + ((g39) & (!g54) & (!g94) & (g95) & (g97)) + ((g39) & (!g54) & (g94) & (!g95) & (!g97)) + ((g39) & (!g54) & (g94) & (!g95) & (g97)) + ((g39) & (!g54) & (g94) & (g95) & (!g97)) + ((g39) & (!g54) & (g94) & (g95) & (g97)) + ((g39) & (g54) & (!g94) & (!g95) & (g97)) + ((g39) & (g54) & (!g94) & (g95) & (!g97)) + ((g39) & (g54) & (!g94) & (g95) & (g97)) + ((g39) & (g54) & (g94) & (!g95) & (!g97)) + ((g39) & (g54) & (g94) & (!g95) & (g97)) + ((g39) & (g54) & (g94) & (g95) & (!g97)) + ((g39) & (g54) & (g94) & (g95) & (g97)));
	assign g99 = (((!g18) & (!g27) & (g92) & (g93) & (g98)) + ((!g18) & (g27) & (g92) & (!g93) & (g98)) + ((!g18) & (g27) & (g92) & (g93) & (!g98)) + ((!g18) & (g27) & (g92) & (g93) & (g98)) + ((g18) & (!g27) & (!g92) & (g93) & (g98)) + ((g18) & (!g27) & (g92) & (!g93) & (!g98)) + ((g18) & (!g27) & (g92) & (!g93) & (g98)) + ((g18) & (!g27) & (g92) & (g93) & (!g98)) + ((g18) & (!g27) & (g92) & (g93) & (g98)) + ((g18) & (g27) & (!g92) & (!g93) & (g98)) + ((g18) & (g27) & (!g92) & (g93) & (!g98)) + ((g18) & (g27) & (!g92) & (g93) & (g98)) + ((g18) & (g27) & (g92) & (!g93) & (!g98)) + ((g18) & (g27) & (g92) & (!g93) & (g98)) + ((g18) & (g27) & (g92) & (g93) & (!g98)) + ((g18) & (g27) & (g92) & (g93) & (g98)));
	assign g100 = (((!g2) & (!g8) & (g90) & (g91) & (g99)) + ((!g2) & (g8) & (g90) & (!g91) & (g99)) + ((!g2) & (g8) & (g90) & (g91) & (!g99)) + ((!g2) & (g8) & (g90) & (g91) & (g99)) + ((g2) & (!g8) & (!g90) & (g91) & (g99)) + ((g2) & (!g8) & (g90) & (!g91) & (!g99)) + ((g2) & (!g8) & (g90) & (!g91) & (g99)) + ((g2) & (!g8) & (g90) & (g91) & (!g99)) + ((g2) & (!g8) & (g90) & (g91) & (g99)) + ((g2) & (g8) & (!g90) & (!g91) & (g99)) + ((g2) & (g8) & (!g90) & (g91) & (!g99)) + ((g2) & (g8) & (!g90) & (g91) & (g99)) + ((g2) & (g8) & (g90) & (!g91) & (!g99)) + ((g2) & (g8) & (g90) & (!g91) & (g99)) + ((g2) & (g8) & (g90) & (g91) & (!g99)) + ((g2) & (g8) & (g90) & (g91) & (g99)));
	assign g101 = (((!g2) & (!g70) & (g80) & (!g87)) + ((!g2) & (g70) & (!g80) & (!g87)) + ((!g2) & (g70) & (!g80) & (g87)) + ((!g2) & (g70) & (g80) & (g87)) + ((g2) & (!g70) & (!g80) & (!g87)) + ((g2) & (g70) & (!g80) & (g87)) + ((g2) & (g70) & (g80) & (!g87)) + ((g2) & (g70) & (g80) & (g87)));
	assign g102 = (((!g1) & (!g69) & (!g83) & (!g85) & (g86)) + ((!g1) & (!g69) & (!g83) & (g85) & (!g86)) + ((!g1) & (!g69) & (!g83) & (g85) & (g86)) + ((!g1) & (g69) & (g83) & (!g85) & (!g86)) + ((!g1) & (g69) & (g83) & (!g85) & (g86)) + ((!g1) & (g69) & (g83) & (g85) & (!g86)) + ((!g1) & (g69) & (g83) & (g85) & (g86)) + ((g1) & (!g69) & (!g83) & (!g85) & (g86)) + ((g1) & (!g69) & (!g83) & (g85) & (g86)) + ((g1) & (g69) & (g83) & (!g85) & (!g86)) + ((g1) & (g69) & (g83) & (!g85) & (g86)) + ((g1) & (g69) & (g83) & (g85) & (!g86)) + ((g1) & (g69) & (g83) & (g85) & (g86)));
	assign g103 = (((!g4) & (!g1) & (!g89) & (!g100) & (!g101) & (!g102)) + ((!g4) & (g1) & (!g89) & (!g100) & (!g101) & (!g102)) + ((!g4) & (g1) & (!g89) & (!g100) & (!g101) & (g102)) + ((!g4) & (g1) & (!g89) & (!g100) & (g101) & (!g102)) + ((!g4) & (g1) & (!g89) & (!g100) & (g101) & (g102)) + ((!g4) & (g1) & (!g89) & (g100) & (!g101) & (!g102)) + ((!g4) & (g1) & (!g89) & (g100) & (!g101) & (g102)) + ((!g4) & (g1) & (!g89) & (g100) & (g101) & (!g102)) + ((!g4) & (g1) & (!g89) & (g100) & (g101) & (g102)) + ((!g4) & (g1) & (g89) & (!g100) & (!g101) & (!g102)) + ((!g4) & (g1) & (g89) & (!g100) & (!g101) & (g102)) + ((g4) & (!g1) & (!g89) & (!g100) & (!g101) & (!g102)) + ((g4) & (!g1) & (!g89) & (!g100) & (g101) & (!g102)) + ((g4) & (!g1) & (!g89) & (g100) & (!g101) & (!g102)) + ((g4) & (g1) & (!g89) & (!g100) & (!g101) & (!g102)) + ((g4) & (g1) & (!g89) & (!g100) & (!g101) & (g102)) + ((g4) & (g1) & (!g89) & (!g100) & (g101) & (!g102)) + ((g4) & (g1) & (!g89) & (!g100) & (g101) & (g102)) + ((g4) & (g1) & (!g89) & (g100) & (!g101) & (!g102)) + ((g4) & (g1) & (!g89) & (g100) & (!g101) & (g102)) + ((g4) & (g1) & (!g89) & (g100) & (g101) & (!g102)) + ((g4) & (g1) & (!g89) & (g100) & (g101) & (g102)) + ((g4) & (g1) & (g89) & (!g100) & (!g101) & (!g102)) + ((g4) & (g1) & (g89) & (!g100) & (!g101) & (g102)) + ((g4) & (g1) & (g89) & (!g100) & (g101) & (!g102)) + ((g4) & (g1) & (g89) & (!g100) & (g101) & (g102)) + ((g4) & (g1) & (g89) & (g100) & (!g101) & (!g102)) + ((g4) & (g1) & (g89) & (g100) & (!g101) & (g102)));
	assign g104 = (((!g88) & (g103)));
	assign g105 = (((!g4) & (!g100) & (!g101) & (!g88) & (!g103)) + ((!g4) & (!g100) & (!g101) & (g88) & (!g103)) + ((!g4) & (!g100) & (!g101) & (g88) & (g103)) + ((!g4) & (!g100) & (g101) & (!g88) & (g103)) + ((!g4) & (g100) & (g101) & (!g88) & (!g103)) + ((!g4) & (g100) & (g101) & (!g88) & (g103)) + ((!g4) & (g100) & (g101) & (g88) & (!g103)) + ((!g4) & (g100) & (g101) & (g88) & (g103)) + ((g4) & (!g100) & (g101) & (!g88) & (!g103)) + ((g4) & (!g100) & (g101) & (!g88) & (g103)) + ((g4) & (!g100) & (g101) & (g88) & (!g103)) + ((g4) & (!g100) & (g101) & (g88) & (g103)) + ((g4) & (g100) & (!g101) & (!g88) & (!g103)) + ((g4) & (g100) & (!g101) & (g88) & (!g103)) + ((g4) & (g100) & (!g101) & (g88) & (g103)) + ((g4) & (g100) & (g101) & (!g88) & (g103)));
	assign g106 = (((!g8) & (!g91) & (g99) & (!g88) & (!g103)) + ((!g8) & (!g91) & (g99) & (g88) & (!g103)) + ((!g8) & (!g91) & (g99) & (g88) & (g103)) + ((!g8) & (g91) & (!g99) & (!g88) & (!g103)) + ((!g8) & (g91) & (!g99) & (!g88) & (g103)) + ((!g8) & (g91) & (!g99) & (g88) & (!g103)) + ((!g8) & (g91) & (!g99) & (g88) & (g103)) + ((!g8) & (g91) & (g99) & (!g88) & (g103)) + ((g8) & (!g91) & (!g99) & (!g88) & (!g103)) + ((g8) & (!g91) & (!g99) & (g88) & (!g103)) + ((g8) & (!g91) & (!g99) & (g88) & (g103)) + ((g8) & (g91) & (!g99) & (!g88) & (g103)) + ((g8) & (g91) & (g99) & (!g88) & (!g103)) + ((g8) & (g91) & (g99) & (!g88) & (g103)) + ((g8) & (g91) & (g99) & (g88) & (!g103)) + ((g8) & (g91) & (g99) & (g88) & (g103)));
	assign g107 = (((!g18) & (!g27) & (g93) & (g98)) + ((!g18) & (g27) & (!g93) & (g98)) + ((!g18) & (g27) & (g93) & (!g98)) + ((!g18) & (g27) & (g93) & (g98)) + ((g18) & (!g27) & (!g93) & (!g98)) + ((g18) & (!g27) & (!g93) & (g98)) + ((g18) & (!g27) & (g93) & (!g98)) + ((g18) & (g27) & (!g93) & (!g98)));
	assign g108 = (((!g92) & (!g88) & (!g103) & (g107)) + ((!g92) & (g88) & (!g103) & (g107)) + ((!g92) & (g88) & (g103) & (g107)) + ((g92) & (!g88) & (!g103) & (!g107)) + ((g92) & (!g88) & (g103) & (!g107)) + ((g92) & (!g88) & (g103) & (g107)) + ((g92) & (g88) & (!g103) & (!g107)) + ((g92) & (g88) & (g103) & (!g107)));
	assign g109 = (((!g27) & (!g93) & (g98) & (!g88) & (!g103)) + ((!g27) & (!g93) & (g98) & (g88) & (!g103)) + ((!g27) & (!g93) & (g98) & (g88) & (g103)) + ((!g27) & (g93) & (!g98) & (!g88) & (!g103)) + ((!g27) & (g93) & (!g98) & (!g88) & (g103)) + ((!g27) & (g93) & (!g98) & (g88) & (!g103)) + ((!g27) & (g93) & (!g98) & (g88) & (g103)) + ((!g27) & (g93) & (g98) & (!g88) & (g103)) + ((g27) & (!g93) & (!g98) & (!g88) & (!g103)) + ((g27) & (!g93) & (!g98) & (g88) & (!g103)) + ((g27) & (!g93) & (!g98) & (g88) & (g103)) + ((g27) & (g93) & (!g98) & (!g88) & (g103)) + ((g27) & (g93) & (g98) & (!g88) & (!g103)) + ((g27) & (g93) & (g98) & (!g88) & (g103)) + ((g27) & (g93) & (g98) & (g88) & (!g103)) + ((g27) & (g93) & (g98) & (g88) & (g103)));
	assign g110 = (((!g39) & (!g54) & (g95) & (g97)) + ((!g39) & (g54) & (!g95) & (g97)) + ((!g39) & (g54) & (g95) & (!g97)) + ((!g39) & (g54) & (g95) & (g97)) + ((g39) & (!g54) & (!g95) & (!g97)) + ((g39) & (!g54) & (!g95) & (g97)) + ((g39) & (!g54) & (g95) & (!g97)) + ((g39) & (g54) & (!g95) & (!g97)));
	assign g111 = (((!g94) & (!g88) & (!g103) & (g110)) + ((!g94) & (g88) & (!g103) & (g110)) + ((!g94) & (g88) & (g103) & (g110)) + ((g94) & (!g88) & (!g103) & (!g110)) + ((g94) & (!g88) & (g103) & (!g110)) + ((g94) & (!g88) & (g103) & (g110)) + ((g94) & (g88) & (!g103) & (!g110)) + ((g94) & (g88) & (g103) & (!g110)));
	assign g112 = (((!g54) & (!g95) & (g97) & (!g88) & (!g103)) + ((!g54) & (!g95) & (g97) & (g88) & (!g103)) + ((!g54) & (!g95) & (g97) & (g88) & (g103)) + ((!g54) & (g95) & (!g97) & (!g88) & (!g103)) + ((!g54) & (g95) & (!g97) & (!g88) & (g103)) + ((!g54) & (g95) & (!g97) & (g88) & (!g103)) + ((!g54) & (g95) & (!g97) & (g88) & (g103)) + ((!g54) & (g95) & (g97) & (!g88) & (g103)) + ((g54) & (!g95) & (!g97) & (!g88) & (!g103)) + ((g54) & (!g95) & (!g97) & (g88) & (!g103)) + ((g54) & (!g95) & (!g97) & (g88) & (g103)) + ((g54) & (g95) & (!g97) & (!g88) & (g103)) + ((g54) & (g95) & (g97) & (!g88) & (!g103)) + ((g54) & (g95) & (g97) & (!g88) & (g103)) + ((g54) & (g95) & (g97) & (g88) & (!g103)) + ((g54) & (g95) & (g97) & (g88) & (g103)));
	assign g113 = (((!g68) & (!ax108x) & (!g87) & (g96)) + ((!g68) & (!ax108x) & (g87) & (g96)) + ((!g68) & (ax108x) & (!g87) & (!g96)) + ((!g68) & (ax108x) & (!g87) & (g96)) + ((g68) & (!ax108x) & (!g87) & (!g96)) + ((g68) & (!ax108x) & (g87) & (!g96)) + ((g68) & (ax108x) & (g87) & (!g96)) + ((g68) & (ax108x) & (g87) & (g96)));
	assign g114 = (((!ax108x) & (!ax109x) & (!g87) & (!g88) & (!g103) & (g113)) + ((!ax108x) & (!ax109x) & (!g87) & (!g88) & (g103) & (!g113)) + ((!ax108x) & (!ax109x) & (!g87) & (!g88) & (g103) & (g113)) + ((!ax108x) & (!ax109x) & (!g87) & (g88) & (!g103) & (g113)) + ((!ax108x) & (!ax109x) & (!g87) & (g88) & (g103) & (g113)) + ((!ax108x) & (!ax109x) & (g87) & (!g88) & (!g103) & (!g113)) + ((!ax108x) & (!ax109x) & (g87) & (g88) & (!g103) & (!g113)) + ((!ax108x) & (!ax109x) & (g87) & (g88) & (g103) & (!g113)) + ((!ax108x) & (ax109x) & (!g87) & (!g88) & (!g103) & (!g113)) + ((!ax108x) & (ax109x) & (!g87) & (g88) & (!g103) & (!g113)) + ((!ax108x) & (ax109x) & (!g87) & (g88) & (g103) & (!g113)) + ((!ax108x) & (ax109x) & (g87) & (!g88) & (!g103) & (g113)) + ((!ax108x) & (ax109x) & (g87) & (!g88) & (g103) & (!g113)) + ((!ax108x) & (ax109x) & (g87) & (!g88) & (g103) & (g113)) + ((!ax108x) & (ax109x) & (g87) & (g88) & (!g103) & (g113)) + ((!ax108x) & (ax109x) & (g87) & (g88) & (g103) & (g113)) + ((ax108x) & (!ax109x) & (!g87) & (!g88) & (!g103) & (!g113)) + ((ax108x) & (!ax109x) & (!g87) & (g88) & (!g103) & (!g113)) + ((ax108x) & (!ax109x) & (!g87) & (g88) & (g103) & (!g113)) + ((ax108x) & (!ax109x) & (g87) & (!g88) & (!g103) & (!g113)) + ((ax108x) & (!ax109x) & (g87) & (g88) & (!g103) & (!g113)) + ((ax108x) & (!ax109x) & (g87) & (g88) & (g103) & (!g113)) + ((ax108x) & (ax109x) & (!g87) & (!g88) & (!g103) & (g113)) + ((ax108x) & (ax109x) & (!g87) & (!g88) & (g103) & (!g113)) + ((ax108x) & (ax109x) & (!g87) & (!g88) & (g103) & (g113)) + ((ax108x) & (ax109x) & (!g87) & (g88) & (!g103) & (g113)) + ((ax108x) & (ax109x) & (!g87) & (g88) & (g103) & (g113)) + ((ax108x) & (ax109x) & (g87) & (!g88) & (!g103) & (g113)) + ((ax108x) & (ax109x) & (g87) & (!g88) & (g103) & (!g113)) + ((ax108x) & (ax109x) & (g87) & (!g88) & (g103) & (g113)) + ((ax108x) & (ax109x) & (g87) & (g88) & (!g103) & (g113)) + ((ax108x) & (ax109x) & (g87) & (g88) & (g103) & (g113)));
	assign g115 = (((!ax108x) & (!g87) & (!g96) & (!g88) & (g103)) + ((!ax108x) & (!g87) & (g96) & (!g88) & (!g103)) + ((!ax108x) & (!g87) & (g96) & (!g88) & (g103)) + ((!ax108x) & (!g87) & (g96) & (g88) & (!g103)) + ((!ax108x) & (!g87) & (g96) & (g88) & (g103)) + ((!ax108x) & (g87) & (g96) & (!g88) & (!g103)) + ((!ax108x) & (g87) & (g96) & (g88) & (!g103)) + ((!ax108x) & (g87) & (g96) & (g88) & (g103)) + ((ax108x) & (!g87) & (!g96) & (!g88) & (!g103)) + ((ax108x) & (!g87) & (!g96) & (g88) & (!g103)) + ((ax108x) & (!g87) & (!g96) & (g88) & (g103)) + ((ax108x) & (g87) & (!g96) & (!g88) & (!g103)) + ((ax108x) & (g87) & (!g96) & (!g88) & (g103)) + ((ax108x) & (g87) & (!g96) & (g88) & (!g103)) + ((ax108x) & (g87) & (!g96) & (g88) & (g103)) + ((ax108x) & (g87) & (g96) & (!g88) & (g103)));
	assign g116 = (((!ax104x) & (!ax105x)));
	assign g117 = (((!g87) & (!ax106x) & (!ax107x) & (!g88) & (!g103) & (!g116)) + ((!g87) & (!ax106x) & (!ax107x) & (g88) & (!g103) & (!g116)) + ((!g87) & (!ax106x) & (!ax107x) & (g88) & (g103) & (!g116)) + ((!g87) & (!ax106x) & (ax107x) & (!g88) & (g103) & (!g116)) + ((!g87) & (ax106x) & (ax107x) & (!g88) & (g103) & (!g116)) + ((!g87) & (ax106x) & (ax107x) & (!g88) & (g103) & (g116)) + ((g87) & (!ax106x) & (!ax107x) & (!g88) & (!g103) & (!g116)) + ((g87) & (!ax106x) & (!ax107x) & (!g88) & (!g103) & (g116)) + ((g87) & (!ax106x) & (!ax107x) & (!g88) & (g103) & (!g116)) + ((g87) & (!ax106x) & (!ax107x) & (g88) & (!g103) & (!g116)) + ((g87) & (!ax106x) & (!ax107x) & (g88) & (!g103) & (g116)) + ((g87) & (!ax106x) & (!ax107x) & (g88) & (g103) & (!g116)) + ((g87) & (!ax106x) & (!ax107x) & (g88) & (g103) & (g116)) + ((g87) & (!ax106x) & (ax107x) & (!g88) & (!g103) & (!g116)) + ((g87) & (!ax106x) & (ax107x) & (!g88) & (g103) & (!g116)) + ((g87) & (!ax106x) & (ax107x) & (!g88) & (g103) & (g116)) + ((g87) & (!ax106x) & (ax107x) & (g88) & (!g103) & (!g116)) + ((g87) & (!ax106x) & (ax107x) & (g88) & (g103) & (!g116)) + ((g87) & (ax106x) & (!ax107x) & (!g88) & (g103) & (!g116)) + ((g87) & (ax106x) & (!ax107x) & (!g88) & (g103) & (g116)) + ((g87) & (ax106x) & (ax107x) & (!g88) & (!g103) & (!g116)) + ((g87) & (ax106x) & (ax107x) & (!g88) & (!g103) & (g116)) + ((g87) & (ax106x) & (ax107x) & (!g88) & (g103) & (!g116)) + ((g87) & (ax106x) & (ax107x) & (!g88) & (g103) & (g116)) + ((g87) & (ax106x) & (ax107x) & (g88) & (!g103) & (!g116)) + ((g87) & (ax106x) & (ax107x) & (g88) & (!g103) & (g116)) + ((g87) & (ax106x) & (ax107x) & (g88) & (g103) & (!g116)) + ((g87) & (ax106x) & (ax107x) & (g88) & (g103) & (g116)));
	assign g118 = (((!g54) & (!g68) & (g114) & (g115) & (g117)) + ((!g54) & (g68) & (g114) & (!g115) & (g117)) + ((!g54) & (g68) & (g114) & (g115) & (!g117)) + ((!g54) & (g68) & (g114) & (g115) & (g117)) + ((g54) & (!g68) & (!g114) & (g115) & (g117)) + ((g54) & (!g68) & (g114) & (!g115) & (!g117)) + ((g54) & (!g68) & (g114) & (!g115) & (g117)) + ((g54) & (!g68) & (g114) & (g115) & (!g117)) + ((g54) & (!g68) & (g114) & (g115) & (g117)) + ((g54) & (g68) & (!g114) & (!g115) & (g117)) + ((g54) & (g68) & (!g114) & (g115) & (!g117)) + ((g54) & (g68) & (!g114) & (g115) & (g117)) + ((g54) & (g68) & (g114) & (!g115) & (!g117)) + ((g54) & (g68) & (g114) & (!g115) & (g117)) + ((g54) & (g68) & (g114) & (g115) & (!g117)) + ((g54) & (g68) & (g114) & (g115) & (g117)));
	assign g119 = (((!g27) & (!g39) & (g111) & (g112) & (g118)) + ((!g27) & (g39) & (g111) & (!g112) & (g118)) + ((!g27) & (g39) & (g111) & (g112) & (!g118)) + ((!g27) & (g39) & (g111) & (g112) & (g118)) + ((g27) & (!g39) & (!g111) & (g112) & (g118)) + ((g27) & (!g39) & (g111) & (!g112) & (!g118)) + ((g27) & (!g39) & (g111) & (!g112) & (g118)) + ((g27) & (!g39) & (g111) & (g112) & (!g118)) + ((g27) & (!g39) & (g111) & (g112) & (g118)) + ((g27) & (g39) & (!g111) & (!g112) & (g118)) + ((g27) & (g39) & (!g111) & (g112) & (!g118)) + ((g27) & (g39) & (!g111) & (g112) & (g118)) + ((g27) & (g39) & (g111) & (!g112) & (!g118)) + ((g27) & (g39) & (g111) & (!g112) & (g118)) + ((g27) & (g39) & (g111) & (g112) & (!g118)) + ((g27) & (g39) & (g111) & (g112) & (g118)));
	assign g120 = (((!g8) & (!g18) & (g108) & (g109) & (g119)) + ((!g8) & (g18) & (g108) & (!g109) & (g119)) + ((!g8) & (g18) & (g108) & (g109) & (!g119)) + ((!g8) & (g18) & (g108) & (g109) & (g119)) + ((g8) & (!g18) & (!g108) & (g109) & (g119)) + ((g8) & (!g18) & (g108) & (!g109) & (!g119)) + ((g8) & (!g18) & (g108) & (!g109) & (g119)) + ((g8) & (!g18) & (g108) & (g109) & (!g119)) + ((g8) & (!g18) & (g108) & (g109) & (g119)) + ((g8) & (g18) & (!g108) & (!g109) & (g119)) + ((g8) & (g18) & (!g108) & (g109) & (!g119)) + ((g8) & (g18) & (!g108) & (g109) & (g119)) + ((g8) & (g18) & (g108) & (!g109) & (!g119)) + ((g8) & (g18) & (g108) & (!g109) & (g119)) + ((g8) & (g18) & (g108) & (g109) & (!g119)) + ((g8) & (g18) & (g108) & (g109) & (g119)));
	assign g121 = (((!g2) & (!g8) & (g91) & (g99)) + ((!g2) & (g8) & (!g91) & (g99)) + ((!g2) & (g8) & (g91) & (!g99)) + ((!g2) & (g8) & (g91) & (g99)) + ((g2) & (!g8) & (!g91) & (!g99)) + ((g2) & (!g8) & (!g91) & (g99)) + ((g2) & (!g8) & (g91) & (!g99)) + ((g2) & (g8) & (!g91) & (!g99)));
	assign g122 = (((!g90) & (!g88) & (!g103) & (g121)) + ((!g90) & (g88) & (!g103) & (g121)) + ((!g90) & (g88) & (g103) & (g121)) + ((g90) & (!g88) & (!g103) & (!g121)) + ((g90) & (!g88) & (g103) & (!g121)) + ((g90) & (!g88) & (g103) & (g121)) + ((g90) & (g88) & (!g103) & (!g121)) + ((g90) & (g88) & (g103) & (!g121)));
	assign g123 = (((!g4) & (!g2) & (!g106) & (!g120) & (g122)) + ((!g4) & (!g2) & (!g106) & (g120) & (g122)) + ((!g4) & (!g2) & (g106) & (!g120) & (g122)) + ((!g4) & (!g2) & (g106) & (g120) & (!g122)) + ((!g4) & (!g2) & (g106) & (g120) & (g122)) + ((!g4) & (g2) & (!g106) & (!g120) & (g122)) + ((!g4) & (g2) & (!g106) & (g120) & (!g122)) + ((!g4) & (g2) & (!g106) & (g120) & (g122)) + ((!g4) & (g2) & (g106) & (!g120) & (!g122)) + ((!g4) & (g2) & (g106) & (!g120) & (g122)) + ((!g4) & (g2) & (g106) & (g120) & (!g122)) + ((!g4) & (g2) & (g106) & (g120) & (g122)) + ((g4) & (!g2) & (g106) & (g120) & (g122)) + ((g4) & (g2) & (!g106) & (g120) & (g122)) + ((g4) & (g2) & (g106) & (!g120) & (g122)) + ((g4) & (g2) & (g106) & (g120) & (g122)));
	assign g124 = (((!g4) & (!g100) & (g101)) + ((!g4) & (g100) & (!g101)) + ((!g4) & (g100) & (g101)) + ((g4) & (g100) & (g101)));
	assign g125 = (((!g89) & (!g124) & (!g88) & (!g103)) + ((!g89) & (!g124) & (g88) & (!g103)) + ((!g89) & (!g124) & (g88) & (g103)) + ((g89) & (g124) & (!g88) & (!g103)) + ((g89) & (g124) & (!g88) & (g103)) + ((g89) & (g124) & (g88) & (!g103)) + ((g89) & (g124) & (g88) & (g103)));
	assign g126 = (((!g1) & (g89) & (!g124) & (!g88) & (g103)) + ((!g1) & (g89) & (g124) & (!g88) & (g103)) + ((g1) & (!g89) & (g124) & (g88) & (!g103)) + ((g1) & (!g89) & (g124) & (g88) & (g103)) + ((g1) & (g89) & (!g124) & (!g88) & (!g103)) + ((g1) & (g89) & (!g124) & (!g88) & (g103)) + ((g1) & (g89) & (!g124) & (g88) & (!g103)) + ((g1) & (g89) & (!g124) & (g88) & (g103)) + ((g1) & (g89) & (g124) & (!g88) & (g103)));
	assign g127 = (((!g1) & (!g105) & (!g123) & (!g125) & (!g126)) + ((g1) & (!g105) & (!g123) & (!g125) & (!g126)) + ((g1) & (!g105) & (!g123) & (g125) & (!g126)) + ((g1) & (!g105) & (g123) & (!g125) & (!g126)) + ((g1) & (!g105) & (g123) & (g125) & (!g126)) + ((g1) & (g105) & (!g123) & (!g125) & (!g126)) + ((g1) & (g105) & (!g123) & (g125) & (!g126)));
	assign g128 = (((g1) & (!g105) & (g123) & (g126)) + ((g1) & (g105) & (!g123) & (!g126)) + ((g1) & (g105) & (!g123) & (g126)));
	assign g129 = (((!g4) & (!g2) & (!g106) & (!g120) & (!g122) & (!g127)) + ((!g4) & (!g2) & (!g106) & (!g120) & (g122) & (g127)) + ((!g4) & (!g2) & (!g106) & (g120) & (!g122) & (!g127)) + ((!g4) & (!g2) & (!g106) & (g120) & (g122) & (g127)) + ((!g4) & (!g2) & (g106) & (!g120) & (!g122) & (!g127)) + ((!g4) & (!g2) & (g106) & (!g120) & (g122) & (g127)) + ((!g4) & (!g2) & (g106) & (g120) & (g122) & (!g127)) + ((!g4) & (!g2) & (g106) & (g120) & (g122) & (g127)) + ((!g4) & (g2) & (!g106) & (!g120) & (!g122) & (!g127)) + ((!g4) & (g2) & (!g106) & (!g120) & (g122) & (g127)) + ((!g4) & (g2) & (!g106) & (g120) & (g122) & (!g127)) + ((!g4) & (g2) & (!g106) & (g120) & (g122) & (g127)) + ((!g4) & (g2) & (g106) & (!g120) & (g122) & (!g127)) + ((!g4) & (g2) & (g106) & (!g120) & (g122) & (g127)) + ((!g4) & (g2) & (g106) & (g120) & (g122) & (!g127)) + ((!g4) & (g2) & (g106) & (g120) & (g122) & (g127)) + ((g4) & (!g2) & (!g106) & (!g120) & (g122) & (!g127)) + ((g4) & (!g2) & (!g106) & (!g120) & (g122) & (g127)) + ((g4) & (!g2) & (!g106) & (g120) & (g122) & (!g127)) + ((g4) & (!g2) & (!g106) & (g120) & (g122) & (g127)) + ((g4) & (!g2) & (g106) & (!g120) & (g122) & (!g127)) + ((g4) & (!g2) & (g106) & (!g120) & (g122) & (g127)) + ((g4) & (!g2) & (g106) & (g120) & (!g122) & (!g127)) + ((g4) & (!g2) & (g106) & (g120) & (g122) & (g127)) + ((g4) & (g2) & (!g106) & (!g120) & (g122) & (!g127)) + ((g4) & (g2) & (!g106) & (!g120) & (g122) & (g127)) + ((g4) & (g2) & (!g106) & (g120) & (!g122) & (!g127)) + ((g4) & (g2) & (!g106) & (g120) & (g122) & (g127)) + ((g4) & (g2) & (g106) & (!g120) & (!g122) & (!g127)) + ((g4) & (g2) & (g106) & (!g120) & (g122) & (g127)) + ((g4) & (g2) & (g106) & (g120) & (!g122) & (!g127)) + ((g4) & (g2) & (g106) & (g120) & (g122) & (g127)));
	assign g130 = (((!g8) & (!g18) & (!g108) & (g109) & (g119) & (!g127)) + ((!g8) & (!g18) & (g108) & (!g109) & (!g119) & (!g127)) + ((!g8) & (!g18) & (g108) & (!g109) & (!g119) & (g127)) + ((!g8) & (!g18) & (g108) & (!g109) & (g119) & (!g127)) + ((!g8) & (!g18) & (g108) & (!g109) & (g119) & (g127)) + ((!g8) & (!g18) & (g108) & (g109) & (!g119) & (!g127)) + ((!g8) & (!g18) & (g108) & (g109) & (!g119) & (g127)) + ((!g8) & (!g18) & (g108) & (g109) & (g119) & (g127)) + ((!g8) & (g18) & (!g108) & (!g109) & (g119) & (!g127)) + ((!g8) & (g18) & (!g108) & (g109) & (!g119) & (!g127)) + ((!g8) & (g18) & (!g108) & (g109) & (g119) & (!g127)) + ((!g8) & (g18) & (g108) & (!g109) & (!g119) & (!g127)) + ((!g8) & (g18) & (g108) & (!g109) & (!g119) & (g127)) + ((!g8) & (g18) & (g108) & (!g109) & (g119) & (g127)) + ((!g8) & (g18) & (g108) & (g109) & (!g119) & (g127)) + ((!g8) & (g18) & (g108) & (g109) & (g119) & (g127)) + ((g8) & (!g18) & (!g108) & (!g109) & (!g119) & (!g127)) + ((g8) & (!g18) & (!g108) & (!g109) & (g119) & (!g127)) + ((g8) & (!g18) & (!g108) & (g109) & (!g119) & (!g127)) + ((g8) & (!g18) & (g108) & (!g109) & (!g119) & (g127)) + ((g8) & (!g18) & (g108) & (!g109) & (g119) & (g127)) + ((g8) & (!g18) & (g108) & (g109) & (!g119) & (g127)) + ((g8) & (!g18) & (g108) & (g109) & (g119) & (!g127)) + ((g8) & (!g18) & (g108) & (g109) & (g119) & (g127)) + ((g8) & (g18) & (!g108) & (!g109) & (!g119) & (!g127)) + ((g8) & (g18) & (g108) & (!g109) & (!g119) & (g127)) + ((g8) & (g18) & (g108) & (!g109) & (g119) & (!g127)) + ((g8) & (g18) & (g108) & (!g109) & (g119) & (g127)) + ((g8) & (g18) & (g108) & (g109) & (!g119) & (!g127)) + ((g8) & (g18) & (g108) & (g109) & (!g119) & (g127)) + ((g8) & (g18) & (g108) & (g109) & (g119) & (!g127)) + ((g8) & (g18) & (g108) & (g109) & (g119) & (g127)));
	assign g131 = (((!g18) & (!g109) & (g119) & (!g127)) + ((!g18) & (g109) & (!g119) & (!g127)) + ((!g18) & (g109) & (!g119) & (g127)) + ((!g18) & (g109) & (g119) & (g127)) + ((g18) & (!g109) & (!g119) & (!g127)) + ((g18) & (g109) & (!g119) & (g127)) + ((g18) & (g109) & (g119) & (!g127)) + ((g18) & (g109) & (g119) & (g127)));
	assign g132 = (((!g27) & (!g39) & (!g111) & (g112) & (g118) & (!g127)) + ((!g27) & (!g39) & (g111) & (!g112) & (!g118) & (!g127)) + ((!g27) & (!g39) & (g111) & (!g112) & (!g118) & (g127)) + ((!g27) & (!g39) & (g111) & (!g112) & (g118) & (!g127)) + ((!g27) & (!g39) & (g111) & (!g112) & (g118) & (g127)) + ((!g27) & (!g39) & (g111) & (g112) & (!g118) & (!g127)) + ((!g27) & (!g39) & (g111) & (g112) & (!g118) & (g127)) + ((!g27) & (!g39) & (g111) & (g112) & (g118) & (g127)) + ((!g27) & (g39) & (!g111) & (!g112) & (g118) & (!g127)) + ((!g27) & (g39) & (!g111) & (g112) & (!g118) & (!g127)) + ((!g27) & (g39) & (!g111) & (g112) & (g118) & (!g127)) + ((!g27) & (g39) & (g111) & (!g112) & (!g118) & (!g127)) + ((!g27) & (g39) & (g111) & (!g112) & (!g118) & (g127)) + ((!g27) & (g39) & (g111) & (!g112) & (g118) & (g127)) + ((!g27) & (g39) & (g111) & (g112) & (!g118) & (g127)) + ((!g27) & (g39) & (g111) & (g112) & (g118) & (g127)) + ((g27) & (!g39) & (!g111) & (!g112) & (!g118) & (!g127)) + ((g27) & (!g39) & (!g111) & (!g112) & (g118) & (!g127)) + ((g27) & (!g39) & (!g111) & (g112) & (!g118) & (!g127)) + ((g27) & (!g39) & (g111) & (!g112) & (!g118) & (g127)) + ((g27) & (!g39) & (g111) & (!g112) & (g118) & (g127)) + ((g27) & (!g39) & (g111) & (g112) & (!g118) & (g127)) + ((g27) & (!g39) & (g111) & (g112) & (g118) & (!g127)) + ((g27) & (!g39) & (g111) & (g112) & (g118) & (g127)) + ((g27) & (g39) & (!g111) & (!g112) & (!g118) & (!g127)) + ((g27) & (g39) & (g111) & (!g112) & (!g118) & (g127)) + ((g27) & (g39) & (g111) & (!g112) & (g118) & (!g127)) + ((g27) & (g39) & (g111) & (!g112) & (g118) & (g127)) + ((g27) & (g39) & (g111) & (g112) & (!g118) & (!g127)) + ((g27) & (g39) & (g111) & (g112) & (!g118) & (g127)) + ((g27) & (g39) & (g111) & (g112) & (g118) & (!g127)) + ((g27) & (g39) & (g111) & (g112) & (g118) & (g127)));
	assign g133 = (((!g39) & (!g112) & (g118) & (!g127)) + ((!g39) & (g112) & (!g118) & (!g127)) + ((!g39) & (g112) & (!g118) & (g127)) + ((!g39) & (g112) & (g118) & (g127)) + ((g39) & (!g112) & (!g118) & (!g127)) + ((g39) & (g112) & (!g118) & (g127)) + ((g39) & (g112) & (g118) & (!g127)) + ((g39) & (g112) & (g118) & (g127)));
	assign g134 = (((!g54) & (!g68) & (!g114) & (g115) & (g117) & (!g127)) + ((!g54) & (!g68) & (g114) & (!g115) & (!g117) & (!g127)) + ((!g54) & (!g68) & (g114) & (!g115) & (!g117) & (g127)) + ((!g54) & (!g68) & (g114) & (!g115) & (g117) & (!g127)) + ((!g54) & (!g68) & (g114) & (!g115) & (g117) & (g127)) + ((!g54) & (!g68) & (g114) & (g115) & (!g117) & (!g127)) + ((!g54) & (!g68) & (g114) & (g115) & (!g117) & (g127)) + ((!g54) & (!g68) & (g114) & (g115) & (g117) & (g127)) + ((!g54) & (g68) & (!g114) & (!g115) & (g117) & (!g127)) + ((!g54) & (g68) & (!g114) & (g115) & (!g117) & (!g127)) + ((!g54) & (g68) & (!g114) & (g115) & (g117) & (!g127)) + ((!g54) & (g68) & (g114) & (!g115) & (!g117) & (!g127)) + ((!g54) & (g68) & (g114) & (!g115) & (!g117) & (g127)) + ((!g54) & (g68) & (g114) & (!g115) & (g117) & (g127)) + ((!g54) & (g68) & (g114) & (g115) & (!g117) & (g127)) + ((!g54) & (g68) & (g114) & (g115) & (g117) & (g127)) + ((g54) & (!g68) & (!g114) & (!g115) & (!g117) & (!g127)) + ((g54) & (!g68) & (!g114) & (!g115) & (g117) & (!g127)) + ((g54) & (!g68) & (!g114) & (g115) & (!g117) & (!g127)) + ((g54) & (!g68) & (g114) & (!g115) & (!g117) & (g127)) + ((g54) & (!g68) & (g114) & (!g115) & (g117) & (g127)) + ((g54) & (!g68) & (g114) & (g115) & (!g117) & (g127)) + ((g54) & (!g68) & (g114) & (g115) & (g117) & (!g127)) + ((g54) & (!g68) & (g114) & (g115) & (g117) & (g127)) + ((g54) & (g68) & (!g114) & (!g115) & (!g117) & (!g127)) + ((g54) & (g68) & (g114) & (!g115) & (!g117) & (g127)) + ((g54) & (g68) & (g114) & (!g115) & (g117) & (!g127)) + ((g54) & (g68) & (g114) & (!g115) & (g117) & (g127)) + ((g54) & (g68) & (g114) & (g115) & (!g117) & (!g127)) + ((g54) & (g68) & (g114) & (g115) & (!g117) & (g127)) + ((g54) & (g68) & (g114) & (g115) & (g117) & (!g127)) + ((g54) & (g68) & (g114) & (g115) & (g117) & (g127)));
	assign g135 = (((!g68) & (!g115) & (g117) & (!g127)) + ((!g68) & (g115) & (!g117) & (!g127)) + ((!g68) & (g115) & (!g117) & (g127)) + ((!g68) & (g115) & (g117) & (g127)) + ((g68) & (!g115) & (!g117) & (!g127)) + ((g68) & (g115) & (!g117) & (g127)) + ((g68) & (g115) & (g117) & (!g127)) + ((g68) & (g115) & (g117) & (g127)));
	assign g136 = (((!g87) & (!ax106x) & (!ax107x) & (!g104) & (!g116) & (g127)) + ((!g87) & (!ax106x) & (!ax107x) & (!g104) & (g116) & (!g127)) + ((!g87) & (!ax106x) & (!ax107x) & (!g104) & (g116) & (g127)) + ((!g87) & (!ax106x) & (!ax107x) & (g104) & (!g116) & (!g127)) + ((!g87) & (!ax106x) & (ax107x) & (!g104) & (!g116) & (!g127)) + ((!g87) & (!ax106x) & (ax107x) & (g104) & (!g116) & (g127)) + ((!g87) & (!ax106x) & (ax107x) & (g104) & (g116) & (!g127)) + ((!g87) & (!ax106x) & (ax107x) & (g104) & (g116) & (g127)) + ((!g87) & (ax106x) & (!ax107x) & (g104) & (!g116) & (!g127)) + ((!g87) & (ax106x) & (!ax107x) & (g104) & (g116) & (!g127)) + ((!g87) & (ax106x) & (ax107x) & (!g104) & (!g116) & (!g127)) + ((!g87) & (ax106x) & (ax107x) & (!g104) & (!g116) & (g127)) + ((!g87) & (ax106x) & (ax107x) & (!g104) & (g116) & (!g127)) + ((!g87) & (ax106x) & (ax107x) & (!g104) & (g116) & (g127)) + ((!g87) & (ax106x) & (ax107x) & (g104) & (!g116) & (g127)) + ((!g87) & (ax106x) & (ax107x) & (g104) & (g116) & (g127)) + ((g87) & (!ax106x) & (!ax107x) & (!g104) & (!g116) & (!g127)) + ((g87) & (!ax106x) & (!ax107x) & (!g104) & (!g116) & (g127)) + ((g87) & (!ax106x) & (!ax107x) & (!g104) & (g116) & (g127)) + ((g87) & (!ax106x) & (!ax107x) & (g104) & (g116) & (!g127)) + ((g87) & (!ax106x) & (ax107x) & (!g104) & (g116) & (!g127)) + ((g87) & (!ax106x) & (ax107x) & (g104) & (!g116) & (!g127)) + ((g87) & (!ax106x) & (ax107x) & (g104) & (!g116) & (g127)) + ((g87) & (!ax106x) & (ax107x) & (g104) & (g116) & (g127)) + ((g87) & (ax106x) & (!ax107x) & (!g104) & (!g116) & (!g127)) + ((g87) & (ax106x) & (!ax107x) & (!g104) & (g116) & (!g127)) + ((g87) & (ax106x) & (ax107x) & (!g104) & (!g116) & (g127)) + ((g87) & (ax106x) & (ax107x) & (!g104) & (g116) & (g127)) + ((g87) & (ax106x) & (ax107x) & (g104) & (!g116) & (!g127)) + ((g87) & (ax106x) & (ax107x) & (g104) & (!g116) & (g127)) + ((g87) & (ax106x) & (ax107x) & (g104) & (g116) & (!g127)) + ((g87) & (ax106x) & (ax107x) & (g104) & (g116) & (g127)));
	assign g137 = (((!ax106x) & (!g104) & (!g116) & (g127)) + ((!ax106x) & (!g104) & (g116) & (!g127)) + ((!ax106x) & (!g104) & (g116) & (g127)) + ((!ax106x) & (g104) & (g116) & (!g127)) + ((ax106x) & (!g104) & (!g116) & (!g127)) + ((ax106x) & (g104) & (!g116) & (!g127)) + ((ax106x) & (g104) & (!g116) & (g127)) + ((ax106x) & (g104) & (g116) & (g127)));
	assign g138 = (((!ax102x) & (!ax103x)));
	assign g139 = (((!g104) & (!ax104x) & (!ax105x) & (!g127) & (!g138)) + ((!g104) & (!ax104x) & (ax105x) & (g127) & (!g138)) + ((!g104) & (ax104x) & (ax105x) & (g127) & (!g138)) + ((!g104) & (ax104x) & (ax105x) & (g127) & (g138)) + ((g104) & (!ax104x) & (!ax105x) & (!g127) & (!g138)) + ((g104) & (!ax104x) & (!ax105x) & (!g127) & (g138)) + ((g104) & (!ax104x) & (!ax105x) & (g127) & (!g138)) + ((g104) & (!ax104x) & (ax105x) & (!g127) & (!g138)) + ((g104) & (!ax104x) & (ax105x) & (g127) & (!g138)) + ((g104) & (!ax104x) & (ax105x) & (g127) & (g138)) + ((g104) & (ax104x) & (!ax105x) & (g127) & (!g138)) + ((g104) & (ax104x) & (!ax105x) & (g127) & (g138)) + ((g104) & (ax104x) & (ax105x) & (!g127) & (!g138)) + ((g104) & (ax104x) & (ax105x) & (!g127) & (g138)) + ((g104) & (ax104x) & (ax105x) & (g127) & (!g138)) + ((g104) & (ax104x) & (ax105x) & (g127) & (g138)));
	assign g140 = (((!g68) & (!g87) & (g136) & (g137) & (g139)) + ((!g68) & (g87) & (g136) & (!g137) & (g139)) + ((!g68) & (g87) & (g136) & (g137) & (!g139)) + ((!g68) & (g87) & (g136) & (g137) & (g139)) + ((g68) & (!g87) & (!g136) & (g137) & (g139)) + ((g68) & (!g87) & (g136) & (!g137) & (!g139)) + ((g68) & (!g87) & (g136) & (!g137) & (g139)) + ((g68) & (!g87) & (g136) & (g137) & (!g139)) + ((g68) & (!g87) & (g136) & (g137) & (g139)) + ((g68) & (g87) & (!g136) & (!g137) & (g139)) + ((g68) & (g87) & (!g136) & (g137) & (!g139)) + ((g68) & (g87) & (!g136) & (g137) & (g139)) + ((g68) & (g87) & (g136) & (!g137) & (!g139)) + ((g68) & (g87) & (g136) & (!g137) & (g139)) + ((g68) & (g87) & (g136) & (g137) & (!g139)) + ((g68) & (g87) & (g136) & (g137) & (g139)));
	assign g141 = (((!g39) & (!g54) & (g134) & (g135) & (g140)) + ((!g39) & (g54) & (g134) & (!g135) & (g140)) + ((!g39) & (g54) & (g134) & (g135) & (!g140)) + ((!g39) & (g54) & (g134) & (g135) & (g140)) + ((g39) & (!g54) & (!g134) & (g135) & (g140)) + ((g39) & (!g54) & (g134) & (!g135) & (!g140)) + ((g39) & (!g54) & (g134) & (!g135) & (g140)) + ((g39) & (!g54) & (g134) & (g135) & (!g140)) + ((g39) & (!g54) & (g134) & (g135) & (g140)) + ((g39) & (g54) & (!g134) & (!g135) & (g140)) + ((g39) & (g54) & (!g134) & (g135) & (!g140)) + ((g39) & (g54) & (!g134) & (g135) & (g140)) + ((g39) & (g54) & (g134) & (!g135) & (!g140)) + ((g39) & (g54) & (g134) & (!g135) & (g140)) + ((g39) & (g54) & (g134) & (g135) & (!g140)) + ((g39) & (g54) & (g134) & (g135) & (g140)));
	assign g142 = (((!g18) & (!g27) & (g132) & (g133) & (g141)) + ((!g18) & (g27) & (g132) & (!g133) & (g141)) + ((!g18) & (g27) & (g132) & (g133) & (!g141)) + ((!g18) & (g27) & (g132) & (g133) & (g141)) + ((g18) & (!g27) & (!g132) & (g133) & (g141)) + ((g18) & (!g27) & (g132) & (!g133) & (!g141)) + ((g18) & (!g27) & (g132) & (!g133) & (g141)) + ((g18) & (!g27) & (g132) & (g133) & (!g141)) + ((g18) & (!g27) & (g132) & (g133) & (g141)) + ((g18) & (g27) & (!g132) & (!g133) & (g141)) + ((g18) & (g27) & (!g132) & (g133) & (!g141)) + ((g18) & (g27) & (!g132) & (g133) & (g141)) + ((g18) & (g27) & (g132) & (!g133) & (!g141)) + ((g18) & (g27) & (g132) & (!g133) & (g141)) + ((g18) & (g27) & (g132) & (g133) & (!g141)) + ((g18) & (g27) & (g132) & (g133) & (g141)));
	assign g143 = (((!g2) & (!g8) & (g130) & (g131) & (g142)) + ((!g2) & (g8) & (g130) & (!g131) & (g142)) + ((!g2) & (g8) & (g130) & (g131) & (!g142)) + ((!g2) & (g8) & (g130) & (g131) & (g142)) + ((g2) & (!g8) & (!g130) & (g131) & (g142)) + ((g2) & (!g8) & (g130) & (!g131) & (!g142)) + ((g2) & (!g8) & (g130) & (!g131) & (g142)) + ((g2) & (!g8) & (g130) & (g131) & (!g142)) + ((g2) & (!g8) & (g130) & (g131) & (g142)) + ((g2) & (g8) & (!g130) & (!g131) & (g142)) + ((g2) & (g8) & (!g130) & (g131) & (!g142)) + ((g2) & (g8) & (!g130) & (g131) & (g142)) + ((g2) & (g8) & (g130) & (!g131) & (!g142)) + ((g2) & (g8) & (g130) & (!g131) & (g142)) + ((g2) & (g8) & (g130) & (g131) & (!g142)) + ((g2) & (g8) & (g130) & (g131) & (g142)));
	assign g144 = (((!g2) & (!g106) & (g120) & (!g127)) + ((!g2) & (g106) & (!g120) & (!g127)) + ((!g2) & (g106) & (!g120) & (g127)) + ((!g2) & (g106) & (g120) & (g127)) + ((g2) & (!g106) & (!g120) & (!g127)) + ((g2) & (g106) & (!g120) & (g127)) + ((g2) & (g106) & (g120) & (!g127)) + ((g2) & (g106) & (g120) & (g127)));
	assign g145 = (((!g1) & (!g105) & (!g123) & (!g125) & (g126)) + ((!g1) & (!g105) & (!g123) & (g125) & (!g126)) + ((!g1) & (!g105) & (!g123) & (g125) & (g126)) + ((!g1) & (g105) & (g123) & (!g125) & (!g126)) + ((!g1) & (g105) & (g123) & (!g125) & (g126)) + ((!g1) & (g105) & (g123) & (g125) & (!g126)) + ((!g1) & (g105) & (g123) & (g125) & (g126)) + ((g1) & (!g105) & (!g123) & (!g125) & (g126)) + ((g1) & (!g105) & (!g123) & (g125) & (g126)) + ((g1) & (g105) & (g123) & (!g125) & (!g126)) + ((g1) & (g105) & (g123) & (!g125) & (g126)) + ((g1) & (g105) & (g123) & (g125) & (!g126)) + ((g1) & (g105) & (g123) & (g125) & (g126)));
	assign g146 = (((!g4) & (!g1) & (!g129) & (!g143) & (!g144) & (!g145)) + ((!g4) & (g1) & (!g129) & (!g143) & (!g144) & (!g145)) + ((!g4) & (g1) & (!g129) & (!g143) & (!g144) & (g145)) + ((!g4) & (g1) & (!g129) & (!g143) & (g144) & (!g145)) + ((!g4) & (g1) & (!g129) & (!g143) & (g144) & (g145)) + ((!g4) & (g1) & (!g129) & (g143) & (!g144) & (!g145)) + ((!g4) & (g1) & (!g129) & (g143) & (!g144) & (g145)) + ((!g4) & (g1) & (!g129) & (g143) & (g144) & (!g145)) + ((!g4) & (g1) & (!g129) & (g143) & (g144) & (g145)) + ((!g4) & (g1) & (g129) & (!g143) & (!g144) & (!g145)) + ((!g4) & (g1) & (g129) & (!g143) & (!g144) & (g145)) + ((g4) & (!g1) & (!g129) & (!g143) & (!g144) & (!g145)) + ((g4) & (!g1) & (!g129) & (!g143) & (g144) & (!g145)) + ((g4) & (!g1) & (!g129) & (g143) & (!g144) & (!g145)) + ((g4) & (g1) & (!g129) & (!g143) & (!g144) & (!g145)) + ((g4) & (g1) & (!g129) & (!g143) & (!g144) & (g145)) + ((g4) & (g1) & (!g129) & (!g143) & (g144) & (!g145)) + ((g4) & (g1) & (!g129) & (!g143) & (g144) & (g145)) + ((g4) & (g1) & (!g129) & (g143) & (!g144) & (!g145)) + ((g4) & (g1) & (!g129) & (g143) & (!g144) & (g145)) + ((g4) & (g1) & (!g129) & (g143) & (g144) & (!g145)) + ((g4) & (g1) & (!g129) & (g143) & (g144) & (g145)) + ((g4) & (g1) & (g129) & (!g143) & (!g144) & (!g145)) + ((g4) & (g1) & (g129) & (!g143) & (!g144) & (g145)) + ((g4) & (g1) & (g129) & (!g143) & (g144) & (!g145)) + ((g4) & (g1) & (g129) & (!g143) & (g144) & (g145)) + ((g4) & (g1) & (g129) & (g143) & (!g144) & (!g145)) + ((g4) & (g1) & (g129) & (g143) & (!g144) & (g145)));
	assign g147 = (((!g128) & (g146)));
	assign g148 = (((!g4) & (!g143) & (!g144) & (!g128) & (!g146)) + ((!g4) & (!g143) & (!g144) & (g128) & (!g146)) + ((!g4) & (!g143) & (!g144) & (g128) & (g146)) + ((!g4) & (!g143) & (g144) & (!g128) & (g146)) + ((!g4) & (g143) & (g144) & (!g128) & (!g146)) + ((!g4) & (g143) & (g144) & (!g128) & (g146)) + ((!g4) & (g143) & (g144) & (g128) & (!g146)) + ((!g4) & (g143) & (g144) & (g128) & (g146)) + ((g4) & (!g143) & (g144) & (!g128) & (!g146)) + ((g4) & (!g143) & (g144) & (!g128) & (g146)) + ((g4) & (!g143) & (g144) & (g128) & (!g146)) + ((g4) & (!g143) & (g144) & (g128) & (g146)) + ((g4) & (g143) & (!g144) & (!g128) & (!g146)) + ((g4) & (g143) & (!g144) & (g128) & (!g146)) + ((g4) & (g143) & (!g144) & (g128) & (g146)) + ((g4) & (g143) & (g144) & (!g128) & (g146)));
	assign g149 = (((!g2) & (!g8) & (g131) & (g142)) + ((!g2) & (g8) & (!g131) & (g142)) + ((!g2) & (g8) & (g131) & (!g142)) + ((!g2) & (g8) & (g131) & (g142)) + ((g2) & (!g8) & (!g131) & (!g142)) + ((g2) & (!g8) & (!g131) & (g142)) + ((g2) & (!g8) & (g131) & (!g142)) + ((g2) & (g8) & (!g131) & (!g142)));
	assign g150 = (((!g130) & (!g128) & (!g146) & (g149)) + ((!g130) & (g128) & (!g146) & (g149)) + ((!g130) & (g128) & (g146) & (g149)) + ((g130) & (!g128) & (!g146) & (!g149)) + ((g130) & (!g128) & (g146) & (!g149)) + ((g130) & (!g128) & (g146) & (g149)) + ((g130) & (g128) & (!g146) & (!g149)) + ((g130) & (g128) & (g146) & (!g149)));
	assign g151 = (((!g8) & (!g131) & (g142) & (!g128) & (!g146)) + ((!g8) & (!g131) & (g142) & (g128) & (!g146)) + ((!g8) & (!g131) & (g142) & (g128) & (g146)) + ((!g8) & (g131) & (!g142) & (!g128) & (!g146)) + ((!g8) & (g131) & (!g142) & (!g128) & (g146)) + ((!g8) & (g131) & (!g142) & (g128) & (!g146)) + ((!g8) & (g131) & (!g142) & (g128) & (g146)) + ((!g8) & (g131) & (g142) & (!g128) & (g146)) + ((g8) & (!g131) & (!g142) & (!g128) & (!g146)) + ((g8) & (!g131) & (!g142) & (g128) & (!g146)) + ((g8) & (!g131) & (!g142) & (g128) & (g146)) + ((g8) & (g131) & (!g142) & (!g128) & (g146)) + ((g8) & (g131) & (g142) & (!g128) & (!g146)) + ((g8) & (g131) & (g142) & (!g128) & (g146)) + ((g8) & (g131) & (g142) & (g128) & (!g146)) + ((g8) & (g131) & (g142) & (g128) & (g146)));
	assign g152 = (((!g18) & (!g27) & (g133) & (g141)) + ((!g18) & (g27) & (!g133) & (g141)) + ((!g18) & (g27) & (g133) & (!g141)) + ((!g18) & (g27) & (g133) & (g141)) + ((g18) & (!g27) & (!g133) & (!g141)) + ((g18) & (!g27) & (!g133) & (g141)) + ((g18) & (!g27) & (g133) & (!g141)) + ((g18) & (g27) & (!g133) & (!g141)));
	assign g153 = (((!g132) & (!g128) & (!g146) & (g152)) + ((!g132) & (g128) & (!g146) & (g152)) + ((!g132) & (g128) & (g146) & (g152)) + ((g132) & (!g128) & (!g146) & (!g152)) + ((g132) & (!g128) & (g146) & (!g152)) + ((g132) & (!g128) & (g146) & (g152)) + ((g132) & (g128) & (!g146) & (!g152)) + ((g132) & (g128) & (g146) & (!g152)));
	assign g154 = (((!g27) & (!g133) & (g141) & (!g128) & (!g146)) + ((!g27) & (!g133) & (g141) & (g128) & (!g146)) + ((!g27) & (!g133) & (g141) & (g128) & (g146)) + ((!g27) & (g133) & (!g141) & (!g128) & (!g146)) + ((!g27) & (g133) & (!g141) & (!g128) & (g146)) + ((!g27) & (g133) & (!g141) & (g128) & (!g146)) + ((!g27) & (g133) & (!g141) & (g128) & (g146)) + ((!g27) & (g133) & (g141) & (!g128) & (g146)) + ((g27) & (!g133) & (!g141) & (!g128) & (!g146)) + ((g27) & (!g133) & (!g141) & (g128) & (!g146)) + ((g27) & (!g133) & (!g141) & (g128) & (g146)) + ((g27) & (g133) & (!g141) & (!g128) & (g146)) + ((g27) & (g133) & (g141) & (!g128) & (!g146)) + ((g27) & (g133) & (g141) & (!g128) & (g146)) + ((g27) & (g133) & (g141) & (g128) & (!g146)) + ((g27) & (g133) & (g141) & (g128) & (g146)));
	assign g155 = (((!g39) & (!g54) & (g135) & (g140)) + ((!g39) & (g54) & (!g135) & (g140)) + ((!g39) & (g54) & (g135) & (!g140)) + ((!g39) & (g54) & (g135) & (g140)) + ((g39) & (!g54) & (!g135) & (!g140)) + ((g39) & (!g54) & (!g135) & (g140)) + ((g39) & (!g54) & (g135) & (!g140)) + ((g39) & (g54) & (!g135) & (!g140)));
	assign g156 = (((!g134) & (!g128) & (!g146) & (g155)) + ((!g134) & (g128) & (!g146) & (g155)) + ((!g134) & (g128) & (g146) & (g155)) + ((g134) & (!g128) & (!g146) & (!g155)) + ((g134) & (!g128) & (g146) & (!g155)) + ((g134) & (!g128) & (g146) & (g155)) + ((g134) & (g128) & (!g146) & (!g155)) + ((g134) & (g128) & (g146) & (!g155)));
	assign g157 = (((!g54) & (!g135) & (g140) & (!g128) & (!g146)) + ((!g54) & (!g135) & (g140) & (g128) & (!g146)) + ((!g54) & (!g135) & (g140) & (g128) & (g146)) + ((!g54) & (g135) & (!g140) & (!g128) & (!g146)) + ((!g54) & (g135) & (!g140) & (!g128) & (g146)) + ((!g54) & (g135) & (!g140) & (g128) & (!g146)) + ((!g54) & (g135) & (!g140) & (g128) & (g146)) + ((!g54) & (g135) & (g140) & (!g128) & (g146)) + ((g54) & (!g135) & (!g140) & (!g128) & (!g146)) + ((g54) & (!g135) & (!g140) & (g128) & (!g146)) + ((g54) & (!g135) & (!g140) & (g128) & (g146)) + ((g54) & (g135) & (!g140) & (!g128) & (g146)) + ((g54) & (g135) & (g140) & (!g128) & (!g146)) + ((g54) & (g135) & (g140) & (!g128) & (g146)) + ((g54) & (g135) & (g140) & (g128) & (!g146)) + ((g54) & (g135) & (g140) & (g128) & (g146)));
	assign g158 = (((!g68) & (!g87) & (g137) & (g139)) + ((!g68) & (g87) & (!g137) & (g139)) + ((!g68) & (g87) & (g137) & (!g139)) + ((!g68) & (g87) & (g137) & (g139)) + ((g68) & (!g87) & (!g137) & (!g139)) + ((g68) & (!g87) & (!g137) & (g139)) + ((g68) & (!g87) & (g137) & (!g139)) + ((g68) & (g87) & (!g137) & (!g139)));
	assign g159 = (((!g136) & (!g128) & (!g146) & (g158)) + ((!g136) & (g128) & (!g146) & (g158)) + ((!g136) & (g128) & (g146) & (g158)) + ((g136) & (!g128) & (!g146) & (!g158)) + ((g136) & (!g128) & (g146) & (!g158)) + ((g136) & (!g128) & (g146) & (g158)) + ((g136) & (g128) & (!g146) & (!g158)) + ((g136) & (g128) & (g146) & (!g158)));
	assign g160 = (((!g87) & (!g137) & (g139) & (!g128) & (!g146)) + ((!g87) & (!g137) & (g139) & (g128) & (!g146)) + ((!g87) & (!g137) & (g139) & (g128) & (g146)) + ((!g87) & (g137) & (!g139) & (!g128) & (!g146)) + ((!g87) & (g137) & (!g139) & (!g128) & (g146)) + ((!g87) & (g137) & (!g139) & (g128) & (!g146)) + ((!g87) & (g137) & (!g139) & (g128) & (g146)) + ((!g87) & (g137) & (g139) & (!g128) & (g146)) + ((g87) & (!g137) & (!g139) & (!g128) & (!g146)) + ((g87) & (!g137) & (!g139) & (g128) & (!g146)) + ((g87) & (!g137) & (!g139) & (g128) & (g146)) + ((g87) & (g137) & (!g139) & (!g128) & (g146)) + ((g87) & (g137) & (g139) & (!g128) & (!g146)) + ((g87) & (g137) & (g139) & (!g128) & (g146)) + ((g87) & (g137) & (g139) & (g128) & (!g146)) + ((g87) & (g137) & (g139) & (g128) & (g146)));
	assign g161 = (((!g104) & (!ax104x) & (!g127) & (g138)) + ((!g104) & (!ax104x) & (g127) & (g138)) + ((!g104) & (ax104x) & (!g127) & (!g138)) + ((!g104) & (ax104x) & (!g127) & (g138)) + ((g104) & (!ax104x) & (!g127) & (!g138)) + ((g104) & (!ax104x) & (g127) & (!g138)) + ((g104) & (ax104x) & (g127) & (!g138)) + ((g104) & (ax104x) & (g127) & (g138)));
	assign g162 = (((!ax104x) & (!ax105x) & (!g127) & (!g128) & (!g146) & (g161)) + ((!ax104x) & (!ax105x) & (!g127) & (!g128) & (g146) & (!g161)) + ((!ax104x) & (!ax105x) & (!g127) & (!g128) & (g146) & (g161)) + ((!ax104x) & (!ax105x) & (!g127) & (g128) & (!g146) & (g161)) + ((!ax104x) & (!ax105x) & (!g127) & (g128) & (g146) & (g161)) + ((!ax104x) & (!ax105x) & (g127) & (!g128) & (!g146) & (!g161)) + ((!ax104x) & (!ax105x) & (g127) & (g128) & (!g146) & (!g161)) + ((!ax104x) & (!ax105x) & (g127) & (g128) & (g146) & (!g161)) + ((!ax104x) & (ax105x) & (!g127) & (!g128) & (!g146) & (!g161)) + ((!ax104x) & (ax105x) & (!g127) & (g128) & (!g146) & (!g161)) + ((!ax104x) & (ax105x) & (!g127) & (g128) & (g146) & (!g161)) + ((!ax104x) & (ax105x) & (g127) & (!g128) & (!g146) & (g161)) + ((!ax104x) & (ax105x) & (g127) & (!g128) & (g146) & (!g161)) + ((!ax104x) & (ax105x) & (g127) & (!g128) & (g146) & (g161)) + ((!ax104x) & (ax105x) & (g127) & (g128) & (!g146) & (g161)) + ((!ax104x) & (ax105x) & (g127) & (g128) & (g146) & (g161)) + ((ax104x) & (!ax105x) & (!g127) & (!g128) & (!g146) & (!g161)) + ((ax104x) & (!ax105x) & (!g127) & (g128) & (!g146) & (!g161)) + ((ax104x) & (!ax105x) & (!g127) & (g128) & (g146) & (!g161)) + ((ax104x) & (!ax105x) & (g127) & (!g128) & (!g146) & (!g161)) + ((ax104x) & (!ax105x) & (g127) & (g128) & (!g146) & (!g161)) + ((ax104x) & (!ax105x) & (g127) & (g128) & (g146) & (!g161)) + ((ax104x) & (ax105x) & (!g127) & (!g128) & (!g146) & (g161)) + ((ax104x) & (ax105x) & (!g127) & (!g128) & (g146) & (!g161)) + ((ax104x) & (ax105x) & (!g127) & (!g128) & (g146) & (g161)) + ((ax104x) & (ax105x) & (!g127) & (g128) & (!g146) & (g161)) + ((ax104x) & (ax105x) & (!g127) & (g128) & (g146) & (g161)) + ((ax104x) & (ax105x) & (g127) & (!g128) & (!g146) & (g161)) + ((ax104x) & (ax105x) & (g127) & (!g128) & (g146) & (!g161)) + ((ax104x) & (ax105x) & (g127) & (!g128) & (g146) & (g161)) + ((ax104x) & (ax105x) & (g127) & (g128) & (!g146) & (g161)) + ((ax104x) & (ax105x) & (g127) & (g128) & (g146) & (g161)));
	assign g163 = (((!ax104x) & (!g127) & (!g138) & (!g128) & (g146)) + ((!ax104x) & (!g127) & (g138) & (!g128) & (!g146)) + ((!ax104x) & (!g127) & (g138) & (!g128) & (g146)) + ((!ax104x) & (!g127) & (g138) & (g128) & (!g146)) + ((!ax104x) & (!g127) & (g138) & (g128) & (g146)) + ((!ax104x) & (g127) & (g138) & (!g128) & (!g146)) + ((!ax104x) & (g127) & (g138) & (g128) & (!g146)) + ((!ax104x) & (g127) & (g138) & (g128) & (g146)) + ((ax104x) & (!g127) & (!g138) & (!g128) & (!g146)) + ((ax104x) & (!g127) & (!g138) & (g128) & (!g146)) + ((ax104x) & (!g127) & (!g138) & (g128) & (g146)) + ((ax104x) & (g127) & (!g138) & (!g128) & (!g146)) + ((ax104x) & (g127) & (!g138) & (!g128) & (g146)) + ((ax104x) & (g127) & (!g138) & (g128) & (!g146)) + ((ax104x) & (g127) & (!g138) & (g128) & (g146)) + ((ax104x) & (g127) & (g138) & (!g128) & (g146)));
	assign g164 = (((!ax100x) & (!ax101x)));
	assign g165 = (((!g127) & (!ax102x) & (!ax103x) & (!g128) & (!g146) & (!g164)) + ((!g127) & (!ax102x) & (!ax103x) & (g128) & (!g146) & (!g164)) + ((!g127) & (!ax102x) & (!ax103x) & (g128) & (g146) & (!g164)) + ((!g127) & (!ax102x) & (ax103x) & (!g128) & (g146) & (!g164)) + ((!g127) & (ax102x) & (ax103x) & (!g128) & (g146) & (!g164)) + ((!g127) & (ax102x) & (ax103x) & (!g128) & (g146) & (g164)) + ((g127) & (!ax102x) & (!ax103x) & (!g128) & (!g146) & (!g164)) + ((g127) & (!ax102x) & (!ax103x) & (!g128) & (!g146) & (g164)) + ((g127) & (!ax102x) & (!ax103x) & (!g128) & (g146) & (!g164)) + ((g127) & (!ax102x) & (!ax103x) & (g128) & (!g146) & (!g164)) + ((g127) & (!ax102x) & (!ax103x) & (g128) & (!g146) & (g164)) + ((g127) & (!ax102x) & (!ax103x) & (g128) & (g146) & (!g164)) + ((g127) & (!ax102x) & (!ax103x) & (g128) & (g146) & (g164)) + ((g127) & (!ax102x) & (ax103x) & (!g128) & (!g146) & (!g164)) + ((g127) & (!ax102x) & (ax103x) & (!g128) & (g146) & (!g164)) + ((g127) & (!ax102x) & (ax103x) & (!g128) & (g146) & (g164)) + ((g127) & (!ax102x) & (ax103x) & (g128) & (!g146) & (!g164)) + ((g127) & (!ax102x) & (ax103x) & (g128) & (g146) & (!g164)) + ((g127) & (ax102x) & (!ax103x) & (!g128) & (g146) & (!g164)) + ((g127) & (ax102x) & (!ax103x) & (!g128) & (g146) & (g164)) + ((g127) & (ax102x) & (ax103x) & (!g128) & (!g146) & (!g164)) + ((g127) & (ax102x) & (ax103x) & (!g128) & (!g146) & (g164)) + ((g127) & (ax102x) & (ax103x) & (!g128) & (g146) & (!g164)) + ((g127) & (ax102x) & (ax103x) & (!g128) & (g146) & (g164)) + ((g127) & (ax102x) & (ax103x) & (g128) & (!g146) & (!g164)) + ((g127) & (ax102x) & (ax103x) & (g128) & (!g146) & (g164)) + ((g127) & (ax102x) & (ax103x) & (g128) & (g146) & (!g164)) + ((g127) & (ax102x) & (ax103x) & (g128) & (g146) & (g164)));
	assign g166 = (((!g87) & (!g104) & (g162) & (g163) & (g165)) + ((!g87) & (g104) & (g162) & (!g163) & (g165)) + ((!g87) & (g104) & (g162) & (g163) & (!g165)) + ((!g87) & (g104) & (g162) & (g163) & (g165)) + ((g87) & (!g104) & (!g162) & (g163) & (g165)) + ((g87) & (!g104) & (g162) & (!g163) & (!g165)) + ((g87) & (!g104) & (g162) & (!g163) & (g165)) + ((g87) & (!g104) & (g162) & (g163) & (!g165)) + ((g87) & (!g104) & (g162) & (g163) & (g165)) + ((g87) & (g104) & (!g162) & (!g163) & (g165)) + ((g87) & (g104) & (!g162) & (g163) & (!g165)) + ((g87) & (g104) & (!g162) & (g163) & (g165)) + ((g87) & (g104) & (g162) & (!g163) & (!g165)) + ((g87) & (g104) & (g162) & (!g163) & (g165)) + ((g87) & (g104) & (g162) & (g163) & (!g165)) + ((g87) & (g104) & (g162) & (g163) & (g165)));
	assign g167 = (((!g54) & (!g68) & (g159) & (g160) & (g166)) + ((!g54) & (g68) & (g159) & (!g160) & (g166)) + ((!g54) & (g68) & (g159) & (g160) & (!g166)) + ((!g54) & (g68) & (g159) & (g160) & (g166)) + ((g54) & (!g68) & (!g159) & (g160) & (g166)) + ((g54) & (!g68) & (g159) & (!g160) & (!g166)) + ((g54) & (!g68) & (g159) & (!g160) & (g166)) + ((g54) & (!g68) & (g159) & (g160) & (!g166)) + ((g54) & (!g68) & (g159) & (g160) & (g166)) + ((g54) & (g68) & (!g159) & (!g160) & (g166)) + ((g54) & (g68) & (!g159) & (g160) & (!g166)) + ((g54) & (g68) & (!g159) & (g160) & (g166)) + ((g54) & (g68) & (g159) & (!g160) & (!g166)) + ((g54) & (g68) & (g159) & (!g160) & (g166)) + ((g54) & (g68) & (g159) & (g160) & (!g166)) + ((g54) & (g68) & (g159) & (g160) & (g166)));
	assign g168 = (((!g27) & (!g39) & (g156) & (g157) & (g167)) + ((!g27) & (g39) & (g156) & (!g157) & (g167)) + ((!g27) & (g39) & (g156) & (g157) & (!g167)) + ((!g27) & (g39) & (g156) & (g157) & (g167)) + ((g27) & (!g39) & (!g156) & (g157) & (g167)) + ((g27) & (!g39) & (g156) & (!g157) & (!g167)) + ((g27) & (!g39) & (g156) & (!g157) & (g167)) + ((g27) & (!g39) & (g156) & (g157) & (!g167)) + ((g27) & (!g39) & (g156) & (g157) & (g167)) + ((g27) & (g39) & (!g156) & (!g157) & (g167)) + ((g27) & (g39) & (!g156) & (g157) & (!g167)) + ((g27) & (g39) & (!g156) & (g157) & (g167)) + ((g27) & (g39) & (g156) & (!g157) & (!g167)) + ((g27) & (g39) & (g156) & (!g157) & (g167)) + ((g27) & (g39) & (g156) & (g157) & (!g167)) + ((g27) & (g39) & (g156) & (g157) & (g167)));
	assign g169 = (((!g8) & (!g18) & (g153) & (g154) & (g168)) + ((!g8) & (g18) & (g153) & (!g154) & (g168)) + ((!g8) & (g18) & (g153) & (g154) & (!g168)) + ((!g8) & (g18) & (g153) & (g154) & (g168)) + ((g8) & (!g18) & (!g153) & (g154) & (g168)) + ((g8) & (!g18) & (g153) & (!g154) & (!g168)) + ((g8) & (!g18) & (g153) & (!g154) & (g168)) + ((g8) & (!g18) & (g153) & (g154) & (!g168)) + ((g8) & (!g18) & (g153) & (g154) & (g168)) + ((g8) & (g18) & (!g153) & (!g154) & (g168)) + ((g8) & (g18) & (!g153) & (g154) & (!g168)) + ((g8) & (g18) & (!g153) & (g154) & (g168)) + ((g8) & (g18) & (g153) & (!g154) & (!g168)) + ((g8) & (g18) & (g153) & (!g154) & (g168)) + ((g8) & (g18) & (g153) & (g154) & (!g168)) + ((g8) & (g18) & (g153) & (g154) & (g168)));
	assign g170 = (((!g4) & (!g2) & (!g150) & (g151) & (g169)) + ((!g4) & (!g2) & (g150) & (!g151) & (!g169)) + ((!g4) & (!g2) & (g150) & (!g151) & (g169)) + ((!g4) & (!g2) & (g150) & (g151) & (!g169)) + ((!g4) & (!g2) & (g150) & (g151) & (g169)) + ((!g4) & (g2) & (!g150) & (!g151) & (g169)) + ((!g4) & (g2) & (!g150) & (g151) & (!g169)) + ((!g4) & (g2) & (!g150) & (g151) & (g169)) + ((!g4) & (g2) & (g150) & (!g151) & (!g169)) + ((!g4) & (g2) & (g150) & (!g151) & (g169)) + ((!g4) & (g2) & (g150) & (g151) & (!g169)) + ((!g4) & (g2) & (g150) & (g151) & (g169)) + ((g4) & (!g2) & (g150) & (g151) & (g169)) + ((g4) & (g2) & (g150) & (!g151) & (g169)) + ((g4) & (g2) & (g150) & (g151) & (!g169)) + ((g4) & (g2) & (g150) & (g151) & (g169)));
	assign g171 = (((!g4) & (!g143) & (g144)) + ((!g4) & (g143) & (!g144)) + ((!g4) & (g143) & (g144)) + ((g4) & (g143) & (g144)));
	assign g172 = (((!g129) & (!g171) & (!g128) & (!g146)) + ((!g129) & (!g171) & (g128) & (!g146)) + ((!g129) & (!g171) & (g128) & (g146)) + ((g129) & (g171) & (!g128) & (!g146)) + ((g129) & (g171) & (!g128) & (g146)) + ((g129) & (g171) & (g128) & (!g146)) + ((g129) & (g171) & (g128) & (g146)));
	assign g173 = (((!g1) & (g129) & (!g171) & (!g128) & (g146)) + ((!g1) & (g129) & (g171) & (!g128) & (g146)) + ((g1) & (!g129) & (g171) & (g128) & (!g146)) + ((g1) & (!g129) & (g171) & (g128) & (g146)) + ((g1) & (g129) & (!g171) & (!g128) & (!g146)) + ((g1) & (g129) & (!g171) & (!g128) & (g146)) + ((g1) & (g129) & (!g171) & (g128) & (!g146)) + ((g1) & (g129) & (!g171) & (g128) & (g146)) + ((g1) & (g129) & (g171) & (!g128) & (g146)));
	assign g174 = (((!g1) & (!g148) & (!g170) & (!g172) & (!g173)) + ((g1) & (!g148) & (!g170) & (!g172) & (!g173)) + ((g1) & (!g148) & (!g170) & (g172) & (!g173)) + ((g1) & (!g148) & (g170) & (!g172) & (!g173)) + ((g1) & (!g148) & (g170) & (g172) & (!g173)) + ((g1) & (g148) & (!g170) & (!g172) & (!g173)) + ((g1) & (g148) & (!g170) & (g172) & (!g173)));
	assign g175 = (((!g4) & (!g2) & (!g150) & (!g151) & (!g169) & (!g174)) + ((!g4) & (!g2) & (!g150) & (!g151) & (g169) & (!g174)) + ((!g4) & (!g2) & (!g150) & (g151) & (!g169) & (!g174)) + ((!g4) & (!g2) & (g150) & (!g151) & (!g169) & (g174)) + ((!g4) & (!g2) & (g150) & (!g151) & (g169) & (g174)) + ((!g4) & (!g2) & (g150) & (g151) & (!g169) & (g174)) + ((!g4) & (!g2) & (g150) & (g151) & (g169) & (!g174)) + ((!g4) & (!g2) & (g150) & (g151) & (g169) & (g174)) + ((!g4) & (g2) & (!g150) & (!g151) & (!g169) & (!g174)) + ((!g4) & (g2) & (g150) & (!g151) & (!g169) & (g174)) + ((!g4) & (g2) & (g150) & (!g151) & (g169) & (!g174)) + ((!g4) & (g2) & (g150) & (!g151) & (g169) & (g174)) + ((!g4) & (g2) & (g150) & (g151) & (!g169) & (!g174)) + ((!g4) & (g2) & (g150) & (g151) & (!g169) & (g174)) + ((!g4) & (g2) & (g150) & (g151) & (g169) & (!g174)) + ((!g4) & (g2) & (g150) & (g151) & (g169) & (g174)) + ((g4) & (!g2) & (!g150) & (g151) & (g169) & (!g174)) + ((g4) & (!g2) & (g150) & (!g151) & (!g169) & (!g174)) + ((g4) & (!g2) & (g150) & (!g151) & (!g169) & (g174)) + ((g4) & (!g2) & (g150) & (!g151) & (g169) & (!g174)) + ((g4) & (!g2) & (g150) & (!g151) & (g169) & (g174)) + ((g4) & (!g2) & (g150) & (g151) & (!g169) & (!g174)) + ((g4) & (!g2) & (g150) & (g151) & (!g169) & (g174)) + ((g4) & (!g2) & (g150) & (g151) & (g169) & (g174)) + ((g4) & (g2) & (!g150) & (!g151) & (g169) & (!g174)) + ((g4) & (g2) & (!g150) & (g151) & (!g169) & (!g174)) + ((g4) & (g2) & (!g150) & (g151) & (g169) & (!g174)) + ((g4) & (g2) & (g150) & (!g151) & (!g169) & (!g174)) + ((g4) & (g2) & (g150) & (!g151) & (!g169) & (g174)) + ((g4) & (g2) & (g150) & (!g151) & (g169) & (g174)) + ((g4) & (g2) & (g150) & (g151) & (!g169) & (g174)) + ((g4) & (g2) & (g150) & (g151) & (g169) & (g174)));
	assign g176 = (((!g8) & (!g18) & (!g153) & (g154) & (g168) & (!g174)) + ((!g8) & (!g18) & (g153) & (!g154) & (!g168) & (!g174)) + ((!g8) & (!g18) & (g153) & (!g154) & (!g168) & (g174)) + ((!g8) & (!g18) & (g153) & (!g154) & (g168) & (!g174)) + ((!g8) & (!g18) & (g153) & (!g154) & (g168) & (g174)) + ((!g8) & (!g18) & (g153) & (g154) & (!g168) & (!g174)) + ((!g8) & (!g18) & (g153) & (g154) & (!g168) & (g174)) + ((!g8) & (!g18) & (g153) & (g154) & (g168) & (g174)) + ((!g8) & (g18) & (!g153) & (!g154) & (g168) & (!g174)) + ((!g8) & (g18) & (!g153) & (g154) & (!g168) & (!g174)) + ((!g8) & (g18) & (!g153) & (g154) & (g168) & (!g174)) + ((!g8) & (g18) & (g153) & (!g154) & (!g168) & (!g174)) + ((!g8) & (g18) & (g153) & (!g154) & (!g168) & (g174)) + ((!g8) & (g18) & (g153) & (!g154) & (g168) & (g174)) + ((!g8) & (g18) & (g153) & (g154) & (!g168) & (g174)) + ((!g8) & (g18) & (g153) & (g154) & (g168) & (g174)) + ((g8) & (!g18) & (!g153) & (!g154) & (!g168) & (!g174)) + ((g8) & (!g18) & (!g153) & (!g154) & (g168) & (!g174)) + ((g8) & (!g18) & (!g153) & (g154) & (!g168) & (!g174)) + ((g8) & (!g18) & (g153) & (!g154) & (!g168) & (g174)) + ((g8) & (!g18) & (g153) & (!g154) & (g168) & (g174)) + ((g8) & (!g18) & (g153) & (g154) & (!g168) & (g174)) + ((g8) & (!g18) & (g153) & (g154) & (g168) & (!g174)) + ((g8) & (!g18) & (g153) & (g154) & (g168) & (g174)) + ((g8) & (g18) & (!g153) & (!g154) & (!g168) & (!g174)) + ((g8) & (g18) & (g153) & (!g154) & (!g168) & (g174)) + ((g8) & (g18) & (g153) & (!g154) & (g168) & (!g174)) + ((g8) & (g18) & (g153) & (!g154) & (g168) & (g174)) + ((g8) & (g18) & (g153) & (g154) & (!g168) & (!g174)) + ((g8) & (g18) & (g153) & (g154) & (!g168) & (g174)) + ((g8) & (g18) & (g153) & (g154) & (g168) & (!g174)) + ((g8) & (g18) & (g153) & (g154) & (g168) & (g174)));
	assign g177 = (((!g18) & (!g154) & (g168) & (!g174)) + ((!g18) & (g154) & (!g168) & (!g174)) + ((!g18) & (g154) & (!g168) & (g174)) + ((!g18) & (g154) & (g168) & (g174)) + ((g18) & (!g154) & (!g168) & (!g174)) + ((g18) & (g154) & (!g168) & (g174)) + ((g18) & (g154) & (g168) & (!g174)) + ((g18) & (g154) & (g168) & (g174)));
	assign g178 = (((!g27) & (!g39) & (!g156) & (g157) & (g167) & (!g174)) + ((!g27) & (!g39) & (g156) & (!g157) & (!g167) & (!g174)) + ((!g27) & (!g39) & (g156) & (!g157) & (!g167) & (g174)) + ((!g27) & (!g39) & (g156) & (!g157) & (g167) & (!g174)) + ((!g27) & (!g39) & (g156) & (!g157) & (g167) & (g174)) + ((!g27) & (!g39) & (g156) & (g157) & (!g167) & (!g174)) + ((!g27) & (!g39) & (g156) & (g157) & (!g167) & (g174)) + ((!g27) & (!g39) & (g156) & (g157) & (g167) & (g174)) + ((!g27) & (g39) & (!g156) & (!g157) & (g167) & (!g174)) + ((!g27) & (g39) & (!g156) & (g157) & (!g167) & (!g174)) + ((!g27) & (g39) & (!g156) & (g157) & (g167) & (!g174)) + ((!g27) & (g39) & (g156) & (!g157) & (!g167) & (!g174)) + ((!g27) & (g39) & (g156) & (!g157) & (!g167) & (g174)) + ((!g27) & (g39) & (g156) & (!g157) & (g167) & (g174)) + ((!g27) & (g39) & (g156) & (g157) & (!g167) & (g174)) + ((!g27) & (g39) & (g156) & (g157) & (g167) & (g174)) + ((g27) & (!g39) & (!g156) & (!g157) & (!g167) & (!g174)) + ((g27) & (!g39) & (!g156) & (!g157) & (g167) & (!g174)) + ((g27) & (!g39) & (!g156) & (g157) & (!g167) & (!g174)) + ((g27) & (!g39) & (g156) & (!g157) & (!g167) & (g174)) + ((g27) & (!g39) & (g156) & (!g157) & (g167) & (g174)) + ((g27) & (!g39) & (g156) & (g157) & (!g167) & (g174)) + ((g27) & (!g39) & (g156) & (g157) & (g167) & (!g174)) + ((g27) & (!g39) & (g156) & (g157) & (g167) & (g174)) + ((g27) & (g39) & (!g156) & (!g157) & (!g167) & (!g174)) + ((g27) & (g39) & (g156) & (!g157) & (!g167) & (g174)) + ((g27) & (g39) & (g156) & (!g157) & (g167) & (!g174)) + ((g27) & (g39) & (g156) & (!g157) & (g167) & (g174)) + ((g27) & (g39) & (g156) & (g157) & (!g167) & (!g174)) + ((g27) & (g39) & (g156) & (g157) & (!g167) & (g174)) + ((g27) & (g39) & (g156) & (g157) & (g167) & (!g174)) + ((g27) & (g39) & (g156) & (g157) & (g167) & (g174)));
	assign g179 = (((!g39) & (!g157) & (g167) & (!g174)) + ((!g39) & (g157) & (!g167) & (!g174)) + ((!g39) & (g157) & (!g167) & (g174)) + ((!g39) & (g157) & (g167) & (g174)) + ((g39) & (!g157) & (!g167) & (!g174)) + ((g39) & (g157) & (!g167) & (g174)) + ((g39) & (g157) & (g167) & (!g174)) + ((g39) & (g157) & (g167) & (g174)));
	assign g180 = (((!g54) & (!g68) & (!g159) & (g160) & (g166) & (!g174)) + ((!g54) & (!g68) & (g159) & (!g160) & (!g166) & (!g174)) + ((!g54) & (!g68) & (g159) & (!g160) & (!g166) & (g174)) + ((!g54) & (!g68) & (g159) & (!g160) & (g166) & (!g174)) + ((!g54) & (!g68) & (g159) & (!g160) & (g166) & (g174)) + ((!g54) & (!g68) & (g159) & (g160) & (!g166) & (!g174)) + ((!g54) & (!g68) & (g159) & (g160) & (!g166) & (g174)) + ((!g54) & (!g68) & (g159) & (g160) & (g166) & (g174)) + ((!g54) & (g68) & (!g159) & (!g160) & (g166) & (!g174)) + ((!g54) & (g68) & (!g159) & (g160) & (!g166) & (!g174)) + ((!g54) & (g68) & (!g159) & (g160) & (g166) & (!g174)) + ((!g54) & (g68) & (g159) & (!g160) & (!g166) & (!g174)) + ((!g54) & (g68) & (g159) & (!g160) & (!g166) & (g174)) + ((!g54) & (g68) & (g159) & (!g160) & (g166) & (g174)) + ((!g54) & (g68) & (g159) & (g160) & (!g166) & (g174)) + ((!g54) & (g68) & (g159) & (g160) & (g166) & (g174)) + ((g54) & (!g68) & (!g159) & (!g160) & (!g166) & (!g174)) + ((g54) & (!g68) & (!g159) & (!g160) & (g166) & (!g174)) + ((g54) & (!g68) & (!g159) & (g160) & (!g166) & (!g174)) + ((g54) & (!g68) & (g159) & (!g160) & (!g166) & (g174)) + ((g54) & (!g68) & (g159) & (!g160) & (g166) & (g174)) + ((g54) & (!g68) & (g159) & (g160) & (!g166) & (g174)) + ((g54) & (!g68) & (g159) & (g160) & (g166) & (!g174)) + ((g54) & (!g68) & (g159) & (g160) & (g166) & (g174)) + ((g54) & (g68) & (!g159) & (!g160) & (!g166) & (!g174)) + ((g54) & (g68) & (g159) & (!g160) & (!g166) & (g174)) + ((g54) & (g68) & (g159) & (!g160) & (g166) & (!g174)) + ((g54) & (g68) & (g159) & (!g160) & (g166) & (g174)) + ((g54) & (g68) & (g159) & (g160) & (!g166) & (!g174)) + ((g54) & (g68) & (g159) & (g160) & (!g166) & (g174)) + ((g54) & (g68) & (g159) & (g160) & (g166) & (!g174)) + ((g54) & (g68) & (g159) & (g160) & (g166) & (g174)));
	assign g181 = (((!g68) & (!g160) & (g166) & (!g174)) + ((!g68) & (g160) & (!g166) & (!g174)) + ((!g68) & (g160) & (!g166) & (g174)) + ((!g68) & (g160) & (g166) & (g174)) + ((g68) & (!g160) & (!g166) & (!g174)) + ((g68) & (g160) & (!g166) & (g174)) + ((g68) & (g160) & (g166) & (!g174)) + ((g68) & (g160) & (g166) & (g174)));
	assign g182 = (((!g87) & (!g104) & (!g162) & (g163) & (g165) & (!g174)) + ((!g87) & (!g104) & (g162) & (!g163) & (!g165) & (!g174)) + ((!g87) & (!g104) & (g162) & (!g163) & (!g165) & (g174)) + ((!g87) & (!g104) & (g162) & (!g163) & (g165) & (!g174)) + ((!g87) & (!g104) & (g162) & (!g163) & (g165) & (g174)) + ((!g87) & (!g104) & (g162) & (g163) & (!g165) & (!g174)) + ((!g87) & (!g104) & (g162) & (g163) & (!g165) & (g174)) + ((!g87) & (!g104) & (g162) & (g163) & (g165) & (g174)) + ((!g87) & (g104) & (!g162) & (!g163) & (g165) & (!g174)) + ((!g87) & (g104) & (!g162) & (g163) & (!g165) & (!g174)) + ((!g87) & (g104) & (!g162) & (g163) & (g165) & (!g174)) + ((!g87) & (g104) & (g162) & (!g163) & (!g165) & (!g174)) + ((!g87) & (g104) & (g162) & (!g163) & (!g165) & (g174)) + ((!g87) & (g104) & (g162) & (!g163) & (g165) & (g174)) + ((!g87) & (g104) & (g162) & (g163) & (!g165) & (g174)) + ((!g87) & (g104) & (g162) & (g163) & (g165) & (g174)) + ((g87) & (!g104) & (!g162) & (!g163) & (!g165) & (!g174)) + ((g87) & (!g104) & (!g162) & (!g163) & (g165) & (!g174)) + ((g87) & (!g104) & (!g162) & (g163) & (!g165) & (!g174)) + ((g87) & (!g104) & (g162) & (!g163) & (!g165) & (g174)) + ((g87) & (!g104) & (g162) & (!g163) & (g165) & (g174)) + ((g87) & (!g104) & (g162) & (g163) & (!g165) & (g174)) + ((g87) & (!g104) & (g162) & (g163) & (g165) & (!g174)) + ((g87) & (!g104) & (g162) & (g163) & (g165) & (g174)) + ((g87) & (g104) & (!g162) & (!g163) & (!g165) & (!g174)) + ((g87) & (g104) & (g162) & (!g163) & (!g165) & (g174)) + ((g87) & (g104) & (g162) & (!g163) & (g165) & (!g174)) + ((g87) & (g104) & (g162) & (!g163) & (g165) & (g174)) + ((g87) & (g104) & (g162) & (g163) & (!g165) & (!g174)) + ((g87) & (g104) & (g162) & (g163) & (!g165) & (g174)) + ((g87) & (g104) & (g162) & (g163) & (g165) & (!g174)) + ((g87) & (g104) & (g162) & (g163) & (g165) & (g174)));
	assign g183 = (((!g104) & (!g163) & (g165) & (!g174)) + ((!g104) & (g163) & (!g165) & (!g174)) + ((!g104) & (g163) & (!g165) & (g174)) + ((!g104) & (g163) & (g165) & (g174)) + ((g104) & (!g163) & (!g165) & (!g174)) + ((g104) & (g163) & (!g165) & (g174)) + ((g104) & (g163) & (g165) & (!g174)) + ((g104) & (g163) & (g165) & (g174)));
	assign g184 = (((!g127) & (!ax102x) & (!ax103x) & (!g147) & (!g164) & (g174)) + ((!g127) & (!ax102x) & (!ax103x) & (!g147) & (g164) & (!g174)) + ((!g127) & (!ax102x) & (!ax103x) & (!g147) & (g164) & (g174)) + ((!g127) & (!ax102x) & (!ax103x) & (g147) & (!g164) & (!g174)) + ((!g127) & (!ax102x) & (ax103x) & (!g147) & (!g164) & (!g174)) + ((!g127) & (!ax102x) & (ax103x) & (g147) & (!g164) & (g174)) + ((!g127) & (!ax102x) & (ax103x) & (g147) & (g164) & (!g174)) + ((!g127) & (!ax102x) & (ax103x) & (g147) & (g164) & (g174)) + ((!g127) & (ax102x) & (!ax103x) & (g147) & (!g164) & (!g174)) + ((!g127) & (ax102x) & (!ax103x) & (g147) & (g164) & (!g174)) + ((!g127) & (ax102x) & (ax103x) & (!g147) & (!g164) & (!g174)) + ((!g127) & (ax102x) & (ax103x) & (!g147) & (!g164) & (g174)) + ((!g127) & (ax102x) & (ax103x) & (!g147) & (g164) & (!g174)) + ((!g127) & (ax102x) & (ax103x) & (!g147) & (g164) & (g174)) + ((!g127) & (ax102x) & (ax103x) & (g147) & (!g164) & (g174)) + ((!g127) & (ax102x) & (ax103x) & (g147) & (g164) & (g174)) + ((g127) & (!ax102x) & (!ax103x) & (!g147) & (!g164) & (!g174)) + ((g127) & (!ax102x) & (!ax103x) & (!g147) & (!g164) & (g174)) + ((g127) & (!ax102x) & (!ax103x) & (!g147) & (g164) & (g174)) + ((g127) & (!ax102x) & (!ax103x) & (g147) & (g164) & (!g174)) + ((g127) & (!ax102x) & (ax103x) & (!g147) & (g164) & (!g174)) + ((g127) & (!ax102x) & (ax103x) & (g147) & (!g164) & (!g174)) + ((g127) & (!ax102x) & (ax103x) & (g147) & (!g164) & (g174)) + ((g127) & (!ax102x) & (ax103x) & (g147) & (g164) & (g174)) + ((g127) & (ax102x) & (!ax103x) & (!g147) & (!g164) & (!g174)) + ((g127) & (ax102x) & (!ax103x) & (!g147) & (g164) & (!g174)) + ((g127) & (ax102x) & (ax103x) & (!g147) & (!g164) & (g174)) + ((g127) & (ax102x) & (ax103x) & (!g147) & (g164) & (g174)) + ((g127) & (ax102x) & (ax103x) & (g147) & (!g164) & (!g174)) + ((g127) & (ax102x) & (ax103x) & (g147) & (!g164) & (g174)) + ((g127) & (ax102x) & (ax103x) & (g147) & (g164) & (!g174)) + ((g127) & (ax102x) & (ax103x) & (g147) & (g164) & (g174)));
	assign g185 = (((!ax102x) & (!g147) & (!g164) & (g174)) + ((!ax102x) & (!g147) & (g164) & (!g174)) + ((!ax102x) & (!g147) & (g164) & (g174)) + ((!ax102x) & (g147) & (g164) & (!g174)) + ((ax102x) & (!g147) & (!g164) & (!g174)) + ((ax102x) & (g147) & (!g164) & (!g174)) + ((ax102x) & (g147) & (!g164) & (g174)) + ((ax102x) & (g147) & (g164) & (g174)));
	assign g186 = (((!ax98x) & (!ax99x)));
	assign g187 = (((!g147) & (!ax100x) & (!ax101x) & (!g174) & (!g186)) + ((!g147) & (!ax100x) & (ax101x) & (g174) & (!g186)) + ((!g147) & (ax100x) & (ax101x) & (g174) & (!g186)) + ((!g147) & (ax100x) & (ax101x) & (g174) & (g186)) + ((g147) & (!ax100x) & (!ax101x) & (!g174) & (!g186)) + ((g147) & (!ax100x) & (!ax101x) & (!g174) & (g186)) + ((g147) & (!ax100x) & (!ax101x) & (g174) & (!g186)) + ((g147) & (!ax100x) & (ax101x) & (!g174) & (!g186)) + ((g147) & (!ax100x) & (ax101x) & (g174) & (!g186)) + ((g147) & (!ax100x) & (ax101x) & (g174) & (g186)) + ((g147) & (ax100x) & (!ax101x) & (g174) & (!g186)) + ((g147) & (ax100x) & (!ax101x) & (g174) & (g186)) + ((g147) & (ax100x) & (ax101x) & (!g174) & (!g186)) + ((g147) & (ax100x) & (ax101x) & (!g174) & (g186)) + ((g147) & (ax100x) & (ax101x) & (g174) & (!g186)) + ((g147) & (ax100x) & (ax101x) & (g174) & (g186)));
	assign g188 = (((!g104) & (!g127) & (g184) & (g185) & (g187)) + ((!g104) & (g127) & (g184) & (!g185) & (g187)) + ((!g104) & (g127) & (g184) & (g185) & (!g187)) + ((!g104) & (g127) & (g184) & (g185) & (g187)) + ((g104) & (!g127) & (!g184) & (g185) & (g187)) + ((g104) & (!g127) & (g184) & (!g185) & (!g187)) + ((g104) & (!g127) & (g184) & (!g185) & (g187)) + ((g104) & (!g127) & (g184) & (g185) & (!g187)) + ((g104) & (!g127) & (g184) & (g185) & (g187)) + ((g104) & (g127) & (!g184) & (!g185) & (g187)) + ((g104) & (g127) & (!g184) & (g185) & (!g187)) + ((g104) & (g127) & (!g184) & (g185) & (g187)) + ((g104) & (g127) & (g184) & (!g185) & (!g187)) + ((g104) & (g127) & (g184) & (!g185) & (g187)) + ((g104) & (g127) & (g184) & (g185) & (!g187)) + ((g104) & (g127) & (g184) & (g185) & (g187)));
	assign g189 = (((!g68) & (!g87) & (g182) & (g183) & (g188)) + ((!g68) & (g87) & (g182) & (!g183) & (g188)) + ((!g68) & (g87) & (g182) & (g183) & (!g188)) + ((!g68) & (g87) & (g182) & (g183) & (g188)) + ((g68) & (!g87) & (!g182) & (g183) & (g188)) + ((g68) & (!g87) & (g182) & (!g183) & (!g188)) + ((g68) & (!g87) & (g182) & (!g183) & (g188)) + ((g68) & (!g87) & (g182) & (g183) & (!g188)) + ((g68) & (!g87) & (g182) & (g183) & (g188)) + ((g68) & (g87) & (!g182) & (!g183) & (g188)) + ((g68) & (g87) & (!g182) & (g183) & (!g188)) + ((g68) & (g87) & (!g182) & (g183) & (g188)) + ((g68) & (g87) & (g182) & (!g183) & (!g188)) + ((g68) & (g87) & (g182) & (!g183) & (g188)) + ((g68) & (g87) & (g182) & (g183) & (!g188)) + ((g68) & (g87) & (g182) & (g183) & (g188)));
	assign g190 = (((!g39) & (!g54) & (g180) & (g181) & (g189)) + ((!g39) & (g54) & (g180) & (!g181) & (g189)) + ((!g39) & (g54) & (g180) & (g181) & (!g189)) + ((!g39) & (g54) & (g180) & (g181) & (g189)) + ((g39) & (!g54) & (!g180) & (g181) & (g189)) + ((g39) & (!g54) & (g180) & (!g181) & (!g189)) + ((g39) & (!g54) & (g180) & (!g181) & (g189)) + ((g39) & (!g54) & (g180) & (g181) & (!g189)) + ((g39) & (!g54) & (g180) & (g181) & (g189)) + ((g39) & (g54) & (!g180) & (!g181) & (g189)) + ((g39) & (g54) & (!g180) & (g181) & (!g189)) + ((g39) & (g54) & (!g180) & (g181) & (g189)) + ((g39) & (g54) & (g180) & (!g181) & (!g189)) + ((g39) & (g54) & (g180) & (!g181) & (g189)) + ((g39) & (g54) & (g180) & (g181) & (!g189)) + ((g39) & (g54) & (g180) & (g181) & (g189)));
	assign g191 = (((!g18) & (!g27) & (g178) & (g179) & (g190)) + ((!g18) & (g27) & (g178) & (!g179) & (g190)) + ((!g18) & (g27) & (g178) & (g179) & (!g190)) + ((!g18) & (g27) & (g178) & (g179) & (g190)) + ((g18) & (!g27) & (!g178) & (g179) & (g190)) + ((g18) & (!g27) & (g178) & (!g179) & (!g190)) + ((g18) & (!g27) & (g178) & (!g179) & (g190)) + ((g18) & (!g27) & (g178) & (g179) & (!g190)) + ((g18) & (!g27) & (g178) & (g179) & (g190)) + ((g18) & (g27) & (!g178) & (!g179) & (g190)) + ((g18) & (g27) & (!g178) & (g179) & (!g190)) + ((g18) & (g27) & (!g178) & (g179) & (g190)) + ((g18) & (g27) & (g178) & (!g179) & (!g190)) + ((g18) & (g27) & (g178) & (!g179) & (g190)) + ((g18) & (g27) & (g178) & (g179) & (!g190)) + ((g18) & (g27) & (g178) & (g179) & (g190)));
	assign g192 = (((!g2) & (!g8) & (g176) & (g177) & (g191)) + ((!g2) & (g8) & (g176) & (!g177) & (g191)) + ((!g2) & (g8) & (g176) & (g177) & (!g191)) + ((!g2) & (g8) & (g176) & (g177) & (g191)) + ((g2) & (!g8) & (!g176) & (g177) & (g191)) + ((g2) & (!g8) & (g176) & (!g177) & (!g191)) + ((g2) & (!g8) & (g176) & (!g177) & (g191)) + ((g2) & (!g8) & (g176) & (g177) & (!g191)) + ((g2) & (!g8) & (g176) & (g177) & (g191)) + ((g2) & (g8) & (!g176) & (!g177) & (g191)) + ((g2) & (g8) & (!g176) & (g177) & (!g191)) + ((g2) & (g8) & (!g176) & (g177) & (g191)) + ((g2) & (g8) & (g176) & (!g177) & (!g191)) + ((g2) & (g8) & (g176) & (!g177) & (g191)) + ((g2) & (g8) & (g176) & (g177) & (!g191)) + ((g2) & (g8) & (g176) & (g177) & (g191)));
	assign g193 = (((!g2) & (!g151) & (g169) & (!g174)) + ((!g2) & (g151) & (!g169) & (!g174)) + ((!g2) & (g151) & (!g169) & (g174)) + ((!g2) & (g151) & (g169) & (g174)) + ((g2) & (!g151) & (!g169) & (!g174)) + ((g2) & (g151) & (!g169) & (g174)) + ((g2) & (g151) & (g169) & (!g174)) + ((g2) & (g151) & (g169) & (g174)));
	assign g194 = (((!g1) & (!g148) & (!g170) & (!g172) & (g173)) + ((!g1) & (!g148) & (!g170) & (g172) & (!g173)) + ((!g1) & (!g148) & (!g170) & (g172) & (g173)) + ((!g1) & (g148) & (g170) & (!g172) & (!g173)) + ((!g1) & (g148) & (g170) & (!g172) & (g173)) + ((!g1) & (g148) & (g170) & (g172) & (!g173)) + ((!g1) & (g148) & (g170) & (g172) & (g173)) + ((g1) & (!g148) & (!g170) & (!g172) & (g173)) + ((g1) & (!g148) & (!g170) & (g172) & (g173)) + ((g1) & (g148) & (g170) & (!g172) & (!g173)) + ((g1) & (g148) & (g170) & (!g172) & (g173)) + ((g1) & (g148) & (g170) & (g172) & (!g173)) + ((g1) & (g148) & (g170) & (g172) & (g173)));
	assign g195 = (((!g4) & (!g1) & (!g175) & (!g192) & (!g193) & (g194)) + ((!g4) & (!g1) & (!g175) & (!g192) & (g193) & (!g194)) + ((!g4) & (!g1) & (!g175) & (!g192) & (g193) & (g194)) + ((!g4) & (!g1) & (!g175) & (g192) & (!g193) & (!g194)) + ((!g4) & (!g1) & (!g175) & (g192) & (!g193) & (g194)) + ((!g4) & (!g1) & (!g175) & (g192) & (g193) & (!g194)) + ((!g4) & (!g1) & (!g175) & (g192) & (g193) & (g194)) + ((!g4) & (!g1) & (g175) & (!g192) & (!g193) & (!g194)) + ((!g4) & (!g1) & (g175) & (!g192) & (!g193) & (g194)) + ((!g4) & (!g1) & (g175) & (!g192) & (g193) & (!g194)) + ((!g4) & (!g1) & (g175) & (!g192) & (g193) & (g194)) + ((!g4) & (!g1) & (g175) & (g192) & (!g193) & (!g194)) + ((!g4) & (!g1) & (g175) & (g192) & (!g193) & (g194)) + ((!g4) & (!g1) & (g175) & (g192) & (g193) & (!g194)) + ((!g4) & (!g1) & (g175) & (g192) & (g193) & (g194)) + ((g4) & (!g1) & (!g175) & (!g192) & (!g193) & (g194)) + ((g4) & (!g1) & (!g175) & (!g192) & (g193) & (g194)) + ((g4) & (!g1) & (!g175) & (g192) & (!g193) & (g194)) + ((g4) & (!g1) & (!g175) & (g192) & (g193) & (!g194)) + ((g4) & (!g1) & (!g175) & (g192) & (g193) & (g194)) + ((g4) & (!g1) & (g175) & (!g192) & (!g193) & (!g194)) + ((g4) & (!g1) & (g175) & (!g192) & (!g193) & (g194)) + ((g4) & (!g1) & (g175) & (!g192) & (g193) & (!g194)) + ((g4) & (!g1) & (g175) & (!g192) & (g193) & (g194)) + ((g4) & (!g1) & (g175) & (g192) & (!g193) & (!g194)) + ((g4) & (!g1) & (g175) & (g192) & (!g193) & (g194)) + ((g4) & (!g1) & (g175) & (g192) & (g193) & (!g194)) + ((g4) & (!g1) & (g175) & (g192) & (g193) & (g194)));
	assign g196 = (((g1) & (!g148) & (g170) & (g173)) + ((g1) & (g148) & (!g170) & (!g173)) + ((g1) & (g148) & (!g170) & (g173)));
	assign g197 = (((!g4) & (!g175) & (!g192) & (!g193) & (!g196)) + ((!g4) & (!g175) & (!g192) & (g193) & (!g196)) + ((!g4) & (!g175) & (g192) & (!g193) & (!g196)) + ((!g4) & (!g175) & (g192) & (g193) & (!g196)) + ((!g4) & (g175) & (!g192) & (!g193) & (!g196)) + ((g4) & (!g175) & (!g192) & (!g193) & (!g196)) + ((g4) & (!g175) & (!g192) & (g193) & (!g196)) + ((g4) & (!g175) & (g192) & (!g193) & (!g196)) + ((g4) & (!g175) & (g192) & (g193) & (!g196)) + ((g4) & (g175) & (!g192) & (!g193) & (!g196)) + ((g4) & (g175) & (!g192) & (g193) & (!g196)) + ((g4) & (g175) & (g192) & (!g193) & (!g196)));
	assign g198 = (((!g195) & (g197)));
	assign g199 = (((!g4) & (!g192) & (!g193) & (!g195) & (!g197)) + ((!g4) & (!g192) & (!g193) & (g195) & (!g197)) + ((!g4) & (!g192) & (!g193) & (g195) & (g197)) + ((!g4) & (!g192) & (g193) & (!g195) & (g197)) + ((!g4) & (g192) & (g193) & (!g195) & (!g197)) + ((!g4) & (g192) & (g193) & (!g195) & (g197)) + ((!g4) & (g192) & (g193) & (g195) & (!g197)) + ((!g4) & (g192) & (g193) & (g195) & (g197)) + ((g4) & (!g192) & (g193) & (!g195) & (!g197)) + ((g4) & (!g192) & (g193) & (!g195) & (g197)) + ((g4) & (!g192) & (g193) & (g195) & (!g197)) + ((g4) & (!g192) & (g193) & (g195) & (g197)) + ((g4) & (g192) & (!g193) & (!g195) & (!g197)) + ((g4) & (g192) & (!g193) & (g195) & (!g197)) + ((g4) & (g192) & (!g193) & (g195) & (g197)) + ((g4) & (g192) & (g193) & (!g195) & (g197)));
	assign g200 = (((!g8) & (!g177) & (g191) & (!g195) & (!g197)) + ((!g8) & (!g177) & (g191) & (g195) & (!g197)) + ((!g8) & (!g177) & (g191) & (g195) & (g197)) + ((!g8) & (g177) & (!g191) & (!g195) & (!g197)) + ((!g8) & (g177) & (!g191) & (!g195) & (g197)) + ((!g8) & (g177) & (!g191) & (g195) & (!g197)) + ((!g8) & (g177) & (!g191) & (g195) & (g197)) + ((!g8) & (g177) & (g191) & (!g195) & (g197)) + ((g8) & (!g177) & (!g191) & (!g195) & (!g197)) + ((g8) & (!g177) & (!g191) & (g195) & (!g197)) + ((g8) & (!g177) & (!g191) & (g195) & (g197)) + ((g8) & (g177) & (!g191) & (!g195) & (g197)) + ((g8) & (g177) & (g191) & (!g195) & (!g197)) + ((g8) & (g177) & (g191) & (!g195) & (g197)) + ((g8) & (g177) & (g191) & (g195) & (!g197)) + ((g8) & (g177) & (g191) & (g195) & (g197)));
	assign g201 = (((!g18) & (!g27) & (g179) & (g190)) + ((!g18) & (g27) & (!g179) & (g190)) + ((!g18) & (g27) & (g179) & (!g190)) + ((!g18) & (g27) & (g179) & (g190)) + ((g18) & (!g27) & (!g179) & (!g190)) + ((g18) & (!g27) & (!g179) & (g190)) + ((g18) & (!g27) & (g179) & (!g190)) + ((g18) & (g27) & (!g179) & (!g190)));
	assign g202 = (((!g178) & (!g195) & (!g197) & (g201)) + ((!g178) & (g195) & (!g197) & (g201)) + ((!g178) & (g195) & (g197) & (g201)) + ((g178) & (!g195) & (!g197) & (!g201)) + ((g178) & (!g195) & (g197) & (!g201)) + ((g178) & (!g195) & (g197) & (g201)) + ((g178) & (g195) & (!g197) & (!g201)) + ((g178) & (g195) & (g197) & (!g201)));
	assign g203 = (((!g27) & (!g179) & (g190) & (!g195) & (!g197)) + ((!g27) & (!g179) & (g190) & (g195) & (!g197)) + ((!g27) & (!g179) & (g190) & (g195) & (g197)) + ((!g27) & (g179) & (!g190) & (!g195) & (!g197)) + ((!g27) & (g179) & (!g190) & (!g195) & (g197)) + ((!g27) & (g179) & (!g190) & (g195) & (!g197)) + ((!g27) & (g179) & (!g190) & (g195) & (g197)) + ((!g27) & (g179) & (g190) & (!g195) & (g197)) + ((g27) & (!g179) & (!g190) & (!g195) & (!g197)) + ((g27) & (!g179) & (!g190) & (g195) & (!g197)) + ((g27) & (!g179) & (!g190) & (g195) & (g197)) + ((g27) & (g179) & (!g190) & (!g195) & (g197)) + ((g27) & (g179) & (g190) & (!g195) & (!g197)) + ((g27) & (g179) & (g190) & (!g195) & (g197)) + ((g27) & (g179) & (g190) & (g195) & (!g197)) + ((g27) & (g179) & (g190) & (g195) & (g197)));
	assign g204 = (((!g39) & (!g54) & (g181) & (g189)) + ((!g39) & (g54) & (!g181) & (g189)) + ((!g39) & (g54) & (g181) & (!g189)) + ((!g39) & (g54) & (g181) & (g189)) + ((g39) & (!g54) & (!g181) & (!g189)) + ((g39) & (!g54) & (!g181) & (g189)) + ((g39) & (!g54) & (g181) & (!g189)) + ((g39) & (g54) & (!g181) & (!g189)));
	assign g205 = (((!g180) & (!g195) & (!g197) & (g204)) + ((!g180) & (g195) & (!g197) & (g204)) + ((!g180) & (g195) & (g197) & (g204)) + ((g180) & (!g195) & (!g197) & (!g204)) + ((g180) & (!g195) & (g197) & (!g204)) + ((g180) & (!g195) & (g197) & (g204)) + ((g180) & (g195) & (!g197) & (!g204)) + ((g180) & (g195) & (g197) & (!g204)));
	assign g206 = (((!g54) & (!g181) & (g189) & (!g195) & (!g197)) + ((!g54) & (!g181) & (g189) & (g195) & (!g197)) + ((!g54) & (!g181) & (g189) & (g195) & (g197)) + ((!g54) & (g181) & (!g189) & (!g195) & (!g197)) + ((!g54) & (g181) & (!g189) & (!g195) & (g197)) + ((!g54) & (g181) & (!g189) & (g195) & (!g197)) + ((!g54) & (g181) & (!g189) & (g195) & (g197)) + ((!g54) & (g181) & (g189) & (!g195) & (g197)) + ((g54) & (!g181) & (!g189) & (!g195) & (!g197)) + ((g54) & (!g181) & (!g189) & (g195) & (!g197)) + ((g54) & (!g181) & (!g189) & (g195) & (g197)) + ((g54) & (g181) & (!g189) & (!g195) & (g197)) + ((g54) & (g181) & (g189) & (!g195) & (!g197)) + ((g54) & (g181) & (g189) & (!g195) & (g197)) + ((g54) & (g181) & (g189) & (g195) & (!g197)) + ((g54) & (g181) & (g189) & (g195) & (g197)));
	assign g207 = (((!g68) & (!g87) & (g183) & (g188)) + ((!g68) & (g87) & (!g183) & (g188)) + ((!g68) & (g87) & (g183) & (!g188)) + ((!g68) & (g87) & (g183) & (g188)) + ((g68) & (!g87) & (!g183) & (!g188)) + ((g68) & (!g87) & (!g183) & (g188)) + ((g68) & (!g87) & (g183) & (!g188)) + ((g68) & (g87) & (!g183) & (!g188)));
	assign g208 = (((!g182) & (!g195) & (!g197) & (g207)) + ((!g182) & (g195) & (!g197) & (g207)) + ((!g182) & (g195) & (g197) & (g207)) + ((g182) & (!g195) & (!g197) & (!g207)) + ((g182) & (!g195) & (g197) & (!g207)) + ((g182) & (!g195) & (g197) & (g207)) + ((g182) & (g195) & (!g197) & (!g207)) + ((g182) & (g195) & (g197) & (!g207)));
	assign g209 = (((!g87) & (!g183) & (g188) & (!g195) & (!g197)) + ((!g87) & (!g183) & (g188) & (g195) & (!g197)) + ((!g87) & (!g183) & (g188) & (g195) & (g197)) + ((!g87) & (g183) & (!g188) & (!g195) & (!g197)) + ((!g87) & (g183) & (!g188) & (!g195) & (g197)) + ((!g87) & (g183) & (!g188) & (g195) & (!g197)) + ((!g87) & (g183) & (!g188) & (g195) & (g197)) + ((!g87) & (g183) & (g188) & (!g195) & (g197)) + ((g87) & (!g183) & (!g188) & (!g195) & (!g197)) + ((g87) & (!g183) & (!g188) & (g195) & (!g197)) + ((g87) & (!g183) & (!g188) & (g195) & (g197)) + ((g87) & (g183) & (!g188) & (!g195) & (g197)) + ((g87) & (g183) & (g188) & (!g195) & (!g197)) + ((g87) & (g183) & (g188) & (!g195) & (g197)) + ((g87) & (g183) & (g188) & (g195) & (!g197)) + ((g87) & (g183) & (g188) & (g195) & (g197)));
	assign g210 = (((!g104) & (!g127) & (g185) & (g187)) + ((!g104) & (g127) & (!g185) & (g187)) + ((!g104) & (g127) & (g185) & (!g187)) + ((!g104) & (g127) & (g185) & (g187)) + ((g104) & (!g127) & (!g185) & (!g187)) + ((g104) & (!g127) & (!g185) & (g187)) + ((g104) & (!g127) & (g185) & (!g187)) + ((g104) & (g127) & (!g185) & (!g187)));
	assign g211 = (((!g184) & (!g195) & (!g197) & (g210)) + ((!g184) & (g195) & (!g197) & (g210)) + ((!g184) & (g195) & (g197) & (g210)) + ((g184) & (!g195) & (!g197) & (!g210)) + ((g184) & (!g195) & (g197) & (!g210)) + ((g184) & (!g195) & (g197) & (g210)) + ((g184) & (g195) & (!g197) & (!g210)) + ((g184) & (g195) & (g197) & (!g210)));
	assign g212 = (((!g127) & (!g185) & (g187) & (!g195) & (!g197)) + ((!g127) & (!g185) & (g187) & (g195) & (!g197)) + ((!g127) & (!g185) & (g187) & (g195) & (g197)) + ((!g127) & (g185) & (!g187) & (!g195) & (!g197)) + ((!g127) & (g185) & (!g187) & (!g195) & (g197)) + ((!g127) & (g185) & (!g187) & (g195) & (!g197)) + ((!g127) & (g185) & (!g187) & (g195) & (g197)) + ((!g127) & (g185) & (g187) & (!g195) & (g197)) + ((g127) & (!g185) & (!g187) & (!g195) & (!g197)) + ((g127) & (!g185) & (!g187) & (g195) & (!g197)) + ((g127) & (!g185) & (!g187) & (g195) & (g197)) + ((g127) & (g185) & (!g187) & (!g195) & (g197)) + ((g127) & (g185) & (g187) & (!g195) & (!g197)) + ((g127) & (g185) & (g187) & (!g195) & (g197)) + ((g127) & (g185) & (g187) & (g195) & (!g197)) + ((g127) & (g185) & (g187) & (g195) & (g197)));
	assign g213 = (((!g147) & (!ax100x) & (!g174) & (g186)) + ((!g147) & (!ax100x) & (g174) & (g186)) + ((!g147) & (ax100x) & (!g174) & (!g186)) + ((!g147) & (ax100x) & (!g174) & (g186)) + ((g147) & (!ax100x) & (!g174) & (!g186)) + ((g147) & (!ax100x) & (g174) & (!g186)) + ((g147) & (ax100x) & (g174) & (!g186)) + ((g147) & (ax100x) & (g174) & (g186)));
	assign g214 = (((!ax100x) & (!ax101x) & (!g174) & (!g195) & (!g197) & (g213)) + ((!ax100x) & (!ax101x) & (!g174) & (!g195) & (g197) & (!g213)) + ((!ax100x) & (!ax101x) & (!g174) & (!g195) & (g197) & (g213)) + ((!ax100x) & (!ax101x) & (!g174) & (g195) & (!g197) & (g213)) + ((!ax100x) & (!ax101x) & (!g174) & (g195) & (g197) & (g213)) + ((!ax100x) & (!ax101x) & (g174) & (!g195) & (!g197) & (!g213)) + ((!ax100x) & (!ax101x) & (g174) & (g195) & (!g197) & (!g213)) + ((!ax100x) & (!ax101x) & (g174) & (g195) & (g197) & (!g213)) + ((!ax100x) & (ax101x) & (!g174) & (!g195) & (!g197) & (!g213)) + ((!ax100x) & (ax101x) & (!g174) & (g195) & (!g197) & (!g213)) + ((!ax100x) & (ax101x) & (!g174) & (g195) & (g197) & (!g213)) + ((!ax100x) & (ax101x) & (g174) & (!g195) & (!g197) & (g213)) + ((!ax100x) & (ax101x) & (g174) & (!g195) & (g197) & (!g213)) + ((!ax100x) & (ax101x) & (g174) & (!g195) & (g197) & (g213)) + ((!ax100x) & (ax101x) & (g174) & (g195) & (!g197) & (g213)) + ((!ax100x) & (ax101x) & (g174) & (g195) & (g197) & (g213)) + ((ax100x) & (!ax101x) & (!g174) & (!g195) & (!g197) & (!g213)) + ((ax100x) & (!ax101x) & (!g174) & (g195) & (!g197) & (!g213)) + ((ax100x) & (!ax101x) & (!g174) & (g195) & (g197) & (!g213)) + ((ax100x) & (!ax101x) & (g174) & (!g195) & (!g197) & (!g213)) + ((ax100x) & (!ax101x) & (g174) & (g195) & (!g197) & (!g213)) + ((ax100x) & (!ax101x) & (g174) & (g195) & (g197) & (!g213)) + ((ax100x) & (ax101x) & (!g174) & (!g195) & (!g197) & (g213)) + ((ax100x) & (ax101x) & (!g174) & (!g195) & (g197) & (!g213)) + ((ax100x) & (ax101x) & (!g174) & (!g195) & (g197) & (g213)) + ((ax100x) & (ax101x) & (!g174) & (g195) & (!g197) & (g213)) + ((ax100x) & (ax101x) & (!g174) & (g195) & (g197) & (g213)) + ((ax100x) & (ax101x) & (g174) & (!g195) & (!g197) & (g213)) + ((ax100x) & (ax101x) & (g174) & (!g195) & (g197) & (!g213)) + ((ax100x) & (ax101x) & (g174) & (!g195) & (g197) & (g213)) + ((ax100x) & (ax101x) & (g174) & (g195) & (!g197) & (g213)) + ((ax100x) & (ax101x) & (g174) & (g195) & (g197) & (g213)));
	assign g215 = (((!ax100x) & (!g174) & (!g186) & (!g195) & (g197)) + ((!ax100x) & (!g174) & (g186) & (!g195) & (!g197)) + ((!ax100x) & (!g174) & (g186) & (!g195) & (g197)) + ((!ax100x) & (!g174) & (g186) & (g195) & (!g197)) + ((!ax100x) & (!g174) & (g186) & (g195) & (g197)) + ((!ax100x) & (g174) & (g186) & (!g195) & (!g197)) + ((!ax100x) & (g174) & (g186) & (g195) & (!g197)) + ((!ax100x) & (g174) & (g186) & (g195) & (g197)) + ((ax100x) & (!g174) & (!g186) & (!g195) & (!g197)) + ((ax100x) & (!g174) & (!g186) & (g195) & (!g197)) + ((ax100x) & (!g174) & (!g186) & (g195) & (g197)) + ((ax100x) & (g174) & (!g186) & (!g195) & (!g197)) + ((ax100x) & (g174) & (!g186) & (!g195) & (g197)) + ((ax100x) & (g174) & (!g186) & (g195) & (!g197)) + ((ax100x) & (g174) & (!g186) & (g195) & (g197)) + ((ax100x) & (g174) & (g186) & (!g195) & (g197)));
	assign g216 = (((!ax96x) & (!ax97x)));
	assign g217 = (((!g174) & (!ax98x) & (!ax99x) & (!g195) & (!g197) & (!g216)) + ((!g174) & (!ax98x) & (!ax99x) & (g195) & (!g197) & (!g216)) + ((!g174) & (!ax98x) & (!ax99x) & (g195) & (g197) & (!g216)) + ((!g174) & (!ax98x) & (ax99x) & (!g195) & (g197) & (!g216)) + ((!g174) & (ax98x) & (ax99x) & (!g195) & (g197) & (!g216)) + ((!g174) & (ax98x) & (ax99x) & (!g195) & (g197) & (g216)) + ((g174) & (!ax98x) & (!ax99x) & (!g195) & (!g197) & (!g216)) + ((g174) & (!ax98x) & (!ax99x) & (!g195) & (!g197) & (g216)) + ((g174) & (!ax98x) & (!ax99x) & (!g195) & (g197) & (!g216)) + ((g174) & (!ax98x) & (!ax99x) & (g195) & (!g197) & (!g216)) + ((g174) & (!ax98x) & (!ax99x) & (g195) & (!g197) & (g216)) + ((g174) & (!ax98x) & (!ax99x) & (g195) & (g197) & (!g216)) + ((g174) & (!ax98x) & (!ax99x) & (g195) & (g197) & (g216)) + ((g174) & (!ax98x) & (ax99x) & (!g195) & (!g197) & (!g216)) + ((g174) & (!ax98x) & (ax99x) & (!g195) & (g197) & (!g216)) + ((g174) & (!ax98x) & (ax99x) & (!g195) & (g197) & (g216)) + ((g174) & (!ax98x) & (ax99x) & (g195) & (!g197) & (!g216)) + ((g174) & (!ax98x) & (ax99x) & (g195) & (g197) & (!g216)) + ((g174) & (ax98x) & (!ax99x) & (!g195) & (g197) & (!g216)) + ((g174) & (ax98x) & (!ax99x) & (!g195) & (g197) & (g216)) + ((g174) & (ax98x) & (ax99x) & (!g195) & (!g197) & (!g216)) + ((g174) & (ax98x) & (ax99x) & (!g195) & (!g197) & (g216)) + ((g174) & (ax98x) & (ax99x) & (!g195) & (g197) & (!g216)) + ((g174) & (ax98x) & (ax99x) & (!g195) & (g197) & (g216)) + ((g174) & (ax98x) & (ax99x) & (g195) & (!g197) & (!g216)) + ((g174) & (ax98x) & (ax99x) & (g195) & (!g197) & (g216)) + ((g174) & (ax98x) & (ax99x) & (g195) & (g197) & (!g216)) + ((g174) & (ax98x) & (ax99x) & (g195) & (g197) & (g216)));
	assign g218 = (((!g127) & (!g147) & (g214) & (g215) & (g217)) + ((!g127) & (g147) & (g214) & (!g215) & (g217)) + ((!g127) & (g147) & (g214) & (g215) & (!g217)) + ((!g127) & (g147) & (g214) & (g215) & (g217)) + ((g127) & (!g147) & (!g214) & (g215) & (g217)) + ((g127) & (!g147) & (g214) & (!g215) & (!g217)) + ((g127) & (!g147) & (g214) & (!g215) & (g217)) + ((g127) & (!g147) & (g214) & (g215) & (!g217)) + ((g127) & (!g147) & (g214) & (g215) & (g217)) + ((g127) & (g147) & (!g214) & (!g215) & (g217)) + ((g127) & (g147) & (!g214) & (g215) & (!g217)) + ((g127) & (g147) & (!g214) & (g215) & (g217)) + ((g127) & (g147) & (g214) & (!g215) & (!g217)) + ((g127) & (g147) & (g214) & (!g215) & (g217)) + ((g127) & (g147) & (g214) & (g215) & (!g217)) + ((g127) & (g147) & (g214) & (g215) & (g217)));
	assign g219 = (((!g87) & (!g104) & (g211) & (g212) & (g218)) + ((!g87) & (g104) & (g211) & (!g212) & (g218)) + ((!g87) & (g104) & (g211) & (g212) & (!g218)) + ((!g87) & (g104) & (g211) & (g212) & (g218)) + ((g87) & (!g104) & (!g211) & (g212) & (g218)) + ((g87) & (!g104) & (g211) & (!g212) & (!g218)) + ((g87) & (!g104) & (g211) & (!g212) & (g218)) + ((g87) & (!g104) & (g211) & (g212) & (!g218)) + ((g87) & (!g104) & (g211) & (g212) & (g218)) + ((g87) & (g104) & (!g211) & (!g212) & (g218)) + ((g87) & (g104) & (!g211) & (g212) & (!g218)) + ((g87) & (g104) & (!g211) & (g212) & (g218)) + ((g87) & (g104) & (g211) & (!g212) & (!g218)) + ((g87) & (g104) & (g211) & (!g212) & (g218)) + ((g87) & (g104) & (g211) & (g212) & (!g218)) + ((g87) & (g104) & (g211) & (g212) & (g218)));
	assign g220 = (((!g54) & (!g68) & (g208) & (g209) & (g219)) + ((!g54) & (g68) & (g208) & (!g209) & (g219)) + ((!g54) & (g68) & (g208) & (g209) & (!g219)) + ((!g54) & (g68) & (g208) & (g209) & (g219)) + ((g54) & (!g68) & (!g208) & (g209) & (g219)) + ((g54) & (!g68) & (g208) & (!g209) & (!g219)) + ((g54) & (!g68) & (g208) & (!g209) & (g219)) + ((g54) & (!g68) & (g208) & (g209) & (!g219)) + ((g54) & (!g68) & (g208) & (g209) & (g219)) + ((g54) & (g68) & (!g208) & (!g209) & (g219)) + ((g54) & (g68) & (!g208) & (g209) & (!g219)) + ((g54) & (g68) & (!g208) & (g209) & (g219)) + ((g54) & (g68) & (g208) & (!g209) & (!g219)) + ((g54) & (g68) & (g208) & (!g209) & (g219)) + ((g54) & (g68) & (g208) & (g209) & (!g219)) + ((g54) & (g68) & (g208) & (g209) & (g219)));
	assign g221 = (((!g27) & (!g39) & (g205) & (g206) & (g220)) + ((!g27) & (g39) & (g205) & (!g206) & (g220)) + ((!g27) & (g39) & (g205) & (g206) & (!g220)) + ((!g27) & (g39) & (g205) & (g206) & (g220)) + ((g27) & (!g39) & (!g205) & (g206) & (g220)) + ((g27) & (!g39) & (g205) & (!g206) & (!g220)) + ((g27) & (!g39) & (g205) & (!g206) & (g220)) + ((g27) & (!g39) & (g205) & (g206) & (!g220)) + ((g27) & (!g39) & (g205) & (g206) & (g220)) + ((g27) & (g39) & (!g205) & (!g206) & (g220)) + ((g27) & (g39) & (!g205) & (g206) & (!g220)) + ((g27) & (g39) & (!g205) & (g206) & (g220)) + ((g27) & (g39) & (g205) & (!g206) & (!g220)) + ((g27) & (g39) & (g205) & (!g206) & (g220)) + ((g27) & (g39) & (g205) & (g206) & (!g220)) + ((g27) & (g39) & (g205) & (g206) & (g220)));
	assign g222 = (((!g8) & (!g18) & (g202) & (g203) & (g221)) + ((!g8) & (g18) & (g202) & (!g203) & (g221)) + ((!g8) & (g18) & (g202) & (g203) & (!g221)) + ((!g8) & (g18) & (g202) & (g203) & (g221)) + ((g8) & (!g18) & (!g202) & (g203) & (g221)) + ((g8) & (!g18) & (g202) & (!g203) & (!g221)) + ((g8) & (!g18) & (g202) & (!g203) & (g221)) + ((g8) & (!g18) & (g202) & (g203) & (!g221)) + ((g8) & (!g18) & (g202) & (g203) & (g221)) + ((g8) & (g18) & (!g202) & (!g203) & (g221)) + ((g8) & (g18) & (!g202) & (g203) & (!g221)) + ((g8) & (g18) & (!g202) & (g203) & (g221)) + ((g8) & (g18) & (g202) & (!g203) & (!g221)) + ((g8) & (g18) & (g202) & (!g203) & (g221)) + ((g8) & (g18) & (g202) & (g203) & (!g221)) + ((g8) & (g18) & (g202) & (g203) & (g221)));
	assign g223 = (((!g2) & (!g8) & (g177) & (g191)) + ((!g2) & (g8) & (!g177) & (g191)) + ((!g2) & (g8) & (g177) & (!g191)) + ((!g2) & (g8) & (g177) & (g191)) + ((g2) & (!g8) & (!g177) & (!g191)) + ((g2) & (!g8) & (!g177) & (g191)) + ((g2) & (!g8) & (g177) & (!g191)) + ((g2) & (g8) & (!g177) & (!g191)));
	assign g224 = (((!g176) & (!g195) & (!g197) & (g223)) + ((!g176) & (g195) & (!g197) & (g223)) + ((!g176) & (g195) & (g197) & (g223)) + ((g176) & (!g195) & (!g197) & (!g223)) + ((g176) & (!g195) & (g197) & (!g223)) + ((g176) & (!g195) & (g197) & (g223)) + ((g176) & (g195) & (!g197) & (!g223)) + ((g176) & (g195) & (g197) & (!g223)));
	assign g225 = (((!g4) & (!g2) & (!g200) & (!g222) & (g224)) + ((!g4) & (!g2) & (!g200) & (g222) & (g224)) + ((!g4) & (!g2) & (g200) & (!g222) & (g224)) + ((!g4) & (!g2) & (g200) & (g222) & (!g224)) + ((!g4) & (!g2) & (g200) & (g222) & (g224)) + ((!g4) & (g2) & (!g200) & (!g222) & (g224)) + ((!g4) & (g2) & (!g200) & (g222) & (!g224)) + ((!g4) & (g2) & (!g200) & (g222) & (g224)) + ((!g4) & (g2) & (g200) & (!g222) & (!g224)) + ((!g4) & (g2) & (g200) & (!g222) & (g224)) + ((!g4) & (g2) & (g200) & (g222) & (!g224)) + ((!g4) & (g2) & (g200) & (g222) & (g224)) + ((g4) & (!g2) & (g200) & (g222) & (g224)) + ((g4) & (g2) & (!g200) & (g222) & (g224)) + ((g4) & (g2) & (g200) & (!g222) & (g224)) + ((g4) & (g2) & (g200) & (g222) & (g224)));
	assign g226 = (((!g4) & (!g192) & (g193)) + ((!g4) & (g192) & (!g193)) + ((!g4) & (g192) & (g193)) + ((g4) & (g192) & (g193)));
	assign g227 = (((!g175) & (!g226) & (!g195) & (!g197)) + ((!g175) & (!g226) & (g195) & (!g197)) + ((!g175) & (!g226) & (g195) & (g197)) + ((g175) & (g226) & (!g195) & (!g197)) + ((g175) & (g226) & (!g195) & (g197)) + ((g175) & (g226) & (g195) & (!g197)) + ((g175) & (g226) & (g195) & (g197)));
	assign g228 = (((!g1) & (g175) & (!g226) & (!g195) & (!g196)) + ((g1) & (!g175) & (g226) & (!g195) & (g196)) + ((g1) & (!g175) & (g226) & (g195) & (g196)) + ((g1) & (g175) & (!g226) & (!g195) & (!g196)) + ((g1) & (g175) & (!g226) & (!g195) & (g196)) + ((g1) & (g175) & (!g226) & (g195) & (!g196)) + ((g1) & (g175) & (!g226) & (g195) & (g196)));
	assign g229 = (((!g1) & (!g199) & (!g225) & (!g227) & (!g228)) + ((g1) & (!g199) & (!g225) & (!g227) & (!g228)) + ((g1) & (!g199) & (!g225) & (g227) & (!g228)) + ((g1) & (!g199) & (g225) & (!g227) & (!g228)) + ((g1) & (!g199) & (g225) & (g227) & (!g228)) + ((g1) & (g199) & (!g225) & (!g227) & (!g228)) + ((g1) & (g199) & (!g225) & (g227) & (!g228)));
	assign g230 = (((g1) & (!g199) & (g225) & (g228)) + ((g1) & (g199) & (!g225) & (!g228)) + ((g1) & (g199) & (!g225) & (g228)));
	assign g231 = (((!g4) & (!g2) & (!g200) & (!g222) & (!g224) & (!g229)) + ((!g4) & (!g2) & (!g200) & (!g222) & (g224) & (g229)) + ((!g4) & (!g2) & (!g200) & (g222) & (!g224) & (!g229)) + ((!g4) & (!g2) & (!g200) & (g222) & (g224) & (g229)) + ((!g4) & (!g2) & (g200) & (!g222) & (!g224) & (!g229)) + ((!g4) & (!g2) & (g200) & (!g222) & (g224) & (g229)) + ((!g4) & (!g2) & (g200) & (g222) & (g224) & (!g229)) + ((!g4) & (!g2) & (g200) & (g222) & (g224) & (g229)) + ((!g4) & (g2) & (!g200) & (!g222) & (!g224) & (!g229)) + ((!g4) & (g2) & (!g200) & (!g222) & (g224) & (g229)) + ((!g4) & (g2) & (!g200) & (g222) & (g224) & (!g229)) + ((!g4) & (g2) & (!g200) & (g222) & (g224) & (g229)) + ((!g4) & (g2) & (g200) & (!g222) & (g224) & (!g229)) + ((!g4) & (g2) & (g200) & (!g222) & (g224) & (g229)) + ((!g4) & (g2) & (g200) & (g222) & (g224) & (!g229)) + ((!g4) & (g2) & (g200) & (g222) & (g224) & (g229)) + ((g4) & (!g2) & (!g200) & (!g222) & (g224) & (!g229)) + ((g4) & (!g2) & (!g200) & (!g222) & (g224) & (g229)) + ((g4) & (!g2) & (!g200) & (g222) & (g224) & (!g229)) + ((g4) & (!g2) & (!g200) & (g222) & (g224) & (g229)) + ((g4) & (!g2) & (g200) & (!g222) & (g224) & (!g229)) + ((g4) & (!g2) & (g200) & (!g222) & (g224) & (g229)) + ((g4) & (!g2) & (g200) & (g222) & (!g224) & (!g229)) + ((g4) & (!g2) & (g200) & (g222) & (g224) & (g229)) + ((g4) & (g2) & (!g200) & (!g222) & (g224) & (!g229)) + ((g4) & (g2) & (!g200) & (!g222) & (g224) & (g229)) + ((g4) & (g2) & (!g200) & (g222) & (!g224) & (!g229)) + ((g4) & (g2) & (!g200) & (g222) & (g224) & (g229)) + ((g4) & (g2) & (g200) & (!g222) & (!g224) & (!g229)) + ((g4) & (g2) & (g200) & (!g222) & (g224) & (g229)) + ((g4) & (g2) & (g200) & (g222) & (!g224) & (!g229)) + ((g4) & (g2) & (g200) & (g222) & (g224) & (g229)));
	assign g232 = (((!g8) & (!g18) & (!g202) & (g203) & (g221) & (!g229)) + ((!g8) & (!g18) & (g202) & (!g203) & (!g221) & (!g229)) + ((!g8) & (!g18) & (g202) & (!g203) & (!g221) & (g229)) + ((!g8) & (!g18) & (g202) & (!g203) & (g221) & (!g229)) + ((!g8) & (!g18) & (g202) & (!g203) & (g221) & (g229)) + ((!g8) & (!g18) & (g202) & (g203) & (!g221) & (!g229)) + ((!g8) & (!g18) & (g202) & (g203) & (!g221) & (g229)) + ((!g8) & (!g18) & (g202) & (g203) & (g221) & (g229)) + ((!g8) & (g18) & (!g202) & (!g203) & (g221) & (!g229)) + ((!g8) & (g18) & (!g202) & (g203) & (!g221) & (!g229)) + ((!g8) & (g18) & (!g202) & (g203) & (g221) & (!g229)) + ((!g8) & (g18) & (g202) & (!g203) & (!g221) & (!g229)) + ((!g8) & (g18) & (g202) & (!g203) & (!g221) & (g229)) + ((!g8) & (g18) & (g202) & (!g203) & (g221) & (g229)) + ((!g8) & (g18) & (g202) & (g203) & (!g221) & (g229)) + ((!g8) & (g18) & (g202) & (g203) & (g221) & (g229)) + ((g8) & (!g18) & (!g202) & (!g203) & (!g221) & (!g229)) + ((g8) & (!g18) & (!g202) & (!g203) & (g221) & (!g229)) + ((g8) & (!g18) & (!g202) & (g203) & (!g221) & (!g229)) + ((g8) & (!g18) & (g202) & (!g203) & (!g221) & (g229)) + ((g8) & (!g18) & (g202) & (!g203) & (g221) & (g229)) + ((g8) & (!g18) & (g202) & (g203) & (!g221) & (g229)) + ((g8) & (!g18) & (g202) & (g203) & (g221) & (!g229)) + ((g8) & (!g18) & (g202) & (g203) & (g221) & (g229)) + ((g8) & (g18) & (!g202) & (!g203) & (!g221) & (!g229)) + ((g8) & (g18) & (g202) & (!g203) & (!g221) & (g229)) + ((g8) & (g18) & (g202) & (!g203) & (g221) & (!g229)) + ((g8) & (g18) & (g202) & (!g203) & (g221) & (g229)) + ((g8) & (g18) & (g202) & (g203) & (!g221) & (!g229)) + ((g8) & (g18) & (g202) & (g203) & (!g221) & (g229)) + ((g8) & (g18) & (g202) & (g203) & (g221) & (!g229)) + ((g8) & (g18) & (g202) & (g203) & (g221) & (g229)));
	assign g233 = (((!g18) & (!g203) & (g221) & (!g229)) + ((!g18) & (g203) & (!g221) & (!g229)) + ((!g18) & (g203) & (!g221) & (g229)) + ((!g18) & (g203) & (g221) & (g229)) + ((g18) & (!g203) & (!g221) & (!g229)) + ((g18) & (g203) & (!g221) & (g229)) + ((g18) & (g203) & (g221) & (!g229)) + ((g18) & (g203) & (g221) & (g229)));
	assign g234 = (((!g27) & (!g39) & (!g205) & (g206) & (g220) & (!g229)) + ((!g27) & (!g39) & (g205) & (!g206) & (!g220) & (!g229)) + ((!g27) & (!g39) & (g205) & (!g206) & (!g220) & (g229)) + ((!g27) & (!g39) & (g205) & (!g206) & (g220) & (!g229)) + ((!g27) & (!g39) & (g205) & (!g206) & (g220) & (g229)) + ((!g27) & (!g39) & (g205) & (g206) & (!g220) & (!g229)) + ((!g27) & (!g39) & (g205) & (g206) & (!g220) & (g229)) + ((!g27) & (!g39) & (g205) & (g206) & (g220) & (g229)) + ((!g27) & (g39) & (!g205) & (!g206) & (g220) & (!g229)) + ((!g27) & (g39) & (!g205) & (g206) & (!g220) & (!g229)) + ((!g27) & (g39) & (!g205) & (g206) & (g220) & (!g229)) + ((!g27) & (g39) & (g205) & (!g206) & (!g220) & (!g229)) + ((!g27) & (g39) & (g205) & (!g206) & (!g220) & (g229)) + ((!g27) & (g39) & (g205) & (!g206) & (g220) & (g229)) + ((!g27) & (g39) & (g205) & (g206) & (!g220) & (g229)) + ((!g27) & (g39) & (g205) & (g206) & (g220) & (g229)) + ((g27) & (!g39) & (!g205) & (!g206) & (!g220) & (!g229)) + ((g27) & (!g39) & (!g205) & (!g206) & (g220) & (!g229)) + ((g27) & (!g39) & (!g205) & (g206) & (!g220) & (!g229)) + ((g27) & (!g39) & (g205) & (!g206) & (!g220) & (g229)) + ((g27) & (!g39) & (g205) & (!g206) & (g220) & (g229)) + ((g27) & (!g39) & (g205) & (g206) & (!g220) & (g229)) + ((g27) & (!g39) & (g205) & (g206) & (g220) & (!g229)) + ((g27) & (!g39) & (g205) & (g206) & (g220) & (g229)) + ((g27) & (g39) & (!g205) & (!g206) & (!g220) & (!g229)) + ((g27) & (g39) & (g205) & (!g206) & (!g220) & (g229)) + ((g27) & (g39) & (g205) & (!g206) & (g220) & (!g229)) + ((g27) & (g39) & (g205) & (!g206) & (g220) & (g229)) + ((g27) & (g39) & (g205) & (g206) & (!g220) & (!g229)) + ((g27) & (g39) & (g205) & (g206) & (!g220) & (g229)) + ((g27) & (g39) & (g205) & (g206) & (g220) & (!g229)) + ((g27) & (g39) & (g205) & (g206) & (g220) & (g229)));
	assign g235 = (((!g39) & (!g206) & (g220) & (!g229)) + ((!g39) & (g206) & (!g220) & (!g229)) + ((!g39) & (g206) & (!g220) & (g229)) + ((!g39) & (g206) & (g220) & (g229)) + ((g39) & (!g206) & (!g220) & (!g229)) + ((g39) & (g206) & (!g220) & (g229)) + ((g39) & (g206) & (g220) & (!g229)) + ((g39) & (g206) & (g220) & (g229)));
	assign g236 = (((!g54) & (!g68) & (!g208) & (g209) & (g219) & (!g229)) + ((!g54) & (!g68) & (g208) & (!g209) & (!g219) & (!g229)) + ((!g54) & (!g68) & (g208) & (!g209) & (!g219) & (g229)) + ((!g54) & (!g68) & (g208) & (!g209) & (g219) & (!g229)) + ((!g54) & (!g68) & (g208) & (!g209) & (g219) & (g229)) + ((!g54) & (!g68) & (g208) & (g209) & (!g219) & (!g229)) + ((!g54) & (!g68) & (g208) & (g209) & (!g219) & (g229)) + ((!g54) & (!g68) & (g208) & (g209) & (g219) & (g229)) + ((!g54) & (g68) & (!g208) & (!g209) & (g219) & (!g229)) + ((!g54) & (g68) & (!g208) & (g209) & (!g219) & (!g229)) + ((!g54) & (g68) & (!g208) & (g209) & (g219) & (!g229)) + ((!g54) & (g68) & (g208) & (!g209) & (!g219) & (!g229)) + ((!g54) & (g68) & (g208) & (!g209) & (!g219) & (g229)) + ((!g54) & (g68) & (g208) & (!g209) & (g219) & (g229)) + ((!g54) & (g68) & (g208) & (g209) & (!g219) & (g229)) + ((!g54) & (g68) & (g208) & (g209) & (g219) & (g229)) + ((g54) & (!g68) & (!g208) & (!g209) & (!g219) & (!g229)) + ((g54) & (!g68) & (!g208) & (!g209) & (g219) & (!g229)) + ((g54) & (!g68) & (!g208) & (g209) & (!g219) & (!g229)) + ((g54) & (!g68) & (g208) & (!g209) & (!g219) & (g229)) + ((g54) & (!g68) & (g208) & (!g209) & (g219) & (g229)) + ((g54) & (!g68) & (g208) & (g209) & (!g219) & (g229)) + ((g54) & (!g68) & (g208) & (g209) & (g219) & (!g229)) + ((g54) & (!g68) & (g208) & (g209) & (g219) & (g229)) + ((g54) & (g68) & (!g208) & (!g209) & (!g219) & (!g229)) + ((g54) & (g68) & (g208) & (!g209) & (!g219) & (g229)) + ((g54) & (g68) & (g208) & (!g209) & (g219) & (!g229)) + ((g54) & (g68) & (g208) & (!g209) & (g219) & (g229)) + ((g54) & (g68) & (g208) & (g209) & (!g219) & (!g229)) + ((g54) & (g68) & (g208) & (g209) & (!g219) & (g229)) + ((g54) & (g68) & (g208) & (g209) & (g219) & (!g229)) + ((g54) & (g68) & (g208) & (g209) & (g219) & (g229)));
	assign g237 = (((!g68) & (!g209) & (g219) & (!g229)) + ((!g68) & (g209) & (!g219) & (!g229)) + ((!g68) & (g209) & (!g219) & (g229)) + ((!g68) & (g209) & (g219) & (g229)) + ((g68) & (!g209) & (!g219) & (!g229)) + ((g68) & (g209) & (!g219) & (g229)) + ((g68) & (g209) & (g219) & (!g229)) + ((g68) & (g209) & (g219) & (g229)));
	assign g238 = (((!g87) & (!g104) & (!g211) & (g212) & (g218) & (!g229)) + ((!g87) & (!g104) & (g211) & (!g212) & (!g218) & (!g229)) + ((!g87) & (!g104) & (g211) & (!g212) & (!g218) & (g229)) + ((!g87) & (!g104) & (g211) & (!g212) & (g218) & (!g229)) + ((!g87) & (!g104) & (g211) & (!g212) & (g218) & (g229)) + ((!g87) & (!g104) & (g211) & (g212) & (!g218) & (!g229)) + ((!g87) & (!g104) & (g211) & (g212) & (!g218) & (g229)) + ((!g87) & (!g104) & (g211) & (g212) & (g218) & (g229)) + ((!g87) & (g104) & (!g211) & (!g212) & (g218) & (!g229)) + ((!g87) & (g104) & (!g211) & (g212) & (!g218) & (!g229)) + ((!g87) & (g104) & (!g211) & (g212) & (g218) & (!g229)) + ((!g87) & (g104) & (g211) & (!g212) & (!g218) & (!g229)) + ((!g87) & (g104) & (g211) & (!g212) & (!g218) & (g229)) + ((!g87) & (g104) & (g211) & (!g212) & (g218) & (g229)) + ((!g87) & (g104) & (g211) & (g212) & (!g218) & (g229)) + ((!g87) & (g104) & (g211) & (g212) & (g218) & (g229)) + ((g87) & (!g104) & (!g211) & (!g212) & (!g218) & (!g229)) + ((g87) & (!g104) & (!g211) & (!g212) & (g218) & (!g229)) + ((g87) & (!g104) & (!g211) & (g212) & (!g218) & (!g229)) + ((g87) & (!g104) & (g211) & (!g212) & (!g218) & (g229)) + ((g87) & (!g104) & (g211) & (!g212) & (g218) & (g229)) + ((g87) & (!g104) & (g211) & (g212) & (!g218) & (g229)) + ((g87) & (!g104) & (g211) & (g212) & (g218) & (!g229)) + ((g87) & (!g104) & (g211) & (g212) & (g218) & (g229)) + ((g87) & (g104) & (!g211) & (!g212) & (!g218) & (!g229)) + ((g87) & (g104) & (g211) & (!g212) & (!g218) & (g229)) + ((g87) & (g104) & (g211) & (!g212) & (g218) & (!g229)) + ((g87) & (g104) & (g211) & (!g212) & (g218) & (g229)) + ((g87) & (g104) & (g211) & (g212) & (!g218) & (!g229)) + ((g87) & (g104) & (g211) & (g212) & (!g218) & (g229)) + ((g87) & (g104) & (g211) & (g212) & (g218) & (!g229)) + ((g87) & (g104) & (g211) & (g212) & (g218) & (g229)));
	assign g239 = (((!g104) & (!g212) & (g218) & (!g229)) + ((!g104) & (g212) & (!g218) & (!g229)) + ((!g104) & (g212) & (!g218) & (g229)) + ((!g104) & (g212) & (g218) & (g229)) + ((g104) & (!g212) & (!g218) & (!g229)) + ((g104) & (g212) & (!g218) & (g229)) + ((g104) & (g212) & (g218) & (!g229)) + ((g104) & (g212) & (g218) & (g229)));
	assign g240 = (((!g127) & (!g147) & (!g214) & (g215) & (g217) & (!g229)) + ((!g127) & (!g147) & (g214) & (!g215) & (!g217) & (!g229)) + ((!g127) & (!g147) & (g214) & (!g215) & (!g217) & (g229)) + ((!g127) & (!g147) & (g214) & (!g215) & (g217) & (!g229)) + ((!g127) & (!g147) & (g214) & (!g215) & (g217) & (g229)) + ((!g127) & (!g147) & (g214) & (g215) & (!g217) & (!g229)) + ((!g127) & (!g147) & (g214) & (g215) & (!g217) & (g229)) + ((!g127) & (!g147) & (g214) & (g215) & (g217) & (g229)) + ((!g127) & (g147) & (!g214) & (!g215) & (g217) & (!g229)) + ((!g127) & (g147) & (!g214) & (g215) & (!g217) & (!g229)) + ((!g127) & (g147) & (!g214) & (g215) & (g217) & (!g229)) + ((!g127) & (g147) & (g214) & (!g215) & (!g217) & (!g229)) + ((!g127) & (g147) & (g214) & (!g215) & (!g217) & (g229)) + ((!g127) & (g147) & (g214) & (!g215) & (g217) & (g229)) + ((!g127) & (g147) & (g214) & (g215) & (!g217) & (g229)) + ((!g127) & (g147) & (g214) & (g215) & (g217) & (g229)) + ((g127) & (!g147) & (!g214) & (!g215) & (!g217) & (!g229)) + ((g127) & (!g147) & (!g214) & (!g215) & (g217) & (!g229)) + ((g127) & (!g147) & (!g214) & (g215) & (!g217) & (!g229)) + ((g127) & (!g147) & (g214) & (!g215) & (!g217) & (g229)) + ((g127) & (!g147) & (g214) & (!g215) & (g217) & (g229)) + ((g127) & (!g147) & (g214) & (g215) & (!g217) & (g229)) + ((g127) & (!g147) & (g214) & (g215) & (g217) & (!g229)) + ((g127) & (!g147) & (g214) & (g215) & (g217) & (g229)) + ((g127) & (g147) & (!g214) & (!g215) & (!g217) & (!g229)) + ((g127) & (g147) & (g214) & (!g215) & (!g217) & (g229)) + ((g127) & (g147) & (g214) & (!g215) & (g217) & (!g229)) + ((g127) & (g147) & (g214) & (!g215) & (g217) & (g229)) + ((g127) & (g147) & (g214) & (g215) & (!g217) & (!g229)) + ((g127) & (g147) & (g214) & (g215) & (!g217) & (g229)) + ((g127) & (g147) & (g214) & (g215) & (g217) & (!g229)) + ((g127) & (g147) & (g214) & (g215) & (g217) & (g229)));
	assign g241 = (((!g147) & (!g215) & (g217) & (!g229)) + ((!g147) & (g215) & (!g217) & (!g229)) + ((!g147) & (g215) & (!g217) & (g229)) + ((!g147) & (g215) & (g217) & (g229)) + ((g147) & (!g215) & (!g217) & (!g229)) + ((g147) & (g215) & (!g217) & (g229)) + ((g147) & (g215) & (g217) & (!g229)) + ((g147) & (g215) & (g217) & (g229)));
	assign g242 = (((!g174) & (!ax98x) & (!ax99x) & (!g198) & (!g216) & (g229)) + ((!g174) & (!ax98x) & (!ax99x) & (!g198) & (g216) & (!g229)) + ((!g174) & (!ax98x) & (!ax99x) & (!g198) & (g216) & (g229)) + ((!g174) & (!ax98x) & (!ax99x) & (g198) & (!g216) & (!g229)) + ((!g174) & (!ax98x) & (ax99x) & (!g198) & (!g216) & (!g229)) + ((!g174) & (!ax98x) & (ax99x) & (g198) & (!g216) & (g229)) + ((!g174) & (!ax98x) & (ax99x) & (g198) & (g216) & (!g229)) + ((!g174) & (!ax98x) & (ax99x) & (g198) & (g216) & (g229)) + ((!g174) & (ax98x) & (!ax99x) & (g198) & (!g216) & (!g229)) + ((!g174) & (ax98x) & (!ax99x) & (g198) & (g216) & (!g229)) + ((!g174) & (ax98x) & (ax99x) & (!g198) & (!g216) & (!g229)) + ((!g174) & (ax98x) & (ax99x) & (!g198) & (!g216) & (g229)) + ((!g174) & (ax98x) & (ax99x) & (!g198) & (g216) & (!g229)) + ((!g174) & (ax98x) & (ax99x) & (!g198) & (g216) & (g229)) + ((!g174) & (ax98x) & (ax99x) & (g198) & (!g216) & (g229)) + ((!g174) & (ax98x) & (ax99x) & (g198) & (g216) & (g229)) + ((g174) & (!ax98x) & (!ax99x) & (!g198) & (!g216) & (!g229)) + ((g174) & (!ax98x) & (!ax99x) & (!g198) & (!g216) & (g229)) + ((g174) & (!ax98x) & (!ax99x) & (!g198) & (g216) & (g229)) + ((g174) & (!ax98x) & (!ax99x) & (g198) & (g216) & (!g229)) + ((g174) & (!ax98x) & (ax99x) & (!g198) & (g216) & (!g229)) + ((g174) & (!ax98x) & (ax99x) & (g198) & (!g216) & (!g229)) + ((g174) & (!ax98x) & (ax99x) & (g198) & (!g216) & (g229)) + ((g174) & (!ax98x) & (ax99x) & (g198) & (g216) & (g229)) + ((g174) & (ax98x) & (!ax99x) & (!g198) & (!g216) & (!g229)) + ((g174) & (ax98x) & (!ax99x) & (!g198) & (g216) & (!g229)) + ((g174) & (ax98x) & (ax99x) & (!g198) & (!g216) & (g229)) + ((g174) & (ax98x) & (ax99x) & (!g198) & (g216) & (g229)) + ((g174) & (ax98x) & (ax99x) & (g198) & (!g216) & (!g229)) + ((g174) & (ax98x) & (ax99x) & (g198) & (!g216) & (g229)) + ((g174) & (ax98x) & (ax99x) & (g198) & (g216) & (!g229)) + ((g174) & (ax98x) & (ax99x) & (g198) & (g216) & (g229)));
	assign g243 = (((!ax98x) & (!g198) & (!g216) & (g229)) + ((!ax98x) & (!g198) & (g216) & (!g229)) + ((!ax98x) & (!g198) & (g216) & (g229)) + ((!ax98x) & (g198) & (g216) & (!g229)) + ((ax98x) & (!g198) & (!g216) & (!g229)) + ((ax98x) & (g198) & (!g216) & (!g229)) + ((ax98x) & (g198) & (!g216) & (g229)) + ((ax98x) & (g198) & (g216) & (g229)));
	assign g244 = (((!ax94x) & (!ax95x)));
	assign g245 = (((!ax96x) & (!ax97x) & (!g198) & (!g229) & (!g244)) + ((!ax96x) & (!ax97x) & (g198) & (!g229) & (!g244)) + ((!ax96x) & (!ax97x) & (g198) & (!g229) & (g244)) + ((!ax96x) & (!ax97x) & (g198) & (g229) & (!g244)) + ((!ax96x) & (ax97x) & (!g198) & (g229) & (!g244)) + ((!ax96x) & (ax97x) & (g198) & (!g229) & (!g244)) + ((!ax96x) & (ax97x) & (g198) & (g229) & (!g244)) + ((!ax96x) & (ax97x) & (g198) & (g229) & (g244)) + ((ax96x) & (!ax97x) & (g198) & (g229) & (!g244)) + ((ax96x) & (!ax97x) & (g198) & (g229) & (g244)) + ((ax96x) & (ax97x) & (!g198) & (g229) & (!g244)) + ((ax96x) & (ax97x) & (!g198) & (g229) & (g244)) + ((ax96x) & (ax97x) & (g198) & (!g229) & (!g244)) + ((ax96x) & (ax97x) & (g198) & (!g229) & (g244)) + ((ax96x) & (ax97x) & (g198) & (g229) & (!g244)) + ((ax96x) & (ax97x) & (g198) & (g229) & (g244)));
	assign g246 = (((!g147) & (!g174) & (g242) & (g243) & (g245)) + ((!g147) & (g174) & (g242) & (!g243) & (g245)) + ((!g147) & (g174) & (g242) & (g243) & (!g245)) + ((!g147) & (g174) & (g242) & (g243) & (g245)) + ((g147) & (!g174) & (!g242) & (g243) & (g245)) + ((g147) & (!g174) & (g242) & (!g243) & (!g245)) + ((g147) & (!g174) & (g242) & (!g243) & (g245)) + ((g147) & (!g174) & (g242) & (g243) & (!g245)) + ((g147) & (!g174) & (g242) & (g243) & (g245)) + ((g147) & (g174) & (!g242) & (!g243) & (g245)) + ((g147) & (g174) & (!g242) & (g243) & (!g245)) + ((g147) & (g174) & (!g242) & (g243) & (g245)) + ((g147) & (g174) & (g242) & (!g243) & (!g245)) + ((g147) & (g174) & (g242) & (!g243) & (g245)) + ((g147) & (g174) & (g242) & (g243) & (!g245)) + ((g147) & (g174) & (g242) & (g243) & (g245)));
	assign g247 = (((!g104) & (!g127) & (g240) & (g241) & (g246)) + ((!g104) & (g127) & (g240) & (!g241) & (g246)) + ((!g104) & (g127) & (g240) & (g241) & (!g246)) + ((!g104) & (g127) & (g240) & (g241) & (g246)) + ((g104) & (!g127) & (!g240) & (g241) & (g246)) + ((g104) & (!g127) & (g240) & (!g241) & (!g246)) + ((g104) & (!g127) & (g240) & (!g241) & (g246)) + ((g104) & (!g127) & (g240) & (g241) & (!g246)) + ((g104) & (!g127) & (g240) & (g241) & (g246)) + ((g104) & (g127) & (!g240) & (!g241) & (g246)) + ((g104) & (g127) & (!g240) & (g241) & (!g246)) + ((g104) & (g127) & (!g240) & (g241) & (g246)) + ((g104) & (g127) & (g240) & (!g241) & (!g246)) + ((g104) & (g127) & (g240) & (!g241) & (g246)) + ((g104) & (g127) & (g240) & (g241) & (!g246)) + ((g104) & (g127) & (g240) & (g241) & (g246)));
	assign g248 = (((!g68) & (!g87) & (g238) & (g239) & (g247)) + ((!g68) & (g87) & (g238) & (!g239) & (g247)) + ((!g68) & (g87) & (g238) & (g239) & (!g247)) + ((!g68) & (g87) & (g238) & (g239) & (g247)) + ((g68) & (!g87) & (!g238) & (g239) & (g247)) + ((g68) & (!g87) & (g238) & (!g239) & (!g247)) + ((g68) & (!g87) & (g238) & (!g239) & (g247)) + ((g68) & (!g87) & (g238) & (g239) & (!g247)) + ((g68) & (!g87) & (g238) & (g239) & (g247)) + ((g68) & (g87) & (!g238) & (!g239) & (g247)) + ((g68) & (g87) & (!g238) & (g239) & (!g247)) + ((g68) & (g87) & (!g238) & (g239) & (g247)) + ((g68) & (g87) & (g238) & (!g239) & (!g247)) + ((g68) & (g87) & (g238) & (!g239) & (g247)) + ((g68) & (g87) & (g238) & (g239) & (!g247)) + ((g68) & (g87) & (g238) & (g239) & (g247)));
	assign g249 = (((!g39) & (!g54) & (g236) & (g237) & (g248)) + ((!g39) & (g54) & (g236) & (!g237) & (g248)) + ((!g39) & (g54) & (g236) & (g237) & (!g248)) + ((!g39) & (g54) & (g236) & (g237) & (g248)) + ((g39) & (!g54) & (!g236) & (g237) & (g248)) + ((g39) & (!g54) & (g236) & (!g237) & (!g248)) + ((g39) & (!g54) & (g236) & (!g237) & (g248)) + ((g39) & (!g54) & (g236) & (g237) & (!g248)) + ((g39) & (!g54) & (g236) & (g237) & (g248)) + ((g39) & (g54) & (!g236) & (!g237) & (g248)) + ((g39) & (g54) & (!g236) & (g237) & (!g248)) + ((g39) & (g54) & (!g236) & (g237) & (g248)) + ((g39) & (g54) & (g236) & (!g237) & (!g248)) + ((g39) & (g54) & (g236) & (!g237) & (g248)) + ((g39) & (g54) & (g236) & (g237) & (!g248)) + ((g39) & (g54) & (g236) & (g237) & (g248)));
	assign g250 = (((!g18) & (!g27) & (g234) & (g235) & (g249)) + ((!g18) & (g27) & (g234) & (!g235) & (g249)) + ((!g18) & (g27) & (g234) & (g235) & (!g249)) + ((!g18) & (g27) & (g234) & (g235) & (g249)) + ((g18) & (!g27) & (!g234) & (g235) & (g249)) + ((g18) & (!g27) & (g234) & (!g235) & (!g249)) + ((g18) & (!g27) & (g234) & (!g235) & (g249)) + ((g18) & (!g27) & (g234) & (g235) & (!g249)) + ((g18) & (!g27) & (g234) & (g235) & (g249)) + ((g18) & (g27) & (!g234) & (!g235) & (g249)) + ((g18) & (g27) & (!g234) & (g235) & (!g249)) + ((g18) & (g27) & (!g234) & (g235) & (g249)) + ((g18) & (g27) & (g234) & (!g235) & (!g249)) + ((g18) & (g27) & (g234) & (!g235) & (g249)) + ((g18) & (g27) & (g234) & (g235) & (!g249)) + ((g18) & (g27) & (g234) & (g235) & (g249)));
	assign g251 = (((!g2) & (!g8) & (g232) & (g233) & (g250)) + ((!g2) & (g8) & (g232) & (!g233) & (g250)) + ((!g2) & (g8) & (g232) & (g233) & (!g250)) + ((!g2) & (g8) & (g232) & (g233) & (g250)) + ((g2) & (!g8) & (!g232) & (g233) & (g250)) + ((g2) & (!g8) & (g232) & (!g233) & (!g250)) + ((g2) & (!g8) & (g232) & (!g233) & (g250)) + ((g2) & (!g8) & (g232) & (g233) & (!g250)) + ((g2) & (!g8) & (g232) & (g233) & (g250)) + ((g2) & (g8) & (!g232) & (!g233) & (g250)) + ((g2) & (g8) & (!g232) & (g233) & (!g250)) + ((g2) & (g8) & (!g232) & (g233) & (g250)) + ((g2) & (g8) & (g232) & (!g233) & (!g250)) + ((g2) & (g8) & (g232) & (!g233) & (g250)) + ((g2) & (g8) & (g232) & (g233) & (!g250)) + ((g2) & (g8) & (g232) & (g233) & (g250)));
	assign g252 = (((!g2) & (!g200) & (g222) & (!g229)) + ((!g2) & (g200) & (!g222) & (!g229)) + ((!g2) & (g200) & (!g222) & (g229)) + ((!g2) & (g200) & (g222) & (g229)) + ((g2) & (!g200) & (!g222) & (!g229)) + ((g2) & (g200) & (!g222) & (g229)) + ((g2) & (g200) & (g222) & (!g229)) + ((g2) & (g200) & (g222) & (g229)));
	assign g253 = (((!g1) & (!g199) & (!g225) & (!g227) & (g228)) + ((!g1) & (!g199) & (!g225) & (g227) & (!g228)) + ((!g1) & (!g199) & (!g225) & (g227) & (g228)) + ((!g1) & (g199) & (g225) & (!g227) & (!g228)) + ((!g1) & (g199) & (g225) & (!g227) & (g228)) + ((!g1) & (g199) & (g225) & (g227) & (!g228)) + ((!g1) & (g199) & (g225) & (g227) & (g228)) + ((g1) & (!g199) & (!g225) & (!g227) & (g228)) + ((g1) & (!g199) & (!g225) & (g227) & (g228)) + ((g1) & (g199) & (g225) & (!g227) & (!g228)) + ((g1) & (g199) & (g225) & (!g227) & (g228)) + ((g1) & (g199) & (g225) & (g227) & (!g228)) + ((g1) & (g199) & (g225) & (g227) & (g228)));
	assign g254 = (((!g4) & (!g1) & (!g231) & (!g251) & (!g252) & (!g253)) + ((!g4) & (g1) & (!g231) & (!g251) & (!g252) & (!g253)) + ((!g4) & (g1) & (!g231) & (!g251) & (!g252) & (g253)) + ((!g4) & (g1) & (!g231) & (!g251) & (g252) & (!g253)) + ((!g4) & (g1) & (!g231) & (!g251) & (g252) & (g253)) + ((!g4) & (g1) & (!g231) & (g251) & (!g252) & (!g253)) + ((!g4) & (g1) & (!g231) & (g251) & (!g252) & (g253)) + ((!g4) & (g1) & (!g231) & (g251) & (g252) & (!g253)) + ((!g4) & (g1) & (!g231) & (g251) & (g252) & (g253)) + ((!g4) & (g1) & (g231) & (!g251) & (!g252) & (!g253)) + ((!g4) & (g1) & (g231) & (!g251) & (!g252) & (g253)) + ((g4) & (!g1) & (!g231) & (!g251) & (!g252) & (!g253)) + ((g4) & (!g1) & (!g231) & (!g251) & (g252) & (!g253)) + ((g4) & (!g1) & (!g231) & (g251) & (!g252) & (!g253)) + ((g4) & (g1) & (!g231) & (!g251) & (!g252) & (!g253)) + ((g4) & (g1) & (!g231) & (!g251) & (!g252) & (g253)) + ((g4) & (g1) & (!g231) & (!g251) & (g252) & (!g253)) + ((g4) & (g1) & (!g231) & (!g251) & (g252) & (g253)) + ((g4) & (g1) & (!g231) & (g251) & (!g252) & (!g253)) + ((g4) & (g1) & (!g231) & (g251) & (!g252) & (g253)) + ((g4) & (g1) & (!g231) & (g251) & (g252) & (!g253)) + ((g4) & (g1) & (!g231) & (g251) & (g252) & (g253)) + ((g4) & (g1) & (g231) & (!g251) & (!g252) & (!g253)) + ((g4) & (g1) & (g231) & (!g251) & (!g252) & (g253)) + ((g4) & (g1) & (g231) & (!g251) & (g252) & (!g253)) + ((g4) & (g1) & (g231) & (!g251) & (g252) & (g253)) + ((g4) & (g1) & (g231) & (g251) & (!g252) & (!g253)) + ((g4) & (g1) & (g231) & (g251) & (!g252) & (g253)));
	assign g255 = (((!g230) & (g254)));
	assign g256 = (((!g4) & (!g251) & (!g252) & (!g230) & (!g254)) + ((!g4) & (!g251) & (!g252) & (g230) & (!g254)) + ((!g4) & (!g251) & (!g252) & (g230) & (g254)) + ((!g4) & (!g251) & (g252) & (!g230) & (g254)) + ((!g4) & (g251) & (g252) & (!g230) & (!g254)) + ((!g4) & (g251) & (g252) & (!g230) & (g254)) + ((!g4) & (g251) & (g252) & (g230) & (!g254)) + ((!g4) & (g251) & (g252) & (g230) & (g254)) + ((g4) & (!g251) & (g252) & (!g230) & (!g254)) + ((g4) & (!g251) & (g252) & (!g230) & (g254)) + ((g4) & (!g251) & (g252) & (g230) & (!g254)) + ((g4) & (!g251) & (g252) & (g230) & (g254)) + ((g4) & (g251) & (!g252) & (!g230) & (!g254)) + ((g4) & (g251) & (!g252) & (g230) & (!g254)) + ((g4) & (g251) & (!g252) & (g230) & (g254)) + ((g4) & (g251) & (g252) & (!g230) & (g254)));
	assign g257 = (((!g8) & (!g233) & (g250) & (!g230) & (!g254)) + ((!g8) & (!g233) & (g250) & (g230) & (!g254)) + ((!g8) & (!g233) & (g250) & (g230) & (g254)) + ((!g8) & (g233) & (!g250) & (!g230) & (!g254)) + ((!g8) & (g233) & (!g250) & (!g230) & (g254)) + ((!g8) & (g233) & (!g250) & (g230) & (!g254)) + ((!g8) & (g233) & (!g250) & (g230) & (g254)) + ((!g8) & (g233) & (g250) & (!g230) & (g254)) + ((g8) & (!g233) & (!g250) & (!g230) & (!g254)) + ((g8) & (!g233) & (!g250) & (g230) & (!g254)) + ((g8) & (!g233) & (!g250) & (g230) & (g254)) + ((g8) & (g233) & (!g250) & (!g230) & (g254)) + ((g8) & (g233) & (g250) & (!g230) & (!g254)) + ((g8) & (g233) & (g250) & (!g230) & (g254)) + ((g8) & (g233) & (g250) & (g230) & (!g254)) + ((g8) & (g233) & (g250) & (g230) & (g254)));
	assign g258 = (((!g18) & (!g27) & (g235) & (g249)) + ((!g18) & (g27) & (!g235) & (g249)) + ((!g18) & (g27) & (g235) & (!g249)) + ((!g18) & (g27) & (g235) & (g249)) + ((g18) & (!g27) & (!g235) & (!g249)) + ((g18) & (!g27) & (!g235) & (g249)) + ((g18) & (!g27) & (g235) & (!g249)) + ((g18) & (g27) & (!g235) & (!g249)));
	assign g259 = (((!g234) & (!g230) & (!g254) & (g258)) + ((!g234) & (g230) & (!g254) & (g258)) + ((!g234) & (g230) & (g254) & (g258)) + ((g234) & (!g230) & (!g254) & (!g258)) + ((g234) & (!g230) & (g254) & (!g258)) + ((g234) & (!g230) & (g254) & (g258)) + ((g234) & (g230) & (!g254) & (!g258)) + ((g234) & (g230) & (g254) & (!g258)));
	assign g260 = (((!g27) & (!g235) & (g249) & (!g230) & (!g254)) + ((!g27) & (!g235) & (g249) & (g230) & (!g254)) + ((!g27) & (!g235) & (g249) & (g230) & (g254)) + ((!g27) & (g235) & (!g249) & (!g230) & (!g254)) + ((!g27) & (g235) & (!g249) & (!g230) & (g254)) + ((!g27) & (g235) & (!g249) & (g230) & (!g254)) + ((!g27) & (g235) & (!g249) & (g230) & (g254)) + ((!g27) & (g235) & (g249) & (!g230) & (g254)) + ((g27) & (!g235) & (!g249) & (!g230) & (!g254)) + ((g27) & (!g235) & (!g249) & (g230) & (!g254)) + ((g27) & (!g235) & (!g249) & (g230) & (g254)) + ((g27) & (g235) & (!g249) & (!g230) & (g254)) + ((g27) & (g235) & (g249) & (!g230) & (!g254)) + ((g27) & (g235) & (g249) & (!g230) & (g254)) + ((g27) & (g235) & (g249) & (g230) & (!g254)) + ((g27) & (g235) & (g249) & (g230) & (g254)));
	assign g261 = (((!g39) & (!g54) & (g237) & (g248)) + ((!g39) & (g54) & (!g237) & (g248)) + ((!g39) & (g54) & (g237) & (!g248)) + ((!g39) & (g54) & (g237) & (g248)) + ((g39) & (!g54) & (!g237) & (!g248)) + ((g39) & (!g54) & (!g237) & (g248)) + ((g39) & (!g54) & (g237) & (!g248)) + ((g39) & (g54) & (!g237) & (!g248)));
	assign g262 = (((!g236) & (!g230) & (!g254) & (g261)) + ((!g236) & (g230) & (!g254) & (g261)) + ((!g236) & (g230) & (g254) & (g261)) + ((g236) & (!g230) & (!g254) & (!g261)) + ((g236) & (!g230) & (g254) & (!g261)) + ((g236) & (!g230) & (g254) & (g261)) + ((g236) & (g230) & (!g254) & (!g261)) + ((g236) & (g230) & (g254) & (!g261)));
	assign g263 = (((!g54) & (!g237) & (g248) & (!g230) & (!g254)) + ((!g54) & (!g237) & (g248) & (g230) & (!g254)) + ((!g54) & (!g237) & (g248) & (g230) & (g254)) + ((!g54) & (g237) & (!g248) & (!g230) & (!g254)) + ((!g54) & (g237) & (!g248) & (!g230) & (g254)) + ((!g54) & (g237) & (!g248) & (g230) & (!g254)) + ((!g54) & (g237) & (!g248) & (g230) & (g254)) + ((!g54) & (g237) & (g248) & (!g230) & (g254)) + ((g54) & (!g237) & (!g248) & (!g230) & (!g254)) + ((g54) & (!g237) & (!g248) & (g230) & (!g254)) + ((g54) & (!g237) & (!g248) & (g230) & (g254)) + ((g54) & (g237) & (!g248) & (!g230) & (g254)) + ((g54) & (g237) & (g248) & (!g230) & (!g254)) + ((g54) & (g237) & (g248) & (!g230) & (g254)) + ((g54) & (g237) & (g248) & (g230) & (!g254)) + ((g54) & (g237) & (g248) & (g230) & (g254)));
	assign g264 = (((!g68) & (!g87) & (g239) & (g247)) + ((!g68) & (g87) & (!g239) & (g247)) + ((!g68) & (g87) & (g239) & (!g247)) + ((!g68) & (g87) & (g239) & (g247)) + ((g68) & (!g87) & (!g239) & (!g247)) + ((g68) & (!g87) & (!g239) & (g247)) + ((g68) & (!g87) & (g239) & (!g247)) + ((g68) & (g87) & (!g239) & (!g247)));
	assign g265 = (((!g238) & (!g230) & (!g254) & (g264)) + ((!g238) & (g230) & (!g254) & (g264)) + ((!g238) & (g230) & (g254) & (g264)) + ((g238) & (!g230) & (!g254) & (!g264)) + ((g238) & (!g230) & (g254) & (!g264)) + ((g238) & (!g230) & (g254) & (g264)) + ((g238) & (g230) & (!g254) & (!g264)) + ((g238) & (g230) & (g254) & (!g264)));
	assign g266 = (((!g87) & (!g239) & (g247) & (!g230) & (!g254)) + ((!g87) & (!g239) & (g247) & (g230) & (!g254)) + ((!g87) & (!g239) & (g247) & (g230) & (g254)) + ((!g87) & (g239) & (!g247) & (!g230) & (!g254)) + ((!g87) & (g239) & (!g247) & (!g230) & (g254)) + ((!g87) & (g239) & (!g247) & (g230) & (!g254)) + ((!g87) & (g239) & (!g247) & (g230) & (g254)) + ((!g87) & (g239) & (g247) & (!g230) & (g254)) + ((g87) & (!g239) & (!g247) & (!g230) & (!g254)) + ((g87) & (!g239) & (!g247) & (g230) & (!g254)) + ((g87) & (!g239) & (!g247) & (g230) & (g254)) + ((g87) & (g239) & (!g247) & (!g230) & (g254)) + ((g87) & (g239) & (g247) & (!g230) & (!g254)) + ((g87) & (g239) & (g247) & (!g230) & (g254)) + ((g87) & (g239) & (g247) & (g230) & (!g254)) + ((g87) & (g239) & (g247) & (g230) & (g254)));
	assign g267 = (((!g104) & (!g127) & (g241) & (g246)) + ((!g104) & (g127) & (!g241) & (g246)) + ((!g104) & (g127) & (g241) & (!g246)) + ((!g104) & (g127) & (g241) & (g246)) + ((g104) & (!g127) & (!g241) & (!g246)) + ((g104) & (!g127) & (!g241) & (g246)) + ((g104) & (!g127) & (g241) & (!g246)) + ((g104) & (g127) & (!g241) & (!g246)));
	assign g268 = (((!g240) & (!g230) & (!g254) & (g267)) + ((!g240) & (g230) & (!g254) & (g267)) + ((!g240) & (g230) & (g254) & (g267)) + ((g240) & (!g230) & (!g254) & (!g267)) + ((g240) & (!g230) & (g254) & (!g267)) + ((g240) & (!g230) & (g254) & (g267)) + ((g240) & (g230) & (!g254) & (!g267)) + ((g240) & (g230) & (g254) & (!g267)));
	assign g269 = (((!g127) & (!g241) & (g246) & (!g230) & (!g254)) + ((!g127) & (!g241) & (g246) & (g230) & (!g254)) + ((!g127) & (!g241) & (g246) & (g230) & (g254)) + ((!g127) & (g241) & (!g246) & (!g230) & (!g254)) + ((!g127) & (g241) & (!g246) & (!g230) & (g254)) + ((!g127) & (g241) & (!g246) & (g230) & (!g254)) + ((!g127) & (g241) & (!g246) & (g230) & (g254)) + ((!g127) & (g241) & (g246) & (!g230) & (g254)) + ((g127) & (!g241) & (!g246) & (!g230) & (!g254)) + ((g127) & (!g241) & (!g246) & (g230) & (!g254)) + ((g127) & (!g241) & (!g246) & (g230) & (g254)) + ((g127) & (g241) & (!g246) & (!g230) & (g254)) + ((g127) & (g241) & (g246) & (!g230) & (!g254)) + ((g127) & (g241) & (g246) & (!g230) & (g254)) + ((g127) & (g241) & (g246) & (g230) & (!g254)) + ((g127) & (g241) & (g246) & (g230) & (g254)));
	assign g270 = (((!g147) & (!g174) & (g243) & (g245)) + ((!g147) & (g174) & (!g243) & (g245)) + ((!g147) & (g174) & (g243) & (!g245)) + ((!g147) & (g174) & (g243) & (g245)) + ((g147) & (!g174) & (!g243) & (!g245)) + ((g147) & (!g174) & (!g243) & (g245)) + ((g147) & (!g174) & (g243) & (!g245)) + ((g147) & (g174) & (!g243) & (!g245)));
	assign g271 = (((!g242) & (!g230) & (!g254) & (g270)) + ((!g242) & (g230) & (!g254) & (g270)) + ((!g242) & (g230) & (g254) & (g270)) + ((g242) & (!g230) & (!g254) & (!g270)) + ((g242) & (!g230) & (g254) & (!g270)) + ((g242) & (!g230) & (g254) & (g270)) + ((g242) & (g230) & (!g254) & (!g270)) + ((g242) & (g230) & (g254) & (!g270)));
	assign g272 = (((!g174) & (!g243) & (g245) & (!g230) & (!g254)) + ((!g174) & (!g243) & (g245) & (g230) & (!g254)) + ((!g174) & (!g243) & (g245) & (g230) & (g254)) + ((!g174) & (g243) & (!g245) & (!g230) & (!g254)) + ((!g174) & (g243) & (!g245) & (!g230) & (g254)) + ((!g174) & (g243) & (!g245) & (g230) & (!g254)) + ((!g174) & (g243) & (!g245) & (g230) & (g254)) + ((!g174) & (g243) & (g245) & (!g230) & (g254)) + ((g174) & (!g243) & (!g245) & (!g230) & (!g254)) + ((g174) & (!g243) & (!g245) & (g230) & (!g254)) + ((g174) & (!g243) & (!g245) & (g230) & (g254)) + ((g174) & (g243) & (!g245) & (!g230) & (g254)) + ((g174) & (g243) & (g245) & (!g230) & (!g254)) + ((g174) & (g243) & (g245) & (!g230) & (g254)) + ((g174) & (g243) & (g245) & (g230) & (!g254)) + ((g174) & (g243) & (g245) & (g230) & (g254)));
	assign g273 = (((!ax96x) & (!g198) & (!g229) & (!g244)) + ((!ax96x) & (!g198) & (g229) & (!g244)) + ((!ax96x) & (g198) & (!g229) & (g244)) + ((!ax96x) & (g198) & (g229) & (g244)) + ((ax96x) & (!g198) & (g229) & (!g244)) + ((ax96x) & (!g198) & (g229) & (g244)) + ((ax96x) & (g198) & (!g229) & (!g244)) + ((ax96x) & (g198) & (!g229) & (g244)));
	assign g274 = (((!ax96x) & (!ax97x) & (!g229) & (!g230) & (!g254) & (!g273)) + ((!ax96x) & (!ax97x) & (!g229) & (!g230) & (g254) & (!g273)) + ((!ax96x) & (!ax97x) & (!g229) & (!g230) & (g254) & (g273)) + ((!ax96x) & (!ax97x) & (!g229) & (g230) & (!g254) & (!g273)) + ((!ax96x) & (!ax97x) & (!g229) & (g230) & (g254) & (!g273)) + ((!ax96x) & (!ax97x) & (g229) & (!g230) & (!g254) & (g273)) + ((!ax96x) & (!ax97x) & (g229) & (g230) & (!g254) & (g273)) + ((!ax96x) & (!ax97x) & (g229) & (g230) & (g254) & (g273)) + ((!ax96x) & (ax97x) & (!g229) & (!g230) & (!g254) & (g273)) + ((!ax96x) & (ax97x) & (!g229) & (g230) & (!g254) & (g273)) + ((!ax96x) & (ax97x) & (!g229) & (g230) & (g254) & (g273)) + ((!ax96x) & (ax97x) & (g229) & (!g230) & (!g254) & (!g273)) + ((!ax96x) & (ax97x) & (g229) & (!g230) & (g254) & (!g273)) + ((!ax96x) & (ax97x) & (g229) & (!g230) & (g254) & (g273)) + ((!ax96x) & (ax97x) & (g229) & (g230) & (!g254) & (!g273)) + ((!ax96x) & (ax97x) & (g229) & (g230) & (g254) & (!g273)) + ((ax96x) & (!ax97x) & (!g229) & (!g230) & (!g254) & (g273)) + ((ax96x) & (!ax97x) & (!g229) & (g230) & (!g254) & (g273)) + ((ax96x) & (!ax97x) & (!g229) & (g230) & (g254) & (g273)) + ((ax96x) & (!ax97x) & (g229) & (!g230) & (!g254) & (g273)) + ((ax96x) & (!ax97x) & (g229) & (g230) & (!g254) & (g273)) + ((ax96x) & (!ax97x) & (g229) & (g230) & (g254) & (g273)) + ((ax96x) & (ax97x) & (!g229) & (!g230) & (!g254) & (!g273)) + ((ax96x) & (ax97x) & (!g229) & (!g230) & (g254) & (!g273)) + ((ax96x) & (ax97x) & (!g229) & (!g230) & (g254) & (g273)) + ((ax96x) & (ax97x) & (!g229) & (g230) & (!g254) & (!g273)) + ((ax96x) & (ax97x) & (!g229) & (g230) & (g254) & (!g273)) + ((ax96x) & (ax97x) & (g229) & (!g230) & (!g254) & (!g273)) + ((ax96x) & (ax97x) & (g229) & (!g230) & (g254) & (!g273)) + ((ax96x) & (ax97x) & (g229) & (!g230) & (g254) & (g273)) + ((ax96x) & (ax97x) & (g229) & (g230) & (!g254) & (!g273)) + ((ax96x) & (ax97x) & (g229) & (g230) & (g254) & (!g273)));
	assign g275 = (((!ax96x) & (!g229) & (!g244) & (!g230) & (g254)) + ((!ax96x) & (!g229) & (g244) & (!g230) & (!g254)) + ((!ax96x) & (!g229) & (g244) & (!g230) & (g254)) + ((!ax96x) & (!g229) & (g244) & (g230) & (!g254)) + ((!ax96x) & (!g229) & (g244) & (g230) & (g254)) + ((!ax96x) & (g229) & (g244) & (!g230) & (!g254)) + ((!ax96x) & (g229) & (g244) & (g230) & (!g254)) + ((!ax96x) & (g229) & (g244) & (g230) & (g254)) + ((ax96x) & (!g229) & (!g244) & (!g230) & (!g254)) + ((ax96x) & (!g229) & (!g244) & (g230) & (!g254)) + ((ax96x) & (!g229) & (!g244) & (g230) & (g254)) + ((ax96x) & (g229) & (!g244) & (!g230) & (!g254)) + ((ax96x) & (g229) & (!g244) & (!g230) & (g254)) + ((ax96x) & (g229) & (!g244) & (g230) & (!g254)) + ((ax96x) & (g229) & (!g244) & (g230) & (g254)) + ((ax96x) & (g229) & (g244) & (!g230) & (g254)));
	assign g276 = (((!ax92x) & (!ax93x)));
	assign g277 = (((!g229) & (!ax94x) & (!ax95x) & (!g230) & (!g254) & (!g276)) + ((!g229) & (!ax94x) & (!ax95x) & (g230) & (!g254) & (!g276)) + ((!g229) & (!ax94x) & (!ax95x) & (g230) & (g254) & (!g276)) + ((!g229) & (!ax94x) & (ax95x) & (!g230) & (g254) & (!g276)) + ((!g229) & (ax94x) & (ax95x) & (!g230) & (g254) & (!g276)) + ((!g229) & (ax94x) & (ax95x) & (!g230) & (g254) & (g276)) + ((g229) & (!ax94x) & (!ax95x) & (!g230) & (!g254) & (!g276)) + ((g229) & (!ax94x) & (!ax95x) & (!g230) & (!g254) & (g276)) + ((g229) & (!ax94x) & (!ax95x) & (!g230) & (g254) & (!g276)) + ((g229) & (!ax94x) & (!ax95x) & (g230) & (!g254) & (!g276)) + ((g229) & (!ax94x) & (!ax95x) & (g230) & (!g254) & (g276)) + ((g229) & (!ax94x) & (!ax95x) & (g230) & (g254) & (!g276)) + ((g229) & (!ax94x) & (!ax95x) & (g230) & (g254) & (g276)) + ((g229) & (!ax94x) & (ax95x) & (!g230) & (!g254) & (!g276)) + ((g229) & (!ax94x) & (ax95x) & (!g230) & (g254) & (!g276)) + ((g229) & (!ax94x) & (ax95x) & (!g230) & (g254) & (g276)) + ((g229) & (!ax94x) & (ax95x) & (g230) & (!g254) & (!g276)) + ((g229) & (!ax94x) & (ax95x) & (g230) & (g254) & (!g276)) + ((g229) & (ax94x) & (!ax95x) & (!g230) & (g254) & (!g276)) + ((g229) & (ax94x) & (!ax95x) & (!g230) & (g254) & (g276)) + ((g229) & (ax94x) & (ax95x) & (!g230) & (!g254) & (!g276)) + ((g229) & (ax94x) & (ax95x) & (!g230) & (!g254) & (g276)) + ((g229) & (ax94x) & (ax95x) & (!g230) & (g254) & (!g276)) + ((g229) & (ax94x) & (ax95x) & (!g230) & (g254) & (g276)) + ((g229) & (ax94x) & (ax95x) & (g230) & (!g254) & (!g276)) + ((g229) & (ax94x) & (ax95x) & (g230) & (!g254) & (g276)) + ((g229) & (ax94x) & (ax95x) & (g230) & (g254) & (!g276)) + ((g229) & (ax94x) & (ax95x) & (g230) & (g254) & (g276)));
	assign g278 = (((!g174) & (!g198) & (g274) & (g275) & (g277)) + ((!g174) & (g198) & (g274) & (!g275) & (g277)) + ((!g174) & (g198) & (g274) & (g275) & (!g277)) + ((!g174) & (g198) & (g274) & (g275) & (g277)) + ((g174) & (!g198) & (!g274) & (g275) & (g277)) + ((g174) & (!g198) & (g274) & (!g275) & (!g277)) + ((g174) & (!g198) & (g274) & (!g275) & (g277)) + ((g174) & (!g198) & (g274) & (g275) & (!g277)) + ((g174) & (!g198) & (g274) & (g275) & (g277)) + ((g174) & (g198) & (!g274) & (!g275) & (g277)) + ((g174) & (g198) & (!g274) & (g275) & (!g277)) + ((g174) & (g198) & (!g274) & (g275) & (g277)) + ((g174) & (g198) & (g274) & (!g275) & (!g277)) + ((g174) & (g198) & (g274) & (!g275) & (g277)) + ((g174) & (g198) & (g274) & (g275) & (!g277)) + ((g174) & (g198) & (g274) & (g275) & (g277)));
	assign g279 = (((!g127) & (!g147) & (g271) & (g272) & (g278)) + ((!g127) & (g147) & (g271) & (!g272) & (g278)) + ((!g127) & (g147) & (g271) & (g272) & (!g278)) + ((!g127) & (g147) & (g271) & (g272) & (g278)) + ((g127) & (!g147) & (!g271) & (g272) & (g278)) + ((g127) & (!g147) & (g271) & (!g272) & (!g278)) + ((g127) & (!g147) & (g271) & (!g272) & (g278)) + ((g127) & (!g147) & (g271) & (g272) & (!g278)) + ((g127) & (!g147) & (g271) & (g272) & (g278)) + ((g127) & (g147) & (!g271) & (!g272) & (g278)) + ((g127) & (g147) & (!g271) & (g272) & (!g278)) + ((g127) & (g147) & (!g271) & (g272) & (g278)) + ((g127) & (g147) & (g271) & (!g272) & (!g278)) + ((g127) & (g147) & (g271) & (!g272) & (g278)) + ((g127) & (g147) & (g271) & (g272) & (!g278)) + ((g127) & (g147) & (g271) & (g272) & (g278)));
	assign g280 = (((!g87) & (!g104) & (g268) & (g269) & (g279)) + ((!g87) & (g104) & (g268) & (!g269) & (g279)) + ((!g87) & (g104) & (g268) & (g269) & (!g279)) + ((!g87) & (g104) & (g268) & (g269) & (g279)) + ((g87) & (!g104) & (!g268) & (g269) & (g279)) + ((g87) & (!g104) & (g268) & (!g269) & (!g279)) + ((g87) & (!g104) & (g268) & (!g269) & (g279)) + ((g87) & (!g104) & (g268) & (g269) & (!g279)) + ((g87) & (!g104) & (g268) & (g269) & (g279)) + ((g87) & (g104) & (!g268) & (!g269) & (g279)) + ((g87) & (g104) & (!g268) & (g269) & (!g279)) + ((g87) & (g104) & (!g268) & (g269) & (g279)) + ((g87) & (g104) & (g268) & (!g269) & (!g279)) + ((g87) & (g104) & (g268) & (!g269) & (g279)) + ((g87) & (g104) & (g268) & (g269) & (!g279)) + ((g87) & (g104) & (g268) & (g269) & (g279)));
	assign g281 = (((!g54) & (!g68) & (g265) & (g266) & (g280)) + ((!g54) & (g68) & (g265) & (!g266) & (g280)) + ((!g54) & (g68) & (g265) & (g266) & (!g280)) + ((!g54) & (g68) & (g265) & (g266) & (g280)) + ((g54) & (!g68) & (!g265) & (g266) & (g280)) + ((g54) & (!g68) & (g265) & (!g266) & (!g280)) + ((g54) & (!g68) & (g265) & (!g266) & (g280)) + ((g54) & (!g68) & (g265) & (g266) & (!g280)) + ((g54) & (!g68) & (g265) & (g266) & (g280)) + ((g54) & (g68) & (!g265) & (!g266) & (g280)) + ((g54) & (g68) & (!g265) & (g266) & (!g280)) + ((g54) & (g68) & (!g265) & (g266) & (g280)) + ((g54) & (g68) & (g265) & (!g266) & (!g280)) + ((g54) & (g68) & (g265) & (!g266) & (g280)) + ((g54) & (g68) & (g265) & (g266) & (!g280)) + ((g54) & (g68) & (g265) & (g266) & (g280)));
	assign g282 = (((!g27) & (!g39) & (g262) & (g263) & (g281)) + ((!g27) & (g39) & (g262) & (!g263) & (g281)) + ((!g27) & (g39) & (g262) & (g263) & (!g281)) + ((!g27) & (g39) & (g262) & (g263) & (g281)) + ((g27) & (!g39) & (!g262) & (g263) & (g281)) + ((g27) & (!g39) & (g262) & (!g263) & (!g281)) + ((g27) & (!g39) & (g262) & (!g263) & (g281)) + ((g27) & (!g39) & (g262) & (g263) & (!g281)) + ((g27) & (!g39) & (g262) & (g263) & (g281)) + ((g27) & (g39) & (!g262) & (!g263) & (g281)) + ((g27) & (g39) & (!g262) & (g263) & (!g281)) + ((g27) & (g39) & (!g262) & (g263) & (g281)) + ((g27) & (g39) & (g262) & (!g263) & (!g281)) + ((g27) & (g39) & (g262) & (!g263) & (g281)) + ((g27) & (g39) & (g262) & (g263) & (!g281)) + ((g27) & (g39) & (g262) & (g263) & (g281)));
	assign g283 = (((!g8) & (!g18) & (g259) & (g260) & (g282)) + ((!g8) & (g18) & (g259) & (!g260) & (g282)) + ((!g8) & (g18) & (g259) & (g260) & (!g282)) + ((!g8) & (g18) & (g259) & (g260) & (g282)) + ((g8) & (!g18) & (!g259) & (g260) & (g282)) + ((g8) & (!g18) & (g259) & (!g260) & (!g282)) + ((g8) & (!g18) & (g259) & (!g260) & (g282)) + ((g8) & (!g18) & (g259) & (g260) & (!g282)) + ((g8) & (!g18) & (g259) & (g260) & (g282)) + ((g8) & (g18) & (!g259) & (!g260) & (g282)) + ((g8) & (g18) & (!g259) & (g260) & (!g282)) + ((g8) & (g18) & (!g259) & (g260) & (g282)) + ((g8) & (g18) & (g259) & (!g260) & (!g282)) + ((g8) & (g18) & (g259) & (!g260) & (g282)) + ((g8) & (g18) & (g259) & (g260) & (!g282)) + ((g8) & (g18) & (g259) & (g260) & (g282)));
	assign g284 = (((!g2) & (!g8) & (g233) & (g250)) + ((!g2) & (g8) & (!g233) & (g250)) + ((!g2) & (g8) & (g233) & (!g250)) + ((!g2) & (g8) & (g233) & (g250)) + ((g2) & (!g8) & (!g233) & (!g250)) + ((g2) & (!g8) & (!g233) & (g250)) + ((g2) & (!g8) & (g233) & (!g250)) + ((g2) & (g8) & (!g233) & (!g250)));
	assign g285 = (((!g232) & (!g230) & (!g254) & (g284)) + ((!g232) & (g230) & (!g254) & (g284)) + ((!g232) & (g230) & (g254) & (g284)) + ((g232) & (!g230) & (!g254) & (!g284)) + ((g232) & (!g230) & (g254) & (!g284)) + ((g232) & (!g230) & (g254) & (g284)) + ((g232) & (g230) & (!g254) & (!g284)) + ((g232) & (g230) & (g254) & (!g284)));
	assign g286 = (((!g4) & (!g2) & (!g257) & (!g283) & (g285)) + ((!g4) & (!g2) & (!g257) & (g283) & (g285)) + ((!g4) & (!g2) & (g257) & (!g283) & (g285)) + ((!g4) & (!g2) & (g257) & (g283) & (!g285)) + ((!g4) & (!g2) & (g257) & (g283) & (g285)) + ((!g4) & (g2) & (!g257) & (!g283) & (g285)) + ((!g4) & (g2) & (!g257) & (g283) & (!g285)) + ((!g4) & (g2) & (!g257) & (g283) & (g285)) + ((!g4) & (g2) & (g257) & (!g283) & (!g285)) + ((!g4) & (g2) & (g257) & (!g283) & (g285)) + ((!g4) & (g2) & (g257) & (g283) & (!g285)) + ((!g4) & (g2) & (g257) & (g283) & (g285)) + ((g4) & (!g2) & (g257) & (g283) & (g285)) + ((g4) & (g2) & (!g257) & (g283) & (g285)) + ((g4) & (g2) & (g257) & (!g283) & (g285)) + ((g4) & (g2) & (g257) & (g283) & (g285)));
	assign g287 = (((!g4) & (!g251) & (g252)) + ((!g4) & (g251) & (!g252)) + ((!g4) & (g251) & (g252)) + ((g4) & (g251) & (g252)));
	assign g288 = (((!g231) & (!g287) & (!g230) & (!g254)) + ((!g231) & (!g287) & (g230) & (!g254)) + ((!g231) & (!g287) & (g230) & (g254)) + ((g231) & (g287) & (!g230) & (!g254)) + ((g231) & (g287) & (!g230) & (g254)) + ((g231) & (g287) & (g230) & (!g254)) + ((g231) & (g287) & (g230) & (g254)));
	assign g289 = (((!g1) & (g231) & (!g287) & (!g230) & (g254)) + ((!g1) & (g231) & (g287) & (!g230) & (g254)) + ((g1) & (!g231) & (g287) & (g230) & (!g254)) + ((g1) & (!g231) & (g287) & (g230) & (g254)) + ((g1) & (g231) & (!g287) & (!g230) & (!g254)) + ((g1) & (g231) & (!g287) & (!g230) & (g254)) + ((g1) & (g231) & (!g287) & (g230) & (!g254)) + ((g1) & (g231) & (!g287) & (g230) & (g254)) + ((g1) & (g231) & (g287) & (!g230) & (g254)));
	assign g290 = (((!g1) & (!g256) & (!g286) & (!g288) & (!g289)) + ((g1) & (!g256) & (!g286) & (!g288) & (!g289)) + ((g1) & (!g256) & (!g286) & (g288) & (!g289)) + ((g1) & (!g256) & (g286) & (!g288) & (!g289)) + ((g1) & (!g256) & (g286) & (g288) & (!g289)) + ((g1) & (g256) & (!g286) & (!g288) & (!g289)) + ((g1) & (g256) & (!g286) & (g288) & (!g289)));
	assign g291 = (((g1) & (!g256) & (g286) & (g289)) + ((g1) & (g256) & (!g286) & (!g289)) + ((g1) & (g256) & (!g286) & (g289)));
	assign g292 = (((!g4) & (!g2) & (!g257) & (!g283) & (!g285) & (!g290)) + ((!g4) & (!g2) & (!g257) & (!g283) & (g285) & (g290)) + ((!g4) & (!g2) & (!g257) & (g283) & (!g285) & (!g290)) + ((!g4) & (!g2) & (!g257) & (g283) & (g285) & (g290)) + ((!g4) & (!g2) & (g257) & (!g283) & (!g285) & (!g290)) + ((!g4) & (!g2) & (g257) & (!g283) & (g285) & (g290)) + ((!g4) & (!g2) & (g257) & (g283) & (g285) & (!g290)) + ((!g4) & (!g2) & (g257) & (g283) & (g285) & (g290)) + ((!g4) & (g2) & (!g257) & (!g283) & (!g285) & (!g290)) + ((!g4) & (g2) & (!g257) & (!g283) & (g285) & (g290)) + ((!g4) & (g2) & (!g257) & (g283) & (g285) & (!g290)) + ((!g4) & (g2) & (!g257) & (g283) & (g285) & (g290)) + ((!g4) & (g2) & (g257) & (!g283) & (g285) & (!g290)) + ((!g4) & (g2) & (g257) & (!g283) & (g285) & (g290)) + ((!g4) & (g2) & (g257) & (g283) & (g285) & (!g290)) + ((!g4) & (g2) & (g257) & (g283) & (g285) & (g290)) + ((g4) & (!g2) & (!g257) & (!g283) & (g285) & (!g290)) + ((g4) & (!g2) & (!g257) & (!g283) & (g285) & (g290)) + ((g4) & (!g2) & (!g257) & (g283) & (g285) & (!g290)) + ((g4) & (!g2) & (!g257) & (g283) & (g285) & (g290)) + ((g4) & (!g2) & (g257) & (!g283) & (g285) & (!g290)) + ((g4) & (!g2) & (g257) & (!g283) & (g285) & (g290)) + ((g4) & (!g2) & (g257) & (g283) & (!g285) & (!g290)) + ((g4) & (!g2) & (g257) & (g283) & (g285) & (g290)) + ((g4) & (g2) & (!g257) & (!g283) & (g285) & (!g290)) + ((g4) & (g2) & (!g257) & (!g283) & (g285) & (g290)) + ((g4) & (g2) & (!g257) & (g283) & (!g285) & (!g290)) + ((g4) & (g2) & (!g257) & (g283) & (g285) & (g290)) + ((g4) & (g2) & (g257) & (!g283) & (!g285) & (!g290)) + ((g4) & (g2) & (g257) & (!g283) & (g285) & (g290)) + ((g4) & (g2) & (g257) & (g283) & (!g285) & (!g290)) + ((g4) & (g2) & (g257) & (g283) & (g285) & (g290)));
	assign g293 = (((!g8) & (!g18) & (!g259) & (g260) & (g282) & (!g290)) + ((!g8) & (!g18) & (g259) & (!g260) & (!g282) & (!g290)) + ((!g8) & (!g18) & (g259) & (!g260) & (!g282) & (g290)) + ((!g8) & (!g18) & (g259) & (!g260) & (g282) & (!g290)) + ((!g8) & (!g18) & (g259) & (!g260) & (g282) & (g290)) + ((!g8) & (!g18) & (g259) & (g260) & (!g282) & (!g290)) + ((!g8) & (!g18) & (g259) & (g260) & (!g282) & (g290)) + ((!g8) & (!g18) & (g259) & (g260) & (g282) & (g290)) + ((!g8) & (g18) & (!g259) & (!g260) & (g282) & (!g290)) + ((!g8) & (g18) & (!g259) & (g260) & (!g282) & (!g290)) + ((!g8) & (g18) & (!g259) & (g260) & (g282) & (!g290)) + ((!g8) & (g18) & (g259) & (!g260) & (!g282) & (!g290)) + ((!g8) & (g18) & (g259) & (!g260) & (!g282) & (g290)) + ((!g8) & (g18) & (g259) & (!g260) & (g282) & (g290)) + ((!g8) & (g18) & (g259) & (g260) & (!g282) & (g290)) + ((!g8) & (g18) & (g259) & (g260) & (g282) & (g290)) + ((g8) & (!g18) & (!g259) & (!g260) & (!g282) & (!g290)) + ((g8) & (!g18) & (!g259) & (!g260) & (g282) & (!g290)) + ((g8) & (!g18) & (!g259) & (g260) & (!g282) & (!g290)) + ((g8) & (!g18) & (g259) & (!g260) & (!g282) & (g290)) + ((g8) & (!g18) & (g259) & (!g260) & (g282) & (g290)) + ((g8) & (!g18) & (g259) & (g260) & (!g282) & (g290)) + ((g8) & (!g18) & (g259) & (g260) & (g282) & (!g290)) + ((g8) & (!g18) & (g259) & (g260) & (g282) & (g290)) + ((g8) & (g18) & (!g259) & (!g260) & (!g282) & (!g290)) + ((g8) & (g18) & (g259) & (!g260) & (!g282) & (g290)) + ((g8) & (g18) & (g259) & (!g260) & (g282) & (!g290)) + ((g8) & (g18) & (g259) & (!g260) & (g282) & (g290)) + ((g8) & (g18) & (g259) & (g260) & (!g282) & (!g290)) + ((g8) & (g18) & (g259) & (g260) & (!g282) & (g290)) + ((g8) & (g18) & (g259) & (g260) & (g282) & (!g290)) + ((g8) & (g18) & (g259) & (g260) & (g282) & (g290)));
	assign g294 = (((!g18) & (!g260) & (g282) & (!g290)) + ((!g18) & (g260) & (!g282) & (!g290)) + ((!g18) & (g260) & (!g282) & (g290)) + ((!g18) & (g260) & (g282) & (g290)) + ((g18) & (!g260) & (!g282) & (!g290)) + ((g18) & (g260) & (!g282) & (g290)) + ((g18) & (g260) & (g282) & (!g290)) + ((g18) & (g260) & (g282) & (g290)));
	assign g295 = (((!g27) & (!g39) & (!g262) & (g263) & (g281) & (!g290)) + ((!g27) & (!g39) & (g262) & (!g263) & (!g281) & (!g290)) + ((!g27) & (!g39) & (g262) & (!g263) & (!g281) & (g290)) + ((!g27) & (!g39) & (g262) & (!g263) & (g281) & (!g290)) + ((!g27) & (!g39) & (g262) & (!g263) & (g281) & (g290)) + ((!g27) & (!g39) & (g262) & (g263) & (!g281) & (!g290)) + ((!g27) & (!g39) & (g262) & (g263) & (!g281) & (g290)) + ((!g27) & (!g39) & (g262) & (g263) & (g281) & (g290)) + ((!g27) & (g39) & (!g262) & (!g263) & (g281) & (!g290)) + ((!g27) & (g39) & (!g262) & (g263) & (!g281) & (!g290)) + ((!g27) & (g39) & (!g262) & (g263) & (g281) & (!g290)) + ((!g27) & (g39) & (g262) & (!g263) & (!g281) & (!g290)) + ((!g27) & (g39) & (g262) & (!g263) & (!g281) & (g290)) + ((!g27) & (g39) & (g262) & (!g263) & (g281) & (g290)) + ((!g27) & (g39) & (g262) & (g263) & (!g281) & (g290)) + ((!g27) & (g39) & (g262) & (g263) & (g281) & (g290)) + ((g27) & (!g39) & (!g262) & (!g263) & (!g281) & (!g290)) + ((g27) & (!g39) & (!g262) & (!g263) & (g281) & (!g290)) + ((g27) & (!g39) & (!g262) & (g263) & (!g281) & (!g290)) + ((g27) & (!g39) & (g262) & (!g263) & (!g281) & (g290)) + ((g27) & (!g39) & (g262) & (!g263) & (g281) & (g290)) + ((g27) & (!g39) & (g262) & (g263) & (!g281) & (g290)) + ((g27) & (!g39) & (g262) & (g263) & (g281) & (!g290)) + ((g27) & (!g39) & (g262) & (g263) & (g281) & (g290)) + ((g27) & (g39) & (!g262) & (!g263) & (!g281) & (!g290)) + ((g27) & (g39) & (g262) & (!g263) & (!g281) & (g290)) + ((g27) & (g39) & (g262) & (!g263) & (g281) & (!g290)) + ((g27) & (g39) & (g262) & (!g263) & (g281) & (g290)) + ((g27) & (g39) & (g262) & (g263) & (!g281) & (!g290)) + ((g27) & (g39) & (g262) & (g263) & (!g281) & (g290)) + ((g27) & (g39) & (g262) & (g263) & (g281) & (!g290)) + ((g27) & (g39) & (g262) & (g263) & (g281) & (g290)));
	assign g296 = (((!g39) & (!g263) & (g281) & (!g290)) + ((!g39) & (g263) & (!g281) & (!g290)) + ((!g39) & (g263) & (!g281) & (g290)) + ((!g39) & (g263) & (g281) & (g290)) + ((g39) & (!g263) & (!g281) & (!g290)) + ((g39) & (g263) & (!g281) & (g290)) + ((g39) & (g263) & (g281) & (!g290)) + ((g39) & (g263) & (g281) & (g290)));
	assign g297 = (((!g54) & (!g68) & (!g265) & (g266) & (g280) & (!g290)) + ((!g54) & (!g68) & (g265) & (!g266) & (!g280) & (!g290)) + ((!g54) & (!g68) & (g265) & (!g266) & (!g280) & (g290)) + ((!g54) & (!g68) & (g265) & (!g266) & (g280) & (!g290)) + ((!g54) & (!g68) & (g265) & (!g266) & (g280) & (g290)) + ((!g54) & (!g68) & (g265) & (g266) & (!g280) & (!g290)) + ((!g54) & (!g68) & (g265) & (g266) & (!g280) & (g290)) + ((!g54) & (!g68) & (g265) & (g266) & (g280) & (g290)) + ((!g54) & (g68) & (!g265) & (!g266) & (g280) & (!g290)) + ((!g54) & (g68) & (!g265) & (g266) & (!g280) & (!g290)) + ((!g54) & (g68) & (!g265) & (g266) & (g280) & (!g290)) + ((!g54) & (g68) & (g265) & (!g266) & (!g280) & (!g290)) + ((!g54) & (g68) & (g265) & (!g266) & (!g280) & (g290)) + ((!g54) & (g68) & (g265) & (!g266) & (g280) & (g290)) + ((!g54) & (g68) & (g265) & (g266) & (!g280) & (g290)) + ((!g54) & (g68) & (g265) & (g266) & (g280) & (g290)) + ((g54) & (!g68) & (!g265) & (!g266) & (!g280) & (!g290)) + ((g54) & (!g68) & (!g265) & (!g266) & (g280) & (!g290)) + ((g54) & (!g68) & (!g265) & (g266) & (!g280) & (!g290)) + ((g54) & (!g68) & (g265) & (!g266) & (!g280) & (g290)) + ((g54) & (!g68) & (g265) & (!g266) & (g280) & (g290)) + ((g54) & (!g68) & (g265) & (g266) & (!g280) & (g290)) + ((g54) & (!g68) & (g265) & (g266) & (g280) & (!g290)) + ((g54) & (!g68) & (g265) & (g266) & (g280) & (g290)) + ((g54) & (g68) & (!g265) & (!g266) & (!g280) & (!g290)) + ((g54) & (g68) & (g265) & (!g266) & (!g280) & (g290)) + ((g54) & (g68) & (g265) & (!g266) & (g280) & (!g290)) + ((g54) & (g68) & (g265) & (!g266) & (g280) & (g290)) + ((g54) & (g68) & (g265) & (g266) & (!g280) & (!g290)) + ((g54) & (g68) & (g265) & (g266) & (!g280) & (g290)) + ((g54) & (g68) & (g265) & (g266) & (g280) & (!g290)) + ((g54) & (g68) & (g265) & (g266) & (g280) & (g290)));
	assign g298 = (((!g68) & (!g266) & (g280) & (!g290)) + ((!g68) & (g266) & (!g280) & (!g290)) + ((!g68) & (g266) & (!g280) & (g290)) + ((!g68) & (g266) & (g280) & (g290)) + ((g68) & (!g266) & (!g280) & (!g290)) + ((g68) & (g266) & (!g280) & (g290)) + ((g68) & (g266) & (g280) & (!g290)) + ((g68) & (g266) & (g280) & (g290)));
	assign g299 = (((!g87) & (!g104) & (!g268) & (g269) & (g279) & (!g290)) + ((!g87) & (!g104) & (g268) & (!g269) & (!g279) & (!g290)) + ((!g87) & (!g104) & (g268) & (!g269) & (!g279) & (g290)) + ((!g87) & (!g104) & (g268) & (!g269) & (g279) & (!g290)) + ((!g87) & (!g104) & (g268) & (!g269) & (g279) & (g290)) + ((!g87) & (!g104) & (g268) & (g269) & (!g279) & (!g290)) + ((!g87) & (!g104) & (g268) & (g269) & (!g279) & (g290)) + ((!g87) & (!g104) & (g268) & (g269) & (g279) & (g290)) + ((!g87) & (g104) & (!g268) & (!g269) & (g279) & (!g290)) + ((!g87) & (g104) & (!g268) & (g269) & (!g279) & (!g290)) + ((!g87) & (g104) & (!g268) & (g269) & (g279) & (!g290)) + ((!g87) & (g104) & (g268) & (!g269) & (!g279) & (!g290)) + ((!g87) & (g104) & (g268) & (!g269) & (!g279) & (g290)) + ((!g87) & (g104) & (g268) & (!g269) & (g279) & (g290)) + ((!g87) & (g104) & (g268) & (g269) & (!g279) & (g290)) + ((!g87) & (g104) & (g268) & (g269) & (g279) & (g290)) + ((g87) & (!g104) & (!g268) & (!g269) & (!g279) & (!g290)) + ((g87) & (!g104) & (!g268) & (!g269) & (g279) & (!g290)) + ((g87) & (!g104) & (!g268) & (g269) & (!g279) & (!g290)) + ((g87) & (!g104) & (g268) & (!g269) & (!g279) & (g290)) + ((g87) & (!g104) & (g268) & (!g269) & (g279) & (g290)) + ((g87) & (!g104) & (g268) & (g269) & (!g279) & (g290)) + ((g87) & (!g104) & (g268) & (g269) & (g279) & (!g290)) + ((g87) & (!g104) & (g268) & (g269) & (g279) & (g290)) + ((g87) & (g104) & (!g268) & (!g269) & (!g279) & (!g290)) + ((g87) & (g104) & (g268) & (!g269) & (!g279) & (g290)) + ((g87) & (g104) & (g268) & (!g269) & (g279) & (!g290)) + ((g87) & (g104) & (g268) & (!g269) & (g279) & (g290)) + ((g87) & (g104) & (g268) & (g269) & (!g279) & (!g290)) + ((g87) & (g104) & (g268) & (g269) & (!g279) & (g290)) + ((g87) & (g104) & (g268) & (g269) & (g279) & (!g290)) + ((g87) & (g104) & (g268) & (g269) & (g279) & (g290)));
	assign g300 = (((!g104) & (!g269) & (g279) & (!g290)) + ((!g104) & (g269) & (!g279) & (!g290)) + ((!g104) & (g269) & (!g279) & (g290)) + ((!g104) & (g269) & (g279) & (g290)) + ((g104) & (!g269) & (!g279) & (!g290)) + ((g104) & (g269) & (!g279) & (g290)) + ((g104) & (g269) & (g279) & (!g290)) + ((g104) & (g269) & (g279) & (g290)));
	assign g301 = (((!g127) & (!g147) & (!g271) & (g272) & (g278) & (!g290)) + ((!g127) & (!g147) & (g271) & (!g272) & (!g278) & (!g290)) + ((!g127) & (!g147) & (g271) & (!g272) & (!g278) & (g290)) + ((!g127) & (!g147) & (g271) & (!g272) & (g278) & (!g290)) + ((!g127) & (!g147) & (g271) & (!g272) & (g278) & (g290)) + ((!g127) & (!g147) & (g271) & (g272) & (!g278) & (!g290)) + ((!g127) & (!g147) & (g271) & (g272) & (!g278) & (g290)) + ((!g127) & (!g147) & (g271) & (g272) & (g278) & (g290)) + ((!g127) & (g147) & (!g271) & (!g272) & (g278) & (!g290)) + ((!g127) & (g147) & (!g271) & (g272) & (!g278) & (!g290)) + ((!g127) & (g147) & (!g271) & (g272) & (g278) & (!g290)) + ((!g127) & (g147) & (g271) & (!g272) & (!g278) & (!g290)) + ((!g127) & (g147) & (g271) & (!g272) & (!g278) & (g290)) + ((!g127) & (g147) & (g271) & (!g272) & (g278) & (g290)) + ((!g127) & (g147) & (g271) & (g272) & (!g278) & (g290)) + ((!g127) & (g147) & (g271) & (g272) & (g278) & (g290)) + ((g127) & (!g147) & (!g271) & (!g272) & (!g278) & (!g290)) + ((g127) & (!g147) & (!g271) & (!g272) & (g278) & (!g290)) + ((g127) & (!g147) & (!g271) & (g272) & (!g278) & (!g290)) + ((g127) & (!g147) & (g271) & (!g272) & (!g278) & (g290)) + ((g127) & (!g147) & (g271) & (!g272) & (g278) & (g290)) + ((g127) & (!g147) & (g271) & (g272) & (!g278) & (g290)) + ((g127) & (!g147) & (g271) & (g272) & (g278) & (!g290)) + ((g127) & (!g147) & (g271) & (g272) & (g278) & (g290)) + ((g127) & (g147) & (!g271) & (!g272) & (!g278) & (!g290)) + ((g127) & (g147) & (g271) & (!g272) & (!g278) & (g290)) + ((g127) & (g147) & (g271) & (!g272) & (g278) & (!g290)) + ((g127) & (g147) & (g271) & (!g272) & (g278) & (g290)) + ((g127) & (g147) & (g271) & (g272) & (!g278) & (!g290)) + ((g127) & (g147) & (g271) & (g272) & (!g278) & (g290)) + ((g127) & (g147) & (g271) & (g272) & (g278) & (!g290)) + ((g127) & (g147) & (g271) & (g272) & (g278) & (g290)));
	assign g302 = (((!g147) & (!g272) & (g278) & (!g290)) + ((!g147) & (g272) & (!g278) & (!g290)) + ((!g147) & (g272) & (!g278) & (g290)) + ((!g147) & (g272) & (g278) & (g290)) + ((g147) & (!g272) & (!g278) & (!g290)) + ((g147) & (g272) & (!g278) & (g290)) + ((g147) & (g272) & (g278) & (!g290)) + ((g147) & (g272) & (g278) & (g290)));
	assign g303 = (((!g174) & (!g198) & (!g274) & (g275) & (g277) & (!g290)) + ((!g174) & (!g198) & (g274) & (!g275) & (!g277) & (!g290)) + ((!g174) & (!g198) & (g274) & (!g275) & (!g277) & (g290)) + ((!g174) & (!g198) & (g274) & (!g275) & (g277) & (!g290)) + ((!g174) & (!g198) & (g274) & (!g275) & (g277) & (g290)) + ((!g174) & (!g198) & (g274) & (g275) & (!g277) & (!g290)) + ((!g174) & (!g198) & (g274) & (g275) & (!g277) & (g290)) + ((!g174) & (!g198) & (g274) & (g275) & (g277) & (g290)) + ((!g174) & (g198) & (!g274) & (!g275) & (g277) & (!g290)) + ((!g174) & (g198) & (!g274) & (g275) & (!g277) & (!g290)) + ((!g174) & (g198) & (!g274) & (g275) & (g277) & (!g290)) + ((!g174) & (g198) & (g274) & (!g275) & (!g277) & (!g290)) + ((!g174) & (g198) & (g274) & (!g275) & (!g277) & (g290)) + ((!g174) & (g198) & (g274) & (!g275) & (g277) & (g290)) + ((!g174) & (g198) & (g274) & (g275) & (!g277) & (g290)) + ((!g174) & (g198) & (g274) & (g275) & (g277) & (g290)) + ((g174) & (!g198) & (!g274) & (!g275) & (!g277) & (!g290)) + ((g174) & (!g198) & (!g274) & (!g275) & (g277) & (!g290)) + ((g174) & (!g198) & (!g274) & (g275) & (!g277) & (!g290)) + ((g174) & (!g198) & (g274) & (!g275) & (!g277) & (g290)) + ((g174) & (!g198) & (g274) & (!g275) & (g277) & (g290)) + ((g174) & (!g198) & (g274) & (g275) & (!g277) & (g290)) + ((g174) & (!g198) & (g274) & (g275) & (g277) & (!g290)) + ((g174) & (!g198) & (g274) & (g275) & (g277) & (g290)) + ((g174) & (g198) & (!g274) & (!g275) & (!g277) & (!g290)) + ((g174) & (g198) & (g274) & (!g275) & (!g277) & (g290)) + ((g174) & (g198) & (g274) & (!g275) & (g277) & (!g290)) + ((g174) & (g198) & (g274) & (!g275) & (g277) & (g290)) + ((g174) & (g198) & (g274) & (g275) & (!g277) & (!g290)) + ((g174) & (g198) & (g274) & (g275) & (!g277) & (g290)) + ((g174) & (g198) & (g274) & (g275) & (g277) & (!g290)) + ((g174) & (g198) & (g274) & (g275) & (g277) & (g290)));
	assign g304 = (((!g198) & (!g275) & (g277) & (!g290)) + ((!g198) & (g275) & (!g277) & (!g290)) + ((!g198) & (g275) & (!g277) & (g290)) + ((!g198) & (g275) & (g277) & (g290)) + ((g198) & (!g275) & (!g277) & (!g290)) + ((g198) & (g275) & (!g277) & (g290)) + ((g198) & (g275) & (g277) & (!g290)) + ((g198) & (g275) & (g277) & (g290)));
	assign g305 = (((!g229) & (!ax94x) & (!ax95x) & (!g255) & (!g276) & (g290)) + ((!g229) & (!ax94x) & (!ax95x) & (!g255) & (g276) & (!g290)) + ((!g229) & (!ax94x) & (!ax95x) & (!g255) & (g276) & (g290)) + ((!g229) & (!ax94x) & (!ax95x) & (g255) & (!g276) & (!g290)) + ((!g229) & (!ax94x) & (ax95x) & (!g255) & (!g276) & (!g290)) + ((!g229) & (!ax94x) & (ax95x) & (g255) & (!g276) & (g290)) + ((!g229) & (!ax94x) & (ax95x) & (g255) & (g276) & (!g290)) + ((!g229) & (!ax94x) & (ax95x) & (g255) & (g276) & (g290)) + ((!g229) & (ax94x) & (!ax95x) & (g255) & (!g276) & (!g290)) + ((!g229) & (ax94x) & (!ax95x) & (g255) & (g276) & (!g290)) + ((!g229) & (ax94x) & (ax95x) & (!g255) & (!g276) & (!g290)) + ((!g229) & (ax94x) & (ax95x) & (!g255) & (!g276) & (g290)) + ((!g229) & (ax94x) & (ax95x) & (!g255) & (g276) & (!g290)) + ((!g229) & (ax94x) & (ax95x) & (!g255) & (g276) & (g290)) + ((!g229) & (ax94x) & (ax95x) & (g255) & (!g276) & (g290)) + ((!g229) & (ax94x) & (ax95x) & (g255) & (g276) & (g290)) + ((g229) & (!ax94x) & (!ax95x) & (!g255) & (!g276) & (!g290)) + ((g229) & (!ax94x) & (!ax95x) & (!g255) & (!g276) & (g290)) + ((g229) & (!ax94x) & (!ax95x) & (!g255) & (g276) & (g290)) + ((g229) & (!ax94x) & (!ax95x) & (g255) & (g276) & (!g290)) + ((g229) & (!ax94x) & (ax95x) & (!g255) & (g276) & (!g290)) + ((g229) & (!ax94x) & (ax95x) & (g255) & (!g276) & (!g290)) + ((g229) & (!ax94x) & (ax95x) & (g255) & (!g276) & (g290)) + ((g229) & (!ax94x) & (ax95x) & (g255) & (g276) & (g290)) + ((g229) & (ax94x) & (!ax95x) & (!g255) & (!g276) & (!g290)) + ((g229) & (ax94x) & (!ax95x) & (!g255) & (g276) & (!g290)) + ((g229) & (ax94x) & (ax95x) & (!g255) & (!g276) & (g290)) + ((g229) & (ax94x) & (ax95x) & (!g255) & (g276) & (g290)) + ((g229) & (ax94x) & (ax95x) & (g255) & (!g276) & (!g290)) + ((g229) & (ax94x) & (ax95x) & (g255) & (!g276) & (g290)) + ((g229) & (ax94x) & (ax95x) & (g255) & (g276) & (!g290)) + ((g229) & (ax94x) & (ax95x) & (g255) & (g276) & (g290)));
	assign g306 = (((!ax94x) & (!g255) & (!g276) & (g290)) + ((!ax94x) & (!g255) & (g276) & (!g290)) + ((!ax94x) & (!g255) & (g276) & (g290)) + ((!ax94x) & (g255) & (g276) & (!g290)) + ((ax94x) & (!g255) & (!g276) & (!g290)) + ((ax94x) & (g255) & (!g276) & (!g290)) + ((ax94x) & (g255) & (!g276) & (g290)) + ((ax94x) & (g255) & (g276) & (g290)));
	assign g307 = (((!ax90x) & (!ax91x)));
	assign g308 = (((!g255) & (!ax92x) & (!ax93x) & (!g290) & (!g307)) + ((!g255) & (!ax92x) & (ax93x) & (g290) & (!g307)) + ((!g255) & (ax92x) & (ax93x) & (g290) & (!g307)) + ((!g255) & (ax92x) & (ax93x) & (g290) & (g307)) + ((g255) & (!ax92x) & (!ax93x) & (!g290) & (!g307)) + ((g255) & (!ax92x) & (!ax93x) & (!g290) & (g307)) + ((g255) & (!ax92x) & (!ax93x) & (g290) & (!g307)) + ((g255) & (!ax92x) & (ax93x) & (!g290) & (!g307)) + ((g255) & (!ax92x) & (ax93x) & (g290) & (!g307)) + ((g255) & (!ax92x) & (ax93x) & (g290) & (g307)) + ((g255) & (ax92x) & (!ax93x) & (g290) & (!g307)) + ((g255) & (ax92x) & (!ax93x) & (g290) & (g307)) + ((g255) & (ax92x) & (ax93x) & (!g290) & (!g307)) + ((g255) & (ax92x) & (ax93x) & (!g290) & (g307)) + ((g255) & (ax92x) & (ax93x) & (g290) & (!g307)) + ((g255) & (ax92x) & (ax93x) & (g290) & (g307)));
	assign g309 = (((!g198) & (!g229) & (g305) & (g306) & (g308)) + ((!g198) & (g229) & (g305) & (!g306) & (g308)) + ((!g198) & (g229) & (g305) & (g306) & (!g308)) + ((!g198) & (g229) & (g305) & (g306) & (g308)) + ((g198) & (!g229) & (!g305) & (g306) & (g308)) + ((g198) & (!g229) & (g305) & (!g306) & (!g308)) + ((g198) & (!g229) & (g305) & (!g306) & (g308)) + ((g198) & (!g229) & (g305) & (g306) & (!g308)) + ((g198) & (!g229) & (g305) & (g306) & (g308)) + ((g198) & (g229) & (!g305) & (!g306) & (g308)) + ((g198) & (g229) & (!g305) & (g306) & (!g308)) + ((g198) & (g229) & (!g305) & (g306) & (g308)) + ((g198) & (g229) & (g305) & (!g306) & (!g308)) + ((g198) & (g229) & (g305) & (!g306) & (g308)) + ((g198) & (g229) & (g305) & (g306) & (!g308)) + ((g198) & (g229) & (g305) & (g306) & (g308)));
	assign g310 = (((!g147) & (!g174) & (g303) & (g304) & (g309)) + ((!g147) & (g174) & (g303) & (!g304) & (g309)) + ((!g147) & (g174) & (g303) & (g304) & (!g309)) + ((!g147) & (g174) & (g303) & (g304) & (g309)) + ((g147) & (!g174) & (!g303) & (g304) & (g309)) + ((g147) & (!g174) & (g303) & (!g304) & (!g309)) + ((g147) & (!g174) & (g303) & (!g304) & (g309)) + ((g147) & (!g174) & (g303) & (g304) & (!g309)) + ((g147) & (!g174) & (g303) & (g304) & (g309)) + ((g147) & (g174) & (!g303) & (!g304) & (g309)) + ((g147) & (g174) & (!g303) & (g304) & (!g309)) + ((g147) & (g174) & (!g303) & (g304) & (g309)) + ((g147) & (g174) & (g303) & (!g304) & (!g309)) + ((g147) & (g174) & (g303) & (!g304) & (g309)) + ((g147) & (g174) & (g303) & (g304) & (!g309)) + ((g147) & (g174) & (g303) & (g304) & (g309)));
	assign g311 = (((!g104) & (!g127) & (g301) & (g302) & (g310)) + ((!g104) & (g127) & (g301) & (!g302) & (g310)) + ((!g104) & (g127) & (g301) & (g302) & (!g310)) + ((!g104) & (g127) & (g301) & (g302) & (g310)) + ((g104) & (!g127) & (!g301) & (g302) & (g310)) + ((g104) & (!g127) & (g301) & (!g302) & (!g310)) + ((g104) & (!g127) & (g301) & (!g302) & (g310)) + ((g104) & (!g127) & (g301) & (g302) & (!g310)) + ((g104) & (!g127) & (g301) & (g302) & (g310)) + ((g104) & (g127) & (!g301) & (!g302) & (g310)) + ((g104) & (g127) & (!g301) & (g302) & (!g310)) + ((g104) & (g127) & (!g301) & (g302) & (g310)) + ((g104) & (g127) & (g301) & (!g302) & (!g310)) + ((g104) & (g127) & (g301) & (!g302) & (g310)) + ((g104) & (g127) & (g301) & (g302) & (!g310)) + ((g104) & (g127) & (g301) & (g302) & (g310)));
	assign g312 = (((!g68) & (!g87) & (g299) & (g300) & (g311)) + ((!g68) & (g87) & (g299) & (!g300) & (g311)) + ((!g68) & (g87) & (g299) & (g300) & (!g311)) + ((!g68) & (g87) & (g299) & (g300) & (g311)) + ((g68) & (!g87) & (!g299) & (g300) & (g311)) + ((g68) & (!g87) & (g299) & (!g300) & (!g311)) + ((g68) & (!g87) & (g299) & (!g300) & (g311)) + ((g68) & (!g87) & (g299) & (g300) & (!g311)) + ((g68) & (!g87) & (g299) & (g300) & (g311)) + ((g68) & (g87) & (!g299) & (!g300) & (g311)) + ((g68) & (g87) & (!g299) & (g300) & (!g311)) + ((g68) & (g87) & (!g299) & (g300) & (g311)) + ((g68) & (g87) & (g299) & (!g300) & (!g311)) + ((g68) & (g87) & (g299) & (!g300) & (g311)) + ((g68) & (g87) & (g299) & (g300) & (!g311)) + ((g68) & (g87) & (g299) & (g300) & (g311)));
	assign g313 = (((!g39) & (!g54) & (g297) & (g298) & (g312)) + ((!g39) & (g54) & (g297) & (!g298) & (g312)) + ((!g39) & (g54) & (g297) & (g298) & (!g312)) + ((!g39) & (g54) & (g297) & (g298) & (g312)) + ((g39) & (!g54) & (!g297) & (g298) & (g312)) + ((g39) & (!g54) & (g297) & (!g298) & (!g312)) + ((g39) & (!g54) & (g297) & (!g298) & (g312)) + ((g39) & (!g54) & (g297) & (g298) & (!g312)) + ((g39) & (!g54) & (g297) & (g298) & (g312)) + ((g39) & (g54) & (!g297) & (!g298) & (g312)) + ((g39) & (g54) & (!g297) & (g298) & (!g312)) + ((g39) & (g54) & (!g297) & (g298) & (g312)) + ((g39) & (g54) & (g297) & (!g298) & (!g312)) + ((g39) & (g54) & (g297) & (!g298) & (g312)) + ((g39) & (g54) & (g297) & (g298) & (!g312)) + ((g39) & (g54) & (g297) & (g298) & (g312)));
	assign g314 = (((!g18) & (!g27) & (g295) & (g296) & (g313)) + ((!g18) & (g27) & (g295) & (!g296) & (g313)) + ((!g18) & (g27) & (g295) & (g296) & (!g313)) + ((!g18) & (g27) & (g295) & (g296) & (g313)) + ((g18) & (!g27) & (!g295) & (g296) & (g313)) + ((g18) & (!g27) & (g295) & (!g296) & (!g313)) + ((g18) & (!g27) & (g295) & (!g296) & (g313)) + ((g18) & (!g27) & (g295) & (g296) & (!g313)) + ((g18) & (!g27) & (g295) & (g296) & (g313)) + ((g18) & (g27) & (!g295) & (!g296) & (g313)) + ((g18) & (g27) & (!g295) & (g296) & (!g313)) + ((g18) & (g27) & (!g295) & (g296) & (g313)) + ((g18) & (g27) & (g295) & (!g296) & (!g313)) + ((g18) & (g27) & (g295) & (!g296) & (g313)) + ((g18) & (g27) & (g295) & (g296) & (!g313)) + ((g18) & (g27) & (g295) & (g296) & (g313)));
	assign g315 = (((!g2) & (!g8) & (g293) & (g294) & (g314)) + ((!g2) & (g8) & (g293) & (!g294) & (g314)) + ((!g2) & (g8) & (g293) & (g294) & (!g314)) + ((!g2) & (g8) & (g293) & (g294) & (g314)) + ((g2) & (!g8) & (!g293) & (g294) & (g314)) + ((g2) & (!g8) & (g293) & (!g294) & (!g314)) + ((g2) & (!g8) & (g293) & (!g294) & (g314)) + ((g2) & (!g8) & (g293) & (g294) & (!g314)) + ((g2) & (!g8) & (g293) & (g294) & (g314)) + ((g2) & (g8) & (!g293) & (!g294) & (g314)) + ((g2) & (g8) & (!g293) & (g294) & (!g314)) + ((g2) & (g8) & (!g293) & (g294) & (g314)) + ((g2) & (g8) & (g293) & (!g294) & (!g314)) + ((g2) & (g8) & (g293) & (!g294) & (g314)) + ((g2) & (g8) & (g293) & (g294) & (!g314)) + ((g2) & (g8) & (g293) & (g294) & (g314)));
	assign g316 = (((!g2) & (!g257) & (g283) & (!g290)) + ((!g2) & (g257) & (!g283) & (!g290)) + ((!g2) & (g257) & (!g283) & (g290)) + ((!g2) & (g257) & (g283) & (g290)) + ((g2) & (!g257) & (!g283) & (!g290)) + ((g2) & (g257) & (!g283) & (g290)) + ((g2) & (g257) & (g283) & (!g290)) + ((g2) & (g257) & (g283) & (g290)));
	assign g317 = (((!g1) & (!g256) & (!g286) & (!g288) & (g289)) + ((!g1) & (!g256) & (!g286) & (g288) & (!g289)) + ((!g1) & (!g256) & (!g286) & (g288) & (g289)) + ((!g1) & (g256) & (g286) & (!g288) & (!g289)) + ((!g1) & (g256) & (g286) & (!g288) & (g289)) + ((!g1) & (g256) & (g286) & (g288) & (!g289)) + ((!g1) & (g256) & (g286) & (g288) & (g289)) + ((g1) & (!g256) & (!g286) & (!g288) & (g289)) + ((g1) & (!g256) & (!g286) & (g288) & (g289)) + ((g1) & (g256) & (g286) & (!g288) & (!g289)) + ((g1) & (g256) & (g286) & (!g288) & (g289)) + ((g1) & (g256) & (g286) & (g288) & (!g289)) + ((g1) & (g256) & (g286) & (g288) & (g289)));
	assign g318 = (((!g4) & (!g1) & (!g292) & (!g315) & (!g316) & (!g317)) + ((!g4) & (g1) & (!g292) & (!g315) & (!g316) & (!g317)) + ((!g4) & (g1) & (!g292) & (!g315) & (!g316) & (g317)) + ((!g4) & (g1) & (!g292) & (!g315) & (g316) & (!g317)) + ((!g4) & (g1) & (!g292) & (!g315) & (g316) & (g317)) + ((!g4) & (g1) & (!g292) & (g315) & (!g316) & (!g317)) + ((!g4) & (g1) & (!g292) & (g315) & (!g316) & (g317)) + ((!g4) & (g1) & (!g292) & (g315) & (g316) & (!g317)) + ((!g4) & (g1) & (!g292) & (g315) & (g316) & (g317)) + ((!g4) & (g1) & (g292) & (!g315) & (!g316) & (!g317)) + ((!g4) & (g1) & (g292) & (!g315) & (!g316) & (g317)) + ((g4) & (!g1) & (!g292) & (!g315) & (!g316) & (!g317)) + ((g4) & (!g1) & (!g292) & (!g315) & (g316) & (!g317)) + ((g4) & (!g1) & (!g292) & (g315) & (!g316) & (!g317)) + ((g4) & (g1) & (!g292) & (!g315) & (!g316) & (!g317)) + ((g4) & (g1) & (!g292) & (!g315) & (!g316) & (g317)) + ((g4) & (g1) & (!g292) & (!g315) & (g316) & (!g317)) + ((g4) & (g1) & (!g292) & (!g315) & (g316) & (g317)) + ((g4) & (g1) & (!g292) & (g315) & (!g316) & (!g317)) + ((g4) & (g1) & (!g292) & (g315) & (!g316) & (g317)) + ((g4) & (g1) & (!g292) & (g315) & (g316) & (!g317)) + ((g4) & (g1) & (!g292) & (g315) & (g316) & (g317)) + ((g4) & (g1) & (g292) & (!g315) & (!g316) & (!g317)) + ((g4) & (g1) & (g292) & (!g315) & (!g316) & (g317)) + ((g4) & (g1) & (g292) & (!g315) & (g316) & (!g317)) + ((g4) & (g1) & (g292) & (!g315) & (g316) & (g317)) + ((g4) & (g1) & (g292) & (g315) & (!g316) & (!g317)) + ((g4) & (g1) & (g292) & (g315) & (!g316) & (g317)));
	assign g319 = (((!g291) & (g318)));
	assign g320 = (((!g4) & (!g315) & (!g316) & (!g291) & (!g318)) + ((!g4) & (!g315) & (!g316) & (g291) & (!g318)) + ((!g4) & (!g315) & (!g316) & (g291) & (g318)) + ((!g4) & (!g315) & (g316) & (!g291) & (g318)) + ((!g4) & (g315) & (g316) & (!g291) & (!g318)) + ((!g4) & (g315) & (g316) & (!g291) & (g318)) + ((!g4) & (g315) & (g316) & (g291) & (!g318)) + ((!g4) & (g315) & (g316) & (g291) & (g318)) + ((g4) & (!g315) & (g316) & (!g291) & (!g318)) + ((g4) & (!g315) & (g316) & (!g291) & (g318)) + ((g4) & (!g315) & (g316) & (g291) & (!g318)) + ((g4) & (!g315) & (g316) & (g291) & (g318)) + ((g4) & (g315) & (!g316) & (!g291) & (!g318)) + ((g4) & (g315) & (!g316) & (g291) & (!g318)) + ((g4) & (g315) & (!g316) & (g291) & (g318)) + ((g4) & (g315) & (g316) & (!g291) & (g318)));
	assign g321 = (((!g8) & (!g294) & (g314) & (!g291) & (!g318)) + ((!g8) & (!g294) & (g314) & (g291) & (!g318)) + ((!g8) & (!g294) & (g314) & (g291) & (g318)) + ((!g8) & (g294) & (!g314) & (!g291) & (!g318)) + ((!g8) & (g294) & (!g314) & (!g291) & (g318)) + ((!g8) & (g294) & (!g314) & (g291) & (!g318)) + ((!g8) & (g294) & (!g314) & (g291) & (g318)) + ((!g8) & (g294) & (g314) & (!g291) & (g318)) + ((g8) & (!g294) & (!g314) & (!g291) & (!g318)) + ((g8) & (!g294) & (!g314) & (g291) & (!g318)) + ((g8) & (!g294) & (!g314) & (g291) & (g318)) + ((g8) & (g294) & (!g314) & (!g291) & (g318)) + ((g8) & (g294) & (g314) & (!g291) & (!g318)) + ((g8) & (g294) & (g314) & (!g291) & (g318)) + ((g8) & (g294) & (g314) & (g291) & (!g318)) + ((g8) & (g294) & (g314) & (g291) & (g318)));
	assign g322 = (((!g18) & (!g27) & (g296) & (g313)) + ((!g18) & (g27) & (!g296) & (g313)) + ((!g18) & (g27) & (g296) & (!g313)) + ((!g18) & (g27) & (g296) & (g313)) + ((g18) & (!g27) & (!g296) & (!g313)) + ((g18) & (!g27) & (!g296) & (g313)) + ((g18) & (!g27) & (g296) & (!g313)) + ((g18) & (g27) & (!g296) & (!g313)));
	assign g323 = (((!g295) & (!g291) & (!g318) & (g322)) + ((!g295) & (g291) & (!g318) & (g322)) + ((!g295) & (g291) & (g318) & (g322)) + ((g295) & (!g291) & (!g318) & (!g322)) + ((g295) & (!g291) & (g318) & (!g322)) + ((g295) & (!g291) & (g318) & (g322)) + ((g295) & (g291) & (!g318) & (!g322)) + ((g295) & (g291) & (g318) & (!g322)));
	assign g324 = (((!g27) & (!g296) & (g313) & (!g291) & (!g318)) + ((!g27) & (!g296) & (g313) & (g291) & (!g318)) + ((!g27) & (!g296) & (g313) & (g291) & (g318)) + ((!g27) & (g296) & (!g313) & (!g291) & (!g318)) + ((!g27) & (g296) & (!g313) & (!g291) & (g318)) + ((!g27) & (g296) & (!g313) & (g291) & (!g318)) + ((!g27) & (g296) & (!g313) & (g291) & (g318)) + ((!g27) & (g296) & (g313) & (!g291) & (g318)) + ((g27) & (!g296) & (!g313) & (!g291) & (!g318)) + ((g27) & (!g296) & (!g313) & (g291) & (!g318)) + ((g27) & (!g296) & (!g313) & (g291) & (g318)) + ((g27) & (g296) & (!g313) & (!g291) & (g318)) + ((g27) & (g296) & (g313) & (!g291) & (!g318)) + ((g27) & (g296) & (g313) & (!g291) & (g318)) + ((g27) & (g296) & (g313) & (g291) & (!g318)) + ((g27) & (g296) & (g313) & (g291) & (g318)));
	assign g325 = (((!g39) & (!g54) & (g298) & (g312)) + ((!g39) & (g54) & (!g298) & (g312)) + ((!g39) & (g54) & (g298) & (!g312)) + ((!g39) & (g54) & (g298) & (g312)) + ((g39) & (!g54) & (!g298) & (!g312)) + ((g39) & (!g54) & (!g298) & (g312)) + ((g39) & (!g54) & (g298) & (!g312)) + ((g39) & (g54) & (!g298) & (!g312)));
	assign g326 = (((!g297) & (!g291) & (!g318) & (g325)) + ((!g297) & (g291) & (!g318) & (g325)) + ((!g297) & (g291) & (g318) & (g325)) + ((g297) & (!g291) & (!g318) & (!g325)) + ((g297) & (!g291) & (g318) & (!g325)) + ((g297) & (!g291) & (g318) & (g325)) + ((g297) & (g291) & (!g318) & (!g325)) + ((g297) & (g291) & (g318) & (!g325)));
	assign g327 = (((!g54) & (!g298) & (g312) & (!g291) & (!g318)) + ((!g54) & (!g298) & (g312) & (g291) & (!g318)) + ((!g54) & (!g298) & (g312) & (g291) & (g318)) + ((!g54) & (g298) & (!g312) & (!g291) & (!g318)) + ((!g54) & (g298) & (!g312) & (!g291) & (g318)) + ((!g54) & (g298) & (!g312) & (g291) & (!g318)) + ((!g54) & (g298) & (!g312) & (g291) & (g318)) + ((!g54) & (g298) & (g312) & (!g291) & (g318)) + ((g54) & (!g298) & (!g312) & (!g291) & (!g318)) + ((g54) & (!g298) & (!g312) & (g291) & (!g318)) + ((g54) & (!g298) & (!g312) & (g291) & (g318)) + ((g54) & (g298) & (!g312) & (!g291) & (g318)) + ((g54) & (g298) & (g312) & (!g291) & (!g318)) + ((g54) & (g298) & (g312) & (!g291) & (g318)) + ((g54) & (g298) & (g312) & (g291) & (!g318)) + ((g54) & (g298) & (g312) & (g291) & (g318)));
	assign g328 = (((!g68) & (!g87) & (g300) & (g311)) + ((!g68) & (g87) & (!g300) & (g311)) + ((!g68) & (g87) & (g300) & (!g311)) + ((!g68) & (g87) & (g300) & (g311)) + ((g68) & (!g87) & (!g300) & (!g311)) + ((g68) & (!g87) & (!g300) & (g311)) + ((g68) & (!g87) & (g300) & (!g311)) + ((g68) & (g87) & (!g300) & (!g311)));
	assign g329 = (((!g299) & (!g291) & (!g318) & (g328)) + ((!g299) & (g291) & (!g318) & (g328)) + ((!g299) & (g291) & (g318) & (g328)) + ((g299) & (!g291) & (!g318) & (!g328)) + ((g299) & (!g291) & (g318) & (!g328)) + ((g299) & (!g291) & (g318) & (g328)) + ((g299) & (g291) & (!g318) & (!g328)) + ((g299) & (g291) & (g318) & (!g328)));
	assign g330 = (((!g87) & (!g300) & (g311) & (!g291) & (!g318)) + ((!g87) & (!g300) & (g311) & (g291) & (!g318)) + ((!g87) & (!g300) & (g311) & (g291) & (g318)) + ((!g87) & (g300) & (!g311) & (!g291) & (!g318)) + ((!g87) & (g300) & (!g311) & (!g291) & (g318)) + ((!g87) & (g300) & (!g311) & (g291) & (!g318)) + ((!g87) & (g300) & (!g311) & (g291) & (g318)) + ((!g87) & (g300) & (g311) & (!g291) & (g318)) + ((g87) & (!g300) & (!g311) & (!g291) & (!g318)) + ((g87) & (!g300) & (!g311) & (g291) & (!g318)) + ((g87) & (!g300) & (!g311) & (g291) & (g318)) + ((g87) & (g300) & (!g311) & (!g291) & (g318)) + ((g87) & (g300) & (g311) & (!g291) & (!g318)) + ((g87) & (g300) & (g311) & (!g291) & (g318)) + ((g87) & (g300) & (g311) & (g291) & (!g318)) + ((g87) & (g300) & (g311) & (g291) & (g318)));
	assign g331 = (((!g104) & (!g127) & (g302) & (g310)) + ((!g104) & (g127) & (!g302) & (g310)) + ((!g104) & (g127) & (g302) & (!g310)) + ((!g104) & (g127) & (g302) & (g310)) + ((g104) & (!g127) & (!g302) & (!g310)) + ((g104) & (!g127) & (!g302) & (g310)) + ((g104) & (!g127) & (g302) & (!g310)) + ((g104) & (g127) & (!g302) & (!g310)));
	assign g332 = (((!g301) & (!g291) & (!g318) & (g331)) + ((!g301) & (g291) & (!g318) & (g331)) + ((!g301) & (g291) & (g318) & (g331)) + ((g301) & (!g291) & (!g318) & (!g331)) + ((g301) & (!g291) & (g318) & (!g331)) + ((g301) & (!g291) & (g318) & (g331)) + ((g301) & (g291) & (!g318) & (!g331)) + ((g301) & (g291) & (g318) & (!g331)));
	assign g333 = (((!g127) & (!g302) & (g310) & (!g291) & (!g318)) + ((!g127) & (!g302) & (g310) & (g291) & (!g318)) + ((!g127) & (!g302) & (g310) & (g291) & (g318)) + ((!g127) & (g302) & (!g310) & (!g291) & (!g318)) + ((!g127) & (g302) & (!g310) & (!g291) & (g318)) + ((!g127) & (g302) & (!g310) & (g291) & (!g318)) + ((!g127) & (g302) & (!g310) & (g291) & (g318)) + ((!g127) & (g302) & (g310) & (!g291) & (g318)) + ((g127) & (!g302) & (!g310) & (!g291) & (!g318)) + ((g127) & (!g302) & (!g310) & (g291) & (!g318)) + ((g127) & (!g302) & (!g310) & (g291) & (g318)) + ((g127) & (g302) & (!g310) & (!g291) & (g318)) + ((g127) & (g302) & (g310) & (!g291) & (!g318)) + ((g127) & (g302) & (g310) & (!g291) & (g318)) + ((g127) & (g302) & (g310) & (g291) & (!g318)) + ((g127) & (g302) & (g310) & (g291) & (g318)));
	assign g334 = (((!g147) & (!g174) & (g304) & (g309)) + ((!g147) & (g174) & (!g304) & (g309)) + ((!g147) & (g174) & (g304) & (!g309)) + ((!g147) & (g174) & (g304) & (g309)) + ((g147) & (!g174) & (!g304) & (!g309)) + ((g147) & (!g174) & (!g304) & (g309)) + ((g147) & (!g174) & (g304) & (!g309)) + ((g147) & (g174) & (!g304) & (!g309)));
	assign g335 = (((!g303) & (!g291) & (!g318) & (g334)) + ((!g303) & (g291) & (!g318) & (g334)) + ((!g303) & (g291) & (g318) & (g334)) + ((g303) & (!g291) & (!g318) & (!g334)) + ((g303) & (!g291) & (g318) & (!g334)) + ((g303) & (!g291) & (g318) & (g334)) + ((g303) & (g291) & (!g318) & (!g334)) + ((g303) & (g291) & (g318) & (!g334)));
	assign g336 = (((!g174) & (!g304) & (g309) & (!g291) & (!g318)) + ((!g174) & (!g304) & (g309) & (g291) & (!g318)) + ((!g174) & (!g304) & (g309) & (g291) & (g318)) + ((!g174) & (g304) & (!g309) & (!g291) & (!g318)) + ((!g174) & (g304) & (!g309) & (!g291) & (g318)) + ((!g174) & (g304) & (!g309) & (g291) & (!g318)) + ((!g174) & (g304) & (!g309) & (g291) & (g318)) + ((!g174) & (g304) & (g309) & (!g291) & (g318)) + ((g174) & (!g304) & (!g309) & (!g291) & (!g318)) + ((g174) & (!g304) & (!g309) & (g291) & (!g318)) + ((g174) & (!g304) & (!g309) & (g291) & (g318)) + ((g174) & (g304) & (!g309) & (!g291) & (g318)) + ((g174) & (g304) & (g309) & (!g291) & (!g318)) + ((g174) & (g304) & (g309) & (!g291) & (g318)) + ((g174) & (g304) & (g309) & (g291) & (!g318)) + ((g174) & (g304) & (g309) & (g291) & (g318)));
	assign g337 = (((!g198) & (!g229) & (g306) & (g308)) + ((!g198) & (g229) & (!g306) & (g308)) + ((!g198) & (g229) & (g306) & (!g308)) + ((!g198) & (g229) & (g306) & (g308)) + ((g198) & (!g229) & (!g306) & (!g308)) + ((g198) & (!g229) & (!g306) & (g308)) + ((g198) & (!g229) & (g306) & (!g308)) + ((g198) & (g229) & (!g306) & (!g308)));
	assign g338 = (((!g305) & (!g291) & (!g318) & (g337)) + ((!g305) & (g291) & (!g318) & (g337)) + ((!g305) & (g291) & (g318) & (g337)) + ((g305) & (!g291) & (!g318) & (!g337)) + ((g305) & (!g291) & (g318) & (!g337)) + ((g305) & (!g291) & (g318) & (g337)) + ((g305) & (g291) & (!g318) & (!g337)) + ((g305) & (g291) & (g318) & (!g337)));
	assign g339 = (((!g229) & (!g306) & (g308) & (!g291) & (!g318)) + ((!g229) & (!g306) & (g308) & (g291) & (!g318)) + ((!g229) & (!g306) & (g308) & (g291) & (g318)) + ((!g229) & (g306) & (!g308) & (!g291) & (!g318)) + ((!g229) & (g306) & (!g308) & (!g291) & (g318)) + ((!g229) & (g306) & (!g308) & (g291) & (!g318)) + ((!g229) & (g306) & (!g308) & (g291) & (g318)) + ((!g229) & (g306) & (g308) & (!g291) & (g318)) + ((g229) & (!g306) & (!g308) & (!g291) & (!g318)) + ((g229) & (!g306) & (!g308) & (g291) & (!g318)) + ((g229) & (!g306) & (!g308) & (g291) & (g318)) + ((g229) & (g306) & (!g308) & (!g291) & (g318)) + ((g229) & (g306) & (g308) & (!g291) & (!g318)) + ((g229) & (g306) & (g308) & (!g291) & (g318)) + ((g229) & (g306) & (g308) & (g291) & (!g318)) + ((g229) & (g306) & (g308) & (g291) & (g318)));
	assign g340 = (((!g255) & (!ax92x) & (!g290) & (g307)) + ((!g255) & (!ax92x) & (g290) & (g307)) + ((!g255) & (ax92x) & (!g290) & (!g307)) + ((!g255) & (ax92x) & (!g290) & (g307)) + ((g255) & (!ax92x) & (!g290) & (!g307)) + ((g255) & (!ax92x) & (g290) & (!g307)) + ((g255) & (ax92x) & (g290) & (!g307)) + ((g255) & (ax92x) & (g290) & (g307)));
	assign g341 = (((!ax92x) & (!ax93x) & (!g290) & (!g291) & (!g318) & (g340)) + ((!ax92x) & (!ax93x) & (!g290) & (!g291) & (g318) & (!g340)) + ((!ax92x) & (!ax93x) & (!g290) & (!g291) & (g318) & (g340)) + ((!ax92x) & (!ax93x) & (!g290) & (g291) & (!g318) & (g340)) + ((!ax92x) & (!ax93x) & (!g290) & (g291) & (g318) & (g340)) + ((!ax92x) & (!ax93x) & (g290) & (!g291) & (!g318) & (!g340)) + ((!ax92x) & (!ax93x) & (g290) & (g291) & (!g318) & (!g340)) + ((!ax92x) & (!ax93x) & (g290) & (g291) & (g318) & (!g340)) + ((!ax92x) & (ax93x) & (!g290) & (!g291) & (!g318) & (!g340)) + ((!ax92x) & (ax93x) & (!g290) & (g291) & (!g318) & (!g340)) + ((!ax92x) & (ax93x) & (!g290) & (g291) & (g318) & (!g340)) + ((!ax92x) & (ax93x) & (g290) & (!g291) & (!g318) & (g340)) + ((!ax92x) & (ax93x) & (g290) & (!g291) & (g318) & (!g340)) + ((!ax92x) & (ax93x) & (g290) & (!g291) & (g318) & (g340)) + ((!ax92x) & (ax93x) & (g290) & (g291) & (!g318) & (g340)) + ((!ax92x) & (ax93x) & (g290) & (g291) & (g318) & (g340)) + ((ax92x) & (!ax93x) & (!g290) & (!g291) & (!g318) & (!g340)) + ((ax92x) & (!ax93x) & (!g290) & (g291) & (!g318) & (!g340)) + ((ax92x) & (!ax93x) & (!g290) & (g291) & (g318) & (!g340)) + ((ax92x) & (!ax93x) & (g290) & (!g291) & (!g318) & (!g340)) + ((ax92x) & (!ax93x) & (g290) & (g291) & (!g318) & (!g340)) + ((ax92x) & (!ax93x) & (g290) & (g291) & (g318) & (!g340)) + ((ax92x) & (ax93x) & (!g290) & (!g291) & (!g318) & (g340)) + ((ax92x) & (ax93x) & (!g290) & (!g291) & (g318) & (!g340)) + ((ax92x) & (ax93x) & (!g290) & (!g291) & (g318) & (g340)) + ((ax92x) & (ax93x) & (!g290) & (g291) & (!g318) & (g340)) + ((ax92x) & (ax93x) & (!g290) & (g291) & (g318) & (g340)) + ((ax92x) & (ax93x) & (g290) & (!g291) & (!g318) & (g340)) + ((ax92x) & (ax93x) & (g290) & (!g291) & (g318) & (!g340)) + ((ax92x) & (ax93x) & (g290) & (!g291) & (g318) & (g340)) + ((ax92x) & (ax93x) & (g290) & (g291) & (!g318) & (g340)) + ((ax92x) & (ax93x) & (g290) & (g291) & (g318) & (g340)));
	assign g342 = (((!ax92x) & (!g290) & (!g307) & (!g291) & (g318)) + ((!ax92x) & (!g290) & (g307) & (!g291) & (!g318)) + ((!ax92x) & (!g290) & (g307) & (!g291) & (g318)) + ((!ax92x) & (!g290) & (g307) & (g291) & (!g318)) + ((!ax92x) & (!g290) & (g307) & (g291) & (g318)) + ((!ax92x) & (g290) & (g307) & (!g291) & (!g318)) + ((!ax92x) & (g290) & (g307) & (g291) & (!g318)) + ((!ax92x) & (g290) & (g307) & (g291) & (g318)) + ((ax92x) & (!g290) & (!g307) & (!g291) & (!g318)) + ((ax92x) & (!g290) & (!g307) & (g291) & (!g318)) + ((ax92x) & (!g290) & (!g307) & (g291) & (g318)) + ((ax92x) & (g290) & (!g307) & (!g291) & (!g318)) + ((ax92x) & (g290) & (!g307) & (!g291) & (g318)) + ((ax92x) & (g290) & (!g307) & (g291) & (!g318)) + ((ax92x) & (g290) & (!g307) & (g291) & (g318)) + ((ax92x) & (g290) & (g307) & (!g291) & (g318)));
	assign g343 = (((!ax88x) & (!ax89x)));
	assign g344 = (((!g290) & (!ax90x) & (!ax91x) & (!g291) & (!g318) & (!g343)) + ((!g290) & (!ax90x) & (!ax91x) & (g291) & (!g318) & (!g343)) + ((!g290) & (!ax90x) & (!ax91x) & (g291) & (g318) & (!g343)) + ((!g290) & (!ax90x) & (ax91x) & (!g291) & (g318) & (!g343)) + ((!g290) & (ax90x) & (ax91x) & (!g291) & (g318) & (!g343)) + ((!g290) & (ax90x) & (ax91x) & (!g291) & (g318) & (g343)) + ((g290) & (!ax90x) & (!ax91x) & (!g291) & (!g318) & (!g343)) + ((g290) & (!ax90x) & (!ax91x) & (!g291) & (!g318) & (g343)) + ((g290) & (!ax90x) & (!ax91x) & (!g291) & (g318) & (!g343)) + ((g290) & (!ax90x) & (!ax91x) & (g291) & (!g318) & (!g343)) + ((g290) & (!ax90x) & (!ax91x) & (g291) & (!g318) & (g343)) + ((g290) & (!ax90x) & (!ax91x) & (g291) & (g318) & (!g343)) + ((g290) & (!ax90x) & (!ax91x) & (g291) & (g318) & (g343)) + ((g290) & (!ax90x) & (ax91x) & (!g291) & (!g318) & (!g343)) + ((g290) & (!ax90x) & (ax91x) & (!g291) & (g318) & (!g343)) + ((g290) & (!ax90x) & (ax91x) & (!g291) & (g318) & (g343)) + ((g290) & (!ax90x) & (ax91x) & (g291) & (!g318) & (!g343)) + ((g290) & (!ax90x) & (ax91x) & (g291) & (g318) & (!g343)) + ((g290) & (ax90x) & (!ax91x) & (!g291) & (g318) & (!g343)) + ((g290) & (ax90x) & (!ax91x) & (!g291) & (g318) & (g343)) + ((g290) & (ax90x) & (ax91x) & (!g291) & (!g318) & (!g343)) + ((g290) & (ax90x) & (ax91x) & (!g291) & (!g318) & (g343)) + ((g290) & (ax90x) & (ax91x) & (!g291) & (g318) & (!g343)) + ((g290) & (ax90x) & (ax91x) & (!g291) & (g318) & (g343)) + ((g290) & (ax90x) & (ax91x) & (g291) & (!g318) & (!g343)) + ((g290) & (ax90x) & (ax91x) & (g291) & (!g318) & (g343)) + ((g290) & (ax90x) & (ax91x) & (g291) & (g318) & (!g343)) + ((g290) & (ax90x) & (ax91x) & (g291) & (g318) & (g343)));
	assign g345 = (((!g229) & (!g255) & (g341) & (g342) & (g344)) + ((!g229) & (g255) & (g341) & (!g342) & (g344)) + ((!g229) & (g255) & (g341) & (g342) & (!g344)) + ((!g229) & (g255) & (g341) & (g342) & (g344)) + ((g229) & (!g255) & (!g341) & (g342) & (g344)) + ((g229) & (!g255) & (g341) & (!g342) & (!g344)) + ((g229) & (!g255) & (g341) & (!g342) & (g344)) + ((g229) & (!g255) & (g341) & (g342) & (!g344)) + ((g229) & (!g255) & (g341) & (g342) & (g344)) + ((g229) & (g255) & (!g341) & (!g342) & (g344)) + ((g229) & (g255) & (!g341) & (g342) & (!g344)) + ((g229) & (g255) & (!g341) & (g342) & (g344)) + ((g229) & (g255) & (g341) & (!g342) & (!g344)) + ((g229) & (g255) & (g341) & (!g342) & (g344)) + ((g229) & (g255) & (g341) & (g342) & (!g344)) + ((g229) & (g255) & (g341) & (g342) & (g344)));
	assign g346 = (((!g174) & (!g198) & (g338) & (g339) & (g345)) + ((!g174) & (g198) & (g338) & (!g339) & (g345)) + ((!g174) & (g198) & (g338) & (g339) & (!g345)) + ((!g174) & (g198) & (g338) & (g339) & (g345)) + ((g174) & (!g198) & (!g338) & (g339) & (g345)) + ((g174) & (!g198) & (g338) & (!g339) & (!g345)) + ((g174) & (!g198) & (g338) & (!g339) & (g345)) + ((g174) & (!g198) & (g338) & (g339) & (!g345)) + ((g174) & (!g198) & (g338) & (g339) & (g345)) + ((g174) & (g198) & (!g338) & (!g339) & (g345)) + ((g174) & (g198) & (!g338) & (g339) & (!g345)) + ((g174) & (g198) & (!g338) & (g339) & (g345)) + ((g174) & (g198) & (g338) & (!g339) & (!g345)) + ((g174) & (g198) & (g338) & (!g339) & (g345)) + ((g174) & (g198) & (g338) & (g339) & (!g345)) + ((g174) & (g198) & (g338) & (g339) & (g345)));
	assign g347 = (((!g127) & (!g147) & (g335) & (g336) & (g346)) + ((!g127) & (g147) & (g335) & (!g336) & (g346)) + ((!g127) & (g147) & (g335) & (g336) & (!g346)) + ((!g127) & (g147) & (g335) & (g336) & (g346)) + ((g127) & (!g147) & (!g335) & (g336) & (g346)) + ((g127) & (!g147) & (g335) & (!g336) & (!g346)) + ((g127) & (!g147) & (g335) & (!g336) & (g346)) + ((g127) & (!g147) & (g335) & (g336) & (!g346)) + ((g127) & (!g147) & (g335) & (g336) & (g346)) + ((g127) & (g147) & (!g335) & (!g336) & (g346)) + ((g127) & (g147) & (!g335) & (g336) & (!g346)) + ((g127) & (g147) & (!g335) & (g336) & (g346)) + ((g127) & (g147) & (g335) & (!g336) & (!g346)) + ((g127) & (g147) & (g335) & (!g336) & (g346)) + ((g127) & (g147) & (g335) & (g336) & (!g346)) + ((g127) & (g147) & (g335) & (g336) & (g346)));
	assign g348 = (((!g87) & (!g104) & (g332) & (g333) & (g347)) + ((!g87) & (g104) & (g332) & (!g333) & (g347)) + ((!g87) & (g104) & (g332) & (g333) & (!g347)) + ((!g87) & (g104) & (g332) & (g333) & (g347)) + ((g87) & (!g104) & (!g332) & (g333) & (g347)) + ((g87) & (!g104) & (g332) & (!g333) & (!g347)) + ((g87) & (!g104) & (g332) & (!g333) & (g347)) + ((g87) & (!g104) & (g332) & (g333) & (!g347)) + ((g87) & (!g104) & (g332) & (g333) & (g347)) + ((g87) & (g104) & (!g332) & (!g333) & (g347)) + ((g87) & (g104) & (!g332) & (g333) & (!g347)) + ((g87) & (g104) & (!g332) & (g333) & (g347)) + ((g87) & (g104) & (g332) & (!g333) & (!g347)) + ((g87) & (g104) & (g332) & (!g333) & (g347)) + ((g87) & (g104) & (g332) & (g333) & (!g347)) + ((g87) & (g104) & (g332) & (g333) & (g347)));
	assign g349 = (((!g54) & (!g68) & (g329) & (g330) & (g348)) + ((!g54) & (g68) & (g329) & (!g330) & (g348)) + ((!g54) & (g68) & (g329) & (g330) & (!g348)) + ((!g54) & (g68) & (g329) & (g330) & (g348)) + ((g54) & (!g68) & (!g329) & (g330) & (g348)) + ((g54) & (!g68) & (g329) & (!g330) & (!g348)) + ((g54) & (!g68) & (g329) & (!g330) & (g348)) + ((g54) & (!g68) & (g329) & (g330) & (!g348)) + ((g54) & (!g68) & (g329) & (g330) & (g348)) + ((g54) & (g68) & (!g329) & (!g330) & (g348)) + ((g54) & (g68) & (!g329) & (g330) & (!g348)) + ((g54) & (g68) & (!g329) & (g330) & (g348)) + ((g54) & (g68) & (g329) & (!g330) & (!g348)) + ((g54) & (g68) & (g329) & (!g330) & (g348)) + ((g54) & (g68) & (g329) & (g330) & (!g348)) + ((g54) & (g68) & (g329) & (g330) & (g348)));
	assign g350 = (((!g27) & (!g39) & (g326) & (g327) & (g349)) + ((!g27) & (g39) & (g326) & (!g327) & (g349)) + ((!g27) & (g39) & (g326) & (g327) & (!g349)) + ((!g27) & (g39) & (g326) & (g327) & (g349)) + ((g27) & (!g39) & (!g326) & (g327) & (g349)) + ((g27) & (!g39) & (g326) & (!g327) & (!g349)) + ((g27) & (!g39) & (g326) & (!g327) & (g349)) + ((g27) & (!g39) & (g326) & (g327) & (!g349)) + ((g27) & (!g39) & (g326) & (g327) & (g349)) + ((g27) & (g39) & (!g326) & (!g327) & (g349)) + ((g27) & (g39) & (!g326) & (g327) & (!g349)) + ((g27) & (g39) & (!g326) & (g327) & (g349)) + ((g27) & (g39) & (g326) & (!g327) & (!g349)) + ((g27) & (g39) & (g326) & (!g327) & (g349)) + ((g27) & (g39) & (g326) & (g327) & (!g349)) + ((g27) & (g39) & (g326) & (g327) & (g349)));
	assign g351 = (((!g8) & (!g18) & (g323) & (g324) & (g350)) + ((!g8) & (g18) & (g323) & (!g324) & (g350)) + ((!g8) & (g18) & (g323) & (g324) & (!g350)) + ((!g8) & (g18) & (g323) & (g324) & (g350)) + ((g8) & (!g18) & (!g323) & (g324) & (g350)) + ((g8) & (!g18) & (g323) & (!g324) & (!g350)) + ((g8) & (!g18) & (g323) & (!g324) & (g350)) + ((g8) & (!g18) & (g323) & (g324) & (!g350)) + ((g8) & (!g18) & (g323) & (g324) & (g350)) + ((g8) & (g18) & (!g323) & (!g324) & (g350)) + ((g8) & (g18) & (!g323) & (g324) & (!g350)) + ((g8) & (g18) & (!g323) & (g324) & (g350)) + ((g8) & (g18) & (g323) & (!g324) & (!g350)) + ((g8) & (g18) & (g323) & (!g324) & (g350)) + ((g8) & (g18) & (g323) & (g324) & (!g350)) + ((g8) & (g18) & (g323) & (g324) & (g350)));
	assign g352 = (((!g2) & (!g8) & (g294) & (g314)) + ((!g2) & (g8) & (!g294) & (g314)) + ((!g2) & (g8) & (g294) & (!g314)) + ((!g2) & (g8) & (g294) & (g314)) + ((g2) & (!g8) & (!g294) & (!g314)) + ((g2) & (!g8) & (!g294) & (g314)) + ((g2) & (!g8) & (g294) & (!g314)) + ((g2) & (g8) & (!g294) & (!g314)));
	assign g353 = (((!g293) & (!g291) & (!g318) & (g352)) + ((!g293) & (g291) & (!g318) & (g352)) + ((!g293) & (g291) & (g318) & (g352)) + ((g293) & (!g291) & (!g318) & (!g352)) + ((g293) & (!g291) & (g318) & (!g352)) + ((g293) & (!g291) & (g318) & (g352)) + ((g293) & (g291) & (!g318) & (!g352)) + ((g293) & (g291) & (g318) & (!g352)));
	assign g354 = (((!g4) & (!g2) & (!g321) & (!g351) & (g353)) + ((!g4) & (!g2) & (!g321) & (g351) & (g353)) + ((!g4) & (!g2) & (g321) & (!g351) & (g353)) + ((!g4) & (!g2) & (g321) & (g351) & (!g353)) + ((!g4) & (!g2) & (g321) & (g351) & (g353)) + ((!g4) & (g2) & (!g321) & (!g351) & (g353)) + ((!g4) & (g2) & (!g321) & (g351) & (!g353)) + ((!g4) & (g2) & (!g321) & (g351) & (g353)) + ((!g4) & (g2) & (g321) & (!g351) & (!g353)) + ((!g4) & (g2) & (g321) & (!g351) & (g353)) + ((!g4) & (g2) & (g321) & (g351) & (!g353)) + ((!g4) & (g2) & (g321) & (g351) & (g353)) + ((g4) & (!g2) & (g321) & (g351) & (g353)) + ((g4) & (g2) & (!g321) & (g351) & (g353)) + ((g4) & (g2) & (g321) & (!g351) & (g353)) + ((g4) & (g2) & (g321) & (g351) & (g353)));
	assign g355 = (((!g4) & (!g315) & (g316)) + ((!g4) & (g315) & (!g316)) + ((!g4) & (g315) & (g316)) + ((g4) & (g315) & (g316)));
	assign g356 = (((!g292) & (!g355) & (!g291) & (!g318)) + ((!g292) & (!g355) & (g291) & (!g318)) + ((!g292) & (!g355) & (g291) & (g318)) + ((g292) & (g355) & (!g291) & (!g318)) + ((g292) & (g355) & (!g291) & (g318)) + ((g292) & (g355) & (g291) & (!g318)) + ((g292) & (g355) & (g291) & (g318)));
	assign g357 = (((!g1) & (g292) & (!g355) & (!g291) & (g318)) + ((!g1) & (g292) & (g355) & (!g291) & (g318)) + ((g1) & (!g292) & (g355) & (g291) & (!g318)) + ((g1) & (!g292) & (g355) & (g291) & (g318)) + ((g1) & (g292) & (!g355) & (!g291) & (!g318)) + ((g1) & (g292) & (!g355) & (!g291) & (g318)) + ((g1) & (g292) & (!g355) & (g291) & (!g318)) + ((g1) & (g292) & (!g355) & (g291) & (g318)) + ((g1) & (g292) & (g355) & (!g291) & (g318)));
	assign g358 = (((!g1) & (!g320) & (!g354) & (!g356) & (!g357)) + ((g1) & (!g320) & (!g354) & (!g356) & (!g357)) + ((g1) & (!g320) & (!g354) & (g356) & (!g357)) + ((g1) & (!g320) & (g354) & (!g356) & (!g357)) + ((g1) & (!g320) & (g354) & (g356) & (!g357)) + ((g1) & (g320) & (!g354) & (!g356) & (!g357)) + ((g1) & (g320) & (!g354) & (g356) & (!g357)));
	assign g359 = (((g1) & (!g320) & (g354) & (g357)) + ((g1) & (g320) & (!g354) & (!g357)) + ((g1) & (g320) & (!g354) & (g357)));
	assign g360 = (((!g4) & (!g2) & (!g321) & (!g351) & (!g353) & (!g358)) + ((!g4) & (!g2) & (!g321) & (!g351) & (g353) & (g358)) + ((!g4) & (!g2) & (!g321) & (g351) & (!g353) & (!g358)) + ((!g4) & (!g2) & (!g321) & (g351) & (g353) & (g358)) + ((!g4) & (!g2) & (g321) & (!g351) & (!g353) & (!g358)) + ((!g4) & (!g2) & (g321) & (!g351) & (g353) & (g358)) + ((!g4) & (!g2) & (g321) & (g351) & (g353) & (!g358)) + ((!g4) & (!g2) & (g321) & (g351) & (g353) & (g358)) + ((!g4) & (g2) & (!g321) & (!g351) & (!g353) & (!g358)) + ((!g4) & (g2) & (!g321) & (!g351) & (g353) & (g358)) + ((!g4) & (g2) & (!g321) & (g351) & (g353) & (!g358)) + ((!g4) & (g2) & (!g321) & (g351) & (g353) & (g358)) + ((!g4) & (g2) & (g321) & (!g351) & (g353) & (!g358)) + ((!g4) & (g2) & (g321) & (!g351) & (g353) & (g358)) + ((!g4) & (g2) & (g321) & (g351) & (g353) & (!g358)) + ((!g4) & (g2) & (g321) & (g351) & (g353) & (g358)) + ((g4) & (!g2) & (!g321) & (!g351) & (g353) & (!g358)) + ((g4) & (!g2) & (!g321) & (!g351) & (g353) & (g358)) + ((g4) & (!g2) & (!g321) & (g351) & (g353) & (!g358)) + ((g4) & (!g2) & (!g321) & (g351) & (g353) & (g358)) + ((g4) & (!g2) & (g321) & (!g351) & (g353) & (!g358)) + ((g4) & (!g2) & (g321) & (!g351) & (g353) & (g358)) + ((g4) & (!g2) & (g321) & (g351) & (!g353) & (!g358)) + ((g4) & (!g2) & (g321) & (g351) & (g353) & (g358)) + ((g4) & (g2) & (!g321) & (!g351) & (g353) & (!g358)) + ((g4) & (g2) & (!g321) & (!g351) & (g353) & (g358)) + ((g4) & (g2) & (!g321) & (g351) & (!g353) & (!g358)) + ((g4) & (g2) & (!g321) & (g351) & (g353) & (g358)) + ((g4) & (g2) & (g321) & (!g351) & (!g353) & (!g358)) + ((g4) & (g2) & (g321) & (!g351) & (g353) & (g358)) + ((g4) & (g2) & (g321) & (g351) & (!g353) & (!g358)) + ((g4) & (g2) & (g321) & (g351) & (g353) & (g358)));
	assign g361 = (((!g8) & (!g18) & (!g323) & (g324) & (g350) & (!g358)) + ((!g8) & (!g18) & (g323) & (!g324) & (!g350) & (!g358)) + ((!g8) & (!g18) & (g323) & (!g324) & (!g350) & (g358)) + ((!g8) & (!g18) & (g323) & (!g324) & (g350) & (!g358)) + ((!g8) & (!g18) & (g323) & (!g324) & (g350) & (g358)) + ((!g8) & (!g18) & (g323) & (g324) & (!g350) & (!g358)) + ((!g8) & (!g18) & (g323) & (g324) & (!g350) & (g358)) + ((!g8) & (!g18) & (g323) & (g324) & (g350) & (g358)) + ((!g8) & (g18) & (!g323) & (!g324) & (g350) & (!g358)) + ((!g8) & (g18) & (!g323) & (g324) & (!g350) & (!g358)) + ((!g8) & (g18) & (!g323) & (g324) & (g350) & (!g358)) + ((!g8) & (g18) & (g323) & (!g324) & (!g350) & (!g358)) + ((!g8) & (g18) & (g323) & (!g324) & (!g350) & (g358)) + ((!g8) & (g18) & (g323) & (!g324) & (g350) & (g358)) + ((!g8) & (g18) & (g323) & (g324) & (!g350) & (g358)) + ((!g8) & (g18) & (g323) & (g324) & (g350) & (g358)) + ((g8) & (!g18) & (!g323) & (!g324) & (!g350) & (!g358)) + ((g8) & (!g18) & (!g323) & (!g324) & (g350) & (!g358)) + ((g8) & (!g18) & (!g323) & (g324) & (!g350) & (!g358)) + ((g8) & (!g18) & (g323) & (!g324) & (!g350) & (g358)) + ((g8) & (!g18) & (g323) & (!g324) & (g350) & (g358)) + ((g8) & (!g18) & (g323) & (g324) & (!g350) & (g358)) + ((g8) & (!g18) & (g323) & (g324) & (g350) & (!g358)) + ((g8) & (!g18) & (g323) & (g324) & (g350) & (g358)) + ((g8) & (g18) & (!g323) & (!g324) & (!g350) & (!g358)) + ((g8) & (g18) & (g323) & (!g324) & (!g350) & (g358)) + ((g8) & (g18) & (g323) & (!g324) & (g350) & (!g358)) + ((g8) & (g18) & (g323) & (!g324) & (g350) & (g358)) + ((g8) & (g18) & (g323) & (g324) & (!g350) & (!g358)) + ((g8) & (g18) & (g323) & (g324) & (!g350) & (g358)) + ((g8) & (g18) & (g323) & (g324) & (g350) & (!g358)) + ((g8) & (g18) & (g323) & (g324) & (g350) & (g358)));
	assign g362 = (((!g18) & (!g324) & (g350) & (!g358)) + ((!g18) & (g324) & (!g350) & (!g358)) + ((!g18) & (g324) & (!g350) & (g358)) + ((!g18) & (g324) & (g350) & (g358)) + ((g18) & (!g324) & (!g350) & (!g358)) + ((g18) & (g324) & (!g350) & (g358)) + ((g18) & (g324) & (g350) & (!g358)) + ((g18) & (g324) & (g350) & (g358)));
	assign g363 = (((!g27) & (!g39) & (!g326) & (g327) & (g349) & (!g358)) + ((!g27) & (!g39) & (g326) & (!g327) & (!g349) & (!g358)) + ((!g27) & (!g39) & (g326) & (!g327) & (!g349) & (g358)) + ((!g27) & (!g39) & (g326) & (!g327) & (g349) & (!g358)) + ((!g27) & (!g39) & (g326) & (!g327) & (g349) & (g358)) + ((!g27) & (!g39) & (g326) & (g327) & (!g349) & (!g358)) + ((!g27) & (!g39) & (g326) & (g327) & (!g349) & (g358)) + ((!g27) & (!g39) & (g326) & (g327) & (g349) & (g358)) + ((!g27) & (g39) & (!g326) & (!g327) & (g349) & (!g358)) + ((!g27) & (g39) & (!g326) & (g327) & (!g349) & (!g358)) + ((!g27) & (g39) & (!g326) & (g327) & (g349) & (!g358)) + ((!g27) & (g39) & (g326) & (!g327) & (!g349) & (!g358)) + ((!g27) & (g39) & (g326) & (!g327) & (!g349) & (g358)) + ((!g27) & (g39) & (g326) & (!g327) & (g349) & (g358)) + ((!g27) & (g39) & (g326) & (g327) & (!g349) & (g358)) + ((!g27) & (g39) & (g326) & (g327) & (g349) & (g358)) + ((g27) & (!g39) & (!g326) & (!g327) & (!g349) & (!g358)) + ((g27) & (!g39) & (!g326) & (!g327) & (g349) & (!g358)) + ((g27) & (!g39) & (!g326) & (g327) & (!g349) & (!g358)) + ((g27) & (!g39) & (g326) & (!g327) & (!g349) & (g358)) + ((g27) & (!g39) & (g326) & (!g327) & (g349) & (g358)) + ((g27) & (!g39) & (g326) & (g327) & (!g349) & (g358)) + ((g27) & (!g39) & (g326) & (g327) & (g349) & (!g358)) + ((g27) & (!g39) & (g326) & (g327) & (g349) & (g358)) + ((g27) & (g39) & (!g326) & (!g327) & (!g349) & (!g358)) + ((g27) & (g39) & (g326) & (!g327) & (!g349) & (g358)) + ((g27) & (g39) & (g326) & (!g327) & (g349) & (!g358)) + ((g27) & (g39) & (g326) & (!g327) & (g349) & (g358)) + ((g27) & (g39) & (g326) & (g327) & (!g349) & (!g358)) + ((g27) & (g39) & (g326) & (g327) & (!g349) & (g358)) + ((g27) & (g39) & (g326) & (g327) & (g349) & (!g358)) + ((g27) & (g39) & (g326) & (g327) & (g349) & (g358)));
	assign g364 = (((!g39) & (!g327) & (g349) & (!g358)) + ((!g39) & (g327) & (!g349) & (!g358)) + ((!g39) & (g327) & (!g349) & (g358)) + ((!g39) & (g327) & (g349) & (g358)) + ((g39) & (!g327) & (!g349) & (!g358)) + ((g39) & (g327) & (!g349) & (g358)) + ((g39) & (g327) & (g349) & (!g358)) + ((g39) & (g327) & (g349) & (g358)));
	assign g365 = (((!g54) & (!g68) & (!g329) & (g330) & (g348) & (!g358)) + ((!g54) & (!g68) & (g329) & (!g330) & (!g348) & (!g358)) + ((!g54) & (!g68) & (g329) & (!g330) & (!g348) & (g358)) + ((!g54) & (!g68) & (g329) & (!g330) & (g348) & (!g358)) + ((!g54) & (!g68) & (g329) & (!g330) & (g348) & (g358)) + ((!g54) & (!g68) & (g329) & (g330) & (!g348) & (!g358)) + ((!g54) & (!g68) & (g329) & (g330) & (!g348) & (g358)) + ((!g54) & (!g68) & (g329) & (g330) & (g348) & (g358)) + ((!g54) & (g68) & (!g329) & (!g330) & (g348) & (!g358)) + ((!g54) & (g68) & (!g329) & (g330) & (!g348) & (!g358)) + ((!g54) & (g68) & (!g329) & (g330) & (g348) & (!g358)) + ((!g54) & (g68) & (g329) & (!g330) & (!g348) & (!g358)) + ((!g54) & (g68) & (g329) & (!g330) & (!g348) & (g358)) + ((!g54) & (g68) & (g329) & (!g330) & (g348) & (g358)) + ((!g54) & (g68) & (g329) & (g330) & (!g348) & (g358)) + ((!g54) & (g68) & (g329) & (g330) & (g348) & (g358)) + ((g54) & (!g68) & (!g329) & (!g330) & (!g348) & (!g358)) + ((g54) & (!g68) & (!g329) & (!g330) & (g348) & (!g358)) + ((g54) & (!g68) & (!g329) & (g330) & (!g348) & (!g358)) + ((g54) & (!g68) & (g329) & (!g330) & (!g348) & (g358)) + ((g54) & (!g68) & (g329) & (!g330) & (g348) & (g358)) + ((g54) & (!g68) & (g329) & (g330) & (!g348) & (g358)) + ((g54) & (!g68) & (g329) & (g330) & (g348) & (!g358)) + ((g54) & (!g68) & (g329) & (g330) & (g348) & (g358)) + ((g54) & (g68) & (!g329) & (!g330) & (!g348) & (!g358)) + ((g54) & (g68) & (g329) & (!g330) & (!g348) & (g358)) + ((g54) & (g68) & (g329) & (!g330) & (g348) & (!g358)) + ((g54) & (g68) & (g329) & (!g330) & (g348) & (g358)) + ((g54) & (g68) & (g329) & (g330) & (!g348) & (!g358)) + ((g54) & (g68) & (g329) & (g330) & (!g348) & (g358)) + ((g54) & (g68) & (g329) & (g330) & (g348) & (!g358)) + ((g54) & (g68) & (g329) & (g330) & (g348) & (g358)));
	assign g366 = (((!g68) & (!g330) & (g348) & (!g358)) + ((!g68) & (g330) & (!g348) & (!g358)) + ((!g68) & (g330) & (!g348) & (g358)) + ((!g68) & (g330) & (g348) & (g358)) + ((g68) & (!g330) & (!g348) & (!g358)) + ((g68) & (g330) & (!g348) & (g358)) + ((g68) & (g330) & (g348) & (!g358)) + ((g68) & (g330) & (g348) & (g358)));
	assign g367 = (((!g87) & (!g104) & (!g332) & (g333) & (g347) & (!g358)) + ((!g87) & (!g104) & (g332) & (!g333) & (!g347) & (!g358)) + ((!g87) & (!g104) & (g332) & (!g333) & (!g347) & (g358)) + ((!g87) & (!g104) & (g332) & (!g333) & (g347) & (!g358)) + ((!g87) & (!g104) & (g332) & (!g333) & (g347) & (g358)) + ((!g87) & (!g104) & (g332) & (g333) & (!g347) & (!g358)) + ((!g87) & (!g104) & (g332) & (g333) & (!g347) & (g358)) + ((!g87) & (!g104) & (g332) & (g333) & (g347) & (g358)) + ((!g87) & (g104) & (!g332) & (!g333) & (g347) & (!g358)) + ((!g87) & (g104) & (!g332) & (g333) & (!g347) & (!g358)) + ((!g87) & (g104) & (!g332) & (g333) & (g347) & (!g358)) + ((!g87) & (g104) & (g332) & (!g333) & (!g347) & (!g358)) + ((!g87) & (g104) & (g332) & (!g333) & (!g347) & (g358)) + ((!g87) & (g104) & (g332) & (!g333) & (g347) & (g358)) + ((!g87) & (g104) & (g332) & (g333) & (!g347) & (g358)) + ((!g87) & (g104) & (g332) & (g333) & (g347) & (g358)) + ((g87) & (!g104) & (!g332) & (!g333) & (!g347) & (!g358)) + ((g87) & (!g104) & (!g332) & (!g333) & (g347) & (!g358)) + ((g87) & (!g104) & (!g332) & (g333) & (!g347) & (!g358)) + ((g87) & (!g104) & (g332) & (!g333) & (!g347) & (g358)) + ((g87) & (!g104) & (g332) & (!g333) & (g347) & (g358)) + ((g87) & (!g104) & (g332) & (g333) & (!g347) & (g358)) + ((g87) & (!g104) & (g332) & (g333) & (g347) & (!g358)) + ((g87) & (!g104) & (g332) & (g333) & (g347) & (g358)) + ((g87) & (g104) & (!g332) & (!g333) & (!g347) & (!g358)) + ((g87) & (g104) & (g332) & (!g333) & (!g347) & (g358)) + ((g87) & (g104) & (g332) & (!g333) & (g347) & (!g358)) + ((g87) & (g104) & (g332) & (!g333) & (g347) & (g358)) + ((g87) & (g104) & (g332) & (g333) & (!g347) & (!g358)) + ((g87) & (g104) & (g332) & (g333) & (!g347) & (g358)) + ((g87) & (g104) & (g332) & (g333) & (g347) & (!g358)) + ((g87) & (g104) & (g332) & (g333) & (g347) & (g358)));
	assign g368 = (((!g104) & (!g333) & (g347) & (!g358)) + ((!g104) & (g333) & (!g347) & (!g358)) + ((!g104) & (g333) & (!g347) & (g358)) + ((!g104) & (g333) & (g347) & (g358)) + ((g104) & (!g333) & (!g347) & (!g358)) + ((g104) & (g333) & (!g347) & (g358)) + ((g104) & (g333) & (g347) & (!g358)) + ((g104) & (g333) & (g347) & (g358)));
	assign g369 = (((!g127) & (!g147) & (!g335) & (g336) & (g346) & (!g358)) + ((!g127) & (!g147) & (g335) & (!g336) & (!g346) & (!g358)) + ((!g127) & (!g147) & (g335) & (!g336) & (!g346) & (g358)) + ((!g127) & (!g147) & (g335) & (!g336) & (g346) & (!g358)) + ((!g127) & (!g147) & (g335) & (!g336) & (g346) & (g358)) + ((!g127) & (!g147) & (g335) & (g336) & (!g346) & (!g358)) + ((!g127) & (!g147) & (g335) & (g336) & (!g346) & (g358)) + ((!g127) & (!g147) & (g335) & (g336) & (g346) & (g358)) + ((!g127) & (g147) & (!g335) & (!g336) & (g346) & (!g358)) + ((!g127) & (g147) & (!g335) & (g336) & (!g346) & (!g358)) + ((!g127) & (g147) & (!g335) & (g336) & (g346) & (!g358)) + ((!g127) & (g147) & (g335) & (!g336) & (!g346) & (!g358)) + ((!g127) & (g147) & (g335) & (!g336) & (!g346) & (g358)) + ((!g127) & (g147) & (g335) & (!g336) & (g346) & (g358)) + ((!g127) & (g147) & (g335) & (g336) & (!g346) & (g358)) + ((!g127) & (g147) & (g335) & (g336) & (g346) & (g358)) + ((g127) & (!g147) & (!g335) & (!g336) & (!g346) & (!g358)) + ((g127) & (!g147) & (!g335) & (!g336) & (g346) & (!g358)) + ((g127) & (!g147) & (!g335) & (g336) & (!g346) & (!g358)) + ((g127) & (!g147) & (g335) & (!g336) & (!g346) & (g358)) + ((g127) & (!g147) & (g335) & (!g336) & (g346) & (g358)) + ((g127) & (!g147) & (g335) & (g336) & (!g346) & (g358)) + ((g127) & (!g147) & (g335) & (g336) & (g346) & (!g358)) + ((g127) & (!g147) & (g335) & (g336) & (g346) & (g358)) + ((g127) & (g147) & (!g335) & (!g336) & (!g346) & (!g358)) + ((g127) & (g147) & (g335) & (!g336) & (!g346) & (g358)) + ((g127) & (g147) & (g335) & (!g336) & (g346) & (!g358)) + ((g127) & (g147) & (g335) & (!g336) & (g346) & (g358)) + ((g127) & (g147) & (g335) & (g336) & (!g346) & (!g358)) + ((g127) & (g147) & (g335) & (g336) & (!g346) & (g358)) + ((g127) & (g147) & (g335) & (g336) & (g346) & (!g358)) + ((g127) & (g147) & (g335) & (g336) & (g346) & (g358)));
	assign g370 = (((!g147) & (!g336) & (g346) & (!g358)) + ((!g147) & (g336) & (!g346) & (!g358)) + ((!g147) & (g336) & (!g346) & (g358)) + ((!g147) & (g336) & (g346) & (g358)) + ((g147) & (!g336) & (!g346) & (!g358)) + ((g147) & (g336) & (!g346) & (g358)) + ((g147) & (g336) & (g346) & (!g358)) + ((g147) & (g336) & (g346) & (g358)));
	assign g371 = (((!g174) & (!g198) & (!g338) & (g339) & (g345) & (!g358)) + ((!g174) & (!g198) & (g338) & (!g339) & (!g345) & (!g358)) + ((!g174) & (!g198) & (g338) & (!g339) & (!g345) & (g358)) + ((!g174) & (!g198) & (g338) & (!g339) & (g345) & (!g358)) + ((!g174) & (!g198) & (g338) & (!g339) & (g345) & (g358)) + ((!g174) & (!g198) & (g338) & (g339) & (!g345) & (!g358)) + ((!g174) & (!g198) & (g338) & (g339) & (!g345) & (g358)) + ((!g174) & (!g198) & (g338) & (g339) & (g345) & (g358)) + ((!g174) & (g198) & (!g338) & (!g339) & (g345) & (!g358)) + ((!g174) & (g198) & (!g338) & (g339) & (!g345) & (!g358)) + ((!g174) & (g198) & (!g338) & (g339) & (g345) & (!g358)) + ((!g174) & (g198) & (g338) & (!g339) & (!g345) & (!g358)) + ((!g174) & (g198) & (g338) & (!g339) & (!g345) & (g358)) + ((!g174) & (g198) & (g338) & (!g339) & (g345) & (g358)) + ((!g174) & (g198) & (g338) & (g339) & (!g345) & (g358)) + ((!g174) & (g198) & (g338) & (g339) & (g345) & (g358)) + ((g174) & (!g198) & (!g338) & (!g339) & (!g345) & (!g358)) + ((g174) & (!g198) & (!g338) & (!g339) & (g345) & (!g358)) + ((g174) & (!g198) & (!g338) & (g339) & (!g345) & (!g358)) + ((g174) & (!g198) & (g338) & (!g339) & (!g345) & (g358)) + ((g174) & (!g198) & (g338) & (!g339) & (g345) & (g358)) + ((g174) & (!g198) & (g338) & (g339) & (!g345) & (g358)) + ((g174) & (!g198) & (g338) & (g339) & (g345) & (!g358)) + ((g174) & (!g198) & (g338) & (g339) & (g345) & (g358)) + ((g174) & (g198) & (!g338) & (!g339) & (!g345) & (!g358)) + ((g174) & (g198) & (g338) & (!g339) & (!g345) & (g358)) + ((g174) & (g198) & (g338) & (!g339) & (g345) & (!g358)) + ((g174) & (g198) & (g338) & (!g339) & (g345) & (g358)) + ((g174) & (g198) & (g338) & (g339) & (!g345) & (!g358)) + ((g174) & (g198) & (g338) & (g339) & (!g345) & (g358)) + ((g174) & (g198) & (g338) & (g339) & (g345) & (!g358)) + ((g174) & (g198) & (g338) & (g339) & (g345) & (g358)));
	assign g372 = (((!g198) & (!g339) & (g345) & (!g358)) + ((!g198) & (g339) & (!g345) & (!g358)) + ((!g198) & (g339) & (!g345) & (g358)) + ((!g198) & (g339) & (g345) & (g358)) + ((g198) & (!g339) & (!g345) & (!g358)) + ((g198) & (g339) & (!g345) & (g358)) + ((g198) & (g339) & (g345) & (!g358)) + ((g198) & (g339) & (g345) & (g358)));
	assign g373 = (((!g229) & (!g255) & (!g341) & (g342) & (g344) & (!g358)) + ((!g229) & (!g255) & (g341) & (!g342) & (!g344) & (!g358)) + ((!g229) & (!g255) & (g341) & (!g342) & (!g344) & (g358)) + ((!g229) & (!g255) & (g341) & (!g342) & (g344) & (!g358)) + ((!g229) & (!g255) & (g341) & (!g342) & (g344) & (g358)) + ((!g229) & (!g255) & (g341) & (g342) & (!g344) & (!g358)) + ((!g229) & (!g255) & (g341) & (g342) & (!g344) & (g358)) + ((!g229) & (!g255) & (g341) & (g342) & (g344) & (g358)) + ((!g229) & (g255) & (!g341) & (!g342) & (g344) & (!g358)) + ((!g229) & (g255) & (!g341) & (g342) & (!g344) & (!g358)) + ((!g229) & (g255) & (!g341) & (g342) & (g344) & (!g358)) + ((!g229) & (g255) & (g341) & (!g342) & (!g344) & (!g358)) + ((!g229) & (g255) & (g341) & (!g342) & (!g344) & (g358)) + ((!g229) & (g255) & (g341) & (!g342) & (g344) & (g358)) + ((!g229) & (g255) & (g341) & (g342) & (!g344) & (g358)) + ((!g229) & (g255) & (g341) & (g342) & (g344) & (g358)) + ((g229) & (!g255) & (!g341) & (!g342) & (!g344) & (!g358)) + ((g229) & (!g255) & (!g341) & (!g342) & (g344) & (!g358)) + ((g229) & (!g255) & (!g341) & (g342) & (!g344) & (!g358)) + ((g229) & (!g255) & (g341) & (!g342) & (!g344) & (g358)) + ((g229) & (!g255) & (g341) & (!g342) & (g344) & (g358)) + ((g229) & (!g255) & (g341) & (g342) & (!g344) & (g358)) + ((g229) & (!g255) & (g341) & (g342) & (g344) & (!g358)) + ((g229) & (!g255) & (g341) & (g342) & (g344) & (g358)) + ((g229) & (g255) & (!g341) & (!g342) & (!g344) & (!g358)) + ((g229) & (g255) & (g341) & (!g342) & (!g344) & (g358)) + ((g229) & (g255) & (g341) & (!g342) & (g344) & (!g358)) + ((g229) & (g255) & (g341) & (!g342) & (g344) & (g358)) + ((g229) & (g255) & (g341) & (g342) & (!g344) & (!g358)) + ((g229) & (g255) & (g341) & (g342) & (!g344) & (g358)) + ((g229) & (g255) & (g341) & (g342) & (g344) & (!g358)) + ((g229) & (g255) & (g341) & (g342) & (g344) & (g358)));
	assign g374 = (((!g255) & (!g342) & (g344) & (!g358)) + ((!g255) & (g342) & (!g344) & (!g358)) + ((!g255) & (g342) & (!g344) & (g358)) + ((!g255) & (g342) & (g344) & (g358)) + ((g255) & (!g342) & (!g344) & (!g358)) + ((g255) & (g342) & (!g344) & (g358)) + ((g255) & (g342) & (g344) & (!g358)) + ((g255) & (g342) & (g344) & (g358)));
	assign g375 = (((!g290) & (!ax90x) & (!ax91x) & (!g319) & (!g343) & (g358)) + ((!g290) & (!ax90x) & (!ax91x) & (!g319) & (g343) & (!g358)) + ((!g290) & (!ax90x) & (!ax91x) & (!g319) & (g343) & (g358)) + ((!g290) & (!ax90x) & (!ax91x) & (g319) & (!g343) & (!g358)) + ((!g290) & (!ax90x) & (ax91x) & (!g319) & (!g343) & (!g358)) + ((!g290) & (!ax90x) & (ax91x) & (g319) & (!g343) & (g358)) + ((!g290) & (!ax90x) & (ax91x) & (g319) & (g343) & (!g358)) + ((!g290) & (!ax90x) & (ax91x) & (g319) & (g343) & (g358)) + ((!g290) & (ax90x) & (!ax91x) & (g319) & (!g343) & (!g358)) + ((!g290) & (ax90x) & (!ax91x) & (g319) & (g343) & (!g358)) + ((!g290) & (ax90x) & (ax91x) & (!g319) & (!g343) & (!g358)) + ((!g290) & (ax90x) & (ax91x) & (!g319) & (!g343) & (g358)) + ((!g290) & (ax90x) & (ax91x) & (!g319) & (g343) & (!g358)) + ((!g290) & (ax90x) & (ax91x) & (!g319) & (g343) & (g358)) + ((!g290) & (ax90x) & (ax91x) & (g319) & (!g343) & (g358)) + ((!g290) & (ax90x) & (ax91x) & (g319) & (g343) & (g358)) + ((g290) & (!ax90x) & (!ax91x) & (!g319) & (!g343) & (!g358)) + ((g290) & (!ax90x) & (!ax91x) & (!g319) & (!g343) & (g358)) + ((g290) & (!ax90x) & (!ax91x) & (!g319) & (g343) & (g358)) + ((g290) & (!ax90x) & (!ax91x) & (g319) & (g343) & (!g358)) + ((g290) & (!ax90x) & (ax91x) & (!g319) & (g343) & (!g358)) + ((g290) & (!ax90x) & (ax91x) & (g319) & (!g343) & (!g358)) + ((g290) & (!ax90x) & (ax91x) & (g319) & (!g343) & (g358)) + ((g290) & (!ax90x) & (ax91x) & (g319) & (g343) & (g358)) + ((g290) & (ax90x) & (!ax91x) & (!g319) & (!g343) & (!g358)) + ((g290) & (ax90x) & (!ax91x) & (!g319) & (g343) & (!g358)) + ((g290) & (ax90x) & (ax91x) & (!g319) & (!g343) & (g358)) + ((g290) & (ax90x) & (ax91x) & (!g319) & (g343) & (g358)) + ((g290) & (ax90x) & (ax91x) & (g319) & (!g343) & (!g358)) + ((g290) & (ax90x) & (ax91x) & (g319) & (!g343) & (g358)) + ((g290) & (ax90x) & (ax91x) & (g319) & (g343) & (!g358)) + ((g290) & (ax90x) & (ax91x) & (g319) & (g343) & (g358)));
	assign g376 = (((!ax90x) & (!g319) & (!g343) & (g358)) + ((!ax90x) & (!g319) & (g343) & (!g358)) + ((!ax90x) & (!g319) & (g343) & (g358)) + ((!ax90x) & (g319) & (g343) & (!g358)) + ((ax90x) & (!g319) & (!g343) & (!g358)) + ((ax90x) & (g319) & (!g343) & (!g358)) + ((ax90x) & (g319) & (!g343) & (g358)) + ((ax90x) & (g319) & (g343) & (g358)));
	assign g377 = (((!ax86x) & (!ax87x)));
	assign g378 = (((!g319) & (!ax88x) & (!ax89x) & (!g358) & (!g377)) + ((!g319) & (!ax88x) & (ax89x) & (g358) & (!g377)) + ((!g319) & (ax88x) & (ax89x) & (g358) & (!g377)) + ((!g319) & (ax88x) & (ax89x) & (g358) & (g377)) + ((g319) & (!ax88x) & (!ax89x) & (!g358) & (!g377)) + ((g319) & (!ax88x) & (!ax89x) & (!g358) & (g377)) + ((g319) & (!ax88x) & (!ax89x) & (g358) & (!g377)) + ((g319) & (!ax88x) & (ax89x) & (!g358) & (!g377)) + ((g319) & (!ax88x) & (ax89x) & (g358) & (!g377)) + ((g319) & (!ax88x) & (ax89x) & (g358) & (g377)) + ((g319) & (ax88x) & (!ax89x) & (g358) & (!g377)) + ((g319) & (ax88x) & (!ax89x) & (g358) & (g377)) + ((g319) & (ax88x) & (ax89x) & (!g358) & (!g377)) + ((g319) & (ax88x) & (ax89x) & (!g358) & (g377)) + ((g319) & (ax88x) & (ax89x) & (g358) & (!g377)) + ((g319) & (ax88x) & (ax89x) & (g358) & (g377)));
	assign g379 = (((!g255) & (!g290) & (g375) & (g376) & (g378)) + ((!g255) & (g290) & (g375) & (!g376) & (g378)) + ((!g255) & (g290) & (g375) & (g376) & (!g378)) + ((!g255) & (g290) & (g375) & (g376) & (g378)) + ((g255) & (!g290) & (!g375) & (g376) & (g378)) + ((g255) & (!g290) & (g375) & (!g376) & (!g378)) + ((g255) & (!g290) & (g375) & (!g376) & (g378)) + ((g255) & (!g290) & (g375) & (g376) & (!g378)) + ((g255) & (!g290) & (g375) & (g376) & (g378)) + ((g255) & (g290) & (!g375) & (!g376) & (g378)) + ((g255) & (g290) & (!g375) & (g376) & (!g378)) + ((g255) & (g290) & (!g375) & (g376) & (g378)) + ((g255) & (g290) & (g375) & (!g376) & (!g378)) + ((g255) & (g290) & (g375) & (!g376) & (g378)) + ((g255) & (g290) & (g375) & (g376) & (!g378)) + ((g255) & (g290) & (g375) & (g376) & (g378)));
	assign g380 = (((!g198) & (!g229) & (g373) & (g374) & (g379)) + ((!g198) & (g229) & (g373) & (!g374) & (g379)) + ((!g198) & (g229) & (g373) & (g374) & (!g379)) + ((!g198) & (g229) & (g373) & (g374) & (g379)) + ((g198) & (!g229) & (!g373) & (g374) & (g379)) + ((g198) & (!g229) & (g373) & (!g374) & (!g379)) + ((g198) & (!g229) & (g373) & (!g374) & (g379)) + ((g198) & (!g229) & (g373) & (g374) & (!g379)) + ((g198) & (!g229) & (g373) & (g374) & (g379)) + ((g198) & (g229) & (!g373) & (!g374) & (g379)) + ((g198) & (g229) & (!g373) & (g374) & (!g379)) + ((g198) & (g229) & (!g373) & (g374) & (g379)) + ((g198) & (g229) & (g373) & (!g374) & (!g379)) + ((g198) & (g229) & (g373) & (!g374) & (g379)) + ((g198) & (g229) & (g373) & (g374) & (!g379)) + ((g198) & (g229) & (g373) & (g374) & (g379)));
	assign g381 = (((!g147) & (!g174) & (g371) & (g372) & (g380)) + ((!g147) & (g174) & (g371) & (!g372) & (g380)) + ((!g147) & (g174) & (g371) & (g372) & (!g380)) + ((!g147) & (g174) & (g371) & (g372) & (g380)) + ((g147) & (!g174) & (!g371) & (g372) & (g380)) + ((g147) & (!g174) & (g371) & (!g372) & (!g380)) + ((g147) & (!g174) & (g371) & (!g372) & (g380)) + ((g147) & (!g174) & (g371) & (g372) & (!g380)) + ((g147) & (!g174) & (g371) & (g372) & (g380)) + ((g147) & (g174) & (!g371) & (!g372) & (g380)) + ((g147) & (g174) & (!g371) & (g372) & (!g380)) + ((g147) & (g174) & (!g371) & (g372) & (g380)) + ((g147) & (g174) & (g371) & (!g372) & (!g380)) + ((g147) & (g174) & (g371) & (!g372) & (g380)) + ((g147) & (g174) & (g371) & (g372) & (!g380)) + ((g147) & (g174) & (g371) & (g372) & (g380)));
	assign g382 = (((!g104) & (!g127) & (g369) & (g370) & (g381)) + ((!g104) & (g127) & (g369) & (!g370) & (g381)) + ((!g104) & (g127) & (g369) & (g370) & (!g381)) + ((!g104) & (g127) & (g369) & (g370) & (g381)) + ((g104) & (!g127) & (!g369) & (g370) & (g381)) + ((g104) & (!g127) & (g369) & (!g370) & (!g381)) + ((g104) & (!g127) & (g369) & (!g370) & (g381)) + ((g104) & (!g127) & (g369) & (g370) & (!g381)) + ((g104) & (!g127) & (g369) & (g370) & (g381)) + ((g104) & (g127) & (!g369) & (!g370) & (g381)) + ((g104) & (g127) & (!g369) & (g370) & (!g381)) + ((g104) & (g127) & (!g369) & (g370) & (g381)) + ((g104) & (g127) & (g369) & (!g370) & (!g381)) + ((g104) & (g127) & (g369) & (!g370) & (g381)) + ((g104) & (g127) & (g369) & (g370) & (!g381)) + ((g104) & (g127) & (g369) & (g370) & (g381)));
	assign g383 = (((!g68) & (!g87) & (g367) & (g368) & (g382)) + ((!g68) & (g87) & (g367) & (!g368) & (g382)) + ((!g68) & (g87) & (g367) & (g368) & (!g382)) + ((!g68) & (g87) & (g367) & (g368) & (g382)) + ((g68) & (!g87) & (!g367) & (g368) & (g382)) + ((g68) & (!g87) & (g367) & (!g368) & (!g382)) + ((g68) & (!g87) & (g367) & (!g368) & (g382)) + ((g68) & (!g87) & (g367) & (g368) & (!g382)) + ((g68) & (!g87) & (g367) & (g368) & (g382)) + ((g68) & (g87) & (!g367) & (!g368) & (g382)) + ((g68) & (g87) & (!g367) & (g368) & (!g382)) + ((g68) & (g87) & (!g367) & (g368) & (g382)) + ((g68) & (g87) & (g367) & (!g368) & (!g382)) + ((g68) & (g87) & (g367) & (!g368) & (g382)) + ((g68) & (g87) & (g367) & (g368) & (!g382)) + ((g68) & (g87) & (g367) & (g368) & (g382)));
	assign g384 = (((!g39) & (!g54) & (g365) & (g366) & (g383)) + ((!g39) & (g54) & (g365) & (!g366) & (g383)) + ((!g39) & (g54) & (g365) & (g366) & (!g383)) + ((!g39) & (g54) & (g365) & (g366) & (g383)) + ((g39) & (!g54) & (!g365) & (g366) & (g383)) + ((g39) & (!g54) & (g365) & (!g366) & (!g383)) + ((g39) & (!g54) & (g365) & (!g366) & (g383)) + ((g39) & (!g54) & (g365) & (g366) & (!g383)) + ((g39) & (!g54) & (g365) & (g366) & (g383)) + ((g39) & (g54) & (!g365) & (!g366) & (g383)) + ((g39) & (g54) & (!g365) & (g366) & (!g383)) + ((g39) & (g54) & (!g365) & (g366) & (g383)) + ((g39) & (g54) & (g365) & (!g366) & (!g383)) + ((g39) & (g54) & (g365) & (!g366) & (g383)) + ((g39) & (g54) & (g365) & (g366) & (!g383)) + ((g39) & (g54) & (g365) & (g366) & (g383)));
	assign g385 = (((!g18) & (!g27) & (g363) & (g364) & (g384)) + ((!g18) & (g27) & (g363) & (!g364) & (g384)) + ((!g18) & (g27) & (g363) & (g364) & (!g384)) + ((!g18) & (g27) & (g363) & (g364) & (g384)) + ((g18) & (!g27) & (!g363) & (g364) & (g384)) + ((g18) & (!g27) & (g363) & (!g364) & (!g384)) + ((g18) & (!g27) & (g363) & (!g364) & (g384)) + ((g18) & (!g27) & (g363) & (g364) & (!g384)) + ((g18) & (!g27) & (g363) & (g364) & (g384)) + ((g18) & (g27) & (!g363) & (!g364) & (g384)) + ((g18) & (g27) & (!g363) & (g364) & (!g384)) + ((g18) & (g27) & (!g363) & (g364) & (g384)) + ((g18) & (g27) & (g363) & (!g364) & (!g384)) + ((g18) & (g27) & (g363) & (!g364) & (g384)) + ((g18) & (g27) & (g363) & (g364) & (!g384)) + ((g18) & (g27) & (g363) & (g364) & (g384)));
	assign g386 = (((!g2) & (!g8) & (g361) & (g362) & (g385)) + ((!g2) & (g8) & (g361) & (!g362) & (g385)) + ((!g2) & (g8) & (g361) & (g362) & (!g385)) + ((!g2) & (g8) & (g361) & (g362) & (g385)) + ((g2) & (!g8) & (!g361) & (g362) & (g385)) + ((g2) & (!g8) & (g361) & (!g362) & (!g385)) + ((g2) & (!g8) & (g361) & (!g362) & (g385)) + ((g2) & (!g8) & (g361) & (g362) & (!g385)) + ((g2) & (!g8) & (g361) & (g362) & (g385)) + ((g2) & (g8) & (!g361) & (!g362) & (g385)) + ((g2) & (g8) & (!g361) & (g362) & (!g385)) + ((g2) & (g8) & (!g361) & (g362) & (g385)) + ((g2) & (g8) & (g361) & (!g362) & (!g385)) + ((g2) & (g8) & (g361) & (!g362) & (g385)) + ((g2) & (g8) & (g361) & (g362) & (!g385)) + ((g2) & (g8) & (g361) & (g362) & (g385)));
	assign g387 = (((!g2) & (!g321) & (g351) & (!g358)) + ((!g2) & (g321) & (!g351) & (!g358)) + ((!g2) & (g321) & (!g351) & (g358)) + ((!g2) & (g321) & (g351) & (g358)) + ((g2) & (!g321) & (!g351) & (!g358)) + ((g2) & (g321) & (!g351) & (g358)) + ((g2) & (g321) & (g351) & (!g358)) + ((g2) & (g321) & (g351) & (g358)));
	assign g388 = (((!g1) & (!g320) & (!g354) & (!g356) & (g357)) + ((!g1) & (!g320) & (!g354) & (g356) & (!g357)) + ((!g1) & (!g320) & (!g354) & (g356) & (g357)) + ((!g1) & (g320) & (g354) & (!g356) & (!g357)) + ((!g1) & (g320) & (g354) & (!g356) & (g357)) + ((!g1) & (g320) & (g354) & (g356) & (!g357)) + ((!g1) & (g320) & (g354) & (g356) & (g357)) + ((g1) & (!g320) & (!g354) & (!g356) & (g357)) + ((g1) & (!g320) & (!g354) & (g356) & (g357)) + ((g1) & (g320) & (g354) & (!g356) & (!g357)) + ((g1) & (g320) & (g354) & (!g356) & (g357)) + ((g1) & (g320) & (g354) & (g356) & (!g357)) + ((g1) & (g320) & (g354) & (g356) & (g357)));
	assign g389 = (((!g4) & (!g1) & (!g360) & (!g386) & (!g387) & (!g388)) + ((!g4) & (g1) & (!g360) & (!g386) & (!g387) & (!g388)) + ((!g4) & (g1) & (!g360) & (!g386) & (!g387) & (g388)) + ((!g4) & (g1) & (!g360) & (!g386) & (g387) & (!g388)) + ((!g4) & (g1) & (!g360) & (!g386) & (g387) & (g388)) + ((!g4) & (g1) & (!g360) & (g386) & (!g387) & (!g388)) + ((!g4) & (g1) & (!g360) & (g386) & (!g387) & (g388)) + ((!g4) & (g1) & (!g360) & (g386) & (g387) & (!g388)) + ((!g4) & (g1) & (!g360) & (g386) & (g387) & (g388)) + ((!g4) & (g1) & (g360) & (!g386) & (!g387) & (!g388)) + ((!g4) & (g1) & (g360) & (!g386) & (!g387) & (g388)) + ((g4) & (!g1) & (!g360) & (!g386) & (!g387) & (!g388)) + ((g4) & (!g1) & (!g360) & (!g386) & (g387) & (!g388)) + ((g4) & (!g1) & (!g360) & (g386) & (!g387) & (!g388)) + ((g4) & (g1) & (!g360) & (!g386) & (!g387) & (!g388)) + ((g4) & (g1) & (!g360) & (!g386) & (!g387) & (g388)) + ((g4) & (g1) & (!g360) & (!g386) & (g387) & (!g388)) + ((g4) & (g1) & (!g360) & (!g386) & (g387) & (g388)) + ((g4) & (g1) & (!g360) & (g386) & (!g387) & (!g388)) + ((g4) & (g1) & (!g360) & (g386) & (!g387) & (g388)) + ((g4) & (g1) & (!g360) & (g386) & (g387) & (!g388)) + ((g4) & (g1) & (!g360) & (g386) & (g387) & (g388)) + ((g4) & (g1) & (g360) & (!g386) & (!g387) & (!g388)) + ((g4) & (g1) & (g360) & (!g386) & (!g387) & (g388)) + ((g4) & (g1) & (g360) & (!g386) & (g387) & (!g388)) + ((g4) & (g1) & (g360) & (!g386) & (g387) & (g388)) + ((g4) & (g1) & (g360) & (g386) & (!g387) & (!g388)) + ((g4) & (g1) & (g360) & (g386) & (!g387) & (g388)));
	assign g390 = (((!g359) & (g389)));
	assign g391 = (((!g4) & (!g386) & (!g387) & (!g359) & (!g389)) + ((!g4) & (!g386) & (!g387) & (g359) & (!g389)) + ((!g4) & (!g386) & (!g387) & (g359) & (g389)) + ((!g4) & (!g386) & (g387) & (!g359) & (g389)) + ((!g4) & (g386) & (g387) & (!g359) & (!g389)) + ((!g4) & (g386) & (g387) & (!g359) & (g389)) + ((!g4) & (g386) & (g387) & (g359) & (!g389)) + ((!g4) & (g386) & (g387) & (g359) & (g389)) + ((g4) & (!g386) & (g387) & (!g359) & (!g389)) + ((g4) & (!g386) & (g387) & (!g359) & (g389)) + ((g4) & (!g386) & (g387) & (g359) & (!g389)) + ((g4) & (!g386) & (g387) & (g359) & (g389)) + ((g4) & (g386) & (!g387) & (!g359) & (!g389)) + ((g4) & (g386) & (!g387) & (g359) & (!g389)) + ((g4) & (g386) & (!g387) & (g359) & (g389)) + ((g4) & (g386) & (g387) & (!g359) & (g389)));
	assign g392 = (((!g8) & (!g362) & (g385) & (!g359) & (!g389)) + ((!g8) & (!g362) & (g385) & (g359) & (!g389)) + ((!g8) & (!g362) & (g385) & (g359) & (g389)) + ((!g8) & (g362) & (!g385) & (!g359) & (!g389)) + ((!g8) & (g362) & (!g385) & (!g359) & (g389)) + ((!g8) & (g362) & (!g385) & (g359) & (!g389)) + ((!g8) & (g362) & (!g385) & (g359) & (g389)) + ((!g8) & (g362) & (g385) & (!g359) & (g389)) + ((g8) & (!g362) & (!g385) & (!g359) & (!g389)) + ((g8) & (!g362) & (!g385) & (g359) & (!g389)) + ((g8) & (!g362) & (!g385) & (g359) & (g389)) + ((g8) & (g362) & (!g385) & (!g359) & (g389)) + ((g8) & (g362) & (g385) & (!g359) & (!g389)) + ((g8) & (g362) & (g385) & (!g359) & (g389)) + ((g8) & (g362) & (g385) & (g359) & (!g389)) + ((g8) & (g362) & (g385) & (g359) & (g389)));
	assign g393 = (((!g18) & (!g27) & (g364) & (g384)) + ((!g18) & (g27) & (!g364) & (g384)) + ((!g18) & (g27) & (g364) & (!g384)) + ((!g18) & (g27) & (g364) & (g384)) + ((g18) & (!g27) & (!g364) & (!g384)) + ((g18) & (!g27) & (!g364) & (g384)) + ((g18) & (!g27) & (g364) & (!g384)) + ((g18) & (g27) & (!g364) & (!g384)));
	assign g394 = (((!g363) & (!g359) & (!g389) & (g393)) + ((!g363) & (g359) & (!g389) & (g393)) + ((!g363) & (g359) & (g389) & (g393)) + ((g363) & (!g359) & (!g389) & (!g393)) + ((g363) & (!g359) & (g389) & (!g393)) + ((g363) & (!g359) & (g389) & (g393)) + ((g363) & (g359) & (!g389) & (!g393)) + ((g363) & (g359) & (g389) & (!g393)));
	assign g395 = (((!g27) & (!g364) & (g384) & (!g359) & (!g389)) + ((!g27) & (!g364) & (g384) & (g359) & (!g389)) + ((!g27) & (!g364) & (g384) & (g359) & (g389)) + ((!g27) & (g364) & (!g384) & (!g359) & (!g389)) + ((!g27) & (g364) & (!g384) & (!g359) & (g389)) + ((!g27) & (g364) & (!g384) & (g359) & (!g389)) + ((!g27) & (g364) & (!g384) & (g359) & (g389)) + ((!g27) & (g364) & (g384) & (!g359) & (g389)) + ((g27) & (!g364) & (!g384) & (!g359) & (!g389)) + ((g27) & (!g364) & (!g384) & (g359) & (!g389)) + ((g27) & (!g364) & (!g384) & (g359) & (g389)) + ((g27) & (g364) & (!g384) & (!g359) & (g389)) + ((g27) & (g364) & (g384) & (!g359) & (!g389)) + ((g27) & (g364) & (g384) & (!g359) & (g389)) + ((g27) & (g364) & (g384) & (g359) & (!g389)) + ((g27) & (g364) & (g384) & (g359) & (g389)));
	assign g396 = (((!g39) & (!g54) & (g366) & (g383)) + ((!g39) & (g54) & (!g366) & (g383)) + ((!g39) & (g54) & (g366) & (!g383)) + ((!g39) & (g54) & (g366) & (g383)) + ((g39) & (!g54) & (!g366) & (!g383)) + ((g39) & (!g54) & (!g366) & (g383)) + ((g39) & (!g54) & (g366) & (!g383)) + ((g39) & (g54) & (!g366) & (!g383)));
	assign g397 = (((!g365) & (!g359) & (!g389) & (g396)) + ((!g365) & (g359) & (!g389) & (g396)) + ((!g365) & (g359) & (g389) & (g396)) + ((g365) & (!g359) & (!g389) & (!g396)) + ((g365) & (!g359) & (g389) & (!g396)) + ((g365) & (!g359) & (g389) & (g396)) + ((g365) & (g359) & (!g389) & (!g396)) + ((g365) & (g359) & (g389) & (!g396)));
	assign g398 = (((!g54) & (!g366) & (g383) & (!g359) & (!g389)) + ((!g54) & (!g366) & (g383) & (g359) & (!g389)) + ((!g54) & (!g366) & (g383) & (g359) & (g389)) + ((!g54) & (g366) & (!g383) & (!g359) & (!g389)) + ((!g54) & (g366) & (!g383) & (!g359) & (g389)) + ((!g54) & (g366) & (!g383) & (g359) & (!g389)) + ((!g54) & (g366) & (!g383) & (g359) & (g389)) + ((!g54) & (g366) & (g383) & (!g359) & (g389)) + ((g54) & (!g366) & (!g383) & (!g359) & (!g389)) + ((g54) & (!g366) & (!g383) & (g359) & (!g389)) + ((g54) & (!g366) & (!g383) & (g359) & (g389)) + ((g54) & (g366) & (!g383) & (!g359) & (g389)) + ((g54) & (g366) & (g383) & (!g359) & (!g389)) + ((g54) & (g366) & (g383) & (!g359) & (g389)) + ((g54) & (g366) & (g383) & (g359) & (!g389)) + ((g54) & (g366) & (g383) & (g359) & (g389)));
	assign g399 = (((!g68) & (!g87) & (g368) & (g382)) + ((!g68) & (g87) & (!g368) & (g382)) + ((!g68) & (g87) & (g368) & (!g382)) + ((!g68) & (g87) & (g368) & (g382)) + ((g68) & (!g87) & (!g368) & (!g382)) + ((g68) & (!g87) & (!g368) & (g382)) + ((g68) & (!g87) & (g368) & (!g382)) + ((g68) & (g87) & (!g368) & (!g382)));
	assign g400 = (((!g367) & (!g359) & (!g389) & (g399)) + ((!g367) & (g359) & (!g389) & (g399)) + ((!g367) & (g359) & (g389) & (g399)) + ((g367) & (!g359) & (!g389) & (!g399)) + ((g367) & (!g359) & (g389) & (!g399)) + ((g367) & (!g359) & (g389) & (g399)) + ((g367) & (g359) & (!g389) & (!g399)) + ((g367) & (g359) & (g389) & (!g399)));
	assign g401 = (((!g87) & (!g368) & (g382) & (!g359) & (!g389)) + ((!g87) & (!g368) & (g382) & (g359) & (!g389)) + ((!g87) & (!g368) & (g382) & (g359) & (g389)) + ((!g87) & (g368) & (!g382) & (!g359) & (!g389)) + ((!g87) & (g368) & (!g382) & (!g359) & (g389)) + ((!g87) & (g368) & (!g382) & (g359) & (!g389)) + ((!g87) & (g368) & (!g382) & (g359) & (g389)) + ((!g87) & (g368) & (g382) & (!g359) & (g389)) + ((g87) & (!g368) & (!g382) & (!g359) & (!g389)) + ((g87) & (!g368) & (!g382) & (g359) & (!g389)) + ((g87) & (!g368) & (!g382) & (g359) & (g389)) + ((g87) & (g368) & (!g382) & (!g359) & (g389)) + ((g87) & (g368) & (g382) & (!g359) & (!g389)) + ((g87) & (g368) & (g382) & (!g359) & (g389)) + ((g87) & (g368) & (g382) & (g359) & (!g389)) + ((g87) & (g368) & (g382) & (g359) & (g389)));
	assign g402 = (((!g104) & (!g127) & (g370) & (g381)) + ((!g104) & (g127) & (!g370) & (g381)) + ((!g104) & (g127) & (g370) & (!g381)) + ((!g104) & (g127) & (g370) & (g381)) + ((g104) & (!g127) & (!g370) & (!g381)) + ((g104) & (!g127) & (!g370) & (g381)) + ((g104) & (!g127) & (g370) & (!g381)) + ((g104) & (g127) & (!g370) & (!g381)));
	assign g403 = (((!g369) & (!g359) & (!g389) & (g402)) + ((!g369) & (g359) & (!g389) & (g402)) + ((!g369) & (g359) & (g389) & (g402)) + ((g369) & (!g359) & (!g389) & (!g402)) + ((g369) & (!g359) & (g389) & (!g402)) + ((g369) & (!g359) & (g389) & (g402)) + ((g369) & (g359) & (!g389) & (!g402)) + ((g369) & (g359) & (g389) & (!g402)));
	assign g404 = (((!g127) & (!g370) & (g381) & (!g359) & (!g389)) + ((!g127) & (!g370) & (g381) & (g359) & (!g389)) + ((!g127) & (!g370) & (g381) & (g359) & (g389)) + ((!g127) & (g370) & (!g381) & (!g359) & (!g389)) + ((!g127) & (g370) & (!g381) & (!g359) & (g389)) + ((!g127) & (g370) & (!g381) & (g359) & (!g389)) + ((!g127) & (g370) & (!g381) & (g359) & (g389)) + ((!g127) & (g370) & (g381) & (!g359) & (g389)) + ((g127) & (!g370) & (!g381) & (!g359) & (!g389)) + ((g127) & (!g370) & (!g381) & (g359) & (!g389)) + ((g127) & (!g370) & (!g381) & (g359) & (g389)) + ((g127) & (g370) & (!g381) & (!g359) & (g389)) + ((g127) & (g370) & (g381) & (!g359) & (!g389)) + ((g127) & (g370) & (g381) & (!g359) & (g389)) + ((g127) & (g370) & (g381) & (g359) & (!g389)) + ((g127) & (g370) & (g381) & (g359) & (g389)));
	assign g405 = (((!g147) & (!g174) & (g372) & (g380)) + ((!g147) & (g174) & (!g372) & (g380)) + ((!g147) & (g174) & (g372) & (!g380)) + ((!g147) & (g174) & (g372) & (g380)) + ((g147) & (!g174) & (!g372) & (!g380)) + ((g147) & (!g174) & (!g372) & (g380)) + ((g147) & (!g174) & (g372) & (!g380)) + ((g147) & (g174) & (!g372) & (!g380)));
	assign g406 = (((!g371) & (!g359) & (!g389) & (g405)) + ((!g371) & (g359) & (!g389) & (g405)) + ((!g371) & (g359) & (g389) & (g405)) + ((g371) & (!g359) & (!g389) & (!g405)) + ((g371) & (!g359) & (g389) & (!g405)) + ((g371) & (!g359) & (g389) & (g405)) + ((g371) & (g359) & (!g389) & (!g405)) + ((g371) & (g359) & (g389) & (!g405)));
	assign g407 = (((!g174) & (!g372) & (g380) & (!g359) & (!g389)) + ((!g174) & (!g372) & (g380) & (g359) & (!g389)) + ((!g174) & (!g372) & (g380) & (g359) & (g389)) + ((!g174) & (g372) & (!g380) & (!g359) & (!g389)) + ((!g174) & (g372) & (!g380) & (!g359) & (g389)) + ((!g174) & (g372) & (!g380) & (g359) & (!g389)) + ((!g174) & (g372) & (!g380) & (g359) & (g389)) + ((!g174) & (g372) & (g380) & (!g359) & (g389)) + ((g174) & (!g372) & (!g380) & (!g359) & (!g389)) + ((g174) & (!g372) & (!g380) & (g359) & (!g389)) + ((g174) & (!g372) & (!g380) & (g359) & (g389)) + ((g174) & (g372) & (!g380) & (!g359) & (g389)) + ((g174) & (g372) & (g380) & (!g359) & (!g389)) + ((g174) & (g372) & (g380) & (!g359) & (g389)) + ((g174) & (g372) & (g380) & (g359) & (!g389)) + ((g174) & (g372) & (g380) & (g359) & (g389)));
	assign g408 = (((!g198) & (!g229) & (g374) & (g379)) + ((!g198) & (g229) & (!g374) & (g379)) + ((!g198) & (g229) & (g374) & (!g379)) + ((!g198) & (g229) & (g374) & (g379)) + ((g198) & (!g229) & (!g374) & (!g379)) + ((g198) & (!g229) & (!g374) & (g379)) + ((g198) & (!g229) & (g374) & (!g379)) + ((g198) & (g229) & (!g374) & (!g379)));
	assign g409 = (((!g373) & (!g359) & (!g389) & (g408)) + ((!g373) & (g359) & (!g389) & (g408)) + ((!g373) & (g359) & (g389) & (g408)) + ((g373) & (!g359) & (!g389) & (!g408)) + ((g373) & (!g359) & (g389) & (!g408)) + ((g373) & (!g359) & (g389) & (g408)) + ((g373) & (g359) & (!g389) & (!g408)) + ((g373) & (g359) & (g389) & (!g408)));
	assign g410 = (((!g229) & (!g374) & (g379) & (!g359) & (!g389)) + ((!g229) & (!g374) & (g379) & (g359) & (!g389)) + ((!g229) & (!g374) & (g379) & (g359) & (g389)) + ((!g229) & (g374) & (!g379) & (!g359) & (!g389)) + ((!g229) & (g374) & (!g379) & (!g359) & (g389)) + ((!g229) & (g374) & (!g379) & (g359) & (!g389)) + ((!g229) & (g374) & (!g379) & (g359) & (g389)) + ((!g229) & (g374) & (g379) & (!g359) & (g389)) + ((g229) & (!g374) & (!g379) & (!g359) & (!g389)) + ((g229) & (!g374) & (!g379) & (g359) & (!g389)) + ((g229) & (!g374) & (!g379) & (g359) & (g389)) + ((g229) & (g374) & (!g379) & (!g359) & (g389)) + ((g229) & (g374) & (g379) & (!g359) & (!g389)) + ((g229) & (g374) & (g379) & (!g359) & (g389)) + ((g229) & (g374) & (g379) & (g359) & (!g389)) + ((g229) & (g374) & (g379) & (g359) & (g389)));
	assign g411 = (((!g255) & (!g290) & (g376) & (g378)) + ((!g255) & (g290) & (!g376) & (g378)) + ((!g255) & (g290) & (g376) & (!g378)) + ((!g255) & (g290) & (g376) & (g378)) + ((g255) & (!g290) & (!g376) & (!g378)) + ((g255) & (!g290) & (!g376) & (g378)) + ((g255) & (!g290) & (g376) & (!g378)) + ((g255) & (g290) & (!g376) & (!g378)));
	assign g412 = (((!g375) & (!g359) & (!g389) & (g411)) + ((!g375) & (g359) & (!g389) & (g411)) + ((!g375) & (g359) & (g389) & (g411)) + ((g375) & (!g359) & (!g389) & (!g411)) + ((g375) & (!g359) & (g389) & (!g411)) + ((g375) & (!g359) & (g389) & (g411)) + ((g375) & (g359) & (!g389) & (!g411)) + ((g375) & (g359) & (g389) & (!g411)));
	assign g413 = (((!g290) & (!g376) & (g378) & (!g359) & (!g389)) + ((!g290) & (!g376) & (g378) & (g359) & (!g389)) + ((!g290) & (!g376) & (g378) & (g359) & (g389)) + ((!g290) & (g376) & (!g378) & (!g359) & (!g389)) + ((!g290) & (g376) & (!g378) & (!g359) & (g389)) + ((!g290) & (g376) & (!g378) & (g359) & (!g389)) + ((!g290) & (g376) & (!g378) & (g359) & (g389)) + ((!g290) & (g376) & (g378) & (!g359) & (g389)) + ((g290) & (!g376) & (!g378) & (!g359) & (!g389)) + ((g290) & (!g376) & (!g378) & (g359) & (!g389)) + ((g290) & (!g376) & (!g378) & (g359) & (g389)) + ((g290) & (g376) & (!g378) & (!g359) & (g389)) + ((g290) & (g376) & (g378) & (!g359) & (!g389)) + ((g290) & (g376) & (g378) & (!g359) & (g389)) + ((g290) & (g376) & (g378) & (g359) & (!g389)) + ((g290) & (g376) & (g378) & (g359) & (g389)));
	assign g414 = (((!g319) & (!ax88x) & (!g358) & (g377)) + ((!g319) & (!ax88x) & (g358) & (g377)) + ((!g319) & (ax88x) & (!g358) & (!g377)) + ((!g319) & (ax88x) & (!g358) & (g377)) + ((g319) & (!ax88x) & (!g358) & (!g377)) + ((g319) & (!ax88x) & (g358) & (!g377)) + ((g319) & (ax88x) & (g358) & (!g377)) + ((g319) & (ax88x) & (g358) & (g377)));
	assign g415 = (((!ax88x) & (!ax89x) & (!g358) & (!g359) & (!g389) & (g414)) + ((!ax88x) & (!ax89x) & (!g358) & (!g359) & (g389) & (!g414)) + ((!ax88x) & (!ax89x) & (!g358) & (!g359) & (g389) & (g414)) + ((!ax88x) & (!ax89x) & (!g358) & (g359) & (!g389) & (g414)) + ((!ax88x) & (!ax89x) & (!g358) & (g359) & (g389) & (g414)) + ((!ax88x) & (!ax89x) & (g358) & (!g359) & (!g389) & (!g414)) + ((!ax88x) & (!ax89x) & (g358) & (g359) & (!g389) & (!g414)) + ((!ax88x) & (!ax89x) & (g358) & (g359) & (g389) & (!g414)) + ((!ax88x) & (ax89x) & (!g358) & (!g359) & (!g389) & (!g414)) + ((!ax88x) & (ax89x) & (!g358) & (g359) & (!g389) & (!g414)) + ((!ax88x) & (ax89x) & (!g358) & (g359) & (g389) & (!g414)) + ((!ax88x) & (ax89x) & (g358) & (!g359) & (!g389) & (g414)) + ((!ax88x) & (ax89x) & (g358) & (!g359) & (g389) & (!g414)) + ((!ax88x) & (ax89x) & (g358) & (!g359) & (g389) & (g414)) + ((!ax88x) & (ax89x) & (g358) & (g359) & (!g389) & (g414)) + ((!ax88x) & (ax89x) & (g358) & (g359) & (g389) & (g414)) + ((ax88x) & (!ax89x) & (!g358) & (!g359) & (!g389) & (!g414)) + ((ax88x) & (!ax89x) & (!g358) & (g359) & (!g389) & (!g414)) + ((ax88x) & (!ax89x) & (!g358) & (g359) & (g389) & (!g414)) + ((ax88x) & (!ax89x) & (g358) & (!g359) & (!g389) & (!g414)) + ((ax88x) & (!ax89x) & (g358) & (g359) & (!g389) & (!g414)) + ((ax88x) & (!ax89x) & (g358) & (g359) & (g389) & (!g414)) + ((ax88x) & (ax89x) & (!g358) & (!g359) & (!g389) & (g414)) + ((ax88x) & (ax89x) & (!g358) & (!g359) & (g389) & (!g414)) + ((ax88x) & (ax89x) & (!g358) & (!g359) & (g389) & (g414)) + ((ax88x) & (ax89x) & (!g358) & (g359) & (!g389) & (g414)) + ((ax88x) & (ax89x) & (!g358) & (g359) & (g389) & (g414)) + ((ax88x) & (ax89x) & (g358) & (!g359) & (!g389) & (g414)) + ((ax88x) & (ax89x) & (g358) & (!g359) & (g389) & (!g414)) + ((ax88x) & (ax89x) & (g358) & (!g359) & (g389) & (g414)) + ((ax88x) & (ax89x) & (g358) & (g359) & (!g389) & (g414)) + ((ax88x) & (ax89x) & (g358) & (g359) & (g389) & (g414)));
	assign g416 = (((!ax88x) & (!g358) & (!g377) & (!g359) & (g389)) + ((!ax88x) & (!g358) & (g377) & (!g359) & (!g389)) + ((!ax88x) & (!g358) & (g377) & (!g359) & (g389)) + ((!ax88x) & (!g358) & (g377) & (g359) & (!g389)) + ((!ax88x) & (!g358) & (g377) & (g359) & (g389)) + ((!ax88x) & (g358) & (g377) & (!g359) & (!g389)) + ((!ax88x) & (g358) & (g377) & (g359) & (!g389)) + ((!ax88x) & (g358) & (g377) & (g359) & (g389)) + ((ax88x) & (!g358) & (!g377) & (!g359) & (!g389)) + ((ax88x) & (!g358) & (!g377) & (g359) & (!g389)) + ((ax88x) & (!g358) & (!g377) & (g359) & (g389)) + ((ax88x) & (g358) & (!g377) & (!g359) & (!g389)) + ((ax88x) & (g358) & (!g377) & (!g359) & (g389)) + ((ax88x) & (g358) & (!g377) & (g359) & (!g389)) + ((ax88x) & (g358) & (!g377) & (g359) & (g389)) + ((ax88x) & (g358) & (g377) & (!g359) & (g389)));
	assign g417 = (((!ax84x) & (!ax85x)));
	assign g418 = (((!g358) & (!ax86x) & (!ax87x) & (!g359) & (!g389) & (!g417)) + ((!g358) & (!ax86x) & (!ax87x) & (g359) & (!g389) & (!g417)) + ((!g358) & (!ax86x) & (!ax87x) & (g359) & (g389) & (!g417)) + ((!g358) & (!ax86x) & (ax87x) & (!g359) & (g389) & (!g417)) + ((!g358) & (ax86x) & (ax87x) & (!g359) & (g389) & (!g417)) + ((!g358) & (ax86x) & (ax87x) & (!g359) & (g389) & (g417)) + ((g358) & (!ax86x) & (!ax87x) & (!g359) & (!g389) & (!g417)) + ((g358) & (!ax86x) & (!ax87x) & (!g359) & (!g389) & (g417)) + ((g358) & (!ax86x) & (!ax87x) & (!g359) & (g389) & (!g417)) + ((g358) & (!ax86x) & (!ax87x) & (g359) & (!g389) & (!g417)) + ((g358) & (!ax86x) & (!ax87x) & (g359) & (!g389) & (g417)) + ((g358) & (!ax86x) & (!ax87x) & (g359) & (g389) & (!g417)) + ((g358) & (!ax86x) & (!ax87x) & (g359) & (g389) & (g417)) + ((g358) & (!ax86x) & (ax87x) & (!g359) & (!g389) & (!g417)) + ((g358) & (!ax86x) & (ax87x) & (!g359) & (g389) & (!g417)) + ((g358) & (!ax86x) & (ax87x) & (!g359) & (g389) & (g417)) + ((g358) & (!ax86x) & (ax87x) & (g359) & (!g389) & (!g417)) + ((g358) & (!ax86x) & (ax87x) & (g359) & (g389) & (!g417)) + ((g358) & (ax86x) & (!ax87x) & (!g359) & (g389) & (!g417)) + ((g358) & (ax86x) & (!ax87x) & (!g359) & (g389) & (g417)) + ((g358) & (ax86x) & (ax87x) & (!g359) & (!g389) & (!g417)) + ((g358) & (ax86x) & (ax87x) & (!g359) & (!g389) & (g417)) + ((g358) & (ax86x) & (ax87x) & (!g359) & (g389) & (!g417)) + ((g358) & (ax86x) & (ax87x) & (!g359) & (g389) & (g417)) + ((g358) & (ax86x) & (ax87x) & (g359) & (!g389) & (!g417)) + ((g358) & (ax86x) & (ax87x) & (g359) & (!g389) & (g417)) + ((g358) & (ax86x) & (ax87x) & (g359) & (g389) & (!g417)) + ((g358) & (ax86x) & (ax87x) & (g359) & (g389) & (g417)));
	assign g419 = (((!g290) & (!g319) & (g415) & (g416) & (g418)) + ((!g290) & (g319) & (g415) & (!g416) & (g418)) + ((!g290) & (g319) & (g415) & (g416) & (!g418)) + ((!g290) & (g319) & (g415) & (g416) & (g418)) + ((g290) & (!g319) & (!g415) & (g416) & (g418)) + ((g290) & (!g319) & (g415) & (!g416) & (!g418)) + ((g290) & (!g319) & (g415) & (!g416) & (g418)) + ((g290) & (!g319) & (g415) & (g416) & (!g418)) + ((g290) & (!g319) & (g415) & (g416) & (g418)) + ((g290) & (g319) & (!g415) & (!g416) & (g418)) + ((g290) & (g319) & (!g415) & (g416) & (!g418)) + ((g290) & (g319) & (!g415) & (g416) & (g418)) + ((g290) & (g319) & (g415) & (!g416) & (!g418)) + ((g290) & (g319) & (g415) & (!g416) & (g418)) + ((g290) & (g319) & (g415) & (g416) & (!g418)) + ((g290) & (g319) & (g415) & (g416) & (g418)));
	assign g420 = (((!g229) & (!g255) & (g412) & (g413) & (g419)) + ((!g229) & (g255) & (g412) & (!g413) & (g419)) + ((!g229) & (g255) & (g412) & (g413) & (!g419)) + ((!g229) & (g255) & (g412) & (g413) & (g419)) + ((g229) & (!g255) & (!g412) & (g413) & (g419)) + ((g229) & (!g255) & (g412) & (!g413) & (!g419)) + ((g229) & (!g255) & (g412) & (!g413) & (g419)) + ((g229) & (!g255) & (g412) & (g413) & (!g419)) + ((g229) & (!g255) & (g412) & (g413) & (g419)) + ((g229) & (g255) & (!g412) & (!g413) & (g419)) + ((g229) & (g255) & (!g412) & (g413) & (!g419)) + ((g229) & (g255) & (!g412) & (g413) & (g419)) + ((g229) & (g255) & (g412) & (!g413) & (!g419)) + ((g229) & (g255) & (g412) & (!g413) & (g419)) + ((g229) & (g255) & (g412) & (g413) & (!g419)) + ((g229) & (g255) & (g412) & (g413) & (g419)));
	assign g421 = (((!g174) & (!g198) & (g409) & (g410) & (g420)) + ((!g174) & (g198) & (g409) & (!g410) & (g420)) + ((!g174) & (g198) & (g409) & (g410) & (!g420)) + ((!g174) & (g198) & (g409) & (g410) & (g420)) + ((g174) & (!g198) & (!g409) & (g410) & (g420)) + ((g174) & (!g198) & (g409) & (!g410) & (!g420)) + ((g174) & (!g198) & (g409) & (!g410) & (g420)) + ((g174) & (!g198) & (g409) & (g410) & (!g420)) + ((g174) & (!g198) & (g409) & (g410) & (g420)) + ((g174) & (g198) & (!g409) & (!g410) & (g420)) + ((g174) & (g198) & (!g409) & (g410) & (!g420)) + ((g174) & (g198) & (!g409) & (g410) & (g420)) + ((g174) & (g198) & (g409) & (!g410) & (!g420)) + ((g174) & (g198) & (g409) & (!g410) & (g420)) + ((g174) & (g198) & (g409) & (g410) & (!g420)) + ((g174) & (g198) & (g409) & (g410) & (g420)));
	assign g422 = (((!g127) & (!g147) & (g406) & (g407) & (g421)) + ((!g127) & (g147) & (g406) & (!g407) & (g421)) + ((!g127) & (g147) & (g406) & (g407) & (!g421)) + ((!g127) & (g147) & (g406) & (g407) & (g421)) + ((g127) & (!g147) & (!g406) & (g407) & (g421)) + ((g127) & (!g147) & (g406) & (!g407) & (!g421)) + ((g127) & (!g147) & (g406) & (!g407) & (g421)) + ((g127) & (!g147) & (g406) & (g407) & (!g421)) + ((g127) & (!g147) & (g406) & (g407) & (g421)) + ((g127) & (g147) & (!g406) & (!g407) & (g421)) + ((g127) & (g147) & (!g406) & (g407) & (!g421)) + ((g127) & (g147) & (!g406) & (g407) & (g421)) + ((g127) & (g147) & (g406) & (!g407) & (!g421)) + ((g127) & (g147) & (g406) & (!g407) & (g421)) + ((g127) & (g147) & (g406) & (g407) & (!g421)) + ((g127) & (g147) & (g406) & (g407) & (g421)));
	assign g423 = (((!g87) & (!g104) & (g403) & (g404) & (g422)) + ((!g87) & (g104) & (g403) & (!g404) & (g422)) + ((!g87) & (g104) & (g403) & (g404) & (!g422)) + ((!g87) & (g104) & (g403) & (g404) & (g422)) + ((g87) & (!g104) & (!g403) & (g404) & (g422)) + ((g87) & (!g104) & (g403) & (!g404) & (!g422)) + ((g87) & (!g104) & (g403) & (!g404) & (g422)) + ((g87) & (!g104) & (g403) & (g404) & (!g422)) + ((g87) & (!g104) & (g403) & (g404) & (g422)) + ((g87) & (g104) & (!g403) & (!g404) & (g422)) + ((g87) & (g104) & (!g403) & (g404) & (!g422)) + ((g87) & (g104) & (!g403) & (g404) & (g422)) + ((g87) & (g104) & (g403) & (!g404) & (!g422)) + ((g87) & (g104) & (g403) & (!g404) & (g422)) + ((g87) & (g104) & (g403) & (g404) & (!g422)) + ((g87) & (g104) & (g403) & (g404) & (g422)));
	assign g424 = (((!g54) & (!g68) & (g400) & (g401) & (g423)) + ((!g54) & (g68) & (g400) & (!g401) & (g423)) + ((!g54) & (g68) & (g400) & (g401) & (!g423)) + ((!g54) & (g68) & (g400) & (g401) & (g423)) + ((g54) & (!g68) & (!g400) & (g401) & (g423)) + ((g54) & (!g68) & (g400) & (!g401) & (!g423)) + ((g54) & (!g68) & (g400) & (!g401) & (g423)) + ((g54) & (!g68) & (g400) & (g401) & (!g423)) + ((g54) & (!g68) & (g400) & (g401) & (g423)) + ((g54) & (g68) & (!g400) & (!g401) & (g423)) + ((g54) & (g68) & (!g400) & (g401) & (!g423)) + ((g54) & (g68) & (!g400) & (g401) & (g423)) + ((g54) & (g68) & (g400) & (!g401) & (!g423)) + ((g54) & (g68) & (g400) & (!g401) & (g423)) + ((g54) & (g68) & (g400) & (g401) & (!g423)) + ((g54) & (g68) & (g400) & (g401) & (g423)));
	assign g425 = (((!g27) & (!g39) & (g397) & (g398) & (g424)) + ((!g27) & (g39) & (g397) & (!g398) & (g424)) + ((!g27) & (g39) & (g397) & (g398) & (!g424)) + ((!g27) & (g39) & (g397) & (g398) & (g424)) + ((g27) & (!g39) & (!g397) & (g398) & (g424)) + ((g27) & (!g39) & (g397) & (!g398) & (!g424)) + ((g27) & (!g39) & (g397) & (!g398) & (g424)) + ((g27) & (!g39) & (g397) & (g398) & (!g424)) + ((g27) & (!g39) & (g397) & (g398) & (g424)) + ((g27) & (g39) & (!g397) & (!g398) & (g424)) + ((g27) & (g39) & (!g397) & (g398) & (!g424)) + ((g27) & (g39) & (!g397) & (g398) & (g424)) + ((g27) & (g39) & (g397) & (!g398) & (!g424)) + ((g27) & (g39) & (g397) & (!g398) & (g424)) + ((g27) & (g39) & (g397) & (g398) & (!g424)) + ((g27) & (g39) & (g397) & (g398) & (g424)));
	assign g426 = (((!g8) & (!g18) & (g394) & (g395) & (g425)) + ((!g8) & (g18) & (g394) & (!g395) & (g425)) + ((!g8) & (g18) & (g394) & (g395) & (!g425)) + ((!g8) & (g18) & (g394) & (g395) & (g425)) + ((g8) & (!g18) & (!g394) & (g395) & (g425)) + ((g8) & (!g18) & (g394) & (!g395) & (!g425)) + ((g8) & (!g18) & (g394) & (!g395) & (g425)) + ((g8) & (!g18) & (g394) & (g395) & (!g425)) + ((g8) & (!g18) & (g394) & (g395) & (g425)) + ((g8) & (g18) & (!g394) & (!g395) & (g425)) + ((g8) & (g18) & (!g394) & (g395) & (!g425)) + ((g8) & (g18) & (!g394) & (g395) & (g425)) + ((g8) & (g18) & (g394) & (!g395) & (!g425)) + ((g8) & (g18) & (g394) & (!g395) & (g425)) + ((g8) & (g18) & (g394) & (g395) & (!g425)) + ((g8) & (g18) & (g394) & (g395) & (g425)));
	assign g427 = (((!g2) & (!g8) & (g362) & (g385)) + ((!g2) & (g8) & (!g362) & (g385)) + ((!g2) & (g8) & (g362) & (!g385)) + ((!g2) & (g8) & (g362) & (g385)) + ((g2) & (!g8) & (!g362) & (!g385)) + ((g2) & (!g8) & (!g362) & (g385)) + ((g2) & (!g8) & (g362) & (!g385)) + ((g2) & (g8) & (!g362) & (!g385)));
	assign g428 = (((!g361) & (!g359) & (!g389) & (g427)) + ((!g361) & (g359) & (!g389) & (g427)) + ((!g361) & (g359) & (g389) & (g427)) + ((g361) & (!g359) & (!g389) & (!g427)) + ((g361) & (!g359) & (g389) & (!g427)) + ((g361) & (!g359) & (g389) & (g427)) + ((g361) & (g359) & (!g389) & (!g427)) + ((g361) & (g359) & (g389) & (!g427)));
	assign g429 = (((!g4) & (!g2) & (!g392) & (!g426) & (g428)) + ((!g4) & (!g2) & (!g392) & (g426) & (g428)) + ((!g4) & (!g2) & (g392) & (!g426) & (g428)) + ((!g4) & (!g2) & (g392) & (g426) & (!g428)) + ((!g4) & (!g2) & (g392) & (g426) & (g428)) + ((!g4) & (g2) & (!g392) & (!g426) & (g428)) + ((!g4) & (g2) & (!g392) & (g426) & (!g428)) + ((!g4) & (g2) & (!g392) & (g426) & (g428)) + ((!g4) & (g2) & (g392) & (!g426) & (!g428)) + ((!g4) & (g2) & (g392) & (!g426) & (g428)) + ((!g4) & (g2) & (g392) & (g426) & (!g428)) + ((!g4) & (g2) & (g392) & (g426) & (g428)) + ((g4) & (!g2) & (g392) & (g426) & (g428)) + ((g4) & (g2) & (!g392) & (g426) & (g428)) + ((g4) & (g2) & (g392) & (!g426) & (g428)) + ((g4) & (g2) & (g392) & (g426) & (g428)));
	assign g430 = (((!g4) & (!g386) & (g387)) + ((!g4) & (g386) & (!g387)) + ((!g4) & (g386) & (g387)) + ((g4) & (g386) & (g387)));
	assign g431 = (((!g360) & (!g430) & (!g359) & (!g389)) + ((!g360) & (!g430) & (g359) & (!g389)) + ((!g360) & (!g430) & (g359) & (g389)) + ((g360) & (g430) & (!g359) & (!g389)) + ((g360) & (g430) & (!g359) & (g389)) + ((g360) & (g430) & (g359) & (!g389)) + ((g360) & (g430) & (g359) & (g389)));
	assign g432 = (((!g1) & (g360) & (!g430) & (!g359) & (g389)) + ((!g1) & (g360) & (g430) & (!g359) & (g389)) + ((g1) & (!g360) & (g430) & (g359) & (!g389)) + ((g1) & (!g360) & (g430) & (g359) & (g389)) + ((g1) & (g360) & (!g430) & (!g359) & (!g389)) + ((g1) & (g360) & (!g430) & (!g359) & (g389)) + ((g1) & (g360) & (!g430) & (g359) & (!g389)) + ((g1) & (g360) & (!g430) & (g359) & (g389)) + ((g1) & (g360) & (g430) & (!g359) & (g389)));
	assign g433 = (((!g1) & (!g391) & (!g429) & (!g431) & (!g432)) + ((g1) & (!g391) & (!g429) & (!g431) & (!g432)) + ((g1) & (!g391) & (!g429) & (g431) & (!g432)) + ((g1) & (!g391) & (g429) & (!g431) & (!g432)) + ((g1) & (!g391) & (g429) & (g431) & (!g432)) + ((g1) & (g391) & (!g429) & (!g431) & (!g432)) + ((g1) & (g391) & (!g429) & (g431) & (!g432)));
	assign g434 = (((g1) & (!g391) & (g429) & (g432)) + ((g1) & (g391) & (!g429) & (!g432)) + ((g1) & (g391) & (!g429) & (g432)));
	assign g435 = (((!g4) & (!g2) & (!g392) & (!g426) & (!g428) & (!g433)) + ((!g4) & (!g2) & (!g392) & (!g426) & (g428) & (g433)) + ((!g4) & (!g2) & (!g392) & (g426) & (!g428) & (!g433)) + ((!g4) & (!g2) & (!g392) & (g426) & (g428) & (g433)) + ((!g4) & (!g2) & (g392) & (!g426) & (!g428) & (!g433)) + ((!g4) & (!g2) & (g392) & (!g426) & (g428) & (g433)) + ((!g4) & (!g2) & (g392) & (g426) & (g428) & (!g433)) + ((!g4) & (!g2) & (g392) & (g426) & (g428) & (g433)) + ((!g4) & (g2) & (!g392) & (!g426) & (!g428) & (!g433)) + ((!g4) & (g2) & (!g392) & (!g426) & (g428) & (g433)) + ((!g4) & (g2) & (!g392) & (g426) & (g428) & (!g433)) + ((!g4) & (g2) & (!g392) & (g426) & (g428) & (g433)) + ((!g4) & (g2) & (g392) & (!g426) & (g428) & (!g433)) + ((!g4) & (g2) & (g392) & (!g426) & (g428) & (g433)) + ((!g4) & (g2) & (g392) & (g426) & (g428) & (!g433)) + ((!g4) & (g2) & (g392) & (g426) & (g428) & (g433)) + ((g4) & (!g2) & (!g392) & (!g426) & (g428) & (!g433)) + ((g4) & (!g2) & (!g392) & (!g426) & (g428) & (g433)) + ((g4) & (!g2) & (!g392) & (g426) & (g428) & (!g433)) + ((g4) & (!g2) & (!g392) & (g426) & (g428) & (g433)) + ((g4) & (!g2) & (g392) & (!g426) & (g428) & (!g433)) + ((g4) & (!g2) & (g392) & (!g426) & (g428) & (g433)) + ((g4) & (!g2) & (g392) & (g426) & (!g428) & (!g433)) + ((g4) & (!g2) & (g392) & (g426) & (g428) & (g433)) + ((g4) & (g2) & (!g392) & (!g426) & (g428) & (!g433)) + ((g4) & (g2) & (!g392) & (!g426) & (g428) & (g433)) + ((g4) & (g2) & (!g392) & (g426) & (!g428) & (!g433)) + ((g4) & (g2) & (!g392) & (g426) & (g428) & (g433)) + ((g4) & (g2) & (g392) & (!g426) & (!g428) & (!g433)) + ((g4) & (g2) & (g392) & (!g426) & (g428) & (g433)) + ((g4) & (g2) & (g392) & (g426) & (!g428) & (!g433)) + ((g4) & (g2) & (g392) & (g426) & (g428) & (g433)));
	assign g436 = (((!g8) & (!g18) & (!g394) & (g395) & (g425) & (!g433)) + ((!g8) & (!g18) & (g394) & (!g395) & (!g425) & (!g433)) + ((!g8) & (!g18) & (g394) & (!g395) & (!g425) & (g433)) + ((!g8) & (!g18) & (g394) & (!g395) & (g425) & (!g433)) + ((!g8) & (!g18) & (g394) & (!g395) & (g425) & (g433)) + ((!g8) & (!g18) & (g394) & (g395) & (!g425) & (!g433)) + ((!g8) & (!g18) & (g394) & (g395) & (!g425) & (g433)) + ((!g8) & (!g18) & (g394) & (g395) & (g425) & (g433)) + ((!g8) & (g18) & (!g394) & (!g395) & (g425) & (!g433)) + ((!g8) & (g18) & (!g394) & (g395) & (!g425) & (!g433)) + ((!g8) & (g18) & (!g394) & (g395) & (g425) & (!g433)) + ((!g8) & (g18) & (g394) & (!g395) & (!g425) & (!g433)) + ((!g8) & (g18) & (g394) & (!g395) & (!g425) & (g433)) + ((!g8) & (g18) & (g394) & (!g395) & (g425) & (g433)) + ((!g8) & (g18) & (g394) & (g395) & (!g425) & (g433)) + ((!g8) & (g18) & (g394) & (g395) & (g425) & (g433)) + ((g8) & (!g18) & (!g394) & (!g395) & (!g425) & (!g433)) + ((g8) & (!g18) & (!g394) & (!g395) & (g425) & (!g433)) + ((g8) & (!g18) & (!g394) & (g395) & (!g425) & (!g433)) + ((g8) & (!g18) & (g394) & (!g395) & (!g425) & (g433)) + ((g8) & (!g18) & (g394) & (!g395) & (g425) & (g433)) + ((g8) & (!g18) & (g394) & (g395) & (!g425) & (g433)) + ((g8) & (!g18) & (g394) & (g395) & (g425) & (!g433)) + ((g8) & (!g18) & (g394) & (g395) & (g425) & (g433)) + ((g8) & (g18) & (!g394) & (!g395) & (!g425) & (!g433)) + ((g8) & (g18) & (g394) & (!g395) & (!g425) & (g433)) + ((g8) & (g18) & (g394) & (!g395) & (g425) & (!g433)) + ((g8) & (g18) & (g394) & (!g395) & (g425) & (g433)) + ((g8) & (g18) & (g394) & (g395) & (!g425) & (!g433)) + ((g8) & (g18) & (g394) & (g395) & (!g425) & (g433)) + ((g8) & (g18) & (g394) & (g395) & (g425) & (!g433)) + ((g8) & (g18) & (g394) & (g395) & (g425) & (g433)));
	assign g437 = (((!g18) & (!g395) & (g425) & (!g433)) + ((!g18) & (g395) & (!g425) & (!g433)) + ((!g18) & (g395) & (!g425) & (g433)) + ((!g18) & (g395) & (g425) & (g433)) + ((g18) & (!g395) & (!g425) & (!g433)) + ((g18) & (g395) & (!g425) & (g433)) + ((g18) & (g395) & (g425) & (!g433)) + ((g18) & (g395) & (g425) & (g433)));
	assign g438 = (((!g27) & (!g39) & (!g397) & (g398) & (g424) & (!g433)) + ((!g27) & (!g39) & (g397) & (!g398) & (!g424) & (!g433)) + ((!g27) & (!g39) & (g397) & (!g398) & (!g424) & (g433)) + ((!g27) & (!g39) & (g397) & (!g398) & (g424) & (!g433)) + ((!g27) & (!g39) & (g397) & (!g398) & (g424) & (g433)) + ((!g27) & (!g39) & (g397) & (g398) & (!g424) & (!g433)) + ((!g27) & (!g39) & (g397) & (g398) & (!g424) & (g433)) + ((!g27) & (!g39) & (g397) & (g398) & (g424) & (g433)) + ((!g27) & (g39) & (!g397) & (!g398) & (g424) & (!g433)) + ((!g27) & (g39) & (!g397) & (g398) & (!g424) & (!g433)) + ((!g27) & (g39) & (!g397) & (g398) & (g424) & (!g433)) + ((!g27) & (g39) & (g397) & (!g398) & (!g424) & (!g433)) + ((!g27) & (g39) & (g397) & (!g398) & (!g424) & (g433)) + ((!g27) & (g39) & (g397) & (!g398) & (g424) & (g433)) + ((!g27) & (g39) & (g397) & (g398) & (!g424) & (g433)) + ((!g27) & (g39) & (g397) & (g398) & (g424) & (g433)) + ((g27) & (!g39) & (!g397) & (!g398) & (!g424) & (!g433)) + ((g27) & (!g39) & (!g397) & (!g398) & (g424) & (!g433)) + ((g27) & (!g39) & (!g397) & (g398) & (!g424) & (!g433)) + ((g27) & (!g39) & (g397) & (!g398) & (!g424) & (g433)) + ((g27) & (!g39) & (g397) & (!g398) & (g424) & (g433)) + ((g27) & (!g39) & (g397) & (g398) & (!g424) & (g433)) + ((g27) & (!g39) & (g397) & (g398) & (g424) & (!g433)) + ((g27) & (!g39) & (g397) & (g398) & (g424) & (g433)) + ((g27) & (g39) & (!g397) & (!g398) & (!g424) & (!g433)) + ((g27) & (g39) & (g397) & (!g398) & (!g424) & (g433)) + ((g27) & (g39) & (g397) & (!g398) & (g424) & (!g433)) + ((g27) & (g39) & (g397) & (!g398) & (g424) & (g433)) + ((g27) & (g39) & (g397) & (g398) & (!g424) & (!g433)) + ((g27) & (g39) & (g397) & (g398) & (!g424) & (g433)) + ((g27) & (g39) & (g397) & (g398) & (g424) & (!g433)) + ((g27) & (g39) & (g397) & (g398) & (g424) & (g433)));
	assign g439 = (((!g39) & (!g398) & (g424) & (!g433)) + ((!g39) & (g398) & (!g424) & (!g433)) + ((!g39) & (g398) & (!g424) & (g433)) + ((!g39) & (g398) & (g424) & (g433)) + ((g39) & (!g398) & (!g424) & (!g433)) + ((g39) & (g398) & (!g424) & (g433)) + ((g39) & (g398) & (g424) & (!g433)) + ((g39) & (g398) & (g424) & (g433)));
	assign g440 = (((!g54) & (!g68) & (!g400) & (g401) & (g423) & (!g433)) + ((!g54) & (!g68) & (g400) & (!g401) & (!g423) & (!g433)) + ((!g54) & (!g68) & (g400) & (!g401) & (!g423) & (g433)) + ((!g54) & (!g68) & (g400) & (!g401) & (g423) & (!g433)) + ((!g54) & (!g68) & (g400) & (!g401) & (g423) & (g433)) + ((!g54) & (!g68) & (g400) & (g401) & (!g423) & (!g433)) + ((!g54) & (!g68) & (g400) & (g401) & (!g423) & (g433)) + ((!g54) & (!g68) & (g400) & (g401) & (g423) & (g433)) + ((!g54) & (g68) & (!g400) & (!g401) & (g423) & (!g433)) + ((!g54) & (g68) & (!g400) & (g401) & (!g423) & (!g433)) + ((!g54) & (g68) & (!g400) & (g401) & (g423) & (!g433)) + ((!g54) & (g68) & (g400) & (!g401) & (!g423) & (!g433)) + ((!g54) & (g68) & (g400) & (!g401) & (!g423) & (g433)) + ((!g54) & (g68) & (g400) & (!g401) & (g423) & (g433)) + ((!g54) & (g68) & (g400) & (g401) & (!g423) & (g433)) + ((!g54) & (g68) & (g400) & (g401) & (g423) & (g433)) + ((g54) & (!g68) & (!g400) & (!g401) & (!g423) & (!g433)) + ((g54) & (!g68) & (!g400) & (!g401) & (g423) & (!g433)) + ((g54) & (!g68) & (!g400) & (g401) & (!g423) & (!g433)) + ((g54) & (!g68) & (g400) & (!g401) & (!g423) & (g433)) + ((g54) & (!g68) & (g400) & (!g401) & (g423) & (g433)) + ((g54) & (!g68) & (g400) & (g401) & (!g423) & (g433)) + ((g54) & (!g68) & (g400) & (g401) & (g423) & (!g433)) + ((g54) & (!g68) & (g400) & (g401) & (g423) & (g433)) + ((g54) & (g68) & (!g400) & (!g401) & (!g423) & (!g433)) + ((g54) & (g68) & (g400) & (!g401) & (!g423) & (g433)) + ((g54) & (g68) & (g400) & (!g401) & (g423) & (!g433)) + ((g54) & (g68) & (g400) & (!g401) & (g423) & (g433)) + ((g54) & (g68) & (g400) & (g401) & (!g423) & (!g433)) + ((g54) & (g68) & (g400) & (g401) & (!g423) & (g433)) + ((g54) & (g68) & (g400) & (g401) & (g423) & (!g433)) + ((g54) & (g68) & (g400) & (g401) & (g423) & (g433)));
	assign g441 = (((!g68) & (!g401) & (g423) & (!g433)) + ((!g68) & (g401) & (!g423) & (!g433)) + ((!g68) & (g401) & (!g423) & (g433)) + ((!g68) & (g401) & (g423) & (g433)) + ((g68) & (!g401) & (!g423) & (!g433)) + ((g68) & (g401) & (!g423) & (g433)) + ((g68) & (g401) & (g423) & (!g433)) + ((g68) & (g401) & (g423) & (g433)));
	assign g442 = (((!g87) & (!g104) & (!g403) & (g404) & (g422) & (!g433)) + ((!g87) & (!g104) & (g403) & (!g404) & (!g422) & (!g433)) + ((!g87) & (!g104) & (g403) & (!g404) & (!g422) & (g433)) + ((!g87) & (!g104) & (g403) & (!g404) & (g422) & (!g433)) + ((!g87) & (!g104) & (g403) & (!g404) & (g422) & (g433)) + ((!g87) & (!g104) & (g403) & (g404) & (!g422) & (!g433)) + ((!g87) & (!g104) & (g403) & (g404) & (!g422) & (g433)) + ((!g87) & (!g104) & (g403) & (g404) & (g422) & (g433)) + ((!g87) & (g104) & (!g403) & (!g404) & (g422) & (!g433)) + ((!g87) & (g104) & (!g403) & (g404) & (!g422) & (!g433)) + ((!g87) & (g104) & (!g403) & (g404) & (g422) & (!g433)) + ((!g87) & (g104) & (g403) & (!g404) & (!g422) & (!g433)) + ((!g87) & (g104) & (g403) & (!g404) & (!g422) & (g433)) + ((!g87) & (g104) & (g403) & (!g404) & (g422) & (g433)) + ((!g87) & (g104) & (g403) & (g404) & (!g422) & (g433)) + ((!g87) & (g104) & (g403) & (g404) & (g422) & (g433)) + ((g87) & (!g104) & (!g403) & (!g404) & (!g422) & (!g433)) + ((g87) & (!g104) & (!g403) & (!g404) & (g422) & (!g433)) + ((g87) & (!g104) & (!g403) & (g404) & (!g422) & (!g433)) + ((g87) & (!g104) & (g403) & (!g404) & (!g422) & (g433)) + ((g87) & (!g104) & (g403) & (!g404) & (g422) & (g433)) + ((g87) & (!g104) & (g403) & (g404) & (!g422) & (g433)) + ((g87) & (!g104) & (g403) & (g404) & (g422) & (!g433)) + ((g87) & (!g104) & (g403) & (g404) & (g422) & (g433)) + ((g87) & (g104) & (!g403) & (!g404) & (!g422) & (!g433)) + ((g87) & (g104) & (g403) & (!g404) & (!g422) & (g433)) + ((g87) & (g104) & (g403) & (!g404) & (g422) & (!g433)) + ((g87) & (g104) & (g403) & (!g404) & (g422) & (g433)) + ((g87) & (g104) & (g403) & (g404) & (!g422) & (!g433)) + ((g87) & (g104) & (g403) & (g404) & (!g422) & (g433)) + ((g87) & (g104) & (g403) & (g404) & (g422) & (!g433)) + ((g87) & (g104) & (g403) & (g404) & (g422) & (g433)));
	assign g443 = (((!g104) & (!g404) & (g422) & (!g433)) + ((!g104) & (g404) & (!g422) & (!g433)) + ((!g104) & (g404) & (!g422) & (g433)) + ((!g104) & (g404) & (g422) & (g433)) + ((g104) & (!g404) & (!g422) & (!g433)) + ((g104) & (g404) & (!g422) & (g433)) + ((g104) & (g404) & (g422) & (!g433)) + ((g104) & (g404) & (g422) & (g433)));
	assign g444 = (((!g127) & (!g147) & (!g406) & (g407) & (g421) & (!g433)) + ((!g127) & (!g147) & (g406) & (!g407) & (!g421) & (!g433)) + ((!g127) & (!g147) & (g406) & (!g407) & (!g421) & (g433)) + ((!g127) & (!g147) & (g406) & (!g407) & (g421) & (!g433)) + ((!g127) & (!g147) & (g406) & (!g407) & (g421) & (g433)) + ((!g127) & (!g147) & (g406) & (g407) & (!g421) & (!g433)) + ((!g127) & (!g147) & (g406) & (g407) & (!g421) & (g433)) + ((!g127) & (!g147) & (g406) & (g407) & (g421) & (g433)) + ((!g127) & (g147) & (!g406) & (!g407) & (g421) & (!g433)) + ((!g127) & (g147) & (!g406) & (g407) & (!g421) & (!g433)) + ((!g127) & (g147) & (!g406) & (g407) & (g421) & (!g433)) + ((!g127) & (g147) & (g406) & (!g407) & (!g421) & (!g433)) + ((!g127) & (g147) & (g406) & (!g407) & (!g421) & (g433)) + ((!g127) & (g147) & (g406) & (!g407) & (g421) & (g433)) + ((!g127) & (g147) & (g406) & (g407) & (!g421) & (g433)) + ((!g127) & (g147) & (g406) & (g407) & (g421) & (g433)) + ((g127) & (!g147) & (!g406) & (!g407) & (!g421) & (!g433)) + ((g127) & (!g147) & (!g406) & (!g407) & (g421) & (!g433)) + ((g127) & (!g147) & (!g406) & (g407) & (!g421) & (!g433)) + ((g127) & (!g147) & (g406) & (!g407) & (!g421) & (g433)) + ((g127) & (!g147) & (g406) & (!g407) & (g421) & (g433)) + ((g127) & (!g147) & (g406) & (g407) & (!g421) & (g433)) + ((g127) & (!g147) & (g406) & (g407) & (g421) & (!g433)) + ((g127) & (!g147) & (g406) & (g407) & (g421) & (g433)) + ((g127) & (g147) & (!g406) & (!g407) & (!g421) & (!g433)) + ((g127) & (g147) & (g406) & (!g407) & (!g421) & (g433)) + ((g127) & (g147) & (g406) & (!g407) & (g421) & (!g433)) + ((g127) & (g147) & (g406) & (!g407) & (g421) & (g433)) + ((g127) & (g147) & (g406) & (g407) & (!g421) & (!g433)) + ((g127) & (g147) & (g406) & (g407) & (!g421) & (g433)) + ((g127) & (g147) & (g406) & (g407) & (g421) & (!g433)) + ((g127) & (g147) & (g406) & (g407) & (g421) & (g433)));
	assign g445 = (((!g147) & (!g407) & (g421) & (!g433)) + ((!g147) & (g407) & (!g421) & (!g433)) + ((!g147) & (g407) & (!g421) & (g433)) + ((!g147) & (g407) & (g421) & (g433)) + ((g147) & (!g407) & (!g421) & (!g433)) + ((g147) & (g407) & (!g421) & (g433)) + ((g147) & (g407) & (g421) & (!g433)) + ((g147) & (g407) & (g421) & (g433)));
	assign g446 = (((!g174) & (!g198) & (!g409) & (g410) & (g420) & (!g433)) + ((!g174) & (!g198) & (g409) & (!g410) & (!g420) & (!g433)) + ((!g174) & (!g198) & (g409) & (!g410) & (!g420) & (g433)) + ((!g174) & (!g198) & (g409) & (!g410) & (g420) & (!g433)) + ((!g174) & (!g198) & (g409) & (!g410) & (g420) & (g433)) + ((!g174) & (!g198) & (g409) & (g410) & (!g420) & (!g433)) + ((!g174) & (!g198) & (g409) & (g410) & (!g420) & (g433)) + ((!g174) & (!g198) & (g409) & (g410) & (g420) & (g433)) + ((!g174) & (g198) & (!g409) & (!g410) & (g420) & (!g433)) + ((!g174) & (g198) & (!g409) & (g410) & (!g420) & (!g433)) + ((!g174) & (g198) & (!g409) & (g410) & (g420) & (!g433)) + ((!g174) & (g198) & (g409) & (!g410) & (!g420) & (!g433)) + ((!g174) & (g198) & (g409) & (!g410) & (!g420) & (g433)) + ((!g174) & (g198) & (g409) & (!g410) & (g420) & (g433)) + ((!g174) & (g198) & (g409) & (g410) & (!g420) & (g433)) + ((!g174) & (g198) & (g409) & (g410) & (g420) & (g433)) + ((g174) & (!g198) & (!g409) & (!g410) & (!g420) & (!g433)) + ((g174) & (!g198) & (!g409) & (!g410) & (g420) & (!g433)) + ((g174) & (!g198) & (!g409) & (g410) & (!g420) & (!g433)) + ((g174) & (!g198) & (g409) & (!g410) & (!g420) & (g433)) + ((g174) & (!g198) & (g409) & (!g410) & (g420) & (g433)) + ((g174) & (!g198) & (g409) & (g410) & (!g420) & (g433)) + ((g174) & (!g198) & (g409) & (g410) & (g420) & (!g433)) + ((g174) & (!g198) & (g409) & (g410) & (g420) & (g433)) + ((g174) & (g198) & (!g409) & (!g410) & (!g420) & (!g433)) + ((g174) & (g198) & (g409) & (!g410) & (!g420) & (g433)) + ((g174) & (g198) & (g409) & (!g410) & (g420) & (!g433)) + ((g174) & (g198) & (g409) & (!g410) & (g420) & (g433)) + ((g174) & (g198) & (g409) & (g410) & (!g420) & (!g433)) + ((g174) & (g198) & (g409) & (g410) & (!g420) & (g433)) + ((g174) & (g198) & (g409) & (g410) & (g420) & (!g433)) + ((g174) & (g198) & (g409) & (g410) & (g420) & (g433)));
	assign g447 = (((!g198) & (!g410) & (g420) & (!g433)) + ((!g198) & (g410) & (!g420) & (!g433)) + ((!g198) & (g410) & (!g420) & (g433)) + ((!g198) & (g410) & (g420) & (g433)) + ((g198) & (!g410) & (!g420) & (!g433)) + ((g198) & (g410) & (!g420) & (g433)) + ((g198) & (g410) & (g420) & (!g433)) + ((g198) & (g410) & (g420) & (g433)));
	assign g448 = (((!g229) & (!g255) & (!g412) & (g413) & (g419) & (!g433)) + ((!g229) & (!g255) & (g412) & (!g413) & (!g419) & (!g433)) + ((!g229) & (!g255) & (g412) & (!g413) & (!g419) & (g433)) + ((!g229) & (!g255) & (g412) & (!g413) & (g419) & (!g433)) + ((!g229) & (!g255) & (g412) & (!g413) & (g419) & (g433)) + ((!g229) & (!g255) & (g412) & (g413) & (!g419) & (!g433)) + ((!g229) & (!g255) & (g412) & (g413) & (!g419) & (g433)) + ((!g229) & (!g255) & (g412) & (g413) & (g419) & (g433)) + ((!g229) & (g255) & (!g412) & (!g413) & (g419) & (!g433)) + ((!g229) & (g255) & (!g412) & (g413) & (!g419) & (!g433)) + ((!g229) & (g255) & (!g412) & (g413) & (g419) & (!g433)) + ((!g229) & (g255) & (g412) & (!g413) & (!g419) & (!g433)) + ((!g229) & (g255) & (g412) & (!g413) & (!g419) & (g433)) + ((!g229) & (g255) & (g412) & (!g413) & (g419) & (g433)) + ((!g229) & (g255) & (g412) & (g413) & (!g419) & (g433)) + ((!g229) & (g255) & (g412) & (g413) & (g419) & (g433)) + ((g229) & (!g255) & (!g412) & (!g413) & (!g419) & (!g433)) + ((g229) & (!g255) & (!g412) & (!g413) & (g419) & (!g433)) + ((g229) & (!g255) & (!g412) & (g413) & (!g419) & (!g433)) + ((g229) & (!g255) & (g412) & (!g413) & (!g419) & (g433)) + ((g229) & (!g255) & (g412) & (!g413) & (g419) & (g433)) + ((g229) & (!g255) & (g412) & (g413) & (!g419) & (g433)) + ((g229) & (!g255) & (g412) & (g413) & (g419) & (!g433)) + ((g229) & (!g255) & (g412) & (g413) & (g419) & (g433)) + ((g229) & (g255) & (!g412) & (!g413) & (!g419) & (!g433)) + ((g229) & (g255) & (g412) & (!g413) & (!g419) & (g433)) + ((g229) & (g255) & (g412) & (!g413) & (g419) & (!g433)) + ((g229) & (g255) & (g412) & (!g413) & (g419) & (g433)) + ((g229) & (g255) & (g412) & (g413) & (!g419) & (!g433)) + ((g229) & (g255) & (g412) & (g413) & (!g419) & (g433)) + ((g229) & (g255) & (g412) & (g413) & (g419) & (!g433)) + ((g229) & (g255) & (g412) & (g413) & (g419) & (g433)));
	assign g449 = (((!g255) & (!g413) & (g419) & (!g433)) + ((!g255) & (g413) & (!g419) & (!g433)) + ((!g255) & (g413) & (!g419) & (g433)) + ((!g255) & (g413) & (g419) & (g433)) + ((g255) & (!g413) & (!g419) & (!g433)) + ((g255) & (g413) & (!g419) & (g433)) + ((g255) & (g413) & (g419) & (!g433)) + ((g255) & (g413) & (g419) & (g433)));
	assign g450 = (((!g290) & (!g319) & (!g415) & (g416) & (g418) & (!g433)) + ((!g290) & (!g319) & (g415) & (!g416) & (!g418) & (!g433)) + ((!g290) & (!g319) & (g415) & (!g416) & (!g418) & (g433)) + ((!g290) & (!g319) & (g415) & (!g416) & (g418) & (!g433)) + ((!g290) & (!g319) & (g415) & (!g416) & (g418) & (g433)) + ((!g290) & (!g319) & (g415) & (g416) & (!g418) & (!g433)) + ((!g290) & (!g319) & (g415) & (g416) & (!g418) & (g433)) + ((!g290) & (!g319) & (g415) & (g416) & (g418) & (g433)) + ((!g290) & (g319) & (!g415) & (!g416) & (g418) & (!g433)) + ((!g290) & (g319) & (!g415) & (g416) & (!g418) & (!g433)) + ((!g290) & (g319) & (!g415) & (g416) & (g418) & (!g433)) + ((!g290) & (g319) & (g415) & (!g416) & (!g418) & (!g433)) + ((!g290) & (g319) & (g415) & (!g416) & (!g418) & (g433)) + ((!g290) & (g319) & (g415) & (!g416) & (g418) & (g433)) + ((!g290) & (g319) & (g415) & (g416) & (!g418) & (g433)) + ((!g290) & (g319) & (g415) & (g416) & (g418) & (g433)) + ((g290) & (!g319) & (!g415) & (!g416) & (!g418) & (!g433)) + ((g290) & (!g319) & (!g415) & (!g416) & (g418) & (!g433)) + ((g290) & (!g319) & (!g415) & (g416) & (!g418) & (!g433)) + ((g290) & (!g319) & (g415) & (!g416) & (!g418) & (g433)) + ((g290) & (!g319) & (g415) & (!g416) & (g418) & (g433)) + ((g290) & (!g319) & (g415) & (g416) & (!g418) & (g433)) + ((g290) & (!g319) & (g415) & (g416) & (g418) & (!g433)) + ((g290) & (!g319) & (g415) & (g416) & (g418) & (g433)) + ((g290) & (g319) & (!g415) & (!g416) & (!g418) & (!g433)) + ((g290) & (g319) & (g415) & (!g416) & (!g418) & (g433)) + ((g290) & (g319) & (g415) & (!g416) & (g418) & (!g433)) + ((g290) & (g319) & (g415) & (!g416) & (g418) & (g433)) + ((g290) & (g319) & (g415) & (g416) & (!g418) & (!g433)) + ((g290) & (g319) & (g415) & (g416) & (!g418) & (g433)) + ((g290) & (g319) & (g415) & (g416) & (g418) & (!g433)) + ((g290) & (g319) & (g415) & (g416) & (g418) & (g433)));
	assign g451 = (((!g319) & (!g416) & (g418) & (!g433)) + ((!g319) & (g416) & (!g418) & (!g433)) + ((!g319) & (g416) & (!g418) & (g433)) + ((!g319) & (g416) & (g418) & (g433)) + ((g319) & (!g416) & (!g418) & (!g433)) + ((g319) & (g416) & (!g418) & (g433)) + ((g319) & (g416) & (g418) & (!g433)) + ((g319) & (g416) & (g418) & (g433)));
	assign g452 = (((!g358) & (!ax86x) & (!ax87x) & (!g390) & (!g417) & (g433)) + ((!g358) & (!ax86x) & (!ax87x) & (!g390) & (g417) & (!g433)) + ((!g358) & (!ax86x) & (!ax87x) & (!g390) & (g417) & (g433)) + ((!g358) & (!ax86x) & (!ax87x) & (g390) & (!g417) & (!g433)) + ((!g358) & (!ax86x) & (ax87x) & (!g390) & (!g417) & (!g433)) + ((!g358) & (!ax86x) & (ax87x) & (g390) & (!g417) & (g433)) + ((!g358) & (!ax86x) & (ax87x) & (g390) & (g417) & (!g433)) + ((!g358) & (!ax86x) & (ax87x) & (g390) & (g417) & (g433)) + ((!g358) & (ax86x) & (!ax87x) & (g390) & (!g417) & (!g433)) + ((!g358) & (ax86x) & (!ax87x) & (g390) & (g417) & (!g433)) + ((!g358) & (ax86x) & (ax87x) & (!g390) & (!g417) & (!g433)) + ((!g358) & (ax86x) & (ax87x) & (!g390) & (!g417) & (g433)) + ((!g358) & (ax86x) & (ax87x) & (!g390) & (g417) & (!g433)) + ((!g358) & (ax86x) & (ax87x) & (!g390) & (g417) & (g433)) + ((!g358) & (ax86x) & (ax87x) & (g390) & (!g417) & (g433)) + ((!g358) & (ax86x) & (ax87x) & (g390) & (g417) & (g433)) + ((g358) & (!ax86x) & (!ax87x) & (!g390) & (!g417) & (!g433)) + ((g358) & (!ax86x) & (!ax87x) & (!g390) & (!g417) & (g433)) + ((g358) & (!ax86x) & (!ax87x) & (!g390) & (g417) & (g433)) + ((g358) & (!ax86x) & (!ax87x) & (g390) & (g417) & (!g433)) + ((g358) & (!ax86x) & (ax87x) & (!g390) & (g417) & (!g433)) + ((g358) & (!ax86x) & (ax87x) & (g390) & (!g417) & (!g433)) + ((g358) & (!ax86x) & (ax87x) & (g390) & (!g417) & (g433)) + ((g358) & (!ax86x) & (ax87x) & (g390) & (g417) & (g433)) + ((g358) & (ax86x) & (!ax87x) & (!g390) & (!g417) & (!g433)) + ((g358) & (ax86x) & (!ax87x) & (!g390) & (g417) & (!g433)) + ((g358) & (ax86x) & (ax87x) & (!g390) & (!g417) & (g433)) + ((g358) & (ax86x) & (ax87x) & (!g390) & (g417) & (g433)) + ((g358) & (ax86x) & (ax87x) & (g390) & (!g417) & (!g433)) + ((g358) & (ax86x) & (ax87x) & (g390) & (!g417) & (g433)) + ((g358) & (ax86x) & (ax87x) & (g390) & (g417) & (!g433)) + ((g358) & (ax86x) & (ax87x) & (g390) & (g417) & (g433)));
	assign g453 = (((!ax86x) & (!g390) & (!g417) & (g433)) + ((!ax86x) & (!g390) & (g417) & (!g433)) + ((!ax86x) & (!g390) & (g417) & (g433)) + ((!ax86x) & (g390) & (g417) & (!g433)) + ((ax86x) & (!g390) & (!g417) & (!g433)) + ((ax86x) & (g390) & (!g417) & (!g433)) + ((ax86x) & (g390) & (!g417) & (g433)) + ((ax86x) & (g390) & (g417) & (g433)));
	assign g454 = (((!ax82x) & (!ax83x)));
	assign g455 = (((!g390) & (!ax84x) & (!ax85x) & (!g433) & (!g454)) + ((!g390) & (!ax84x) & (ax85x) & (g433) & (!g454)) + ((!g390) & (ax84x) & (ax85x) & (g433) & (!g454)) + ((!g390) & (ax84x) & (ax85x) & (g433) & (g454)) + ((g390) & (!ax84x) & (!ax85x) & (!g433) & (!g454)) + ((g390) & (!ax84x) & (!ax85x) & (!g433) & (g454)) + ((g390) & (!ax84x) & (!ax85x) & (g433) & (!g454)) + ((g390) & (!ax84x) & (ax85x) & (!g433) & (!g454)) + ((g390) & (!ax84x) & (ax85x) & (g433) & (!g454)) + ((g390) & (!ax84x) & (ax85x) & (g433) & (g454)) + ((g390) & (ax84x) & (!ax85x) & (g433) & (!g454)) + ((g390) & (ax84x) & (!ax85x) & (g433) & (g454)) + ((g390) & (ax84x) & (ax85x) & (!g433) & (!g454)) + ((g390) & (ax84x) & (ax85x) & (!g433) & (g454)) + ((g390) & (ax84x) & (ax85x) & (g433) & (!g454)) + ((g390) & (ax84x) & (ax85x) & (g433) & (g454)));
	assign g456 = (((!g319) & (!g358) & (g452) & (g453) & (g455)) + ((!g319) & (g358) & (g452) & (!g453) & (g455)) + ((!g319) & (g358) & (g452) & (g453) & (!g455)) + ((!g319) & (g358) & (g452) & (g453) & (g455)) + ((g319) & (!g358) & (!g452) & (g453) & (g455)) + ((g319) & (!g358) & (g452) & (!g453) & (!g455)) + ((g319) & (!g358) & (g452) & (!g453) & (g455)) + ((g319) & (!g358) & (g452) & (g453) & (!g455)) + ((g319) & (!g358) & (g452) & (g453) & (g455)) + ((g319) & (g358) & (!g452) & (!g453) & (g455)) + ((g319) & (g358) & (!g452) & (g453) & (!g455)) + ((g319) & (g358) & (!g452) & (g453) & (g455)) + ((g319) & (g358) & (g452) & (!g453) & (!g455)) + ((g319) & (g358) & (g452) & (!g453) & (g455)) + ((g319) & (g358) & (g452) & (g453) & (!g455)) + ((g319) & (g358) & (g452) & (g453) & (g455)));
	assign g457 = (((!g255) & (!g290) & (g450) & (g451) & (g456)) + ((!g255) & (g290) & (g450) & (!g451) & (g456)) + ((!g255) & (g290) & (g450) & (g451) & (!g456)) + ((!g255) & (g290) & (g450) & (g451) & (g456)) + ((g255) & (!g290) & (!g450) & (g451) & (g456)) + ((g255) & (!g290) & (g450) & (!g451) & (!g456)) + ((g255) & (!g290) & (g450) & (!g451) & (g456)) + ((g255) & (!g290) & (g450) & (g451) & (!g456)) + ((g255) & (!g290) & (g450) & (g451) & (g456)) + ((g255) & (g290) & (!g450) & (!g451) & (g456)) + ((g255) & (g290) & (!g450) & (g451) & (!g456)) + ((g255) & (g290) & (!g450) & (g451) & (g456)) + ((g255) & (g290) & (g450) & (!g451) & (!g456)) + ((g255) & (g290) & (g450) & (!g451) & (g456)) + ((g255) & (g290) & (g450) & (g451) & (!g456)) + ((g255) & (g290) & (g450) & (g451) & (g456)));
	assign g458 = (((!g198) & (!g229) & (g448) & (g449) & (g457)) + ((!g198) & (g229) & (g448) & (!g449) & (g457)) + ((!g198) & (g229) & (g448) & (g449) & (!g457)) + ((!g198) & (g229) & (g448) & (g449) & (g457)) + ((g198) & (!g229) & (!g448) & (g449) & (g457)) + ((g198) & (!g229) & (g448) & (!g449) & (!g457)) + ((g198) & (!g229) & (g448) & (!g449) & (g457)) + ((g198) & (!g229) & (g448) & (g449) & (!g457)) + ((g198) & (!g229) & (g448) & (g449) & (g457)) + ((g198) & (g229) & (!g448) & (!g449) & (g457)) + ((g198) & (g229) & (!g448) & (g449) & (!g457)) + ((g198) & (g229) & (!g448) & (g449) & (g457)) + ((g198) & (g229) & (g448) & (!g449) & (!g457)) + ((g198) & (g229) & (g448) & (!g449) & (g457)) + ((g198) & (g229) & (g448) & (g449) & (!g457)) + ((g198) & (g229) & (g448) & (g449) & (g457)));
	assign g459 = (((!g147) & (!g174) & (g446) & (g447) & (g458)) + ((!g147) & (g174) & (g446) & (!g447) & (g458)) + ((!g147) & (g174) & (g446) & (g447) & (!g458)) + ((!g147) & (g174) & (g446) & (g447) & (g458)) + ((g147) & (!g174) & (!g446) & (g447) & (g458)) + ((g147) & (!g174) & (g446) & (!g447) & (!g458)) + ((g147) & (!g174) & (g446) & (!g447) & (g458)) + ((g147) & (!g174) & (g446) & (g447) & (!g458)) + ((g147) & (!g174) & (g446) & (g447) & (g458)) + ((g147) & (g174) & (!g446) & (!g447) & (g458)) + ((g147) & (g174) & (!g446) & (g447) & (!g458)) + ((g147) & (g174) & (!g446) & (g447) & (g458)) + ((g147) & (g174) & (g446) & (!g447) & (!g458)) + ((g147) & (g174) & (g446) & (!g447) & (g458)) + ((g147) & (g174) & (g446) & (g447) & (!g458)) + ((g147) & (g174) & (g446) & (g447) & (g458)));
	assign g460 = (((!g104) & (!g127) & (g444) & (g445) & (g459)) + ((!g104) & (g127) & (g444) & (!g445) & (g459)) + ((!g104) & (g127) & (g444) & (g445) & (!g459)) + ((!g104) & (g127) & (g444) & (g445) & (g459)) + ((g104) & (!g127) & (!g444) & (g445) & (g459)) + ((g104) & (!g127) & (g444) & (!g445) & (!g459)) + ((g104) & (!g127) & (g444) & (!g445) & (g459)) + ((g104) & (!g127) & (g444) & (g445) & (!g459)) + ((g104) & (!g127) & (g444) & (g445) & (g459)) + ((g104) & (g127) & (!g444) & (!g445) & (g459)) + ((g104) & (g127) & (!g444) & (g445) & (!g459)) + ((g104) & (g127) & (!g444) & (g445) & (g459)) + ((g104) & (g127) & (g444) & (!g445) & (!g459)) + ((g104) & (g127) & (g444) & (!g445) & (g459)) + ((g104) & (g127) & (g444) & (g445) & (!g459)) + ((g104) & (g127) & (g444) & (g445) & (g459)));
	assign g461 = (((!g68) & (!g87) & (g442) & (g443) & (g460)) + ((!g68) & (g87) & (g442) & (!g443) & (g460)) + ((!g68) & (g87) & (g442) & (g443) & (!g460)) + ((!g68) & (g87) & (g442) & (g443) & (g460)) + ((g68) & (!g87) & (!g442) & (g443) & (g460)) + ((g68) & (!g87) & (g442) & (!g443) & (!g460)) + ((g68) & (!g87) & (g442) & (!g443) & (g460)) + ((g68) & (!g87) & (g442) & (g443) & (!g460)) + ((g68) & (!g87) & (g442) & (g443) & (g460)) + ((g68) & (g87) & (!g442) & (!g443) & (g460)) + ((g68) & (g87) & (!g442) & (g443) & (!g460)) + ((g68) & (g87) & (!g442) & (g443) & (g460)) + ((g68) & (g87) & (g442) & (!g443) & (!g460)) + ((g68) & (g87) & (g442) & (!g443) & (g460)) + ((g68) & (g87) & (g442) & (g443) & (!g460)) + ((g68) & (g87) & (g442) & (g443) & (g460)));
	assign g462 = (((!g39) & (!g54) & (g440) & (g441) & (g461)) + ((!g39) & (g54) & (g440) & (!g441) & (g461)) + ((!g39) & (g54) & (g440) & (g441) & (!g461)) + ((!g39) & (g54) & (g440) & (g441) & (g461)) + ((g39) & (!g54) & (!g440) & (g441) & (g461)) + ((g39) & (!g54) & (g440) & (!g441) & (!g461)) + ((g39) & (!g54) & (g440) & (!g441) & (g461)) + ((g39) & (!g54) & (g440) & (g441) & (!g461)) + ((g39) & (!g54) & (g440) & (g441) & (g461)) + ((g39) & (g54) & (!g440) & (!g441) & (g461)) + ((g39) & (g54) & (!g440) & (g441) & (!g461)) + ((g39) & (g54) & (!g440) & (g441) & (g461)) + ((g39) & (g54) & (g440) & (!g441) & (!g461)) + ((g39) & (g54) & (g440) & (!g441) & (g461)) + ((g39) & (g54) & (g440) & (g441) & (!g461)) + ((g39) & (g54) & (g440) & (g441) & (g461)));
	assign g463 = (((!g18) & (!g27) & (g438) & (g439) & (g462)) + ((!g18) & (g27) & (g438) & (!g439) & (g462)) + ((!g18) & (g27) & (g438) & (g439) & (!g462)) + ((!g18) & (g27) & (g438) & (g439) & (g462)) + ((g18) & (!g27) & (!g438) & (g439) & (g462)) + ((g18) & (!g27) & (g438) & (!g439) & (!g462)) + ((g18) & (!g27) & (g438) & (!g439) & (g462)) + ((g18) & (!g27) & (g438) & (g439) & (!g462)) + ((g18) & (!g27) & (g438) & (g439) & (g462)) + ((g18) & (g27) & (!g438) & (!g439) & (g462)) + ((g18) & (g27) & (!g438) & (g439) & (!g462)) + ((g18) & (g27) & (!g438) & (g439) & (g462)) + ((g18) & (g27) & (g438) & (!g439) & (!g462)) + ((g18) & (g27) & (g438) & (!g439) & (g462)) + ((g18) & (g27) & (g438) & (g439) & (!g462)) + ((g18) & (g27) & (g438) & (g439) & (g462)));
	assign g464 = (((!g2) & (!g8) & (g436) & (g437) & (g463)) + ((!g2) & (g8) & (g436) & (!g437) & (g463)) + ((!g2) & (g8) & (g436) & (g437) & (!g463)) + ((!g2) & (g8) & (g436) & (g437) & (g463)) + ((g2) & (!g8) & (!g436) & (g437) & (g463)) + ((g2) & (!g8) & (g436) & (!g437) & (!g463)) + ((g2) & (!g8) & (g436) & (!g437) & (g463)) + ((g2) & (!g8) & (g436) & (g437) & (!g463)) + ((g2) & (!g8) & (g436) & (g437) & (g463)) + ((g2) & (g8) & (!g436) & (!g437) & (g463)) + ((g2) & (g8) & (!g436) & (g437) & (!g463)) + ((g2) & (g8) & (!g436) & (g437) & (g463)) + ((g2) & (g8) & (g436) & (!g437) & (!g463)) + ((g2) & (g8) & (g436) & (!g437) & (g463)) + ((g2) & (g8) & (g436) & (g437) & (!g463)) + ((g2) & (g8) & (g436) & (g437) & (g463)));
	assign g465 = (((!g2) & (!g392) & (g426) & (!g433)) + ((!g2) & (g392) & (!g426) & (!g433)) + ((!g2) & (g392) & (!g426) & (g433)) + ((!g2) & (g392) & (g426) & (g433)) + ((g2) & (!g392) & (!g426) & (!g433)) + ((g2) & (g392) & (!g426) & (g433)) + ((g2) & (g392) & (g426) & (!g433)) + ((g2) & (g392) & (g426) & (g433)));
	assign g466 = (((!g1) & (!g391) & (!g429) & (!g431) & (g432)) + ((!g1) & (!g391) & (!g429) & (g431) & (!g432)) + ((!g1) & (!g391) & (!g429) & (g431) & (g432)) + ((!g1) & (g391) & (g429) & (!g431) & (!g432)) + ((!g1) & (g391) & (g429) & (!g431) & (g432)) + ((!g1) & (g391) & (g429) & (g431) & (!g432)) + ((!g1) & (g391) & (g429) & (g431) & (g432)) + ((g1) & (!g391) & (!g429) & (!g431) & (g432)) + ((g1) & (!g391) & (!g429) & (g431) & (g432)) + ((g1) & (g391) & (g429) & (!g431) & (!g432)) + ((g1) & (g391) & (g429) & (!g431) & (g432)) + ((g1) & (g391) & (g429) & (g431) & (!g432)) + ((g1) & (g391) & (g429) & (g431) & (g432)));
	assign g467 = (((!g4) & (!g1) & (!g435) & (!g464) & (!g465) & (!g466)) + ((!g4) & (g1) & (!g435) & (!g464) & (!g465) & (!g466)) + ((!g4) & (g1) & (!g435) & (!g464) & (!g465) & (g466)) + ((!g4) & (g1) & (!g435) & (!g464) & (g465) & (!g466)) + ((!g4) & (g1) & (!g435) & (!g464) & (g465) & (g466)) + ((!g4) & (g1) & (!g435) & (g464) & (!g465) & (!g466)) + ((!g4) & (g1) & (!g435) & (g464) & (!g465) & (g466)) + ((!g4) & (g1) & (!g435) & (g464) & (g465) & (!g466)) + ((!g4) & (g1) & (!g435) & (g464) & (g465) & (g466)) + ((!g4) & (g1) & (g435) & (!g464) & (!g465) & (!g466)) + ((!g4) & (g1) & (g435) & (!g464) & (!g465) & (g466)) + ((g4) & (!g1) & (!g435) & (!g464) & (!g465) & (!g466)) + ((g4) & (!g1) & (!g435) & (!g464) & (g465) & (!g466)) + ((g4) & (!g1) & (!g435) & (g464) & (!g465) & (!g466)) + ((g4) & (g1) & (!g435) & (!g464) & (!g465) & (!g466)) + ((g4) & (g1) & (!g435) & (!g464) & (!g465) & (g466)) + ((g4) & (g1) & (!g435) & (!g464) & (g465) & (!g466)) + ((g4) & (g1) & (!g435) & (!g464) & (g465) & (g466)) + ((g4) & (g1) & (!g435) & (g464) & (!g465) & (!g466)) + ((g4) & (g1) & (!g435) & (g464) & (!g465) & (g466)) + ((g4) & (g1) & (!g435) & (g464) & (g465) & (!g466)) + ((g4) & (g1) & (!g435) & (g464) & (g465) & (g466)) + ((g4) & (g1) & (g435) & (!g464) & (!g465) & (!g466)) + ((g4) & (g1) & (g435) & (!g464) & (!g465) & (g466)) + ((g4) & (g1) & (g435) & (!g464) & (g465) & (!g466)) + ((g4) & (g1) & (g435) & (!g464) & (g465) & (g466)) + ((g4) & (g1) & (g435) & (g464) & (!g465) & (!g466)) + ((g4) & (g1) & (g435) & (g464) & (!g465) & (g466)));
	assign g468 = (((!g434) & (g467)));
	assign g469 = (((!g4) & (!g464) & (!g465) & (!g434) & (!g467)) + ((!g4) & (!g464) & (!g465) & (g434) & (!g467)) + ((!g4) & (!g464) & (!g465) & (g434) & (g467)) + ((!g4) & (!g464) & (g465) & (!g434) & (g467)) + ((!g4) & (g464) & (g465) & (!g434) & (!g467)) + ((!g4) & (g464) & (g465) & (!g434) & (g467)) + ((!g4) & (g464) & (g465) & (g434) & (!g467)) + ((!g4) & (g464) & (g465) & (g434) & (g467)) + ((g4) & (!g464) & (g465) & (!g434) & (!g467)) + ((g4) & (!g464) & (g465) & (!g434) & (g467)) + ((g4) & (!g464) & (g465) & (g434) & (!g467)) + ((g4) & (!g464) & (g465) & (g434) & (g467)) + ((g4) & (g464) & (!g465) & (!g434) & (!g467)) + ((g4) & (g464) & (!g465) & (g434) & (!g467)) + ((g4) & (g464) & (!g465) & (g434) & (g467)) + ((g4) & (g464) & (g465) & (!g434) & (g467)));
	assign g470 = (((!g8) & (!g437) & (g463) & (!g434) & (!g467)) + ((!g8) & (!g437) & (g463) & (g434) & (!g467)) + ((!g8) & (!g437) & (g463) & (g434) & (g467)) + ((!g8) & (g437) & (!g463) & (!g434) & (!g467)) + ((!g8) & (g437) & (!g463) & (!g434) & (g467)) + ((!g8) & (g437) & (!g463) & (g434) & (!g467)) + ((!g8) & (g437) & (!g463) & (g434) & (g467)) + ((!g8) & (g437) & (g463) & (!g434) & (g467)) + ((g8) & (!g437) & (!g463) & (!g434) & (!g467)) + ((g8) & (!g437) & (!g463) & (g434) & (!g467)) + ((g8) & (!g437) & (!g463) & (g434) & (g467)) + ((g8) & (g437) & (!g463) & (!g434) & (g467)) + ((g8) & (g437) & (g463) & (!g434) & (!g467)) + ((g8) & (g437) & (g463) & (!g434) & (g467)) + ((g8) & (g437) & (g463) & (g434) & (!g467)) + ((g8) & (g437) & (g463) & (g434) & (g467)));
	assign g471 = (((!g18) & (!g27) & (g439) & (g462)) + ((!g18) & (g27) & (!g439) & (g462)) + ((!g18) & (g27) & (g439) & (!g462)) + ((!g18) & (g27) & (g439) & (g462)) + ((g18) & (!g27) & (!g439) & (!g462)) + ((g18) & (!g27) & (!g439) & (g462)) + ((g18) & (!g27) & (g439) & (!g462)) + ((g18) & (g27) & (!g439) & (!g462)));
	assign g472 = (((!g438) & (!g434) & (!g467) & (g471)) + ((!g438) & (g434) & (!g467) & (g471)) + ((!g438) & (g434) & (g467) & (g471)) + ((g438) & (!g434) & (!g467) & (!g471)) + ((g438) & (!g434) & (g467) & (!g471)) + ((g438) & (!g434) & (g467) & (g471)) + ((g438) & (g434) & (!g467) & (!g471)) + ((g438) & (g434) & (g467) & (!g471)));
	assign g473 = (((!g27) & (!g439) & (g462) & (!g434) & (!g467)) + ((!g27) & (!g439) & (g462) & (g434) & (!g467)) + ((!g27) & (!g439) & (g462) & (g434) & (g467)) + ((!g27) & (g439) & (!g462) & (!g434) & (!g467)) + ((!g27) & (g439) & (!g462) & (!g434) & (g467)) + ((!g27) & (g439) & (!g462) & (g434) & (!g467)) + ((!g27) & (g439) & (!g462) & (g434) & (g467)) + ((!g27) & (g439) & (g462) & (!g434) & (g467)) + ((g27) & (!g439) & (!g462) & (!g434) & (!g467)) + ((g27) & (!g439) & (!g462) & (g434) & (!g467)) + ((g27) & (!g439) & (!g462) & (g434) & (g467)) + ((g27) & (g439) & (!g462) & (!g434) & (g467)) + ((g27) & (g439) & (g462) & (!g434) & (!g467)) + ((g27) & (g439) & (g462) & (!g434) & (g467)) + ((g27) & (g439) & (g462) & (g434) & (!g467)) + ((g27) & (g439) & (g462) & (g434) & (g467)));
	assign g474 = (((!g39) & (!g54) & (g441) & (g461)) + ((!g39) & (g54) & (!g441) & (g461)) + ((!g39) & (g54) & (g441) & (!g461)) + ((!g39) & (g54) & (g441) & (g461)) + ((g39) & (!g54) & (!g441) & (!g461)) + ((g39) & (!g54) & (!g441) & (g461)) + ((g39) & (!g54) & (g441) & (!g461)) + ((g39) & (g54) & (!g441) & (!g461)));
	assign g475 = (((!g440) & (!g434) & (!g467) & (g474)) + ((!g440) & (g434) & (!g467) & (g474)) + ((!g440) & (g434) & (g467) & (g474)) + ((g440) & (!g434) & (!g467) & (!g474)) + ((g440) & (!g434) & (g467) & (!g474)) + ((g440) & (!g434) & (g467) & (g474)) + ((g440) & (g434) & (!g467) & (!g474)) + ((g440) & (g434) & (g467) & (!g474)));
	assign g476 = (((!g54) & (!g441) & (g461) & (!g434) & (!g467)) + ((!g54) & (!g441) & (g461) & (g434) & (!g467)) + ((!g54) & (!g441) & (g461) & (g434) & (g467)) + ((!g54) & (g441) & (!g461) & (!g434) & (!g467)) + ((!g54) & (g441) & (!g461) & (!g434) & (g467)) + ((!g54) & (g441) & (!g461) & (g434) & (!g467)) + ((!g54) & (g441) & (!g461) & (g434) & (g467)) + ((!g54) & (g441) & (g461) & (!g434) & (g467)) + ((g54) & (!g441) & (!g461) & (!g434) & (!g467)) + ((g54) & (!g441) & (!g461) & (g434) & (!g467)) + ((g54) & (!g441) & (!g461) & (g434) & (g467)) + ((g54) & (g441) & (!g461) & (!g434) & (g467)) + ((g54) & (g441) & (g461) & (!g434) & (!g467)) + ((g54) & (g441) & (g461) & (!g434) & (g467)) + ((g54) & (g441) & (g461) & (g434) & (!g467)) + ((g54) & (g441) & (g461) & (g434) & (g467)));
	assign g477 = (((!g68) & (!g87) & (g443) & (g460)) + ((!g68) & (g87) & (!g443) & (g460)) + ((!g68) & (g87) & (g443) & (!g460)) + ((!g68) & (g87) & (g443) & (g460)) + ((g68) & (!g87) & (!g443) & (!g460)) + ((g68) & (!g87) & (!g443) & (g460)) + ((g68) & (!g87) & (g443) & (!g460)) + ((g68) & (g87) & (!g443) & (!g460)));
	assign g478 = (((!g442) & (!g434) & (!g467) & (g477)) + ((!g442) & (g434) & (!g467) & (g477)) + ((!g442) & (g434) & (g467) & (g477)) + ((g442) & (!g434) & (!g467) & (!g477)) + ((g442) & (!g434) & (g467) & (!g477)) + ((g442) & (!g434) & (g467) & (g477)) + ((g442) & (g434) & (!g467) & (!g477)) + ((g442) & (g434) & (g467) & (!g477)));
	assign g479 = (((!g87) & (!g443) & (g460) & (!g434) & (!g467)) + ((!g87) & (!g443) & (g460) & (g434) & (!g467)) + ((!g87) & (!g443) & (g460) & (g434) & (g467)) + ((!g87) & (g443) & (!g460) & (!g434) & (!g467)) + ((!g87) & (g443) & (!g460) & (!g434) & (g467)) + ((!g87) & (g443) & (!g460) & (g434) & (!g467)) + ((!g87) & (g443) & (!g460) & (g434) & (g467)) + ((!g87) & (g443) & (g460) & (!g434) & (g467)) + ((g87) & (!g443) & (!g460) & (!g434) & (!g467)) + ((g87) & (!g443) & (!g460) & (g434) & (!g467)) + ((g87) & (!g443) & (!g460) & (g434) & (g467)) + ((g87) & (g443) & (!g460) & (!g434) & (g467)) + ((g87) & (g443) & (g460) & (!g434) & (!g467)) + ((g87) & (g443) & (g460) & (!g434) & (g467)) + ((g87) & (g443) & (g460) & (g434) & (!g467)) + ((g87) & (g443) & (g460) & (g434) & (g467)));
	assign g480 = (((!g104) & (!g127) & (g445) & (g459)) + ((!g104) & (g127) & (!g445) & (g459)) + ((!g104) & (g127) & (g445) & (!g459)) + ((!g104) & (g127) & (g445) & (g459)) + ((g104) & (!g127) & (!g445) & (!g459)) + ((g104) & (!g127) & (!g445) & (g459)) + ((g104) & (!g127) & (g445) & (!g459)) + ((g104) & (g127) & (!g445) & (!g459)));
	assign g481 = (((!g444) & (!g434) & (!g467) & (g480)) + ((!g444) & (g434) & (!g467) & (g480)) + ((!g444) & (g434) & (g467) & (g480)) + ((g444) & (!g434) & (!g467) & (!g480)) + ((g444) & (!g434) & (g467) & (!g480)) + ((g444) & (!g434) & (g467) & (g480)) + ((g444) & (g434) & (!g467) & (!g480)) + ((g444) & (g434) & (g467) & (!g480)));
	assign g482 = (((!g127) & (!g445) & (g459) & (!g434) & (!g467)) + ((!g127) & (!g445) & (g459) & (g434) & (!g467)) + ((!g127) & (!g445) & (g459) & (g434) & (g467)) + ((!g127) & (g445) & (!g459) & (!g434) & (!g467)) + ((!g127) & (g445) & (!g459) & (!g434) & (g467)) + ((!g127) & (g445) & (!g459) & (g434) & (!g467)) + ((!g127) & (g445) & (!g459) & (g434) & (g467)) + ((!g127) & (g445) & (g459) & (!g434) & (g467)) + ((g127) & (!g445) & (!g459) & (!g434) & (!g467)) + ((g127) & (!g445) & (!g459) & (g434) & (!g467)) + ((g127) & (!g445) & (!g459) & (g434) & (g467)) + ((g127) & (g445) & (!g459) & (!g434) & (g467)) + ((g127) & (g445) & (g459) & (!g434) & (!g467)) + ((g127) & (g445) & (g459) & (!g434) & (g467)) + ((g127) & (g445) & (g459) & (g434) & (!g467)) + ((g127) & (g445) & (g459) & (g434) & (g467)));
	assign g483 = (((!g147) & (!g174) & (g447) & (g458)) + ((!g147) & (g174) & (!g447) & (g458)) + ((!g147) & (g174) & (g447) & (!g458)) + ((!g147) & (g174) & (g447) & (g458)) + ((g147) & (!g174) & (!g447) & (!g458)) + ((g147) & (!g174) & (!g447) & (g458)) + ((g147) & (!g174) & (g447) & (!g458)) + ((g147) & (g174) & (!g447) & (!g458)));
	assign g484 = (((!g446) & (!g434) & (!g467) & (g483)) + ((!g446) & (g434) & (!g467) & (g483)) + ((!g446) & (g434) & (g467) & (g483)) + ((g446) & (!g434) & (!g467) & (!g483)) + ((g446) & (!g434) & (g467) & (!g483)) + ((g446) & (!g434) & (g467) & (g483)) + ((g446) & (g434) & (!g467) & (!g483)) + ((g446) & (g434) & (g467) & (!g483)));
	assign g485 = (((!g174) & (!g447) & (g458) & (!g434) & (!g467)) + ((!g174) & (!g447) & (g458) & (g434) & (!g467)) + ((!g174) & (!g447) & (g458) & (g434) & (g467)) + ((!g174) & (g447) & (!g458) & (!g434) & (!g467)) + ((!g174) & (g447) & (!g458) & (!g434) & (g467)) + ((!g174) & (g447) & (!g458) & (g434) & (!g467)) + ((!g174) & (g447) & (!g458) & (g434) & (g467)) + ((!g174) & (g447) & (g458) & (!g434) & (g467)) + ((g174) & (!g447) & (!g458) & (!g434) & (!g467)) + ((g174) & (!g447) & (!g458) & (g434) & (!g467)) + ((g174) & (!g447) & (!g458) & (g434) & (g467)) + ((g174) & (g447) & (!g458) & (!g434) & (g467)) + ((g174) & (g447) & (g458) & (!g434) & (!g467)) + ((g174) & (g447) & (g458) & (!g434) & (g467)) + ((g174) & (g447) & (g458) & (g434) & (!g467)) + ((g174) & (g447) & (g458) & (g434) & (g467)));
	assign g486 = (((!g198) & (!g229) & (g449) & (g457)) + ((!g198) & (g229) & (!g449) & (g457)) + ((!g198) & (g229) & (g449) & (!g457)) + ((!g198) & (g229) & (g449) & (g457)) + ((g198) & (!g229) & (!g449) & (!g457)) + ((g198) & (!g229) & (!g449) & (g457)) + ((g198) & (!g229) & (g449) & (!g457)) + ((g198) & (g229) & (!g449) & (!g457)));
	assign g487 = (((!g448) & (!g434) & (!g467) & (g486)) + ((!g448) & (g434) & (!g467) & (g486)) + ((!g448) & (g434) & (g467) & (g486)) + ((g448) & (!g434) & (!g467) & (!g486)) + ((g448) & (!g434) & (g467) & (!g486)) + ((g448) & (!g434) & (g467) & (g486)) + ((g448) & (g434) & (!g467) & (!g486)) + ((g448) & (g434) & (g467) & (!g486)));
	assign g488 = (((!g229) & (!g449) & (g457) & (!g434) & (!g467)) + ((!g229) & (!g449) & (g457) & (g434) & (!g467)) + ((!g229) & (!g449) & (g457) & (g434) & (g467)) + ((!g229) & (g449) & (!g457) & (!g434) & (!g467)) + ((!g229) & (g449) & (!g457) & (!g434) & (g467)) + ((!g229) & (g449) & (!g457) & (g434) & (!g467)) + ((!g229) & (g449) & (!g457) & (g434) & (g467)) + ((!g229) & (g449) & (g457) & (!g434) & (g467)) + ((g229) & (!g449) & (!g457) & (!g434) & (!g467)) + ((g229) & (!g449) & (!g457) & (g434) & (!g467)) + ((g229) & (!g449) & (!g457) & (g434) & (g467)) + ((g229) & (g449) & (!g457) & (!g434) & (g467)) + ((g229) & (g449) & (g457) & (!g434) & (!g467)) + ((g229) & (g449) & (g457) & (!g434) & (g467)) + ((g229) & (g449) & (g457) & (g434) & (!g467)) + ((g229) & (g449) & (g457) & (g434) & (g467)));
	assign g489 = (((!g255) & (!g290) & (g451) & (g456)) + ((!g255) & (g290) & (!g451) & (g456)) + ((!g255) & (g290) & (g451) & (!g456)) + ((!g255) & (g290) & (g451) & (g456)) + ((g255) & (!g290) & (!g451) & (!g456)) + ((g255) & (!g290) & (!g451) & (g456)) + ((g255) & (!g290) & (g451) & (!g456)) + ((g255) & (g290) & (!g451) & (!g456)));
	assign g490 = (((!g450) & (!g434) & (!g467) & (g489)) + ((!g450) & (g434) & (!g467) & (g489)) + ((!g450) & (g434) & (g467) & (g489)) + ((g450) & (!g434) & (!g467) & (!g489)) + ((g450) & (!g434) & (g467) & (!g489)) + ((g450) & (!g434) & (g467) & (g489)) + ((g450) & (g434) & (!g467) & (!g489)) + ((g450) & (g434) & (g467) & (!g489)));
	assign g491 = (((!g290) & (!g451) & (g456) & (!g434) & (!g467)) + ((!g290) & (!g451) & (g456) & (g434) & (!g467)) + ((!g290) & (!g451) & (g456) & (g434) & (g467)) + ((!g290) & (g451) & (!g456) & (!g434) & (!g467)) + ((!g290) & (g451) & (!g456) & (!g434) & (g467)) + ((!g290) & (g451) & (!g456) & (g434) & (!g467)) + ((!g290) & (g451) & (!g456) & (g434) & (g467)) + ((!g290) & (g451) & (g456) & (!g434) & (g467)) + ((g290) & (!g451) & (!g456) & (!g434) & (!g467)) + ((g290) & (!g451) & (!g456) & (g434) & (!g467)) + ((g290) & (!g451) & (!g456) & (g434) & (g467)) + ((g290) & (g451) & (!g456) & (!g434) & (g467)) + ((g290) & (g451) & (g456) & (!g434) & (!g467)) + ((g290) & (g451) & (g456) & (!g434) & (g467)) + ((g290) & (g451) & (g456) & (g434) & (!g467)) + ((g290) & (g451) & (g456) & (g434) & (g467)));
	assign g492 = (((!g319) & (!g358) & (g453) & (g455)) + ((!g319) & (g358) & (!g453) & (g455)) + ((!g319) & (g358) & (g453) & (!g455)) + ((!g319) & (g358) & (g453) & (g455)) + ((g319) & (!g358) & (!g453) & (!g455)) + ((g319) & (!g358) & (!g453) & (g455)) + ((g319) & (!g358) & (g453) & (!g455)) + ((g319) & (g358) & (!g453) & (!g455)));
	assign g493 = (((!g452) & (!g434) & (!g467) & (g492)) + ((!g452) & (g434) & (!g467) & (g492)) + ((!g452) & (g434) & (g467) & (g492)) + ((g452) & (!g434) & (!g467) & (!g492)) + ((g452) & (!g434) & (g467) & (!g492)) + ((g452) & (!g434) & (g467) & (g492)) + ((g452) & (g434) & (!g467) & (!g492)) + ((g452) & (g434) & (g467) & (!g492)));
	assign g494 = (((!g358) & (!g453) & (g455) & (!g434) & (!g467)) + ((!g358) & (!g453) & (g455) & (g434) & (!g467)) + ((!g358) & (!g453) & (g455) & (g434) & (g467)) + ((!g358) & (g453) & (!g455) & (!g434) & (!g467)) + ((!g358) & (g453) & (!g455) & (!g434) & (g467)) + ((!g358) & (g453) & (!g455) & (g434) & (!g467)) + ((!g358) & (g453) & (!g455) & (g434) & (g467)) + ((!g358) & (g453) & (g455) & (!g434) & (g467)) + ((g358) & (!g453) & (!g455) & (!g434) & (!g467)) + ((g358) & (!g453) & (!g455) & (g434) & (!g467)) + ((g358) & (!g453) & (!g455) & (g434) & (g467)) + ((g358) & (g453) & (!g455) & (!g434) & (g467)) + ((g358) & (g453) & (g455) & (!g434) & (!g467)) + ((g358) & (g453) & (g455) & (!g434) & (g467)) + ((g358) & (g453) & (g455) & (g434) & (!g467)) + ((g358) & (g453) & (g455) & (g434) & (g467)));
	assign g495 = (((!g390) & (!ax84x) & (!g433) & (g454)) + ((!g390) & (!ax84x) & (g433) & (g454)) + ((!g390) & (ax84x) & (!g433) & (!g454)) + ((!g390) & (ax84x) & (!g433) & (g454)) + ((g390) & (!ax84x) & (!g433) & (!g454)) + ((g390) & (!ax84x) & (g433) & (!g454)) + ((g390) & (ax84x) & (g433) & (!g454)) + ((g390) & (ax84x) & (g433) & (g454)));
	assign g496 = (((!ax84x) & (!ax85x) & (!g433) & (!g434) & (!g467) & (g495)) + ((!ax84x) & (!ax85x) & (!g433) & (!g434) & (g467) & (!g495)) + ((!ax84x) & (!ax85x) & (!g433) & (!g434) & (g467) & (g495)) + ((!ax84x) & (!ax85x) & (!g433) & (g434) & (!g467) & (g495)) + ((!ax84x) & (!ax85x) & (!g433) & (g434) & (g467) & (g495)) + ((!ax84x) & (!ax85x) & (g433) & (!g434) & (!g467) & (!g495)) + ((!ax84x) & (!ax85x) & (g433) & (g434) & (!g467) & (!g495)) + ((!ax84x) & (!ax85x) & (g433) & (g434) & (g467) & (!g495)) + ((!ax84x) & (ax85x) & (!g433) & (!g434) & (!g467) & (!g495)) + ((!ax84x) & (ax85x) & (!g433) & (g434) & (!g467) & (!g495)) + ((!ax84x) & (ax85x) & (!g433) & (g434) & (g467) & (!g495)) + ((!ax84x) & (ax85x) & (g433) & (!g434) & (!g467) & (g495)) + ((!ax84x) & (ax85x) & (g433) & (!g434) & (g467) & (!g495)) + ((!ax84x) & (ax85x) & (g433) & (!g434) & (g467) & (g495)) + ((!ax84x) & (ax85x) & (g433) & (g434) & (!g467) & (g495)) + ((!ax84x) & (ax85x) & (g433) & (g434) & (g467) & (g495)) + ((ax84x) & (!ax85x) & (!g433) & (!g434) & (!g467) & (!g495)) + ((ax84x) & (!ax85x) & (!g433) & (g434) & (!g467) & (!g495)) + ((ax84x) & (!ax85x) & (!g433) & (g434) & (g467) & (!g495)) + ((ax84x) & (!ax85x) & (g433) & (!g434) & (!g467) & (!g495)) + ((ax84x) & (!ax85x) & (g433) & (g434) & (!g467) & (!g495)) + ((ax84x) & (!ax85x) & (g433) & (g434) & (g467) & (!g495)) + ((ax84x) & (ax85x) & (!g433) & (!g434) & (!g467) & (g495)) + ((ax84x) & (ax85x) & (!g433) & (!g434) & (g467) & (!g495)) + ((ax84x) & (ax85x) & (!g433) & (!g434) & (g467) & (g495)) + ((ax84x) & (ax85x) & (!g433) & (g434) & (!g467) & (g495)) + ((ax84x) & (ax85x) & (!g433) & (g434) & (g467) & (g495)) + ((ax84x) & (ax85x) & (g433) & (!g434) & (!g467) & (g495)) + ((ax84x) & (ax85x) & (g433) & (!g434) & (g467) & (!g495)) + ((ax84x) & (ax85x) & (g433) & (!g434) & (g467) & (g495)) + ((ax84x) & (ax85x) & (g433) & (g434) & (!g467) & (g495)) + ((ax84x) & (ax85x) & (g433) & (g434) & (g467) & (g495)));
	assign g497 = (((!ax84x) & (!g433) & (!g454) & (!g434) & (g467)) + ((!ax84x) & (!g433) & (g454) & (!g434) & (!g467)) + ((!ax84x) & (!g433) & (g454) & (!g434) & (g467)) + ((!ax84x) & (!g433) & (g454) & (g434) & (!g467)) + ((!ax84x) & (!g433) & (g454) & (g434) & (g467)) + ((!ax84x) & (g433) & (g454) & (!g434) & (!g467)) + ((!ax84x) & (g433) & (g454) & (g434) & (!g467)) + ((!ax84x) & (g433) & (g454) & (g434) & (g467)) + ((ax84x) & (!g433) & (!g454) & (!g434) & (!g467)) + ((ax84x) & (!g433) & (!g454) & (g434) & (!g467)) + ((ax84x) & (!g433) & (!g454) & (g434) & (g467)) + ((ax84x) & (g433) & (!g454) & (!g434) & (!g467)) + ((ax84x) & (g433) & (!g454) & (!g434) & (g467)) + ((ax84x) & (g433) & (!g454) & (g434) & (!g467)) + ((ax84x) & (g433) & (!g454) & (g434) & (g467)) + ((ax84x) & (g433) & (g454) & (!g434) & (g467)));
	assign g498 = (((!ax80x) & (!ax81x)));
	assign g499 = (((!g433) & (!ax82x) & (!ax83x) & (!g434) & (!g467) & (!g498)) + ((!g433) & (!ax82x) & (!ax83x) & (g434) & (!g467) & (!g498)) + ((!g433) & (!ax82x) & (!ax83x) & (g434) & (g467) & (!g498)) + ((!g433) & (!ax82x) & (ax83x) & (!g434) & (g467) & (!g498)) + ((!g433) & (ax82x) & (ax83x) & (!g434) & (g467) & (!g498)) + ((!g433) & (ax82x) & (ax83x) & (!g434) & (g467) & (g498)) + ((g433) & (!ax82x) & (!ax83x) & (!g434) & (!g467) & (!g498)) + ((g433) & (!ax82x) & (!ax83x) & (!g434) & (!g467) & (g498)) + ((g433) & (!ax82x) & (!ax83x) & (!g434) & (g467) & (!g498)) + ((g433) & (!ax82x) & (!ax83x) & (g434) & (!g467) & (!g498)) + ((g433) & (!ax82x) & (!ax83x) & (g434) & (!g467) & (g498)) + ((g433) & (!ax82x) & (!ax83x) & (g434) & (g467) & (!g498)) + ((g433) & (!ax82x) & (!ax83x) & (g434) & (g467) & (g498)) + ((g433) & (!ax82x) & (ax83x) & (!g434) & (!g467) & (!g498)) + ((g433) & (!ax82x) & (ax83x) & (!g434) & (g467) & (!g498)) + ((g433) & (!ax82x) & (ax83x) & (!g434) & (g467) & (g498)) + ((g433) & (!ax82x) & (ax83x) & (g434) & (!g467) & (!g498)) + ((g433) & (!ax82x) & (ax83x) & (g434) & (g467) & (!g498)) + ((g433) & (ax82x) & (!ax83x) & (!g434) & (g467) & (!g498)) + ((g433) & (ax82x) & (!ax83x) & (!g434) & (g467) & (g498)) + ((g433) & (ax82x) & (ax83x) & (!g434) & (!g467) & (!g498)) + ((g433) & (ax82x) & (ax83x) & (!g434) & (!g467) & (g498)) + ((g433) & (ax82x) & (ax83x) & (!g434) & (g467) & (!g498)) + ((g433) & (ax82x) & (ax83x) & (!g434) & (g467) & (g498)) + ((g433) & (ax82x) & (ax83x) & (g434) & (!g467) & (!g498)) + ((g433) & (ax82x) & (ax83x) & (g434) & (!g467) & (g498)) + ((g433) & (ax82x) & (ax83x) & (g434) & (g467) & (!g498)) + ((g433) & (ax82x) & (ax83x) & (g434) & (g467) & (g498)));
	assign g500 = (((!g358) & (!g390) & (g496) & (g497) & (g499)) + ((!g358) & (g390) & (g496) & (!g497) & (g499)) + ((!g358) & (g390) & (g496) & (g497) & (!g499)) + ((!g358) & (g390) & (g496) & (g497) & (g499)) + ((g358) & (!g390) & (!g496) & (g497) & (g499)) + ((g358) & (!g390) & (g496) & (!g497) & (!g499)) + ((g358) & (!g390) & (g496) & (!g497) & (g499)) + ((g358) & (!g390) & (g496) & (g497) & (!g499)) + ((g358) & (!g390) & (g496) & (g497) & (g499)) + ((g358) & (g390) & (!g496) & (!g497) & (g499)) + ((g358) & (g390) & (!g496) & (g497) & (!g499)) + ((g358) & (g390) & (!g496) & (g497) & (g499)) + ((g358) & (g390) & (g496) & (!g497) & (!g499)) + ((g358) & (g390) & (g496) & (!g497) & (g499)) + ((g358) & (g390) & (g496) & (g497) & (!g499)) + ((g358) & (g390) & (g496) & (g497) & (g499)));
	assign g501 = (((!g290) & (!g319) & (g493) & (g494) & (g500)) + ((!g290) & (g319) & (g493) & (!g494) & (g500)) + ((!g290) & (g319) & (g493) & (g494) & (!g500)) + ((!g290) & (g319) & (g493) & (g494) & (g500)) + ((g290) & (!g319) & (!g493) & (g494) & (g500)) + ((g290) & (!g319) & (g493) & (!g494) & (!g500)) + ((g290) & (!g319) & (g493) & (!g494) & (g500)) + ((g290) & (!g319) & (g493) & (g494) & (!g500)) + ((g290) & (!g319) & (g493) & (g494) & (g500)) + ((g290) & (g319) & (!g493) & (!g494) & (g500)) + ((g290) & (g319) & (!g493) & (g494) & (!g500)) + ((g290) & (g319) & (!g493) & (g494) & (g500)) + ((g290) & (g319) & (g493) & (!g494) & (!g500)) + ((g290) & (g319) & (g493) & (!g494) & (g500)) + ((g290) & (g319) & (g493) & (g494) & (!g500)) + ((g290) & (g319) & (g493) & (g494) & (g500)));
	assign g502 = (((!g229) & (!g255) & (g490) & (g491) & (g501)) + ((!g229) & (g255) & (g490) & (!g491) & (g501)) + ((!g229) & (g255) & (g490) & (g491) & (!g501)) + ((!g229) & (g255) & (g490) & (g491) & (g501)) + ((g229) & (!g255) & (!g490) & (g491) & (g501)) + ((g229) & (!g255) & (g490) & (!g491) & (!g501)) + ((g229) & (!g255) & (g490) & (!g491) & (g501)) + ((g229) & (!g255) & (g490) & (g491) & (!g501)) + ((g229) & (!g255) & (g490) & (g491) & (g501)) + ((g229) & (g255) & (!g490) & (!g491) & (g501)) + ((g229) & (g255) & (!g490) & (g491) & (!g501)) + ((g229) & (g255) & (!g490) & (g491) & (g501)) + ((g229) & (g255) & (g490) & (!g491) & (!g501)) + ((g229) & (g255) & (g490) & (!g491) & (g501)) + ((g229) & (g255) & (g490) & (g491) & (!g501)) + ((g229) & (g255) & (g490) & (g491) & (g501)));
	assign g503 = (((!g174) & (!g198) & (g487) & (g488) & (g502)) + ((!g174) & (g198) & (g487) & (!g488) & (g502)) + ((!g174) & (g198) & (g487) & (g488) & (!g502)) + ((!g174) & (g198) & (g487) & (g488) & (g502)) + ((g174) & (!g198) & (!g487) & (g488) & (g502)) + ((g174) & (!g198) & (g487) & (!g488) & (!g502)) + ((g174) & (!g198) & (g487) & (!g488) & (g502)) + ((g174) & (!g198) & (g487) & (g488) & (!g502)) + ((g174) & (!g198) & (g487) & (g488) & (g502)) + ((g174) & (g198) & (!g487) & (!g488) & (g502)) + ((g174) & (g198) & (!g487) & (g488) & (!g502)) + ((g174) & (g198) & (!g487) & (g488) & (g502)) + ((g174) & (g198) & (g487) & (!g488) & (!g502)) + ((g174) & (g198) & (g487) & (!g488) & (g502)) + ((g174) & (g198) & (g487) & (g488) & (!g502)) + ((g174) & (g198) & (g487) & (g488) & (g502)));
	assign g504 = (((!g127) & (!g147) & (g484) & (g485) & (g503)) + ((!g127) & (g147) & (g484) & (!g485) & (g503)) + ((!g127) & (g147) & (g484) & (g485) & (!g503)) + ((!g127) & (g147) & (g484) & (g485) & (g503)) + ((g127) & (!g147) & (!g484) & (g485) & (g503)) + ((g127) & (!g147) & (g484) & (!g485) & (!g503)) + ((g127) & (!g147) & (g484) & (!g485) & (g503)) + ((g127) & (!g147) & (g484) & (g485) & (!g503)) + ((g127) & (!g147) & (g484) & (g485) & (g503)) + ((g127) & (g147) & (!g484) & (!g485) & (g503)) + ((g127) & (g147) & (!g484) & (g485) & (!g503)) + ((g127) & (g147) & (!g484) & (g485) & (g503)) + ((g127) & (g147) & (g484) & (!g485) & (!g503)) + ((g127) & (g147) & (g484) & (!g485) & (g503)) + ((g127) & (g147) & (g484) & (g485) & (!g503)) + ((g127) & (g147) & (g484) & (g485) & (g503)));
	assign g505 = (((!g87) & (!g104) & (g481) & (g482) & (g504)) + ((!g87) & (g104) & (g481) & (!g482) & (g504)) + ((!g87) & (g104) & (g481) & (g482) & (!g504)) + ((!g87) & (g104) & (g481) & (g482) & (g504)) + ((g87) & (!g104) & (!g481) & (g482) & (g504)) + ((g87) & (!g104) & (g481) & (!g482) & (!g504)) + ((g87) & (!g104) & (g481) & (!g482) & (g504)) + ((g87) & (!g104) & (g481) & (g482) & (!g504)) + ((g87) & (!g104) & (g481) & (g482) & (g504)) + ((g87) & (g104) & (!g481) & (!g482) & (g504)) + ((g87) & (g104) & (!g481) & (g482) & (!g504)) + ((g87) & (g104) & (!g481) & (g482) & (g504)) + ((g87) & (g104) & (g481) & (!g482) & (!g504)) + ((g87) & (g104) & (g481) & (!g482) & (g504)) + ((g87) & (g104) & (g481) & (g482) & (!g504)) + ((g87) & (g104) & (g481) & (g482) & (g504)));
	assign g506 = (((!g54) & (!g68) & (g478) & (g479) & (g505)) + ((!g54) & (g68) & (g478) & (!g479) & (g505)) + ((!g54) & (g68) & (g478) & (g479) & (!g505)) + ((!g54) & (g68) & (g478) & (g479) & (g505)) + ((g54) & (!g68) & (!g478) & (g479) & (g505)) + ((g54) & (!g68) & (g478) & (!g479) & (!g505)) + ((g54) & (!g68) & (g478) & (!g479) & (g505)) + ((g54) & (!g68) & (g478) & (g479) & (!g505)) + ((g54) & (!g68) & (g478) & (g479) & (g505)) + ((g54) & (g68) & (!g478) & (!g479) & (g505)) + ((g54) & (g68) & (!g478) & (g479) & (!g505)) + ((g54) & (g68) & (!g478) & (g479) & (g505)) + ((g54) & (g68) & (g478) & (!g479) & (!g505)) + ((g54) & (g68) & (g478) & (!g479) & (g505)) + ((g54) & (g68) & (g478) & (g479) & (!g505)) + ((g54) & (g68) & (g478) & (g479) & (g505)));
	assign g507 = (((!g27) & (!g39) & (g475) & (g476) & (g506)) + ((!g27) & (g39) & (g475) & (!g476) & (g506)) + ((!g27) & (g39) & (g475) & (g476) & (!g506)) + ((!g27) & (g39) & (g475) & (g476) & (g506)) + ((g27) & (!g39) & (!g475) & (g476) & (g506)) + ((g27) & (!g39) & (g475) & (!g476) & (!g506)) + ((g27) & (!g39) & (g475) & (!g476) & (g506)) + ((g27) & (!g39) & (g475) & (g476) & (!g506)) + ((g27) & (!g39) & (g475) & (g476) & (g506)) + ((g27) & (g39) & (!g475) & (!g476) & (g506)) + ((g27) & (g39) & (!g475) & (g476) & (!g506)) + ((g27) & (g39) & (!g475) & (g476) & (g506)) + ((g27) & (g39) & (g475) & (!g476) & (!g506)) + ((g27) & (g39) & (g475) & (!g476) & (g506)) + ((g27) & (g39) & (g475) & (g476) & (!g506)) + ((g27) & (g39) & (g475) & (g476) & (g506)));
	assign g508 = (((!g8) & (!g18) & (g472) & (g473) & (g507)) + ((!g8) & (g18) & (g472) & (!g473) & (g507)) + ((!g8) & (g18) & (g472) & (g473) & (!g507)) + ((!g8) & (g18) & (g472) & (g473) & (g507)) + ((g8) & (!g18) & (!g472) & (g473) & (g507)) + ((g8) & (!g18) & (g472) & (!g473) & (!g507)) + ((g8) & (!g18) & (g472) & (!g473) & (g507)) + ((g8) & (!g18) & (g472) & (g473) & (!g507)) + ((g8) & (!g18) & (g472) & (g473) & (g507)) + ((g8) & (g18) & (!g472) & (!g473) & (g507)) + ((g8) & (g18) & (!g472) & (g473) & (!g507)) + ((g8) & (g18) & (!g472) & (g473) & (g507)) + ((g8) & (g18) & (g472) & (!g473) & (!g507)) + ((g8) & (g18) & (g472) & (!g473) & (g507)) + ((g8) & (g18) & (g472) & (g473) & (!g507)) + ((g8) & (g18) & (g472) & (g473) & (g507)));
	assign g509 = (((!g2) & (!g8) & (g437) & (g463)) + ((!g2) & (g8) & (!g437) & (g463)) + ((!g2) & (g8) & (g437) & (!g463)) + ((!g2) & (g8) & (g437) & (g463)) + ((g2) & (!g8) & (!g437) & (!g463)) + ((g2) & (!g8) & (!g437) & (g463)) + ((g2) & (!g8) & (g437) & (!g463)) + ((g2) & (g8) & (!g437) & (!g463)));
	assign g510 = (((!g436) & (!g434) & (!g467) & (g509)) + ((!g436) & (g434) & (!g467) & (g509)) + ((!g436) & (g434) & (g467) & (g509)) + ((g436) & (!g434) & (!g467) & (!g509)) + ((g436) & (!g434) & (g467) & (!g509)) + ((g436) & (!g434) & (g467) & (g509)) + ((g436) & (g434) & (!g467) & (!g509)) + ((g436) & (g434) & (g467) & (!g509)));
	assign g511 = (((!g4) & (!g2) & (!g470) & (!g508) & (g510)) + ((!g4) & (!g2) & (!g470) & (g508) & (g510)) + ((!g4) & (!g2) & (g470) & (!g508) & (g510)) + ((!g4) & (!g2) & (g470) & (g508) & (!g510)) + ((!g4) & (!g2) & (g470) & (g508) & (g510)) + ((!g4) & (g2) & (!g470) & (!g508) & (g510)) + ((!g4) & (g2) & (!g470) & (g508) & (!g510)) + ((!g4) & (g2) & (!g470) & (g508) & (g510)) + ((!g4) & (g2) & (g470) & (!g508) & (!g510)) + ((!g4) & (g2) & (g470) & (!g508) & (g510)) + ((!g4) & (g2) & (g470) & (g508) & (!g510)) + ((!g4) & (g2) & (g470) & (g508) & (g510)) + ((g4) & (!g2) & (g470) & (g508) & (g510)) + ((g4) & (g2) & (!g470) & (g508) & (g510)) + ((g4) & (g2) & (g470) & (!g508) & (g510)) + ((g4) & (g2) & (g470) & (g508) & (g510)));
	assign g512 = (((!g4) & (!g464) & (g465)) + ((!g4) & (g464) & (!g465)) + ((!g4) & (g464) & (g465)) + ((g4) & (g464) & (g465)));
	assign g513 = (((!g435) & (!g512) & (!g434) & (!g467)) + ((!g435) & (!g512) & (g434) & (!g467)) + ((!g435) & (!g512) & (g434) & (g467)) + ((g435) & (g512) & (!g434) & (!g467)) + ((g435) & (g512) & (!g434) & (g467)) + ((g435) & (g512) & (g434) & (!g467)) + ((g435) & (g512) & (g434) & (g467)));
	assign g514 = (((!g1) & (g435) & (!g512) & (!g434) & (g467)) + ((!g1) & (g435) & (g512) & (!g434) & (g467)) + ((g1) & (!g435) & (g512) & (g434) & (!g467)) + ((g1) & (!g435) & (g512) & (g434) & (g467)) + ((g1) & (g435) & (!g512) & (!g434) & (!g467)) + ((g1) & (g435) & (!g512) & (!g434) & (g467)) + ((g1) & (g435) & (!g512) & (g434) & (!g467)) + ((g1) & (g435) & (!g512) & (g434) & (g467)) + ((g1) & (g435) & (g512) & (!g434) & (g467)));
	assign g515 = (((!g1) & (!g469) & (!g511) & (!g513) & (!g514)) + ((g1) & (!g469) & (!g511) & (!g513) & (!g514)) + ((g1) & (!g469) & (!g511) & (g513) & (!g514)) + ((g1) & (!g469) & (g511) & (!g513) & (!g514)) + ((g1) & (!g469) & (g511) & (g513) & (!g514)) + ((g1) & (g469) & (!g511) & (!g513) & (!g514)) + ((g1) & (g469) & (!g511) & (g513) & (!g514)));
	assign g516 = (((g1) & (!g469) & (g511) & (g514)) + ((g1) & (g469) & (!g511) & (!g514)) + ((g1) & (g469) & (!g511) & (g514)));
	assign g517 = (((!g4) & (!g2) & (!g470) & (!g508) & (!g510) & (!g515)) + ((!g4) & (!g2) & (!g470) & (!g508) & (g510) & (g515)) + ((!g4) & (!g2) & (!g470) & (g508) & (!g510) & (!g515)) + ((!g4) & (!g2) & (!g470) & (g508) & (g510) & (g515)) + ((!g4) & (!g2) & (g470) & (!g508) & (!g510) & (!g515)) + ((!g4) & (!g2) & (g470) & (!g508) & (g510) & (g515)) + ((!g4) & (!g2) & (g470) & (g508) & (g510) & (!g515)) + ((!g4) & (!g2) & (g470) & (g508) & (g510) & (g515)) + ((!g4) & (g2) & (!g470) & (!g508) & (!g510) & (!g515)) + ((!g4) & (g2) & (!g470) & (!g508) & (g510) & (g515)) + ((!g4) & (g2) & (!g470) & (g508) & (g510) & (!g515)) + ((!g4) & (g2) & (!g470) & (g508) & (g510) & (g515)) + ((!g4) & (g2) & (g470) & (!g508) & (g510) & (!g515)) + ((!g4) & (g2) & (g470) & (!g508) & (g510) & (g515)) + ((!g4) & (g2) & (g470) & (g508) & (g510) & (!g515)) + ((!g4) & (g2) & (g470) & (g508) & (g510) & (g515)) + ((g4) & (!g2) & (!g470) & (!g508) & (g510) & (!g515)) + ((g4) & (!g2) & (!g470) & (!g508) & (g510) & (g515)) + ((g4) & (!g2) & (!g470) & (g508) & (g510) & (!g515)) + ((g4) & (!g2) & (!g470) & (g508) & (g510) & (g515)) + ((g4) & (!g2) & (g470) & (!g508) & (g510) & (!g515)) + ((g4) & (!g2) & (g470) & (!g508) & (g510) & (g515)) + ((g4) & (!g2) & (g470) & (g508) & (!g510) & (!g515)) + ((g4) & (!g2) & (g470) & (g508) & (g510) & (g515)) + ((g4) & (g2) & (!g470) & (!g508) & (g510) & (!g515)) + ((g4) & (g2) & (!g470) & (!g508) & (g510) & (g515)) + ((g4) & (g2) & (!g470) & (g508) & (!g510) & (!g515)) + ((g4) & (g2) & (!g470) & (g508) & (g510) & (g515)) + ((g4) & (g2) & (g470) & (!g508) & (!g510) & (!g515)) + ((g4) & (g2) & (g470) & (!g508) & (g510) & (g515)) + ((g4) & (g2) & (g470) & (g508) & (!g510) & (!g515)) + ((g4) & (g2) & (g470) & (g508) & (g510) & (g515)));
	assign g518 = (((!g8) & (!g18) & (!g472) & (g473) & (g507) & (!g515)) + ((!g8) & (!g18) & (g472) & (!g473) & (!g507) & (!g515)) + ((!g8) & (!g18) & (g472) & (!g473) & (!g507) & (g515)) + ((!g8) & (!g18) & (g472) & (!g473) & (g507) & (!g515)) + ((!g8) & (!g18) & (g472) & (!g473) & (g507) & (g515)) + ((!g8) & (!g18) & (g472) & (g473) & (!g507) & (!g515)) + ((!g8) & (!g18) & (g472) & (g473) & (!g507) & (g515)) + ((!g8) & (!g18) & (g472) & (g473) & (g507) & (g515)) + ((!g8) & (g18) & (!g472) & (!g473) & (g507) & (!g515)) + ((!g8) & (g18) & (!g472) & (g473) & (!g507) & (!g515)) + ((!g8) & (g18) & (!g472) & (g473) & (g507) & (!g515)) + ((!g8) & (g18) & (g472) & (!g473) & (!g507) & (!g515)) + ((!g8) & (g18) & (g472) & (!g473) & (!g507) & (g515)) + ((!g8) & (g18) & (g472) & (!g473) & (g507) & (g515)) + ((!g8) & (g18) & (g472) & (g473) & (!g507) & (g515)) + ((!g8) & (g18) & (g472) & (g473) & (g507) & (g515)) + ((g8) & (!g18) & (!g472) & (!g473) & (!g507) & (!g515)) + ((g8) & (!g18) & (!g472) & (!g473) & (g507) & (!g515)) + ((g8) & (!g18) & (!g472) & (g473) & (!g507) & (!g515)) + ((g8) & (!g18) & (g472) & (!g473) & (!g507) & (g515)) + ((g8) & (!g18) & (g472) & (!g473) & (g507) & (g515)) + ((g8) & (!g18) & (g472) & (g473) & (!g507) & (g515)) + ((g8) & (!g18) & (g472) & (g473) & (g507) & (!g515)) + ((g8) & (!g18) & (g472) & (g473) & (g507) & (g515)) + ((g8) & (g18) & (!g472) & (!g473) & (!g507) & (!g515)) + ((g8) & (g18) & (g472) & (!g473) & (!g507) & (g515)) + ((g8) & (g18) & (g472) & (!g473) & (g507) & (!g515)) + ((g8) & (g18) & (g472) & (!g473) & (g507) & (g515)) + ((g8) & (g18) & (g472) & (g473) & (!g507) & (!g515)) + ((g8) & (g18) & (g472) & (g473) & (!g507) & (g515)) + ((g8) & (g18) & (g472) & (g473) & (g507) & (!g515)) + ((g8) & (g18) & (g472) & (g473) & (g507) & (g515)));
	assign g519 = (((!g18) & (!g473) & (g507) & (!g515)) + ((!g18) & (g473) & (!g507) & (!g515)) + ((!g18) & (g473) & (!g507) & (g515)) + ((!g18) & (g473) & (g507) & (g515)) + ((g18) & (!g473) & (!g507) & (!g515)) + ((g18) & (g473) & (!g507) & (g515)) + ((g18) & (g473) & (g507) & (!g515)) + ((g18) & (g473) & (g507) & (g515)));
	assign g520 = (((!g27) & (!g39) & (!g475) & (g476) & (g506) & (!g515)) + ((!g27) & (!g39) & (g475) & (!g476) & (!g506) & (!g515)) + ((!g27) & (!g39) & (g475) & (!g476) & (!g506) & (g515)) + ((!g27) & (!g39) & (g475) & (!g476) & (g506) & (!g515)) + ((!g27) & (!g39) & (g475) & (!g476) & (g506) & (g515)) + ((!g27) & (!g39) & (g475) & (g476) & (!g506) & (!g515)) + ((!g27) & (!g39) & (g475) & (g476) & (!g506) & (g515)) + ((!g27) & (!g39) & (g475) & (g476) & (g506) & (g515)) + ((!g27) & (g39) & (!g475) & (!g476) & (g506) & (!g515)) + ((!g27) & (g39) & (!g475) & (g476) & (!g506) & (!g515)) + ((!g27) & (g39) & (!g475) & (g476) & (g506) & (!g515)) + ((!g27) & (g39) & (g475) & (!g476) & (!g506) & (!g515)) + ((!g27) & (g39) & (g475) & (!g476) & (!g506) & (g515)) + ((!g27) & (g39) & (g475) & (!g476) & (g506) & (g515)) + ((!g27) & (g39) & (g475) & (g476) & (!g506) & (g515)) + ((!g27) & (g39) & (g475) & (g476) & (g506) & (g515)) + ((g27) & (!g39) & (!g475) & (!g476) & (!g506) & (!g515)) + ((g27) & (!g39) & (!g475) & (!g476) & (g506) & (!g515)) + ((g27) & (!g39) & (!g475) & (g476) & (!g506) & (!g515)) + ((g27) & (!g39) & (g475) & (!g476) & (!g506) & (g515)) + ((g27) & (!g39) & (g475) & (!g476) & (g506) & (g515)) + ((g27) & (!g39) & (g475) & (g476) & (!g506) & (g515)) + ((g27) & (!g39) & (g475) & (g476) & (g506) & (!g515)) + ((g27) & (!g39) & (g475) & (g476) & (g506) & (g515)) + ((g27) & (g39) & (!g475) & (!g476) & (!g506) & (!g515)) + ((g27) & (g39) & (g475) & (!g476) & (!g506) & (g515)) + ((g27) & (g39) & (g475) & (!g476) & (g506) & (!g515)) + ((g27) & (g39) & (g475) & (!g476) & (g506) & (g515)) + ((g27) & (g39) & (g475) & (g476) & (!g506) & (!g515)) + ((g27) & (g39) & (g475) & (g476) & (!g506) & (g515)) + ((g27) & (g39) & (g475) & (g476) & (g506) & (!g515)) + ((g27) & (g39) & (g475) & (g476) & (g506) & (g515)));
	assign g521 = (((!g39) & (!g476) & (g506) & (!g515)) + ((!g39) & (g476) & (!g506) & (!g515)) + ((!g39) & (g476) & (!g506) & (g515)) + ((!g39) & (g476) & (g506) & (g515)) + ((g39) & (!g476) & (!g506) & (!g515)) + ((g39) & (g476) & (!g506) & (g515)) + ((g39) & (g476) & (g506) & (!g515)) + ((g39) & (g476) & (g506) & (g515)));
	assign g522 = (((!g54) & (!g68) & (!g478) & (g479) & (g505) & (!g515)) + ((!g54) & (!g68) & (g478) & (!g479) & (!g505) & (!g515)) + ((!g54) & (!g68) & (g478) & (!g479) & (!g505) & (g515)) + ((!g54) & (!g68) & (g478) & (!g479) & (g505) & (!g515)) + ((!g54) & (!g68) & (g478) & (!g479) & (g505) & (g515)) + ((!g54) & (!g68) & (g478) & (g479) & (!g505) & (!g515)) + ((!g54) & (!g68) & (g478) & (g479) & (!g505) & (g515)) + ((!g54) & (!g68) & (g478) & (g479) & (g505) & (g515)) + ((!g54) & (g68) & (!g478) & (!g479) & (g505) & (!g515)) + ((!g54) & (g68) & (!g478) & (g479) & (!g505) & (!g515)) + ((!g54) & (g68) & (!g478) & (g479) & (g505) & (!g515)) + ((!g54) & (g68) & (g478) & (!g479) & (!g505) & (!g515)) + ((!g54) & (g68) & (g478) & (!g479) & (!g505) & (g515)) + ((!g54) & (g68) & (g478) & (!g479) & (g505) & (g515)) + ((!g54) & (g68) & (g478) & (g479) & (!g505) & (g515)) + ((!g54) & (g68) & (g478) & (g479) & (g505) & (g515)) + ((g54) & (!g68) & (!g478) & (!g479) & (!g505) & (!g515)) + ((g54) & (!g68) & (!g478) & (!g479) & (g505) & (!g515)) + ((g54) & (!g68) & (!g478) & (g479) & (!g505) & (!g515)) + ((g54) & (!g68) & (g478) & (!g479) & (!g505) & (g515)) + ((g54) & (!g68) & (g478) & (!g479) & (g505) & (g515)) + ((g54) & (!g68) & (g478) & (g479) & (!g505) & (g515)) + ((g54) & (!g68) & (g478) & (g479) & (g505) & (!g515)) + ((g54) & (!g68) & (g478) & (g479) & (g505) & (g515)) + ((g54) & (g68) & (!g478) & (!g479) & (!g505) & (!g515)) + ((g54) & (g68) & (g478) & (!g479) & (!g505) & (g515)) + ((g54) & (g68) & (g478) & (!g479) & (g505) & (!g515)) + ((g54) & (g68) & (g478) & (!g479) & (g505) & (g515)) + ((g54) & (g68) & (g478) & (g479) & (!g505) & (!g515)) + ((g54) & (g68) & (g478) & (g479) & (!g505) & (g515)) + ((g54) & (g68) & (g478) & (g479) & (g505) & (!g515)) + ((g54) & (g68) & (g478) & (g479) & (g505) & (g515)));
	assign g523 = (((!g68) & (!g479) & (g505) & (!g515)) + ((!g68) & (g479) & (!g505) & (!g515)) + ((!g68) & (g479) & (!g505) & (g515)) + ((!g68) & (g479) & (g505) & (g515)) + ((g68) & (!g479) & (!g505) & (!g515)) + ((g68) & (g479) & (!g505) & (g515)) + ((g68) & (g479) & (g505) & (!g515)) + ((g68) & (g479) & (g505) & (g515)));
	assign g524 = (((!g87) & (!g104) & (!g481) & (g482) & (g504) & (!g515)) + ((!g87) & (!g104) & (g481) & (!g482) & (!g504) & (!g515)) + ((!g87) & (!g104) & (g481) & (!g482) & (!g504) & (g515)) + ((!g87) & (!g104) & (g481) & (!g482) & (g504) & (!g515)) + ((!g87) & (!g104) & (g481) & (!g482) & (g504) & (g515)) + ((!g87) & (!g104) & (g481) & (g482) & (!g504) & (!g515)) + ((!g87) & (!g104) & (g481) & (g482) & (!g504) & (g515)) + ((!g87) & (!g104) & (g481) & (g482) & (g504) & (g515)) + ((!g87) & (g104) & (!g481) & (!g482) & (g504) & (!g515)) + ((!g87) & (g104) & (!g481) & (g482) & (!g504) & (!g515)) + ((!g87) & (g104) & (!g481) & (g482) & (g504) & (!g515)) + ((!g87) & (g104) & (g481) & (!g482) & (!g504) & (!g515)) + ((!g87) & (g104) & (g481) & (!g482) & (!g504) & (g515)) + ((!g87) & (g104) & (g481) & (!g482) & (g504) & (g515)) + ((!g87) & (g104) & (g481) & (g482) & (!g504) & (g515)) + ((!g87) & (g104) & (g481) & (g482) & (g504) & (g515)) + ((g87) & (!g104) & (!g481) & (!g482) & (!g504) & (!g515)) + ((g87) & (!g104) & (!g481) & (!g482) & (g504) & (!g515)) + ((g87) & (!g104) & (!g481) & (g482) & (!g504) & (!g515)) + ((g87) & (!g104) & (g481) & (!g482) & (!g504) & (g515)) + ((g87) & (!g104) & (g481) & (!g482) & (g504) & (g515)) + ((g87) & (!g104) & (g481) & (g482) & (!g504) & (g515)) + ((g87) & (!g104) & (g481) & (g482) & (g504) & (!g515)) + ((g87) & (!g104) & (g481) & (g482) & (g504) & (g515)) + ((g87) & (g104) & (!g481) & (!g482) & (!g504) & (!g515)) + ((g87) & (g104) & (g481) & (!g482) & (!g504) & (g515)) + ((g87) & (g104) & (g481) & (!g482) & (g504) & (!g515)) + ((g87) & (g104) & (g481) & (!g482) & (g504) & (g515)) + ((g87) & (g104) & (g481) & (g482) & (!g504) & (!g515)) + ((g87) & (g104) & (g481) & (g482) & (!g504) & (g515)) + ((g87) & (g104) & (g481) & (g482) & (g504) & (!g515)) + ((g87) & (g104) & (g481) & (g482) & (g504) & (g515)));
	assign g525 = (((!g104) & (!g482) & (g504) & (!g515)) + ((!g104) & (g482) & (!g504) & (!g515)) + ((!g104) & (g482) & (!g504) & (g515)) + ((!g104) & (g482) & (g504) & (g515)) + ((g104) & (!g482) & (!g504) & (!g515)) + ((g104) & (g482) & (!g504) & (g515)) + ((g104) & (g482) & (g504) & (!g515)) + ((g104) & (g482) & (g504) & (g515)));
	assign g526 = (((!g127) & (!g147) & (!g484) & (g485) & (g503) & (!g515)) + ((!g127) & (!g147) & (g484) & (!g485) & (!g503) & (!g515)) + ((!g127) & (!g147) & (g484) & (!g485) & (!g503) & (g515)) + ((!g127) & (!g147) & (g484) & (!g485) & (g503) & (!g515)) + ((!g127) & (!g147) & (g484) & (!g485) & (g503) & (g515)) + ((!g127) & (!g147) & (g484) & (g485) & (!g503) & (!g515)) + ((!g127) & (!g147) & (g484) & (g485) & (!g503) & (g515)) + ((!g127) & (!g147) & (g484) & (g485) & (g503) & (g515)) + ((!g127) & (g147) & (!g484) & (!g485) & (g503) & (!g515)) + ((!g127) & (g147) & (!g484) & (g485) & (!g503) & (!g515)) + ((!g127) & (g147) & (!g484) & (g485) & (g503) & (!g515)) + ((!g127) & (g147) & (g484) & (!g485) & (!g503) & (!g515)) + ((!g127) & (g147) & (g484) & (!g485) & (!g503) & (g515)) + ((!g127) & (g147) & (g484) & (!g485) & (g503) & (g515)) + ((!g127) & (g147) & (g484) & (g485) & (!g503) & (g515)) + ((!g127) & (g147) & (g484) & (g485) & (g503) & (g515)) + ((g127) & (!g147) & (!g484) & (!g485) & (!g503) & (!g515)) + ((g127) & (!g147) & (!g484) & (!g485) & (g503) & (!g515)) + ((g127) & (!g147) & (!g484) & (g485) & (!g503) & (!g515)) + ((g127) & (!g147) & (g484) & (!g485) & (!g503) & (g515)) + ((g127) & (!g147) & (g484) & (!g485) & (g503) & (g515)) + ((g127) & (!g147) & (g484) & (g485) & (!g503) & (g515)) + ((g127) & (!g147) & (g484) & (g485) & (g503) & (!g515)) + ((g127) & (!g147) & (g484) & (g485) & (g503) & (g515)) + ((g127) & (g147) & (!g484) & (!g485) & (!g503) & (!g515)) + ((g127) & (g147) & (g484) & (!g485) & (!g503) & (g515)) + ((g127) & (g147) & (g484) & (!g485) & (g503) & (!g515)) + ((g127) & (g147) & (g484) & (!g485) & (g503) & (g515)) + ((g127) & (g147) & (g484) & (g485) & (!g503) & (!g515)) + ((g127) & (g147) & (g484) & (g485) & (!g503) & (g515)) + ((g127) & (g147) & (g484) & (g485) & (g503) & (!g515)) + ((g127) & (g147) & (g484) & (g485) & (g503) & (g515)));
	assign g527 = (((!g147) & (!g485) & (g503) & (!g515)) + ((!g147) & (g485) & (!g503) & (!g515)) + ((!g147) & (g485) & (!g503) & (g515)) + ((!g147) & (g485) & (g503) & (g515)) + ((g147) & (!g485) & (!g503) & (!g515)) + ((g147) & (g485) & (!g503) & (g515)) + ((g147) & (g485) & (g503) & (!g515)) + ((g147) & (g485) & (g503) & (g515)));
	assign g528 = (((!g174) & (!g198) & (!g487) & (g488) & (g502) & (!g515)) + ((!g174) & (!g198) & (g487) & (!g488) & (!g502) & (!g515)) + ((!g174) & (!g198) & (g487) & (!g488) & (!g502) & (g515)) + ((!g174) & (!g198) & (g487) & (!g488) & (g502) & (!g515)) + ((!g174) & (!g198) & (g487) & (!g488) & (g502) & (g515)) + ((!g174) & (!g198) & (g487) & (g488) & (!g502) & (!g515)) + ((!g174) & (!g198) & (g487) & (g488) & (!g502) & (g515)) + ((!g174) & (!g198) & (g487) & (g488) & (g502) & (g515)) + ((!g174) & (g198) & (!g487) & (!g488) & (g502) & (!g515)) + ((!g174) & (g198) & (!g487) & (g488) & (!g502) & (!g515)) + ((!g174) & (g198) & (!g487) & (g488) & (g502) & (!g515)) + ((!g174) & (g198) & (g487) & (!g488) & (!g502) & (!g515)) + ((!g174) & (g198) & (g487) & (!g488) & (!g502) & (g515)) + ((!g174) & (g198) & (g487) & (!g488) & (g502) & (g515)) + ((!g174) & (g198) & (g487) & (g488) & (!g502) & (g515)) + ((!g174) & (g198) & (g487) & (g488) & (g502) & (g515)) + ((g174) & (!g198) & (!g487) & (!g488) & (!g502) & (!g515)) + ((g174) & (!g198) & (!g487) & (!g488) & (g502) & (!g515)) + ((g174) & (!g198) & (!g487) & (g488) & (!g502) & (!g515)) + ((g174) & (!g198) & (g487) & (!g488) & (!g502) & (g515)) + ((g174) & (!g198) & (g487) & (!g488) & (g502) & (g515)) + ((g174) & (!g198) & (g487) & (g488) & (!g502) & (g515)) + ((g174) & (!g198) & (g487) & (g488) & (g502) & (!g515)) + ((g174) & (!g198) & (g487) & (g488) & (g502) & (g515)) + ((g174) & (g198) & (!g487) & (!g488) & (!g502) & (!g515)) + ((g174) & (g198) & (g487) & (!g488) & (!g502) & (g515)) + ((g174) & (g198) & (g487) & (!g488) & (g502) & (!g515)) + ((g174) & (g198) & (g487) & (!g488) & (g502) & (g515)) + ((g174) & (g198) & (g487) & (g488) & (!g502) & (!g515)) + ((g174) & (g198) & (g487) & (g488) & (!g502) & (g515)) + ((g174) & (g198) & (g487) & (g488) & (g502) & (!g515)) + ((g174) & (g198) & (g487) & (g488) & (g502) & (g515)));
	assign g529 = (((!g198) & (!g488) & (g502) & (!g515)) + ((!g198) & (g488) & (!g502) & (!g515)) + ((!g198) & (g488) & (!g502) & (g515)) + ((!g198) & (g488) & (g502) & (g515)) + ((g198) & (!g488) & (!g502) & (!g515)) + ((g198) & (g488) & (!g502) & (g515)) + ((g198) & (g488) & (g502) & (!g515)) + ((g198) & (g488) & (g502) & (g515)));
	assign g530 = (((!g229) & (!g255) & (!g490) & (g491) & (g501) & (!g515)) + ((!g229) & (!g255) & (g490) & (!g491) & (!g501) & (!g515)) + ((!g229) & (!g255) & (g490) & (!g491) & (!g501) & (g515)) + ((!g229) & (!g255) & (g490) & (!g491) & (g501) & (!g515)) + ((!g229) & (!g255) & (g490) & (!g491) & (g501) & (g515)) + ((!g229) & (!g255) & (g490) & (g491) & (!g501) & (!g515)) + ((!g229) & (!g255) & (g490) & (g491) & (!g501) & (g515)) + ((!g229) & (!g255) & (g490) & (g491) & (g501) & (g515)) + ((!g229) & (g255) & (!g490) & (!g491) & (g501) & (!g515)) + ((!g229) & (g255) & (!g490) & (g491) & (!g501) & (!g515)) + ((!g229) & (g255) & (!g490) & (g491) & (g501) & (!g515)) + ((!g229) & (g255) & (g490) & (!g491) & (!g501) & (!g515)) + ((!g229) & (g255) & (g490) & (!g491) & (!g501) & (g515)) + ((!g229) & (g255) & (g490) & (!g491) & (g501) & (g515)) + ((!g229) & (g255) & (g490) & (g491) & (!g501) & (g515)) + ((!g229) & (g255) & (g490) & (g491) & (g501) & (g515)) + ((g229) & (!g255) & (!g490) & (!g491) & (!g501) & (!g515)) + ((g229) & (!g255) & (!g490) & (!g491) & (g501) & (!g515)) + ((g229) & (!g255) & (!g490) & (g491) & (!g501) & (!g515)) + ((g229) & (!g255) & (g490) & (!g491) & (!g501) & (g515)) + ((g229) & (!g255) & (g490) & (!g491) & (g501) & (g515)) + ((g229) & (!g255) & (g490) & (g491) & (!g501) & (g515)) + ((g229) & (!g255) & (g490) & (g491) & (g501) & (!g515)) + ((g229) & (!g255) & (g490) & (g491) & (g501) & (g515)) + ((g229) & (g255) & (!g490) & (!g491) & (!g501) & (!g515)) + ((g229) & (g255) & (g490) & (!g491) & (!g501) & (g515)) + ((g229) & (g255) & (g490) & (!g491) & (g501) & (!g515)) + ((g229) & (g255) & (g490) & (!g491) & (g501) & (g515)) + ((g229) & (g255) & (g490) & (g491) & (!g501) & (!g515)) + ((g229) & (g255) & (g490) & (g491) & (!g501) & (g515)) + ((g229) & (g255) & (g490) & (g491) & (g501) & (!g515)) + ((g229) & (g255) & (g490) & (g491) & (g501) & (g515)));
	assign g531 = (((!g255) & (!g491) & (g501) & (!g515)) + ((!g255) & (g491) & (!g501) & (!g515)) + ((!g255) & (g491) & (!g501) & (g515)) + ((!g255) & (g491) & (g501) & (g515)) + ((g255) & (!g491) & (!g501) & (!g515)) + ((g255) & (g491) & (!g501) & (g515)) + ((g255) & (g491) & (g501) & (!g515)) + ((g255) & (g491) & (g501) & (g515)));
	assign g532 = (((!g290) & (!g319) & (!g493) & (g494) & (g500) & (!g515)) + ((!g290) & (!g319) & (g493) & (!g494) & (!g500) & (!g515)) + ((!g290) & (!g319) & (g493) & (!g494) & (!g500) & (g515)) + ((!g290) & (!g319) & (g493) & (!g494) & (g500) & (!g515)) + ((!g290) & (!g319) & (g493) & (!g494) & (g500) & (g515)) + ((!g290) & (!g319) & (g493) & (g494) & (!g500) & (!g515)) + ((!g290) & (!g319) & (g493) & (g494) & (!g500) & (g515)) + ((!g290) & (!g319) & (g493) & (g494) & (g500) & (g515)) + ((!g290) & (g319) & (!g493) & (!g494) & (g500) & (!g515)) + ((!g290) & (g319) & (!g493) & (g494) & (!g500) & (!g515)) + ((!g290) & (g319) & (!g493) & (g494) & (g500) & (!g515)) + ((!g290) & (g319) & (g493) & (!g494) & (!g500) & (!g515)) + ((!g290) & (g319) & (g493) & (!g494) & (!g500) & (g515)) + ((!g290) & (g319) & (g493) & (!g494) & (g500) & (g515)) + ((!g290) & (g319) & (g493) & (g494) & (!g500) & (g515)) + ((!g290) & (g319) & (g493) & (g494) & (g500) & (g515)) + ((g290) & (!g319) & (!g493) & (!g494) & (!g500) & (!g515)) + ((g290) & (!g319) & (!g493) & (!g494) & (g500) & (!g515)) + ((g290) & (!g319) & (!g493) & (g494) & (!g500) & (!g515)) + ((g290) & (!g319) & (g493) & (!g494) & (!g500) & (g515)) + ((g290) & (!g319) & (g493) & (!g494) & (g500) & (g515)) + ((g290) & (!g319) & (g493) & (g494) & (!g500) & (g515)) + ((g290) & (!g319) & (g493) & (g494) & (g500) & (!g515)) + ((g290) & (!g319) & (g493) & (g494) & (g500) & (g515)) + ((g290) & (g319) & (!g493) & (!g494) & (!g500) & (!g515)) + ((g290) & (g319) & (g493) & (!g494) & (!g500) & (g515)) + ((g290) & (g319) & (g493) & (!g494) & (g500) & (!g515)) + ((g290) & (g319) & (g493) & (!g494) & (g500) & (g515)) + ((g290) & (g319) & (g493) & (g494) & (!g500) & (!g515)) + ((g290) & (g319) & (g493) & (g494) & (!g500) & (g515)) + ((g290) & (g319) & (g493) & (g494) & (g500) & (!g515)) + ((g290) & (g319) & (g493) & (g494) & (g500) & (g515)));
	assign g533 = (((!g319) & (!g494) & (g500) & (!g515)) + ((!g319) & (g494) & (!g500) & (!g515)) + ((!g319) & (g494) & (!g500) & (g515)) + ((!g319) & (g494) & (g500) & (g515)) + ((g319) & (!g494) & (!g500) & (!g515)) + ((g319) & (g494) & (!g500) & (g515)) + ((g319) & (g494) & (g500) & (!g515)) + ((g319) & (g494) & (g500) & (g515)));
	assign g534 = (((!g358) & (!g390) & (!g496) & (g497) & (g499) & (!g515)) + ((!g358) & (!g390) & (g496) & (!g497) & (!g499) & (!g515)) + ((!g358) & (!g390) & (g496) & (!g497) & (!g499) & (g515)) + ((!g358) & (!g390) & (g496) & (!g497) & (g499) & (!g515)) + ((!g358) & (!g390) & (g496) & (!g497) & (g499) & (g515)) + ((!g358) & (!g390) & (g496) & (g497) & (!g499) & (!g515)) + ((!g358) & (!g390) & (g496) & (g497) & (!g499) & (g515)) + ((!g358) & (!g390) & (g496) & (g497) & (g499) & (g515)) + ((!g358) & (g390) & (!g496) & (!g497) & (g499) & (!g515)) + ((!g358) & (g390) & (!g496) & (g497) & (!g499) & (!g515)) + ((!g358) & (g390) & (!g496) & (g497) & (g499) & (!g515)) + ((!g358) & (g390) & (g496) & (!g497) & (!g499) & (!g515)) + ((!g358) & (g390) & (g496) & (!g497) & (!g499) & (g515)) + ((!g358) & (g390) & (g496) & (!g497) & (g499) & (g515)) + ((!g358) & (g390) & (g496) & (g497) & (!g499) & (g515)) + ((!g358) & (g390) & (g496) & (g497) & (g499) & (g515)) + ((g358) & (!g390) & (!g496) & (!g497) & (!g499) & (!g515)) + ((g358) & (!g390) & (!g496) & (!g497) & (g499) & (!g515)) + ((g358) & (!g390) & (!g496) & (g497) & (!g499) & (!g515)) + ((g358) & (!g390) & (g496) & (!g497) & (!g499) & (g515)) + ((g358) & (!g390) & (g496) & (!g497) & (g499) & (g515)) + ((g358) & (!g390) & (g496) & (g497) & (!g499) & (g515)) + ((g358) & (!g390) & (g496) & (g497) & (g499) & (!g515)) + ((g358) & (!g390) & (g496) & (g497) & (g499) & (g515)) + ((g358) & (g390) & (!g496) & (!g497) & (!g499) & (!g515)) + ((g358) & (g390) & (g496) & (!g497) & (!g499) & (g515)) + ((g358) & (g390) & (g496) & (!g497) & (g499) & (!g515)) + ((g358) & (g390) & (g496) & (!g497) & (g499) & (g515)) + ((g358) & (g390) & (g496) & (g497) & (!g499) & (!g515)) + ((g358) & (g390) & (g496) & (g497) & (!g499) & (g515)) + ((g358) & (g390) & (g496) & (g497) & (g499) & (!g515)) + ((g358) & (g390) & (g496) & (g497) & (g499) & (g515)));
	assign g535 = (((!g390) & (!g497) & (g499) & (!g515)) + ((!g390) & (g497) & (!g499) & (!g515)) + ((!g390) & (g497) & (!g499) & (g515)) + ((!g390) & (g497) & (g499) & (g515)) + ((g390) & (!g497) & (!g499) & (!g515)) + ((g390) & (g497) & (!g499) & (g515)) + ((g390) & (g497) & (g499) & (!g515)) + ((g390) & (g497) & (g499) & (g515)));
	assign g536 = (((!g433) & (!ax82x) & (!ax83x) & (!g468) & (!g498) & (g515)) + ((!g433) & (!ax82x) & (!ax83x) & (!g468) & (g498) & (!g515)) + ((!g433) & (!ax82x) & (!ax83x) & (!g468) & (g498) & (g515)) + ((!g433) & (!ax82x) & (!ax83x) & (g468) & (!g498) & (!g515)) + ((!g433) & (!ax82x) & (ax83x) & (!g468) & (!g498) & (!g515)) + ((!g433) & (!ax82x) & (ax83x) & (g468) & (!g498) & (g515)) + ((!g433) & (!ax82x) & (ax83x) & (g468) & (g498) & (!g515)) + ((!g433) & (!ax82x) & (ax83x) & (g468) & (g498) & (g515)) + ((!g433) & (ax82x) & (!ax83x) & (g468) & (!g498) & (!g515)) + ((!g433) & (ax82x) & (!ax83x) & (g468) & (g498) & (!g515)) + ((!g433) & (ax82x) & (ax83x) & (!g468) & (!g498) & (!g515)) + ((!g433) & (ax82x) & (ax83x) & (!g468) & (!g498) & (g515)) + ((!g433) & (ax82x) & (ax83x) & (!g468) & (g498) & (!g515)) + ((!g433) & (ax82x) & (ax83x) & (!g468) & (g498) & (g515)) + ((!g433) & (ax82x) & (ax83x) & (g468) & (!g498) & (g515)) + ((!g433) & (ax82x) & (ax83x) & (g468) & (g498) & (g515)) + ((g433) & (!ax82x) & (!ax83x) & (!g468) & (!g498) & (!g515)) + ((g433) & (!ax82x) & (!ax83x) & (!g468) & (!g498) & (g515)) + ((g433) & (!ax82x) & (!ax83x) & (!g468) & (g498) & (g515)) + ((g433) & (!ax82x) & (!ax83x) & (g468) & (g498) & (!g515)) + ((g433) & (!ax82x) & (ax83x) & (!g468) & (g498) & (!g515)) + ((g433) & (!ax82x) & (ax83x) & (g468) & (!g498) & (!g515)) + ((g433) & (!ax82x) & (ax83x) & (g468) & (!g498) & (g515)) + ((g433) & (!ax82x) & (ax83x) & (g468) & (g498) & (g515)) + ((g433) & (ax82x) & (!ax83x) & (!g468) & (!g498) & (!g515)) + ((g433) & (ax82x) & (!ax83x) & (!g468) & (g498) & (!g515)) + ((g433) & (ax82x) & (ax83x) & (!g468) & (!g498) & (g515)) + ((g433) & (ax82x) & (ax83x) & (!g468) & (g498) & (g515)) + ((g433) & (ax82x) & (ax83x) & (g468) & (!g498) & (!g515)) + ((g433) & (ax82x) & (ax83x) & (g468) & (!g498) & (g515)) + ((g433) & (ax82x) & (ax83x) & (g468) & (g498) & (!g515)) + ((g433) & (ax82x) & (ax83x) & (g468) & (g498) & (g515)));
	assign g537 = (((!ax82x) & (!g468) & (!g498) & (g515)) + ((!ax82x) & (!g468) & (g498) & (!g515)) + ((!ax82x) & (!g468) & (g498) & (g515)) + ((!ax82x) & (g468) & (g498) & (!g515)) + ((ax82x) & (!g468) & (!g498) & (!g515)) + ((ax82x) & (g468) & (!g498) & (!g515)) + ((ax82x) & (g468) & (!g498) & (g515)) + ((ax82x) & (g468) & (g498) & (g515)));
	assign g538 = (((!ax78x) & (!ax79x)));
	assign g539 = (((!g468) & (!ax80x) & (!ax81x) & (!g515) & (!g538)) + ((!g468) & (!ax80x) & (ax81x) & (g515) & (!g538)) + ((!g468) & (ax80x) & (ax81x) & (g515) & (!g538)) + ((!g468) & (ax80x) & (ax81x) & (g515) & (g538)) + ((g468) & (!ax80x) & (!ax81x) & (!g515) & (!g538)) + ((g468) & (!ax80x) & (!ax81x) & (!g515) & (g538)) + ((g468) & (!ax80x) & (!ax81x) & (g515) & (!g538)) + ((g468) & (!ax80x) & (ax81x) & (!g515) & (!g538)) + ((g468) & (!ax80x) & (ax81x) & (g515) & (!g538)) + ((g468) & (!ax80x) & (ax81x) & (g515) & (g538)) + ((g468) & (ax80x) & (!ax81x) & (g515) & (!g538)) + ((g468) & (ax80x) & (!ax81x) & (g515) & (g538)) + ((g468) & (ax80x) & (ax81x) & (!g515) & (!g538)) + ((g468) & (ax80x) & (ax81x) & (!g515) & (g538)) + ((g468) & (ax80x) & (ax81x) & (g515) & (!g538)) + ((g468) & (ax80x) & (ax81x) & (g515) & (g538)));
	assign g540 = (((!g390) & (!g433) & (g536) & (g537) & (g539)) + ((!g390) & (g433) & (g536) & (!g537) & (g539)) + ((!g390) & (g433) & (g536) & (g537) & (!g539)) + ((!g390) & (g433) & (g536) & (g537) & (g539)) + ((g390) & (!g433) & (!g536) & (g537) & (g539)) + ((g390) & (!g433) & (g536) & (!g537) & (!g539)) + ((g390) & (!g433) & (g536) & (!g537) & (g539)) + ((g390) & (!g433) & (g536) & (g537) & (!g539)) + ((g390) & (!g433) & (g536) & (g537) & (g539)) + ((g390) & (g433) & (!g536) & (!g537) & (g539)) + ((g390) & (g433) & (!g536) & (g537) & (!g539)) + ((g390) & (g433) & (!g536) & (g537) & (g539)) + ((g390) & (g433) & (g536) & (!g537) & (!g539)) + ((g390) & (g433) & (g536) & (!g537) & (g539)) + ((g390) & (g433) & (g536) & (g537) & (!g539)) + ((g390) & (g433) & (g536) & (g537) & (g539)));
	assign g541 = (((!g319) & (!g358) & (g534) & (g535) & (g540)) + ((!g319) & (g358) & (g534) & (!g535) & (g540)) + ((!g319) & (g358) & (g534) & (g535) & (!g540)) + ((!g319) & (g358) & (g534) & (g535) & (g540)) + ((g319) & (!g358) & (!g534) & (g535) & (g540)) + ((g319) & (!g358) & (g534) & (!g535) & (!g540)) + ((g319) & (!g358) & (g534) & (!g535) & (g540)) + ((g319) & (!g358) & (g534) & (g535) & (!g540)) + ((g319) & (!g358) & (g534) & (g535) & (g540)) + ((g319) & (g358) & (!g534) & (!g535) & (g540)) + ((g319) & (g358) & (!g534) & (g535) & (!g540)) + ((g319) & (g358) & (!g534) & (g535) & (g540)) + ((g319) & (g358) & (g534) & (!g535) & (!g540)) + ((g319) & (g358) & (g534) & (!g535) & (g540)) + ((g319) & (g358) & (g534) & (g535) & (!g540)) + ((g319) & (g358) & (g534) & (g535) & (g540)));
	assign g542 = (((!g255) & (!g290) & (g532) & (g533) & (g541)) + ((!g255) & (g290) & (g532) & (!g533) & (g541)) + ((!g255) & (g290) & (g532) & (g533) & (!g541)) + ((!g255) & (g290) & (g532) & (g533) & (g541)) + ((g255) & (!g290) & (!g532) & (g533) & (g541)) + ((g255) & (!g290) & (g532) & (!g533) & (!g541)) + ((g255) & (!g290) & (g532) & (!g533) & (g541)) + ((g255) & (!g290) & (g532) & (g533) & (!g541)) + ((g255) & (!g290) & (g532) & (g533) & (g541)) + ((g255) & (g290) & (!g532) & (!g533) & (g541)) + ((g255) & (g290) & (!g532) & (g533) & (!g541)) + ((g255) & (g290) & (!g532) & (g533) & (g541)) + ((g255) & (g290) & (g532) & (!g533) & (!g541)) + ((g255) & (g290) & (g532) & (!g533) & (g541)) + ((g255) & (g290) & (g532) & (g533) & (!g541)) + ((g255) & (g290) & (g532) & (g533) & (g541)));
	assign g543 = (((!g198) & (!g229) & (g530) & (g531) & (g542)) + ((!g198) & (g229) & (g530) & (!g531) & (g542)) + ((!g198) & (g229) & (g530) & (g531) & (!g542)) + ((!g198) & (g229) & (g530) & (g531) & (g542)) + ((g198) & (!g229) & (!g530) & (g531) & (g542)) + ((g198) & (!g229) & (g530) & (!g531) & (!g542)) + ((g198) & (!g229) & (g530) & (!g531) & (g542)) + ((g198) & (!g229) & (g530) & (g531) & (!g542)) + ((g198) & (!g229) & (g530) & (g531) & (g542)) + ((g198) & (g229) & (!g530) & (!g531) & (g542)) + ((g198) & (g229) & (!g530) & (g531) & (!g542)) + ((g198) & (g229) & (!g530) & (g531) & (g542)) + ((g198) & (g229) & (g530) & (!g531) & (!g542)) + ((g198) & (g229) & (g530) & (!g531) & (g542)) + ((g198) & (g229) & (g530) & (g531) & (!g542)) + ((g198) & (g229) & (g530) & (g531) & (g542)));
	assign g544 = (((!g147) & (!g174) & (g528) & (g529) & (g543)) + ((!g147) & (g174) & (g528) & (!g529) & (g543)) + ((!g147) & (g174) & (g528) & (g529) & (!g543)) + ((!g147) & (g174) & (g528) & (g529) & (g543)) + ((g147) & (!g174) & (!g528) & (g529) & (g543)) + ((g147) & (!g174) & (g528) & (!g529) & (!g543)) + ((g147) & (!g174) & (g528) & (!g529) & (g543)) + ((g147) & (!g174) & (g528) & (g529) & (!g543)) + ((g147) & (!g174) & (g528) & (g529) & (g543)) + ((g147) & (g174) & (!g528) & (!g529) & (g543)) + ((g147) & (g174) & (!g528) & (g529) & (!g543)) + ((g147) & (g174) & (!g528) & (g529) & (g543)) + ((g147) & (g174) & (g528) & (!g529) & (!g543)) + ((g147) & (g174) & (g528) & (!g529) & (g543)) + ((g147) & (g174) & (g528) & (g529) & (!g543)) + ((g147) & (g174) & (g528) & (g529) & (g543)));
	assign g545 = (((!g104) & (!g127) & (g526) & (g527) & (g544)) + ((!g104) & (g127) & (g526) & (!g527) & (g544)) + ((!g104) & (g127) & (g526) & (g527) & (!g544)) + ((!g104) & (g127) & (g526) & (g527) & (g544)) + ((g104) & (!g127) & (!g526) & (g527) & (g544)) + ((g104) & (!g127) & (g526) & (!g527) & (!g544)) + ((g104) & (!g127) & (g526) & (!g527) & (g544)) + ((g104) & (!g127) & (g526) & (g527) & (!g544)) + ((g104) & (!g127) & (g526) & (g527) & (g544)) + ((g104) & (g127) & (!g526) & (!g527) & (g544)) + ((g104) & (g127) & (!g526) & (g527) & (!g544)) + ((g104) & (g127) & (!g526) & (g527) & (g544)) + ((g104) & (g127) & (g526) & (!g527) & (!g544)) + ((g104) & (g127) & (g526) & (!g527) & (g544)) + ((g104) & (g127) & (g526) & (g527) & (!g544)) + ((g104) & (g127) & (g526) & (g527) & (g544)));
	assign g546 = (((!g68) & (!g87) & (g524) & (g525) & (g545)) + ((!g68) & (g87) & (g524) & (!g525) & (g545)) + ((!g68) & (g87) & (g524) & (g525) & (!g545)) + ((!g68) & (g87) & (g524) & (g525) & (g545)) + ((g68) & (!g87) & (!g524) & (g525) & (g545)) + ((g68) & (!g87) & (g524) & (!g525) & (!g545)) + ((g68) & (!g87) & (g524) & (!g525) & (g545)) + ((g68) & (!g87) & (g524) & (g525) & (!g545)) + ((g68) & (!g87) & (g524) & (g525) & (g545)) + ((g68) & (g87) & (!g524) & (!g525) & (g545)) + ((g68) & (g87) & (!g524) & (g525) & (!g545)) + ((g68) & (g87) & (!g524) & (g525) & (g545)) + ((g68) & (g87) & (g524) & (!g525) & (!g545)) + ((g68) & (g87) & (g524) & (!g525) & (g545)) + ((g68) & (g87) & (g524) & (g525) & (!g545)) + ((g68) & (g87) & (g524) & (g525) & (g545)));
	assign g547 = (((!g39) & (!g54) & (g522) & (g523) & (g546)) + ((!g39) & (g54) & (g522) & (!g523) & (g546)) + ((!g39) & (g54) & (g522) & (g523) & (!g546)) + ((!g39) & (g54) & (g522) & (g523) & (g546)) + ((g39) & (!g54) & (!g522) & (g523) & (g546)) + ((g39) & (!g54) & (g522) & (!g523) & (!g546)) + ((g39) & (!g54) & (g522) & (!g523) & (g546)) + ((g39) & (!g54) & (g522) & (g523) & (!g546)) + ((g39) & (!g54) & (g522) & (g523) & (g546)) + ((g39) & (g54) & (!g522) & (!g523) & (g546)) + ((g39) & (g54) & (!g522) & (g523) & (!g546)) + ((g39) & (g54) & (!g522) & (g523) & (g546)) + ((g39) & (g54) & (g522) & (!g523) & (!g546)) + ((g39) & (g54) & (g522) & (!g523) & (g546)) + ((g39) & (g54) & (g522) & (g523) & (!g546)) + ((g39) & (g54) & (g522) & (g523) & (g546)));
	assign g548 = (((!g18) & (!g27) & (g520) & (g521) & (g547)) + ((!g18) & (g27) & (g520) & (!g521) & (g547)) + ((!g18) & (g27) & (g520) & (g521) & (!g547)) + ((!g18) & (g27) & (g520) & (g521) & (g547)) + ((g18) & (!g27) & (!g520) & (g521) & (g547)) + ((g18) & (!g27) & (g520) & (!g521) & (!g547)) + ((g18) & (!g27) & (g520) & (!g521) & (g547)) + ((g18) & (!g27) & (g520) & (g521) & (!g547)) + ((g18) & (!g27) & (g520) & (g521) & (g547)) + ((g18) & (g27) & (!g520) & (!g521) & (g547)) + ((g18) & (g27) & (!g520) & (g521) & (!g547)) + ((g18) & (g27) & (!g520) & (g521) & (g547)) + ((g18) & (g27) & (g520) & (!g521) & (!g547)) + ((g18) & (g27) & (g520) & (!g521) & (g547)) + ((g18) & (g27) & (g520) & (g521) & (!g547)) + ((g18) & (g27) & (g520) & (g521) & (g547)));
	assign g549 = (((!g2) & (!g8) & (g518) & (g519) & (g548)) + ((!g2) & (g8) & (g518) & (!g519) & (g548)) + ((!g2) & (g8) & (g518) & (g519) & (!g548)) + ((!g2) & (g8) & (g518) & (g519) & (g548)) + ((g2) & (!g8) & (!g518) & (g519) & (g548)) + ((g2) & (!g8) & (g518) & (!g519) & (!g548)) + ((g2) & (!g8) & (g518) & (!g519) & (g548)) + ((g2) & (!g8) & (g518) & (g519) & (!g548)) + ((g2) & (!g8) & (g518) & (g519) & (g548)) + ((g2) & (g8) & (!g518) & (!g519) & (g548)) + ((g2) & (g8) & (!g518) & (g519) & (!g548)) + ((g2) & (g8) & (!g518) & (g519) & (g548)) + ((g2) & (g8) & (g518) & (!g519) & (!g548)) + ((g2) & (g8) & (g518) & (!g519) & (g548)) + ((g2) & (g8) & (g518) & (g519) & (!g548)) + ((g2) & (g8) & (g518) & (g519) & (g548)));
	assign g550 = (((!g2) & (!g470) & (g508) & (!g515)) + ((!g2) & (g470) & (!g508) & (!g515)) + ((!g2) & (g470) & (!g508) & (g515)) + ((!g2) & (g470) & (g508) & (g515)) + ((g2) & (!g470) & (!g508) & (!g515)) + ((g2) & (g470) & (!g508) & (g515)) + ((g2) & (g470) & (g508) & (!g515)) + ((g2) & (g470) & (g508) & (g515)));
	assign g551 = (((!g1) & (!g469) & (!g511) & (!g513) & (g514)) + ((!g1) & (!g469) & (!g511) & (g513) & (!g514)) + ((!g1) & (!g469) & (!g511) & (g513) & (g514)) + ((!g1) & (g469) & (g511) & (!g513) & (!g514)) + ((!g1) & (g469) & (g511) & (!g513) & (g514)) + ((!g1) & (g469) & (g511) & (g513) & (!g514)) + ((!g1) & (g469) & (g511) & (g513) & (g514)) + ((g1) & (!g469) & (!g511) & (!g513) & (g514)) + ((g1) & (!g469) & (!g511) & (g513) & (g514)) + ((g1) & (g469) & (g511) & (!g513) & (!g514)) + ((g1) & (g469) & (g511) & (!g513) & (g514)) + ((g1) & (g469) & (g511) & (g513) & (!g514)) + ((g1) & (g469) & (g511) & (g513) & (g514)));
	assign g552 = (((!g4) & (!g1) & (!g517) & (!g549) & (!g550) & (!g551)) + ((!g4) & (g1) & (!g517) & (!g549) & (!g550) & (!g551)) + ((!g4) & (g1) & (!g517) & (!g549) & (!g550) & (g551)) + ((!g4) & (g1) & (!g517) & (!g549) & (g550) & (!g551)) + ((!g4) & (g1) & (!g517) & (!g549) & (g550) & (g551)) + ((!g4) & (g1) & (!g517) & (g549) & (!g550) & (!g551)) + ((!g4) & (g1) & (!g517) & (g549) & (!g550) & (g551)) + ((!g4) & (g1) & (!g517) & (g549) & (g550) & (!g551)) + ((!g4) & (g1) & (!g517) & (g549) & (g550) & (g551)) + ((!g4) & (g1) & (g517) & (!g549) & (!g550) & (!g551)) + ((!g4) & (g1) & (g517) & (!g549) & (!g550) & (g551)) + ((g4) & (!g1) & (!g517) & (!g549) & (!g550) & (!g551)) + ((g4) & (!g1) & (!g517) & (!g549) & (g550) & (!g551)) + ((g4) & (!g1) & (!g517) & (g549) & (!g550) & (!g551)) + ((g4) & (g1) & (!g517) & (!g549) & (!g550) & (!g551)) + ((g4) & (g1) & (!g517) & (!g549) & (!g550) & (g551)) + ((g4) & (g1) & (!g517) & (!g549) & (g550) & (!g551)) + ((g4) & (g1) & (!g517) & (!g549) & (g550) & (g551)) + ((g4) & (g1) & (!g517) & (g549) & (!g550) & (!g551)) + ((g4) & (g1) & (!g517) & (g549) & (!g550) & (g551)) + ((g4) & (g1) & (!g517) & (g549) & (g550) & (!g551)) + ((g4) & (g1) & (!g517) & (g549) & (g550) & (g551)) + ((g4) & (g1) & (g517) & (!g549) & (!g550) & (!g551)) + ((g4) & (g1) & (g517) & (!g549) & (!g550) & (g551)) + ((g4) & (g1) & (g517) & (!g549) & (g550) & (!g551)) + ((g4) & (g1) & (g517) & (!g549) & (g550) & (g551)) + ((g4) & (g1) & (g517) & (g549) & (!g550) & (!g551)) + ((g4) & (g1) & (g517) & (g549) & (!g550) & (g551)));
	assign g553 = (((!g516) & (g552)));
	assign g554 = (((!g4) & (!g549) & (!g550) & (!g516) & (!g552)) + ((!g4) & (!g549) & (!g550) & (g516) & (!g552)) + ((!g4) & (!g549) & (!g550) & (g516) & (g552)) + ((!g4) & (!g549) & (g550) & (!g516) & (g552)) + ((!g4) & (g549) & (g550) & (!g516) & (!g552)) + ((!g4) & (g549) & (g550) & (!g516) & (g552)) + ((!g4) & (g549) & (g550) & (g516) & (!g552)) + ((!g4) & (g549) & (g550) & (g516) & (g552)) + ((g4) & (!g549) & (g550) & (!g516) & (!g552)) + ((g4) & (!g549) & (g550) & (!g516) & (g552)) + ((g4) & (!g549) & (g550) & (g516) & (!g552)) + ((g4) & (!g549) & (g550) & (g516) & (g552)) + ((g4) & (g549) & (!g550) & (!g516) & (!g552)) + ((g4) & (g549) & (!g550) & (g516) & (!g552)) + ((g4) & (g549) & (!g550) & (g516) & (g552)) + ((g4) & (g549) & (g550) & (!g516) & (g552)));
	assign g555 = (((!g8) & (!g519) & (g548) & (!g516) & (!g552)) + ((!g8) & (!g519) & (g548) & (g516) & (!g552)) + ((!g8) & (!g519) & (g548) & (g516) & (g552)) + ((!g8) & (g519) & (!g548) & (!g516) & (!g552)) + ((!g8) & (g519) & (!g548) & (!g516) & (g552)) + ((!g8) & (g519) & (!g548) & (g516) & (!g552)) + ((!g8) & (g519) & (!g548) & (g516) & (g552)) + ((!g8) & (g519) & (g548) & (!g516) & (g552)) + ((g8) & (!g519) & (!g548) & (!g516) & (!g552)) + ((g8) & (!g519) & (!g548) & (g516) & (!g552)) + ((g8) & (!g519) & (!g548) & (g516) & (g552)) + ((g8) & (g519) & (!g548) & (!g516) & (g552)) + ((g8) & (g519) & (g548) & (!g516) & (!g552)) + ((g8) & (g519) & (g548) & (!g516) & (g552)) + ((g8) & (g519) & (g548) & (g516) & (!g552)) + ((g8) & (g519) & (g548) & (g516) & (g552)));
	assign g556 = (((!g18) & (!g27) & (g521) & (g547)) + ((!g18) & (g27) & (!g521) & (g547)) + ((!g18) & (g27) & (g521) & (!g547)) + ((!g18) & (g27) & (g521) & (g547)) + ((g18) & (!g27) & (!g521) & (!g547)) + ((g18) & (!g27) & (!g521) & (g547)) + ((g18) & (!g27) & (g521) & (!g547)) + ((g18) & (g27) & (!g521) & (!g547)));
	assign g557 = (((!g520) & (!g516) & (!g552) & (g556)) + ((!g520) & (g516) & (!g552) & (g556)) + ((!g520) & (g516) & (g552) & (g556)) + ((g520) & (!g516) & (!g552) & (!g556)) + ((g520) & (!g516) & (g552) & (!g556)) + ((g520) & (!g516) & (g552) & (g556)) + ((g520) & (g516) & (!g552) & (!g556)) + ((g520) & (g516) & (g552) & (!g556)));
	assign g558 = (((!g27) & (!g521) & (g547) & (!g516) & (!g552)) + ((!g27) & (!g521) & (g547) & (g516) & (!g552)) + ((!g27) & (!g521) & (g547) & (g516) & (g552)) + ((!g27) & (g521) & (!g547) & (!g516) & (!g552)) + ((!g27) & (g521) & (!g547) & (!g516) & (g552)) + ((!g27) & (g521) & (!g547) & (g516) & (!g552)) + ((!g27) & (g521) & (!g547) & (g516) & (g552)) + ((!g27) & (g521) & (g547) & (!g516) & (g552)) + ((g27) & (!g521) & (!g547) & (!g516) & (!g552)) + ((g27) & (!g521) & (!g547) & (g516) & (!g552)) + ((g27) & (!g521) & (!g547) & (g516) & (g552)) + ((g27) & (g521) & (!g547) & (!g516) & (g552)) + ((g27) & (g521) & (g547) & (!g516) & (!g552)) + ((g27) & (g521) & (g547) & (!g516) & (g552)) + ((g27) & (g521) & (g547) & (g516) & (!g552)) + ((g27) & (g521) & (g547) & (g516) & (g552)));
	assign g559 = (((!g39) & (!g54) & (g523) & (g546)) + ((!g39) & (g54) & (!g523) & (g546)) + ((!g39) & (g54) & (g523) & (!g546)) + ((!g39) & (g54) & (g523) & (g546)) + ((g39) & (!g54) & (!g523) & (!g546)) + ((g39) & (!g54) & (!g523) & (g546)) + ((g39) & (!g54) & (g523) & (!g546)) + ((g39) & (g54) & (!g523) & (!g546)));
	assign g560 = (((!g522) & (!g516) & (!g552) & (g559)) + ((!g522) & (g516) & (!g552) & (g559)) + ((!g522) & (g516) & (g552) & (g559)) + ((g522) & (!g516) & (!g552) & (!g559)) + ((g522) & (!g516) & (g552) & (!g559)) + ((g522) & (!g516) & (g552) & (g559)) + ((g522) & (g516) & (!g552) & (!g559)) + ((g522) & (g516) & (g552) & (!g559)));
	assign g561 = (((!g54) & (!g523) & (g546) & (!g516) & (!g552)) + ((!g54) & (!g523) & (g546) & (g516) & (!g552)) + ((!g54) & (!g523) & (g546) & (g516) & (g552)) + ((!g54) & (g523) & (!g546) & (!g516) & (!g552)) + ((!g54) & (g523) & (!g546) & (!g516) & (g552)) + ((!g54) & (g523) & (!g546) & (g516) & (!g552)) + ((!g54) & (g523) & (!g546) & (g516) & (g552)) + ((!g54) & (g523) & (g546) & (!g516) & (g552)) + ((g54) & (!g523) & (!g546) & (!g516) & (!g552)) + ((g54) & (!g523) & (!g546) & (g516) & (!g552)) + ((g54) & (!g523) & (!g546) & (g516) & (g552)) + ((g54) & (g523) & (!g546) & (!g516) & (g552)) + ((g54) & (g523) & (g546) & (!g516) & (!g552)) + ((g54) & (g523) & (g546) & (!g516) & (g552)) + ((g54) & (g523) & (g546) & (g516) & (!g552)) + ((g54) & (g523) & (g546) & (g516) & (g552)));
	assign g562 = (((!g68) & (!g87) & (g525) & (g545)) + ((!g68) & (g87) & (!g525) & (g545)) + ((!g68) & (g87) & (g525) & (!g545)) + ((!g68) & (g87) & (g525) & (g545)) + ((g68) & (!g87) & (!g525) & (!g545)) + ((g68) & (!g87) & (!g525) & (g545)) + ((g68) & (!g87) & (g525) & (!g545)) + ((g68) & (g87) & (!g525) & (!g545)));
	assign g563 = (((!g524) & (!g516) & (!g552) & (g562)) + ((!g524) & (g516) & (!g552) & (g562)) + ((!g524) & (g516) & (g552) & (g562)) + ((g524) & (!g516) & (!g552) & (!g562)) + ((g524) & (!g516) & (g552) & (!g562)) + ((g524) & (!g516) & (g552) & (g562)) + ((g524) & (g516) & (!g552) & (!g562)) + ((g524) & (g516) & (g552) & (!g562)));
	assign g564 = (((!g87) & (!g525) & (g545) & (!g516) & (!g552)) + ((!g87) & (!g525) & (g545) & (g516) & (!g552)) + ((!g87) & (!g525) & (g545) & (g516) & (g552)) + ((!g87) & (g525) & (!g545) & (!g516) & (!g552)) + ((!g87) & (g525) & (!g545) & (!g516) & (g552)) + ((!g87) & (g525) & (!g545) & (g516) & (!g552)) + ((!g87) & (g525) & (!g545) & (g516) & (g552)) + ((!g87) & (g525) & (g545) & (!g516) & (g552)) + ((g87) & (!g525) & (!g545) & (!g516) & (!g552)) + ((g87) & (!g525) & (!g545) & (g516) & (!g552)) + ((g87) & (!g525) & (!g545) & (g516) & (g552)) + ((g87) & (g525) & (!g545) & (!g516) & (g552)) + ((g87) & (g525) & (g545) & (!g516) & (!g552)) + ((g87) & (g525) & (g545) & (!g516) & (g552)) + ((g87) & (g525) & (g545) & (g516) & (!g552)) + ((g87) & (g525) & (g545) & (g516) & (g552)));
	assign g565 = (((!g104) & (!g127) & (g527) & (g544)) + ((!g104) & (g127) & (!g527) & (g544)) + ((!g104) & (g127) & (g527) & (!g544)) + ((!g104) & (g127) & (g527) & (g544)) + ((g104) & (!g127) & (!g527) & (!g544)) + ((g104) & (!g127) & (!g527) & (g544)) + ((g104) & (!g127) & (g527) & (!g544)) + ((g104) & (g127) & (!g527) & (!g544)));
	assign g566 = (((!g526) & (!g516) & (!g552) & (g565)) + ((!g526) & (g516) & (!g552) & (g565)) + ((!g526) & (g516) & (g552) & (g565)) + ((g526) & (!g516) & (!g552) & (!g565)) + ((g526) & (!g516) & (g552) & (!g565)) + ((g526) & (!g516) & (g552) & (g565)) + ((g526) & (g516) & (!g552) & (!g565)) + ((g526) & (g516) & (g552) & (!g565)));
	assign g567 = (((!g127) & (!g527) & (g544) & (!g516) & (!g552)) + ((!g127) & (!g527) & (g544) & (g516) & (!g552)) + ((!g127) & (!g527) & (g544) & (g516) & (g552)) + ((!g127) & (g527) & (!g544) & (!g516) & (!g552)) + ((!g127) & (g527) & (!g544) & (!g516) & (g552)) + ((!g127) & (g527) & (!g544) & (g516) & (!g552)) + ((!g127) & (g527) & (!g544) & (g516) & (g552)) + ((!g127) & (g527) & (g544) & (!g516) & (g552)) + ((g127) & (!g527) & (!g544) & (!g516) & (!g552)) + ((g127) & (!g527) & (!g544) & (g516) & (!g552)) + ((g127) & (!g527) & (!g544) & (g516) & (g552)) + ((g127) & (g527) & (!g544) & (!g516) & (g552)) + ((g127) & (g527) & (g544) & (!g516) & (!g552)) + ((g127) & (g527) & (g544) & (!g516) & (g552)) + ((g127) & (g527) & (g544) & (g516) & (!g552)) + ((g127) & (g527) & (g544) & (g516) & (g552)));
	assign g568 = (((!g147) & (!g174) & (g529) & (g543)) + ((!g147) & (g174) & (!g529) & (g543)) + ((!g147) & (g174) & (g529) & (!g543)) + ((!g147) & (g174) & (g529) & (g543)) + ((g147) & (!g174) & (!g529) & (!g543)) + ((g147) & (!g174) & (!g529) & (g543)) + ((g147) & (!g174) & (g529) & (!g543)) + ((g147) & (g174) & (!g529) & (!g543)));
	assign g569 = (((!g528) & (!g516) & (!g552) & (g568)) + ((!g528) & (g516) & (!g552) & (g568)) + ((!g528) & (g516) & (g552) & (g568)) + ((g528) & (!g516) & (!g552) & (!g568)) + ((g528) & (!g516) & (g552) & (!g568)) + ((g528) & (!g516) & (g552) & (g568)) + ((g528) & (g516) & (!g552) & (!g568)) + ((g528) & (g516) & (g552) & (!g568)));
	assign g570 = (((!g174) & (!g529) & (g543) & (!g516) & (!g552)) + ((!g174) & (!g529) & (g543) & (g516) & (!g552)) + ((!g174) & (!g529) & (g543) & (g516) & (g552)) + ((!g174) & (g529) & (!g543) & (!g516) & (!g552)) + ((!g174) & (g529) & (!g543) & (!g516) & (g552)) + ((!g174) & (g529) & (!g543) & (g516) & (!g552)) + ((!g174) & (g529) & (!g543) & (g516) & (g552)) + ((!g174) & (g529) & (g543) & (!g516) & (g552)) + ((g174) & (!g529) & (!g543) & (!g516) & (!g552)) + ((g174) & (!g529) & (!g543) & (g516) & (!g552)) + ((g174) & (!g529) & (!g543) & (g516) & (g552)) + ((g174) & (g529) & (!g543) & (!g516) & (g552)) + ((g174) & (g529) & (g543) & (!g516) & (!g552)) + ((g174) & (g529) & (g543) & (!g516) & (g552)) + ((g174) & (g529) & (g543) & (g516) & (!g552)) + ((g174) & (g529) & (g543) & (g516) & (g552)));
	assign g571 = (((!g198) & (!g229) & (g531) & (g542)) + ((!g198) & (g229) & (!g531) & (g542)) + ((!g198) & (g229) & (g531) & (!g542)) + ((!g198) & (g229) & (g531) & (g542)) + ((g198) & (!g229) & (!g531) & (!g542)) + ((g198) & (!g229) & (!g531) & (g542)) + ((g198) & (!g229) & (g531) & (!g542)) + ((g198) & (g229) & (!g531) & (!g542)));
	assign g572 = (((!g530) & (!g516) & (!g552) & (g571)) + ((!g530) & (g516) & (!g552) & (g571)) + ((!g530) & (g516) & (g552) & (g571)) + ((g530) & (!g516) & (!g552) & (!g571)) + ((g530) & (!g516) & (g552) & (!g571)) + ((g530) & (!g516) & (g552) & (g571)) + ((g530) & (g516) & (!g552) & (!g571)) + ((g530) & (g516) & (g552) & (!g571)));
	assign g573 = (((!g229) & (!g531) & (g542) & (!g516) & (!g552)) + ((!g229) & (!g531) & (g542) & (g516) & (!g552)) + ((!g229) & (!g531) & (g542) & (g516) & (g552)) + ((!g229) & (g531) & (!g542) & (!g516) & (!g552)) + ((!g229) & (g531) & (!g542) & (!g516) & (g552)) + ((!g229) & (g531) & (!g542) & (g516) & (!g552)) + ((!g229) & (g531) & (!g542) & (g516) & (g552)) + ((!g229) & (g531) & (g542) & (!g516) & (g552)) + ((g229) & (!g531) & (!g542) & (!g516) & (!g552)) + ((g229) & (!g531) & (!g542) & (g516) & (!g552)) + ((g229) & (!g531) & (!g542) & (g516) & (g552)) + ((g229) & (g531) & (!g542) & (!g516) & (g552)) + ((g229) & (g531) & (g542) & (!g516) & (!g552)) + ((g229) & (g531) & (g542) & (!g516) & (g552)) + ((g229) & (g531) & (g542) & (g516) & (!g552)) + ((g229) & (g531) & (g542) & (g516) & (g552)));
	assign g574 = (((!g255) & (!g290) & (g533) & (g541)) + ((!g255) & (g290) & (!g533) & (g541)) + ((!g255) & (g290) & (g533) & (!g541)) + ((!g255) & (g290) & (g533) & (g541)) + ((g255) & (!g290) & (!g533) & (!g541)) + ((g255) & (!g290) & (!g533) & (g541)) + ((g255) & (!g290) & (g533) & (!g541)) + ((g255) & (g290) & (!g533) & (!g541)));
	assign g575 = (((!g532) & (!g516) & (!g552) & (g574)) + ((!g532) & (g516) & (!g552) & (g574)) + ((!g532) & (g516) & (g552) & (g574)) + ((g532) & (!g516) & (!g552) & (!g574)) + ((g532) & (!g516) & (g552) & (!g574)) + ((g532) & (!g516) & (g552) & (g574)) + ((g532) & (g516) & (!g552) & (!g574)) + ((g532) & (g516) & (g552) & (!g574)));
	assign g576 = (((!g290) & (!g533) & (g541) & (!g516) & (!g552)) + ((!g290) & (!g533) & (g541) & (g516) & (!g552)) + ((!g290) & (!g533) & (g541) & (g516) & (g552)) + ((!g290) & (g533) & (!g541) & (!g516) & (!g552)) + ((!g290) & (g533) & (!g541) & (!g516) & (g552)) + ((!g290) & (g533) & (!g541) & (g516) & (!g552)) + ((!g290) & (g533) & (!g541) & (g516) & (g552)) + ((!g290) & (g533) & (g541) & (!g516) & (g552)) + ((g290) & (!g533) & (!g541) & (!g516) & (!g552)) + ((g290) & (!g533) & (!g541) & (g516) & (!g552)) + ((g290) & (!g533) & (!g541) & (g516) & (g552)) + ((g290) & (g533) & (!g541) & (!g516) & (g552)) + ((g290) & (g533) & (g541) & (!g516) & (!g552)) + ((g290) & (g533) & (g541) & (!g516) & (g552)) + ((g290) & (g533) & (g541) & (g516) & (!g552)) + ((g290) & (g533) & (g541) & (g516) & (g552)));
	assign g577 = (((!g319) & (!g358) & (g535) & (g540)) + ((!g319) & (g358) & (!g535) & (g540)) + ((!g319) & (g358) & (g535) & (!g540)) + ((!g319) & (g358) & (g535) & (g540)) + ((g319) & (!g358) & (!g535) & (!g540)) + ((g319) & (!g358) & (!g535) & (g540)) + ((g319) & (!g358) & (g535) & (!g540)) + ((g319) & (g358) & (!g535) & (!g540)));
	assign g578 = (((!g534) & (!g516) & (!g552) & (g577)) + ((!g534) & (g516) & (!g552) & (g577)) + ((!g534) & (g516) & (g552) & (g577)) + ((g534) & (!g516) & (!g552) & (!g577)) + ((g534) & (!g516) & (g552) & (!g577)) + ((g534) & (!g516) & (g552) & (g577)) + ((g534) & (g516) & (!g552) & (!g577)) + ((g534) & (g516) & (g552) & (!g577)));
	assign g579 = (((!g358) & (!g535) & (g540) & (!g516) & (!g552)) + ((!g358) & (!g535) & (g540) & (g516) & (!g552)) + ((!g358) & (!g535) & (g540) & (g516) & (g552)) + ((!g358) & (g535) & (!g540) & (!g516) & (!g552)) + ((!g358) & (g535) & (!g540) & (!g516) & (g552)) + ((!g358) & (g535) & (!g540) & (g516) & (!g552)) + ((!g358) & (g535) & (!g540) & (g516) & (g552)) + ((!g358) & (g535) & (g540) & (!g516) & (g552)) + ((g358) & (!g535) & (!g540) & (!g516) & (!g552)) + ((g358) & (!g535) & (!g540) & (g516) & (!g552)) + ((g358) & (!g535) & (!g540) & (g516) & (g552)) + ((g358) & (g535) & (!g540) & (!g516) & (g552)) + ((g358) & (g535) & (g540) & (!g516) & (!g552)) + ((g358) & (g535) & (g540) & (!g516) & (g552)) + ((g358) & (g535) & (g540) & (g516) & (!g552)) + ((g358) & (g535) & (g540) & (g516) & (g552)));
	assign g580 = (((!g390) & (!g433) & (g537) & (g539)) + ((!g390) & (g433) & (!g537) & (g539)) + ((!g390) & (g433) & (g537) & (!g539)) + ((!g390) & (g433) & (g537) & (g539)) + ((g390) & (!g433) & (!g537) & (!g539)) + ((g390) & (!g433) & (!g537) & (g539)) + ((g390) & (!g433) & (g537) & (!g539)) + ((g390) & (g433) & (!g537) & (!g539)));
	assign g581 = (((!g536) & (!g516) & (!g552) & (g580)) + ((!g536) & (g516) & (!g552) & (g580)) + ((!g536) & (g516) & (g552) & (g580)) + ((g536) & (!g516) & (!g552) & (!g580)) + ((g536) & (!g516) & (g552) & (!g580)) + ((g536) & (!g516) & (g552) & (g580)) + ((g536) & (g516) & (!g552) & (!g580)) + ((g536) & (g516) & (g552) & (!g580)));
	assign g582 = (((!g433) & (!g537) & (g539) & (!g516) & (!g552)) + ((!g433) & (!g537) & (g539) & (g516) & (!g552)) + ((!g433) & (!g537) & (g539) & (g516) & (g552)) + ((!g433) & (g537) & (!g539) & (!g516) & (!g552)) + ((!g433) & (g537) & (!g539) & (!g516) & (g552)) + ((!g433) & (g537) & (!g539) & (g516) & (!g552)) + ((!g433) & (g537) & (!g539) & (g516) & (g552)) + ((!g433) & (g537) & (g539) & (!g516) & (g552)) + ((g433) & (!g537) & (!g539) & (!g516) & (!g552)) + ((g433) & (!g537) & (!g539) & (g516) & (!g552)) + ((g433) & (!g537) & (!g539) & (g516) & (g552)) + ((g433) & (g537) & (!g539) & (!g516) & (g552)) + ((g433) & (g537) & (g539) & (!g516) & (!g552)) + ((g433) & (g537) & (g539) & (!g516) & (g552)) + ((g433) & (g537) & (g539) & (g516) & (!g552)) + ((g433) & (g537) & (g539) & (g516) & (g552)));
	assign g583 = (((!g468) & (!ax80x) & (!g515) & (g538)) + ((!g468) & (!ax80x) & (g515) & (g538)) + ((!g468) & (ax80x) & (!g515) & (!g538)) + ((!g468) & (ax80x) & (!g515) & (g538)) + ((g468) & (!ax80x) & (!g515) & (!g538)) + ((g468) & (!ax80x) & (g515) & (!g538)) + ((g468) & (ax80x) & (g515) & (!g538)) + ((g468) & (ax80x) & (g515) & (g538)));
	assign g584 = (((!ax80x) & (!ax81x) & (!g515) & (!g516) & (!g552) & (g583)) + ((!ax80x) & (!ax81x) & (!g515) & (!g516) & (g552) & (!g583)) + ((!ax80x) & (!ax81x) & (!g515) & (!g516) & (g552) & (g583)) + ((!ax80x) & (!ax81x) & (!g515) & (g516) & (!g552) & (g583)) + ((!ax80x) & (!ax81x) & (!g515) & (g516) & (g552) & (g583)) + ((!ax80x) & (!ax81x) & (g515) & (!g516) & (!g552) & (!g583)) + ((!ax80x) & (!ax81x) & (g515) & (g516) & (!g552) & (!g583)) + ((!ax80x) & (!ax81x) & (g515) & (g516) & (g552) & (!g583)) + ((!ax80x) & (ax81x) & (!g515) & (!g516) & (!g552) & (!g583)) + ((!ax80x) & (ax81x) & (!g515) & (g516) & (!g552) & (!g583)) + ((!ax80x) & (ax81x) & (!g515) & (g516) & (g552) & (!g583)) + ((!ax80x) & (ax81x) & (g515) & (!g516) & (!g552) & (g583)) + ((!ax80x) & (ax81x) & (g515) & (!g516) & (g552) & (!g583)) + ((!ax80x) & (ax81x) & (g515) & (!g516) & (g552) & (g583)) + ((!ax80x) & (ax81x) & (g515) & (g516) & (!g552) & (g583)) + ((!ax80x) & (ax81x) & (g515) & (g516) & (g552) & (g583)) + ((ax80x) & (!ax81x) & (!g515) & (!g516) & (!g552) & (!g583)) + ((ax80x) & (!ax81x) & (!g515) & (g516) & (!g552) & (!g583)) + ((ax80x) & (!ax81x) & (!g515) & (g516) & (g552) & (!g583)) + ((ax80x) & (!ax81x) & (g515) & (!g516) & (!g552) & (!g583)) + ((ax80x) & (!ax81x) & (g515) & (g516) & (!g552) & (!g583)) + ((ax80x) & (!ax81x) & (g515) & (g516) & (g552) & (!g583)) + ((ax80x) & (ax81x) & (!g515) & (!g516) & (!g552) & (g583)) + ((ax80x) & (ax81x) & (!g515) & (!g516) & (g552) & (!g583)) + ((ax80x) & (ax81x) & (!g515) & (!g516) & (g552) & (g583)) + ((ax80x) & (ax81x) & (!g515) & (g516) & (!g552) & (g583)) + ((ax80x) & (ax81x) & (!g515) & (g516) & (g552) & (g583)) + ((ax80x) & (ax81x) & (g515) & (!g516) & (!g552) & (g583)) + ((ax80x) & (ax81x) & (g515) & (!g516) & (g552) & (!g583)) + ((ax80x) & (ax81x) & (g515) & (!g516) & (g552) & (g583)) + ((ax80x) & (ax81x) & (g515) & (g516) & (!g552) & (g583)) + ((ax80x) & (ax81x) & (g515) & (g516) & (g552) & (g583)));
	assign g585 = (((!ax80x) & (!g515) & (!g538) & (!g516) & (g552)) + ((!ax80x) & (!g515) & (g538) & (!g516) & (!g552)) + ((!ax80x) & (!g515) & (g538) & (!g516) & (g552)) + ((!ax80x) & (!g515) & (g538) & (g516) & (!g552)) + ((!ax80x) & (!g515) & (g538) & (g516) & (g552)) + ((!ax80x) & (g515) & (g538) & (!g516) & (!g552)) + ((!ax80x) & (g515) & (g538) & (g516) & (!g552)) + ((!ax80x) & (g515) & (g538) & (g516) & (g552)) + ((ax80x) & (!g515) & (!g538) & (!g516) & (!g552)) + ((ax80x) & (!g515) & (!g538) & (g516) & (!g552)) + ((ax80x) & (!g515) & (!g538) & (g516) & (g552)) + ((ax80x) & (g515) & (!g538) & (!g516) & (!g552)) + ((ax80x) & (g515) & (!g538) & (!g516) & (g552)) + ((ax80x) & (g515) & (!g538) & (g516) & (!g552)) + ((ax80x) & (g515) & (!g538) & (g516) & (g552)) + ((ax80x) & (g515) & (g538) & (!g516) & (g552)));
	assign g586 = (((!ax76x) & (!ax77x)));
	assign g587 = (((!g515) & (!ax78x) & (!ax79x) & (!g516) & (!g552) & (!g586)) + ((!g515) & (!ax78x) & (!ax79x) & (g516) & (!g552) & (!g586)) + ((!g515) & (!ax78x) & (!ax79x) & (g516) & (g552) & (!g586)) + ((!g515) & (!ax78x) & (ax79x) & (!g516) & (g552) & (!g586)) + ((!g515) & (ax78x) & (ax79x) & (!g516) & (g552) & (!g586)) + ((!g515) & (ax78x) & (ax79x) & (!g516) & (g552) & (g586)) + ((g515) & (!ax78x) & (!ax79x) & (!g516) & (!g552) & (!g586)) + ((g515) & (!ax78x) & (!ax79x) & (!g516) & (!g552) & (g586)) + ((g515) & (!ax78x) & (!ax79x) & (!g516) & (g552) & (!g586)) + ((g515) & (!ax78x) & (!ax79x) & (g516) & (!g552) & (!g586)) + ((g515) & (!ax78x) & (!ax79x) & (g516) & (!g552) & (g586)) + ((g515) & (!ax78x) & (!ax79x) & (g516) & (g552) & (!g586)) + ((g515) & (!ax78x) & (!ax79x) & (g516) & (g552) & (g586)) + ((g515) & (!ax78x) & (ax79x) & (!g516) & (!g552) & (!g586)) + ((g515) & (!ax78x) & (ax79x) & (!g516) & (g552) & (!g586)) + ((g515) & (!ax78x) & (ax79x) & (!g516) & (g552) & (g586)) + ((g515) & (!ax78x) & (ax79x) & (g516) & (!g552) & (!g586)) + ((g515) & (!ax78x) & (ax79x) & (g516) & (g552) & (!g586)) + ((g515) & (ax78x) & (!ax79x) & (!g516) & (g552) & (!g586)) + ((g515) & (ax78x) & (!ax79x) & (!g516) & (g552) & (g586)) + ((g515) & (ax78x) & (ax79x) & (!g516) & (!g552) & (!g586)) + ((g515) & (ax78x) & (ax79x) & (!g516) & (!g552) & (g586)) + ((g515) & (ax78x) & (ax79x) & (!g516) & (g552) & (!g586)) + ((g515) & (ax78x) & (ax79x) & (!g516) & (g552) & (g586)) + ((g515) & (ax78x) & (ax79x) & (g516) & (!g552) & (!g586)) + ((g515) & (ax78x) & (ax79x) & (g516) & (!g552) & (g586)) + ((g515) & (ax78x) & (ax79x) & (g516) & (g552) & (!g586)) + ((g515) & (ax78x) & (ax79x) & (g516) & (g552) & (g586)));
	assign g588 = (((!g433) & (!g468) & (g584) & (g585) & (g587)) + ((!g433) & (g468) & (g584) & (!g585) & (g587)) + ((!g433) & (g468) & (g584) & (g585) & (!g587)) + ((!g433) & (g468) & (g584) & (g585) & (g587)) + ((g433) & (!g468) & (!g584) & (g585) & (g587)) + ((g433) & (!g468) & (g584) & (!g585) & (!g587)) + ((g433) & (!g468) & (g584) & (!g585) & (g587)) + ((g433) & (!g468) & (g584) & (g585) & (!g587)) + ((g433) & (!g468) & (g584) & (g585) & (g587)) + ((g433) & (g468) & (!g584) & (!g585) & (g587)) + ((g433) & (g468) & (!g584) & (g585) & (!g587)) + ((g433) & (g468) & (!g584) & (g585) & (g587)) + ((g433) & (g468) & (g584) & (!g585) & (!g587)) + ((g433) & (g468) & (g584) & (!g585) & (g587)) + ((g433) & (g468) & (g584) & (g585) & (!g587)) + ((g433) & (g468) & (g584) & (g585) & (g587)));
	assign g589 = (((!g358) & (!g390) & (g581) & (g582) & (g588)) + ((!g358) & (g390) & (g581) & (!g582) & (g588)) + ((!g358) & (g390) & (g581) & (g582) & (!g588)) + ((!g358) & (g390) & (g581) & (g582) & (g588)) + ((g358) & (!g390) & (!g581) & (g582) & (g588)) + ((g358) & (!g390) & (g581) & (!g582) & (!g588)) + ((g358) & (!g390) & (g581) & (!g582) & (g588)) + ((g358) & (!g390) & (g581) & (g582) & (!g588)) + ((g358) & (!g390) & (g581) & (g582) & (g588)) + ((g358) & (g390) & (!g581) & (!g582) & (g588)) + ((g358) & (g390) & (!g581) & (g582) & (!g588)) + ((g358) & (g390) & (!g581) & (g582) & (g588)) + ((g358) & (g390) & (g581) & (!g582) & (!g588)) + ((g358) & (g390) & (g581) & (!g582) & (g588)) + ((g358) & (g390) & (g581) & (g582) & (!g588)) + ((g358) & (g390) & (g581) & (g582) & (g588)));
	assign g590 = (((!g290) & (!g319) & (g578) & (g579) & (g589)) + ((!g290) & (g319) & (g578) & (!g579) & (g589)) + ((!g290) & (g319) & (g578) & (g579) & (!g589)) + ((!g290) & (g319) & (g578) & (g579) & (g589)) + ((g290) & (!g319) & (!g578) & (g579) & (g589)) + ((g290) & (!g319) & (g578) & (!g579) & (!g589)) + ((g290) & (!g319) & (g578) & (!g579) & (g589)) + ((g290) & (!g319) & (g578) & (g579) & (!g589)) + ((g290) & (!g319) & (g578) & (g579) & (g589)) + ((g290) & (g319) & (!g578) & (!g579) & (g589)) + ((g290) & (g319) & (!g578) & (g579) & (!g589)) + ((g290) & (g319) & (!g578) & (g579) & (g589)) + ((g290) & (g319) & (g578) & (!g579) & (!g589)) + ((g290) & (g319) & (g578) & (!g579) & (g589)) + ((g290) & (g319) & (g578) & (g579) & (!g589)) + ((g290) & (g319) & (g578) & (g579) & (g589)));
	assign g591 = (((!g229) & (!g255) & (g575) & (g576) & (g590)) + ((!g229) & (g255) & (g575) & (!g576) & (g590)) + ((!g229) & (g255) & (g575) & (g576) & (!g590)) + ((!g229) & (g255) & (g575) & (g576) & (g590)) + ((g229) & (!g255) & (!g575) & (g576) & (g590)) + ((g229) & (!g255) & (g575) & (!g576) & (!g590)) + ((g229) & (!g255) & (g575) & (!g576) & (g590)) + ((g229) & (!g255) & (g575) & (g576) & (!g590)) + ((g229) & (!g255) & (g575) & (g576) & (g590)) + ((g229) & (g255) & (!g575) & (!g576) & (g590)) + ((g229) & (g255) & (!g575) & (g576) & (!g590)) + ((g229) & (g255) & (!g575) & (g576) & (g590)) + ((g229) & (g255) & (g575) & (!g576) & (!g590)) + ((g229) & (g255) & (g575) & (!g576) & (g590)) + ((g229) & (g255) & (g575) & (g576) & (!g590)) + ((g229) & (g255) & (g575) & (g576) & (g590)));
	assign g592 = (((!g174) & (!g198) & (g572) & (g573) & (g591)) + ((!g174) & (g198) & (g572) & (!g573) & (g591)) + ((!g174) & (g198) & (g572) & (g573) & (!g591)) + ((!g174) & (g198) & (g572) & (g573) & (g591)) + ((g174) & (!g198) & (!g572) & (g573) & (g591)) + ((g174) & (!g198) & (g572) & (!g573) & (!g591)) + ((g174) & (!g198) & (g572) & (!g573) & (g591)) + ((g174) & (!g198) & (g572) & (g573) & (!g591)) + ((g174) & (!g198) & (g572) & (g573) & (g591)) + ((g174) & (g198) & (!g572) & (!g573) & (g591)) + ((g174) & (g198) & (!g572) & (g573) & (!g591)) + ((g174) & (g198) & (!g572) & (g573) & (g591)) + ((g174) & (g198) & (g572) & (!g573) & (!g591)) + ((g174) & (g198) & (g572) & (!g573) & (g591)) + ((g174) & (g198) & (g572) & (g573) & (!g591)) + ((g174) & (g198) & (g572) & (g573) & (g591)));
	assign g593 = (((!g127) & (!g147) & (g569) & (g570) & (g592)) + ((!g127) & (g147) & (g569) & (!g570) & (g592)) + ((!g127) & (g147) & (g569) & (g570) & (!g592)) + ((!g127) & (g147) & (g569) & (g570) & (g592)) + ((g127) & (!g147) & (!g569) & (g570) & (g592)) + ((g127) & (!g147) & (g569) & (!g570) & (!g592)) + ((g127) & (!g147) & (g569) & (!g570) & (g592)) + ((g127) & (!g147) & (g569) & (g570) & (!g592)) + ((g127) & (!g147) & (g569) & (g570) & (g592)) + ((g127) & (g147) & (!g569) & (!g570) & (g592)) + ((g127) & (g147) & (!g569) & (g570) & (!g592)) + ((g127) & (g147) & (!g569) & (g570) & (g592)) + ((g127) & (g147) & (g569) & (!g570) & (!g592)) + ((g127) & (g147) & (g569) & (!g570) & (g592)) + ((g127) & (g147) & (g569) & (g570) & (!g592)) + ((g127) & (g147) & (g569) & (g570) & (g592)));
	assign g594 = (((!g87) & (!g104) & (g566) & (g567) & (g593)) + ((!g87) & (g104) & (g566) & (!g567) & (g593)) + ((!g87) & (g104) & (g566) & (g567) & (!g593)) + ((!g87) & (g104) & (g566) & (g567) & (g593)) + ((g87) & (!g104) & (!g566) & (g567) & (g593)) + ((g87) & (!g104) & (g566) & (!g567) & (!g593)) + ((g87) & (!g104) & (g566) & (!g567) & (g593)) + ((g87) & (!g104) & (g566) & (g567) & (!g593)) + ((g87) & (!g104) & (g566) & (g567) & (g593)) + ((g87) & (g104) & (!g566) & (!g567) & (g593)) + ((g87) & (g104) & (!g566) & (g567) & (!g593)) + ((g87) & (g104) & (!g566) & (g567) & (g593)) + ((g87) & (g104) & (g566) & (!g567) & (!g593)) + ((g87) & (g104) & (g566) & (!g567) & (g593)) + ((g87) & (g104) & (g566) & (g567) & (!g593)) + ((g87) & (g104) & (g566) & (g567) & (g593)));
	assign g595 = (((!g54) & (!g68) & (g563) & (g564) & (g594)) + ((!g54) & (g68) & (g563) & (!g564) & (g594)) + ((!g54) & (g68) & (g563) & (g564) & (!g594)) + ((!g54) & (g68) & (g563) & (g564) & (g594)) + ((g54) & (!g68) & (!g563) & (g564) & (g594)) + ((g54) & (!g68) & (g563) & (!g564) & (!g594)) + ((g54) & (!g68) & (g563) & (!g564) & (g594)) + ((g54) & (!g68) & (g563) & (g564) & (!g594)) + ((g54) & (!g68) & (g563) & (g564) & (g594)) + ((g54) & (g68) & (!g563) & (!g564) & (g594)) + ((g54) & (g68) & (!g563) & (g564) & (!g594)) + ((g54) & (g68) & (!g563) & (g564) & (g594)) + ((g54) & (g68) & (g563) & (!g564) & (!g594)) + ((g54) & (g68) & (g563) & (!g564) & (g594)) + ((g54) & (g68) & (g563) & (g564) & (!g594)) + ((g54) & (g68) & (g563) & (g564) & (g594)));
	assign g596 = (((!g27) & (!g39) & (g560) & (g561) & (g595)) + ((!g27) & (g39) & (g560) & (!g561) & (g595)) + ((!g27) & (g39) & (g560) & (g561) & (!g595)) + ((!g27) & (g39) & (g560) & (g561) & (g595)) + ((g27) & (!g39) & (!g560) & (g561) & (g595)) + ((g27) & (!g39) & (g560) & (!g561) & (!g595)) + ((g27) & (!g39) & (g560) & (!g561) & (g595)) + ((g27) & (!g39) & (g560) & (g561) & (!g595)) + ((g27) & (!g39) & (g560) & (g561) & (g595)) + ((g27) & (g39) & (!g560) & (!g561) & (g595)) + ((g27) & (g39) & (!g560) & (g561) & (!g595)) + ((g27) & (g39) & (!g560) & (g561) & (g595)) + ((g27) & (g39) & (g560) & (!g561) & (!g595)) + ((g27) & (g39) & (g560) & (!g561) & (g595)) + ((g27) & (g39) & (g560) & (g561) & (!g595)) + ((g27) & (g39) & (g560) & (g561) & (g595)));
	assign g597 = (((!g8) & (!g18) & (g557) & (g558) & (g596)) + ((!g8) & (g18) & (g557) & (!g558) & (g596)) + ((!g8) & (g18) & (g557) & (g558) & (!g596)) + ((!g8) & (g18) & (g557) & (g558) & (g596)) + ((g8) & (!g18) & (!g557) & (g558) & (g596)) + ((g8) & (!g18) & (g557) & (!g558) & (!g596)) + ((g8) & (!g18) & (g557) & (!g558) & (g596)) + ((g8) & (!g18) & (g557) & (g558) & (!g596)) + ((g8) & (!g18) & (g557) & (g558) & (g596)) + ((g8) & (g18) & (!g557) & (!g558) & (g596)) + ((g8) & (g18) & (!g557) & (g558) & (!g596)) + ((g8) & (g18) & (!g557) & (g558) & (g596)) + ((g8) & (g18) & (g557) & (!g558) & (!g596)) + ((g8) & (g18) & (g557) & (!g558) & (g596)) + ((g8) & (g18) & (g557) & (g558) & (!g596)) + ((g8) & (g18) & (g557) & (g558) & (g596)));
	assign g598 = (((!g2) & (!g8) & (g519) & (g548)) + ((!g2) & (g8) & (!g519) & (g548)) + ((!g2) & (g8) & (g519) & (!g548)) + ((!g2) & (g8) & (g519) & (g548)) + ((g2) & (!g8) & (!g519) & (!g548)) + ((g2) & (!g8) & (!g519) & (g548)) + ((g2) & (!g8) & (g519) & (!g548)) + ((g2) & (g8) & (!g519) & (!g548)));
	assign g599 = (((!g518) & (!g516) & (!g552) & (g598)) + ((!g518) & (g516) & (!g552) & (g598)) + ((!g518) & (g516) & (g552) & (g598)) + ((g518) & (!g516) & (!g552) & (!g598)) + ((g518) & (!g516) & (g552) & (!g598)) + ((g518) & (!g516) & (g552) & (g598)) + ((g518) & (g516) & (!g552) & (!g598)) + ((g518) & (g516) & (g552) & (!g598)));
	assign g600 = (((!g4) & (!g2) & (!g555) & (!g597) & (g599)) + ((!g4) & (!g2) & (!g555) & (g597) & (g599)) + ((!g4) & (!g2) & (g555) & (!g597) & (g599)) + ((!g4) & (!g2) & (g555) & (g597) & (!g599)) + ((!g4) & (!g2) & (g555) & (g597) & (g599)) + ((!g4) & (g2) & (!g555) & (!g597) & (g599)) + ((!g4) & (g2) & (!g555) & (g597) & (!g599)) + ((!g4) & (g2) & (!g555) & (g597) & (g599)) + ((!g4) & (g2) & (g555) & (!g597) & (!g599)) + ((!g4) & (g2) & (g555) & (!g597) & (g599)) + ((!g4) & (g2) & (g555) & (g597) & (!g599)) + ((!g4) & (g2) & (g555) & (g597) & (g599)) + ((g4) & (!g2) & (g555) & (g597) & (g599)) + ((g4) & (g2) & (!g555) & (g597) & (g599)) + ((g4) & (g2) & (g555) & (!g597) & (g599)) + ((g4) & (g2) & (g555) & (g597) & (g599)));
	assign g601 = (((!g4) & (!g549) & (g550)) + ((!g4) & (g549) & (!g550)) + ((!g4) & (g549) & (g550)) + ((g4) & (g549) & (g550)));
	assign g602 = (((!g517) & (!g601) & (!g516) & (!g552)) + ((!g517) & (!g601) & (g516) & (!g552)) + ((!g517) & (!g601) & (g516) & (g552)) + ((g517) & (g601) & (!g516) & (!g552)) + ((g517) & (g601) & (!g516) & (g552)) + ((g517) & (g601) & (g516) & (!g552)) + ((g517) & (g601) & (g516) & (g552)));
	assign g603 = (((!g1) & (g517) & (!g601) & (!g516) & (g552)) + ((!g1) & (g517) & (g601) & (!g516) & (g552)) + ((g1) & (!g517) & (g601) & (g516) & (!g552)) + ((g1) & (!g517) & (g601) & (g516) & (g552)) + ((g1) & (g517) & (!g601) & (!g516) & (!g552)) + ((g1) & (g517) & (!g601) & (!g516) & (g552)) + ((g1) & (g517) & (!g601) & (g516) & (!g552)) + ((g1) & (g517) & (!g601) & (g516) & (g552)) + ((g1) & (g517) & (g601) & (!g516) & (g552)));
	assign g604 = (((!g1) & (!g554) & (!g600) & (!g602) & (!g603)) + ((g1) & (!g554) & (!g600) & (!g602) & (!g603)) + ((g1) & (!g554) & (!g600) & (g602) & (!g603)) + ((g1) & (!g554) & (g600) & (!g602) & (!g603)) + ((g1) & (!g554) & (g600) & (g602) & (!g603)) + ((g1) & (g554) & (!g600) & (!g602) & (!g603)) + ((g1) & (g554) & (!g600) & (g602) & (!g603)));
	assign g605 = (((g1) & (!g554) & (g600) & (g603)) + ((g1) & (g554) & (!g600) & (!g603)) + ((g1) & (g554) & (!g600) & (g603)));
	assign g606 = (((!g4) & (!g2) & (!g555) & (!g597) & (!g599) & (!g604)) + ((!g4) & (!g2) & (!g555) & (!g597) & (g599) & (g604)) + ((!g4) & (!g2) & (!g555) & (g597) & (!g599) & (!g604)) + ((!g4) & (!g2) & (!g555) & (g597) & (g599) & (g604)) + ((!g4) & (!g2) & (g555) & (!g597) & (!g599) & (!g604)) + ((!g4) & (!g2) & (g555) & (!g597) & (g599) & (g604)) + ((!g4) & (!g2) & (g555) & (g597) & (g599) & (!g604)) + ((!g4) & (!g2) & (g555) & (g597) & (g599) & (g604)) + ((!g4) & (g2) & (!g555) & (!g597) & (!g599) & (!g604)) + ((!g4) & (g2) & (!g555) & (!g597) & (g599) & (g604)) + ((!g4) & (g2) & (!g555) & (g597) & (g599) & (!g604)) + ((!g4) & (g2) & (!g555) & (g597) & (g599) & (g604)) + ((!g4) & (g2) & (g555) & (!g597) & (g599) & (!g604)) + ((!g4) & (g2) & (g555) & (!g597) & (g599) & (g604)) + ((!g4) & (g2) & (g555) & (g597) & (g599) & (!g604)) + ((!g4) & (g2) & (g555) & (g597) & (g599) & (g604)) + ((g4) & (!g2) & (!g555) & (!g597) & (g599) & (!g604)) + ((g4) & (!g2) & (!g555) & (!g597) & (g599) & (g604)) + ((g4) & (!g2) & (!g555) & (g597) & (g599) & (!g604)) + ((g4) & (!g2) & (!g555) & (g597) & (g599) & (g604)) + ((g4) & (!g2) & (g555) & (!g597) & (g599) & (!g604)) + ((g4) & (!g2) & (g555) & (!g597) & (g599) & (g604)) + ((g4) & (!g2) & (g555) & (g597) & (!g599) & (!g604)) + ((g4) & (!g2) & (g555) & (g597) & (g599) & (g604)) + ((g4) & (g2) & (!g555) & (!g597) & (g599) & (!g604)) + ((g4) & (g2) & (!g555) & (!g597) & (g599) & (g604)) + ((g4) & (g2) & (!g555) & (g597) & (!g599) & (!g604)) + ((g4) & (g2) & (!g555) & (g597) & (g599) & (g604)) + ((g4) & (g2) & (g555) & (!g597) & (!g599) & (!g604)) + ((g4) & (g2) & (g555) & (!g597) & (g599) & (g604)) + ((g4) & (g2) & (g555) & (g597) & (!g599) & (!g604)) + ((g4) & (g2) & (g555) & (g597) & (g599) & (g604)));
	assign g607 = (((!g8) & (!g18) & (!g557) & (g558) & (g596) & (!g604)) + ((!g8) & (!g18) & (g557) & (!g558) & (!g596) & (!g604)) + ((!g8) & (!g18) & (g557) & (!g558) & (!g596) & (g604)) + ((!g8) & (!g18) & (g557) & (!g558) & (g596) & (!g604)) + ((!g8) & (!g18) & (g557) & (!g558) & (g596) & (g604)) + ((!g8) & (!g18) & (g557) & (g558) & (!g596) & (!g604)) + ((!g8) & (!g18) & (g557) & (g558) & (!g596) & (g604)) + ((!g8) & (!g18) & (g557) & (g558) & (g596) & (g604)) + ((!g8) & (g18) & (!g557) & (!g558) & (g596) & (!g604)) + ((!g8) & (g18) & (!g557) & (g558) & (!g596) & (!g604)) + ((!g8) & (g18) & (!g557) & (g558) & (g596) & (!g604)) + ((!g8) & (g18) & (g557) & (!g558) & (!g596) & (!g604)) + ((!g8) & (g18) & (g557) & (!g558) & (!g596) & (g604)) + ((!g8) & (g18) & (g557) & (!g558) & (g596) & (g604)) + ((!g8) & (g18) & (g557) & (g558) & (!g596) & (g604)) + ((!g8) & (g18) & (g557) & (g558) & (g596) & (g604)) + ((g8) & (!g18) & (!g557) & (!g558) & (!g596) & (!g604)) + ((g8) & (!g18) & (!g557) & (!g558) & (g596) & (!g604)) + ((g8) & (!g18) & (!g557) & (g558) & (!g596) & (!g604)) + ((g8) & (!g18) & (g557) & (!g558) & (!g596) & (g604)) + ((g8) & (!g18) & (g557) & (!g558) & (g596) & (g604)) + ((g8) & (!g18) & (g557) & (g558) & (!g596) & (g604)) + ((g8) & (!g18) & (g557) & (g558) & (g596) & (!g604)) + ((g8) & (!g18) & (g557) & (g558) & (g596) & (g604)) + ((g8) & (g18) & (!g557) & (!g558) & (!g596) & (!g604)) + ((g8) & (g18) & (g557) & (!g558) & (!g596) & (g604)) + ((g8) & (g18) & (g557) & (!g558) & (g596) & (!g604)) + ((g8) & (g18) & (g557) & (!g558) & (g596) & (g604)) + ((g8) & (g18) & (g557) & (g558) & (!g596) & (!g604)) + ((g8) & (g18) & (g557) & (g558) & (!g596) & (g604)) + ((g8) & (g18) & (g557) & (g558) & (g596) & (!g604)) + ((g8) & (g18) & (g557) & (g558) & (g596) & (g604)));
	assign g608 = (((!g18) & (!g558) & (g596) & (!g604)) + ((!g18) & (g558) & (!g596) & (!g604)) + ((!g18) & (g558) & (!g596) & (g604)) + ((!g18) & (g558) & (g596) & (g604)) + ((g18) & (!g558) & (!g596) & (!g604)) + ((g18) & (g558) & (!g596) & (g604)) + ((g18) & (g558) & (g596) & (!g604)) + ((g18) & (g558) & (g596) & (g604)));
	assign g609 = (((!g27) & (!g39) & (!g560) & (g561) & (g595) & (!g604)) + ((!g27) & (!g39) & (g560) & (!g561) & (!g595) & (!g604)) + ((!g27) & (!g39) & (g560) & (!g561) & (!g595) & (g604)) + ((!g27) & (!g39) & (g560) & (!g561) & (g595) & (!g604)) + ((!g27) & (!g39) & (g560) & (!g561) & (g595) & (g604)) + ((!g27) & (!g39) & (g560) & (g561) & (!g595) & (!g604)) + ((!g27) & (!g39) & (g560) & (g561) & (!g595) & (g604)) + ((!g27) & (!g39) & (g560) & (g561) & (g595) & (g604)) + ((!g27) & (g39) & (!g560) & (!g561) & (g595) & (!g604)) + ((!g27) & (g39) & (!g560) & (g561) & (!g595) & (!g604)) + ((!g27) & (g39) & (!g560) & (g561) & (g595) & (!g604)) + ((!g27) & (g39) & (g560) & (!g561) & (!g595) & (!g604)) + ((!g27) & (g39) & (g560) & (!g561) & (!g595) & (g604)) + ((!g27) & (g39) & (g560) & (!g561) & (g595) & (g604)) + ((!g27) & (g39) & (g560) & (g561) & (!g595) & (g604)) + ((!g27) & (g39) & (g560) & (g561) & (g595) & (g604)) + ((g27) & (!g39) & (!g560) & (!g561) & (!g595) & (!g604)) + ((g27) & (!g39) & (!g560) & (!g561) & (g595) & (!g604)) + ((g27) & (!g39) & (!g560) & (g561) & (!g595) & (!g604)) + ((g27) & (!g39) & (g560) & (!g561) & (!g595) & (g604)) + ((g27) & (!g39) & (g560) & (!g561) & (g595) & (g604)) + ((g27) & (!g39) & (g560) & (g561) & (!g595) & (g604)) + ((g27) & (!g39) & (g560) & (g561) & (g595) & (!g604)) + ((g27) & (!g39) & (g560) & (g561) & (g595) & (g604)) + ((g27) & (g39) & (!g560) & (!g561) & (!g595) & (!g604)) + ((g27) & (g39) & (g560) & (!g561) & (!g595) & (g604)) + ((g27) & (g39) & (g560) & (!g561) & (g595) & (!g604)) + ((g27) & (g39) & (g560) & (!g561) & (g595) & (g604)) + ((g27) & (g39) & (g560) & (g561) & (!g595) & (!g604)) + ((g27) & (g39) & (g560) & (g561) & (!g595) & (g604)) + ((g27) & (g39) & (g560) & (g561) & (g595) & (!g604)) + ((g27) & (g39) & (g560) & (g561) & (g595) & (g604)));
	assign g610 = (((!g39) & (!g561) & (g595) & (!g604)) + ((!g39) & (g561) & (!g595) & (!g604)) + ((!g39) & (g561) & (!g595) & (g604)) + ((!g39) & (g561) & (g595) & (g604)) + ((g39) & (!g561) & (!g595) & (!g604)) + ((g39) & (g561) & (!g595) & (g604)) + ((g39) & (g561) & (g595) & (!g604)) + ((g39) & (g561) & (g595) & (g604)));
	assign g611 = (((!g54) & (!g68) & (!g563) & (g564) & (g594) & (!g604)) + ((!g54) & (!g68) & (g563) & (!g564) & (!g594) & (!g604)) + ((!g54) & (!g68) & (g563) & (!g564) & (!g594) & (g604)) + ((!g54) & (!g68) & (g563) & (!g564) & (g594) & (!g604)) + ((!g54) & (!g68) & (g563) & (!g564) & (g594) & (g604)) + ((!g54) & (!g68) & (g563) & (g564) & (!g594) & (!g604)) + ((!g54) & (!g68) & (g563) & (g564) & (!g594) & (g604)) + ((!g54) & (!g68) & (g563) & (g564) & (g594) & (g604)) + ((!g54) & (g68) & (!g563) & (!g564) & (g594) & (!g604)) + ((!g54) & (g68) & (!g563) & (g564) & (!g594) & (!g604)) + ((!g54) & (g68) & (!g563) & (g564) & (g594) & (!g604)) + ((!g54) & (g68) & (g563) & (!g564) & (!g594) & (!g604)) + ((!g54) & (g68) & (g563) & (!g564) & (!g594) & (g604)) + ((!g54) & (g68) & (g563) & (!g564) & (g594) & (g604)) + ((!g54) & (g68) & (g563) & (g564) & (!g594) & (g604)) + ((!g54) & (g68) & (g563) & (g564) & (g594) & (g604)) + ((g54) & (!g68) & (!g563) & (!g564) & (!g594) & (!g604)) + ((g54) & (!g68) & (!g563) & (!g564) & (g594) & (!g604)) + ((g54) & (!g68) & (!g563) & (g564) & (!g594) & (!g604)) + ((g54) & (!g68) & (g563) & (!g564) & (!g594) & (g604)) + ((g54) & (!g68) & (g563) & (!g564) & (g594) & (g604)) + ((g54) & (!g68) & (g563) & (g564) & (!g594) & (g604)) + ((g54) & (!g68) & (g563) & (g564) & (g594) & (!g604)) + ((g54) & (!g68) & (g563) & (g564) & (g594) & (g604)) + ((g54) & (g68) & (!g563) & (!g564) & (!g594) & (!g604)) + ((g54) & (g68) & (g563) & (!g564) & (!g594) & (g604)) + ((g54) & (g68) & (g563) & (!g564) & (g594) & (!g604)) + ((g54) & (g68) & (g563) & (!g564) & (g594) & (g604)) + ((g54) & (g68) & (g563) & (g564) & (!g594) & (!g604)) + ((g54) & (g68) & (g563) & (g564) & (!g594) & (g604)) + ((g54) & (g68) & (g563) & (g564) & (g594) & (!g604)) + ((g54) & (g68) & (g563) & (g564) & (g594) & (g604)));
	assign g612 = (((!g68) & (!g564) & (g594) & (!g604)) + ((!g68) & (g564) & (!g594) & (!g604)) + ((!g68) & (g564) & (!g594) & (g604)) + ((!g68) & (g564) & (g594) & (g604)) + ((g68) & (!g564) & (!g594) & (!g604)) + ((g68) & (g564) & (!g594) & (g604)) + ((g68) & (g564) & (g594) & (!g604)) + ((g68) & (g564) & (g594) & (g604)));
	assign g613 = (((!g87) & (!g104) & (!g566) & (g567) & (g593) & (!g604)) + ((!g87) & (!g104) & (g566) & (!g567) & (!g593) & (!g604)) + ((!g87) & (!g104) & (g566) & (!g567) & (!g593) & (g604)) + ((!g87) & (!g104) & (g566) & (!g567) & (g593) & (!g604)) + ((!g87) & (!g104) & (g566) & (!g567) & (g593) & (g604)) + ((!g87) & (!g104) & (g566) & (g567) & (!g593) & (!g604)) + ((!g87) & (!g104) & (g566) & (g567) & (!g593) & (g604)) + ((!g87) & (!g104) & (g566) & (g567) & (g593) & (g604)) + ((!g87) & (g104) & (!g566) & (!g567) & (g593) & (!g604)) + ((!g87) & (g104) & (!g566) & (g567) & (!g593) & (!g604)) + ((!g87) & (g104) & (!g566) & (g567) & (g593) & (!g604)) + ((!g87) & (g104) & (g566) & (!g567) & (!g593) & (!g604)) + ((!g87) & (g104) & (g566) & (!g567) & (!g593) & (g604)) + ((!g87) & (g104) & (g566) & (!g567) & (g593) & (g604)) + ((!g87) & (g104) & (g566) & (g567) & (!g593) & (g604)) + ((!g87) & (g104) & (g566) & (g567) & (g593) & (g604)) + ((g87) & (!g104) & (!g566) & (!g567) & (!g593) & (!g604)) + ((g87) & (!g104) & (!g566) & (!g567) & (g593) & (!g604)) + ((g87) & (!g104) & (!g566) & (g567) & (!g593) & (!g604)) + ((g87) & (!g104) & (g566) & (!g567) & (!g593) & (g604)) + ((g87) & (!g104) & (g566) & (!g567) & (g593) & (g604)) + ((g87) & (!g104) & (g566) & (g567) & (!g593) & (g604)) + ((g87) & (!g104) & (g566) & (g567) & (g593) & (!g604)) + ((g87) & (!g104) & (g566) & (g567) & (g593) & (g604)) + ((g87) & (g104) & (!g566) & (!g567) & (!g593) & (!g604)) + ((g87) & (g104) & (g566) & (!g567) & (!g593) & (g604)) + ((g87) & (g104) & (g566) & (!g567) & (g593) & (!g604)) + ((g87) & (g104) & (g566) & (!g567) & (g593) & (g604)) + ((g87) & (g104) & (g566) & (g567) & (!g593) & (!g604)) + ((g87) & (g104) & (g566) & (g567) & (!g593) & (g604)) + ((g87) & (g104) & (g566) & (g567) & (g593) & (!g604)) + ((g87) & (g104) & (g566) & (g567) & (g593) & (g604)));
	assign g614 = (((!g104) & (!g567) & (g593) & (!g604)) + ((!g104) & (g567) & (!g593) & (!g604)) + ((!g104) & (g567) & (!g593) & (g604)) + ((!g104) & (g567) & (g593) & (g604)) + ((g104) & (!g567) & (!g593) & (!g604)) + ((g104) & (g567) & (!g593) & (g604)) + ((g104) & (g567) & (g593) & (!g604)) + ((g104) & (g567) & (g593) & (g604)));
	assign g615 = (((!g127) & (!g147) & (!g569) & (g570) & (g592) & (!g604)) + ((!g127) & (!g147) & (g569) & (!g570) & (!g592) & (!g604)) + ((!g127) & (!g147) & (g569) & (!g570) & (!g592) & (g604)) + ((!g127) & (!g147) & (g569) & (!g570) & (g592) & (!g604)) + ((!g127) & (!g147) & (g569) & (!g570) & (g592) & (g604)) + ((!g127) & (!g147) & (g569) & (g570) & (!g592) & (!g604)) + ((!g127) & (!g147) & (g569) & (g570) & (!g592) & (g604)) + ((!g127) & (!g147) & (g569) & (g570) & (g592) & (g604)) + ((!g127) & (g147) & (!g569) & (!g570) & (g592) & (!g604)) + ((!g127) & (g147) & (!g569) & (g570) & (!g592) & (!g604)) + ((!g127) & (g147) & (!g569) & (g570) & (g592) & (!g604)) + ((!g127) & (g147) & (g569) & (!g570) & (!g592) & (!g604)) + ((!g127) & (g147) & (g569) & (!g570) & (!g592) & (g604)) + ((!g127) & (g147) & (g569) & (!g570) & (g592) & (g604)) + ((!g127) & (g147) & (g569) & (g570) & (!g592) & (g604)) + ((!g127) & (g147) & (g569) & (g570) & (g592) & (g604)) + ((g127) & (!g147) & (!g569) & (!g570) & (!g592) & (!g604)) + ((g127) & (!g147) & (!g569) & (!g570) & (g592) & (!g604)) + ((g127) & (!g147) & (!g569) & (g570) & (!g592) & (!g604)) + ((g127) & (!g147) & (g569) & (!g570) & (!g592) & (g604)) + ((g127) & (!g147) & (g569) & (!g570) & (g592) & (g604)) + ((g127) & (!g147) & (g569) & (g570) & (!g592) & (g604)) + ((g127) & (!g147) & (g569) & (g570) & (g592) & (!g604)) + ((g127) & (!g147) & (g569) & (g570) & (g592) & (g604)) + ((g127) & (g147) & (!g569) & (!g570) & (!g592) & (!g604)) + ((g127) & (g147) & (g569) & (!g570) & (!g592) & (g604)) + ((g127) & (g147) & (g569) & (!g570) & (g592) & (!g604)) + ((g127) & (g147) & (g569) & (!g570) & (g592) & (g604)) + ((g127) & (g147) & (g569) & (g570) & (!g592) & (!g604)) + ((g127) & (g147) & (g569) & (g570) & (!g592) & (g604)) + ((g127) & (g147) & (g569) & (g570) & (g592) & (!g604)) + ((g127) & (g147) & (g569) & (g570) & (g592) & (g604)));
	assign g616 = (((!g147) & (!g570) & (g592) & (!g604)) + ((!g147) & (g570) & (!g592) & (!g604)) + ((!g147) & (g570) & (!g592) & (g604)) + ((!g147) & (g570) & (g592) & (g604)) + ((g147) & (!g570) & (!g592) & (!g604)) + ((g147) & (g570) & (!g592) & (g604)) + ((g147) & (g570) & (g592) & (!g604)) + ((g147) & (g570) & (g592) & (g604)));
	assign g617 = (((!g174) & (!g198) & (!g572) & (g573) & (g591) & (!g604)) + ((!g174) & (!g198) & (g572) & (!g573) & (!g591) & (!g604)) + ((!g174) & (!g198) & (g572) & (!g573) & (!g591) & (g604)) + ((!g174) & (!g198) & (g572) & (!g573) & (g591) & (!g604)) + ((!g174) & (!g198) & (g572) & (!g573) & (g591) & (g604)) + ((!g174) & (!g198) & (g572) & (g573) & (!g591) & (!g604)) + ((!g174) & (!g198) & (g572) & (g573) & (!g591) & (g604)) + ((!g174) & (!g198) & (g572) & (g573) & (g591) & (g604)) + ((!g174) & (g198) & (!g572) & (!g573) & (g591) & (!g604)) + ((!g174) & (g198) & (!g572) & (g573) & (!g591) & (!g604)) + ((!g174) & (g198) & (!g572) & (g573) & (g591) & (!g604)) + ((!g174) & (g198) & (g572) & (!g573) & (!g591) & (!g604)) + ((!g174) & (g198) & (g572) & (!g573) & (!g591) & (g604)) + ((!g174) & (g198) & (g572) & (!g573) & (g591) & (g604)) + ((!g174) & (g198) & (g572) & (g573) & (!g591) & (g604)) + ((!g174) & (g198) & (g572) & (g573) & (g591) & (g604)) + ((g174) & (!g198) & (!g572) & (!g573) & (!g591) & (!g604)) + ((g174) & (!g198) & (!g572) & (!g573) & (g591) & (!g604)) + ((g174) & (!g198) & (!g572) & (g573) & (!g591) & (!g604)) + ((g174) & (!g198) & (g572) & (!g573) & (!g591) & (g604)) + ((g174) & (!g198) & (g572) & (!g573) & (g591) & (g604)) + ((g174) & (!g198) & (g572) & (g573) & (!g591) & (g604)) + ((g174) & (!g198) & (g572) & (g573) & (g591) & (!g604)) + ((g174) & (!g198) & (g572) & (g573) & (g591) & (g604)) + ((g174) & (g198) & (!g572) & (!g573) & (!g591) & (!g604)) + ((g174) & (g198) & (g572) & (!g573) & (!g591) & (g604)) + ((g174) & (g198) & (g572) & (!g573) & (g591) & (!g604)) + ((g174) & (g198) & (g572) & (!g573) & (g591) & (g604)) + ((g174) & (g198) & (g572) & (g573) & (!g591) & (!g604)) + ((g174) & (g198) & (g572) & (g573) & (!g591) & (g604)) + ((g174) & (g198) & (g572) & (g573) & (g591) & (!g604)) + ((g174) & (g198) & (g572) & (g573) & (g591) & (g604)));
	assign g618 = (((!g198) & (!g573) & (g591) & (!g604)) + ((!g198) & (g573) & (!g591) & (!g604)) + ((!g198) & (g573) & (!g591) & (g604)) + ((!g198) & (g573) & (g591) & (g604)) + ((g198) & (!g573) & (!g591) & (!g604)) + ((g198) & (g573) & (!g591) & (g604)) + ((g198) & (g573) & (g591) & (!g604)) + ((g198) & (g573) & (g591) & (g604)));
	assign g619 = (((!g229) & (!g255) & (!g575) & (g576) & (g590) & (!g604)) + ((!g229) & (!g255) & (g575) & (!g576) & (!g590) & (!g604)) + ((!g229) & (!g255) & (g575) & (!g576) & (!g590) & (g604)) + ((!g229) & (!g255) & (g575) & (!g576) & (g590) & (!g604)) + ((!g229) & (!g255) & (g575) & (!g576) & (g590) & (g604)) + ((!g229) & (!g255) & (g575) & (g576) & (!g590) & (!g604)) + ((!g229) & (!g255) & (g575) & (g576) & (!g590) & (g604)) + ((!g229) & (!g255) & (g575) & (g576) & (g590) & (g604)) + ((!g229) & (g255) & (!g575) & (!g576) & (g590) & (!g604)) + ((!g229) & (g255) & (!g575) & (g576) & (!g590) & (!g604)) + ((!g229) & (g255) & (!g575) & (g576) & (g590) & (!g604)) + ((!g229) & (g255) & (g575) & (!g576) & (!g590) & (!g604)) + ((!g229) & (g255) & (g575) & (!g576) & (!g590) & (g604)) + ((!g229) & (g255) & (g575) & (!g576) & (g590) & (g604)) + ((!g229) & (g255) & (g575) & (g576) & (!g590) & (g604)) + ((!g229) & (g255) & (g575) & (g576) & (g590) & (g604)) + ((g229) & (!g255) & (!g575) & (!g576) & (!g590) & (!g604)) + ((g229) & (!g255) & (!g575) & (!g576) & (g590) & (!g604)) + ((g229) & (!g255) & (!g575) & (g576) & (!g590) & (!g604)) + ((g229) & (!g255) & (g575) & (!g576) & (!g590) & (g604)) + ((g229) & (!g255) & (g575) & (!g576) & (g590) & (g604)) + ((g229) & (!g255) & (g575) & (g576) & (!g590) & (g604)) + ((g229) & (!g255) & (g575) & (g576) & (g590) & (!g604)) + ((g229) & (!g255) & (g575) & (g576) & (g590) & (g604)) + ((g229) & (g255) & (!g575) & (!g576) & (!g590) & (!g604)) + ((g229) & (g255) & (g575) & (!g576) & (!g590) & (g604)) + ((g229) & (g255) & (g575) & (!g576) & (g590) & (!g604)) + ((g229) & (g255) & (g575) & (!g576) & (g590) & (g604)) + ((g229) & (g255) & (g575) & (g576) & (!g590) & (!g604)) + ((g229) & (g255) & (g575) & (g576) & (!g590) & (g604)) + ((g229) & (g255) & (g575) & (g576) & (g590) & (!g604)) + ((g229) & (g255) & (g575) & (g576) & (g590) & (g604)));
	assign g620 = (((!g255) & (!g576) & (g590) & (!g604)) + ((!g255) & (g576) & (!g590) & (!g604)) + ((!g255) & (g576) & (!g590) & (g604)) + ((!g255) & (g576) & (g590) & (g604)) + ((g255) & (!g576) & (!g590) & (!g604)) + ((g255) & (g576) & (!g590) & (g604)) + ((g255) & (g576) & (g590) & (!g604)) + ((g255) & (g576) & (g590) & (g604)));
	assign g621 = (((!g290) & (!g319) & (!g578) & (g579) & (g589) & (!g604)) + ((!g290) & (!g319) & (g578) & (!g579) & (!g589) & (!g604)) + ((!g290) & (!g319) & (g578) & (!g579) & (!g589) & (g604)) + ((!g290) & (!g319) & (g578) & (!g579) & (g589) & (!g604)) + ((!g290) & (!g319) & (g578) & (!g579) & (g589) & (g604)) + ((!g290) & (!g319) & (g578) & (g579) & (!g589) & (!g604)) + ((!g290) & (!g319) & (g578) & (g579) & (!g589) & (g604)) + ((!g290) & (!g319) & (g578) & (g579) & (g589) & (g604)) + ((!g290) & (g319) & (!g578) & (!g579) & (g589) & (!g604)) + ((!g290) & (g319) & (!g578) & (g579) & (!g589) & (!g604)) + ((!g290) & (g319) & (!g578) & (g579) & (g589) & (!g604)) + ((!g290) & (g319) & (g578) & (!g579) & (!g589) & (!g604)) + ((!g290) & (g319) & (g578) & (!g579) & (!g589) & (g604)) + ((!g290) & (g319) & (g578) & (!g579) & (g589) & (g604)) + ((!g290) & (g319) & (g578) & (g579) & (!g589) & (g604)) + ((!g290) & (g319) & (g578) & (g579) & (g589) & (g604)) + ((g290) & (!g319) & (!g578) & (!g579) & (!g589) & (!g604)) + ((g290) & (!g319) & (!g578) & (!g579) & (g589) & (!g604)) + ((g290) & (!g319) & (!g578) & (g579) & (!g589) & (!g604)) + ((g290) & (!g319) & (g578) & (!g579) & (!g589) & (g604)) + ((g290) & (!g319) & (g578) & (!g579) & (g589) & (g604)) + ((g290) & (!g319) & (g578) & (g579) & (!g589) & (g604)) + ((g290) & (!g319) & (g578) & (g579) & (g589) & (!g604)) + ((g290) & (!g319) & (g578) & (g579) & (g589) & (g604)) + ((g290) & (g319) & (!g578) & (!g579) & (!g589) & (!g604)) + ((g290) & (g319) & (g578) & (!g579) & (!g589) & (g604)) + ((g290) & (g319) & (g578) & (!g579) & (g589) & (!g604)) + ((g290) & (g319) & (g578) & (!g579) & (g589) & (g604)) + ((g290) & (g319) & (g578) & (g579) & (!g589) & (!g604)) + ((g290) & (g319) & (g578) & (g579) & (!g589) & (g604)) + ((g290) & (g319) & (g578) & (g579) & (g589) & (!g604)) + ((g290) & (g319) & (g578) & (g579) & (g589) & (g604)));
	assign g622 = (((!g319) & (!g579) & (g589) & (!g604)) + ((!g319) & (g579) & (!g589) & (!g604)) + ((!g319) & (g579) & (!g589) & (g604)) + ((!g319) & (g579) & (g589) & (g604)) + ((g319) & (!g579) & (!g589) & (!g604)) + ((g319) & (g579) & (!g589) & (g604)) + ((g319) & (g579) & (g589) & (!g604)) + ((g319) & (g579) & (g589) & (g604)));
	assign g623 = (((!g358) & (!g390) & (!g581) & (g582) & (g588) & (!g604)) + ((!g358) & (!g390) & (g581) & (!g582) & (!g588) & (!g604)) + ((!g358) & (!g390) & (g581) & (!g582) & (!g588) & (g604)) + ((!g358) & (!g390) & (g581) & (!g582) & (g588) & (!g604)) + ((!g358) & (!g390) & (g581) & (!g582) & (g588) & (g604)) + ((!g358) & (!g390) & (g581) & (g582) & (!g588) & (!g604)) + ((!g358) & (!g390) & (g581) & (g582) & (!g588) & (g604)) + ((!g358) & (!g390) & (g581) & (g582) & (g588) & (g604)) + ((!g358) & (g390) & (!g581) & (!g582) & (g588) & (!g604)) + ((!g358) & (g390) & (!g581) & (g582) & (!g588) & (!g604)) + ((!g358) & (g390) & (!g581) & (g582) & (g588) & (!g604)) + ((!g358) & (g390) & (g581) & (!g582) & (!g588) & (!g604)) + ((!g358) & (g390) & (g581) & (!g582) & (!g588) & (g604)) + ((!g358) & (g390) & (g581) & (!g582) & (g588) & (g604)) + ((!g358) & (g390) & (g581) & (g582) & (!g588) & (g604)) + ((!g358) & (g390) & (g581) & (g582) & (g588) & (g604)) + ((g358) & (!g390) & (!g581) & (!g582) & (!g588) & (!g604)) + ((g358) & (!g390) & (!g581) & (!g582) & (g588) & (!g604)) + ((g358) & (!g390) & (!g581) & (g582) & (!g588) & (!g604)) + ((g358) & (!g390) & (g581) & (!g582) & (!g588) & (g604)) + ((g358) & (!g390) & (g581) & (!g582) & (g588) & (g604)) + ((g358) & (!g390) & (g581) & (g582) & (!g588) & (g604)) + ((g358) & (!g390) & (g581) & (g582) & (g588) & (!g604)) + ((g358) & (!g390) & (g581) & (g582) & (g588) & (g604)) + ((g358) & (g390) & (!g581) & (!g582) & (!g588) & (!g604)) + ((g358) & (g390) & (g581) & (!g582) & (!g588) & (g604)) + ((g358) & (g390) & (g581) & (!g582) & (g588) & (!g604)) + ((g358) & (g390) & (g581) & (!g582) & (g588) & (g604)) + ((g358) & (g390) & (g581) & (g582) & (!g588) & (!g604)) + ((g358) & (g390) & (g581) & (g582) & (!g588) & (g604)) + ((g358) & (g390) & (g581) & (g582) & (g588) & (!g604)) + ((g358) & (g390) & (g581) & (g582) & (g588) & (g604)));
	assign g624 = (((!g390) & (!g582) & (g588) & (!g604)) + ((!g390) & (g582) & (!g588) & (!g604)) + ((!g390) & (g582) & (!g588) & (g604)) + ((!g390) & (g582) & (g588) & (g604)) + ((g390) & (!g582) & (!g588) & (!g604)) + ((g390) & (g582) & (!g588) & (g604)) + ((g390) & (g582) & (g588) & (!g604)) + ((g390) & (g582) & (g588) & (g604)));
	assign g625 = (((!g433) & (!g468) & (!g584) & (g585) & (g587) & (!g604)) + ((!g433) & (!g468) & (g584) & (!g585) & (!g587) & (!g604)) + ((!g433) & (!g468) & (g584) & (!g585) & (!g587) & (g604)) + ((!g433) & (!g468) & (g584) & (!g585) & (g587) & (!g604)) + ((!g433) & (!g468) & (g584) & (!g585) & (g587) & (g604)) + ((!g433) & (!g468) & (g584) & (g585) & (!g587) & (!g604)) + ((!g433) & (!g468) & (g584) & (g585) & (!g587) & (g604)) + ((!g433) & (!g468) & (g584) & (g585) & (g587) & (g604)) + ((!g433) & (g468) & (!g584) & (!g585) & (g587) & (!g604)) + ((!g433) & (g468) & (!g584) & (g585) & (!g587) & (!g604)) + ((!g433) & (g468) & (!g584) & (g585) & (g587) & (!g604)) + ((!g433) & (g468) & (g584) & (!g585) & (!g587) & (!g604)) + ((!g433) & (g468) & (g584) & (!g585) & (!g587) & (g604)) + ((!g433) & (g468) & (g584) & (!g585) & (g587) & (g604)) + ((!g433) & (g468) & (g584) & (g585) & (!g587) & (g604)) + ((!g433) & (g468) & (g584) & (g585) & (g587) & (g604)) + ((g433) & (!g468) & (!g584) & (!g585) & (!g587) & (!g604)) + ((g433) & (!g468) & (!g584) & (!g585) & (g587) & (!g604)) + ((g433) & (!g468) & (!g584) & (g585) & (!g587) & (!g604)) + ((g433) & (!g468) & (g584) & (!g585) & (!g587) & (g604)) + ((g433) & (!g468) & (g584) & (!g585) & (g587) & (g604)) + ((g433) & (!g468) & (g584) & (g585) & (!g587) & (g604)) + ((g433) & (!g468) & (g584) & (g585) & (g587) & (!g604)) + ((g433) & (!g468) & (g584) & (g585) & (g587) & (g604)) + ((g433) & (g468) & (!g584) & (!g585) & (!g587) & (!g604)) + ((g433) & (g468) & (g584) & (!g585) & (!g587) & (g604)) + ((g433) & (g468) & (g584) & (!g585) & (g587) & (!g604)) + ((g433) & (g468) & (g584) & (!g585) & (g587) & (g604)) + ((g433) & (g468) & (g584) & (g585) & (!g587) & (!g604)) + ((g433) & (g468) & (g584) & (g585) & (!g587) & (g604)) + ((g433) & (g468) & (g584) & (g585) & (g587) & (!g604)) + ((g433) & (g468) & (g584) & (g585) & (g587) & (g604)));
	assign g626 = (((!g468) & (!g585) & (g587) & (!g604)) + ((!g468) & (g585) & (!g587) & (!g604)) + ((!g468) & (g585) & (!g587) & (g604)) + ((!g468) & (g585) & (g587) & (g604)) + ((g468) & (!g585) & (!g587) & (!g604)) + ((g468) & (g585) & (!g587) & (g604)) + ((g468) & (g585) & (g587) & (!g604)) + ((g468) & (g585) & (g587) & (g604)));
	assign g627 = (((!g515) & (!ax78x) & (!ax79x) & (!g553) & (!g586) & (g604)) + ((!g515) & (!ax78x) & (!ax79x) & (!g553) & (g586) & (!g604)) + ((!g515) & (!ax78x) & (!ax79x) & (!g553) & (g586) & (g604)) + ((!g515) & (!ax78x) & (!ax79x) & (g553) & (!g586) & (!g604)) + ((!g515) & (!ax78x) & (ax79x) & (!g553) & (!g586) & (!g604)) + ((!g515) & (!ax78x) & (ax79x) & (g553) & (!g586) & (g604)) + ((!g515) & (!ax78x) & (ax79x) & (g553) & (g586) & (!g604)) + ((!g515) & (!ax78x) & (ax79x) & (g553) & (g586) & (g604)) + ((!g515) & (ax78x) & (!ax79x) & (g553) & (!g586) & (!g604)) + ((!g515) & (ax78x) & (!ax79x) & (g553) & (g586) & (!g604)) + ((!g515) & (ax78x) & (ax79x) & (!g553) & (!g586) & (!g604)) + ((!g515) & (ax78x) & (ax79x) & (!g553) & (!g586) & (g604)) + ((!g515) & (ax78x) & (ax79x) & (!g553) & (g586) & (!g604)) + ((!g515) & (ax78x) & (ax79x) & (!g553) & (g586) & (g604)) + ((!g515) & (ax78x) & (ax79x) & (g553) & (!g586) & (g604)) + ((!g515) & (ax78x) & (ax79x) & (g553) & (g586) & (g604)) + ((g515) & (!ax78x) & (!ax79x) & (!g553) & (!g586) & (!g604)) + ((g515) & (!ax78x) & (!ax79x) & (!g553) & (!g586) & (g604)) + ((g515) & (!ax78x) & (!ax79x) & (!g553) & (g586) & (g604)) + ((g515) & (!ax78x) & (!ax79x) & (g553) & (g586) & (!g604)) + ((g515) & (!ax78x) & (ax79x) & (!g553) & (g586) & (!g604)) + ((g515) & (!ax78x) & (ax79x) & (g553) & (!g586) & (!g604)) + ((g515) & (!ax78x) & (ax79x) & (g553) & (!g586) & (g604)) + ((g515) & (!ax78x) & (ax79x) & (g553) & (g586) & (g604)) + ((g515) & (ax78x) & (!ax79x) & (!g553) & (!g586) & (!g604)) + ((g515) & (ax78x) & (!ax79x) & (!g553) & (g586) & (!g604)) + ((g515) & (ax78x) & (ax79x) & (!g553) & (!g586) & (g604)) + ((g515) & (ax78x) & (ax79x) & (!g553) & (g586) & (g604)) + ((g515) & (ax78x) & (ax79x) & (g553) & (!g586) & (!g604)) + ((g515) & (ax78x) & (ax79x) & (g553) & (!g586) & (g604)) + ((g515) & (ax78x) & (ax79x) & (g553) & (g586) & (!g604)) + ((g515) & (ax78x) & (ax79x) & (g553) & (g586) & (g604)));
	assign g628 = (((!ax78x) & (!g553) & (!g586) & (g604)) + ((!ax78x) & (!g553) & (g586) & (!g604)) + ((!ax78x) & (!g553) & (g586) & (g604)) + ((!ax78x) & (g553) & (g586) & (!g604)) + ((ax78x) & (!g553) & (!g586) & (!g604)) + ((ax78x) & (g553) & (!g586) & (!g604)) + ((ax78x) & (g553) & (!g586) & (g604)) + ((ax78x) & (g553) & (g586) & (g604)));
	assign g629 = (((!ax74x) & (!ax75x)));
	assign g630 = (((!g553) & (!ax76x) & (!ax77x) & (!g604) & (!g629)) + ((!g553) & (!ax76x) & (ax77x) & (g604) & (!g629)) + ((!g553) & (ax76x) & (ax77x) & (g604) & (!g629)) + ((!g553) & (ax76x) & (ax77x) & (g604) & (g629)) + ((g553) & (!ax76x) & (!ax77x) & (!g604) & (!g629)) + ((g553) & (!ax76x) & (!ax77x) & (!g604) & (g629)) + ((g553) & (!ax76x) & (!ax77x) & (g604) & (!g629)) + ((g553) & (!ax76x) & (ax77x) & (!g604) & (!g629)) + ((g553) & (!ax76x) & (ax77x) & (g604) & (!g629)) + ((g553) & (!ax76x) & (ax77x) & (g604) & (g629)) + ((g553) & (ax76x) & (!ax77x) & (g604) & (!g629)) + ((g553) & (ax76x) & (!ax77x) & (g604) & (g629)) + ((g553) & (ax76x) & (ax77x) & (!g604) & (!g629)) + ((g553) & (ax76x) & (ax77x) & (!g604) & (g629)) + ((g553) & (ax76x) & (ax77x) & (g604) & (!g629)) + ((g553) & (ax76x) & (ax77x) & (g604) & (g629)));
	assign g631 = (((!g468) & (!g515) & (g627) & (g628) & (g630)) + ((!g468) & (g515) & (g627) & (!g628) & (g630)) + ((!g468) & (g515) & (g627) & (g628) & (!g630)) + ((!g468) & (g515) & (g627) & (g628) & (g630)) + ((g468) & (!g515) & (!g627) & (g628) & (g630)) + ((g468) & (!g515) & (g627) & (!g628) & (!g630)) + ((g468) & (!g515) & (g627) & (!g628) & (g630)) + ((g468) & (!g515) & (g627) & (g628) & (!g630)) + ((g468) & (!g515) & (g627) & (g628) & (g630)) + ((g468) & (g515) & (!g627) & (!g628) & (g630)) + ((g468) & (g515) & (!g627) & (g628) & (!g630)) + ((g468) & (g515) & (!g627) & (g628) & (g630)) + ((g468) & (g515) & (g627) & (!g628) & (!g630)) + ((g468) & (g515) & (g627) & (!g628) & (g630)) + ((g468) & (g515) & (g627) & (g628) & (!g630)) + ((g468) & (g515) & (g627) & (g628) & (g630)));
	assign g632 = (((!g390) & (!g433) & (g625) & (g626) & (g631)) + ((!g390) & (g433) & (g625) & (!g626) & (g631)) + ((!g390) & (g433) & (g625) & (g626) & (!g631)) + ((!g390) & (g433) & (g625) & (g626) & (g631)) + ((g390) & (!g433) & (!g625) & (g626) & (g631)) + ((g390) & (!g433) & (g625) & (!g626) & (!g631)) + ((g390) & (!g433) & (g625) & (!g626) & (g631)) + ((g390) & (!g433) & (g625) & (g626) & (!g631)) + ((g390) & (!g433) & (g625) & (g626) & (g631)) + ((g390) & (g433) & (!g625) & (!g626) & (g631)) + ((g390) & (g433) & (!g625) & (g626) & (!g631)) + ((g390) & (g433) & (!g625) & (g626) & (g631)) + ((g390) & (g433) & (g625) & (!g626) & (!g631)) + ((g390) & (g433) & (g625) & (!g626) & (g631)) + ((g390) & (g433) & (g625) & (g626) & (!g631)) + ((g390) & (g433) & (g625) & (g626) & (g631)));
	assign g633 = (((!g319) & (!g358) & (g623) & (g624) & (g632)) + ((!g319) & (g358) & (g623) & (!g624) & (g632)) + ((!g319) & (g358) & (g623) & (g624) & (!g632)) + ((!g319) & (g358) & (g623) & (g624) & (g632)) + ((g319) & (!g358) & (!g623) & (g624) & (g632)) + ((g319) & (!g358) & (g623) & (!g624) & (!g632)) + ((g319) & (!g358) & (g623) & (!g624) & (g632)) + ((g319) & (!g358) & (g623) & (g624) & (!g632)) + ((g319) & (!g358) & (g623) & (g624) & (g632)) + ((g319) & (g358) & (!g623) & (!g624) & (g632)) + ((g319) & (g358) & (!g623) & (g624) & (!g632)) + ((g319) & (g358) & (!g623) & (g624) & (g632)) + ((g319) & (g358) & (g623) & (!g624) & (!g632)) + ((g319) & (g358) & (g623) & (!g624) & (g632)) + ((g319) & (g358) & (g623) & (g624) & (!g632)) + ((g319) & (g358) & (g623) & (g624) & (g632)));
	assign g634 = (((!g255) & (!g290) & (g621) & (g622) & (g633)) + ((!g255) & (g290) & (g621) & (!g622) & (g633)) + ((!g255) & (g290) & (g621) & (g622) & (!g633)) + ((!g255) & (g290) & (g621) & (g622) & (g633)) + ((g255) & (!g290) & (!g621) & (g622) & (g633)) + ((g255) & (!g290) & (g621) & (!g622) & (!g633)) + ((g255) & (!g290) & (g621) & (!g622) & (g633)) + ((g255) & (!g290) & (g621) & (g622) & (!g633)) + ((g255) & (!g290) & (g621) & (g622) & (g633)) + ((g255) & (g290) & (!g621) & (!g622) & (g633)) + ((g255) & (g290) & (!g621) & (g622) & (!g633)) + ((g255) & (g290) & (!g621) & (g622) & (g633)) + ((g255) & (g290) & (g621) & (!g622) & (!g633)) + ((g255) & (g290) & (g621) & (!g622) & (g633)) + ((g255) & (g290) & (g621) & (g622) & (!g633)) + ((g255) & (g290) & (g621) & (g622) & (g633)));
	assign g635 = (((!g198) & (!g229) & (g619) & (g620) & (g634)) + ((!g198) & (g229) & (g619) & (!g620) & (g634)) + ((!g198) & (g229) & (g619) & (g620) & (!g634)) + ((!g198) & (g229) & (g619) & (g620) & (g634)) + ((g198) & (!g229) & (!g619) & (g620) & (g634)) + ((g198) & (!g229) & (g619) & (!g620) & (!g634)) + ((g198) & (!g229) & (g619) & (!g620) & (g634)) + ((g198) & (!g229) & (g619) & (g620) & (!g634)) + ((g198) & (!g229) & (g619) & (g620) & (g634)) + ((g198) & (g229) & (!g619) & (!g620) & (g634)) + ((g198) & (g229) & (!g619) & (g620) & (!g634)) + ((g198) & (g229) & (!g619) & (g620) & (g634)) + ((g198) & (g229) & (g619) & (!g620) & (!g634)) + ((g198) & (g229) & (g619) & (!g620) & (g634)) + ((g198) & (g229) & (g619) & (g620) & (!g634)) + ((g198) & (g229) & (g619) & (g620) & (g634)));
	assign g636 = (((!g147) & (!g174) & (g617) & (g618) & (g635)) + ((!g147) & (g174) & (g617) & (!g618) & (g635)) + ((!g147) & (g174) & (g617) & (g618) & (!g635)) + ((!g147) & (g174) & (g617) & (g618) & (g635)) + ((g147) & (!g174) & (!g617) & (g618) & (g635)) + ((g147) & (!g174) & (g617) & (!g618) & (!g635)) + ((g147) & (!g174) & (g617) & (!g618) & (g635)) + ((g147) & (!g174) & (g617) & (g618) & (!g635)) + ((g147) & (!g174) & (g617) & (g618) & (g635)) + ((g147) & (g174) & (!g617) & (!g618) & (g635)) + ((g147) & (g174) & (!g617) & (g618) & (!g635)) + ((g147) & (g174) & (!g617) & (g618) & (g635)) + ((g147) & (g174) & (g617) & (!g618) & (!g635)) + ((g147) & (g174) & (g617) & (!g618) & (g635)) + ((g147) & (g174) & (g617) & (g618) & (!g635)) + ((g147) & (g174) & (g617) & (g618) & (g635)));
	assign g637 = (((!g104) & (!g127) & (g615) & (g616) & (g636)) + ((!g104) & (g127) & (g615) & (!g616) & (g636)) + ((!g104) & (g127) & (g615) & (g616) & (!g636)) + ((!g104) & (g127) & (g615) & (g616) & (g636)) + ((g104) & (!g127) & (!g615) & (g616) & (g636)) + ((g104) & (!g127) & (g615) & (!g616) & (!g636)) + ((g104) & (!g127) & (g615) & (!g616) & (g636)) + ((g104) & (!g127) & (g615) & (g616) & (!g636)) + ((g104) & (!g127) & (g615) & (g616) & (g636)) + ((g104) & (g127) & (!g615) & (!g616) & (g636)) + ((g104) & (g127) & (!g615) & (g616) & (!g636)) + ((g104) & (g127) & (!g615) & (g616) & (g636)) + ((g104) & (g127) & (g615) & (!g616) & (!g636)) + ((g104) & (g127) & (g615) & (!g616) & (g636)) + ((g104) & (g127) & (g615) & (g616) & (!g636)) + ((g104) & (g127) & (g615) & (g616) & (g636)));
	assign g638 = (((!g68) & (!g87) & (g613) & (g614) & (g637)) + ((!g68) & (g87) & (g613) & (!g614) & (g637)) + ((!g68) & (g87) & (g613) & (g614) & (!g637)) + ((!g68) & (g87) & (g613) & (g614) & (g637)) + ((g68) & (!g87) & (!g613) & (g614) & (g637)) + ((g68) & (!g87) & (g613) & (!g614) & (!g637)) + ((g68) & (!g87) & (g613) & (!g614) & (g637)) + ((g68) & (!g87) & (g613) & (g614) & (!g637)) + ((g68) & (!g87) & (g613) & (g614) & (g637)) + ((g68) & (g87) & (!g613) & (!g614) & (g637)) + ((g68) & (g87) & (!g613) & (g614) & (!g637)) + ((g68) & (g87) & (!g613) & (g614) & (g637)) + ((g68) & (g87) & (g613) & (!g614) & (!g637)) + ((g68) & (g87) & (g613) & (!g614) & (g637)) + ((g68) & (g87) & (g613) & (g614) & (!g637)) + ((g68) & (g87) & (g613) & (g614) & (g637)));
	assign g639 = (((!g39) & (!g54) & (g611) & (g612) & (g638)) + ((!g39) & (g54) & (g611) & (!g612) & (g638)) + ((!g39) & (g54) & (g611) & (g612) & (!g638)) + ((!g39) & (g54) & (g611) & (g612) & (g638)) + ((g39) & (!g54) & (!g611) & (g612) & (g638)) + ((g39) & (!g54) & (g611) & (!g612) & (!g638)) + ((g39) & (!g54) & (g611) & (!g612) & (g638)) + ((g39) & (!g54) & (g611) & (g612) & (!g638)) + ((g39) & (!g54) & (g611) & (g612) & (g638)) + ((g39) & (g54) & (!g611) & (!g612) & (g638)) + ((g39) & (g54) & (!g611) & (g612) & (!g638)) + ((g39) & (g54) & (!g611) & (g612) & (g638)) + ((g39) & (g54) & (g611) & (!g612) & (!g638)) + ((g39) & (g54) & (g611) & (!g612) & (g638)) + ((g39) & (g54) & (g611) & (g612) & (!g638)) + ((g39) & (g54) & (g611) & (g612) & (g638)));
	assign g640 = (((!g18) & (!g27) & (g609) & (g610) & (g639)) + ((!g18) & (g27) & (g609) & (!g610) & (g639)) + ((!g18) & (g27) & (g609) & (g610) & (!g639)) + ((!g18) & (g27) & (g609) & (g610) & (g639)) + ((g18) & (!g27) & (!g609) & (g610) & (g639)) + ((g18) & (!g27) & (g609) & (!g610) & (!g639)) + ((g18) & (!g27) & (g609) & (!g610) & (g639)) + ((g18) & (!g27) & (g609) & (g610) & (!g639)) + ((g18) & (!g27) & (g609) & (g610) & (g639)) + ((g18) & (g27) & (!g609) & (!g610) & (g639)) + ((g18) & (g27) & (!g609) & (g610) & (!g639)) + ((g18) & (g27) & (!g609) & (g610) & (g639)) + ((g18) & (g27) & (g609) & (!g610) & (!g639)) + ((g18) & (g27) & (g609) & (!g610) & (g639)) + ((g18) & (g27) & (g609) & (g610) & (!g639)) + ((g18) & (g27) & (g609) & (g610) & (g639)));
	assign g641 = (((!g2) & (!g8) & (g607) & (g608) & (g640)) + ((!g2) & (g8) & (g607) & (!g608) & (g640)) + ((!g2) & (g8) & (g607) & (g608) & (!g640)) + ((!g2) & (g8) & (g607) & (g608) & (g640)) + ((g2) & (!g8) & (!g607) & (g608) & (g640)) + ((g2) & (!g8) & (g607) & (!g608) & (!g640)) + ((g2) & (!g8) & (g607) & (!g608) & (g640)) + ((g2) & (!g8) & (g607) & (g608) & (!g640)) + ((g2) & (!g8) & (g607) & (g608) & (g640)) + ((g2) & (g8) & (!g607) & (!g608) & (g640)) + ((g2) & (g8) & (!g607) & (g608) & (!g640)) + ((g2) & (g8) & (!g607) & (g608) & (g640)) + ((g2) & (g8) & (g607) & (!g608) & (!g640)) + ((g2) & (g8) & (g607) & (!g608) & (g640)) + ((g2) & (g8) & (g607) & (g608) & (!g640)) + ((g2) & (g8) & (g607) & (g608) & (g640)));
	assign g642 = (((!g2) & (!g555) & (g597) & (!g604)) + ((!g2) & (g555) & (!g597) & (!g604)) + ((!g2) & (g555) & (!g597) & (g604)) + ((!g2) & (g555) & (g597) & (g604)) + ((g2) & (!g555) & (!g597) & (!g604)) + ((g2) & (g555) & (!g597) & (g604)) + ((g2) & (g555) & (g597) & (!g604)) + ((g2) & (g555) & (g597) & (g604)));
	assign g643 = (((!g1) & (!g554) & (!g600) & (!g602) & (g603)) + ((!g1) & (!g554) & (!g600) & (g602) & (!g603)) + ((!g1) & (!g554) & (!g600) & (g602) & (g603)) + ((!g1) & (g554) & (g600) & (!g602) & (!g603)) + ((!g1) & (g554) & (g600) & (!g602) & (g603)) + ((!g1) & (g554) & (g600) & (g602) & (!g603)) + ((!g1) & (g554) & (g600) & (g602) & (g603)) + ((g1) & (!g554) & (!g600) & (!g602) & (g603)) + ((g1) & (!g554) & (!g600) & (g602) & (g603)) + ((g1) & (g554) & (g600) & (!g602) & (!g603)) + ((g1) & (g554) & (g600) & (!g602) & (g603)) + ((g1) & (g554) & (g600) & (g602) & (!g603)) + ((g1) & (g554) & (g600) & (g602) & (g603)));
	assign g644 = (((!g4) & (!g1) & (!g606) & (!g641) & (!g642) & (!g643)) + ((!g4) & (g1) & (!g606) & (!g641) & (!g642) & (!g643)) + ((!g4) & (g1) & (!g606) & (!g641) & (!g642) & (g643)) + ((!g4) & (g1) & (!g606) & (!g641) & (g642) & (!g643)) + ((!g4) & (g1) & (!g606) & (!g641) & (g642) & (g643)) + ((!g4) & (g1) & (!g606) & (g641) & (!g642) & (!g643)) + ((!g4) & (g1) & (!g606) & (g641) & (!g642) & (g643)) + ((!g4) & (g1) & (!g606) & (g641) & (g642) & (!g643)) + ((!g4) & (g1) & (!g606) & (g641) & (g642) & (g643)) + ((!g4) & (g1) & (g606) & (!g641) & (!g642) & (!g643)) + ((!g4) & (g1) & (g606) & (!g641) & (!g642) & (g643)) + ((g4) & (!g1) & (!g606) & (!g641) & (!g642) & (!g643)) + ((g4) & (!g1) & (!g606) & (!g641) & (g642) & (!g643)) + ((g4) & (!g1) & (!g606) & (g641) & (!g642) & (!g643)) + ((g4) & (g1) & (!g606) & (!g641) & (!g642) & (!g643)) + ((g4) & (g1) & (!g606) & (!g641) & (!g642) & (g643)) + ((g4) & (g1) & (!g606) & (!g641) & (g642) & (!g643)) + ((g4) & (g1) & (!g606) & (!g641) & (g642) & (g643)) + ((g4) & (g1) & (!g606) & (g641) & (!g642) & (!g643)) + ((g4) & (g1) & (!g606) & (g641) & (!g642) & (g643)) + ((g4) & (g1) & (!g606) & (g641) & (g642) & (!g643)) + ((g4) & (g1) & (!g606) & (g641) & (g642) & (g643)) + ((g4) & (g1) & (g606) & (!g641) & (!g642) & (!g643)) + ((g4) & (g1) & (g606) & (!g641) & (!g642) & (g643)) + ((g4) & (g1) & (g606) & (!g641) & (g642) & (!g643)) + ((g4) & (g1) & (g606) & (!g641) & (g642) & (g643)) + ((g4) & (g1) & (g606) & (g641) & (!g642) & (!g643)) + ((g4) & (g1) & (g606) & (g641) & (!g642) & (g643)));
	assign g645 = (((!g605) & (g644)));
	assign g646 = (((!g4) & (!g641) & (!g642) & (!g605) & (!g644)) + ((!g4) & (!g641) & (!g642) & (g605) & (!g644)) + ((!g4) & (!g641) & (!g642) & (g605) & (g644)) + ((!g4) & (!g641) & (g642) & (!g605) & (g644)) + ((!g4) & (g641) & (g642) & (!g605) & (!g644)) + ((!g4) & (g641) & (g642) & (!g605) & (g644)) + ((!g4) & (g641) & (g642) & (g605) & (!g644)) + ((!g4) & (g641) & (g642) & (g605) & (g644)) + ((g4) & (!g641) & (g642) & (!g605) & (!g644)) + ((g4) & (!g641) & (g642) & (!g605) & (g644)) + ((g4) & (!g641) & (g642) & (g605) & (!g644)) + ((g4) & (!g641) & (g642) & (g605) & (g644)) + ((g4) & (g641) & (!g642) & (!g605) & (!g644)) + ((g4) & (g641) & (!g642) & (g605) & (!g644)) + ((g4) & (g641) & (!g642) & (g605) & (g644)) + ((g4) & (g641) & (g642) & (!g605) & (g644)));
	assign g647 = (((!g8) & (!g608) & (g640) & (!g605) & (!g644)) + ((!g8) & (!g608) & (g640) & (g605) & (!g644)) + ((!g8) & (!g608) & (g640) & (g605) & (g644)) + ((!g8) & (g608) & (!g640) & (!g605) & (!g644)) + ((!g8) & (g608) & (!g640) & (!g605) & (g644)) + ((!g8) & (g608) & (!g640) & (g605) & (!g644)) + ((!g8) & (g608) & (!g640) & (g605) & (g644)) + ((!g8) & (g608) & (g640) & (!g605) & (g644)) + ((g8) & (!g608) & (!g640) & (!g605) & (!g644)) + ((g8) & (!g608) & (!g640) & (g605) & (!g644)) + ((g8) & (!g608) & (!g640) & (g605) & (g644)) + ((g8) & (g608) & (!g640) & (!g605) & (g644)) + ((g8) & (g608) & (g640) & (!g605) & (!g644)) + ((g8) & (g608) & (g640) & (!g605) & (g644)) + ((g8) & (g608) & (g640) & (g605) & (!g644)) + ((g8) & (g608) & (g640) & (g605) & (g644)));
	assign g648 = (((!g18) & (!g27) & (g610) & (g639)) + ((!g18) & (g27) & (!g610) & (g639)) + ((!g18) & (g27) & (g610) & (!g639)) + ((!g18) & (g27) & (g610) & (g639)) + ((g18) & (!g27) & (!g610) & (!g639)) + ((g18) & (!g27) & (!g610) & (g639)) + ((g18) & (!g27) & (g610) & (!g639)) + ((g18) & (g27) & (!g610) & (!g639)));
	assign g649 = (((!g609) & (!g605) & (!g644) & (g648)) + ((!g609) & (g605) & (!g644) & (g648)) + ((!g609) & (g605) & (g644) & (g648)) + ((g609) & (!g605) & (!g644) & (!g648)) + ((g609) & (!g605) & (g644) & (!g648)) + ((g609) & (!g605) & (g644) & (g648)) + ((g609) & (g605) & (!g644) & (!g648)) + ((g609) & (g605) & (g644) & (!g648)));
	assign g650 = (((!g27) & (!g610) & (g639) & (!g605) & (!g644)) + ((!g27) & (!g610) & (g639) & (g605) & (!g644)) + ((!g27) & (!g610) & (g639) & (g605) & (g644)) + ((!g27) & (g610) & (!g639) & (!g605) & (!g644)) + ((!g27) & (g610) & (!g639) & (!g605) & (g644)) + ((!g27) & (g610) & (!g639) & (g605) & (!g644)) + ((!g27) & (g610) & (!g639) & (g605) & (g644)) + ((!g27) & (g610) & (g639) & (!g605) & (g644)) + ((g27) & (!g610) & (!g639) & (!g605) & (!g644)) + ((g27) & (!g610) & (!g639) & (g605) & (!g644)) + ((g27) & (!g610) & (!g639) & (g605) & (g644)) + ((g27) & (g610) & (!g639) & (!g605) & (g644)) + ((g27) & (g610) & (g639) & (!g605) & (!g644)) + ((g27) & (g610) & (g639) & (!g605) & (g644)) + ((g27) & (g610) & (g639) & (g605) & (!g644)) + ((g27) & (g610) & (g639) & (g605) & (g644)));
	assign g651 = (((!g39) & (!g54) & (g612) & (g638)) + ((!g39) & (g54) & (!g612) & (g638)) + ((!g39) & (g54) & (g612) & (!g638)) + ((!g39) & (g54) & (g612) & (g638)) + ((g39) & (!g54) & (!g612) & (!g638)) + ((g39) & (!g54) & (!g612) & (g638)) + ((g39) & (!g54) & (g612) & (!g638)) + ((g39) & (g54) & (!g612) & (!g638)));
	assign g652 = (((!g611) & (!g605) & (!g644) & (g651)) + ((!g611) & (g605) & (!g644) & (g651)) + ((!g611) & (g605) & (g644) & (g651)) + ((g611) & (!g605) & (!g644) & (!g651)) + ((g611) & (!g605) & (g644) & (!g651)) + ((g611) & (!g605) & (g644) & (g651)) + ((g611) & (g605) & (!g644) & (!g651)) + ((g611) & (g605) & (g644) & (!g651)));
	assign g653 = (((!g54) & (!g612) & (g638) & (!g605) & (!g644)) + ((!g54) & (!g612) & (g638) & (g605) & (!g644)) + ((!g54) & (!g612) & (g638) & (g605) & (g644)) + ((!g54) & (g612) & (!g638) & (!g605) & (!g644)) + ((!g54) & (g612) & (!g638) & (!g605) & (g644)) + ((!g54) & (g612) & (!g638) & (g605) & (!g644)) + ((!g54) & (g612) & (!g638) & (g605) & (g644)) + ((!g54) & (g612) & (g638) & (!g605) & (g644)) + ((g54) & (!g612) & (!g638) & (!g605) & (!g644)) + ((g54) & (!g612) & (!g638) & (g605) & (!g644)) + ((g54) & (!g612) & (!g638) & (g605) & (g644)) + ((g54) & (g612) & (!g638) & (!g605) & (g644)) + ((g54) & (g612) & (g638) & (!g605) & (!g644)) + ((g54) & (g612) & (g638) & (!g605) & (g644)) + ((g54) & (g612) & (g638) & (g605) & (!g644)) + ((g54) & (g612) & (g638) & (g605) & (g644)));
	assign g654 = (((!g68) & (!g87) & (g614) & (g637)) + ((!g68) & (g87) & (!g614) & (g637)) + ((!g68) & (g87) & (g614) & (!g637)) + ((!g68) & (g87) & (g614) & (g637)) + ((g68) & (!g87) & (!g614) & (!g637)) + ((g68) & (!g87) & (!g614) & (g637)) + ((g68) & (!g87) & (g614) & (!g637)) + ((g68) & (g87) & (!g614) & (!g637)));
	assign g655 = (((!g613) & (!g605) & (!g644) & (g654)) + ((!g613) & (g605) & (!g644) & (g654)) + ((!g613) & (g605) & (g644) & (g654)) + ((g613) & (!g605) & (!g644) & (!g654)) + ((g613) & (!g605) & (g644) & (!g654)) + ((g613) & (!g605) & (g644) & (g654)) + ((g613) & (g605) & (!g644) & (!g654)) + ((g613) & (g605) & (g644) & (!g654)));
	assign g656 = (((!g87) & (!g614) & (g637) & (!g605) & (!g644)) + ((!g87) & (!g614) & (g637) & (g605) & (!g644)) + ((!g87) & (!g614) & (g637) & (g605) & (g644)) + ((!g87) & (g614) & (!g637) & (!g605) & (!g644)) + ((!g87) & (g614) & (!g637) & (!g605) & (g644)) + ((!g87) & (g614) & (!g637) & (g605) & (!g644)) + ((!g87) & (g614) & (!g637) & (g605) & (g644)) + ((!g87) & (g614) & (g637) & (!g605) & (g644)) + ((g87) & (!g614) & (!g637) & (!g605) & (!g644)) + ((g87) & (!g614) & (!g637) & (g605) & (!g644)) + ((g87) & (!g614) & (!g637) & (g605) & (g644)) + ((g87) & (g614) & (!g637) & (!g605) & (g644)) + ((g87) & (g614) & (g637) & (!g605) & (!g644)) + ((g87) & (g614) & (g637) & (!g605) & (g644)) + ((g87) & (g614) & (g637) & (g605) & (!g644)) + ((g87) & (g614) & (g637) & (g605) & (g644)));
	assign g657 = (((!g104) & (!g127) & (g616) & (g636)) + ((!g104) & (g127) & (!g616) & (g636)) + ((!g104) & (g127) & (g616) & (!g636)) + ((!g104) & (g127) & (g616) & (g636)) + ((g104) & (!g127) & (!g616) & (!g636)) + ((g104) & (!g127) & (!g616) & (g636)) + ((g104) & (!g127) & (g616) & (!g636)) + ((g104) & (g127) & (!g616) & (!g636)));
	assign g658 = (((!g615) & (!g605) & (!g644) & (g657)) + ((!g615) & (g605) & (!g644) & (g657)) + ((!g615) & (g605) & (g644) & (g657)) + ((g615) & (!g605) & (!g644) & (!g657)) + ((g615) & (!g605) & (g644) & (!g657)) + ((g615) & (!g605) & (g644) & (g657)) + ((g615) & (g605) & (!g644) & (!g657)) + ((g615) & (g605) & (g644) & (!g657)));
	assign g659 = (((!g127) & (!g616) & (g636) & (!g605) & (!g644)) + ((!g127) & (!g616) & (g636) & (g605) & (!g644)) + ((!g127) & (!g616) & (g636) & (g605) & (g644)) + ((!g127) & (g616) & (!g636) & (!g605) & (!g644)) + ((!g127) & (g616) & (!g636) & (!g605) & (g644)) + ((!g127) & (g616) & (!g636) & (g605) & (!g644)) + ((!g127) & (g616) & (!g636) & (g605) & (g644)) + ((!g127) & (g616) & (g636) & (!g605) & (g644)) + ((g127) & (!g616) & (!g636) & (!g605) & (!g644)) + ((g127) & (!g616) & (!g636) & (g605) & (!g644)) + ((g127) & (!g616) & (!g636) & (g605) & (g644)) + ((g127) & (g616) & (!g636) & (!g605) & (g644)) + ((g127) & (g616) & (g636) & (!g605) & (!g644)) + ((g127) & (g616) & (g636) & (!g605) & (g644)) + ((g127) & (g616) & (g636) & (g605) & (!g644)) + ((g127) & (g616) & (g636) & (g605) & (g644)));
	assign g660 = (((!g147) & (!g174) & (g618) & (g635)) + ((!g147) & (g174) & (!g618) & (g635)) + ((!g147) & (g174) & (g618) & (!g635)) + ((!g147) & (g174) & (g618) & (g635)) + ((g147) & (!g174) & (!g618) & (!g635)) + ((g147) & (!g174) & (!g618) & (g635)) + ((g147) & (!g174) & (g618) & (!g635)) + ((g147) & (g174) & (!g618) & (!g635)));
	assign g661 = (((!g617) & (!g605) & (!g644) & (g660)) + ((!g617) & (g605) & (!g644) & (g660)) + ((!g617) & (g605) & (g644) & (g660)) + ((g617) & (!g605) & (!g644) & (!g660)) + ((g617) & (!g605) & (g644) & (!g660)) + ((g617) & (!g605) & (g644) & (g660)) + ((g617) & (g605) & (!g644) & (!g660)) + ((g617) & (g605) & (g644) & (!g660)));
	assign g662 = (((!g174) & (!g618) & (g635) & (!g605) & (!g644)) + ((!g174) & (!g618) & (g635) & (g605) & (!g644)) + ((!g174) & (!g618) & (g635) & (g605) & (g644)) + ((!g174) & (g618) & (!g635) & (!g605) & (!g644)) + ((!g174) & (g618) & (!g635) & (!g605) & (g644)) + ((!g174) & (g618) & (!g635) & (g605) & (!g644)) + ((!g174) & (g618) & (!g635) & (g605) & (g644)) + ((!g174) & (g618) & (g635) & (!g605) & (g644)) + ((g174) & (!g618) & (!g635) & (!g605) & (!g644)) + ((g174) & (!g618) & (!g635) & (g605) & (!g644)) + ((g174) & (!g618) & (!g635) & (g605) & (g644)) + ((g174) & (g618) & (!g635) & (!g605) & (g644)) + ((g174) & (g618) & (g635) & (!g605) & (!g644)) + ((g174) & (g618) & (g635) & (!g605) & (g644)) + ((g174) & (g618) & (g635) & (g605) & (!g644)) + ((g174) & (g618) & (g635) & (g605) & (g644)));
	assign g663 = (((!g198) & (!g229) & (g620) & (g634)) + ((!g198) & (g229) & (!g620) & (g634)) + ((!g198) & (g229) & (g620) & (!g634)) + ((!g198) & (g229) & (g620) & (g634)) + ((g198) & (!g229) & (!g620) & (!g634)) + ((g198) & (!g229) & (!g620) & (g634)) + ((g198) & (!g229) & (g620) & (!g634)) + ((g198) & (g229) & (!g620) & (!g634)));
	assign g664 = (((!g619) & (!g605) & (!g644) & (g663)) + ((!g619) & (g605) & (!g644) & (g663)) + ((!g619) & (g605) & (g644) & (g663)) + ((g619) & (!g605) & (!g644) & (!g663)) + ((g619) & (!g605) & (g644) & (!g663)) + ((g619) & (!g605) & (g644) & (g663)) + ((g619) & (g605) & (!g644) & (!g663)) + ((g619) & (g605) & (g644) & (!g663)));
	assign g665 = (((!g229) & (!g620) & (g634) & (!g605) & (!g644)) + ((!g229) & (!g620) & (g634) & (g605) & (!g644)) + ((!g229) & (!g620) & (g634) & (g605) & (g644)) + ((!g229) & (g620) & (!g634) & (!g605) & (!g644)) + ((!g229) & (g620) & (!g634) & (!g605) & (g644)) + ((!g229) & (g620) & (!g634) & (g605) & (!g644)) + ((!g229) & (g620) & (!g634) & (g605) & (g644)) + ((!g229) & (g620) & (g634) & (!g605) & (g644)) + ((g229) & (!g620) & (!g634) & (!g605) & (!g644)) + ((g229) & (!g620) & (!g634) & (g605) & (!g644)) + ((g229) & (!g620) & (!g634) & (g605) & (g644)) + ((g229) & (g620) & (!g634) & (!g605) & (g644)) + ((g229) & (g620) & (g634) & (!g605) & (!g644)) + ((g229) & (g620) & (g634) & (!g605) & (g644)) + ((g229) & (g620) & (g634) & (g605) & (!g644)) + ((g229) & (g620) & (g634) & (g605) & (g644)));
	assign g666 = (((!g255) & (!g290) & (g622) & (g633)) + ((!g255) & (g290) & (!g622) & (g633)) + ((!g255) & (g290) & (g622) & (!g633)) + ((!g255) & (g290) & (g622) & (g633)) + ((g255) & (!g290) & (!g622) & (!g633)) + ((g255) & (!g290) & (!g622) & (g633)) + ((g255) & (!g290) & (g622) & (!g633)) + ((g255) & (g290) & (!g622) & (!g633)));
	assign g667 = (((!g621) & (!g605) & (!g644) & (g666)) + ((!g621) & (g605) & (!g644) & (g666)) + ((!g621) & (g605) & (g644) & (g666)) + ((g621) & (!g605) & (!g644) & (!g666)) + ((g621) & (!g605) & (g644) & (!g666)) + ((g621) & (!g605) & (g644) & (g666)) + ((g621) & (g605) & (!g644) & (!g666)) + ((g621) & (g605) & (g644) & (!g666)));
	assign g668 = (((!g290) & (!g622) & (g633) & (!g605) & (!g644)) + ((!g290) & (!g622) & (g633) & (g605) & (!g644)) + ((!g290) & (!g622) & (g633) & (g605) & (g644)) + ((!g290) & (g622) & (!g633) & (!g605) & (!g644)) + ((!g290) & (g622) & (!g633) & (!g605) & (g644)) + ((!g290) & (g622) & (!g633) & (g605) & (!g644)) + ((!g290) & (g622) & (!g633) & (g605) & (g644)) + ((!g290) & (g622) & (g633) & (!g605) & (g644)) + ((g290) & (!g622) & (!g633) & (!g605) & (!g644)) + ((g290) & (!g622) & (!g633) & (g605) & (!g644)) + ((g290) & (!g622) & (!g633) & (g605) & (g644)) + ((g290) & (g622) & (!g633) & (!g605) & (g644)) + ((g290) & (g622) & (g633) & (!g605) & (!g644)) + ((g290) & (g622) & (g633) & (!g605) & (g644)) + ((g290) & (g622) & (g633) & (g605) & (!g644)) + ((g290) & (g622) & (g633) & (g605) & (g644)));
	assign g669 = (((!g319) & (!g358) & (g624) & (g632)) + ((!g319) & (g358) & (!g624) & (g632)) + ((!g319) & (g358) & (g624) & (!g632)) + ((!g319) & (g358) & (g624) & (g632)) + ((g319) & (!g358) & (!g624) & (!g632)) + ((g319) & (!g358) & (!g624) & (g632)) + ((g319) & (!g358) & (g624) & (!g632)) + ((g319) & (g358) & (!g624) & (!g632)));
	assign g670 = (((!g623) & (!g605) & (!g644) & (g669)) + ((!g623) & (g605) & (!g644) & (g669)) + ((!g623) & (g605) & (g644) & (g669)) + ((g623) & (!g605) & (!g644) & (!g669)) + ((g623) & (!g605) & (g644) & (!g669)) + ((g623) & (!g605) & (g644) & (g669)) + ((g623) & (g605) & (!g644) & (!g669)) + ((g623) & (g605) & (g644) & (!g669)));
	assign g671 = (((!g358) & (!g624) & (g632) & (!g605) & (!g644)) + ((!g358) & (!g624) & (g632) & (g605) & (!g644)) + ((!g358) & (!g624) & (g632) & (g605) & (g644)) + ((!g358) & (g624) & (!g632) & (!g605) & (!g644)) + ((!g358) & (g624) & (!g632) & (!g605) & (g644)) + ((!g358) & (g624) & (!g632) & (g605) & (!g644)) + ((!g358) & (g624) & (!g632) & (g605) & (g644)) + ((!g358) & (g624) & (g632) & (!g605) & (g644)) + ((g358) & (!g624) & (!g632) & (!g605) & (!g644)) + ((g358) & (!g624) & (!g632) & (g605) & (!g644)) + ((g358) & (!g624) & (!g632) & (g605) & (g644)) + ((g358) & (g624) & (!g632) & (!g605) & (g644)) + ((g358) & (g624) & (g632) & (!g605) & (!g644)) + ((g358) & (g624) & (g632) & (!g605) & (g644)) + ((g358) & (g624) & (g632) & (g605) & (!g644)) + ((g358) & (g624) & (g632) & (g605) & (g644)));
	assign g672 = (((!g390) & (!g433) & (g626) & (g631)) + ((!g390) & (g433) & (!g626) & (g631)) + ((!g390) & (g433) & (g626) & (!g631)) + ((!g390) & (g433) & (g626) & (g631)) + ((g390) & (!g433) & (!g626) & (!g631)) + ((g390) & (!g433) & (!g626) & (g631)) + ((g390) & (!g433) & (g626) & (!g631)) + ((g390) & (g433) & (!g626) & (!g631)));
	assign g673 = (((!g625) & (!g605) & (!g644) & (g672)) + ((!g625) & (g605) & (!g644) & (g672)) + ((!g625) & (g605) & (g644) & (g672)) + ((g625) & (!g605) & (!g644) & (!g672)) + ((g625) & (!g605) & (g644) & (!g672)) + ((g625) & (!g605) & (g644) & (g672)) + ((g625) & (g605) & (!g644) & (!g672)) + ((g625) & (g605) & (g644) & (!g672)));
	assign g674 = (((!g433) & (!g626) & (g631) & (!g605) & (!g644)) + ((!g433) & (!g626) & (g631) & (g605) & (!g644)) + ((!g433) & (!g626) & (g631) & (g605) & (g644)) + ((!g433) & (g626) & (!g631) & (!g605) & (!g644)) + ((!g433) & (g626) & (!g631) & (!g605) & (g644)) + ((!g433) & (g626) & (!g631) & (g605) & (!g644)) + ((!g433) & (g626) & (!g631) & (g605) & (g644)) + ((!g433) & (g626) & (g631) & (!g605) & (g644)) + ((g433) & (!g626) & (!g631) & (!g605) & (!g644)) + ((g433) & (!g626) & (!g631) & (g605) & (!g644)) + ((g433) & (!g626) & (!g631) & (g605) & (g644)) + ((g433) & (g626) & (!g631) & (!g605) & (g644)) + ((g433) & (g626) & (g631) & (!g605) & (!g644)) + ((g433) & (g626) & (g631) & (!g605) & (g644)) + ((g433) & (g626) & (g631) & (g605) & (!g644)) + ((g433) & (g626) & (g631) & (g605) & (g644)));
	assign g675 = (((!g468) & (!g515) & (g628) & (g630)) + ((!g468) & (g515) & (!g628) & (g630)) + ((!g468) & (g515) & (g628) & (!g630)) + ((!g468) & (g515) & (g628) & (g630)) + ((g468) & (!g515) & (!g628) & (!g630)) + ((g468) & (!g515) & (!g628) & (g630)) + ((g468) & (!g515) & (g628) & (!g630)) + ((g468) & (g515) & (!g628) & (!g630)));
	assign g676 = (((!g627) & (!g605) & (!g644) & (g675)) + ((!g627) & (g605) & (!g644) & (g675)) + ((!g627) & (g605) & (g644) & (g675)) + ((g627) & (!g605) & (!g644) & (!g675)) + ((g627) & (!g605) & (g644) & (!g675)) + ((g627) & (!g605) & (g644) & (g675)) + ((g627) & (g605) & (!g644) & (!g675)) + ((g627) & (g605) & (g644) & (!g675)));
	assign g677 = (((!g515) & (!g628) & (g630) & (!g605) & (!g644)) + ((!g515) & (!g628) & (g630) & (g605) & (!g644)) + ((!g515) & (!g628) & (g630) & (g605) & (g644)) + ((!g515) & (g628) & (!g630) & (!g605) & (!g644)) + ((!g515) & (g628) & (!g630) & (!g605) & (g644)) + ((!g515) & (g628) & (!g630) & (g605) & (!g644)) + ((!g515) & (g628) & (!g630) & (g605) & (g644)) + ((!g515) & (g628) & (g630) & (!g605) & (g644)) + ((g515) & (!g628) & (!g630) & (!g605) & (!g644)) + ((g515) & (!g628) & (!g630) & (g605) & (!g644)) + ((g515) & (!g628) & (!g630) & (g605) & (g644)) + ((g515) & (g628) & (!g630) & (!g605) & (g644)) + ((g515) & (g628) & (g630) & (!g605) & (!g644)) + ((g515) & (g628) & (g630) & (!g605) & (g644)) + ((g515) & (g628) & (g630) & (g605) & (!g644)) + ((g515) & (g628) & (g630) & (g605) & (g644)));
	assign g678 = (((!g553) & (!ax76x) & (!g604) & (g629)) + ((!g553) & (!ax76x) & (g604) & (g629)) + ((!g553) & (ax76x) & (!g604) & (!g629)) + ((!g553) & (ax76x) & (!g604) & (g629)) + ((g553) & (!ax76x) & (!g604) & (!g629)) + ((g553) & (!ax76x) & (g604) & (!g629)) + ((g553) & (ax76x) & (g604) & (!g629)) + ((g553) & (ax76x) & (g604) & (g629)));
	assign g679 = (((!ax76x) & (!ax77x) & (!g604) & (!g605) & (!g644) & (g678)) + ((!ax76x) & (!ax77x) & (!g604) & (!g605) & (g644) & (!g678)) + ((!ax76x) & (!ax77x) & (!g604) & (!g605) & (g644) & (g678)) + ((!ax76x) & (!ax77x) & (!g604) & (g605) & (!g644) & (g678)) + ((!ax76x) & (!ax77x) & (!g604) & (g605) & (g644) & (g678)) + ((!ax76x) & (!ax77x) & (g604) & (!g605) & (!g644) & (!g678)) + ((!ax76x) & (!ax77x) & (g604) & (g605) & (!g644) & (!g678)) + ((!ax76x) & (!ax77x) & (g604) & (g605) & (g644) & (!g678)) + ((!ax76x) & (ax77x) & (!g604) & (!g605) & (!g644) & (!g678)) + ((!ax76x) & (ax77x) & (!g604) & (g605) & (!g644) & (!g678)) + ((!ax76x) & (ax77x) & (!g604) & (g605) & (g644) & (!g678)) + ((!ax76x) & (ax77x) & (g604) & (!g605) & (!g644) & (g678)) + ((!ax76x) & (ax77x) & (g604) & (!g605) & (g644) & (!g678)) + ((!ax76x) & (ax77x) & (g604) & (!g605) & (g644) & (g678)) + ((!ax76x) & (ax77x) & (g604) & (g605) & (!g644) & (g678)) + ((!ax76x) & (ax77x) & (g604) & (g605) & (g644) & (g678)) + ((ax76x) & (!ax77x) & (!g604) & (!g605) & (!g644) & (!g678)) + ((ax76x) & (!ax77x) & (!g604) & (g605) & (!g644) & (!g678)) + ((ax76x) & (!ax77x) & (!g604) & (g605) & (g644) & (!g678)) + ((ax76x) & (!ax77x) & (g604) & (!g605) & (!g644) & (!g678)) + ((ax76x) & (!ax77x) & (g604) & (g605) & (!g644) & (!g678)) + ((ax76x) & (!ax77x) & (g604) & (g605) & (g644) & (!g678)) + ((ax76x) & (ax77x) & (!g604) & (!g605) & (!g644) & (g678)) + ((ax76x) & (ax77x) & (!g604) & (!g605) & (g644) & (!g678)) + ((ax76x) & (ax77x) & (!g604) & (!g605) & (g644) & (g678)) + ((ax76x) & (ax77x) & (!g604) & (g605) & (!g644) & (g678)) + ((ax76x) & (ax77x) & (!g604) & (g605) & (g644) & (g678)) + ((ax76x) & (ax77x) & (g604) & (!g605) & (!g644) & (g678)) + ((ax76x) & (ax77x) & (g604) & (!g605) & (g644) & (!g678)) + ((ax76x) & (ax77x) & (g604) & (!g605) & (g644) & (g678)) + ((ax76x) & (ax77x) & (g604) & (g605) & (!g644) & (g678)) + ((ax76x) & (ax77x) & (g604) & (g605) & (g644) & (g678)));
	assign g680 = (((!ax76x) & (!g604) & (!g629) & (!g605) & (g644)) + ((!ax76x) & (!g604) & (g629) & (!g605) & (!g644)) + ((!ax76x) & (!g604) & (g629) & (!g605) & (g644)) + ((!ax76x) & (!g604) & (g629) & (g605) & (!g644)) + ((!ax76x) & (!g604) & (g629) & (g605) & (g644)) + ((!ax76x) & (g604) & (g629) & (!g605) & (!g644)) + ((!ax76x) & (g604) & (g629) & (g605) & (!g644)) + ((!ax76x) & (g604) & (g629) & (g605) & (g644)) + ((ax76x) & (!g604) & (!g629) & (!g605) & (!g644)) + ((ax76x) & (!g604) & (!g629) & (g605) & (!g644)) + ((ax76x) & (!g604) & (!g629) & (g605) & (g644)) + ((ax76x) & (g604) & (!g629) & (!g605) & (!g644)) + ((ax76x) & (g604) & (!g629) & (!g605) & (g644)) + ((ax76x) & (g604) & (!g629) & (g605) & (!g644)) + ((ax76x) & (g604) & (!g629) & (g605) & (g644)) + ((ax76x) & (g604) & (g629) & (!g605) & (g644)));
	assign g681 = (((!ax72x) & (!ax73x)));
	assign g682 = (((!g604) & (!ax74x) & (!ax75x) & (!g605) & (!g644) & (!g681)) + ((!g604) & (!ax74x) & (!ax75x) & (g605) & (!g644) & (!g681)) + ((!g604) & (!ax74x) & (!ax75x) & (g605) & (g644) & (!g681)) + ((!g604) & (!ax74x) & (ax75x) & (!g605) & (g644) & (!g681)) + ((!g604) & (ax74x) & (ax75x) & (!g605) & (g644) & (!g681)) + ((!g604) & (ax74x) & (ax75x) & (!g605) & (g644) & (g681)) + ((g604) & (!ax74x) & (!ax75x) & (!g605) & (!g644) & (!g681)) + ((g604) & (!ax74x) & (!ax75x) & (!g605) & (!g644) & (g681)) + ((g604) & (!ax74x) & (!ax75x) & (!g605) & (g644) & (!g681)) + ((g604) & (!ax74x) & (!ax75x) & (g605) & (!g644) & (!g681)) + ((g604) & (!ax74x) & (!ax75x) & (g605) & (!g644) & (g681)) + ((g604) & (!ax74x) & (!ax75x) & (g605) & (g644) & (!g681)) + ((g604) & (!ax74x) & (!ax75x) & (g605) & (g644) & (g681)) + ((g604) & (!ax74x) & (ax75x) & (!g605) & (!g644) & (!g681)) + ((g604) & (!ax74x) & (ax75x) & (!g605) & (g644) & (!g681)) + ((g604) & (!ax74x) & (ax75x) & (!g605) & (g644) & (g681)) + ((g604) & (!ax74x) & (ax75x) & (g605) & (!g644) & (!g681)) + ((g604) & (!ax74x) & (ax75x) & (g605) & (g644) & (!g681)) + ((g604) & (ax74x) & (!ax75x) & (!g605) & (g644) & (!g681)) + ((g604) & (ax74x) & (!ax75x) & (!g605) & (g644) & (g681)) + ((g604) & (ax74x) & (ax75x) & (!g605) & (!g644) & (!g681)) + ((g604) & (ax74x) & (ax75x) & (!g605) & (!g644) & (g681)) + ((g604) & (ax74x) & (ax75x) & (!g605) & (g644) & (!g681)) + ((g604) & (ax74x) & (ax75x) & (!g605) & (g644) & (g681)) + ((g604) & (ax74x) & (ax75x) & (g605) & (!g644) & (!g681)) + ((g604) & (ax74x) & (ax75x) & (g605) & (!g644) & (g681)) + ((g604) & (ax74x) & (ax75x) & (g605) & (g644) & (!g681)) + ((g604) & (ax74x) & (ax75x) & (g605) & (g644) & (g681)));
	assign g683 = (((!g515) & (!g553) & (g679) & (g680) & (g682)) + ((!g515) & (g553) & (g679) & (!g680) & (g682)) + ((!g515) & (g553) & (g679) & (g680) & (!g682)) + ((!g515) & (g553) & (g679) & (g680) & (g682)) + ((g515) & (!g553) & (!g679) & (g680) & (g682)) + ((g515) & (!g553) & (g679) & (!g680) & (!g682)) + ((g515) & (!g553) & (g679) & (!g680) & (g682)) + ((g515) & (!g553) & (g679) & (g680) & (!g682)) + ((g515) & (!g553) & (g679) & (g680) & (g682)) + ((g515) & (g553) & (!g679) & (!g680) & (g682)) + ((g515) & (g553) & (!g679) & (g680) & (!g682)) + ((g515) & (g553) & (!g679) & (g680) & (g682)) + ((g515) & (g553) & (g679) & (!g680) & (!g682)) + ((g515) & (g553) & (g679) & (!g680) & (g682)) + ((g515) & (g553) & (g679) & (g680) & (!g682)) + ((g515) & (g553) & (g679) & (g680) & (g682)));
	assign g684 = (((!g433) & (!g468) & (g676) & (g677) & (g683)) + ((!g433) & (g468) & (g676) & (!g677) & (g683)) + ((!g433) & (g468) & (g676) & (g677) & (!g683)) + ((!g433) & (g468) & (g676) & (g677) & (g683)) + ((g433) & (!g468) & (!g676) & (g677) & (g683)) + ((g433) & (!g468) & (g676) & (!g677) & (!g683)) + ((g433) & (!g468) & (g676) & (!g677) & (g683)) + ((g433) & (!g468) & (g676) & (g677) & (!g683)) + ((g433) & (!g468) & (g676) & (g677) & (g683)) + ((g433) & (g468) & (!g676) & (!g677) & (g683)) + ((g433) & (g468) & (!g676) & (g677) & (!g683)) + ((g433) & (g468) & (!g676) & (g677) & (g683)) + ((g433) & (g468) & (g676) & (!g677) & (!g683)) + ((g433) & (g468) & (g676) & (!g677) & (g683)) + ((g433) & (g468) & (g676) & (g677) & (!g683)) + ((g433) & (g468) & (g676) & (g677) & (g683)));
	assign g685 = (((!g358) & (!g390) & (g673) & (g674) & (g684)) + ((!g358) & (g390) & (g673) & (!g674) & (g684)) + ((!g358) & (g390) & (g673) & (g674) & (!g684)) + ((!g358) & (g390) & (g673) & (g674) & (g684)) + ((g358) & (!g390) & (!g673) & (g674) & (g684)) + ((g358) & (!g390) & (g673) & (!g674) & (!g684)) + ((g358) & (!g390) & (g673) & (!g674) & (g684)) + ((g358) & (!g390) & (g673) & (g674) & (!g684)) + ((g358) & (!g390) & (g673) & (g674) & (g684)) + ((g358) & (g390) & (!g673) & (!g674) & (g684)) + ((g358) & (g390) & (!g673) & (g674) & (!g684)) + ((g358) & (g390) & (!g673) & (g674) & (g684)) + ((g358) & (g390) & (g673) & (!g674) & (!g684)) + ((g358) & (g390) & (g673) & (!g674) & (g684)) + ((g358) & (g390) & (g673) & (g674) & (!g684)) + ((g358) & (g390) & (g673) & (g674) & (g684)));
	assign g686 = (((!g290) & (!g319) & (g670) & (g671) & (g685)) + ((!g290) & (g319) & (g670) & (!g671) & (g685)) + ((!g290) & (g319) & (g670) & (g671) & (!g685)) + ((!g290) & (g319) & (g670) & (g671) & (g685)) + ((g290) & (!g319) & (!g670) & (g671) & (g685)) + ((g290) & (!g319) & (g670) & (!g671) & (!g685)) + ((g290) & (!g319) & (g670) & (!g671) & (g685)) + ((g290) & (!g319) & (g670) & (g671) & (!g685)) + ((g290) & (!g319) & (g670) & (g671) & (g685)) + ((g290) & (g319) & (!g670) & (!g671) & (g685)) + ((g290) & (g319) & (!g670) & (g671) & (!g685)) + ((g290) & (g319) & (!g670) & (g671) & (g685)) + ((g290) & (g319) & (g670) & (!g671) & (!g685)) + ((g290) & (g319) & (g670) & (!g671) & (g685)) + ((g290) & (g319) & (g670) & (g671) & (!g685)) + ((g290) & (g319) & (g670) & (g671) & (g685)));
	assign g687 = (((!g229) & (!g255) & (g667) & (g668) & (g686)) + ((!g229) & (g255) & (g667) & (!g668) & (g686)) + ((!g229) & (g255) & (g667) & (g668) & (!g686)) + ((!g229) & (g255) & (g667) & (g668) & (g686)) + ((g229) & (!g255) & (!g667) & (g668) & (g686)) + ((g229) & (!g255) & (g667) & (!g668) & (!g686)) + ((g229) & (!g255) & (g667) & (!g668) & (g686)) + ((g229) & (!g255) & (g667) & (g668) & (!g686)) + ((g229) & (!g255) & (g667) & (g668) & (g686)) + ((g229) & (g255) & (!g667) & (!g668) & (g686)) + ((g229) & (g255) & (!g667) & (g668) & (!g686)) + ((g229) & (g255) & (!g667) & (g668) & (g686)) + ((g229) & (g255) & (g667) & (!g668) & (!g686)) + ((g229) & (g255) & (g667) & (!g668) & (g686)) + ((g229) & (g255) & (g667) & (g668) & (!g686)) + ((g229) & (g255) & (g667) & (g668) & (g686)));
	assign g688 = (((!g174) & (!g198) & (g664) & (g665) & (g687)) + ((!g174) & (g198) & (g664) & (!g665) & (g687)) + ((!g174) & (g198) & (g664) & (g665) & (!g687)) + ((!g174) & (g198) & (g664) & (g665) & (g687)) + ((g174) & (!g198) & (!g664) & (g665) & (g687)) + ((g174) & (!g198) & (g664) & (!g665) & (!g687)) + ((g174) & (!g198) & (g664) & (!g665) & (g687)) + ((g174) & (!g198) & (g664) & (g665) & (!g687)) + ((g174) & (!g198) & (g664) & (g665) & (g687)) + ((g174) & (g198) & (!g664) & (!g665) & (g687)) + ((g174) & (g198) & (!g664) & (g665) & (!g687)) + ((g174) & (g198) & (!g664) & (g665) & (g687)) + ((g174) & (g198) & (g664) & (!g665) & (!g687)) + ((g174) & (g198) & (g664) & (!g665) & (g687)) + ((g174) & (g198) & (g664) & (g665) & (!g687)) + ((g174) & (g198) & (g664) & (g665) & (g687)));
	assign g689 = (((!g127) & (!g147) & (g661) & (g662) & (g688)) + ((!g127) & (g147) & (g661) & (!g662) & (g688)) + ((!g127) & (g147) & (g661) & (g662) & (!g688)) + ((!g127) & (g147) & (g661) & (g662) & (g688)) + ((g127) & (!g147) & (!g661) & (g662) & (g688)) + ((g127) & (!g147) & (g661) & (!g662) & (!g688)) + ((g127) & (!g147) & (g661) & (!g662) & (g688)) + ((g127) & (!g147) & (g661) & (g662) & (!g688)) + ((g127) & (!g147) & (g661) & (g662) & (g688)) + ((g127) & (g147) & (!g661) & (!g662) & (g688)) + ((g127) & (g147) & (!g661) & (g662) & (!g688)) + ((g127) & (g147) & (!g661) & (g662) & (g688)) + ((g127) & (g147) & (g661) & (!g662) & (!g688)) + ((g127) & (g147) & (g661) & (!g662) & (g688)) + ((g127) & (g147) & (g661) & (g662) & (!g688)) + ((g127) & (g147) & (g661) & (g662) & (g688)));
	assign g690 = (((!g87) & (!g104) & (g658) & (g659) & (g689)) + ((!g87) & (g104) & (g658) & (!g659) & (g689)) + ((!g87) & (g104) & (g658) & (g659) & (!g689)) + ((!g87) & (g104) & (g658) & (g659) & (g689)) + ((g87) & (!g104) & (!g658) & (g659) & (g689)) + ((g87) & (!g104) & (g658) & (!g659) & (!g689)) + ((g87) & (!g104) & (g658) & (!g659) & (g689)) + ((g87) & (!g104) & (g658) & (g659) & (!g689)) + ((g87) & (!g104) & (g658) & (g659) & (g689)) + ((g87) & (g104) & (!g658) & (!g659) & (g689)) + ((g87) & (g104) & (!g658) & (g659) & (!g689)) + ((g87) & (g104) & (!g658) & (g659) & (g689)) + ((g87) & (g104) & (g658) & (!g659) & (!g689)) + ((g87) & (g104) & (g658) & (!g659) & (g689)) + ((g87) & (g104) & (g658) & (g659) & (!g689)) + ((g87) & (g104) & (g658) & (g659) & (g689)));
	assign g691 = (((!g54) & (!g68) & (g655) & (g656) & (g690)) + ((!g54) & (g68) & (g655) & (!g656) & (g690)) + ((!g54) & (g68) & (g655) & (g656) & (!g690)) + ((!g54) & (g68) & (g655) & (g656) & (g690)) + ((g54) & (!g68) & (!g655) & (g656) & (g690)) + ((g54) & (!g68) & (g655) & (!g656) & (!g690)) + ((g54) & (!g68) & (g655) & (!g656) & (g690)) + ((g54) & (!g68) & (g655) & (g656) & (!g690)) + ((g54) & (!g68) & (g655) & (g656) & (g690)) + ((g54) & (g68) & (!g655) & (!g656) & (g690)) + ((g54) & (g68) & (!g655) & (g656) & (!g690)) + ((g54) & (g68) & (!g655) & (g656) & (g690)) + ((g54) & (g68) & (g655) & (!g656) & (!g690)) + ((g54) & (g68) & (g655) & (!g656) & (g690)) + ((g54) & (g68) & (g655) & (g656) & (!g690)) + ((g54) & (g68) & (g655) & (g656) & (g690)));
	assign g692 = (((!g27) & (!g39) & (g652) & (g653) & (g691)) + ((!g27) & (g39) & (g652) & (!g653) & (g691)) + ((!g27) & (g39) & (g652) & (g653) & (!g691)) + ((!g27) & (g39) & (g652) & (g653) & (g691)) + ((g27) & (!g39) & (!g652) & (g653) & (g691)) + ((g27) & (!g39) & (g652) & (!g653) & (!g691)) + ((g27) & (!g39) & (g652) & (!g653) & (g691)) + ((g27) & (!g39) & (g652) & (g653) & (!g691)) + ((g27) & (!g39) & (g652) & (g653) & (g691)) + ((g27) & (g39) & (!g652) & (!g653) & (g691)) + ((g27) & (g39) & (!g652) & (g653) & (!g691)) + ((g27) & (g39) & (!g652) & (g653) & (g691)) + ((g27) & (g39) & (g652) & (!g653) & (!g691)) + ((g27) & (g39) & (g652) & (!g653) & (g691)) + ((g27) & (g39) & (g652) & (g653) & (!g691)) + ((g27) & (g39) & (g652) & (g653) & (g691)));
	assign g693 = (((!g8) & (!g18) & (g649) & (g650) & (g692)) + ((!g8) & (g18) & (g649) & (!g650) & (g692)) + ((!g8) & (g18) & (g649) & (g650) & (!g692)) + ((!g8) & (g18) & (g649) & (g650) & (g692)) + ((g8) & (!g18) & (!g649) & (g650) & (g692)) + ((g8) & (!g18) & (g649) & (!g650) & (!g692)) + ((g8) & (!g18) & (g649) & (!g650) & (g692)) + ((g8) & (!g18) & (g649) & (g650) & (!g692)) + ((g8) & (!g18) & (g649) & (g650) & (g692)) + ((g8) & (g18) & (!g649) & (!g650) & (g692)) + ((g8) & (g18) & (!g649) & (g650) & (!g692)) + ((g8) & (g18) & (!g649) & (g650) & (g692)) + ((g8) & (g18) & (g649) & (!g650) & (!g692)) + ((g8) & (g18) & (g649) & (!g650) & (g692)) + ((g8) & (g18) & (g649) & (g650) & (!g692)) + ((g8) & (g18) & (g649) & (g650) & (g692)));
	assign g694 = (((!g2) & (!g8) & (g608) & (g640)) + ((!g2) & (g8) & (!g608) & (g640)) + ((!g2) & (g8) & (g608) & (!g640)) + ((!g2) & (g8) & (g608) & (g640)) + ((g2) & (!g8) & (!g608) & (!g640)) + ((g2) & (!g8) & (!g608) & (g640)) + ((g2) & (!g8) & (g608) & (!g640)) + ((g2) & (g8) & (!g608) & (!g640)));
	assign g695 = (((!g607) & (!g605) & (!g644) & (g694)) + ((!g607) & (g605) & (!g644) & (g694)) + ((!g607) & (g605) & (g644) & (g694)) + ((g607) & (!g605) & (!g644) & (!g694)) + ((g607) & (!g605) & (g644) & (!g694)) + ((g607) & (!g605) & (g644) & (g694)) + ((g607) & (g605) & (!g644) & (!g694)) + ((g607) & (g605) & (g644) & (!g694)));
	assign g696 = (((!g4) & (!g2) & (!g647) & (!g693) & (g695)) + ((!g4) & (!g2) & (!g647) & (g693) & (g695)) + ((!g4) & (!g2) & (g647) & (!g693) & (g695)) + ((!g4) & (!g2) & (g647) & (g693) & (!g695)) + ((!g4) & (!g2) & (g647) & (g693) & (g695)) + ((!g4) & (g2) & (!g647) & (!g693) & (g695)) + ((!g4) & (g2) & (!g647) & (g693) & (!g695)) + ((!g4) & (g2) & (!g647) & (g693) & (g695)) + ((!g4) & (g2) & (g647) & (!g693) & (!g695)) + ((!g4) & (g2) & (g647) & (!g693) & (g695)) + ((!g4) & (g2) & (g647) & (g693) & (!g695)) + ((!g4) & (g2) & (g647) & (g693) & (g695)) + ((g4) & (!g2) & (g647) & (g693) & (g695)) + ((g4) & (g2) & (!g647) & (g693) & (g695)) + ((g4) & (g2) & (g647) & (!g693) & (g695)) + ((g4) & (g2) & (g647) & (g693) & (g695)));
	assign g697 = (((!g4) & (!g641) & (g642)) + ((!g4) & (g641) & (!g642)) + ((!g4) & (g641) & (g642)) + ((g4) & (g641) & (g642)));
	assign g698 = (((!g606) & (!g697) & (!g605) & (!g644)) + ((!g606) & (!g697) & (g605) & (!g644)) + ((!g606) & (!g697) & (g605) & (g644)) + ((g606) & (g697) & (!g605) & (!g644)) + ((g606) & (g697) & (!g605) & (g644)) + ((g606) & (g697) & (g605) & (!g644)) + ((g606) & (g697) & (g605) & (g644)));
	assign g699 = (((!g1) & (g606) & (!g697) & (!g605) & (g644)) + ((!g1) & (g606) & (g697) & (!g605) & (g644)) + ((g1) & (!g606) & (g697) & (g605) & (!g644)) + ((g1) & (!g606) & (g697) & (g605) & (g644)) + ((g1) & (g606) & (!g697) & (!g605) & (!g644)) + ((g1) & (g606) & (!g697) & (!g605) & (g644)) + ((g1) & (g606) & (!g697) & (g605) & (!g644)) + ((g1) & (g606) & (!g697) & (g605) & (g644)) + ((g1) & (g606) & (g697) & (!g605) & (g644)));
	assign g700 = (((!g1) & (!g646) & (!g696) & (!g698) & (!g699)) + ((g1) & (!g646) & (!g696) & (!g698) & (!g699)) + ((g1) & (!g646) & (!g696) & (g698) & (!g699)) + ((g1) & (!g646) & (g696) & (!g698) & (!g699)) + ((g1) & (!g646) & (g696) & (g698) & (!g699)) + ((g1) & (g646) & (!g696) & (!g698) & (!g699)) + ((g1) & (g646) & (!g696) & (g698) & (!g699)));
	assign g701 = (((g1) & (!g646) & (g696) & (g699)) + ((g1) & (g646) & (!g696) & (!g699)) + ((g1) & (g646) & (!g696) & (g699)));
	assign g702 = (((!g4) & (!g2) & (!g647) & (!g693) & (!g695) & (!g700)) + ((!g4) & (!g2) & (!g647) & (!g693) & (g695) & (g700)) + ((!g4) & (!g2) & (!g647) & (g693) & (!g695) & (!g700)) + ((!g4) & (!g2) & (!g647) & (g693) & (g695) & (g700)) + ((!g4) & (!g2) & (g647) & (!g693) & (!g695) & (!g700)) + ((!g4) & (!g2) & (g647) & (!g693) & (g695) & (g700)) + ((!g4) & (!g2) & (g647) & (g693) & (g695) & (!g700)) + ((!g4) & (!g2) & (g647) & (g693) & (g695) & (g700)) + ((!g4) & (g2) & (!g647) & (!g693) & (!g695) & (!g700)) + ((!g4) & (g2) & (!g647) & (!g693) & (g695) & (g700)) + ((!g4) & (g2) & (!g647) & (g693) & (g695) & (!g700)) + ((!g4) & (g2) & (!g647) & (g693) & (g695) & (g700)) + ((!g4) & (g2) & (g647) & (!g693) & (g695) & (!g700)) + ((!g4) & (g2) & (g647) & (!g693) & (g695) & (g700)) + ((!g4) & (g2) & (g647) & (g693) & (g695) & (!g700)) + ((!g4) & (g2) & (g647) & (g693) & (g695) & (g700)) + ((g4) & (!g2) & (!g647) & (!g693) & (g695) & (!g700)) + ((g4) & (!g2) & (!g647) & (!g693) & (g695) & (g700)) + ((g4) & (!g2) & (!g647) & (g693) & (g695) & (!g700)) + ((g4) & (!g2) & (!g647) & (g693) & (g695) & (g700)) + ((g4) & (!g2) & (g647) & (!g693) & (g695) & (!g700)) + ((g4) & (!g2) & (g647) & (!g693) & (g695) & (g700)) + ((g4) & (!g2) & (g647) & (g693) & (!g695) & (!g700)) + ((g4) & (!g2) & (g647) & (g693) & (g695) & (g700)) + ((g4) & (g2) & (!g647) & (!g693) & (g695) & (!g700)) + ((g4) & (g2) & (!g647) & (!g693) & (g695) & (g700)) + ((g4) & (g2) & (!g647) & (g693) & (!g695) & (!g700)) + ((g4) & (g2) & (!g647) & (g693) & (g695) & (g700)) + ((g4) & (g2) & (g647) & (!g693) & (!g695) & (!g700)) + ((g4) & (g2) & (g647) & (!g693) & (g695) & (g700)) + ((g4) & (g2) & (g647) & (g693) & (!g695) & (!g700)) + ((g4) & (g2) & (g647) & (g693) & (g695) & (g700)));
	assign g703 = (((!g8) & (!g18) & (!g649) & (g650) & (g692) & (!g700)) + ((!g8) & (!g18) & (g649) & (!g650) & (!g692) & (!g700)) + ((!g8) & (!g18) & (g649) & (!g650) & (!g692) & (g700)) + ((!g8) & (!g18) & (g649) & (!g650) & (g692) & (!g700)) + ((!g8) & (!g18) & (g649) & (!g650) & (g692) & (g700)) + ((!g8) & (!g18) & (g649) & (g650) & (!g692) & (!g700)) + ((!g8) & (!g18) & (g649) & (g650) & (!g692) & (g700)) + ((!g8) & (!g18) & (g649) & (g650) & (g692) & (g700)) + ((!g8) & (g18) & (!g649) & (!g650) & (g692) & (!g700)) + ((!g8) & (g18) & (!g649) & (g650) & (!g692) & (!g700)) + ((!g8) & (g18) & (!g649) & (g650) & (g692) & (!g700)) + ((!g8) & (g18) & (g649) & (!g650) & (!g692) & (!g700)) + ((!g8) & (g18) & (g649) & (!g650) & (!g692) & (g700)) + ((!g8) & (g18) & (g649) & (!g650) & (g692) & (g700)) + ((!g8) & (g18) & (g649) & (g650) & (!g692) & (g700)) + ((!g8) & (g18) & (g649) & (g650) & (g692) & (g700)) + ((g8) & (!g18) & (!g649) & (!g650) & (!g692) & (!g700)) + ((g8) & (!g18) & (!g649) & (!g650) & (g692) & (!g700)) + ((g8) & (!g18) & (!g649) & (g650) & (!g692) & (!g700)) + ((g8) & (!g18) & (g649) & (!g650) & (!g692) & (g700)) + ((g8) & (!g18) & (g649) & (!g650) & (g692) & (g700)) + ((g8) & (!g18) & (g649) & (g650) & (!g692) & (g700)) + ((g8) & (!g18) & (g649) & (g650) & (g692) & (!g700)) + ((g8) & (!g18) & (g649) & (g650) & (g692) & (g700)) + ((g8) & (g18) & (!g649) & (!g650) & (!g692) & (!g700)) + ((g8) & (g18) & (g649) & (!g650) & (!g692) & (g700)) + ((g8) & (g18) & (g649) & (!g650) & (g692) & (!g700)) + ((g8) & (g18) & (g649) & (!g650) & (g692) & (g700)) + ((g8) & (g18) & (g649) & (g650) & (!g692) & (!g700)) + ((g8) & (g18) & (g649) & (g650) & (!g692) & (g700)) + ((g8) & (g18) & (g649) & (g650) & (g692) & (!g700)) + ((g8) & (g18) & (g649) & (g650) & (g692) & (g700)));
	assign g704 = (((!g18) & (!g650) & (g692) & (!g700)) + ((!g18) & (g650) & (!g692) & (!g700)) + ((!g18) & (g650) & (!g692) & (g700)) + ((!g18) & (g650) & (g692) & (g700)) + ((g18) & (!g650) & (!g692) & (!g700)) + ((g18) & (g650) & (!g692) & (g700)) + ((g18) & (g650) & (g692) & (!g700)) + ((g18) & (g650) & (g692) & (g700)));
	assign g705 = (((!g27) & (!g39) & (!g652) & (g653) & (g691) & (!g700)) + ((!g27) & (!g39) & (g652) & (!g653) & (!g691) & (!g700)) + ((!g27) & (!g39) & (g652) & (!g653) & (!g691) & (g700)) + ((!g27) & (!g39) & (g652) & (!g653) & (g691) & (!g700)) + ((!g27) & (!g39) & (g652) & (!g653) & (g691) & (g700)) + ((!g27) & (!g39) & (g652) & (g653) & (!g691) & (!g700)) + ((!g27) & (!g39) & (g652) & (g653) & (!g691) & (g700)) + ((!g27) & (!g39) & (g652) & (g653) & (g691) & (g700)) + ((!g27) & (g39) & (!g652) & (!g653) & (g691) & (!g700)) + ((!g27) & (g39) & (!g652) & (g653) & (!g691) & (!g700)) + ((!g27) & (g39) & (!g652) & (g653) & (g691) & (!g700)) + ((!g27) & (g39) & (g652) & (!g653) & (!g691) & (!g700)) + ((!g27) & (g39) & (g652) & (!g653) & (!g691) & (g700)) + ((!g27) & (g39) & (g652) & (!g653) & (g691) & (g700)) + ((!g27) & (g39) & (g652) & (g653) & (!g691) & (g700)) + ((!g27) & (g39) & (g652) & (g653) & (g691) & (g700)) + ((g27) & (!g39) & (!g652) & (!g653) & (!g691) & (!g700)) + ((g27) & (!g39) & (!g652) & (!g653) & (g691) & (!g700)) + ((g27) & (!g39) & (!g652) & (g653) & (!g691) & (!g700)) + ((g27) & (!g39) & (g652) & (!g653) & (!g691) & (g700)) + ((g27) & (!g39) & (g652) & (!g653) & (g691) & (g700)) + ((g27) & (!g39) & (g652) & (g653) & (!g691) & (g700)) + ((g27) & (!g39) & (g652) & (g653) & (g691) & (!g700)) + ((g27) & (!g39) & (g652) & (g653) & (g691) & (g700)) + ((g27) & (g39) & (!g652) & (!g653) & (!g691) & (!g700)) + ((g27) & (g39) & (g652) & (!g653) & (!g691) & (g700)) + ((g27) & (g39) & (g652) & (!g653) & (g691) & (!g700)) + ((g27) & (g39) & (g652) & (!g653) & (g691) & (g700)) + ((g27) & (g39) & (g652) & (g653) & (!g691) & (!g700)) + ((g27) & (g39) & (g652) & (g653) & (!g691) & (g700)) + ((g27) & (g39) & (g652) & (g653) & (g691) & (!g700)) + ((g27) & (g39) & (g652) & (g653) & (g691) & (g700)));
	assign g706 = (((!g39) & (!g653) & (g691) & (!g700)) + ((!g39) & (g653) & (!g691) & (!g700)) + ((!g39) & (g653) & (!g691) & (g700)) + ((!g39) & (g653) & (g691) & (g700)) + ((g39) & (!g653) & (!g691) & (!g700)) + ((g39) & (g653) & (!g691) & (g700)) + ((g39) & (g653) & (g691) & (!g700)) + ((g39) & (g653) & (g691) & (g700)));
	assign g707 = (((!g54) & (!g68) & (!g655) & (g656) & (g690) & (!g700)) + ((!g54) & (!g68) & (g655) & (!g656) & (!g690) & (!g700)) + ((!g54) & (!g68) & (g655) & (!g656) & (!g690) & (g700)) + ((!g54) & (!g68) & (g655) & (!g656) & (g690) & (!g700)) + ((!g54) & (!g68) & (g655) & (!g656) & (g690) & (g700)) + ((!g54) & (!g68) & (g655) & (g656) & (!g690) & (!g700)) + ((!g54) & (!g68) & (g655) & (g656) & (!g690) & (g700)) + ((!g54) & (!g68) & (g655) & (g656) & (g690) & (g700)) + ((!g54) & (g68) & (!g655) & (!g656) & (g690) & (!g700)) + ((!g54) & (g68) & (!g655) & (g656) & (!g690) & (!g700)) + ((!g54) & (g68) & (!g655) & (g656) & (g690) & (!g700)) + ((!g54) & (g68) & (g655) & (!g656) & (!g690) & (!g700)) + ((!g54) & (g68) & (g655) & (!g656) & (!g690) & (g700)) + ((!g54) & (g68) & (g655) & (!g656) & (g690) & (g700)) + ((!g54) & (g68) & (g655) & (g656) & (!g690) & (g700)) + ((!g54) & (g68) & (g655) & (g656) & (g690) & (g700)) + ((g54) & (!g68) & (!g655) & (!g656) & (!g690) & (!g700)) + ((g54) & (!g68) & (!g655) & (!g656) & (g690) & (!g700)) + ((g54) & (!g68) & (!g655) & (g656) & (!g690) & (!g700)) + ((g54) & (!g68) & (g655) & (!g656) & (!g690) & (g700)) + ((g54) & (!g68) & (g655) & (!g656) & (g690) & (g700)) + ((g54) & (!g68) & (g655) & (g656) & (!g690) & (g700)) + ((g54) & (!g68) & (g655) & (g656) & (g690) & (!g700)) + ((g54) & (!g68) & (g655) & (g656) & (g690) & (g700)) + ((g54) & (g68) & (!g655) & (!g656) & (!g690) & (!g700)) + ((g54) & (g68) & (g655) & (!g656) & (!g690) & (g700)) + ((g54) & (g68) & (g655) & (!g656) & (g690) & (!g700)) + ((g54) & (g68) & (g655) & (!g656) & (g690) & (g700)) + ((g54) & (g68) & (g655) & (g656) & (!g690) & (!g700)) + ((g54) & (g68) & (g655) & (g656) & (!g690) & (g700)) + ((g54) & (g68) & (g655) & (g656) & (g690) & (!g700)) + ((g54) & (g68) & (g655) & (g656) & (g690) & (g700)));
	assign g708 = (((!g68) & (!g656) & (g690) & (!g700)) + ((!g68) & (g656) & (!g690) & (!g700)) + ((!g68) & (g656) & (!g690) & (g700)) + ((!g68) & (g656) & (g690) & (g700)) + ((g68) & (!g656) & (!g690) & (!g700)) + ((g68) & (g656) & (!g690) & (g700)) + ((g68) & (g656) & (g690) & (!g700)) + ((g68) & (g656) & (g690) & (g700)));
	assign g709 = (((!g87) & (!g104) & (!g658) & (g659) & (g689) & (!g700)) + ((!g87) & (!g104) & (g658) & (!g659) & (!g689) & (!g700)) + ((!g87) & (!g104) & (g658) & (!g659) & (!g689) & (g700)) + ((!g87) & (!g104) & (g658) & (!g659) & (g689) & (!g700)) + ((!g87) & (!g104) & (g658) & (!g659) & (g689) & (g700)) + ((!g87) & (!g104) & (g658) & (g659) & (!g689) & (!g700)) + ((!g87) & (!g104) & (g658) & (g659) & (!g689) & (g700)) + ((!g87) & (!g104) & (g658) & (g659) & (g689) & (g700)) + ((!g87) & (g104) & (!g658) & (!g659) & (g689) & (!g700)) + ((!g87) & (g104) & (!g658) & (g659) & (!g689) & (!g700)) + ((!g87) & (g104) & (!g658) & (g659) & (g689) & (!g700)) + ((!g87) & (g104) & (g658) & (!g659) & (!g689) & (!g700)) + ((!g87) & (g104) & (g658) & (!g659) & (!g689) & (g700)) + ((!g87) & (g104) & (g658) & (!g659) & (g689) & (g700)) + ((!g87) & (g104) & (g658) & (g659) & (!g689) & (g700)) + ((!g87) & (g104) & (g658) & (g659) & (g689) & (g700)) + ((g87) & (!g104) & (!g658) & (!g659) & (!g689) & (!g700)) + ((g87) & (!g104) & (!g658) & (!g659) & (g689) & (!g700)) + ((g87) & (!g104) & (!g658) & (g659) & (!g689) & (!g700)) + ((g87) & (!g104) & (g658) & (!g659) & (!g689) & (g700)) + ((g87) & (!g104) & (g658) & (!g659) & (g689) & (g700)) + ((g87) & (!g104) & (g658) & (g659) & (!g689) & (g700)) + ((g87) & (!g104) & (g658) & (g659) & (g689) & (!g700)) + ((g87) & (!g104) & (g658) & (g659) & (g689) & (g700)) + ((g87) & (g104) & (!g658) & (!g659) & (!g689) & (!g700)) + ((g87) & (g104) & (g658) & (!g659) & (!g689) & (g700)) + ((g87) & (g104) & (g658) & (!g659) & (g689) & (!g700)) + ((g87) & (g104) & (g658) & (!g659) & (g689) & (g700)) + ((g87) & (g104) & (g658) & (g659) & (!g689) & (!g700)) + ((g87) & (g104) & (g658) & (g659) & (!g689) & (g700)) + ((g87) & (g104) & (g658) & (g659) & (g689) & (!g700)) + ((g87) & (g104) & (g658) & (g659) & (g689) & (g700)));
	assign g710 = (((!g104) & (!g659) & (g689) & (!g700)) + ((!g104) & (g659) & (!g689) & (!g700)) + ((!g104) & (g659) & (!g689) & (g700)) + ((!g104) & (g659) & (g689) & (g700)) + ((g104) & (!g659) & (!g689) & (!g700)) + ((g104) & (g659) & (!g689) & (g700)) + ((g104) & (g659) & (g689) & (!g700)) + ((g104) & (g659) & (g689) & (g700)));
	assign g711 = (((!g127) & (!g147) & (!g661) & (g662) & (g688) & (!g700)) + ((!g127) & (!g147) & (g661) & (!g662) & (!g688) & (!g700)) + ((!g127) & (!g147) & (g661) & (!g662) & (!g688) & (g700)) + ((!g127) & (!g147) & (g661) & (!g662) & (g688) & (!g700)) + ((!g127) & (!g147) & (g661) & (!g662) & (g688) & (g700)) + ((!g127) & (!g147) & (g661) & (g662) & (!g688) & (!g700)) + ((!g127) & (!g147) & (g661) & (g662) & (!g688) & (g700)) + ((!g127) & (!g147) & (g661) & (g662) & (g688) & (g700)) + ((!g127) & (g147) & (!g661) & (!g662) & (g688) & (!g700)) + ((!g127) & (g147) & (!g661) & (g662) & (!g688) & (!g700)) + ((!g127) & (g147) & (!g661) & (g662) & (g688) & (!g700)) + ((!g127) & (g147) & (g661) & (!g662) & (!g688) & (!g700)) + ((!g127) & (g147) & (g661) & (!g662) & (!g688) & (g700)) + ((!g127) & (g147) & (g661) & (!g662) & (g688) & (g700)) + ((!g127) & (g147) & (g661) & (g662) & (!g688) & (g700)) + ((!g127) & (g147) & (g661) & (g662) & (g688) & (g700)) + ((g127) & (!g147) & (!g661) & (!g662) & (!g688) & (!g700)) + ((g127) & (!g147) & (!g661) & (!g662) & (g688) & (!g700)) + ((g127) & (!g147) & (!g661) & (g662) & (!g688) & (!g700)) + ((g127) & (!g147) & (g661) & (!g662) & (!g688) & (g700)) + ((g127) & (!g147) & (g661) & (!g662) & (g688) & (g700)) + ((g127) & (!g147) & (g661) & (g662) & (!g688) & (g700)) + ((g127) & (!g147) & (g661) & (g662) & (g688) & (!g700)) + ((g127) & (!g147) & (g661) & (g662) & (g688) & (g700)) + ((g127) & (g147) & (!g661) & (!g662) & (!g688) & (!g700)) + ((g127) & (g147) & (g661) & (!g662) & (!g688) & (g700)) + ((g127) & (g147) & (g661) & (!g662) & (g688) & (!g700)) + ((g127) & (g147) & (g661) & (!g662) & (g688) & (g700)) + ((g127) & (g147) & (g661) & (g662) & (!g688) & (!g700)) + ((g127) & (g147) & (g661) & (g662) & (!g688) & (g700)) + ((g127) & (g147) & (g661) & (g662) & (g688) & (!g700)) + ((g127) & (g147) & (g661) & (g662) & (g688) & (g700)));
	assign g712 = (((!g147) & (!g662) & (g688) & (!g700)) + ((!g147) & (g662) & (!g688) & (!g700)) + ((!g147) & (g662) & (!g688) & (g700)) + ((!g147) & (g662) & (g688) & (g700)) + ((g147) & (!g662) & (!g688) & (!g700)) + ((g147) & (g662) & (!g688) & (g700)) + ((g147) & (g662) & (g688) & (!g700)) + ((g147) & (g662) & (g688) & (g700)));
	assign g713 = (((!g174) & (!g198) & (!g664) & (g665) & (g687) & (!g700)) + ((!g174) & (!g198) & (g664) & (!g665) & (!g687) & (!g700)) + ((!g174) & (!g198) & (g664) & (!g665) & (!g687) & (g700)) + ((!g174) & (!g198) & (g664) & (!g665) & (g687) & (!g700)) + ((!g174) & (!g198) & (g664) & (!g665) & (g687) & (g700)) + ((!g174) & (!g198) & (g664) & (g665) & (!g687) & (!g700)) + ((!g174) & (!g198) & (g664) & (g665) & (!g687) & (g700)) + ((!g174) & (!g198) & (g664) & (g665) & (g687) & (g700)) + ((!g174) & (g198) & (!g664) & (!g665) & (g687) & (!g700)) + ((!g174) & (g198) & (!g664) & (g665) & (!g687) & (!g700)) + ((!g174) & (g198) & (!g664) & (g665) & (g687) & (!g700)) + ((!g174) & (g198) & (g664) & (!g665) & (!g687) & (!g700)) + ((!g174) & (g198) & (g664) & (!g665) & (!g687) & (g700)) + ((!g174) & (g198) & (g664) & (!g665) & (g687) & (g700)) + ((!g174) & (g198) & (g664) & (g665) & (!g687) & (g700)) + ((!g174) & (g198) & (g664) & (g665) & (g687) & (g700)) + ((g174) & (!g198) & (!g664) & (!g665) & (!g687) & (!g700)) + ((g174) & (!g198) & (!g664) & (!g665) & (g687) & (!g700)) + ((g174) & (!g198) & (!g664) & (g665) & (!g687) & (!g700)) + ((g174) & (!g198) & (g664) & (!g665) & (!g687) & (g700)) + ((g174) & (!g198) & (g664) & (!g665) & (g687) & (g700)) + ((g174) & (!g198) & (g664) & (g665) & (!g687) & (g700)) + ((g174) & (!g198) & (g664) & (g665) & (g687) & (!g700)) + ((g174) & (!g198) & (g664) & (g665) & (g687) & (g700)) + ((g174) & (g198) & (!g664) & (!g665) & (!g687) & (!g700)) + ((g174) & (g198) & (g664) & (!g665) & (!g687) & (g700)) + ((g174) & (g198) & (g664) & (!g665) & (g687) & (!g700)) + ((g174) & (g198) & (g664) & (!g665) & (g687) & (g700)) + ((g174) & (g198) & (g664) & (g665) & (!g687) & (!g700)) + ((g174) & (g198) & (g664) & (g665) & (!g687) & (g700)) + ((g174) & (g198) & (g664) & (g665) & (g687) & (!g700)) + ((g174) & (g198) & (g664) & (g665) & (g687) & (g700)));
	assign g714 = (((!g198) & (!g665) & (g687) & (!g700)) + ((!g198) & (g665) & (!g687) & (!g700)) + ((!g198) & (g665) & (!g687) & (g700)) + ((!g198) & (g665) & (g687) & (g700)) + ((g198) & (!g665) & (!g687) & (!g700)) + ((g198) & (g665) & (!g687) & (g700)) + ((g198) & (g665) & (g687) & (!g700)) + ((g198) & (g665) & (g687) & (g700)));
	assign g715 = (((!g229) & (!g255) & (!g667) & (g668) & (g686) & (!g700)) + ((!g229) & (!g255) & (g667) & (!g668) & (!g686) & (!g700)) + ((!g229) & (!g255) & (g667) & (!g668) & (!g686) & (g700)) + ((!g229) & (!g255) & (g667) & (!g668) & (g686) & (!g700)) + ((!g229) & (!g255) & (g667) & (!g668) & (g686) & (g700)) + ((!g229) & (!g255) & (g667) & (g668) & (!g686) & (!g700)) + ((!g229) & (!g255) & (g667) & (g668) & (!g686) & (g700)) + ((!g229) & (!g255) & (g667) & (g668) & (g686) & (g700)) + ((!g229) & (g255) & (!g667) & (!g668) & (g686) & (!g700)) + ((!g229) & (g255) & (!g667) & (g668) & (!g686) & (!g700)) + ((!g229) & (g255) & (!g667) & (g668) & (g686) & (!g700)) + ((!g229) & (g255) & (g667) & (!g668) & (!g686) & (!g700)) + ((!g229) & (g255) & (g667) & (!g668) & (!g686) & (g700)) + ((!g229) & (g255) & (g667) & (!g668) & (g686) & (g700)) + ((!g229) & (g255) & (g667) & (g668) & (!g686) & (g700)) + ((!g229) & (g255) & (g667) & (g668) & (g686) & (g700)) + ((g229) & (!g255) & (!g667) & (!g668) & (!g686) & (!g700)) + ((g229) & (!g255) & (!g667) & (!g668) & (g686) & (!g700)) + ((g229) & (!g255) & (!g667) & (g668) & (!g686) & (!g700)) + ((g229) & (!g255) & (g667) & (!g668) & (!g686) & (g700)) + ((g229) & (!g255) & (g667) & (!g668) & (g686) & (g700)) + ((g229) & (!g255) & (g667) & (g668) & (!g686) & (g700)) + ((g229) & (!g255) & (g667) & (g668) & (g686) & (!g700)) + ((g229) & (!g255) & (g667) & (g668) & (g686) & (g700)) + ((g229) & (g255) & (!g667) & (!g668) & (!g686) & (!g700)) + ((g229) & (g255) & (g667) & (!g668) & (!g686) & (g700)) + ((g229) & (g255) & (g667) & (!g668) & (g686) & (!g700)) + ((g229) & (g255) & (g667) & (!g668) & (g686) & (g700)) + ((g229) & (g255) & (g667) & (g668) & (!g686) & (!g700)) + ((g229) & (g255) & (g667) & (g668) & (!g686) & (g700)) + ((g229) & (g255) & (g667) & (g668) & (g686) & (!g700)) + ((g229) & (g255) & (g667) & (g668) & (g686) & (g700)));
	assign g716 = (((!g255) & (!g668) & (g686) & (!g700)) + ((!g255) & (g668) & (!g686) & (!g700)) + ((!g255) & (g668) & (!g686) & (g700)) + ((!g255) & (g668) & (g686) & (g700)) + ((g255) & (!g668) & (!g686) & (!g700)) + ((g255) & (g668) & (!g686) & (g700)) + ((g255) & (g668) & (g686) & (!g700)) + ((g255) & (g668) & (g686) & (g700)));
	assign g717 = (((!g290) & (!g319) & (!g670) & (g671) & (g685) & (!g700)) + ((!g290) & (!g319) & (g670) & (!g671) & (!g685) & (!g700)) + ((!g290) & (!g319) & (g670) & (!g671) & (!g685) & (g700)) + ((!g290) & (!g319) & (g670) & (!g671) & (g685) & (!g700)) + ((!g290) & (!g319) & (g670) & (!g671) & (g685) & (g700)) + ((!g290) & (!g319) & (g670) & (g671) & (!g685) & (!g700)) + ((!g290) & (!g319) & (g670) & (g671) & (!g685) & (g700)) + ((!g290) & (!g319) & (g670) & (g671) & (g685) & (g700)) + ((!g290) & (g319) & (!g670) & (!g671) & (g685) & (!g700)) + ((!g290) & (g319) & (!g670) & (g671) & (!g685) & (!g700)) + ((!g290) & (g319) & (!g670) & (g671) & (g685) & (!g700)) + ((!g290) & (g319) & (g670) & (!g671) & (!g685) & (!g700)) + ((!g290) & (g319) & (g670) & (!g671) & (!g685) & (g700)) + ((!g290) & (g319) & (g670) & (!g671) & (g685) & (g700)) + ((!g290) & (g319) & (g670) & (g671) & (!g685) & (g700)) + ((!g290) & (g319) & (g670) & (g671) & (g685) & (g700)) + ((g290) & (!g319) & (!g670) & (!g671) & (!g685) & (!g700)) + ((g290) & (!g319) & (!g670) & (!g671) & (g685) & (!g700)) + ((g290) & (!g319) & (!g670) & (g671) & (!g685) & (!g700)) + ((g290) & (!g319) & (g670) & (!g671) & (!g685) & (g700)) + ((g290) & (!g319) & (g670) & (!g671) & (g685) & (g700)) + ((g290) & (!g319) & (g670) & (g671) & (!g685) & (g700)) + ((g290) & (!g319) & (g670) & (g671) & (g685) & (!g700)) + ((g290) & (!g319) & (g670) & (g671) & (g685) & (g700)) + ((g290) & (g319) & (!g670) & (!g671) & (!g685) & (!g700)) + ((g290) & (g319) & (g670) & (!g671) & (!g685) & (g700)) + ((g290) & (g319) & (g670) & (!g671) & (g685) & (!g700)) + ((g290) & (g319) & (g670) & (!g671) & (g685) & (g700)) + ((g290) & (g319) & (g670) & (g671) & (!g685) & (!g700)) + ((g290) & (g319) & (g670) & (g671) & (!g685) & (g700)) + ((g290) & (g319) & (g670) & (g671) & (g685) & (!g700)) + ((g290) & (g319) & (g670) & (g671) & (g685) & (g700)));
	assign g718 = (((!g319) & (!g671) & (g685) & (!g700)) + ((!g319) & (g671) & (!g685) & (!g700)) + ((!g319) & (g671) & (!g685) & (g700)) + ((!g319) & (g671) & (g685) & (g700)) + ((g319) & (!g671) & (!g685) & (!g700)) + ((g319) & (g671) & (!g685) & (g700)) + ((g319) & (g671) & (g685) & (!g700)) + ((g319) & (g671) & (g685) & (g700)));
	assign g719 = (((!g358) & (!g390) & (!g673) & (g674) & (g684) & (!g700)) + ((!g358) & (!g390) & (g673) & (!g674) & (!g684) & (!g700)) + ((!g358) & (!g390) & (g673) & (!g674) & (!g684) & (g700)) + ((!g358) & (!g390) & (g673) & (!g674) & (g684) & (!g700)) + ((!g358) & (!g390) & (g673) & (!g674) & (g684) & (g700)) + ((!g358) & (!g390) & (g673) & (g674) & (!g684) & (!g700)) + ((!g358) & (!g390) & (g673) & (g674) & (!g684) & (g700)) + ((!g358) & (!g390) & (g673) & (g674) & (g684) & (g700)) + ((!g358) & (g390) & (!g673) & (!g674) & (g684) & (!g700)) + ((!g358) & (g390) & (!g673) & (g674) & (!g684) & (!g700)) + ((!g358) & (g390) & (!g673) & (g674) & (g684) & (!g700)) + ((!g358) & (g390) & (g673) & (!g674) & (!g684) & (!g700)) + ((!g358) & (g390) & (g673) & (!g674) & (!g684) & (g700)) + ((!g358) & (g390) & (g673) & (!g674) & (g684) & (g700)) + ((!g358) & (g390) & (g673) & (g674) & (!g684) & (g700)) + ((!g358) & (g390) & (g673) & (g674) & (g684) & (g700)) + ((g358) & (!g390) & (!g673) & (!g674) & (!g684) & (!g700)) + ((g358) & (!g390) & (!g673) & (!g674) & (g684) & (!g700)) + ((g358) & (!g390) & (!g673) & (g674) & (!g684) & (!g700)) + ((g358) & (!g390) & (g673) & (!g674) & (!g684) & (g700)) + ((g358) & (!g390) & (g673) & (!g674) & (g684) & (g700)) + ((g358) & (!g390) & (g673) & (g674) & (!g684) & (g700)) + ((g358) & (!g390) & (g673) & (g674) & (g684) & (!g700)) + ((g358) & (!g390) & (g673) & (g674) & (g684) & (g700)) + ((g358) & (g390) & (!g673) & (!g674) & (!g684) & (!g700)) + ((g358) & (g390) & (g673) & (!g674) & (!g684) & (g700)) + ((g358) & (g390) & (g673) & (!g674) & (g684) & (!g700)) + ((g358) & (g390) & (g673) & (!g674) & (g684) & (g700)) + ((g358) & (g390) & (g673) & (g674) & (!g684) & (!g700)) + ((g358) & (g390) & (g673) & (g674) & (!g684) & (g700)) + ((g358) & (g390) & (g673) & (g674) & (g684) & (!g700)) + ((g358) & (g390) & (g673) & (g674) & (g684) & (g700)));
	assign g720 = (((!g390) & (!g674) & (g684) & (!g700)) + ((!g390) & (g674) & (!g684) & (!g700)) + ((!g390) & (g674) & (!g684) & (g700)) + ((!g390) & (g674) & (g684) & (g700)) + ((g390) & (!g674) & (!g684) & (!g700)) + ((g390) & (g674) & (!g684) & (g700)) + ((g390) & (g674) & (g684) & (!g700)) + ((g390) & (g674) & (g684) & (g700)));
	assign g721 = (((!g433) & (!g468) & (!g676) & (g677) & (g683) & (!g700)) + ((!g433) & (!g468) & (g676) & (!g677) & (!g683) & (!g700)) + ((!g433) & (!g468) & (g676) & (!g677) & (!g683) & (g700)) + ((!g433) & (!g468) & (g676) & (!g677) & (g683) & (!g700)) + ((!g433) & (!g468) & (g676) & (!g677) & (g683) & (g700)) + ((!g433) & (!g468) & (g676) & (g677) & (!g683) & (!g700)) + ((!g433) & (!g468) & (g676) & (g677) & (!g683) & (g700)) + ((!g433) & (!g468) & (g676) & (g677) & (g683) & (g700)) + ((!g433) & (g468) & (!g676) & (!g677) & (g683) & (!g700)) + ((!g433) & (g468) & (!g676) & (g677) & (!g683) & (!g700)) + ((!g433) & (g468) & (!g676) & (g677) & (g683) & (!g700)) + ((!g433) & (g468) & (g676) & (!g677) & (!g683) & (!g700)) + ((!g433) & (g468) & (g676) & (!g677) & (!g683) & (g700)) + ((!g433) & (g468) & (g676) & (!g677) & (g683) & (g700)) + ((!g433) & (g468) & (g676) & (g677) & (!g683) & (g700)) + ((!g433) & (g468) & (g676) & (g677) & (g683) & (g700)) + ((g433) & (!g468) & (!g676) & (!g677) & (!g683) & (!g700)) + ((g433) & (!g468) & (!g676) & (!g677) & (g683) & (!g700)) + ((g433) & (!g468) & (!g676) & (g677) & (!g683) & (!g700)) + ((g433) & (!g468) & (g676) & (!g677) & (!g683) & (g700)) + ((g433) & (!g468) & (g676) & (!g677) & (g683) & (g700)) + ((g433) & (!g468) & (g676) & (g677) & (!g683) & (g700)) + ((g433) & (!g468) & (g676) & (g677) & (g683) & (!g700)) + ((g433) & (!g468) & (g676) & (g677) & (g683) & (g700)) + ((g433) & (g468) & (!g676) & (!g677) & (!g683) & (!g700)) + ((g433) & (g468) & (g676) & (!g677) & (!g683) & (g700)) + ((g433) & (g468) & (g676) & (!g677) & (g683) & (!g700)) + ((g433) & (g468) & (g676) & (!g677) & (g683) & (g700)) + ((g433) & (g468) & (g676) & (g677) & (!g683) & (!g700)) + ((g433) & (g468) & (g676) & (g677) & (!g683) & (g700)) + ((g433) & (g468) & (g676) & (g677) & (g683) & (!g700)) + ((g433) & (g468) & (g676) & (g677) & (g683) & (g700)));
	assign g722 = (((!g468) & (!g677) & (g683) & (!g700)) + ((!g468) & (g677) & (!g683) & (!g700)) + ((!g468) & (g677) & (!g683) & (g700)) + ((!g468) & (g677) & (g683) & (g700)) + ((g468) & (!g677) & (!g683) & (!g700)) + ((g468) & (g677) & (!g683) & (g700)) + ((g468) & (g677) & (g683) & (!g700)) + ((g468) & (g677) & (g683) & (g700)));
	assign g723 = (((!g515) & (!g553) & (!g679) & (g680) & (g682) & (!g700)) + ((!g515) & (!g553) & (g679) & (!g680) & (!g682) & (!g700)) + ((!g515) & (!g553) & (g679) & (!g680) & (!g682) & (g700)) + ((!g515) & (!g553) & (g679) & (!g680) & (g682) & (!g700)) + ((!g515) & (!g553) & (g679) & (!g680) & (g682) & (g700)) + ((!g515) & (!g553) & (g679) & (g680) & (!g682) & (!g700)) + ((!g515) & (!g553) & (g679) & (g680) & (!g682) & (g700)) + ((!g515) & (!g553) & (g679) & (g680) & (g682) & (g700)) + ((!g515) & (g553) & (!g679) & (!g680) & (g682) & (!g700)) + ((!g515) & (g553) & (!g679) & (g680) & (!g682) & (!g700)) + ((!g515) & (g553) & (!g679) & (g680) & (g682) & (!g700)) + ((!g515) & (g553) & (g679) & (!g680) & (!g682) & (!g700)) + ((!g515) & (g553) & (g679) & (!g680) & (!g682) & (g700)) + ((!g515) & (g553) & (g679) & (!g680) & (g682) & (g700)) + ((!g515) & (g553) & (g679) & (g680) & (!g682) & (g700)) + ((!g515) & (g553) & (g679) & (g680) & (g682) & (g700)) + ((g515) & (!g553) & (!g679) & (!g680) & (!g682) & (!g700)) + ((g515) & (!g553) & (!g679) & (!g680) & (g682) & (!g700)) + ((g515) & (!g553) & (!g679) & (g680) & (!g682) & (!g700)) + ((g515) & (!g553) & (g679) & (!g680) & (!g682) & (g700)) + ((g515) & (!g553) & (g679) & (!g680) & (g682) & (g700)) + ((g515) & (!g553) & (g679) & (g680) & (!g682) & (g700)) + ((g515) & (!g553) & (g679) & (g680) & (g682) & (!g700)) + ((g515) & (!g553) & (g679) & (g680) & (g682) & (g700)) + ((g515) & (g553) & (!g679) & (!g680) & (!g682) & (!g700)) + ((g515) & (g553) & (g679) & (!g680) & (!g682) & (g700)) + ((g515) & (g553) & (g679) & (!g680) & (g682) & (!g700)) + ((g515) & (g553) & (g679) & (!g680) & (g682) & (g700)) + ((g515) & (g553) & (g679) & (g680) & (!g682) & (!g700)) + ((g515) & (g553) & (g679) & (g680) & (!g682) & (g700)) + ((g515) & (g553) & (g679) & (g680) & (g682) & (!g700)) + ((g515) & (g553) & (g679) & (g680) & (g682) & (g700)));
	assign g724 = (((!g553) & (!g680) & (g682) & (!g700)) + ((!g553) & (g680) & (!g682) & (!g700)) + ((!g553) & (g680) & (!g682) & (g700)) + ((!g553) & (g680) & (g682) & (g700)) + ((g553) & (!g680) & (!g682) & (!g700)) + ((g553) & (g680) & (!g682) & (g700)) + ((g553) & (g680) & (g682) & (!g700)) + ((g553) & (g680) & (g682) & (g700)));
	assign g725 = (((!g604) & (!ax74x) & (!ax75x) & (!g645) & (!g681) & (g700)) + ((!g604) & (!ax74x) & (!ax75x) & (!g645) & (g681) & (!g700)) + ((!g604) & (!ax74x) & (!ax75x) & (!g645) & (g681) & (g700)) + ((!g604) & (!ax74x) & (!ax75x) & (g645) & (!g681) & (!g700)) + ((!g604) & (!ax74x) & (ax75x) & (!g645) & (!g681) & (!g700)) + ((!g604) & (!ax74x) & (ax75x) & (g645) & (!g681) & (g700)) + ((!g604) & (!ax74x) & (ax75x) & (g645) & (g681) & (!g700)) + ((!g604) & (!ax74x) & (ax75x) & (g645) & (g681) & (g700)) + ((!g604) & (ax74x) & (!ax75x) & (g645) & (!g681) & (!g700)) + ((!g604) & (ax74x) & (!ax75x) & (g645) & (g681) & (!g700)) + ((!g604) & (ax74x) & (ax75x) & (!g645) & (!g681) & (!g700)) + ((!g604) & (ax74x) & (ax75x) & (!g645) & (!g681) & (g700)) + ((!g604) & (ax74x) & (ax75x) & (!g645) & (g681) & (!g700)) + ((!g604) & (ax74x) & (ax75x) & (!g645) & (g681) & (g700)) + ((!g604) & (ax74x) & (ax75x) & (g645) & (!g681) & (g700)) + ((!g604) & (ax74x) & (ax75x) & (g645) & (g681) & (g700)) + ((g604) & (!ax74x) & (!ax75x) & (!g645) & (!g681) & (!g700)) + ((g604) & (!ax74x) & (!ax75x) & (!g645) & (!g681) & (g700)) + ((g604) & (!ax74x) & (!ax75x) & (!g645) & (g681) & (g700)) + ((g604) & (!ax74x) & (!ax75x) & (g645) & (g681) & (!g700)) + ((g604) & (!ax74x) & (ax75x) & (!g645) & (g681) & (!g700)) + ((g604) & (!ax74x) & (ax75x) & (g645) & (!g681) & (!g700)) + ((g604) & (!ax74x) & (ax75x) & (g645) & (!g681) & (g700)) + ((g604) & (!ax74x) & (ax75x) & (g645) & (g681) & (g700)) + ((g604) & (ax74x) & (!ax75x) & (!g645) & (!g681) & (!g700)) + ((g604) & (ax74x) & (!ax75x) & (!g645) & (g681) & (!g700)) + ((g604) & (ax74x) & (ax75x) & (!g645) & (!g681) & (g700)) + ((g604) & (ax74x) & (ax75x) & (!g645) & (g681) & (g700)) + ((g604) & (ax74x) & (ax75x) & (g645) & (!g681) & (!g700)) + ((g604) & (ax74x) & (ax75x) & (g645) & (!g681) & (g700)) + ((g604) & (ax74x) & (ax75x) & (g645) & (g681) & (!g700)) + ((g604) & (ax74x) & (ax75x) & (g645) & (g681) & (g700)));
	assign g726 = (((!ax74x) & (!g645) & (!g681) & (g700)) + ((!ax74x) & (!g645) & (g681) & (!g700)) + ((!ax74x) & (!g645) & (g681) & (g700)) + ((!ax74x) & (g645) & (g681) & (!g700)) + ((ax74x) & (!g645) & (!g681) & (!g700)) + ((ax74x) & (g645) & (!g681) & (!g700)) + ((ax74x) & (g645) & (!g681) & (g700)) + ((ax74x) & (g645) & (g681) & (g700)));
	assign g727 = (((!ax70x) & (!ax71x)));
	assign g728 = (((!g645) & (!ax72x) & (!ax73x) & (!g700) & (!g727)) + ((!g645) & (!ax72x) & (ax73x) & (g700) & (!g727)) + ((!g645) & (ax72x) & (ax73x) & (g700) & (!g727)) + ((!g645) & (ax72x) & (ax73x) & (g700) & (g727)) + ((g645) & (!ax72x) & (!ax73x) & (!g700) & (!g727)) + ((g645) & (!ax72x) & (!ax73x) & (!g700) & (g727)) + ((g645) & (!ax72x) & (!ax73x) & (g700) & (!g727)) + ((g645) & (!ax72x) & (ax73x) & (!g700) & (!g727)) + ((g645) & (!ax72x) & (ax73x) & (g700) & (!g727)) + ((g645) & (!ax72x) & (ax73x) & (g700) & (g727)) + ((g645) & (ax72x) & (!ax73x) & (g700) & (!g727)) + ((g645) & (ax72x) & (!ax73x) & (g700) & (g727)) + ((g645) & (ax72x) & (ax73x) & (!g700) & (!g727)) + ((g645) & (ax72x) & (ax73x) & (!g700) & (g727)) + ((g645) & (ax72x) & (ax73x) & (g700) & (!g727)) + ((g645) & (ax72x) & (ax73x) & (g700) & (g727)));
	assign g729 = (((!g553) & (!g604) & (g725) & (g726) & (g728)) + ((!g553) & (g604) & (g725) & (!g726) & (g728)) + ((!g553) & (g604) & (g725) & (g726) & (!g728)) + ((!g553) & (g604) & (g725) & (g726) & (g728)) + ((g553) & (!g604) & (!g725) & (g726) & (g728)) + ((g553) & (!g604) & (g725) & (!g726) & (!g728)) + ((g553) & (!g604) & (g725) & (!g726) & (g728)) + ((g553) & (!g604) & (g725) & (g726) & (!g728)) + ((g553) & (!g604) & (g725) & (g726) & (g728)) + ((g553) & (g604) & (!g725) & (!g726) & (g728)) + ((g553) & (g604) & (!g725) & (g726) & (!g728)) + ((g553) & (g604) & (!g725) & (g726) & (g728)) + ((g553) & (g604) & (g725) & (!g726) & (!g728)) + ((g553) & (g604) & (g725) & (!g726) & (g728)) + ((g553) & (g604) & (g725) & (g726) & (!g728)) + ((g553) & (g604) & (g725) & (g726) & (g728)));
	assign g730 = (((!g468) & (!g515) & (g723) & (g724) & (g729)) + ((!g468) & (g515) & (g723) & (!g724) & (g729)) + ((!g468) & (g515) & (g723) & (g724) & (!g729)) + ((!g468) & (g515) & (g723) & (g724) & (g729)) + ((g468) & (!g515) & (!g723) & (g724) & (g729)) + ((g468) & (!g515) & (g723) & (!g724) & (!g729)) + ((g468) & (!g515) & (g723) & (!g724) & (g729)) + ((g468) & (!g515) & (g723) & (g724) & (!g729)) + ((g468) & (!g515) & (g723) & (g724) & (g729)) + ((g468) & (g515) & (!g723) & (!g724) & (g729)) + ((g468) & (g515) & (!g723) & (g724) & (!g729)) + ((g468) & (g515) & (!g723) & (g724) & (g729)) + ((g468) & (g515) & (g723) & (!g724) & (!g729)) + ((g468) & (g515) & (g723) & (!g724) & (g729)) + ((g468) & (g515) & (g723) & (g724) & (!g729)) + ((g468) & (g515) & (g723) & (g724) & (g729)));
	assign g731 = (((!g390) & (!g433) & (g721) & (g722) & (g730)) + ((!g390) & (g433) & (g721) & (!g722) & (g730)) + ((!g390) & (g433) & (g721) & (g722) & (!g730)) + ((!g390) & (g433) & (g721) & (g722) & (g730)) + ((g390) & (!g433) & (!g721) & (g722) & (g730)) + ((g390) & (!g433) & (g721) & (!g722) & (!g730)) + ((g390) & (!g433) & (g721) & (!g722) & (g730)) + ((g390) & (!g433) & (g721) & (g722) & (!g730)) + ((g390) & (!g433) & (g721) & (g722) & (g730)) + ((g390) & (g433) & (!g721) & (!g722) & (g730)) + ((g390) & (g433) & (!g721) & (g722) & (!g730)) + ((g390) & (g433) & (!g721) & (g722) & (g730)) + ((g390) & (g433) & (g721) & (!g722) & (!g730)) + ((g390) & (g433) & (g721) & (!g722) & (g730)) + ((g390) & (g433) & (g721) & (g722) & (!g730)) + ((g390) & (g433) & (g721) & (g722) & (g730)));
	assign g732 = (((!g319) & (!g358) & (g719) & (g720) & (g731)) + ((!g319) & (g358) & (g719) & (!g720) & (g731)) + ((!g319) & (g358) & (g719) & (g720) & (!g731)) + ((!g319) & (g358) & (g719) & (g720) & (g731)) + ((g319) & (!g358) & (!g719) & (g720) & (g731)) + ((g319) & (!g358) & (g719) & (!g720) & (!g731)) + ((g319) & (!g358) & (g719) & (!g720) & (g731)) + ((g319) & (!g358) & (g719) & (g720) & (!g731)) + ((g319) & (!g358) & (g719) & (g720) & (g731)) + ((g319) & (g358) & (!g719) & (!g720) & (g731)) + ((g319) & (g358) & (!g719) & (g720) & (!g731)) + ((g319) & (g358) & (!g719) & (g720) & (g731)) + ((g319) & (g358) & (g719) & (!g720) & (!g731)) + ((g319) & (g358) & (g719) & (!g720) & (g731)) + ((g319) & (g358) & (g719) & (g720) & (!g731)) + ((g319) & (g358) & (g719) & (g720) & (g731)));
	assign g733 = (((!g255) & (!g290) & (g717) & (g718) & (g732)) + ((!g255) & (g290) & (g717) & (!g718) & (g732)) + ((!g255) & (g290) & (g717) & (g718) & (!g732)) + ((!g255) & (g290) & (g717) & (g718) & (g732)) + ((g255) & (!g290) & (!g717) & (g718) & (g732)) + ((g255) & (!g290) & (g717) & (!g718) & (!g732)) + ((g255) & (!g290) & (g717) & (!g718) & (g732)) + ((g255) & (!g290) & (g717) & (g718) & (!g732)) + ((g255) & (!g290) & (g717) & (g718) & (g732)) + ((g255) & (g290) & (!g717) & (!g718) & (g732)) + ((g255) & (g290) & (!g717) & (g718) & (!g732)) + ((g255) & (g290) & (!g717) & (g718) & (g732)) + ((g255) & (g290) & (g717) & (!g718) & (!g732)) + ((g255) & (g290) & (g717) & (!g718) & (g732)) + ((g255) & (g290) & (g717) & (g718) & (!g732)) + ((g255) & (g290) & (g717) & (g718) & (g732)));
	assign g734 = (((!g198) & (!g229) & (g715) & (g716) & (g733)) + ((!g198) & (g229) & (g715) & (!g716) & (g733)) + ((!g198) & (g229) & (g715) & (g716) & (!g733)) + ((!g198) & (g229) & (g715) & (g716) & (g733)) + ((g198) & (!g229) & (!g715) & (g716) & (g733)) + ((g198) & (!g229) & (g715) & (!g716) & (!g733)) + ((g198) & (!g229) & (g715) & (!g716) & (g733)) + ((g198) & (!g229) & (g715) & (g716) & (!g733)) + ((g198) & (!g229) & (g715) & (g716) & (g733)) + ((g198) & (g229) & (!g715) & (!g716) & (g733)) + ((g198) & (g229) & (!g715) & (g716) & (!g733)) + ((g198) & (g229) & (!g715) & (g716) & (g733)) + ((g198) & (g229) & (g715) & (!g716) & (!g733)) + ((g198) & (g229) & (g715) & (!g716) & (g733)) + ((g198) & (g229) & (g715) & (g716) & (!g733)) + ((g198) & (g229) & (g715) & (g716) & (g733)));
	assign g735 = (((!g147) & (!g174) & (g713) & (g714) & (g734)) + ((!g147) & (g174) & (g713) & (!g714) & (g734)) + ((!g147) & (g174) & (g713) & (g714) & (!g734)) + ((!g147) & (g174) & (g713) & (g714) & (g734)) + ((g147) & (!g174) & (!g713) & (g714) & (g734)) + ((g147) & (!g174) & (g713) & (!g714) & (!g734)) + ((g147) & (!g174) & (g713) & (!g714) & (g734)) + ((g147) & (!g174) & (g713) & (g714) & (!g734)) + ((g147) & (!g174) & (g713) & (g714) & (g734)) + ((g147) & (g174) & (!g713) & (!g714) & (g734)) + ((g147) & (g174) & (!g713) & (g714) & (!g734)) + ((g147) & (g174) & (!g713) & (g714) & (g734)) + ((g147) & (g174) & (g713) & (!g714) & (!g734)) + ((g147) & (g174) & (g713) & (!g714) & (g734)) + ((g147) & (g174) & (g713) & (g714) & (!g734)) + ((g147) & (g174) & (g713) & (g714) & (g734)));
	assign g736 = (((!g104) & (!g127) & (g711) & (g712) & (g735)) + ((!g104) & (g127) & (g711) & (!g712) & (g735)) + ((!g104) & (g127) & (g711) & (g712) & (!g735)) + ((!g104) & (g127) & (g711) & (g712) & (g735)) + ((g104) & (!g127) & (!g711) & (g712) & (g735)) + ((g104) & (!g127) & (g711) & (!g712) & (!g735)) + ((g104) & (!g127) & (g711) & (!g712) & (g735)) + ((g104) & (!g127) & (g711) & (g712) & (!g735)) + ((g104) & (!g127) & (g711) & (g712) & (g735)) + ((g104) & (g127) & (!g711) & (!g712) & (g735)) + ((g104) & (g127) & (!g711) & (g712) & (!g735)) + ((g104) & (g127) & (!g711) & (g712) & (g735)) + ((g104) & (g127) & (g711) & (!g712) & (!g735)) + ((g104) & (g127) & (g711) & (!g712) & (g735)) + ((g104) & (g127) & (g711) & (g712) & (!g735)) + ((g104) & (g127) & (g711) & (g712) & (g735)));
	assign g737 = (((!g68) & (!g87) & (g709) & (g710) & (g736)) + ((!g68) & (g87) & (g709) & (!g710) & (g736)) + ((!g68) & (g87) & (g709) & (g710) & (!g736)) + ((!g68) & (g87) & (g709) & (g710) & (g736)) + ((g68) & (!g87) & (!g709) & (g710) & (g736)) + ((g68) & (!g87) & (g709) & (!g710) & (!g736)) + ((g68) & (!g87) & (g709) & (!g710) & (g736)) + ((g68) & (!g87) & (g709) & (g710) & (!g736)) + ((g68) & (!g87) & (g709) & (g710) & (g736)) + ((g68) & (g87) & (!g709) & (!g710) & (g736)) + ((g68) & (g87) & (!g709) & (g710) & (!g736)) + ((g68) & (g87) & (!g709) & (g710) & (g736)) + ((g68) & (g87) & (g709) & (!g710) & (!g736)) + ((g68) & (g87) & (g709) & (!g710) & (g736)) + ((g68) & (g87) & (g709) & (g710) & (!g736)) + ((g68) & (g87) & (g709) & (g710) & (g736)));
	assign g738 = (((!g39) & (!g54) & (g707) & (g708) & (g737)) + ((!g39) & (g54) & (g707) & (!g708) & (g737)) + ((!g39) & (g54) & (g707) & (g708) & (!g737)) + ((!g39) & (g54) & (g707) & (g708) & (g737)) + ((g39) & (!g54) & (!g707) & (g708) & (g737)) + ((g39) & (!g54) & (g707) & (!g708) & (!g737)) + ((g39) & (!g54) & (g707) & (!g708) & (g737)) + ((g39) & (!g54) & (g707) & (g708) & (!g737)) + ((g39) & (!g54) & (g707) & (g708) & (g737)) + ((g39) & (g54) & (!g707) & (!g708) & (g737)) + ((g39) & (g54) & (!g707) & (g708) & (!g737)) + ((g39) & (g54) & (!g707) & (g708) & (g737)) + ((g39) & (g54) & (g707) & (!g708) & (!g737)) + ((g39) & (g54) & (g707) & (!g708) & (g737)) + ((g39) & (g54) & (g707) & (g708) & (!g737)) + ((g39) & (g54) & (g707) & (g708) & (g737)));
	assign g739 = (((!g18) & (!g27) & (g705) & (g706) & (g738)) + ((!g18) & (g27) & (g705) & (!g706) & (g738)) + ((!g18) & (g27) & (g705) & (g706) & (!g738)) + ((!g18) & (g27) & (g705) & (g706) & (g738)) + ((g18) & (!g27) & (!g705) & (g706) & (g738)) + ((g18) & (!g27) & (g705) & (!g706) & (!g738)) + ((g18) & (!g27) & (g705) & (!g706) & (g738)) + ((g18) & (!g27) & (g705) & (g706) & (!g738)) + ((g18) & (!g27) & (g705) & (g706) & (g738)) + ((g18) & (g27) & (!g705) & (!g706) & (g738)) + ((g18) & (g27) & (!g705) & (g706) & (!g738)) + ((g18) & (g27) & (!g705) & (g706) & (g738)) + ((g18) & (g27) & (g705) & (!g706) & (!g738)) + ((g18) & (g27) & (g705) & (!g706) & (g738)) + ((g18) & (g27) & (g705) & (g706) & (!g738)) + ((g18) & (g27) & (g705) & (g706) & (g738)));
	assign g740 = (((!g2) & (!g8) & (g703) & (g704) & (g739)) + ((!g2) & (g8) & (g703) & (!g704) & (g739)) + ((!g2) & (g8) & (g703) & (g704) & (!g739)) + ((!g2) & (g8) & (g703) & (g704) & (g739)) + ((g2) & (!g8) & (!g703) & (g704) & (g739)) + ((g2) & (!g8) & (g703) & (!g704) & (!g739)) + ((g2) & (!g8) & (g703) & (!g704) & (g739)) + ((g2) & (!g8) & (g703) & (g704) & (!g739)) + ((g2) & (!g8) & (g703) & (g704) & (g739)) + ((g2) & (g8) & (!g703) & (!g704) & (g739)) + ((g2) & (g8) & (!g703) & (g704) & (!g739)) + ((g2) & (g8) & (!g703) & (g704) & (g739)) + ((g2) & (g8) & (g703) & (!g704) & (!g739)) + ((g2) & (g8) & (g703) & (!g704) & (g739)) + ((g2) & (g8) & (g703) & (g704) & (!g739)) + ((g2) & (g8) & (g703) & (g704) & (g739)));
	assign g741 = (((!g2) & (!g647) & (g693) & (!g700)) + ((!g2) & (g647) & (!g693) & (!g700)) + ((!g2) & (g647) & (!g693) & (g700)) + ((!g2) & (g647) & (g693) & (g700)) + ((g2) & (!g647) & (!g693) & (!g700)) + ((g2) & (g647) & (!g693) & (g700)) + ((g2) & (g647) & (g693) & (!g700)) + ((g2) & (g647) & (g693) & (g700)));
	assign g742 = (((!g1) & (!g646) & (!g696) & (!g698) & (g699)) + ((!g1) & (!g646) & (!g696) & (g698) & (!g699)) + ((!g1) & (!g646) & (!g696) & (g698) & (g699)) + ((!g1) & (g646) & (g696) & (!g698) & (!g699)) + ((!g1) & (g646) & (g696) & (!g698) & (g699)) + ((!g1) & (g646) & (g696) & (g698) & (!g699)) + ((!g1) & (g646) & (g696) & (g698) & (g699)) + ((g1) & (!g646) & (!g696) & (!g698) & (g699)) + ((g1) & (!g646) & (!g696) & (g698) & (g699)) + ((g1) & (g646) & (g696) & (!g698) & (!g699)) + ((g1) & (g646) & (g696) & (!g698) & (g699)) + ((g1) & (g646) & (g696) & (g698) & (!g699)) + ((g1) & (g646) & (g696) & (g698) & (g699)));
	assign g743 = (((!g4) & (!g1) & (!g702) & (!g740) & (!g741) & (!g742)) + ((!g4) & (g1) & (!g702) & (!g740) & (!g741) & (!g742)) + ((!g4) & (g1) & (!g702) & (!g740) & (!g741) & (g742)) + ((!g4) & (g1) & (!g702) & (!g740) & (g741) & (!g742)) + ((!g4) & (g1) & (!g702) & (!g740) & (g741) & (g742)) + ((!g4) & (g1) & (!g702) & (g740) & (!g741) & (!g742)) + ((!g4) & (g1) & (!g702) & (g740) & (!g741) & (g742)) + ((!g4) & (g1) & (!g702) & (g740) & (g741) & (!g742)) + ((!g4) & (g1) & (!g702) & (g740) & (g741) & (g742)) + ((!g4) & (g1) & (g702) & (!g740) & (!g741) & (!g742)) + ((!g4) & (g1) & (g702) & (!g740) & (!g741) & (g742)) + ((g4) & (!g1) & (!g702) & (!g740) & (!g741) & (!g742)) + ((g4) & (!g1) & (!g702) & (!g740) & (g741) & (!g742)) + ((g4) & (!g1) & (!g702) & (g740) & (!g741) & (!g742)) + ((g4) & (g1) & (!g702) & (!g740) & (!g741) & (!g742)) + ((g4) & (g1) & (!g702) & (!g740) & (!g741) & (g742)) + ((g4) & (g1) & (!g702) & (!g740) & (g741) & (!g742)) + ((g4) & (g1) & (!g702) & (!g740) & (g741) & (g742)) + ((g4) & (g1) & (!g702) & (g740) & (!g741) & (!g742)) + ((g4) & (g1) & (!g702) & (g740) & (!g741) & (g742)) + ((g4) & (g1) & (!g702) & (g740) & (g741) & (!g742)) + ((g4) & (g1) & (!g702) & (g740) & (g741) & (g742)) + ((g4) & (g1) & (g702) & (!g740) & (!g741) & (!g742)) + ((g4) & (g1) & (g702) & (!g740) & (!g741) & (g742)) + ((g4) & (g1) & (g702) & (!g740) & (g741) & (!g742)) + ((g4) & (g1) & (g702) & (!g740) & (g741) & (g742)) + ((g4) & (g1) & (g702) & (g740) & (!g741) & (!g742)) + ((g4) & (g1) & (g702) & (g740) & (!g741) & (g742)));
	assign g744 = (((!g701) & (g743)));
	assign g745 = (((!g4) & (!g740) & (!g741) & (!g701) & (!g743)) + ((!g4) & (!g740) & (!g741) & (g701) & (!g743)) + ((!g4) & (!g740) & (!g741) & (g701) & (g743)) + ((!g4) & (!g740) & (g741) & (!g701) & (g743)) + ((!g4) & (g740) & (g741) & (!g701) & (!g743)) + ((!g4) & (g740) & (g741) & (!g701) & (g743)) + ((!g4) & (g740) & (g741) & (g701) & (!g743)) + ((!g4) & (g740) & (g741) & (g701) & (g743)) + ((g4) & (!g740) & (g741) & (!g701) & (!g743)) + ((g4) & (!g740) & (g741) & (!g701) & (g743)) + ((g4) & (!g740) & (g741) & (g701) & (!g743)) + ((g4) & (!g740) & (g741) & (g701) & (g743)) + ((g4) & (g740) & (!g741) & (!g701) & (!g743)) + ((g4) & (g740) & (!g741) & (g701) & (!g743)) + ((g4) & (g740) & (!g741) & (g701) & (g743)) + ((g4) & (g740) & (g741) & (!g701) & (g743)));
	assign g746 = (((!g2) & (!g8) & (g704) & (g739)) + ((!g2) & (g8) & (!g704) & (g739)) + ((!g2) & (g8) & (g704) & (!g739)) + ((!g2) & (g8) & (g704) & (g739)) + ((g2) & (!g8) & (!g704) & (!g739)) + ((g2) & (!g8) & (!g704) & (g739)) + ((g2) & (!g8) & (g704) & (!g739)) + ((g2) & (g8) & (!g704) & (!g739)));
	assign g747 = (((!g703) & (!g701) & (!g743) & (g746)) + ((!g703) & (g701) & (!g743) & (g746)) + ((!g703) & (g701) & (g743) & (g746)) + ((g703) & (!g701) & (!g743) & (!g746)) + ((g703) & (!g701) & (g743) & (!g746)) + ((g703) & (!g701) & (g743) & (g746)) + ((g703) & (g701) & (!g743) & (!g746)) + ((g703) & (g701) & (g743) & (!g746)));
	assign g748 = (((!g8) & (!g704) & (g739) & (!g701) & (!g743)) + ((!g8) & (!g704) & (g739) & (g701) & (!g743)) + ((!g8) & (!g704) & (g739) & (g701) & (g743)) + ((!g8) & (g704) & (!g739) & (!g701) & (!g743)) + ((!g8) & (g704) & (!g739) & (!g701) & (g743)) + ((!g8) & (g704) & (!g739) & (g701) & (!g743)) + ((!g8) & (g704) & (!g739) & (g701) & (g743)) + ((!g8) & (g704) & (g739) & (!g701) & (g743)) + ((g8) & (!g704) & (!g739) & (!g701) & (!g743)) + ((g8) & (!g704) & (!g739) & (g701) & (!g743)) + ((g8) & (!g704) & (!g739) & (g701) & (g743)) + ((g8) & (g704) & (!g739) & (!g701) & (g743)) + ((g8) & (g704) & (g739) & (!g701) & (!g743)) + ((g8) & (g704) & (g739) & (!g701) & (g743)) + ((g8) & (g704) & (g739) & (g701) & (!g743)) + ((g8) & (g704) & (g739) & (g701) & (g743)));
	assign g749 = (((!g18) & (!g27) & (g706) & (g738)) + ((!g18) & (g27) & (!g706) & (g738)) + ((!g18) & (g27) & (g706) & (!g738)) + ((!g18) & (g27) & (g706) & (g738)) + ((g18) & (!g27) & (!g706) & (!g738)) + ((g18) & (!g27) & (!g706) & (g738)) + ((g18) & (!g27) & (g706) & (!g738)) + ((g18) & (g27) & (!g706) & (!g738)));
	assign g750 = (((!g705) & (!g701) & (!g743) & (g749)) + ((!g705) & (g701) & (!g743) & (g749)) + ((!g705) & (g701) & (g743) & (g749)) + ((g705) & (!g701) & (!g743) & (!g749)) + ((g705) & (!g701) & (g743) & (!g749)) + ((g705) & (!g701) & (g743) & (g749)) + ((g705) & (g701) & (!g743) & (!g749)) + ((g705) & (g701) & (g743) & (!g749)));
	assign g751 = (((!g27) & (!g706) & (g738) & (!g701) & (!g743)) + ((!g27) & (!g706) & (g738) & (g701) & (!g743)) + ((!g27) & (!g706) & (g738) & (g701) & (g743)) + ((!g27) & (g706) & (!g738) & (!g701) & (!g743)) + ((!g27) & (g706) & (!g738) & (!g701) & (g743)) + ((!g27) & (g706) & (!g738) & (g701) & (!g743)) + ((!g27) & (g706) & (!g738) & (g701) & (g743)) + ((!g27) & (g706) & (g738) & (!g701) & (g743)) + ((g27) & (!g706) & (!g738) & (!g701) & (!g743)) + ((g27) & (!g706) & (!g738) & (g701) & (!g743)) + ((g27) & (!g706) & (!g738) & (g701) & (g743)) + ((g27) & (g706) & (!g738) & (!g701) & (g743)) + ((g27) & (g706) & (g738) & (!g701) & (!g743)) + ((g27) & (g706) & (g738) & (!g701) & (g743)) + ((g27) & (g706) & (g738) & (g701) & (!g743)) + ((g27) & (g706) & (g738) & (g701) & (g743)));
	assign g752 = (((!g39) & (!g54) & (g708) & (g737)) + ((!g39) & (g54) & (!g708) & (g737)) + ((!g39) & (g54) & (g708) & (!g737)) + ((!g39) & (g54) & (g708) & (g737)) + ((g39) & (!g54) & (!g708) & (!g737)) + ((g39) & (!g54) & (!g708) & (g737)) + ((g39) & (!g54) & (g708) & (!g737)) + ((g39) & (g54) & (!g708) & (!g737)));
	assign g753 = (((!g707) & (!g701) & (!g743) & (g752)) + ((!g707) & (g701) & (!g743) & (g752)) + ((!g707) & (g701) & (g743) & (g752)) + ((g707) & (!g701) & (!g743) & (!g752)) + ((g707) & (!g701) & (g743) & (!g752)) + ((g707) & (!g701) & (g743) & (g752)) + ((g707) & (g701) & (!g743) & (!g752)) + ((g707) & (g701) & (g743) & (!g752)));
	assign g754 = (((!g54) & (!g708) & (g737) & (!g701) & (!g743)) + ((!g54) & (!g708) & (g737) & (g701) & (!g743)) + ((!g54) & (!g708) & (g737) & (g701) & (g743)) + ((!g54) & (g708) & (!g737) & (!g701) & (!g743)) + ((!g54) & (g708) & (!g737) & (!g701) & (g743)) + ((!g54) & (g708) & (!g737) & (g701) & (!g743)) + ((!g54) & (g708) & (!g737) & (g701) & (g743)) + ((!g54) & (g708) & (g737) & (!g701) & (g743)) + ((g54) & (!g708) & (!g737) & (!g701) & (!g743)) + ((g54) & (!g708) & (!g737) & (g701) & (!g743)) + ((g54) & (!g708) & (!g737) & (g701) & (g743)) + ((g54) & (g708) & (!g737) & (!g701) & (g743)) + ((g54) & (g708) & (g737) & (!g701) & (!g743)) + ((g54) & (g708) & (g737) & (!g701) & (g743)) + ((g54) & (g708) & (g737) & (g701) & (!g743)) + ((g54) & (g708) & (g737) & (g701) & (g743)));
	assign g755 = (((!g68) & (!g87) & (g710) & (g736)) + ((!g68) & (g87) & (!g710) & (g736)) + ((!g68) & (g87) & (g710) & (!g736)) + ((!g68) & (g87) & (g710) & (g736)) + ((g68) & (!g87) & (!g710) & (!g736)) + ((g68) & (!g87) & (!g710) & (g736)) + ((g68) & (!g87) & (g710) & (!g736)) + ((g68) & (g87) & (!g710) & (!g736)));
	assign g756 = (((!g709) & (!g701) & (!g743) & (g755)) + ((!g709) & (g701) & (!g743) & (g755)) + ((!g709) & (g701) & (g743) & (g755)) + ((g709) & (!g701) & (!g743) & (!g755)) + ((g709) & (!g701) & (g743) & (!g755)) + ((g709) & (!g701) & (g743) & (g755)) + ((g709) & (g701) & (!g743) & (!g755)) + ((g709) & (g701) & (g743) & (!g755)));
	assign g757 = (((!g87) & (!g710) & (g736) & (!g701) & (!g743)) + ((!g87) & (!g710) & (g736) & (g701) & (!g743)) + ((!g87) & (!g710) & (g736) & (g701) & (g743)) + ((!g87) & (g710) & (!g736) & (!g701) & (!g743)) + ((!g87) & (g710) & (!g736) & (!g701) & (g743)) + ((!g87) & (g710) & (!g736) & (g701) & (!g743)) + ((!g87) & (g710) & (!g736) & (g701) & (g743)) + ((!g87) & (g710) & (g736) & (!g701) & (g743)) + ((g87) & (!g710) & (!g736) & (!g701) & (!g743)) + ((g87) & (!g710) & (!g736) & (g701) & (!g743)) + ((g87) & (!g710) & (!g736) & (g701) & (g743)) + ((g87) & (g710) & (!g736) & (!g701) & (g743)) + ((g87) & (g710) & (g736) & (!g701) & (!g743)) + ((g87) & (g710) & (g736) & (!g701) & (g743)) + ((g87) & (g710) & (g736) & (g701) & (!g743)) + ((g87) & (g710) & (g736) & (g701) & (g743)));
	assign g758 = (((!g104) & (!g127) & (g712) & (g735)) + ((!g104) & (g127) & (!g712) & (g735)) + ((!g104) & (g127) & (g712) & (!g735)) + ((!g104) & (g127) & (g712) & (g735)) + ((g104) & (!g127) & (!g712) & (!g735)) + ((g104) & (!g127) & (!g712) & (g735)) + ((g104) & (!g127) & (g712) & (!g735)) + ((g104) & (g127) & (!g712) & (!g735)));
	assign g759 = (((!g711) & (!g701) & (!g743) & (g758)) + ((!g711) & (g701) & (!g743) & (g758)) + ((!g711) & (g701) & (g743) & (g758)) + ((g711) & (!g701) & (!g743) & (!g758)) + ((g711) & (!g701) & (g743) & (!g758)) + ((g711) & (!g701) & (g743) & (g758)) + ((g711) & (g701) & (!g743) & (!g758)) + ((g711) & (g701) & (g743) & (!g758)));
	assign g760 = (((!g127) & (!g712) & (g735) & (!g701) & (!g743)) + ((!g127) & (!g712) & (g735) & (g701) & (!g743)) + ((!g127) & (!g712) & (g735) & (g701) & (g743)) + ((!g127) & (g712) & (!g735) & (!g701) & (!g743)) + ((!g127) & (g712) & (!g735) & (!g701) & (g743)) + ((!g127) & (g712) & (!g735) & (g701) & (!g743)) + ((!g127) & (g712) & (!g735) & (g701) & (g743)) + ((!g127) & (g712) & (g735) & (!g701) & (g743)) + ((g127) & (!g712) & (!g735) & (!g701) & (!g743)) + ((g127) & (!g712) & (!g735) & (g701) & (!g743)) + ((g127) & (!g712) & (!g735) & (g701) & (g743)) + ((g127) & (g712) & (!g735) & (!g701) & (g743)) + ((g127) & (g712) & (g735) & (!g701) & (!g743)) + ((g127) & (g712) & (g735) & (!g701) & (g743)) + ((g127) & (g712) & (g735) & (g701) & (!g743)) + ((g127) & (g712) & (g735) & (g701) & (g743)));
	assign g761 = (((!g147) & (!g174) & (g714) & (g734)) + ((!g147) & (g174) & (!g714) & (g734)) + ((!g147) & (g174) & (g714) & (!g734)) + ((!g147) & (g174) & (g714) & (g734)) + ((g147) & (!g174) & (!g714) & (!g734)) + ((g147) & (!g174) & (!g714) & (g734)) + ((g147) & (!g174) & (g714) & (!g734)) + ((g147) & (g174) & (!g714) & (!g734)));
	assign g762 = (((!g713) & (!g701) & (!g743) & (g761)) + ((!g713) & (g701) & (!g743) & (g761)) + ((!g713) & (g701) & (g743) & (g761)) + ((g713) & (!g701) & (!g743) & (!g761)) + ((g713) & (!g701) & (g743) & (!g761)) + ((g713) & (!g701) & (g743) & (g761)) + ((g713) & (g701) & (!g743) & (!g761)) + ((g713) & (g701) & (g743) & (!g761)));
	assign g763 = (((!g174) & (!g714) & (g734) & (!g701) & (!g743)) + ((!g174) & (!g714) & (g734) & (g701) & (!g743)) + ((!g174) & (!g714) & (g734) & (g701) & (g743)) + ((!g174) & (g714) & (!g734) & (!g701) & (!g743)) + ((!g174) & (g714) & (!g734) & (!g701) & (g743)) + ((!g174) & (g714) & (!g734) & (g701) & (!g743)) + ((!g174) & (g714) & (!g734) & (g701) & (g743)) + ((!g174) & (g714) & (g734) & (!g701) & (g743)) + ((g174) & (!g714) & (!g734) & (!g701) & (!g743)) + ((g174) & (!g714) & (!g734) & (g701) & (!g743)) + ((g174) & (!g714) & (!g734) & (g701) & (g743)) + ((g174) & (g714) & (!g734) & (!g701) & (g743)) + ((g174) & (g714) & (g734) & (!g701) & (!g743)) + ((g174) & (g714) & (g734) & (!g701) & (g743)) + ((g174) & (g714) & (g734) & (g701) & (!g743)) + ((g174) & (g714) & (g734) & (g701) & (g743)));
	assign g764 = (((!g198) & (!g229) & (g716) & (g733)) + ((!g198) & (g229) & (!g716) & (g733)) + ((!g198) & (g229) & (g716) & (!g733)) + ((!g198) & (g229) & (g716) & (g733)) + ((g198) & (!g229) & (!g716) & (!g733)) + ((g198) & (!g229) & (!g716) & (g733)) + ((g198) & (!g229) & (g716) & (!g733)) + ((g198) & (g229) & (!g716) & (!g733)));
	assign g765 = (((!g715) & (!g701) & (!g743) & (g764)) + ((!g715) & (g701) & (!g743) & (g764)) + ((!g715) & (g701) & (g743) & (g764)) + ((g715) & (!g701) & (!g743) & (!g764)) + ((g715) & (!g701) & (g743) & (!g764)) + ((g715) & (!g701) & (g743) & (g764)) + ((g715) & (g701) & (!g743) & (!g764)) + ((g715) & (g701) & (g743) & (!g764)));
	assign g766 = (((!g229) & (!g716) & (g733) & (!g701) & (!g743)) + ((!g229) & (!g716) & (g733) & (g701) & (!g743)) + ((!g229) & (!g716) & (g733) & (g701) & (g743)) + ((!g229) & (g716) & (!g733) & (!g701) & (!g743)) + ((!g229) & (g716) & (!g733) & (!g701) & (g743)) + ((!g229) & (g716) & (!g733) & (g701) & (!g743)) + ((!g229) & (g716) & (!g733) & (g701) & (g743)) + ((!g229) & (g716) & (g733) & (!g701) & (g743)) + ((g229) & (!g716) & (!g733) & (!g701) & (!g743)) + ((g229) & (!g716) & (!g733) & (g701) & (!g743)) + ((g229) & (!g716) & (!g733) & (g701) & (g743)) + ((g229) & (g716) & (!g733) & (!g701) & (g743)) + ((g229) & (g716) & (g733) & (!g701) & (!g743)) + ((g229) & (g716) & (g733) & (!g701) & (g743)) + ((g229) & (g716) & (g733) & (g701) & (!g743)) + ((g229) & (g716) & (g733) & (g701) & (g743)));
	assign g767 = (((!g255) & (!g290) & (g718) & (g732)) + ((!g255) & (g290) & (!g718) & (g732)) + ((!g255) & (g290) & (g718) & (!g732)) + ((!g255) & (g290) & (g718) & (g732)) + ((g255) & (!g290) & (!g718) & (!g732)) + ((g255) & (!g290) & (!g718) & (g732)) + ((g255) & (!g290) & (g718) & (!g732)) + ((g255) & (g290) & (!g718) & (!g732)));
	assign g768 = (((!g717) & (!g701) & (!g743) & (g767)) + ((!g717) & (g701) & (!g743) & (g767)) + ((!g717) & (g701) & (g743) & (g767)) + ((g717) & (!g701) & (!g743) & (!g767)) + ((g717) & (!g701) & (g743) & (!g767)) + ((g717) & (!g701) & (g743) & (g767)) + ((g717) & (g701) & (!g743) & (!g767)) + ((g717) & (g701) & (g743) & (!g767)));
	assign g769 = (((!g290) & (!g718) & (g732) & (!g701) & (!g743)) + ((!g290) & (!g718) & (g732) & (g701) & (!g743)) + ((!g290) & (!g718) & (g732) & (g701) & (g743)) + ((!g290) & (g718) & (!g732) & (!g701) & (!g743)) + ((!g290) & (g718) & (!g732) & (!g701) & (g743)) + ((!g290) & (g718) & (!g732) & (g701) & (!g743)) + ((!g290) & (g718) & (!g732) & (g701) & (g743)) + ((!g290) & (g718) & (g732) & (!g701) & (g743)) + ((g290) & (!g718) & (!g732) & (!g701) & (!g743)) + ((g290) & (!g718) & (!g732) & (g701) & (!g743)) + ((g290) & (!g718) & (!g732) & (g701) & (g743)) + ((g290) & (g718) & (!g732) & (!g701) & (g743)) + ((g290) & (g718) & (g732) & (!g701) & (!g743)) + ((g290) & (g718) & (g732) & (!g701) & (g743)) + ((g290) & (g718) & (g732) & (g701) & (!g743)) + ((g290) & (g718) & (g732) & (g701) & (g743)));
	assign g770 = (((!g319) & (!g358) & (g720) & (g731)) + ((!g319) & (g358) & (!g720) & (g731)) + ((!g319) & (g358) & (g720) & (!g731)) + ((!g319) & (g358) & (g720) & (g731)) + ((g319) & (!g358) & (!g720) & (!g731)) + ((g319) & (!g358) & (!g720) & (g731)) + ((g319) & (!g358) & (g720) & (!g731)) + ((g319) & (g358) & (!g720) & (!g731)));
	assign g771 = (((!g719) & (!g701) & (!g743) & (g770)) + ((!g719) & (g701) & (!g743) & (g770)) + ((!g719) & (g701) & (g743) & (g770)) + ((g719) & (!g701) & (!g743) & (!g770)) + ((g719) & (!g701) & (g743) & (!g770)) + ((g719) & (!g701) & (g743) & (g770)) + ((g719) & (g701) & (!g743) & (!g770)) + ((g719) & (g701) & (g743) & (!g770)));
	assign g772 = (((!g358) & (!g720) & (g731) & (!g701) & (!g743)) + ((!g358) & (!g720) & (g731) & (g701) & (!g743)) + ((!g358) & (!g720) & (g731) & (g701) & (g743)) + ((!g358) & (g720) & (!g731) & (!g701) & (!g743)) + ((!g358) & (g720) & (!g731) & (!g701) & (g743)) + ((!g358) & (g720) & (!g731) & (g701) & (!g743)) + ((!g358) & (g720) & (!g731) & (g701) & (g743)) + ((!g358) & (g720) & (g731) & (!g701) & (g743)) + ((g358) & (!g720) & (!g731) & (!g701) & (!g743)) + ((g358) & (!g720) & (!g731) & (g701) & (!g743)) + ((g358) & (!g720) & (!g731) & (g701) & (g743)) + ((g358) & (g720) & (!g731) & (!g701) & (g743)) + ((g358) & (g720) & (g731) & (!g701) & (!g743)) + ((g358) & (g720) & (g731) & (!g701) & (g743)) + ((g358) & (g720) & (g731) & (g701) & (!g743)) + ((g358) & (g720) & (g731) & (g701) & (g743)));
	assign g773 = (((!g390) & (!g433) & (g722) & (g730)) + ((!g390) & (g433) & (!g722) & (g730)) + ((!g390) & (g433) & (g722) & (!g730)) + ((!g390) & (g433) & (g722) & (g730)) + ((g390) & (!g433) & (!g722) & (!g730)) + ((g390) & (!g433) & (!g722) & (g730)) + ((g390) & (!g433) & (g722) & (!g730)) + ((g390) & (g433) & (!g722) & (!g730)));
	assign g774 = (((!g721) & (!g701) & (!g743) & (g773)) + ((!g721) & (g701) & (!g743) & (g773)) + ((!g721) & (g701) & (g743) & (g773)) + ((g721) & (!g701) & (!g743) & (!g773)) + ((g721) & (!g701) & (g743) & (!g773)) + ((g721) & (!g701) & (g743) & (g773)) + ((g721) & (g701) & (!g743) & (!g773)) + ((g721) & (g701) & (g743) & (!g773)));
	assign g775 = (((!g433) & (!g722) & (g730) & (!g701) & (!g743)) + ((!g433) & (!g722) & (g730) & (g701) & (!g743)) + ((!g433) & (!g722) & (g730) & (g701) & (g743)) + ((!g433) & (g722) & (!g730) & (!g701) & (!g743)) + ((!g433) & (g722) & (!g730) & (!g701) & (g743)) + ((!g433) & (g722) & (!g730) & (g701) & (!g743)) + ((!g433) & (g722) & (!g730) & (g701) & (g743)) + ((!g433) & (g722) & (g730) & (!g701) & (g743)) + ((g433) & (!g722) & (!g730) & (!g701) & (!g743)) + ((g433) & (!g722) & (!g730) & (g701) & (!g743)) + ((g433) & (!g722) & (!g730) & (g701) & (g743)) + ((g433) & (g722) & (!g730) & (!g701) & (g743)) + ((g433) & (g722) & (g730) & (!g701) & (!g743)) + ((g433) & (g722) & (g730) & (!g701) & (g743)) + ((g433) & (g722) & (g730) & (g701) & (!g743)) + ((g433) & (g722) & (g730) & (g701) & (g743)));
	assign g776 = (((!g468) & (!g515) & (g724) & (g729)) + ((!g468) & (g515) & (!g724) & (g729)) + ((!g468) & (g515) & (g724) & (!g729)) + ((!g468) & (g515) & (g724) & (g729)) + ((g468) & (!g515) & (!g724) & (!g729)) + ((g468) & (!g515) & (!g724) & (g729)) + ((g468) & (!g515) & (g724) & (!g729)) + ((g468) & (g515) & (!g724) & (!g729)));
	assign g777 = (((!g723) & (!g701) & (!g743) & (g776)) + ((!g723) & (g701) & (!g743) & (g776)) + ((!g723) & (g701) & (g743) & (g776)) + ((g723) & (!g701) & (!g743) & (!g776)) + ((g723) & (!g701) & (g743) & (!g776)) + ((g723) & (!g701) & (g743) & (g776)) + ((g723) & (g701) & (!g743) & (!g776)) + ((g723) & (g701) & (g743) & (!g776)));
	assign g778 = (((!g515) & (!g724) & (g729) & (!g701) & (!g743)) + ((!g515) & (!g724) & (g729) & (g701) & (!g743)) + ((!g515) & (!g724) & (g729) & (g701) & (g743)) + ((!g515) & (g724) & (!g729) & (!g701) & (!g743)) + ((!g515) & (g724) & (!g729) & (!g701) & (g743)) + ((!g515) & (g724) & (!g729) & (g701) & (!g743)) + ((!g515) & (g724) & (!g729) & (g701) & (g743)) + ((!g515) & (g724) & (g729) & (!g701) & (g743)) + ((g515) & (!g724) & (!g729) & (!g701) & (!g743)) + ((g515) & (!g724) & (!g729) & (g701) & (!g743)) + ((g515) & (!g724) & (!g729) & (g701) & (g743)) + ((g515) & (g724) & (!g729) & (!g701) & (g743)) + ((g515) & (g724) & (g729) & (!g701) & (!g743)) + ((g515) & (g724) & (g729) & (!g701) & (g743)) + ((g515) & (g724) & (g729) & (g701) & (!g743)) + ((g515) & (g724) & (g729) & (g701) & (g743)));
	assign g779 = (((!g553) & (!g604) & (g726) & (g728)) + ((!g553) & (g604) & (!g726) & (g728)) + ((!g553) & (g604) & (g726) & (!g728)) + ((!g553) & (g604) & (g726) & (g728)) + ((g553) & (!g604) & (!g726) & (!g728)) + ((g553) & (!g604) & (!g726) & (g728)) + ((g553) & (!g604) & (g726) & (!g728)) + ((g553) & (g604) & (!g726) & (!g728)));
	assign g780 = (((!g725) & (!g701) & (!g743) & (g779)) + ((!g725) & (g701) & (!g743) & (g779)) + ((!g725) & (g701) & (g743) & (g779)) + ((g725) & (!g701) & (!g743) & (!g779)) + ((g725) & (!g701) & (g743) & (!g779)) + ((g725) & (!g701) & (g743) & (g779)) + ((g725) & (g701) & (!g743) & (!g779)) + ((g725) & (g701) & (g743) & (!g779)));
	assign g781 = (((!g604) & (!g726) & (g728) & (!g701) & (!g743)) + ((!g604) & (!g726) & (g728) & (g701) & (!g743)) + ((!g604) & (!g726) & (g728) & (g701) & (g743)) + ((!g604) & (g726) & (!g728) & (!g701) & (!g743)) + ((!g604) & (g726) & (!g728) & (!g701) & (g743)) + ((!g604) & (g726) & (!g728) & (g701) & (!g743)) + ((!g604) & (g726) & (!g728) & (g701) & (g743)) + ((!g604) & (g726) & (g728) & (!g701) & (g743)) + ((g604) & (!g726) & (!g728) & (!g701) & (!g743)) + ((g604) & (!g726) & (!g728) & (g701) & (!g743)) + ((g604) & (!g726) & (!g728) & (g701) & (g743)) + ((g604) & (g726) & (!g728) & (!g701) & (g743)) + ((g604) & (g726) & (g728) & (!g701) & (!g743)) + ((g604) & (g726) & (g728) & (!g701) & (g743)) + ((g604) & (g726) & (g728) & (g701) & (!g743)) + ((g604) & (g726) & (g728) & (g701) & (g743)));
	assign g782 = (((!g645) & (!ax72x) & (!g700) & (g727)) + ((!g645) & (!ax72x) & (g700) & (g727)) + ((!g645) & (ax72x) & (!g700) & (!g727)) + ((!g645) & (ax72x) & (!g700) & (g727)) + ((g645) & (!ax72x) & (!g700) & (!g727)) + ((g645) & (!ax72x) & (g700) & (!g727)) + ((g645) & (ax72x) & (g700) & (!g727)) + ((g645) & (ax72x) & (g700) & (g727)));
	assign g783 = (((!ax72x) & (!ax73x) & (!g700) & (!g701) & (!g743) & (g782)) + ((!ax72x) & (!ax73x) & (!g700) & (!g701) & (g743) & (!g782)) + ((!ax72x) & (!ax73x) & (!g700) & (!g701) & (g743) & (g782)) + ((!ax72x) & (!ax73x) & (!g700) & (g701) & (!g743) & (g782)) + ((!ax72x) & (!ax73x) & (!g700) & (g701) & (g743) & (g782)) + ((!ax72x) & (!ax73x) & (g700) & (!g701) & (!g743) & (!g782)) + ((!ax72x) & (!ax73x) & (g700) & (g701) & (!g743) & (!g782)) + ((!ax72x) & (!ax73x) & (g700) & (g701) & (g743) & (!g782)) + ((!ax72x) & (ax73x) & (!g700) & (!g701) & (!g743) & (!g782)) + ((!ax72x) & (ax73x) & (!g700) & (g701) & (!g743) & (!g782)) + ((!ax72x) & (ax73x) & (!g700) & (g701) & (g743) & (!g782)) + ((!ax72x) & (ax73x) & (g700) & (!g701) & (!g743) & (g782)) + ((!ax72x) & (ax73x) & (g700) & (!g701) & (g743) & (!g782)) + ((!ax72x) & (ax73x) & (g700) & (!g701) & (g743) & (g782)) + ((!ax72x) & (ax73x) & (g700) & (g701) & (!g743) & (g782)) + ((!ax72x) & (ax73x) & (g700) & (g701) & (g743) & (g782)) + ((ax72x) & (!ax73x) & (!g700) & (!g701) & (!g743) & (!g782)) + ((ax72x) & (!ax73x) & (!g700) & (g701) & (!g743) & (!g782)) + ((ax72x) & (!ax73x) & (!g700) & (g701) & (g743) & (!g782)) + ((ax72x) & (!ax73x) & (g700) & (!g701) & (!g743) & (!g782)) + ((ax72x) & (!ax73x) & (g700) & (g701) & (!g743) & (!g782)) + ((ax72x) & (!ax73x) & (g700) & (g701) & (g743) & (!g782)) + ((ax72x) & (ax73x) & (!g700) & (!g701) & (!g743) & (g782)) + ((ax72x) & (ax73x) & (!g700) & (!g701) & (g743) & (!g782)) + ((ax72x) & (ax73x) & (!g700) & (!g701) & (g743) & (g782)) + ((ax72x) & (ax73x) & (!g700) & (g701) & (!g743) & (g782)) + ((ax72x) & (ax73x) & (!g700) & (g701) & (g743) & (g782)) + ((ax72x) & (ax73x) & (g700) & (!g701) & (!g743) & (g782)) + ((ax72x) & (ax73x) & (g700) & (!g701) & (g743) & (!g782)) + ((ax72x) & (ax73x) & (g700) & (!g701) & (g743) & (g782)) + ((ax72x) & (ax73x) & (g700) & (g701) & (!g743) & (g782)) + ((ax72x) & (ax73x) & (g700) & (g701) & (g743) & (g782)));
	assign g784 = (((!ax72x) & (!g700) & (!g727) & (!g701) & (g743)) + ((!ax72x) & (!g700) & (g727) & (!g701) & (!g743)) + ((!ax72x) & (!g700) & (g727) & (!g701) & (g743)) + ((!ax72x) & (!g700) & (g727) & (g701) & (!g743)) + ((!ax72x) & (!g700) & (g727) & (g701) & (g743)) + ((!ax72x) & (g700) & (g727) & (!g701) & (!g743)) + ((!ax72x) & (g700) & (g727) & (g701) & (!g743)) + ((!ax72x) & (g700) & (g727) & (g701) & (g743)) + ((ax72x) & (!g700) & (!g727) & (!g701) & (!g743)) + ((ax72x) & (!g700) & (!g727) & (g701) & (!g743)) + ((ax72x) & (!g700) & (!g727) & (g701) & (g743)) + ((ax72x) & (g700) & (!g727) & (!g701) & (!g743)) + ((ax72x) & (g700) & (!g727) & (!g701) & (g743)) + ((ax72x) & (g700) & (!g727) & (g701) & (!g743)) + ((ax72x) & (g700) & (!g727) & (g701) & (g743)) + ((ax72x) & (g700) & (g727) & (!g701) & (g743)));
	assign g785 = (((!ax68x) & (!ax69x)));
	assign g786 = (((!g700) & (!ax70x) & (!ax71x) & (!g701) & (!g743) & (!g785)) + ((!g700) & (!ax70x) & (!ax71x) & (g701) & (!g743) & (!g785)) + ((!g700) & (!ax70x) & (!ax71x) & (g701) & (g743) & (!g785)) + ((!g700) & (!ax70x) & (ax71x) & (!g701) & (g743) & (!g785)) + ((!g700) & (ax70x) & (ax71x) & (!g701) & (g743) & (!g785)) + ((!g700) & (ax70x) & (ax71x) & (!g701) & (g743) & (g785)) + ((g700) & (!ax70x) & (!ax71x) & (!g701) & (!g743) & (!g785)) + ((g700) & (!ax70x) & (!ax71x) & (!g701) & (!g743) & (g785)) + ((g700) & (!ax70x) & (!ax71x) & (!g701) & (g743) & (!g785)) + ((g700) & (!ax70x) & (!ax71x) & (g701) & (!g743) & (!g785)) + ((g700) & (!ax70x) & (!ax71x) & (g701) & (!g743) & (g785)) + ((g700) & (!ax70x) & (!ax71x) & (g701) & (g743) & (!g785)) + ((g700) & (!ax70x) & (!ax71x) & (g701) & (g743) & (g785)) + ((g700) & (!ax70x) & (ax71x) & (!g701) & (!g743) & (!g785)) + ((g700) & (!ax70x) & (ax71x) & (!g701) & (g743) & (!g785)) + ((g700) & (!ax70x) & (ax71x) & (!g701) & (g743) & (g785)) + ((g700) & (!ax70x) & (ax71x) & (g701) & (!g743) & (!g785)) + ((g700) & (!ax70x) & (ax71x) & (g701) & (g743) & (!g785)) + ((g700) & (ax70x) & (!ax71x) & (!g701) & (g743) & (!g785)) + ((g700) & (ax70x) & (!ax71x) & (!g701) & (g743) & (g785)) + ((g700) & (ax70x) & (ax71x) & (!g701) & (!g743) & (!g785)) + ((g700) & (ax70x) & (ax71x) & (!g701) & (!g743) & (g785)) + ((g700) & (ax70x) & (ax71x) & (!g701) & (g743) & (!g785)) + ((g700) & (ax70x) & (ax71x) & (!g701) & (g743) & (g785)) + ((g700) & (ax70x) & (ax71x) & (g701) & (!g743) & (!g785)) + ((g700) & (ax70x) & (ax71x) & (g701) & (!g743) & (g785)) + ((g700) & (ax70x) & (ax71x) & (g701) & (g743) & (!g785)) + ((g700) & (ax70x) & (ax71x) & (g701) & (g743) & (g785)));
	assign g787 = (((!g604) & (!g645) & (g783) & (g784) & (g786)) + ((!g604) & (g645) & (g783) & (!g784) & (g786)) + ((!g604) & (g645) & (g783) & (g784) & (!g786)) + ((!g604) & (g645) & (g783) & (g784) & (g786)) + ((g604) & (!g645) & (!g783) & (g784) & (g786)) + ((g604) & (!g645) & (g783) & (!g784) & (!g786)) + ((g604) & (!g645) & (g783) & (!g784) & (g786)) + ((g604) & (!g645) & (g783) & (g784) & (!g786)) + ((g604) & (!g645) & (g783) & (g784) & (g786)) + ((g604) & (g645) & (!g783) & (!g784) & (g786)) + ((g604) & (g645) & (!g783) & (g784) & (!g786)) + ((g604) & (g645) & (!g783) & (g784) & (g786)) + ((g604) & (g645) & (g783) & (!g784) & (!g786)) + ((g604) & (g645) & (g783) & (!g784) & (g786)) + ((g604) & (g645) & (g783) & (g784) & (!g786)) + ((g604) & (g645) & (g783) & (g784) & (g786)));
	assign g788 = (((!g515) & (!g553) & (g780) & (g781) & (g787)) + ((!g515) & (g553) & (g780) & (!g781) & (g787)) + ((!g515) & (g553) & (g780) & (g781) & (!g787)) + ((!g515) & (g553) & (g780) & (g781) & (g787)) + ((g515) & (!g553) & (!g780) & (g781) & (g787)) + ((g515) & (!g553) & (g780) & (!g781) & (!g787)) + ((g515) & (!g553) & (g780) & (!g781) & (g787)) + ((g515) & (!g553) & (g780) & (g781) & (!g787)) + ((g515) & (!g553) & (g780) & (g781) & (g787)) + ((g515) & (g553) & (!g780) & (!g781) & (g787)) + ((g515) & (g553) & (!g780) & (g781) & (!g787)) + ((g515) & (g553) & (!g780) & (g781) & (g787)) + ((g515) & (g553) & (g780) & (!g781) & (!g787)) + ((g515) & (g553) & (g780) & (!g781) & (g787)) + ((g515) & (g553) & (g780) & (g781) & (!g787)) + ((g515) & (g553) & (g780) & (g781) & (g787)));
	assign g789 = (((!g433) & (!g468) & (g777) & (g778) & (g788)) + ((!g433) & (g468) & (g777) & (!g778) & (g788)) + ((!g433) & (g468) & (g777) & (g778) & (!g788)) + ((!g433) & (g468) & (g777) & (g778) & (g788)) + ((g433) & (!g468) & (!g777) & (g778) & (g788)) + ((g433) & (!g468) & (g777) & (!g778) & (!g788)) + ((g433) & (!g468) & (g777) & (!g778) & (g788)) + ((g433) & (!g468) & (g777) & (g778) & (!g788)) + ((g433) & (!g468) & (g777) & (g778) & (g788)) + ((g433) & (g468) & (!g777) & (!g778) & (g788)) + ((g433) & (g468) & (!g777) & (g778) & (!g788)) + ((g433) & (g468) & (!g777) & (g778) & (g788)) + ((g433) & (g468) & (g777) & (!g778) & (!g788)) + ((g433) & (g468) & (g777) & (!g778) & (g788)) + ((g433) & (g468) & (g777) & (g778) & (!g788)) + ((g433) & (g468) & (g777) & (g778) & (g788)));
	assign g790 = (((!g358) & (!g390) & (g774) & (g775) & (g789)) + ((!g358) & (g390) & (g774) & (!g775) & (g789)) + ((!g358) & (g390) & (g774) & (g775) & (!g789)) + ((!g358) & (g390) & (g774) & (g775) & (g789)) + ((g358) & (!g390) & (!g774) & (g775) & (g789)) + ((g358) & (!g390) & (g774) & (!g775) & (!g789)) + ((g358) & (!g390) & (g774) & (!g775) & (g789)) + ((g358) & (!g390) & (g774) & (g775) & (!g789)) + ((g358) & (!g390) & (g774) & (g775) & (g789)) + ((g358) & (g390) & (!g774) & (!g775) & (g789)) + ((g358) & (g390) & (!g774) & (g775) & (!g789)) + ((g358) & (g390) & (!g774) & (g775) & (g789)) + ((g358) & (g390) & (g774) & (!g775) & (!g789)) + ((g358) & (g390) & (g774) & (!g775) & (g789)) + ((g358) & (g390) & (g774) & (g775) & (!g789)) + ((g358) & (g390) & (g774) & (g775) & (g789)));
	assign g791 = (((!g290) & (!g319) & (g771) & (g772) & (g790)) + ((!g290) & (g319) & (g771) & (!g772) & (g790)) + ((!g290) & (g319) & (g771) & (g772) & (!g790)) + ((!g290) & (g319) & (g771) & (g772) & (g790)) + ((g290) & (!g319) & (!g771) & (g772) & (g790)) + ((g290) & (!g319) & (g771) & (!g772) & (!g790)) + ((g290) & (!g319) & (g771) & (!g772) & (g790)) + ((g290) & (!g319) & (g771) & (g772) & (!g790)) + ((g290) & (!g319) & (g771) & (g772) & (g790)) + ((g290) & (g319) & (!g771) & (!g772) & (g790)) + ((g290) & (g319) & (!g771) & (g772) & (!g790)) + ((g290) & (g319) & (!g771) & (g772) & (g790)) + ((g290) & (g319) & (g771) & (!g772) & (!g790)) + ((g290) & (g319) & (g771) & (!g772) & (g790)) + ((g290) & (g319) & (g771) & (g772) & (!g790)) + ((g290) & (g319) & (g771) & (g772) & (g790)));
	assign g792 = (((!g229) & (!g255) & (g768) & (g769) & (g791)) + ((!g229) & (g255) & (g768) & (!g769) & (g791)) + ((!g229) & (g255) & (g768) & (g769) & (!g791)) + ((!g229) & (g255) & (g768) & (g769) & (g791)) + ((g229) & (!g255) & (!g768) & (g769) & (g791)) + ((g229) & (!g255) & (g768) & (!g769) & (!g791)) + ((g229) & (!g255) & (g768) & (!g769) & (g791)) + ((g229) & (!g255) & (g768) & (g769) & (!g791)) + ((g229) & (!g255) & (g768) & (g769) & (g791)) + ((g229) & (g255) & (!g768) & (!g769) & (g791)) + ((g229) & (g255) & (!g768) & (g769) & (!g791)) + ((g229) & (g255) & (!g768) & (g769) & (g791)) + ((g229) & (g255) & (g768) & (!g769) & (!g791)) + ((g229) & (g255) & (g768) & (!g769) & (g791)) + ((g229) & (g255) & (g768) & (g769) & (!g791)) + ((g229) & (g255) & (g768) & (g769) & (g791)));
	assign g793 = (((!g174) & (!g198) & (g765) & (g766) & (g792)) + ((!g174) & (g198) & (g765) & (!g766) & (g792)) + ((!g174) & (g198) & (g765) & (g766) & (!g792)) + ((!g174) & (g198) & (g765) & (g766) & (g792)) + ((g174) & (!g198) & (!g765) & (g766) & (g792)) + ((g174) & (!g198) & (g765) & (!g766) & (!g792)) + ((g174) & (!g198) & (g765) & (!g766) & (g792)) + ((g174) & (!g198) & (g765) & (g766) & (!g792)) + ((g174) & (!g198) & (g765) & (g766) & (g792)) + ((g174) & (g198) & (!g765) & (!g766) & (g792)) + ((g174) & (g198) & (!g765) & (g766) & (!g792)) + ((g174) & (g198) & (!g765) & (g766) & (g792)) + ((g174) & (g198) & (g765) & (!g766) & (!g792)) + ((g174) & (g198) & (g765) & (!g766) & (g792)) + ((g174) & (g198) & (g765) & (g766) & (!g792)) + ((g174) & (g198) & (g765) & (g766) & (g792)));
	assign g794 = (((!g127) & (!g147) & (g762) & (g763) & (g793)) + ((!g127) & (g147) & (g762) & (!g763) & (g793)) + ((!g127) & (g147) & (g762) & (g763) & (!g793)) + ((!g127) & (g147) & (g762) & (g763) & (g793)) + ((g127) & (!g147) & (!g762) & (g763) & (g793)) + ((g127) & (!g147) & (g762) & (!g763) & (!g793)) + ((g127) & (!g147) & (g762) & (!g763) & (g793)) + ((g127) & (!g147) & (g762) & (g763) & (!g793)) + ((g127) & (!g147) & (g762) & (g763) & (g793)) + ((g127) & (g147) & (!g762) & (!g763) & (g793)) + ((g127) & (g147) & (!g762) & (g763) & (!g793)) + ((g127) & (g147) & (!g762) & (g763) & (g793)) + ((g127) & (g147) & (g762) & (!g763) & (!g793)) + ((g127) & (g147) & (g762) & (!g763) & (g793)) + ((g127) & (g147) & (g762) & (g763) & (!g793)) + ((g127) & (g147) & (g762) & (g763) & (g793)));
	assign g795 = (((!g87) & (!g104) & (g759) & (g760) & (g794)) + ((!g87) & (g104) & (g759) & (!g760) & (g794)) + ((!g87) & (g104) & (g759) & (g760) & (!g794)) + ((!g87) & (g104) & (g759) & (g760) & (g794)) + ((g87) & (!g104) & (!g759) & (g760) & (g794)) + ((g87) & (!g104) & (g759) & (!g760) & (!g794)) + ((g87) & (!g104) & (g759) & (!g760) & (g794)) + ((g87) & (!g104) & (g759) & (g760) & (!g794)) + ((g87) & (!g104) & (g759) & (g760) & (g794)) + ((g87) & (g104) & (!g759) & (!g760) & (g794)) + ((g87) & (g104) & (!g759) & (g760) & (!g794)) + ((g87) & (g104) & (!g759) & (g760) & (g794)) + ((g87) & (g104) & (g759) & (!g760) & (!g794)) + ((g87) & (g104) & (g759) & (!g760) & (g794)) + ((g87) & (g104) & (g759) & (g760) & (!g794)) + ((g87) & (g104) & (g759) & (g760) & (g794)));
	assign g796 = (((!g54) & (!g68) & (g756) & (g757) & (g795)) + ((!g54) & (g68) & (g756) & (!g757) & (g795)) + ((!g54) & (g68) & (g756) & (g757) & (!g795)) + ((!g54) & (g68) & (g756) & (g757) & (g795)) + ((g54) & (!g68) & (!g756) & (g757) & (g795)) + ((g54) & (!g68) & (g756) & (!g757) & (!g795)) + ((g54) & (!g68) & (g756) & (!g757) & (g795)) + ((g54) & (!g68) & (g756) & (g757) & (!g795)) + ((g54) & (!g68) & (g756) & (g757) & (g795)) + ((g54) & (g68) & (!g756) & (!g757) & (g795)) + ((g54) & (g68) & (!g756) & (g757) & (!g795)) + ((g54) & (g68) & (!g756) & (g757) & (g795)) + ((g54) & (g68) & (g756) & (!g757) & (!g795)) + ((g54) & (g68) & (g756) & (!g757) & (g795)) + ((g54) & (g68) & (g756) & (g757) & (!g795)) + ((g54) & (g68) & (g756) & (g757) & (g795)));
	assign g797 = (((!g27) & (!g39) & (g753) & (g754) & (g796)) + ((!g27) & (g39) & (g753) & (!g754) & (g796)) + ((!g27) & (g39) & (g753) & (g754) & (!g796)) + ((!g27) & (g39) & (g753) & (g754) & (g796)) + ((g27) & (!g39) & (!g753) & (g754) & (g796)) + ((g27) & (!g39) & (g753) & (!g754) & (!g796)) + ((g27) & (!g39) & (g753) & (!g754) & (g796)) + ((g27) & (!g39) & (g753) & (g754) & (!g796)) + ((g27) & (!g39) & (g753) & (g754) & (g796)) + ((g27) & (g39) & (!g753) & (!g754) & (g796)) + ((g27) & (g39) & (!g753) & (g754) & (!g796)) + ((g27) & (g39) & (!g753) & (g754) & (g796)) + ((g27) & (g39) & (g753) & (!g754) & (!g796)) + ((g27) & (g39) & (g753) & (!g754) & (g796)) + ((g27) & (g39) & (g753) & (g754) & (!g796)) + ((g27) & (g39) & (g753) & (g754) & (g796)));
	assign g798 = (((!g8) & (!g18) & (g750) & (g751) & (g797)) + ((!g8) & (g18) & (g750) & (!g751) & (g797)) + ((!g8) & (g18) & (g750) & (g751) & (!g797)) + ((!g8) & (g18) & (g750) & (g751) & (g797)) + ((g8) & (!g18) & (!g750) & (g751) & (g797)) + ((g8) & (!g18) & (g750) & (!g751) & (!g797)) + ((g8) & (!g18) & (g750) & (!g751) & (g797)) + ((g8) & (!g18) & (g750) & (g751) & (!g797)) + ((g8) & (!g18) & (g750) & (g751) & (g797)) + ((g8) & (g18) & (!g750) & (!g751) & (g797)) + ((g8) & (g18) & (!g750) & (g751) & (!g797)) + ((g8) & (g18) & (!g750) & (g751) & (g797)) + ((g8) & (g18) & (g750) & (!g751) & (!g797)) + ((g8) & (g18) & (g750) & (!g751) & (g797)) + ((g8) & (g18) & (g750) & (g751) & (!g797)) + ((g8) & (g18) & (g750) & (g751) & (g797)));
	assign g799 = (((!g4) & (!g2) & (!g747) & (g748) & (g798)) + ((!g4) & (!g2) & (g747) & (!g748) & (!g798)) + ((!g4) & (!g2) & (g747) & (!g748) & (g798)) + ((!g4) & (!g2) & (g747) & (g748) & (!g798)) + ((!g4) & (!g2) & (g747) & (g748) & (g798)) + ((!g4) & (g2) & (!g747) & (!g748) & (g798)) + ((!g4) & (g2) & (!g747) & (g748) & (!g798)) + ((!g4) & (g2) & (!g747) & (g748) & (g798)) + ((!g4) & (g2) & (g747) & (!g748) & (!g798)) + ((!g4) & (g2) & (g747) & (!g748) & (g798)) + ((!g4) & (g2) & (g747) & (g748) & (!g798)) + ((!g4) & (g2) & (g747) & (g748) & (g798)) + ((g4) & (!g2) & (g747) & (g748) & (g798)) + ((g4) & (g2) & (g747) & (!g748) & (g798)) + ((g4) & (g2) & (g747) & (g748) & (!g798)) + ((g4) & (g2) & (g747) & (g748) & (g798)));
	assign g800 = (((!g4) & (!g740) & (g741)) + ((!g4) & (g740) & (!g741)) + ((!g4) & (g740) & (g741)) + ((g4) & (g740) & (g741)));
	assign g801 = (((!g702) & (!g800) & (!g701) & (!g743)) + ((!g702) & (!g800) & (g701) & (!g743)) + ((!g702) & (!g800) & (g701) & (g743)) + ((g702) & (g800) & (!g701) & (!g743)) + ((g702) & (g800) & (!g701) & (g743)) + ((g702) & (g800) & (g701) & (!g743)) + ((g702) & (g800) & (g701) & (g743)));
	assign g802 = (((!g1) & (g702) & (!g800) & (!g701) & (g743)) + ((!g1) & (g702) & (g800) & (!g701) & (g743)) + ((g1) & (!g702) & (g800) & (g701) & (!g743)) + ((g1) & (!g702) & (g800) & (g701) & (g743)) + ((g1) & (g702) & (!g800) & (!g701) & (!g743)) + ((g1) & (g702) & (!g800) & (!g701) & (g743)) + ((g1) & (g702) & (!g800) & (g701) & (!g743)) + ((g1) & (g702) & (!g800) & (g701) & (g743)) + ((g1) & (g702) & (g800) & (!g701) & (g743)));
	assign g803 = (((!g1) & (!g745) & (!g799) & (!g801) & (!g802)) + ((g1) & (!g745) & (!g799) & (!g801) & (!g802)) + ((g1) & (!g745) & (!g799) & (g801) & (!g802)) + ((g1) & (!g745) & (g799) & (!g801) & (!g802)) + ((g1) & (!g745) & (g799) & (g801) & (!g802)) + ((g1) & (g745) & (!g799) & (!g801) & (!g802)) + ((g1) & (g745) & (!g799) & (g801) & (!g802)));
	assign g804 = (((!g4) & (!g2) & (!g747) & (!g748) & (!g798) & (!g803)) + ((!g4) & (!g2) & (!g747) & (!g748) & (g798) & (!g803)) + ((!g4) & (!g2) & (!g747) & (g748) & (!g798) & (!g803)) + ((!g4) & (!g2) & (g747) & (!g748) & (!g798) & (g803)) + ((!g4) & (!g2) & (g747) & (!g748) & (g798) & (g803)) + ((!g4) & (!g2) & (g747) & (g748) & (!g798) & (g803)) + ((!g4) & (!g2) & (g747) & (g748) & (g798) & (!g803)) + ((!g4) & (!g2) & (g747) & (g748) & (g798) & (g803)) + ((!g4) & (g2) & (!g747) & (!g748) & (!g798) & (!g803)) + ((!g4) & (g2) & (g747) & (!g748) & (!g798) & (g803)) + ((!g4) & (g2) & (g747) & (!g748) & (g798) & (!g803)) + ((!g4) & (g2) & (g747) & (!g748) & (g798) & (g803)) + ((!g4) & (g2) & (g747) & (g748) & (!g798) & (!g803)) + ((!g4) & (g2) & (g747) & (g748) & (!g798) & (g803)) + ((!g4) & (g2) & (g747) & (g748) & (g798) & (!g803)) + ((!g4) & (g2) & (g747) & (g748) & (g798) & (g803)) + ((g4) & (!g2) & (!g747) & (g748) & (g798) & (!g803)) + ((g4) & (!g2) & (g747) & (!g748) & (!g798) & (!g803)) + ((g4) & (!g2) & (g747) & (!g748) & (!g798) & (g803)) + ((g4) & (!g2) & (g747) & (!g748) & (g798) & (!g803)) + ((g4) & (!g2) & (g747) & (!g748) & (g798) & (g803)) + ((g4) & (!g2) & (g747) & (g748) & (!g798) & (!g803)) + ((g4) & (!g2) & (g747) & (g748) & (!g798) & (g803)) + ((g4) & (!g2) & (g747) & (g748) & (g798) & (g803)) + ((g4) & (g2) & (!g747) & (!g748) & (g798) & (!g803)) + ((g4) & (g2) & (!g747) & (g748) & (!g798) & (!g803)) + ((g4) & (g2) & (!g747) & (g748) & (g798) & (!g803)) + ((g4) & (g2) & (g747) & (!g748) & (!g798) & (!g803)) + ((g4) & (g2) & (g747) & (!g748) & (!g798) & (g803)) + ((g4) & (g2) & (g747) & (!g748) & (g798) & (g803)) + ((g4) & (g2) & (g747) & (g748) & (!g798) & (g803)) + ((g4) & (g2) & (g747) & (g748) & (g798) & (g803)));
	assign g805 = (((!g8) & (!g18) & (!g750) & (g751) & (g797) & (!g803)) + ((!g8) & (!g18) & (g750) & (!g751) & (!g797) & (!g803)) + ((!g8) & (!g18) & (g750) & (!g751) & (!g797) & (g803)) + ((!g8) & (!g18) & (g750) & (!g751) & (g797) & (!g803)) + ((!g8) & (!g18) & (g750) & (!g751) & (g797) & (g803)) + ((!g8) & (!g18) & (g750) & (g751) & (!g797) & (!g803)) + ((!g8) & (!g18) & (g750) & (g751) & (!g797) & (g803)) + ((!g8) & (!g18) & (g750) & (g751) & (g797) & (g803)) + ((!g8) & (g18) & (!g750) & (!g751) & (g797) & (!g803)) + ((!g8) & (g18) & (!g750) & (g751) & (!g797) & (!g803)) + ((!g8) & (g18) & (!g750) & (g751) & (g797) & (!g803)) + ((!g8) & (g18) & (g750) & (!g751) & (!g797) & (!g803)) + ((!g8) & (g18) & (g750) & (!g751) & (!g797) & (g803)) + ((!g8) & (g18) & (g750) & (!g751) & (g797) & (g803)) + ((!g8) & (g18) & (g750) & (g751) & (!g797) & (g803)) + ((!g8) & (g18) & (g750) & (g751) & (g797) & (g803)) + ((g8) & (!g18) & (!g750) & (!g751) & (!g797) & (!g803)) + ((g8) & (!g18) & (!g750) & (!g751) & (g797) & (!g803)) + ((g8) & (!g18) & (!g750) & (g751) & (!g797) & (!g803)) + ((g8) & (!g18) & (g750) & (!g751) & (!g797) & (g803)) + ((g8) & (!g18) & (g750) & (!g751) & (g797) & (g803)) + ((g8) & (!g18) & (g750) & (g751) & (!g797) & (g803)) + ((g8) & (!g18) & (g750) & (g751) & (g797) & (!g803)) + ((g8) & (!g18) & (g750) & (g751) & (g797) & (g803)) + ((g8) & (g18) & (!g750) & (!g751) & (!g797) & (!g803)) + ((g8) & (g18) & (g750) & (!g751) & (!g797) & (g803)) + ((g8) & (g18) & (g750) & (!g751) & (g797) & (!g803)) + ((g8) & (g18) & (g750) & (!g751) & (g797) & (g803)) + ((g8) & (g18) & (g750) & (g751) & (!g797) & (!g803)) + ((g8) & (g18) & (g750) & (g751) & (!g797) & (g803)) + ((g8) & (g18) & (g750) & (g751) & (g797) & (!g803)) + ((g8) & (g18) & (g750) & (g751) & (g797) & (g803)));
	assign g806 = (((!g18) & (!g751) & (g797) & (!g803)) + ((!g18) & (g751) & (!g797) & (!g803)) + ((!g18) & (g751) & (!g797) & (g803)) + ((!g18) & (g751) & (g797) & (g803)) + ((g18) & (!g751) & (!g797) & (!g803)) + ((g18) & (g751) & (!g797) & (g803)) + ((g18) & (g751) & (g797) & (!g803)) + ((g18) & (g751) & (g797) & (g803)));
	assign g807 = (((!g27) & (!g39) & (!g753) & (g754) & (g796) & (!g803)) + ((!g27) & (!g39) & (g753) & (!g754) & (!g796) & (!g803)) + ((!g27) & (!g39) & (g753) & (!g754) & (!g796) & (g803)) + ((!g27) & (!g39) & (g753) & (!g754) & (g796) & (!g803)) + ((!g27) & (!g39) & (g753) & (!g754) & (g796) & (g803)) + ((!g27) & (!g39) & (g753) & (g754) & (!g796) & (!g803)) + ((!g27) & (!g39) & (g753) & (g754) & (!g796) & (g803)) + ((!g27) & (!g39) & (g753) & (g754) & (g796) & (g803)) + ((!g27) & (g39) & (!g753) & (!g754) & (g796) & (!g803)) + ((!g27) & (g39) & (!g753) & (g754) & (!g796) & (!g803)) + ((!g27) & (g39) & (!g753) & (g754) & (g796) & (!g803)) + ((!g27) & (g39) & (g753) & (!g754) & (!g796) & (!g803)) + ((!g27) & (g39) & (g753) & (!g754) & (!g796) & (g803)) + ((!g27) & (g39) & (g753) & (!g754) & (g796) & (g803)) + ((!g27) & (g39) & (g753) & (g754) & (!g796) & (g803)) + ((!g27) & (g39) & (g753) & (g754) & (g796) & (g803)) + ((g27) & (!g39) & (!g753) & (!g754) & (!g796) & (!g803)) + ((g27) & (!g39) & (!g753) & (!g754) & (g796) & (!g803)) + ((g27) & (!g39) & (!g753) & (g754) & (!g796) & (!g803)) + ((g27) & (!g39) & (g753) & (!g754) & (!g796) & (g803)) + ((g27) & (!g39) & (g753) & (!g754) & (g796) & (g803)) + ((g27) & (!g39) & (g753) & (g754) & (!g796) & (g803)) + ((g27) & (!g39) & (g753) & (g754) & (g796) & (!g803)) + ((g27) & (!g39) & (g753) & (g754) & (g796) & (g803)) + ((g27) & (g39) & (!g753) & (!g754) & (!g796) & (!g803)) + ((g27) & (g39) & (g753) & (!g754) & (!g796) & (g803)) + ((g27) & (g39) & (g753) & (!g754) & (g796) & (!g803)) + ((g27) & (g39) & (g753) & (!g754) & (g796) & (g803)) + ((g27) & (g39) & (g753) & (g754) & (!g796) & (!g803)) + ((g27) & (g39) & (g753) & (g754) & (!g796) & (g803)) + ((g27) & (g39) & (g753) & (g754) & (g796) & (!g803)) + ((g27) & (g39) & (g753) & (g754) & (g796) & (g803)));
	assign g808 = (((!g39) & (!g754) & (g796) & (!g803)) + ((!g39) & (g754) & (!g796) & (!g803)) + ((!g39) & (g754) & (!g796) & (g803)) + ((!g39) & (g754) & (g796) & (g803)) + ((g39) & (!g754) & (!g796) & (!g803)) + ((g39) & (g754) & (!g796) & (g803)) + ((g39) & (g754) & (g796) & (!g803)) + ((g39) & (g754) & (g796) & (g803)));
	assign g809 = (((!g54) & (!g68) & (!g756) & (g757) & (g795) & (!g803)) + ((!g54) & (!g68) & (g756) & (!g757) & (!g795) & (!g803)) + ((!g54) & (!g68) & (g756) & (!g757) & (!g795) & (g803)) + ((!g54) & (!g68) & (g756) & (!g757) & (g795) & (!g803)) + ((!g54) & (!g68) & (g756) & (!g757) & (g795) & (g803)) + ((!g54) & (!g68) & (g756) & (g757) & (!g795) & (!g803)) + ((!g54) & (!g68) & (g756) & (g757) & (!g795) & (g803)) + ((!g54) & (!g68) & (g756) & (g757) & (g795) & (g803)) + ((!g54) & (g68) & (!g756) & (!g757) & (g795) & (!g803)) + ((!g54) & (g68) & (!g756) & (g757) & (!g795) & (!g803)) + ((!g54) & (g68) & (!g756) & (g757) & (g795) & (!g803)) + ((!g54) & (g68) & (g756) & (!g757) & (!g795) & (!g803)) + ((!g54) & (g68) & (g756) & (!g757) & (!g795) & (g803)) + ((!g54) & (g68) & (g756) & (!g757) & (g795) & (g803)) + ((!g54) & (g68) & (g756) & (g757) & (!g795) & (g803)) + ((!g54) & (g68) & (g756) & (g757) & (g795) & (g803)) + ((g54) & (!g68) & (!g756) & (!g757) & (!g795) & (!g803)) + ((g54) & (!g68) & (!g756) & (!g757) & (g795) & (!g803)) + ((g54) & (!g68) & (!g756) & (g757) & (!g795) & (!g803)) + ((g54) & (!g68) & (g756) & (!g757) & (!g795) & (g803)) + ((g54) & (!g68) & (g756) & (!g757) & (g795) & (g803)) + ((g54) & (!g68) & (g756) & (g757) & (!g795) & (g803)) + ((g54) & (!g68) & (g756) & (g757) & (g795) & (!g803)) + ((g54) & (!g68) & (g756) & (g757) & (g795) & (g803)) + ((g54) & (g68) & (!g756) & (!g757) & (!g795) & (!g803)) + ((g54) & (g68) & (g756) & (!g757) & (!g795) & (g803)) + ((g54) & (g68) & (g756) & (!g757) & (g795) & (!g803)) + ((g54) & (g68) & (g756) & (!g757) & (g795) & (g803)) + ((g54) & (g68) & (g756) & (g757) & (!g795) & (!g803)) + ((g54) & (g68) & (g756) & (g757) & (!g795) & (g803)) + ((g54) & (g68) & (g756) & (g757) & (g795) & (!g803)) + ((g54) & (g68) & (g756) & (g757) & (g795) & (g803)));
	assign g810 = (((!g68) & (!g757) & (g795) & (!g803)) + ((!g68) & (g757) & (!g795) & (!g803)) + ((!g68) & (g757) & (!g795) & (g803)) + ((!g68) & (g757) & (g795) & (g803)) + ((g68) & (!g757) & (!g795) & (!g803)) + ((g68) & (g757) & (!g795) & (g803)) + ((g68) & (g757) & (g795) & (!g803)) + ((g68) & (g757) & (g795) & (g803)));
	assign g811 = (((!g87) & (!g104) & (!g759) & (g760) & (g794) & (!g803)) + ((!g87) & (!g104) & (g759) & (!g760) & (!g794) & (!g803)) + ((!g87) & (!g104) & (g759) & (!g760) & (!g794) & (g803)) + ((!g87) & (!g104) & (g759) & (!g760) & (g794) & (!g803)) + ((!g87) & (!g104) & (g759) & (!g760) & (g794) & (g803)) + ((!g87) & (!g104) & (g759) & (g760) & (!g794) & (!g803)) + ((!g87) & (!g104) & (g759) & (g760) & (!g794) & (g803)) + ((!g87) & (!g104) & (g759) & (g760) & (g794) & (g803)) + ((!g87) & (g104) & (!g759) & (!g760) & (g794) & (!g803)) + ((!g87) & (g104) & (!g759) & (g760) & (!g794) & (!g803)) + ((!g87) & (g104) & (!g759) & (g760) & (g794) & (!g803)) + ((!g87) & (g104) & (g759) & (!g760) & (!g794) & (!g803)) + ((!g87) & (g104) & (g759) & (!g760) & (!g794) & (g803)) + ((!g87) & (g104) & (g759) & (!g760) & (g794) & (g803)) + ((!g87) & (g104) & (g759) & (g760) & (!g794) & (g803)) + ((!g87) & (g104) & (g759) & (g760) & (g794) & (g803)) + ((g87) & (!g104) & (!g759) & (!g760) & (!g794) & (!g803)) + ((g87) & (!g104) & (!g759) & (!g760) & (g794) & (!g803)) + ((g87) & (!g104) & (!g759) & (g760) & (!g794) & (!g803)) + ((g87) & (!g104) & (g759) & (!g760) & (!g794) & (g803)) + ((g87) & (!g104) & (g759) & (!g760) & (g794) & (g803)) + ((g87) & (!g104) & (g759) & (g760) & (!g794) & (g803)) + ((g87) & (!g104) & (g759) & (g760) & (g794) & (!g803)) + ((g87) & (!g104) & (g759) & (g760) & (g794) & (g803)) + ((g87) & (g104) & (!g759) & (!g760) & (!g794) & (!g803)) + ((g87) & (g104) & (g759) & (!g760) & (!g794) & (g803)) + ((g87) & (g104) & (g759) & (!g760) & (g794) & (!g803)) + ((g87) & (g104) & (g759) & (!g760) & (g794) & (g803)) + ((g87) & (g104) & (g759) & (g760) & (!g794) & (!g803)) + ((g87) & (g104) & (g759) & (g760) & (!g794) & (g803)) + ((g87) & (g104) & (g759) & (g760) & (g794) & (!g803)) + ((g87) & (g104) & (g759) & (g760) & (g794) & (g803)));
	assign g812 = (((!g104) & (!g760) & (g794) & (!g803)) + ((!g104) & (g760) & (!g794) & (!g803)) + ((!g104) & (g760) & (!g794) & (g803)) + ((!g104) & (g760) & (g794) & (g803)) + ((g104) & (!g760) & (!g794) & (!g803)) + ((g104) & (g760) & (!g794) & (g803)) + ((g104) & (g760) & (g794) & (!g803)) + ((g104) & (g760) & (g794) & (g803)));
	assign g813 = (((!g127) & (!g147) & (!g762) & (g763) & (g793) & (!g803)) + ((!g127) & (!g147) & (g762) & (!g763) & (!g793) & (!g803)) + ((!g127) & (!g147) & (g762) & (!g763) & (!g793) & (g803)) + ((!g127) & (!g147) & (g762) & (!g763) & (g793) & (!g803)) + ((!g127) & (!g147) & (g762) & (!g763) & (g793) & (g803)) + ((!g127) & (!g147) & (g762) & (g763) & (!g793) & (!g803)) + ((!g127) & (!g147) & (g762) & (g763) & (!g793) & (g803)) + ((!g127) & (!g147) & (g762) & (g763) & (g793) & (g803)) + ((!g127) & (g147) & (!g762) & (!g763) & (g793) & (!g803)) + ((!g127) & (g147) & (!g762) & (g763) & (!g793) & (!g803)) + ((!g127) & (g147) & (!g762) & (g763) & (g793) & (!g803)) + ((!g127) & (g147) & (g762) & (!g763) & (!g793) & (!g803)) + ((!g127) & (g147) & (g762) & (!g763) & (!g793) & (g803)) + ((!g127) & (g147) & (g762) & (!g763) & (g793) & (g803)) + ((!g127) & (g147) & (g762) & (g763) & (!g793) & (g803)) + ((!g127) & (g147) & (g762) & (g763) & (g793) & (g803)) + ((g127) & (!g147) & (!g762) & (!g763) & (!g793) & (!g803)) + ((g127) & (!g147) & (!g762) & (!g763) & (g793) & (!g803)) + ((g127) & (!g147) & (!g762) & (g763) & (!g793) & (!g803)) + ((g127) & (!g147) & (g762) & (!g763) & (!g793) & (g803)) + ((g127) & (!g147) & (g762) & (!g763) & (g793) & (g803)) + ((g127) & (!g147) & (g762) & (g763) & (!g793) & (g803)) + ((g127) & (!g147) & (g762) & (g763) & (g793) & (!g803)) + ((g127) & (!g147) & (g762) & (g763) & (g793) & (g803)) + ((g127) & (g147) & (!g762) & (!g763) & (!g793) & (!g803)) + ((g127) & (g147) & (g762) & (!g763) & (!g793) & (g803)) + ((g127) & (g147) & (g762) & (!g763) & (g793) & (!g803)) + ((g127) & (g147) & (g762) & (!g763) & (g793) & (g803)) + ((g127) & (g147) & (g762) & (g763) & (!g793) & (!g803)) + ((g127) & (g147) & (g762) & (g763) & (!g793) & (g803)) + ((g127) & (g147) & (g762) & (g763) & (g793) & (!g803)) + ((g127) & (g147) & (g762) & (g763) & (g793) & (g803)));
	assign g814 = (((!g147) & (!g763) & (g793) & (!g803)) + ((!g147) & (g763) & (!g793) & (!g803)) + ((!g147) & (g763) & (!g793) & (g803)) + ((!g147) & (g763) & (g793) & (g803)) + ((g147) & (!g763) & (!g793) & (!g803)) + ((g147) & (g763) & (!g793) & (g803)) + ((g147) & (g763) & (g793) & (!g803)) + ((g147) & (g763) & (g793) & (g803)));
	assign g815 = (((!g174) & (!g198) & (!g765) & (g766) & (g792) & (!g803)) + ((!g174) & (!g198) & (g765) & (!g766) & (!g792) & (!g803)) + ((!g174) & (!g198) & (g765) & (!g766) & (!g792) & (g803)) + ((!g174) & (!g198) & (g765) & (!g766) & (g792) & (!g803)) + ((!g174) & (!g198) & (g765) & (!g766) & (g792) & (g803)) + ((!g174) & (!g198) & (g765) & (g766) & (!g792) & (!g803)) + ((!g174) & (!g198) & (g765) & (g766) & (!g792) & (g803)) + ((!g174) & (!g198) & (g765) & (g766) & (g792) & (g803)) + ((!g174) & (g198) & (!g765) & (!g766) & (g792) & (!g803)) + ((!g174) & (g198) & (!g765) & (g766) & (!g792) & (!g803)) + ((!g174) & (g198) & (!g765) & (g766) & (g792) & (!g803)) + ((!g174) & (g198) & (g765) & (!g766) & (!g792) & (!g803)) + ((!g174) & (g198) & (g765) & (!g766) & (!g792) & (g803)) + ((!g174) & (g198) & (g765) & (!g766) & (g792) & (g803)) + ((!g174) & (g198) & (g765) & (g766) & (!g792) & (g803)) + ((!g174) & (g198) & (g765) & (g766) & (g792) & (g803)) + ((g174) & (!g198) & (!g765) & (!g766) & (!g792) & (!g803)) + ((g174) & (!g198) & (!g765) & (!g766) & (g792) & (!g803)) + ((g174) & (!g198) & (!g765) & (g766) & (!g792) & (!g803)) + ((g174) & (!g198) & (g765) & (!g766) & (!g792) & (g803)) + ((g174) & (!g198) & (g765) & (!g766) & (g792) & (g803)) + ((g174) & (!g198) & (g765) & (g766) & (!g792) & (g803)) + ((g174) & (!g198) & (g765) & (g766) & (g792) & (!g803)) + ((g174) & (!g198) & (g765) & (g766) & (g792) & (g803)) + ((g174) & (g198) & (!g765) & (!g766) & (!g792) & (!g803)) + ((g174) & (g198) & (g765) & (!g766) & (!g792) & (g803)) + ((g174) & (g198) & (g765) & (!g766) & (g792) & (!g803)) + ((g174) & (g198) & (g765) & (!g766) & (g792) & (g803)) + ((g174) & (g198) & (g765) & (g766) & (!g792) & (!g803)) + ((g174) & (g198) & (g765) & (g766) & (!g792) & (g803)) + ((g174) & (g198) & (g765) & (g766) & (g792) & (!g803)) + ((g174) & (g198) & (g765) & (g766) & (g792) & (g803)));
	assign g816 = (((!g198) & (!g766) & (g792) & (!g803)) + ((!g198) & (g766) & (!g792) & (!g803)) + ((!g198) & (g766) & (!g792) & (g803)) + ((!g198) & (g766) & (g792) & (g803)) + ((g198) & (!g766) & (!g792) & (!g803)) + ((g198) & (g766) & (!g792) & (g803)) + ((g198) & (g766) & (g792) & (!g803)) + ((g198) & (g766) & (g792) & (g803)));
	assign g817 = (((!g229) & (!g255) & (!g768) & (g769) & (g791) & (!g803)) + ((!g229) & (!g255) & (g768) & (!g769) & (!g791) & (!g803)) + ((!g229) & (!g255) & (g768) & (!g769) & (!g791) & (g803)) + ((!g229) & (!g255) & (g768) & (!g769) & (g791) & (!g803)) + ((!g229) & (!g255) & (g768) & (!g769) & (g791) & (g803)) + ((!g229) & (!g255) & (g768) & (g769) & (!g791) & (!g803)) + ((!g229) & (!g255) & (g768) & (g769) & (!g791) & (g803)) + ((!g229) & (!g255) & (g768) & (g769) & (g791) & (g803)) + ((!g229) & (g255) & (!g768) & (!g769) & (g791) & (!g803)) + ((!g229) & (g255) & (!g768) & (g769) & (!g791) & (!g803)) + ((!g229) & (g255) & (!g768) & (g769) & (g791) & (!g803)) + ((!g229) & (g255) & (g768) & (!g769) & (!g791) & (!g803)) + ((!g229) & (g255) & (g768) & (!g769) & (!g791) & (g803)) + ((!g229) & (g255) & (g768) & (!g769) & (g791) & (g803)) + ((!g229) & (g255) & (g768) & (g769) & (!g791) & (g803)) + ((!g229) & (g255) & (g768) & (g769) & (g791) & (g803)) + ((g229) & (!g255) & (!g768) & (!g769) & (!g791) & (!g803)) + ((g229) & (!g255) & (!g768) & (!g769) & (g791) & (!g803)) + ((g229) & (!g255) & (!g768) & (g769) & (!g791) & (!g803)) + ((g229) & (!g255) & (g768) & (!g769) & (!g791) & (g803)) + ((g229) & (!g255) & (g768) & (!g769) & (g791) & (g803)) + ((g229) & (!g255) & (g768) & (g769) & (!g791) & (g803)) + ((g229) & (!g255) & (g768) & (g769) & (g791) & (!g803)) + ((g229) & (!g255) & (g768) & (g769) & (g791) & (g803)) + ((g229) & (g255) & (!g768) & (!g769) & (!g791) & (!g803)) + ((g229) & (g255) & (g768) & (!g769) & (!g791) & (g803)) + ((g229) & (g255) & (g768) & (!g769) & (g791) & (!g803)) + ((g229) & (g255) & (g768) & (!g769) & (g791) & (g803)) + ((g229) & (g255) & (g768) & (g769) & (!g791) & (!g803)) + ((g229) & (g255) & (g768) & (g769) & (!g791) & (g803)) + ((g229) & (g255) & (g768) & (g769) & (g791) & (!g803)) + ((g229) & (g255) & (g768) & (g769) & (g791) & (g803)));
	assign g818 = (((!g255) & (!g769) & (g791) & (!g803)) + ((!g255) & (g769) & (!g791) & (!g803)) + ((!g255) & (g769) & (!g791) & (g803)) + ((!g255) & (g769) & (g791) & (g803)) + ((g255) & (!g769) & (!g791) & (!g803)) + ((g255) & (g769) & (!g791) & (g803)) + ((g255) & (g769) & (g791) & (!g803)) + ((g255) & (g769) & (g791) & (g803)));
	assign g819 = (((!g290) & (!g319) & (!g771) & (g772) & (g790) & (!g803)) + ((!g290) & (!g319) & (g771) & (!g772) & (!g790) & (!g803)) + ((!g290) & (!g319) & (g771) & (!g772) & (!g790) & (g803)) + ((!g290) & (!g319) & (g771) & (!g772) & (g790) & (!g803)) + ((!g290) & (!g319) & (g771) & (!g772) & (g790) & (g803)) + ((!g290) & (!g319) & (g771) & (g772) & (!g790) & (!g803)) + ((!g290) & (!g319) & (g771) & (g772) & (!g790) & (g803)) + ((!g290) & (!g319) & (g771) & (g772) & (g790) & (g803)) + ((!g290) & (g319) & (!g771) & (!g772) & (g790) & (!g803)) + ((!g290) & (g319) & (!g771) & (g772) & (!g790) & (!g803)) + ((!g290) & (g319) & (!g771) & (g772) & (g790) & (!g803)) + ((!g290) & (g319) & (g771) & (!g772) & (!g790) & (!g803)) + ((!g290) & (g319) & (g771) & (!g772) & (!g790) & (g803)) + ((!g290) & (g319) & (g771) & (!g772) & (g790) & (g803)) + ((!g290) & (g319) & (g771) & (g772) & (!g790) & (g803)) + ((!g290) & (g319) & (g771) & (g772) & (g790) & (g803)) + ((g290) & (!g319) & (!g771) & (!g772) & (!g790) & (!g803)) + ((g290) & (!g319) & (!g771) & (!g772) & (g790) & (!g803)) + ((g290) & (!g319) & (!g771) & (g772) & (!g790) & (!g803)) + ((g290) & (!g319) & (g771) & (!g772) & (!g790) & (g803)) + ((g290) & (!g319) & (g771) & (!g772) & (g790) & (g803)) + ((g290) & (!g319) & (g771) & (g772) & (!g790) & (g803)) + ((g290) & (!g319) & (g771) & (g772) & (g790) & (!g803)) + ((g290) & (!g319) & (g771) & (g772) & (g790) & (g803)) + ((g290) & (g319) & (!g771) & (!g772) & (!g790) & (!g803)) + ((g290) & (g319) & (g771) & (!g772) & (!g790) & (g803)) + ((g290) & (g319) & (g771) & (!g772) & (g790) & (!g803)) + ((g290) & (g319) & (g771) & (!g772) & (g790) & (g803)) + ((g290) & (g319) & (g771) & (g772) & (!g790) & (!g803)) + ((g290) & (g319) & (g771) & (g772) & (!g790) & (g803)) + ((g290) & (g319) & (g771) & (g772) & (g790) & (!g803)) + ((g290) & (g319) & (g771) & (g772) & (g790) & (g803)));
	assign g820 = (((!g319) & (!g772) & (g790) & (!g803)) + ((!g319) & (g772) & (!g790) & (!g803)) + ((!g319) & (g772) & (!g790) & (g803)) + ((!g319) & (g772) & (g790) & (g803)) + ((g319) & (!g772) & (!g790) & (!g803)) + ((g319) & (g772) & (!g790) & (g803)) + ((g319) & (g772) & (g790) & (!g803)) + ((g319) & (g772) & (g790) & (g803)));
	assign g821 = (((!g358) & (!g390) & (!g774) & (g775) & (g789) & (!g803)) + ((!g358) & (!g390) & (g774) & (!g775) & (!g789) & (!g803)) + ((!g358) & (!g390) & (g774) & (!g775) & (!g789) & (g803)) + ((!g358) & (!g390) & (g774) & (!g775) & (g789) & (!g803)) + ((!g358) & (!g390) & (g774) & (!g775) & (g789) & (g803)) + ((!g358) & (!g390) & (g774) & (g775) & (!g789) & (!g803)) + ((!g358) & (!g390) & (g774) & (g775) & (!g789) & (g803)) + ((!g358) & (!g390) & (g774) & (g775) & (g789) & (g803)) + ((!g358) & (g390) & (!g774) & (!g775) & (g789) & (!g803)) + ((!g358) & (g390) & (!g774) & (g775) & (!g789) & (!g803)) + ((!g358) & (g390) & (!g774) & (g775) & (g789) & (!g803)) + ((!g358) & (g390) & (g774) & (!g775) & (!g789) & (!g803)) + ((!g358) & (g390) & (g774) & (!g775) & (!g789) & (g803)) + ((!g358) & (g390) & (g774) & (!g775) & (g789) & (g803)) + ((!g358) & (g390) & (g774) & (g775) & (!g789) & (g803)) + ((!g358) & (g390) & (g774) & (g775) & (g789) & (g803)) + ((g358) & (!g390) & (!g774) & (!g775) & (!g789) & (!g803)) + ((g358) & (!g390) & (!g774) & (!g775) & (g789) & (!g803)) + ((g358) & (!g390) & (!g774) & (g775) & (!g789) & (!g803)) + ((g358) & (!g390) & (g774) & (!g775) & (!g789) & (g803)) + ((g358) & (!g390) & (g774) & (!g775) & (g789) & (g803)) + ((g358) & (!g390) & (g774) & (g775) & (!g789) & (g803)) + ((g358) & (!g390) & (g774) & (g775) & (g789) & (!g803)) + ((g358) & (!g390) & (g774) & (g775) & (g789) & (g803)) + ((g358) & (g390) & (!g774) & (!g775) & (!g789) & (!g803)) + ((g358) & (g390) & (g774) & (!g775) & (!g789) & (g803)) + ((g358) & (g390) & (g774) & (!g775) & (g789) & (!g803)) + ((g358) & (g390) & (g774) & (!g775) & (g789) & (g803)) + ((g358) & (g390) & (g774) & (g775) & (!g789) & (!g803)) + ((g358) & (g390) & (g774) & (g775) & (!g789) & (g803)) + ((g358) & (g390) & (g774) & (g775) & (g789) & (!g803)) + ((g358) & (g390) & (g774) & (g775) & (g789) & (g803)));
	assign g822 = (((!g390) & (!g775) & (g789) & (!g803)) + ((!g390) & (g775) & (!g789) & (!g803)) + ((!g390) & (g775) & (!g789) & (g803)) + ((!g390) & (g775) & (g789) & (g803)) + ((g390) & (!g775) & (!g789) & (!g803)) + ((g390) & (g775) & (!g789) & (g803)) + ((g390) & (g775) & (g789) & (!g803)) + ((g390) & (g775) & (g789) & (g803)));
	assign g823 = (((!g433) & (!g468) & (!g777) & (g778) & (g788) & (!g803)) + ((!g433) & (!g468) & (g777) & (!g778) & (!g788) & (!g803)) + ((!g433) & (!g468) & (g777) & (!g778) & (!g788) & (g803)) + ((!g433) & (!g468) & (g777) & (!g778) & (g788) & (!g803)) + ((!g433) & (!g468) & (g777) & (!g778) & (g788) & (g803)) + ((!g433) & (!g468) & (g777) & (g778) & (!g788) & (!g803)) + ((!g433) & (!g468) & (g777) & (g778) & (!g788) & (g803)) + ((!g433) & (!g468) & (g777) & (g778) & (g788) & (g803)) + ((!g433) & (g468) & (!g777) & (!g778) & (g788) & (!g803)) + ((!g433) & (g468) & (!g777) & (g778) & (!g788) & (!g803)) + ((!g433) & (g468) & (!g777) & (g778) & (g788) & (!g803)) + ((!g433) & (g468) & (g777) & (!g778) & (!g788) & (!g803)) + ((!g433) & (g468) & (g777) & (!g778) & (!g788) & (g803)) + ((!g433) & (g468) & (g777) & (!g778) & (g788) & (g803)) + ((!g433) & (g468) & (g777) & (g778) & (!g788) & (g803)) + ((!g433) & (g468) & (g777) & (g778) & (g788) & (g803)) + ((g433) & (!g468) & (!g777) & (!g778) & (!g788) & (!g803)) + ((g433) & (!g468) & (!g777) & (!g778) & (g788) & (!g803)) + ((g433) & (!g468) & (!g777) & (g778) & (!g788) & (!g803)) + ((g433) & (!g468) & (g777) & (!g778) & (!g788) & (g803)) + ((g433) & (!g468) & (g777) & (!g778) & (g788) & (g803)) + ((g433) & (!g468) & (g777) & (g778) & (!g788) & (g803)) + ((g433) & (!g468) & (g777) & (g778) & (g788) & (!g803)) + ((g433) & (!g468) & (g777) & (g778) & (g788) & (g803)) + ((g433) & (g468) & (!g777) & (!g778) & (!g788) & (!g803)) + ((g433) & (g468) & (g777) & (!g778) & (!g788) & (g803)) + ((g433) & (g468) & (g777) & (!g778) & (g788) & (!g803)) + ((g433) & (g468) & (g777) & (!g778) & (g788) & (g803)) + ((g433) & (g468) & (g777) & (g778) & (!g788) & (!g803)) + ((g433) & (g468) & (g777) & (g778) & (!g788) & (g803)) + ((g433) & (g468) & (g777) & (g778) & (g788) & (!g803)) + ((g433) & (g468) & (g777) & (g778) & (g788) & (g803)));
	assign g824 = (((!g468) & (!g778) & (g788) & (!g803)) + ((!g468) & (g778) & (!g788) & (!g803)) + ((!g468) & (g778) & (!g788) & (g803)) + ((!g468) & (g778) & (g788) & (g803)) + ((g468) & (!g778) & (!g788) & (!g803)) + ((g468) & (g778) & (!g788) & (g803)) + ((g468) & (g778) & (g788) & (!g803)) + ((g468) & (g778) & (g788) & (g803)));
	assign g825 = (((!g515) & (!g553) & (!g780) & (g781) & (g787) & (!g803)) + ((!g515) & (!g553) & (g780) & (!g781) & (!g787) & (!g803)) + ((!g515) & (!g553) & (g780) & (!g781) & (!g787) & (g803)) + ((!g515) & (!g553) & (g780) & (!g781) & (g787) & (!g803)) + ((!g515) & (!g553) & (g780) & (!g781) & (g787) & (g803)) + ((!g515) & (!g553) & (g780) & (g781) & (!g787) & (!g803)) + ((!g515) & (!g553) & (g780) & (g781) & (!g787) & (g803)) + ((!g515) & (!g553) & (g780) & (g781) & (g787) & (g803)) + ((!g515) & (g553) & (!g780) & (!g781) & (g787) & (!g803)) + ((!g515) & (g553) & (!g780) & (g781) & (!g787) & (!g803)) + ((!g515) & (g553) & (!g780) & (g781) & (g787) & (!g803)) + ((!g515) & (g553) & (g780) & (!g781) & (!g787) & (!g803)) + ((!g515) & (g553) & (g780) & (!g781) & (!g787) & (g803)) + ((!g515) & (g553) & (g780) & (!g781) & (g787) & (g803)) + ((!g515) & (g553) & (g780) & (g781) & (!g787) & (g803)) + ((!g515) & (g553) & (g780) & (g781) & (g787) & (g803)) + ((g515) & (!g553) & (!g780) & (!g781) & (!g787) & (!g803)) + ((g515) & (!g553) & (!g780) & (!g781) & (g787) & (!g803)) + ((g515) & (!g553) & (!g780) & (g781) & (!g787) & (!g803)) + ((g515) & (!g553) & (g780) & (!g781) & (!g787) & (g803)) + ((g515) & (!g553) & (g780) & (!g781) & (g787) & (g803)) + ((g515) & (!g553) & (g780) & (g781) & (!g787) & (g803)) + ((g515) & (!g553) & (g780) & (g781) & (g787) & (!g803)) + ((g515) & (!g553) & (g780) & (g781) & (g787) & (g803)) + ((g515) & (g553) & (!g780) & (!g781) & (!g787) & (!g803)) + ((g515) & (g553) & (g780) & (!g781) & (!g787) & (g803)) + ((g515) & (g553) & (g780) & (!g781) & (g787) & (!g803)) + ((g515) & (g553) & (g780) & (!g781) & (g787) & (g803)) + ((g515) & (g553) & (g780) & (g781) & (!g787) & (!g803)) + ((g515) & (g553) & (g780) & (g781) & (!g787) & (g803)) + ((g515) & (g553) & (g780) & (g781) & (g787) & (!g803)) + ((g515) & (g553) & (g780) & (g781) & (g787) & (g803)));
	assign g826 = (((!g553) & (!g781) & (g787) & (!g803)) + ((!g553) & (g781) & (!g787) & (!g803)) + ((!g553) & (g781) & (!g787) & (g803)) + ((!g553) & (g781) & (g787) & (g803)) + ((g553) & (!g781) & (!g787) & (!g803)) + ((g553) & (g781) & (!g787) & (g803)) + ((g553) & (g781) & (g787) & (!g803)) + ((g553) & (g781) & (g787) & (g803)));
	assign g827 = (((!g604) & (!g645) & (!g783) & (g784) & (g786) & (!g803)) + ((!g604) & (!g645) & (g783) & (!g784) & (!g786) & (!g803)) + ((!g604) & (!g645) & (g783) & (!g784) & (!g786) & (g803)) + ((!g604) & (!g645) & (g783) & (!g784) & (g786) & (!g803)) + ((!g604) & (!g645) & (g783) & (!g784) & (g786) & (g803)) + ((!g604) & (!g645) & (g783) & (g784) & (!g786) & (!g803)) + ((!g604) & (!g645) & (g783) & (g784) & (!g786) & (g803)) + ((!g604) & (!g645) & (g783) & (g784) & (g786) & (g803)) + ((!g604) & (g645) & (!g783) & (!g784) & (g786) & (!g803)) + ((!g604) & (g645) & (!g783) & (g784) & (!g786) & (!g803)) + ((!g604) & (g645) & (!g783) & (g784) & (g786) & (!g803)) + ((!g604) & (g645) & (g783) & (!g784) & (!g786) & (!g803)) + ((!g604) & (g645) & (g783) & (!g784) & (!g786) & (g803)) + ((!g604) & (g645) & (g783) & (!g784) & (g786) & (g803)) + ((!g604) & (g645) & (g783) & (g784) & (!g786) & (g803)) + ((!g604) & (g645) & (g783) & (g784) & (g786) & (g803)) + ((g604) & (!g645) & (!g783) & (!g784) & (!g786) & (!g803)) + ((g604) & (!g645) & (!g783) & (!g784) & (g786) & (!g803)) + ((g604) & (!g645) & (!g783) & (g784) & (!g786) & (!g803)) + ((g604) & (!g645) & (g783) & (!g784) & (!g786) & (g803)) + ((g604) & (!g645) & (g783) & (!g784) & (g786) & (g803)) + ((g604) & (!g645) & (g783) & (g784) & (!g786) & (g803)) + ((g604) & (!g645) & (g783) & (g784) & (g786) & (!g803)) + ((g604) & (!g645) & (g783) & (g784) & (g786) & (g803)) + ((g604) & (g645) & (!g783) & (!g784) & (!g786) & (!g803)) + ((g604) & (g645) & (g783) & (!g784) & (!g786) & (g803)) + ((g604) & (g645) & (g783) & (!g784) & (g786) & (!g803)) + ((g604) & (g645) & (g783) & (!g784) & (g786) & (g803)) + ((g604) & (g645) & (g783) & (g784) & (!g786) & (!g803)) + ((g604) & (g645) & (g783) & (g784) & (!g786) & (g803)) + ((g604) & (g645) & (g783) & (g784) & (g786) & (!g803)) + ((g604) & (g645) & (g783) & (g784) & (g786) & (g803)));
	assign g828 = (((!g645) & (!g784) & (g786) & (!g803)) + ((!g645) & (g784) & (!g786) & (!g803)) + ((!g645) & (g784) & (!g786) & (g803)) + ((!g645) & (g784) & (g786) & (g803)) + ((g645) & (!g784) & (!g786) & (!g803)) + ((g645) & (g784) & (!g786) & (g803)) + ((g645) & (g784) & (g786) & (!g803)) + ((g645) & (g784) & (g786) & (g803)));
	assign g829 = (((!g700) & (!ax70x) & (!ax71x) & (!g744) & (!g785) & (g803)) + ((!g700) & (!ax70x) & (!ax71x) & (!g744) & (g785) & (!g803)) + ((!g700) & (!ax70x) & (!ax71x) & (!g744) & (g785) & (g803)) + ((!g700) & (!ax70x) & (!ax71x) & (g744) & (!g785) & (!g803)) + ((!g700) & (!ax70x) & (ax71x) & (!g744) & (!g785) & (!g803)) + ((!g700) & (!ax70x) & (ax71x) & (g744) & (!g785) & (g803)) + ((!g700) & (!ax70x) & (ax71x) & (g744) & (g785) & (!g803)) + ((!g700) & (!ax70x) & (ax71x) & (g744) & (g785) & (g803)) + ((!g700) & (ax70x) & (!ax71x) & (g744) & (!g785) & (!g803)) + ((!g700) & (ax70x) & (!ax71x) & (g744) & (g785) & (!g803)) + ((!g700) & (ax70x) & (ax71x) & (!g744) & (!g785) & (!g803)) + ((!g700) & (ax70x) & (ax71x) & (!g744) & (!g785) & (g803)) + ((!g700) & (ax70x) & (ax71x) & (!g744) & (g785) & (!g803)) + ((!g700) & (ax70x) & (ax71x) & (!g744) & (g785) & (g803)) + ((!g700) & (ax70x) & (ax71x) & (g744) & (!g785) & (g803)) + ((!g700) & (ax70x) & (ax71x) & (g744) & (g785) & (g803)) + ((g700) & (!ax70x) & (!ax71x) & (!g744) & (!g785) & (!g803)) + ((g700) & (!ax70x) & (!ax71x) & (!g744) & (!g785) & (g803)) + ((g700) & (!ax70x) & (!ax71x) & (!g744) & (g785) & (g803)) + ((g700) & (!ax70x) & (!ax71x) & (g744) & (g785) & (!g803)) + ((g700) & (!ax70x) & (ax71x) & (!g744) & (g785) & (!g803)) + ((g700) & (!ax70x) & (ax71x) & (g744) & (!g785) & (!g803)) + ((g700) & (!ax70x) & (ax71x) & (g744) & (!g785) & (g803)) + ((g700) & (!ax70x) & (ax71x) & (g744) & (g785) & (g803)) + ((g700) & (ax70x) & (!ax71x) & (!g744) & (!g785) & (!g803)) + ((g700) & (ax70x) & (!ax71x) & (!g744) & (g785) & (!g803)) + ((g700) & (ax70x) & (ax71x) & (!g744) & (!g785) & (g803)) + ((g700) & (ax70x) & (ax71x) & (!g744) & (g785) & (g803)) + ((g700) & (ax70x) & (ax71x) & (g744) & (!g785) & (!g803)) + ((g700) & (ax70x) & (ax71x) & (g744) & (!g785) & (g803)) + ((g700) & (ax70x) & (ax71x) & (g744) & (g785) & (!g803)) + ((g700) & (ax70x) & (ax71x) & (g744) & (g785) & (g803)));
	assign g830 = (((!ax70x) & (!g744) & (!g785) & (g803)) + ((!ax70x) & (!g744) & (g785) & (!g803)) + ((!ax70x) & (!g744) & (g785) & (g803)) + ((!ax70x) & (g744) & (g785) & (!g803)) + ((ax70x) & (!g744) & (!g785) & (!g803)) + ((ax70x) & (g744) & (!g785) & (!g803)) + ((ax70x) & (g744) & (!g785) & (g803)) + ((ax70x) & (g744) & (g785) & (g803)));
	assign g831 = (((!ax66x) & (!ax67x)));
	assign g832 = (((!g744) & (!ax68x) & (!ax69x) & (!g803) & (!g831)) + ((!g744) & (!ax68x) & (ax69x) & (g803) & (!g831)) + ((!g744) & (ax68x) & (ax69x) & (g803) & (!g831)) + ((!g744) & (ax68x) & (ax69x) & (g803) & (g831)) + ((g744) & (!ax68x) & (!ax69x) & (!g803) & (!g831)) + ((g744) & (!ax68x) & (!ax69x) & (!g803) & (g831)) + ((g744) & (!ax68x) & (!ax69x) & (g803) & (!g831)) + ((g744) & (!ax68x) & (ax69x) & (!g803) & (!g831)) + ((g744) & (!ax68x) & (ax69x) & (g803) & (!g831)) + ((g744) & (!ax68x) & (ax69x) & (g803) & (g831)) + ((g744) & (ax68x) & (!ax69x) & (g803) & (!g831)) + ((g744) & (ax68x) & (!ax69x) & (g803) & (g831)) + ((g744) & (ax68x) & (ax69x) & (!g803) & (!g831)) + ((g744) & (ax68x) & (ax69x) & (!g803) & (g831)) + ((g744) & (ax68x) & (ax69x) & (g803) & (!g831)) + ((g744) & (ax68x) & (ax69x) & (g803) & (g831)));
	assign g833 = (((!g645) & (!g700) & (g829) & (g830) & (g832)) + ((!g645) & (g700) & (g829) & (!g830) & (g832)) + ((!g645) & (g700) & (g829) & (g830) & (!g832)) + ((!g645) & (g700) & (g829) & (g830) & (g832)) + ((g645) & (!g700) & (!g829) & (g830) & (g832)) + ((g645) & (!g700) & (g829) & (!g830) & (!g832)) + ((g645) & (!g700) & (g829) & (!g830) & (g832)) + ((g645) & (!g700) & (g829) & (g830) & (!g832)) + ((g645) & (!g700) & (g829) & (g830) & (g832)) + ((g645) & (g700) & (!g829) & (!g830) & (g832)) + ((g645) & (g700) & (!g829) & (g830) & (!g832)) + ((g645) & (g700) & (!g829) & (g830) & (g832)) + ((g645) & (g700) & (g829) & (!g830) & (!g832)) + ((g645) & (g700) & (g829) & (!g830) & (g832)) + ((g645) & (g700) & (g829) & (g830) & (!g832)) + ((g645) & (g700) & (g829) & (g830) & (g832)));
	assign g834 = (((!g553) & (!g604) & (g827) & (g828) & (g833)) + ((!g553) & (g604) & (g827) & (!g828) & (g833)) + ((!g553) & (g604) & (g827) & (g828) & (!g833)) + ((!g553) & (g604) & (g827) & (g828) & (g833)) + ((g553) & (!g604) & (!g827) & (g828) & (g833)) + ((g553) & (!g604) & (g827) & (!g828) & (!g833)) + ((g553) & (!g604) & (g827) & (!g828) & (g833)) + ((g553) & (!g604) & (g827) & (g828) & (!g833)) + ((g553) & (!g604) & (g827) & (g828) & (g833)) + ((g553) & (g604) & (!g827) & (!g828) & (g833)) + ((g553) & (g604) & (!g827) & (g828) & (!g833)) + ((g553) & (g604) & (!g827) & (g828) & (g833)) + ((g553) & (g604) & (g827) & (!g828) & (!g833)) + ((g553) & (g604) & (g827) & (!g828) & (g833)) + ((g553) & (g604) & (g827) & (g828) & (!g833)) + ((g553) & (g604) & (g827) & (g828) & (g833)));
	assign g835 = (((!g468) & (!g515) & (g825) & (g826) & (g834)) + ((!g468) & (g515) & (g825) & (!g826) & (g834)) + ((!g468) & (g515) & (g825) & (g826) & (!g834)) + ((!g468) & (g515) & (g825) & (g826) & (g834)) + ((g468) & (!g515) & (!g825) & (g826) & (g834)) + ((g468) & (!g515) & (g825) & (!g826) & (!g834)) + ((g468) & (!g515) & (g825) & (!g826) & (g834)) + ((g468) & (!g515) & (g825) & (g826) & (!g834)) + ((g468) & (!g515) & (g825) & (g826) & (g834)) + ((g468) & (g515) & (!g825) & (!g826) & (g834)) + ((g468) & (g515) & (!g825) & (g826) & (!g834)) + ((g468) & (g515) & (!g825) & (g826) & (g834)) + ((g468) & (g515) & (g825) & (!g826) & (!g834)) + ((g468) & (g515) & (g825) & (!g826) & (g834)) + ((g468) & (g515) & (g825) & (g826) & (!g834)) + ((g468) & (g515) & (g825) & (g826) & (g834)));
	assign g836 = (((!g390) & (!g433) & (g823) & (g824) & (g835)) + ((!g390) & (g433) & (g823) & (!g824) & (g835)) + ((!g390) & (g433) & (g823) & (g824) & (!g835)) + ((!g390) & (g433) & (g823) & (g824) & (g835)) + ((g390) & (!g433) & (!g823) & (g824) & (g835)) + ((g390) & (!g433) & (g823) & (!g824) & (!g835)) + ((g390) & (!g433) & (g823) & (!g824) & (g835)) + ((g390) & (!g433) & (g823) & (g824) & (!g835)) + ((g390) & (!g433) & (g823) & (g824) & (g835)) + ((g390) & (g433) & (!g823) & (!g824) & (g835)) + ((g390) & (g433) & (!g823) & (g824) & (!g835)) + ((g390) & (g433) & (!g823) & (g824) & (g835)) + ((g390) & (g433) & (g823) & (!g824) & (!g835)) + ((g390) & (g433) & (g823) & (!g824) & (g835)) + ((g390) & (g433) & (g823) & (g824) & (!g835)) + ((g390) & (g433) & (g823) & (g824) & (g835)));
	assign g837 = (((!g319) & (!g358) & (g821) & (g822) & (g836)) + ((!g319) & (g358) & (g821) & (!g822) & (g836)) + ((!g319) & (g358) & (g821) & (g822) & (!g836)) + ((!g319) & (g358) & (g821) & (g822) & (g836)) + ((g319) & (!g358) & (!g821) & (g822) & (g836)) + ((g319) & (!g358) & (g821) & (!g822) & (!g836)) + ((g319) & (!g358) & (g821) & (!g822) & (g836)) + ((g319) & (!g358) & (g821) & (g822) & (!g836)) + ((g319) & (!g358) & (g821) & (g822) & (g836)) + ((g319) & (g358) & (!g821) & (!g822) & (g836)) + ((g319) & (g358) & (!g821) & (g822) & (!g836)) + ((g319) & (g358) & (!g821) & (g822) & (g836)) + ((g319) & (g358) & (g821) & (!g822) & (!g836)) + ((g319) & (g358) & (g821) & (!g822) & (g836)) + ((g319) & (g358) & (g821) & (g822) & (!g836)) + ((g319) & (g358) & (g821) & (g822) & (g836)));
	assign g838 = (((!g255) & (!g290) & (g819) & (g820) & (g837)) + ((!g255) & (g290) & (g819) & (!g820) & (g837)) + ((!g255) & (g290) & (g819) & (g820) & (!g837)) + ((!g255) & (g290) & (g819) & (g820) & (g837)) + ((g255) & (!g290) & (!g819) & (g820) & (g837)) + ((g255) & (!g290) & (g819) & (!g820) & (!g837)) + ((g255) & (!g290) & (g819) & (!g820) & (g837)) + ((g255) & (!g290) & (g819) & (g820) & (!g837)) + ((g255) & (!g290) & (g819) & (g820) & (g837)) + ((g255) & (g290) & (!g819) & (!g820) & (g837)) + ((g255) & (g290) & (!g819) & (g820) & (!g837)) + ((g255) & (g290) & (!g819) & (g820) & (g837)) + ((g255) & (g290) & (g819) & (!g820) & (!g837)) + ((g255) & (g290) & (g819) & (!g820) & (g837)) + ((g255) & (g290) & (g819) & (g820) & (!g837)) + ((g255) & (g290) & (g819) & (g820) & (g837)));
	assign g839 = (((!g198) & (!g229) & (g817) & (g818) & (g838)) + ((!g198) & (g229) & (g817) & (!g818) & (g838)) + ((!g198) & (g229) & (g817) & (g818) & (!g838)) + ((!g198) & (g229) & (g817) & (g818) & (g838)) + ((g198) & (!g229) & (!g817) & (g818) & (g838)) + ((g198) & (!g229) & (g817) & (!g818) & (!g838)) + ((g198) & (!g229) & (g817) & (!g818) & (g838)) + ((g198) & (!g229) & (g817) & (g818) & (!g838)) + ((g198) & (!g229) & (g817) & (g818) & (g838)) + ((g198) & (g229) & (!g817) & (!g818) & (g838)) + ((g198) & (g229) & (!g817) & (g818) & (!g838)) + ((g198) & (g229) & (!g817) & (g818) & (g838)) + ((g198) & (g229) & (g817) & (!g818) & (!g838)) + ((g198) & (g229) & (g817) & (!g818) & (g838)) + ((g198) & (g229) & (g817) & (g818) & (!g838)) + ((g198) & (g229) & (g817) & (g818) & (g838)));
	assign g840 = (((!g147) & (!g174) & (g815) & (g816) & (g839)) + ((!g147) & (g174) & (g815) & (!g816) & (g839)) + ((!g147) & (g174) & (g815) & (g816) & (!g839)) + ((!g147) & (g174) & (g815) & (g816) & (g839)) + ((g147) & (!g174) & (!g815) & (g816) & (g839)) + ((g147) & (!g174) & (g815) & (!g816) & (!g839)) + ((g147) & (!g174) & (g815) & (!g816) & (g839)) + ((g147) & (!g174) & (g815) & (g816) & (!g839)) + ((g147) & (!g174) & (g815) & (g816) & (g839)) + ((g147) & (g174) & (!g815) & (!g816) & (g839)) + ((g147) & (g174) & (!g815) & (g816) & (!g839)) + ((g147) & (g174) & (!g815) & (g816) & (g839)) + ((g147) & (g174) & (g815) & (!g816) & (!g839)) + ((g147) & (g174) & (g815) & (!g816) & (g839)) + ((g147) & (g174) & (g815) & (g816) & (!g839)) + ((g147) & (g174) & (g815) & (g816) & (g839)));
	assign g841 = (((!g104) & (!g127) & (g813) & (g814) & (g840)) + ((!g104) & (g127) & (g813) & (!g814) & (g840)) + ((!g104) & (g127) & (g813) & (g814) & (!g840)) + ((!g104) & (g127) & (g813) & (g814) & (g840)) + ((g104) & (!g127) & (!g813) & (g814) & (g840)) + ((g104) & (!g127) & (g813) & (!g814) & (!g840)) + ((g104) & (!g127) & (g813) & (!g814) & (g840)) + ((g104) & (!g127) & (g813) & (g814) & (!g840)) + ((g104) & (!g127) & (g813) & (g814) & (g840)) + ((g104) & (g127) & (!g813) & (!g814) & (g840)) + ((g104) & (g127) & (!g813) & (g814) & (!g840)) + ((g104) & (g127) & (!g813) & (g814) & (g840)) + ((g104) & (g127) & (g813) & (!g814) & (!g840)) + ((g104) & (g127) & (g813) & (!g814) & (g840)) + ((g104) & (g127) & (g813) & (g814) & (!g840)) + ((g104) & (g127) & (g813) & (g814) & (g840)));
	assign g842 = (((!g68) & (!g87) & (g811) & (g812) & (g841)) + ((!g68) & (g87) & (g811) & (!g812) & (g841)) + ((!g68) & (g87) & (g811) & (g812) & (!g841)) + ((!g68) & (g87) & (g811) & (g812) & (g841)) + ((g68) & (!g87) & (!g811) & (g812) & (g841)) + ((g68) & (!g87) & (g811) & (!g812) & (!g841)) + ((g68) & (!g87) & (g811) & (!g812) & (g841)) + ((g68) & (!g87) & (g811) & (g812) & (!g841)) + ((g68) & (!g87) & (g811) & (g812) & (g841)) + ((g68) & (g87) & (!g811) & (!g812) & (g841)) + ((g68) & (g87) & (!g811) & (g812) & (!g841)) + ((g68) & (g87) & (!g811) & (g812) & (g841)) + ((g68) & (g87) & (g811) & (!g812) & (!g841)) + ((g68) & (g87) & (g811) & (!g812) & (g841)) + ((g68) & (g87) & (g811) & (g812) & (!g841)) + ((g68) & (g87) & (g811) & (g812) & (g841)));
	assign g843 = (((!g39) & (!g54) & (g809) & (g810) & (g842)) + ((!g39) & (g54) & (g809) & (!g810) & (g842)) + ((!g39) & (g54) & (g809) & (g810) & (!g842)) + ((!g39) & (g54) & (g809) & (g810) & (g842)) + ((g39) & (!g54) & (!g809) & (g810) & (g842)) + ((g39) & (!g54) & (g809) & (!g810) & (!g842)) + ((g39) & (!g54) & (g809) & (!g810) & (g842)) + ((g39) & (!g54) & (g809) & (g810) & (!g842)) + ((g39) & (!g54) & (g809) & (g810) & (g842)) + ((g39) & (g54) & (!g809) & (!g810) & (g842)) + ((g39) & (g54) & (!g809) & (g810) & (!g842)) + ((g39) & (g54) & (!g809) & (g810) & (g842)) + ((g39) & (g54) & (g809) & (!g810) & (!g842)) + ((g39) & (g54) & (g809) & (!g810) & (g842)) + ((g39) & (g54) & (g809) & (g810) & (!g842)) + ((g39) & (g54) & (g809) & (g810) & (g842)));
	assign g844 = (((!g18) & (!g27) & (g807) & (g808) & (g843)) + ((!g18) & (g27) & (g807) & (!g808) & (g843)) + ((!g18) & (g27) & (g807) & (g808) & (!g843)) + ((!g18) & (g27) & (g807) & (g808) & (g843)) + ((g18) & (!g27) & (!g807) & (g808) & (g843)) + ((g18) & (!g27) & (g807) & (!g808) & (!g843)) + ((g18) & (!g27) & (g807) & (!g808) & (g843)) + ((g18) & (!g27) & (g807) & (g808) & (!g843)) + ((g18) & (!g27) & (g807) & (g808) & (g843)) + ((g18) & (g27) & (!g807) & (!g808) & (g843)) + ((g18) & (g27) & (!g807) & (g808) & (!g843)) + ((g18) & (g27) & (!g807) & (g808) & (g843)) + ((g18) & (g27) & (g807) & (!g808) & (!g843)) + ((g18) & (g27) & (g807) & (!g808) & (g843)) + ((g18) & (g27) & (g807) & (g808) & (!g843)) + ((g18) & (g27) & (g807) & (g808) & (g843)));
	assign g845 = (((!g2) & (!g8) & (g805) & (g806) & (g844)) + ((!g2) & (g8) & (g805) & (!g806) & (g844)) + ((!g2) & (g8) & (g805) & (g806) & (!g844)) + ((!g2) & (g8) & (g805) & (g806) & (g844)) + ((g2) & (!g8) & (!g805) & (g806) & (g844)) + ((g2) & (!g8) & (g805) & (!g806) & (!g844)) + ((g2) & (!g8) & (g805) & (!g806) & (g844)) + ((g2) & (!g8) & (g805) & (g806) & (!g844)) + ((g2) & (!g8) & (g805) & (g806) & (g844)) + ((g2) & (g8) & (!g805) & (!g806) & (g844)) + ((g2) & (g8) & (!g805) & (g806) & (!g844)) + ((g2) & (g8) & (!g805) & (g806) & (g844)) + ((g2) & (g8) & (g805) & (!g806) & (!g844)) + ((g2) & (g8) & (g805) & (!g806) & (g844)) + ((g2) & (g8) & (g805) & (g806) & (!g844)) + ((g2) & (g8) & (g805) & (g806) & (g844)));
	assign g846 = (((!g2) & (!g748) & (g798) & (!g803)) + ((!g2) & (g748) & (!g798) & (!g803)) + ((!g2) & (g748) & (!g798) & (g803)) + ((!g2) & (g748) & (g798) & (g803)) + ((g2) & (!g748) & (!g798) & (!g803)) + ((g2) & (g748) & (!g798) & (g803)) + ((g2) & (g748) & (g798) & (!g803)) + ((g2) & (g748) & (g798) & (g803)));
	assign g847 = (((!g1) & (!g745) & (!g799) & (!g801) & (g802)) + ((!g1) & (!g745) & (!g799) & (g801) & (!g802)) + ((!g1) & (!g745) & (!g799) & (g801) & (g802)) + ((!g1) & (g745) & (g799) & (!g801) & (!g802)) + ((!g1) & (g745) & (g799) & (!g801) & (g802)) + ((!g1) & (g745) & (g799) & (g801) & (!g802)) + ((!g1) & (g745) & (g799) & (g801) & (g802)) + ((g1) & (!g745) & (!g799) & (!g801) & (g802)) + ((g1) & (!g745) & (!g799) & (g801) & (g802)) + ((g1) & (g745) & (g799) & (!g801) & (!g802)) + ((g1) & (g745) & (g799) & (!g801) & (g802)) + ((g1) & (g745) & (g799) & (g801) & (!g802)) + ((g1) & (g745) & (g799) & (g801) & (g802)));
	assign g848 = (((!g4) & (!g1) & (!g804) & (!g845) & (!g846) & (g847)) + ((!g4) & (!g1) & (!g804) & (!g845) & (g846) & (!g847)) + ((!g4) & (!g1) & (!g804) & (!g845) & (g846) & (g847)) + ((!g4) & (!g1) & (!g804) & (g845) & (!g846) & (!g847)) + ((!g4) & (!g1) & (!g804) & (g845) & (!g846) & (g847)) + ((!g4) & (!g1) & (!g804) & (g845) & (g846) & (!g847)) + ((!g4) & (!g1) & (!g804) & (g845) & (g846) & (g847)) + ((!g4) & (!g1) & (g804) & (!g845) & (!g846) & (!g847)) + ((!g4) & (!g1) & (g804) & (!g845) & (!g846) & (g847)) + ((!g4) & (!g1) & (g804) & (!g845) & (g846) & (!g847)) + ((!g4) & (!g1) & (g804) & (!g845) & (g846) & (g847)) + ((!g4) & (!g1) & (g804) & (g845) & (!g846) & (!g847)) + ((!g4) & (!g1) & (g804) & (g845) & (!g846) & (g847)) + ((!g4) & (!g1) & (g804) & (g845) & (g846) & (!g847)) + ((!g4) & (!g1) & (g804) & (g845) & (g846) & (g847)) + ((g4) & (!g1) & (!g804) & (!g845) & (!g846) & (g847)) + ((g4) & (!g1) & (!g804) & (!g845) & (g846) & (g847)) + ((g4) & (!g1) & (!g804) & (g845) & (!g846) & (g847)) + ((g4) & (!g1) & (!g804) & (g845) & (g846) & (!g847)) + ((g4) & (!g1) & (!g804) & (g845) & (g846) & (g847)) + ((g4) & (!g1) & (g804) & (!g845) & (!g846) & (!g847)) + ((g4) & (!g1) & (g804) & (!g845) & (!g846) & (g847)) + ((g4) & (!g1) & (g804) & (!g845) & (g846) & (!g847)) + ((g4) & (!g1) & (g804) & (!g845) & (g846) & (g847)) + ((g4) & (!g1) & (g804) & (g845) & (!g846) & (!g847)) + ((g4) & (!g1) & (g804) & (g845) & (!g846) & (g847)) + ((g4) & (!g1) & (g804) & (g845) & (g846) & (!g847)) + ((g4) & (!g1) & (g804) & (g845) & (g846) & (g847)));
	assign g849 = (((g1) & (!g745) & (g799) & (g802)) + ((g1) & (g745) & (!g799) & (!g802)) + ((g1) & (g745) & (!g799) & (g802)));
	assign g850 = (((!g4) & (!g804) & (!g845) & (!g846) & (!g849)) + ((!g4) & (!g804) & (!g845) & (g846) & (!g849)) + ((!g4) & (!g804) & (g845) & (!g846) & (!g849)) + ((!g4) & (!g804) & (g845) & (g846) & (!g849)) + ((!g4) & (g804) & (!g845) & (!g846) & (!g849)) + ((g4) & (!g804) & (!g845) & (!g846) & (!g849)) + ((g4) & (!g804) & (!g845) & (g846) & (!g849)) + ((g4) & (!g804) & (g845) & (!g846) & (!g849)) + ((g4) & (!g804) & (g845) & (g846) & (!g849)) + ((g4) & (g804) & (!g845) & (!g846) & (!g849)) + ((g4) & (g804) & (!g845) & (g846) & (!g849)) + ((g4) & (g804) & (g845) & (!g846) & (!g849)));
	assign g851 = (((!g848) & (g850)));
	assign g852 = (((!g4) & (!g845) & (!g846) & (!g848) & (!g850)) + ((!g4) & (!g845) & (!g846) & (g848) & (!g850)) + ((!g4) & (!g845) & (!g846) & (g848) & (g850)) + ((!g4) & (!g845) & (g846) & (!g848) & (g850)) + ((!g4) & (g845) & (g846) & (!g848) & (!g850)) + ((!g4) & (g845) & (g846) & (!g848) & (g850)) + ((!g4) & (g845) & (g846) & (g848) & (!g850)) + ((!g4) & (g845) & (g846) & (g848) & (g850)) + ((g4) & (!g845) & (g846) & (!g848) & (!g850)) + ((g4) & (!g845) & (g846) & (!g848) & (g850)) + ((g4) & (!g845) & (g846) & (g848) & (!g850)) + ((g4) & (!g845) & (g846) & (g848) & (g850)) + ((g4) & (g845) & (!g846) & (!g848) & (!g850)) + ((g4) & (g845) & (!g846) & (g848) & (!g850)) + ((g4) & (g845) & (!g846) & (g848) & (g850)) + ((g4) & (g845) & (g846) & (!g848) & (g850)));
	assign g853 = (((!g8) & (!g806) & (g844) & (!g848) & (!g850)) + ((!g8) & (!g806) & (g844) & (g848) & (!g850)) + ((!g8) & (!g806) & (g844) & (g848) & (g850)) + ((!g8) & (g806) & (!g844) & (!g848) & (!g850)) + ((!g8) & (g806) & (!g844) & (!g848) & (g850)) + ((!g8) & (g806) & (!g844) & (g848) & (!g850)) + ((!g8) & (g806) & (!g844) & (g848) & (g850)) + ((!g8) & (g806) & (g844) & (!g848) & (g850)) + ((g8) & (!g806) & (!g844) & (!g848) & (!g850)) + ((g8) & (!g806) & (!g844) & (g848) & (!g850)) + ((g8) & (!g806) & (!g844) & (g848) & (g850)) + ((g8) & (g806) & (!g844) & (!g848) & (g850)) + ((g8) & (g806) & (g844) & (!g848) & (!g850)) + ((g8) & (g806) & (g844) & (!g848) & (g850)) + ((g8) & (g806) & (g844) & (g848) & (!g850)) + ((g8) & (g806) & (g844) & (g848) & (g850)));
	assign g854 = (((!g18) & (!g27) & (g808) & (g843)) + ((!g18) & (g27) & (!g808) & (g843)) + ((!g18) & (g27) & (g808) & (!g843)) + ((!g18) & (g27) & (g808) & (g843)) + ((g18) & (!g27) & (!g808) & (!g843)) + ((g18) & (!g27) & (!g808) & (g843)) + ((g18) & (!g27) & (g808) & (!g843)) + ((g18) & (g27) & (!g808) & (!g843)));
	assign g855 = (((!g807) & (!g848) & (!g850) & (g854)) + ((!g807) & (g848) & (!g850) & (g854)) + ((!g807) & (g848) & (g850) & (g854)) + ((g807) & (!g848) & (!g850) & (!g854)) + ((g807) & (!g848) & (g850) & (!g854)) + ((g807) & (!g848) & (g850) & (g854)) + ((g807) & (g848) & (!g850) & (!g854)) + ((g807) & (g848) & (g850) & (!g854)));
	assign g856 = (((!g27) & (!g808) & (g843) & (!g848) & (!g850)) + ((!g27) & (!g808) & (g843) & (g848) & (!g850)) + ((!g27) & (!g808) & (g843) & (g848) & (g850)) + ((!g27) & (g808) & (!g843) & (!g848) & (!g850)) + ((!g27) & (g808) & (!g843) & (!g848) & (g850)) + ((!g27) & (g808) & (!g843) & (g848) & (!g850)) + ((!g27) & (g808) & (!g843) & (g848) & (g850)) + ((!g27) & (g808) & (g843) & (!g848) & (g850)) + ((g27) & (!g808) & (!g843) & (!g848) & (!g850)) + ((g27) & (!g808) & (!g843) & (g848) & (!g850)) + ((g27) & (!g808) & (!g843) & (g848) & (g850)) + ((g27) & (g808) & (!g843) & (!g848) & (g850)) + ((g27) & (g808) & (g843) & (!g848) & (!g850)) + ((g27) & (g808) & (g843) & (!g848) & (g850)) + ((g27) & (g808) & (g843) & (g848) & (!g850)) + ((g27) & (g808) & (g843) & (g848) & (g850)));
	assign g857 = (((!g39) & (!g54) & (g810) & (g842)) + ((!g39) & (g54) & (!g810) & (g842)) + ((!g39) & (g54) & (g810) & (!g842)) + ((!g39) & (g54) & (g810) & (g842)) + ((g39) & (!g54) & (!g810) & (!g842)) + ((g39) & (!g54) & (!g810) & (g842)) + ((g39) & (!g54) & (g810) & (!g842)) + ((g39) & (g54) & (!g810) & (!g842)));
	assign g858 = (((!g809) & (!g848) & (!g850) & (g857)) + ((!g809) & (g848) & (!g850) & (g857)) + ((!g809) & (g848) & (g850) & (g857)) + ((g809) & (!g848) & (!g850) & (!g857)) + ((g809) & (!g848) & (g850) & (!g857)) + ((g809) & (!g848) & (g850) & (g857)) + ((g809) & (g848) & (!g850) & (!g857)) + ((g809) & (g848) & (g850) & (!g857)));
	assign g859 = (((!g54) & (!g810) & (g842) & (!g848) & (!g850)) + ((!g54) & (!g810) & (g842) & (g848) & (!g850)) + ((!g54) & (!g810) & (g842) & (g848) & (g850)) + ((!g54) & (g810) & (!g842) & (!g848) & (!g850)) + ((!g54) & (g810) & (!g842) & (!g848) & (g850)) + ((!g54) & (g810) & (!g842) & (g848) & (!g850)) + ((!g54) & (g810) & (!g842) & (g848) & (g850)) + ((!g54) & (g810) & (g842) & (!g848) & (g850)) + ((g54) & (!g810) & (!g842) & (!g848) & (!g850)) + ((g54) & (!g810) & (!g842) & (g848) & (!g850)) + ((g54) & (!g810) & (!g842) & (g848) & (g850)) + ((g54) & (g810) & (!g842) & (!g848) & (g850)) + ((g54) & (g810) & (g842) & (!g848) & (!g850)) + ((g54) & (g810) & (g842) & (!g848) & (g850)) + ((g54) & (g810) & (g842) & (g848) & (!g850)) + ((g54) & (g810) & (g842) & (g848) & (g850)));
	assign g860 = (((!g68) & (!g87) & (g812) & (g841)) + ((!g68) & (g87) & (!g812) & (g841)) + ((!g68) & (g87) & (g812) & (!g841)) + ((!g68) & (g87) & (g812) & (g841)) + ((g68) & (!g87) & (!g812) & (!g841)) + ((g68) & (!g87) & (!g812) & (g841)) + ((g68) & (!g87) & (g812) & (!g841)) + ((g68) & (g87) & (!g812) & (!g841)));
	assign g861 = (((!g811) & (!g848) & (!g850) & (g860)) + ((!g811) & (g848) & (!g850) & (g860)) + ((!g811) & (g848) & (g850) & (g860)) + ((g811) & (!g848) & (!g850) & (!g860)) + ((g811) & (!g848) & (g850) & (!g860)) + ((g811) & (!g848) & (g850) & (g860)) + ((g811) & (g848) & (!g850) & (!g860)) + ((g811) & (g848) & (g850) & (!g860)));
	assign g862 = (((!g87) & (!g812) & (g841) & (!g848) & (!g850)) + ((!g87) & (!g812) & (g841) & (g848) & (!g850)) + ((!g87) & (!g812) & (g841) & (g848) & (g850)) + ((!g87) & (g812) & (!g841) & (!g848) & (!g850)) + ((!g87) & (g812) & (!g841) & (!g848) & (g850)) + ((!g87) & (g812) & (!g841) & (g848) & (!g850)) + ((!g87) & (g812) & (!g841) & (g848) & (g850)) + ((!g87) & (g812) & (g841) & (!g848) & (g850)) + ((g87) & (!g812) & (!g841) & (!g848) & (!g850)) + ((g87) & (!g812) & (!g841) & (g848) & (!g850)) + ((g87) & (!g812) & (!g841) & (g848) & (g850)) + ((g87) & (g812) & (!g841) & (!g848) & (g850)) + ((g87) & (g812) & (g841) & (!g848) & (!g850)) + ((g87) & (g812) & (g841) & (!g848) & (g850)) + ((g87) & (g812) & (g841) & (g848) & (!g850)) + ((g87) & (g812) & (g841) & (g848) & (g850)));
	assign g863 = (((!g104) & (!g127) & (g814) & (g840)) + ((!g104) & (g127) & (!g814) & (g840)) + ((!g104) & (g127) & (g814) & (!g840)) + ((!g104) & (g127) & (g814) & (g840)) + ((g104) & (!g127) & (!g814) & (!g840)) + ((g104) & (!g127) & (!g814) & (g840)) + ((g104) & (!g127) & (g814) & (!g840)) + ((g104) & (g127) & (!g814) & (!g840)));
	assign g864 = (((!g813) & (!g848) & (!g850) & (g863)) + ((!g813) & (g848) & (!g850) & (g863)) + ((!g813) & (g848) & (g850) & (g863)) + ((g813) & (!g848) & (!g850) & (!g863)) + ((g813) & (!g848) & (g850) & (!g863)) + ((g813) & (!g848) & (g850) & (g863)) + ((g813) & (g848) & (!g850) & (!g863)) + ((g813) & (g848) & (g850) & (!g863)));
	assign g865 = (((!g127) & (!g814) & (g840) & (!g848) & (!g850)) + ((!g127) & (!g814) & (g840) & (g848) & (!g850)) + ((!g127) & (!g814) & (g840) & (g848) & (g850)) + ((!g127) & (g814) & (!g840) & (!g848) & (!g850)) + ((!g127) & (g814) & (!g840) & (!g848) & (g850)) + ((!g127) & (g814) & (!g840) & (g848) & (!g850)) + ((!g127) & (g814) & (!g840) & (g848) & (g850)) + ((!g127) & (g814) & (g840) & (!g848) & (g850)) + ((g127) & (!g814) & (!g840) & (!g848) & (!g850)) + ((g127) & (!g814) & (!g840) & (g848) & (!g850)) + ((g127) & (!g814) & (!g840) & (g848) & (g850)) + ((g127) & (g814) & (!g840) & (!g848) & (g850)) + ((g127) & (g814) & (g840) & (!g848) & (!g850)) + ((g127) & (g814) & (g840) & (!g848) & (g850)) + ((g127) & (g814) & (g840) & (g848) & (!g850)) + ((g127) & (g814) & (g840) & (g848) & (g850)));
	assign g866 = (((!g147) & (!g174) & (g816) & (g839)) + ((!g147) & (g174) & (!g816) & (g839)) + ((!g147) & (g174) & (g816) & (!g839)) + ((!g147) & (g174) & (g816) & (g839)) + ((g147) & (!g174) & (!g816) & (!g839)) + ((g147) & (!g174) & (!g816) & (g839)) + ((g147) & (!g174) & (g816) & (!g839)) + ((g147) & (g174) & (!g816) & (!g839)));
	assign g867 = (((!g815) & (!g848) & (!g850) & (g866)) + ((!g815) & (g848) & (!g850) & (g866)) + ((!g815) & (g848) & (g850) & (g866)) + ((g815) & (!g848) & (!g850) & (!g866)) + ((g815) & (!g848) & (g850) & (!g866)) + ((g815) & (!g848) & (g850) & (g866)) + ((g815) & (g848) & (!g850) & (!g866)) + ((g815) & (g848) & (g850) & (!g866)));
	assign g868 = (((!g174) & (!g816) & (g839) & (!g848) & (!g850)) + ((!g174) & (!g816) & (g839) & (g848) & (!g850)) + ((!g174) & (!g816) & (g839) & (g848) & (g850)) + ((!g174) & (g816) & (!g839) & (!g848) & (!g850)) + ((!g174) & (g816) & (!g839) & (!g848) & (g850)) + ((!g174) & (g816) & (!g839) & (g848) & (!g850)) + ((!g174) & (g816) & (!g839) & (g848) & (g850)) + ((!g174) & (g816) & (g839) & (!g848) & (g850)) + ((g174) & (!g816) & (!g839) & (!g848) & (!g850)) + ((g174) & (!g816) & (!g839) & (g848) & (!g850)) + ((g174) & (!g816) & (!g839) & (g848) & (g850)) + ((g174) & (g816) & (!g839) & (!g848) & (g850)) + ((g174) & (g816) & (g839) & (!g848) & (!g850)) + ((g174) & (g816) & (g839) & (!g848) & (g850)) + ((g174) & (g816) & (g839) & (g848) & (!g850)) + ((g174) & (g816) & (g839) & (g848) & (g850)));
	assign g869 = (((!g198) & (!g229) & (g818) & (g838)) + ((!g198) & (g229) & (!g818) & (g838)) + ((!g198) & (g229) & (g818) & (!g838)) + ((!g198) & (g229) & (g818) & (g838)) + ((g198) & (!g229) & (!g818) & (!g838)) + ((g198) & (!g229) & (!g818) & (g838)) + ((g198) & (!g229) & (g818) & (!g838)) + ((g198) & (g229) & (!g818) & (!g838)));
	assign g870 = (((!g817) & (!g848) & (!g850) & (g869)) + ((!g817) & (g848) & (!g850) & (g869)) + ((!g817) & (g848) & (g850) & (g869)) + ((g817) & (!g848) & (!g850) & (!g869)) + ((g817) & (!g848) & (g850) & (!g869)) + ((g817) & (!g848) & (g850) & (g869)) + ((g817) & (g848) & (!g850) & (!g869)) + ((g817) & (g848) & (g850) & (!g869)));
	assign g871 = (((!g229) & (!g818) & (g838) & (!g848) & (!g850)) + ((!g229) & (!g818) & (g838) & (g848) & (!g850)) + ((!g229) & (!g818) & (g838) & (g848) & (g850)) + ((!g229) & (g818) & (!g838) & (!g848) & (!g850)) + ((!g229) & (g818) & (!g838) & (!g848) & (g850)) + ((!g229) & (g818) & (!g838) & (g848) & (!g850)) + ((!g229) & (g818) & (!g838) & (g848) & (g850)) + ((!g229) & (g818) & (g838) & (!g848) & (g850)) + ((g229) & (!g818) & (!g838) & (!g848) & (!g850)) + ((g229) & (!g818) & (!g838) & (g848) & (!g850)) + ((g229) & (!g818) & (!g838) & (g848) & (g850)) + ((g229) & (g818) & (!g838) & (!g848) & (g850)) + ((g229) & (g818) & (g838) & (!g848) & (!g850)) + ((g229) & (g818) & (g838) & (!g848) & (g850)) + ((g229) & (g818) & (g838) & (g848) & (!g850)) + ((g229) & (g818) & (g838) & (g848) & (g850)));
	assign g872 = (((!g255) & (!g290) & (g820) & (g837)) + ((!g255) & (g290) & (!g820) & (g837)) + ((!g255) & (g290) & (g820) & (!g837)) + ((!g255) & (g290) & (g820) & (g837)) + ((g255) & (!g290) & (!g820) & (!g837)) + ((g255) & (!g290) & (!g820) & (g837)) + ((g255) & (!g290) & (g820) & (!g837)) + ((g255) & (g290) & (!g820) & (!g837)));
	assign g873 = (((!g819) & (!g848) & (!g850) & (g872)) + ((!g819) & (g848) & (!g850) & (g872)) + ((!g819) & (g848) & (g850) & (g872)) + ((g819) & (!g848) & (!g850) & (!g872)) + ((g819) & (!g848) & (g850) & (!g872)) + ((g819) & (!g848) & (g850) & (g872)) + ((g819) & (g848) & (!g850) & (!g872)) + ((g819) & (g848) & (g850) & (!g872)));
	assign g874 = (((!g290) & (!g820) & (g837) & (!g848) & (!g850)) + ((!g290) & (!g820) & (g837) & (g848) & (!g850)) + ((!g290) & (!g820) & (g837) & (g848) & (g850)) + ((!g290) & (g820) & (!g837) & (!g848) & (!g850)) + ((!g290) & (g820) & (!g837) & (!g848) & (g850)) + ((!g290) & (g820) & (!g837) & (g848) & (!g850)) + ((!g290) & (g820) & (!g837) & (g848) & (g850)) + ((!g290) & (g820) & (g837) & (!g848) & (g850)) + ((g290) & (!g820) & (!g837) & (!g848) & (!g850)) + ((g290) & (!g820) & (!g837) & (g848) & (!g850)) + ((g290) & (!g820) & (!g837) & (g848) & (g850)) + ((g290) & (g820) & (!g837) & (!g848) & (g850)) + ((g290) & (g820) & (g837) & (!g848) & (!g850)) + ((g290) & (g820) & (g837) & (!g848) & (g850)) + ((g290) & (g820) & (g837) & (g848) & (!g850)) + ((g290) & (g820) & (g837) & (g848) & (g850)));
	assign g875 = (((!g319) & (!g358) & (g822) & (g836)) + ((!g319) & (g358) & (!g822) & (g836)) + ((!g319) & (g358) & (g822) & (!g836)) + ((!g319) & (g358) & (g822) & (g836)) + ((g319) & (!g358) & (!g822) & (!g836)) + ((g319) & (!g358) & (!g822) & (g836)) + ((g319) & (!g358) & (g822) & (!g836)) + ((g319) & (g358) & (!g822) & (!g836)));
	assign g876 = (((!g821) & (!g848) & (!g850) & (g875)) + ((!g821) & (g848) & (!g850) & (g875)) + ((!g821) & (g848) & (g850) & (g875)) + ((g821) & (!g848) & (!g850) & (!g875)) + ((g821) & (!g848) & (g850) & (!g875)) + ((g821) & (!g848) & (g850) & (g875)) + ((g821) & (g848) & (!g850) & (!g875)) + ((g821) & (g848) & (g850) & (!g875)));
	assign g877 = (((!g358) & (!g822) & (g836) & (!g848) & (!g850)) + ((!g358) & (!g822) & (g836) & (g848) & (!g850)) + ((!g358) & (!g822) & (g836) & (g848) & (g850)) + ((!g358) & (g822) & (!g836) & (!g848) & (!g850)) + ((!g358) & (g822) & (!g836) & (!g848) & (g850)) + ((!g358) & (g822) & (!g836) & (g848) & (!g850)) + ((!g358) & (g822) & (!g836) & (g848) & (g850)) + ((!g358) & (g822) & (g836) & (!g848) & (g850)) + ((g358) & (!g822) & (!g836) & (!g848) & (!g850)) + ((g358) & (!g822) & (!g836) & (g848) & (!g850)) + ((g358) & (!g822) & (!g836) & (g848) & (g850)) + ((g358) & (g822) & (!g836) & (!g848) & (g850)) + ((g358) & (g822) & (g836) & (!g848) & (!g850)) + ((g358) & (g822) & (g836) & (!g848) & (g850)) + ((g358) & (g822) & (g836) & (g848) & (!g850)) + ((g358) & (g822) & (g836) & (g848) & (g850)));
	assign g878 = (((!g390) & (!g433) & (g824) & (g835)) + ((!g390) & (g433) & (!g824) & (g835)) + ((!g390) & (g433) & (g824) & (!g835)) + ((!g390) & (g433) & (g824) & (g835)) + ((g390) & (!g433) & (!g824) & (!g835)) + ((g390) & (!g433) & (!g824) & (g835)) + ((g390) & (!g433) & (g824) & (!g835)) + ((g390) & (g433) & (!g824) & (!g835)));
	assign g879 = (((!g823) & (!g848) & (!g850) & (g878)) + ((!g823) & (g848) & (!g850) & (g878)) + ((!g823) & (g848) & (g850) & (g878)) + ((g823) & (!g848) & (!g850) & (!g878)) + ((g823) & (!g848) & (g850) & (!g878)) + ((g823) & (!g848) & (g850) & (g878)) + ((g823) & (g848) & (!g850) & (!g878)) + ((g823) & (g848) & (g850) & (!g878)));
	assign g880 = (((!g433) & (!g824) & (g835) & (!g848) & (!g850)) + ((!g433) & (!g824) & (g835) & (g848) & (!g850)) + ((!g433) & (!g824) & (g835) & (g848) & (g850)) + ((!g433) & (g824) & (!g835) & (!g848) & (!g850)) + ((!g433) & (g824) & (!g835) & (!g848) & (g850)) + ((!g433) & (g824) & (!g835) & (g848) & (!g850)) + ((!g433) & (g824) & (!g835) & (g848) & (g850)) + ((!g433) & (g824) & (g835) & (!g848) & (g850)) + ((g433) & (!g824) & (!g835) & (!g848) & (!g850)) + ((g433) & (!g824) & (!g835) & (g848) & (!g850)) + ((g433) & (!g824) & (!g835) & (g848) & (g850)) + ((g433) & (g824) & (!g835) & (!g848) & (g850)) + ((g433) & (g824) & (g835) & (!g848) & (!g850)) + ((g433) & (g824) & (g835) & (!g848) & (g850)) + ((g433) & (g824) & (g835) & (g848) & (!g850)) + ((g433) & (g824) & (g835) & (g848) & (g850)));
	assign g881 = (((!g468) & (!g515) & (g826) & (g834)) + ((!g468) & (g515) & (!g826) & (g834)) + ((!g468) & (g515) & (g826) & (!g834)) + ((!g468) & (g515) & (g826) & (g834)) + ((g468) & (!g515) & (!g826) & (!g834)) + ((g468) & (!g515) & (!g826) & (g834)) + ((g468) & (!g515) & (g826) & (!g834)) + ((g468) & (g515) & (!g826) & (!g834)));
	assign g882 = (((!g825) & (!g848) & (!g850) & (g881)) + ((!g825) & (g848) & (!g850) & (g881)) + ((!g825) & (g848) & (g850) & (g881)) + ((g825) & (!g848) & (!g850) & (!g881)) + ((g825) & (!g848) & (g850) & (!g881)) + ((g825) & (!g848) & (g850) & (g881)) + ((g825) & (g848) & (!g850) & (!g881)) + ((g825) & (g848) & (g850) & (!g881)));
	assign g883 = (((!g515) & (!g826) & (g834) & (!g848) & (!g850)) + ((!g515) & (!g826) & (g834) & (g848) & (!g850)) + ((!g515) & (!g826) & (g834) & (g848) & (g850)) + ((!g515) & (g826) & (!g834) & (!g848) & (!g850)) + ((!g515) & (g826) & (!g834) & (!g848) & (g850)) + ((!g515) & (g826) & (!g834) & (g848) & (!g850)) + ((!g515) & (g826) & (!g834) & (g848) & (g850)) + ((!g515) & (g826) & (g834) & (!g848) & (g850)) + ((g515) & (!g826) & (!g834) & (!g848) & (!g850)) + ((g515) & (!g826) & (!g834) & (g848) & (!g850)) + ((g515) & (!g826) & (!g834) & (g848) & (g850)) + ((g515) & (g826) & (!g834) & (!g848) & (g850)) + ((g515) & (g826) & (g834) & (!g848) & (!g850)) + ((g515) & (g826) & (g834) & (!g848) & (g850)) + ((g515) & (g826) & (g834) & (g848) & (!g850)) + ((g515) & (g826) & (g834) & (g848) & (g850)));
	assign g884 = (((!g553) & (!g604) & (g828) & (g833)) + ((!g553) & (g604) & (!g828) & (g833)) + ((!g553) & (g604) & (g828) & (!g833)) + ((!g553) & (g604) & (g828) & (g833)) + ((g553) & (!g604) & (!g828) & (!g833)) + ((g553) & (!g604) & (!g828) & (g833)) + ((g553) & (!g604) & (g828) & (!g833)) + ((g553) & (g604) & (!g828) & (!g833)));
	assign g885 = (((!g827) & (!g848) & (!g850) & (g884)) + ((!g827) & (g848) & (!g850) & (g884)) + ((!g827) & (g848) & (g850) & (g884)) + ((g827) & (!g848) & (!g850) & (!g884)) + ((g827) & (!g848) & (g850) & (!g884)) + ((g827) & (!g848) & (g850) & (g884)) + ((g827) & (g848) & (!g850) & (!g884)) + ((g827) & (g848) & (g850) & (!g884)));
	assign g886 = (((!g604) & (!g828) & (g833) & (!g848) & (!g850)) + ((!g604) & (!g828) & (g833) & (g848) & (!g850)) + ((!g604) & (!g828) & (g833) & (g848) & (g850)) + ((!g604) & (g828) & (!g833) & (!g848) & (!g850)) + ((!g604) & (g828) & (!g833) & (!g848) & (g850)) + ((!g604) & (g828) & (!g833) & (g848) & (!g850)) + ((!g604) & (g828) & (!g833) & (g848) & (g850)) + ((!g604) & (g828) & (g833) & (!g848) & (g850)) + ((g604) & (!g828) & (!g833) & (!g848) & (!g850)) + ((g604) & (!g828) & (!g833) & (g848) & (!g850)) + ((g604) & (!g828) & (!g833) & (g848) & (g850)) + ((g604) & (g828) & (!g833) & (!g848) & (g850)) + ((g604) & (g828) & (g833) & (!g848) & (!g850)) + ((g604) & (g828) & (g833) & (!g848) & (g850)) + ((g604) & (g828) & (g833) & (g848) & (!g850)) + ((g604) & (g828) & (g833) & (g848) & (g850)));
	assign g887 = (((!g645) & (!g700) & (g830) & (g832)) + ((!g645) & (g700) & (!g830) & (g832)) + ((!g645) & (g700) & (g830) & (!g832)) + ((!g645) & (g700) & (g830) & (g832)) + ((g645) & (!g700) & (!g830) & (!g832)) + ((g645) & (!g700) & (!g830) & (g832)) + ((g645) & (!g700) & (g830) & (!g832)) + ((g645) & (g700) & (!g830) & (!g832)));
	assign g888 = (((!g829) & (!g848) & (!g850) & (g887)) + ((!g829) & (g848) & (!g850) & (g887)) + ((!g829) & (g848) & (g850) & (g887)) + ((g829) & (!g848) & (!g850) & (!g887)) + ((g829) & (!g848) & (g850) & (!g887)) + ((g829) & (!g848) & (g850) & (g887)) + ((g829) & (g848) & (!g850) & (!g887)) + ((g829) & (g848) & (g850) & (!g887)));
	assign g889 = (((!g700) & (!g830) & (g832) & (!g848) & (!g850)) + ((!g700) & (!g830) & (g832) & (g848) & (!g850)) + ((!g700) & (!g830) & (g832) & (g848) & (g850)) + ((!g700) & (g830) & (!g832) & (!g848) & (!g850)) + ((!g700) & (g830) & (!g832) & (!g848) & (g850)) + ((!g700) & (g830) & (!g832) & (g848) & (!g850)) + ((!g700) & (g830) & (!g832) & (g848) & (g850)) + ((!g700) & (g830) & (g832) & (!g848) & (g850)) + ((g700) & (!g830) & (!g832) & (!g848) & (!g850)) + ((g700) & (!g830) & (!g832) & (g848) & (!g850)) + ((g700) & (!g830) & (!g832) & (g848) & (g850)) + ((g700) & (g830) & (!g832) & (!g848) & (g850)) + ((g700) & (g830) & (g832) & (!g848) & (!g850)) + ((g700) & (g830) & (g832) & (!g848) & (g850)) + ((g700) & (g830) & (g832) & (g848) & (!g850)) + ((g700) & (g830) & (g832) & (g848) & (g850)));
	assign g890 = (((!g744) & (!ax68x) & (!g803) & (g831)) + ((!g744) & (!ax68x) & (g803) & (g831)) + ((!g744) & (ax68x) & (!g803) & (!g831)) + ((!g744) & (ax68x) & (!g803) & (g831)) + ((g744) & (!ax68x) & (!g803) & (!g831)) + ((g744) & (!ax68x) & (g803) & (!g831)) + ((g744) & (ax68x) & (g803) & (!g831)) + ((g744) & (ax68x) & (g803) & (g831)));
	assign g891 = (((!ax68x) & (!ax69x) & (!g803) & (!g848) & (!g850) & (g890)) + ((!ax68x) & (!ax69x) & (!g803) & (!g848) & (g850) & (!g890)) + ((!ax68x) & (!ax69x) & (!g803) & (!g848) & (g850) & (g890)) + ((!ax68x) & (!ax69x) & (!g803) & (g848) & (!g850) & (g890)) + ((!ax68x) & (!ax69x) & (!g803) & (g848) & (g850) & (g890)) + ((!ax68x) & (!ax69x) & (g803) & (!g848) & (!g850) & (!g890)) + ((!ax68x) & (!ax69x) & (g803) & (g848) & (!g850) & (!g890)) + ((!ax68x) & (!ax69x) & (g803) & (g848) & (g850) & (!g890)) + ((!ax68x) & (ax69x) & (!g803) & (!g848) & (!g850) & (!g890)) + ((!ax68x) & (ax69x) & (!g803) & (g848) & (!g850) & (!g890)) + ((!ax68x) & (ax69x) & (!g803) & (g848) & (g850) & (!g890)) + ((!ax68x) & (ax69x) & (g803) & (!g848) & (!g850) & (g890)) + ((!ax68x) & (ax69x) & (g803) & (!g848) & (g850) & (!g890)) + ((!ax68x) & (ax69x) & (g803) & (!g848) & (g850) & (g890)) + ((!ax68x) & (ax69x) & (g803) & (g848) & (!g850) & (g890)) + ((!ax68x) & (ax69x) & (g803) & (g848) & (g850) & (g890)) + ((ax68x) & (!ax69x) & (!g803) & (!g848) & (!g850) & (!g890)) + ((ax68x) & (!ax69x) & (!g803) & (g848) & (!g850) & (!g890)) + ((ax68x) & (!ax69x) & (!g803) & (g848) & (g850) & (!g890)) + ((ax68x) & (!ax69x) & (g803) & (!g848) & (!g850) & (!g890)) + ((ax68x) & (!ax69x) & (g803) & (g848) & (!g850) & (!g890)) + ((ax68x) & (!ax69x) & (g803) & (g848) & (g850) & (!g890)) + ((ax68x) & (ax69x) & (!g803) & (!g848) & (!g850) & (g890)) + ((ax68x) & (ax69x) & (!g803) & (!g848) & (g850) & (!g890)) + ((ax68x) & (ax69x) & (!g803) & (!g848) & (g850) & (g890)) + ((ax68x) & (ax69x) & (!g803) & (g848) & (!g850) & (g890)) + ((ax68x) & (ax69x) & (!g803) & (g848) & (g850) & (g890)) + ((ax68x) & (ax69x) & (g803) & (!g848) & (!g850) & (g890)) + ((ax68x) & (ax69x) & (g803) & (!g848) & (g850) & (!g890)) + ((ax68x) & (ax69x) & (g803) & (!g848) & (g850) & (g890)) + ((ax68x) & (ax69x) & (g803) & (g848) & (!g850) & (g890)) + ((ax68x) & (ax69x) & (g803) & (g848) & (g850) & (g890)));
	assign g892 = (((!ax68x) & (!g803) & (!g831) & (!g848) & (g850)) + ((!ax68x) & (!g803) & (g831) & (!g848) & (!g850)) + ((!ax68x) & (!g803) & (g831) & (!g848) & (g850)) + ((!ax68x) & (!g803) & (g831) & (g848) & (!g850)) + ((!ax68x) & (!g803) & (g831) & (g848) & (g850)) + ((!ax68x) & (g803) & (g831) & (!g848) & (!g850)) + ((!ax68x) & (g803) & (g831) & (g848) & (!g850)) + ((!ax68x) & (g803) & (g831) & (g848) & (g850)) + ((ax68x) & (!g803) & (!g831) & (!g848) & (!g850)) + ((ax68x) & (!g803) & (!g831) & (g848) & (!g850)) + ((ax68x) & (!g803) & (!g831) & (g848) & (g850)) + ((ax68x) & (g803) & (!g831) & (!g848) & (!g850)) + ((ax68x) & (g803) & (!g831) & (!g848) & (g850)) + ((ax68x) & (g803) & (!g831) & (g848) & (!g850)) + ((ax68x) & (g803) & (!g831) & (g848) & (g850)) + ((ax68x) & (g803) & (g831) & (!g848) & (g850)));
	assign g893 = (((!ax64x) & (!ax65x)));
	assign g894 = (((!g803) & (!ax66x) & (!ax67x) & (!g848) & (!g850) & (!g893)) + ((!g803) & (!ax66x) & (!ax67x) & (g848) & (!g850) & (!g893)) + ((!g803) & (!ax66x) & (!ax67x) & (g848) & (g850) & (!g893)) + ((!g803) & (!ax66x) & (ax67x) & (!g848) & (g850) & (!g893)) + ((!g803) & (ax66x) & (ax67x) & (!g848) & (g850) & (!g893)) + ((!g803) & (ax66x) & (ax67x) & (!g848) & (g850) & (g893)) + ((g803) & (!ax66x) & (!ax67x) & (!g848) & (!g850) & (!g893)) + ((g803) & (!ax66x) & (!ax67x) & (!g848) & (!g850) & (g893)) + ((g803) & (!ax66x) & (!ax67x) & (!g848) & (g850) & (!g893)) + ((g803) & (!ax66x) & (!ax67x) & (g848) & (!g850) & (!g893)) + ((g803) & (!ax66x) & (!ax67x) & (g848) & (!g850) & (g893)) + ((g803) & (!ax66x) & (!ax67x) & (g848) & (g850) & (!g893)) + ((g803) & (!ax66x) & (!ax67x) & (g848) & (g850) & (g893)) + ((g803) & (!ax66x) & (ax67x) & (!g848) & (!g850) & (!g893)) + ((g803) & (!ax66x) & (ax67x) & (!g848) & (g850) & (!g893)) + ((g803) & (!ax66x) & (ax67x) & (!g848) & (g850) & (g893)) + ((g803) & (!ax66x) & (ax67x) & (g848) & (!g850) & (!g893)) + ((g803) & (!ax66x) & (ax67x) & (g848) & (g850) & (!g893)) + ((g803) & (ax66x) & (!ax67x) & (!g848) & (g850) & (!g893)) + ((g803) & (ax66x) & (!ax67x) & (!g848) & (g850) & (g893)) + ((g803) & (ax66x) & (ax67x) & (!g848) & (!g850) & (!g893)) + ((g803) & (ax66x) & (ax67x) & (!g848) & (!g850) & (g893)) + ((g803) & (ax66x) & (ax67x) & (!g848) & (g850) & (!g893)) + ((g803) & (ax66x) & (ax67x) & (!g848) & (g850) & (g893)) + ((g803) & (ax66x) & (ax67x) & (g848) & (!g850) & (!g893)) + ((g803) & (ax66x) & (ax67x) & (g848) & (!g850) & (g893)) + ((g803) & (ax66x) & (ax67x) & (g848) & (g850) & (!g893)) + ((g803) & (ax66x) & (ax67x) & (g848) & (g850) & (g893)));
	assign g895 = (((!g700) & (!g744) & (g891) & (g892) & (g894)) + ((!g700) & (g744) & (g891) & (!g892) & (g894)) + ((!g700) & (g744) & (g891) & (g892) & (!g894)) + ((!g700) & (g744) & (g891) & (g892) & (g894)) + ((g700) & (!g744) & (!g891) & (g892) & (g894)) + ((g700) & (!g744) & (g891) & (!g892) & (!g894)) + ((g700) & (!g744) & (g891) & (!g892) & (g894)) + ((g700) & (!g744) & (g891) & (g892) & (!g894)) + ((g700) & (!g744) & (g891) & (g892) & (g894)) + ((g700) & (g744) & (!g891) & (!g892) & (g894)) + ((g700) & (g744) & (!g891) & (g892) & (!g894)) + ((g700) & (g744) & (!g891) & (g892) & (g894)) + ((g700) & (g744) & (g891) & (!g892) & (!g894)) + ((g700) & (g744) & (g891) & (!g892) & (g894)) + ((g700) & (g744) & (g891) & (g892) & (!g894)) + ((g700) & (g744) & (g891) & (g892) & (g894)));
	assign g896 = (((!g604) & (!g645) & (g888) & (g889) & (g895)) + ((!g604) & (g645) & (g888) & (!g889) & (g895)) + ((!g604) & (g645) & (g888) & (g889) & (!g895)) + ((!g604) & (g645) & (g888) & (g889) & (g895)) + ((g604) & (!g645) & (!g888) & (g889) & (g895)) + ((g604) & (!g645) & (g888) & (!g889) & (!g895)) + ((g604) & (!g645) & (g888) & (!g889) & (g895)) + ((g604) & (!g645) & (g888) & (g889) & (!g895)) + ((g604) & (!g645) & (g888) & (g889) & (g895)) + ((g604) & (g645) & (!g888) & (!g889) & (g895)) + ((g604) & (g645) & (!g888) & (g889) & (!g895)) + ((g604) & (g645) & (!g888) & (g889) & (g895)) + ((g604) & (g645) & (g888) & (!g889) & (!g895)) + ((g604) & (g645) & (g888) & (!g889) & (g895)) + ((g604) & (g645) & (g888) & (g889) & (!g895)) + ((g604) & (g645) & (g888) & (g889) & (g895)));
	assign g897 = (((!g515) & (!g553) & (g885) & (g886) & (g896)) + ((!g515) & (g553) & (g885) & (!g886) & (g896)) + ((!g515) & (g553) & (g885) & (g886) & (!g896)) + ((!g515) & (g553) & (g885) & (g886) & (g896)) + ((g515) & (!g553) & (!g885) & (g886) & (g896)) + ((g515) & (!g553) & (g885) & (!g886) & (!g896)) + ((g515) & (!g553) & (g885) & (!g886) & (g896)) + ((g515) & (!g553) & (g885) & (g886) & (!g896)) + ((g515) & (!g553) & (g885) & (g886) & (g896)) + ((g515) & (g553) & (!g885) & (!g886) & (g896)) + ((g515) & (g553) & (!g885) & (g886) & (!g896)) + ((g515) & (g553) & (!g885) & (g886) & (g896)) + ((g515) & (g553) & (g885) & (!g886) & (!g896)) + ((g515) & (g553) & (g885) & (!g886) & (g896)) + ((g515) & (g553) & (g885) & (g886) & (!g896)) + ((g515) & (g553) & (g885) & (g886) & (g896)));
	assign g898 = (((!g433) & (!g468) & (g882) & (g883) & (g897)) + ((!g433) & (g468) & (g882) & (!g883) & (g897)) + ((!g433) & (g468) & (g882) & (g883) & (!g897)) + ((!g433) & (g468) & (g882) & (g883) & (g897)) + ((g433) & (!g468) & (!g882) & (g883) & (g897)) + ((g433) & (!g468) & (g882) & (!g883) & (!g897)) + ((g433) & (!g468) & (g882) & (!g883) & (g897)) + ((g433) & (!g468) & (g882) & (g883) & (!g897)) + ((g433) & (!g468) & (g882) & (g883) & (g897)) + ((g433) & (g468) & (!g882) & (!g883) & (g897)) + ((g433) & (g468) & (!g882) & (g883) & (!g897)) + ((g433) & (g468) & (!g882) & (g883) & (g897)) + ((g433) & (g468) & (g882) & (!g883) & (!g897)) + ((g433) & (g468) & (g882) & (!g883) & (g897)) + ((g433) & (g468) & (g882) & (g883) & (!g897)) + ((g433) & (g468) & (g882) & (g883) & (g897)));
	assign g899 = (((!g358) & (!g390) & (g879) & (g880) & (g898)) + ((!g358) & (g390) & (g879) & (!g880) & (g898)) + ((!g358) & (g390) & (g879) & (g880) & (!g898)) + ((!g358) & (g390) & (g879) & (g880) & (g898)) + ((g358) & (!g390) & (!g879) & (g880) & (g898)) + ((g358) & (!g390) & (g879) & (!g880) & (!g898)) + ((g358) & (!g390) & (g879) & (!g880) & (g898)) + ((g358) & (!g390) & (g879) & (g880) & (!g898)) + ((g358) & (!g390) & (g879) & (g880) & (g898)) + ((g358) & (g390) & (!g879) & (!g880) & (g898)) + ((g358) & (g390) & (!g879) & (g880) & (!g898)) + ((g358) & (g390) & (!g879) & (g880) & (g898)) + ((g358) & (g390) & (g879) & (!g880) & (!g898)) + ((g358) & (g390) & (g879) & (!g880) & (g898)) + ((g358) & (g390) & (g879) & (g880) & (!g898)) + ((g358) & (g390) & (g879) & (g880) & (g898)));
	assign g900 = (((!g290) & (!g319) & (g876) & (g877) & (g899)) + ((!g290) & (g319) & (g876) & (!g877) & (g899)) + ((!g290) & (g319) & (g876) & (g877) & (!g899)) + ((!g290) & (g319) & (g876) & (g877) & (g899)) + ((g290) & (!g319) & (!g876) & (g877) & (g899)) + ((g290) & (!g319) & (g876) & (!g877) & (!g899)) + ((g290) & (!g319) & (g876) & (!g877) & (g899)) + ((g290) & (!g319) & (g876) & (g877) & (!g899)) + ((g290) & (!g319) & (g876) & (g877) & (g899)) + ((g290) & (g319) & (!g876) & (!g877) & (g899)) + ((g290) & (g319) & (!g876) & (g877) & (!g899)) + ((g290) & (g319) & (!g876) & (g877) & (g899)) + ((g290) & (g319) & (g876) & (!g877) & (!g899)) + ((g290) & (g319) & (g876) & (!g877) & (g899)) + ((g290) & (g319) & (g876) & (g877) & (!g899)) + ((g290) & (g319) & (g876) & (g877) & (g899)));
	assign g901 = (((!g229) & (!g255) & (g873) & (g874) & (g900)) + ((!g229) & (g255) & (g873) & (!g874) & (g900)) + ((!g229) & (g255) & (g873) & (g874) & (!g900)) + ((!g229) & (g255) & (g873) & (g874) & (g900)) + ((g229) & (!g255) & (!g873) & (g874) & (g900)) + ((g229) & (!g255) & (g873) & (!g874) & (!g900)) + ((g229) & (!g255) & (g873) & (!g874) & (g900)) + ((g229) & (!g255) & (g873) & (g874) & (!g900)) + ((g229) & (!g255) & (g873) & (g874) & (g900)) + ((g229) & (g255) & (!g873) & (!g874) & (g900)) + ((g229) & (g255) & (!g873) & (g874) & (!g900)) + ((g229) & (g255) & (!g873) & (g874) & (g900)) + ((g229) & (g255) & (g873) & (!g874) & (!g900)) + ((g229) & (g255) & (g873) & (!g874) & (g900)) + ((g229) & (g255) & (g873) & (g874) & (!g900)) + ((g229) & (g255) & (g873) & (g874) & (g900)));
	assign g902 = (((!g174) & (!g198) & (g870) & (g871) & (g901)) + ((!g174) & (g198) & (g870) & (!g871) & (g901)) + ((!g174) & (g198) & (g870) & (g871) & (!g901)) + ((!g174) & (g198) & (g870) & (g871) & (g901)) + ((g174) & (!g198) & (!g870) & (g871) & (g901)) + ((g174) & (!g198) & (g870) & (!g871) & (!g901)) + ((g174) & (!g198) & (g870) & (!g871) & (g901)) + ((g174) & (!g198) & (g870) & (g871) & (!g901)) + ((g174) & (!g198) & (g870) & (g871) & (g901)) + ((g174) & (g198) & (!g870) & (!g871) & (g901)) + ((g174) & (g198) & (!g870) & (g871) & (!g901)) + ((g174) & (g198) & (!g870) & (g871) & (g901)) + ((g174) & (g198) & (g870) & (!g871) & (!g901)) + ((g174) & (g198) & (g870) & (!g871) & (g901)) + ((g174) & (g198) & (g870) & (g871) & (!g901)) + ((g174) & (g198) & (g870) & (g871) & (g901)));
	assign g903 = (((!g127) & (!g147) & (g867) & (g868) & (g902)) + ((!g127) & (g147) & (g867) & (!g868) & (g902)) + ((!g127) & (g147) & (g867) & (g868) & (!g902)) + ((!g127) & (g147) & (g867) & (g868) & (g902)) + ((g127) & (!g147) & (!g867) & (g868) & (g902)) + ((g127) & (!g147) & (g867) & (!g868) & (!g902)) + ((g127) & (!g147) & (g867) & (!g868) & (g902)) + ((g127) & (!g147) & (g867) & (g868) & (!g902)) + ((g127) & (!g147) & (g867) & (g868) & (g902)) + ((g127) & (g147) & (!g867) & (!g868) & (g902)) + ((g127) & (g147) & (!g867) & (g868) & (!g902)) + ((g127) & (g147) & (!g867) & (g868) & (g902)) + ((g127) & (g147) & (g867) & (!g868) & (!g902)) + ((g127) & (g147) & (g867) & (!g868) & (g902)) + ((g127) & (g147) & (g867) & (g868) & (!g902)) + ((g127) & (g147) & (g867) & (g868) & (g902)));
	assign g904 = (((!g87) & (!g104) & (g864) & (g865) & (g903)) + ((!g87) & (g104) & (g864) & (!g865) & (g903)) + ((!g87) & (g104) & (g864) & (g865) & (!g903)) + ((!g87) & (g104) & (g864) & (g865) & (g903)) + ((g87) & (!g104) & (!g864) & (g865) & (g903)) + ((g87) & (!g104) & (g864) & (!g865) & (!g903)) + ((g87) & (!g104) & (g864) & (!g865) & (g903)) + ((g87) & (!g104) & (g864) & (g865) & (!g903)) + ((g87) & (!g104) & (g864) & (g865) & (g903)) + ((g87) & (g104) & (!g864) & (!g865) & (g903)) + ((g87) & (g104) & (!g864) & (g865) & (!g903)) + ((g87) & (g104) & (!g864) & (g865) & (g903)) + ((g87) & (g104) & (g864) & (!g865) & (!g903)) + ((g87) & (g104) & (g864) & (!g865) & (g903)) + ((g87) & (g104) & (g864) & (g865) & (!g903)) + ((g87) & (g104) & (g864) & (g865) & (g903)));
	assign g905 = (((!g54) & (!g68) & (g861) & (g862) & (g904)) + ((!g54) & (g68) & (g861) & (!g862) & (g904)) + ((!g54) & (g68) & (g861) & (g862) & (!g904)) + ((!g54) & (g68) & (g861) & (g862) & (g904)) + ((g54) & (!g68) & (!g861) & (g862) & (g904)) + ((g54) & (!g68) & (g861) & (!g862) & (!g904)) + ((g54) & (!g68) & (g861) & (!g862) & (g904)) + ((g54) & (!g68) & (g861) & (g862) & (!g904)) + ((g54) & (!g68) & (g861) & (g862) & (g904)) + ((g54) & (g68) & (!g861) & (!g862) & (g904)) + ((g54) & (g68) & (!g861) & (g862) & (!g904)) + ((g54) & (g68) & (!g861) & (g862) & (g904)) + ((g54) & (g68) & (g861) & (!g862) & (!g904)) + ((g54) & (g68) & (g861) & (!g862) & (g904)) + ((g54) & (g68) & (g861) & (g862) & (!g904)) + ((g54) & (g68) & (g861) & (g862) & (g904)));
	assign g906 = (((!g27) & (!g39) & (g858) & (g859) & (g905)) + ((!g27) & (g39) & (g858) & (!g859) & (g905)) + ((!g27) & (g39) & (g858) & (g859) & (!g905)) + ((!g27) & (g39) & (g858) & (g859) & (g905)) + ((g27) & (!g39) & (!g858) & (g859) & (g905)) + ((g27) & (!g39) & (g858) & (!g859) & (!g905)) + ((g27) & (!g39) & (g858) & (!g859) & (g905)) + ((g27) & (!g39) & (g858) & (g859) & (!g905)) + ((g27) & (!g39) & (g858) & (g859) & (g905)) + ((g27) & (g39) & (!g858) & (!g859) & (g905)) + ((g27) & (g39) & (!g858) & (g859) & (!g905)) + ((g27) & (g39) & (!g858) & (g859) & (g905)) + ((g27) & (g39) & (g858) & (!g859) & (!g905)) + ((g27) & (g39) & (g858) & (!g859) & (g905)) + ((g27) & (g39) & (g858) & (g859) & (!g905)) + ((g27) & (g39) & (g858) & (g859) & (g905)));
	assign g907 = (((!g8) & (!g18) & (g855) & (g856) & (g906)) + ((!g8) & (g18) & (g855) & (!g856) & (g906)) + ((!g8) & (g18) & (g855) & (g856) & (!g906)) + ((!g8) & (g18) & (g855) & (g856) & (g906)) + ((g8) & (!g18) & (!g855) & (g856) & (g906)) + ((g8) & (!g18) & (g855) & (!g856) & (!g906)) + ((g8) & (!g18) & (g855) & (!g856) & (g906)) + ((g8) & (!g18) & (g855) & (g856) & (!g906)) + ((g8) & (!g18) & (g855) & (g856) & (g906)) + ((g8) & (g18) & (!g855) & (!g856) & (g906)) + ((g8) & (g18) & (!g855) & (g856) & (!g906)) + ((g8) & (g18) & (!g855) & (g856) & (g906)) + ((g8) & (g18) & (g855) & (!g856) & (!g906)) + ((g8) & (g18) & (g855) & (!g856) & (g906)) + ((g8) & (g18) & (g855) & (g856) & (!g906)) + ((g8) & (g18) & (g855) & (g856) & (g906)));
	assign g908 = (((!g2) & (!g8) & (g806) & (g844)) + ((!g2) & (g8) & (!g806) & (g844)) + ((!g2) & (g8) & (g806) & (!g844)) + ((!g2) & (g8) & (g806) & (g844)) + ((g2) & (!g8) & (!g806) & (!g844)) + ((g2) & (!g8) & (!g806) & (g844)) + ((g2) & (!g8) & (g806) & (!g844)) + ((g2) & (g8) & (!g806) & (!g844)));
	assign g909 = (((!g805) & (!g848) & (!g850) & (g908)) + ((!g805) & (g848) & (!g850) & (g908)) + ((!g805) & (g848) & (g850) & (g908)) + ((g805) & (!g848) & (!g850) & (!g908)) + ((g805) & (!g848) & (g850) & (!g908)) + ((g805) & (!g848) & (g850) & (g908)) + ((g805) & (g848) & (!g850) & (!g908)) + ((g805) & (g848) & (g850) & (!g908)));
	assign g910 = (((!g4) & (!g2) & (!g853) & (!g907) & (g909)) + ((!g4) & (!g2) & (!g853) & (g907) & (g909)) + ((!g4) & (!g2) & (g853) & (!g907) & (g909)) + ((!g4) & (!g2) & (g853) & (g907) & (!g909)) + ((!g4) & (!g2) & (g853) & (g907) & (g909)) + ((!g4) & (g2) & (!g853) & (!g907) & (g909)) + ((!g4) & (g2) & (!g853) & (g907) & (!g909)) + ((!g4) & (g2) & (!g853) & (g907) & (g909)) + ((!g4) & (g2) & (g853) & (!g907) & (!g909)) + ((!g4) & (g2) & (g853) & (!g907) & (g909)) + ((!g4) & (g2) & (g853) & (g907) & (!g909)) + ((!g4) & (g2) & (g853) & (g907) & (g909)) + ((g4) & (!g2) & (g853) & (g907) & (g909)) + ((g4) & (g2) & (!g853) & (g907) & (g909)) + ((g4) & (g2) & (g853) & (!g907) & (g909)) + ((g4) & (g2) & (g853) & (g907) & (g909)));
	assign g911 = (((!g4) & (!g845) & (g846)) + ((!g4) & (g845) & (!g846)) + ((!g4) & (g845) & (g846)) + ((g4) & (g845) & (g846)));
	assign g912 = (((!g804) & (!g911) & (!g848) & (!g850)) + ((!g804) & (!g911) & (g848) & (!g850)) + ((!g804) & (!g911) & (g848) & (g850)) + ((g804) & (g911) & (!g848) & (!g850)) + ((g804) & (g911) & (!g848) & (g850)) + ((g804) & (g911) & (g848) & (!g850)) + ((g804) & (g911) & (g848) & (g850)));
	assign g913 = (((!g1) & (g804) & (!g911) & (!g848) & (!g849)) + ((g1) & (!g804) & (g911) & (!g848) & (g849)) + ((g1) & (!g804) & (g911) & (g848) & (g849)) + ((g1) & (g804) & (!g911) & (!g848) & (!g849)) + ((g1) & (g804) & (!g911) & (!g848) & (g849)) + ((g1) & (g804) & (!g911) & (g848) & (!g849)) + ((g1) & (g804) & (!g911) & (g848) & (g849)));
	assign g914 = (((!g1) & (!g852) & (!g910) & (!g912) & (!g913)) + ((g1) & (!g852) & (!g910) & (!g912) & (!g913)) + ((g1) & (!g852) & (!g910) & (g912) & (!g913)) + ((g1) & (!g852) & (g910) & (!g912) & (!g913)) + ((g1) & (!g852) & (g910) & (g912) & (!g913)) + ((g1) & (g852) & (!g910) & (!g912) & (!g913)) + ((g1) & (g852) & (!g910) & (g912) & (!g913)));
	assign g915 = (((!ax62x) & (!ax63x)));
	assign g916 = (((g1) & (!g852) & (g910) & (g913)) + ((g1) & (g852) & (!g910) & (!g913)) + ((g1) & (g852) & (!g910) & (g913)));
	assign g917 = (((!g4) & (!g2) & (!g853) & (!g907) & (!g909) & (!g914)) + ((!g4) & (!g2) & (!g853) & (!g907) & (g909) & (g914)) + ((!g4) & (!g2) & (!g853) & (g907) & (!g909) & (!g914)) + ((!g4) & (!g2) & (!g853) & (g907) & (g909) & (g914)) + ((!g4) & (!g2) & (g853) & (!g907) & (!g909) & (!g914)) + ((!g4) & (!g2) & (g853) & (!g907) & (g909) & (g914)) + ((!g4) & (!g2) & (g853) & (g907) & (g909) & (!g914)) + ((!g4) & (!g2) & (g853) & (g907) & (g909) & (g914)) + ((!g4) & (g2) & (!g853) & (!g907) & (!g909) & (!g914)) + ((!g4) & (g2) & (!g853) & (!g907) & (g909) & (g914)) + ((!g4) & (g2) & (!g853) & (g907) & (g909) & (!g914)) + ((!g4) & (g2) & (!g853) & (g907) & (g909) & (g914)) + ((!g4) & (g2) & (g853) & (!g907) & (g909) & (!g914)) + ((!g4) & (g2) & (g853) & (!g907) & (g909) & (g914)) + ((!g4) & (g2) & (g853) & (g907) & (g909) & (!g914)) + ((!g4) & (g2) & (g853) & (g907) & (g909) & (g914)) + ((g4) & (!g2) & (!g853) & (!g907) & (g909) & (!g914)) + ((g4) & (!g2) & (!g853) & (!g907) & (g909) & (g914)) + ((g4) & (!g2) & (!g853) & (g907) & (g909) & (!g914)) + ((g4) & (!g2) & (!g853) & (g907) & (g909) & (g914)) + ((g4) & (!g2) & (g853) & (!g907) & (g909) & (!g914)) + ((g4) & (!g2) & (g853) & (!g907) & (g909) & (g914)) + ((g4) & (!g2) & (g853) & (g907) & (!g909) & (!g914)) + ((g4) & (!g2) & (g853) & (g907) & (g909) & (g914)) + ((g4) & (g2) & (!g853) & (!g907) & (g909) & (!g914)) + ((g4) & (g2) & (!g853) & (!g907) & (g909) & (g914)) + ((g4) & (g2) & (!g853) & (g907) & (!g909) & (!g914)) + ((g4) & (g2) & (!g853) & (g907) & (g909) & (g914)) + ((g4) & (g2) & (g853) & (!g907) & (!g909) & (!g914)) + ((g4) & (g2) & (g853) & (!g907) & (g909) & (g914)) + ((g4) & (g2) & (g853) & (g907) & (!g909) & (!g914)) + ((g4) & (g2) & (g853) & (g907) & (g909) & (g914)));
	assign g918 = (((!g8) & (!g18) & (!g855) & (g856) & (g906) & (!g914)) + ((!g8) & (!g18) & (g855) & (!g856) & (!g906) & (!g914)) + ((!g8) & (!g18) & (g855) & (!g856) & (!g906) & (g914)) + ((!g8) & (!g18) & (g855) & (!g856) & (g906) & (!g914)) + ((!g8) & (!g18) & (g855) & (!g856) & (g906) & (g914)) + ((!g8) & (!g18) & (g855) & (g856) & (!g906) & (!g914)) + ((!g8) & (!g18) & (g855) & (g856) & (!g906) & (g914)) + ((!g8) & (!g18) & (g855) & (g856) & (g906) & (g914)) + ((!g8) & (g18) & (!g855) & (!g856) & (g906) & (!g914)) + ((!g8) & (g18) & (!g855) & (g856) & (!g906) & (!g914)) + ((!g8) & (g18) & (!g855) & (g856) & (g906) & (!g914)) + ((!g8) & (g18) & (g855) & (!g856) & (!g906) & (!g914)) + ((!g8) & (g18) & (g855) & (!g856) & (!g906) & (g914)) + ((!g8) & (g18) & (g855) & (!g856) & (g906) & (g914)) + ((!g8) & (g18) & (g855) & (g856) & (!g906) & (g914)) + ((!g8) & (g18) & (g855) & (g856) & (g906) & (g914)) + ((g8) & (!g18) & (!g855) & (!g856) & (!g906) & (!g914)) + ((g8) & (!g18) & (!g855) & (!g856) & (g906) & (!g914)) + ((g8) & (!g18) & (!g855) & (g856) & (!g906) & (!g914)) + ((g8) & (!g18) & (g855) & (!g856) & (!g906) & (g914)) + ((g8) & (!g18) & (g855) & (!g856) & (g906) & (g914)) + ((g8) & (!g18) & (g855) & (g856) & (!g906) & (g914)) + ((g8) & (!g18) & (g855) & (g856) & (g906) & (!g914)) + ((g8) & (!g18) & (g855) & (g856) & (g906) & (g914)) + ((g8) & (g18) & (!g855) & (!g856) & (!g906) & (!g914)) + ((g8) & (g18) & (g855) & (!g856) & (!g906) & (g914)) + ((g8) & (g18) & (g855) & (!g856) & (g906) & (!g914)) + ((g8) & (g18) & (g855) & (!g856) & (g906) & (g914)) + ((g8) & (g18) & (g855) & (g856) & (!g906) & (!g914)) + ((g8) & (g18) & (g855) & (g856) & (!g906) & (g914)) + ((g8) & (g18) & (g855) & (g856) & (g906) & (!g914)) + ((g8) & (g18) & (g855) & (g856) & (g906) & (g914)));
	assign g919 = (((!g18) & (!g856) & (g906) & (!g914)) + ((!g18) & (g856) & (!g906) & (!g914)) + ((!g18) & (g856) & (!g906) & (g914)) + ((!g18) & (g856) & (g906) & (g914)) + ((g18) & (!g856) & (!g906) & (!g914)) + ((g18) & (g856) & (!g906) & (g914)) + ((g18) & (g856) & (g906) & (!g914)) + ((g18) & (g856) & (g906) & (g914)));
	assign g920 = (((!g27) & (!g39) & (!g858) & (g859) & (g905) & (!g914)) + ((!g27) & (!g39) & (g858) & (!g859) & (!g905) & (!g914)) + ((!g27) & (!g39) & (g858) & (!g859) & (!g905) & (g914)) + ((!g27) & (!g39) & (g858) & (!g859) & (g905) & (!g914)) + ((!g27) & (!g39) & (g858) & (!g859) & (g905) & (g914)) + ((!g27) & (!g39) & (g858) & (g859) & (!g905) & (!g914)) + ((!g27) & (!g39) & (g858) & (g859) & (!g905) & (g914)) + ((!g27) & (!g39) & (g858) & (g859) & (g905) & (g914)) + ((!g27) & (g39) & (!g858) & (!g859) & (g905) & (!g914)) + ((!g27) & (g39) & (!g858) & (g859) & (!g905) & (!g914)) + ((!g27) & (g39) & (!g858) & (g859) & (g905) & (!g914)) + ((!g27) & (g39) & (g858) & (!g859) & (!g905) & (!g914)) + ((!g27) & (g39) & (g858) & (!g859) & (!g905) & (g914)) + ((!g27) & (g39) & (g858) & (!g859) & (g905) & (g914)) + ((!g27) & (g39) & (g858) & (g859) & (!g905) & (g914)) + ((!g27) & (g39) & (g858) & (g859) & (g905) & (g914)) + ((g27) & (!g39) & (!g858) & (!g859) & (!g905) & (!g914)) + ((g27) & (!g39) & (!g858) & (!g859) & (g905) & (!g914)) + ((g27) & (!g39) & (!g858) & (g859) & (!g905) & (!g914)) + ((g27) & (!g39) & (g858) & (!g859) & (!g905) & (g914)) + ((g27) & (!g39) & (g858) & (!g859) & (g905) & (g914)) + ((g27) & (!g39) & (g858) & (g859) & (!g905) & (g914)) + ((g27) & (!g39) & (g858) & (g859) & (g905) & (!g914)) + ((g27) & (!g39) & (g858) & (g859) & (g905) & (g914)) + ((g27) & (g39) & (!g858) & (!g859) & (!g905) & (!g914)) + ((g27) & (g39) & (g858) & (!g859) & (!g905) & (g914)) + ((g27) & (g39) & (g858) & (!g859) & (g905) & (!g914)) + ((g27) & (g39) & (g858) & (!g859) & (g905) & (g914)) + ((g27) & (g39) & (g858) & (g859) & (!g905) & (!g914)) + ((g27) & (g39) & (g858) & (g859) & (!g905) & (g914)) + ((g27) & (g39) & (g858) & (g859) & (g905) & (!g914)) + ((g27) & (g39) & (g858) & (g859) & (g905) & (g914)));
	assign g921 = (((!g39) & (!g859) & (g905) & (!g914)) + ((!g39) & (g859) & (!g905) & (!g914)) + ((!g39) & (g859) & (!g905) & (g914)) + ((!g39) & (g859) & (g905) & (g914)) + ((g39) & (!g859) & (!g905) & (!g914)) + ((g39) & (g859) & (!g905) & (g914)) + ((g39) & (g859) & (g905) & (!g914)) + ((g39) & (g859) & (g905) & (g914)));
	assign g922 = (((!g54) & (!g68) & (!g861) & (g862) & (g904) & (!g914)) + ((!g54) & (!g68) & (g861) & (!g862) & (!g904) & (!g914)) + ((!g54) & (!g68) & (g861) & (!g862) & (!g904) & (g914)) + ((!g54) & (!g68) & (g861) & (!g862) & (g904) & (!g914)) + ((!g54) & (!g68) & (g861) & (!g862) & (g904) & (g914)) + ((!g54) & (!g68) & (g861) & (g862) & (!g904) & (!g914)) + ((!g54) & (!g68) & (g861) & (g862) & (!g904) & (g914)) + ((!g54) & (!g68) & (g861) & (g862) & (g904) & (g914)) + ((!g54) & (g68) & (!g861) & (!g862) & (g904) & (!g914)) + ((!g54) & (g68) & (!g861) & (g862) & (!g904) & (!g914)) + ((!g54) & (g68) & (!g861) & (g862) & (g904) & (!g914)) + ((!g54) & (g68) & (g861) & (!g862) & (!g904) & (!g914)) + ((!g54) & (g68) & (g861) & (!g862) & (!g904) & (g914)) + ((!g54) & (g68) & (g861) & (!g862) & (g904) & (g914)) + ((!g54) & (g68) & (g861) & (g862) & (!g904) & (g914)) + ((!g54) & (g68) & (g861) & (g862) & (g904) & (g914)) + ((g54) & (!g68) & (!g861) & (!g862) & (!g904) & (!g914)) + ((g54) & (!g68) & (!g861) & (!g862) & (g904) & (!g914)) + ((g54) & (!g68) & (!g861) & (g862) & (!g904) & (!g914)) + ((g54) & (!g68) & (g861) & (!g862) & (!g904) & (g914)) + ((g54) & (!g68) & (g861) & (!g862) & (g904) & (g914)) + ((g54) & (!g68) & (g861) & (g862) & (!g904) & (g914)) + ((g54) & (!g68) & (g861) & (g862) & (g904) & (!g914)) + ((g54) & (!g68) & (g861) & (g862) & (g904) & (g914)) + ((g54) & (g68) & (!g861) & (!g862) & (!g904) & (!g914)) + ((g54) & (g68) & (g861) & (!g862) & (!g904) & (g914)) + ((g54) & (g68) & (g861) & (!g862) & (g904) & (!g914)) + ((g54) & (g68) & (g861) & (!g862) & (g904) & (g914)) + ((g54) & (g68) & (g861) & (g862) & (!g904) & (!g914)) + ((g54) & (g68) & (g861) & (g862) & (!g904) & (g914)) + ((g54) & (g68) & (g861) & (g862) & (g904) & (!g914)) + ((g54) & (g68) & (g861) & (g862) & (g904) & (g914)));
	assign g923 = (((!g68) & (!g862) & (g904) & (!g914)) + ((!g68) & (g862) & (!g904) & (!g914)) + ((!g68) & (g862) & (!g904) & (g914)) + ((!g68) & (g862) & (g904) & (g914)) + ((g68) & (!g862) & (!g904) & (!g914)) + ((g68) & (g862) & (!g904) & (g914)) + ((g68) & (g862) & (g904) & (!g914)) + ((g68) & (g862) & (g904) & (g914)));
	assign g924 = (((!g87) & (!g104) & (!g864) & (g865) & (g903) & (!g914)) + ((!g87) & (!g104) & (g864) & (!g865) & (!g903) & (!g914)) + ((!g87) & (!g104) & (g864) & (!g865) & (!g903) & (g914)) + ((!g87) & (!g104) & (g864) & (!g865) & (g903) & (!g914)) + ((!g87) & (!g104) & (g864) & (!g865) & (g903) & (g914)) + ((!g87) & (!g104) & (g864) & (g865) & (!g903) & (!g914)) + ((!g87) & (!g104) & (g864) & (g865) & (!g903) & (g914)) + ((!g87) & (!g104) & (g864) & (g865) & (g903) & (g914)) + ((!g87) & (g104) & (!g864) & (!g865) & (g903) & (!g914)) + ((!g87) & (g104) & (!g864) & (g865) & (!g903) & (!g914)) + ((!g87) & (g104) & (!g864) & (g865) & (g903) & (!g914)) + ((!g87) & (g104) & (g864) & (!g865) & (!g903) & (!g914)) + ((!g87) & (g104) & (g864) & (!g865) & (!g903) & (g914)) + ((!g87) & (g104) & (g864) & (!g865) & (g903) & (g914)) + ((!g87) & (g104) & (g864) & (g865) & (!g903) & (g914)) + ((!g87) & (g104) & (g864) & (g865) & (g903) & (g914)) + ((g87) & (!g104) & (!g864) & (!g865) & (!g903) & (!g914)) + ((g87) & (!g104) & (!g864) & (!g865) & (g903) & (!g914)) + ((g87) & (!g104) & (!g864) & (g865) & (!g903) & (!g914)) + ((g87) & (!g104) & (g864) & (!g865) & (!g903) & (g914)) + ((g87) & (!g104) & (g864) & (!g865) & (g903) & (g914)) + ((g87) & (!g104) & (g864) & (g865) & (!g903) & (g914)) + ((g87) & (!g104) & (g864) & (g865) & (g903) & (!g914)) + ((g87) & (!g104) & (g864) & (g865) & (g903) & (g914)) + ((g87) & (g104) & (!g864) & (!g865) & (!g903) & (!g914)) + ((g87) & (g104) & (g864) & (!g865) & (!g903) & (g914)) + ((g87) & (g104) & (g864) & (!g865) & (g903) & (!g914)) + ((g87) & (g104) & (g864) & (!g865) & (g903) & (g914)) + ((g87) & (g104) & (g864) & (g865) & (!g903) & (!g914)) + ((g87) & (g104) & (g864) & (g865) & (!g903) & (g914)) + ((g87) & (g104) & (g864) & (g865) & (g903) & (!g914)) + ((g87) & (g104) & (g864) & (g865) & (g903) & (g914)));
	assign g925 = (((!g104) & (!g865) & (g903) & (!g914)) + ((!g104) & (g865) & (!g903) & (!g914)) + ((!g104) & (g865) & (!g903) & (g914)) + ((!g104) & (g865) & (g903) & (g914)) + ((g104) & (!g865) & (!g903) & (!g914)) + ((g104) & (g865) & (!g903) & (g914)) + ((g104) & (g865) & (g903) & (!g914)) + ((g104) & (g865) & (g903) & (g914)));
	assign g926 = (((!g127) & (!g147) & (!g867) & (g868) & (g902) & (!g914)) + ((!g127) & (!g147) & (g867) & (!g868) & (!g902) & (!g914)) + ((!g127) & (!g147) & (g867) & (!g868) & (!g902) & (g914)) + ((!g127) & (!g147) & (g867) & (!g868) & (g902) & (!g914)) + ((!g127) & (!g147) & (g867) & (!g868) & (g902) & (g914)) + ((!g127) & (!g147) & (g867) & (g868) & (!g902) & (!g914)) + ((!g127) & (!g147) & (g867) & (g868) & (!g902) & (g914)) + ((!g127) & (!g147) & (g867) & (g868) & (g902) & (g914)) + ((!g127) & (g147) & (!g867) & (!g868) & (g902) & (!g914)) + ((!g127) & (g147) & (!g867) & (g868) & (!g902) & (!g914)) + ((!g127) & (g147) & (!g867) & (g868) & (g902) & (!g914)) + ((!g127) & (g147) & (g867) & (!g868) & (!g902) & (!g914)) + ((!g127) & (g147) & (g867) & (!g868) & (!g902) & (g914)) + ((!g127) & (g147) & (g867) & (!g868) & (g902) & (g914)) + ((!g127) & (g147) & (g867) & (g868) & (!g902) & (g914)) + ((!g127) & (g147) & (g867) & (g868) & (g902) & (g914)) + ((g127) & (!g147) & (!g867) & (!g868) & (!g902) & (!g914)) + ((g127) & (!g147) & (!g867) & (!g868) & (g902) & (!g914)) + ((g127) & (!g147) & (!g867) & (g868) & (!g902) & (!g914)) + ((g127) & (!g147) & (g867) & (!g868) & (!g902) & (g914)) + ((g127) & (!g147) & (g867) & (!g868) & (g902) & (g914)) + ((g127) & (!g147) & (g867) & (g868) & (!g902) & (g914)) + ((g127) & (!g147) & (g867) & (g868) & (g902) & (!g914)) + ((g127) & (!g147) & (g867) & (g868) & (g902) & (g914)) + ((g127) & (g147) & (!g867) & (!g868) & (!g902) & (!g914)) + ((g127) & (g147) & (g867) & (!g868) & (!g902) & (g914)) + ((g127) & (g147) & (g867) & (!g868) & (g902) & (!g914)) + ((g127) & (g147) & (g867) & (!g868) & (g902) & (g914)) + ((g127) & (g147) & (g867) & (g868) & (!g902) & (!g914)) + ((g127) & (g147) & (g867) & (g868) & (!g902) & (g914)) + ((g127) & (g147) & (g867) & (g868) & (g902) & (!g914)) + ((g127) & (g147) & (g867) & (g868) & (g902) & (g914)));
	assign g927 = (((!g147) & (!g868) & (g902) & (!g914)) + ((!g147) & (g868) & (!g902) & (!g914)) + ((!g147) & (g868) & (!g902) & (g914)) + ((!g147) & (g868) & (g902) & (g914)) + ((g147) & (!g868) & (!g902) & (!g914)) + ((g147) & (g868) & (!g902) & (g914)) + ((g147) & (g868) & (g902) & (!g914)) + ((g147) & (g868) & (g902) & (g914)));
	assign g928 = (((!g174) & (!g198) & (!g870) & (g871) & (g901) & (!g914)) + ((!g174) & (!g198) & (g870) & (!g871) & (!g901) & (!g914)) + ((!g174) & (!g198) & (g870) & (!g871) & (!g901) & (g914)) + ((!g174) & (!g198) & (g870) & (!g871) & (g901) & (!g914)) + ((!g174) & (!g198) & (g870) & (!g871) & (g901) & (g914)) + ((!g174) & (!g198) & (g870) & (g871) & (!g901) & (!g914)) + ((!g174) & (!g198) & (g870) & (g871) & (!g901) & (g914)) + ((!g174) & (!g198) & (g870) & (g871) & (g901) & (g914)) + ((!g174) & (g198) & (!g870) & (!g871) & (g901) & (!g914)) + ((!g174) & (g198) & (!g870) & (g871) & (!g901) & (!g914)) + ((!g174) & (g198) & (!g870) & (g871) & (g901) & (!g914)) + ((!g174) & (g198) & (g870) & (!g871) & (!g901) & (!g914)) + ((!g174) & (g198) & (g870) & (!g871) & (!g901) & (g914)) + ((!g174) & (g198) & (g870) & (!g871) & (g901) & (g914)) + ((!g174) & (g198) & (g870) & (g871) & (!g901) & (g914)) + ((!g174) & (g198) & (g870) & (g871) & (g901) & (g914)) + ((g174) & (!g198) & (!g870) & (!g871) & (!g901) & (!g914)) + ((g174) & (!g198) & (!g870) & (!g871) & (g901) & (!g914)) + ((g174) & (!g198) & (!g870) & (g871) & (!g901) & (!g914)) + ((g174) & (!g198) & (g870) & (!g871) & (!g901) & (g914)) + ((g174) & (!g198) & (g870) & (!g871) & (g901) & (g914)) + ((g174) & (!g198) & (g870) & (g871) & (!g901) & (g914)) + ((g174) & (!g198) & (g870) & (g871) & (g901) & (!g914)) + ((g174) & (!g198) & (g870) & (g871) & (g901) & (g914)) + ((g174) & (g198) & (!g870) & (!g871) & (!g901) & (!g914)) + ((g174) & (g198) & (g870) & (!g871) & (!g901) & (g914)) + ((g174) & (g198) & (g870) & (!g871) & (g901) & (!g914)) + ((g174) & (g198) & (g870) & (!g871) & (g901) & (g914)) + ((g174) & (g198) & (g870) & (g871) & (!g901) & (!g914)) + ((g174) & (g198) & (g870) & (g871) & (!g901) & (g914)) + ((g174) & (g198) & (g870) & (g871) & (g901) & (!g914)) + ((g174) & (g198) & (g870) & (g871) & (g901) & (g914)));
	assign g929 = (((!g198) & (!g871) & (g901) & (!g914)) + ((!g198) & (g871) & (!g901) & (!g914)) + ((!g198) & (g871) & (!g901) & (g914)) + ((!g198) & (g871) & (g901) & (g914)) + ((g198) & (!g871) & (!g901) & (!g914)) + ((g198) & (g871) & (!g901) & (g914)) + ((g198) & (g871) & (g901) & (!g914)) + ((g198) & (g871) & (g901) & (g914)));
	assign g930 = (((!g229) & (!g255) & (!g873) & (g874) & (g900) & (!g914)) + ((!g229) & (!g255) & (g873) & (!g874) & (!g900) & (!g914)) + ((!g229) & (!g255) & (g873) & (!g874) & (!g900) & (g914)) + ((!g229) & (!g255) & (g873) & (!g874) & (g900) & (!g914)) + ((!g229) & (!g255) & (g873) & (!g874) & (g900) & (g914)) + ((!g229) & (!g255) & (g873) & (g874) & (!g900) & (!g914)) + ((!g229) & (!g255) & (g873) & (g874) & (!g900) & (g914)) + ((!g229) & (!g255) & (g873) & (g874) & (g900) & (g914)) + ((!g229) & (g255) & (!g873) & (!g874) & (g900) & (!g914)) + ((!g229) & (g255) & (!g873) & (g874) & (!g900) & (!g914)) + ((!g229) & (g255) & (!g873) & (g874) & (g900) & (!g914)) + ((!g229) & (g255) & (g873) & (!g874) & (!g900) & (!g914)) + ((!g229) & (g255) & (g873) & (!g874) & (!g900) & (g914)) + ((!g229) & (g255) & (g873) & (!g874) & (g900) & (g914)) + ((!g229) & (g255) & (g873) & (g874) & (!g900) & (g914)) + ((!g229) & (g255) & (g873) & (g874) & (g900) & (g914)) + ((g229) & (!g255) & (!g873) & (!g874) & (!g900) & (!g914)) + ((g229) & (!g255) & (!g873) & (!g874) & (g900) & (!g914)) + ((g229) & (!g255) & (!g873) & (g874) & (!g900) & (!g914)) + ((g229) & (!g255) & (g873) & (!g874) & (!g900) & (g914)) + ((g229) & (!g255) & (g873) & (!g874) & (g900) & (g914)) + ((g229) & (!g255) & (g873) & (g874) & (!g900) & (g914)) + ((g229) & (!g255) & (g873) & (g874) & (g900) & (!g914)) + ((g229) & (!g255) & (g873) & (g874) & (g900) & (g914)) + ((g229) & (g255) & (!g873) & (!g874) & (!g900) & (!g914)) + ((g229) & (g255) & (g873) & (!g874) & (!g900) & (g914)) + ((g229) & (g255) & (g873) & (!g874) & (g900) & (!g914)) + ((g229) & (g255) & (g873) & (!g874) & (g900) & (g914)) + ((g229) & (g255) & (g873) & (g874) & (!g900) & (!g914)) + ((g229) & (g255) & (g873) & (g874) & (!g900) & (g914)) + ((g229) & (g255) & (g873) & (g874) & (g900) & (!g914)) + ((g229) & (g255) & (g873) & (g874) & (g900) & (g914)));
	assign g931 = (((!g255) & (!g874) & (g900) & (!g914)) + ((!g255) & (g874) & (!g900) & (!g914)) + ((!g255) & (g874) & (!g900) & (g914)) + ((!g255) & (g874) & (g900) & (g914)) + ((g255) & (!g874) & (!g900) & (!g914)) + ((g255) & (g874) & (!g900) & (g914)) + ((g255) & (g874) & (g900) & (!g914)) + ((g255) & (g874) & (g900) & (g914)));
	assign g932 = (((!g290) & (!g319) & (!g876) & (g877) & (g899) & (!g914)) + ((!g290) & (!g319) & (g876) & (!g877) & (!g899) & (!g914)) + ((!g290) & (!g319) & (g876) & (!g877) & (!g899) & (g914)) + ((!g290) & (!g319) & (g876) & (!g877) & (g899) & (!g914)) + ((!g290) & (!g319) & (g876) & (!g877) & (g899) & (g914)) + ((!g290) & (!g319) & (g876) & (g877) & (!g899) & (!g914)) + ((!g290) & (!g319) & (g876) & (g877) & (!g899) & (g914)) + ((!g290) & (!g319) & (g876) & (g877) & (g899) & (g914)) + ((!g290) & (g319) & (!g876) & (!g877) & (g899) & (!g914)) + ((!g290) & (g319) & (!g876) & (g877) & (!g899) & (!g914)) + ((!g290) & (g319) & (!g876) & (g877) & (g899) & (!g914)) + ((!g290) & (g319) & (g876) & (!g877) & (!g899) & (!g914)) + ((!g290) & (g319) & (g876) & (!g877) & (!g899) & (g914)) + ((!g290) & (g319) & (g876) & (!g877) & (g899) & (g914)) + ((!g290) & (g319) & (g876) & (g877) & (!g899) & (g914)) + ((!g290) & (g319) & (g876) & (g877) & (g899) & (g914)) + ((g290) & (!g319) & (!g876) & (!g877) & (!g899) & (!g914)) + ((g290) & (!g319) & (!g876) & (!g877) & (g899) & (!g914)) + ((g290) & (!g319) & (!g876) & (g877) & (!g899) & (!g914)) + ((g290) & (!g319) & (g876) & (!g877) & (!g899) & (g914)) + ((g290) & (!g319) & (g876) & (!g877) & (g899) & (g914)) + ((g290) & (!g319) & (g876) & (g877) & (!g899) & (g914)) + ((g290) & (!g319) & (g876) & (g877) & (g899) & (!g914)) + ((g290) & (!g319) & (g876) & (g877) & (g899) & (g914)) + ((g290) & (g319) & (!g876) & (!g877) & (!g899) & (!g914)) + ((g290) & (g319) & (g876) & (!g877) & (!g899) & (g914)) + ((g290) & (g319) & (g876) & (!g877) & (g899) & (!g914)) + ((g290) & (g319) & (g876) & (!g877) & (g899) & (g914)) + ((g290) & (g319) & (g876) & (g877) & (!g899) & (!g914)) + ((g290) & (g319) & (g876) & (g877) & (!g899) & (g914)) + ((g290) & (g319) & (g876) & (g877) & (g899) & (!g914)) + ((g290) & (g319) & (g876) & (g877) & (g899) & (g914)));
	assign g933 = (((!g319) & (!g877) & (g899) & (!g914)) + ((!g319) & (g877) & (!g899) & (!g914)) + ((!g319) & (g877) & (!g899) & (g914)) + ((!g319) & (g877) & (g899) & (g914)) + ((g319) & (!g877) & (!g899) & (!g914)) + ((g319) & (g877) & (!g899) & (g914)) + ((g319) & (g877) & (g899) & (!g914)) + ((g319) & (g877) & (g899) & (g914)));
	assign g934 = (((!g358) & (!g390) & (!g879) & (g880) & (g898) & (!g914)) + ((!g358) & (!g390) & (g879) & (!g880) & (!g898) & (!g914)) + ((!g358) & (!g390) & (g879) & (!g880) & (!g898) & (g914)) + ((!g358) & (!g390) & (g879) & (!g880) & (g898) & (!g914)) + ((!g358) & (!g390) & (g879) & (!g880) & (g898) & (g914)) + ((!g358) & (!g390) & (g879) & (g880) & (!g898) & (!g914)) + ((!g358) & (!g390) & (g879) & (g880) & (!g898) & (g914)) + ((!g358) & (!g390) & (g879) & (g880) & (g898) & (g914)) + ((!g358) & (g390) & (!g879) & (!g880) & (g898) & (!g914)) + ((!g358) & (g390) & (!g879) & (g880) & (!g898) & (!g914)) + ((!g358) & (g390) & (!g879) & (g880) & (g898) & (!g914)) + ((!g358) & (g390) & (g879) & (!g880) & (!g898) & (!g914)) + ((!g358) & (g390) & (g879) & (!g880) & (!g898) & (g914)) + ((!g358) & (g390) & (g879) & (!g880) & (g898) & (g914)) + ((!g358) & (g390) & (g879) & (g880) & (!g898) & (g914)) + ((!g358) & (g390) & (g879) & (g880) & (g898) & (g914)) + ((g358) & (!g390) & (!g879) & (!g880) & (!g898) & (!g914)) + ((g358) & (!g390) & (!g879) & (!g880) & (g898) & (!g914)) + ((g358) & (!g390) & (!g879) & (g880) & (!g898) & (!g914)) + ((g358) & (!g390) & (g879) & (!g880) & (!g898) & (g914)) + ((g358) & (!g390) & (g879) & (!g880) & (g898) & (g914)) + ((g358) & (!g390) & (g879) & (g880) & (!g898) & (g914)) + ((g358) & (!g390) & (g879) & (g880) & (g898) & (!g914)) + ((g358) & (!g390) & (g879) & (g880) & (g898) & (g914)) + ((g358) & (g390) & (!g879) & (!g880) & (!g898) & (!g914)) + ((g358) & (g390) & (g879) & (!g880) & (!g898) & (g914)) + ((g358) & (g390) & (g879) & (!g880) & (g898) & (!g914)) + ((g358) & (g390) & (g879) & (!g880) & (g898) & (g914)) + ((g358) & (g390) & (g879) & (g880) & (!g898) & (!g914)) + ((g358) & (g390) & (g879) & (g880) & (!g898) & (g914)) + ((g358) & (g390) & (g879) & (g880) & (g898) & (!g914)) + ((g358) & (g390) & (g879) & (g880) & (g898) & (g914)));
	assign g935 = (((!g390) & (!g880) & (g898) & (!g914)) + ((!g390) & (g880) & (!g898) & (!g914)) + ((!g390) & (g880) & (!g898) & (g914)) + ((!g390) & (g880) & (g898) & (g914)) + ((g390) & (!g880) & (!g898) & (!g914)) + ((g390) & (g880) & (!g898) & (g914)) + ((g390) & (g880) & (g898) & (!g914)) + ((g390) & (g880) & (g898) & (g914)));
	assign g936 = (((!g433) & (!g468) & (!g882) & (g883) & (g897) & (!g914)) + ((!g433) & (!g468) & (g882) & (!g883) & (!g897) & (!g914)) + ((!g433) & (!g468) & (g882) & (!g883) & (!g897) & (g914)) + ((!g433) & (!g468) & (g882) & (!g883) & (g897) & (!g914)) + ((!g433) & (!g468) & (g882) & (!g883) & (g897) & (g914)) + ((!g433) & (!g468) & (g882) & (g883) & (!g897) & (!g914)) + ((!g433) & (!g468) & (g882) & (g883) & (!g897) & (g914)) + ((!g433) & (!g468) & (g882) & (g883) & (g897) & (g914)) + ((!g433) & (g468) & (!g882) & (!g883) & (g897) & (!g914)) + ((!g433) & (g468) & (!g882) & (g883) & (!g897) & (!g914)) + ((!g433) & (g468) & (!g882) & (g883) & (g897) & (!g914)) + ((!g433) & (g468) & (g882) & (!g883) & (!g897) & (!g914)) + ((!g433) & (g468) & (g882) & (!g883) & (!g897) & (g914)) + ((!g433) & (g468) & (g882) & (!g883) & (g897) & (g914)) + ((!g433) & (g468) & (g882) & (g883) & (!g897) & (g914)) + ((!g433) & (g468) & (g882) & (g883) & (g897) & (g914)) + ((g433) & (!g468) & (!g882) & (!g883) & (!g897) & (!g914)) + ((g433) & (!g468) & (!g882) & (!g883) & (g897) & (!g914)) + ((g433) & (!g468) & (!g882) & (g883) & (!g897) & (!g914)) + ((g433) & (!g468) & (g882) & (!g883) & (!g897) & (g914)) + ((g433) & (!g468) & (g882) & (!g883) & (g897) & (g914)) + ((g433) & (!g468) & (g882) & (g883) & (!g897) & (g914)) + ((g433) & (!g468) & (g882) & (g883) & (g897) & (!g914)) + ((g433) & (!g468) & (g882) & (g883) & (g897) & (g914)) + ((g433) & (g468) & (!g882) & (!g883) & (!g897) & (!g914)) + ((g433) & (g468) & (g882) & (!g883) & (!g897) & (g914)) + ((g433) & (g468) & (g882) & (!g883) & (g897) & (!g914)) + ((g433) & (g468) & (g882) & (!g883) & (g897) & (g914)) + ((g433) & (g468) & (g882) & (g883) & (!g897) & (!g914)) + ((g433) & (g468) & (g882) & (g883) & (!g897) & (g914)) + ((g433) & (g468) & (g882) & (g883) & (g897) & (!g914)) + ((g433) & (g468) & (g882) & (g883) & (g897) & (g914)));
	assign g937 = (((!g468) & (!g883) & (g897) & (!g914)) + ((!g468) & (g883) & (!g897) & (!g914)) + ((!g468) & (g883) & (!g897) & (g914)) + ((!g468) & (g883) & (g897) & (g914)) + ((g468) & (!g883) & (!g897) & (!g914)) + ((g468) & (g883) & (!g897) & (g914)) + ((g468) & (g883) & (g897) & (!g914)) + ((g468) & (g883) & (g897) & (g914)));
	assign g938 = (((!g515) & (!g553) & (!g885) & (g886) & (g896) & (!g914)) + ((!g515) & (!g553) & (g885) & (!g886) & (!g896) & (!g914)) + ((!g515) & (!g553) & (g885) & (!g886) & (!g896) & (g914)) + ((!g515) & (!g553) & (g885) & (!g886) & (g896) & (!g914)) + ((!g515) & (!g553) & (g885) & (!g886) & (g896) & (g914)) + ((!g515) & (!g553) & (g885) & (g886) & (!g896) & (!g914)) + ((!g515) & (!g553) & (g885) & (g886) & (!g896) & (g914)) + ((!g515) & (!g553) & (g885) & (g886) & (g896) & (g914)) + ((!g515) & (g553) & (!g885) & (!g886) & (g896) & (!g914)) + ((!g515) & (g553) & (!g885) & (g886) & (!g896) & (!g914)) + ((!g515) & (g553) & (!g885) & (g886) & (g896) & (!g914)) + ((!g515) & (g553) & (g885) & (!g886) & (!g896) & (!g914)) + ((!g515) & (g553) & (g885) & (!g886) & (!g896) & (g914)) + ((!g515) & (g553) & (g885) & (!g886) & (g896) & (g914)) + ((!g515) & (g553) & (g885) & (g886) & (!g896) & (g914)) + ((!g515) & (g553) & (g885) & (g886) & (g896) & (g914)) + ((g515) & (!g553) & (!g885) & (!g886) & (!g896) & (!g914)) + ((g515) & (!g553) & (!g885) & (!g886) & (g896) & (!g914)) + ((g515) & (!g553) & (!g885) & (g886) & (!g896) & (!g914)) + ((g515) & (!g553) & (g885) & (!g886) & (!g896) & (g914)) + ((g515) & (!g553) & (g885) & (!g886) & (g896) & (g914)) + ((g515) & (!g553) & (g885) & (g886) & (!g896) & (g914)) + ((g515) & (!g553) & (g885) & (g886) & (g896) & (!g914)) + ((g515) & (!g553) & (g885) & (g886) & (g896) & (g914)) + ((g515) & (g553) & (!g885) & (!g886) & (!g896) & (!g914)) + ((g515) & (g553) & (g885) & (!g886) & (!g896) & (g914)) + ((g515) & (g553) & (g885) & (!g886) & (g896) & (!g914)) + ((g515) & (g553) & (g885) & (!g886) & (g896) & (g914)) + ((g515) & (g553) & (g885) & (g886) & (!g896) & (!g914)) + ((g515) & (g553) & (g885) & (g886) & (!g896) & (g914)) + ((g515) & (g553) & (g885) & (g886) & (g896) & (!g914)) + ((g515) & (g553) & (g885) & (g886) & (g896) & (g914)));
	assign g939 = (((!g553) & (!g886) & (g896) & (!g914)) + ((!g553) & (g886) & (!g896) & (!g914)) + ((!g553) & (g886) & (!g896) & (g914)) + ((!g553) & (g886) & (g896) & (g914)) + ((g553) & (!g886) & (!g896) & (!g914)) + ((g553) & (g886) & (!g896) & (g914)) + ((g553) & (g886) & (g896) & (!g914)) + ((g553) & (g886) & (g896) & (g914)));
	assign g940 = (((!g604) & (!g645) & (!g888) & (g889) & (g895) & (!g914)) + ((!g604) & (!g645) & (g888) & (!g889) & (!g895) & (!g914)) + ((!g604) & (!g645) & (g888) & (!g889) & (!g895) & (g914)) + ((!g604) & (!g645) & (g888) & (!g889) & (g895) & (!g914)) + ((!g604) & (!g645) & (g888) & (!g889) & (g895) & (g914)) + ((!g604) & (!g645) & (g888) & (g889) & (!g895) & (!g914)) + ((!g604) & (!g645) & (g888) & (g889) & (!g895) & (g914)) + ((!g604) & (!g645) & (g888) & (g889) & (g895) & (g914)) + ((!g604) & (g645) & (!g888) & (!g889) & (g895) & (!g914)) + ((!g604) & (g645) & (!g888) & (g889) & (!g895) & (!g914)) + ((!g604) & (g645) & (!g888) & (g889) & (g895) & (!g914)) + ((!g604) & (g645) & (g888) & (!g889) & (!g895) & (!g914)) + ((!g604) & (g645) & (g888) & (!g889) & (!g895) & (g914)) + ((!g604) & (g645) & (g888) & (!g889) & (g895) & (g914)) + ((!g604) & (g645) & (g888) & (g889) & (!g895) & (g914)) + ((!g604) & (g645) & (g888) & (g889) & (g895) & (g914)) + ((g604) & (!g645) & (!g888) & (!g889) & (!g895) & (!g914)) + ((g604) & (!g645) & (!g888) & (!g889) & (g895) & (!g914)) + ((g604) & (!g645) & (!g888) & (g889) & (!g895) & (!g914)) + ((g604) & (!g645) & (g888) & (!g889) & (!g895) & (g914)) + ((g604) & (!g645) & (g888) & (!g889) & (g895) & (g914)) + ((g604) & (!g645) & (g888) & (g889) & (!g895) & (g914)) + ((g604) & (!g645) & (g888) & (g889) & (g895) & (!g914)) + ((g604) & (!g645) & (g888) & (g889) & (g895) & (g914)) + ((g604) & (g645) & (!g888) & (!g889) & (!g895) & (!g914)) + ((g604) & (g645) & (g888) & (!g889) & (!g895) & (g914)) + ((g604) & (g645) & (g888) & (!g889) & (g895) & (!g914)) + ((g604) & (g645) & (g888) & (!g889) & (g895) & (g914)) + ((g604) & (g645) & (g888) & (g889) & (!g895) & (!g914)) + ((g604) & (g645) & (g888) & (g889) & (!g895) & (g914)) + ((g604) & (g645) & (g888) & (g889) & (g895) & (!g914)) + ((g604) & (g645) & (g888) & (g889) & (g895) & (g914)));
	assign g941 = (((!g645) & (!g889) & (g895) & (!g914)) + ((!g645) & (g889) & (!g895) & (!g914)) + ((!g645) & (g889) & (!g895) & (g914)) + ((!g645) & (g889) & (g895) & (g914)) + ((g645) & (!g889) & (!g895) & (!g914)) + ((g645) & (g889) & (!g895) & (g914)) + ((g645) & (g889) & (g895) & (!g914)) + ((g645) & (g889) & (g895) & (g914)));
	assign g942 = (((!g700) & (!g744) & (!g891) & (g892) & (g894) & (!g914)) + ((!g700) & (!g744) & (g891) & (!g892) & (!g894) & (!g914)) + ((!g700) & (!g744) & (g891) & (!g892) & (!g894) & (g914)) + ((!g700) & (!g744) & (g891) & (!g892) & (g894) & (!g914)) + ((!g700) & (!g744) & (g891) & (!g892) & (g894) & (g914)) + ((!g700) & (!g744) & (g891) & (g892) & (!g894) & (!g914)) + ((!g700) & (!g744) & (g891) & (g892) & (!g894) & (g914)) + ((!g700) & (!g744) & (g891) & (g892) & (g894) & (g914)) + ((!g700) & (g744) & (!g891) & (!g892) & (g894) & (!g914)) + ((!g700) & (g744) & (!g891) & (g892) & (!g894) & (!g914)) + ((!g700) & (g744) & (!g891) & (g892) & (g894) & (!g914)) + ((!g700) & (g744) & (g891) & (!g892) & (!g894) & (!g914)) + ((!g700) & (g744) & (g891) & (!g892) & (!g894) & (g914)) + ((!g700) & (g744) & (g891) & (!g892) & (g894) & (g914)) + ((!g700) & (g744) & (g891) & (g892) & (!g894) & (g914)) + ((!g700) & (g744) & (g891) & (g892) & (g894) & (g914)) + ((g700) & (!g744) & (!g891) & (!g892) & (!g894) & (!g914)) + ((g700) & (!g744) & (!g891) & (!g892) & (g894) & (!g914)) + ((g700) & (!g744) & (!g891) & (g892) & (!g894) & (!g914)) + ((g700) & (!g744) & (g891) & (!g892) & (!g894) & (g914)) + ((g700) & (!g744) & (g891) & (!g892) & (g894) & (g914)) + ((g700) & (!g744) & (g891) & (g892) & (!g894) & (g914)) + ((g700) & (!g744) & (g891) & (g892) & (g894) & (!g914)) + ((g700) & (!g744) & (g891) & (g892) & (g894) & (g914)) + ((g700) & (g744) & (!g891) & (!g892) & (!g894) & (!g914)) + ((g700) & (g744) & (g891) & (!g892) & (!g894) & (g914)) + ((g700) & (g744) & (g891) & (!g892) & (g894) & (!g914)) + ((g700) & (g744) & (g891) & (!g892) & (g894) & (g914)) + ((g700) & (g744) & (g891) & (g892) & (!g894) & (!g914)) + ((g700) & (g744) & (g891) & (g892) & (!g894) & (g914)) + ((g700) & (g744) & (g891) & (g892) & (g894) & (!g914)) + ((g700) & (g744) & (g891) & (g892) & (g894) & (g914)));
	assign g943 = (((!g744) & (!g892) & (g894) & (!g914)) + ((!g744) & (g892) & (!g894) & (!g914)) + ((!g744) & (g892) & (!g894) & (g914)) + ((!g744) & (g892) & (g894) & (g914)) + ((g744) & (!g892) & (!g894) & (!g914)) + ((g744) & (g892) & (!g894) & (g914)) + ((g744) & (g892) & (g894) & (!g914)) + ((g744) & (g892) & (g894) & (g914)));
	assign g944 = (((!g803) & (!ax66x) & (!ax67x) & (!g851) & (!g893) & (g914)) + ((!g803) & (!ax66x) & (!ax67x) & (!g851) & (g893) & (!g914)) + ((!g803) & (!ax66x) & (!ax67x) & (!g851) & (g893) & (g914)) + ((!g803) & (!ax66x) & (!ax67x) & (g851) & (!g893) & (!g914)) + ((!g803) & (!ax66x) & (ax67x) & (!g851) & (!g893) & (!g914)) + ((!g803) & (!ax66x) & (ax67x) & (g851) & (!g893) & (g914)) + ((!g803) & (!ax66x) & (ax67x) & (g851) & (g893) & (!g914)) + ((!g803) & (!ax66x) & (ax67x) & (g851) & (g893) & (g914)) + ((!g803) & (ax66x) & (!ax67x) & (g851) & (!g893) & (!g914)) + ((!g803) & (ax66x) & (!ax67x) & (g851) & (g893) & (!g914)) + ((!g803) & (ax66x) & (ax67x) & (!g851) & (!g893) & (!g914)) + ((!g803) & (ax66x) & (ax67x) & (!g851) & (!g893) & (g914)) + ((!g803) & (ax66x) & (ax67x) & (!g851) & (g893) & (!g914)) + ((!g803) & (ax66x) & (ax67x) & (!g851) & (g893) & (g914)) + ((!g803) & (ax66x) & (ax67x) & (g851) & (!g893) & (g914)) + ((!g803) & (ax66x) & (ax67x) & (g851) & (g893) & (g914)) + ((g803) & (!ax66x) & (!ax67x) & (!g851) & (!g893) & (!g914)) + ((g803) & (!ax66x) & (!ax67x) & (!g851) & (!g893) & (g914)) + ((g803) & (!ax66x) & (!ax67x) & (!g851) & (g893) & (g914)) + ((g803) & (!ax66x) & (!ax67x) & (g851) & (g893) & (!g914)) + ((g803) & (!ax66x) & (ax67x) & (!g851) & (g893) & (!g914)) + ((g803) & (!ax66x) & (ax67x) & (g851) & (!g893) & (!g914)) + ((g803) & (!ax66x) & (ax67x) & (g851) & (!g893) & (g914)) + ((g803) & (!ax66x) & (ax67x) & (g851) & (g893) & (g914)) + ((g803) & (ax66x) & (!ax67x) & (!g851) & (!g893) & (!g914)) + ((g803) & (ax66x) & (!ax67x) & (!g851) & (g893) & (!g914)) + ((g803) & (ax66x) & (ax67x) & (!g851) & (!g893) & (g914)) + ((g803) & (ax66x) & (ax67x) & (!g851) & (g893) & (g914)) + ((g803) & (ax66x) & (ax67x) & (g851) & (!g893) & (!g914)) + ((g803) & (ax66x) & (ax67x) & (g851) & (!g893) & (g914)) + ((g803) & (ax66x) & (ax67x) & (g851) & (g893) & (!g914)) + ((g803) & (ax66x) & (ax67x) & (g851) & (g893) & (g914)));
	assign g945 = (((!ax66x) & (!g851) & (!g893) & (g914)) + ((!ax66x) & (!g851) & (g893) & (!g914)) + ((!ax66x) & (!g851) & (g893) & (g914)) + ((!ax66x) & (g851) & (g893) & (!g914)) + ((ax66x) & (!g851) & (!g893) & (!g914)) + ((ax66x) & (g851) & (!g893) & (!g914)) + ((ax66x) & (g851) & (!g893) & (g914)) + ((ax66x) & (g851) & (g893) & (g914)));
	assign g946 = (((!ax64x) & (!ax65x) & (!g851) & (!g914) & (!g915)) + ((!ax64x) & (!ax65x) & (g851) & (!g914) & (!g915)) + ((!ax64x) & (!ax65x) & (g851) & (!g914) & (g915)) + ((!ax64x) & (!ax65x) & (g851) & (g914) & (!g915)) + ((!ax64x) & (ax65x) & (!g851) & (g914) & (!g915)) + ((!ax64x) & (ax65x) & (g851) & (!g914) & (!g915)) + ((!ax64x) & (ax65x) & (g851) & (g914) & (!g915)) + ((!ax64x) & (ax65x) & (g851) & (g914) & (g915)) + ((ax64x) & (!ax65x) & (g851) & (g914) & (!g915)) + ((ax64x) & (!ax65x) & (g851) & (g914) & (g915)) + ((ax64x) & (ax65x) & (!g851) & (g914) & (!g915)) + ((ax64x) & (ax65x) & (!g851) & (g914) & (g915)) + ((ax64x) & (ax65x) & (g851) & (!g914) & (!g915)) + ((ax64x) & (ax65x) & (g851) & (!g914) & (g915)) + ((ax64x) & (ax65x) & (g851) & (g914) & (!g915)) + ((ax64x) & (ax65x) & (g851) & (g914) & (g915)));
	assign g947 = (((!g744) & (!g803) & (g944) & (g945) & (g946)) + ((!g744) & (g803) & (g944) & (!g945) & (g946)) + ((!g744) & (g803) & (g944) & (g945) & (!g946)) + ((!g744) & (g803) & (g944) & (g945) & (g946)) + ((g744) & (!g803) & (!g944) & (g945) & (g946)) + ((g744) & (!g803) & (g944) & (!g945) & (!g946)) + ((g744) & (!g803) & (g944) & (!g945) & (g946)) + ((g744) & (!g803) & (g944) & (g945) & (!g946)) + ((g744) & (!g803) & (g944) & (g945) & (g946)) + ((g744) & (g803) & (!g944) & (!g945) & (g946)) + ((g744) & (g803) & (!g944) & (g945) & (!g946)) + ((g744) & (g803) & (!g944) & (g945) & (g946)) + ((g744) & (g803) & (g944) & (!g945) & (!g946)) + ((g744) & (g803) & (g944) & (!g945) & (g946)) + ((g744) & (g803) & (g944) & (g945) & (!g946)) + ((g744) & (g803) & (g944) & (g945) & (g946)));
	assign g948 = (((!g645) & (!g700) & (g942) & (g943) & (g947)) + ((!g645) & (g700) & (g942) & (!g943) & (g947)) + ((!g645) & (g700) & (g942) & (g943) & (!g947)) + ((!g645) & (g700) & (g942) & (g943) & (g947)) + ((g645) & (!g700) & (!g942) & (g943) & (g947)) + ((g645) & (!g700) & (g942) & (!g943) & (!g947)) + ((g645) & (!g700) & (g942) & (!g943) & (g947)) + ((g645) & (!g700) & (g942) & (g943) & (!g947)) + ((g645) & (!g700) & (g942) & (g943) & (g947)) + ((g645) & (g700) & (!g942) & (!g943) & (g947)) + ((g645) & (g700) & (!g942) & (g943) & (!g947)) + ((g645) & (g700) & (!g942) & (g943) & (g947)) + ((g645) & (g700) & (g942) & (!g943) & (!g947)) + ((g645) & (g700) & (g942) & (!g943) & (g947)) + ((g645) & (g700) & (g942) & (g943) & (!g947)) + ((g645) & (g700) & (g942) & (g943) & (g947)));
	assign g949 = (((!g553) & (!g604) & (g940) & (g941) & (g948)) + ((!g553) & (g604) & (g940) & (!g941) & (g948)) + ((!g553) & (g604) & (g940) & (g941) & (!g948)) + ((!g553) & (g604) & (g940) & (g941) & (g948)) + ((g553) & (!g604) & (!g940) & (g941) & (g948)) + ((g553) & (!g604) & (g940) & (!g941) & (!g948)) + ((g553) & (!g604) & (g940) & (!g941) & (g948)) + ((g553) & (!g604) & (g940) & (g941) & (!g948)) + ((g553) & (!g604) & (g940) & (g941) & (g948)) + ((g553) & (g604) & (!g940) & (!g941) & (g948)) + ((g553) & (g604) & (!g940) & (g941) & (!g948)) + ((g553) & (g604) & (!g940) & (g941) & (g948)) + ((g553) & (g604) & (g940) & (!g941) & (!g948)) + ((g553) & (g604) & (g940) & (!g941) & (g948)) + ((g553) & (g604) & (g940) & (g941) & (!g948)) + ((g553) & (g604) & (g940) & (g941) & (g948)));
	assign g950 = (((!g468) & (!g515) & (g938) & (g939) & (g949)) + ((!g468) & (g515) & (g938) & (!g939) & (g949)) + ((!g468) & (g515) & (g938) & (g939) & (!g949)) + ((!g468) & (g515) & (g938) & (g939) & (g949)) + ((g468) & (!g515) & (!g938) & (g939) & (g949)) + ((g468) & (!g515) & (g938) & (!g939) & (!g949)) + ((g468) & (!g515) & (g938) & (!g939) & (g949)) + ((g468) & (!g515) & (g938) & (g939) & (!g949)) + ((g468) & (!g515) & (g938) & (g939) & (g949)) + ((g468) & (g515) & (!g938) & (!g939) & (g949)) + ((g468) & (g515) & (!g938) & (g939) & (!g949)) + ((g468) & (g515) & (!g938) & (g939) & (g949)) + ((g468) & (g515) & (g938) & (!g939) & (!g949)) + ((g468) & (g515) & (g938) & (!g939) & (g949)) + ((g468) & (g515) & (g938) & (g939) & (!g949)) + ((g468) & (g515) & (g938) & (g939) & (g949)));
	assign g951 = (((!g390) & (!g433) & (g936) & (g937) & (g950)) + ((!g390) & (g433) & (g936) & (!g937) & (g950)) + ((!g390) & (g433) & (g936) & (g937) & (!g950)) + ((!g390) & (g433) & (g936) & (g937) & (g950)) + ((g390) & (!g433) & (!g936) & (g937) & (g950)) + ((g390) & (!g433) & (g936) & (!g937) & (!g950)) + ((g390) & (!g433) & (g936) & (!g937) & (g950)) + ((g390) & (!g433) & (g936) & (g937) & (!g950)) + ((g390) & (!g433) & (g936) & (g937) & (g950)) + ((g390) & (g433) & (!g936) & (!g937) & (g950)) + ((g390) & (g433) & (!g936) & (g937) & (!g950)) + ((g390) & (g433) & (!g936) & (g937) & (g950)) + ((g390) & (g433) & (g936) & (!g937) & (!g950)) + ((g390) & (g433) & (g936) & (!g937) & (g950)) + ((g390) & (g433) & (g936) & (g937) & (!g950)) + ((g390) & (g433) & (g936) & (g937) & (g950)));
	assign g952 = (((!g319) & (!g358) & (g934) & (g935) & (g951)) + ((!g319) & (g358) & (g934) & (!g935) & (g951)) + ((!g319) & (g358) & (g934) & (g935) & (!g951)) + ((!g319) & (g358) & (g934) & (g935) & (g951)) + ((g319) & (!g358) & (!g934) & (g935) & (g951)) + ((g319) & (!g358) & (g934) & (!g935) & (!g951)) + ((g319) & (!g358) & (g934) & (!g935) & (g951)) + ((g319) & (!g358) & (g934) & (g935) & (!g951)) + ((g319) & (!g358) & (g934) & (g935) & (g951)) + ((g319) & (g358) & (!g934) & (!g935) & (g951)) + ((g319) & (g358) & (!g934) & (g935) & (!g951)) + ((g319) & (g358) & (!g934) & (g935) & (g951)) + ((g319) & (g358) & (g934) & (!g935) & (!g951)) + ((g319) & (g358) & (g934) & (!g935) & (g951)) + ((g319) & (g358) & (g934) & (g935) & (!g951)) + ((g319) & (g358) & (g934) & (g935) & (g951)));
	assign g953 = (((!g255) & (!g290) & (g932) & (g933) & (g952)) + ((!g255) & (g290) & (g932) & (!g933) & (g952)) + ((!g255) & (g290) & (g932) & (g933) & (!g952)) + ((!g255) & (g290) & (g932) & (g933) & (g952)) + ((g255) & (!g290) & (!g932) & (g933) & (g952)) + ((g255) & (!g290) & (g932) & (!g933) & (!g952)) + ((g255) & (!g290) & (g932) & (!g933) & (g952)) + ((g255) & (!g290) & (g932) & (g933) & (!g952)) + ((g255) & (!g290) & (g932) & (g933) & (g952)) + ((g255) & (g290) & (!g932) & (!g933) & (g952)) + ((g255) & (g290) & (!g932) & (g933) & (!g952)) + ((g255) & (g290) & (!g932) & (g933) & (g952)) + ((g255) & (g290) & (g932) & (!g933) & (!g952)) + ((g255) & (g290) & (g932) & (!g933) & (g952)) + ((g255) & (g290) & (g932) & (g933) & (!g952)) + ((g255) & (g290) & (g932) & (g933) & (g952)));
	assign g954 = (((!g198) & (!g229) & (g930) & (g931) & (g953)) + ((!g198) & (g229) & (g930) & (!g931) & (g953)) + ((!g198) & (g229) & (g930) & (g931) & (!g953)) + ((!g198) & (g229) & (g930) & (g931) & (g953)) + ((g198) & (!g229) & (!g930) & (g931) & (g953)) + ((g198) & (!g229) & (g930) & (!g931) & (!g953)) + ((g198) & (!g229) & (g930) & (!g931) & (g953)) + ((g198) & (!g229) & (g930) & (g931) & (!g953)) + ((g198) & (!g229) & (g930) & (g931) & (g953)) + ((g198) & (g229) & (!g930) & (!g931) & (g953)) + ((g198) & (g229) & (!g930) & (g931) & (!g953)) + ((g198) & (g229) & (!g930) & (g931) & (g953)) + ((g198) & (g229) & (g930) & (!g931) & (!g953)) + ((g198) & (g229) & (g930) & (!g931) & (g953)) + ((g198) & (g229) & (g930) & (g931) & (!g953)) + ((g198) & (g229) & (g930) & (g931) & (g953)));
	assign g955 = (((!g147) & (!g174) & (g928) & (g929) & (g954)) + ((!g147) & (g174) & (g928) & (!g929) & (g954)) + ((!g147) & (g174) & (g928) & (g929) & (!g954)) + ((!g147) & (g174) & (g928) & (g929) & (g954)) + ((g147) & (!g174) & (!g928) & (g929) & (g954)) + ((g147) & (!g174) & (g928) & (!g929) & (!g954)) + ((g147) & (!g174) & (g928) & (!g929) & (g954)) + ((g147) & (!g174) & (g928) & (g929) & (!g954)) + ((g147) & (!g174) & (g928) & (g929) & (g954)) + ((g147) & (g174) & (!g928) & (!g929) & (g954)) + ((g147) & (g174) & (!g928) & (g929) & (!g954)) + ((g147) & (g174) & (!g928) & (g929) & (g954)) + ((g147) & (g174) & (g928) & (!g929) & (!g954)) + ((g147) & (g174) & (g928) & (!g929) & (g954)) + ((g147) & (g174) & (g928) & (g929) & (!g954)) + ((g147) & (g174) & (g928) & (g929) & (g954)));
	assign g956 = (((!g104) & (!g127) & (g926) & (g927) & (g955)) + ((!g104) & (g127) & (g926) & (!g927) & (g955)) + ((!g104) & (g127) & (g926) & (g927) & (!g955)) + ((!g104) & (g127) & (g926) & (g927) & (g955)) + ((g104) & (!g127) & (!g926) & (g927) & (g955)) + ((g104) & (!g127) & (g926) & (!g927) & (!g955)) + ((g104) & (!g127) & (g926) & (!g927) & (g955)) + ((g104) & (!g127) & (g926) & (g927) & (!g955)) + ((g104) & (!g127) & (g926) & (g927) & (g955)) + ((g104) & (g127) & (!g926) & (!g927) & (g955)) + ((g104) & (g127) & (!g926) & (g927) & (!g955)) + ((g104) & (g127) & (!g926) & (g927) & (g955)) + ((g104) & (g127) & (g926) & (!g927) & (!g955)) + ((g104) & (g127) & (g926) & (!g927) & (g955)) + ((g104) & (g127) & (g926) & (g927) & (!g955)) + ((g104) & (g127) & (g926) & (g927) & (g955)));
	assign g957 = (((!g68) & (!g87) & (g924) & (g925) & (g956)) + ((!g68) & (g87) & (g924) & (!g925) & (g956)) + ((!g68) & (g87) & (g924) & (g925) & (!g956)) + ((!g68) & (g87) & (g924) & (g925) & (g956)) + ((g68) & (!g87) & (!g924) & (g925) & (g956)) + ((g68) & (!g87) & (g924) & (!g925) & (!g956)) + ((g68) & (!g87) & (g924) & (!g925) & (g956)) + ((g68) & (!g87) & (g924) & (g925) & (!g956)) + ((g68) & (!g87) & (g924) & (g925) & (g956)) + ((g68) & (g87) & (!g924) & (!g925) & (g956)) + ((g68) & (g87) & (!g924) & (g925) & (!g956)) + ((g68) & (g87) & (!g924) & (g925) & (g956)) + ((g68) & (g87) & (g924) & (!g925) & (!g956)) + ((g68) & (g87) & (g924) & (!g925) & (g956)) + ((g68) & (g87) & (g924) & (g925) & (!g956)) + ((g68) & (g87) & (g924) & (g925) & (g956)));
	assign g958 = (((!g39) & (!g54) & (g922) & (g923) & (g957)) + ((!g39) & (g54) & (g922) & (!g923) & (g957)) + ((!g39) & (g54) & (g922) & (g923) & (!g957)) + ((!g39) & (g54) & (g922) & (g923) & (g957)) + ((g39) & (!g54) & (!g922) & (g923) & (g957)) + ((g39) & (!g54) & (g922) & (!g923) & (!g957)) + ((g39) & (!g54) & (g922) & (!g923) & (g957)) + ((g39) & (!g54) & (g922) & (g923) & (!g957)) + ((g39) & (!g54) & (g922) & (g923) & (g957)) + ((g39) & (g54) & (!g922) & (!g923) & (g957)) + ((g39) & (g54) & (!g922) & (g923) & (!g957)) + ((g39) & (g54) & (!g922) & (g923) & (g957)) + ((g39) & (g54) & (g922) & (!g923) & (!g957)) + ((g39) & (g54) & (g922) & (!g923) & (g957)) + ((g39) & (g54) & (g922) & (g923) & (!g957)) + ((g39) & (g54) & (g922) & (g923) & (g957)));
	assign g959 = (((!g18) & (!g27) & (g920) & (g921) & (g958)) + ((!g18) & (g27) & (g920) & (!g921) & (g958)) + ((!g18) & (g27) & (g920) & (g921) & (!g958)) + ((!g18) & (g27) & (g920) & (g921) & (g958)) + ((g18) & (!g27) & (!g920) & (g921) & (g958)) + ((g18) & (!g27) & (g920) & (!g921) & (!g958)) + ((g18) & (!g27) & (g920) & (!g921) & (g958)) + ((g18) & (!g27) & (g920) & (g921) & (!g958)) + ((g18) & (!g27) & (g920) & (g921) & (g958)) + ((g18) & (g27) & (!g920) & (!g921) & (g958)) + ((g18) & (g27) & (!g920) & (g921) & (!g958)) + ((g18) & (g27) & (!g920) & (g921) & (g958)) + ((g18) & (g27) & (g920) & (!g921) & (!g958)) + ((g18) & (g27) & (g920) & (!g921) & (g958)) + ((g18) & (g27) & (g920) & (g921) & (!g958)) + ((g18) & (g27) & (g920) & (g921) & (g958)));
	assign g960 = (((!g2) & (!g8) & (g918) & (g919) & (g959)) + ((!g2) & (g8) & (g918) & (!g919) & (g959)) + ((!g2) & (g8) & (g918) & (g919) & (!g959)) + ((!g2) & (g8) & (g918) & (g919) & (g959)) + ((g2) & (!g8) & (!g918) & (g919) & (g959)) + ((g2) & (!g8) & (g918) & (!g919) & (!g959)) + ((g2) & (!g8) & (g918) & (!g919) & (g959)) + ((g2) & (!g8) & (g918) & (g919) & (!g959)) + ((g2) & (!g8) & (g918) & (g919) & (g959)) + ((g2) & (g8) & (!g918) & (!g919) & (g959)) + ((g2) & (g8) & (!g918) & (g919) & (!g959)) + ((g2) & (g8) & (!g918) & (g919) & (g959)) + ((g2) & (g8) & (g918) & (!g919) & (!g959)) + ((g2) & (g8) & (g918) & (!g919) & (g959)) + ((g2) & (g8) & (g918) & (g919) & (!g959)) + ((g2) & (g8) & (g918) & (g919) & (g959)));
	assign g961 = (((!g2) & (!g853) & (g907) & (!g914)) + ((!g2) & (g853) & (!g907) & (!g914)) + ((!g2) & (g853) & (!g907) & (g914)) + ((!g2) & (g853) & (g907) & (g914)) + ((g2) & (!g853) & (!g907) & (!g914)) + ((g2) & (g853) & (!g907) & (g914)) + ((g2) & (g853) & (g907) & (!g914)) + ((g2) & (g853) & (g907) & (g914)));
	assign g962 = (((!g1) & (!g852) & (!g910) & (!g912) & (g913)) + ((!g1) & (!g852) & (!g910) & (g912) & (!g913)) + ((!g1) & (!g852) & (!g910) & (g912) & (g913)) + ((!g1) & (g852) & (g910) & (!g912) & (!g913)) + ((!g1) & (g852) & (g910) & (!g912) & (g913)) + ((!g1) & (g852) & (g910) & (g912) & (!g913)) + ((!g1) & (g852) & (g910) & (g912) & (g913)) + ((g1) & (!g852) & (!g910) & (!g912) & (g913)) + ((g1) & (!g852) & (!g910) & (g912) & (g913)) + ((g1) & (g852) & (g910) & (!g912) & (!g913)) + ((g1) & (g852) & (g910) & (!g912) & (g913)) + ((g1) & (g852) & (g910) & (g912) & (!g913)) + ((g1) & (g852) & (g910) & (g912) & (g913)));
	assign g963 = (((!g4) & (!g1) & (!g917) & (!g960) & (!g961) & (!g962)) + ((!g4) & (g1) & (!g917) & (!g960) & (!g961) & (!g962)) + ((!g4) & (g1) & (!g917) & (!g960) & (!g961) & (g962)) + ((!g4) & (g1) & (!g917) & (!g960) & (g961) & (!g962)) + ((!g4) & (g1) & (!g917) & (!g960) & (g961) & (g962)) + ((!g4) & (g1) & (!g917) & (g960) & (!g961) & (!g962)) + ((!g4) & (g1) & (!g917) & (g960) & (!g961) & (g962)) + ((!g4) & (g1) & (!g917) & (g960) & (g961) & (!g962)) + ((!g4) & (g1) & (!g917) & (g960) & (g961) & (g962)) + ((!g4) & (g1) & (g917) & (!g960) & (!g961) & (!g962)) + ((!g4) & (g1) & (g917) & (!g960) & (!g961) & (g962)) + ((g4) & (!g1) & (!g917) & (!g960) & (!g961) & (!g962)) + ((g4) & (!g1) & (!g917) & (!g960) & (g961) & (!g962)) + ((g4) & (!g1) & (!g917) & (g960) & (!g961) & (!g962)) + ((g4) & (g1) & (!g917) & (!g960) & (!g961) & (!g962)) + ((g4) & (g1) & (!g917) & (!g960) & (!g961) & (g962)) + ((g4) & (g1) & (!g917) & (!g960) & (g961) & (!g962)) + ((g4) & (g1) & (!g917) & (!g960) & (g961) & (g962)) + ((g4) & (g1) & (!g917) & (g960) & (!g961) & (!g962)) + ((g4) & (g1) & (!g917) & (g960) & (!g961) & (g962)) + ((g4) & (g1) & (!g917) & (g960) & (g961) & (!g962)) + ((g4) & (g1) & (!g917) & (g960) & (g961) & (g962)) + ((g4) & (g1) & (g917) & (!g960) & (!g961) & (!g962)) + ((g4) & (g1) & (g917) & (!g960) & (!g961) & (g962)) + ((g4) & (g1) & (g917) & (!g960) & (g961) & (!g962)) + ((g4) & (g1) & (g917) & (!g960) & (g961) & (g962)) + ((g4) & (g1) & (g917) & (g960) & (!g961) & (!g962)) + ((g4) & (g1) & (g917) & (g960) & (!g961) & (g962)));
	assign g964 = (((!ax64x) & (!g914) & (!g915) & (!g916) & (g963)) + ((!ax64x) & (!g914) & (g915) & (!g916) & (!g963)) + ((!ax64x) & (!g914) & (g915) & (!g916) & (g963)) + ((!ax64x) & (!g914) & (g915) & (g916) & (!g963)) + ((!ax64x) & (!g914) & (g915) & (g916) & (g963)) + ((!ax64x) & (g914) & (g915) & (!g916) & (!g963)) + ((!ax64x) & (g914) & (g915) & (g916) & (!g963)) + ((!ax64x) & (g914) & (g915) & (g916) & (g963)) + ((ax64x) & (!g914) & (!g915) & (!g916) & (!g963)) + ((ax64x) & (!g914) & (!g915) & (g916) & (!g963)) + ((ax64x) & (!g914) & (!g915) & (g916) & (g963)) + ((ax64x) & (g914) & (!g915) & (!g916) & (!g963)) + ((ax64x) & (g914) & (!g915) & (!g916) & (g963)) + ((ax64x) & (g914) & (!g915) & (g916) & (!g963)) + ((ax64x) & (g914) & (!g915) & (g916) & (g963)) + ((ax64x) & (g914) & (g915) & (!g916) & (g963)));
	assign g965 = (((!ax60x) & (!ax61x)));
	assign g966 = (((!g914) & (!ax62x) & (!ax63x) & (!g916) & (!g963) & (!g965)) + ((!g914) & (!ax62x) & (!ax63x) & (g916) & (!g963) & (!g965)) + ((!g914) & (!ax62x) & (!ax63x) & (g916) & (g963) & (!g965)) + ((!g914) & (!ax62x) & (ax63x) & (!g916) & (g963) & (!g965)) + ((!g914) & (ax62x) & (ax63x) & (!g916) & (g963) & (!g965)) + ((!g914) & (ax62x) & (ax63x) & (!g916) & (g963) & (g965)) + ((g914) & (!ax62x) & (!ax63x) & (!g916) & (!g963) & (!g965)) + ((g914) & (!ax62x) & (!ax63x) & (!g916) & (!g963) & (g965)) + ((g914) & (!ax62x) & (!ax63x) & (!g916) & (g963) & (!g965)) + ((g914) & (!ax62x) & (!ax63x) & (g916) & (!g963) & (!g965)) + ((g914) & (!ax62x) & (!ax63x) & (g916) & (!g963) & (g965)) + ((g914) & (!ax62x) & (!ax63x) & (g916) & (g963) & (!g965)) + ((g914) & (!ax62x) & (!ax63x) & (g916) & (g963) & (g965)) + ((g914) & (!ax62x) & (ax63x) & (!g916) & (!g963) & (!g965)) + ((g914) & (!ax62x) & (ax63x) & (!g916) & (g963) & (!g965)) + ((g914) & (!ax62x) & (ax63x) & (!g916) & (g963) & (g965)) + ((g914) & (!ax62x) & (ax63x) & (g916) & (!g963) & (!g965)) + ((g914) & (!ax62x) & (ax63x) & (g916) & (g963) & (!g965)) + ((g914) & (ax62x) & (!ax63x) & (!g916) & (g963) & (!g965)) + ((g914) & (ax62x) & (!ax63x) & (!g916) & (g963) & (g965)) + ((g914) & (ax62x) & (ax63x) & (!g916) & (!g963) & (!g965)) + ((g914) & (ax62x) & (ax63x) & (!g916) & (!g963) & (g965)) + ((g914) & (ax62x) & (ax63x) & (!g916) & (g963) & (!g965)) + ((g914) & (ax62x) & (ax63x) & (!g916) & (g963) & (g965)) + ((g914) & (ax62x) & (ax63x) & (g916) & (!g963) & (!g965)) + ((g914) & (ax62x) & (ax63x) & (g916) & (!g963) & (g965)) + ((g914) & (ax62x) & (ax63x) & (g916) & (g963) & (!g965)) + ((g914) & (ax62x) & (ax63x) & (g916) & (g963) & (g965)));
	assign g967 = (((!g4) & (!g960) & (!g961) & (!g916) & (!g963)) + ((!g4) & (!g960) & (!g961) & (g916) & (!g963)) + ((!g4) & (!g960) & (!g961) & (g916) & (g963)) + ((!g4) & (!g960) & (g961) & (!g916) & (g963)) + ((!g4) & (g960) & (g961) & (!g916) & (!g963)) + ((!g4) & (g960) & (g961) & (!g916) & (g963)) + ((!g4) & (g960) & (g961) & (g916) & (!g963)) + ((!g4) & (g960) & (g961) & (g916) & (g963)) + ((g4) & (!g960) & (g961) & (!g916) & (!g963)) + ((g4) & (!g960) & (g961) & (!g916) & (g963)) + ((g4) & (!g960) & (g961) & (g916) & (!g963)) + ((g4) & (!g960) & (g961) & (g916) & (g963)) + ((g4) & (g960) & (!g961) & (!g916) & (!g963)) + ((g4) & (g960) & (!g961) & (g916) & (!g963)) + ((g4) & (g960) & (!g961) & (g916) & (g963)) + ((g4) & (g960) & (g961) & (!g916) & (g963)));
	assign g968 = (((!g8) & (!g919) & (g959) & (!g916) & (!g963)) + ((!g8) & (!g919) & (g959) & (g916) & (!g963)) + ((!g8) & (!g919) & (g959) & (g916) & (g963)) + ((!g8) & (g919) & (!g959) & (!g916) & (!g963)) + ((!g8) & (g919) & (!g959) & (!g916) & (g963)) + ((!g8) & (g919) & (!g959) & (g916) & (!g963)) + ((!g8) & (g919) & (!g959) & (g916) & (g963)) + ((!g8) & (g919) & (g959) & (!g916) & (g963)) + ((g8) & (!g919) & (!g959) & (!g916) & (!g963)) + ((g8) & (!g919) & (!g959) & (g916) & (!g963)) + ((g8) & (!g919) & (!g959) & (g916) & (g963)) + ((g8) & (g919) & (!g959) & (!g916) & (g963)) + ((g8) & (g919) & (g959) & (!g916) & (!g963)) + ((g8) & (g919) & (g959) & (!g916) & (g963)) + ((g8) & (g919) & (g959) & (g916) & (!g963)) + ((g8) & (g919) & (g959) & (g916) & (g963)));
	assign g969 = (((!g18) & (!g27) & (g921) & (g958)) + ((!g18) & (g27) & (!g921) & (g958)) + ((!g18) & (g27) & (g921) & (!g958)) + ((!g18) & (g27) & (g921) & (g958)) + ((g18) & (!g27) & (!g921) & (!g958)) + ((g18) & (!g27) & (!g921) & (g958)) + ((g18) & (!g27) & (g921) & (!g958)) + ((g18) & (g27) & (!g921) & (!g958)));
	assign g970 = (((!g920) & (!g916) & (!g963) & (g969)) + ((!g920) & (g916) & (!g963) & (g969)) + ((!g920) & (g916) & (g963) & (g969)) + ((g920) & (!g916) & (!g963) & (!g969)) + ((g920) & (!g916) & (g963) & (!g969)) + ((g920) & (!g916) & (g963) & (g969)) + ((g920) & (g916) & (!g963) & (!g969)) + ((g920) & (g916) & (g963) & (!g969)));
	assign g971 = (((!g27) & (!g921) & (g958) & (!g916) & (!g963)) + ((!g27) & (!g921) & (g958) & (g916) & (!g963)) + ((!g27) & (!g921) & (g958) & (g916) & (g963)) + ((!g27) & (g921) & (!g958) & (!g916) & (!g963)) + ((!g27) & (g921) & (!g958) & (!g916) & (g963)) + ((!g27) & (g921) & (!g958) & (g916) & (!g963)) + ((!g27) & (g921) & (!g958) & (g916) & (g963)) + ((!g27) & (g921) & (g958) & (!g916) & (g963)) + ((g27) & (!g921) & (!g958) & (!g916) & (!g963)) + ((g27) & (!g921) & (!g958) & (g916) & (!g963)) + ((g27) & (!g921) & (!g958) & (g916) & (g963)) + ((g27) & (g921) & (!g958) & (!g916) & (g963)) + ((g27) & (g921) & (g958) & (!g916) & (!g963)) + ((g27) & (g921) & (g958) & (!g916) & (g963)) + ((g27) & (g921) & (g958) & (g916) & (!g963)) + ((g27) & (g921) & (g958) & (g916) & (g963)));
	assign g972 = (((!g39) & (!g54) & (g923) & (g957)) + ((!g39) & (g54) & (!g923) & (g957)) + ((!g39) & (g54) & (g923) & (!g957)) + ((!g39) & (g54) & (g923) & (g957)) + ((g39) & (!g54) & (!g923) & (!g957)) + ((g39) & (!g54) & (!g923) & (g957)) + ((g39) & (!g54) & (g923) & (!g957)) + ((g39) & (g54) & (!g923) & (!g957)));
	assign g973 = (((!g922) & (!g916) & (!g963) & (g972)) + ((!g922) & (g916) & (!g963) & (g972)) + ((!g922) & (g916) & (g963) & (g972)) + ((g922) & (!g916) & (!g963) & (!g972)) + ((g922) & (!g916) & (g963) & (!g972)) + ((g922) & (!g916) & (g963) & (g972)) + ((g922) & (g916) & (!g963) & (!g972)) + ((g922) & (g916) & (g963) & (!g972)));
	assign g974 = (((!g54) & (!g923) & (g957) & (!g916) & (!g963)) + ((!g54) & (!g923) & (g957) & (g916) & (!g963)) + ((!g54) & (!g923) & (g957) & (g916) & (g963)) + ((!g54) & (g923) & (!g957) & (!g916) & (!g963)) + ((!g54) & (g923) & (!g957) & (!g916) & (g963)) + ((!g54) & (g923) & (!g957) & (g916) & (!g963)) + ((!g54) & (g923) & (!g957) & (g916) & (g963)) + ((!g54) & (g923) & (g957) & (!g916) & (g963)) + ((g54) & (!g923) & (!g957) & (!g916) & (!g963)) + ((g54) & (!g923) & (!g957) & (g916) & (!g963)) + ((g54) & (!g923) & (!g957) & (g916) & (g963)) + ((g54) & (g923) & (!g957) & (!g916) & (g963)) + ((g54) & (g923) & (g957) & (!g916) & (!g963)) + ((g54) & (g923) & (g957) & (!g916) & (g963)) + ((g54) & (g923) & (g957) & (g916) & (!g963)) + ((g54) & (g923) & (g957) & (g916) & (g963)));
	assign g975 = (((!g68) & (!g87) & (g925) & (g956)) + ((!g68) & (g87) & (!g925) & (g956)) + ((!g68) & (g87) & (g925) & (!g956)) + ((!g68) & (g87) & (g925) & (g956)) + ((g68) & (!g87) & (!g925) & (!g956)) + ((g68) & (!g87) & (!g925) & (g956)) + ((g68) & (!g87) & (g925) & (!g956)) + ((g68) & (g87) & (!g925) & (!g956)));
	assign g976 = (((!g924) & (!g916) & (!g963) & (g975)) + ((!g924) & (g916) & (!g963) & (g975)) + ((!g924) & (g916) & (g963) & (g975)) + ((g924) & (!g916) & (!g963) & (!g975)) + ((g924) & (!g916) & (g963) & (!g975)) + ((g924) & (!g916) & (g963) & (g975)) + ((g924) & (g916) & (!g963) & (!g975)) + ((g924) & (g916) & (g963) & (!g975)));
	assign g977 = (((!g87) & (!g925) & (g956) & (!g916) & (!g963)) + ((!g87) & (!g925) & (g956) & (g916) & (!g963)) + ((!g87) & (!g925) & (g956) & (g916) & (g963)) + ((!g87) & (g925) & (!g956) & (!g916) & (!g963)) + ((!g87) & (g925) & (!g956) & (!g916) & (g963)) + ((!g87) & (g925) & (!g956) & (g916) & (!g963)) + ((!g87) & (g925) & (!g956) & (g916) & (g963)) + ((!g87) & (g925) & (g956) & (!g916) & (g963)) + ((g87) & (!g925) & (!g956) & (!g916) & (!g963)) + ((g87) & (!g925) & (!g956) & (g916) & (!g963)) + ((g87) & (!g925) & (!g956) & (g916) & (g963)) + ((g87) & (g925) & (!g956) & (!g916) & (g963)) + ((g87) & (g925) & (g956) & (!g916) & (!g963)) + ((g87) & (g925) & (g956) & (!g916) & (g963)) + ((g87) & (g925) & (g956) & (g916) & (!g963)) + ((g87) & (g925) & (g956) & (g916) & (g963)));
	assign g978 = (((!g104) & (!g127) & (g927) & (g955)) + ((!g104) & (g127) & (!g927) & (g955)) + ((!g104) & (g127) & (g927) & (!g955)) + ((!g104) & (g127) & (g927) & (g955)) + ((g104) & (!g127) & (!g927) & (!g955)) + ((g104) & (!g127) & (!g927) & (g955)) + ((g104) & (!g127) & (g927) & (!g955)) + ((g104) & (g127) & (!g927) & (!g955)));
	assign g979 = (((!g926) & (!g916) & (!g963) & (g978)) + ((!g926) & (g916) & (!g963) & (g978)) + ((!g926) & (g916) & (g963) & (g978)) + ((g926) & (!g916) & (!g963) & (!g978)) + ((g926) & (!g916) & (g963) & (!g978)) + ((g926) & (!g916) & (g963) & (g978)) + ((g926) & (g916) & (!g963) & (!g978)) + ((g926) & (g916) & (g963) & (!g978)));
	assign g980 = (((!g127) & (!g927) & (g955) & (!g916) & (!g963)) + ((!g127) & (!g927) & (g955) & (g916) & (!g963)) + ((!g127) & (!g927) & (g955) & (g916) & (g963)) + ((!g127) & (g927) & (!g955) & (!g916) & (!g963)) + ((!g127) & (g927) & (!g955) & (!g916) & (g963)) + ((!g127) & (g927) & (!g955) & (g916) & (!g963)) + ((!g127) & (g927) & (!g955) & (g916) & (g963)) + ((!g127) & (g927) & (g955) & (!g916) & (g963)) + ((g127) & (!g927) & (!g955) & (!g916) & (!g963)) + ((g127) & (!g927) & (!g955) & (g916) & (!g963)) + ((g127) & (!g927) & (!g955) & (g916) & (g963)) + ((g127) & (g927) & (!g955) & (!g916) & (g963)) + ((g127) & (g927) & (g955) & (!g916) & (!g963)) + ((g127) & (g927) & (g955) & (!g916) & (g963)) + ((g127) & (g927) & (g955) & (g916) & (!g963)) + ((g127) & (g927) & (g955) & (g916) & (g963)));
	assign g981 = (((!g147) & (!g174) & (g929) & (g954)) + ((!g147) & (g174) & (!g929) & (g954)) + ((!g147) & (g174) & (g929) & (!g954)) + ((!g147) & (g174) & (g929) & (g954)) + ((g147) & (!g174) & (!g929) & (!g954)) + ((g147) & (!g174) & (!g929) & (g954)) + ((g147) & (!g174) & (g929) & (!g954)) + ((g147) & (g174) & (!g929) & (!g954)));
	assign g982 = (((!g928) & (!g916) & (!g963) & (g981)) + ((!g928) & (g916) & (!g963) & (g981)) + ((!g928) & (g916) & (g963) & (g981)) + ((g928) & (!g916) & (!g963) & (!g981)) + ((g928) & (!g916) & (g963) & (!g981)) + ((g928) & (!g916) & (g963) & (g981)) + ((g928) & (g916) & (!g963) & (!g981)) + ((g928) & (g916) & (g963) & (!g981)));
	assign g983 = (((!g174) & (!g929) & (g954) & (!g916) & (!g963)) + ((!g174) & (!g929) & (g954) & (g916) & (!g963)) + ((!g174) & (!g929) & (g954) & (g916) & (g963)) + ((!g174) & (g929) & (!g954) & (!g916) & (!g963)) + ((!g174) & (g929) & (!g954) & (!g916) & (g963)) + ((!g174) & (g929) & (!g954) & (g916) & (!g963)) + ((!g174) & (g929) & (!g954) & (g916) & (g963)) + ((!g174) & (g929) & (g954) & (!g916) & (g963)) + ((g174) & (!g929) & (!g954) & (!g916) & (!g963)) + ((g174) & (!g929) & (!g954) & (g916) & (!g963)) + ((g174) & (!g929) & (!g954) & (g916) & (g963)) + ((g174) & (g929) & (!g954) & (!g916) & (g963)) + ((g174) & (g929) & (g954) & (!g916) & (!g963)) + ((g174) & (g929) & (g954) & (!g916) & (g963)) + ((g174) & (g929) & (g954) & (g916) & (!g963)) + ((g174) & (g929) & (g954) & (g916) & (g963)));
	assign g984 = (((!g198) & (!g229) & (g931) & (g953)) + ((!g198) & (g229) & (!g931) & (g953)) + ((!g198) & (g229) & (g931) & (!g953)) + ((!g198) & (g229) & (g931) & (g953)) + ((g198) & (!g229) & (!g931) & (!g953)) + ((g198) & (!g229) & (!g931) & (g953)) + ((g198) & (!g229) & (g931) & (!g953)) + ((g198) & (g229) & (!g931) & (!g953)));
	assign g985 = (((!g930) & (!g916) & (!g963) & (g984)) + ((!g930) & (g916) & (!g963) & (g984)) + ((!g930) & (g916) & (g963) & (g984)) + ((g930) & (!g916) & (!g963) & (!g984)) + ((g930) & (!g916) & (g963) & (!g984)) + ((g930) & (!g916) & (g963) & (g984)) + ((g930) & (g916) & (!g963) & (!g984)) + ((g930) & (g916) & (g963) & (!g984)));
	assign g986 = (((!g229) & (!g931) & (g953) & (!g916) & (!g963)) + ((!g229) & (!g931) & (g953) & (g916) & (!g963)) + ((!g229) & (!g931) & (g953) & (g916) & (g963)) + ((!g229) & (g931) & (!g953) & (!g916) & (!g963)) + ((!g229) & (g931) & (!g953) & (!g916) & (g963)) + ((!g229) & (g931) & (!g953) & (g916) & (!g963)) + ((!g229) & (g931) & (!g953) & (g916) & (g963)) + ((!g229) & (g931) & (g953) & (!g916) & (g963)) + ((g229) & (!g931) & (!g953) & (!g916) & (!g963)) + ((g229) & (!g931) & (!g953) & (g916) & (!g963)) + ((g229) & (!g931) & (!g953) & (g916) & (g963)) + ((g229) & (g931) & (!g953) & (!g916) & (g963)) + ((g229) & (g931) & (g953) & (!g916) & (!g963)) + ((g229) & (g931) & (g953) & (!g916) & (g963)) + ((g229) & (g931) & (g953) & (g916) & (!g963)) + ((g229) & (g931) & (g953) & (g916) & (g963)));
	assign g987 = (((!g255) & (!g290) & (g933) & (g952)) + ((!g255) & (g290) & (!g933) & (g952)) + ((!g255) & (g290) & (g933) & (!g952)) + ((!g255) & (g290) & (g933) & (g952)) + ((g255) & (!g290) & (!g933) & (!g952)) + ((g255) & (!g290) & (!g933) & (g952)) + ((g255) & (!g290) & (g933) & (!g952)) + ((g255) & (g290) & (!g933) & (!g952)));
	assign g988 = (((!g932) & (!g916) & (!g963) & (g987)) + ((!g932) & (g916) & (!g963) & (g987)) + ((!g932) & (g916) & (g963) & (g987)) + ((g932) & (!g916) & (!g963) & (!g987)) + ((g932) & (!g916) & (g963) & (!g987)) + ((g932) & (!g916) & (g963) & (g987)) + ((g932) & (g916) & (!g963) & (!g987)) + ((g932) & (g916) & (g963) & (!g987)));
	assign g989 = (((!g290) & (!g933) & (g952) & (!g916) & (!g963)) + ((!g290) & (!g933) & (g952) & (g916) & (!g963)) + ((!g290) & (!g933) & (g952) & (g916) & (g963)) + ((!g290) & (g933) & (!g952) & (!g916) & (!g963)) + ((!g290) & (g933) & (!g952) & (!g916) & (g963)) + ((!g290) & (g933) & (!g952) & (g916) & (!g963)) + ((!g290) & (g933) & (!g952) & (g916) & (g963)) + ((!g290) & (g933) & (g952) & (!g916) & (g963)) + ((g290) & (!g933) & (!g952) & (!g916) & (!g963)) + ((g290) & (!g933) & (!g952) & (g916) & (!g963)) + ((g290) & (!g933) & (!g952) & (g916) & (g963)) + ((g290) & (g933) & (!g952) & (!g916) & (g963)) + ((g290) & (g933) & (g952) & (!g916) & (!g963)) + ((g290) & (g933) & (g952) & (!g916) & (g963)) + ((g290) & (g933) & (g952) & (g916) & (!g963)) + ((g290) & (g933) & (g952) & (g916) & (g963)));
	assign g990 = (((!g319) & (!g358) & (g935) & (g951)) + ((!g319) & (g358) & (!g935) & (g951)) + ((!g319) & (g358) & (g935) & (!g951)) + ((!g319) & (g358) & (g935) & (g951)) + ((g319) & (!g358) & (!g935) & (!g951)) + ((g319) & (!g358) & (!g935) & (g951)) + ((g319) & (!g358) & (g935) & (!g951)) + ((g319) & (g358) & (!g935) & (!g951)));
	assign g991 = (((!g934) & (!g916) & (!g963) & (g990)) + ((!g934) & (g916) & (!g963) & (g990)) + ((!g934) & (g916) & (g963) & (g990)) + ((g934) & (!g916) & (!g963) & (!g990)) + ((g934) & (!g916) & (g963) & (!g990)) + ((g934) & (!g916) & (g963) & (g990)) + ((g934) & (g916) & (!g963) & (!g990)) + ((g934) & (g916) & (g963) & (!g990)));
	assign g992 = (((!g358) & (!g935) & (g951) & (!g916) & (!g963)) + ((!g358) & (!g935) & (g951) & (g916) & (!g963)) + ((!g358) & (!g935) & (g951) & (g916) & (g963)) + ((!g358) & (g935) & (!g951) & (!g916) & (!g963)) + ((!g358) & (g935) & (!g951) & (!g916) & (g963)) + ((!g358) & (g935) & (!g951) & (g916) & (!g963)) + ((!g358) & (g935) & (!g951) & (g916) & (g963)) + ((!g358) & (g935) & (g951) & (!g916) & (g963)) + ((g358) & (!g935) & (!g951) & (!g916) & (!g963)) + ((g358) & (!g935) & (!g951) & (g916) & (!g963)) + ((g358) & (!g935) & (!g951) & (g916) & (g963)) + ((g358) & (g935) & (!g951) & (!g916) & (g963)) + ((g358) & (g935) & (g951) & (!g916) & (!g963)) + ((g358) & (g935) & (g951) & (!g916) & (g963)) + ((g358) & (g935) & (g951) & (g916) & (!g963)) + ((g358) & (g935) & (g951) & (g916) & (g963)));
	assign g993 = (((!g390) & (!g433) & (g937) & (g950)) + ((!g390) & (g433) & (!g937) & (g950)) + ((!g390) & (g433) & (g937) & (!g950)) + ((!g390) & (g433) & (g937) & (g950)) + ((g390) & (!g433) & (!g937) & (!g950)) + ((g390) & (!g433) & (!g937) & (g950)) + ((g390) & (!g433) & (g937) & (!g950)) + ((g390) & (g433) & (!g937) & (!g950)));
	assign g994 = (((!g936) & (!g916) & (!g963) & (g993)) + ((!g936) & (g916) & (!g963) & (g993)) + ((!g936) & (g916) & (g963) & (g993)) + ((g936) & (!g916) & (!g963) & (!g993)) + ((g936) & (!g916) & (g963) & (!g993)) + ((g936) & (!g916) & (g963) & (g993)) + ((g936) & (g916) & (!g963) & (!g993)) + ((g936) & (g916) & (g963) & (!g993)));
	assign g995 = (((!g433) & (!g937) & (g950) & (!g916) & (!g963)) + ((!g433) & (!g937) & (g950) & (g916) & (!g963)) + ((!g433) & (!g937) & (g950) & (g916) & (g963)) + ((!g433) & (g937) & (!g950) & (!g916) & (!g963)) + ((!g433) & (g937) & (!g950) & (!g916) & (g963)) + ((!g433) & (g937) & (!g950) & (g916) & (!g963)) + ((!g433) & (g937) & (!g950) & (g916) & (g963)) + ((!g433) & (g937) & (g950) & (!g916) & (g963)) + ((g433) & (!g937) & (!g950) & (!g916) & (!g963)) + ((g433) & (!g937) & (!g950) & (g916) & (!g963)) + ((g433) & (!g937) & (!g950) & (g916) & (g963)) + ((g433) & (g937) & (!g950) & (!g916) & (g963)) + ((g433) & (g937) & (g950) & (!g916) & (!g963)) + ((g433) & (g937) & (g950) & (!g916) & (g963)) + ((g433) & (g937) & (g950) & (g916) & (!g963)) + ((g433) & (g937) & (g950) & (g916) & (g963)));
	assign g996 = (((!g468) & (!g515) & (g939) & (g949)) + ((!g468) & (g515) & (!g939) & (g949)) + ((!g468) & (g515) & (g939) & (!g949)) + ((!g468) & (g515) & (g939) & (g949)) + ((g468) & (!g515) & (!g939) & (!g949)) + ((g468) & (!g515) & (!g939) & (g949)) + ((g468) & (!g515) & (g939) & (!g949)) + ((g468) & (g515) & (!g939) & (!g949)));
	assign g997 = (((!g938) & (!g916) & (!g963) & (g996)) + ((!g938) & (g916) & (!g963) & (g996)) + ((!g938) & (g916) & (g963) & (g996)) + ((g938) & (!g916) & (!g963) & (!g996)) + ((g938) & (!g916) & (g963) & (!g996)) + ((g938) & (!g916) & (g963) & (g996)) + ((g938) & (g916) & (!g963) & (!g996)) + ((g938) & (g916) & (g963) & (!g996)));
	assign g998 = (((!g515) & (!g939) & (g949) & (!g916) & (!g963)) + ((!g515) & (!g939) & (g949) & (g916) & (!g963)) + ((!g515) & (!g939) & (g949) & (g916) & (g963)) + ((!g515) & (g939) & (!g949) & (!g916) & (!g963)) + ((!g515) & (g939) & (!g949) & (!g916) & (g963)) + ((!g515) & (g939) & (!g949) & (g916) & (!g963)) + ((!g515) & (g939) & (!g949) & (g916) & (g963)) + ((!g515) & (g939) & (g949) & (!g916) & (g963)) + ((g515) & (!g939) & (!g949) & (!g916) & (!g963)) + ((g515) & (!g939) & (!g949) & (g916) & (!g963)) + ((g515) & (!g939) & (!g949) & (g916) & (g963)) + ((g515) & (g939) & (!g949) & (!g916) & (g963)) + ((g515) & (g939) & (g949) & (!g916) & (!g963)) + ((g515) & (g939) & (g949) & (!g916) & (g963)) + ((g515) & (g939) & (g949) & (g916) & (!g963)) + ((g515) & (g939) & (g949) & (g916) & (g963)));
	assign g999 = (((!g553) & (!g604) & (g941) & (g948)) + ((!g553) & (g604) & (!g941) & (g948)) + ((!g553) & (g604) & (g941) & (!g948)) + ((!g553) & (g604) & (g941) & (g948)) + ((g553) & (!g604) & (!g941) & (!g948)) + ((g553) & (!g604) & (!g941) & (g948)) + ((g553) & (!g604) & (g941) & (!g948)) + ((g553) & (g604) & (!g941) & (!g948)));
	assign g1000 = (((!g940) & (!g916) & (!g963) & (g999)) + ((!g940) & (g916) & (!g963) & (g999)) + ((!g940) & (g916) & (g963) & (g999)) + ((g940) & (!g916) & (!g963) & (!g999)) + ((g940) & (!g916) & (g963) & (!g999)) + ((g940) & (!g916) & (g963) & (g999)) + ((g940) & (g916) & (!g963) & (!g999)) + ((g940) & (g916) & (g963) & (!g999)));
	assign g1001 = (((!g604) & (!g941) & (g948) & (!g916) & (!g963)) + ((!g604) & (!g941) & (g948) & (g916) & (!g963)) + ((!g604) & (!g941) & (g948) & (g916) & (g963)) + ((!g604) & (g941) & (!g948) & (!g916) & (!g963)) + ((!g604) & (g941) & (!g948) & (!g916) & (g963)) + ((!g604) & (g941) & (!g948) & (g916) & (!g963)) + ((!g604) & (g941) & (!g948) & (g916) & (g963)) + ((!g604) & (g941) & (g948) & (!g916) & (g963)) + ((g604) & (!g941) & (!g948) & (!g916) & (!g963)) + ((g604) & (!g941) & (!g948) & (g916) & (!g963)) + ((g604) & (!g941) & (!g948) & (g916) & (g963)) + ((g604) & (g941) & (!g948) & (!g916) & (g963)) + ((g604) & (g941) & (g948) & (!g916) & (!g963)) + ((g604) & (g941) & (g948) & (!g916) & (g963)) + ((g604) & (g941) & (g948) & (g916) & (!g963)) + ((g604) & (g941) & (g948) & (g916) & (g963)));
	assign g1002 = (((!g645) & (!g700) & (g943) & (g947)) + ((!g645) & (g700) & (!g943) & (g947)) + ((!g645) & (g700) & (g943) & (!g947)) + ((!g645) & (g700) & (g943) & (g947)) + ((g645) & (!g700) & (!g943) & (!g947)) + ((g645) & (!g700) & (!g943) & (g947)) + ((g645) & (!g700) & (g943) & (!g947)) + ((g645) & (g700) & (!g943) & (!g947)));
	assign g1003 = (((!g942) & (!g916) & (!g963) & (g1002)) + ((!g942) & (g916) & (!g963) & (g1002)) + ((!g942) & (g916) & (g963) & (g1002)) + ((g942) & (!g916) & (!g963) & (!g1002)) + ((g942) & (!g916) & (g963) & (!g1002)) + ((g942) & (!g916) & (g963) & (g1002)) + ((g942) & (g916) & (!g963) & (!g1002)) + ((g942) & (g916) & (g963) & (!g1002)));
	assign g1004 = (((!g700) & (!g943) & (g947) & (!g916) & (!g963)) + ((!g700) & (!g943) & (g947) & (g916) & (!g963)) + ((!g700) & (!g943) & (g947) & (g916) & (g963)) + ((!g700) & (g943) & (!g947) & (!g916) & (!g963)) + ((!g700) & (g943) & (!g947) & (!g916) & (g963)) + ((!g700) & (g943) & (!g947) & (g916) & (!g963)) + ((!g700) & (g943) & (!g947) & (g916) & (g963)) + ((!g700) & (g943) & (g947) & (!g916) & (g963)) + ((g700) & (!g943) & (!g947) & (!g916) & (!g963)) + ((g700) & (!g943) & (!g947) & (g916) & (!g963)) + ((g700) & (!g943) & (!g947) & (g916) & (g963)) + ((g700) & (g943) & (!g947) & (!g916) & (g963)) + ((g700) & (g943) & (g947) & (!g916) & (!g963)) + ((g700) & (g943) & (g947) & (!g916) & (g963)) + ((g700) & (g943) & (g947) & (g916) & (!g963)) + ((g700) & (g943) & (g947) & (g916) & (g963)));
	assign g1005 = (((!g744) & (!g803) & (g945) & (g946)) + ((!g744) & (g803) & (!g945) & (g946)) + ((!g744) & (g803) & (g945) & (!g946)) + ((!g744) & (g803) & (g945) & (g946)) + ((g744) & (!g803) & (!g945) & (!g946)) + ((g744) & (!g803) & (!g945) & (g946)) + ((g744) & (!g803) & (g945) & (!g946)) + ((g744) & (g803) & (!g945) & (!g946)));
	assign g1006 = (((!g944) & (!g916) & (!g963) & (g1005)) + ((!g944) & (g916) & (!g963) & (g1005)) + ((!g944) & (g916) & (g963) & (g1005)) + ((g944) & (!g916) & (!g963) & (!g1005)) + ((g944) & (!g916) & (g963) & (!g1005)) + ((g944) & (!g916) & (g963) & (g1005)) + ((g944) & (g916) & (!g963) & (!g1005)) + ((g944) & (g916) & (g963) & (!g1005)));
	assign g1007 = (((!g803) & (!g945) & (g946) & (!g916) & (!g963)) + ((!g803) & (!g945) & (g946) & (g916) & (!g963)) + ((!g803) & (!g945) & (g946) & (g916) & (g963)) + ((!g803) & (g945) & (!g946) & (!g916) & (!g963)) + ((!g803) & (g945) & (!g946) & (!g916) & (g963)) + ((!g803) & (g945) & (!g946) & (g916) & (!g963)) + ((!g803) & (g945) & (!g946) & (g916) & (g963)) + ((!g803) & (g945) & (g946) & (!g916) & (g963)) + ((g803) & (!g945) & (!g946) & (!g916) & (!g963)) + ((g803) & (!g945) & (!g946) & (g916) & (!g963)) + ((g803) & (!g945) & (!g946) & (g916) & (g963)) + ((g803) & (g945) & (!g946) & (!g916) & (g963)) + ((g803) & (g945) & (g946) & (!g916) & (!g963)) + ((g803) & (g945) & (g946) & (!g916) & (g963)) + ((g803) & (g945) & (g946) & (g916) & (!g963)) + ((g803) & (g945) & (g946) & (g916) & (g963)));
	assign g1008 = (((!ax64x) & (!g851) & (!g914) & (!g915)) + ((!ax64x) & (!g851) & (g914) & (!g915)) + ((!ax64x) & (g851) & (!g914) & (g915)) + ((!ax64x) & (g851) & (g914) & (g915)) + ((ax64x) & (!g851) & (g914) & (!g915)) + ((ax64x) & (!g851) & (g914) & (g915)) + ((ax64x) & (g851) & (!g914) & (!g915)) + ((ax64x) & (g851) & (!g914) & (g915)));
	assign g1009 = (((!ax64x) & (!ax65x) & (!g914) & (!g916) & (!g963) & (!g1008)) + ((!ax64x) & (!ax65x) & (!g914) & (!g916) & (g963) & (!g1008)) + ((!ax64x) & (!ax65x) & (!g914) & (!g916) & (g963) & (g1008)) + ((!ax64x) & (!ax65x) & (!g914) & (g916) & (!g963) & (!g1008)) + ((!ax64x) & (!ax65x) & (!g914) & (g916) & (g963) & (!g1008)) + ((!ax64x) & (!ax65x) & (g914) & (!g916) & (!g963) & (g1008)) + ((!ax64x) & (!ax65x) & (g914) & (g916) & (!g963) & (g1008)) + ((!ax64x) & (!ax65x) & (g914) & (g916) & (g963) & (g1008)) + ((!ax64x) & (ax65x) & (!g914) & (!g916) & (!g963) & (g1008)) + ((!ax64x) & (ax65x) & (!g914) & (g916) & (!g963) & (g1008)) + ((!ax64x) & (ax65x) & (!g914) & (g916) & (g963) & (g1008)) + ((!ax64x) & (ax65x) & (g914) & (!g916) & (!g963) & (!g1008)) + ((!ax64x) & (ax65x) & (g914) & (!g916) & (g963) & (!g1008)) + ((!ax64x) & (ax65x) & (g914) & (!g916) & (g963) & (g1008)) + ((!ax64x) & (ax65x) & (g914) & (g916) & (!g963) & (!g1008)) + ((!ax64x) & (ax65x) & (g914) & (g916) & (g963) & (!g1008)) + ((ax64x) & (!ax65x) & (!g914) & (!g916) & (!g963) & (g1008)) + ((ax64x) & (!ax65x) & (!g914) & (g916) & (!g963) & (g1008)) + ((ax64x) & (!ax65x) & (!g914) & (g916) & (g963) & (g1008)) + ((ax64x) & (!ax65x) & (g914) & (!g916) & (!g963) & (g1008)) + ((ax64x) & (!ax65x) & (g914) & (g916) & (!g963) & (g1008)) + ((ax64x) & (!ax65x) & (g914) & (g916) & (g963) & (g1008)) + ((ax64x) & (ax65x) & (!g914) & (!g916) & (!g963) & (!g1008)) + ((ax64x) & (ax65x) & (!g914) & (!g916) & (g963) & (!g1008)) + ((ax64x) & (ax65x) & (!g914) & (!g916) & (g963) & (g1008)) + ((ax64x) & (ax65x) & (!g914) & (g916) & (!g963) & (!g1008)) + ((ax64x) & (ax65x) & (!g914) & (g916) & (g963) & (!g1008)) + ((ax64x) & (ax65x) & (g914) & (!g916) & (!g963) & (!g1008)) + ((ax64x) & (ax65x) & (g914) & (!g916) & (g963) & (!g1008)) + ((ax64x) & (ax65x) & (g914) & (!g916) & (g963) & (g1008)) + ((ax64x) & (ax65x) & (g914) & (g916) & (!g963) & (!g1008)) + ((ax64x) & (ax65x) & (g914) & (g916) & (g963) & (!g1008)));
	assign g1010 = (((!g803) & (!g851) & (g1009) & (g964) & (g966)) + ((!g803) & (g851) & (g1009) & (!g964) & (g966)) + ((!g803) & (g851) & (g1009) & (g964) & (!g966)) + ((!g803) & (g851) & (g1009) & (g964) & (g966)) + ((g803) & (!g851) & (!g1009) & (g964) & (g966)) + ((g803) & (!g851) & (g1009) & (!g964) & (!g966)) + ((g803) & (!g851) & (g1009) & (!g964) & (g966)) + ((g803) & (!g851) & (g1009) & (g964) & (!g966)) + ((g803) & (!g851) & (g1009) & (g964) & (g966)) + ((g803) & (g851) & (!g1009) & (!g964) & (g966)) + ((g803) & (g851) & (!g1009) & (g964) & (!g966)) + ((g803) & (g851) & (!g1009) & (g964) & (g966)) + ((g803) & (g851) & (g1009) & (!g964) & (!g966)) + ((g803) & (g851) & (g1009) & (!g964) & (g966)) + ((g803) & (g851) & (g1009) & (g964) & (!g966)) + ((g803) & (g851) & (g1009) & (g964) & (g966)));
	assign g1011 = (((!g700) & (!g744) & (g1006) & (g1007) & (g1010)) + ((!g700) & (g744) & (g1006) & (!g1007) & (g1010)) + ((!g700) & (g744) & (g1006) & (g1007) & (!g1010)) + ((!g700) & (g744) & (g1006) & (g1007) & (g1010)) + ((g700) & (!g744) & (!g1006) & (g1007) & (g1010)) + ((g700) & (!g744) & (g1006) & (!g1007) & (!g1010)) + ((g700) & (!g744) & (g1006) & (!g1007) & (g1010)) + ((g700) & (!g744) & (g1006) & (g1007) & (!g1010)) + ((g700) & (!g744) & (g1006) & (g1007) & (g1010)) + ((g700) & (g744) & (!g1006) & (!g1007) & (g1010)) + ((g700) & (g744) & (!g1006) & (g1007) & (!g1010)) + ((g700) & (g744) & (!g1006) & (g1007) & (g1010)) + ((g700) & (g744) & (g1006) & (!g1007) & (!g1010)) + ((g700) & (g744) & (g1006) & (!g1007) & (g1010)) + ((g700) & (g744) & (g1006) & (g1007) & (!g1010)) + ((g700) & (g744) & (g1006) & (g1007) & (g1010)));
	assign g1012 = (((!g604) & (!g645) & (g1003) & (g1004) & (g1011)) + ((!g604) & (g645) & (g1003) & (!g1004) & (g1011)) + ((!g604) & (g645) & (g1003) & (g1004) & (!g1011)) + ((!g604) & (g645) & (g1003) & (g1004) & (g1011)) + ((g604) & (!g645) & (!g1003) & (g1004) & (g1011)) + ((g604) & (!g645) & (g1003) & (!g1004) & (!g1011)) + ((g604) & (!g645) & (g1003) & (!g1004) & (g1011)) + ((g604) & (!g645) & (g1003) & (g1004) & (!g1011)) + ((g604) & (!g645) & (g1003) & (g1004) & (g1011)) + ((g604) & (g645) & (!g1003) & (!g1004) & (g1011)) + ((g604) & (g645) & (!g1003) & (g1004) & (!g1011)) + ((g604) & (g645) & (!g1003) & (g1004) & (g1011)) + ((g604) & (g645) & (g1003) & (!g1004) & (!g1011)) + ((g604) & (g645) & (g1003) & (!g1004) & (g1011)) + ((g604) & (g645) & (g1003) & (g1004) & (!g1011)) + ((g604) & (g645) & (g1003) & (g1004) & (g1011)));
	assign g1013 = (((!g515) & (!g553) & (g1000) & (g1001) & (g1012)) + ((!g515) & (g553) & (g1000) & (!g1001) & (g1012)) + ((!g515) & (g553) & (g1000) & (g1001) & (!g1012)) + ((!g515) & (g553) & (g1000) & (g1001) & (g1012)) + ((g515) & (!g553) & (!g1000) & (g1001) & (g1012)) + ((g515) & (!g553) & (g1000) & (!g1001) & (!g1012)) + ((g515) & (!g553) & (g1000) & (!g1001) & (g1012)) + ((g515) & (!g553) & (g1000) & (g1001) & (!g1012)) + ((g515) & (!g553) & (g1000) & (g1001) & (g1012)) + ((g515) & (g553) & (!g1000) & (!g1001) & (g1012)) + ((g515) & (g553) & (!g1000) & (g1001) & (!g1012)) + ((g515) & (g553) & (!g1000) & (g1001) & (g1012)) + ((g515) & (g553) & (g1000) & (!g1001) & (!g1012)) + ((g515) & (g553) & (g1000) & (!g1001) & (g1012)) + ((g515) & (g553) & (g1000) & (g1001) & (!g1012)) + ((g515) & (g553) & (g1000) & (g1001) & (g1012)));
	assign g1014 = (((!g433) & (!g468) & (g997) & (g998) & (g1013)) + ((!g433) & (g468) & (g997) & (!g998) & (g1013)) + ((!g433) & (g468) & (g997) & (g998) & (!g1013)) + ((!g433) & (g468) & (g997) & (g998) & (g1013)) + ((g433) & (!g468) & (!g997) & (g998) & (g1013)) + ((g433) & (!g468) & (g997) & (!g998) & (!g1013)) + ((g433) & (!g468) & (g997) & (!g998) & (g1013)) + ((g433) & (!g468) & (g997) & (g998) & (!g1013)) + ((g433) & (!g468) & (g997) & (g998) & (g1013)) + ((g433) & (g468) & (!g997) & (!g998) & (g1013)) + ((g433) & (g468) & (!g997) & (g998) & (!g1013)) + ((g433) & (g468) & (!g997) & (g998) & (g1013)) + ((g433) & (g468) & (g997) & (!g998) & (!g1013)) + ((g433) & (g468) & (g997) & (!g998) & (g1013)) + ((g433) & (g468) & (g997) & (g998) & (!g1013)) + ((g433) & (g468) & (g997) & (g998) & (g1013)));
	assign g1015 = (((!g358) & (!g390) & (g994) & (g995) & (g1014)) + ((!g358) & (g390) & (g994) & (!g995) & (g1014)) + ((!g358) & (g390) & (g994) & (g995) & (!g1014)) + ((!g358) & (g390) & (g994) & (g995) & (g1014)) + ((g358) & (!g390) & (!g994) & (g995) & (g1014)) + ((g358) & (!g390) & (g994) & (!g995) & (!g1014)) + ((g358) & (!g390) & (g994) & (!g995) & (g1014)) + ((g358) & (!g390) & (g994) & (g995) & (!g1014)) + ((g358) & (!g390) & (g994) & (g995) & (g1014)) + ((g358) & (g390) & (!g994) & (!g995) & (g1014)) + ((g358) & (g390) & (!g994) & (g995) & (!g1014)) + ((g358) & (g390) & (!g994) & (g995) & (g1014)) + ((g358) & (g390) & (g994) & (!g995) & (!g1014)) + ((g358) & (g390) & (g994) & (!g995) & (g1014)) + ((g358) & (g390) & (g994) & (g995) & (!g1014)) + ((g358) & (g390) & (g994) & (g995) & (g1014)));
	assign g1016 = (((!g290) & (!g319) & (g991) & (g992) & (g1015)) + ((!g290) & (g319) & (g991) & (!g992) & (g1015)) + ((!g290) & (g319) & (g991) & (g992) & (!g1015)) + ((!g290) & (g319) & (g991) & (g992) & (g1015)) + ((g290) & (!g319) & (!g991) & (g992) & (g1015)) + ((g290) & (!g319) & (g991) & (!g992) & (!g1015)) + ((g290) & (!g319) & (g991) & (!g992) & (g1015)) + ((g290) & (!g319) & (g991) & (g992) & (!g1015)) + ((g290) & (!g319) & (g991) & (g992) & (g1015)) + ((g290) & (g319) & (!g991) & (!g992) & (g1015)) + ((g290) & (g319) & (!g991) & (g992) & (!g1015)) + ((g290) & (g319) & (!g991) & (g992) & (g1015)) + ((g290) & (g319) & (g991) & (!g992) & (!g1015)) + ((g290) & (g319) & (g991) & (!g992) & (g1015)) + ((g290) & (g319) & (g991) & (g992) & (!g1015)) + ((g290) & (g319) & (g991) & (g992) & (g1015)));
	assign g1017 = (((!g229) & (!g255) & (g988) & (g989) & (g1016)) + ((!g229) & (g255) & (g988) & (!g989) & (g1016)) + ((!g229) & (g255) & (g988) & (g989) & (!g1016)) + ((!g229) & (g255) & (g988) & (g989) & (g1016)) + ((g229) & (!g255) & (!g988) & (g989) & (g1016)) + ((g229) & (!g255) & (g988) & (!g989) & (!g1016)) + ((g229) & (!g255) & (g988) & (!g989) & (g1016)) + ((g229) & (!g255) & (g988) & (g989) & (!g1016)) + ((g229) & (!g255) & (g988) & (g989) & (g1016)) + ((g229) & (g255) & (!g988) & (!g989) & (g1016)) + ((g229) & (g255) & (!g988) & (g989) & (!g1016)) + ((g229) & (g255) & (!g988) & (g989) & (g1016)) + ((g229) & (g255) & (g988) & (!g989) & (!g1016)) + ((g229) & (g255) & (g988) & (!g989) & (g1016)) + ((g229) & (g255) & (g988) & (g989) & (!g1016)) + ((g229) & (g255) & (g988) & (g989) & (g1016)));
	assign g1018 = (((!g174) & (!g198) & (g985) & (g986) & (g1017)) + ((!g174) & (g198) & (g985) & (!g986) & (g1017)) + ((!g174) & (g198) & (g985) & (g986) & (!g1017)) + ((!g174) & (g198) & (g985) & (g986) & (g1017)) + ((g174) & (!g198) & (!g985) & (g986) & (g1017)) + ((g174) & (!g198) & (g985) & (!g986) & (!g1017)) + ((g174) & (!g198) & (g985) & (!g986) & (g1017)) + ((g174) & (!g198) & (g985) & (g986) & (!g1017)) + ((g174) & (!g198) & (g985) & (g986) & (g1017)) + ((g174) & (g198) & (!g985) & (!g986) & (g1017)) + ((g174) & (g198) & (!g985) & (g986) & (!g1017)) + ((g174) & (g198) & (!g985) & (g986) & (g1017)) + ((g174) & (g198) & (g985) & (!g986) & (!g1017)) + ((g174) & (g198) & (g985) & (!g986) & (g1017)) + ((g174) & (g198) & (g985) & (g986) & (!g1017)) + ((g174) & (g198) & (g985) & (g986) & (g1017)));
	assign g1019 = (((!g127) & (!g147) & (g982) & (g983) & (g1018)) + ((!g127) & (g147) & (g982) & (!g983) & (g1018)) + ((!g127) & (g147) & (g982) & (g983) & (!g1018)) + ((!g127) & (g147) & (g982) & (g983) & (g1018)) + ((g127) & (!g147) & (!g982) & (g983) & (g1018)) + ((g127) & (!g147) & (g982) & (!g983) & (!g1018)) + ((g127) & (!g147) & (g982) & (!g983) & (g1018)) + ((g127) & (!g147) & (g982) & (g983) & (!g1018)) + ((g127) & (!g147) & (g982) & (g983) & (g1018)) + ((g127) & (g147) & (!g982) & (!g983) & (g1018)) + ((g127) & (g147) & (!g982) & (g983) & (!g1018)) + ((g127) & (g147) & (!g982) & (g983) & (g1018)) + ((g127) & (g147) & (g982) & (!g983) & (!g1018)) + ((g127) & (g147) & (g982) & (!g983) & (g1018)) + ((g127) & (g147) & (g982) & (g983) & (!g1018)) + ((g127) & (g147) & (g982) & (g983) & (g1018)));
	assign g1020 = (((!g87) & (!g104) & (g979) & (g980) & (g1019)) + ((!g87) & (g104) & (g979) & (!g980) & (g1019)) + ((!g87) & (g104) & (g979) & (g980) & (!g1019)) + ((!g87) & (g104) & (g979) & (g980) & (g1019)) + ((g87) & (!g104) & (!g979) & (g980) & (g1019)) + ((g87) & (!g104) & (g979) & (!g980) & (!g1019)) + ((g87) & (!g104) & (g979) & (!g980) & (g1019)) + ((g87) & (!g104) & (g979) & (g980) & (!g1019)) + ((g87) & (!g104) & (g979) & (g980) & (g1019)) + ((g87) & (g104) & (!g979) & (!g980) & (g1019)) + ((g87) & (g104) & (!g979) & (g980) & (!g1019)) + ((g87) & (g104) & (!g979) & (g980) & (g1019)) + ((g87) & (g104) & (g979) & (!g980) & (!g1019)) + ((g87) & (g104) & (g979) & (!g980) & (g1019)) + ((g87) & (g104) & (g979) & (g980) & (!g1019)) + ((g87) & (g104) & (g979) & (g980) & (g1019)));
	assign g1021 = (((!g54) & (!g68) & (g976) & (g977) & (g1020)) + ((!g54) & (g68) & (g976) & (!g977) & (g1020)) + ((!g54) & (g68) & (g976) & (g977) & (!g1020)) + ((!g54) & (g68) & (g976) & (g977) & (g1020)) + ((g54) & (!g68) & (!g976) & (g977) & (g1020)) + ((g54) & (!g68) & (g976) & (!g977) & (!g1020)) + ((g54) & (!g68) & (g976) & (!g977) & (g1020)) + ((g54) & (!g68) & (g976) & (g977) & (!g1020)) + ((g54) & (!g68) & (g976) & (g977) & (g1020)) + ((g54) & (g68) & (!g976) & (!g977) & (g1020)) + ((g54) & (g68) & (!g976) & (g977) & (!g1020)) + ((g54) & (g68) & (!g976) & (g977) & (g1020)) + ((g54) & (g68) & (g976) & (!g977) & (!g1020)) + ((g54) & (g68) & (g976) & (!g977) & (g1020)) + ((g54) & (g68) & (g976) & (g977) & (!g1020)) + ((g54) & (g68) & (g976) & (g977) & (g1020)));
	assign g1022 = (((!g27) & (!g39) & (g973) & (g974) & (g1021)) + ((!g27) & (g39) & (g973) & (!g974) & (g1021)) + ((!g27) & (g39) & (g973) & (g974) & (!g1021)) + ((!g27) & (g39) & (g973) & (g974) & (g1021)) + ((g27) & (!g39) & (!g973) & (g974) & (g1021)) + ((g27) & (!g39) & (g973) & (!g974) & (!g1021)) + ((g27) & (!g39) & (g973) & (!g974) & (g1021)) + ((g27) & (!g39) & (g973) & (g974) & (!g1021)) + ((g27) & (!g39) & (g973) & (g974) & (g1021)) + ((g27) & (g39) & (!g973) & (!g974) & (g1021)) + ((g27) & (g39) & (!g973) & (g974) & (!g1021)) + ((g27) & (g39) & (!g973) & (g974) & (g1021)) + ((g27) & (g39) & (g973) & (!g974) & (!g1021)) + ((g27) & (g39) & (g973) & (!g974) & (g1021)) + ((g27) & (g39) & (g973) & (g974) & (!g1021)) + ((g27) & (g39) & (g973) & (g974) & (g1021)));
	assign g1023 = (((!g8) & (!g18) & (g970) & (g971) & (g1022)) + ((!g8) & (g18) & (g970) & (!g971) & (g1022)) + ((!g8) & (g18) & (g970) & (g971) & (!g1022)) + ((!g8) & (g18) & (g970) & (g971) & (g1022)) + ((g8) & (!g18) & (!g970) & (g971) & (g1022)) + ((g8) & (!g18) & (g970) & (!g971) & (!g1022)) + ((g8) & (!g18) & (g970) & (!g971) & (g1022)) + ((g8) & (!g18) & (g970) & (g971) & (!g1022)) + ((g8) & (!g18) & (g970) & (g971) & (g1022)) + ((g8) & (g18) & (!g970) & (!g971) & (g1022)) + ((g8) & (g18) & (!g970) & (g971) & (!g1022)) + ((g8) & (g18) & (!g970) & (g971) & (g1022)) + ((g8) & (g18) & (g970) & (!g971) & (!g1022)) + ((g8) & (g18) & (g970) & (!g971) & (g1022)) + ((g8) & (g18) & (g970) & (g971) & (!g1022)) + ((g8) & (g18) & (g970) & (g971) & (g1022)));
	assign g1024 = (((!g2) & (!g8) & (g919) & (g959)) + ((!g2) & (g8) & (!g919) & (g959)) + ((!g2) & (g8) & (g919) & (!g959)) + ((!g2) & (g8) & (g919) & (g959)) + ((g2) & (!g8) & (!g919) & (!g959)) + ((g2) & (!g8) & (!g919) & (g959)) + ((g2) & (!g8) & (g919) & (!g959)) + ((g2) & (g8) & (!g919) & (!g959)));
	assign g1025 = (((!g918) & (!g916) & (!g963) & (g1024)) + ((!g918) & (g916) & (!g963) & (g1024)) + ((!g918) & (g916) & (g963) & (g1024)) + ((g918) & (!g916) & (!g963) & (!g1024)) + ((g918) & (!g916) & (g963) & (!g1024)) + ((g918) & (!g916) & (g963) & (g1024)) + ((g918) & (g916) & (!g963) & (!g1024)) + ((g918) & (g916) & (g963) & (!g1024)));
	assign g1026 = (((!g4) & (!g2) & (!g968) & (!g1023) & (g1025)) + ((!g4) & (!g2) & (!g968) & (g1023) & (g1025)) + ((!g4) & (!g2) & (g968) & (!g1023) & (g1025)) + ((!g4) & (!g2) & (g968) & (g1023) & (!g1025)) + ((!g4) & (!g2) & (g968) & (g1023) & (g1025)) + ((!g4) & (g2) & (!g968) & (!g1023) & (g1025)) + ((!g4) & (g2) & (!g968) & (g1023) & (!g1025)) + ((!g4) & (g2) & (!g968) & (g1023) & (g1025)) + ((!g4) & (g2) & (g968) & (!g1023) & (!g1025)) + ((!g4) & (g2) & (g968) & (!g1023) & (g1025)) + ((!g4) & (g2) & (g968) & (g1023) & (!g1025)) + ((!g4) & (g2) & (g968) & (g1023) & (g1025)) + ((g4) & (!g2) & (g968) & (g1023) & (g1025)) + ((g4) & (g2) & (!g968) & (g1023) & (g1025)) + ((g4) & (g2) & (g968) & (!g1023) & (g1025)) + ((g4) & (g2) & (g968) & (g1023) & (g1025)));
	assign g1027 = (((!g4) & (!g960) & (g961)) + ((!g4) & (g960) & (!g961)) + ((!g4) & (g960) & (g961)) + ((g4) & (g960) & (g961)));
	assign g1028 = (((!g917) & (!g1027) & (!g916) & (!g963)) + ((!g917) & (!g1027) & (g916) & (!g963)) + ((!g917) & (!g1027) & (g916) & (g963)) + ((g917) & (g1027) & (!g916) & (!g963)) + ((g917) & (g1027) & (!g916) & (g963)) + ((g917) & (g1027) & (g916) & (!g963)) + ((g917) & (g1027) & (g916) & (g963)));
	assign g1029 = (((!g1) & (g917) & (!g1027) & (!g916) & (g963)) + ((!g1) & (g917) & (g1027) & (!g916) & (g963)) + ((g1) & (!g917) & (g1027) & (g916) & (!g963)) + ((g1) & (!g917) & (g1027) & (g916) & (g963)) + ((g1) & (g917) & (!g1027) & (!g916) & (!g963)) + ((g1) & (g917) & (!g1027) & (!g916) & (g963)) + ((g1) & (g917) & (!g1027) & (g916) & (!g963)) + ((g1) & (g917) & (!g1027) & (g916) & (g963)) + ((g1) & (g917) & (g1027) & (!g916) & (g963)));
	assign g1030 = (((!g1) & (!g967) & (!g1026) & (!g1028) & (!g1029)) + ((g1) & (!g967) & (!g1026) & (!g1028) & (!g1029)) + ((g1) & (!g967) & (!g1026) & (g1028) & (!g1029)) + ((g1) & (!g967) & (g1026) & (!g1028) & (!g1029)) + ((g1) & (!g967) & (g1026) & (g1028) & (!g1029)) + ((g1) & (g967) & (!g1026) & (!g1028) & (!g1029)) + ((g1) & (g967) & (!g1026) & (g1028) & (!g1029)));
	assign g1031 = (((!g851) & (!g964) & (g966) & (!g1030)) + ((!g851) & (g964) & (!g966) & (!g1030)) + ((!g851) & (g964) & (!g966) & (g1030)) + ((!g851) & (g964) & (g966) & (g1030)) + ((g851) & (!g964) & (!g966) & (!g1030)) + ((g851) & (g964) & (!g966) & (g1030)) + ((g851) & (g964) & (g966) & (!g1030)) + ((g851) & (g964) & (g966) & (g1030)));
	assign g1032 = (((!g916) & (g963)));
	assign g1033 = (((!g914) & (!ax62x) & (!ax63x) & (!g1032) & (!g965) & (g1030)) + ((!g914) & (!ax62x) & (!ax63x) & (!g1032) & (g965) & (!g1030)) + ((!g914) & (!ax62x) & (!ax63x) & (!g1032) & (g965) & (g1030)) + ((!g914) & (!ax62x) & (!ax63x) & (g1032) & (!g965) & (!g1030)) + ((!g914) & (!ax62x) & (ax63x) & (!g1032) & (!g965) & (!g1030)) + ((!g914) & (!ax62x) & (ax63x) & (g1032) & (!g965) & (g1030)) + ((!g914) & (!ax62x) & (ax63x) & (g1032) & (g965) & (!g1030)) + ((!g914) & (!ax62x) & (ax63x) & (g1032) & (g965) & (g1030)) + ((!g914) & (ax62x) & (!ax63x) & (g1032) & (!g965) & (!g1030)) + ((!g914) & (ax62x) & (!ax63x) & (g1032) & (g965) & (!g1030)) + ((!g914) & (ax62x) & (ax63x) & (!g1032) & (!g965) & (!g1030)) + ((!g914) & (ax62x) & (ax63x) & (!g1032) & (!g965) & (g1030)) + ((!g914) & (ax62x) & (ax63x) & (!g1032) & (g965) & (!g1030)) + ((!g914) & (ax62x) & (ax63x) & (!g1032) & (g965) & (g1030)) + ((!g914) & (ax62x) & (ax63x) & (g1032) & (!g965) & (g1030)) + ((!g914) & (ax62x) & (ax63x) & (g1032) & (g965) & (g1030)) + ((g914) & (!ax62x) & (!ax63x) & (!g1032) & (!g965) & (!g1030)) + ((g914) & (!ax62x) & (!ax63x) & (!g1032) & (!g965) & (g1030)) + ((g914) & (!ax62x) & (!ax63x) & (!g1032) & (g965) & (g1030)) + ((g914) & (!ax62x) & (!ax63x) & (g1032) & (g965) & (!g1030)) + ((g914) & (!ax62x) & (ax63x) & (!g1032) & (g965) & (!g1030)) + ((g914) & (!ax62x) & (ax63x) & (g1032) & (!g965) & (!g1030)) + ((g914) & (!ax62x) & (ax63x) & (g1032) & (!g965) & (g1030)) + ((g914) & (!ax62x) & (ax63x) & (g1032) & (g965) & (g1030)) + ((g914) & (ax62x) & (!ax63x) & (!g1032) & (!g965) & (!g1030)) + ((g914) & (ax62x) & (!ax63x) & (!g1032) & (g965) & (!g1030)) + ((g914) & (ax62x) & (ax63x) & (!g1032) & (!g965) & (g1030)) + ((g914) & (ax62x) & (ax63x) & (!g1032) & (g965) & (g1030)) + ((g914) & (ax62x) & (ax63x) & (g1032) & (!g965) & (!g1030)) + ((g914) & (ax62x) & (ax63x) & (g1032) & (!g965) & (g1030)) + ((g914) & (ax62x) & (ax63x) & (g1032) & (g965) & (!g1030)) + ((g914) & (ax62x) & (ax63x) & (g1032) & (g965) & (g1030)));
	assign g1034 = (((!ax62x) & (!g1032) & (!g965) & (g1030)) + ((!ax62x) & (!g1032) & (g965) & (!g1030)) + ((!ax62x) & (!g1032) & (g965) & (g1030)) + ((!ax62x) & (g1032) & (g965) & (!g1030)) + ((ax62x) & (!g1032) & (!g965) & (!g1030)) + ((ax62x) & (g1032) & (!g965) & (!g1030)) + ((ax62x) & (g1032) & (!g965) & (g1030)) + ((ax62x) & (g1032) & (g965) & (g1030)));
	assign g1035 = (((!ax58x) & (!ax59x)));
	assign g1036 = (((!g1032) & (!ax60x) & (!ax61x) & (!g1030) & (!g1035)) + ((!g1032) & (!ax60x) & (ax61x) & (g1030) & (!g1035)) + ((!g1032) & (ax60x) & (ax61x) & (g1030) & (!g1035)) + ((!g1032) & (ax60x) & (ax61x) & (g1030) & (g1035)) + ((g1032) & (!ax60x) & (!ax61x) & (!g1030) & (!g1035)) + ((g1032) & (!ax60x) & (!ax61x) & (!g1030) & (g1035)) + ((g1032) & (!ax60x) & (!ax61x) & (g1030) & (!g1035)) + ((g1032) & (!ax60x) & (ax61x) & (!g1030) & (!g1035)) + ((g1032) & (!ax60x) & (ax61x) & (g1030) & (!g1035)) + ((g1032) & (!ax60x) & (ax61x) & (g1030) & (g1035)) + ((g1032) & (ax60x) & (!ax61x) & (g1030) & (!g1035)) + ((g1032) & (ax60x) & (!ax61x) & (g1030) & (g1035)) + ((g1032) & (ax60x) & (ax61x) & (!g1030) & (!g1035)) + ((g1032) & (ax60x) & (ax61x) & (!g1030) & (g1035)) + ((g1032) & (ax60x) & (ax61x) & (g1030) & (!g1035)) + ((g1032) & (ax60x) & (ax61x) & (g1030) & (g1035)));
	assign g1037 = (((!g851) & (!g914) & (g1033) & (g1034) & (g1036)) + ((!g851) & (g914) & (g1033) & (!g1034) & (g1036)) + ((!g851) & (g914) & (g1033) & (g1034) & (!g1036)) + ((!g851) & (g914) & (g1033) & (g1034) & (g1036)) + ((g851) & (!g914) & (!g1033) & (g1034) & (g1036)) + ((g851) & (!g914) & (g1033) & (!g1034) & (!g1036)) + ((g851) & (!g914) & (g1033) & (!g1034) & (g1036)) + ((g851) & (!g914) & (g1033) & (g1034) & (!g1036)) + ((g851) & (!g914) & (g1033) & (g1034) & (g1036)) + ((g851) & (g914) & (!g1033) & (!g1034) & (g1036)) + ((g851) & (g914) & (!g1033) & (g1034) & (!g1036)) + ((g851) & (g914) & (!g1033) & (g1034) & (g1036)) + ((g851) & (g914) & (g1033) & (!g1034) & (!g1036)) + ((g851) & (g914) & (g1033) & (!g1034) & (g1036)) + ((g851) & (g914) & (g1033) & (g1034) & (!g1036)) + ((g851) & (g914) & (g1033) & (g1034) & (g1036)));
	assign g1038 = (((g1) & (!g967) & (g1026) & (g1029)) + ((g1) & (g967) & (!g1026) & (!g1029)) + ((g1) & (g967) & (!g1026) & (g1029)));
	assign g1039 = (((!g4) & (!g2) & (!g968) & (!g1023) & (!g1025) & (!g1030)) + ((!g4) & (!g2) & (!g968) & (!g1023) & (g1025) & (g1030)) + ((!g4) & (!g2) & (!g968) & (g1023) & (!g1025) & (!g1030)) + ((!g4) & (!g2) & (!g968) & (g1023) & (g1025) & (g1030)) + ((!g4) & (!g2) & (g968) & (!g1023) & (!g1025) & (!g1030)) + ((!g4) & (!g2) & (g968) & (!g1023) & (g1025) & (g1030)) + ((!g4) & (!g2) & (g968) & (g1023) & (g1025) & (!g1030)) + ((!g4) & (!g2) & (g968) & (g1023) & (g1025) & (g1030)) + ((!g4) & (g2) & (!g968) & (!g1023) & (!g1025) & (!g1030)) + ((!g4) & (g2) & (!g968) & (!g1023) & (g1025) & (g1030)) + ((!g4) & (g2) & (!g968) & (g1023) & (g1025) & (!g1030)) + ((!g4) & (g2) & (!g968) & (g1023) & (g1025) & (g1030)) + ((!g4) & (g2) & (g968) & (!g1023) & (g1025) & (!g1030)) + ((!g4) & (g2) & (g968) & (!g1023) & (g1025) & (g1030)) + ((!g4) & (g2) & (g968) & (g1023) & (g1025) & (!g1030)) + ((!g4) & (g2) & (g968) & (g1023) & (g1025) & (g1030)) + ((g4) & (!g2) & (!g968) & (!g1023) & (g1025) & (!g1030)) + ((g4) & (!g2) & (!g968) & (!g1023) & (g1025) & (g1030)) + ((g4) & (!g2) & (!g968) & (g1023) & (g1025) & (!g1030)) + ((g4) & (!g2) & (!g968) & (g1023) & (g1025) & (g1030)) + ((g4) & (!g2) & (g968) & (!g1023) & (g1025) & (!g1030)) + ((g4) & (!g2) & (g968) & (!g1023) & (g1025) & (g1030)) + ((g4) & (!g2) & (g968) & (g1023) & (!g1025) & (!g1030)) + ((g4) & (!g2) & (g968) & (g1023) & (g1025) & (g1030)) + ((g4) & (g2) & (!g968) & (!g1023) & (g1025) & (!g1030)) + ((g4) & (g2) & (!g968) & (!g1023) & (g1025) & (g1030)) + ((g4) & (g2) & (!g968) & (g1023) & (!g1025) & (!g1030)) + ((g4) & (g2) & (!g968) & (g1023) & (g1025) & (g1030)) + ((g4) & (g2) & (g968) & (!g1023) & (!g1025) & (!g1030)) + ((g4) & (g2) & (g968) & (!g1023) & (g1025) & (g1030)) + ((g4) & (g2) & (g968) & (g1023) & (!g1025) & (!g1030)) + ((g4) & (g2) & (g968) & (g1023) & (g1025) & (g1030)));
	assign g1040 = (((!g8) & (!g18) & (!g970) & (g971) & (g1022) & (!g1030)) + ((!g8) & (!g18) & (g970) & (!g971) & (!g1022) & (!g1030)) + ((!g8) & (!g18) & (g970) & (!g971) & (!g1022) & (g1030)) + ((!g8) & (!g18) & (g970) & (!g971) & (g1022) & (!g1030)) + ((!g8) & (!g18) & (g970) & (!g971) & (g1022) & (g1030)) + ((!g8) & (!g18) & (g970) & (g971) & (!g1022) & (!g1030)) + ((!g8) & (!g18) & (g970) & (g971) & (!g1022) & (g1030)) + ((!g8) & (!g18) & (g970) & (g971) & (g1022) & (g1030)) + ((!g8) & (g18) & (!g970) & (!g971) & (g1022) & (!g1030)) + ((!g8) & (g18) & (!g970) & (g971) & (!g1022) & (!g1030)) + ((!g8) & (g18) & (!g970) & (g971) & (g1022) & (!g1030)) + ((!g8) & (g18) & (g970) & (!g971) & (!g1022) & (!g1030)) + ((!g8) & (g18) & (g970) & (!g971) & (!g1022) & (g1030)) + ((!g8) & (g18) & (g970) & (!g971) & (g1022) & (g1030)) + ((!g8) & (g18) & (g970) & (g971) & (!g1022) & (g1030)) + ((!g8) & (g18) & (g970) & (g971) & (g1022) & (g1030)) + ((g8) & (!g18) & (!g970) & (!g971) & (!g1022) & (!g1030)) + ((g8) & (!g18) & (!g970) & (!g971) & (g1022) & (!g1030)) + ((g8) & (!g18) & (!g970) & (g971) & (!g1022) & (!g1030)) + ((g8) & (!g18) & (g970) & (!g971) & (!g1022) & (g1030)) + ((g8) & (!g18) & (g970) & (!g971) & (g1022) & (g1030)) + ((g8) & (!g18) & (g970) & (g971) & (!g1022) & (g1030)) + ((g8) & (!g18) & (g970) & (g971) & (g1022) & (!g1030)) + ((g8) & (!g18) & (g970) & (g971) & (g1022) & (g1030)) + ((g8) & (g18) & (!g970) & (!g971) & (!g1022) & (!g1030)) + ((g8) & (g18) & (g970) & (!g971) & (!g1022) & (g1030)) + ((g8) & (g18) & (g970) & (!g971) & (g1022) & (!g1030)) + ((g8) & (g18) & (g970) & (!g971) & (g1022) & (g1030)) + ((g8) & (g18) & (g970) & (g971) & (!g1022) & (!g1030)) + ((g8) & (g18) & (g970) & (g971) & (!g1022) & (g1030)) + ((g8) & (g18) & (g970) & (g971) & (g1022) & (!g1030)) + ((g8) & (g18) & (g970) & (g971) & (g1022) & (g1030)));
	assign g1041 = (((!g18) & (!g971) & (g1022) & (!g1030)) + ((!g18) & (g971) & (!g1022) & (!g1030)) + ((!g18) & (g971) & (!g1022) & (g1030)) + ((!g18) & (g971) & (g1022) & (g1030)) + ((g18) & (!g971) & (!g1022) & (!g1030)) + ((g18) & (g971) & (!g1022) & (g1030)) + ((g18) & (g971) & (g1022) & (!g1030)) + ((g18) & (g971) & (g1022) & (g1030)));
	assign g1042 = (((!g27) & (!g39) & (!g973) & (g974) & (g1021) & (!g1030)) + ((!g27) & (!g39) & (g973) & (!g974) & (!g1021) & (!g1030)) + ((!g27) & (!g39) & (g973) & (!g974) & (!g1021) & (g1030)) + ((!g27) & (!g39) & (g973) & (!g974) & (g1021) & (!g1030)) + ((!g27) & (!g39) & (g973) & (!g974) & (g1021) & (g1030)) + ((!g27) & (!g39) & (g973) & (g974) & (!g1021) & (!g1030)) + ((!g27) & (!g39) & (g973) & (g974) & (!g1021) & (g1030)) + ((!g27) & (!g39) & (g973) & (g974) & (g1021) & (g1030)) + ((!g27) & (g39) & (!g973) & (!g974) & (g1021) & (!g1030)) + ((!g27) & (g39) & (!g973) & (g974) & (!g1021) & (!g1030)) + ((!g27) & (g39) & (!g973) & (g974) & (g1021) & (!g1030)) + ((!g27) & (g39) & (g973) & (!g974) & (!g1021) & (!g1030)) + ((!g27) & (g39) & (g973) & (!g974) & (!g1021) & (g1030)) + ((!g27) & (g39) & (g973) & (!g974) & (g1021) & (g1030)) + ((!g27) & (g39) & (g973) & (g974) & (!g1021) & (g1030)) + ((!g27) & (g39) & (g973) & (g974) & (g1021) & (g1030)) + ((g27) & (!g39) & (!g973) & (!g974) & (!g1021) & (!g1030)) + ((g27) & (!g39) & (!g973) & (!g974) & (g1021) & (!g1030)) + ((g27) & (!g39) & (!g973) & (g974) & (!g1021) & (!g1030)) + ((g27) & (!g39) & (g973) & (!g974) & (!g1021) & (g1030)) + ((g27) & (!g39) & (g973) & (!g974) & (g1021) & (g1030)) + ((g27) & (!g39) & (g973) & (g974) & (!g1021) & (g1030)) + ((g27) & (!g39) & (g973) & (g974) & (g1021) & (!g1030)) + ((g27) & (!g39) & (g973) & (g974) & (g1021) & (g1030)) + ((g27) & (g39) & (!g973) & (!g974) & (!g1021) & (!g1030)) + ((g27) & (g39) & (g973) & (!g974) & (!g1021) & (g1030)) + ((g27) & (g39) & (g973) & (!g974) & (g1021) & (!g1030)) + ((g27) & (g39) & (g973) & (!g974) & (g1021) & (g1030)) + ((g27) & (g39) & (g973) & (g974) & (!g1021) & (!g1030)) + ((g27) & (g39) & (g973) & (g974) & (!g1021) & (g1030)) + ((g27) & (g39) & (g973) & (g974) & (g1021) & (!g1030)) + ((g27) & (g39) & (g973) & (g974) & (g1021) & (g1030)));
	assign g1043 = (((!g39) & (!g974) & (g1021) & (!g1030)) + ((!g39) & (g974) & (!g1021) & (!g1030)) + ((!g39) & (g974) & (!g1021) & (g1030)) + ((!g39) & (g974) & (g1021) & (g1030)) + ((g39) & (!g974) & (!g1021) & (!g1030)) + ((g39) & (g974) & (!g1021) & (g1030)) + ((g39) & (g974) & (g1021) & (!g1030)) + ((g39) & (g974) & (g1021) & (g1030)));
	assign g1044 = (((!g54) & (!g68) & (!g976) & (g977) & (g1020) & (!g1030)) + ((!g54) & (!g68) & (g976) & (!g977) & (!g1020) & (!g1030)) + ((!g54) & (!g68) & (g976) & (!g977) & (!g1020) & (g1030)) + ((!g54) & (!g68) & (g976) & (!g977) & (g1020) & (!g1030)) + ((!g54) & (!g68) & (g976) & (!g977) & (g1020) & (g1030)) + ((!g54) & (!g68) & (g976) & (g977) & (!g1020) & (!g1030)) + ((!g54) & (!g68) & (g976) & (g977) & (!g1020) & (g1030)) + ((!g54) & (!g68) & (g976) & (g977) & (g1020) & (g1030)) + ((!g54) & (g68) & (!g976) & (!g977) & (g1020) & (!g1030)) + ((!g54) & (g68) & (!g976) & (g977) & (!g1020) & (!g1030)) + ((!g54) & (g68) & (!g976) & (g977) & (g1020) & (!g1030)) + ((!g54) & (g68) & (g976) & (!g977) & (!g1020) & (!g1030)) + ((!g54) & (g68) & (g976) & (!g977) & (!g1020) & (g1030)) + ((!g54) & (g68) & (g976) & (!g977) & (g1020) & (g1030)) + ((!g54) & (g68) & (g976) & (g977) & (!g1020) & (g1030)) + ((!g54) & (g68) & (g976) & (g977) & (g1020) & (g1030)) + ((g54) & (!g68) & (!g976) & (!g977) & (!g1020) & (!g1030)) + ((g54) & (!g68) & (!g976) & (!g977) & (g1020) & (!g1030)) + ((g54) & (!g68) & (!g976) & (g977) & (!g1020) & (!g1030)) + ((g54) & (!g68) & (g976) & (!g977) & (!g1020) & (g1030)) + ((g54) & (!g68) & (g976) & (!g977) & (g1020) & (g1030)) + ((g54) & (!g68) & (g976) & (g977) & (!g1020) & (g1030)) + ((g54) & (!g68) & (g976) & (g977) & (g1020) & (!g1030)) + ((g54) & (!g68) & (g976) & (g977) & (g1020) & (g1030)) + ((g54) & (g68) & (!g976) & (!g977) & (!g1020) & (!g1030)) + ((g54) & (g68) & (g976) & (!g977) & (!g1020) & (g1030)) + ((g54) & (g68) & (g976) & (!g977) & (g1020) & (!g1030)) + ((g54) & (g68) & (g976) & (!g977) & (g1020) & (g1030)) + ((g54) & (g68) & (g976) & (g977) & (!g1020) & (!g1030)) + ((g54) & (g68) & (g976) & (g977) & (!g1020) & (g1030)) + ((g54) & (g68) & (g976) & (g977) & (g1020) & (!g1030)) + ((g54) & (g68) & (g976) & (g977) & (g1020) & (g1030)));
	assign g1045 = (((!g68) & (!g977) & (g1020) & (!g1030)) + ((!g68) & (g977) & (!g1020) & (!g1030)) + ((!g68) & (g977) & (!g1020) & (g1030)) + ((!g68) & (g977) & (g1020) & (g1030)) + ((g68) & (!g977) & (!g1020) & (!g1030)) + ((g68) & (g977) & (!g1020) & (g1030)) + ((g68) & (g977) & (g1020) & (!g1030)) + ((g68) & (g977) & (g1020) & (g1030)));
	assign g1046 = (((!g87) & (!g104) & (!g979) & (g980) & (g1019) & (!g1030)) + ((!g87) & (!g104) & (g979) & (!g980) & (!g1019) & (!g1030)) + ((!g87) & (!g104) & (g979) & (!g980) & (!g1019) & (g1030)) + ((!g87) & (!g104) & (g979) & (!g980) & (g1019) & (!g1030)) + ((!g87) & (!g104) & (g979) & (!g980) & (g1019) & (g1030)) + ((!g87) & (!g104) & (g979) & (g980) & (!g1019) & (!g1030)) + ((!g87) & (!g104) & (g979) & (g980) & (!g1019) & (g1030)) + ((!g87) & (!g104) & (g979) & (g980) & (g1019) & (g1030)) + ((!g87) & (g104) & (!g979) & (!g980) & (g1019) & (!g1030)) + ((!g87) & (g104) & (!g979) & (g980) & (!g1019) & (!g1030)) + ((!g87) & (g104) & (!g979) & (g980) & (g1019) & (!g1030)) + ((!g87) & (g104) & (g979) & (!g980) & (!g1019) & (!g1030)) + ((!g87) & (g104) & (g979) & (!g980) & (!g1019) & (g1030)) + ((!g87) & (g104) & (g979) & (!g980) & (g1019) & (g1030)) + ((!g87) & (g104) & (g979) & (g980) & (!g1019) & (g1030)) + ((!g87) & (g104) & (g979) & (g980) & (g1019) & (g1030)) + ((g87) & (!g104) & (!g979) & (!g980) & (!g1019) & (!g1030)) + ((g87) & (!g104) & (!g979) & (!g980) & (g1019) & (!g1030)) + ((g87) & (!g104) & (!g979) & (g980) & (!g1019) & (!g1030)) + ((g87) & (!g104) & (g979) & (!g980) & (!g1019) & (g1030)) + ((g87) & (!g104) & (g979) & (!g980) & (g1019) & (g1030)) + ((g87) & (!g104) & (g979) & (g980) & (!g1019) & (g1030)) + ((g87) & (!g104) & (g979) & (g980) & (g1019) & (!g1030)) + ((g87) & (!g104) & (g979) & (g980) & (g1019) & (g1030)) + ((g87) & (g104) & (!g979) & (!g980) & (!g1019) & (!g1030)) + ((g87) & (g104) & (g979) & (!g980) & (!g1019) & (g1030)) + ((g87) & (g104) & (g979) & (!g980) & (g1019) & (!g1030)) + ((g87) & (g104) & (g979) & (!g980) & (g1019) & (g1030)) + ((g87) & (g104) & (g979) & (g980) & (!g1019) & (!g1030)) + ((g87) & (g104) & (g979) & (g980) & (!g1019) & (g1030)) + ((g87) & (g104) & (g979) & (g980) & (g1019) & (!g1030)) + ((g87) & (g104) & (g979) & (g980) & (g1019) & (g1030)));
	assign g1047 = (((!g104) & (!g980) & (g1019) & (!g1030)) + ((!g104) & (g980) & (!g1019) & (!g1030)) + ((!g104) & (g980) & (!g1019) & (g1030)) + ((!g104) & (g980) & (g1019) & (g1030)) + ((g104) & (!g980) & (!g1019) & (!g1030)) + ((g104) & (g980) & (!g1019) & (g1030)) + ((g104) & (g980) & (g1019) & (!g1030)) + ((g104) & (g980) & (g1019) & (g1030)));
	assign g1048 = (((!g127) & (!g147) & (!g982) & (g983) & (g1018) & (!g1030)) + ((!g127) & (!g147) & (g982) & (!g983) & (!g1018) & (!g1030)) + ((!g127) & (!g147) & (g982) & (!g983) & (!g1018) & (g1030)) + ((!g127) & (!g147) & (g982) & (!g983) & (g1018) & (!g1030)) + ((!g127) & (!g147) & (g982) & (!g983) & (g1018) & (g1030)) + ((!g127) & (!g147) & (g982) & (g983) & (!g1018) & (!g1030)) + ((!g127) & (!g147) & (g982) & (g983) & (!g1018) & (g1030)) + ((!g127) & (!g147) & (g982) & (g983) & (g1018) & (g1030)) + ((!g127) & (g147) & (!g982) & (!g983) & (g1018) & (!g1030)) + ((!g127) & (g147) & (!g982) & (g983) & (!g1018) & (!g1030)) + ((!g127) & (g147) & (!g982) & (g983) & (g1018) & (!g1030)) + ((!g127) & (g147) & (g982) & (!g983) & (!g1018) & (!g1030)) + ((!g127) & (g147) & (g982) & (!g983) & (!g1018) & (g1030)) + ((!g127) & (g147) & (g982) & (!g983) & (g1018) & (g1030)) + ((!g127) & (g147) & (g982) & (g983) & (!g1018) & (g1030)) + ((!g127) & (g147) & (g982) & (g983) & (g1018) & (g1030)) + ((g127) & (!g147) & (!g982) & (!g983) & (!g1018) & (!g1030)) + ((g127) & (!g147) & (!g982) & (!g983) & (g1018) & (!g1030)) + ((g127) & (!g147) & (!g982) & (g983) & (!g1018) & (!g1030)) + ((g127) & (!g147) & (g982) & (!g983) & (!g1018) & (g1030)) + ((g127) & (!g147) & (g982) & (!g983) & (g1018) & (g1030)) + ((g127) & (!g147) & (g982) & (g983) & (!g1018) & (g1030)) + ((g127) & (!g147) & (g982) & (g983) & (g1018) & (!g1030)) + ((g127) & (!g147) & (g982) & (g983) & (g1018) & (g1030)) + ((g127) & (g147) & (!g982) & (!g983) & (!g1018) & (!g1030)) + ((g127) & (g147) & (g982) & (!g983) & (!g1018) & (g1030)) + ((g127) & (g147) & (g982) & (!g983) & (g1018) & (!g1030)) + ((g127) & (g147) & (g982) & (!g983) & (g1018) & (g1030)) + ((g127) & (g147) & (g982) & (g983) & (!g1018) & (!g1030)) + ((g127) & (g147) & (g982) & (g983) & (!g1018) & (g1030)) + ((g127) & (g147) & (g982) & (g983) & (g1018) & (!g1030)) + ((g127) & (g147) & (g982) & (g983) & (g1018) & (g1030)));
	assign g1049 = (((!g147) & (!g983) & (g1018) & (!g1030)) + ((!g147) & (g983) & (!g1018) & (!g1030)) + ((!g147) & (g983) & (!g1018) & (g1030)) + ((!g147) & (g983) & (g1018) & (g1030)) + ((g147) & (!g983) & (!g1018) & (!g1030)) + ((g147) & (g983) & (!g1018) & (g1030)) + ((g147) & (g983) & (g1018) & (!g1030)) + ((g147) & (g983) & (g1018) & (g1030)));
	assign g1050 = (((!g174) & (!g198) & (!g985) & (g986) & (g1017) & (!g1030)) + ((!g174) & (!g198) & (g985) & (!g986) & (!g1017) & (!g1030)) + ((!g174) & (!g198) & (g985) & (!g986) & (!g1017) & (g1030)) + ((!g174) & (!g198) & (g985) & (!g986) & (g1017) & (!g1030)) + ((!g174) & (!g198) & (g985) & (!g986) & (g1017) & (g1030)) + ((!g174) & (!g198) & (g985) & (g986) & (!g1017) & (!g1030)) + ((!g174) & (!g198) & (g985) & (g986) & (!g1017) & (g1030)) + ((!g174) & (!g198) & (g985) & (g986) & (g1017) & (g1030)) + ((!g174) & (g198) & (!g985) & (!g986) & (g1017) & (!g1030)) + ((!g174) & (g198) & (!g985) & (g986) & (!g1017) & (!g1030)) + ((!g174) & (g198) & (!g985) & (g986) & (g1017) & (!g1030)) + ((!g174) & (g198) & (g985) & (!g986) & (!g1017) & (!g1030)) + ((!g174) & (g198) & (g985) & (!g986) & (!g1017) & (g1030)) + ((!g174) & (g198) & (g985) & (!g986) & (g1017) & (g1030)) + ((!g174) & (g198) & (g985) & (g986) & (!g1017) & (g1030)) + ((!g174) & (g198) & (g985) & (g986) & (g1017) & (g1030)) + ((g174) & (!g198) & (!g985) & (!g986) & (!g1017) & (!g1030)) + ((g174) & (!g198) & (!g985) & (!g986) & (g1017) & (!g1030)) + ((g174) & (!g198) & (!g985) & (g986) & (!g1017) & (!g1030)) + ((g174) & (!g198) & (g985) & (!g986) & (!g1017) & (g1030)) + ((g174) & (!g198) & (g985) & (!g986) & (g1017) & (g1030)) + ((g174) & (!g198) & (g985) & (g986) & (!g1017) & (g1030)) + ((g174) & (!g198) & (g985) & (g986) & (g1017) & (!g1030)) + ((g174) & (!g198) & (g985) & (g986) & (g1017) & (g1030)) + ((g174) & (g198) & (!g985) & (!g986) & (!g1017) & (!g1030)) + ((g174) & (g198) & (g985) & (!g986) & (!g1017) & (g1030)) + ((g174) & (g198) & (g985) & (!g986) & (g1017) & (!g1030)) + ((g174) & (g198) & (g985) & (!g986) & (g1017) & (g1030)) + ((g174) & (g198) & (g985) & (g986) & (!g1017) & (!g1030)) + ((g174) & (g198) & (g985) & (g986) & (!g1017) & (g1030)) + ((g174) & (g198) & (g985) & (g986) & (g1017) & (!g1030)) + ((g174) & (g198) & (g985) & (g986) & (g1017) & (g1030)));
	assign g1051 = (((!g198) & (!g986) & (g1017) & (!g1030)) + ((!g198) & (g986) & (!g1017) & (!g1030)) + ((!g198) & (g986) & (!g1017) & (g1030)) + ((!g198) & (g986) & (g1017) & (g1030)) + ((g198) & (!g986) & (!g1017) & (!g1030)) + ((g198) & (g986) & (!g1017) & (g1030)) + ((g198) & (g986) & (g1017) & (!g1030)) + ((g198) & (g986) & (g1017) & (g1030)));
	assign g1052 = (((!g229) & (!g255) & (!g988) & (g989) & (g1016) & (!g1030)) + ((!g229) & (!g255) & (g988) & (!g989) & (!g1016) & (!g1030)) + ((!g229) & (!g255) & (g988) & (!g989) & (!g1016) & (g1030)) + ((!g229) & (!g255) & (g988) & (!g989) & (g1016) & (!g1030)) + ((!g229) & (!g255) & (g988) & (!g989) & (g1016) & (g1030)) + ((!g229) & (!g255) & (g988) & (g989) & (!g1016) & (!g1030)) + ((!g229) & (!g255) & (g988) & (g989) & (!g1016) & (g1030)) + ((!g229) & (!g255) & (g988) & (g989) & (g1016) & (g1030)) + ((!g229) & (g255) & (!g988) & (!g989) & (g1016) & (!g1030)) + ((!g229) & (g255) & (!g988) & (g989) & (!g1016) & (!g1030)) + ((!g229) & (g255) & (!g988) & (g989) & (g1016) & (!g1030)) + ((!g229) & (g255) & (g988) & (!g989) & (!g1016) & (!g1030)) + ((!g229) & (g255) & (g988) & (!g989) & (!g1016) & (g1030)) + ((!g229) & (g255) & (g988) & (!g989) & (g1016) & (g1030)) + ((!g229) & (g255) & (g988) & (g989) & (!g1016) & (g1030)) + ((!g229) & (g255) & (g988) & (g989) & (g1016) & (g1030)) + ((g229) & (!g255) & (!g988) & (!g989) & (!g1016) & (!g1030)) + ((g229) & (!g255) & (!g988) & (!g989) & (g1016) & (!g1030)) + ((g229) & (!g255) & (!g988) & (g989) & (!g1016) & (!g1030)) + ((g229) & (!g255) & (g988) & (!g989) & (!g1016) & (g1030)) + ((g229) & (!g255) & (g988) & (!g989) & (g1016) & (g1030)) + ((g229) & (!g255) & (g988) & (g989) & (!g1016) & (g1030)) + ((g229) & (!g255) & (g988) & (g989) & (g1016) & (!g1030)) + ((g229) & (!g255) & (g988) & (g989) & (g1016) & (g1030)) + ((g229) & (g255) & (!g988) & (!g989) & (!g1016) & (!g1030)) + ((g229) & (g255) & (g988) & (!g989) & (!g1016) & (g1030)) + ((g229) & (g255) & (g988) & (!g989) & (g1016) & (!g1030)) + ((g229) & (g255) & (g988) & (!g989) & (g1016) & (g1030)) + ((g229) & (g255) & (g988) & (g989) & (!g1016) & (!g1030)) + ((g229) & (g255) & (g988) & (g989) & (!g1016) & (g1030)) + ((g229) & (g255) & (g988) & (g989) & (g1016) & (!g1030)) + ((g229) & (g255) & (g988) & (g989) & (g1016) & (g1030)));
	assign g1053 = (((!g255) & (!g989) & (g1016) & (!g1030)) + ((!g255) & (g989) & (!g1016) & (!g1030)) + ((!g255) & (g989) & (!g1016) & (g1030)) + ((!g255) & (g989) & (g1016) & (g1030)) + ((g255) & (!g989) & (!g1016) & (!g1030)) + ((g255) & (g989) & (!g1016) & (g1030)) + ((g255) & (g989) & (g1016) & (!g1030)) + ((g255) & (g989) & (g1016) & (g1030)));
	assign g1054 = (((!g290) & (!g319) & (!g991) & (g992) & (g1015) & (!g1030)) + ((!g290) & (!g319) & (g991) & (!g992) & (!g1015) & (!g1030)) + ((!g290) & (!g319) & (g991) & (!g992) & (!g1015) & (g1030)) + ((!g290) & (!g319) & (g991) & (!g992) & (g1015) & (!g1030)) + ((!g290) & (!g319) & (g991) & (!g992) & (g1015) & (g1030)) + ((!g290) & (!g319) & (g991) & (g992) & (!g1015) & (!g1030)) + ((!g290) & (!g319) & (g991) & (g992) & (!g1015) & (g1030)) + ((!g290) & (!g319) & (g991) & (g992) & (g1015) & (g1030)) + ((!g290) & (g319) & (!g991) & (!g992) & (g1015) & (!g1030)) + ((!g290) & (g319) & (!g991) & (g992) & (!g1015) & (!g1030)) + ((!g290) & (g319) & (!g991) & (g992) & (g1015) & (!g1030)) + ((!g290) & (g319) & (g991) & (!g992) & (!g1015) & (!g1030)) + ((!g290) & (g319) & (g991) & (!g992) & (!g1015) & (g1030)) + ((!g290) & (g319) & (g991) & (!g992) & (g1015) & (g1030)) + ((!g290) & (g319) & (g991) & (g992) & (!g1015) & (g1030)) + ((!g290) & (g319) & (g991) & (g992) & (g1015) & (g1030)) + ((g290) & (!g319) & (!g991) & (!g992) & (!g1015) & (!g1030)) + ((g290) & (!g319) & (!g991) & (!g992) & (g1015) & (!g1030)) + ((g290) & (!g319) & (!g991) & (g992) & (!g1015) & (!g1030)) + ((g290) & (!g319) & (g991) & (!g992) & (!g1015) & (g1030)) + ((g290) & (!g319) & (g991) & (!g992) & (g1015) & (g1030)) + ((g290) & (!g319) & (g991) & (g992) & (!g1015) & (g1030)) + ((g290) & (!g319) & (g991) & (g992) & (g1015) & (!g1030)) + ((g290) & (!g319) & (g991) & (g992) & (g1015) & (g1030)) + ((g290) & (g319) & (!g991) & (!g992) & (!g1015) & (!g1030)) + ((g290) & (g319) & (g991) & (!g992) & (!g1015) & (g1030)) + ((g290) & (g319) & (g991) & (!g992) & (g1015) & (!g1030)) + ((g290) & (g319) & (g991) & (!g992) & (g1015) & (g1030)) + ((g290) & (g319) & (g991) & (g992) & (!g1015) & (!g1030)) + ((g290) & (g319) & (g991) & (g992) & (!g1015) & (g1030)) + ((g290) & (g319) & (g991) & (g992) & (g1015) & (!g1030)) + ((g290) & (g319) & (g991) & (g992) & (g1015) & (g1030)));
	assign g1055 = (((!g319) & (!g992) & (g1015) & (!g1030)) + ((!g319) & (g992) & (!g1015) & (!g1030)) + ((!g319) & (g992) & (!g1015) & (g1030)) + ((!g319) & (g992) & (g1015) & (g1030)) + ((g319) & (!g992) & (!g1015) & (!g1030)) + ((g319) & (g992) & (!g1015) & (g1030)) + ((g319) & (g992) & (g1015) & (!g1030)) + ((g319) & (g992) & (g1015) & (g1030)));
	assign g1056 = (((!g358) & (!g390) & (!g994) & (g995) & (g1014) & (!g1030)) + ((!g358) & (!g390) & (g994) & (!g995) & (!g1014) & (!g1030)) + ((!g358) & (!g390) & (g994) & (!g995) & (!g1014) & (g1030)) + ((!g358) & (!g390) & (g994) & (!g995) & (g1014) & (!g1030)) + ((!g358) & (!g390) & (g994) & (!g995) & (g1014) & (g1030)) + ((!g358) & (!g390) & (g994) & (g995) & (!g1014) & (!g1030)) + ((!g358) & (!g390) & (g994) & (g995) & (!g1014) & (g1030)) + ((!g358) & (!g390) & (g994) & (g995) & (g1014) & (g1030)) + ((!g358) & (g390) & (!g994) & (!g995) & (g1014) & (!g1030)) + ((!g358) & (g390) & (!g994) & (g995) & (!g1014) & (!g1030)) + ((!g358) & (g390) & (!g994) & (g995) & (g1014) & (!g1030)) + ((!g358) & (g390) & (g994) & (!g995) & (!g1014) & (!g1030)) + ((!g358) & (g390) & (g994) & (!g995) & (!g1014) & (g1030)) + ((!g358) & (g390) & (g994) & (!g995) & (g1014) & (g1030)) + ((!g358) & (g390) & (g994) & (g995) & (!g1014) & (g1030)) + ((!g358) & (g390) & (g994) & (g995) & (g1014) & (g1030)) + ((g358) & (!g390) & (!g994) & (!g995) & (!g1014) & (!g1030)) + ((g358) & (!g390) & (!g994) & (!g995) & (g1014) & (!g1030)) + ((g358) & (!g390) & (!g994) & (g995) & (!g1014) & (!g1030)) + ((g358) & (!g390) & (g994) & (!g995) & (!g1014) & (g1030)) + ((g358) & (!g390) & (g994) & (!g995) & (g1014) & (g1030)) + ((g358) & (!g390) & (g994) & (g995) & (!g1014) & (g1030)) + ((g358) & (!g390) & (g994) & (g995) & (g1014) & (!g1030)) + ((g358) & (!g390) & (g994) & (g995) & (g1014) & (g1030)) + ((g358) & (g390) & (!g994) & (!g995) & (!g1014) & (!g1030)) + ((g358) & (g390) & (g994) & (!g995) & (!g1014) & (g1030)) + ((g358) & (g390) & (g994) & (!g995) & (g1014) & (!g1030)) + ((g358) & (g390) & (g994) & (!g995) & (g1014) & (g1030)) + ((g358) & (g390) & (g994) & (g995) & (!g1014) & (!g1030)) + ((g358) & (g390) & (g994) & (g995) & (!g1014) & (g1030)) + ((g358) & (g390) & (g994) & (g995) & (g1014) & (!g1030)) + ((g358) & (g390) & (g994) & (g995) & (g1014) & (g1030)));
	assign g1057 = (((!g390) & (!g995) & (g1014) & (!g1030)) + ((!g390) & (g995) & (!g1014) & (!g1030)) + ((!g390) & (g995) & (!g1014) & (g1030)) + ((!g390) & (g995) & (g1014) & (g1030)) + ((g390) & (!g995) & (!g1014) & (!g1030)) + ((g390) & (g995) & (!g1014) & (g1030)) + ((g390) & (g995) & (g1014) & (!g1030)) + ((g390) & (g995) & (g1014) & (g1030)));
	assign g1058 = (((!g433) & (!g468) & (!g997) & (g998) & (g1013) & (!g1030)) + ((!g433) & (!g468) & (g997) & (!g998) & (!g1013) & (!g1030)) + ((!g433) & (!g468) & (g997) & (!g998) & (!g1013) & (g1030)) + ((!g433) & (!g468) & (g997) & (!g998) & (g1013) & (!g1030)) + ((!g433) & (!g468) & (g997) & (!g998) & (g1013) & (g1030)) + ((!g433) & (!g468) & (g997) & (g998) & (!g1013) & (!g1030)) + ((!g433) & (!g468) & (g997) & (g998) & (!g1013) & (g1030)) + ((!g433) & (!g468) & (g997) & (g998) & (g1013) & (g1030)) + ((!g433) & (g468) & (!g997) & (!g998) & (g1013) & (!g1030)) + ((!g433) & (g468) & (!g997) & (g998) & (!g1013) & (!g1030)) + ((!g433) & (g468) & (!g997) & (g998) & (g1013) & (!g1030)) + ((!g433) & (g468) & (g997) & (!g998) & (!g1013) & (!g1030)) + ((!g433) & (g468) & (g997) & (!g998) & (!g1013) & (g1030)) + ((!g433) & (g468) & (g997) & (!g998) & (g1013) & (g1030)) + ((!g433) & (g468) & (g997) & (g998) & (!g1013) & (g1030)) + ((!g433) & (g468) & (g997) & (g998) & (g1013) & (g1030)) + ((g433) & (!g468) & (!g997) & (!g998) & (!g1013) & (!g1030)) + ((g433) & (!g468) & (!g997) & (!g998) & (g1013) & (!g1030)) + ((g433) & (!g468) & (!g997) & (g998) & (!g1013) & (!g1030)) + ((g433) & (!g468) & (g997) & (!g998) & (!g1013) & (g1030)) + ((g433) & (!g468) & (g997) & (!g998) & (g1013) & (g1030)) + ((g433) & (!g468) & (g997) & (g998) & (!g1013) & (g1030)) + ((g433) & (!g468) & (g997) & (g998) & (g1013) & (!g1030)) + ((g433) & (!g468) & (g997) & (g998) & (g1013) & (g1030)) + ((g433) & (g468) & (!g997) & (!g998) & (!g1013) & (!g1030)) + ((g433) & (g468) & (g997) & (!g998) & (!g1013) & (g1030)) + ((g433) & (g468) & (g997) & (!g998) & (g1013) & (!g1030)) + ((g433) & (g468) & (g997) & (!g998) & (g1013) & (g1030)) + ((g433) & (g468) & (g997) & (g998) & (!g1013) & (!g1030)) + ((g433) & (g468) & (g997) & (g998) & (!g1013) & (g1030)) + ((g433) & (g468) & (g997) & (g998) & (g1013) & (!g1030)) + ((g433) & (g468) & (g997) & (g998) & (g1013) & (g1030)));
	assign g1059 = (((!g468) & (!g998) & (g1013) & (!g1030)) + ((!g468) & (g998) & (!g1013) & (!g1030)) + ((!g468) & (g998) & (!g1013) & (g1030)) + ((!g468) & (g998) & (g1013) & (g1030)) + ((g468) & (!g998) & (!g1013) & (!g1030)) + ((g468) & (g998) & (!g1013) & (g1030)) + ((g468) & (g998) & (g1013) & (!g1030)) + ((g468) & (g998) & (g1013) & (g1030)));
	assign g1060 = (((!g515) & (!g553) & (!g1000) & (g1001) & (g1012) & (!g1030)) + ((!g515) & (!g553) & (g1000) & (!g1001) & (!g1012) & (!g1030)) + ((!g515) & (!g553) & (g1000) & (!g1001) & (!g1012) & (g1030)) + ((!g515) & (!g553) & (g1000) & (!g1001) & (g1012) & (!g1030)) + ((!g515) & (!g553) & (g1000) & (!g1001) & (g1012) & (g1030)) + ((!g515) & (!g553) & (g1000) & (g1001) & (!g1012) & (!g1030)) + ((!g515) & (!g553) & (g1000) & (g1001) & (!g1012) & (g1030)) + ((!g515) & (!g553) & (g1000) & (g1001) & (g1012) & (g1030)) + ((!g515) & (g553) & (!g1000) & (!g1001) & (g1012) & (!g1030)) + ((!g515) & (g553) & (!g1000) & (g1001) & (!g1012) & (!g1030)) + ((!g515) & (g553) & (!g1000) & (g1001) & (g1012) & (!g1030)) + ((!g515) & (g553) & (g1000) & (!g1001) & (!g1012) & (!g1030)) + ((!g515) & (g553) & (g1000) & (!g1001) & (!g1012) & (g1030)) + ((!g515) & (g553) & (g1000) & (!g1001) & (g1012) & (g1030)) + ((!g515) & (g553) & (g1000) & (g1001) & (!g1012) & (g1030)) + ((!g515) & (g553) & (g1000) & (g1001) & (g1012) & (g1030)) + ((g515) & (!g553) & (!g1000) & (!g1001) & (!g1012) & (!g1030)) + ((g515) & (!g553) & (!g1000) & (!g1001) & (g1012) & (!g1030)) + ((g515) & (!g553) & (!g1000) & (g1001) & (!g1012) & (!g1030)) + ((g515) & (!g553) & (g1000) & (!g1001) & (!g1012) & (g1030)) + ((g515) & (!g553) & (g1000) & (!g1001) & (g1012) & (g1030)) + ((g515) & (!g553) & (g1000) & (g1001) & (!g1012) & (g1030)) + ((g515) & (!g553) & (g1000) & (g1001) & (g1012) & (!g1030)) + ((g515) & (!g553) & (g1000) & (g1001) & (g1012) & (g1030)) + ((g515) & (g553) & (!g1000) & (!g1001) & (!g1012) & (!g1030)) + ((g515) & (g553) & (g1000) & (!g1001) & (!g1012) & (g1030)) + ((g515) & (g553) & (g1000) & (!g1001) & (g1012) & (!g1030)) + ((g515) & (g553) & (g1000) & (!g1001) & (g1012) & (g1030)) + ((g515) & (g553) & (g1000) & (g1001) & (!g1012) & (!g1030)) + ((g515) & (g553) & (g1000) & (g1001) & (!g1012) & (g1030)) + ((g515) & (g553) & (g1000) & (g1001) & (g1012) & (!g1030)) + ((g515) & (g553) & (g1000) & (g1001) & (g1012) & (g1030)));
	assign g1061 = (((!g553) & (!g1001) & (g1012) & (!g1030)) + ((!g553) & (g1001) & (!g1012) & (!g1030)) + ((!g553) & (g1001) & (!g1012) & (g1030)) + ((!g553) & (g1001) & (g1012) & (g1030)) + ((g553) & (!g1001) & (!g1012) & (!g1030)) + ((g553) & (g1001) & (!g1012) & (g1030)) + ((g553) & (g1001) & (g1012) & (!g1030)) + ((g553) & (g1001) & (g1012) & (g1030)));
	assign g1062 = (((!g604) & (!g645) & (!g1003) & (g1004) & (g1011) & (!g1030)) + ((!g604) & (!g645) & (g1003) & (!g1004) & (!g1011) & (!g1030)) + ((!g604) & (!g645) & (g1003) & (!g1004) & (!g1011) & (g1030)) + ((!g604) & (!g645) & (g1003) & (!g1004) & (g1011) & (!g1030)) + ((!g604) & (!g645) & (g1003) & (!g1004) & (g1011) & (g1030)) + ((!g604) & (!g645) & (g1003) & (g1004) & (!g1011) & (!g1030)) + ((!g604) & (!g645) & (g1003) & (g1004) & (!g1011) & (g1030)) + ((!g604) & (!g645) & (g1003) & (g1004) & (g1011) & (g1030)) + ((!g604) & (g645) & (!g1003) & (!g1004) & (g1011) & (!g1030)) + ((!g604) & (g645) & (!g1003) & (g1004) & (!g1011) & (!g1030)) + ((!g604) & (g645) & (!g1003) & (g1004) & (g1011) & (!g1030)) + ((!g604) & (g645) & (g1003) & (!g1004) & (!g1011) & (!g1030)) + ((!g604) & (g645) & (g1003) & (!g1004) & (!g1011) & (g1030)) + ((!g604) & (g645) & (g1003) & (!g1004) & (g1011) & (g1030)) + ((!g604) & (g645) & (g1003) & (g1004) & (!g1011) & (g1030)) + ((!g604) & (g645) & (g1003) & (g1004) & (g1011) & (g1030)) + ((g604) & (!g645) & (!g1003) & (!g1004) & (!g1011) & (!g1030)) + ((g604) & (!g645) & (!g1003) & (!g1004) & (g1011) & (!g1030)) + ((g604) & (!g645) & (!g1003) & (g1004) & (!g1011) & (!g1030)) + ((g604) & (!g645) & (g1003) & (!g1004) & (!g1011) & (g1030)) + ((g604) & (!g645) & (g1003) & (!g1004) & (g1011) & (g1030)) + ((g604) & (!g645) & (g1003) & (g1004) & (!g1011) & (g1030)) + ((g604) & (!g645) & (g1003) & (g1004) & (g1011) & (!g1030)) + ((g604) & (!g645) & (g1003) & (g1004) & (g1011) & (g1030)) + ((g604) & (g645) & (!g1003) & (!g1004) & (!g1011) & (!g1030)) + ((g604) & (g645) & (g1003) & (!g1004) & (!g1011) & (g1030)) + ((g604) & (g645) & (g1003) & (!g1004) & (g1011) & (!g1030)) + ((g604) & (g645) & (g1003) & (!g1004) & (g1011) & (g1030)) + ((g604) & (g645) & (g1003) & (g1004) & (!g1011) & (!g1030)) + ((g604) & (g645) & (g1003) & (g1004) & (!g1011) & (g1030)) + ((g604) & (g645) & (g1003) & (g1004) & (g1011) & (!g1030)) + ((g604) & (g645) & (g1003) & (g1004) & (g1011) & (g1030)));
	assign g1063 = (((!g645) & (!g1004) & (g1011) & (!g1030)) + ((!g645) & (g1004) & (!g1011) & (!g1030)) + ((!g645) & (g1004) & (!g1011) & (g1030)) + ((!g645) & (g1004) & (g1011) & (g1030)) + ((g645) & (!g1004) & (!g1011) & (!g1030)) + ((g645) & (g1004) & (!g1011) & (g1030)) + ((g645) & (g1004) & (g1011) & (!g1030)) + ((g645) & (g1004) & (g1011) & (g1030)));
	assign g1064 = (((!g700) & (!g744) & (!g1006) & (g1007) & (g1010) & (!g1030)) + ((!g700) & (!g744) & (g1006) & (!g1007) & (!g1010) & (!g1030)) + ((!g700) & (!g744) & (g1006) & (!g1007) & (!g1010) & (g1030)) + ((!g700) & (!g744) & (g1006) & (!g1007) & (g1010) & (!g1030)) + ((!g700) & (!g744) & (g1006) & (!g1007) & (g1010) & (g1030)) + ((!g700) & (!g744) & (g1006) & (g1007) & (!g1010) & (!g1030)) + ((!g700) & (!g744) & (g1006) & (g1007) & (!g1010) & (g1030)) + ((!g700) & (!g744) & (g1006) & (g1007) & (g1010) & (g1030)) + ((!g700) & (g744) & (!g1006) & (!g1007) & (g1010) & (!g1030)) + ((!g700) & (g744) & (!g1006) & (g1007) & (!g1010) & (!g1030)) + ((!g700) & (g744) & (!g1006) & (g1007) & (g1010) & (!g1030)) + ((!g700) & (g744) & (g1006) & (!g1007) & (!g1010) & (!g1030)) + ((!g700) & (g744) & (g1006) & (!g1007) & (!g1010) & (g1030)) + ((!g700) & (g744) & (g1006) & (!g1007) & (g1010) & (g1030)) + ((!g700) & (g744) & (g1006) & (g1007) & (!g1010) & (g1030)) + ((!g700) & (g744) & (g1006) & (g1007) & (g1010) & (g1030)) + ((g700) & (!g744) & (!g1006) & (!g1007) & (!g1010) & (!g1030)) + ((g700) & (!g744) & (!g1006) & (!g1007) & (g1010) & (!g1030)) + ((g700) & (!g744) & (!g1006) & (g1007) & (!g1010) & (!g1030)) + ((g700) & (!g744) & (g1006) & (!g1007) & (!g1010) & (g1030)) + ((g700) & (!g744) & (g1006) & (!g1007) & (g1010) & (g1030)) + ((g700) & (!g744) & (g1006) & (g1007) & (!g1010) & (g1030)) + ((g700) & (!g744) & (g1006) & (g1007) & (g1010) & (!g1030)) + ((g700) & (!g744) & (g1006) & (g1007) & (g1010) & (g1030)) + ((g700) & (g744) & (!g1006) & (!g1007) & (!g1010) & (!g1030)) + ((g700) & (g744) & (g1006) & (!g1007) & (!g1010) & (g1030)) + ((g700) & (g744) & (g1006) & (!g1007) & (g1010) & (!g1030)) + ((g700) & (g744) & (g1006) & (!g1007) & (g1010) & (g1030)) + ((g700) & (g744) & (g1006) & (g1007) & (!g1010) & (!g1030)) + ((g700) & (g744) & (g1006) & (g1007) & (!g1010) & (g1030)) + ((g700) & (g744) & (g1006) & (g1007) & (g1010) & (!g1030)) + ((g700) & (g744) & (g1006) & (g1007) & (g1010) & (g1030)));
	assign g1065 = (((!g744) & (!g1007) & (g1010) & (!g1030)) + ((!g744) & (g1007) & (!g1010) & (!g1030)) + ((!g744) & (g1007) & (!g1010) & (g1030)) + ((!g744) & (g1007) & (g1010) & (g1030)) + ((g744) & (!g1007) & (!g1010) & (!g1030)) + ((g744) & (g1007) & (!g1010) & (g1030)) + ((g744) & (g1007) & (g1010) & (!g1030)) + ((g744) & (g1007) & (g1010) & (g1030)));
	assign g1066 = (((!g803) & (!g851) & (!g1009) & (g964) & (g966) & (!g1030)) + ((!g803) & (!g851) & (g1009) & (!g964) & (!g966) & (!g1030)) + ((!g803) & (!g851) & (g1009) & (!g964) & (!g966) & (g1030)) + ((!g803) & (!g851) & (g1009) & (!g964) & (g966) & (!g1030)) + ((!g803) & (!g851) & (g1009) & (!g964) & (g966) & (g1030)) + ((!g803) & (!g851) & (g1009) & (g964) & (!g966) & (!g1030)) + ((!g803) & (!g851) & (g1009) & (g964) & (!g966) & (g1030)) + ((!g803) & (!g851) & (g1009) & (g964) & (g966) & (g1030)) + ((!g803) & (g851) & (!g1009) & (!g964) & (g966) & (!g1030)) + ((!g803) & (g851) & (!g1009) & (g964) & (!g966) & (!g1030)) + ((!g803) & (g851) & (!g1009) & (g964) & (g966) & (!g1030)) + ((!g803) & (g851) & (g1009) & (!g964) & (!g966) & (!g1030)) + ((!g803) & (g851) & (g1009) & (!g964) & (!g966) & (g1030)) + ((!g803) & (g851) & (g1009) & (!g964) & (g966) & (g1030)) + ((!g803) & (g851) & (g1009) & (g964) & (!g966) & (g1030)) + ((!g803) & (g851) & (g1009) & (g964) & (g966) & (g1030)) + ((g803) & (!g851) & (!g1009) & (!g964) & (!g966) & (!g1030)) + ((g803) & (!g851) & (!g1009) & (!g964) & (g966) & (!g1030)) + ((g803) & (!g851) & (!g1009) & (g964) & (!g966) & (!g1030)) + ((g803) & (!g851) & (g1009) & (!g964) & (!g966) & (g1030)) + ((g803) & (!g851) & (g1009) & (!g964) & (g966) & (g1030)) + ((g803) & (!g851) & (g1009) & (g964) & (!g966) & (g1030)) + ((g803) & (!g851) & (g1009) & (g964) & (g966) & (!g1030)) + ((g803) & (!g851) & (g1009) & (g964) & (g966) & (g1030)) + ((g803) & (g851) & (!g1009) & (!g964) & (!g966) & (!g1030)) + ((g803) & (g851) & (g1009) & (!g964) & (!g966) & (g1030)) + ((g803) & (g851) & (g1009) & (!g964) & (g966) & (!g1030)) + ((g803) & (g851) & (g1009) & (!g964) & (g966) & (g1030)) + ((g803) & (g851) & (g1009) & (g964) & (!g966) & (!g1030)) + ((g803) & (g851) & (g1009) & (g964) & (!g966) & (g1030)) + ((g803) & (g851) & (g1009) & (g964) & (g966) & (!g1030)) + ((g803) & (g851) & (g1009) & (g964) & (g966) & (g1030)));
	assign g1067 = (((!g744) & (!g803) & (g1066) & (g1031) & (g1037)) + ((!g744) & (g803) & (g1066) & (!g1031) & (g1037)) + ((!g744) & (g803) & (g1066) & (g1031) & (!g1037)) + ((!g744) & (g803) & (g1066) & (g1031) & (g1037)) + ((g744) & (!g803) & (!g1066) & (g1031) & (g1037)) + ((g744) & (!g803) & (g1066) & (!g1031) & (!g1037)) + ((g744) & (!g803) & (g1066) & (!g1031) & (g1037)) + ((g744) & (!g803) & (g1066) & (g1031) & (!g1037)) + ((g744) & (!g803) & (g1066) & (g1031) & (g1037)) + ((g744) & (g803) & (!g1066) & (!g1031) & (g1037)) + ((g744) & (g803) & (!g1066) & (g1031) & (!g1037)) + ((g744) & (g803) & (!g1066) & (g1031) & (g1037)) + ((g744) & (g803) & (g1066) & (!g1031) & (!g1037)) + ((g744) & (g803) & (g1066) & (!g1031) & (g1037)) + ((g744) & (g803) & (g1066) & (g1031) & (!g1037)) + ((g744) & (g803) & (g1066) & (g1031) & (g1037)));
	assign g1068 = (((!g645) & (!g700) & (g1064) & (g1065) & (g1067)) + ((!g645) & (g700) & (g1064) & (!g1065) & (g1067)) + ((!g645) & (g700) & (g1064) & (g1065) & (!g1067)) + ((!g645) & (g700) & (g1064) & (g1065) & (g1067)) + ((g645) & (!g700) & (!g1064) & (g1065) & (g1067)) + ((g645) & (!g700) & (g1064) & (!g1065) & (!g1067)) + ((g645) & (!g700) & (g1064) & (!g1065) & (g1067)) + ((g645) & (!g700) & (g1064) & (g1065) & (!g1067)) + ((g645) & (!g700) & (g1064) & (g1065) & (g1067)) + ((g645) & (g700) & (!g1064) & (!g1065) & (g1067)) + ((g645) & (g700) & (!g1064) & (g1065) & (!g1067)) + ((g645) & (g700) & (!g1064) & (g1065) & (g1067)) + ((g645) & (g700) & (g1064) & (!g1065) & (!g1067)) + ((g645) & (g700) & (g1064) & (!g1065) & (g1067)) + ((g645) & (g700) & (g1064) & (g1065) & (!g1067)) + ((g645) & (g700) & (g1064) & (g1065) & (g1067)));
	assign g1069 = (((!g553) & (!g604) & (g1062) & (g1063) & (g1068)) + ((!g553) & (g604) & (g1062) & (!g1063) & (g1068)) + ((!g553) & (g604) & (g1062) & (g1063) & (!g1068)) + ((!g553) & (g604) & (g1062) & (g1063) & (g1068)) + ((g553) & (!g604) & (!g1062) & (g1063) & (g1068)) + ((g553) & (!g604) & (g1062) & (!g1063) & (!g1068)) + ((g553) & (!g604) & (g1062) & (!g1063) & (g1068)) + ((g553) & (!g604) & (g1062) & (g1063) & (!g1068)) + ((g553) & (!g604) & (g1062) & (g1063) & (g1068)) + ((g553) & (g604) & (!g1062) & (!g1063) & (g1068)) + ((g553) & (g604) & (!g1062) & (g1063) & (!g1068)) + ((g553) & (g604) & (!g1062) & (g1063) & (g1068)) + ((g553) & (g604) & (g1062) & (!g1063) & (!g1068)) + ((g553) & (g604) & (g1062) & (!g1063) & (g1068)) + ((g553) & (g604) & (g1062) & (g1063) & (!g1068)) + ((g553) & (g604) & (g1062) & (g1063) & (g1068)));
	assign g1070 = (((!g468) & (!g515) & (g1060) & (g1061) & (g1069)) + ((!g468) & (g515) & (g1060) & (!g1061) & (g1069)) + ((!g468) & (g515) & (g1060) & (g1061) & (!g1069)) + ((!g468) & (g515) & (g1060) & (g1061) & (g1069)) + ((g468) & (!g515) & (!g1060) & (g1061) & (g1069)) + ((g468) & (!g515) & (g1060) & (!g1061) & (!g1069)) + ((g468) & (!g515) & (g1060) & (!g1061) & (g1069)) + ((g468) & (!g515) & (g1060) & (g1061) & (!g1069)) + ((g468) & (!g515) & (g1060) & (g1061) & (g1069)) + ((g468) & (g515) & (!g1060) & (!g1061) & (g1069)) + ((g468) & (g515) & (!g1060) & (g1061) & (!g1069)) + ((g468) & (g515) & (!g1060) & (g1061) & (g1069)) + ((g468) & (g515) & (g1060) & (!g1061) & (!g1069)) + ((g468) & (g515) & (g1060) & (!g1061) & (g1069)) + ((g468) & (g515) & (g1060) & (g1061) & (!g1069)) + ((g468) & (g515) & (g1060) & (g1061) & (g1069)));
	assign g1071 = (((!g390) & (!g433) & (g1058) & (g1059) & (g1070)) + ((!g390) & (g433) & (g1058) & (!g1059) & (g1070)) + ((!g390) & (g433) & (g1058) & (g1059) & (!g1070)) + ((!g390) & (g433) & (g1058) & (g1059) & (g1070)) + ((g390) & (!g433) & (!g1058) & (g1059) & (g1070)) + ((g390) & (!g433) & (g1058) & (!g1059) & (!g1070)) + ((g390) & (!g433) & (g1058) & (!g1059) & (g1070)) + ((g390) & (!g433) & (g1058) & (g1059) & (!g1070)) + ((g390) & (!g433) & (g1058) & (g1059) & (g1070)) + ((g390) & (g433) & (!g1058) & (!g1059) & (g1070)) + ((g390) & (g433) & (!g1058) & (g1059) & (!g1070)) + ((g390) & (g433) & (!g1058) & (g1059) & (g1070)) + ((g390) & (g433) & (g1058) & (!g1059) & (!g1070)) + ((g390) & (g433) & (g1058) & (!g1059) & (g1070)) + ((g390) & (g433) & (g1058) & (g1059) & (!g1070)) + ((g390) & (g433) & (g1058) & (g1059) & (g1070)));
	assign g1072 = (((!g319) & (!g358) & (g1056) & (g1057) & (g1071)) + ((!g319) & (g358) & (g1056) & (!g1057) & (g1071)) + ((!g319) & (g358) & (g1056) & (g1057) & (!g1071)) + ((!g319) & (g358) & (g1056) & (g1057) & (g1071)) + ((g319) & (!g358) & (!g1056) & (g1057) & (g1071)) + ((g319) & (!g358) & (g1056) & (!g1057) & (!g1071)) + ((g319) & (!g358) & (g1056) & (!g1057) & (g1071)) + ((g319) & (!g358) & (g1056) & (g1057) & (!g1071)) + ((g319) & (!g358) & (g1056) & (g1057) & (g1071)) + ((g319) & (g358) & (!g1056) & (!g1057) & (g1071)) + ((g319) & (g358) & (!g1056) & (g1057) & (!g1071)) + ((g319) & (g358) & (!g1056) & (g1057) & (g1071)) + ((g319) & (g358) & (g1056) & (!g1057) & (!g1071)) + ((g319) & (g358) & (g1056) & (!g1057) & (g1071)) + ((g319) & (g358) & (g1056) & (g1057) & (!g1071)) + ((g319) & (g358) & (g1056) & (g1057) & (g1071)));
	assign g1073 = (((!g255) & (!g290) & (g1054) & (g1055) & (g1072)) + ((!g255) & (g290) & (g1054) & (!g1055) & (g1072)) + ((!g255) & (g290) & (g1054) & (g1055) & (!g1072)) + ((!g255) & (g290) & (g1054) & (g1055) & (g1072)) + ((g255) & (!g290) & (!g1054) & (g1055) & (g1072)) + ((g255) & (!g290) & (g1054) & (!g1055) & (!g1072)) + ((g255) & (!g290) & (g1054) & (!g1055) & (g1072)) + ((g255) & (!g290) & (g1054) & (g1055) & (!g1072)) + ((g255) & (!g290) & (g1054) & (g1055) & (g1072)) + ((g255) & (g290) & (!g1054) & (!g1055) & (g1072)) + ((g255) & (g290) & (!g1054) & (g1055) & (!g1072)) + ((g255) & (g290) & (!g1054) & (g1055) & (g1072)) + ((g255) & (g290) & (g1054) & (!g1055) & (!g1072)) + ((g255) & (g290) & (g1054) & (!g1055) & (g1072)) + ((g255) & (g290) & (g1054) & (g1055) & (!g1072)) + ((g255) & (g290) & (g1054) & (g1055) & (g1072)));
	assign g1074 = (((!g198) & (!g229) & (g1052) & (g1053) & (g1073)) + ((!g198) & (g229) & (g1052) & (!g1053) & (g1073)) + ((!g198) & (g229) & (g1052) & (g1053) & (!g1073)) + ((!g198) & (g229) & (g1052) & (g1053) & (g1073)) + ((g198) & (!g229) & (!g1052) & (g1053) & (g1073)) + ((g198) & (!g229) & (g1052) & (!g1053) & (!g1073)) + ((g198) & (!g229) & (g1052) & (!g1053) & (g1073)) + ((g198) & (!g229) & (g1052) & (g1053) & (!g1073)) + ((g198) & (!g229) & (g1052) & (g1053) & (g1073)) + ((g198) & (g229) & (!g1052) & (!g1053) & (g1073)) + ((g198) & (g229) & (!g1052) & (g1053) & (!g1073)) + ((g198) & (g229) & (!g1052) & (g1053) & (g1073)) + ((g198) & (g229) & (g1052) & (!g1053) & (!g1073)) + ((g198) & (g229) & (g1052) & (!g1053) & (g1073)) + ((g198) & (g229) & (g1052) & (g1053) & (!g1073)) + ((g198) & (g229) & (g1052) & (g1053) & (g1073)));
	assign g1075 = (((!g147) & (!g174) & (g1050) & (g1051) & (g1074)) + ((!g147) & (g174) & (g1050) & (!g1051) & (g1074)) + ((!g147) & (g174) & (g1050) & (g1051) & (!g1074)) + ((!g147) & (g174) & (g1050) & (g1051) & (g1074)) + ((g147) & (!g174) & (!g1050) & (g1051) & (g1074)) + ((g147) & (!g174) & (g1050) & (!g1051) & (!g1074)) + ((g147) & (!g174) & (g1050) & (!g1051) & (g1074)) + ((g147) & (!g174) & (g1050) & (g1051) & (!g1074)) + ((g147) & (!g174) & (g1050) & (g1051) & (g1074)) + ((g147) & (g174) & (!g1050) & (!g1051) & (g1074)) + ((g147) & (g174) & (!g1050) & (g1051) & (!g1074)) + ((g147) & (g174) & (!g1050) & (g1051) & (g1074)) + ((g147) & (g174) & (g1050) & (!g1051) & (!g1074)) + ((g147) & (g174) & (g1050) & (!g1051) & (g1074)) + ((g147) & (g174) & (g1050) & (g1051) & (!g1074)) + ((g147) & (g174) & (g1050) & (g1051) & (g1074)));
	assign g1076 = (((!g104) & (!g127) & (g1048) & (g1049) & (g1075)) + ((!g104) & (g127) & (g1048) & (!g1049) & (g1075)) + ((!g104) & (g127) & (g1048) & (g1049) & (!g1075)) + ((!g104) & (g127) & (g1048) & (g1049) & (g1075)) + ((g104) & (!g127) & (!g1048) & (g1049) & (g1075)) + ((g104) & (!g127) & (g1048) & (!g1049) & (!g1075)) + ((g104) & (!g127) & (g1048) & (!g1049) & (g1075)) + ((g104) & (!g127) & (g1048) & (g1049) & (!g1075)) + ((g104) & (!g127) & (g1048) & (g1049) & (g1075)) + ((g104) & (g127) & (!g1048) & (!g1049) & (g1075)) + ((g104) & (g127) & (!g1048) & (g1049) & (!g1075)) + ((g104) & (g127) & (!g1048) & (g1049) & (g1075)) + ((g104) & (g127) & (g1048) & (!g1049) & (!g1075)) + ((g104) & (g127) & (g1048) & (!g1049) & (g1075)) + ((g104) & (g127) & (g1048) & (g1049) & (!g1075)) + ((g104) & (g127) & (g1048) & (g1049) & (g1075)));
	assign g1077 = (((!g68) & (!g87) & (g1046) & (g1047) & (g1076)) + ((!g68) & (g87) & (g1046) & (!g1047) & (g1076)) + ((!g68) & (g87) & (g1046) & (g1047) & (!g1076)) + ((!g68) & (g87) & (g1046) & (g1047) & (g1076)) + ((g68) & (!g87) & (!g1046) & (g1047) & (g1076)) + ((g68) & (!g87) & (g1046) & (!g1047) & (!g1076)) + ((g68) & (!g87) & (g1046) & (!g1047) & (g1076)) + ((g68) & (!g87) & (g1046) & (g1047) & (!g1076)) + ((g68) & (!g87) & (g1046) & (g1047) & (g1076)) + ((g68) & (g87) & (!g1046) & (!g1047) & (g1076)) + ((g68) & (g87) & (!g1046) & (g1047) & (!g1076)) + ((g68) & (g87) & (!g1046) & (g1047) & (g1076)) + ((g68) & (g87) & (g1046) & (!g1047) & (!g1076)) + ((g68) & (g87) & (g1046) & (!g1047) & (g1076)) + ((g68) & (g87) & (g1046) & (g1047) & (!g1076)) + ((g68) & (g87) & (g1046) & (g1047) & (g1076)));
	assign g1078 = (((!g39) & (!g54) & (g1044) & (g1045) & (g1077)) + ((!g39) & (g54) & (g1044) & (!g1045) & (g1077)) + ((!g39) & (g54) & (g1044) & (g1045) & (!g1077)) + ((!g39) & (g54) & (g1044) & (g1045) & (g1077)) + ((g39) & (!g54) & (!g1044) & (g1045) & (g1077)) + ((g39) & (!g54) & (g1044) & (!g1045) & (!g1077)) + ((g39) & (!g54) & (g1044) & (!g1045) & (g1077)) + ((g39) & (!g54) & (g1044) & (g1045) & (!g1077)) + ((g39) & (!g54) & (g1044) & (g1045) & (g1077)) + ((g39) & (g54) & (!g1044) & (!g1045) & (g1077)) + ((g39) & (g54) & (!g1044) & (g1045) & (!g1077)) + ((g39) & (g54) & (!g1044) & (g1045) & (g1077)) + ((g39) & (g54) & (g1044) & (!g1045) & (!g1077)) + ((g39) & (g54) & (g1044) & (!g1045) & (g1077)) + ((g39) & (g54) & (g1044) & (g1045) & (!g1077)) + ((g39) & (g54) & (g1044) & (g1045) & (g1077)));
	assign g1079 = (((!g18) & (!g27) & (g1042) & (g1043) & (g1078)) + ((!g18) & (g27) & (g1042) & (!g1043) & (g1078)) + ((!g18) & (g27) & (g1042) & (g1043) & (!g1078)) + ((!g18) & (g27) & (g1042) & (g1043) & (g1078)) + ((g18) & (!g27) & (!g1042) & (g1043) & (g1078)) + ((g18) & (!g27) & (g1042) & (!g1043) & (!g1078)) + ((g18) & (!g27) & (g1042) & (!g1043) & (g1078)) + ((g18) & (!g27) & (g1042) & (g1043) & (!g1078)) + ((g18) & (!g27) & (g1042) & (g1043) & (g1078)) + ((g18) & (g27) & (!g1042) & (!g1043) & (g1078)) + ((g18) & (g27) & (!g1042) & (g1043) & (!g1078)) + ((g18) & (g27) & (!g1042) & (g1043) & (g1078)) + ((g18) & (g27) & (g1042) & (!g1043) & (!g1078)) + ((g18) & (g27) & (g1042) & (!g1043) & (g1078)) + ((g18) & (g27) & (g1042) & (g1043) & (!g1078)) + ((g18) & (g27) & (g1042) & (g1043) & (g1078)));
	assign g1080 = (((!g2) & (!g8) & (g1040) & (g1041) & (g1079)) + ((!g2) & (g8) & (g1040) & (!g1041) & (g1079)) + ((!g2) & (g8) & (g1040) & (g1041) & (!g1079)) + ((!g2) & (g8) & (g1040) & (g1041) & (g1079)) + ((g2) & (!g8) & (!g1040) & (g1041) & (g1079)) + ((g2) & (!g8) & (g1040) & (!g1041) & (!g1079)) + ((g2) & (!g8) & (g1040) & (!g1041) & (g1079)) + ((g2) & (!g8) & (g1040) & (g1041) & (!g1079)) + ((g2) & (!g8) & (g1040) & (g1041) & (g1079)) + ((g2) & (g8) & (!g1040) & (!g1041) & (g1079)) + ((g2) & (g8) & (!g1040) & (g1041) & (!g1079)) + ((g2) & (g8) & (!g1040) & (g1041) & (g1079)) + ((g2) & (g8) & (g1040) & (!g1041) & (!g1079)) + ((g2) & (g8) & (g1040) & (!g1041) & (g1079)) + ((g2) & (g8) & (g1040) & (g1041) & (!g1079)) + ((g2) & (g8) & (g1040) & (g1041) & (g1079)));
	assign g1081 = (((!g2) & (!g968) & (g1023) & (!g1030)) + ((!g2) & (g968) & (!g1023) & (!g1030)) + ((!g2) & (g968) & (!g1023) & (g1030)) + ((!g2) & (g968) & (g1023) & (g1030)) + ((g2) & (!g968) & (!g1023) & (!g1030)) + ((g2) & (g968) & (!g1023) & (g1030)) + ((g2) & (g968) & (g1023) & (!g1030)) + ((g2) & (g968) & (g1023) & (g1030)));
	assign g1082 = (((!g1) & (!g967) & (!g1026) & (!g1028) & (g1029)) + ((!g1) & (!g967) & (!g1026) & (g1028) & (!g1029)) + ((!g1) & (!g967) & (!g1026) & (g1028) & (g1029)) + ((!g1) & (g967) & (g1026) & (!g1028) & (!g1029)) + ((!g1) & (g967) & (g1026) & (!g1028) & (g1029)) + ((!g1) & (g967) & (g1026) & (g1028) & (!g1029)) + ((!g1) & (g967) & (g1026) & (g1028) & (g1029)) + ((g1) & (!g967) & (!g1026) & (!g1028) & (g1029)) + ((g1) & (!g967) & (!g1026) & (g1028) & (g1029)) + ((g1) & (g967) & (g1026) & (!g1028) & (!g1029)) + ((g1) & (g967) & (g1026) & (!g1028) & (g1029)) + ((g1) & (g967) & (g1026) & (g1028) & (!g1029)) + ((g1) & (g967) & (g1026) & (g1028) & (g1029)));
	assign g1083 = (((!g4) & (!g1) & (!g1039) & (!g1080) & (!g1081) & (!g1082)) + ((!g4) & (g1) & (!g1039) & (!g1080) & (!g1081) & (!g1082)) + ((!g4) & (g1) & (!g1039) & (!g1080) & (!g1081) & (g1082)) + ((!g4) & (g1) & (!g1039) & (!g1080) & (g1081) & (!g1082)) + ((!g4) & (g1) & (!g1039) & (!g1080) & (g1081) & (g1082)) + ((!g4) & (g1) & (!g1039) & (g1080) & (!g1081) & (!g1082)) + ((!g4) & (g1) & (!g1039) & (g1080) & (!g1081) & (g1082)) + ((!g4) & (g1) & (!g1039) & (g1080) & (g1081) & (!g1082)) + ((!g4) & (g1) & (!g1039) & (g1080) & (g1081) & (g1082)) + ((!g4) & (g1) & (g1039) & (!g1080) & (!g1081) & (!g1082)) + ((!g4) & (g1) & (g1039) & (!g1080) & (!g1081) & (g1082)) + ((g4) & (!g1) & (!g1039) & (!g1080) & (!g1081) & (!g1082)) + ((g4) & (!g1) & (!g1039) & (!g1080) & (g1081) & (!g1082)) + ((g4) & (!g1) & (!g1039) & (g1080) & (!g1081) & (!g1082)) + ((g4) & (g1) & (!g1039) & (!g1080) & (!g1081) & (!g1082)) + ((g4) & (g1) & (!g1039) & (!g1080) & (!g1081) & (g1082)) + ((g4) & (g1) & (!g1039) & (!g1080) & (g1081) & (!g1082)) + ((g4) & (g1) & (!g1039) & (!g1080) & (g1081) & (g1082)) + ((g4) & (g1) & (!g1039) & (g1080) & (!g1081) & (!g1082)) + ((g4) & (g1) & (!g1039) & (g1080) & (!g1081) & (g1082)) + ((g4) & (g1) & (!g1039) & (g1080) & (g1081) & (!g1082)) + ((g4) & (g1) & (!g1039) & (g1080) & (g1081) & (g1082)) + ((g4) & (g1) & (g1039) & (!g1080) & (!g1081) & (!g1082)) + ((g4) & (g1) & (g1039) & (!g1080) & (!g1081) & (g1082)) + ((g4) & (g1) & (g1039) & (!g1080) & (g1081) & (!g1082)) + ((g4) & (g1) & (g1039) & (!g1080) & (g1081) & (g1082)) + ((g4) & (g1) & (g1039) & (g1080) & (!g1081) & (!g1082)) + ((g4) & (g1) & (g1039) & (g1080) & (!g1081) & (g1082)));
	assign g1084 = (((!g803) & (!g1031) & (g1037) & (!g1038) & (!g1083)) + ((!g803) & (!g1031) & (g1037) & (g1038) & (!g1083)) + ((!g803) & (!g1031) & (g1037) & (g1038) & (g1083)) + ((!g803) & (g1031) & (!g1037) & (!g1038) & (!g1083)) + ((!g803) & (g1031) & (!g1037) & (!g1038) & (g1083)) + ((!g803) & (g1031) & (!g1037) & (g1038) & (!g1083)) + ((!g803) & (g1031) & (!g1037) & (g1038) & (g1083)) + ((!g803) & (g1031) & (g1037) & (!g1038) & (g1083)) + ((g803) & (!g1031) & (!g1037) & (!g1038) & (!g1083)) + ((g803) & (!g1031) & (!g1037) & (g1038) & (!g1083)) + ((g803) & (!g1031) & (!g1037) & (g1038) & (g1083)) + ((g803) & (g1031) & (!g1037) & (!g1038) & (g1083)) + ((g803) & (g1031) & (g1037) & (!g1038) & (!g1083)) + ((g803) & (g1031) & (g1037) & (!g1038) & (g1083)) + ((g803) & (g1031) & (g1037) & (g1038) & (!g1083)) + ((g803) & (g1031) & (g1037) & (g1038) & (g1083)));
	assign g1085 = (((!g851) & (!g914) & (g1034) & (g1036)) + ((!g851) & (g914) & (!g1034) & (g1036)) + ((!g851) & (g914) & (g1034) & (!g1036)) + ((!g851) & (g914) & (g1034) & (g1036)) + ((g851) & (!g914) & (!g1034) & (!g1036)) + ((g851) & (!g914) & (!g1034) & (g1036)) + ((g851) & (!g914) & (g1034) & (!g1036)) + ((g851) & (g914) & (!g1034) & (!g1036)));
	assign g1086 = (((!g1033) & (!g1038) & (!g1083) & (g1085)) + ((!g1033) & (g1038) & (!g1083) & (g1085)) + ((!g1033) & (g1038) & (g1083) & (g1085)) + ((g1033) & (!g1038) & (!g1083) & (!g1085)) + ((g1033) & (!g1038) & (g1083) & (!g1085)) + ((g1033) & (!g1038) & (g1083) & (g1085)) + ((g1033) & (g1038) & (!g1083) & (!g1085)) + ((g1033) & (g1038) & (g1083) & (!g1085)));
	assign g1087 = (((!g914) & (!g1034) & (g1036) & (!g1038) & (!g1083)) + ((!g914) & (!g1034) & (g1036) & (g1038) & (!g1083)) + ((!g914) & (!g1034) & (g1036) & (g1038) & (g1083)) + ((!g914) & (g1034) & (!g1036) & (!g1038) & (!g1083)) + ((!g914) & (g1034) & (!g1036) & (!g1038) & (g1083)) + ((!g914) & (g1034) & (!g1036) & (g1038) & (!g1083)) + ((!g914) & (g1034) & (!g1036) & (g1038) & (g1083)) + ((!g914) & (g1034) & (g1036) & (!g1038) & (g1083)) + ((g914) & (!g1034) & (!g1036) & (!g1038) & (!g1083)) + ((g914) & (!g1034) & (!g1036) & (g1038) & (!g1083)) + ((g914) & (!g1034) & (!g1036) & (g1038) & (g1083)) + ((g914) & (g1034) & (!g1036) & (!g1038) & (g1083)) + ((g914) & (g1034) & (g1036) & (!g1038) & (!g1083)) + ((g914) & (g1034) & (g1036) & (!g1038) & (g1083)) + ((g914) & (g1034) & (g1036) & (g1038) & (!g1083)) + ((g914) & (g1034) & (g1036) & (g1038) & (g1083)));
	assign g1088 = (((!g1032) & (!ax60x) & (!g1030) & (g1035)) + ((!g1032) & (!ax60x) & (g1030) & (g1035)) + ((!g1032) & (ax60x) & (!g1030) & (!g1035)) + ((!g1032) & (ax60x) & (!g1030) & (g1035)) + ((g1032) & (!ax60x) & (!g1030) & (!g1035)) + ((g1032) & (!ax60x) & (g1030) & (!g1035)) + ((g1032) & (ax60x) & (g1030) & (!g1035)) + ((g1032) & (ax60x) & (g1030) & (g1035)));
	assign g1089 = (((!ax60x) & (!ax61x) & (!g1030) & (!g1038) & (!g1083) & (g1088)) + ((!ax60x) & (!ax61x) & (!g1030) & (!g1038) & (g1083) & (!g1088)) + ((!ax60x) & (!ax61x) & (!g1030) & (!g1038) & (g1083) & (g1088)) + ((!ax60x) & (!ax61x) & (!g1030) & (g1038) & (!g1083) & (g1088)) + ((!ax60x) & (!ax61x) & (!g1030) & (g1038) & (g1083) & (g1088)) + ((!ax60x) & (!ax61x) & (g1030) & (!g1038) & (!g1083) & (!g1088)) + ((!ax60x) & (!ax61x) & (g1030) & (g1038) & (!g1083) & (!g1088)) + ((!ax60x) & (!ax61x) & (g1030) & (g1038) & (g1083) & (!g1088)) + ((!ax60x) & (ax61x) & (!g1030) & (!g1038) & (!g1083) & (!g1088)) + ((!ax60x) & (ax61x) & (!g1030) & (g1038) & (!g1083) & (!g1088)) + ((!ax60x) & (ax61x) & (!g1030) & (g1038) & (g1083) & (!g1088)) + ((!ax60x) & (ax61x) & (g1030) & (!g1038) & (!g1083) & (g1088)) + ((!ax60x) & (ax61x) & (g1030) & (!g1038) & (g1083) & (!g1088)) + ((!ax60x) & (ax61x) & (g1030) & (!g1038) & (g1083) & (g1088)) + ((!ax60x) & (ax61x) & (g1030) & (g1038) & (!g1083) & (g1088)) + ((!ax60x) & (ax61x) & (g1030) & (g1038) & (g1083) & (g1088)) + ((ax60x) & (!ax61x) & (!g1030) & (!g1038) & (!g1083) & (!g1088)) + ((ax60x) & (!ax61x) & (!g1030) & (g1038) & (!g1083) & (!g1088)) + ((ax60x) & (!ax61x) & (!g1030) & (g1038) & (g1083) & (!g1088)) + ((ax60x) & (!ax61x) & (g1030) & (!g1038) & (!g1083) & (!g1088)) + ((ax60x) & (!ax61x) & (g1030) & (g1038) & (!g1083) & (!g1088)) + ((ax60x) & (!ax61x) & (g1030) & (g1038) & (g1083) & (!g1088)) + ((ax60x) & (ax61x) & (!g1030) & (!g1038) & (!g1083) & (g1088)) + ((ax60x) & (ax61x) & (!g1030) & (!g1038) & (g1083) & (!g1088)) + ((ax60x) & (ax61x) & (!g1030) & (!g1038) & (g1083) & (g1088)) + ((ax60x) & (ax61x) & (!g1030) & (g1038) & (!g1083) & (g1088)) + ((ax60x) & (ax61x) & (!g1030) & (g1038) & (g1083) & (g1088)) + ((ax60x) & (ax61x) & (g1030) & (!g1038) & (!g1083) & (g1088)) + ((ax60x) & (ax61x) & (g1030) & (!g1038) & (g1083) & (!g1088)) + ((ax60x) & (ax61x) & (g1030) & (!g1038) & (g1083) & (g1088)) + ((ax60x) & (ax61x) & (g1030) & (g1038) & (!g1083) & (g1088)) + ((ax60x) & (ax61x) & (g1030) & (g1038) & (g1083) & (g1088)));
	assign g1090 = (((!ax60x) & (!g1030) & (!g1035) & (!g1038) & (g1083)) + ((!ax60x) & (!g1030) & (g1035) & (!g1038) & (!g1083)) + ((!ax60x) & (!g1030) & (g1035) & (!g1038) & (g1083)) + ((!ax60x) & (!g1030) & (g1035) & (g1038) & (!g1083)) + ((!ax60x) & (!g1030) & (g1035) & (g1038) & (g1083)) + ((!ax60x) & (g1030) & (g1035) & (!g1038) & (!g1083)) + ((!ax60x) & (g1030) & (g1035) & (g1038) & (!g1083)) + ((!ax60x) & (g1030) & (g1035) & (g1038) & (g1083)) + ((ax60x) & (!g1030) & (!g1035) & (!g1038) & (!g1083)) + ((ax60x) & (!g1030) & (!g1035) & (g1038) & (!g1083)) + ((ax60x) & (!g1030) & (!g1035) & (g1038) & (g1083)) + ((ax60x) & (g1030) & (!g1035) & (!g1038) & (!g1083)) + ((ax60x) & (g1030) & (!g1035) & (!g1038) & (g1083)) + ((ax60x) & (g1030) & (!g1035) & (g1038) & (!g1083)) + ((ax60x) & (g1030) & (!g1035) & (g1038) & (g1083)) + ((ax60x) & (g1030) & (g1035) & (!g1038) & (g1083)));
	assign g1091 = (((!ax56x) & (!ax57x)));
	assign g1092 = (((!g1030) & (!ax58x) & (!ax59x) & (!g1038) & (!g1083) & (!g1091)) + ((!g1030) & (!ax58x) & (!ax59x) & (g1038) & (!g1083) & (!g1091)) + ((!g1030) & (!ax58x) & (!ax59x) & (g1038) & (g1083) & (!g1091)) + ((!g1030) & (!ax58x) & (ax59x) & (!g1038) & (g1083) & (!g1091)) + ((!g1030) & (ax58x) & (ax59x) & (!g1038) & (g1083) & (!g1091)) + ((!g1030) & (ax58x) & (ax59x) & (!g1038) & (g1083) & (g1091)) + ((g1030) & (!ax58x) & (!ax59x) & (!g1038) & (!g1083) & (!g1091)) + ((g1030) & (!ax58x) & (!ax59x) & (!g1038) & (!g1083) & (g1091)) + ((g1030) & (!ax58x) & (!ax59x) & (!g1038) & (g1083) & (!g1091)) + ((g1030) & (!ax58x) & (!ax59x) & (g1038) & (!g1083) & (!g1091)) + ((g1030) & (!ax58x) & (!ax59x) & (g1038) & (!g1083) & (g1091)) + ((g1030) & (!ax58x) & (!ax59x) & (g1038) & (g1083) & (!g1091)) + ((g1030) & (!ax58x) & (!ax59x) & (g1038) & (g1083) & (g1091)) + ((g1030) & (!ax58x) & (ax59x) & (!g1038) & (!g1083) & (!g1091)) + ((g1030) & (!ax58x) & (ax59x) & (!g1038) & (g1083) & (!g1091)) + ((g1030) & (!ax58x) & (ax59x) & (!g1038) & (g1083) & (g1091)) + ((g1030) & (!ax58x) & (ax59x) & (g1038) & (!g1083) & (!g1091)) + ((g1030) & (!ax58x) & (ax59x) & (g1038) & (g1083) & (!g1091)) + ((g1030) & (ax58x) & (!ax59x) & (!g1038) & (g1083) & (!g1091)) + ((g1030) & (ax58x) & (!ax59x) & (!g1038) & (g1083) & (g1091)) + ((g1030) & (ax58x) & (ax59x) & (!g1038) & (!g1083) & (!g1091)) + ((g1030) & (ax58x) & (ax59x) & (!g1038) & (!g1083) & (g1091)) + ((g1030) & (ax58x) & (ax59x) & (!g1038) & (g1083) & (!g1091)) + ((g1030) & (ax58x) & (ax59x) & (!g1038) & (g1083) & (g1091)) + ((g1030) & (ax58x) & (ax59x) & (g1038) & (!g1083) & (!g1091)) + ((g1030) & (ax58x) & (ax59x) & (g1038) & (!g1083) & (g1091)) + ((g1030) & (ax58x) & (ax59x) & (g1038) & (g1083) & (!g1091)) + ((g1030) & (ax58x) & (ax59x) & (g1038) & (g1083) & (g1091)));
	assign g1093 = (((!g914) & (!g1032) & (g1089) & (g1090) & (g1092)) + ((!g914) & (g1032) & (g1089) & (!g1090) & (g1092)) + ((!g914) & (g1032) & (g1089) & (g1090) & (!g1092)) + ((!g914) & (g1032) & (g1089) & (g1090) & (g1092)) + ((g914) & (!g1032) & (!g1089) & (g1090) & (g1092)) + ((g914) & (!g1032) & (g1089) & (!g1090) & (!g1092)) + ((g914) & (!g1032) & (g1089) & (!g1090) & (g1092)) + ((g914) & (!g1032) & (g1089) & (g1090) & (!g1092)) + ((g914) & (!g1032) & (g1089) & (g1090) & (g1092)) + ((g914) & (g1032) & (!g1089) & (!g1090) & (g1092)) + ((g914) & (g1032) & (!g1089) & (g1090) & (!g1092)) + ((g914) & (g1032) & (!g1089) & (g1090) & (g1092)) + ((g914) & (g1032) & (g1089) & (!g1090) & (!g1092)) + ((g914) & (g1032) & (g1089) & (!g1090) & (g1092)) + ((g914) & (g1032) & (g1089) & (g1090) & (!g1092)) + ((g914) & (g1032) & (g1089) & (g1090) & (g1092)));
	assign g1094 = (((!g803) & (!g851) & (g1086) & (g1087) & (g1093)) + ((!g803) & (g851) & (g1086) & (!g1087) & (g1093)) + ((!g803) & (g851) & (g1086) & (g1087) & (!g1093)) + ((!g803) & (g851) & (g1086) & (g1087) & (g1093)) + ((g803) & (!g851) & (!g1086) & (g1087) & (g1093)) + ((g803) & (!g851) & (g1086) & (!g1087) & (!g1093)) + ((g803) & (!g851) & (g1086) & (!g1087) & (g1093)) + ((g803) & (!g851) & (g1086) & (g1087) & (!g1093)) + ((g803) & (!g851) & (g1086) & (g1087) & (g1093)) + ((g803) & (g851) & (!g1086) & (!g1087) & (g1093)) + ((g803) & (g851) & (!g1086) & (g1087) & (!g1093)) + ((g803) & (g851) & (!g1086) & (g1087) & (g1093)) + ((g803) & (g851) & (g1086) & (!g1087) & (!g1093)) + ((g803) & (g851) & (g1086) & (!g1087) & (g1093)) + ((g803) & (g851) & (g1086) & (g1087) & (!g1093)) + ((g803) & (g851) & (g1086) & (g1087) & (g1093)));
	assign g1095 = (((!g4) & (!g1080) & (!g1081) & (!g1038) & (!g1083)) + ((!g4) & (!g1080) & (!g1081) & (g1038) & (!g1083)) + ((!g4) & (!g1080) & (!g1081) & (g1038) & (g1083)) + ((!g4) & (!g1080) & (g1081) & (!g1038) & (g1083)) + ((!g4) & (g1080) & (g1081) & (!g1038) & (!g1083)) + ((!g4) & (g1080) & (g1081) & (!g1038) & (g1083)) + ((!g4) & (g1080) & (g1081) & (g1038) & (!g1083)) + ((!g4) & (g1080) & (g1081) & (g1038) & (g1083)) + ((g4) & (!g1080) & (g1081) & (!g1038) & (!g1083)) + ((g4) & (!g1080) & (g1081) & (!g1038) & (g1083)) + ((g4) & (!g1080) & (g1081) & (g1038) & (!g1083)) + ((g4) & (!g1080) & (g1081) & (g1038) & (g1083)) + ((g4) & (g1080) & (!g1081) & (!g1038) & (!g1083)) + ((g4) & (g1080) & (!g1081) & (g1038) & (!g1083)) + ((g4) & (g1080) & (!g1081) & (g1038) & (g1083)) + ((g4) & (g1080) & (g1081) & (!g1038) & (g1083)));
	assign g1096 = (((!g8) & (!g1041) & (g1079) & (!g1038) & (!g1083)) + ((!g8) & (!g1041) & (g1079) & (g1038) & (!g1083)) + ((!g8) & (!g1041) & (g1079) & (g1038) & (g1083)) + ((!g8) & (g1041) & (!g1079) & (!g1038) & (!g1083)) + ((!g8) & (g1041) & (!g1079) & (!g1038) & (g1083)) + ((!g8) & (g1041) & (!g1079) & (g1038) & (!g1083)) + ((!g8) & (g1041) & (!g1079) & (g1038) & (g1083)) + ((!g8) & (g1041) & (g1079) & (!g1038) & (g1083)) + ((g8) & (!g1041) & (!g1079) & (!g1038) & (!g1083)) + ((g8) & (!g1041) & (!g1079) & (g1038) & (!g1083)) + ((g8) & (!g1041) & (!g1079) & (g1038) & (g1083)) + ((g8) & (g1041) & (!g1079) & (!g1038) & (g1083)) + ((g8) & (g1041) & (g1079) & (!g1038) & (!g1083)) + ((g8) & (g1041) & (g1079) & (!g1038) & (g1083)) + ((g8) & (g1041) & (g1079) & (g1038) & (!g1083)) + ((g8) & (g1041) & (g1079) & (g1038) & (g1083)));
	assign g1097 = (((!g18) & (!g27) & (g1043) & (g1078)) + ((!g18) & (g27) & (!g1043) & (g1078)) + ((!g18) & (g27) & (g1043) & (!g1078)) + ((!g18) & (g27) & (g1043) & (g1078)) + ((g18) & (!g27) & (!g1043) & (!g1078)) + ((g18) & (!g27) & (!g1043) & (g1078)) + ((g18) & (!g27) & (g1043) & (!g1078)) + ((g18) & (g27) & (!g1043) & (!g1078)));
	assign g1098 = (((!g1042) & (!g1038) & (!g1083) & (g1097)) + ((!g1042) & (g1038) & (!g1083) & (g1097)) + ((!g1042) & (g1038) & (g1083) & (g1097)) + ((g1042) & (!g1038) & (!g1083) & (!g1097)) + ((g1042) & (!g1038) & (g1083) & (!g1097)) + ((g1042) & (!g1038) & (g1083) & (g1097)) + ((g1042) & (g1038) & (!g1083) & (!g1097)) + ((g1042) & (g1038) & (g1083) & (!g1097)));
	assign g1099 = (((!g27) & (!g1043) & (g1078) & (!g1038) & (!g1083)) + ((!g27) & (!g1043) & (g1078) & (g1038) & (!g1083)) + ((!g27) & (!g1043) & (g1078) & (g1038) & (g1083)) + ((!g27) & (g1043) & (!g1078) & (!g1038) & (!g1083)) + ((!g27) & (g1043) & (!g1078) & (!g1038) & (g1083)) + ((!g27) & (g1043) & (!g1078) & (g1038) & (!g1083)) + ((!g27) & (g1043) & (!g1078) & (g1038) & (g1083)) + ((!g27) & (g1043) & (g1078) & (!g1038) & (g1083)) + ((g27) & (!g1043) & (!g1078) & (!g1038) & (!g1083)) + ((g27) & (!g1043) & (!g1078) & (g1038) & (!g1083)) + ((g27) & (!g1043) & (!g1078) & (g1038) & (g1083)) + ((g27) & (g1043) & (!g1078) & (!g1038) & (g1083)) + ((g27) & (g1043) & (g1078) & (!g1038) & (!g1083)) + ((g27) & (g1043) & (g1078) & (!g1038) & (g1083)) + ((g27) & (g1043) & (g1078) & (g1038) & (!g1083)) + ((g27) & (g1043) & (g1078) & (g1038) & (g1083)));
	assign g1100 = (((!g39) & (!g54) & (g1045) & (g1077)) + ((!g39) & (g54) & (!g1045) & (g1077)) + ((!g39) & (g54) & (g1045) & (!g1077)) + ((!g39) & (g54) & (g1045) & (g1077)) + ((g39) & (!g54) & (!g1045) & (!g1077)) + ((g39) & (!g54) & (!g1045) & (g1077)) + ((g39) & (!g54) & (g1045) & (!g1077)) + ((g39) & (g54) & (!g1045) & (!g1077)));
	assign g1101 = (((!g1044) & (!g1038) & (!g1083) & (g1100)) + ((!g1044) & (g1038) & (!g1083) & (g1100)) + ((!g1044) & (g1038) & (g1083) & (g1100)) + ((g1044) & (!g1038) & (!g1083) & (!g1100)) + ((g1044) & (!g1038) & (g1083) & (!g1100)) + ((g1044) & (!g1038) & (g1083) & (g1100)) + ((g1044) & (g1038) & (!g1083) & (!g1100)) + ((g1044) & (g1038) & (g1083) & (!g1100)));
	assign g1102 = (((!g54) & (!g1045) & (g1077) & (!g1038) & (!g1083)) + ((!g54) & (!g1045) & (g1077) & (g1038) & (!g1083)) + ((!g54) & (!g1045) & (g1077) & (g1038) & (g1083)) + ((!g54) & (g1045) & (!g1077) & (!g1038) & (!g1083)) + ((!g54) & (g1045) & (!g1077) & (!g1038) & (g1083)) + ((!g54) & (g1045) & (!g1077) & (g1038) & (!g1083)) + ((!g54) & (g1045) & (!g1077) & (g1038) & (g1083)) + ((!g54) & (g1045) & (g1077) & (!g1038) & (g1083)) + ((g54) & (!g1045) & (!g1077) & (!g1038) & (!g1083)) + ((g54) & (!g1045) & (!g1077) & (g1038) & (!g1083)) + ((g54) & (!g1045) & (!g1077) & (g1038) & (g1083)) + ((g54) & (g1045) & (!g1077) & (!g1038) & (g1083)) + ((g54) & (g1045) & (g1077) & (!g1038) & (!g1083)) + ((g54) & (g1045) & (g1077) & (!g1038) & (g1083)) + ((g54) & (g1045) & (g1077) & (g1038) & (!g1083)) + ((g54) & (g1045) & (g1077) & (g1038) & (g1083)));
	assign g1103 = (((!g68) & (!g87) & (g1047) & (g1076)) + ((!g68) & (g87) & (!g1047) & (g1076)) + ((!g68) & (g87) & (g1047) & (!g1076)) + ((!g68) & (g87) & (g1047) & (g1076)) + ((g68) & (!g87) & (!g1047) & (!g1076)) + ((g68) & (!g87) & (!g1047) & (g1076)) + ((g68) & (!g87) & (g1047) & (!g1076)) + ((g68) & (g87) & (!g1047) & (!g1076)));
	assign g1104 = (((!g1046) & (!g1038) & (!g1083) & (g1103)) + ((!g1046) & (g1038) & (!g1083) & (g1103)) + ((!g1046) & (g1038) & (g1083) & (g1103)) + ((g1046) & (!g1038) & (!g1083) & (!g1103)) + ((g1046) & (!g1038) & (g1083) & (!g1103)) + ((g1046) & (!g1038) & (g1083) & (g1103)) + ((g1046) & (g1038) & (!g1083) & (!g1103)) + ((g1046) & (g1038) & (g1083) & (!g1103)));
	assign g1105 = (((!g87) & (!g1047) & (g1076) & (!g1038) & (!g1083)) + ((!g87) & (!g1047) & (g1076) & (g1038) & (!g1083)) + ((!g87) & (!g1047) & (g1076) & (g1038) & (g1083)) + ((!g87) & (g1047) & (!g1076) & (!g1038) & (!g1083)) + ((!g87) & (g1047) & (!g1076) & (!g1038) & (g1083)) + ((!g87) & (g1047) & (!g1076) & (g1038) & (!g1083)) + ((!g87) & (g1047) & (!g1076) & (g1038) & (g1083)) + ((!g87) & (g1047) & (g1076) & (!g1038) & (g1083)) + ((g87) & (!g1047) & (!g1076) & (!g1038) & (!g1083)) + ((g87) & (!g1047) & (!g1076) & (g1038) & (!g1083)) + ((g87) & (!g1047) & (!g1076) & (g1038) & (g1083)) + ((g87) & (g1047) & (!g1076) & (!g1038) & (g1083)) + ((g87) & (g1047) & (g1076) & (!g1038) & (!g1083)) + ((g87) & (g1047) & (g1076) & (!g1038) & (g1083)) + ((g87) & (g1047) & (g1076) & (g1038) & (!g1083)) + ((g87) & (g1047) & (g1076) & (g1038) & (g1083)));
	assign g1106 = (((!g104) & (!g127) & (g1049) & (g1075)) + ((!g104) & (g127) & (!g1049) & (g1075)) + ((!g104) & (g127) & (g1049) & (!g1075)) + ((!g104) & (g127) & (g1049) & (g1075)) + ((g104) & (!g127) & (!g1049) & (!g1075)) + ((g104) & (!g127) & (!g1049) & (g1075)) + ((g104) & (!g127) & (g1049) & (!g1075)) + ((g104) & (g127) & (!g1049) & (!g1075)));
	assign g1107 = (((!g1048) & (!g1038) & (!g1083) & (g1106)) + ((!g1048) & (g1038) & (!g1083) & (g1106)) + ((!g1048) & (g1038) & (g1083) & (g1106)) + ((g1048) & (!g1038) & (!g1083) & (!g1106)) + ((g1048) & (!g1038) & (g1083) & (!g1106)) + ((g1048) & (!g1038) & (g1083) & (g1106)) + ((g1048) & (g1038) & (!g1083) & (!g1106)) + ((g1048) & (g1038) & (g1083) & (!g1106)));
	assign g1108 = (((!g127) & (!g1049) & (g1075) & (!g1038) & (!g1083)) + ((!g127) & (!g1049) & (g1075) & (g1038) & (!g1083)) + ((!g127) & (!g1049) & (g1075) & (g1038) & (g1083)) + ((!g127) & (g1049) & (!g1075) & (!g1038) & (!g1083)) + ((!g127) & (g1049) & (!g1075) & (!g1038) & (g1083)) + ((!g127) & (g1049) & (!g1075) & (g1038) & (!g1083)) + ((!g127) & (g1049) & (!g1075) & (g1038) & (g1083)) + ((!g127) & (g1049) & (g1075) & (!g1038) & (g1083)) + ((g127) & (!g1049) & (!g1075) & (!g1038) & (!g1083)) + ((g127) & (!g1049) & (!g1075) & (g1038) & (!g1083)) + ((g127) & (!g1049) & (!g1075) & (g1038) & (g1083)) + ((g127) & (g1049) & (!g1075) & (!g1038) & (g1083)) + ((g127) & (g1049) & (g1075) & (!g1038) & (!g1083)) + ((g127) & (g1049) & (g1075) & (!g1038) & (g1083)) + ((g127) & (g1049) & (g1075) & (g1038) & (!g1083)) + ((g127) & (g1049) & (g1075) & (g1038) & (g1083)));
	assign g1109 = (((!g147) & (!g174) & (g1051) & (g1074)) + ((!g147) & (g174) & (!g1051) & (g1074)) + ((!g147) & (g174) & (g1051) & (!g1074)) + ((!g147) & (g174) & (g1051) & (g1074)) + ((g147) & (!g174) & (!g1051) & (!g1074)) + ((g147) & (!g174) & (!g1051) & (g1074)) + ((g147) & (!g174) & (g1051) & (!g1074)) + ((g147) & (g174) & (!g1051) & (!g1074)));
	assign g1110 = (((!g1050) & (!g1038) & (!g1083) & (g1109)) + ((!g1050) & (g1038) & (!g1083) & (g1109)) + ((!g1050) & (g1038) & (g1083) & (g1109)) + ((g1050) & (!g1038) & (!g1083) & (!g1109)) + ((g1050) & (!g1038) & (g1083) & (!g1109)) + ((g1050) & (!g1038) & (g1083) & (g1109)) + ((g1050) & (g1038) & (!g1083) & (!g1109)) + ((g1050) & (g1038) & (g1083) & (!g1109)));
	assign g1111 = (((!g174) & (!g1051) & (g1074) & (!g1038) & (!g1083)) + ((!g174) & (!g1051) & (g1074) & (g1038) & (!g1083)) + ((!g174) & (!g1051) & (g1074) & (g1038) & (g1083)) + ((!g174) & (g1051) & (!g1074) & (!g1038) & (!g1083)) + ((!g174) & (g1051) & (!g1074) & (!g1038) & (g1083)) + ((!g174) & (g1051) & (!g1074) & (g1038) & (!g1083)) + ((!g174) & (g1051) & (!g1074) & (g1038) & (g1083)) + ((!g174) & (g1051) & (g1074) & (!g1038) & (g1083)) + ((g174) & (!g1051) & (!g1074) & (!g1038) & (!g1083)) + ((g174) & (!g1051) & (!g1074) & (g1038) & (!g1083)) + ((g174) & (!g1051) & (!g1074) & (g1038) & (g1083)) + ((g174) & (g1051) & (!g1074) & (!g1038) & (g1083)) + ((g174) & (g1051) & (g1074) & (!g1038) & (!g1083)) + ((g174) & (g1051) & (g1074) & (!g1038) & (g1083)) + ((g174) & (g1051) & (g1074) & (g1038) & (!g1083)) + ((g174) & (g1051) & (g1074) & (g1038) & (g1083)));
	assign g1112 = (((!g198) & (!g229) & (g1053) & (g1073)) + ((!g198) & (g229) & (!g1053) & (g1073)) + ((!g198) & (g229) & (g1053) & (!g1073)) + ((!g198) & (g229) & (g1053) & (g1073)) + ((g198) & (!g229) & (!g1053) & (!g1073)) + ((g198) & (!g229) & (!g1053) & (g1073)) + ((g198) & (!g229) & (g1053) & (!g1073)) + ((g198) & (g229) & (!g1053) & (!g1073)));
	assign g1113 = (((!g1052) & (!g1038) & (!g1083) & (g1112)) + ((!g1052) & (g1038) & (!g1083) & (g1112)) + ((!g1052) & (g1038) & (g1083) & (g1112)) + ((g1052) & (!g1038) & (!g1083) & (!g1112)) + ((g1052) & (!g1038) & (g1083) & (!g1112)) + ((g1052) & (!g1038) & (g1083) & (g1112)) + ((g1052) & (g1038) & (!g1083) & (!g1112)) + ((g1052) & (g1038) & (g1083) & (!g1112)));
	assign g1114 = (((!g229) & (!g1053) & (g1073) & (!g1038) & (!g1083)) + ((!g229) & (!g1053) & (g1073) & (g1038) & (!g1083)) + ((!g229) & (!g1053) & (g1073) & (g1038) & (g1083)) + ((!g229) & (g1053) & (!g1073) & (!g1038) & (!g1083)) + ((!g229) & (g1053) & (!g1073) & (!g1038) & (g1083)) + ((!g229) & (g1053) & (!g1073) & (g1038) & (!g1083)) + ((!g229) & (g1053) & (!g1073) & (g1038) & (g1083)) + ((!g229) & (g1053) & (g1073) & (!g1038) & (g1083)) + ((g229) & (!g1053) & (!g1073) & (!g1038) & (!g1083)) + ((g229) & (!g1053) & (!g1073) & (g1038) & (!g1083)) + ((g229) & (!g1053) & (!g1073) & (g1038) & (g1083)) + ((g229) & (g1053) & (!g1073) & (!g1038) & (g1083)) + ((g229) & (g1053) & (g1073) & (!g1038) & (!g1083)) + ((g229) & (g1053) & (g1073) & (!g1038) & (g1083)) + ((g229) & (g1053) & (g1073) & (g1038) & (!g1083)) + ((g229) & (g1053) & (g1073) & (g1038) & (g1083)));
	assign g1115 = (((!g255) & (!g290) & (g1055) & (g1072)) + ((!g255) & (g290) & (!g1055) & (g1072)) + ((!g255) & (g290) & (g1055) & (!g1072)) + ((!g255) & (g290) & (g1055) & (g1072)) + ((g255) & (!g290) & (!g1055) & (!g1072)) + ((g255) & (!g290) & (!g1055) & (g1072)) + ((g255) & (!g290) & (g1055) & (!g1072)) + ((g255) & (g290) & (!g1055) & (!g1072)));
	assign g1116 = (((!g1054) & (!g1038) & (!g1083) & (g1115)) + ((!g1054) & (g1038) & (!g1083) & (g1115)) + ((!g1054) & (g1038) & (g1083) & (g1115)) + ((g1054) & (!g1038) & (!g1083) & (!g1115)) + ((g1054) & (!g1038) & (g1083) & (!g1115)) + ((g1054) & (!g1038) & (g1083) & (g1115)) + ((g1054) & (g1038) & (!g1083) & (!g1115)) + ((g1054) & (g1038) & (g1083) & (!g1115)));
	assign g1117 = (((!g290) & (!g1055) & (g1072) & (!g1038) & (!g1083)) + ((!g290) & (!g1055) & (g1072) & (g1038) & (!g1083)) + ((!g290) & (!g1055) & (g1072) & (g1038) & (g1083)) + ((!g290) & (g1055) & (!g1072) & (!g1038) & (!g1083)) + ((!g290) & (g1055) & (!g1072) & (!g1038) & (g1083)) + ((!g290) & (g1055) & (!g1072) & (g1038) & (!g1083)) + ((!g290) & (g1055) & (!g1072) & (g1038) & (g1083)) + ((!g290) & (g1055) & (g1072) & (!g1038) & (g1083)) + ((g290) & (!g1055) & (!g1072) & (!g1038) & (!g1083)) + ((g290) & (!g1055) & (!g1072) & (g1038) & (!g1083)) + ((g290) & (!g1055) & (!g1072) & (g1038) & (g1083)) + ((g290) & (g1055) & (!g1072) & (!g1038) & (g1083)) + ((g290) & (g1055) & (g1072) & (!g1038) & (!g1083)) + ((g290) & (g1055) & (g1072) & (!g1038) & (g1083)) + ((g290) & (g1055) & (g1072) & (g1038) & (!g1083)) + ((g290) & (g1055) & (g1072) & (g1038) & (g1083)));
	assign g1118 = (((!g319) & (!g358) & (g1057) & (g1071)) + ((!g319) & (g358) & (!g1057) & (g1071)) + ((!g319) & (g358) & (g1057) & (!g1071)) + ((!g319) & (g358) & (g1057) & (g1071)) + ((g319) & (!g358) & (!g1057) & (!g1071)) + ((g319) & (!g358) & (!g1057) & (g1071)) + ((g319) & (!g358) & (g1057) & (!g1071)) + ((g319) & (g358) & (!g1057) & (!g1071)));
	assign g1119 = (((!g1056) & (!g1038) & (!g1083) & (g1118)) + ((!g1056) & (g1038) & (!g1083) & (g1118)) + ((!g1056) & (g1038) & (g1083) & (g1118)) + ((g1056) & (!g1038) & (!g1083) & (!g1118)) + ((g1056) & (!g1038) & (g1083) & (!g1118)) + ((g1056) & (!g1038) & (g1083) & (g1118)) + ((g1056) & (g1038) & (!g1083) & (!g1118)) + ((g1056) & (g1038) & (g1083) & (!g1118)));
	assign g1120 = (((!g358) & (!g1057) & (g1071) & (!g1038) & (!g1083)) + ((!g358) & (!g1057) & (g1071) & (g1038) & (!g1083)) + ((!g358) & (!g1057) & (g1071) & (g1038) & (g1083)) + ((!g358) & (g1057) & (!g1071) & (!g1038) & (!g1083)) + ((!g358) & (g1057) & (!g1071) & (!g1038) & (g1083)) + ((!g358) & (g1057) & (!g1071) & (g1038) & (!g1083)) + ((!g358) & (g1057) & (!g1071) & (g1038) & (g1083)) + ((!g358) & (g1057) & (g1071) & (!g1038) & (g1083)) + ((g358) & (!g1057) & (!g1071) & (!g1038) & (!g1083)) + ((g358) & (!g1057) & (!g1071) & (g1038) & (!g1083)) + ((g358) & (!g1057) & (!g1071) & (g1038) & (g1083)) + ((g358) & (g1057) & (!g1071) & (!g1038) & (g1083)) + ((g358) & (g1057) & (g1071) & (!g1038) & (!g1083)) + ((g358) & (g1057) & (g1071) & (!g1038) & (g1083)) + ((g358) & (g1057) & (g1071) & (g1038) & (!g1083)) + ((g358) & (g1057) & (g1071) & (g1038) & (g1083)));
	assign g1121 = (((!g390) & (!g433) & (g1059) & (g1070)) + ((!g390) & (g433) & (!g1059) & (g1070)) + ((!g390) & (g433) & (g1059) & (!g1070)) + ((!g390) & (g433) & (g1059) & (g1070)) + ((g390) & (!g433) & (!g1059) & (!g1070)) + ((g390) & (!g433) & (!g1059) & (g1070)) + ((g390) & (!g433) & (g1059) & (!g1070)) + ((g390) & (g433) & (!g1059) & (!g1070)));
	assign g1122 = (((!g1058) & (!g1038) & (!g1083) & (g1121)) + ((!g1058) & (g1038) & (!g1083) & (g1121)) + ((!g1058) & (g1038) & (g1083) & (g1121)) + ((g1058) & (!g1038) & (!g1083) & (!g1121)) + ((g1058) & (!g1038) & (g1083) & (!g1121)) + ((g1058) & (!g1038) & (g1083) & (g1121)) + ((g1058) & (g1038) & (!g1083) & (!g1121)) + ((g1058) & (g1038) & (g1083) & (!g1121)));
	assign g1123 = (((!g433) & (!g1059) & (g1070) & (!g1038) & (!g1083)) + ((!g433) & (!g1059) & (g1070) & (g1038) & (!g1083)) + ((!g433) & (!g1059) & (g1070) & (g1038) & (g1083)) + ((!g433) & (g1059) & (!g1070) & (!g1038) & (!g1083)) + ((!g433) & (g1059) & (!g1070) & (!g1038) & (g1083)) + ((!g433) & (g1059) & (!g1070) & (g1038) & (!g1083)) + ((!g433) & (g1059) & (!g1070) & (g1038) & (g1083)) + ((!g433) & (g1059) & (g1070) & (!g1038) & (g1083)) + ((g433) & (!g1059) & (!g1070) & (!g1038) & (!g1083)) + ((g433) & (!g1059) & (!g1070) & (g1038) & (!g1083)) + ((g433) & (!g1059) & (!g1070) & (g1038) & (g1083)) + ((g433) & (g1059) & (!g1070) & (!g1038) & (g1083)) + ((g433) & (g1059) & (g1070) & (!g1038) & (!g1083)) + ((g433) & (g1059) & (g1070) & (!g1038) & (g1083)) + ((g433) & (g1059) & (g1070) & (g1038) & (!g1083)) + ((g433) & (g1059) & (g1070) & (g1038) & (g1083)));
	assign g1124 = (((!g468) & (!g515) & (g1061) & (g1069)) + ((!g468) & (g515) & (!g1061) & (g1069)) + ((!g468) & (g515) & (g1061) & (!g1069)) + ((!g468) & (g515) & (g1061) & (g1069)) + ((g468) & (!g515) & (!g1061) & (!g1069)) + ((g468) & (!g515) & (!g1061) & (g1069)) + ((g468) & (!g515) & (g1061) & (!g1069)) + ((g468) & (g515) & (!g1061) & (!g1069)));
	assign g1125 = (((!g1060) & (!g1038) & (!g1083) & (g1124)) + ((!g1060) & (g1038) & (!g1083) & (g1124)) + ((!g1060) & (g1038) & (g1083) & (g1124)) + ((g1060) & (!g1038) & (!g1083) & (!g1124)) + ((g1060) & (!g1038) & (g1083) & (!g1124)) + ((g1060) & (!g1038) & (g1083) & (g1124)) + ((g1060) & (g1038) & (!g1083) & (!g1124)) + ((g1060) & (g1038) & (g1083) & (!g1124)));
	assign g1126 = (((!g515) & (!g1061) & (g1069) & (!g1038) & (!g1083)) + ((!g515) & (!g1061) & (g1069) & (g1038) & (!g1083)) + ((!g515) & (!g1061) & (g1069) & (g1038) & (g1083)) + ((!g515) & (g1061) & (!g1069) & (!g1038) & (!g1083)) + ((!g515) & (g1061) & (!g1069) & (!g1038) & (g1083)) + ((!g515) & (g1061) & (!g1069) & (g1038) & (!g1083)) + ((!g515) & (g1061) & (!g1069) & (g1038) & (g1083)) + ((!g515) & (g1061) & (g1069) & (!g1038) & (g1083)) + ((g515) & (!g1061) & (!g1069) & (!g1038) & (!g1083)) + ((g515) & (!g1061) & (!g1069) & (g1038) & (!g1083)) + ((g515) & (!g1061) & (!g1069) & (g1038) & (g1083)) + ((g515) & (g1061) & (!g1069) & (!g1038) & (g1083)) + ((g515) & (g1061) & (g1069) & (!g1038) & (!g1083)) + ((g515) & (g1061) & (g1069) & (!g1038) & (g1083)) + ((g515) & (g1061) & (g1069) & (g1038) & (!g1083)) + ((g515) & (g1061) & (g1069) & (g1038) & (g1083)));
	assign g1127 = (((!g553) & (!g604) & (g1063) & (g1068)) + ((!g553) & (g604) & (!g1063) & (g1068)) + ((!g553) & (g604) & (g1063) & (!g1068)) + ((!g553) & (g604) & (g1063) & (g1068)) + ((g553) & (!g604) & (!g1063) & (!g1068)) + ((g553) & (!g604) & (!g1063) & (g1068)) + ((g553) & (!g604) & (g1063) & (!g1068)) + ((g553) & (g604) & (!g1063) & (!g1068)));
	assign g1128 = (((!g1062) & (!g1038) & (!g1083) & (g1127)) + ((!g1062) & (g1038) & (!g1083) & (g1127)) + ((!g1062) & (g1038) & (g1083) & (g1127)) + ((g1062) & (!g1038) & (!g1083) & (!g1127)) + ((g1062) & (!g1038) & (g1083) & (!g1127)) + ((g1062) & (!g1038) & (g1083) & (g1127)) + ((g1062) & (g1038) & (!g1083) & (!g1127)) + ((g1062) & (g1038) & (g1083) & (!g1127)));
	assign g1129 = (((!g604) & (!g1063) & (g1068) & (!g1038) & (!g1083)) + ((!g604) & (!g1063) & (g1068) & (g1038) & (!g1083)) + ((!g604) & (!g1063) & (g1068) & (g1038) & (g1083)) + ((!g604) & (g1063) & (!g1068) & (!g1038) & (!g1083)) + ((!g604) & (g1063) & (!g1068) & (!g1038) & (g1083)) + ((!g604) & (g1063) & (!g1068) & (g1038) & (!g1083)) + ((!g604) & (g1063) & (!g1068) & (g1038) & (g1083)) + ((!g604) & (g1063) & (g1068) & (!g1038) & (g1083)) + ((g604) & (!g1063) & (!g1068) & (!g1038) & (!g1083)) + ((g604) & (!g1063) & (!g1068) & (g1038) & (!g1083)) + ((g604) & (!g1063) & (!g1068) & (g1038) & (g1083)) + ((g604) & (g1063) & (!g1068) & (!g1038) & (g1083)) + ((g604) & (g1063) & (g1068) & (!g1038) & (!g1083)) + ((g604) & (g1063) & (g1068) & (!g1038) & (g1083)) + ((g604) & (g1063) & (g1068) & (g1038) & (!g1083)) + ((g604) & (g1063) & (g1068) & (g1038) & (g1083)));
	assign g1130 = (((!g645) & (!g700) & (g1065) & (g1067)) + ((!g645) & (g700) & (!g1065) & (g1067)) + ((!g645) & (g700) & (g1065) & (!g1067)) + ((!g645) & (g700) & (g1065) & (g1067)) + ((g645) & (!g700) & (!g1065) & (!g1067)) + ((g645) & (!g700) & (!g1065) & (g1067)) + ((g645) & (!g700) & (g1065) & (!g1067)) + ((g645) & (g700) & (!g1065) & (!g1067)));
	assign g1131 = (((!g1064) & (!g1038) & (!g1083) & (g1130)) + ((!g1064) & (g1038) & (!g1083) & (g1130)) + ((!g1064) & (g1038) & (g1083) & (g1130)) + ((g1064) & (!g1038) & (!g1083) & (!g1130)) + ((g1064) & (!g1038) & (g1083) & (!g1130)) + ((g1064) & (!g1038) & (g1083) & (g1130)) + ((g1064) & (g1038) & (!g1083) & (!g1130)) + ((g1064) & (g1038) & (g1083) & (!g1130)));
	assign g1132 = (((!g700) & (!g1065) & (g1067) & (!g1038) & (!g1083)) + ((!g700) & (!g1065) & (g1067) & (g1038) & (!g1083)) + ((!g700) & (!g1065) & (g1067) & (g1038) & (g1083)) + ((!g700) & (g1065) & (!g1067) & (!g1038) & (!g1083)) + ((!g700) & (g1065) & (!g1067) & (!g1038) & (g1083)) + ((!g700) & (g1065) & (!g1067) & (g1038) & (!g1083)) + ((!g700) & (g1065) & (!g1067) & (g1038) & (g1083)) + ((!g700) & (g1065) & (g1067) & (!g1038) & (g1083)) + ((g700) & (!g1065) & (!g1067) & (!g1038) & (!g1083)) + ((g700) & (!g1065) & (!g1067) & (g1038) & (!g1083)) + ((g700) & (!g1065) & (!g1067) & (g1038) & (g1083)) + ((g700) & (g1065) & (!g1067) & (!g1038) & (g1083)) + ((g700) & (g1065) & (g1067) & (!g1038) & (!g1083)) + ((g700) & (g1065) & (g1067) & (!g1038) & (g1083)) + ((g700) & (g1065) & (g1067) & (g1038) & (!g1083)) + ((g700) & (g1065) & (g1067) & (g1038) & (g1083)));
	assign g1133 = (((!g744) & (!g803) & (g1031) & (g1037)) + ((!g744) & (g803) & (!g1031) & (g1037)) + ((!g744) & (g803) & (g1031) & (!g1037)) + ((!g744) & (g803) & (g1031) & (g1037)) + ((g744) & (!g803) & (!g1031) & (!g1037)) + ((g744) & (!g803) & (!g1031) & (g1037)) + ((g744) & (!g803) & (g1031) & (!g1037)) + ((g744) & (g803) & (!g1031) & (!g1037)));
	assign g1134 = (((!g1066) & (!g1038) & (!g1083) & (g1133)) + ((!g1066) & (g1038) & (!g1083) & (g1133)) + ((!g1066) & (g1038) & (g1083) & (g1133)) + ((g1066) & (!g1038) & (!g1083) & (!g1133)) + ((g1066) & (!g1038) & (g1083) & (!g1133)) + ((g1066) & (!g1038) & (g1083) & (g1133)) + ((g1066) & (g1038) & (!g1083) & (!g1133)) + ((g1066) & (g1038) & (g1083) & (!g1133)));
	assign g1135 = (((!g700) & (!g744) & (g1134) & (g1084) & (g1094)) + ((!g700) & (g744) & (g1134) & (!g1084) & (g1094)) + ((!g700) & (g744) & (g1134) & (g1084) & (!g1094)) + ((!g700) & (g744) & (g1134) & (g1084) & (g1094)) + ((g700) & (!g744) & (!g1134) & (g1084) & (g1094)) + ((g700) & (!g744) & (g1134) & (!g1084) & (!g1094)) + ((g700) & (!g744) & (g1134) & (!g1084) & (g1094)) + ((g700) & (!g744) & (g1134) & (g1084) & (!g1094)) + ((g700) & (!g744) & (g1134) & (g1084) & (g1094)) + ((g700) & (g744) & (!g1134) & (!g1084) & (g1094)) + ((g700) & (g744) & (!g1134) & (g1084) & (!g1094)) + ((g700) & (g744) & (!g1134) & (g1084) & (g1094)) + ((g700) & (g744) & (g1134) & (!g1084) & (!g1094)) + ((g700) & (g744) & (g1134) & (!g1084) & (g1094)) + ((g700) & (g744) & (g1134) & (g1084) & (!g1094)) + ((g700) & (g744) & (g1134) & (g1084) & (g1094)));
	assign g1136 = (((!g604) & (!g645) & (g1131) & (g1132) & (g1135)) + ((!g604) & (g645) & (g1131) & (!g1132) & (g1135)) + ((!g604) & (g645) & (g1131) & (g1132) & (!g1135)) + ((!g604) & (g645) & (g1131) & (g1132) & (g1135)) + ((g604) & (!g645) & (!g1131) & (g1132) & (g1135)) + ((g604) & (!g645) & (g1131) & (!g1132) & (!g1135)) + ((g604) & (!g645) & (g1131) & (!g1132) & (g1135)) + ((g604) & (!g645) & (g1131) & (g1132) & (!g1135)) + ((g604) & (!g645) & (g1131) & (g1132) & (g1135)) + ((g604) & (g645) & (!g1131) & (!g1132) & (g1135)) + ((g604) & (g645) & (!g1131) & (g1132) & (!g1135)) + ((g604) & (g645) & (!g1131) & (g1132) & (g1135)) + ((g604) & (g645) & (g1131) & (!g1132) & (!g1135)) + ((g604) & (g645) & (g1131) & (!g1132) & (g1135)) + ((g604) & (g645) & (g1131) & (g1132) & (!g1135)) + ((g604) & (g645) & (g1131) & (g1132) & (g1135)));
	assign g1137 = (((!g515) & (!g553) & (g1128) & (g1129) & (g1136)) + ((!g515) & (g553) & (g1128) & (!g1129) & (g1136)) + ((!g515) & (g553) & (g1128) & (g1129) & (!g1136)) + ((!g515) & (g553) & (g1128) & (g1129) & (g1136)) + ((g515) & (!g553) & (!g1128) & (g1129) & (g1136)) + ((g515) & (!g553) & (g1128) & (!g1129) & (!g1136)) + ((g515) & (!g553) & (g1128) & (!g1129) & (g1136)) + ((g515) & (!g553) & (g1128) & (g1129) & (!g1136)) + ((g515) & (!g553) & (g1128) & (g1129) & (g1136)) + ((g515) & (g553) & (!g1128) & (!g1129) & (g1136)) + ((g515) & (g553) & (!g1128) & (g1129) & (!g1136)) + ((g515) & (g553) & (!g1128) & (g1129) & (g1136)) + ((g515) & (g553) & (g1128) & (!g1129) & (!g1136)) + ((g515) & (g553) & (g1128) & (!g1129) & (g1136)) + ((g515) & (g553) & (g1128) & (g1129) & (!g1136)) + ((g515) & (g553) & (g1128) & (g1129) & (g1136)));
	assign g1138 = (((!g433) & (!g468) & (g1125) & (g1126) & (g1137)) + ((!g433) & (g468) & (g1125) & (!g1126) & (g1137)) + ((!g433) & (g468) & (g1125) & (g1126) & (!g1137)) + ((!g433) & (g468) & (g1125) & (g1126) & (g1137)) + ((g433) & (!g468) & (!g1125) & (g1126) & (g1137)) + ((g433) & (!g468) & (g1125) & (!g1126) & (!g1137)) + ((g433) & (!g468) & (g1125) & (!g1126) & (g1137)) + ((g433) & (!g468) & (g1125) & (g1126) & (!g1137)) + ((g433) & (!g468) & (g1125) & (g1126) & (g1137)) + ((g433) & (g468) & (!g1125) & (!g1126) & (g1137)) + ((g433) & (g468) & (!g1125) & (g1126) & (!g1137)) + ((g433) & (g468) & (!g1125) & (g1126) & (g1137)) + ((g433) & (g468) & (g1125) & (!g1126) & (!g1137)) + ((g433) & (g468) & (g1125) & (!g1126) & (g1137)) + ((g433) & (g468) & (g1125) & (g1126) & (!g1137)) + ((g433) & (g468) & (g1125) & (g1126) & (g1137)));
	assign g1139 = (((!g358) & (!g390) & (g1122) & (g1123) & (g1138)) + ((!g358) & (g390) & (g1122) & (!g1123) & (g1138)) + ((!g358) & (g390) & (g1122) & (g1123) & (!g1138)) + ((!g358) & (g390) & (g1122) & (g1123) & (g1138)) + ((g358) & (!g390) & (!g1122) & (g1123) & (g1138)) + ((g358) & (!g390) & (g1122) & (!g1123) & (!g1138)) + ((g358) & (!g390) & (g1122) & (!g1123) & (g1138)) + ((g358) & (!g390) & (g1122) & (g1123) & (!g1138)) + ((g358) & (!g390) & (g1122) & (g1123) & (g1138)) + ((g358) & (g390) & (!g1122) & (!g1123) & (g1138)) + ((g358) & (g390) & (!g1122) & (g1123) & (!g1138)) + ((g358) & (g390) & (!g1122) & (g1123) & (g1138)) + ((g358) & (g390) & (g1122) & (!g1123) & (!g1138)) + ((g358) & (g390) & (g1122) & (!g1123) & (g1138)) + ((g358) & (g390) & (g1122) & (g1123) & (!g1138)) + ((g358) & (g390) & (g1122) & (g1123) & (g1138)));
	assign g1140 = (((!g290) & (!g319) & (g1119) & (g1120) & (g1139)) + ((!g290) & (g319) & (g1119) & (!g1120) & (g1139)) + ((!g290) & (g319) & (g1119) & (g1120) & (!g1139)) + ((!g290) & (g319) & (g1119) & (g1120) & (g1139)) + ((g290) & (!g319) & (!g1119) & (g1120) & (g1139)) + ((g290) & (!g319) & (g1119) & (!g1120) & (!g1139)) + ((g290) & (!g319) & (g1119) & (!g1120) & (g1139)) + ((g290) & (!g319) & (g1119) & (g1120) & (!g1139)) + ((g290) & (!g319) & (g1119) & (g1120) & (g1139)) + ((g290) & (g319) & (!g1119) & (!g1120) & (g1139)) + ((g290) & (g319) & (!g1119) & (g1120) & (!g1139)) + ((g290) & (g319) & (!g1119) & (g1120) & (g1139)) + ((g290) & (g319) & (g1119) & (!g1120) & (!g1139)) + ((g290) & (g319) & (g1119) & (!g1120) & (g1139)) + ((g290) & (g319) & (g1119) & (g1120) & (!g1139)) + ((g290) & (g319) & (g1119) & (g1120) & (g1139)));
	assign g1141 = (((!g229) & (!g255) & (g1116) & (g1117) & (g1140)) + ((!g229) & (g255) & (g1116) & (!g1117) & (g1140)) + ((!g229) & (g255) & (g1116) & (g1117) & (!g1140)) + ((!g229) & (g255) & (g1116) & (g1117) & (g1140)) + ((g229) & (!g255) & (!g1116) & (g1117) & (g1140)) + ((g229) & (!g255) & (g1116) & (!g1117) & (!g1140)) + ((g229) & (!g255) & (g1116) & (!g1117) & (g1140)) + ((g229) & (!g255) & (g1116) & (g1117) & (!g1140)) + ((g229) & (!g255) & (g1116) & (g1117) & (g1140)) + ((g229) & (g255) & (!g1116) & (!g1117) & (g1140)) + ((g229) & (g255) & (!g1116) & (g1117) & (!g1140)) + ((g229) & (g255) & (!g1116) & (g1117) & (g1140)) + ((g229) & (g255) & (g1116) & (!g1117) & (!g1140)) + ((g229) & (g255) & (g1116) & (!g1117) & (g1140)) + ((g229) & (g255) & (g1116) & (g1117) & (!g1140)) + ((g229) & (g255) & (g1116) & (g1117) & (g1140)));
	assign g1142 = (((!g174) & (!g198) & (g1113) & (g1114) & (g1141)) + ((!g174) & (g198) & (g1113) & (!g1114) & (g1141)) + ((!g174) & (g198) & (g1113) & (g1114) & (!g1141)) + ((!g174) & (g198) & (g1113) & (g1114) & (g1141)) + ((g174) & (!g198) & (!g1113) & (g1114) & (g1141)) + ((g174) & (!g198) & (g1113) & (!g1114) & (!g1141)) + ((g174) & (!g198) & (g1113) & (!g1114) & (g1141)) + ((g174) & (!g198) & (g1113) & (g1114) & (!g1141)) + ((g174) & (!g198) & (g1113) & (g1114) & (g1141)) + ((g174) & (g198) & (!g1113) & (!g1114) & (g1141)) + ((g174) & (g198) & (!g1113) & (g1114) & (!g1141)) + ((g174) & (g198) & (!g1113) & (g1114) & (g1141)) + ((g174) & (g198) & (g1113) & (!g1114) & (!g1141)) + ((g174) & (g198) & (g1113) & (!g1114) & (g1141)) + ((g174) & (g198) & (g1113) & (g1114) & (!g1141)) + ((g174) & (g198) & (g1113) & (g1114) & (g1141)));
	assign g1143 = (((!g127) & (!g147) & (g1110) & (g1111) & (g1142)) + ((!g127) & (g147) & (g1110) & (!g1111) & (g1142)) + ((!g127) & (g147) & (g1110) & (g1111) & (!g1142)) + ((!g127) & (g147) & (g1110) & (g1111) & (g1142)) + ((g127) & (!g147) & (!g1110) & (g1111) & (g1142)) + ((g127) & (!g147) & (g1110) & (!g1111) & (!g1142)) + ((g127) & (!g147) & (g1110) & (!g1111) & (g1142)) + ((g127) & (!g147) & (g1110) & (g1111) & (!g1142)) + ((g127) & (!g147) & (g1110) & (g1111) & (g1142)) + ((g127) & (g147) & (!g1110) & (!g1111) & (g1142)) + ((g127) & (g147) & (!g1110) & (g1111) & (!g1142)) + ((g127) & (g147) & (!g1110) & (g1111) & (g1142)) + ((g127) & (g147) & (g1110) & (!g1111) & (!g1142)) + ((g127) & (g147) & (g1110) & (!g1111) & (g1142)) + ((g127) & (g147) & (g1110) & (g1111) & (!g1142)) + ((g127) & (g147) & (g1110) & (g1111) & (g1142)));
	assign g1144 = (((!g87) & (!g104) & (g1107) & (g1108) & (g1143)) + ((!g87) & (g104) & (g1107) & (!g1108) & (g1143)) + ((!g87) & (g104) & (g1107) & (g1108) & (!g1143)) + ((!g87) & (g104) & (g1107) & (g1108) & (g1143)) + ((g87) & (!g104) & (!g1107) & (g1108) & (g1143)) + ((g87) & (!g104) & (g1107) & (!g1108) & (!g1143)) + ((g87) & (!g104) & (g1107) & (!g1108) & (g1143)) + ((g87) & (!g104) & (g1107) & (g1108) & (!g1143)) + ((g87) & (!g104) & (g1107) & (g1108) & (g1143)) + ((g87) & (g104) & (!g1107) & (!g1108) & (g1143)) + ((g87) & (g104) & (!g1107) & (g1108) & (!g1143)) + ((g87) & (g104) & (!g1107) & (g1108) & (g1143)) + ((g87) & (g104) & (g1107) & (!g1108) & (!g1143)) + ((g87) & (g104) & (g1107) & (!g1108) & (g1143)) + ((g87) & (g104) & (g1107) & (g1108) & (!g1143)) + ((g87) & (g104) & (g1107) & (g1108) & (g1143)));
	assign g1145 = (((!g54) & (!g68) & (g1104) & (g1105) & (g1144)) + ((!g54) & (g68) & (g1104) & (!g1105) & (g1144)) + ((!g54) & (g68) & (g1104) & (g1105) & (!g1144)) + ((!g54) & (g68) & (g1104) & (g1105) & (g1144)) + ((g54) & (!g68) & (!g1104) & (g1105) & (g1144)) + ((g54) & (!g68) & (g1104) & (!g1105) & (!g1144)) + ((g54) & (!g68) & (g1104) & (!g1105) & (g1144)) + ((g54) & (!g68) & (g1104) & (g1105) & (!g1144)) + ((g54) & (!g68) & (g1104) & (g1105) & (g1144)) + ((g54) & (g68) & (!g1104) & (!g1105) & (g1144)) + ((g54) & (g68) & (!g1104) & (g1105) & (!g1144)) + ((g54) & (g68) & (!g1104) & (g1105) & (g1144)) + ((g54) & (g68) & (g1104) & (!g1105) & (!g1144)) + ((g54) & (g68) & (g1104) & (!g1105) & (g1144)) + ((g54) & (g68) & (g1104) & (g1105) & (!g1144)) + ((g54) & (g68) & (g1104) & (g1105) & (g1144)));
	assign g1146 = (((!g27) & (!g39) & (g1101) & (g1102) & (g1145)) + ((!g27) & (g39) & (g1101) & (!g1102) & (g1145)) + ((!g27) & (g39) & (g1101) & (g1102) & (!g1145)) + ((!g27) & (g39) & (g1101) & (g1102) & (g1145)) + ((g27) & (!g39) & (!g1101) & (g1102) & (g1145)) + ((g27) & (!g39) & (g1101) & (!g1102) & (!g1145)) + ((g27) & (!g39) & (g1101) & (!g1102) & (g1145)) + ((g27) & (!g39) & (g1101) & (g1102) & (!g1145)) + ((g27) & (!g39) & (g1101) & (g1102) & (g1145)) + ((g27) & (g39) & (!g1101) & (!g1102) & (g1145)) + ((g27) & (g39) & (!g1101) & (g1102) & (!g1145)) + ((g27) & (g39) & (!g1101) & (g1102) & (g1145)) + ((g27) & (g39) & (g1101) & (!g1102) & (!g1145)) + ((g27) & (g39) & (g1101) & (!g1102) & (g1145)) + ((g27) & (g39) & (g1101) & (g1102) & (!g1145)) + ((g27) & (g39) & (g1101) & (g1102) & (g1145)));
	assign g1147 = (((!g8) & (!g18) & (g1098) & (g1099) & (g1146)) + ((!g8) & (g18) & (g1098) & (!g1099) & (g1146)) + ((!g8) & (g18) & (g1098) & (g1099) & (!g1146)) + ((!g8) & (g18) & (g1098) & (g1099) & (g1146)) + ((g8) & (!g18) & (!g1098) & (g1099) & (g1146)) + ((g8) & (!g18) & (g1098) & (!g1099) & (!g1146)) + ((g8) & (!g18) & (g1098) & (!g1099) & (g1146)) + ((g8) & (!g18) & (g1098) & (g1099) & (!g1146)) + ((g8) & (!g18) & (g1098) & (g1099) & (g1146)) + ((g8) & (g18) & (!g1098) & (!g1099) & (g1146)) + ((g8) & (g18) & (!g1098) & (g1099) & (!g1146)) + ((g8) & (g18) & (!g1098) & (g1099) & (g1146)) + ((g8) & (g18) & (g1098) & (!g1099) & (!g1146)) + ((g8) & (g18) & (g1098) & (!g1099) & (g1146)) + ((g8) & (g18) & (g1098) & (g1099) & (!g1146)) + ((g8) & (g18) & (g1098) & (g1099) & (g1146)));
	assign g1148 = (((!g2) & (!g8) & (g1041) & (g1079)) + ((!g2) & (g8) & (!g1041) & (g1079)) + ((!g2) & (g8) & (g1041) & (!g1079)) + ((!g2) & (g8) & (g1041) & (g1079)) + ((g2) & (!g8) & (!g1041) & (!g1079)) + ((g2) & (!g8) & (!g1041) & (g1079)) + ((g2) & (!g8) & (g1041) & (!g1079)) + ((g2) & (g8) & (!g1041) & (!g1079)));
	assign g1149 = (((!g1040) & (!g1038) & (!g1083) & (g1148)) + ((!g1040) & (g1038) & (!g1083) & (g1148)) + ((!g1040) & (g1038) & (g1083) & (g1148)) + ((g1040) & (!g1038) & (!g1083) & (!g1148)) + ((g1040) & (!g1038) & (g1083) & (!g1148)) + ((g1040) & (!g1038) & (g1083) & (g1148)) + ((g1040) & (g1038) & (!g1083) & (!g1148)) + ((g1040) & (g1038) & (g1083) & (!g1148)));
	assign g1150 = (((!g4) & (!g2) & (!g1096) & (!g1147) & (g1149)) + ((!g4) & (!g2) & (!g1096) & (g1147) & (g1149)) + ((!g4) & (!g2) & (g1096) & (!g1147) & (g1149)) + ((!g4) & (!g2) & (g1096) & (g1147) & (!g1149)) + ((!g4) & (!g2) & (g1096) & (g1147) & (g1149)) + ((!g4) & (g2) & (!g1096) & (!g1147) & (g1149)) + ((!g4) & (g2) & (!g1096) & (g1147) & (!g1149)) + ((!g4) & (g2) & (!g1096) & (g1147) & (g1149)) + ((!g4) & (g2) & (g1096) & (!g1147) & (!g1149)) + ((!g4) & (g2) & (g1096) & (!g1147) & (g1149)) + ((!g4) & (g2) & (g1096) & (g1147) & (!g1149)) + ((!g4) & (g2) & (g1096) & (g1147) & (g1149)) + ((g4) & (!g2) & (g1096) & (g1147) & (g1149)) + ((g4) & (g2) & (!g1096) & (g1147) & (g1149)) + ((g4) & (g2) & (g1096) & (!g1147) & (g1149)) + ((g4) & (g2) & (g1096) & (g1147) & (g1149)));
	assign g1151 = (((!g4) & (!g1080) & (g1081)) + ((!g4) & (g1080) & (!g1081)) + ((!g4) & (g1080) & (g1081)) + ((g4) & (g1080) & (g1081)));
	assign g1152 = (((!g1039) & (!g1151) & (!g1038) & (!g1083)) + ((!g1039) & (!g1151) & (g1038) & (!g1083)) + ((!g1039) & (!g1151) & (g1038) & (g1083)) + ((g1039) & (g1151) & (!g1038) & (!g1083)) + ((g1039) & (g1151) & (!g1038) & (g1083)) + ((g1039) & (g1151) & (g1038) & (!g1083)) + ((g1039) & (g1151) & (g1038) & (g1083)));
	assign g1153 = (((!g1) & (g1039) & (!g1151) & (!g1038) & (g1083)) + ((!g1) & (g1039) & (g1151) & (!g1038) & (g1083)) + ((g1) & (!g1039) & (g1151) & (g1038) & (!g1083)) + ((g1) & (!g1039) & (g1151) & (g1038) & (g1083)) + ((g1) & (g1039) & (!g1151) & (!g1038) & (!g1083)) + ((g1) & (g1039) & (!g1151) & (!g1038) & (g1083)) + ((g1) & (g1039) & (!g1151) & (g1038) & (!g1083)) + ((g1) & (g1039) & (!g1151) & (g1038) & (g1083)) + ((g1) & (g1039) & (g1151) & (!g1038) & (g1083)));
	assign g1154 = (((!g1) & (!g1095) & (!g1150) & (!g1152) & (!g1153)) + ((g1) & (!g1095) & (!g1150) & (!g1152) & (!g1153)) + ((g1) & (!g1095) & (!g1150) & (g1152) & (!g1153)) + ((g1) & (!g1095) & (g1150) & (!g1152) & (!g1153)) + ((g1) & (!g1095) & (g1150) & (g1152) & (!g1153)) + ((g1) & (g1095) & (!g1150) & (!g1152) & (!g1153)) + ((g1) & (g1095) & (!g1150) & (g1152) & (!g1153)));
	assign g1155 = (((!g744) & (!g1084) & (g1094) & (!g1154)) + ((!g744) & (g1084) & (!g1094) & (!g1154)) + ((!g744) & (g1084) & (!g1094) & (g1154)) + ((!g744) & (g1084) & (g1094) & (g1154)) + ((g744) & (!g1084) & (!g1094) & (!g1154)) + ((g744) & (g1084) & (!g1094) & (g1154)) + ((g744) & (g1084) & (g1094) & (!g1154)) + ((g744) & (g1084) & (g1094) & (g1154)));
	assign g1156 = (((!g803) & (!g851) & (!g1086) & (g1087) & (g1093) & (!g1154)) + ((!g803) & (!g851) & (g1086) & (!g1087) & (!g1093) & (!g1154)) + ((!g803) & (!g851) & (g1086) & (!g1087) & (!g1093) & (g1154)) + ((!g803) & (!g851) & (g1086) & (!g1087) & (g1093) & (!g1154)) + ((!g803) & (!g851) & (g1086) & (!g1087) & (g1093) & (g1154)) + ((!g803) & (!g851) & (g1086) & (g1087) & (!g1093) & (!g1154)) + ((!g803) & (!g851) & (g1086) & (g1087) & (!g1093) & (g1154)) + ((!g803) & (!g851) & (g1086) & (g1087) & (g1093) & (g1154)) + ((!g803) & (g851) & (!g1086) & (!g1087) & (g1093) & (!g1154)) + ((!g803) & (g851) & (!g1086) & (g1087) & (!g1093) & (!g1154)) + ((!g803) & (g851) & (!g1086) & (g1087) & (g1093) & (!g1154)) + ((!g803) & (g851) & (g1086) & (!g1087) & (!g1093) & (!g1154)) + ((!g803) & (g851) & (g1086) & (!g1087) & (!g1093) & (g1154)) + ((!g803) & (g851) & (g1086) & (!g1087) & (g1093) & (g1154)) + ((!g803) & (g851) & (g1086) & (g1087) & (!g1093) & (g1154)) + ((!g803) & (g851) & (g1086) & (g1087) & (g1093) & (g1154)) + ((g803) & (!g851) & (!g1086) & (!g1087) & (!g1093) & (!g1154)) + ((g803) & (!g851) & (!g1086) & (!g1087) & (g1093) & (!g1154)) + ((g803) & (!g851) & (!g1086) & (g1087) & (!g1093) & (!g1154)) + ((g803) & (!g851) & (g1086) & (!g1087) & (!g1093) & (g1154)) + ((g803) & (!g851) & (g1086) & (!g1087) & (g1093) & (g1154)) + ((g803) & (!g851) & (g1086) & (g1087) & (!g1093) & (g1154)) + ((g803) & (!g851) & (g1086) & (g1087) & (g1093) & (!g1154)) + ((g803) & (!g851) & (g1086) & (g1087) & (g1093) & (g1154)) + ((g803) & (g851) & (!g1086) & (!g1087) & (!g1093) & (!g1154)) + ((g803) & (g851) & (g1086) & (!g1087) & (!g1093) & (g1154)) + ((g803) & (g851) & (g1086) & (!g1087) & (g1093) & (!g1154)) + ((g803) & (g851) & (g1086) & (!g1087) & (g1093) & (g1154)) + ((g803) & (g851) & (g1086) & (g1087) & (!g1093) & (!g1154)) + ((g803) & (g851) & (g1086) & (g1087) & (!g1093) & (g1154)) + ((g803) & (g851) & (g1086) & (g1087) & (g1093) & (!g1154)) + ((g803) & (g851) & (g1086) & (g1087) & (g1093) & (g1154)));
	assign g1157 = (((!g851) & (!g1087) & (g1093) & (!g1154)) + ((!g851) & (g1087) & (!g1093) & (!g1154)) + ((!g851) & (g1087) & (!g1093) & (g1154)) + ((!g851) & (g1087) & (g1093) & (g1154)) + ((g851) & (!g1087) & (!g1093) & (!g1154)) + ((g851) & (g1087) & (!g1093) & (g1154)) + ((g851) & (g1087) & (g1093) & (!g1154)) + ((g851) & (g1087) & (g1093) & (g1154)));
	assign g1158 = (((!g914) & (!g1032) & (!g1089) & (g1090) & (g1092) & (!g1154)) + ((!g914) & (!g1032) & (g1089) & (!g1090) & (!g1092) & (!g1154)) + ((!g914) & (!g1032) & (g1089) & (!g1090) & (!g1092) & (g1154)) + ((!g914) & (!g1032) & (g1089) & (!g1090) & (g1092) & (!g1154)) + ((!g914) & (!g1032) & (g1089) & (!g1090) & (g1092) & (g1154)) + ((!g914) & (!g1032) & (g1089) & (g1090) & (!g1092) & (!g1154)) + ((!g914) & (!g1032) & (g1089) & (g1090) & (!g1092) & (g1154)) + ((!g914) & (!g1032) & (g1089) & (g1090) & (g1092) & (g1154)) + ((!g914) & (g1032) & (!g1089) & (!g1090) & (g1092) & (!g1154)) + ((!g914) & (g1032) & (!g1089) & (g1090) & (!g1092) & (!g1154)) + ((!g914) & (g1032) & (!g1089) & (g1090) & (g1092) & (!g1154)) + ((!g914) & (g1032) & (g1089) & (!g1090) & (!g1092) & (!g1154)) + ((!g914) & (g1032) & (g1089) & (!g1090) & (!g1092) & (g1154)) + ((!g914) & (g1032) & (g1089) & (!g1090) & (g1092) & (g1154)) + ((!g914) & (g1032) & (g1089) & (g1090) & (!g1092) & (g1154)) + ((!g914) & (g1032) & (g1089) & (g1090) & (g1092) & (g1154)) + ((g914) & (!g1032) & (!g1089) & (!g1090) & (!g1092) & (!g1154)) + ((g914) & (!g1032) & (!g1089) & (!g1090) & (g1092) & (!g1154)) + ((g914) & (!g1032) & (!g1089) & (g1090) & (!g1092) & (!g1154)) + ((g914) & (!g1032) & (g1089) & (!g1090) & (!g1092) & (g1154)) + ((g914) & (!g1032) & (g1089) & (!g1090) & (g1092) & (g1154)) + ((g914) & (!g1032) & (g1089) & (g1090) & (!g1092) & (g1154)) + ((g914) & (!g1032) & (g1089) & (g1090) & (g1092) & (!g1154)) + ((g914) & (!g1032) & (g1089) & (g1090) & (g1092) & (g1154)) + ((g914) & (g1032) & (!g1089) & (!g1090) & (!g1092) & (!g1154)) + ((g914) & (g1032) & (g1089) & (!g1090) & (!g1092) & (g1154)) + ((g914) & (g1032) & (g1089) & (!g1090) & (g1092) & (!g1154)) + ((g914) & (g1032) & (g1089) & (!g1090) & (g1092) & (g1154)) + ((g914) & (g1032) & (g1089) & (g1090) & (!g1092) & (!g1154)) + ((g914) & (g1032) & (g1089) & (g1090) & (!g1092) & (g1154)) + ((g914) & (g1032) & (g1089) & (g1090) & (g1092) & (!g1154)) + ((g914) & (g1032) & (g1089) & (g1090) & (g1092) & (g1154)));
	assign g1159 = (((!g1032) & (!g1090) & (g1092) & (!g1154)) + ((!g1032) & (g1090) & (!g1092) & (!g1154)) + ((!g1032) & (g1090) & (!g1092) & (g1154)) + ((!g1032) & (g1090) & (g1092) & (g1154)) + ((g1032) & (!g1090) & (!g1092) & (!g1154)) + ((g1032) & (g1090) & (!g1092) & (g1154)) + ((g1032) & (g1090) & (g1092) & (!g1154)) + ((g1032) & (g1090) & (g1092) & (g1154)));
	assign g1160 = (((!g1038) & (g1083)));
	assign g1161 = (((!g1030) & (!ax58x) & (!ax59x) & (!g1160) & (!g1091) & (g1154)) + ((!g1030) & (!ax58x) & (!ax59x) & (!g1160) & (g1091) & (!g1154)) + ((!g1030) & (!ax58x) & (!ax59x) & (!g1160) & (g1091) & (g1154)) + ((!g1030) & (!ax58x) & (!ax59x) & (g1160) & (!g1091) & (!g1154)) + ((!g1030) & (!ax58x) & (ax59x) & (!g1160) & (!g1091) & (!g1154)) + ((!g1030) & (!ax58x) & (ax59x) & (g1160) & (!g1091) & (g1154)) + ((!g1030) & (!ax58x) & (ax59x) & (g1160) & (g1091) & (!g1154)) + ((!g1030) & (!ax58x) & (ax59x) & (g1160) & (g1091) & (g1154)) + ((!g1030) & (ax58x) & (!ax59x) & (g1160) & (!g1091) & (!g1154)) + ((!g1030) & (ax58x) & (!ax59x) & (g1160) & (g1091) & (!g1154)) + ((!g1030) & (ax58x) & (ax59x) & (!g1160) & (!g1091) & (!g1154)) + ((!g1030) & (ax58x) & (ax59x) & (!g1160) & (!g1091) & (g1154)) + ((!g1030) & (ax58x) & (ax59x) & (!g1160) & (g1091) & (!g1154)) + ((!g1030) & (ax58x) & (ax59x) & (!g1160) & (g1091) & (g1154)) + ((!g1030) & (ax58x) & (ax59x) & (g1160) & (!g1091) & (g1154)) + ((!g1030) & (ax58x) & (ax59x) & (g1160) & (g1091) & (g1154)) + ((g1030) & (!ax58x) & (!ax59x) & (!g1160) & (!g1091) & (!g1154)) + ((g1030) & (!ax58x) & (!ax59x) & (!g1160) & (!g1091) & (g1154)) + ((g1030) & (!ax58x) & (!ax59x) & (!g1160) & (g1091) & (g1154)) + ((g1030) & (!ax58x) & (!ax59x) & (g1160) & (g1091) & (!g1154)) + ((g1030) & (!ax58x) & (ax59x) & (!g1160) & (g1091) & (!g1154)) + ((g1030) & (!ax58x) & (ax59x) & (g1160) & (!g1091) & (!g1154)) + ((g1030) & (!ax58x) & (ax59x) & (g1160) & (!g1091) & (g1154)) + ((g1030) & (!ax58x) & (ax59x) & (g1160) & (g1091) & (g1154)) + ((g1030) & (ax58x) & (!ax59x) & (!g1160) & (!g1091) & (!g1154)) + ((g1030) & (ax58x) & (!ax59x) & (!g1160) & (g1091) & (!g1154)) + ((g1030) & (ax58x) & (ax59x) & (!g1160) & (!g1091) & (g1154)) + ((g1030) & (ax58x) & (ax59x) & (!g1160) & (g1091) & (g1154)) + ((g1030) & (ax58x) & (ax59x) & (g1160) & (!g1091) & (!g1154)) + ((g1030) & (ax58x) & (ax59x) & (g1160) & (!g1091) & (g1154)) + ((g1030) & (ax58x) & (ax59x) & (g1160) & (g1091) & (!g1154)) + ((g1030) & (ax58x) & (ax59x) & (g1160) & (g1091) & (g1154)));
	assign g1162 = (((!ax58x) & (!g1160) & (!g1091) & (g1154)) + ((!ax58x) & (!g1160) & (g1091) & (!g1154)) + ((!ax58x) & (!g1160) & (g1091) & (g1154)) + ((!ax58x) & (g1160) & (g1091) & (!g1154)) + ((ax58x) & (!g1160) & (!g1091) & (!g1154)) + ((ax58x) & (g1160) & (!g1091) & (!g1154)) + ((ax58x) & (g1160) & (!g1091) & (g1154)) + ((ax58x) & (g1160) & (g1091) & (g1154)));
	assign g1163 = (((!ax54x) & (!ax55x)));
	assign g1164 = (((!g1160) & (!ax56x) & (!ax57x) & (!g1154) & (!g1163)) + ((!g1160) & (!ax56x) & (ax57x) & (g1154) & (!g1163)) + ((!g1160) & (ax56x) & (ax57x) & (g1154) & (!g1163)) + ((!g1160) & (ax56x) & (ax57x) & (g1154) & (g1163)) + ((g1160) & (!ax56x) & (!ax57x) & (!g1154) & (!g1163)) + ((g1160) & (!ax56x) & (!ax57x) & (!g1154) & (g1163)) + ((g1160) & (!ax56x) & (!ax57x) & (g1154) & (!g1163)) + ((g1160) & (!ax56x) & (ax57x) & (!g1154) & (!g1163)) + ((g1160) & (!ax56x) & (ax57x) & (g1154) & (!g1163)) + ((g1160) & (!ax56x) & (ax57x) & (g1154) & (g1163)) + ((g1160) & (ax56x) & (!ax57x) & (g1154) & (!g1163)) + ((g1160) & (ax56x) & (!ax57x) & (g1154) & (g1163)) + ((g1160) & (ax56x) & (ax57x) & (!g1154) & (!g1163)) + ((g1160) & (ax56x) & (ax57x) & (!g1154) & (g1163)) + ((g1160) & (ax56x) & (ax57x) & (g1154) & (!g1163)) + ((g1160) & (ax56x) & (ax57x) & (g1154) & (g1163)));
	assign g1165 = (((!g1032) & (!g1030) & (g1161) & (g1162) & (g1164)) + ((!g1032) & (g1030) & (g1161) & (!g1162) & (g1164)) + ((!g1032) & (g1030) & (g1161) & (g1162) & (!g1164)) + ((!g1032) & (g1030) & (g1161) & (g1162) & (g1164)) + ((g1032) & (!g1030) & (!g1161) & (g1162) & (g1164)) + ((g1032) & (!g1030) & (g1161) & (!g1162) & (!g1164)) + ((g1032) & (!g1030) & (g1161) & (!g1162) & (g1164)) + ((g1032) & (!g1030) & (g1161) & (g1162) & (!g1164)) + ((g1032) & (!g1030) & (g1161) & (g1162) & (g1164)) + ((g1032) & (g1030) & (!g1161) & (!g1162) & (g1164)) + ((g1032) & (g1030) & (!g1161) & (g1162) & (!g1164)) + ((g1032) & (g1030) & (!g1161) & (g1162) & (g1164)) + ((g1032) & (g1030) & (g1161) & (!g1162) & (!g1164)) + ((g1032) & (g1030) & (g1161) & (!g1162) & (g1164)) + ((g1032) & (g1030) & (g1161) & (g1162) & (!g1164)) + ((g1032) & (g1030) & (g1161) & (g1162) & (g1164)));
	assign g1166 = (((!g851) & (!g914) & (g1158) & (g1159) & (g1165)) + ((!g851) & (g914) & (g1158) & (!g1159) & (g1165)) + ((!g851) & (g914) & (g1158) & (g1159) & (!g1165)) + ((!g851) & (g914) & (g1158) & (g1159) & (g1165)) + ((g851) & (!g914) & (!g1158) & (g1159) & (g1165)) + ((g851) & (!g914) & (g1158) & (!g1159) & (!g1165)) + ((g851) & (!g914) & (g1158) & (!g1159) & (g1165)) + ((g851) & (!g914) & (g1158) & (g1159) & (!g1165)) + ((g851) & (!g914) & (g1158) & (g1159) & (g1165)) + ((g851) & (g914) & (!g1158) & (!g1159) & (g1165)) + ((g851) & (g914) & (!g1158) & (g1159) & (!g1165)) + ((g851) & (g914) & (!g1158) & (g1159) & (g1165)) + ((g851) & (g914) & (g1158) & (!g1159) & (!g1165)) + ((g851) & (g914) & (g1158) & (!g1159) & (g1165)) + ((g851) & (g914) & (g1158) & (g1159) & (!g1165)) + ((g851) & (g914) & (g1158) & (g1159) & (g1165)));
	assign g1167 = (((!g744) & (!g803) & (g1156) & (g1157) & (g1166)) + ((!g744) & (g803) & (g1156) & (!g1157) & (g1166)) + ((!g744) & (g803) & (g1156) & (g1157) & (!g1166)) + ((!g744) & (g803) & (g1156) & (g1157) & (g1166)) + ((g744) & (!g803) & (!g1156) & (g1157) & (g1166)) + ((g744) & (!g803) & (g1156) & (!g1157) & (!g1166)) + ((g744) & (!g803) & (g1156) & (!g1157) & (g1166)) + ((g744) & (!g803) & (g1156) & (g1157) & (!g1166)) + ((g744) & (!g803) & (g1156) & (g1157) & (g1166)) + ((g744) & (g803) & (!g1156) & (!g1157) & (g1166)) + ((g744) & (g803) & (!g1156) & (g1157) & (!g1166)) + ((g744) & (g803) & (!g1156) & (g1157) & (g1166)) + ((g744) & (g803) & (g1156) & (!g1157) & (!g1166)) + ((g744) & (g803) & (g1156) & (!g1157) & (g1166)) + ((g744) & (g803) & (g1156) & (g1157) & (!g1166)) + ((g744) & (g803) & (g1156) & (g1157) & (g1166)));
	assign g1168 = (((g1) & (!g1095) & (g1150) & (g1153)) + ((g1) & (g1095) & (!g1150) & (!g1153)) + ((g1) & (g1095) & (!g1150) & (g1153)));
	assign g1169 = (((!g4) & (!g2) & (!g1096) & (!g1147) & (!g1149) & (!g1154)) + ((!g4) & (!g2) & (!g1096) & (!g1147) & (g1149) & (g1154)) + ((!g4) & (!g2) & (!g1096) & (g1147) & (!g1149) & (!g1154)) + ((!g4) & (!g2) & (!g1096) & (g1147) & (g1149) & (g1154)) + ((!g4) & (!g2) & (g1096) & (!g1147) & (!g1149) & (!g1154)) + ((!g4) & (!g2) & (g1096) & (!g1147) & (g1149) & (g1154)) + ((!g4) & (!g2) & (g1096) & (g1147) & (g1149) & (!g1154)) + ((!g4) & (!g2) & (g1096) & (g1147) & (g1149) & (g1154)) + ((!g4) & (g2) & (!g1096) & (!g1147) & (!g1149) & (!g1154)) + ((!g4) & (g2) & (!g1096) & (!g1147) & (g1149) & (g1154)) + ((!g4) & (g2) & (!g1096) & (g1147) & (g1149) & (!g1154)) + ((!g4) & (g2) & (!g1096) & (g1147) & (g1149) & (g1154)) + ((!g4) & (g2) & (g1096) & (!g1147) & (g1149) & (!g1154)) + ((!g4) & (g2) & (g1096) & (!g1147) & (g1149) & (g1154)) + ((!g4) & (g2) & (g1096) & (g1147) & (g1149) & (!g1154)) + ((!g4) & (g2) & (g1096) & (g1147) & (g1149) & (g1154)) + ((g4) & (!g2) & (!g1096) & (!g1147) & (g1149) & (!g1154)) + ((g4) & (!g2) & (!g1096) & (!g1147) & (g1149) & (g1154)) + ((g4) & (!g2) & (!g1096) & (g1147) & (g1149) & (!g1154)) + ((g4) & (!g2) & (!g1096) & (g1147) & (g1149) & (g1154)) + ((g4) & (!g2) & (g1096) & (!g1147) & (g1149) & (!g1154)) + ((g4) & (!g2) & (g1096) & (!g1147) & (g1149) & (g1154)) + ((g4) & (!g2) & (g1096) & (g1147) & (!g1149) & (!g1154)) + ((g4) & (!g2) & (g1096) & (g1147) & (g1149) & (g1154)) + ((g4) & (g2) & (!g1096) & (!g1147) & (g1149) & (!g1154)) + ((g4) & (g2) & (!g1096) & (!g1147) & (g1149) & (g1154)) + ((g4) & (g2) & (!g1096) & (g1147) & (!g1149) & (!g1154)) + ((g4) & (g2) & (!g1096) & (g1147) & (g1149) & (g1154)) + ((g4) & (g2) & (g1096) & (!g1147) & (!g1149) & (!g1154)) + ((g4) & (g2) & (g1096) & (!g1147) & (g1149) & (g1154)) + ((g4) & (g2) & (g1096) & (g1147) & (!g1149) & (!g1154)) + ((g4) & (g2) & (g1096) & (g1147) & (g1149) & (g1154)));
	assign g1170 = (((!g8) & (!g18) & (!g1098) & (g1099) & (g1146) & (!g1154)) + ((!g8) & (!g18) & (g1098) & (!g1099) & (!g1146) & (!g1154)) + ((!g8) & (!g18) & (g1098) & (!g1099) & (!g1146) & (g1154)) + ((!g8) & (!g18) & (g1098) & (!g1099) & (g1146) & (!g1154)) + ((!g8) & (!g18) & (g1098) & (!g1099) & (g1146) & (g1154)) + ((!g8) & (!g18) & (g1098) & (g1099) & (!g1146) & (!g1154)) + ((!g8) & (!g18) & (g1098) & (g1099) & (!g1146) & (g1154)) + ((!g8) & (!g18) & (g1098) & (g1099) & (g1146) & (g1154)) + ((!g8) & (g18) & (!g1098) & (!g1099) & (g1146) & (!g1154)) + ((!g8) & (g18) & (!g1098) & (g1099) & (!g1146) & (!g1154)) + ((!g8) & (g18) & (!g1098) & (g1099) & (g1146) & (!g1154)) + ((!g8) & (g18) & (g1098) & (!g1099) & (!g1146) & (!g1154)) + ((!g8) & (g18) & (g1098) & (!g1099) & (!g1146) & (g1154)) + ((!g8) & (g18) & (g1098) & (!g1099) & (g1146) & (g1154)) + ((!g8) & (g18) & (g1098) & (g1099) & (!g1146) & (g1154)) + ((!g8) & (g18) & (g1098) & (g1099) & (g1146) & (g1154)) + ((g8) & (!g18) & (!g1098) & (!g1099) & (!g1146) & (!g1154)) + ((g8) & (!g18) & (!g1098) & (!g1099) & (g1146) & (!g1154)) + ((g8) & (!g18) & (!g1098) & (g1099) & (!g1146) & (!g1154)) + ((g8) & (!g18) & (g1098) & (!g1099) & (!g1146) & (g1154)) + ((g8) & (!g18) & (g1098) & (!g1099) & (g1146) & (g1154)) + ((g8) & (!g18) & (g1098) & (g1099) & (!g1146) & (g1154)) + ((g8) & (!g18) & (g1098) & (g1099) & (g1146) & (!g1154)) + ((g8) & (!g18) & (g1098) & (g1099) & (g1146) & (g1154)) + ((g8) & (g18) & (!g1098) & (!g1099) & (!g1146) & (!g1154)) + ((g8) & (g18) & (g1098) & (!g1099) & (!g1146) & (g1154)) + ((g8) & (g18) & (g1098) & (!g1099) & (g1146) & (!g1154)) + ((g8) & (g18) & (g1098) & (!g1099) & (g1146) & (g1154)) + ((g8) & (g18) & (g1098) & (g1099) & (!g1146) & (!g1154)) + ((g8) & (g18) & (g1098) & (g1099) & (!g1146) & (g1154)) + ((g8) & (g18) & (g1098) & (g1099) & (g1146) & (!g1154)) + ((g8) & (g18) & (g1098) & (g1099) & (g1146) & (g1154)));
	assign g1171 = (((!g18) & (!g1099) & (g1146) & (!g1154)) + ((!g18) & (g1099) & (!g1146) & (!g1154)) + ((!g18) & (g1099) & (!g1146) & (g1154)) + ((!g18) & (g1099) & (g1146) & (g1154)) + ((g18) & (!g1099) & (!g1146) & (!g1154)) + ((g18) & (g1099) & (!g1146) & (g1154)) + ((g18) & (g1099) & (g1146) & (!g1154)) + ((g18) & (g1099) & (g1146) & (g1154)));
	assign g1172 = (((!g27) & (!g39) & (!g1101) & (g1102) & (g1145) & (!g1154)) + ((!g27) & (!g39) & (g1101) & (!g1102) & (!g1145) & (!g1154)) + ((!g27) & (!g39) & (g1101) & (!g1102) & (!g1145) & (g1154)) + ((!g27) & (!g39) & (g1101) & (!g1102) & (g1145) & (!g1154)) + ((!g27) & (!g39) & (g1101) & (!g1102) & (g1145) & (g1154)) + ((!g27) & (!g39) & (g1101) & (g1102) & (!g1145) & (!g1154)) + ((!g27) & (!g39) & (g1101) & (g1102) & (!g1145) & (g1154)) + ((!g27) & (!g39) & (g1101) & (g1102) & (g1145) & (g1154)) + ((!g27) & (g39) & (!g1101) & (!g1102) & (g1145) & (!g1154)) + ((!g27) & (g39) & (!g1101) & (g1102) & (!g1145) & (!g1154)) + ((!g27) & (g39) & (!g1101) & (g1102) & (g1145) & (!g1154)) + ((!g27) & (g39) & (g1101) & (!g1102) & (!g1145) & (!g1154)) + ((!g27) & (g39) & (g1101) & (!g1102) & (!g1145) & (g1154)) + ((!g27) & (g39) & (g1101) & (!g1102) & (g1145) & (g1154)) + ((!g27) & (g39) & (g1101) & (g1102) & (!g1145) & (g1154)) + ((!g27) & (g39) & (g1101) & (g1102) & (g1145) & (g1154)) + ((g27) & (!g39) & (!g1101) & (!g1102) & (!g1145) & (!g1154)) + ((g27) & (!g39) & (!g1101) & (!g1102) & (g1145) & (!g1154)) + ((g27) & (!g39) & (!g1101) & (g1102) & (!g1145) & (!g1154)) + ((g27) & (!g39) & (g1101) & (!g1102) & (!g1145) & (g1154)) + ((g27) & (!g39) & (g1101) & (!g1102) & (g1145) & (g1154)) + ((g27) & (!g39) & (g1101) & (g1102) & (!g1145) & (g1154)) + ((g27) & (!g39) & (g1101) & (g1102) & (g1145) & (!g1154)) + ((g27) & (!g39) & (g1101) & (g1102) & (g1145) & (g1154)) + ((g27) & (g39) & (!g1101) & (!g1102) & (!g1145) & (!g1154)) + ((g27) & (g39) & (g1101) & (!g1102) & (!g1145) & (g1154)) + ((g27) & (g39) & (g1101) & (!g1102) & (g1145) & (!g1154)) + ((g27) & (g39) & (g1101) & (!g1102) & (g1145) & (g1154)) + ((g27) & (g39) & (g1101) & (g1102) & (!g1145) & (!g1154)) + ((g27) & (g39) & (g1101) & (g1102) & (!g1145) & (g1154)) + ((g27) & (g39) & (g1101) & (g1102) & (g1145) & (!g1154)) + ((g27) & (g39) & (g1101) & (g1102) & (g1145) & (g1154)));
	assign g1173 = (((!g39) & (!g1102) & (g1145) & (!g1154)) + ((!g39) & (g1102) & (!g1145) & (!g1154)) + ((!g39) & (g1102) & (!g1145) & (g1154)) + ((!g39) & (g1102) & (g1145) & (g1154)) + ((g39) & (!g1102) & (!g1145) & (!g1154)) + ((g39) & (g1102) & (!g1145) & (g1154)) + ((g39) & (g1102) & (g1145) & (!g1154)) + ((g39) & (g1102) & (g1145) & (g1154)));
	assign g1174 = (((!g54) & (!g68) & (!g1104) & (g1105) & (g1144) & (!g1154)) + ((!g54) & (!g68) & (g1104) & (!g1105) & (!g1144) & (!g1154)) + ((!g54) & (!g68) & (g1104) & (!g1105) & (!g1144) & (g1154)) + ((!g54) & (!g68) & (g1104) & (!g1105) & (g1144) & (!g1154)) + ((!g54) & (!g68) & (g1104) & (!g1105) & (g1144) & (g1154)) + ((!g54) & (!g68) & (g1104) & (g1105) & (!g1144) & (!g1154)) + ((!g54) & (!g68) & (g1104) & (g1105) & (!g1144) & (g1154)) + ((!g54) & (!g68) & (g1104) & (g1105) & (g1144) & (g1154)) + ((!g54) & (g68) & (!g1104) & (!g1105) & (g1144) & (!g1154)) + ((!g54) & (g68) & (!g1104) & (g1105) & (!g1144) & (!g1154)) + ((!g54) & (g68) & (!g1104) & (g1105) & (g1144) & (!g1154)) + ((!g54) & (g68) & (g1104) & (!g1105) & (!g1144) & (!g1154)) + ((!g54) & (g68) & (g1104) & (!g1105) & (!g1144) & (g1154)) + ((!g54) & (g68) & (g1104) & (!g1105) & (g1144) & (g1154)) + ((!g54) & (g68) & (g1104) & (g1105) & (!g1144) & (g1154)) + ((!g54) & (g68) & (g1104) & (g1105) & (g1144) & (g1154)) + ((g54) & (!g68) & (!g1104) & (!g1105) & (!g1144) & (!g1154)) + ((g54) & (!g68) & (!g1104) & (!g1105) & (g1144) & (!g1154)) + ((g54) & (!g68) & (!g1104) & (g1105) & (!g1144) & (!g1154)) + ((g54) & (!g68) & (g1104) & (!g1105) & (!g1144) & (g1154)) + ((g54) & (!g68) & (g1104) & (!g1105) & (g1144) & (g1154)) + ((g54) & (!g68) & (g1104) & (g1105) & (!g1144) & (g1154)) + ((g54) & (!g68) & (g1104) & (g1105) & (g1144) & (!g1154)) + ((g54) & (!g68) & (g1104) & (g1105) & (g1144) & (g1154)) + ((g54) & (g68) & (!g1104) & (!g1105) & (!g1144) & (!g1154)) + ((g54) & (g68) & (g1104) & (!g1105) & (!g1144) & (g1154)) + ((g54) & (g68) & (g1104) & (!g1105) & (g1144) & (!g1154)) + ((g54) & (g68) & (g1104) & (!g1105) & (g1144) & (g1154)) + ((g54) & (g68) & (g1104) & (g1105) & (!g1144) & (!g1154)) + ((g54) & (g68) & (g1104) & (g1105) & (!g1144) & (g1154)) + ((g54) & (g68) & (g1104) & (g1105) & (g1144) & (!g1154)) + ((g54) & (g68) & (g1104) & (g1105) & (g1144) & (g1154)));
	assign g1175 = (((!g68) & (!g1105) & (g1144) & (!g1154)) + ((!g68) & (g1105) & (!g1144) & (!g1154)) + ((!g68) & (g1105) & (!g1144) & (g1154)) + ((!g68) & (g1105) & (g1144) & (g1154)) + ((g68) & (!g1105) & (!g1144) & (!g1154)) + ((g68) & (g1105) & (!g1144) & (g1154)) + ((g68) & (g1105) & (g1144) & (!g1154)) + ((g68) & (g1105) & (g1144) & (g1154)));
	assign g1176 = (((!g87) & (!g104) & (!g1107) & (g1108) & (g1143) & (!g1154)) + ((!g87) & (!g104) & (g1107) & (!g1108) & (!g1143) & (!g1154)) + ((!g87) & (!g104) & (g1107) & (!g1108) & (!g1143) & (g1154)) + ((!g87) & (!g104) & (g1107) & (!g1108) & (g1143) & (!g1154)) + ((!g87) & (!g104) & (g1107) & (!g1108) & (g1143) & (g1154)) + ((!g87) & (!g104) & (g1107) & (g1108) & (!g1143) & (!g1154)) + ((!g87) & (!g104) & (g1107) & (g1108) & (!g1143) & (g1154)) + ((!g87) & (!g104) & (g1107) & (g1108) & (g1143) & (g1154)) + ((!g87) & (g104) & (!g1107) & (!g1108) & (g1143) & (!g1154)) + ((!g87) & (g104) & (!g1107) & (g1108) & (!g1143) & (!g1154)) + ((!g87) & (g104) & (!g1107) & (g1108) & (g1143) & (!g1154)) + ((!g87) & (g104) & (g1107) & (!g1108) & (!g1143) & (!g1154)) + ((!g87) & (g104) & (g1107) & (!g1108) & (!g1143) & (g1154)) + ((!g87) & (g104) & (g1107) & (!g1108) & (g1143) & (g1154)) + ((!g87) & (g104) & (g1107) & (g1108) & (!g1143) & (g1154)) + ((!g87) & (g104) & (g1107) & (g1108) & (g1143) & (g1154)) + ((g87) & (!g104) & (!g1107) & (!g1108) & (!g1143) & (!g1154)) + ((g87) & (!g104) & (!g1107) & (!g1108) & (g1143) & (!g1154)) + ((g87) & (!g104) & (!g1107) & (g1108) & (!g1143) & (!g1154)) + ((g87) & (!g104) & (g1107) & (!g1108) & (!g1143) & (g1154)) + ((g87) & (!g104) & (g1107) & (!g1108) & (g1143) & (g1154)) + ((g87) & (!g104) & (g1107) & (g1108) & (!g1143) & (g1154)) + ((g87) & (!g104) & (g1107) & (g1108) & (g1143) & (!g1154)) + ((g87) & (!g104) & (g1107) & (g1108) & (g1143) & (g1154)) + ((g87) & (g104) & (!g1107) & (!g1108) & (!g1143) & (!g1154)) + ((g87) & (g104) & (g1107) & (!g1108) & (!g1143) & (g1154)) + ((g87) & (g104) & (g1107) & (!g1108) & (g1143) & (!g1154)) + ((g87) & (g104) & (g1107) & (!g1108) & (g1143) & (g1154)) + ((g87) & (g104) & (g1107) & (g1108) & (!g1143) & (!g1154)) + ((g87) & (g104) & (g1107) & (g1108) & (!g1143) & (g1154)) + ((g87) & (g104) & (g1107) & (g1108) & (g1143) & (!g1154)) + ((g87) & (g104) & (g1107) & (g1108) & (g1143) & (g1154)));
	assign g1177 = (((!g104) & (!g1108) & (g1143) & (!g1154)) + ((!g104) & (g1108) & (!g1143) & (!g1154)) + ((!g104) & (g1108) & (!g1143) & (g1154)) + ((!g104) & (g1108) & (g1143) & (g1154)) + ((g104) & (!g1108) & (!g1143) & (!g1154)) + ((g104) & (g1108) & (!g1143) & (g1154)) + ((g104) & (g1108) & (g1143) & (!g1154)) + ((g104) & (g1108) & (g1143) & (g1154)));
	assign g1178 = (((!g127) & (!g147) & (!g1110) & (g1111) & (g1142) & (!g1154)) + ((!g127) & (!g147) & (g1110) & (!g1111) & (!g1142) & (!g1154)) + ((!g127) & (!g147) & (g1110) & (!g1111) & (!g1142) & (g1154)) + ((!g127) & (!g147) & (g1110) & (!g1111) & (g1142) & (!g1154)) + ((!g127) & (!g147) & (g1110) & (!g1111) & (g1142) & (g1154)) + ((!g127) & (!g147) & (g1110) & (g1111) & (!g1142) & (!g1154)) + ((!g127) & (!g147) & (g1110) & (g1111) & (!g1142) & (g1154)) + ((!g127) & (!g147) & (g1110) & (g1111) & (g1142) & (g1154)) + ((!g127) & (g147) & (!g1110) & (!g1111) & (g1142) & (!g1154)) + ((!g127) & (g147) & (!g1110) & (g1111) & (!g1142) & (!g1154)) + ((!g127) & (g147) & (!g1110) & (g1111) & (g1142) & (!g1154)) + ((!g127) & (g147) & (g1110) & (!g1111) & (!g1142) & (!g1154)) + ((!g127) & (g147) & (g1110) & (!g1111) & (!g1142) & (g1154)) + ((!g127) & (g147) & (g1110) & (!g1111) & (g1142) & (g1154)) + ((!g127) & (g147) & (g1110) & (g1111) & (!g1142) & (g1154)) + ((!g127) & (g147) & (g1110) & (g1111) & (g1142) & (g1154)) + ((g127) & (!g147) & (!g1110) & (!g1111) & (!g1142) & (!g1154)) + ((g127) & (!g147) & (!g1110) & (!g1111) & (g1142) & (!g1154)) + ((g127) & (!g147) & (!g1110) & (g1111) & (!g1142) & (!g1154)) + ((g127) & (!g147) & (g1110) & (!g1111) & (!g1142) & (g1154)) + ((g127) & (!g147) & (g1110) & (!g1111) & (g1142) & (g1154)) + ((g127) & (!g147) & (g1110) & (g1111) & (!g1142) & (g1154)) + ((g127) & (!g147) & (g1110) & (g1111) & (g1142) & (!g1154)) + ((g127) & (!g147) & (g1110) & (g1111) & (g1142) & (g1154)) + ((g127) & (g147) & (!g1110) & (!g1111) & (!g1142) & (!g1154)) + ((g127) & (g147) & (g1110) & (!g1111) & (!g1142) & (g1154)) + ((g127) & (g147) & (g1110) & (!g1111) & (g1142) & (!g1154)) + ((g127) & (g147) & (g1110) & (!g1111) & (g1142) & (g1154)) + ((g127) & (g147) & (g1110) & (g1111) & (!g1142) & (!g1154)) + ((g127) & (g147) & (g1110) & (g1111) & (!g1142) & (g1154)) + ((g127) & (g147) & (g1110) & (g1111) & (g1142) & (!g1154)) + ((g127) & (g147) & (g1110) & (g1111) & (g1142) & (g1154)));
	assign g1179 = (((!g147) & (!g1111) & (g1142) & (!g1154)) + ((!g147) & (g1111) & (!g1142) & (!g1154)) + ((!g147) & (g1111) & (!g1142) & (g1154)) + ((!g147) & (g1111) & (g1142) & (g1154)) + ((g147) & (!g1111) & (!g1142) & (!g1154)) + ((g147) & (g1111) & (!g1142) & (g1154)) + ((g147) & (g1111) & (g1142) & (!g1154)) + ((g147) & (g1111) & (g1142) & (g1154)));
	assign g1180 = (((!g174) & (!g198) & (!g1113) & (g1114) & (g1141) & (!g1154)) + ((!g174) & (!g198) & (g1113) & (!g1114) & (!g1141) & (!g1154)) + ((!g174) & (!g198) & (g1113) & (!g1114) & (!g1141) & (g1154)) + ((!g174) & (!g198) & (g1113) & (!g1114) & (g1141) & (!g1154)) + ((!g174) & (!g198) & (g1113) & (!g1114) & (g1141) & (g1154)) + ((!g174) & (!g198) & (g1113) & (g1114) & (!g1141) & (!g1154)) + ((!g174) & (!g198) & (g1113) & (g1114) & (!g1141) & (g1154)) + ((!g174) & (!g198) & (g1113) & (g1114) & (g1141) & (g1154)) + ((!g174) & (g198) & (!g1113) & (!g1114) & (g1141) & (!g1154)) + ((!g174) & (g198) & (!g1113) & (g1114) & (!g1141) & (!g1154)) + ((!g174) & (g198) & (!g1113) & (g1114) & (g1141) & (!g1154)) + ((!g174) & (g198) & (g1113) & (!g1114) & (!g1141) & (!g1154)) + ((!g174) & (g198) & (g1113) & (!g1114) & (!g1141) & (g1154)) + ((!g174) & (g198) & (g1113) & (!g1114) & (g1141) & (g1154)) + ((!g174) & (g198) & (g1113) & (g1114) & (!g1141) & (g1154)) + ((!g174) & (g198) & (g1113) & (g1114) & (g1141) & (g1154)) + ((g174) & (!g198) & (!g1113) & (!g1114) & (!g1141) & (!g1154)) + ((g174) & (!g198) & (!g1113) & (!g1114) & (g1141) & (!g1154)) + ((g174) & (!g198) & (!g1113) & (g1114) & (!g1141) & (!g1154)) + ((g174) & (!g198) & (g1113) & (!g1114) & (!g1141) & (g1154)) + ((g174) & (!g198) & (g1113) & (!g1114) & (g1141) & (g1154)) + ((g174) & (!g198) & (g1113) & (g1114) & (!g1141) & (g1154)) + ((g174) & (!g198) & (g1113) & (g1114) & (g1141) & (!g1154)) + ((g174) & (!g198) & (g1113) & (g1114) & (g1141) & (g1154)) + ((g174) & (g198) & (!g1113) & (!g1114) & (!g1141) & (!g1154)) + ((g174) & (g198) & (g1113) & (!g1114) & (!g1141) & (g1154)) + ((g174) & (g198) & (g1113) & (!g1114) & (g1141) & (!g1154)) + ((g174) & (g198) & (g1113) & (!g1114) & (g1141) & (g1154)) + ((g174) & (g198) & (g1113) & (g1114) & (!g1141) & (!g1154)) + ((g174) & (g198) & (g1113) & (g1114) & (!g1141) & (g1154)) + ((g174) & (g198) & (g1113) & (g1114) & (g1141) & (!g1154)) + ((g174) & (g198) & (g1113) & (g1114) & (g1141) & (g1154)));
	assign g1181 = (((!g198) & (!g1114) & (g1141) & (!g1154)) + ((!g198) & (g1114) & (!g1141) & (!g1154)) + ((!g198) & (g1114) & (!g1141) & (g1154)) + ((!g198) & (g1114) & (g1141) & (g1154)) + ((g198) & (!g1114) & (!g1141) & (!g1154)) + ((g198) & (g1114) & (!g1141) & (g1154)) + ((g198) & (g1114) & (g1141) & (!g1154)) + ((g198) & (g1114) & (g1141) & (g1154)));
	assign g1182 = (((!g229) & (!g255) & (!g1116) & (g1117) & (g1140) & (!g1154)) + ((!g229) & (!g255) & (g1116) & (!g1117) & (!g1140) & (!g1154)) + ((!g229) & (!g255) & (g1116) & (!g1117) & (!g1140) & (g1154)) + ((!g229) & (!g255) & (g1116) & (!g1117) & (g1140) & (!g1154)) + ((!g229) & (!g255) & (g1116) & (!g1117) & (g1140) & (g1154)) + ((!g229) & (!g255) & (g1116) & (g1117) & (!g1140) & (!g1154)) + ((!g229) & (!g255) & (g1116) & (g1117) & (!g1140) & (g1154)) + ((!g229) & (!g255) & (g1116) & (g1117) & (g1140) & (g1154)) + ((!g229) & (g255) & (!g1116) & (!g1117) & (g1140) & (!g1154)) + ((!g229) & (g255) & (!g1116) & (g1117) & (!g1140) & (!g1154)) + ((!g229) & (g255) & (!g1116) & (g1117) & (g1140) & (!g1154)) + ((!g229) & (g255) & (g1116) & (!g1117) & (!g1140) & (!g1154)) + ((!g229) & (g255) & (g1116) & (!g1117) & (!g1140) & (g1154)) + ((!g229) & (g255) & (g1116) & (!g1117) & (g1140) & (g1154)) + ((!g229) & (g255) & (g1116) & (g1117) & (!g1140) & (g1154)) + ((!g229) & (g255) & (g1116) & (g1117) & (g1140) & (g1154)) + ((g229) & (!g255) & (!g1116) & (!g1117) & (!g1140) & (!g1154)) + ((g229) & (!g255) & (!g1116) & (!g1117) & (g1140) & (!g1154)) + ((g229) & (!g255) & (!g1116) & (g1117) & (!g1140) & (!g1154)) + ((g229) & (!g255) & (g1116) & (!g1117) & (!g1140) & (g1154)) + ((g229) & (!g255) & (g1116) & (!g1117) & (g1140) & (g1154)) + ((g229) & (!g255) & (g1116) & (g1117) & (!g1140) & (g1154)) + ((g229) & (!g255) & (g1116) & (g1117) & (g1140) & (!g1154)) + ((g229) & (!g255) & (g1116) & (g1117) & (g1140) & (g1154)) + ((g229) & (g255) & (!g1116) & (!g1117) & (!g1140) & (!g1154)) + ((g229) & (g255) & (g1116) & (!g1117) & (!g1140) & (g1154)) + ((g229) & (g255) & (g1116) & (!g1117) & (g1140) & (!g1154)) + ((g229) & (g255) & (g1116) & (!g1117) & (g1140) & (g1154)) + ((g229) & (g255) & (g1116) & (g1117) & (!g1140) & (!g1154)) + ((g229) & (g255) & (g1116) & (g1117) & (!g1140) & (g1154)) + ((g229) & (g255) & (g1116) & (g1117) & (g1140) & (!g1154)) + ((g229) & (g255) & (g1116) & (g1117) & (g1140) & (g1154)));
	assign g1183 = (((!g255) & (!g1117) & (g1140) & (!g1154)) + ((!g255) & (g1117) & (!g1140) & (!g1154)) + ((!g255) & (g1117) & (!g1140) & (g1154)) + ((!g255) & (g1117) & (g1140) & (g1154)) + ((g255) & (!g1117) & (!g1140) & (!g1154)) + ((g255) & (g1117) & (!g1140) & (g1154)) + ((g255) & (g1117) & (g1140) & (!g1154)) + ((g255) & (g1117) & (g1140) & (g1154)));
	assign g1184 = (((!g290) & (!g319) & (!g1119) & (g1120) & (g1139) & (!g1154)) + ((!g290) & (!g319) & (g1119) & (!g1120) & (!g1139) & (!g1154)) + ((!g290) & (!g319) & (g1119) & (!g1120) & (!g1139) & (g1154)) + ((!g290) & (!g319) & (g1119) & (!g1120) & (g1139) & (!g1154)) + ((!g290) & (!g319) & (g1119) & (!g1120) & (g1139) & (g1154)) + ((!g290) & (!g319) & (g1119) & (g1120) & (!g1139) & (!g1154)) + ((!g290) & (!g319) & (g1119) & (g1120) & (!g1139) & (g1154)) + ((!g290) & (!g319) & (g1119) & (g1120) & (g1139) & (g1154)) + ((!g290) & (g319) & (!g1119) & (!g1120) & (g1139) & (!g1154)) + ((!g290) & (g319) & (!g1119) & (g1120) & (!g1139) & (!g1154)) + ((!g290) & (g319) & (!g1119) & (g1120) & (g1139) & (!g1154)) + ((!g290) & (g319) & (g1119) & (!g1120) & (!g1139) & (!g1154)) + ((!g290) & (g319) & (g1119) & (!g1120) & (!g1139) & (g1154)) + ((!g290) & (g319) & (g1119) & (!g1120) & (g1139) & (g1154)) + ((!g290) & (g319) & (g1119) & (g1120) & (!g1139) & (g1154)) + ((!g290) & (g319) & (g1119) & (g1120) & (g1139) & (g1154)) + ((g290) & (!g319) & (!g1119) & (!g1120) & (!g1139) & (!g1154)) + ((g290) & (!g319) & (!g1119) & (!g1120) & (g1139) & (!g1154)) + ((g290) & (!g319) & (!g1119) & (g1120) & (!g1139) & (!g1154)) + ((g290) & (!g319) & (g1119) & (!g1120) & (!g1139) & (g1154)) + ((g290) & (!g319) & (g1119) & (!g1120) & (g1139) & (g1154)) + ((g290) & (!g319) & (g1119) & (g1120) & (!g1139) & (g1154)) + ((g290) & (!g319) & (g1119) & (g1120) & (g1139) & (!g1154)) + ((g290) & (!g319) & (g1119) & (g1120) & (g1139) & (g1154)) + ((g290) & (g319) & (!g1119) & (!g1120) & (!g1139) & (!g1154)) + ((g290) & (g319) & (g1119) & (!g1120) & (!g1139) & (g1154)) + ((g290) & (g319) & (g1119) & (!g1120) & (g1139) & (!g1154)) + ((g290) & (g319) & (g1119) & (!g1120) & (g1139) & (g1154)) + ((g290) & (g319) & (g1119) & (g1120) & (!g1139) & (!g1154)) + ((g290) & (g319) & (g1119) & (g1120) & (!g1139) & (g1154)) + ((g290) & (g319) & (g1119) & (g1120) & (g1139) & (!g1154)) + ((g290) & (g319) & (g1119) & (g1120) & (g1139) & (g1154)));
	assign g1185 = (((!g319) & (!g1120) & (g1139) & (!g1154)) + ((!g319) & (g1120) & (!g1139) & (!g1154)) + ((!g319) & (g1120) & (!g1139) & (g1154)) + ((!g319) & (g1120) & (g1139) & (g1154)) + ((g319) & (!g1120) & (!g1139) & (!g1154)) + ((g319) & (g1120) & (!g1139) & (g1154)) + ((g319) & (g1120) & (g1139) & (!g1154)) + ((g319) & (g1120) & (g1139) & (g1154)));
	assign g1186 = (((!g358) & (!g390) & (!g1122) & (g1123) & (g1138) & (!g1154)) + ((!g358) & (!g390) & (g1122) & (!g1123) & (!g1138) & (!g1154)) + ((!g358) & (!g390) & (g1122) & (!g1123) & (!g1138) & (g1154)) + ((!g358) & (!g390) & (g1122) & (!g1123) & (g1138) & (!g1154)) + ((!g358) & (!g390) & (g1122) & (!g1123) & (g1138) & (g1154)) + ((!g358) & (!g390) & (g1122) & (g1123) & (!g1138) & (!g1154)) + ((!g358) & (!g390) & (g1122) & (g1123) & (!g1138) & (g1154)) + ((!g358) & (!g390) & (g1122) & (g1123) & (g1138) & (g1154)) + ((!g358) & (g390) & (!g1122) & (!g1123) & (g1138) & (!g1154)) + ((!g358) & (g390) & (!g1122) & (g1123) & (!g1138) & (!g1154)) + ((!g358) & (g390) & (!g1122) & (g1123) & (g1138) & (!g1154)) + ((!g358) & (g390) & (g1122) & (!g1123) & (!g1138) & (!g1154)) + ((!g358) & (g390) & (g1122) & (!g1123) & (!g1138) & (g1154)) + ((!g358) & (g390) & (g1122) & (!g1123) & (g1138) & (g1154)) + ((!g358) & (g390) & (g1122) & (g1123) & (!g1138) & (g1154)) + ((!g358) & (g390) & (g1122) & (g1123) & (g1138) & (g1154)) + ((g358) & (!g390) & (!g1122) & (!g1123) & (!g1138) & (!g1154)) + ((g358) & (!g390) & (!g1122) & (!g1123) & (g1138) & (!g1154)) + ((g358) & (!g390) & (!g1122) & (g1123) & (!g1138) & (!g1154)) + ((g358) & (!g390) & (g1122) & (!g1123) & (!g1138) & (g1154)) + ((g358) & (!g390) & (g1122) & (!g1123) & (g1138) & (g1154)) + ((g358) & (!g390) & (g1122) & (g1123) & (!g1138) & (g1154)) + ((g358) & (!g390) & (g1122) & (g1123) & (g1138) & (!g1154)) + ((g358) & (!g390) & (g1122) & (g1123) & (g1138) & (g1154)) + ((g358) & (g390) & (!g1122) & (!g1123) & (!g1138) & (!g1154)) + ((g358) & (g390) & (g1122) & (!g1123) & (!g1138) & (g1154)) + ((g358) & (g390) & (g1122) & (!g1123) & (g1138) & (!g1154)) + ((g358) & (g390) & (g1122) & (!g1123) & (g1138) & (g1154)) + ((g358) & (g390) & (g1122) & (g1123) & (!g1138) & (!g1154)) + ((g358) & (g390) & (g1122) & (g1123) & (!g1138) & (g1154)) + ((g358) & (g390) & (g1122) & (g1123) & (g1138) & (!g1154)) + ((g358) & (g390) & (g1122) & (g1123) & (g1138) & (g1154)));
	assign g1187 = (((!g390) & (!g1123) & (g1138) & (!g1154)) + ((!g390) & (g1123) & (!g1138) & (!g1154)) + ((!g390) & (g1123) & (!g1138) & (g1154)) + ((!g390) & (g1123) & (g1138) & (g1154)) + ((g390) & (!g1123) & (!g1138) & (!g1154)) + ((g390) & (g1123) & (!g1138) & (g1154)) + ((g390) & (g1123) & (g1138) & (!g1154)) + ((g390) & (g1123) & (g1138) & (g1154)));
	assign g1188 = (((!g433) & (!g468) & (!g1125) & (g1126) & (g1137) & (!g1154)) + ((!g433) & (!g468) & (g1125) & (!g1126) & (!g1137) & (!g1154)) + ((!g433) & (!g468) & (g1125) & (!g1126) & (!g1137) & (g1154)) + ((!g433) & (!g468) & (g1125) & (!g1126) & (g1137) & (!g1154)) + ((!g433) & (!g468) & (g1125) & (!g1126) & (g1137) & (g1154)) + ((!g433) & (!g468) & (g1125) & (g1126) & (!g1137) & (!g1154)) + ((!g433) & (!g468) & (g1125) & (g1126) & (!g1137) & (g1154)) + ((!g433) & (!g468) & (g1125) & (g1126) & (g1137) & (g1154)) + ((!g433) & (g468) & (!g1125) & (!g1126) & (g1137) & (!g1154)) + ((!g433) & (g468) & (!g1125) & (g1126) & (!g1137) & (!g1154)) + ((!g433) & (g468) & (!g1125) & (g1126) & (g1137) & (!g1154)) + ((!g433) & (g468) & (g1125) & (!g1126) & (!g1137) & (!g1154)) + ((!g433) & (g468) & (g1125) & (!g1126) & (!g1137) & (g1154)) + ((!g433) & (g468) & (g1125) & (!g1126) & (g1137) & (g1154)) + ((!g433) & (g468) & (g1125) & (g1126) & (!g1137) & (g1154)) + ((!g433) & (g468) & (g1125) & (g1126) & (g1137) & (g1154)) + ((g433) & (!g468) & (!g1125) & (!g1126) & (!g1137) & (!g1154)) + ((g433) & (!g468) & (!g1125) & (!g1126) & (g1137) & (!g1154)) + ((g433) & (!g468) & (!g1125) & (g1126) & (!g1137) & (!g1154)) + ((g433) & (!g468) & (g1125) & (!g1126) & (!g1137) & (g1154)) + ((g433) & (!g468) & (g1125) & (!g1126) & (g1137) & (g1154)) + ((g433) & (!g468) & (g1125) & (g1126) & (!g1137) & (g1154)) + ((g433) & (!g468) & (g1125) & (g1126) & (g1137) & (!g1154)) + ((g433) & (!g468) & (g1125) & (g1126) & (g1137) & (g1154)) + ((g433) & (g468) & (!g1125) & (!g1126) & (!g1137) & (!g1154)) + ((g433) & (g468) & (g1125) & (!g1126) & (!g1137) & (g1154)) + ((g433) & (g468) & (g1125) & (!g1126) & (g1137) & (!g1154)) + ((g433) & (g468) & (g1125) & (!g1126) & (g1137) & (g1154)) + ((g433) & (g468) & (g1125) & (g1126) & (!g1137) & (!g1154)) + ((g433) & (g468) & (g1125) & (g1126) & (!g1137) & (g1154)) + ((g433) & (g468) & (g1125) & (g1126) & (g1137) & (!g1154)) + ((g433) & (g468) & (g1125) & (g1126) & (g1137) & (g1154)));
	assign g1189 = (((!g468) & (!g1126) & (g1137) & (!g1154)) + ((!g468) & (g1126) & (!g1137) & (!g1154)) + ((!g468) & (g1126) & (!g1137) & (g1154)) + ((!g468) & (g1126) & (g1137) & (g1154)) + ((g468) & (!g1126) & (!g1137) & (!g1154)) + ((g468) & (g1126) & (!g1137) & (g1154)) + ((g468) & (g1126) & (g1137) & (!g1154)) + ((g468) & (g1126) & (g1137) & (g1154)));
	assign g1190 = (((!g515) & (!g553) & (!g1128) & (g1129) & (g1136) & (!g1154)) + ((!g515) & (!g553) & (g1128) & (!g1129) & (!g1136) & (!g1154)) + ((!g515) & (!g553) & (g1128) & (!g1129) & (!g1136) & (g1154)) + ((!g515) & (!g553) & (g1128) & (!g1129) & (g1136) & (!g1154)) + ((!g515) & (!g553) & (g1128) & (!g1129) & (g1136) & (g1154)) + ((!g515) & (!g553) & (g1128) & (g1129) & (!g1136) & (!g1154)) + ((!g515) & (!g553) & (g1128) & (g1129) & (!g1136) & (g1154)) + ((!g515) & (!g553) & (g1128) & (g1129) & (g1136) & (g1154)) + ((!g515) & (g553) & (!g1128) & (!g1129) & (g1136) & (!g1154)) + ((!g515) & (g553) & (!g1128) & (g1129) & (!g1136) & (!g1154)) + ((!g515) & (g553) & (!g1128) & (g1129) & (g1136) & (!g1154)) + ((!g515) & (g553) & (g1128) & (!g1129) & (!g1136) & (!g1154)) + ((!g515) & (g553) & (g1128) & (!g1129) & (!g1136) & (g1154)) + ((!g515) & (g553) & (g1128) & (!g1129) & (g1136) & (g1154)) + ((!g515) & (g553) & (g1128) & (g1129) & (!g1136) & (g1154)) + ((!g515) & (g553) & (g1128) & (g1129) & (g1136) & (g1154)) + ((g515) & (!g553) & (!g1128) & (!g1129) & (!g1136) & (!g1154)) + ((g515) & (!g553) & (!g1128) & (!g1129) & (g1136) & (!g1154)) + ((g515) & (!g553) & (!g1128) & (g1129) & (!g1136) & (!g1154)) + ((g515) & (!g553) & (g1128) & (!g1129) & (!g1136) & (g1154)) + ((g515) & (!g553) & (g1128) & (!g1129) & (g1136) & (g1154)) + ((g515) & (!g553) & (g1128) & (g1129) & (!g1136) & (g1154)) + ((g515) & (!g553) & (g1128) & (g1129) & (g1136) & (!g1154)) + ((g515) & (!g553) & (g1128) & (g1129) & (g1136) & (g1154)) + ((g515) & (g553) & (!g1128) & (!g1129) & (!g1136) & (!g1154)) + ((g515) & (g553) & (g1128) & (!g1129) & (!g1136) & (g1154)) + ((g515) & (g553) & (g1128) & (!g1129) & (g1136) & (!g1154)) + ((g515) & (g553) & (g1128) & (!g1129) & (g1136) & (g1154)) + ((g515) & (g553) & (g1128) & (g1129) & (!g1136) & (!g1154)) + ((g515) & (g553) & (g1128) & (g1129) & (!g1136) & (g1154)) + ((g515) & (g553) & (g1128) & (g1129) & (g1136) & (!g1154)) + ((g515) & (g553) & (g1128) & (g1129) & (g1136) & (g1154)));
	assign g1191 = (((!g553) & (!g1129) & (g1136) & (!g1154)) + ((!g553) & (g1129) & (!g1136) & (!g1154)) + ((!g553) & (g1129) & (!g1136) & (g1154)) + ((!g553) & (g1129) & (g1136) & (g1154)) + ((g553) & (!g1129) & (!g1136) & (!g1154)) + ((g553) & (g1129) & (!g1136) & (g1154)) + ((g553) & (g1129) & (g1136) & (!g1154)) + ((g553) & (g1129) & (g1136) & (g1154)));
	assign g1192 = (((!g604) & (!g645) & (!g1131) & (g1132) & (g1135) & (!g1154)) + ((!g604) & (!g645) & (g1131) & (!g1132) & (!g1135) & (!g1154)) + ((!g604) & (!g645) & (g1131) & (!g1132) & (!g1135) & (g1154)) + ((!g604) & (!g645) & (g1131) & (!g1132) & (g1135) & (!g1154)) + ((!g604) & (!g645) & (g1131) & (!g1132) & (g1135) & (g1154)) + ((!g604) & (!g645) & (g1131) & (g1132) & (!g1135) & (!g1154)) + ((!g604) & (!g645) & (g1131) & (g1132) & (!g1135) & (g1154)) + ((!g604) & (!g645) & (g1131) & (g1132) & (g1135) & (g1154)) + ((!g604) & (g645) & (!g1131) & (!g1132) & (g1135) & (!g1154)) + ((!g604) & (g645) & (!g1131) & (g1132) & (!g1135) & (!g1154)) + ((!g604) & (g645) & (!g1131) & (g1132) & (g1135) & (!g1154)) + ((!g604) & (g645) & (g1131) & (!g1132) & (!g1135) & (!g1154)) + ((!g604) & (g645) & (g1131) & (!g1132) & (!g1135) & (g1154)) + ((!g604) & (g645) & (g1131) & (!g1132) & (g1135) & (g1154)) + ((!g604) & (g645) & (g1131) & (g1132) & (!g1135) & (g1154)) + ((!g604) & (g645) & (g1131) & (g1132) & (g1135) & (g1154)) + ((g604) & (!g645) & (!g1131) & (!g1132) & (!g1135) & (!g1154)) + ((g604) & (!g645) & (!g1131) & (!g1132) & (g1135) & (!g1154)) + ((g604) & (!g645) & (!g1131) & (g1132) & (!g1135) & (!g1154)) + ((g604) & (!g645) & (g1131) & (!g1132) & (!g1135) & (g1154)) + ((g604) & (!g645) & (g1131) & (!g1132) & (g1135) & (g1154)) + ((g604) & (!g645) & (g1131) & (g1132) & (!g1135) & (g1154)) + ((g604) & (!g645) & (g1131) & (g1132) & (g1135) & (!g1154)) + ((g604) & (!g645) & (g1131) & (g1132) & (g1135) & (g1154)) + ((g604) & (g645) & (!g1131) & (!g1132) & (!g1135) & (!g1154)) + ((g604) & (g645) & (g1131) & (!g1132) & (!g1135) & (g1154)) + ((g604) & (g645) & (g1131) & (!g1132) & (g1135) & (!g1154)) + ((g604) & (g645) & (g1131) & (!g1132) & (g1135) & (g1154)) + ((g604) & (g645) & (g1131) & (g1132) & (!g1135) & (!g1154)) + ((g604) & (g645) & (g1131) & (g1132) & (!g1135) & (g1154)) + ((g604) & (g645) & (g1131) & (g1132) & (g1135) & (!g1154)) + ((g604) & (g645) & (g1131) & (g1132) & (g1135) & (g1154)));
	assign g1193 = (((!g645) & (!g1132) & (g1135) & (!g1154)) + ((!g645) & (g1132) & (!g1135) & (!g1154)) + ((!g645) & (g1132) & (!g1135) & (g1154)) + ((!g645) & (g1132) & (g1135) & (g1154)) + ((g645) & (!g1132) & (!g1135) & (!g1154)) + ((g645) & (g1132) & (!g1135) & (g1154)) + ((g645) & (g1132) & (g1135) & (!g1154)) + ((g645) & (g1132) & (g1135) & (g1154)));
	assign g1194 = (((!g700) & (!g744) & (!g1134) & (g1084) & (g1094) & (!g1154)) + ((!g700) & (!g744) & (g1134) & (!g1084) & (!g1094) & (!g1154)) + ((!g700) & (!g744) & (g1134) & (!g1084) & (!g1094) & (g1154)) + ((!g700) & (!g744) & (g1134) & (!g1084) & (g1094) & (!g1154)) + ((!g700) & (!g744) & (g1134) & (!g1084) & (g1094) & (g1154)) + ((!g700) & (!g744) & (g1134) & (g1084) & (!g1094) & (!g1154)) + ((!g700) & (!g744) & (g1134) & (g1084) & (!g1094) & (g1154)) + ((!g700) & (!g744) & (g1134) & (g1084) & (g1094) & (g1154)) + ((!g700) & (g744) & (!g1134) & (!g1084) & (g1094) & (!g1154)) + ((!g700) & (g744) & (!g1134) & (g1084) & (!g1094) & (!g1154)) + ((!g700) & (g744) & (!g1134) & (g1084) & (g1094) & (!g1154)) + ((!g700) & (g744) & (g1134) & (!g1084) & (!g1094) & (!g1154)) + ((!g700) & (g744) & (g1134) & (!g1084) & (!g1094) & (g1154)) + ((!g700) & (g744) & (g1134) & (!g1084) & (g1094) & (g1154)) + ((!g700) & (g744) & (g1134) & (g1084) & (!g1094) & (g1154)) + ((!g700) & (g744) & (g1134) & (g1084) & (g1094) & (g1154)) + ((g700) & (!g744) & (!g1134) & (!g1084) & (!g1094) & (!g1154)) + ((g700) & (!g744) & (!g1134) & (!g1084) & (g1094) & (!g1154)) + ((g700) & (!g744) & (!g1134) & (g1084) & (!g1094) & (!g1154)) + ((g700) & (!g744) & (g1134) & (!g1084) & (!g1094) & (g1154)) + ((g700) & (!g744) & (g1134) & (!g1084) & (g1094) & (g1154)) + ((g700) & (!g744) & (g1134) & (g1084) & (!g1094) & (g1154)) + ((g700) & (!g744) & (g1134) & (g1084) & (g1094) & (!g1154)) + ((g700) & (!g744) & (g1134) & (g1084) & (g1094) & (g1154)) + ((g700) & (g744) & (!g1134) & (!g1084) & (!g1094) & (!g1154)) + ((g700) & (g744) & (g1134) & (!g1084) & (!g1094) & (g1154)) + ((g700) & (g744) & (g1134) & (!g1084) & (g1094) & (!g1154)) + ((g700) & (g744) & (g1134) & (!g1084) & (g1094) & (g1154)) + ((g700) & (g744) & (g1134) & (g1084) & (!g1094) & (!g1154)) + ((g700) & (g744) & (g1134) & (g1084) & (!g1094) & (g1154)) + ((g700) & (g744) & (g1134) & (g1084) & (g1094) & (!g1154)) + ((g700) & (g744) & (g1134) & (g1084) & (g1094) & (g1154)));
	assign g1195 = (((!g645) & (!g700) & (g1194) & (g1155) & (g1167)) + ((!g645) & (g700) & (g1194) & (!g1155) & (g1167)) + ((!g645) & (g700) & (g1194) & (g1155) & (!g1167)) + ((!g645) & (g700) & (g1194) & (g1155) & (g1167)) + ((g645) & (!g700) & (!g1194) & (g1155) & (g1167)) + ((g645) & (!g700) & (g1194) & (!g1155) & (!g1167)) + ((g645) & (!g700) & (g1194) & (!g1155) & (g1167)) + ((g645) & (!g700) & (g1194) & (g1155) & (!g1167)) + ((g645) & (!g700) & (g1194) & (g1155) & (g1167)) + ((g645) & (g700) & (!g1194) & (!g1155) & (g1167)) + ((g645) & (g700) & (!g1194) & (g1155) & (!g1167)) + ((g645) & (g700) & (!g1194) & (g1155) & (g1167)) + ((g645) & (g700) & (g1194) & (!g1155) & (!g1167)) + ((g645) & (g700) & (g1194) & (!g1155) & (g1167)) + ((g645) & (g700) & (g1194) & (g1155) & (!g1167)) + ((g645) & (g700) & (g1194) & (g1155) & (g1167)));
	assign g1196 = (((!g553) & (!g604) & (g1192) & (g1193) & (g1195)) + ((!g553) & (g604) & (g1192) & (!g1193) & (g1195)) + ((!g553) & (g604) & (g1192) & (g1193) & (!g1195)) + ((!g553) & (g604) & (g1192) & (g1193) & (g1195)) + ((g553) & (!g604) & (!g1192) & (g1193) & (g1195)) + ((g553) & (!g604) & (g1192) & (!g1193) & (!g1195)) + ((g553) & (!g604) & (g1192) & (!g1193) & (g1195)) + ((g553) & (!g604) & (g1192) & (g1193) & (!g1195)) + ((g553) & (!g604) & (g1192) & (g1193) & (g1195)) + ((g553) & (g604) & (!g1192) & (!g1193) & (g1195)) + ((g553) & (g604) & (!g1192) & (g1193) & (!g1195)) + ((g553) & (g604) & (!g1192) & (g1193) & (g1195)) + ((g553) & (g604) & (g1192) & (!g1193) & (!g1195)) + ((g553) & (g604) & (g1192) & (!g1193) & (g1195)) + ((g553) & (g604) & (g1192) & (g1193) & (!g1195)) + ((g553) & (g604) & (g1192) & (g1193) & (g1195)));
	assign g1197 = (((!g468) & (!g515) & (g1190) & (g1191) & (g1196)) + ((!g468) & (g515) & (g1190) & (!g1191) & (g1196)) + ((!g468) & (g515) & (g1190) & (g1191) & (!g1196)) + ((!g468) & (g515) & (g1190) & (g1191) & (g1196)) + ((g468) & (!g515) & (!g1190) & (g1191) & (g1196)) + ((g468) & (!g515) & (g1190) & (!g1191) & (!g1196)) + ((g468) & (!g515) & (g1190) & (!g1191) & (g1196)) + ((g468) & (!g515) & (g1190) & (g1191) & (!g1196)) + ((g468) & (!g515) & (g1190) & (g1191) & (g1196)) + ((g468) & (g515) & (!g1190) & (!g1191) & (g1196)) + ((g468) & (g515) & (!g1190) & (g1191) & (!g1196)) + ((g468) & (g515) & (!g1190) & (g1191) & (g1196)) + ((g468) & (g515) & (g1190) & (!g1191) & (!g1196)) + ((g468) & (g515) & (g1190) & (!g1191) & (g1196)) + ((g468) & (g515) & (g1190) & (g1191) & (!g1196)) + ((g468) & (g515) & (g1190) & (g1191) & (g1196)));
	assign g1198 = (((!g390) & (!g433) & (g1188) & (g1189) & (g1197)) + ((!g390) & (g433) & (g1188) & (!g1189) & (g1197)) + ((!g390) & (g433) & (g1188) & (g1189) & (!g1197)) + ((!g390) & (g433) & (g1188) & (g1189) & (g1197)) + ((g390) & (!g433) & (!g1188) & (g1189) & (g1197)) + ((g390) & (!g433) & (g1188) & (!g1189) & (!g1197)) + ((g390) & (!g433) & (g1188) & (!g1189) & (g1197)) + ((g390) & (!g433) & (g1188) & (g1189) & (!g1197)) + ((g390) & (!g433) & (g1188) & (g1189) & (g1197)) + ((g390) & (g433) & (!g1188) & (!g1189) & (g1197)) + ((g390) & (g433) & (!g1188) & (g1189) & (!g1197)) + ((g390) & (g433) & (!g1188) & (g1189) & (g1197)) + ((g390) & (g433) & (g1188) & (!g1189) & (!g1197)) + ((g390) & (g433) & (g1188) & (!g1189) & (g1197)) + ((g390) & (g433) & (g1188) & (g1189) & (!g1197)) + ((g390) & (g433) & (g1188) & (g1189) & (g1197)));
	assign g1199 = (((!g319) & (!g358) & (g1186) & (g1187) & (g1198)) + ((!g319) & (g358) & (g1186) & (!g1187) & (g1198)) + ((!g319) & (g358) & (g1186) & (g1187) & (!g1198)) + ((!g319) & (g358) & (g1186) & (g1187) & (g1198)) + ((g319) & (!g358) & (!g1186) & (g1187) & (g1198)) + ((g319) & (!g358) & (g1186) & (!g1187) & (!g1198)) + ((g319) & (!g358) & (g1186) & (!g1187) & (g1198)) + ((g319) & (!g358) & (g1186) & (g1187) & (!g1198)) + ((g319) & (!g358) & (g1186) & (g1187) & (g1198)) + ((g319) & (g358) & (!g1186) & (!g1187) & (g1198)) + ((g319) & (g358) & (!g1186) & (g1187) & (!g1198)) + ((g319) & (g358) & (!g1186) & (g1187) & (g1198)) + ((g319) & (g358) & (g1186) & (!g1187) & (!g1198)) + ((g319) & (g358) & (g1186) & (!g1187) & (g1198)) + ((g319) & (g358) & (g1186) & (g1187) & (!g1198)) + ((g319) & (g358) & (g1186) & (g1187) & (g1198)));
	assign g1200 = (((!g255) & (!g290) & (g1184) & (g1185) & (g1199)) + ((!g255) & (g290) & (g1184) & (!g1185) & (g1199)) + ((!g255) & (g290) & (g1184) & (g1185) & (!g1199)) + ((!g255) & (g290) & (g1184) & (g1185) & (g1199)) + ((g255) & (!g290) & (!g1184) & (g1185) & (g1199)) + ((g255) & (!g290) & (g1184) & (!g1185) & (!g1199)) + ((g255) & (!g290) & (g1184) & (!g1185) & (g1199)) + ((g255) & (!g290) & (g1184) & (g1185) & (!g1199)) + ((g255) & (!g290) & (g1184) & (g1185) & (g1199)) + ((g255) & (g290) & (!g1184) & (!g1185) & (g1199)) + ((g255) & (g290) & (!g1184) & (g1185) & (!g1199)) + ((g255) & (g290) & (!g1184) & (g1185) & (g1199)) + ((g255) & (g290) & (g1184) & (!g1185) & (!g1199)) + ((g255) & (g290) & (g1184) & (!g1185) & (g1199)) + ((g255) & (g290) & (g1184) & (g1185) & (!g1199)) + ((g255) & (g290) & (g1184) & (g1185) & (g1199)));
	assign g1201 = (((!g198) & (!g229) & (g1182) & (g1183) & (g1200)) + ((!g198) & (g229) & (g1182) & (!g1183) & (g1200)) + ((!g198) & (g229) & (g1182) & (g1183) & (!g1200)) + ((!g198) & (g229) & (g1182) & (g1183) & (g1200)) + ((g198) & (!g229) & (!g1182) & (g1183) & (g1200)) + ((g198) & (!g229) & (g1182) & (!g1183) & (!g1200)) + ((g198) & (!g229) & (g1182) & (!g1183) & (g1200)) + ((g198) & (!g229) & (g1182) & (g1183) & (!g1200)) + ((g198) & (!g229) & (g1182) & (g1183) & (g1200)) + ((g198) & (g229) & (!g1182) & (!g1183) & (g1200)) + ((g198) & (g229) & (!g1182) & (g1183) & (!g1200)) + ((g198) & (g229) & (!g1182) & (g1183) & (g1200)) + ((g198) & (g229) & (g1182) & (!g1183) & (!g1200)) + ((g198) & (g229) & (g1182) & (!g1183) & (g1200)) + ((g198) & (g229) & (g1182) & (g1183) & (!g1200)) + ((g198) & (g229) & (g1182) & (g1183) & (g1200)));
	assign g1202 = (((!g147) & (!g174) & (g1180) & (g1181) & (g1201)) + ((!g147) & (g174) & (g1180) & (!g1181) & (g1201)) + ((!g147) & (g174) & (g1180) & (g1181) & (!g1201)) + ((!g147) & (g174) & (g1180) & (g1181) & (g1201)) + ((g147) & (!g174) & (!g1180) & (g1181) & (g1201)) + ((g147) & (!g174) & (g1180) & (!g1181) & (!g1201)) + ((g147) & (!g174) & (g1180) & (!g1181) & (g1201)) + ((g147) & (!g174) & (g1180) & (g1181) & (!g1201)) + ((g147) & (!g174) & (g1180) & (g1181) & (g1201)) + ((g147) & (g174) & (!g1180) & (!g1181) & (g1201)) + ((g147) & (g174) & (!g1180) & (g1181) & (!g1201)) + ((g147) & (g174) & (!g1180) & (g1181) & (g1201)) + ((g147) & (g174) & (g1180) & (!g1181) & (!g1201)) + ((g147) & (g174) & (g1180) & (!g1181) & (g1201)) + ((g147) & (g174) & (g1180) & (g1181) & (!g1201)) + ((g147) & (g174) & (g1180) & (g1181) & (g1201)));
	assign g1203 = (((!g104) & (!g127) & (g1178) & (g1179) & (g1202)) + ((!g104) & (g127) & (g1178) & (!g1179) & (g1202)) + ((!g104) & (g127) & (g1178) & (g1179) & (!g1202)) + ((!g104) & (g127) & (g1178) & (g1179) & (g1202)) + ((g104) & (!g127) & (!g1178) & (g1179) & (g1202)) + ((g104) & (!g127) & (g1178) & (!g1179) & (!g1202)) + ((g104) & (!g127) & (g1178) & (!g1179) & (g1202)) + ((g104) & (!g127) & (g1178) & (g1179) & (!g1202)) + ((g104) & (!g127) & (g1178) & (g1179) & (g1202)) + ((g104) & (g127) & (!g1178) & (!g1179) & (g1202)) + ((g104) & (g127) & (!g1178) & (g1179) & (!g1202)) + ((g104) & (g127) & (!g1178) & (g1179) & (g1202)) + ((g104) & (g127) & (g1178) & (!g1179) & (!g1202)) + ((g104) & (g127) & (g1178) & (!g1179) & (g1202)) + ((g104) & (g127) & (g1178) & (g1179) & (!g1202)) + ((g104) & (g127) & (g1178) & (g1179) & (g1202)));
	assign g1204 = (((!g68) & (!g87) & (g1176) & (g1177) & (g1203)) + ((!g68) & (g87) & (g1176) & (!g1177) & (g1203)) + ((!g68) & (g87) & (g1176) & (g1177) & (!g1203)) + ((!g68) & (g87) & (g1176) & (g1177) & (g1203)) + ((g68) & (!g87) & (!g1176) & (g1177) & (g1203)) + ((g68) & (!g87) & (g1176) & (!g1177) & (!g1203)) + ((g68) & (!g87) & (g1176) & (!g1177) & (g1203)) + ((g68) & (!g87) & (g1176) & (g1177) & (!g1203)) + ((g68) & (!g87) & (g1176) & (g1177) & (g1203)) + ((g68) & (g87) & (!g1176) & (!g1177) & (g1203)) + ((g68) & (g87) & (!g1176) & (g1177) & (!g1203)) + ((g68) & (g87) & (!g1176) & (g1177) & (g1203)) + ((g68) & (g87) & (g1176) & (!g1177) & (!g1203)) + ((g68) & (g87) & (g1176) & (!g1177) & (g1203)) + ((g68) & (g87) & (g1176) & (g1177) & (!g1203)) + ((g68) & (g87) & (g1176) & (g1177) & (g1203)));
	assign g1205 = (((!g39) & (!g54) & (g1174) & (g1175) & (g1204)) + ((!g39) & (g54) & (g1174) & (!g1175) & (g1204)) + ((!g39) & (g54) & (g1174) & (g1175) & (!g1204)) + ((!g39) & (g54) & (g1174) & (g1175) & (g1204)) + ((g39) & (!g54) & (!g1174) & (g1175) & (g1204)) + ((g39) & (!g54) & (g1174) & (!g1175) & (!g1204)) + ((g39) & (!g54) & (g1174) & (!g1175) & (g1204)) + ((g39) & (!g54) & (g1174) & (g1175) & (!g1204)) + ((g39) & (!g54) & (g1174) & (g1175) & (g1204)) + ((g39) & (g54) & (!g1174) & (!g1175) & (g1204)) + ((g39) & (g54) & (!g1174) & (g1175) & (!g1204)) + ((g39) & (g54) & (!g1174) & (g1175) & (g1204)) + ((g39) & (g54) & (g1174) & (!g1175) & (!g1204)) + ((g39) & (g54) & (g1174) & (!g1175) & (g1204)) + ((g39) & (g54) & (g1174) & (g1175) & (!g1204)) + ((g39) & (g54) & (g1174) & (g1175) & (g1204)));
	assign g1206 = (((!g18) & (!g27) & (g1172) & (g1173) & (g1205)) + ((!g18) & (g27) & (g1172) & (!g1173) & (g1205)) + ((!g18) & (g27) & (g1172) & (g1173) & (!g1205)) + ((!g18) & (g27) & (g1172) & (g1173) & (g1205)) + ((g18) & (!g27) & (!g1172) & (g1173) & (g1205)) + ((g18) & (!g27) & (g1172) & (!g1173) & (!g1205)) + ((g18) & (!g27) & (g1172) & (!g1173) & (g1205)) + ((g18) & (!g27) & (g1172) & (g1173) & (!g1205)) + ((g18) & (!g27) & (g1172) & (g1173) & (g1205)) + ((g18) & (g27) & (!g1172) & (!g1173) & (g1205)) + ((g18) & (g27) & (!g1172) & (g1173) & (!g1205)) + ((g18) & (g27) & (!g1172) & (g1173) & (g1205)) + ((g18) & (g27) & (g1172) & (!g1173) & (!g1205)) + ((g18) & (g27) & (g1172) & (!g1173) & (g1205)) + ((g18) & (g27) & (g1172) & (g1173) & (!g1205)) + ((g18) & (g27) & (g1172) & (g1173) & (g1205)));
	assign g1207 = (((!g2) & (!g8) & (g1170) & (g1171) & (g1206)) + ((!g2) & (g8) & (g1170) & (!g1171) & (g1206)) + ((!g2) & (g8) & (g1170) & (g1171) & (!g1206)) + ((!g2) & (g8) & (g1170) & (g1171) & (g1206)) + ((g2) & (!g8) & (!g1170) & (g1171) & (g1206)) + ((g2) & (!g8) & (g1170) & (!g1171) & (!g1206)) + ((g2) & (!g8) & (g1170) & (!g1171) & (g1206)) + ((g2) & (!g8) & (g1170) & (g1171) & (!g1206)) + ((g2) & (!g8) & (g1170) & (g1171) & (g1206)) + ((g2) & (g8) & (!g1170) & (!g1171) & (g1206)) + ((g2) & (g8) & (!g1170) & (g1171) & (!g1206)) + ((g2) & (g8) & (!g1170) & (g1171) & (g1206)) + ((g2) & (g8) & (g1170) & (!g1171) & (!g1206)) + ((g2) & (g8) & (g1170) & (!g1171) & (g1206)) + ((g2) & (g8) & (g1170) & (g1171) & (!g1206)) + ((g2) & (g8) & (g1170) & (g1171) & (g1206)));
	assign g1208 = (((!g2) & (!g1096) & (g1147) & (!g1154)) + ((!g2) & (g1096) & (!g1147) & (!g1154)) + ((!g2) & (g1096) & (!g1147) & (g1154)) + ((!g2) & (g1096) & (g1147) & (g1154)) + ((g2) & (!g1096) & (!g1147) & (!g1154)) + ((g2) & (g1096) & (!g1147) & (g1154)) + ((g2) & (g1096) & (g1147) & (!g1154)) + ((g2) & (g1096) & (g1147) & (g1154)));
	assign g1209 = (((!g1) & (!g1095) & (!g1150) & (!g1152) & (g1153)) + ((!g1) & (!g1095) & (!g1150) & (g1152) & (!g1153)) + ((!g1) & (!g1095) & (!g1150) & (g1152) & (g1153)) + ((!g1) & (g1095) & (g1150) & (!g1152) & (!g1153)) + ((!g1) & (g1095) & (g1150) & (!g1152) & (g1153)) + ((!g1) & (g1095) & (g1150) & (g1152) & (!g1153)) + ((!g1) & (g1095) & (g1150) & (g1152) & (g1153)) + ((g1) & (!g1095) & (!g1150) & (!g1152) & (g1153)) + ((g1) & (!g1095) & (!g1150) & (g1152) & (g1153)) + ((g1) & (g1095) & (g1150) & (!g1152) & (!g1153)) + ((g1) & (g1095) & (g1150) & (!g1152) & (g1153)) + ((g1) & (g1095) & (g1150) & (g1152) & (!g1153)) + ((g1) & (g1095) & (g1150) & (g1152) & (g1153)));
	assign g1210 = (((!g4) & (!g1) & (!g1169) & (!g1207) & (!g1208) & (!g1209)) + ((!g4) & (g1) & (!g1169) & (!g1207) & (!g1208) & (!g1209)) + ((!g4) & (g1) & (!g1169) & (!g1207) & (!g1208) & (g1209)) + ((!g4) & (g1) & (!g1169) & (!g1207) & (g1208) & (!g1209)) + ((!g4) & (g1) & (!g1169) & (!g1207) & (g1208) & (g1209)) + ((!g4) & (g1) & (!g1169) & (g1207) & (!g1208) & (!g1209)) + ((!g4) & (g1) & (!g1169) & (g1207) & (!g1208) & (g1209)) + ((!g4) & (g1) & (!g1169) & (g1207) & (g1208) & (!g1209)) + ((!g4) & (g1) & (!g1169) & (g1207) & (g1208) & (g1209)) + ((!g4) & (g1) & (g1169) & (!g1207) & (!g1208) & (!g1209)) + ((!g4) & (g1) & (g1169) & (!g1207) & (!g1208) & (g1209)) + ((g4) & (!g1) & (!g1169) & (!g1207) & (!g1208) & (!g1209)) + ((g4) & (!g1) & (!g1169) & (!g1207) & (g1208) & (!g1209)) + ((g4) & (!g1) & (!g1169) & (g1207) & (!g1208) & (!g1209)) + ((g4) & (g1) & (!g1169) & (!g1207) & (!g1208) & (!g1209)) + ((g4) & (g1) & (!g1169) & (!g1207) & (!g1208) & (g1209)) + ((g4) & (g1) & (!g1169) & (!g1207) & (g1208) & (!g1209)) + ((g4) & (g1) & (!g1169) & (!g1207) & (g1208) & (g1209)) + ((g4) & (g1) & (!g1169) & (g1207) & (!g1208) & (!g1209)) + ((g4) & (g1) & (!g1169) & (g1207) & (!g1208) & (g1209)) + ((g4) & (g1) & (!g1169) & (g1207) & (g1208) & (!g1209)) + ((g4) & (g1) & (!g1169) & (g1207) & (g1208) & (g1209)) + ((g4) & (g1) & (g1169) & (!g1207) & (!g1208) & (!g1209)) + ((g4) & (g1) & (g1169) & (!g1207) & (!g1208) & (g1209)) + ((g4) & (g1) & (g1169) & (!g1207) & (g1208) & (!g1209)) + ((g4) & (g1) & (g1169) & (!g1207) & (g1208) & (g1209)) + ((g4) & (g1) & (g1169) & (g1207) & (!g1208) & (!g1209)) + ((g4) & (g1) & (g1169) & (g1207) & (!g1208) & (g1209)));
	assign g1211 = (((!g700) & (!g1155) & (g1167) & (!g1168) & (!g1210)) + ((!g700) & (!g1155) & (g1167) & (g1168) & (!g1210)) + ((!g700) & (!g1155) & (g1167) & (g1168) & (g1210)) + ((!g700) & (g1155) & (!g1167) & (!g1168) & (!g1210)) + ((!g700) & (g1155) & (!g1167) & (!g1168) & (g1210)) + ((!g700) & (g1155) & (!g1167) & (g1168) & (!g1210)) + ((!g700) & (g1155) & (!g1167) & (g1168) & (g1210)) + ((!g700) & (g1155) & (g1167) & (!g1168) & (g1210)) + ((g700) & (!g1155) & (!g1167) & (!g1168) & (!g1210)) + ((g700) & (!g1155) & (!g1167) & (g1168) & (!g1210)) + ((g700) & (!g1155) & (!g1167) & (g1168) & (g1210)) + ((g700) & (g1155) & (!g1167) & (!g1168) & (g1210)) + ((g700) & (g1155) & (g1167) & (!g1168) & (!g1210)) + ((g700) & (g1155) & (g1167) & (!g1168) & (g1210)) + ((g700) & (g1155) & (g1167) & (g1168) & (!g1210)) + ((g700) & (g1155) & (g1167) & (g1168) & (g1210)));
	assign g1212 = (((!g744) & (!g803) & (g1157) & (g1166)) + ((!g744) & (g803) & (!g1157) & (g1166)) + ((!g744) & (g803) & (g1157) & (!g1166)) + ((!g744) & (g803) & (g1157) & (g1166)) + ((g744) & (!g803) & (!g1157) & (!g1166)) + ((g744) & (!g803) & (!g1157) & (g1166)) + ((g744) & (!g803) & (g1157) & (!g1166)) + ((g744) & (g803) & (!g1157) & (!g1166)));
	assign g1213 = (((!g1156) & (!g1168) & (!g1210) & (g1212)) + ((!g1156) & (g1168) & (!g1210) & (g1212)) + ((!g1156) & (g1168) & (g1210) & (g1212)) + ((g1156) & (!g1168) & (!g1210) & (!g1212)) + ((g1156) & (!g1168) & (g1210) & (!g1212)) + ((g1156) & (!g1168) & (g1210) & (g1212)) + ((g1156) & (g1168) & (!g1210) & (!g1212)) + ((g1156) & (g1168) & (g1210) & (!g1212)));
	assign g1214 = (((!g803) & (!g1157) & (g1166) & (!g1168) & (!g1210)) + ((!g803) & (!g1157) & (g1166) & (g1168) & (!g1210)) + ((!g803) & (!g1157) & (g1166) & (g1168) & (g1210)) + ((!g803) & (g1157) & (!g1166) & (!g1168) & (!g1210)) + ((!g803) & (g1157) & (!g1166) & (!g1168) & (g1210)) + ((!g803) & (g1157) & (!g1166) & (g1168) & (!g1210)) + ((!g803) & (g1157) & (!g1166) & (g1168) & (g1210)) + ((!g803) & (g1157) & (g1166) & (!g1168) & (g1210)) + ((g803) & (!g1157) & (!g1166) & (!g1168) & (!g1210)) + ((g803) & (!g1157) & (!g1166) & (g1168) & (!g1210)) + ((g803) & (!g1157) & (!g1166) & (g1168) & (g1210)) + ((g803) & (g1157) & (!g1166) & (!g1168) & (g1210)) + ((g803) & (g1157) & (g1166) & (!g1168) & (!g1210)) + ((g803) & (g1157) & (g1166) & (!g1168) & (g1210)) + ((g803) & (g1157) & (g1166) & (g1168) & (!g1210)) + ((g803) & (g1157) & (g1166) & (g1168) & (g1210)));
	assign g1215 = (((!g851) & (!g914) & (g1159) & (g1165)) + ((!g851) & (g914) & (!g1159) & (g1165)) + ((!g851) & (g914) & (g1159) & (!g1165)) + ((!g851) & (g914) & (g1159) & (g1165)) + ((g851) & (!g914) & (!g1159) & (!g1165)) + ((g851) & (!g914) & (!g1159) & (g1165)) + ((g851) & (!g914) & (g1159) & (!g1165)) + ((g851) & (g914) & (!g1159) & (!g1165)));
	assign g1216 = (((!g1158) & (!g1168) & (!g1210) & (g1215)) + ((!g1158) & (g1168) & (!g1210) & (g1215)) + ((!g1158) & (g1168) & (g1210) & (g1215)) + ((g1158) & (!g1168) & (!g1210) & (!g1215)) + ((g1158) & (!g1168) & (g1210) & (!g1215)) + ((g1158) & (!g1168) & (g1210) & (g1215)) + ((g1158) & (g1168) & (!g1210) & (!g1215)) + ((g1158) & (g1168) & (g1210) & (!g1215)));
	assign g1217 = (((!g914) & (!g1159) & (g1165) & (!g1168) & (!g1210)) + ((!g914) & (!g1159) & (g1165) & (g1168) & (!g1210)) + ((!g914) & (!g1159) & (g1165) & (g1168) & (g1210)) + ((!g914) & (g1159) & (!g1165) & (!g1168) & (!g1210)) + ((!g914) & (g1159) & (!g1165) & (!g1168) & (g1210)) + ((!g914) & (g1159) & (!g1165) & (g1168) & (!g1210)) + ((!g914) & (g1159) & (!g1165) & (g1168) & (g1210)) + ((!g914) & (g1159) & (g1165) & (!g1168) & (g1210)) + ((g914) & (!g1159) & (!g1165) & (!g1168) & (!g1210)) + ((g914) & (!g1159) & (!g1165) & (g1168) & (!g1210)) + ((g914) & (!g1159) & (!g1165) & (g1168) & (g1210)) + ((g914) & (g1159) & (!g1165) & (!g1168) & (g1210)) + ((g914) & (g1159) & (g1165) & (!g1168) & (!g1210)) + ((g914) & (g1159) & (g1165) & (!g1168) & (g1210)) + ((g914) & (g1159) & (g1165) & (g1168) & (!g1210)) + ((g914) & (g1159) & (g1165) & (g1168) & (g1210)));
	assign g1218 = (((!g1032) & (!g1030) & (g1162) & (g1164)) + ((!g1032) & (g1030) & (!g1162) & (g1164)) + ((!g1032) & (g1030) & (g1162) & (!g1164)) + ((!g1032) & (g1030) & (g1162) & (g1164)) + ((g1032) & (!g1030) & (!g1162) & (!g1164)) + ((g1032) & (!g1030) & (!g1162) & (g1164)) + ((g1032) & (!g1030) & (g1162) & (!g1164)) + ((g1032) & (g1030) & (!g1162) & (!g1164)));
	assign g1219 = (((!g1161) & (!g1168) & (!g1210) & (g1218)) + ((!g1161) & (g1168) & (!g1210) & (g1218)) + ((!g1161) & (g1168) & (g1210) & (g1218)) + ((g1161) & (!g1168) & (!g1210) & (!g1218)) + ((g1161) & (!g1168) & (g1210) & (!g1218)) + ((g1161) & (!g1168) & (g1210) & (g1218)) + ((g1161) & (g1168) & (!g1210) & (!g1218)) + ((g1161) & (g1168) & (g1210) & (!g1218)));
	assign g1220 = (((!g1030) & (!g1162) & (g1164) & (!g1168) & (!g1210)) + ((!g1030) & (!g1162) & (g1164) & (g1168) & (!g1210)) + ((!g1030) & (!g1162) & (g1164) & (g1168) & (g1210)) + ((!g1030) & (g1162) & (!g1164) & (!g1168) & (!g1210)) + ((!g1030) & (g1162) & (!g1164) & (!g1168) & (g1210)) + ((!g1030) & (g1162) & (!g1164) & (g1168) & (!g1210)) + ((!g1030) & (g1162) & (!g1164) & (g1168) & (g1210)) + ((!g1030) & (g1162) & (g1164) & (!g1168) & (g1210)) + ((g1030) & (!g1162) & (!g1164) & (!g1168) & (!g1210)) + ((g1030) & (!g1162) & (!g1164) & (g1168) & (!g1210)) + ((g1030) & (!g1162) & (!g1164) & (g1168) & (g1210)) + ((g1030) & (g1162) & (!g1164) & (!g1168) & (g1210)) + ((g1030) & (g1162) & (g1164) & (!g1168) & (!g1210)) + ((g1030) & (g1162) & (g1164) & (!g1168) & (g1210)) + ((g1030) & (g1162) & (g1164) & (g1168) & (!g1210)) + ((g1030) & (g1162) & (g1164) & (g1168) & (g1210)));
	assign g1221 = (((!g1160) & (!ax56x) & (!g1154) & (g1163)) + ((!g1160) & (!ax56x) & (g1154) & (g1163)) + ((!g1160) & (ax56x) & (!g1154) & (!g1163)) + ((!g1160) & (ax56x) & (!g1154) & (g1163)) + ((g1160) & (!ax56x) & (!g1154) & (!g1163)) + ((g1160) & (!ax56x) & (g1154) & (!g1163)) + ((g1160) & (ax56x) & (g1154) & (!g1163)) + ((g1160) & (ax56x) & (g1154) & (g1163)));
	assign g1222 = (((!ax56x) & (!ax57x) & (!g1154) & (!g1168) & (!g1210) & (g1221)) + ((!ax56x) & (!ax57x) & (!g1154) & (!g1168) & (g1210) & (!g1221)) + ((!ax56x) & (!ax57x) & (!g1154) & (!g1168) & (g1210) & (g1221)) + ((!ax56x) & (!ax57x) & (!g1154) & (g1168) & (!g1210) & (g1221)) + ((!ax56x) & (!ax57x) & (!g1154) & (g1168) & (g1210) & (g1221)) + ((!ax56x) & (!ax57x) & (g1154) & (!g1168) & (!g1210) & (!g1221)) + ((!ax56x) & (!ax57x) & (g1154) & (g1168) & (!g1210) & (!g1221)) + ((!ax56x) & (!ax57x) & (g1154) & (g1168) & (g1210) & (!g1221)) + ((!ax56x) & (ax57x) & (!g1154) & (!g1168) & (!g1210) & (!g1221)) + ((!ax56x) & (ax57x) & (!g1154) & (g1168) & (!g1210) & (!g1221)) + ((!ax56x) & (ax57x) & (!g1154) & (g1168) & (g1210) & (!g1221)) + ((!ax56x) & (ax57x) & (g1154) & (!g1168) & (!g1210) & (g1221)) + ((!ax56x) & (ax57x) & (g1154) & (!g1168) & (g1210) & (!g1221)) + ((!ax56x) & (ax57x) & (g1154) & (!g1168) & (g1210) & (g1221)) + ((!ax56x) & (ax57x) & (g1154) & (g1168) & (!g1210) & (g1221)) + ((!ax56x) & (ax57x) & (g1154) & (g1168) & (g1210) & (g1221)) + ((ax56x) & (!ax57x) & (!g1154) & (!g1168) & (!g1210) & (!g1221)) + ((ax56x) & (!ax57x) & (!g1154) & (g1168) & (!g1210) & (!g1221)) + ((ax56x) & (!ax57x) & (!g1154) & (g1168) & (g1210) & (!g1221)) + ((ax56x) & (!ax57x) & (g1154) & (!g1168) & (!g1210) & (!g1221)) + ((ax56x) & (!ax57x) & (g1154) & (g1168) & (!g1210) & (!g1221)) + ((ax56x) & (!ax57x) & (g1154) & (g1168) & (g1210) & (!g1221)) + ((ax56x) & (ax57x) & (!g1154) & (!g1168) & (!g1210) & (g1221)) + ((ax56x) & (ax57x) & (!g1154) & (!g1168) & (g1210) & (!g1221)) + ((ax56x) & (ax57x) & (!g1154) & (!g1168) & (g1210) & (g1221)) + ((ax56x) & (ax57x) & (!g1154) & (g1168) & (!g1210) & (g1221)) + ((ax56x) & (ax57x) & (!g1154) & (g1168) & (g1210) & (g1221)) + ((ax56x) & (ax57x) & (g1154) & (!g1168) & (!g1210) & (g1221)) + ((ax56x) & (ax57x) & (g1154) & (!g1168) & (g1210) & (!g1221)) + ((ax56x) & (ax57x) & (g1154) & (!g1168) & (g1210) & (g1221)) + ((ax56x) & (ax57x) & (g1154) & (g1168) & (!g1210) & (g1221)) + ((ax56x) & (ax57x) & (g1154) & (g1168) & (g1210) & (g1221)));
	assign g1223 = (((!ax56x) & (!g1154) & (!g1163) & (!g1168) & (g1210)) + ((!ax56x) & (!g1154) & (g1163) & (!g1168) & (!g1210)) + ((!ax56x) & (!g1154) & (g1163) & (!g1168) & (g1210)) + ((!ax56x) & (!g1154) & (g1163) & (g1168) & (!g1210)) + ((!ax56x) & (!g1154) & (g1163) & (g1168) & (g1210)) + ((!ax56x) & (g1154) & (g1163) & (!g1168) & (!g1210)) + ((!ax56x) & (g1154) & (g1163) & (g1168) & (!g1210)) + ((!ax56x) & (g1154) & (g1163) & (g1168) & (g1210)) + ((ax56x) & (!g1154) & (!g1163) & (!g1168) & (!g1210)) + ((ax56x) & (!g1154) & (!g1163) & (g1168) & (!g1210)) + ((ax56x) & (!g1154) & (!g1163) & (g1168) & (g1210)) + ((ax56x) & (g1154) & (!g1163) & (!g1168) & (!g1210)) + ((ax56x) & (g1154) & (!g1163) & (!g1168) & (g1210)) + ((ax56x) & (g1154) & (!g1163) & (g1168) & (!g1210)) + ((ax56x) & (g1154) & (!g1163) & (g1168) & (g1210)) + ((ax56x) & (g1154) & (g1163) & (!g1168) & (g1210)));
	assign g1224 = (((!ax52x) & (!ax53x)));
	assign g1225 = (((!g1154) & (!ax54x) & (!ax55x) & (!g1168) & (!g1210) & (!g1224)) + ((!g1154) & (!ax54x) & (!ax55x) & (g1168) & (!g1210) & (!g1224)) + ((!g1154) & (!ax54x) & (!ax55x) & (g1168) & (g1210) & (!g1224)) + ((!g1154) & (!ax54x) & (ax55x) & (!g1168) & (g1210) & (!g1224)) + ((!g1154) & (ax54x) & (ax55x) & (!g1168) & (g1210) & (!g1224)) + ((!g1154) & (ax54x) & (ax55x) & (!g1168) & (g1210) & (g1224)) + ((g1154) & (!ax54x) & (!ax55x) & (!g1168) & (!g1210) & (!g1224)) + ((g1154) & (!ax54x) & (!ax55x) & (!g1168) & (!g1210) & (g1224)) + ((g1154) & (!ax54x) & (!ax55x) & (!g1168) & (g1210) & (!g1224)) + ((g1154) & (!ax54x) & (!ax55x) & (g1168) & (!g1210) & (!g1224)) + ((g1154) & (!ax54x) & (!ax55x) & (g1168) & (!g1210) & (g1224)) + ((g1154) & (!ax54x) & (!ax55x) & (g1168) & (g1210) & (!g1224)) + ((g1154) & (!ax54x) & (!ax55x) & (g1168) & (g1210) & (g1224)) + ((g1154) & (!ax54x) & (ax55x) & (!g1168) & (!g1210) & (!g1224)) + ((g1154) & (!ax54x) & (ax55x) & (!g1168) & (g1210) & (!g1224)) + ((g1154) & (!ax54x) & (ax55x) & (!g1168) & (g1210) & (g1224)) + ((g1154) & (!ax54x) & (ax55x) & (g1168) & (!g1210) & (!g1224)) + ((g1154) & (!ax54x) & (ax55x) & (g1168) & (g1210) & (!g1224)) + ((g1154) & (ax54x) & (!ax55x) & (!g1168) & (g1210) & (!g1224)) + ((g1154) & (ax54x) & (!ax55x) & (!g1168) & (g1210) & (g1224)) + ((g1154) & (ax54x) & (ax55x) & (!g1168) & (!g1210) & (!g1224)) + ((g1154) & (ax54x) & (ax55x) & (!g1168) & (!g1210) & (g1224)) + ((g1154) & (ax54x) & (ax55x) & (!g1168) & (g1210) & (!g1224)) + ((g1154) & (ax54x) & (ax55x) & (!g1168) & (g1210) & (g1224)) + ((g1154) & (ax54x) & (ax55x) & (g1168) & (!g1210) & (!g1224)) + ((g1154) & (ax54x) & (ax55x) & (g1168) & (!g1210) & (g1224)) + ((g1154) & (ax54x) & (ax55x) & (g1168) & (g1210) & (!g1224)) + ((g1154) & (ax54x) & (ax55x) & (g1168) & (g1210) & (g1224)));
	assign g1226 = (((!g1030) & (!g1160) & (g1222) & (g1223) & (g1225)) + ((!g1030) & (g1160) & (g1222) & (!g1223) & (g1225)) + ((!g1030) & (g1160) & (g1222) & (g1223) & (!g1225)) + ((!g1030) & (g1160) & (g1222) & (g1223) & (g1225)) + ((g1030) & (!g1160) & (!g1222) & (g1223) & (g1225)) + ((g1030) & (!g1160) & (g1222) & (!g1223) & (!g1225)) + ((g1030) & (!g1160) & (g1222) & (!g1223) & (g1225)) + ((g1030) & (!g1160) & (g1222) & (g1223) & (!g1225)) + ((g1030) & (!g1160) & (g1222) & (g1223) & (g1225)) + ((g1030) & (g1160) & (!g1222) & (!g1223) & (g1225)) + ((g1030) & (g1160) & (!g1222) & (g1223) & (!g1225)) + ((g1030) & (g1160) & (!g1222) & (g1223) & (g1225)) + ((g1030) & (g1160) & (g1222) & (!g1223) & (!g1225)) + ((g1030) & (g1160) & (g1222) & (!g1223) & (g1225)) + ((g1030) & (g1160) & (g1222) & (g1223) & (!g1225)) + ((g1030) & (g1160) & (g1222) & (g1223) & (g1225)));
	assign g1227 = (((!g914) & (!g1032) & (g1219) & (g1220) & (g1226)) + ((!g914) & (g1032) & (g1219) & (!g1220) & (g1226)) + ((!g914) & (g1032) & (g1219) & (g1220) & (!g1226)) + ((!g914) & (g1032) & (g1219) & (g1220) & (g1226)) + ((g914) & (!g1032) & (!g1219) & (g1220) & (g1226)) + ((g914) & (!g1032) & (g1219) & (!g1220) & (!g1226)) + ((g914) & (!g1032) & (g1219) & (!g1220) & (g1226)) + ((g914) & (!g1032) & (g1219) & (g1220) & (!g1226)) + ((g914) & (!g1032) & (g1219) & (g1220) & (g1226)) + ((g914) & (g1032) & (!g1219) & (!g1220) & (g1226)) + ((g914) & (g1032) & (!g1219) & (g1220) & (!g1226)) + ((g914) & (g1032) & (!g1219) & (g1220) & (g1226)) + ((g914) & (g1032) & (g1219) & (!g1220) & (!g1226)) + ((g914) & (g1032) & (g1219) & (!g1220) & (g1226)) + ((g914) & (g1032) & (g1219) & (g1220) & (!g1226)) + ((g914) & (g1032) & (g1219) & (g1220) & (g1226)));
	assign g1228 = (((!g803) & (!g851) & (g1216) & (g1217) & (g1227)) + ((!g803) & (g851) & (g1216) & (!g1217) & (g1227)) + ((!g803) & (g851) & (g1216) & (g1217) & (!g1227)) + ((!g803) & (g851) & (g1216) & (g1217) & (g1227)) + ((g803) & (!g851) & (!g1216) & (g1217) & (g1227)) + ((g803) & (!g851) & (g1216) & (!g1217) & (!g1227)) + ((g803) & (!g851) & (g1216) & (!g1217) & (g1227)) + ((g803) & (!g851) & (g1216) & (g1217) & (!g1227)) + ((g803) & (!g851) & (g1216) & (g1217) & (g1227)) + ((g803) & (g851) & (!g1216) & (!g1217) & (g1227)) + ((g803) & (g851) & (!g1216) & (g1217) & (!g1227)) + ((g803) & (g851) & (!g1216) & (g1217) & (g1227)) + ((g803) & (g851) & (g1216) & (!g1217) & (!g1227)) + ((g803) & (g851) & (g1216) & (!g1217) & (g1227)) + ((g803) & (g851) & (g1216) & (g1217) & (!g1227)) + ((g803) & (g851) & (g1216) & (g1217) & (g1227)));
	assign g1229 = (((!g700) & (!g744) & (g1213) & (g1214) & (g1228)) + ((!g700) & (g744) & (g1213) & (!g1214) & (g1228)) + ((!g700) & (g744) & (g1213) & (g1214) & (!g1228)) + ((!g700) & (g744) & (g1213) & (g1214) & (g1228)) + ((g700) & (!g744) & (!g1213) & (g1214) & (g1228)) + ((g700) & (!g744) & (g1213) & (!g1214) & (!g1228)) + ((g700) & (!g744) & (g1213) & (!g1214) & (g1228)) + ((g700) & (!g744) & (g1213) & (g1214) & (!g1228)) + ((g700) & (!g744) & (g1213) & (g1214) & (g1228)) + ((g700) & (g744) & (!g1213) & (!g1214) & (g1228)) + ((g700) & (g744) & (!g1213) & (g1214) & (!g1228)) + ((g700) & (g744) & (!g1213) & (g1214) & (g1228)) + ((g700) & (g744) & (g1213) & (!g1214) & (!g1228)) + ((g700) & (g744) & (g1213) & (!g1214) & (g1228)) + ((g700) & (g744) & (g1213) & (g1214) & (!g1228)) + ((g700) & (g744) & (g1213) & (g1214) & (g1228)));
	assign g1230 = (((!g4) & (!g1207) & (!g1208) & (!g1168) & (!g1210)) + ((!g4) & (!g1207) & (!g1208) & (g1168) & (!g1210)) + ((!g4) & (!g1207) & (!g1208) & (g1168) & (g1210)) + ((!g4) & (!g1207) & (g1208) & (!g1168) & (g1210)) + ((!g4) & (g1207) & (g1208) & (!g1168) & (!g1210)) + ((!g4) & (g1207) & (g1208) & (!g1168) & (g1210)) + ((!g4) & (g1207) & (g1208) & (g1168) & (!g1210)) + ((!g4) & (g1207) & (g1208) & (g1168) & (g1210)) + ((g4) & (!g1207) & (g1208) & (!g1168) & (!g1210)) + ((g4) & (!g1207) & (g1208) & (!g1168) & (g1210)) + ((g4) & (!g1207) & (g1208) & (g1168) & (!g1210)) + ((g4) & (!g1207) & (g1208) & (g1168) & (g1210)) + ((g4) & (g1207) & (!g1208) & (!g1168) & (!g1210)) + ((g4) & (g1207) & (!g1208) & (g1168) & (!g1210)) + ((g4) & (g1207) & (!g1208) & (g1168) & (g1210)) + ((g4) & (g1207) & (g1208) & (!g1168) & (g1210)));
	assign g1231 = (((!g8) & (!g1171) & (g1206) & (!g1168) & (!g1210)) + ((!g8) & (!g1171) & (g1206) & (g1168) & (!g1210)) + ((!g8) & (!g1171) & (g1206) & (g1168) & (g1210)) + ((!g8) & (g1171) & (!g1206) & (!g1168) & (!g1210)) + ((!g8) & (g1171) & (!g1206) & (!g1168) & (g1210)) + ((!g8) & (g1171) & (!g1206) & (g1168) & (!g1210)) + ((!g8) & (g1171) & (!g1206) & (g1168) & (g1210)) + ((!g8) & (g1171) & (g1206) & (!g1168) & (g1210)) + ((g8) & (!g1171) & (!g1206) & (!g1168) & (!g1210)) + ((g8) & (!g1171) & (!g1206) & (g1168) & (!g1210)) + ((g8) & (!g1171) & (!g1206) & (g1168) & (g1210)) + ((g8) & (g1171) & (!g1206) & (!g1168) & (g1210)) + ((g8) & (g1171) & (g1206) & (!g1168) & (!g1210)) + ((g8) & (g1171) & (g1206) & (!g1168) & (g1210)) + ((g8) & (g1171) & (g1206) & (g1168) & (!g1210)) + ((g8) & (g1171) & (g1206) & (g1168) & (g1210)));
	assign g1232 = (((!g18) & (!g27) & (g1173) & (g1205)) + ((!g18) & (g27) & (!g1173) & (g1205)) + ((!g18) & (g27) & (g1173) & (!g1205)) + ((!g18) & (g27) & (g1173) & (g1205)) + ((g18) & (!g27) & (!g1173) & (!g1205)) + ((g18) & (!g27) & (!g1173) & (g1205)) + ((g18) & (!g27) & (g1173) & (!g1205)) + ((g18) & (g27) & (!g1173) & (!g1205)));
	assign g1233 = (((!g1172) & (!g1168) & (!g1210) & (g1232)) + ((!g1172) & (g1168) & (!g1210) & (g1232)) + ((!g1172) & (g1168) & (g1210) & (g1232)) + ((g1172) & (!g1168) & (!g1210) & (!g1232)) + ((g1172) & (!g1168) & (g1210) & (!g1232)) + ((g1172) & (!g1168) & (g1210) & (g1232)) + ((g1172) & (g1168) & (!g1210) & (!g1232)) + ((g1172) & (g1168) & (g1210) & (!g1232)));
	assign g1234 = (((!g27) & (!g1173) & (g1205) & (!g1168) & (!g1210)) + ((!g27) & (!g1173) & (g1205) & (g1168) & (!g1210)) + ((!g27) & (!g1173) & (g1205) & (g1168) & (g1210)) + ((!g27) & (g1173) & (!g1205) & (!g1168) & (!g1210)) + ((!g27) & (g1173) & (!g1205) & (!g1168) & (g1210)) + ((!g27) & (g1173) & (!g1205) & (g1168) & (!g1210)) + ((!g27) & (g1173) & (!g1205) & (g1168) & (g1210)) + ((!g27) & (g1173) & (g1205) & (!g1168) & (g1210)) + ((g27) & (!g1173) & (!g1205) & (!g1168) & (!g1210)) + ((g27) & (!g1173) & (!g1205) & (g1168) & (!g1210)) + ((g27) & (!g1173) & (!g1205) & (g1168) & (g1210)) + ((g27) & (g1173) & (!g1205) & (!g1168) & (g1210)) + ((g27) & (g1173) & (g1205) & (!g1168) & (!g1210)) + ((g27) & (g1173) & (g1205) & (!g1168) & (g1210)) + ((g27) & (g1173) & (g1205) & (g1168) & (!g1210)) + ((g27) & (g1173) & (g1205) & (g1168) & (g1210)));
	assign g1235 = (((!g39) & (!g54) & (g1175) & (g1204)) + ((!g39) & (g54) & (!g1175) & (g1204)) + ((!g39) & (g54) & (g1175) & (!g1204)) + ((!g39) & (g54) & (g1175) & (g1204)) + ((g39) & (!g54) & (!g1175) & (!g1204)) + ((g39) & (!g54) & (!g1175) & (g1204)) + ((g39) & (!g54) & (g1175) & (!g1204)) + ((g39) & (g54) & (!g1175) & (!g1204)));
	assign g1236 = (((!g1174) & (!g1168) & (!g1210) & (g1235)) + ((!g1174) & (g1168) & (!g1210) & (g1235)) + ((!g1174) & (g1168) & (g1210) & (g1235)) + ((g1174) & (!g1168) & (!g1210) & (!g1235)) + ((g1174) & (!g1168) & (g1210) & (!g1235)) + ((g1174) & (!g1168) & (g1210) & (g1235)) + ((g1174) & (g1168) & (!g1210) & (!g1235)) + ((g1174) & (g1168) & (g1210) & (!g1235)));
	assign g1237 = (((!g54) & (!g1175) & (g1204) & (!g1168) & (!g1210)) + ((!g54) & (!g1175) & (g1204) & (g1168) & (!g1210)) + ((!g54) & (!g1175) & (g1204) & (g1168) & (g1210)) + ((!g54) & (g1175) & (!g1204) & (!g1168) & (!g1210)) + ((!g54) & (g1175) & (!g1204) & (!g1168) & (g1210)) + ((!g54) & (g1175) & (!g1204) & (g1168) & (!g1210)) + ((!g54) & (g1175) & (!g1204) & (g1168) & (g1210)) + ((!g54) & (g1175) & (g1204) & (!g1168) & (g1210)) + ((g54) & (!g1175) & (!g1204) & (!g1168) & (!g1210)) + ((g54) & (!g1175) & (!g1204) & (g1168) & (!g1210)) + ((g54) & (!g1175) & (!g1204) & (g1168) & (g1210)) + ((g54) & (g1175) & (!g1204) & (!g1168) & (g1210)) + ((g54) & (g1175) & (g1204) & (!g1168) & (!g1210)) + ((g54) & (g1175) & (g1204) & (!g1168) & (g1210)) + ((g54) & (g1175) & (g1204) & (g1168) & (!g1210)) + ((g54) & (g1175) & (g1204) & (g1168) & (g1210)));
	assign g1238 = (((!g68) & (!g87) & (g1177) & (g1203)) + ((!g68) & (g87) & (!g1177) & (g1203)) + ((!g68) & (g87) & (g1177) & (!g1203)) + ((!g68) & (g87) & (g1177) & (g1203)) + ((g68) & (!g87) & (!g1177) & (!g1203)) + ((g68) & (!g87) & (!g1177) & (g1203)) + ((g68) & (!g87) & (g1177) & (!g1203)) + ((g68) & (g87) & (!g1177) & (!g1203)));
	assign g1239 = (((!g1176) & (!g1168) & (!g1210) & (g1238)) + ((!g1176) & (g1168) & (!g1210) & (g1238)) + ((!g1176) & (g1168) & (g1210) & (g1238)) + ((g1176) & (!g1168) & (!g1210) & (!g1238)) + ((g1176) & (!g1168) & (g1210) & (!g1238)) + ((g1176) & (!g1168) & (g1210) & (g1238)) + ((g1176) & (g1168) & (!g1210) & (!g1238)) + ((g1176) & (g1168) & (g1210) & (!g1238)));
	assign g1240 = (((!g87) & (!g1177) & (g1203) & (!g1168) & (!g1210)) + ((!g87) & (!g1177) & (g1203) & (g1168) & (!g1210)) + ((!g87) & (!g1177) & (g1203) & (g1168) & (g1210)) + ((!g87) & (g1177) & (!g1203) & (!g1168) & (!g1210)) + ((!g87) & (g1177) & (!g1203) & (!g1168) & (g1210)) + ((!g87) & (g1177) & (!g1203) & (g1168) & (!g1210)) + ((!g87) & (g1177) & (!g1203) & (g1168) & (g1210)) + ((!g87) & (g1177) & (g1203) & (!g1168) & (g1210)) + ((g87) & (!g1177) & (!g1203) & (!g1168) & (!g1210)) + ((g87) & (!g1177) & (!g1203) & (g1168) & (!g1210)) + ((g87) & (!g1177) & (!g1203) & (g1168) & (g1210)) + ((g87) & (g1177) & (!g1203) & (!g1168) & (g1210)) + ((g87) & (g1177) & (g1203) & (!g1168) & (!g1210)) + ((g87) & (g1177) & (g1203) & (!g1168) & (g1210)) + ((g87) & (g1177) & (g1203) & (g1168) & (!g1210)) + ((g87) & (g1177) & (g1203) & (g1168) & (g1210)));
	assign g1241 = (((!g104) & (!g127) & (g1179) & (g1202)) + ((!g104) & (g127) & (!g1179) & (g1202)) + ((!g104) & (g127) & (g1179) & (!g1202)) + ((!g104) & (g127) & (g1179) & (g1202)) + ((g104) & (!g127) & (!g1179) & (!g1202)) + ((g104) & (!g127) & (!g1179) & (g1202)) + ((g104) & (!g127) & (g1179) & (!g1202)) + ((g104) & (g127) & (!g1179) & (!g1202)));
	assign g1242 = (((!g1178) & (!g1168) & (!g1210) & (g1241)) + ((!g1178) & (g1168) & (!g1210) & (g1241)) + ((!g1178) & (g1168) & (g1210) & (g1241)) + ((g1178) & (!g1168) & (!g1210) & (!g1241)) + ((g1178) & (!g1168) & (g1210) & (!g1241)) + ((g1178) & (!g1168) & (g1210) & (g1241)) + ((g1178) & (g1168) & (!g1210) & (!g1241)) + ((g1178) & (g1168) & (g1210) & (!g1241)));
	assign g1243 = (((!g127) & (!g1179) & (g1202) & (!g1168) & (!g1210)) + ((!g127) & (!g1179) & (g1202) & (g1168) & (!g1210)) + ((!g127) & (!g1179) & (g1202) & (g1168) & (g1210)) + ((!g127) & (g1179) & (!g1202) & (!g1168) & (!g1210)) + ((!g127) & (g1179) & (!g1202) & (!g1168) & (g1210)) + ((!g127) & (g1179) & (!g1202) & (g1168) & (!g1210)) + ((!g127) & (g1179) & (!g1202) & (g1168) & (g1210)) + ((!g127) & (g1179) & (g1202) & (!g1168) & (g1210)) + ((g127) & (!g1179) & (!g1202) & (!g1168) & (!g1210)) + ((g127) & (!g1179) & (!g1202) & (g1168) & (!g1210)) + ((g127) & (!g1179) & (!g1202) & (g1168) & (g1210)) + ((g127) & (g1179) & (!g1202) & (!g1168) & (g1210)) + ((g127) & (g1179) & (g1202) & (!g1168) & (!g1210)) + ((g127) & (g1179) & (g1202) & (!g1168) & (g1210)) + ((g127) & (g1179) & (g1202) & (g1168) & (!g1210)) + ((g127) & (g1179) & (g1202) & (g1168) & (g1210)));
	assign g1244 = (((!g147) & (!g174) & (g1181) & (g1201)) + ((!g147) & (g174) & (!g1181) & (g1201)) + ((!g147) & (g174) & (g1181) & (!g1201)) + ((!g147) & (g174) & (g1181) & (g1201)) + ((g147) & (!g174) & (!g1181) & (!g1201)) + ((g147) & (!g174) & (!g1181) & (g1201)) + ((g147) & (!g174) & (g1181) & (!g1201)) + ((g147) & (g174) & (!g1181) & (!g1201)));
	assign g1245 = (((!g1180) & (!g1168) & (!g1210) & (g1244)) + ((!g1180) & (g1168) & (!g1210) & (g1244)) + ((!g1180) & (g1168) & (g1210) & (g1244)) + ((g1180) & (!g1168) & (!g1210) & (!g1244)) + ((g1180) & (!g1168) & (g1210) & (!g1244)) + ((g1180) & (!g1168) & (g1210) & (g1244)) + ((g1180) & (g1168) & (!g1210) & (!g1244)) + ((g1180) & (g1168) & (g1210) & (!g1244)));
	assign g1246 = (((!g174) & (!g1181) & (g1201) & (!g1168) & (!g1210)) + ((!g174) & (!g1181) & (g1201) & (g1168) & (!g1210)) + ((!g174) & (!g1181) & (g1201) & (g1168) & (g1210)) + ((!g174) & (g1181) & (!g1201) & (!g1168) & (!g1210)) + ((!g174) & (g1181) & (!g1201) & (!g1168) & (g1210)) + ((!g174) & (g1181) & (!g1201) & (g1168) & (!g1210)) + ((!g174) & (g1181) & (!g1201) & (g1168) & (g1210)) + ((!g174) & (g1181) & (g1201) & (!g1168) & (g1210)) + ((g174) & (!g1181) & (!g1201) & (!g1168) & (!g1210)) + ((g174) & (!g1181) & (!g1201) & (g1168) & (!g1210)) + ((g174) & (!g1181) & (!g1201) & (g1168) & (g1210)) + ((g174) & (g1181) & (!g1201) & (!g1168) & (g1210)) + ((g174) & (g1181) & (g1201) & (!g1168) & (!g1210)) + ((g174) & (g1181) & (g1201) & (!g1168) & (g1210)) + ((g174) & (g1181) & (g1201) & (g1168) & (!g1210)) + ((g174) & (g1181) & (g1201) & (g1168) & (g1210)));
	assign g1247 = (((!g198) & (!g229) & (g1183) & (g1200)) + ((!g198) & (g229) & (!g1183) & (g1200)) + ((!g198) & (g229) & (g1183) & (!g1200)) + ((!g198) & (g229) & (g1183) & (g1200)) + ((g198) & (!g229) & (!g1183) & (!g1200)) + ((g198) & (!g229) & (!g1183) & (g1200)) + ((g198) & (!g229) & (g1183) & (!g1200)) + ((g198) & (g229) & (!g1183) & (!g1200)));
	assign g1248 = (((!g1182) & (!g1168) & (!g1210) & (g1247)) + ((!g1182) & (g1168) & (!g1210) & (g1247)) + ((!g1182) & (g1168) & (g1210) & (g1247)) + ((g1182) & (!g1168) & (!g1210) & (!g1247)) + ((g1182) & (!g1168) & (g1210) & (!g1247)) + ((g1182) & (!g1168) & (g1210) & (g1247)) + ((g1182) & (g1168) & (!g1210) & (!g1247)) + ((g1182) & (g1168) & (g1210) & (!g1247)));
	assign g1249 = (((!g229) & (!g1183) & (g1200) & (!g1168) & (!g1210)) + ((!g229) & (!g1183) & (g1200) & (g1168) & (!g1210)) + ((!g229) & (!g1183) & (g1200) & (g1168) & (g1210)) + ((!g229) & (g1183) & (!g1200) & (!g1168) & (!g1210)) + ((!g229) & (g1183) & (!g1200) & (!g1168) & (g1210)) + ((!g229) & (g1183) & (!g1200) & (g1168) & (!g1210)) + ((!g229) & (g1183) & (!g1200) & (g1168) & (g1210)) + ((!g229) & (g1183) & (g1200) & (!g1168) & (g1210)) + ((g229) & (!g1183) & (!g1200) & (!g1168) & (!g1210)) + ((g229) & (!g1183) & (!g1200) & (g1168) & (!g1210)) + ((g229) & (!g1183) & (!g1200) & (g1168) & (g1210)) + ((g229) & (g1183) & (!g1200) & (!g1168) & (g1210)) + ((g229) & (g1183) & (g1200) & (!g1168) & (!g1210)) + ((g229) & (g1183) & (g1200) & (!g1168) & (g1210)) + ((g229) & (g1183) & (g1200) & (g1168) & (!g1210)) + ((g229) & (g1183) & (g1200) & (g1168) & (g1210)));
	assign g1250 = (((!g255) & (!g290) & (g1185) & (g1199)) + ((!g255) & (g290) & (!g1185) & (g1199)) + ((!g255) & (g290) & (g1185) & (!g1199)) + ((!g255) & (g290) & (g1185) & (g1199)) + ((g255) & (!g290) & (!g1185) & (!g1199)) + ((g255) & (!g290) & (!g1185) & (g1199)) + ((g255) & (!g290) & (g1185) & (!g1199)) + ((g255) & (g290) & (!g1185) & (!g1199)));
	assign g1251 = (((!g1184) & (!g1168) & (!g1210) & (g1250)) + ((!g1184) & (g1168) & (!g1210) & (g1250)) + ((!g1184) & (g1168) & (g1210) & (g1250)) + ((g1184) & (!g1168) & (!g1210) & (!g1250)) + ((g1184) & (!g1168) & (g1210) & (!g1250)) + ((g1184) & (!g1168) & (g1210) & (g1250)) + ((g1184) & (g1168) & (!g1210) & (!g1250)) + ((g1184) & (g1168) & (g1210) & (!g1250)));
	assign g1252 = (((!g290) & (!g1185) & (g1199) & (!g1168) & (!g1210)) + ((!g290) & (!g1185) & (g1199) & (g1168) & (!g1210)) + ((!g290) & (!g1185) & (g1199) & (g1168) & (g1210)) + ((!g290) & (g1185) & (!g1199) & (!g1168) & (!g1210)) + ((!g290) & (g1185) & (!g1199) & (!g1168) & (g1210)) + ((!g290) & (g1185) & (!g1199) & (g1168) & (!g1210)) + ((!g290) & (g1185) & (!g1199) & (g1168) & (g1210)) + ((!g290) & (g1185) & (g1199) & (!g1168) & (g1210)) + ((g290) & (!g1185) & (!g1199) & (!g1168) & (!g1210)) + ((g290) & (!g1185) & (!g1199) & (g1168) & (!g1210)) + ((g290) & (!g1185) & (!g1199) & (g1168) & (g1210)) + ((g290) & (g1185) & (!g1199) & (!g1168) & (g1210)) + ((g290) & (g1185) & (g1199) & (!g1168) & (!g1210)) + ((g290) & (g1185) & (g1199) & (!g1168) & (g1210)) + ((g290) & (g1185) & (g1199) & (g1168) & (!g1210)) + ((g290) & (g1185) & (g1199) & (g1168) & (g1210)));
	assign g1253 = (((!g319) & (!g358) & (g1187) & (g1198)) + ((!g319) & (g358) & (!g1187) & (g1198)) + ((!g319) & (g358) & (g1187) & (!g1198)) + ((!g319) & (g358) & (g1187) & (g1198)) + ((g319) & (!g358) & (!g1187) & (!g1198)) + ((g319) & (!g358) & (!g1187) & (g1198)) + ((g319) & (!g358) & (g1187) & (!g1198)) + ((g319) & (g358) & (!g1187) & (!g1198)));
	assign g1254 = (((!g1186) & (!g1168) & (!g1210) & (g1253)) + ((!g1186) & (g1168) & (!g1210) & (g1253)) + ((!g1186) & (g1168) & (g1210) & (g1253)) + ((g1186) & (!g1168) & (!g1210) & (!g1253)) + ((g1186) & (!g1168) & (g1210) & (!g1253)) + ((g1186) & (!g1168) & (g1210) & (g1253)) + ((g1186) & (g1168) & (!g1210) & (!g1253)) + ((g1186) & (g1168) & (g1210) & (!g1253)));
	assign g1255 = (((!g358) & (!g1187) & (g1198) & (!g1168) & (!g1210)) + ((!g358) & (!g1187) & (g1198) & (g1168) & (!g1210)) + ((!g358) & (!g1187) & (g1198) & (g1168) & (g1210)) + ((!g358) & (g1187) & (!g1198) & (!g1168) & (!g1210)) + ((!g358) & (g1187) & (!g1198) & (!g1168) & (g1210)) + ((!g358) & (g1187) & (!g1198) & (g1168) & (!g1210)) + ((!g358) & (g1187) & (!g1198) & (g1168) & (g1210)) + ((!g358) & (g1187) & (g1198) & (!g1168) & (g1210)) + ((g358) & (!g1187) & (!g1198) & (!g1168) & (!g1210)) + ((g358) & (!g1187) & (!g1198) & (g1168) & (!g1210)) + ((g358) & (!g1187) & (!g1198) & (g1168) & (g1210)) + ((g358) & (g1187) & (!g1198) & (!g1168) & (g1210)) + ((g358) & (g1187) & (g1198) & (!g1168) & (!g1210)) + ((g358) & (g1187) & (g1198) & (!g1168) & (g1210)) + ((g358) & (g1187) & (g1198) & (g1168) & (!g1210)) + ((g358) & (g1187) & (g1198) & (g1168) & (g1210)));
	assign g1256 = (((!g390) & (!g433) & (g1189) & (g1197)) + ((!g390) & (g433) & (!g1189) & (g1197)) + ((!g390) & (g433) & (g1189) & (!g1197)) + ((!g390) & (g433) & (g1189) & (g1197)) + ((g390) & (!g433) & (!g1189) & (!g1197)) + ((g390) & (!g433) & (!g1189) & (g1197)) + ((g390) & (!g433) & (g1189) & (!g1197)) + ((g390) & (g433) & (!g1189) & (!g1197)));
	assign g1257 = (((!g1188) & (!g1168) & (!g1210) & (g1256)) + ((!g1188) & (g1168) & (!g1210) & (g1256)) + ((!g1188) & (g1168) & (g1210) & (g1256)) + ((g1188) & (!g1168) & (!g1210) & (!g1256)) + ((g1188) & (!g1168) & (g1210) & (!g1256)) + ((g1188) & (!g1168) & (g1210) & (g1256)) + ((g1188) & (g1168) & (!g1210) & (!g1256)) + ((g1188) & (g1168) & (g1210) & (!g1256)));
	assign g1258 = (((!g433) & (!g1189) & (g1197) & (!g1168) & (!g1210)) + ((!g433) & (!g1189) & (g1197) & (g1168) & (!g1210)) + ((!g433) & (!g1189) & (g1197) & (g1168) & (g1210)) + ((!g433) & (g1189) & (!g1197) & (!g1168) & (!g1210)) + ((!g433) & (g1189) & (!g1197) & (!g1168) & (g1210)) + ((!g433) & (g1189) & (!g1197) & (g1168) & (!g1210)) + ((!g433) & (g1189) & (!g1197) & (g1168) & (g1210)) + ((!g433) & (g1189) & (g1197) & (!g1168) & (g1210)) + ((g433) & (!g1189) & (!g1197) & (!g1168) & (!g1210)) + ((g433) & (!g1189) & (!g1197) & (g1168) & (!g1210)) + ((g433) & (!g1189) & (!g1197) & (g1168) & (g1210)) + ((g433) & (g1189) & (!g1197) & (!g1168) & (g1210)) + ((g433) & (g1189) & (g1197) & (!g1168) & (!g1210)) + ((g433) & (g1189) & (g1197) & (!g1168) & (g1210)) + ((g433) & (g1189) & (g1197) & (g1168) & (!g1210)) + ((g433) & (g1189) & (g1197) & (g1168) & (g1210)));
	assign g1259 = (((!g468) & (!g515) & (g1191) & (g1196)) + ((!g468) & (g515) & (!g1191) & (g1196)) + ((!g468) & (g515) & (g1191) & (!g1196)) + ((!g468) & (g515) & (g1191) & (g1196)) + ((g468) & (!g515) & (!g1191) & (!g1196)) + ((g468) & (!g515) & (!g1191) & (g1196)) + ((g468) & (!g515) & (g1191) & (!g1196)) + ((g468) & (g515) & (!g1191) & (!g1196)));
	assign g1260 = (((!g1190) & (!g1168) & (!g1210) & (g1259)) + ((!g1190) & (g1168) & (!g1210) & (g1259)) + ((!g1190) & (g1168) & (g1210) & (g1259)) + ((g1190) & (!g1168) & (!g1210) & (!g1259)) + ((g1190) & (!g1168) & (g1210) & (!g1259)) + ((g1190) & (!g1168) & (g1210) & (g1259)) + ((g1190) & (g1168) & (!g1210) & (!g1259)) + ((g1190) & (g1168) & (g1210) & (!g1259)));
	assign g1261 = (((!g515) & (!g1191) & (g1196) & (!g1168) & (!g1210)) + ((!g515) & (!g1191) & (g1196) & (g1168) & (!g1210)) + ((!g515) & (!g1191) & (g1196) & (g1168) & (g1210)) + ((!g515) & (g1191) & (!g1196) & (!g1168) & (!g1210)) + ((!g515) & (g1191) & (!g1196) & (!g1168) & (g1210)) + ((!g515) & (g1191) & (!g1196) & (g1168) & (!g1210)) + ((!g515) & (g1191) & (!g1196) & (g1168) & (g1210)) + ((!g515) & (g1191) & (g1196) & (!g1168) & (g1210)) + ((g515) & (!g1191) & (!g1196) & (!g1168) & (!g1210)) + ((g515) & (!g1191) & (!g1196) & (g1168) & (!g1210)) + ((g515) & (!g1191) & (!g1196) & (g1168) & (g1210)) + ((g515) & (g1191) & (!g1196) & (!g1168) & (g1210)) + ((g515) & (g1191) & (g1196) & (!g1168) & (!g1210)) + ((g515) & (g1191) & (g1196) & (!g1168) & (g1210)) + ((g515) & (g1191) & (g1196) & (g1168) & (!g1210)) + ((g515) & (g1191) & (g1196) & (g1168) & (g1210)));
	assign g1262 = (((!g553) & (!g604) & (g1193) & (g1195)) + ((!g553) & (g604) & (!g1193) & (g1195)) + ((!g553) & (g604) & (g1193) & (!g1195)) + ((!g553) & (g604) & (g1193) & (g1195)) + ((g553) & (!g604) & (!g1193) & (!g1195)) + ((g553) & (!g604) & (!g1193) & (g1195)) + ((g553) & (!g604) & (g1193) & (!g1195)) + ((g553) & (g604) & (!g1193) & (!g1195)));
	assign g1263 = (((!g1192) & (!g1168) & (!g1210) & (g1262)) + ((!g1192) & (g1168) & (!g1210) & (g1262)) + ((!g1192) & (g1168) & (g1210) & (g1262)) + ((g1192) & (!g1168) & (!g1210) & (!g1262)) + ((g1192) & (!g1168) & (g1210) & (!g1262)) + ((g1192) & (!g1168) & (g1210) & (g1262)) + ((g1192) & (g1168) & (!g1210) & (!g1262)) + ((g1192) & (g1168) & (g1210) & (!g1262)));
	assign g1264 = (((!g604) & (!g1193) & (g1195) & (!g1168) & (!g1210)) + ((!g604) & (!g1193) & (g1195) & (g1168) & (!g1210)) + ((!g604) & (!g1193) & (g1195) & (g1168) & (g1210)) + ((!g604) & (g1193) & (!g1195) & (!g1168) & (!g1210)) + ((!g604) & (g1193) & (!g1195) & (!g1168) & (g1210)) + ((!g604) & (g1193) & (!g1195) & (g1168) & (!g1210)) + ((!g604) & (g1193) & (!g1195) & (g1168) & (g1210)) + ((!g604) & (g1193) & (g1195) & (!g1168) & (g1210)) + ((g604) & (!g1193) & (!g1195) & (!g1168) & (!g1210)) + ((g604) & (!g1193) & (!g1195) & (g1168) & (!g1210)) + ((g604) & (!g1193) & (!g1195) & (g1168) & (g1210)) + ((g604) & (g1193) & (!g1195) & (!g1168) & (g1210)) + ((g604) & (g1193) & (g1195) & (!g1168) & (!g1210)) + ((g604) & (g1193) & (g1195) & (!g1168) & (g1210)) + ((g604) & (g1193) & (g1195) & (g1168) & (!g1210)) + ((g604) & (g1193) & (g1195) & (g1168) & (g1210)));
	assign g1265 = (((!g645) & (!g700) & (g1155) & (g1167)) + ((!g645) & (g700) & (!g1155) & (g1167)) + ((!g645) & (g700) & (g1155) & (!g1167)) + ((!g645) & (g700) & (g1155) & (g1167)) + ((g645) & (!g700) & (!g1155) & (!g1167)) + ((g645) & (!g700) & (!g1155) & (g1167)) + ((g645) & (!g700) & (g1155) & (!g1167)) + ((g645) & (g700) & (!g1155) & (!g1167)));
	assign g1266 = (((!g1194) & (!g1168) & (!g1210) & (g1265)) + ((!g1194) & (g1168) & (!g1210) & (g1265)) + ((!g1194) & (g1168) & (g1210) & (g1265)) + ((g1194) & (!g1168) & (!g1210) & (!g1265)) + ((g1194) & (!g1168) & (g1210) & (!g1265)) + ((g1194) & (!g1168) & (g1210) & (g1265)) + ((g1194) & (g1168) & (!g1210) & (!g1265)) + ((g1194) & (g1168) & (g1210) & (!g1265)));
	assign g1267 = (((!g604) & (!g645) & (g1266) & (g1211) & (g1229)) + ((!g604) & (g645) & (g1266) & (!g1211) & (g1229)) + ((!g604) & (g645) & (g1266) & (g1211) & (!g1229)) + ((!g604) & (g645) & (g1266) & (g1211) & (g1229)) + ((g604) & (!g645) & (!g1266) & (g1211) & (g1229)) + ((g604) & (!g645) & (g1266) & (!g1211) & (!g1229)) + ((g604) & (!g645) & (g1266) & (!g1211) & (g1229)) + ((g604) & (!g645) & (g1266) & (g1211) & (!g1229)) + ((g604) & (!g645) & (g1266) & (g1211) & (g1229)) + ((g604) & (g645) & (!g1266) & (!g1211) & (g1229)) + ((g604) & (g645) & (!g1266) & (g1211) & (!g1229)) + ((g604) & (g645) & (!g1266) & (g1211) & (g1229)) + ((g604) & (g645) & (g1266) & (!g1211) & (!g1229)) + ((g604) & (g645) & (g1266) & (!g1211) & (g1229)) + ((g604) & (g645) & (g1266) & (g1211) & (!g1229)) + ((g604) & (g645) & (g1266) & (g1211) & (g1229)));
	assign g1268 = (((!g515) & (!g553) & (g1263) & (g1264) & (g1267)) + ((!g515) & (g553) & (g1263) & (!g1264) & (g1267)) + ((!g515) & (g553) & (g1263) & (g1264) & (!g1267)) + ((!g515) & (g553) & (g1263) & (g1264) & (g1267)) + ((g515) & (!g553) & (!g1263) & (g1264) & (g1267)) + ((g515) & (!g553) & (g1263) & (!g1264) & (!g1267)) + ((g515) & (!g553) & (g1263) & (!g1264) & (g1267)) + ((g515) & (!g553) & (g1263) & (g1264) & (!g1267)) + ((g515) & (!g553) & (g1263) & (g1264) & (g1267)) + ((g515) & (g553) & (!g1263) & (!g1264) & (g1267)) + ((g515) & (g553) & (!g1263) & (g1264) & (!g1267)) + ((g515) & (g553) & (!g1263) & (g1264) & (g1267)) + ((g515) & (g553) & (g1263) & (!g1264) & (!g1267)) + ((g515) & (g553) & (g1263) & (!g1264) & (g1267)) + ((g515) & (g553) & (g1263) & (g1264) & (!g1267)) + ((g515) & (g553) & (g1263) & (g1264) & (g1267)));
	assign g1269 = (((!g433) & (!g468) & (g1260) & (g1261) & (g1268)) + ((!g433) & (g468) & (g1260) & (!g1261) & (g1268)) + ((!g433) & (g468) & (g1260) & (g1261) & (!g1268)) + ((!g433) & (g468) & (g1260) & (g1261) & (g1268)) + ((g433) & (!g468) & (!g1260) & (g1261) & (g1268)) + ((g433) & (!g468) & (g1260) & (!g1261) & (!g1268)) + ((g433) & (!g468) & (g1260) & (!g1261) & (g1268)) + ((g433) & (!g468) & (g1260) & (g1261) & (!g1268)) + ((g433) & (!g468) & (g1260) & (g1261) & (g1268)) + ((g433) & (g468) & (!g1260) & (!g1261) & (g1268)) + ((g433) & (g468) & (!g1260) & (g1261) & (!g1268)) + ((g433) & (g468) & (!g1260) & (g1261) & (g1268)) + ((g433) & (g468) & (g1260) & (!g1261) & (!g1268)) + ((g433) & (g468) & (g1260) & (!g1261) & (g1268)) + ((g433) & (g468) & (g1260) & (g1261) & (!g1268)) + ((g433) & (g468) & (g1260) & (g1261) & (g1268)));
	assign g1270 = (((!g358) & (!g390) & (g1257) & (g1258) & (g1269)) + ((!g358) & (g390) & (g1257) & (!g1258) & (g1269)) + ((!g358) & (g390) & (g1257) & (g1258) & (!g1269)) + ((!g358) & (g390) & (g1257) & (g1258) & (g1269)) + ((g358) & (!g390) & (!g1257) & (g1258) & (g1269)) + ((g358) & (!g390) & (g1257) & (!g1258) & (!g1269)) + ((g358) & (!g390) & (g1257) & (!g1258) & (g1269)) + ((g358) & (!g390) & (g1257) & (g1258) & (!g1269)) + ((g358) & (!g390) & (g1257) & (g1258) & (g1269)) + ((g358) & (g390) & (!g1257) & (!g1258) & (g1269)) + ((g358) & (g390) & (!g1257) & (g1258) & (!g1269)) + ((g358) & (g390) & (!g1257) & (g1258) & (g1269)) + ((g358) & (g390) & (g1257) & (!g1258) & (!g1269)) + ((g358) & (g390) & (g1257) & (!g1258) & (g1269)) + ((g358) & (g390) & (g1257) & (g1258) & (!g1269)) + ((g358) & (g390) & (g1257) & (g1258) & (g1269)));
	assign g1271 = (((!g290) & (!g319) & (g1254) & (g1255) & (g1270)) + ((!g290) & (g319) & (g1254) & (!g1255) & (g1270)) + ((!g290) & (g319) & (g1254) & (g1255) & (!g1270)) + ((!g290) & (g319) & (g1254) & (g1255) & (g1270)) + ((g290) & (!g319) & (!g1254) & (g1255) & (g1270)) + ((g290) & (!g319) & (g1254) & (!g1255) & (!g1270)) + ((g290) & (!g319) & (g1254) & (!g1255) & (g1270)) + ((g290) & (!g319) & (g1254) & (g1255) & (!g1270)) + ((g290) & (!g319) & (g1254) & (g1255) & (g1270)) + ((g290) & (g319) & (!g1254) & (!g1255) & (g1270)) + ((g290) & (g319) & (!g1254) & (g1255) & (!g1270)) + ((g290) & (g319) & (!g1254) & (g1255) & (g1270)) + ((g290) & (g319) & (g1254) & (!g1255) & (!g1270)) + ((g290) & (g319) & (g1254) & (!g1255) & (g1270)) + ((g290) & (g319) & (g1254) & (g1255) & (!g1270)) + ((g290) & (g319) & (g1254) & (g1255) & (g1270)));
	assign g1272 = (((!g229) & (!g255) & (g1251) & (g1252) & (g1271)) + ((!g229) & (g255) & (g1251) & (!g1252) & (g1271)) + ((!g229) & (g255) & (g1251) & (g1252) & (!g1271)) + ((!g229) & (g255) & (g1251) & (g1252) & (g1271)) + ((g229) & (!g255) & (!g1251) & (g1252) & (g1271)) + ((g229) & (!g255) & (g1251) & (!g1252) & (!g1271)) + ((g229) & (!g255) & (g1251) & (!g1252) & (g1271)) + ((g229) & (!g255) & (g1251) & (g1252) & (!g1271)) + ((g229) & (!g255) & (g1251) & (g1252) & (g1271)) + ((g229) & (g255) & (!g1251) & (!g1252) & (g1271)) + ((g229) & (g255) & (!g1251) & (g1252) & (!g1271)) + ((g229) & (g255) & (!g1251) & (g1252) & (g1271)) + ((g229) & (g255) & (g1251) & (!g1252) & (!g1271)) + ((g229) & (g255) & (g1251) & (!g1252) & (g1271)) + ((g229) & (g255) & (g1251) & (g1252) & (!g1271)) + ((g229) & (g255) & (g1251) & (g1252) & (g1271)));
	assign g1273 = (((!g174) & (!g198) & (g1248) & (g1249) & (g1272)) + ((!g174) & (g198) & (g1248) & (!g1249) & (g1272)) + ((!g174) & (g198) & (g1248) & (g1249) & (!g1272)) + ((!g174) & (g198) & (g1248) & (g1249) & (g1272)) + ((g174) & (!g198) & (!g1248) & (g1249) & (g1272)) + ((g174) & (!g198) & (g1248) & (!g1249) & (!g1272)) + ((g174) & (!g198) & (g1248) & (!g1249) & (g1272)) + ((g174) & (!g198) & (g1248) & (g1249) & (!g1272)) + ((g174) & (!g198) & (g1248) & (g1249) & (g1272)) + ((g174) & (g198) & (!g1248) & (!g1249) & (g1272)) + ((g174) & (g198) & (!g1248) & (g1249) & (!g1272)) + ((g174) & (g198) & (!g1248) & (g1249) & (g1272)) + ((g174) & (g198) & (g1248) & (!g1249) & (!g1272)) + ((g174) & (g198) & (g1248) & (!g1249) & (g1272)) + ((g174) & (g198) & (g1248) & (g1249) & (!g1272)) + ((g174) & (g198) & (g1248) & (g1249) & (g1272)));
	assign g1274 = (((!g127) & (!g147) & (g1245) & (g1246) & (g1273)) + ((!g127) & (g147) & (g1245) & (!g1246) & (g1273)) + ((!g127) & (g147) & (g1245) & (g1246) & (!g1273)) + ((!g127) & (g147) & (g1245) & (g1246) & (g1273)) + ((g127) & (!g147) & (!g1245) & (g1246) & (g1273)) + ((g127) & (!g147) & (g1245) & (!g1246) & (!g1273)) + ((g127) & (!g147) & (g1245) & (!g1246) & (g1273)) + ((g127) & (!g147) & (g1245) & (g1246) & (!g1273)) + ((g127) & (!g147) & (g1245) & (g1246) & (g1273)) + ((g127) & (g147) & (!g1245) & (!g1246) & (g1273)) + ((g127) & (g147) & (!g1245) & (g1246) & (!g1273)) + ((g127) & (g147) & (!g1245) & (g1246) & (g1273)) + ((g127) & (g147) & (g1245) & (!g1246) & (!g1273)) + ((g127) & (g147) & (g1245) & (!g1246) & (g1273)) + ((g127) & (g147) & (g1245) & (g1246) & (!g1273)) + ((g127) & (g147) & (g1245) & (g1246) & (g1273)));
	assign g1275 = (((!g87) & (!g104) & (g1242) & (g1243) & (g1274)) + ((!g87) & (g104) & (g1242) & (!g1243) & (g1274)) + ((!g87) & (g104) & (g1242) & (g1243) & (!g1274)) + ((!g87) & (g104) & (g1242) & (g1243) & (g1274)) + ((g87) & (!g104) & (!g1242) & (g1243) & (g1274)) + ((g87) & (!g104) & (g1242) & (!g1243) & (!g1274)) + ((g87) & (!g104) & (g1242) & (!g1243) & (g1274)) + ((g87) & (!g104) & (g1242) & (g1243) & (!g1274)) + ((g87) & (!g104) & (g1242) & (g1243) & (g1274)) + ((g87) & (g104) & (!g1242) & (!g1243) & (g1274)) + ((g87) & (g104) & (!g1242) & (g1243) & (!g1274)) + ((g87) & (g104) & (!g1242) & (g1243) & (g1274)) + ((g87) & (g104) & (g1242) & (!g1243) & (!g1274)) + ((g87) & (g104) & (g1242) & (!g1243) & (g1274)) + ((g87) & (g104) & (g1242) & (g1243) & (!g1274)) + ((g87) & (g104) & (g1242) & (g1243) & (g1274)));
	assign g1276 = (((!g54) & (!g68) & (g1239) & (g1240) & (g1275)) + ((!g54) & (g68) & (g1239) & (!g1240) & (g1275)) + ((!g54) & (g68) & (g1239) & (g1240) & (!g1275)) + ((!g54) & (g68) & (g1239) & (g1240) & (g1275)) + ((g54) & (!g68) & (!g1239) & (g1240) & (g1275)) + ((g54) & (!g68) & (g1239) & (!g1240) & (!g1275)) + ((g54) & (!g68) & (g1239) & (!g1240) & (g1275)) + ((g54) & (!g68) & (g1239) & (g1240) & (!g1275)) + ((g54) & (!g68) & (g1239) & (g1240) & (g1275)) + ((g54) & (g68) & (!g1239) & (!g1240) & (g1275)) + ((g54) & (g68) & (!g1239) & (g1240) & (!g1275)) + ((g54) & (g68) & (!g1239) & (g1240) & (g1275)) + ((g54) & (g68) & (g1239) & (!g1240) & (!g1275)) + ((g54) & (g68) & (g1239) & (!g1240) & (g1275)) + ((g54) & (g68) & (g1239) & (g1240) & (!g1275)) + ((g54) & (g68) & (g1239) & (g1240) & (g1275)));
	assign g1277 = (((!g27) & (!g39) & (g1236) & (g1237) & (g1276)) + ((!g27) & (g39) & (g1236) & (!g1237) & (g1276)) + ((!g27) & (g39) & (g1236) & (g1237) & (!g1276)) + ((!g27) & (g39) & (g1236) & (g1237) & (g1276)) + ((g27) & (!g39) & (!g1236) & (g1237) & (g1276)) + ((g27) & (!g39) & (g1236) & (!g1237) & (!g1276)) + ((g27) & (!g39) & (g1236) & (!g1237) & (g1276)) + ((g27) & (!g39) & (g1236) & (g1237) & (!g1276)) + ((g27) & (!g39) & (g1236) & (g1237) & (g1276)) + ((g27) & (g39) & (!g1236) & (!g1237) & (g1276)) + ((g27) & (g39) & (!g1236) & (g1237) & (!g1276)) + ((g27) & (g39) & (!g1236) & (g1237) & (g1276)) + ((g27) & (g39) & (g1236) & (!g1237) & (!g1276)) + ((g27) & (g39) & (g1236) & (!g1237) & (g1276)) + ((g27) & (g39) & (g1236) & (g1237) & (!g1276)) + ((g27) & (g39) & (g1236) & (g1237) & (g1276)));
	assign g1278 = (((!g8) & (!g18) & (g1233) & (g1234) & (g1277)) + ((!g8) & (g18) & (g1233) & (!g1234) & (g1277)) + ((!g8) & (g18) & (g1233) & (g1234) & (!g1277)) + ((!g8) & (g18) & (g1233) & (g1234) & (g1277)) + ((g8) & (!g18) & (!g1233) & (g1234) & (g1277)) + ((g8) & (!g18) & (g1233) & (!g1234) & (!g1277)) + ((g8) & (!g18) & (g1233) & (!g1234) & (g1277)) + ((g8) & (!g18) & (g1233) & (g1234) & (!g1277)) + ((g8) & (!g18) & (g1233) & (g1234) & (g1277)) + ((g8) & (g18) & (!g1233) & (!g1234) & (g1277)) + ((g8) & (g18) & (!g1233) & (g1234) & (!g1277)) + ((g8) & (g18) & (!g1233) & (g1234) & (g1277)) + ((g8) & (g18) & (g1233) & (!g1234) & (!g1277)) + ((g8) & (g18) & (g1233) & (!g1234) & (g1277)) + ((g8) & (g18) & (g1233) & (g1234) & (!g1277)) + ((g8) & (g18) & (g1233) & (g1234) & (g1277)));
	assign g1279 = (((!g2) & (!g8) & (g1171) & (g1206)) + ((!g2) & (g8) & (!g1171) & (g1206)) + ((!g2) & (g8) & (g1171) & (!g1206)) + ((!g2) & (g8) & (g1171) & (g1206)) + ((g2) & (!g8) & (!g1171) & (!g1206)) + ((g2) & (!g8) & (!g1171) & (g1206)) + ((g2) & (!g8) & (g1171) & (!g1206)) + ((g2) & (g8) & (!g1171) & (!g1206)));
	assign g1280 = (((!g1170) & (!g1168) & (!g1210) & (g1279)) + ((!g1170) & (g1168) & (!g1210) & (g1279)) + ((!g1170) & (g1168) & (g1210) & (g1279)) + ((g1170) & (!g1168) & (!g1210) & (!g1279)) + ((g1170) & (!g1168) & (g1210) & (!g1279)) + ((g1170) & (!g1168) & (g1210) & (g1279)) + ((g1170) & (g1168) & (!g1210) & (!g1279)) + ((g1170) & (g1168) & (g1210) & (!g1279)));
	assign g1281 = (((!g4) & (!g2) & (!g1231) & (!g1278) & (g1280)) + ((!g4) & (!g2) & (!g1231) & (g1278) & (g1280)) + ((!g4) & (!g2) & (g1231) & (!g1278) & (g1280)) + ((!g4) & (!g2) & (g1231) & (g1278) & (!g1280)) + ((!g4) & (!g2) & (g1231) & (g1278) & (g1280)) + ((!g4) & (g2) & (!g1231) & (!g1278) & (g1280)) + ((!g4) & (g2) & (!g1231) & (g1278) & (!g1280)) + ((!g4) & (g2) & (!g1231) & (g1278) & (g1280)) + ((!g4) & (g2) & (g1231) & (!g1278) & (!g1280)) + ((!g4) & (g2) & (g1231) & (!g1278) & (g1280)) + ((!g4) & (g2) & (g1231) & (g1278) & (!g1280)) + ((!g4) & (g2) & (g1231) & (g1278) & (g1280)) + ((g4) & (!g2) & (g1231) & (g1278) & (g1280)) + ((g4) & (g2) & (!g1231) & (g1278) & (g1280)) + ((g4) & (g2) & (g1231) & (!g1278) & (g1280)) + ((g4) & (g2) & (g1231) & (g1278) & (g1280)));
	assign g1282 = (((!g4) & (!g1207) & (g1208)) + ((!g4) & (g1207) & (!g1208)) + ((!g4) & (g1207) & (g1208)) + ((g4) & (g1207) & (g1208)));
	assign g1283 = (((!g1169) & (!g1282) & (!g1168) & (!g1210)) + ((!g1169) & (!g1282) & (g1168) & (!g1210)) + ((!g1169) & (!g1282) & (g1168) & (g1210)) + ((g1169) & (g1282) & (!g1168) & (!g1210)) + ((g1169) & (g1282) & (!g1168) & (g1210)) + ((g1169) & (g1282) & (g1168) & (!g1210)) + ((g1169) & (g1282) & (g1168) & (g1210)));
	assign g1284 = (((!g1) & (g1169) & (!g1282) & (!g1168) & (g1210)) + ((!g1) & (g1169) & (g1282) & (!g1168) & (g1210)) + ((g1) & (!g1169) & (g1282) & (g1168) & (!g1210)) + ((g1) & (!g1169) & (g1282) & (g1168) & (g1210)) + ((g1) & (g1169) & (!g1282) & (!g1168) & (!g1210)) + ((g1) & (g1169) & (!g1282) & (!g1168) & (g1210)) + ((g1) & (g1169) & (!g1282) & (g1168) & (!g1210)) + ((g1) & (g1169) & (!g1282) & (g1168) & (g1210)) + ((g1) & (g1169) & (g1282) & (!g1168) & (g1210)));
	assign g1285 = (((!g1) & (!g1230) & (!g1281) & (!g1283) & (!g1284)) + ((g1) & (!g1230) & (!g1281) & (!g1283) & (!g1284)) + ((g1) & (!g1230) & (!g1281) & (g1283) & (!g1284)) + ((g1) & (!g1230) & (g1281) & (!g1283) & (!g1284)) + ((g1) & (!g1230) & (g1281) & (g1283) & (!g1284)) + ((g1) & (g1230) & (!g1281) & (!g1283) & (!g1284)) + ((g1) & (g1230) & (!g1281) & (g1283) & (!g1284)));
	assign g1286 = (((!g645) & (!g1211) & (g1229) & (!g1285)) + ((!g645) & (g1211) & (!g1229) & (!g1285)) + ((!g645) & (g1211) & (!g1229) & (g1285)) + ((!g645) & (g1211) & (g1229) & (g1285)) + ((g645) & (!g1211) & (!g1229) & (!g1285)) + ((g645) & (g1211) & (!g1229) & (g1285)) + ((g645) & (g1211) & (g1229) & (!g1285)) + ((g645) & (g1211) & (g1229) & (g1285)));
	assign g1287 = (((!g700) & (!g744) & (!g1213) & (g1214) & (g1228) & (!g1285)) + ((!g700) & (!g744) & (g1213) & (!g1214) & (!g1228) & (!g1285)) + ((!g700) & (!g744) & (g1213) & (!g1214) & (!g1228) & (g1285)) + ((!g700) & (!g744) & (g1213) & (!g1214) & (g1228) & (!g1285)) + ((!g700) & (!g744) & (g1213) & (!g1214) & (g1228) & (g1285)) + ((!g700) & (!g744) & (g1213) & (g1214) & (!g1228) & (!g1285)) + ((!g700) & (!g744) & (g1213) & (g1214) & (!g1228) & (g1285)) + ((!g700) & (!g744) & (g1213) & (g1214) & (g1228) & (g1285)) + ((!g700) & (g744) & (!g1213) & (!g1214) & (g1228) & (!g1285)) + ((!g700) & (g744) & (!g1213) & (g1214) & (!g1228) & (!g1285)) + ((!g700) & (g744) & (!g1213) & (g1214) & (g1228) & (!g1285)) + ((!g700) & (g744) & (g1213) & (!g1214) & (!g1228) & (!g1285)) + ((!g700) & (g744) & (g1213) & (!g1214) & (!g1228) & (g1285)) + ((!g700) & (g744) & (g1213) & (!g1214) & (g1228) & (g1285)) + ((!g700) & (g744) & (g1213) & (g1214) & (!g1228) & (g1285)) + ((!g700) & (g744) & (g1213) & (g1214) & (g1228) & (g1285)) + ((g700) & (!g744) & (!g1213) & (!g1214) & (!g1228) & (!g1285)) + ((g700) & (!g744) & (!g1213) & (!g1214) & (g1228) & (!g1285)) + ((g700) & (!g744) & (!g1213) & (g1214) & (!g1228) & (!g1285)) + ((g700) & (!g744) & (g1213) & (!g1214) & (!g1228) & (g1285)) + ((g700) & (!g744) & (g1213) & (!g1214) & (g1228) & (g1285)) + ((g700) & (!g744) & (g1213) & (g1214) & (!g1228) & (g1285)) + ((g700) & (!g744) & (g1213) & (g1214) & (g1228) & (!g1285)) + ((g700) & (!g744) & (g1213) & (g1214) & (g1228) & (g1285)) + ((g700) & (g744) & (!g1213) & (!g1214) & (!g1228) & (!g1285)) + ((g700) & (g744) & (g1213) & (!g1214) & (!g1228) & (g1285)) + ((g700) & (g744) & (g1213) & (!g1214) & (g1228) & (!g1285)) + ((g700) & (g744) & (g1213) & (!g1214) & (g1228) & (g1285)) + ((g700) & (g744) & (g1213) & (g1214) & (!g1228) & (!g1285)) + ((g700) & (g744) & (g1213) & (g1214) & (!g1228) & (g1285)) + ((g700) & (g744) & (g1213) & (g1214) & (g1228) & (!g1285)) + ((g700) & (g744) & (g1213) & (g1214) & (g1228) & (g1285)));
	assign g1288 = (((!g744) & (!g1214) & (g1228) & (!g1285)) + ((!g744) & (g1214) & (!g1228) & (!g1285)) + ((!g744) & (g1214) & (!g1228) & (g1285)) + ((!g744) & (g1214) & (g1228) & (g1285)) + ((g744) & (!g1214) & (!g1228) & (!g1285)) + ((g744) & (g1214) & (!g1228) & (g1285)) + ((g744) & (g1214) & (g1228) & (!g1285)) + ((g744) & (g1214) & (g1228) & (g1285)));
	assign g1289 = (((!g803) & (!g851) & (!g1216) & (g1217) & (g1227) & (!g1285)) + ((!g803) & (!g851) & (g1216) & (!g1217) & (!g1227) & (!g1285)) + ((!g803) & (!g851) & (g1216) & (!g1217) & (!g1227) & (g1285)) + ((!g803) & (!g851) & (g1216) & (!g1217) & (g1227) & (!g1285)) + ((!g803) & (!g851) & (g1216) & (!g1217) & (g1227) & (g1285)) + ((!g803) & (!g851) & (g1216) & (g1217) & (!g1227) & (!g1285)) + ((!g803) & (!g851) & (g1216) & (g1217) & (!g1227) & (g1285)) + ((!g803) & (!g851) & (g1216) & (g1217) & (g1227) & (g1285)) + ((!g803) & (g851) & (!g1216) & (!g1217) & (g1227) & (!g1285)) + ((!g803) & (g851) & (!g1216) & (g1217) & (!g1227) & (!g1285)) + ((!g803) & (g851) & (!g1216) & (g1217) & (g1227) & (!g1285)) + ((!g803) & (g851) & (g1216) & (!g1217) & (!g1227) & (!g1285)) + ((!g803) & (g851) & (g1216) & (!g1217) & (!g1227) & (g1285)) + ((!g803) & (g851) & (g1216) & (!g1217) & (g1227) & (g1285)) + ((!g803) & (g851) & (g1216) & (g1217) & (!g1227) & (g1285)) + ((!g803) & (g851) & (g1216) & (g1217) & (g1227) & (g1285)) + ((g803) & (!g851) & (!g1216) & (!g1217) & (!g1227) & (!g1285)) + ((g803) & (!g851) & (!g1216) & (!g1217) & (g1227) & (!g1285)) + ((g803) & (!g851) & (!g1216) & (g1217) & (!g1227) & (!g1285)) + ((g803) & (!g851) & (g1216) & (!g1217) & (!g1227) & (g1285)) + ((g803) & (!g851) & (g1216) & (!g1217) & (g1227) & (g1285)) + ((g803) & (!g851) & (g1216) & (g1217) & (!g1227) & (g1285)) + ((g803) & (!g851) & (g1216) & (g1217) & (g1227) & (!g1285)) + ((g803) & (!g851) & (g1216) & (g1217) & (g1227) & (g1285)) + ((g803) & (g851) & (!g1216) & (!g1217) & (!g1227) & (!g1285)) + ((g803) & (g851) & (g1216) & (!g1217) & (!g1227) & (g1285)) + ((g803) & (g851) & (g1216) & (!g1217) & (g1227) & (!g1285)) + ((g803) & (g851) & (g1216) & (!g1217) & (g1227) & (g1285)) + ((g803) & (g851) & (g1216) & (g1217) & (!g1227) & (!g1285)) + ((g803) & (g851) & (g1216) & (g1217) & (!g1227) & (g1285)) + ((g803) & (g851) & (g1216) & (g1217) & (g1227) & (!g1285)) + ((g803) & (g851) & (g1216) & (g1217) & (g1227) & (g1285)));
	assign g1290 = (((!g851) & (!g1217) & (g1227) & (!g1285)) + ((!g851) & (g1217) & (!g1227) & (!g1285)) + ((!g851) & (g1217) & (!g1227) & (g1285)) + ((!g851) & (g1217) & (g1227) & (g1285)) + ((g851) & (!g1217) & (!g1227) & (!g1285)) + ((g851) & (g1217) & (!g1227) & (g1285)) + ((g851) & (g1217) & (g1227) & (!g1285)) + ((g851) & (g1217) & (g1227) & (g1285)));
	assign g1291 = (((!g914) & (!g1032) & (!g1219) & (g1220) & (g1226) & (!g1285)) + ((!g914) & (!g1032) & (g1219) & (!g1220) & (!g1226) & (!g1285)) + ((!g914) & (!g1032) & (g1219) & (!g1220) & (!g1226) & (g1285)) + ((!g914) & (!g1032) & (g1219) & (!g1220) & (g1226) & (!g1285)) + ((!g914) & (!g1032) & (g1219) & (!g1220) & (g1226) & (g1285)) + ((!g914) & (!g1032) & (g1219) & (g1220) & (!g1226) & (!g1285)) + ((!g914) & (!g1032) & (g1219) & (g1220) & (!g1226) & (g1285)) + ((!g914) & (!g1032) & (g1219) & (g1220) & (g1226) & (g1285)) + ((!g914) & (g1032) & (!g1219) & (!g1220) & (g1226) & (!g1285)) + ((!g914) & (g1032) & (!g1219) & (g1220) & (!g1226) & (!g1285)) + ((!g914) & (g1032) & (!g1219) & (g1220) & (g1226) & (!g1285)) + ((!g914) & (g1032) & (g1219) & (!g1220) & (!g1226) & (!g1285)) + ((!g914) & (g1032) & (g1219) & (!g1220) & (!g1226) & (g1285)) + ((!g914) & (g1032) & (g1219) & (!g1220) & (g1226) & (g1285)) + ((!g914) & (g1032) & (g1219) & (g1220) & (!g1226) & (g1285)) + ((!g914) & (g1032) & (g1219) & (g1220) & (g1226) & (g1285)) + ((g914) & (!g1032) & (!g1219) & (!g1220) & (!g1226) & (!g1285)) + ((g914) & (!g1032) & (!g1219) & (!g1220) & (g1226) & (!g1285)) + ((g914) & (!g1032) & (!g1219) & (g1220) & (!g1226) & (!g1285)) + ((g914) & (!g1032) & (g1219) & (!g1220) & (!g1226) & (g1285)) + ((g914) & (!g1032) & (g1219) & (!g1220) & (g1226) & (g1285)) + ((g914) & (!g1032) & (g1219) & (g1220) & (!g1226) & (g1285)) + ((g914) & (!g1032) & (g1219) & (g1220) & (g1226) & (!g1285)) + ((g914) & (!g1032) & (g1219) & (g1220) & (g1226) & (g1285)) + ((g914) & (g1032) & (!g1219) & (!g1220) & (!g1226) & (!g1285)) + ((g914) & (g1032) & (g1219) & (!g1220) & (!g1226) & (g1285)) + ((g914) & (g1032) & (g1219) & (!g1220) & (g1226) & (!g1285)) + ((g914) & (g1032) & (g1219) & (!g1220) & (g1226) & (g1285)) + ((g914) & (g1032) & (g1219) & (g1220) & (!g1226) & (!g1285)) + ((g914) & (g1032) & (g1219) & (g1220) & (!g1226) & (g1285)) + ((g914) & (g1032) & (g1219) & (g1220) & (g1226) & (!g1285)) + ((g914) & (g1032) & (g1219) & (g1220) & (g1226) & (g1285)));
	assign g1292 = (((!g1032) & (!g1220) & (g1226) & (!g1285)) + ((!g1032) & (g1220) & (!g1226) & (!g1285)) + ((!g1032) & (g1220) & (!g1226) & (g1285)) + ((!g1032) & (g1220) & (g1226) & (g1285)) + ((g1032) & (!g1220) & (!g1226) & (!g1285)) + ((g1032) & (g1220) & (!g1226) & (g1285)) + ((g1032) & (g1220) & (g1226) & (!g1285)) + ((g1032) & (g1220) & (g1226) & (g1285)));
	assign g1293 = (((!g1030) & (!g1160) & (!g1222) & (g1223) & (g1225) & (!g1285)) + ((!g1030) & (!g1160) & (g1222) & (!g1223) & (!g1225) & (!g1285)) + ((!g1030) & (!g1160) & (g1222) & (!g1223) & (!g1225) & (g1285)) + ((!g1030) & (!g1160) & (g1222) & (!g1223) & (g1225) & (!g1285)) + ((!g1030) & (!g1160) & (g1222) & (!g1223) & (g1225) & (g1285)) + ((!g1030) & (!g1160) & (g1222) & (g1223) & (!g1225) & (!g1285)) + ((!g1030) & (!g1160) & (g1222) & (g1223) & (!g1225) & (g1285)) + ((!g1030) & (!g1160) & (g1222) & (g1223) & (g1225) & (g1285)) + ((!g1030) & (g1160) & (!g1222) & (!g1223) & (g1225) & (!g1285)) + ((!g1030) & (g1160) & (!g1222) & (g1223) & (!g1225) & (!g1285)) + ((!g1030) & (g1160) & (!g1222) & (g1223) & (g1225) & (!g1285)) + ((!g1030) & (g1160) & (g1222) & (!g1223) & (!g1225) & (!g1285)) + ((!g1030) & (g1160) & (g1222) & (!g1223) & (!g1225) & (g1285)) + ((!g1030) & (g1160) & (g1222) & (!g1223) & (g1225) & (g1285)) + ((!g1030) & (g1160) & (g1222) & (g1223) & (!g1225) & (g1285)) + ((!g1030) & (g1160) & (g1222) & (g1223) & (g1225) & (g1285)) + ((g1030) & (!g1160) & (!g1222) & (!g1223) & (!g1225) & (!g1285)) + ((g1030) & (!g1160) & (!g1222) & (!g1223) & (g1225) & (!g1285)) + ((g1030) & (!g1160) & (!g1222) & (g1223) & (!g1225) & (!g1285)) + ((g1030) & (!g1160) & (g1222) & (!g1223) & (!g1225) & (g1285)) + ((g1030) & (!g1160) & (g1222) & (!g1223) & (g1225) & (g1285)) + ((g1030) & (!g1160) & (g1222) & (g1223) & (!g1225) & (g1285)) + ((g1030) & (!g1160) & (g1222) & (g1223) & (g1225) & (!g1285)) + ((g1030) & (!g1160) & (g1222) & (g1223) & (g1225) & (g1285)) + ((g1030) & (g1160) & (!g1222) & (!g1223) & (!g1225) & (!g1285)) + ((g1030) & (g1160) & (g1222) & (!g1223) & (!g1225) & (g1285)) + ((g1030) & (g1160) & (g1222) & (!g1223) & (g1225) & (!g1285)) + ((g1030) & (g1160) & (g1222) & (!g1223) & (g1225) & (g1285)) + ((g1030) & (g1160) & (g1222) & (g1223) & (!g1225) & (!g1285)) + ((g1030) & (g1160) & (g1222) & (g1223) & (!g1225) & (g1285)) + ((g1030) & (g1160) & (g1222) & (g1223) & (g1225) & (!g1285)) + ((g1030) & (g1160) & (g1222) & (g1223) & (g1225) & (g1285)));
	assign g1294 = (((!g1160) & (!g1223) & (g1225) & (!g1285)) + ((!g1160) & (g1223) & (!g1225) & (!g1285)) + ((!g1160) & (g1223) & (!g1225) & (g1285)) + ((!g1160) & (g1223) & (g1225) & (g1285)) + ((g1160) & (!g1223) & (!g1225) & (!g1285)) + ((g1160) & (g1223) & (!g1225) & (g1285)) + ((g1160) & (g1223) & (g1225) & (!g1285)) + ((g1160) & (g1223) & (g1225) & (g1285)));
	assign g1295 = (((!g1168) & (g1210)));
	assign g1296 = (((!g1154) & (!ax54x) & (!ax55x) & (!g1295) & (!g1224) & (g1285)) + ((!g1154) & (!ax54x) & (!ax55x) & (!g1295) & (g1224) & (!g1285)) + ((!g1154) & (!ax54x) & (!ax55x) & (!g1295) & (g1224) & (g1285)) + ((!g1154) & (!ax54x) & (!ax55x) & (g1295) & (!g1224) & (!g1285)) + ((!g1154) & (!ax54x) & (ax55x) & (!g1295) & (!g1224) & (!g1285)) + ((!g1154) & (!ax54x) & (ax55x) & (g1295) & (!g1224) & (g1285)) + ((!g1154) & (!ax54x) & (ax55x) & (g1295) & (g1224) & (!g1285)) + ((!g1154) & (!ax54x) & (ax55x) & (g1295) & (g1224) & (g1285)) + ((!g1154) & (ax54x) & (!ax55x) & (g1295) & (!g1224) & (!g1285)) + ((!g1154) & (ax54x) & (!ax55x) & (g1295) & (g1224) & (!g1285)) + ((!g1154) & (ax54x) & (ax55x) & (!g1295) & (!g1224) & (!g1285)) + ((!g1154) & (ax54x) & (ax55x) & (!g1295) & (!g1224) & (g1285)) + ((!g1154) & (ax54x) & (ax55x) & (!g1295) & (g1224) & (!g1285)) + ((!g1154) & (ax54x) & (ax55x) & (!g1295) & (g1224) & (g1285)) + ((!g1154) & (ax54x) & (ax55x) & (g1295) & (!g1224) & (g1285)) + ((!g1154) & (ax54x) & (ax55x) & (g1295) & (g1224) & (g1285)) + ((g1154) & (!ax54x) & (!ax55x) & (!g1295) & (!g1224) & (!g1285)) + ((g1154) & (!ax54x) & (!ax55x) & (!g1295) & (!g1224) & (g1285)) + ((g1154) & (!ax54x) & (!ax55x) & (!g1295) & (g1224) & (g1285)) + ((g1154) & (!ax54x) & (!ax55x) & (g1295) & (g1224) & (!g1285)) + ((g1154) & (!ax54x) & (ax55x) & (!g1295) & (g1224) & (!g1285)) + ((g1154) & (!ax54x) & (ax55x) & (g1295) & (!g1224) & (!g1285)) + ((g1154) & (!ax54x) & (ax55x) & (g1295) & (!g1224) & (g1285)) + ((g1154) & (!ax54x) & (ax55x) & (g1295) & (g1224) & (g1285)) + ((g1154) & (ax54x) & (!ax55x) & (!g1295) & (!g1224) & (!g1285)) + ((g1154) & (ax54x) & (!ax55x) & (!g1295) & (g1224) & (!g1285)) + ((g1154) & (ax54x) & (ax55x) & (!g1295) & (!g1224) & (g1285)) + ((g1154) & (ax54x) & (ax55x) & (!g1295) & (g1224) & (g1285)) + ((g1154) & (ax54x) & (ax55x) & (g1295) & (!g1224) & (!g1285)) + ((g1154) & (ax54x) & (ax55x) & (g1295) & (!g1224) & (g1285)) + ((g1154) & (ax54x) & (ax55x) & (g1295) & (g1224) & (!g1285)) + ((g1154) & (ax54x) & (ax55x) & (g1295) & (g1224) & (g1285)));
	assign g1297 = (((!ax54x) & (!g1295) & (!g1224) & (g1285)) + ((!ax54x) & (!g1295) & (g1224) & (!g1285)) + ((!ax54x) & (!g1295) & (g1224) & (g1285)) + ((!ax54x) & (g1295) & (g1224) & (!g1285)) + ((ax54x) & (!g1295) & (!g1224) & (!g1285)) + ((ax54x) & (g1295) & (!g1224) & (!g1285)) + ((ax54x) & (g1295) & (!g1224) & (g1285)) + ((ax54x) & (g1295) & (g1224) & (g1285)));
	assign g1298 = (((!ax50x) & (!ax51x)));
	assign g1299 = (((!g1295) & (!ax52x) & (!ax53x) & (!g1285) & (!g1298)) + ((!g1295) & (!ax52x) & (ax53x) & (g1285) & (!g1298)) + ((!g1295) & (ax52x) & (ax53x) & (g1285) & (!g1298)) + ((!g1295) & (ax52x) & (ax53x) & (g1285) & (g1298)) + ((g1295) & (!ax52x) & (!ax53x) & (!g1285) & (!g1298)) + ((g1295) & (!ax52x) & (!ax53x) & (!g1285) & (g1298)) + ((g1295) & (!ax52x) & (!ax53x) & (g1285) & (!g1298)) + ((g1295) & (!ax52x) & (ax53x) & (!g1285) & (!g1298)) + ((g1295) & (!ax52x) & (ax53x) & (g1285) & (!g1298)) + ((g1295) & (!ax52x) & (ax53x) & (g1285) & (g1298)) + ((g1295) & (ax52x) & (!ax53x) & (g1285) & (!g1298)) + ((g1295) & (ax52x) & (!ax53x) & (g1285) & (g1298)) + ((g1295) & (ax52x) & (ax53x) & (!g1285) & (!g1298)) + ((g1295) & (ax52x) & (ax53x) & (!g1285) & (g1298)) + ((g1295) & (ax52x) & (ax53x) & (g1285) & (!g1298)) + ((g1295) & (ax52x) & (ax53x) & (g1285) & (g1298)));
	assign g1300 = (((!g1160) & (!g1154) & (g1296) & (g1297) & (g1299)) + ((!g1160) & (g1154) & (g1296) & (!g1297) & (g1299)) + ((!g1160) & (g1154) & (g1296) & (g1297) & (!g1299)) + ((!g1160) & (g1154) & (g1296) & (g1297) & (g1299)) + ((g1160) & (!g1154) & (!g1296) & (g1297) & (g1299)) + ((g1160) & (!g1154) & (g1296) & (!g1297) & (!g1299)) + ((g1160) & (!g1154) & (g1296) & (!g1297) & (g1299)) + ((g1160) & (!g1154) & (g1296) & (g1297) & (!g1299)) + ((g1160) & (!g1154) & (g1296) & (g1297) & (g1299)) + ((g1160) & (g1154) & (!g1296) & (!g1297) & (g1299)) + ((g1160) & (g1154) & (!g1296) & (g1297) & (!g1299)) + ((g1160) & (g1154) & (!g1296) & (g1297) & (g1299)) + ((g1160) & (g1154) & (g1296) & (!g1297) & (!g1299)) + ((g1160) & (g1154) & (g1296) & (!g1297) & (g1299)) + ((g1160) & (g1154) & (g1296) & (g1297) & (!g1299)) + ((g1160) & (g1154) & (g1296) & (g1297) & (g1299)));
	assign g1301 = (((!g1032) & (!g1030) & (g1293) & (g1294) & (g1300)) + ((!g1032) & (g1030) & (g1293) & (!g1294) & (g1300)) + ((!g1032) & (g1030) & (g1293) & (g1294) & (!g1300)) + ((!g1032) & (g1030) & (g1293) & (g1294) & (g1300)) + ((g1032) & (!g1030) & (!g1293) & (g1294) & (g1300)) + ((g1032) & (!g1030) & (g1293) & (!g1294) & (!g1300)) + ((g1032) & (!g1030) & (g1293) & (!g1294) & (g1300)) + ((g1032) & (!g1030) & (g1293) & (g1294) & (!g1300)) + ((g1032) & (!g1030) & (g1293) & (g1294) & (g1300)) + ((g1032) & (g1030) & (!g1293) & (!g1294) & (g1300)) + ((g1032) & (g1030) & (!g1293) & (g1294) & (!g1300)) + ((g1032) & (g1030) & (!g1293) & (g1294) & (g1300)) + ((g1032) & (g1030) & (g1293) & (!g1294) & (!g1300)) + ((g1032) & (g1030) & (g1293) & (!g1294) & (g1300)) + ((g1032) & (g1030) & (g1293) & (g1294) & (!g1300)) + ((g1032) & (g1030) & (g1293) & (g1294) & (g1300)));
	assign g1302 = (((!g851) & (!g914) & (g1291) & (g1292) & (g1301)) + ((!g851) & (g914) & (g1291) & (!g1292) & (g1301)) + ((!g851) & (g914) & (g1291) & (g1292) & (!g1301)) + ((!g851) & (g914) & (g1291) & (g1292) & (g1301)) + ((g851) & (!g914) & (!g1291) & (g1292) & (g1301)) + ((g851) & (!g914) & (g1291) & (!g1292) & (!g1301)) + ((g851) & (!g914) & (g1291) & (!g1292) & (g1301)) + ((g851) & (!g914) & (g1291) & (g1292) & (!g1301)) + ((g851) & (!g914) & (g1291) & (g1292) & (g1301)) + ((g851) & (g914) & (!g1291) & (!g1292) & (g1301)) + ((g851) & (g914) & (!g1291) & (g1292) & (!g1301)) + ((g851) & (g914) & (!g1291) & (g1292) & (g1301)) + ((g851) & (g914) & (g1291) & (!g1292) & (!g1301)) + ((g851) & (g914) & (g1291) & (!g1292) & (g1301)) + ((g851) & (g914) & (g1291) & (g1292) & (!g1301)) + ((g851) & (g914) & (g1291) & (g1292) & (g1301)));
	assign g1303 = (((!g744) & (!g803) & (g1289) & (g1290) & (g1302)) + ((!g744) & (g803) & (g1289) & (!g1290) & (g1302)) + ((!g744) & (g803) & (g1289) & (g1290) & (!g1302)) + ((!g744) & (g803) & (g1289) & (g1290) & (g1302)) + ((g744) & (!g803) & (!g1289) & (g1290) & (g1302)) + ((g744) & (!g803) & (g1289) & (!g1290) & (!g1302)) + ((g744) & (!g803) & (g1289) & (!g1290) & (g1302)) + ((g744) & (!g803) & (g1289) & (g1290) & (!g1302)) + ((g744) & (!g803) & (g1289) & (g1290) & (g1302)) + ((g744) & (g803) & (!g1289) & (!g1290) & (g1302)) + ((g744) & (g803) & (!g1289) & (g1290) & (!g1302)) + ((g744) & (g803) & (!g1289) & (g1290) & (g1302)) + ((g744) & (g803) & (g1289) & (!g1290) & (!g1302)) + ((g744) & (g803) & (g1289) & (!g1290) & (g1302)) + ((g744) & (g803) & (g1289) & (g1290) & (!g1302)) + ((g744) & (g803) & (g1289) & (g1290) & (g1302)));
	assign g1304 = (((!g645) & (!g700) & (g1287) & (g1288) & (g1303)) + ((!g645) & (g700) & (g1287) & (!g1288) & (g1303)) + ((!g645) & (g700) & (g1287) & (g1288) & (!g1303)) + ((!g645) & (g700) & (g1287) & (g1288) & (g1303)) + ((g645) & (!g700) & (!g1287) & (g1288) & (g1303)) + ((g645) & (!g700) & (g1287) & (!g1288) & (!g1303)) + ((g645) & (!g700) & (g1287) & (!g1288) & (g1303)) + ((g645) & (!g700) & (g1287) & (g1288) & (!g1303)) + ((g645) & (!g700) & (g1287) & (g1288) & (g1303)) + ((g645) & (g700) & (!g1287) & (!g1288) & (g1303)) + ((g645) & (g700) & (!g1287) & (g1288) & (!g1303)) + ((g645) & (g700) & (!g1287) & (g1288) & (g1303)) + ((g645) & (g700) & (g1287) & (!g1288) & (!g1303)) + ((g645) & (g700) & (g1287) & (!g1288) & (g1303)) + ((g645) & (g700) & (g1287) & (g1288) & (!g1303)) + ((g645) & (g700) & (g1287) & (g1288) & (g1303)));
	assign g1305 = (((g1) & (!g1230) & (g1281) & (g1284)) + ((g1) & (g1230) & (!g1281) & (!g1284)) + ((g1) & (g1230) & (!g1281) & (g1284)));
	assign g1306 = (((!g4) & (!g2) & (!g1231) & (!g1278) & (!g1280) & (!g1285)) + ((!g4) & (!g2) & (!g1231) & (!g1278) & (g1280) & (g1285)) + ((!g4) & (!g2) & (!g1231) & (g1278) & (!g1280) & (!g1285)) + ((!g4) & (!g2) & (!g1231) & (g1278) & (g1280) & (g1285)) + ((!g4) & (!g2) & (g1231) & (!g1278) & (!g1280) & (!g1285)) + ((!g4) & (!g2) & (g1231) & (!g1278) & (g1280) & (g1285)) + ((!g4) & (!g2) & (g1231) & (g1278) & (g1280) & (!g1285)) + ((!g4) & (!g2) & (g1231) & (g1278) & (g1280) & (g1285)) + ((!g4) & (g2) & (!g1231) & (!g1278) & (!g1280) & (!g1285)) + ((!g4) & (g2) & (!g1231) & (!g1278) & (g1280) & (g1285)) + ((!g4) & (g2) & (!g1231) & (g1278) & (g1280) & (!g1285)) + ((!g4) & (g2) & (!g1231) & (g1278) & (g1280) & (g1285)) + ((!g4) & (g2) & (g1231) & (!g1278) & (g1280) & (!g1285)) + ((!g4) & (g2) & (g1231) & (!g1278) & (g1280) & (g1285)) + ((!g4) & (g2) & (g1231) & (g1278) & (g1280) & (!g1285)) + ((!g4) & (g2) & (g1231) & (g1278) & (g1280) & (g1285)) + ((g4) & (!g2) & (!g1231) & (!g1278) & (g1280) & (!g1285)) + ((g4) & (!g2) & (!g1231) & (!g1278) & (g1280) & (g1285)) + ((g4) & (!g2) & (!g1231) & (g1278) & (g1280) & (!g1285)) + ((g4) & (!g2) & (!g1231) & (g1278) & (g1280) & (g1285)) + ((g4) & (!g2) & (g1231) & (!g1278) & (g1280) & (!g1285)) + ((g4) & (!g2) & (g1231) & (!g1278) & (g1280) & (g1285)) + ((g4) & (!g2) & (g1231) & (g1278) & (!g1280) & (!g1285)) + ((g4) & (!g2) & (g1231) & (g1278) & (g1280) & (g1285)) + ((g4) & (g2) & (!g1231) & (!g1278) & (g1280) & (!g1285)) + ((g4) & (g2) & (!g1231) & (!g1278) & (g1280) & (g1285)) + ((g4) & (g2) & (!g1231) & (g1278) & (!g1280) & (!g1285)) + ((g4) & (g2) & (!g1231) & (g1278) & (g1280) & (g1285)) + ((g4) & (g2) & (g1231) & (!g1278) & (!g1280) & (!g1285)) + ((g4) & (g2) & (g1231) & (!g1278) & (g1280) & (g1285)) + ((g4) & (g2) & (g1231) & (g1278) & (!g1280) & (!g1285)) + ((g4) & (g2) & (g1231) & (g1278) & (g1280) & (g1285)));
	assign g1307 = (((!g8) & (!g18) & (!g1233) & (g1234) & (g1277) & (!g1285)) + ((!g8) & (!g18) & (g1233) & (!g1234) & (!g1277) & (!g1285)) + ((!g8) & (!g18) & (g1233) & (!g1234) & (!g1277) & (g1285)) + ((!g8) & (!g18) & (g1233) & (!g1234) & (g1277) & (!g1285)) + ((!g8) & (!g18) & (g1233) & (!g1234) & (g1277) & (g1285)) + ((!g8) & (!g18) & (g1233) & (g1234) & (!g1277) & (!g1285)) + ((!g8) & (!g18) & (g1233) & (g1234) & (!g1277) & (g1285)) + ((!g8) & (!g18) & (g1233) & (g1234) & (g1277) & (g1285)) + ((!g8) & (g18) & (!g1233) & (!g1234) & (g1277) & (!g1285)) + ((!g8) & (g18) & (!g1233) & (g1234) & (!g1277) & (!g1285)) + ((!g8) & (g18) & (!g1233) & (g1234) & (g1277) & (!g1285)) + ((!g8) & (g18) & (g1233) & (!g1234) & (!g1277) & (!g1285)) + ((!g8) & (g18) & (g1233) & (!g1234) & (!g1277) & (g1285)) + ((!g8) & (g18) & (g1233) & (!g1234) & (g1277) & (g1285)) + ((!g8) & (g18) & (g1233) & (g1234) & (!g1277) & (g1285)) + ((!g8) & (g18) & (g1233) & (g1234) & (g1277) & (g1285)) + ((g8) & (!g18) & (!g1233) & (!g1234) & (!g1277) & (!g1285)) + ((g8) & (!g18) & (!g1233) & (!g1234) & (g1277) & (!g1285)) + ((g8) & (!g18) & (!g1233) & (g1234) & (!g1277) & (!g1285)) + ((g8) & (!g18) & (g1233) & (!g1234) & (!g1277) & (g1285)) + ((g8) & (!g18) & (g1233) & (!g1234) & (g1277) & (g1285)) + ((g8) & (!g18) & (g1233) & (g1234) & (!g1277) & (g1285)) + ((g8) & (!g18) & (g1233) & (g1234) & (g1277) & (!g1285)) + ((g8) & (!g18) & (g1233) & (g1234) & (g1277) & (g1285)) + ((g8) & (g18) & (!g1233) & (!g1234) & (!g1277) & (!g1285)) + ((g8) & (g18) & (g1233) & (!g1234) & (!g1277) & (g1285)) + ((g8) & (g18) & (g1233) & (!g1234) & (g1277) & (!g1285)) + ((g8) & (g18) & (g1233) & (!g1234) & (g1277) & (g1285)) + ((g8) & (g18) & (g1233) & (g1234) & (!g1277) & (!g1285)) + ((g8) & (g18) & (g1233) & (g1234) & (!g1277) & (g1285)) + ((g8) & (g18) & (g1233) & (g1234) & (g1277) & (!g1285)) + ((g8) & (g18) & (g1233) & (g1234) & (g1277) & (g1285)));
	assign g1308 = (((!g18) & (!g1234) & (g1277) & (!g1285)) + ((!g18) & (g1234) & (!g1277) & (!g1285)) + ((!g18) & (g1234) & (!g1277) & (g1285)) + ((!g18) & (g1234) & (g1277) & (g1285)) + ((g18) & (!g1234) & (!g1277) & (!g1285)) + ((g18) & (g1234) & (!g1277) & (g1285)) + ((g18) & (g1234) & (g1277) & (!g1285)) + ((g18) & (g1234) & (g1277) & (g1285)));
	assign g1309 = (((!g27) & (!g39) & (!g1236) & (g1237) & (g1276) & (!g1285)) + ((!g27) & (!g39) & (g1236) & (!g1237) & (!g1276) & (!g1285)) + ((!g27) & (!g39) & (g1236) & (!g1237) & (!g1276) & (g1285)) + ((!g27) & (!g39) & (g1236) & (!g1237) & (g1276) & (!g1285)) + ((!g27) & (!g39) & (g1236) & (!g1237) & (g1276) & (g1285)) + ((!g27) & (!g39) & (g1236) & (g1237) & (!g1276) & (!g1285)) + ((!g27) & (!g39) & (g1236) & (g1237) & (!g1276) & (g1285)) + ((!g27) & (!g39) & (g1236) & (g1237) & (g1276) & (g1285)) + ((!g27) & (g39) & (!g1236) & (!g1237) & (g1276) & (!g1285)) + ((!g27) & (g39) & (!g1236) & (g1237) & (!g1276) & (!g1285)) + ((!g27) & (g39) & (!g1236) & (g1237) & (g1276) & (!g1285)) + ((!g27) & (g39) & (g1236) & (!g1237) & (!g1276) & (!g1285)) + ((!g27) & (g39) & (g1236) & (!g1237) & (!g1276) & (g1285)) + ((!g27) & (g39) & (g1236) & (!g1237) & (g1276) & (g1285)) + ((!g27) & (g39) & (g1236) & (g1237) & (!g1276) & (g1285)) + ((!g27) & (g39) & (g1236) & (g1237) & (g1276) & (g1285)) + ((g27) & (!g39) & (!g1236) & (!g1237) & (!g1276) & (!g1285)) + ((g27) & (!g39) & (!g1236) & (!g1237) & (g1276) & (!g1285)) + ((g27) & (!g39) & (!g1236) & (g1237) & (!g1276) & (!g1285)) + ((g27) & (!g39) & (g1236) & (!g1237) & (!g1276) & (g1285)) + ((g27) & (!g39) & (g1236) & (!g1237) & (g1276) & (g1285)) + ((g27) & (!g39) & (g1236) & (g1237) & (!g1276) & (g1285)) + ((g27) & (!g39) & (g1236) & (g1237) & (g1276) & (!g1285)) + ((g27) & (!g39) & (g1236) & (g1237) & (g1276) & (g1285)) + ((g27) & (g39) & (!g1236) & (!g1237) & (!g1276) & (!g1285)) + ((g27) & (g39) & (g1236) & (!g1237) & (!g1276) & (g1285)) + ((g27) & (g39) & (g1236) & (!g1237) & (g1276) & (!g1285)) + ((g27) & (g39) & (g1236) & (!g1237) & (g1276) & (g1285)) + ((g27) & (g39) & (g1236) & (g1237) & (!g1276) & (!g1285)) + ((g27) & (g39) & (g1236) & (g1237) & (!g1276) & (g1285)) + ((g27) & (g39) & (g1236) & (g1237) & (g1276) & (!g1285)) + ((g27) & (g39) & (g1236) & (g1237) & (g1276) & (g1285)));
	assign g1310 = (((!g39) & (!g1237) & (g1276) & (!g1285)) + ((!g39) & (g1237) & (!g1276) & (!g1285)) + ((!g39) & (g1237) & (!g1276) & (g1285)) + ((!g39) & (g1237) & (g1276) & (g1285)) + ((g39) & (!g1237) & (!g1276) & (!g1285)) + ((g39) & (g1237) & (!g1276) & (g1285)) + ((g39) & (g1237) & (g1276) & (!g1285)) + ((g39) & (g1237) & (g1276) & (g1285)));
	assign g1311 = (((!g54) & (!g68) & (!g1239) & (g1240) & (g1275) & (!g1285)) + ((!g54) & (!g68) & (g1239) & (!g1240) & (!g1275) & (!g1285)) + ((!g54) & (!g68) & (g1239) & (!g1240) & (!g1275) & (g1285)) + ((!g54) & (!g68) & (g1239) & (!g1240) & (g1275) & (!g1285)) + ((!g54) & (!g68) & (g1239) & (!g1240) & (g1275) & (g1285)) + ((!g54) & (!g68) & (g1239) & (g1240) & (!g1275) & (!g1285)) + ((!g54) & (!g68) & (g1239) & (g1240) & (!g1275) & (g1285)) + ((!g54) & (!g68) & (g1239) & (g1240) & (g1275) & (g1285)) + ((!g54) & (g68) & (!g1239) & (!g1240) & (g1275) & (!g1285)) + ((!g54) & (g68) & (!g1239) & (g1240) & (!g1275) & (!g1285)) + ((!g54) & (g68) & (!g1239) & (g1240) & (g1275) & (!g1285)) + ((!g54) & (g68) & (g1239) & (!g1240) & (!g1275) & (!g1285)) + ((!g54) & (g68) & (g1239) & (!g1240) & (!g1275) & (g1285)) + ((!g54) & (g68) & (g1239) & (!g1240) & (g1275) & (g1285)) + ((!g54) & (g68) & (g1239) & (g1240) & (!g1275) & (g1285)) + ((!g54) & (g68) & (g1239) & (g1240) & (g1275) & (g1285)) + ((g54) & (!g68) & (!g1239) & (!g1240) & (!g1275) & (!g1285)) + ((g54) & (!g68) & (!g1239) & (!g1240) & (g1275) & (!g1285)) + ((g54) & (!g68) & (!g1239) & (g1240) & (!g1275) & (!g1285)) + ((g54) & (!g68) & (g1239) & (!g1240) & (!g1275) & (g1285)) + ((g54) & (!g68) & (g1239) & (!g1240) & (g1275) & (g1285)) + ((g54) & (!g68) & (g1239) & (g1240) & (!g1275) & (g1285)) + ((g54) & (!g68) & (g1239) & (g1240) & (g1275) & (!g1285)) + ((g54) & (!g68) & (g1239) & (g1240) & (g1275) & (g1285)) + ((g54) & (g68) & (!g1239) & (!g1240) & (!g1275) & (!g1285)) + ((g54) & (g68) & (g1239) & (!g1240) & (!g1275) & (g1285)) + ((g54) & (g68) & (g1239) & (!g1240) & (g1275) & (!g1285)) + ((g54) & (g68) & (g1239) & (!g1240) & (g1275) & (g1285)) + ((g54) & (g68) & (g1239) & (g1240) & (!g1275) & (!g1285)) + ((g54) & (g68) & (g1239) & (g1240) & (!g1275) & (g1285)) + ((g54) & (g68) & (g1239) & (g1240) & (g1275) & (!g1285)) + ((g54) & (g68) & (g1239) & (g1240) & (g1275) & (g1285)));
	assign g1312 = (((!g68) & (!g1240) & (g1275) & (!g1285)) + ((!g68) & (g1240) & (!g1275) & (!g1285)) + ((!g68) & (g1240) & (!g1275) & (g1285)) + ((!g68) & (g1240) & (g1275) & (g1285)) + ((g68) & (!g1240) & (!g1275) & (!g1285)) + ((g68) & (g1240) & (!g1275) & (g1285)) + ((g68) & (g1240) & (g1275) & (!g1285)) + ((g68) & (g1240) & (g1275) & (g1285)));
	assign g1313 = (((!g87) & (!g104) & (!g1242) & (g1243) & (g1274) & (!g1285)) + ((!g87) & (!g104) & (g1242) & (!g1243) & (!g1274) & (!g1285)) + ((!g87) & (!g104) & (g1242) & (!g1243) & (!g1274) & (g1285)) + ((!g87) & (!g104) & (g1242) & (!g1243) & (g1274) & (!g1285)) + ((!g87) & (!g104) & (g1242) & (!g1243) & (g1274) & (g1285)) + ((!g87) & (!g104) & (g1242) & (g1243) & (!g1274) & (!g1285)) + ((!g87) & (!g104) & (g1242) & (g1243) & (!g1274) & (g1285)) + ((!g87) & (!g104) & (g1242) & (g1243) & (g1274) & (g1285)) + ((!g87) & (g104) & (!g1242) & (!g1243) & (g1274) & (!g1285)) + ((!g87) & (g104) & (!g1242) & (g1243) & (!g1274) & (!g1285)) + ((!g87) & (g104) & (!g1242) & (g1243) & (g1274) & (!g1285)) + ((!g87) & (g104) & (g1242) & (!g1243) & (!g1274) & (!g1285)) + ((!g87) & (g104) & (g1242) & (!g1243) & (!g1274) & (g1285)) + ((!g87) & (g104) & (g1242) & (!g1243) & (g1274) & (g1285)) + ((!g87) & (g104) & (g1242) & (g1243) & (!g1274) & (g1285)) + ((!g87) & (g104) & (g1242) & (g1243) & (g1274) & (g1285)) + ((g87) & (!g104) & (!g1242) & (!g1243) & (!g1274) & (!g1285)) + ((g87) & (!g104) & (!g1242) & (!g1243) & (g1274) & (!g1285)) + ((g87) & (!g104) & (!g1242) & (g1243) & (!g1274) & (!g1285)) + ((g87) & (!g104) & (g1242) & (!g1243) & (!g1274) & (g1285)) + ((g87) & (!g104) & (g1242) & (!g1243) & (g1274) & (g1285)) + ((g87) & (!g104) & (g1242) & (g1243) & (!g1274) & (g1285)) + ((g87) & (!g104) & (g1242) & (g1243) & (g1274) & (!g1285)) + ((g87) & (!g104) & (g1242) & (g1243) & (g1274) & (g1285)) + ((g87) & (g104) & (!g1242) & (!g1243) & (!g1274) & (!g1285)) + ((g87) & (g104) & (g1242) & (!g1243) & (!g1274) & (g1285)) + ((g87) & (g104) & (g1242) & (!g1243) & (g1274) & (!g1285)) + ((g87) & (g104) & (g1242) & (!g1243) & (g1274) & (g1285)) + ((g87) & (g104) & (g1242) & (g1243) & (!g1274) & (!g1285)) + ((g87) & (g104) & (g1242) & (g1243) & (!g1274) & (g1285)) + ((g87) & (g104) & (g1242) & (g1243) & (g1274) & (!g1285)) + ((g87) & (g104) & (g1242) & (g1243) & (g1274) & (g1285)));
	assign g1314 = (((!g104) & (!g1243) & (g1274) & (!g1285)) + ((!g104) & (g1243) & (!g1274) & (!g1285)) + ((!g104) & (g1243) & (!g1274) & (g1285)) + ((!g104) & (g1243) & (g1274) & (g1285)) + ((g104) & (!g1243) & (!g1274) & (!g1285)) + ((g104) & (g1243) & (!g1274) & (g1285)) + ((g104) & (g1243) & (g1274) & (!g1285)) + ((g104) & (g1243) & (g1274) & (g1285)));
	assign g1315 = (((!g127) & (!g147) & (!g1245) & (g1246) & (g1273) & (!g1285)) + ((!g127) & (!g147) & (g1245) & (!g1246) & (!g1273) & (!g1285)) + ((!g127) & (!g147) & (g1245) & (!g1246) & (!g1273) & (g1285)) + ((!g127) & (!g147) & (g1245) & (!g1246) & (g1273) & (!g1285)) + ((!g127) & (!g147) & (g1245) & (!g1246) & (g1273) & (g1285)) + ((!g127) & (!g147) & (g1245) & (g1246) & (!g1273) & (!g1285)) + ((!g127) & (!g147) & (g1245) & (g1246) & (!g1273) & (g1285)) + ((!g127) & (!g147) & (g1245) & (g1246) & (g1273) & (g1285)) + ((!g127) & (g147) & (!g1245) & (!g1246) & (g1273) & (!g1285)) + ((!g127) & (g147) & (!g1245) & (g1246) & (!g1273) & (!g1285)) + ((!g127) & (g147) & (!g1245) & (g1246) & (g1273) & (!g1285)) + ((!g127) & (g147) & (g1245) & (!g1246) & (!g1273) & (!g1285)) + ((!g127) & (g147) & (g1245) & (!g1246) & (!g1273) & (g1285)) + ((!g127) & (g147) & (g1245) & (!g1246) & (g1273) & (g1285)) + ((!g127) & (g147) & (g1245) & (g1246) & (!g1273) & (g1285)) + ((!g127) & (g147) & (g1245) & (g1246) & (g1273) & (g1285)) + ((g127) & (!g147) & (!g1245) & (!g1246) & (!g1273) & (!g1285)) + ((g127) & (!g147) & (!g1245) & (!g1246) & (g1273) & (!g1285)) + ((g127) & (!g147) & (!g1245) & (g1246) & (!g1273) & (!g1285)) + ((g127) & (!g147) & (g1245) & (!g1246) & (!g1273) & (g1285)) + ((g127) & (!g147) & (g1245) & (!g1246) & (g1273) & (g1285)) + ((g127) & (!g147) & (g1245) & (g1246) & (!g1273) & (g1285)) + ((g127) & (!g147) & (g1245) & (g1246) & (g1273) & (!g1285)) + ((g127) & (!g147) & (g1245) & (g1246) & (g1273) & (g1285)) + ((g127) & (g147) & (!g1245) & (!g1246) & (!g1273) & (!g1285)) + ((g127) & (g147) & (g1245) & (!g1246) & (!g1273) & (g1285)) + ((g127) & (g147) & (g1245) & (!g1246) & (g1273) & (!g1285)) + ((g127) & (g147) & (g1245) & (!g1246) & (g1273) & (g1285)) + ((g127) & (g147) & (g1245) & (g1246) & (!g1273) & (!g1285)) + ((g127) & (g147) & (g1245) & (g1246) & (!g1273) & (g1285)) + ((g127) & (g147) & (g1245) & (g1246) & (g1273) & (!g1285)) + ((g127) & (g147) & (g1245) & (g1246) & (g1273) & (g1285)));
	assign g1316 = (((!g147) & (!g1246) & (g1273) & (!g1285)) + ((!g147) & (g1246) & (!g1273) & (!g1285)) + ((!g147) & (g1246) & (!g1273) & (g1285)) + ((!g147) & (g1246) & (g1273) & (g1285)) + ((g147) & (!g1246) & (!g1273) & (!g1285)) + ((g147) & (g1246) & (!g1273) & (g1285)) + ((g147) & (g1246) & (g1273) & (!g1285)) + ((g147) & (g1246) & (g1273) & (g1285)));
	assign g1317 = (((!g174) & (!g198) & (!g1248) & (g1249) & (g1272) & (!g1285)) + ((!g174) & (!g198) & (g1248) & (!g1249) & (!g1272) & (!g1285)) + ((!g174) & (!g198) & (g1248) & (!g1249) & (!g1272) & (g1285)) + ((!g174) & (!g198) & (g1248) & (!g1249) & (g1272) & (!g1285)) + ((!g174) & (!g198) & (g1248) & (!g1249) & (g1272) & (g1285)) + ((!g174) & (!g198) & (g1248) & (g1249) & (!g1272) & (!g1285)) + ((!g174) & (!g198) & (g1248) & (g1249) & (!g1272) & (g1285)) + ((!g174) & (!g198) & (g1248) & (g1249) & (g1272) & (g1285)) + ((!g174) & (g198) & (!g1248) & (!g1249) & (g1272) & (!g1285)) + ((!g174) & (g198) & (!g1248) & (g1249) & (!g1272) & (!g1285)) + ((!g174) & (g198) & (!g1248) & (g1249) & (g1272) & (!g1285)) + ((!g174) & (g198) & (g1248) & (!g1249) & (!g1272) & (!g1285)) + ((!g174) & (g198) & (g1248) & (!g1249) & (!g1272) & (g1285)) + ((!g174) & (g198) & (g1248) & (!g1249) & (g1272) & (g1285)) + ((!g174) & (g198) & (g1248) & (g1249) & (!g1272) & (g1285)) + ((!g174) & (g198) & (g1248) & (g1249) & (g1272) & (g1285)) + ((g174) & (!g198) & (!g1248) & (!g1249) & (!g1272) & (!g1285)) + ((g174) & (!g198) & (!g1248) & (!g1249) & (g1272) & (!g1285)) + ((g174) & (!g198) & (!g1248) & (g1249) & (!g1272) & (!g1285)) + ((g174) & (!g198) & (g1248) & (!g1249) & (!g1272) & (g1285)) + ((g174) & (!g198) & (g1248) & (!g1249) & (g1272) & (g1285)) + ((g174) & (!g198) & (g1248) & (g1249) & (!g1272) & (g1285)) + ((g174) & (!g198) & (g1248) & (g1249) & (g1272) & (!g1285)) + ((g174) & (!g198) & (g1248) & (g1249) & (g1272) & (g1285)) + ((g174) & (g198) & (!g1248) & (!g1249) & (!g1272) & (!g1285)) + ((g174) & (g198) & (g1248) & (!g1249) & (!g1272) & (g1285)) + ((g174) & (g198) & (g1248) & (!g1249) & (g1272) & (!g1285)) + ((g174) & (g198) & (g1248) & (!g1249) & (g1272) & (g1285)) + ((g174) & (g198) & (g1248) & (g1249) & (!g1272) & (!g1285)) + ((g174) & (g198) & (g1248) & (g1249) & (!g1272) & (g1285)) + ((g174) & (g198) & (g1248) & (g1249) & (g1272) & (!g1285)) + ((g174) & (g198) & (g1248) & (g1249) & (g1272) & (g1285)));
	assign g1318 = (((!g198) & (!g1249) & (g1272) & (!g1285)) + ((!g198) & (g1249) & (!g1272) & (!g1285)) + ((!g198) & (g1249) & (!g1272) & (g1285)) + ((!g198) & (g1249) & (g1272) & (g1285)) + ((g198) & (!g1249) & (!g1272) & (!g1285)) + ((g198) & (g1249) & (!g1272) & (g1285)) + ((g198) & (g1249) & (g1272) & (!g1285)) + ((g198) & (g1249) & (g1272) & (g1285)));
	assign g1319 = (((!g229) & (!g255) & (!g1251) & (g1252) & (g1271) & (!g1285)) + ((!g229) & (!g255) & (g1251) & (!g1252) & (!g1271) & (!g1285)) + ((!g229) & (!g255) & (g1251) & (!g1252) & (!g1271) & (g1285)) + ((!g229) & (!g255) & (g1251) & (!g1252) & (g1271) & (!g1285)) + ((!g229) & (!g255) & (g1251) & (!g1252) & (g1271) & (g1285)) + ((!g229) & (!g255) & (g1251) & (g1252) & (!g1271) & (!g1285)) + ((!g229) & (!g255) & (g1251) & (g1252) & (!g1271) & (g1285)) + ((!g229) & (!g255) & (g1251) & (g1252) & (g1271) & (g1285)) + ((!g229) & (g255) & (!g1251) & (!g1252) & (g1271) & (!g1285)) + ((!g229) & (g255) & (!g1251) & (g1252) & (!g1271) & (!g1285)) + ((!g229) & (g255) & (!g1251) & (g1252) & (g1271) & (!g1285)) + ((!g229) & (g255) & (g1251) & (!g1252) & (!g1271) & (!g1285)) + ((!g229) & (g255) & (g1251) & (!g1252) & (!g1271) & (g1285)) + ((!g229) & (g255) & (g1251) & (!g1252) & (g1271) & (g1285)) + ((!g229) & (g255) & (g1251) & (g1252) & (!g1271) & (g1285)) + ((!g229) & (g255) & (g1251) & (g1252) & (g1271) & (g1285)) + ((g229) & (!g255) & (!g1251) & (!g1252) & (!g1271) & (!g1285)) + ((g229) & (!g255) & (!g1251) & (!g1252) & (g1271) & (!g1285)) + ((g229) & (!g255) & (!g1251) & (g1252) & (!g1271) & (!g1285)) + ((g229) & (!g255) & (g1251) & (!g1252) & (!g1271) & (g1285)) + ((g229) & (!g255) & (g1251) & (!g1252) & (g1271) & (g1285)) + ((g229) & (!g255) & (g1251) & (g1252) & (!g1271) & (g1285)) + ((g229) & (!g255) & (g1251) & (g1252) & (g1271) & (!g1285)) + ((g229) & (!g255) & (g1251) & (g1252) & (g1271) & (g1285)) + ((g229) & (g255) & (!g1251) & (!g1252) & (!g1271) & (!g1285)) + ((g229) & (g255) & (g1251) & (!g1252) & (!g1271) & (g1285)) + ((g229) & (g255) & (g1251) & (!g1252) & (g1271) & (!g1285)) + ((g229) & (g255) & (g1251) & (!g1252) & (g1271) & (g1285)) + ((g229) & (g255) & (g1251) & (g1252) & (!g1271) & (!g1285)) + ((g229) & (g255) & (g1251) & (g1252) & (!g1271) & (g1285)) + ((g229) & (g255) & (g1251) & (g1252) & (g1271) & (!g1285)) + ((g229) & (g255) & (g1251) & (g1252) & (g1271) & (g1285)));
	assign g1320 = (((!g255) & (!g1252) & (g1271) & (!g1285)) + ((!g255) & (g1252) & (!g1271) & (!g1285)) + ((!g255) & (g1252) & (!g1271) & (g1285)) + ((!g255) & (g1252) & (g1271) & (g1285)) + ((g255) & (!g1252) & (!g1271) & (!g1285)) + ((g255) & (g1252) & (!g1271) & (g1285)) + ((g255) & (g1252) & (g1271) & (!g1285)) + ((g255) & (g1252) & (g1271) & (g1285)));
	assign g1321 = (((!g290) & (!g319) & (!g1254) & (g1255) & (g1270) & (!g1285)) + ((!g290) & (!g319) & (g1254) & (!g1255) & (!g1270) & (!g1285)) + ((!g290) & (!g319) & (g1254) & (!g1255) & (!g1270) & (g1285)) + ((!g290) & (!g319) & (g1254) & (!g1255) & (g1270) & (!g1285)) + ((!g290) & (!g319) & (g1254) & (!g1255) & (g1270) & (g1285)) + ((!g290) & (!g319) & (g1254) & (g1255) & (!g1270) & (!g1285)) + ((!g290) & (!g319) & (g1254) & (g1255) & (!g1270) & (g1285)) + ((!g290) & (!g319) & (g1254) & (g1255) & (g1270) & (g1285)) + ((!g290) & (g319) & (!g1254) & (!g1255) & (g1270) & (!g1285)) + ((!g290) & (g319) & (!g1254) & (g1255) & (!g1270) & (!g1285)) + ((!g290) & (g319) & (!g1254) & (g1255) & (g1270) & (!g1285)) + ((!g290) & (g319) & (g1254) & (!g1255) & (!g1270) & (!g1285)) + ((!g290) & (g319) & (g1254) & (!g1255) & (!g1270) & (g1285)) + ((!g290) & (g319) & (g1254) & (!g1255) & (g1270) & (g1285)) + ((!g290) & (g319) & (g1254) & (g1255) & (!g1270) & (g1285)) + ((!g290) & (g319) & (g1254) & (g1255) & (g1270) & (g1285)) + ((g290) & (!g319) & (!g1254) & (!g1255) & (!g1270) & (!g1285)) + ((g290) & (!g319) & (!g1254) & (!g1255) & (g1270) & (!g1285)) + ((g290) & (!g319) & (!g1254) & (g1255) & (!g1270) & (!g1285)) + ((g290) & (!g319) & (g1254) & (!g1255) & (!g1270) & (g1285)) + ((g290) & (!g319) & (g1254) & (!g1255) & (g1270) & (g1285)) + ((g290) & (!g319) & (g1254) & (g1255) & (!g1270) & (g1285)) + ((g290) & (!g319) & (g1254) & (g1255) & (g1270) & (!g1285)) + ((g290) & (!g319) & (g1254) & (g1255) & (g1270) & (g1285)) + ((g290) & (g319) & (!g1254) & (!g1255) & (!g1270) & (!g1285)) + ((g290) & (g319) & (g1254) & (!g1255) & (!g1270) & (g1285)) + ((g290) & (g319) & (g1254) & (!g1255) & (g1270) & (!g1285)) + ((g290) & (g319) & (g1254) & (!g1255) & (g1270) & (g1285)) + ((g290) & (g319) & (g1254) & (g1255) & (!g1270) & (!g1285)) + ((g290) & (g319) & (g1254) & (g1255) & (!g1270) & (g1285)) + ((g290) & (g319) & (g1254) & (g1255) & (g1270) & (!g1285)) + ((g290) & (g319) & (g1254) & (g1255) & (g1270) & (g1285)));
	assign g1322 = (((!g319) & (!g1255) & (g1270) & (!g1285)) + ((!g319) & (g1255) & (!g1270) & (!g1285)) + ((!g319) & (g1255) & (!g1270) & (g1285)) + ((!g319) & (g1255) & (g1270) & (g1285)) + ((g319) & (!g1255) & (!g1270) & (!g1285)) + ((g319) & (g1255) & (!g1270) & (g1285)) + ((g319) & (g1255) & (g1270) & (!g1285)) + ((g319) & (g1255) & (g1270) & (g1285)));
	assign g1323 = (((!g358) & (!g390) & (!g1257) & (g1258) & (g1269) & (!g1285)) + ((!g358) & (!g390) & (g1257) & (!g1258) & (!g1269) & (!g1285)) + ((!g358) & (!g390) & (g1257) & (!g1258) & (!g1269) & (g1285)) + ((!g358) & (!g390) & (g1257) & (!g1258) & (g1269) & (!g1285)) + ((!g358) & (!g390) & (g1257) & (!g1258) & (g1269) & (g1285)) + ((!g358) & (!g390) & (g1257) & (g1258) & (!g1269) & (!g1285)) + ((!g358) & (!g390) & (g1257) & (g1258) & (!g1269) & (g1285)) + ((!g358) & (!g390) & (g1257) & (g1258) & (g1269) & (g1285)) + ((!g358) & (g390) & (!g1257) & (!g1258) & (g1269) & (!g1285)) + ((!g358) & (g390) & (!g1257) & (g1258) & (!g1269) & (!g1285)) + ((!g358) & (g390) & (!g1257) & (g1258) & (g1269) & (!g1285)) + ((!g358) & (g390) & (g1257) & (!g1258) & (!g1269) & (!g1285)) + ((!g358) & (g390) & (g1257) & (!g1258) & (!g1269) & (g1285)) + ((!g358) & (g390) & (g1257) & (!g1258) & (g1269) & (g1285)) + ((!g358) & (g390) & (g1257) & (g1258) & (!g1269) & (g1285)) + ((!g358) & (g390) & (g1257) & (g1258) & (g1269) & (g1285)) + ((g358) & (!g390) & (!g1257) & (!g1258) & (!g1269) & (!g1285)) + ((g358) & (!g390) & (!g1257) & (!g1258) & (g1269) & (!g1285)) + ((g358) & (!g390) & (!g1257) & (g1258) & (!g1269) & (!g1285)) + ((g358) & (!g390) & (g1257) & (!g1258) & (!g1269) & (g1285)) + ((g358) & (!g390) & (g1257) & (!g1258) & (g1269) & (g1285)) + ((g358) & (!g390) & (g1257) & (g1258) & (!g1269) & (g1285)) + ((g358) & (!g390) & (g1257) & (g1258) & (g1269) & (!g1285)) + ((g358) & (!g390) & (g1257) & (g1258) & (g1269) & (g1285)) + ((g358) & (g390) & (!g1257) & (!g1258) & (!g1269) & (!g1285)) + ((g358) & (g390) & (g1257) & (!g1258) & (!g1269) & (g1285)) + ((g358) & (g390) & (g1257) & (!g1258) & (g1269) & (!g1285)) + ((g358) & (g390) & (g1257) & (!g1258) & (g1269) & (g1285)) + ((g358) & (g390) & (g1257) & (g1258) & (!g1269) & (!g1285)) + ((g358) & (g390) & (g1257) & (g1258) & (!g1269) & (g1285)) + ((g358) & (g390) & (g1257) & (g1258) & (g1269) & (!g1285)) + ((g358) & (g390) & (g1257) & (g1258) & (g1269) & (g1285)));
	assign g1324 = (((!g390) & (!g1258) & (g1269) & (!g1285)) + ((!g390) & (g1258) & (!g1269) & (!g1285)) + ((!g390) & (g1258) & (!g1269) & (g1285)) + ((!g390) & (g1258) & (g1269) & (g1285)) + ((g390) & (!g1258) & (!g1269) & (!g1285)) + ((g390) & (g1258) & (!g1269) & (g1285)) + ((g390) & (g1258) & (g1269) & (!g1285)) + ((g390) & (g1258) & (g1269) & (g1285)));
	assign g1325 = (((!g433) & (!g468) & (!g1260) & (g1261) & (g1268) & (!g1285)) + ((!g433) & (!g468) & (g1260) & (!g1261) & (!g1268) & (!g1285)) + ((!g433) & (!g468) & (g1260) & (!g1261) & (!g1268) & (g1285)) + ((!g433) & (!g468) & (g1260) & (!g1261) & (g1268) & (!g1285)) + ((!g433) & (!g468) & (g1260) & (!g1261) & (g1268) & (g1285)) + ((!g433) & (!g468) & (g1260) & (g1261) & (!g1268) & (!g1285)) + ((!g433) & (!g468) & (g1260) & (g1261) & (!g1268) & (g1285)) + ((!g433) & (!g468) & (g1260) & (g1261) & (g1268) & (g1285)) + ((!g433) & (g468) & (!g1260) & (!g1261) & (g1268) & (!g1285)) + ((!g433) & (g468) & (!g1260) & (g1261) & (!g1268) & (!g1285)) + ((!g433) & (g468) & (!g1260) & (g1261) & (g1268) & (!g1285)) + ((!g433) & (g468) & (g1260) & (!g1261) & (!g1268) & (!g1285)) + ((!g433) & (g468) & (g1260) & (!g1261) & (!g1268) & (g1285)) + ((!g433) & (g468) & (g1260) & (!g1261) & (g1268) & (g1285)) + ((!g433) & (g468) & (g1260) & (g1261) & (!g1268) & (g1285)) + ((!g433) & (g468) & (g1260) & (g1261) & (g1268) & (g1285)) + ((g433) & (!g468) & (!g1260) & (!g1261) & (!g1268) & (!g1285)) + ((g433) & (!g468) & (!g1260) & (!g1261) & (g1268) & (!g1285)) + ((g433) & (!g468) & (!g1260) & (g1261) & (!g1268) & (!g1285)) + ((g433) & (!g468) & (g1260) & (!g1261) & (!g1268) & (g1285)) + ((g433) & (!g468) & (g1260) & (!g1261) & (g1268) & (g1285)) + ((g433) & (!g468) & (g1260) & (g1261) & (!g1268) & (g1285)) + ((g433) & (!g468) & (g1260) & (g1261) & (g1268) & (!g1285)) + ((g433) & (!g468) & (g1260) & (g1261) & (g1268) & (g1285)) + ((g433) & (g468) & (!g1260) & (!g1261) & (!g1268) & (!g1285)) + ((g433) & (g468) & (g1260) & (!g1261) & (!g1268) & (g1285)) + ((g433) & (g468) & (g1260) & (!g1261) & (g1268) & (!g1285)) + ((g433) & (g468) & (g1260) & (!g1261) & (g1268) & (g1285)) + ((g433) & (g468) & (g1260) & (g1261) & (!g1268) & (!g1285)) + ((g433) & (g468) & (g1260) & (g1261) & (!g1268) & (g1285)) + ((g433) & (g468) & (g1260) & (g1261) & (g1268) & (!g1285)) + ((g433) & (g468) & (g1260) & (g1261) & (g1268) & (g1285)));
	assign g1326 = (((!g468) & (!g1261) & (g1268) & (!g1285)) + ((!g468) & (g1261) & (!g1268) & (!g1285)) + ((!g468) & (g1261) & (!g1268) & (g1285)) + ((!g468) & (g1261) & (g1268) & (g1285)) + ((g468) & (!g1261) & (!g1268) & (!g1285)) + ((g468) & (g1261) & (!g1268) & (g1285)) + ((g468) & (g1261) & (g1268) & (!g1285)) + ((g468) & (g1261) & (g1268) & (g1285)));
	assign g1327 = (((!g515) & (!g553) & (!g1263) & (g1264) & (g1267) & (!g1285)) + ((!g515) & (!g553) & (g1263) & (!g1264) & (!g1267) & (!g1285)) + ((!g515) & (!g553) & (g1263) & (!g1264) & (!g1267) & (g1285)) + ((!g515) & (!g553) & (g1263) & (!g1264) & (g1267) & (!g1285)) + ((!g515) & (!g553) & (g1263) & (!g1264) & (g1267) & (g1285)) + ((!g515) & (!g553) & (g1263) & (g1264) & (!g1267) & (!g1285)) + ((!g515) & (!g553) & (g1263) & (g1264) & (!g1267) & (g1285)) + ((!g515) & (!g553) & (g1263) & (g1264) & (g1267) & (g1285)) + ((!g515) & (g553) & (!g1263) & (!g1264) & (g1267) & (!g1285)) + ((!g515) & (g553) & (!g1263) & (g1264) & (!g1267) & (!g1285)) + ((!g515) & (g553) & (!g1263) & (g1264) & (g1267) & (!g1285)) + ((!g515) & (g553) & (g1263) & (!g1264) & (!g1267) & (!g1285)) + ((!g515) & (g553) & (g1263) & (!g1264) & (!g1267) & (g1285)) + ((!g515) & (g553) & (g1263) & (!g1264) & (g1267) & (g1285)) + ((!g515) & (g553) & (g1263) & (g1264) & (!g1267) & (g1285)) + ((!g515) & (g553) & (g1263) & (g1264) & (g1267) & (g1285)) + ((g515) & (!g553) & (!g1263) & (!g1264) & (!g1267) & (!g1285)) + ((g515) & (!g553) & (!g1263) & (!g1264) & (g1267) & (!g1285)) + ((g515) & (!g553) & (!g1263) & (g1264) & (!g1267) & (!g1285)) + ((g515) & (!g553) & (g1263) & (!g1264) & (!g1267) & (g1285)) + ((g515) & (!g553) & (g1263) & (!g1264) & (g1267) & (g1285)) + ((g515) & (!g553) & (g1263) & (g1264) & (!g1267) & (g1285)) + ((g515) & (!g553) & (g1263) & (g1264) & (g1267) & (!g1285)) + ((g515) & (!g553) & (g1263) & (g1264) & (g1267) & (g1285)) + ((g515) & (g553) & (!g1263) & (!g1264) & (!g1267) & (!g1285)) + ((g515) & (g553) & (g1263) & (!g1264) & (!g1267) & (g1285)) + ((g515) & (g553) & (g1263) & (!g1264) & (g1267) & (!g1285)) + ((g515) & (g553) & (g1263) & (!g1264) & (g1267) & (g1285)) + ((g515) & (g553) & (g1263) & (g1264) & (!g1267) & (!g1285)) + ((g515) & (g553) & (g1263) & (g1264) & (!g1267) & (g1285)) + ((g515) & (g553) & (g1263) & (g1264) & (g1267) & (!g1285)) + ((g515) & (g553) & (g1263) & (g1264) & (g1267) & (g1285)));
	assign g1328 = (((!g553) & (!g1264) & (g1267) & (!g1285)) + ((!g553) & (g1264) & (!g1267) & (!g1285)) + ((!g553) & (g1264) & (!g1267) & (g1285)) + ((!g553) & (g1264) & (g1267) & (g1285)) + ((g553) & (!g1264) & (!g1267) & (!g1285)) + ((g553) & (g1264) & (!g1267) & (g1285)) + ((g553) & (g1264) & (g1267) & (!g1285)) + ((g553) & (g1264) & (g1267) & (g1285)));
	assign g1329 = (((!g604) & (!g645) & (!g1266) & (g1211) & (g1229) & (!g1285)) + ((!g604) & (!g645) & (g1266) & (!g1211) & (!g1229) & (!g1285)) + ((!g604) & (!g645) & (g1266) & (!g1211) & (!g1229) & (g1285)) + ((!g604) & (!g645) & (g1266) & (!g1211) & (g1229) & (!g1285)) + ((!g604) & (!g645) & (g1266) & (!g1211) & (g1229) & (g1285)) + ((!g604) & (!g645) & (g1266) & (g1211) & (!g1229) & (!g1285)) + ((!g604) & (!g645) & (g1266) & (g1211) & (!g1229) & (g1285)) + ((!g604) & (!g645) & (g1266) & (g1211) & (g1229) & (g1285)) + ((!g604) & (g645) & (!g1266) & (!g1211) & (g1229) & (!g1285)) + ((!g604) & (g645) & (!g1266) & (g1211) & (!g1229) & (!g1285)) + ((!g604) & (g645) & (!g1266) & (g1211) & (g1229) & (!g1285)) + ((!g604) & (g645) & (g1266) & (!g1211) & (!g1229) & (!g1285)) + ((!g604) & (g645) & (g1266) & (!g1211) & (!g1229) & (g1285)) + ((!g604) & (g645) & (g1266) & (!g1211) & (g1229) & (g1285)) + ((!g604) & (g645) & (g1266) & (g1211) & (!g1229) & (g1285)) + ((!g604) & (g645) & (g1266) & (g1211) & (g1229) & (g1285)) + ((g604) & (!g645) & (!g1266) & (!g1211) & (!g1229) & (!g1285)) + ((g604) & (!g645) & (!g1266) & (!g1211) & (g1229) & (!g1285)) + ((g604) & (!g645) & (!g1266) & (g1211) & (!g1229) & (!g1285)) + ((g604) & (!g645) & (g1266) & (!g1211) & (!g1229) & (g1285)) + ((g604) & (!g645) & (g1266) & (!g1211) & (g1229) & (g1285)) + ((g604) & (!g645) & (g1266) & (g1211) & (!g1229) & (g1285)) + ((g604) & (!g645) & (g1266) & (g1211) & (g1229) & (!g1285)) + ((g604) & (!g645) & (g1266) & (g1211) & (g1229) & (g1285)) + ((g604) & (g645) & (!g1266) & (!g1211) & (!g1229) & (!g1285)) + ((g604) & (g645) & (g1266) & (!g1211) & (!g1229) & (g1285)) + ((g604) & (g645) & (g1266) & (!g1211) & (g1229) & (!g1285)) + ((g604) & (g645) & (g1266) & (!g1211) & (g1229) & (g1285)) + ((g604) & (g645) & (g1266) & (g1211) & (!g1229) & (!g1285)) + ((g604) & (g645) & (g1266) & (g1211) & (!g1229) & (g1285)) + ((g604) & (g645) & (g1266) & (g1211) & (g1229) & (!g1285)) + ((g604) & (g645) & (g1266) & (g1211) & (g1229) & (g1285)));
	assign g1330 = (((!g553) & (!g604) & (g1329) & (g1286) & (g1304)) + ((!g553) & (g604) & (g1329) & (!g1286) & (g1304)) + ((!g553) & (g604) & (g1329) & (g1286) & (!g1304)) + ((!g553) & (g604) & (g1329) & (g1286) & (g1304)) + ((g553) & (!g604) & (!g1329) & (g1286) & (g1304)) + ((g553) & (!g604) & (g1329) & (!g1286) & (!g1304)) + ((g553) & (!g604) & (g1329) & (!g1286) & (g1304)) + ((g553) & (!g604) & (g1329) & (g1286) & (!g1304)) + ((g553) & (!g604) & (g1329) & (g1286) & (g1304)) + ((g553) & (g604) & (!g1329) & (!g1286) & (g1304)) + ((g553) & (g604) & (!g1329) & (g1286) & (!g1304)) + ((g553) & (g604) & (!g1329) & (g1286) & (g1304)) + ((g553) & (g604) & (g1329) & (!g1286) & (!g1304)) + ((g553) & (g604) & (g1329) & (!g1286) & (g1304)) + ((g553) & (g604) & (g1329) & (g1286) & (!g1304)) + ((g553) & (g604) & (g1329) & (g1286) & (g1304)));
	assign g1331 = (((!g468) & (!g515) & (g1327) & (g1328) & (g1330)) + ((!g468) & (g515) & (g1327) & (!g1328) & (g1330)) + ((!g468) & (g515) & (g1327) & (g1328) & (!g1330)) + ((!g468) & (g515) & (g1327) & (g1328) & (g1330)) + ((g468) & (!g515) & (!g1327) & (g1328) & (g1330)) + ((g468) & (!g515) & (g1327) & (!g1328) & (!g1330)) + ((g468) & (!g515) & (g1327) & (!g1328) & (g1330)) + ((g468) & (!g515) & (g1327) & (g1328) & (!g1330)) + ((g468) & (!g515) & (g1327) & (g1328) & (g1330)) + ((g468) & (g515) & (!g1327) & (!g1328) & (g1330)) + ((g468) & (g515) & (!g1327) & (g1328) & (!g1330)) + ((g468) & (g515) & (!g1327) & (g1328) & (g1330)) + ((g468) & (g515) & (g1327) & (!g1328) & (!g1330)) + ((g468) & (g515) & (g1327) & (!g1328) & (g1330)) + ((g468) & (g515) & (g1327) & (g1328) & (!g1330)) + ((g468) & (g515) & (g1327) & (g1328) & (g1330)));
	assign g1332 = (((!g390) & (!g433) & (g1325) & (g1326) & (g1331)) + ((!g390) & (g433) & (g1325) & (!g1326) & (g1331)) + ((!g390) & (g433) & (g1325) & (g1326) & (!g1331)) + ((!g390) & (g433) & (g1325) & (g1326) & (g1331)) + ((g390) & (!g433) & (!g1325) & (g1326) & (g1331)) + ((g390) & (!g433) & (g1325) & (!g1326) & (!g1331)) + ((g390) & (!g433) & (g1325) & (!g1326) & (g1331)) + ((g390) & (!g433) & (g1325) & (g1326) & (!g1331)) + ((g390) & (!g433) & (g1325) & (g1326) & (g1331)) + ((g390) & (g433) & (!g1325) & (!g1326) & (g1331)) + ((g390) & (g433) & (!g1325) & (g1326) & (!g1331)) + ((g390) & (g433) & (!g1325) & (g1326) & (g1331)) + ((g390) & (g433) & (g1325) & (!g1326) & (!g1331)) + ((g390) & (g433) & (g1325) & (!g1326) & (g1331)) + ((g390) & (g433) & (g1325) & (g1326) & (!g1331)) + ((g390) & (g433) & (g1325) & (g1326) & (g1331)));
	assign g1333 = (((!g319) & (!g358) & (g1323) & (g1324) & (g1332)) + ((!g319) & (g358) & (g1323) & (!g1324) & (g1332)) + ((!g319) & (g358) & (g1323) & (g1324) & (!g1332)) + ((!g319) & (g358) & (g1323) & (g1324) & (g1332)) + ((g319) & (!g358) & (!g1323) & (g1324) & (g1332)) + ((g319) & (!g358) & (g1323) & (!g1324) & (!g1332)) + ((g319) & (!g358) & (g1323) & (!g1324) & (g1332)) + ((g319) & (!g358) & (g1323) & (g1324) & (!g1332)) + ((g319) & (!g358) & (g1323) & (g1324) & (g1332)) + ((g319) & (g358) & (!g1323) & (!g1324) & (g1332)) + ((g319) & (g358) & (!g1323) & (g1324) & (!g1332)) + ((g319) & (g358) & (!g1323) & (g1324) & (g1332)) + ((g319) & (g358) & (g1323) & (!g1324) & (!g1332)) + ((g319) & (g358) & (g1323) & (!g1324) & (g1332)) + ((g319) & (g358) & (g1323) & (g1324) & (!g1332)) + ((g319) & (g358) & (g1323) & (g1324) & (g1332)));
	assign g1334 = (((!g255) & (!g290) & (g1321) & (g1322) & (g1333)) + ((!g255) & (g290) & (g1321) & (!g1322) & (g1333)) + ((!g255) & (g290) & (g1321) & (g1322) & (!g1333)) + ((!g255) & (g290) & (g1321) & (g1322) & (g1333)) + ((g255) & (!g290) & (!g1321) & (g1322) & (g1333)) + ((g255) & (!g290) & (g1321) & (!g1322) & (!g1333)) + ((g255) & (!g290) & (g1321) & (!g1322) & (g1333)) + ((g255) & (!g290) & (g1321) & (g1322) & (!g1333)) + ((g255) & (!g290) & (g1321) & (g1322) & (g1333)) + ((g255) & (g290) & (!g1321) & (!g1322) & (g1333)) + ((g255) & (g290) & (!g1321) & (g1322) & (!g1333)) + ((g255) & (g290) & (!g1321) & (g1322) & (g1333)) + ((g255) & (g290) & (g1321) & (!g1322) & (!g1333)) + ((g255) & (g290) & (g1321) & (!g1322) & (g1333)) + ((g255) & (g290) & (g1321) & (g1322) & (!g1333)) + ((g255) & (g290) & (g1321) & (g1322) & (g1333)));
	assign g1335 = (((!g198) & (!g229) & (g1319) & (g1320) & (g1334)) + ((!g198) & (g229) & (g1319) & (!g1320) & (g1334)) + ((!g198) & (g229) & (g1319) & (g1320) & (!g1334)) + ((!g198) & (g229) & (g1319) & (g1320) & (g1334)) + ((g198) & (!g229) & (!g1319) & (g1320) & (g1334)) + ((g198) & (!g229) & (g1319) & (!g1320) & (!g1334)) + ((g198) & (!g229) & (g1319) & (!g1320) & (g1334)) + ((g198) & (!g229) & (g1319) & (g1320) & (!g1334)) + ((g198) & (!g229) & (g1319) & (g1320) & (g1334)) + ((g198) & (g229) & (!g1319) & (!g1320) & (g1334)) + ((g198) & (g229) & (!g1319) & (g1320) & (!g1334)) + ((g198) & (g229) & (!g1319) & (g1320) & (g1334)) + ((g198) & (g229) & (g1319) & (!g1320) & (!g1334)) + ((g198) & (g229) & (g1319) & (!g1320) & (g1334)) + ((g198) & (g229) & (g1319) & (g1320) & (!g1334)) + ((g198) & (g229) & (g1319) & (g1320) & (g1334)));
	assign g1336 = (((!g147) & (!g174) & (g1317) & (g1318) & (g1335)) + ((!g147) & (g174) & (g1317) & (!g1318) & (g1335)) + ((!g147) & (g174) & (g1317) & (g1318) & (!g1335)) + ((!g147) & (g174) & (g1317) & (g1318) & (g1335)) + ((g147) & (!g174) & (!g1317) & (g1318) & (g1335)) + ((g147) & (!g174) & (g1317) & (!g1318) & (!g1335)) + ((g147) & (!g174) & (g1317) & (!g1318) & (g1335)) + ((g147) & (!g174) & (g1317) & (g1318) & (!g1335)) + ((g147) & (!g174) & (g1317) & (g1318) & (g1335)) + ((g147) & (g174) & (!g1317) & (!g1318) & (g1335)) + ((g147) & (g174) & (!g1317) & (g1318) & (!g1335)) + ((g147) & (g174) & (!g1317) & (g1318) & (g1335)) + ((g147) & (g174) & (g1317) & (!g1318) & (!g1335)) + ((g147) & (g174) & (g1317) & (!g1318) & (g1335)) + ((g147) & (g174) & (g1317) & (g1318) & (!g1335)) + ((g147) & (g174) & (g1317) & (g1318) & (g1335)));
	assign g1337 = (((!g104) & (!g127) & (g1315) & (g1316) & (g1336)) + ((!g104) & (g127) & (g1315) & (!g1316) & (g1336)) + ((!g104) & (g127) & (g1315) & (g1316) & (!g1336)) + ((!g104) & (g127) & (g1315) & (g1316) & (g1336)) + ((g104) & (!g127) & (!g1315) & (g1316) & (g1336)) + ((g104) & (!g127) & (g1315) & (!g1316) & (!g1336)) + ((g104) & (!g127) & (g1315) & (!g1316) & (g1336)) + ((g104) & (!g127) & (g1315) & (g1316) & (!g1336)) + ((g104) & (!g127) & (g1315) & (g1316) & (g1336)) + ((g104) & (g127) & (!g1315) & (!g1316) & (g1336)) + ((g104) & (g127) & (!g1315) & (g1316) & (!g1336)) + ((g104) & (g127) & (!g1315) & (g1316) & (g1336)) + ((g104) & (g127) & (g1315) & (!g1316) & (!g1336)) + ((g104) & (g127) & (g1315) & (!g1316) & (g1336)) + ((g104) & (g127) & (g1315) & (g1316) & (!g1336)) + ((g104) & (g127) & (g1315) & (g1316) & (g1336)));
	assign g1338 = (((!g68) & (!g87) & (g1313) & (g1314) & (g1337)) + ((!g68) & (g87) & (g1313) & (!g1314) & (g1337)) + ((!g68) & (g87) & (g1313) & (g1314) & (!g1337)) + ((!g68) & (g87) & (g1313) & (g1314) & (g1337)) + ((g68) & (!g87) & (!g1313) & (g1314) & (g1337)) + ((g68) & (!g87) & (g1313) & (!g1314) & (!g1337)) + ((g68) & (!g87) & (g1313) & (!g1314) & (g1337)) + ((g68) & (!g87) & (g1313) & (g1314) & (!g1337)) + ((g68) & (!g87) & (g1313) & (g1314) & (g1337)) + ((g68) & (g87) & (!g1313) & (!g1314) & (g1337)) + ((g68) & (g87) & (!g1313) & (g1314) & (!g1337)) + ((g68) & (g87) & (!g1313) & (g1314) & (g1337)) + ((g68) & (g87) & (g1313) & (!g1314) & (!g1337)) + ((g68) & (g87) & (g1313) & (!g1314) & (g1337)) + ((g68) & (g87) & (g1313) & (g1314) & (!g1337)) + ((g68) & (g87) & (g1313) & (g1314) & (g1337)));
	assign g1339 = (((!g39) & (!g54) & (g1311) & (g1312) & (g1338)) + ((!g39) & (g54) & (g1311) & (!g1312) & (g1338)) + ((!g39) & (g54) & (g1311) & (g1312) & (!g1338)) + ((!g39) & (g54) & (g1311) & (g1312) & (g1338)) + ((g39) & (!g54) & (!g1311) & (g1312) & (g1338)) + ((g39) & (!g54) & (g1311) & (!g1312) & (!g1338)) + ((g39) & (!g54) & (g1311) & (!g1312) & (g1338)) + ((g39) & (!g54) & (g1311) & (g1312) & (!g1338)) + ((g39) & (!g54) & (g1311) & (g1312) & (g1338)) + ((g39) & (g54) & (!g1311) & (!g1312) & (g1338)) + ((g39) & (g54) & (!g1311) & (g1312) & (!g1338)) + ((g39) & (g54) & (!g1311) & (g1312) & (g1338)) + ((g39) & (g54) & (g1311) & (!g1312) & (!g1338)) + ((g39) & (g54) & (g1311) & (!g1312) & (g1338)) + ((g39) & (g54) & (g1311) & (g1312) & (!g1338)) + ((g39) & (g54) & (g1311) & (g1312) & (g1338)));
	assign g1340 = (((!g18) & (!g27) & (g1309) & (g1310) & (g1339)) + ((!g18) & (g27) & (g1309) & (!g1310) & (g1339)) + ((!g18) & (g27) & (g1309) & (g1310) & (!g1339)) + ((!g18) & (g27) & (g1309) & (g1310) & (g1339)) + ((g18) & (!g27) & (!g1309) & (g1310) & (g1339)) + ((g18) & (!g27) & (g1309) & (!g1310) & (!g1339)) + ((g18) & (!g27) & (g1309) & (!g1310) & (g1339)) + ((g18) & (!g27) & (g1309) & (g1310) & (!g1339)) + ((g18) & (!g27) & (g1309) & (g1310) & (g1339)) + ((g18) & (g27) & (!g1309) & (!g1310) & (g1339)) + ((g18) & (g27) & (!g1309) & (g1310) & (!g1339)) + ((g18) & (g27) & (!g1309) & (g1310) & (g1339)) + ((g18) & (g27) & (g1309) & (!g1310) & (!g1339)) + ((g18) & (g27) & (g1309) & (!g1310) & (g1339)) + ((g18) & (g27) & (g1309) & (g1310) & (!g1339)) + ((g18) & (g27) & (g1309) & (g1310) & (g1339)));
	assign g1341 = (((!g2) & (!g8) & (g1307) & (g1308) & (g1340)) + ((!g2) & (g8) & (g1307) & (!g1308) & (g1340)) + ((!g2) & (g8) & (g1307) & (g1308) & (!g1340)) + ((!g2) & (g8) & (g1307) & (g1308) & (g1340)) + ((g2) & (!g8) & (!g1307) & (g1308) & (g1340)) + ((g2) & (!g8) & (g1307) & (!g1308) & (!g1340)) + ((g2) & (!g8) & (g1307) & (!g1308) & (g1340)) + ((g2) & (!g8) & (g1307) & (g1308) & (!g1340)) + ((g2) & (!g8) & (g1307) & (g1308) & (g1340)) + ((g2) & (g8) & (!g1307) & (!g1308) & (g1340)) + ((g2) & (g8) & (!g1307) & (g1308) & (!g1340)) + ((g2) & (g8) & (!g1307) & (g1308) & (g1340)) + ((g2) & (g8) & (g1307) & (!g1308) & (!g1340)) + ((g2) & (g8) & (g1307) & (!g1308) & (g1340)) + ((g2) & (g8) & (g1307) & (g1308) & (!g1340)) + ((g2) & (g8) & (g1307) & (g1308) & (g1340)));
	assign g1342 = (((!g2) & (!g1231) & (g1278) & (!g1285)) + ((!g2) & (g1231) & (!g1278) & (!g1285)) + ((!g2) & (g1231) & (!g1278) & (g1285)) + ((!g2) & (g1231) & (g1278) & (g1285)) + ((g2) & (!g1231) & (!g1278) & (!g1285)) + ((g2) & (g1231) & (!g1278) & (g1285)) + ((g2) & (g1231) & (g1278) & (!g1285)) + ((g2) & (g1231) & (g1278) & (g1285)));
	assign g1343 = (((!g1) & (!g1230) & (!g1281) & (!g1283) & (g1284)) + ((!g1) & (!g1230) & (!g1281) & (g1283) & (!g1284)) + ((!g1) & (!g1230) & (!g1281) & (g1283) & (g1284)) + ((!g1) & (g1230) & (g1281) & (!g1283) & (!g1284)) + ((!g1) & (g1230) & (g1281) & (!g1283) & (g1284)) + ((!g1) & (g1230) & (g1281) & (g1283) & (!g1284)) + ((!g1) & (g1230) & (g1281) & (g1283) & (g1284)) + ((g1) & (!g1230) & (!g1281) & (!g1283) & (g1284)) + ((g1) & (!g1230) & (!g1281) & (g1283) & (g1284)) + ((g1) & (g1230) & (g1281) & (!g1283) & (!g1284)) + ((g1) & (g1230) & (g1281) & (!g1283) & (g1284)) + ((g1) & (g1230) & (g1281) & (g1283) & (!g1284)) + ((g1) & (g1230) & (g1281) & (g1283) & (g1284)));
	assign g1344 = (((!g4) & (!g1) & (!g1306) & (!g1341) & (!g1342) & (!g1343)) + ((!g4) & (g1) & (!g1306) & (!g1341) & (!g1342) & (!g1343)) + ((!g4) & (g1) & (!g1306) & (!g1341) & (!g1342) & (g1343)) + ((!g4) & (g1) & (!g1306) & (!g1341) & (g1342) & (!g1343)) + ((!g4) & (g1) & (!g1306) & (!g1341) & (g1342) & (g1343)) + ((!g4) & (g1) & (!g1306) & (g1341) & (!g1342) & (!g1343)) + ((!g4) & (g1) & (!g1306) & (g1341) & (!g1342) & (g1343)) + ((!g4) & (g1) & (!g1306) & (g1341) & (g1342) & (!g1343)) + ((!g4) & (g1) & (!g1306) & (g1341) & (g1342) & (g1343)) + ((!g4) & (g1) & (g1306) & (!g1341) & (!g1342) & (!g1343)) + ((!g4) & (g1) & (g1306) & (!g1341) & (!g1342) & (g1343)) + ((g4) & (!g1) & (!g1306) & (!g1341) & (!g1342) & (!g1343)) + ((g4) & (!g1) & (!g1306) & (!g1341) & (g1342) & (!g1343)) + ((g4) & (!g1) & (!g1306) & (g1341) & (!g1342) & (!g1343)) + ((g4) & (g1) & (!g1306) & (!g1341) & (!g1342) & (!g1343)) + ((g4) & (g1) & (!g1306) & (!g1341) & (!g1342) & (g1343)) + ((g4) & (g1) & (!g1306) & (!g1341) & (g1342) & (!g1343)) + ((g4) & (g1) & (!g1306) & (!g1341) & (g1342) & (g1343)) + ((g4) & (g1) & (!g1306) & (g1341) & (!g1342) & (!g1343)) + ((g4) & (g1) & (!g1306) & (g1341) & (!g1342) & (g1343)) + ((g4) & (g1) & (!g1306) & (g1341) & (g1342) & (!g1343)) + ((g4) & (g1) & (!g1306) & (g1341) & (g1342) & (g1343)) + ((g4) & (g1) & (g1306) & (!g1341) & (!g1342) & (!g1343)) + ((g4) & (g1) & (g1306) & (!g1341) & (!g1342) & (g1343)) + ((g4) & (g1) & (g1306) & (!g1341) & (g1342) & (!g1343)) + ((g4) & (g1) & (g1306) & (!g1341) & (g1342) & (g1343)) + ((g4) & (g1) & (g1306) & (g1341) & (!g1342) & (!g1343)) + ((g4) & (g1) & (g1306) & (g1341) & (!g1342) & (g1343)));
	assign g1345 = (((!g604) & (!g1286) & (g1304) & (!g1305) & (!g1344)) + ((!g604) & (!g1286) & (g1304) & (g1305) & (!g1344)) + ((!g604) & (!g1286) & (g1304) & (g1305) & (g1344)) + ((!g604) & (g1286) & (!g1304) & (!g1305) & (!g1344)) + ((!g604) & (g1286) & (!g1304) & (!g1305) & (g1344)) + ((!g604) & (g1286) & (!g1304) & (g1305) & (!g1344)) + ((!g604) & (g1286) & (!g1304) & (g1305) & (g1344)) + ((!g604) & (g1286) & (g1304) & (!g1305) & (g1344)) + ((g604) & (!g1286) & (!g1304) & (!g1305) & (!g1344)) + ((g604) & (!g1286) & (!g1304) & (g1305) & (!g1344)) + ((g604) & (!g1286) & (!g1304) & (g1305) & (g1344)) + ((g604) & (g1286) & (!g1304) & (!g1305) & (g1344)) + ((g604) & (g1286) & (g1304) & (!g1305) & (!g1344)) + ((g604) & (g1286) & (g1304) & (!g1305) & (g1344)) + ((g604) & (g1286) & (g1304) & (g1305) & (!g1344)) + ((g604) & (g1286) & (g1304) & (g1305) & (g1344)));
	assign g1346 = (((!g645) & (!g700) & (g1288) & (g1303)) + ((!g645) & (g700) & (!g1288) & (g1303)) + ((!g645) & (g700) & (g1288) & (!g1303)) + ((!g645) & (g700) & (g1288) & (g1303)) + ((g645) & (!g700) & (!g1288) & (!g1303)) + ((g645) & (!g700) & (!g1288) & (g1303)) + ((g645) & (!g700) & (g1288) & (!g1303)) + ((g645) & (g700) & (!g1288) & (!g1303)));
	assign g1347 = (((!g1287) & (!g1305) & (!g1344) & (g1346)) + ((!g1287) & (g1305) & (!g1344) & (g1346)) + ((!g1287) & (g1305) & (g1344) & (g1346)) + ((g1287) & (!g1305) & (!g1344) & (!g1346)) + ((g1287) & (!g1305) & (g1344) & (!g1346)) + ((g1287) & (!g1305) & (g1344) & (g1346)) + ((g1287) & (g1305) & (!g1344) & (!g1346)) + ((g1287) & (g1305) & (g1344) & (!g1346)));
	assign g1348 = (((!g700) & (!g1288) & (g1303) & (!g1305) & (!g1344)) + ((!g700) & (!g1288) & (g1303) & (g1305) & (!g1344)) + ((!g700) & (!g1288) & (g1303) & (g1305) & (g1344)) + ((!g700) & (g1288) & (!g1303) & (!g1305) & (!g1344)) + ((!g700) & (g1288) & (!g1303) & (!g1305) & (g1344)) + ((!g700) & (g1288) & (!g1303) & (g1305) & (!g1344)) + ((!g700) & (g1288) & (!g1303) & (g1305) & (g1344)) + ((!g700) & (g1288) & (g1303) & (!g1305) & (g1344)) + ((g700) & (!g1288) & (!g1303) & (!g1305) & (!g1344)) + ((g700) & (!g1288) & (!g1303) & (g1305) & (!g1344)) + ((g700) & (!g1288) & (!g1303) & (g1305) & (g1344)) + ((g700) & (g1288) & (!g1303) & (!g1305) & (g1344)) + ((g700) & (g1288) & (g1303) & (!g1305) & (!g1344)) + ((g700) & (g1288) & (g1303) & (!g1305) & (g1344)) + ((g700) & (g1288) & (g1303) & (g1305) & (!g1344)) + ((g700) & (g1288) & (g1303) & (g1305) & (g1344)));
	assign g1349 = (((!g744) & (!g803) & (g1290) & (g1302)) + ((!g744) & (g803) & (!g1290) & (g1302)) + ((!g744) & (g803) & (g1290) & (!g1302)) + ((!g744) & (g803) & (g1290) & (g1302)) + ((g744) & (!g803) & (!g1290) & (!g1302)) + ((g744) & (!g803) & (!g1290) & (g1302)) + ((g744) & (!g803) & (g1290) & (!g1302)) + ((g744) & (g803) & (!g1290) & (!g1302)));
	assign g1350 = (((!g1289) & (!g1305) & (!g1344) & (g1349)) + ((!g1289) & (g1305) & (!g1344) & (g1349)) + ((!g1289) & (g1305) & (g1344) & (g1349)) + ((g1289) & (!g1305) & (!g1344) & (!g1349)) + ((g1289) & (!g1305) & (g1344) & (!g1349)) + ((g1289) & (!g1305) & (g1344) & (g1349)) + ((g1289) & (g1305) & (!g1344) & (!g1349)) + ((g1289) & (g1305) & (g1344) & (!g1349)));
	assign g1351 = (((!g803) & (!g1290) & (g1302) & (!g1305) & (!g1344)) + ((!g803) & (!g1290) & (g1302) & (g1305) & (!g1344)) + ((!g803) & (!g1290) & (g1302) & (g1305) & (g1344)) + ((!g803) & (g1290) & (!g1302) & (!g1305) & (!g1344)) + ((!g803) & (g1290) & (!g1302) & (!g1305) & (g1344)) + ((!g803) & (g1290) & (!g1302) & (g1305) & (!g1344)) + ((!g803) & (g1290) & (!g1302) & (g1305) & (g1344)) + ((!g803) & (g1290) & (g1302) & (!g1305) & (g1344)) + ((g803) & (!g1290) & (!g1302) & (!g1305) & (!g1344)) + ((g803) & (!g1290) & (!g1302) & (g1305) & (!g1344)) + ((g803) & (!g1290) & (!g1302) & (g1305) & (g1344)) + ((g803) & (g1290) & (!g1302) & (!g1305) & (g1344)) + ((g803) & (g1290) & (g1302) & (!g1305) & (!g1344)) + ((g803) & (g1290) & (g1302) & (!g1305) & (g1344)) + ((g803) & (g1290) & (g1302) & (g1305) & (!g1344)) + ((g803) & (g1290) & (g1302) & (g1305) & (g1344)));
	assign g1352 = (((!g851) & (!g914) & (g1292) & (g1301)) + ((!g851) & (g914) & (!g1292) & (g1301)) + ((!g851) & (g914) & (g1292) & (!g1301)) + ((!g851) & (g914) & (g1292) & (g1301)) + ((g851) & (!g914) & (!g1292) & (!g1301)) + ((g851) & (!g914) & (!g1292) & (g1301)) + ((g851) & (!g914) & (g1292) & (!g1301)) + ((g851) & (g914) & (!g1292) & (!g1301)));
	assign g1353 = (((!g1291) & (!g1305) & (!g1344) & (g1352)) + ((!g1291) & (g1305) & (!g1344) & (g1352)) + ((!g1291) & (g1305) & (g1344) & (g1352)) + ((g1291) & (!g1305) & (!g1344) & (!g1352)) + ((g1291) & (!g1305) & (g1344) & (!g1352)) + ((g1291) & (!g1305) & (g1344) & (g1352)) + ((g1291) & (g1305) & (!g1344) & (!g1352)) + ((g1291) & (g1305) & (g1344) & (!g1352)));
	assign g1354 = (((!g914) & (!g1292) & (g1301) & (!g1305) & (!g1344)) + ((!g914) & (!g1292) & (g1301) & (g1305) & (!g1344)) + ((!g914) & (!g1292) & (g1301) & (g1305) & (g1344)) + ((!g914) & (g1292) & (!g1301) & (!g1305) & (!g1344)) + ((!g914) & (g1292) & (!g1301) & (!g1305) & (g1344)) + ((!g914) & (g1292) & (!g1301) & (g1305) & (!g1344)) + ((!g914) & (g1292) & (!g1301) & (g1305) & (g1344)) + ((!g914) & (g1292) & (g1301) & (!g1305) & (g1344)) + ((g914) & (!g1292) & (!g1301) & (!g1305) & (!g1344)) + ((g914) & (!g1292) & (!g1301) & (g1305) & (!g1344)) + ((g914) & (!g1292) & (!g1301) & (g1305) & (g1344)) + ((g914) & (g1292) & (!g1301) & (!g1305) & (g1344)) + ((g914) & (g1292) & (g1301) & (!g1305) & (!g1344)) + ((g914) & (g1292) & (g1301) & (!g1305) & (g1344)) + ((g914) & (g1292) & (g1301) & (g1305) & (!g1344)) + ((g914) & (g1292) & (g1301) & (g1305) & (g1344)));
	assign g1355 = (((!g1032) & (!g1030) & (g1294) & (g1300)) + ((!g1032) & (g1030) & (!g1294) & (g1300)) + ((!g1032) & (g1030) & (g1294) & (!g1300)) + ((!g1032) & (g1030) & (g1294) & (g1300)) + ((g1032) & (!g1030) & (!g1294) & (!g1300)) + ((g1032) & (!g1030) & (!g1294) & (g1300)) + ((g1032) & (!g1030) & (g1294) & (!g1300)) + ((g1032) & (g1030) & (!g1294) & (!g1300)));
	assign g1356 = (((!g1293) & (!g1305) & (!g1344) & (g1355)) + ((!g1293) & (g1305) & (!g1344) & (g1355)) + ((!g1293) & (g1305) & (g1344) & (g1355)) + ((g1293) & (!g1305) & (!g1344) & (!g1355)) + ((g1293) & (!g1305) & (g1344) & (!g1355)) + ((g1293) & (!g1305) & (g1344) & (g1355)) + ((g1293) & (g1305) & (!g1344) & (!g1355)) + ((g1293) & (g1305) & (g1344) & (!g1355)));
	assign g1357 = (((!g1030) & (!g1294) & (g1300) & (!g1305) & (!g1344)) + ((!g1030) & (!g1294) & (g1300) & (g1305) & (!g1344)) + ((!g1030) & (!g1294) & (g1300) & (g1305) & (g1344)) + ((!g1030) & (g1294) & (!g1300) & (!g1305) & (!g1344)) + ((!g1030) & (g1294) & (!g1300) & (!g1305) & (g1344)) + ((!g1030) & (g1294) & (!g1300) & (g1305) & (!g1344)) + ((!g1030) & (g1294) & (!g1300) & (g1305) & (g1344)) + ((!g1030) & (g1294) & (g1300) & (!g1305) & (g1344)) + ((g1030) & (!g1294) & (!g1300) & (!g1305) & (!g1344)) + ((g1030) & (!g1294) & (!g1300) & (g1305) & (!g1344)) + ((g1030) & (!g1294) & (!g1300) & (g1305) & (g1344)) + ((g1030) & (g1294) & (!g1300) & (!g1305) & (g1344)) + ((g1030) & (g1294) & (g1300) & (!g1305) & (!g1344)) + ((g1030) & (g1294) & (g1300) & (!g1305) & (g1344)) + ((g1030) & (g1294) & (g1300) & (g1305) & (!g1344)) + ((g1030) & (g1294) & (g1300) & (g1305) & (g1344)));
	assign g1358 = (((!g1160) & (!g1154) & (g1297) & (g1299)) + ((!g1160) & (g1154) & (!g1297) & (g1299)) + ((!g1160) & (g1154) & (g1297) & (!g1299)) + ((!g1160) & (g1154) & (g1297) & (g1299)) + ((g1160) & (!g1154) & (!g1297) & (!g1299)) + ((g1160) & (!g1154) & (!g1297) & (g1299)) + ((g1160) & (!g1154) & (g1297) & (!g1299)) + ((g1160) & (g1154) & (!g1297) & (!g1299)));
	assign g1359 = (((!g1296) & (!g1305) & (!g1344) & (g1358)) + ((!g1296) & (g1305) & (!g1344) & (g1358)) + ((!g1296) & (g1305) & (g1344) & (g1358)) + ((g1296) & (!g1305) & (!g1344) & (!g1358)) + ((g1296) & (!g1305) & (g1344) & (!g1358)) + ((g1296) & (!g1305) & (g1344) & (g1358)) + ((g1296) & (g1305) & (!g1344) & (!g1358)) + ((g1296) & (g1305) & (g1344) & (!g1358)));
	assign g1360 = (((!g1154) & (!g1297) & (g1299) & (!g1305) & (!g1344)) + ((!g1154) & (!g1297) & (g1299) & (g1305) & (!g1344)) + ((!g1154) & (!g1297) & (g1299) & (g1305) & (g1344)) + ((!g1154) & (g1297) & (!g1299) & (!g1305) & (!g1344)) + ((!g1154) & (g1297) & (!g1299) & (!g1305) & (g1344)) + ((!g1154) & (g1297) & (!g1299) & (g1305) & (!g1344)) + ((!g1154) & (g1297) & (!g1299) & (g1305) & (g1344)) + ((!g1154) & (g1297) & (g1299) & (!g1305) & (g1344)) + ((g1154) & (!g1297) & (!g1299) & (!g1305) & (!g1344)) + ((g1154) & (!g1297) & (!g1299) & (g1305) & (!g1344)) + ((g1154) & (!g1297) & (!g1299) & (g1305) & (g1344)) + ((g1154) & (g1297) & (!g1299) & (!g1305) & (g1344)) + ((g1154) & (g1297) & (g1299) & (!g1305) & (!g1344)) + ((g1154) & (g1297) & (g1299) & (!g1305) & (g1344)) + ((g1154) & (g1297) & (g1299) & (g1305) & (!g1344)) + ((g1154) & (g1297) & (g1299) & (g1305) & (g1344)));
	assign g1361 = (((!g1295) & (!ax52x) & (!g1285) & (g1298)) + ((!g1295) & (!ax52x) & (g1285) & (g1298)) + ((!g1295) & (ax52x) & (!g1285) & (!g1298)) + ((!g1295) & (ax52x) & (!g1285) & (g1298)) + ((g1295) & (!ax52x) & (!g1285) & (!g1298)) + ((g1295) & (!ax52x) & (g1285) & (!g1298)) + ((g1295) & (ax52x) & (g1285) & (!g1298)) + ((g1295) & (ax52x) & (g1285) & (g1298)));
	assign g1362 = (((!ax52x) & (!ax53x) & (!g1285) & (!g1305) & (!g1344) & (g1361)) + ((!ax52x) & (!ax53x) & (!g1285) & (!g1305) & (g1344) & (!g1361)) + ((!ax52x) & (!ax53x) & (!g1285) & (!g1305) & (g1344) & (g1361)) + ((!ax52x) & (!ax53x) & (!g1285) & (g1305) & (!g1344) & (g1361)) + ((!ax52x) & (!ax53x) & (!g1285) & (g1305) & (g1344) & (g1361)) + ((!ax52x) & (!ax53x) & (g1285) & (!g1305) & (!g1344) & (!g1361)) + ((!ax52x) & (!ax53x) & (g1285) & (g1305) & (!g1344) & (!g1361)) + ((!ax52x) & (!ax53x) & (g1285) & (g1305) & (g1344) & (!g1361)) + ((!ax52x) & (ax53x) & (!g1285) & (!g1305) & (!g1344) & (!g1361)) + ((!ax52x) & (ax53x) & (!g1285) & (g1305) & (!g1344) & (!g1361)) + ((!ax52x) & (ax53x) & (!g1285) & (g1305) & (g1344) & (!g1361)) + ((!ax52x) & (ax53x) & (g1285) & (!g1305) & (!g1344) & (g1361)) + ((!ax52x) & (ax53x) & (g1285) & (!g1305) & (g1344) & (!g1361)) + ((!ax52x) & (ax53x) & (g1285) & (!g1305) & (g1344) & (g1361)) + ((!ax52x) & (ax53x) & (g1285) & (g1305) & (!g1344) & (g1361)) + ((!ax52x) & (ax53x) & (g1285) & (g1305) & (g1344) & (g1361)) + ((ax52x) & (!ax53x) & (!g1285) & (!g1305) & (!g1344) & (!g1361)) + ((ax52x) & (!ax53x) & (!g1285) & (g1305) & (!g1344) & (!g1361)) + ((ax52x) & (!ax53x) & (!g1285) & (g1305) & (g1344) & (!g1361)) + ((ax52x) & (!ax53x) & (g1285) & (!g1305) & (!g1344) & (!g1361)) + ((ax52x) & (!ax53x) & (g1285) & (g1305) & (!g1344) & (!g1361)) + ((ax52x) & (!ax53x) & (g1285) & (g1305) & (g1344) & (!g1361)) + ((ax52x) & (ax53x) & (!g1285) & (!g1305) & (!g1344) & (g1361)) + ((ax52x) & (ax53x) & (!g1285) & (!g1305) & (g1344) & (!g1361)) + ((ax52x) & (ax53x) & (!g1285) & (!g1305) & (g1344) & (g1361)) + ((ax52x) & (ax53x) & (!g1285) & (g1305) & (!g1344) & (g1361)) + ((ax52x) & (ax53x) & (!g1285) & (g1305) & (g1344) & (g1361)) + ((ax52x) & (ax53x) & (g1285) & (!g1305) & (!g1344) & (g1361)) + ((ax52x) & (ax53x) & (g1285) & (!g1305) & (g1344) & (!g1361)) + ((ax52x) & (ax53x) & (g1285) & (!g1305) & (g1344) & (g1361)) + ((ax52x) & (ax53x) & (g1285) & (g1305) & (!g1344) & (g1361)) + ((ax52x) & (ax53x) & (g1285) & (g1305) & (g1344) & (g1361)));
	assign g1363 = (((!ax52x) & (!g1285) & (!g1298) & (!g1305) & (g1344)) + ((!ax52x) & (!g1285) & (g1298) & (!g1305) & (!g1344)) + ((!ax52x) & (!g1285) & (g1298) & (!g1305) & (g1344)) + ((!ax52x) & (!g1285) & (g1298) & (g1305) & (!g1344)) + ((!ax52x) & (!g1285) & (g1298) & (g1305) & (g1344)) + ((!ax52x) & (g1285) & (g1298) & (!g1305) & (!g1344)) + ((!ax52x) & (g1285) & (g1298) & (g1305) & (!g1344)) + ((!ax52x) & (g1285) & (g1298) & (g1305) & (g1344)) + ((ax52x) & (!g1285) & (!g1298) & (!g1305) & (!g1344)) + ((ax52x) & (!g1285) & (!g1298) & (g1305) & (!g1344)) + ((ax52x) & (!g1285) & (!g1298) & (g1305) & (g1344)) + ((ax52x) & (g1285) & (!g1298) & (!g1305) & (!g1344)) + ((ax52x) & (g1285) & (!g1298) & (!g1305) & (g1344)) + ((ax52x) & (g1285) & (!g1298) & (g1305) & (!g1344)) + ((ax52x) & (g1285) & (!g1298) & (g1305) & (g1344)) + ((ax52x) & (g1285) & (g1298) & (!g1305) & (g1344)));
	assign g1364 = (((!ax48x) & (!ax49x)));
	assign g1365 = (((!g1285) & (!ax50x) & (!ax51x) & (!g1305) & (!g1344) & (!g1364)) + ((!g1285) & (!ax50x) & (!ax51x) & (g1305) & (!g1344) & (!g1364)) + ((!g1285) & (!ax50x) & (!ax51x) & (g1305) & (g1344) & (!g1364)) + ((!g1285) & (!ax50x) & (ax51x) & (!g1305) & (g1344) & (!g1364)) + ((!g1285) & (ax50x) & (ax51x) & (!g1305) & (g1344) & (!g1364)) + ((!g1285) & (ax50x) & (ax51x) & (!g1305) & (g1344) & (g1364)) + ((g1285) & (!ax50x) & (!ax51x) & (!g1305) & (!g1344) & (!g1364)) + ((g1285) & (!ax50x) & (!ax51x) & (!g1305) & (!g1344) & (g1364)) + ((g1285) & (!ax50x) & (!ax51x) & (!g1305) & (g1344) & (!g1364)) + ((g1285) & (!ax50x) & (!ax51x) & (g1305) & (!g1344) & (!g1364)) + ((g1285) & (!ax50x) & (!ax51x) & (g1305) & (!g1344) & (g1364)) + ((g1285) & (!ax50x) & (!ax51x) & (g1305) & (g1344) & (!g1364)) + ((g1285) & (!ax50x) & (!ax51x) & (g1305) & (g1344) & (g1364)) + ((g1285) & (!ax50x) & (ax51x) & (!g1305) & (!g1344) & (!g1364)) + ((g1285) & (!ax50x) & (ax51x) & (!g1305) & (g1344) & (!g1364)) + ((g1285) & (!ax50x) & (ax51x) & (!g1305) & (g1344) & (g1364)) + ((g1285) & (!ax50x) & (ax51x) & (g1305) & (!g1344) & (!g1364)) + ((g1285) & (!ax50x) & (ax51x) & (g1305) & (g1344) & (!g1364)) + ((g1285) & (ax50x) & (!ax51x) & (!g1305) & (g1344) & (!g1364)) + ((g1285) & (ax50x) & (!ax51x) & (!g1305) & (g1344) & (g1364)) + ((g1285) & (ax50x) & (ax51x) & (!g1305) & (!g1344) & (!g1364)) + ((g1285) & (ax50x) & (ax51x) & (!g1305) & (!g1344) & (g1364)) + ((g1285) & (ax50x) & (ax51x) & (!g1305) & (g1344) & (!g1364)) + ((g1285) & (ax50x) & (ax51x) & (!g1305) & (g1344) & (g1364)) + ((g1285) & (ax50x) & (ax51x) & (g1305) & (!g1344) & (!g1364)) + ((g1285) & (ax50x) & (ax51x) & (g1305) & (!g1344) & (g1364)) + ((g1285) & (ax50x) & (ax51x) & (g1305) & (g1344) & (!g1364)) + ((g1285) & (ax50x) & (ax51x) & (g1305) & (g1344) & (g1364)));
	assign g1366 = (((!g1154) & (!g1295) & (g1362) & (g1363) & (g1365)) + ((!g1154) & (g1295) & (g1362) & (!g1363) & (g1365)) + ((!g1154) & (g1295) & (g1362) & (g1363) & (!g1365)) + ((!g1154) & (g1295) & (g1362) & (g1363) & (g1365)) + ((g1154) & (!g1295) & (!g1362) & (g1363) & (g1365)) + ((g1154) & (!g1295) & (g1362) & (!g1363) & (!g1365)) + ((g1154) & (!g1295) & (g1362) & (!g1363) & (g1365)) + ((g1154) & (!g1295) & (g1362) & (g1363) & (!g1365)) + ((g1154) & (!g1295) & (g1362) & (g1363) & (g1365)) + ((g1154) & (g1295) & (!g1362) & (!g1363) & (g1365)) + ((g1154) & (g1295) & (!g1362) & (g1363) & (!g1365)) + ((g1154) & (g1295) & (!g1362) & (g1363) & (g1365)) + ((g1154) & (g1295) & (g1362) & (!g1363) & (!g1365)) + ((g1154) & (g1295) & (g1362) & (!g1363) & (g1365)) + ((g1154) & (g1295) & (g1362) & (g1363) & (!g1365)) + ((g1154) & (g1295) & (g1362) & (g1363) & (g1365)));
	assign g1367 = (((!g1030) & (!g1160) & (g1359) & (g1360) & (g1366)) + ((!g1030) & (g1160) & (g1359) & (!g1360) & (g1366)) + ((!g1030) & (g1160) & (g1359) & (g1360) & (!g1366)) + ((!g1030) & (g1160) & (g1359) & (g1360) & (g1366)) + ((g1030) & (!g1160) & (!g1359) & (g1360) & (g1366)) + ((g1030) & (!g1160) & (g1359) & (!g1360) & (!g1366)) + ((g1030) & (!g1160) & (g1359) & (!g1360) & (g1366)) + ((g1030) & (!g1160) & (g1359) & (g1360) & (!g1366)) + ((g1030) & (!g1160) & (g1359) & (g1360) & (g1366)) + ((g1030) & (g1160) & (!g1359) & (!g1360) & (g1366)) + ((g1030) & (g1160) & (!g1359) & (g1360) & (!g1366)) + ((g1030) & (g1160) & (!g1359) & (g1360) & (g1366)) + ((g1030) & (g1160) & (g1359) & (!g1360) & (!g1366)) + ((g1030) & (g1160) & (g1359) & (!g1360) & (g1366)) + ((g1030) & (g1160) & (g1359) & (g1360) & (!g1366)) + ((g1030) & (g1160) & (g1359) & (g1360) & (g1366)));
	assign g1368 = (((!g914) & (!g1032) & (g1356) & (g1357) & (g1367)) + ((!g914) & (g1032) & (g1356) & (!g1357) & (g1367)) + ((!g914) & (g1032) & (g1356) & (g1357) & (!g1367)) + ((!g914) & (g1032) & (g1356) & (g1357) & (g1367)) + ((g914) & (!g1032) & (!g1356) & (g1357) & (g1367)) + ((g914) & (!g1032) & (g1356) & (!g1357) & (!g1367)) + ((g914) & (!g1032) & (g1356) & (!g1357) & (g1367)) + ((g914) & (!g1032) & (g1356) & (g1357) & (!g1367)) + ((g914) & (!g1032) & (g1356) & (g1357) & (g1367)) + ((g914) & (g1032) & (!g1356) & (!g1357) & (g1367)) + ((g914) & (g1032) & (!g1356) & (g1357) & (!g1367)) + ((g914) & (g1032) & (!g1356) & (g1357) & (g1367)) + ((g914) & (g1032) & (g1356) & (!g1357) & (!g1367)) + ((g914) & (g1032) & (g1356) & (!g1357) & (g1367)) + ((g914) & (g1032) & (g1356) & (g1357) & (!g1367)) + ((g914) & (g1032) & (g1356) & (g1357) & (g1367)));
	assign g1369 = (((!g803) & (!g851) & (g1353) & (g1354) & (g1368)) + ((!g803) & (g851) & (g1353) & (!g1354) & (g1368)) + ((!g803) & (g851) & (g1353) & (g1354) & (!g1368)) + ((!g803) & (g851) & (g1353) & (g1354) & (g1368)) + ((g803) & (!g851) & (!g1353) & (g1354) & (g1368)) + ((g803) & (!g851) & (g1353) & (!g1354) & (!g1368)) + ((g803) & (!g851) & (g1353) & (!g1354) & (g1368)) + ((g803) & (!g851) & (g1353) & (g1354) & (!g1368)) + ((g803) & (!g851) & (g1353) & (g1354) & (g1368)) + ((g803) & (g851) & (!g1353) & (!g1354) & (g1368)) + ((g803) & (g851) & (!g1353) & (g1354) & (!g1368)) + ((g803) & (g851) & (!g1353) & (g1354) & (g1368)) + ((g803) & (g851) & (g1353) & (!g1354) & (!g1368)) + ((g803) & (g851) & (g1353) & (!g1354) & (g1368)) + ((g803) & (g851) & (g1353) & (g1354) & (!g1368)) + ((g803) & (g851) & (g1353) & (g1354) & (g1368)));
	assign g1370 = (((!g700) & (!g744) & (g1350) & (g1351) & (g1369)) + ((!g700) & (g744) & (g1350) & (!g1351) & (g1369)) + ((!g700) & (g744) & (g1350) & (g1351) & (!g1369)) + ((!g700) & (g744) & (g1350) & (g1351) & (g1369)) + ((g700) & (!g744) & (!g1350) & (g1351) & (g1369)) + ((g700) & (!g744) & (g1350) & (!g1351) & (!g1369)) + ((g700) & (!g744) & (g1350) & (!g1351) & (g1369)) + ((g700) & (!g744) & (g1350) & (g1351) & (!g1369)) + ((g700) & (!g744) & (g1350) & (g1351) & (g1369)) + ((g700) & (g744) & (!g1350) & (!g1351) & (g1369)) + ((g700) & (g744) & (!g1350) & (g1351) & (!g1369)) + ((g700) & (g744) & (!g1350) & (g1351) & (g1369)) + ((g700) & (g744) & (g1350) & (!g1351) & (!g1369)) + ((g700) & (g744) & (g1350) & (!g1351) & (g1369)) + ((g700) & (g744) & (g1350) & (g1351) & (!g1369)) + ((g700) & (g744) & (g1350) & (g1351) & (g1369)));
	assign g1371 = (((!g604) & (!g645) & (g1347) & (g1348) & (g1370)) + ((!g604) & (g645) & (g1347) & (!g1348) & (g1370)) + ((!g604) & (g645) & (g1347) & (g1348) & (!g1370)) + ((!g604) & (g645) & (g1347) & (g1348) & (g1370)) + ((g604) & (!g645) & (!g1347) & (g1348) & (g1370)) + ((g604) & (!g645) & (g1347) & (!g1348) & (!g1370)) + ((g604) & (!g645) & (g1347) & (!g1348) & (g1370)) + ((g604) & (!g645) & (g1347) & (g1348) & (!g1370)) + ((g604) & (!g645) & (g1347) & (g1348) & (g1370)) + ((g604) & (g645) & (!g1347) & (!g1348) & (g1370)) + ((g604) & (g645) & (!g1347) & (g1348) & (!g1370)) + ((g604) & (g645) & (!g1347) & (g1348) & (g1370)) + ((g604) & (g645) & (g1347) & (!g1348) & (!g1370)) + ((g604) & (g645) & (g1347) & (!g1348) & (g1370)) + ((g604) & (g645) & (g1347) & (g1348) & (!g1370)) + ((g604) & (g645) & (g1347) & (g1348) & (g1370)));
	assign g1372 = (((!g4) & (!g1341) & (!g1342) & (!g1305) & (!g1344)) + ((!g4) & (!g1341) & (!g1342) & (g1305) & (!g1344)) + ((!g4) & (!g1341) & (!g1342) & (g1305) & (g1344)) + ((!g4) & (!g1341) & (g1342) & (!g1305) & (g1344)) + ((!g4) & (g1341) & (g1342) & (!g1305) & (!g1344)) + ((!g4) & (g1341) & (g1342) & (!g1305) & (g1344)) + ((!g4) & (g1341) & (g1342) & (g1305) & (!g1344)) + ((!g4) & (g1341) & (g1342) & (g1305) & (g1344)) + ((g4) & (!g1341) & (g1342) & (!g1305) & (!g1344)) + ((g4) & (!g1341) & (g1342) & (!g1305) & (g1344)) + ((g4) & (!g1341) & (g1342) & (g1305) & (!g1344)) + ((g4) & (!g1341) & (g1342) & (g1305) & (g1344)) + ((g4) & (g1341) & (!g1342) & (!g1305) & (!g1344)) + ((g4) & (g1341) & (!g1342) & (g1305) & (!g1344)) + ((g4) & (g1341) & (!g1342) & (g1305) & (g1344)) + ((g4) & (g1341) & (g1342) & (!g1305) & (g1344)));
	assign g1373 = (((!g8) & (!g1308) & (g1340) & (!g1305) & (!g1344)) + ((!g8) & (!g1308) & (g1340) & (g1305) & (!g1344)) + ((!g8) & (!g1308) & (g1340) & (g1305) & (g1344)) + ((!g8) & (g1308) & (!g1340) & (!g1305) & (!g1344)) + ((!g8) & (g1308) & (!g1340) & (!g1305) & (g1344)) + ((!g8) & (g1308) & (!g1340) & (g1305) & (!g1344)) + ((!g8) & (g1308) & (!g1340) & (g1305) & (g1344)) + ((!g8) & (g1308) & (g1340) & (!g1305) & (g1344)) + ((g8) & (!g1308) & (!g1340) & (!g1305) & (!g1344)) + ((g8) & (!g1308) & (!g1340) & (g1305) & (!g1344)) + ((g8) & (!g1308) & (!g1340) & (g1305) & (g1344)) + ((g8) & (g1308) & (!g1340) & (!g1305) & (g1344)) + ((g8) & (g1308) & (g1340) & (!g1305) & (!g1344)) + ((g8) & (g1308) & (g1340) & (!g1305) & (g1344)) + ((g8) & (g1308) & (g1340) & (g1305) & (!g1344)) + ((g8) & (g1308) & (g1340) & (g1305) & (g1344)));
	assign g1374 = (((!g18) & (!g27) & (g1310) & (g1339)) + ((!g18) & (g27) & (!g1310) & (g1339)) + ((!g18) & (g27) & (g1310) & (!g1339)) + ((!g18) & (g27) & (g1310) & (g1339)) + ((g18) & (!g27) & (!g1310) & (!g1339)) + ((g18) & (!g27) & (!g1310) & (g1339)) + ((g18) & (!g27) & (g1310) & (!g1339)) + ((g18) & (g27) & (!g1310) & (!g1339)));
	assign g1375 = (((!g1309) & (!g1305) & (!g1344) & (g1374)) + ((!g1309) & (g1305) & (!g1344) & (g1374)) + ((!g1309) & (g1305) & (g1344) & (g1374)) + ((g1309) & (!g1305) & (!g1344) & (!g1374)) + ((g1309) & (!g1305) & (g1344) & (!g1374)) + ((g1309) & (!g1305) & (g1344) & (g1374)) + ((g1309) & (g1305) & (!g1344) & (!g1374)) + ((g1309) & (g1305) & (g1344) & (!g1374)));
	assign g1376 = (((!g27) & (!g1310) & (g1339) & (!g1305) & (!g1344)) + ((!g27) & (!g1310) & (g1339) & (g1305) & (!g1344)) + ((!g27) & (!g1310) & (g1339) & (g1305) & (g1344)) + ((!g27) & (g1310) & (!g1339) & (!g1305) & (!g1344)) + ((!g27) & (g1310) & (!g1339) & (!g1305) & (g1344)) + ((!g27) & (g1310) & (!g1339) & (g1305) & (!g1344)) + ((!g27) & (g1310) & (!g1339) & (g1305) & (g1344)) + ((!g27) & (g1310) & (g1339) & (!g1305) & (g1344)) + ((g27) & (!g1310) & (!g1339) & (!g1305) & (!g1344)) + ((g27) & (!g1310) & (!g1339) & (g1305) & (!g1344)) + ((g27) & (!g1310) & (!g1339) & (g1305) & (g1344)) + ((g27) & (g1310) & (!g1339) & (!g1305) & (g1344)) + ((g27) & (g1310) & (g1339) & (!g1305) & (!g1344)) + ((g27) & (g1310) & (g1339) & (!g1305) & (g1344)) + ((g27) & (g1310) & (g1339) & (g1305) & (!g1344)) + ((g27) & (g1310) & (g1339) & (g1305) & (g1344)));
	assign g1377 = (((!g39) & (!g54) & (g1312) & (g1338)) + ((!g39) & (g54) & (!g1312) & (g1338)) + ((!g39) & (g54) & (g1312) & (!g1338)) + ((!g39) & (g54) & (g1312) & (g1338)) + ((g39) & (!g54) & (!g1312) & (!g1338)) + ((g39) & (!g54) & (!g1312) & (g1338)) + ((g39) & (!g54) & (g1312) & (!g1338)) + ((g39) & (g54) & (!g1312) & (!g1338)));
	assign g1378 = (((!g1311) & (!g1305) & (!g1344) & (g1377)) + ((!g1311) & (g1305) & (!g1344) & (g1377)) + ((!g1311) & (g1305) & (g1344) & (g1377)) + ((g1311) & (!g1305) & (!g1344) & (!g1377)) + ((g1311) & (!g1305) & (g1344) & (!g1377)) + ((g1311) & (!g1305) & (g1344) & (g1377)) + ((g1311) & (g1305) & (!g1344) & (!g1377)) + ((g1311) & (g1305) & (g1344) & (!g1377)));
	assign g1379 = (((!g54) & (!g1312) & (g1338) & (!g1305) & (!g1344)) + ((!g54) & (!g1312) & (g1338) & (g1305) & (!g1344)) + ((!g54) & (!g1312) & (g1338) & (g1305) & (g1344)) + ((!g54) & (g1312) & (!g1338) & (!g1305) & (!g1344)) + ((!g54) & (g1312) & (!g1338) & (!g1305) & (g1344)) + ((!g54) & (g1312) & (!g1338) & (g1305) & (!g1344)) + ((!g54) & (g1312) & (!g1338) & (g1305) & (g1344)) + ((!g54) & (g1312) & (g1338) & (!g1305) & (g1344)) + ((g54) & (!g1312) & (!g1338) & (!g1305) & (!g1344)) + ((g54) & (!g1312) & (!g1338) & (g1305) & (!g1344)) + ((g54) & (!g1312) & (!g1338) & (g1305) & (g1344)) + ((g54) & (g1312) & (!g1338) & (!g1305) & (g1344)) + ((g54) & (g1312) & (g1338) & (!g1305) & (!g1344)) + ((g54) & (g1312) & (g1338) & (!g1305) & (g1344)) + ((g54) & (g1312) & (g1338) & (g1305) & (!g1344)) + ((g54) & (g1312) & (g1338) & (g1305) & (g1344)));
	assign g1380 = (((!g68) & (!g87) & (g1314) & (g1337)) + ((!g68) & (g87) & (!g1314) & (g1337)) + ((!g68) & (g87) & (g1314) & (!g1337)) + ((!g68) & (g87) & (g1314) & (g1337)) + ((g68) & (!g87) & (!g1314) & (!g1337)) + ((g68) & (!g87) & (!g1314) & (g1337)) + ((g68) & (!g87) & (g1314) & (!g1337)) + ((g68) & (g87) & (!g1314) & (!g1337)));
	assign g1381 = (((!g1313) & (!g1305) & (!g1344) & (g1380)) + ((!g1313) & (g1305) & (!g1344) & (g1380)) + ((!g1313) & (g1305) & (g1344) & (g1380)) + ((g1313) & (!g1305) & (!g1344) & (!g1380)) + ((g1313) & (!g1305) & (g1344) & (!g1380)) + ((g1313) & (!g1305) & (g1344) & (g1380)) + ((g1313) & (g1305) & (!g1344) & (!g1380)) + ((g1313) & (g1305) & (g1344) & (!g1380)));
	assign g1382 = (((!g87) & (!g1314) & (g1337) & (!g1305) & (!g1344)) + ((!g87) & (!g1314) & (g1337) & (g1305) & (!g1344)) + ((!g87) & (!g1314) & (g1337) & (g1305) & (g1344)) + ((!g87) & (g1314) & (!g1337) & (!g1305) & (!g1344)) + ((!g87) & (g1314) & (!g1337) & (!g1305) & (g1344)) + ((!g87) & (g1314) & (!g1337) & (g1305) & (!g1344)) + ((!g87) & (g1314) & (!g1337) & (g1305) & (g1344)) + ((!g87) & (g1314) & (g1337) & (!g1305) & (g1344)) + ((g87) & (!g1314) & (!g1337) & (!g1305) & (!g1344)) + ((g87) & (!g1314) & (!g1337) & (g1305) & (!g1344)) + ((g87) & (!g1314) & (!g1337) & (g1305) & (g1344)) + ((g87) & (g1314) & (!g1337) & (!g1305) & (g1344)) + ((g87) & (g1314) & (g1337) & (!g1305) & (!g1344)) + ((g87) & (g1314) & (g1337) & (!g1305) & (g1344)) + ((g87) & (g1314) & (g1337) & (g1305) & (!g1344)) + ((g87) & (g1314) & (g1337) & (g1305) & (g1344)));
	assign g1383 = (((!g104) & (!g127) & (g1316) & (g1336)) + ((!g104) & (g127) & (!g1316) & (g1336)) + ((!g104) & (g127) & (g1316) & (!g1336)) + ((!g104) & (g127) & (g1316) & (g1336)) + ((g104) & (!g127) & (!g1316) & (!g1336)) + ((g104) & (!g127) & (!g1316) & (g1336)) + ((g104) & (!g127) & (g1316) & (!g1336)) + ((g104) & (g127) & (!g1316) & (!g1336)));
	assign g1384 = (((!g1315) & (!g1305) & (!g1344) & (g1383)) + ((!g1315) & (g1305) & (!g1344) & (g1383)) + ((!g1315) & (g1305) & (g1344) & (g1383)) + ((g1315) & (!g1305) & (!g1344) & (!g1383)) + ((g1315) & (!g1305) & (g1344) & (!g1383)) + ((g1315) & (!g1305) & (g1344) & (g1383)) + ((g1315) & (g1305) & (!g1344) & (!g1383)) + ((g1315) & (g1305) & (g1344) & (!g1383)));
	assign g1385 = (((!g127) & (!g1316) & (g1336) & (!g1305) & (!g1344)) + ((!g127) & (!g1316) & (g1336) & (g1305) & (!g1344)) + ((!g127) & (!g1316) & (g1336) & (g1305) & (g1344)) + ((!g127) & (g1316) & (!g1336) & (!g1305) & (!g1344)) + ((!g127) & (g1316) & (!g1336) & (!g1305) & (g1344)) + ((!g127) & (g1316) & (!g1336) & (g1305) & (!g1344)) + ((!g127) & (g1316) & (!g1336) & (g1305) & (g1344)) + ((!g127) & (g1316) & (g1336) & (!g1305) & (g1344)) + ((g127) & (!g1316) & (!g1336) & (!g1305) & (!g1344)) + ((g127) & (!g1316) & (!g1336) & (g1305) & (!g1344)) + ((g127) & (!g1316) & (!g1336) & (g1305) & (g1344)) + ((g127) & (g1316) & (!g1336) & (!g1305) & (g1344)) + ((g127) & (g1316) & (g1336) & (!g1305) & (!g1344)) + ((g127) & (g1316) & (g1336) & (!g1305) & (g1344)) + ((g127) & (g1316) & (g1336) & (g1305) & (!g1344)) + ((g127) & (g1316) & (g1336) & (g1305) & (g1344)));
	assign g1386 = (((!g147) & (!g174) & (g1318) & (g1335)) + ((!g147) & (g174) & (!g1318) & (g1335)) + ((!g147) & (g174) & (g1318) & (!g1335)) + ((!g147) & (g174) & (g1318) & (g1335)) + ((g147) & (!g174) & (!g1318) & (!g1335)) + ((g147) & (!g174) & (!g1318) & (g1335)) + ((g147) & (!g174) & (g1318) & (!g1335)) + ((g147) & (g174) & (!g1318) & (!g1335)));
	assign g1387 = (((!g1317) & (!g1305) & (!g1344) & (g1386)) + ((!g1317) & (g1305) & (!g1344) & (g1386)) + ((!g1317) & (g1305) & (g1344) & (g1386)) + ((g1317) & (!g1305) & (!g1344) & (!g1386)) + ((g1317) & (!g1305) & (g1344) & (!g1386)) + ((g1317) & (!g1305) & (g1344) & (g1386)) + ((g1317) & (g1305) & (!g1344) & (!g1386)) + ((g1317) & (g1305) & (g1344) & (!g1386)));
	assign g1388 = (((!g174) & (!g1318) & (g1335) & (!g1305) & (!g1344)) + ((!g174) & (!g1318) & (g1335) & (g1305) & (!g1344)) + ((!g174) & (!g1318) & (g1335) & (g1305) & (g1344)) + ((!g174) & (g1318) & (!g1335) & (!g1305) & (!g1344)) + ((!g174) & (g1318) & (!g1335) & (!g1305) & (g1344)) + ((!g174) & (g1318) & (!g1335) & (g1305) & (!g1344)) + ((!g174) & (g1318) & (!g1335) & (g1305) & (g1344)) + ((!g174) & (g1318) & (g1335) & (!g1305) & (g1344)) + ((g174) & (!g1318) & (!g1335) & (!g1305) & (!g1344)) + ((g174) & (!g1318) & (!g1335) & (g1305) & (!g1344)) + ((g174) & (!g1318) & (!g1335) & (g1305) & (g1344)) + ((g174) & (g1318) & (!g1335) & (!g1305) & (g1344)) + ((g174) & (g1318) & (g1335) & (!g1305) & (!g1344)) + ((g174) & (g1318) & (g1335) & (!g1305) & (g1344)) + ((g174) & (g1318) & (g1335) & (g1305) & (!g1344)) + ((g174) & (g1318) & (g1335) & (g1305) & (g1344)));
	assign g1389 = (((!g198) & (!g229) & (g1320) & (g1334)) + ((!g198) & (g229) & (!g1320) & (g1334)) + ((!g198) & (g229) & (g1320) & (!g1334)) + ((!g198) & (g229) & (g1320) & (g1334)) + ((g198) & (!g229) & (!g1320) & (!g1334)) + ((g198) & (!g229) & (!g1320) & (g1334)) + ((g198) & (!g229) & (g1320) & (!g1334)) + ((g198) & (g229) & (!g1320) & (!g1334)));
	assign g1390 = (((!g1319) & (!g1305) & (!g1344) & (g1389)) + ((!g1319) & (g1305) & (!g1344) & (g1389)) + ((!g1319) & (g1305) & (g1344) & (g1389)) + ((g1319) & (!g1305) & (!g1344) & (!g1389)) + ((g1319) & (!g1305) & (g1344) & (!g1389)) + ((g1319) & (!g1305) & (g1344) & (g1389)) + ((g1319) & (g1305) & (!g1344) & (!g1389)) + ((g1319) & (g1305) & (g1344) & (!g1389)));
	assign g1391 = (((!g229) & (!g1320) & (g1334) & (!g1305) & (!g1344)) + ((!g229) & (!g1320) & (g1334) & (g1305) & (!g1344)) + ((!g229) & (!g1320) & (g1334) & (g1305) & (g1344)) + ((!g229) & (g1320) & (!g1334) & (!g1305) & (!g1344)) + ((!g229) & (g1320) & (!g1334) & (!g1305) & (g1344)) + ((!g229) & (g1320) & (!g1334) & (g1305) & (!g1344)) + ((!g229) & (g1320) & (!g1334) & (g1305) & (g1344)) + ((!g229) & (g1320) & (g1334) & (!g1305) & (g1344)) + ((g229) & (!g1320) & (!g1334) & (!g1305) & (!g1344)) + ((g229) & (!g1320) & (!g1334) & (g1305) & (!g1344)) + ((g229) & (!g1320) & (!g1334) & (g1305) & (g1344)) + ((g229) & (g1320) & (!g1334) & (!g1305) & (g1344)) + ((g229) & (g1320) & (g1334) & (!g1305) & (!g1344)) + ((g229) & (g1320) & (g1334) & (!g1305) & (g1344)) + ((g229) & (g1320) & (g1334) & (g1305) & (!g1344)) + ((g229) & (g1320) & (g1334) & (g1305) & (g1344)));
	assign g1392 = (((!g255) & (!g290) & (g1322) & (g1333)) + ((!g255) & (g290) & (!g1322) & (g1333)) + ((!g255) & (g290) & (g1322) & (!g1333)) + ((!g255) & (g290) & (g1322) & (g1333)) + ((g255) & (!g290) & (!g1322) & (!g1333)) + ((g255) & (!g290) & (!g1322) & (g1333)) + ((g255) & (!g290) & (g1322) & (!g1333)) + ((g255) & (g290) & (!g1322) & (!g1333)));
	assign g1393 = (((!g1321) & (!g1305) & (!g1344) & (g1392)) + ((!g1321) & (g1305) & (!g1344) & (g1392)) + ((!g1321) & (g1305) & (g1344) & (g1392)) + ((g1321) & (!g1305) & (!g1344) & (!g1392)) + ((g1321) & (!g1305) & (g1344) & (!g1392)) + ((g1321) & (!g1305) & (g1344) & (g1392)) + ((g1321) & (g1305) & (!g1344) & (!g1392)) + ((g1321) & (g1305) & (g1344) & (!g1392)));
	assign g1394 = (((!g290) & (!g1322) & (g1333) & (!g1305) & (!g1344)) + ((!g290) & (!g1322) & (g1333) & (g1305) & (!g1344)) + ((!g290) & (!g1322) & (g1333) & (g1305) & (g1344)) + ((!g290) & (g1322) & (!g1333) & (!g1305) & (!g1344)) + ((!g290) & (g1322) & (!g1333) & (!g1305) & (g1344)) + ((!g290) & (g1322) & (!g1333) & (g1305) & (!g1344)) + ((!g290) & (g1322) & (!g1333) & (g1305) & (g1344)) + ((!g290) & (g1322) & (g1333) & (!g1305) & (g1344)) + ((g290) & (!g1322) & (!g1333) & (!g1305) & (!g1344)) + ((g290) & (!g1322) & (!g1333) & (g1305) & (!g1344)) + ((g290) & (!g1322) & (!g1333) & (g1305) & (g1344)) + ((g290) & (g1322) & (!g1333) & (!g1305) & (g1344)) + ((g290) & (g1322) & (g1333) & (!g1305) & (!g1344)) + ((g290) & (g1322) & (g1333) & (!g1305) & (g1344)) + ((g290) & (g1322) & (g1333) & (g1305) & (!g1344)) + ((g290) & (g1322) & (g1333) & (g1305) & (g1344)));
	assign g1395 = (((!g319) & (!g358) & (g1324) & (g1332)) + ((!g319) & (g358) & (!g1324) & (g1332)) + ((!g319) & (g358) & (g1324) & (!g1332)) + ((!g319) & (g358) & (g1324) & (g1332)) + ((g319) & (!g358) & (!g1324) & (!g1332)) + ((g319) & (!g358) & (!g1324) & (g1332)) + ((g319) & (!g358) & (g1324) & (!g1332)) + ((g319) & (g358) & (!g1324) & (!g1332)));
	assign g1396 = (((!g1323) & (!g1305) & (!g1344) & (g1395)) + ((!g1323) & (g1305) & (!g1344) & (g1395)) + ((!g1323) & (g1305) & (g1344) & (g1395)) + ((g1323) & (!g1305) & (!g1344) & (!g1395)) + ((g1323) & (!g1305) & (g1344) & (!g1395)) + ((g1323) & (!g1305) & (g1344) & (g1395)) + ((g1323) & (g1305) & (!g1344) & (!g1395)) + ((g1323) & (g1305) & (g1344) & (!g1395)));
	assign g1397 = (((!g358) & (!g1324) & (g1332) & (!g1305) & (!g1344)) + ((!g358) & (!g1324) & (g1332) & (g1305) & (!g1344)) + ((!g358) & (!g1324) & (g1332) & (g1305) & (g1344)) + ((!g358) & (g1324) & (!g1332) & (!g1305) & (!g1344)) + ((!g358) & (g1324) & (!g1332) & (!g1305) & (g1344)) + ((!g358) & (g1324) & (!g1332) & (g1305) & (!g1344)) + ((!g358) & (g1324) & (!g1332) & (g1305) & (g1344)) + ((!g358) & (g1324) & (g1332) & (!g1305) & (g1344)) + ((g358) & (!g1324) & (!g1332) & (!g1305) & (!g1344)) + ((g358) & (!g1324) & (!g1332) & (g1305) & (!g1344)) + ((g358) & (!g1324) & (!g1332) & (g1305) & (g1344)) + ((g358) & (g1324) & (!g1332) & (!g1305) & (g1344)) + ((g358) & (g1324) & (g1332) & (!g1305) & (!g1344)) + ((g358) & (g1324) & (g1332) & (!g1305) & (g1344)) + ((g358) & (g1324) & (g1332) & (g1305) & (!g1344)) + ((g358) & (g1324) & (g1332) & (g1305) & (g1344)));
	assign g1398 = (((!g390) & (!g433) & (g1326) & (g1331)) + ((!g390) & (g433) & (!g1326) & (g1331)) + ((!g390) & (g433) & (g1326) & (!g1331)) + ((!g390) & (g433) & (g1326) & (g1331)) + ((g390) & (!g433) & (!g1326) & (!g1331)) + ((g390) & (!g433) & (!g1326) & (g1331)) + ((g390) & (!g433) & (g1326) & (!g1331)) + ((g390) & (g433) & (!g1326) & (!g1331)));
	assign g1399 = (((!g1325) & (!g1305) & (!g1344) & (g1398)) + ((!g1325) & (g1305) & (!g1344) & (g1398)) + ((!g1325) & (g1305) & (g1344) & (g1398)) + ((g1325) & (!g1305) & (!g1344) & (!g1398)) + ((g1325) & (!g1305) & (g1344) & (!g1398)) + ((g1325) & (!g1305) & (g1344) & (g1398)) + ((g1325) & (g1305) & (!g1344) & (!g1398)) + ((g1325) & (g1305) & (g1344) & (!g1398)));
	assign g1400 = (((!g433) & (!g1326) & (g1331) & (!g1305) & (!g1344)) + ((!g433) & (!g1326) & (g1331) & (g1305) & (!g1344)) + ((!g433) & (!g1326) & (g1331) & (g1305) & (g1344)) + ((!g433) & (g1326) & (!g1331) & (!g1305) & (!g1344)) + ((!g433) & (g1326) & (!g1331) & (!g1305) & (g1344)) + ((!g433) & (g1326) & (!g1331) & (g1305) & (!g1344)) + ((!g433) & (g1326) & (!g1331) & (g1305) & (g1344)) + ((!g433) & (g1326) & (g1331) & (!g1305) & (g1344)) + ((g433) & (!g1326) & (!g1331) & (!g1305) & (!g1344)) + ((g433) & (!g1326) & (!g1331) & (g1305) & (!g1344)) + ((g433) & (!g1326) & (!g1331) & (g1305) & (g1344)) + ((g433) & (g1326) & (!g1331) & (!g1305) & (g1344)) + ((g433) & (g1326) & (g1331) & (!g1305) & (!g1344)) + ((g433) & (g1326) & (g1331) & (!g1305) & (g1344)) + ((g433) & (g1326) & (g1331) & (g1305) & (!g1344)) + ((g433) & (g1326) & (g1331) & (g1305) & (g1344)));
	assign g1401 = (((!g468) & (!g515) & (g1328) & (g1330)) + ((!g468) & (g515) & (!g1328) & (g1330)) + ((!g468) & (g515) & (g1328) & (!g1330)) + ((!g468) & (g515) & (g1328) & (g1330)) + ((g468) & (!g515) & (!g1328) & (!g1330)) + ((g468) & (!g515) & (!g1328) & (g1330)) + ((g468) & (!g515) & (g1328) & (!g1330)) + ((g468) & (g515) & (!g1328) & (!g1330)));
	assign g1402 = (((!g1327) & (!g1305) & (!g1344) & (g1401)) + ((!g1327) & (g1305) & (!g1344) & (g1401)) + ((!g1327) & (g1305) & (g1344) & (g1401)) + ((g1327) & (!g1305) & (!g1344) & (!g1401)) + ((g1327) & (!g1305) & (g1344) & (!g1401)) + ((g1327) & (!g1305) & (g1344) & (g1401)) + ((g1327) & (g1305) & (!g1344) & (!g1401)) + ((g1327) & (g1305) & (g1344) & (!g1401)));
	assign g1403 = (((!g515) & (!g1328) & (g1330) & (!g1305) & (!g1344)) + ((!g515) & (!g1328) & (g1330) & (g1305) & (!g1344)) + ((!g515) & (!g1328) & (g1330) & (g1305) & (g1344)) + ((!g515) & (g1328) & (!g1330) & (!g1305) & (!g1344)) + ((!g515) & (g1328) & (!g1330) & (!g1305) & (g1344)) + ((!g515) & (g1328) & (!g1330) & (g1305) & (!g1344)) + ((!g515) & (g1328) & (!g1330) & (g1305) & (g1344)) + ((!g515) & (g1328) & (g1330) & (!g1305) & (g1344)) + ((g515) & (!g1328) & (!g1330) & (!g1305) & (!g1344)) + ((g515) & (!g1328) & (!g1330) & (g1305) & (!g1344)) + ((g515) & (!g1328) & (!g1330) & (g1305) & (g1344)) + ((g515) & (g1328) & (!g1330) & (!g1305) & (g1344)) + ((g515) & (g1328) & (g1330) & (!g1305) & (!g1344)) + ((g515) & (g1328) & (g1330) & (!g1305) & (g1344)) + ((g515) & (g1328) & (g1330) & (g1305) & (!g1344)) + ((g515) & (g1328) & (g1330) & (g1305) & (g1344)));
	assign g1404 = (((!g553) & (!g604) & (g1286) & (g1304)) + ((!g553) & (g604) & (!g1286) & (g1304)) + ((!g553) & (g604) & (g1286) & (!g1304)) + ((!g553) & (g604) & (g1286) & (g1304)) + ((g553) & (!g604) & (!g1286) & (!g1304)) + ((g553) & (!g604) & (!g1286) & (g1304)) + ((g553) & (!g604) & (g1286) & (!g1304)) + ((g553) & (g604) & (!g1286) & (!g1304)));
	assign g1405 = (((!g1329) & (!g1305) & (!g1344) & (g1404)) + ((!g1329) & (g1305) & (!g1344) & (g1404)) + ((!g1329) & (g1305) & (g1344) & (g1404)) + ((g1329) & (!g1305) & (!g1344) & (!g1404)) + ((g1329) & (!g1305) & (g1344) & (!g1404)) + ((g1329) & (!g1305) & (g1344) & (g1404)) + ((g1329) & (g1305) & (!g1344) & (!g1404)) + ((g1329) & (g1305) & (g1344) & (!g1404)));
	assign g1406 = (((!g515) & (!g553) & (g1405) & (g1345) & (g1371)) + ((!g515) & (g553) & (g1405) & (!g1345) & (g1371)) + ((!g515) & (g553) & (g1405) & (g1345) & (!g1371)) + ((!g515) & (g553) & (g1405) & (g1345) & (g1371)) + ((g515) & (!g553) & (!g1405) & (g1345) & (g1371)) + ((g515) & (!g553) & (g1405) & (!g1345) & (!g1371)) + ((g515) & (!g553) & (g1405) & (!g1345) & (g1371)) + ((g515) & (!g553) & (g1405) & (g1345) & (!g1371)) + ((g515) & (!g553) & (g1405) & (g1345) & (g1371)) + ((g515) & (g553) & (!g1405) & (!g1345) & (g1371)) + ((g515) & (g553) & (!g1405) & (g1345) & (!g1371)) + ((g515) & (g553) & (!g1405) & (g1345) & (g1371)) + ((g515) & (g553) & (g1405) & (!g1345) & (!g1371)) + ((g515) & (g553) & (g1405) & (!g1345) & (g1371)) + ((g515) & (g553) & (g1405) & (g1345) & (!g1371)) + ((g515) & (g553) & (g1405) & (g1345) & (g1371)));
	assign g1407 = (((!g433) & (!g468) & (g1402) & (g1403) & (g1406)) + ((!g433) & (g468) & (g1402) & (!g1403) & (g1406)) + ((!g433) & (g468) & (g1402) & (g1403) & (!g1406)) + ((!g433) & (g468) & (g1402) & (g1403) & (g1406)) + ((g433) & (!g468) & (!g1402) & (g1403) & (g1406)) + ((g433) & (!g468) & (g1402) & (!g1403) & (!g1406)) + ((g433) & (!g468) & (g1402) & (!g1403) & (g1406)) + ((g433) & (!g468) & (g1402) & (g1403) & (!g1406)) + ((g433) & (!g468) & (g1402) & (g1403) & (g1406)) + ((g433) & (g468) & (!g1402) & (!g1403) & (g1406)) + ((g433) & (g468) & (!g1402) & (g1403) & (!g1406)) + ((g433) & (g468) & (!g1402) & (g1403) & (g1406)) + ((g433) & (g468) & (g1402) & (!g1403) & (!g1406)) + ((g433) & (g468) & (g1402) & (!g1403) & (g1406)) + ((g433) & (g468) & (g1402) & (g1403) & (!g1406)) + ((g433) & (g468) & (g1402) & (g1403) & (g1406)));
	assign g1408 = (((!g358) & (!g390) & (g1399) & (g1400) & (g1407)) + ((!g358) & (g390) & (g1399) & (!g1400) & (g1407)) + ((!g358) & (g390) & (g1399) & (g1400) & (!g1407)) + ((!g358) & (g390) & (g1399) & (g1400) & (g1407)) + ((g358) & (!g390) & (!g1399) & (g1400) & (g1407)) + ((g358) & (!g390) & (g1399) & (!g1400) & (!g1407)) + ((g358) & (!g390) & (g1399) & (!g1400) & (g1407)) + ((g358) & (!g390) & (g1399) & (g1400) & (!g1407)) + ((g358) & (!g390) & (g1399) & (g1400) & (g1407)) + ((g358) & (g390) & (!g1399) & (!g1400) & (g1407)) + ((g358) & (g390) & (!g1399) & (g1400) & (!g1407)) + ((g358) & (g390) & (!g1399) & (g1400) & (g1407)) + ((g358) & (g390) & (g1399) & (!g1400) & (!g1407)) + ((g358) & (g390) & (g1399) & (!g1400) & (g1407)) + ((g358) & (g390) & (g1399) & (g1400) & (!g1407)) + ((g358) & (g390) & (g1399) & (g1400) & (g1407)));
	assign g1409 = (((!g290) & (!g319) & (g1396) & (g1397) & (g1408)) + ((!g290) & (g319) & (g1396) & (!g1397) & (g1408)) + ((!g290) & (g319) & (g1396) & (g1397) & (!g1408)) + ((!g290) & (g319) & (g1396) & (g1397) & (g1408)) + ((g290) & (!g319) & (!g1396) & (g1397) & (g1408)) + ((g290) & (!g319) & (g1396) & (!g1397) & (!g1408)) + ((g290) & (!g319) & (g1396) & (!g1397) & (g1408)) + ((g290) & (!g319) & (g1396) & (g1397) & (!g1408)) + ((g290) & (!g319) & (g1396) & (g1397) & (g1408)) + ((g290) & (g319) & (!g1396) & (!g1397) & (g1408)) + ((g290) & (g319) & (!g1396) & (g1397) & (!g1408)) + ((g290) & (g319) & (!g1396) & (g1397) & (g1408)) + ((g290) & (g319) & (g1396) & (!g1397) & (!g1408)) + ((g290) & (g319) & (g1396) & (!g1397) & (g1408)) + ((g290) & (g319) & (g1396) & (g1397) & (!g1408)) + ((g290) & (g319) & (g1396) & (g1397) & (g1408)));
	assign g1410 = (((!g229) & (!g255) & (g1393) & (g1394) & (g1409)) + ((!g229) & (g255) & (g1393) & (!g1394) & (g1409)) + ((!g229) & (g255) & (g1393) & (g1394) & (!g1409)) + ((!g229) & (g255) & (g1393) & (g1394) & (g1409)) + ((g229) & (!g255) & (!g1393) & (g1394) & (g1409)) + ((g229) & (!g255) & (g1393) & (!g1394) & (!g1409)) + ((g229) & (!g255) & (g1393) & (!g1394) & (g1409)) + ((g229) & (!g255) & (g1393) & (g1394) & (!g1409)) + ((g229) & (!g255) & (g1393) & (g1394) & (g1409)) + ((g229) & (g255) & (!g1393) & (!g1394) & (g1409)) + ((g229) & (g255) & (!g1393) & (g1394) & (!g1409)) + ((g229) & (g255) & (!g1393) & (g1394) & (g1409)) + ((g229) & (g255) & (g1393) & (!g1394) & (!g1409)) + ((g229) & (g255) & (g1393) & (!g1394) & (g1409)) + ((g229) & (g255) & (g1393) & (g1394) & (!g1409)) + ((g229) & (g255) & (g1393) & (g1394) & (g1409)));
	assign g1411 = (((!g174) & (!g198) & (g1390) & (g1391) & (g1410)) + ((!g174) & (g198) & (g1390) & (!g1391) & (g1410)) + ((!g174) & (g198) & (g1390) & (g1391) & (!g1410)) + ((!g174) & (g198) & (g1390) & (g1391) & (g1410)) + ((g174) & (!g198) & (!g1390) & (g1391) & (g1410)) + ((g174) & (!g198) & (g1390) & (!g1391) & (!g1410)) + ((g174) & (!g198) & (g1390) & (!g1391) & (g1410)) + ((g174) & (!g198) & (g1390) & (g1391) & (!g1410)) + ((g174) & (!g198) & (g1390) & (g1391) & (g1410)) + ((g174) & (g198) & (!g1390) & (!g1391) & (g1410)) + ((g174) & (g198) & (!g1390) & (g1391) & (!g1410)) + ((g174) & (g198) & (!g1390) & (g1391) & (g1410)) + ((g174) & (g198) & (g1390) & (!g1391) & (!g1410)) + ((g174) & (g198) & (g1390) & (!g1391) & (g1410)) + ((g174) & (g198) & (g1390) & (g1391) & (!g1410)) + ((g174) & (g198) & (g1390) & (g1391) & (g1410)));
	assign g1412 = (((!g127) & (!g147) & (g1387) & (g1388) & (g1411)) + ((!g127) & (g147) & (g1387) & (!g1388) & (g1411)) + ((!g127) & (g147) & (g1387) & (g1388) & (!g1411)) + ((!g127) & (g147) & (g1387) & (g1388) & (g1411)) + ((g127) & (!g147) & (!g1387) & (g1388) & (g1411)) + ((g127) & (!g147) & (g1387) & (!g1388) & (!g1411)) + ((g127) & (!g147) & (g1387) & (!g1388) & (g1411)) + ((g127) & (!g147) & (g1387) & (g1388) & (!g1411)) + ((g127) & (!g147) & (g1387) & (g1388) & (g1411)) + ((g127) & (g147) & (!g1387) & (!g1388) & (g1411)) + ((g127) & (g147) & (!g1387) & (g1388) & (!g1411)) + ((g127) & (g147) & (!g1387) & (g1388) & (g1411)) + ((g127) & (g147) & (g1387) & (!g1388) & (!g1411)) + ((g127) & (g147) & (g1387) & (!g1388) & (g1411)) + ((g127) & (g147) & (g1387) & (g1388) & (!g1411)) + ((g127) & (g147) & (g1387) & (g1388) & (g1411)));
	assign g1413 = (((!g87) & (!g104) & (g1384) & (g1385) & (g1412)) + ((!g87) & (g104) & (g1384) & (!g1385) & (g1412)) + ((!g87) & (g104) & (g1384) & (g1385) & (!g1412)) + ((!g87) & (g104) & (g1384) & (g1385) & (g1412)) + ((g87) & (!g104) & (!g1384) & (g1385) & (g1412)) + ((g87) & (!g104) & (g1384) & (!g1385) & (!g1412)) + ((g87) & (!g104) & (g1384) & (!g1385) & (g1412)) + ((g87) & (!g104) & (g1384) & (g1385) & (!g1412)) + ((g87) & (!g104) & (g1384) & (g1385) & (g1412)) + ((g87) & (g104) & (!g1384) & (!g1385) & (g1412)) + ((g87) & (g104) & (!g1384) & (g1385) & (!g1412)) + ((g87) & (g104) & (!g1384) & (g1385) & (g1412)) + ((g87) & (g104) & (g1384) & (!g1385) & (!g1412)) + ((g87) & (g104) & (g1384) & (!g1385) & (g1412)) + ((g87) & (g104) & (g1384) & (g1385) & (!g1412)) + ((g87) & (g104) & (g1384) & (g1385) & (g1412)));
	assign g1414 = (((!g54) & (!g68) & (g1381) & (g1382) & (g1413)) + ((!g54) & (g68) & (g1381) & (!g1382) & (g1413)) + ((!g54) & (g68) & (g1381) & (g1382) & (!g1413)) + ((!g54) & (g68) & (g1381) & (g1382) & (g1413)) + ((g54) & (!g68) & (!g1381) & (g1382) & (g1413)) + ((g54) & (!g68) & (g1381) & (!g1382) & (!g1413)) + ((g54) & (!g68) & (g1381) & (!g1382) & (g1413)) + ((g54) & (!g68) & (g1381) & (g1382) & (!g1413)) + ((g54) & (!g68) & (g1381) & (g1382) & (g1413)) + ((g54) & (g68) & (!g1381) & (!g1382) & (g1413)) + ((g54) & (g68) & (!g1381) & (g1382) & (!g1413)) + ((g54) & (g68) & (!g1381) & (g1382) & (g1413)) + ((g54) & (g68) & (g1381) & (!g1382) & (!g1413)) + ((g54) & (g68) & (g1381) & (!g1382) & (g1413)) + ((g54) & (g68) & (g1381) & (g1382) & (!g1413)) + ((g54) & (g68) & (g1381) & (g1382) & (g1413)));
	assign g1415 = (((!g27) & (!g39) & (g1378) & (g1379) & (g1414)) + ((!g27) & (g39) & (g1378) & (!g1379) & (g1414)) + ((!g27) & (g39) & (g1378) & (g1379) & (!g1414)) + ((!g27) & (g39) & (g1378) & (g1379) & (g1414)) + ((g27) & (!g39) & (!g1378) & (g1379) & (g1414)) + ((g27) & (!g39) & (g1378) & (!g1379) & (!g1414)) + ((g27) & (!g39) & (g1378) & (!g1379) & (g1414)) + ((g27) & (!g39) & (g1378) & (g1379) & (!g1414)) + ((g27) & (!g39) & (g1378) & (g1379) & (g1414)) + ((g27) & (g39) & (!g1378) & (!g1379) & (g1414)) + ((g27) & (g39) & (!g1378) & (g1379) & (!g1414)) + ((g27) & (g39) & (!g1378) & (g1379) & (g1414)) + ((g27) & (g39) & (g1378) & (!g1379) & (!g1414)) + ((g27) & (g39) & (g1378) & (!g1379) & (g1414)) + ((g27) & (g39) & (g1378) & (g1379) & (!g1414)) + ((g27) & (g39) & (g1378) & (g1379) & (g1414)));
	assign g1416 = (((!g8) & (!g18) & (g1375) & (g1376) & (g1415)) + ((!g8) & (g18) & (g1375) & (!g1376) & (g1415)) + ((!g8) & (g18) & (g1375) & (g1376) & (!g1415)) + ((!g8) & (g18) & (g1375) & (g1376) & (g1415)) + ((g8) & (!g18) & (!g1375) & (g1376) & (g1415)) + ((g8) & (!g18) & (g1375) & (!g1376) & (!g1415)) + ((g8) & (!g18) & (g1375) & (!g1376) & (g1415)) + ((g8) & (!g18) & (g1375) & (g1376) & (!g1415)) + ((g8) & (!g18) & (g1375) & (g1376) & (g1415)) + ((g8) & (g18) & (!g1375) & (!g1376) & (g1415)) + ((g8) & (g18) & (!g1375) & (g1376) & (!g1415)) + ((g8) & (g18) & (!g1375) & (g1376) & (g1415)) + ((g8) & (g18) & (g1375) & (!g1376) & (!g1415)) + ((g8) & (g18) & (g1375) & (!g1376) & (g1415)) + ((g8) & (g18) & (g1375) & (g1376) & (!g1415)) + ((g8) & (g18) & (g1375) & (g1376) & (g1415)));
	assign g1417 = (((!g2) & (!g8) & (g1308) & (g1340)) + ((!g2) & (g8) & (!g1308) & (g1340)) + ((!g2) & (g8) & (g1308) & (!g1340)) + ((!g2) & (g8) & (g1308) & (g1340)) + ((g2) & (!g8) & (!g1308) & (!g1340)) + ((g2) & (!g8) & (!g1308) & (g1340)) + ((g2) & (!g8) & (g1308) & (!g1340)) + ((g2) & (g8) & (!g1308) & (!g1340)));
	assign g1418 = (((!g1307) & (!g1305) & (!g1344) & (g1417)) + ((!g1307) & (g1305) & (!g1344) & (g1417)) + ((!g1307) & (g1305) & (g1344) & (g1417)) + ((g1307) & (!g1305) & (!g1344) & (!g1417)) + ((g1307) & (!g1305) & (g1344) & (!g1417)) + ((g1307) & (!g1305) & (g1344) & (g1417)) + ((g1307) & (g1305) & (!g1344) & (!g1417)) + ((g1307) & (g1305) & (g1344) & (!g1417)));
	assign g1419 = (((!g4) & (!g2) & (!g1373) & (!g1416) & (g1418)) + ((!g4) & (!g2) & (!g1373) & (g1416) & (g1418)) + ((!g4) & (!g2) & (g1373) & (!g1416) & (g1418)) + ((!g4) & (!g2) & (g1373) & (g1416) & (!g1418)) + ((!g4) & (!g2) & (g1373) & (g1416) & (g1418)) + ((!g4) & (g2) & (!g1373) & (!g1416) & (g1418)) + ((!g4) & (g2) & (!g1373) & (g1416) & (!g1418)) + ((!g4) & (g2) & (!g1373) & (g1416) & (g1418)) + ((!g4) & (g2) & (g1373) & (!g1416) & (!g1418)) + ((!g4) & (g2) & (g1373) & (!g1416) & (g1418)) + ((!g4) & (g2) & (g1373) & (g1416) & (!g1418)) + ((!g4) & (g2) & (g1373) & (g1416) & (g1418)) + ((g4) & (!g2) & (g1373) & (g1416) & (g1418)) + ((g4) & (g2) & (!g1373) & (g1416) & (g1418)) + ((g4) & (g2) & (g1373) & (!g1416) & (g1418)) + ((g4) & (g2) & (g1373) & (g1416) & (g1418)));
	assign g1420 = (((!g4) & (!g1341) & (g1342)) + ((!g4) & (g1341) & (!g1342)) + ((!g4) & (g1341) & (g1342)) + ((g4) & (g1341) & (g1342)));
	assign g1421 = (((!g1306) & (!g1420) & (!g1305) & (!g1344)) + ((!g1306) & (!g1420) & (g1305) & (!g1344)) + ((!g1306) & (!g1420) & (g1305) & (g1344)) + ((g1306) & (g1420) & (!g1305) & (!g1344)) + ((g1306) & (g1420) & (!g1305) & (g1344)) + ((g1306) & (g1420) & (g1305) & (!g1344)) + ((g1306) & (g1420) & (g1305) & (g1344)));
	assign g1422 = (((!g1) & (g1306) & (!g1420) & (!g1305) & (g1344)) + ((!g1) & (g1306) & (g1420) & (!g1305) & (g1344)) + ((g1) & (!g1306) & (g1420) & (g1305) & (!g1344)) + ((g1) & (!g1306) & (g1420) & (g1305) & (g1344)) + ((g1) & (g1306) & (!g1420) & (!g1305) & (!g1344)) + ((g1) & (g1306) & (!g1420) & (!g1305) & (g1344)) + ((g1) & (g1306) & (!g1420) & (g1305) & (!g1344)) + ((g1) & (g1306) & (!g1420) & (g1305) & (g1344)) + ((g1) & (g1306) & (g1420) & (!g1305) & (g1344)));
	assign g1423 = (((!g1) & (!g1372) & (!g1419) & (!g1421) & (!g1422)) + ((g1) & (!g1372) & (!g1419) & (!g1421) & (!g1422)) + ((g1) & (!g1372) & (!g1419) & (g1421) & (!g1422)) + ((g1) & (!g1372) & (g1419) & (!g1421) & (!g1422)) + ((g1) & (!g1372) & (g1419) & (g1421) & (!g1422)) + ((g1) & (g1372) & (!g1419) & (!g1421) & (!g1422)) + ((g1) & (g1372) & (!g1419) & (g1421) & (!g1422)));
	assign g1424 = (((!g553) & (!g1345) & (g1371) & (!g1423)) + ((!g553) & (g1345) & (!g1371) & (!g1423)) + ((!g553) & (g1345) & (!g1371) & (g1423)) + ((!g553) & (g1345) & (g1371) & (g1423)) + ((g553) & (!g1345) & (!g1371) & (!g1423)) + ((g553) & (g1345) & (!g1371) & (g1423)) + ((g553) & (g1345) & (g1371) & (!g1423)) + ((g553) & (g1345) & (g1371) & (g1423)));
	assign g1425 = (((!g604) & (!g645) & (!g1347) & (g1348) & (g1370) & (!g1423)) + ((!g604) & (!g645) & (g1347) & (!g1348) & (!g1370) & (!g1423)) + ((!g604) & (!g645) & (g1347) & (!g1348) & (!g1370) & (g1423)) + ((!g604) & (!g645) & (g1347) & (!g1348) & (g1370) & (!g1423)) + ((!g604) & (!g645) & (g1347) & (!g1348) & (g1370) & (g1423)) + ((!g604) & (!g645) & (g1347) & (g1348) & (!g1370) & (!g1423)) + ((!g604) & (!g645) & (g1347) & (g1348) & (!g1370) & (g1423)) + ((!g604) & (!g645) & (g1347) & (g1348) & (g1370) & (g1423)) + ((!g604) & (g645) & (!g1347) & (!g1348) & (g1370) & (!g1423)) + ((!g604) & (g645) & (!g1347) & (g1348) & (!g1370) & (!g1423)) + ((!g604) & (g645) & (!g1347) & (g1348) & (g1370) & (!g1423)) + ((!g604) & (g645) & (g1347) & (!g1348) & (!g1370) & (!g1423)) + ((!g604) & (g645) & (g1347) & (!g1348) & (!g1370) & (g1423)) + ((!g604) & (g645) & (g1347) & (!g1348) & (g1370) & (g1423)) + ((!g604) & (g645) & (g1347) & (g1348) & (!g1370) & (g1423)) + ((!g604) & (g645) & (g1347) & (g1348) & (g1370) & (g1423)) + ((g604) & (!g645) & (!g1347) & (!g1348) & (!g1370) & (!g1423)) + ((g604) & (!g645) & (!g1347) & (!g1348) & (g1370) & (!g1423)) + ((g604) & (!g645) & (!g1347) & (g1348) & (!g1370) & (!g1423)) + ((g604) & (!g645) & (g1347) & (!g1348) & (!g1370) & (g1423)) + ((g604) & (!g645) & (g1347) & (!g1348) & (g1370) & (g1423)) + ((g604) & (!g645) & (g1347) & (g1348) & (!g1370) & (g1423)) + ((g604) & (!g645) & (g1347) & (g1348) & (g1370) & (!g1423)) + ((g604) & (!g645) & (g1347) & (g1348) & (g1370) & (g1423)) + ((g604) & (g645) & (!g1347) & (!g1348) & (!g1370) & (!g1423)) + ((g604) & (g645) & (g1347) & (!g1348) & (!g1370) & (g1423)) + ((g604) & (g645) & (g1347) & (!g1348) & (g1370) & (!g1423)) + ((g604) & (g645) & (g1347) & (!g1348) & (g1370) & (g1423)) + ((g604) & (g645) & (g1347) & (g1348) & (!g1370) & (!g1423)) + ((g604) & (g645) & (g1347) & (g1348) & (!g1370) & (g1423)) + ((g604) & (g645) & (g1347) & (g1348) & (g1370) & (!g1423)) + ((g604) & (g645) & (g1347) & (g1348) & (g1370) & (g1423)));
	assign g1426 = (((!g645) & (!g1348) & (g1370) & (!g1423)) + ((!g645) & (g1348) & (!g1370) & (!g1423)) + ((!g645) & (g1348) & (!g1370) & (g1423)) + ((!g645) & (g1348) & (g1370) & (g1423)) + ((g645) & (!g1348) & (!g1370) & (!g1423)) + ((g645) & (g1348) & (!g1370) & (g1423)) + ((g645) & (g1348) & (g1370) & (!g1423)) + ((g645) & (g1348) & (g1370) & (g1423)));
	assign g1427 = (((!g700) & (!g744) & (!g1350) & (g1351) & (g1369) & (!g1423)) + ((!g700) & (!g744) & (g1350) & (!g1351) & (!g1369) & (!g1423)) + ((!g700) & (!g744) & (g1350) & (!g1351) & (!g1369) & (g1423)) + ((!g700) & (!g744) & (g1350) & (!g1351) & (g1369) & (!g1423)) + ((!g700) & (!g744) & (g1350) & (!g1351) & (g1369) & (g1423)) + ((!g700) & (!g744) & (g1350) & (g1351) & (!g1369) & (!g1423)) + ((!g700) & (!g744) & (g1350) & (g1351) & (!g1369) & (g1423)) + ((!g700) & (!g744) & (g1350) & (g1351) & (g1369) & (g1423)) + ((!g700) & (g744) & (!g1350) & (!g1351) & (g1369) & (!g1423)) + ((!g700) & (g744) & (!g1350) & (g1351) & (!g1369) & (!g1423)) + ((!g700) & (g744) & (!g1350) & (g1351) & (g1369) & (!g1423)) + ((!g700) & (g744) & (g1350) & (!g1351) & (!g1369) & (!g1423)) + ((!g700) & (g744) & (g1350) & (!g1351) & (!g1369) & (g1423)) + ((!g700) & (g744) & (g1350) & (!g1351) & (g1369) & (g1423)) + ((!g700) & (g744) & (g1350) & (g1351) & (!g1369) & (g1423)) + ((!g700) & (g744) & (g1350) & (g1351) & (g1369) & (g1423)) + ((g700) & (!g744) & (!g1350) & (!g1351) & (!g1369) & (!g1423)) + ((g700) & (!g744) & (!g1350) & (!g1351) & (g1369) & (!g1423)) + ((g700) & (!g744) & (!g1350) & (g1351) & (!g1369) & (!g1423)) + ((g700) & (!g744) & (g1350) & (!g1351) & (!g1369) & (g1423)) + ((g700) & (!g744) & (g1350) & (!g1351) & (g1369) & (g1423)) + ((g700) & (!g744) & (g1350) & (g1351) & (!g1369) & (g1423)) + ((g700) & (!g744) & (g1350) & (g1351) & (g1369) & (!g1423)) + ((g700) & (!g744) & (g1350) & (g1351) & (g1369) & (g1423)) + ((g700) & (g744) & (!g1350) & (!g1351) & (!g1369) & (!g1423)) + ((g700) & (g744) & (g1350) & (!g1351) & (!g1369) & (g1423)) + ((g700) & (g744) & (g1350) & (!g1351) & (g1369) & (!g1423)) + ((g700) & (g744) & (g1350) & (!g1351) & (g1369) & (g1423)) + ((g700) & (g744) & (g1350) & (g1351) & (!g1369) & (!g1423)) + ((g700) & (g744) & (g1350) & (g1351) & (!g1369) & (g1423)) + ((g700) & (g744) & (g1350) & (g1351) & (g1369) & (!g1423)) + ((g700) & (g744) & (g1350) & (g1351) & (g1369) & (g1423)));
	assign g1428 = (((!g744) & (!g1351) & (g1369) & (!g1423)) + ((!g744) & (g1351) & (!g1369) & (!g1423)) + ((!g744) & (g1351) & (!g1369) & (g1423)) + ((!g744) & (g1351) & (g1369) & (g1423)) + ((g744) & (!g1351) & (!g1369) & (!g1423)) + ((g744) & (g1351) & (!g1369) & (g1423)) + ((g744) & (g1351) & (g1369) & (!g1423)) + ((g744) & (g1351) & (g1369) & (g1423)));
	assign g1429 = (((!g803) & (!g851) & (!g1353) & (g1354) & (g1368) & (!g1423)) + ((!g803) & (!g851) & (g1353) & (!g1354) & (!g1368) & (!g1423)) + ((!g803) & (!g851) & (g1353) & (!g1354) & (!g1368) & (g1423)) + ((!g803) & (!g851) & (g1353) & (!g1354) & (g1368) & (!g1423)) + ((!g803) & (!g851) & (g1353) & (!g1354) & (g1368) & (g1423)) + ((!g803) & (!g851) & (g1353) & (g1354) & (!g1368) & (!g1423)) + ((!g803) & (!g851) & (g1353) & (g1354) & (!g1368) & (g1423)) + ((!g803) & (!g851) & (g1353) & (g1354) & (g1368) & (g1423)) + ((!g803) & (g851) & (!g1353) & (!g1354) & (g1368) & (!g1423)) + ((!g803) & (g851) & (!g1353) & (g1354) & (!g1368) & (!g1423)) + ((!g803) & (g851) & (!g1353) & (g1354) & (g1368) & (!g1423)) + ((!g803) & (g851) & (g1353) & (!g1354) & (!g1368) & (!g1423)) + ((!g803) & (g851) & (g1353) & (!g1354) & (!g1368) & (g1423)) + ((!g803) & (g851) & (g1353) & (!g1354) & (g1368) & (g1423)) + ((!g803) & (g851) & (g1353) & (g1354) & (!g1368) & (g1423)) + ((!g803) & (g851) & (g1353) & (g1354) & (g1368) & (g1423)) + ((g803) & (!g851) & (!g1353) & (!g1354) & (!g1368) & (!g1423)) + ((g803) & (!g851) & (!g1353) & (!g1354) & (g1368) & (!g1423)) + ((g803) & (!g851) & (!g1353) & (g1354) & (!g1368) & (!g1423)) + ((g803) & (!g851) & (g1353) & (!g1354) & (!g1368) & (g1423)) + ((g803) & (!g851) & (g1353) & (!g1354) & (g1368) & (g1423)) + ((g803) & (!g851) & (g1353) & (g1354) & (!g1368) & (g1423)) + ((g803) & (!g851) & (g1353) & (g1354) & (g1368) & (!g1423)) + ((g803) & (!g851) & (g1353) & (g1354) & (g1368) & (g1423)) + ((g803) & (g851) & (!g1353) & (!g1354) & (!g1368) & (!g1423)) + ((g803) & (g851) & (g1353) & (!g1354) & (!g1368) & (g1423)) + ((g803) & (g851) & (g1353) & (!g1354) & (g1368) & (!g1423)) + ((g803) & (g851) & (g1353) & (!g1354) & (g1368) & (g1423)) + ((g803) & (g851) & (g1353) & (g1354) & (!g1368) & (!g1423)) + ((g803) & (g851) & (g1353) & (g1354) & (!g1368) & (g1423)) + ((g803) & (g851) & (g1353) & (g1354) & (g1368) & (!g1423)) + ((g803) & (g851) & (g1353) & (g1354) & (g1368) & (g1423)));
	assign g1430 = (((!g851) & (!g1354) & (g1368) & (!g1423)) + ((!g851) & (g1354) & (!g1368) & (!g1423)) + ((!g851) & (g1354) & (!g1368) & (g1423)) + ((!g851) & (g1354) & (g1368) & (g1423)) + ((g851) & (!g1354) & (!g1368) & (!g1423)) + ((g851) & (g1354) & (!g1368) & (g1423)) + ((g851) & (g1354) & (g1368) & (!g1423)) + ((g851) & (g1354) & (g1368) & (g1423)));
	assign g1431 = (((!g914) & (!g1032) & (!g1356) & (g1357) & (g1367) & (!g1423)) + ((!g914) & (!g1032) & (g1356) & (!g1357) & (!g1367) & (!g1423)) + ((!g914) & (!g1032) & (g1356) & (!g1357) & (!g1367) & (g1423)) + ((!g914) & (!g1032) & (g1356) & (!g1357) & (g1367) & (!g1423)) + ((!g914) & (!g1032) & (g1356) & (!g1357) & (g1367) & (g1423)) + ((!g914) & (!g1032) & (g1356) & (g1357) & (!g1367) & (!g1423)) + ((!g914) & (!g1032) & (g1356) & (g1357) & (!g1367) & (g1423)) + ((!g914) & (!g1032) & (g1356) & (g1357) & (g1367) & (g1423)) + ((!g914) & (g1032) & (!g1356) & (!g1357) & (g1367) & (!g1423)) + ((!g914) & (g1032) & (!g1356) & (g1357) & (!g1367) & (!g1423)) + ((!g914) & (g1032) & (!g1356) & (g1357) & (g1367) & (!g1423)) + ((!g914) & (g1032) & (g1356) & (!g1357) & (!g1367) & (!g1423)) + ((!g914) & (g1032) & (g1356) & (!g1357) & (!g1367) & (g1423)) + ((!g914) & (g1032) & (g1356) & (!g1357) & (g1367) & (g1423)) + ((!g914) & (g1032) & (g1356) & (g1357) & (!g1367) & (g1423)) + ((!g914) & (g1032) & (g1356) & (g1357) & (g1367) & (g1423)) + ((g914) & (!g1032) & (!g1356) & (!g1357) & (!g1367) & (!g1423)) + ((g914) & (!g1032) & (!g1356) & (!g1357) & (g1367) & (!g1423)) + ((g914) & (!g1032) & (!g1356) & (g1357) & (!g1367) & (!g1423)) + ((g914) & (!g1032) & (g1356) & (!g1357) & (!g1367) & (g1423)) + ((g914) & (!g1032) & (g1356) & (!g1357) & (g1367) & (g1423)) + ((g914) & (!g1032) & (g1356) & (g1357) & (!g1367) & (g1423)) + ((g914) & (!g1032) & (g1356) & (g1357) & (g1367) & (!g1423)) + ((g914) & (!g1032) & (g1356) & (g1357) & (g1367) & (g1423)) + ((g914) & (g1032) & (!g1356) & (!g1357) & (!g1367) & (!g1423)) + ((g914) & (g1032) & (g1356) & (!g1357) & (!g1367) & (g1423)) + ((g914) & (g1032) & (g1356) & (!g1357) & (g1367) & (!g1423)) + ((g914) & (g1032) & (g1356) & (!g1357) & (g1367) & (g1423)) + ((g914) & (g1032) & (g1356) & (g1357) & (!g1367) & (!g1423)) + ((g914) & (g1032) & (g1356) & (g1357) & (!g1367) & (g1423)) + ((g914) & (g1032) & (g1356) & (g1357) & (g1367) & (!g1423)) + ((g914) & (g1032) & (g1356) & (g1357) & (g1367) & (g1423)));
	assign g1432 = (((!g1032) & (!g1357) & (g1367) & (!g1423)) + ((!g1032) & (g1357) & (!g1367) & (!g1423)) + ((!g1032) & (g1357) & (!g1367) & (g1423)) + ((!g1032) & (g1357) & (g1367) & (g1423)) + ((g1032) & (!g1357) & (!g1367) & (!g1423)) + ((g1032) & (g1357) & (!g1367) & (g1423)) + ((g1032) & (g1357) & (g1367) & (!g1423)) + ((g1032) & (g1357) & (g1367) & (g1423)));
	assign g1433 = (((!g1030) & (!g1160) & (!g1359) & (g1360) & (g1366) & (!g1423)) + ((!g1030) & (!g1160) & (g1359) & (!g1360) & (!g1366) & (!g1423)) + ((!g1030) & (!g1160) & (g1359) & (!g1360) & (!g1366) & (g1423)) + ((!g1030) & (!g1160) & (g1359) & (!g1360) & (g1366) & (!g1423)) + ((!g1030) & (!g1160) & (g1359) & (!g1360) & (g1366) & (g1423)) + ((!g1030) & (!g1160) & (g1359) & (g1360) & (!g1366) & (!g1423)) + ((!g1030) & (!g1160) & (g1359) & (g1360) & (!g1366) & (g1423)) + ((!g1030) & (!g1160) & (g1359) & (g1360) & (g1366) & (g1423)) + ((!g1030) & (g1160) & (!g1359) & (!g1360) & (g1366) & (!g1423)) + ((!g1030) & (g1160) & (!g1359) & (g1360) & (!g1366) & (!g1423)) + ((!g1030) & (g1160) & (!g1359) & (g1360) & (g1366) & (!g1423)) + ((!g1030) & (g1160) & (g1359) & (!g1360) & (!g1366) & (!g1423)) + ((!g1030) & (g1160) & (g1359) & (!g1360) & (!g1366) & (g1423)) + ((!g1030) & (g1160) & (g1359) & (!g1360) & (g1366) & (g1423)) + ((!g1030) & (g1160) & (g1359) & (g1360) & (!g1366) & (g1423)) + ((!g1030) & (g1160) & (g1359) & (g1360) & (g1366) & (g1423)) + ((g1030) & (!g1160) & (!g1359) & (!g1360) & (!g1366) & (!g1423)) + ((g1030) & (!g1160) & (!g1359) & (!g1360) & (g1366) & (!g1423)) + ((g1030) & (!g1160) & (!g1359) & (g1360) & (!g1366) & (!g1423)) + ((g1030) & (!g1160) & (g1359) & (!g1360) & (!g1366) & (g1423)) + ((g1030) & (!g1160) & (g1359) & (!g1360) & (g1366) & (g1423)) + ((g1030) & (!g1160) & (g1359) & (g1360) & (!g1366) & (g1423)) + ((g1030) & (!g1160) & (g1359) & (g1360) & (g1366) & (!g1423)) + ((g1030) & (!g1160) & (g1359) & (g1360) & (g1366) & (g1423)) + ((g1030) & (g1160) & (!g1359) & (!g1360) & (!g1366) & (!g1423)) + ((g1030) & (g1160) & (g1359) & (!g1360) & (!g1366) & (g1423)) + ((g1030) & (g1160) & (g1359) & (!g1360) & (g1366) & (!g1423)) + ((g1030) & (g1160) & (g1359) & (!g1360) & (g1366) & (g1423)) + ((g1030) & (g1160) & (g1359) & (g1360) & (!g1366) & (!g1423)) + ((g1030) & (g1160) & (g1359) & (g1360) & (!g1366) & (g1423)) + ((g1030) & (g1160) & (g1359) & (g1360) & (g1366) & (!g1423)) + ((g1030) & (g1160) & (g1359) & (g1360) & (g1366) & (g1423)));
	assign g1434 = (((!g1160) & (!g1360) & (g1366) & (!g1423)) + ((!g1160) & (g1360) & (!g1366) & (!g1423)) + ((!g1160) & (g1360) & (!g1366) & (g1423)) + ((!g1160) & (g1360) & (g1366) & (g1423)) + ((g1160) & (!g1360) & (!g1366) & (!g1423)) + ((g1160) & (g1360) & (!g1366) & (g1423)) + ((g1160) & (g1360) & (g1366) & (!g1423)) + ((g1160) & (g1360) & (g1366) & (g1423)));
	assign g1435 = (((!g1154) & (!g1295) & (!g1362) & (g1363) & (g1365) & (!g1423)) + ((!g1154) & (!g1295) & (g1362) & (!g1363) & (!g1365) & (!g1423)) + ((!g1154) & (!g1295) & (g1362) & (!g1363) & (!g1365) & (g1423)) + ((!g1154) & (!g1295) & (g1362) & (!g1363) & (g1365) & (!g1423)) + ((!g1154) & (!g1295) & (g1362) & (!g1363) & (g1365) & (g1423)) + ((!g1154) & (!g1295) & (g1362) & (g1363) & (!g1365) & (!g1423)) + ((!g1154) & (!g1295) & (g1362) & (g1363) & (!g1365) & (g1423)) + ((!g1154) & (!g1295) & (g1362) & (g1363) & (g1365) & (g1423)) + ((!g1154) & (g1295) & (!g1362) & (!g1363) & (g1365) & (!g1423)) + ((!g1154) & (g1295) & (!g1362) & (g1363) & (!g1365) & (!g1423)) + ((!g1154) & (g1295) & (!g1362) & (g1363) & (g1365) & (!g1423)) + ((!g1154) & (g1295) & (g1362) & (!g1363) & (!g1365) & (!g1423)) + ((!g1154) & (g1295) & (g1362) & (!g1363) & (!g1365) & (g1423)) + ((!g1154) & (g1295) & (g1362) & (!g1363) & (g1365) & (g1423)) + ((!g1154) & (g1295) & (g1362) & (g1363) & (!g1365) & (g1423)) + ((!g1154) & (g1295) & (g1362) & (g1363) & (g1365) & (g1423)) + ((g1154) & (!g1295) & (!g1362) & (!g1363) & (!g1365) & (!g1423)) + ((g1154) & (!g1295) & (!g1362) & (!g1363) & (g1365) & (!g1423)) + ((g1154) & (!g1295) & (!g1362) & (g1363) & (!g1365) & (!g1423)) + ((g1154) & (!g1295) & (g1362) & (!g1363) & (!g1365) & (g1423)) + ((g1154) & (!g1295) & (g1362) & (!g1363) & (g1365) & (g1423)) + ((g1154) & (!g1295) & (g1362) & (g1363) & (!g1365) & (g1423)) + ((g1154) & (!g1295) & (g1362) & (g1363) & (g1365) & (!g1423)) + ((g1154) & (!g1295) & (g1362) & (g1363) & (g1365) & (g1423)) + ((g1154) & (g1295) & (!g1362) & (!g1363) & (!g1365) & (!g1423)) + ((g1154) & (g1295) & (g1362) & (!g1363) & (!g1365) & (g1423)) + ((g1154) & (g1295) & (g1362) & (!g1363) & (g1365) & (!g1423)) + ((g1154) & (g1295) & (g1362) & (!g1363) & (g1365) & (g1423)) + ((g1154) & (g1295) & (g1362) & (g1363) & (!g1365) & (!g1423)) + ((g1154) & (g1295) & (g1362) & (g1363) & (!g1365) & (g1423)) + ((g1154) & (g1295) & (g1362) & (g1363) & (g1365) & (!g1423)) + ((g1154) & (g1295) & (g1362) & (g1363) & (g1365) & (g1423)));
	assign g1436 = (((!g1295) & (!g1363) & (g1365) & (!g1423)) + ((!g1295) & (g1363) & (!g1365) & (!g1423)) + ((!g1295) & (g1363) & (!g1365) & (g1423)) + ((!g1295) & (g1363) & (g1365) & (g1423)) + ((g1295) & (!g1363) & (!g1365) & (!g1423)) + ((g1295) & (g1363) & (!g1365) & (g1423)) + ((g1295) & (g1363) & (g1365) & (!g1423)) + ((g1295) & (g1363) & (g1365) & (g1423)));
	assign g1437 = (((!g1305) & (g1344)));
	assign g1438 = (((!g1285) & (!ax50x) & (!ax51x) & (!g1437) & (!g1364) & (g1423)) + ((!g1285) & (!ax50x) & (!ax51x) & (!g1437) & (g1364) & (!g1423)) + ((!g1285) & (!ax50x) & (!ax51x) & (!g1437) & (g1364) & (g1423)) + ((!g1285) & (!ax50x) & (!ax51x) & (g1437) & (!g1364) & (!g1423)) + ((!g1285) & (!ax50x) & (ax51x) & (!g1437) & (!g1364) & (!g1423)) + ((!g1285) & (!ax50x) & (ax51x) & (g1437) & (!g1364) & (g1423)) + ((!g1285) & (!ax50x) & (ax51x) & (g1437) & (g1364) & (!g1423)) + ((!g1285) & (!ax50x) & (ax51x) & (g1437) & (g1364) & (g1423)) + ((!g1285) & (ax50x) & (!ax51x) & (g1437) & (!g1364) & (!g1423)) + ((!g1285) & (ax50x) & (!ax51x) & (g1437) & (g1364) & (!g1423)) + ((!g1285) & (ax50x) & (ax51x) & (!g1437) & (!g1364) & (!g1423)) + ((!g1285) & (ax50x) & (ax51x) & (!g1437) & (!g1364) & (g1423)) + ((!g1285) & (ax50x) & (ax51x) & (!g1437) & (g1364) & (!g1423)) + ((!g1285) & (ax50x) & (ax51x) & (!g1437) & (g1364) & (g1423)) + ((!g1285) & (ax50x) & (ax51x) & (g1437) & (!g1364) & (g1423)) + ((!g1285) & (ax50x) & (ax51x) & (g1437) & (g1364) & (g1423)) + ((g1285) & (!ax50x) & (!ax51x) & (!g1437) & (!g1364) & (!g1423)) + ((g1285) & (!ax50x) & (!ax51x) & (!g1437) & (!g1364) & (g1423)) + ((g1285) & (!ax50x) & (!ax51x) & (!g1437) & (g1364) & (g1423)) + ((g1285) & (!ax50x) & (!ax51x) & (g1437) & (g1364) & (!g1423)) + ((g1285) & (!ax50x) & (ax51x) & (!g1437) & (g1364) & (!g1423)) + ((g1285) & (!ax50x) & (ax51x) & (g1437) & (!g1364) & (!g1423)) + ((g1285) & (!ax50x) & (ax51x) & (g1437) & (!g1364) & (g1423)) + ((g1285) & (!ax50x) & (ax51x) & (g1437) & (g1364) & (g1423)) + ((g1285) & (ax50x) & (!ax51x) & (!g1437) & (!g1364) & (!g1423)) + ((g1285) & (ax50x) & (!ax51x) & (!g1437) & (g1364) & (!g1423)) + ((g1285) & (ax50x) & (ax51x) & (!g1437) & (!g1364) & (g1423)) + ((g1285) & (ax50x) & (ax51x) & (!g1437) & (g1364) & (g1423)) + ((g1285) & (ax50x) & (ax51x) & (g1437) & (!g1364) & (!g1423)) + ((g1285) & (ax50x) & (ax51x) & (g1437) & (!g1364) & (g1423)) + ((g1285) & (ax50x) & (ax51x) & (g1437) & (g1364) & (!g1423)) + ((g1285) & (ax50x) & (ax51x) & (g1437) & (g1364) & (g1423)));
	assign g1439 = (((!ax50x) & (!g1437) & (!g1364) & (g1423)) + ((!ax50x) & (!g1437) & (g1364) & (!g1423)) + ((!ax50x) & (!g1437) & (g1364) & (g1423)) + ((!ax50x) & (g1437) & (g1364) & (!g1423)) + ((ax50x) & (!g1437) & (!g1364) & (!g1423)) + ((ax50x) & (g1437) & (!g1364) & (!g1423)) + ((ax50x) & (g1437) & (!g1364) & (g1423)) + ((ax50x) & (g1437) & (g1364) & (g1423)));
	assign g1440 = (((!ax46x) & (!ax47x)));
	assign g1441 = (((!g1437) & (!ax48x) & (!ax49x) & (!g1423) & (!g1440)) + ((!g1437) & (!ax48x) & (ax49x) & (g1423) & (!g1440)) + ((!g1437) & (ax48x) & (ax49x) & (g1423) & (!g1440)) + ((!g1437) & (ax48x) & (ax49x) & (g1423) & (g1440)) + ((g1437) & (!ax48x) & (!ax49x) & (!g1423) & (!g1440)) + ((g1437) & (!ax48x) & (!ax49x) & (!g1423) & (g1440)) + ((g1437) & (!ax48x) & (!ax49x) & (g1423) & (!g1440)) + ((g1437) & (!ax48x) & (ax49x) & (!g1423) & (!g1440)) + ((g1437) & (!ax48x) & (ax49x) & (g1423) & (!g1440)) + ((g1437) & (!ax48x) & (ax49x) & (g1423) & (g1440)) + ((g1437) & (ax48x) & (!ax49x) & (g1423) & (!g1440)) + ((g1437) & (ax48x) & (!ax49x) & (g1423) & (g1440)) + ((g1437) & (ax48x) & (ax49x) & (!g1423) & (!g1440)) + ((g1437) & (ax48x) & (ax49x) & (!g1423) & (g1440)) + ((g1437) & (ax48x) & (ax49x) & (g1423) & (!g1440)) + ((g1437) & (ax48x) & (ax49x) & (g1423) & (g1440)));
	assign g1442 = (((!g1295) & (!g1285) & (g1438) & (g1439) & (g1441)) + ((!g1295) & (g1285) & (g1438) & (!g1439) & (g1441)) + ((!g1295) & (g1285) & (g1438) & (g1439) & (!g1441)) + ((!g1295) & (g1285) & (g1438) & (g1439) & (g1441)) + ((g1295) & (!g1285) & (!g1438) & (g1439) & (g1441)) + ((g1295) & (!g1285) & (g1438) & (!g1439) & (!g1441)) + ((g1295) & (!g1285) & (g1438) & (!g1439) & (g1441)) + ((g1295) & (!g1285) & (g1438) & (g1439) & (!g1441)) + ((g1295) & (!g1285) & (g1438) & (g1439) & (g1441)) + ((g1295) & (g1285) & (!g1438) & (!g1439) & (g1441)) + ((g1295) & (g1285) & (!g1438) & (g1439) & (!g1441)) + ((g1295) & (g1285) & (!g1438) & (g1439) & (g1441)) + ((g1295) & (g1285) & (g1438) & (!g1439) & (!g1441)) + ((g1295) & (g1285) & (g1438) & (!g1439) & (g1441)) + ((g1295) & (g1285) & (g1438) & (g1439) & (!g1441)) + ((g1295) & (g1285) & (g1438) & (g1439) & (g1441)));
	assign g1443 = (((!g1160) & (!g1154) & (g1435) & (g1436) & (g1442)) + ((!g1160) & (g1154) & (g1435) & (!g1436) & (g1442)) + ((!g1160) & (g1154) & (g1435) & (g1436) & (!g1442)) + ((!g1160) & (g1154) & (g1435) & (g1436) & (g1442)) + ((g1160) & (!g1154) & (!g1435) & (g1436) & (g1442)) + ((g1160) & (!g1154) & (g1435) & (!g1436) & (!g1442)) + ((g1160) & (!g1154) & (g1435) & (!g1436) & (g1442)) + ((g1160) & (!g1154) & (g1435) & (g1436) & (!g1442)) + ((g1160) & (!g1154) & (g1435) & (g1436) & (g1442)) + ((g1160) & (g1154) & (!g1435) & (!g1436) & (g1442)) + ((g1160) & (g1154) & (!g1435) & (g1436) & (!g1442)) + ((g1160) & (g1154) & (!g1435) & (g1436) & (g1442)) + ((g1160) & (g1154) & (g1435) & (!g1436) & (!g1442)) + ((g1160) & (g1154) & (g1435) & (!g1436) & (g1442)) + ((g1160) & (g1154) & (g1435) & (g1436) & (!g1442)) + ((g1160) & (g1154) & (g1435) & (g1436) & (g1442)));
	assign g1444 = (((!g1032) & (!g1030) & (g1433) & (g1434) & (g1443)) + ((!g1032) & (g1030) & (g1433) & (!g1434) & (g1443)) + ((!g1032) & (g1030) & (g1433) & (g1434) & (!g1443)) + ((!g1032) & (g1030) & (g1433) & (g1434) & (g1443)) + ((g1032) & (!g1030) & (!g1433) & (g1434) & (g1443)) + ((g1032) & (!g1030) & (g1433) & (!g1434) & (!g1443)) + ((g1032) & (!g1030) & (g1433) & (!g1434) & (g1443)) + ((g1032) & (!g1030) & (g1433) & (g1434) & (!g1443)) + ((g1032) & (!g1030) & (g1433) & (g1434) & (g1443)) + ((g1032) & (g1030) & (!g1433) & (!g1434) & (g1443)) + ((g1032) & (g1030) & (!g1433) & (g1434) & (!g1443)) + ((g1032) & (g1030) & (!g1433) & (g1434) & (g1443)) + ((g1032) & (g1030) & (g1433) & (!g1434) & (!g1443)) + ((g1032) & (g1030) & (g1433) & (!g1434) & (g1443)) + ((g1032) & (g1030) & (g1433) & (g1434) & (!g1443)) + ((g1032) & (g1030) & (g1433) & (g1434) & (g1443)));
	assign g1445 = (((!g851) & (!g914) & (g1431) & (g1432) & (g1444)) + ((!g851) & (g914) & (g1431) & (!g1432) & (g1444)) + ((!g851) & (g914) & (g1431) & (g1432) & (!g1444)) + ((!g851) & (g914) & (g1431) & (g1432) & (g1444)) + ((g851) & (!g914) & (!g1431) & (g1432) & (g1444)) + ((g851) & (!g914) & (g1431) & (!g1432) & (!g1444)) + ((g851) & (!g914) & (g1431) & (!g1432) & (g1444)) + ((g851) & (!g914) & (g1431) & (g1432) & (!g1444)) + ((g851) & (!g914) & (g1431) & (g1432) & (g1444)) + ((g851) & (g914) & (!g1431) & (!g1432) & (g1444)) + ((g851) & (g914) & (!g1431) & (g1432) & (!g1444)) + ((g851) & (g914) & (!g1431) & (g1432) & (g1444)) + ((g851) & (g914) & (g1431) & (!g1432) & (!g1444)) + ((g851) & (g914) & (g1431) & (!g1432) & (g1444)) + ((g851) & (g914) & (g1431) & (g1432) & (!g1444)) + ((g851) & (g914) & (g1431) & (g1432) & (g1444)));
	assign g1446 = (((!g744) & (!g803) & (g1429) & (g1430) & (g1445)) + ((!g744) & (g803) & (g1429) & (!g1430) & (g1445)) + ((!g744) & (g803) & (g1429) & (g1430) & (!g1445)) + ((!g744) & (g803) & (g1429) & (g1430) & (g1445)) + ((g744) & (!g803) & (!g1429) & (g1430) & (g1445)) + ((g744) & (!g803) & (g1429) & (!g1430) & (!g1445)) + ((g744) & (!g803) & (g1429) & (!g1430) & (g1445)) + ((g744) & (!g803) & (g1429) & (g1430) & (!g1445)) + ((g744) & (!g803) & (g1429) & (g1430) & (g1445)) + ((g744) & (g803) & (!g1429) & (!g1430) & (g1445)) + ((g744) & (g803) & (!g1429) & (g1430) & (!g1445)) + ((g744) & (g803) & (!g1429) & (g1430) & (g1445)) + ((g744) & (g803) & (g1429) & (!g1430) & (!g1445)) + ((g744) & (g803) & (g1429) & (!g1430) & (g1445)) + ((g744) & (g803) & (g1429) & (g1430) & (!g1445)) + ((g744) & (g803) & (g1429) & (g1430) & (g1445)));
	assign g1447 = (((!g645) & (!g700) & (g1427) & (g1428) & (g1446)) + ((!g645) & (g700) & (g1427) & (!g1428) & (g1446)) + ((!g645) & (g700) & (g1427) & (g1428) & (!g1446)) + ((!g645) & (g700) & (g1427) & (g1428) & (g1446)) + ((g645) & (!g700) & (!g1427) & (g1428) & (g1446)) + ((g645) & (!g700) & (g1427) & (!g1428) & (!g1446)) + ((g645) & (!g700) & (g1427) & (!g1428) & (g1446)) + ((g645) & (!g700) & (g1427) & (g1428) & (!g1446)) + ((g645) & (!g700) & (g1427) & (g1428) & (g1446)) + ((g645) & (g700) & (!g1427) & (!g1428) & (g1446)) + ((g645) & (g700) & (!g1427) & (g1428) & (!g1446)) + ((g645) & (g700) & (!g1427) & (g1428) & (g1446)) + ((g645) & (g700) & (g1427) & (!g1428) & (!g1446)) + ((g645) & (g700) & (g1427) & (!g1428) & (g1446)) + ((g645) & (g700) & (g1427) & (g1428) & (!g1446)) + ((g645) & (g700) & (g1427) & (g1428) & (g1446)));
	assign g1448 = (((!g553) & (!g604) & (g1425) & (g1426) & (g1447)) + ((!g553) & (g604) & (g1425) & (!g1426) & (g1447)) + ((!g553) & (g604) & (g1425) & (g1426) & (!g1447)) + ((!g553) & (g604) & (g1425) & (g1426) & (g1447)) + ((g553) & (!g604) & (!g1425) & (g1426) & (g1447)) + ((g553) & (!g604) & (g1425) & (!g1426) & (!g1447)) + ((g553) & (!g604) & (g1425) & (!g1426) & (g1447)) + ((g553) & (!g604) & (g1425) & (g1426) & (!g1447)) + ((g553) & (!g604) & (g1425) & (g1426) & (g1447)) + ((g553) & (g604) & (!g1425) & (!g1426) & (g1447)) + ((g553) & (g604) & (!g1425) & (g1426) & (!g1447)) + ((g553) & (g604) & (!g1425) & (g1426) & (g1447)) + ((g553) & (g604) & (g1425) & (!g1426) & (!g1447)) + ((g553) & (g604) & (g1425) & (!g1426) & (g1447)) + ((g553) & (g604) & (g1425) & (g1426) & (!g1447)) + ((g553) & (g604) & (g1425) & (g1426) & (g1447)));
	assign g1449 = (((g1) & (!g1372) & (g1419) & (g1422)) + ((g1) & (g1372) & (!g1419) & (!g1422)) + ((g1) & (g1372) & (!g1419) & (g1422)));
	assign g1450 = (((!g4) & (!g2) & (!g1373) & (!g1416) & (!g1418) & (!g1423)) + ((!g4) & (!g2) & (!g1373) & (!g1416) & (g1418) & (g1423)) + ((!g4) & (!g2) & (!g1373) & (g1416) & (!g1418) & (!g1423)) + ((!g4) & (!g2) & (!g1373) & (g1416) & (g1418) & (g1423)) + ((!g4) & (!g2) & (g1373) & (!g1416) & (!g1418) & (!g1423)) + ((!g4) & (!g2) & (g1373) & (!g1416) & (g1418) & (g1423)) + ((!g4) & (!g2) & (g1373) & (g1416) & (g1418) & (!g1423)) + ((!g4) & (!g2) & (g1373) & (g1416) & (g1418) & (g1423)) + ((!g4) & (g2) & (!g1373) & (!g1416) & (!g1418) & (!g1423)) + ((!g4) & (g2) & (!g1373) & (!g1416) & (g1418) & (g1423)) + ((!g4) & (g2) & (!g1373) & (g1416) & (g1418) & (!g1423)) + ((!g4) & (g2) & (!g1373) & (g1416) & (g1418) & (g1423)) + ((!g4) & (g2) & (g1373) & (!g1416) & (g1418) & (!g1423)) + ((!g4) & (g2) & (g1373) & (!g1416) & (g1418) & (g1423)) + ((!g4) & (g2) & (g1373) & (g1416) & (g1418) & (!g1423)) + ((!g4) & (g2) & (g1373) & (g1416) & (g1418) & (g1423)) + ((g4) & (!g2) & (!g1373) & (!g1416) & (g1418) & (!g1423)) + ((g4) & (!g2) & (!g1373) & (!g1416) & (g1418) & (g1423)) + ((g4) & (!g2) & (!g1373) & (g1416) & (g1418) & (!g1423)) + ((g4) & (!g2) & (!g1373) & (g1416) & (g1418) & (g1423)) + ((g4) & (!g2) & (g1373) & (!g1416) & (g1418) & (!g1423)) + ((g4) & (!g2) & (g1373) & (!g1416) & (g1418) & (g1423)) + ((g4) & (!g2) & (g1373) & (g1416) & (!g1418) & (!g1423)) + ((g4) & (!g2) & (g1373) & (g1416) & (g1418) & (g1423)) + ((g4) & (g2) & (!g1373) & (!g1416) & (g1418) & (!g1423)) + ((g4) & (g2) & (!g1373) & (!g1416) & (g1418) & (g1423)) + ((g4) & (g2) & (!g1373) & (g1416) & (!g1418) & (!g1423)) + ((g4) & (g2) & (!g1373) & (g1416) & (g1418) & (g1423)) + ((g4) & (g2) & (g1373) & (!g1416) & (!g1418) & (!g1423)) + ((g4) & (g2) & (g1373) & (!g1416) & (g1418) & (g1423)) + ((g4) & (g2) & (g1373) & (g1416) & (!g1418) & (!g1423)) + ((g4) & (g2) & (g1373) & (g1416) & (g1418) & (g1423)));
	assign g1451 = (((!g8) & (!g18) & (!g1375) & (g1376) & (g1415) & (!g1423)) + ((!g8) & (!g18) & (g1375) & (!g1376) & (!g1415) & (!g1423)) + ((!g8) & (!g18) & (g1375) & (!g1376) & (!g1415) & (g1423)) + ((!g8) & (!g18) & (g1375) & (!g1376) & (g1415) & (!g1423)) + ((!g8) & (!g18) & (g1375) & (!g1376) & (g1415) & (g1423)) + ((!g8) & (!g18) & (g1375) & (g1376) & (!g1415) & (!g1423)) + ((!g8) & (!g18) & (g1375) & (g1376) & (!g1415) & (g1423)) + ((!g8) & (!g18) & (g1375) & (g1376) & (g1415) & (g1423)) + ((!g8) & (g18) & (!g1375) & (!g1376) & (g1415) & (!g1423)) + ((!g8) & (g18) & (!g1375) & (g1376) & (!g1415) & (!g1423)) + ((!g8) & (g18) & (!g1375) & (g1376) & (g1415) & (!g1423)) + ((!g8) & (g18) & (g1375) & (!g1376) & (!g1415) & (!g1423)) + ((!g8) & (g18) & (g1375) & (!g1376) & (!g1415) & (g1423)) + ((!g8) & (g18) & (g1375) & (!g1376) & (g1415) & (g1423)) + ((!g8) & (g18) & (g1375) & (g1376) & (!g1415) & (g1423)) + ((!g8) & (g18) & (g1375) & (g1376) & (g1415) & (g1423)) + ((g8) & (!g18) & (!g1375) & (!g1376) & (!g1415) & (!g1423)) + ((g8) & (!g18) & (!g1375) & (!g1376) & (g1415) & (!g1423)) + ((g8) & (!g18) & (!g1375) & (g1376) & (!g1415) & (!g1423)) + ((g8) & (!g18) & (g1375) & (!g1376) & (!g1415) & (g1423)) + ((g8) & (!g18) & (g1375) & (!g1376) & (g1415) & (g1423)) + ((g8) & (!g18) & (g1375) & (g1376) & (!g1415) & (g1423)) + ((g8) & (!g18) & (g1375) & (g1376) & (g1415) & (!g1423)) + ((g8) & (!g18) & (g1375) & (g1376) & (g1415) & (g1423)) + ((g8) & (g18) & (!g1375) & (!g1376) & (!g1415) & (!g1423)) + ((g8) & (g18) & (g1375) & (!g1376) & (!g1415) & (g1423)) + ((g8) & (g18) & (g1375) & (!g1376) & (g1415) & (!g1423)) + ((g8) & (g18) & (g1375) & (!g1376) & (g1415) & (g1423)) + ((g8) & (g18) & (g1375) & (g1376) & (!g1415) & (!g1423)) + ((g8) & (g18) & (g1375) & (g1376) & (!g1415) & (g1423)) + ((g8) & (g18) & (g1375) & (g1376) & (g1415) & (!g1423)) + ((g8) & (g18) & (g1375) & (g1376) & (g1415) & (g1423)));
	assign g1452 = (((!g18) & (!g1376) & (g1415) & (!g1423)) + ((!g18) & (g1376) & (!g1415) & (!g1423)) + ((!g18) & (g1376) & (!g1415) & (g1423)) + ((!g18) & (g1376) & (g1415) & (g1423)) + ((g18) & (!g1376) & (!g1415) & (!g1423)) + ((g18) & (g1376) & (!g1415) & (g1423)) + ((g18) & (g1376) & (g1415) & (!g1423)) + ((g18) & (g1376) & (g1415) & (g1423)));
	assign g1453 = (((!g27) & (!g39) & (!g1378) & (g1379) & (g1414) & (!g1423)) + ((!g27) & (!g39) & (g1378) & (!g1379) & (!g1414) & (!g1423)) + ((!g27) & (!g39) & (g1378) & (!g1379) & (!g1414) & (g1423)) + ((!g27) & (!g39) & (g1378) & (!g1379) & (g1414) & (!g1423)) + ((!g27) & (!g39) & (g1378) & (!g1379) & (g1414) & (g1423)) + ((!g27) & (!g39) & (g1378) & (g1379) & (!g1414) & (!g1423)) + ((!g27) & (!g39) & (g1378) & (g1379) & (!g1414) & (g1423)) + ((!g27) & (!g39) & (g1378) & (g1379) & (g1414) & (g1423)) + ((!g27) & (g39) & (!g1378) & (!g1379) & (g1414) & (!g1423)) + ((!g27) & (g39) & (!g1378) & (g1379) & (!g1414) & (!g1423)) + ((!g27) & (g39) & (!g1378) & (g1379) & (g1414) & (!g1423)) + ((!g27) & (g39) & (g1378) & (!g1379) & (!g1414) & (!g1423)) + ((!g27) & (g39) & (g1378) & (!g1379) & (!g1414) & (g1423)) + ((!g27) & (g39) & (g1378) & (!g1379) & (g1414) & (g1423)) + ((!g27) & (g39) & (g1378) & (g1379) & (!g1414) & (g1423)) + ((!g27) & (g39) & (g1378) & (g1379) & (g1414) & (g1423)) + ((g27) & (!g39) & (!g1378) & (!g1379) & (!g1414) & (!g1423)) + ((g27) & (!g39) & (!g1378) & (!g1379) & (g1414) & (!g1423)) + ((g27) & (!g39) & (!g1378) & (g1379) & (!g1414) & (!g1423)) + ((g27) & (!g39) & (g1378) & (!g1379) & (!g1414) & (g1423)) + ((g27) & (!g39) & (g1378) & (!g1379) & (g1414) & (g1423)) + ((g27) & (!g39) & (g1378) & (g1379) & (!g1414) & (g1423)) + ((g27) & (!g39) & (g1378) & (g1379) & (g1414) & (!g1423)) + ((g27) & (!g39) & (g1378) & (g1379) & (g1414) & (g1423)) + ((g27) & (g39) & (!g1378) & (!g1379) & (!g1414) & (!g1423)) + ((g27) & (g39) & (g1378) & (!g1379) & (!g1414) & (g1423)) + ((g27) & (g39) & (g1378) & (!g1379) & (g1414) & (!g1423)) + ((g27) & (g39) & (g1378) & (!g1379) & (g1414) & (g1423)) + ((g27) & (g39) & (g1378) & (g1379) & (!g1414) & (!g1423)) + ((g27) & (g39) & (g1378) & (g1379) & (!g1414) & (g1423)) + ((g27) & (g39) & (g1378) & (g1379) & (g1414) & (!g1423)) + ((g27) & (g39) & (g1378) & (g1379) & (g1414) & (g1423)));
	assign g1454 = (((!g39) & (!g1379) & (g1414) & (!g1423)) + ((!g39) & (g1379) & (!g1414) & (!g1423)) + ((!g39) & (g1379) & (!g1414) & (g1423)) + ((!g39) & (g1379) & (g1414) & (g1423)) + ((g39) & (!g1379) & (!g1414) & (!g1423)) + ((g39) & (g1379) & (!g1414) & (g1423)) + ((g39) & (g1379) & (g1414) & (!g1423)) + ((g39) & (g1379) & (g1414) & (g1423)));
	assign g1455 = (((!g54) & (!g68) & (!g1381) & (g1382) & (g1413) & (!g1423)) + ((!g54) & (!g68) & (g1381) & (!g1382) & (!g1413) & (!g1423)) + ((!g54) & (!g68) & (g1381) & (!g1382) & (!g1413) & (g1423)) + ((!g54) & (!g68) & (g1381) & (!g1382) & (g1413) & (!g1423)) + ((!g54) & (!g68) & (g1381) & (!g1382) & (g1413) & (g1423)) + ((!g54) & (!g68) & (g1381) & (g1382) & (!g1413) & (!g1423)) + ((!g54) & (!g68) & (g1381) & (g1382) & (!g1413) & (g1423)) + ((!g54) & (!g68) & (g1381) & (g1382) & (g1413) & (g1423)) + ((!g54) & (g68) & (!g1381) & (!g1382) & (g1413) & (!g1423)) + ((!g54) & (g68) & (!g1381) & (g1382) & (!g1413) & (!g1423)) + ((!g54) & (g68) & (!g1381) & (g1382) & (g1413) & (!g1423)) + ((!g54) & (g68) & (g1381) & (!g1382) & (!g1413) & (!g1423)) + ((!g54) & (g68) & (g1381) & (!g1382) & (!g1413) & (g1423)) + ((!g54) & (g68) & (g1381) & (!g1382) & (g1413) & (g1423)) + ((!g54) & (g68) & (g1381) & (g1382) & (!g1413) & (g1423)) + ((!g54) & (g68) & (g1381) & (g1382) & (g1413) & (g1423)) + ((g54) & (!g68) & (!g1381) & (!g1382) & (!g1413) & (!g1423)) + ((g54) & (!g68) & (!g1381) & (!g1382) & (g1413) & (!g1423)) + ((g54) & (!g68) & (!g1381) & (g1382) & (!g1413) & (!g1423)) + ((g54) & (!g68) & (g1381) & (!g1382) & (!g1413) & (g1423)) + ((g54) & (!g68) & (g1381) & (!g1382) & (g1413) & (g1423)) + ((g54) & (!g68) & (g1381) & (g1382) & (!g1413) & (g1423)) + ((g54) & (!g68) & (g1381) & (g1382) & (g1413) & (!g1423)) + ((g54) & (!g68) & (g1381) & (g1382) & (g1413) & (g1423)) + ((g54) & (g68) & (!g1381) & (!g1382) & (!g1413) & (!g1423)) + ((g54) & (g68) & (g1381) & (!g1382) & (!g1413) & (g1423)) + ((g54) & (g68) & (g1381) & (!g1382) & (g1413) & (!g1423)) + ((g54) & (g68) & (g1381) & (!g1382) & (g1413) & (g1423)) + ((g54) & (g68) & (g1381) & (g1382) & (!g1413) & (!g1423)) + ((g54) & (g68) & (g1381) & (g1382) & (!g1413) & (g1423)) + ((g54) & (g68) & (g1381) & (g1382) & (g1413) & (!g1423)) + ((g54) & (g68) & (g1381) & (g1382) & (g1413) & (g1423)));
	assign g1456 = (((!g68) & (!g1382) & (g1413) & (!g1423)) + ((!g68) & (g1382) & (!g1413) & (!g1423)) + ((!g68) & (g1382) & (!g1413) & (g1423)) + ((!g68) & (g1382) & (g1413) & (g1423)) + ((g68) & (!g1382) & (!g1413) & (!g1423)) + ((g68) & (g1382) & (!g1413) & (g1423)) + ((g68) & (g1382) & (g1413) & (!g1423)) + ((g68) & (g1382) & (g1413) & (g1423)));
	assign g1457 = (((!g87) & (!g104) & (!g1384) & (g1385) & (g1412) & (!g1423)) + ((!g87) & (!g104) & (g1384) & (!g1385) & (!g1412) & (!g1423)) + ((!g87) & (!g104) & (g1384) & (!g1385) & (!g1412) & (g1423)) + ((!g87) & (!g104) & (g1384) & (!g1385) & (g1412) & (!g1423)) + ((!g87) & (!g104) & (g1384) & (!g1385) & (g1412) & (g1423)) + ((!g87) & (!g104) & (g1384) & (g1385) & (!g1412) & (!g1423)) + ((!g87) & (!g104) & (g1384) & (g1385) & (!g1412) & (g1423)) + ((!g87) & (!g104) & (g1384) & (g1385) & (g1412) & (g1423)) + ((!g87) & (g104) & (!g1384) & (!g1385) & (g1412) & (!g1423)) + ((!g87) & (g104) & (!g1384) & (g1385) & (!g1412) & (!g1423)) + ((!g87) & (g104) & (!g1384) & (g1385) & (g1412) & (!g1423)) + ((!g87) & (g104) & (g1384) & (!g1385) & (!g1412) & (!g1423)) + ((!g87) & (g104) & (g1384) & (!g1385) & (!g1412) & (g1423)) + ((!g87) & (g104) & (g1384) & (!g1385) & (g1412) & (g1423)) + ((!g87) & (g104) & (g1384) & (g1385) & (!g1412) & (g1423)) + ((!g87) & (g104) & (g1384) & (g1385) & (g1412) & (g1423)) + ((g87) & (!g104) & (!g1384) & (!g1385) & (!g1412) & (!g1423)) + ((g87) & (!g104) & (!g1384) & (!g1385) & (g1412) & (!g1423)) + ((g87) & (!g104) & (!g1384) & (g1385) & (!g1412) & (!g1423)) + ((g87) & (!g104) & (g1384) & (!g1385) & (!g1412) & (g1423)) + ((g87) & (!g104) & (g1384) & (!g1385) & (g1412) & (g1423)) + ((g87) & (!g104) & (g1384) & (g1385) & (!g1412) & (g1423)) + ((g87) & (!g104) & (g1384) & (g1385) & (g1412) & (!g1423)) + ((g87) & (!g104) & (g1384) & (g1385) & (g1412) & (g1423)) + ((g87) & (g104) & (!g1384) & (!g1385) & (!g1412) & (!g1423)) + ((g87) & (g104) & (g1384) & (!g1385) & (!g1412) & (g1423)) + ((g87) & (g104) & (g1384) & (!g1385) & (g1412) & (!g1423)) + ((g87) & (g104) & (g1384) & (!g1385) & (g1412) & (g1423)) + ((g87) & (g104) & (g1384) & (g1385) & (!g1412) & (!g1423)) + ((g87) & (g104) & (g1384) & (g1385) & (!g1412) & (g1423)) + ((g87) & (g104) & (g1384) & (g1385) & (g1412) & (!g1423)) + ((g87) & (g104) & (g1384) & (g1385) & (g1412) & (g1423)));
	assign g1458 = (((!g104) & (!g1385) & (g1412) & (!g1423)) + ((!g104) & (g1385) & (!g1412) & (!g1423)) + ((!g104) & (g1385) & (!g1412) & (g1423)) + ((!g104) & (g1385) & (g1412) & (g1423)) + ((g104) & (!g1385) & (!g1412) & (!g1423)) + ((g104) & (g1385) & (!g1412) & (g1423)) + ((g104) & (g1385) & (g1412) & (!g1423)) + ((g104) & (g1385) & (g1412) & (g1423)));
	assign g1459 = (((!g127) & (!g147) & (!g1387) & (g1388) & (g1411) & (!g1423)) + ((!g127) & (!g147) & (g1387) & (!g1388) & (!g1411) & (!g1423)) + ((!g127) & (!g147) & (g1387) & (!g1388) & (!g1411) & (g1423)) + ((!g127) & (!g147) & (g1387) & (!g1388) & (g1411) & (!g1423)) + ((!g127) & (!g147) & (g1387) & (!g1388) & (g1411) & (g1423)) + ((!g127) & (!g147) & (g1387) & (g1388) & (!g1411) & (!g1423)) + ((!g127) & (!g147) & (g1387) & (g1388) & (!g1411) & (g1423)) + ((!g127) & (!g147) & (g1387) & (g1388) & (g1411) & (g1423)) + ((!g127) & (g147) & (!g1387) & (!g1388) & (g1411) & (!g1423)) + ((!g127) & (g147) & (!g1387) & (g1388) & (!g1411) & (!g1423)) + ((!g127) & (g147) & (!g1387) & (g1388) & (g1411) & (!g1423)) + ((!g127) & (g147) & (g1387) & (!g1388) & (!g1411) & (!g1423)) + ((!g127) & (g147) & (g1387) & (!g1388) & (!g1411) & (g1423)) + ((!g127) & (g147) & (g1387) & (!g1388) & (g1411) & (g1423)) + ((!g127) & (g147) & (g1387) & (g1388) & (!g1411) & (g1423)) + ((!g127) & (g147) & (g1387) & (g1388) & (g1411) & (g1423)) + ((g127) & (!g147) & (!g1387) & (!g1388) & (!g1411) & (!g1423)) + ((g127) & (!g147) & (!g1387) & (!g1388) & (g1411) & (!g1423)) + ((g127) & (!g147) & (!g1387) & (g1388) & (!g1411) & (!g1423)) + ((g127) & (!g147) & (g1387) & (!g1388) & (!g1411) & (g1423)) + ((g127) & (!g147) & (g1387) & (!g1388) & (g1411) & (g1423)) + ((g127) & (!g147) & (g1387) & (g1388) & (!g1411) & (g1423)) + ((g127) & (!g147) & (g1387) & (g1388) & (g1411) & (!g1423)) + ((g127) & (!g147) & (g1387) & (g1388) & (g1411) & (g1423)) + ((g127) & (g147) & (!g1387) & (!g1388) & (!g1411) & (!g1423)) + ((g127) & (g147) & (g1387) & (!g1388) & (!g1411) & (g1423)) + ((g127) & (g147) & (g1387) & (!g1388) & (g1411) & (!g1423)) + ((g127) & (g147) & (g1387) & (!g1388) & (g1411) & (g1423)) + ((g127) & (g147) & (g1387) & (g1388) & (!g1411) & (!g1423)) + ((g127) & (g147) & (g1387) & (g1388) & (!g1411) & (g1423)) + ((g127) & (g147) & (g1387) & (g1388) & (g1411) & (!g1423)) + ((g127) & (g147) & (g1387) & (g1388) & (g1411) & (g1423)));
	assign g1460 = (((!g147) & (!g1388) & (g1411) & (!g1423)) + ((!g147) & (g1388) & (!g1411) & (!g1423)) + ((!g147) & (g1388) & (!g1411) & (g1423)) + ((!g147) & (g1388) & (g1411) & (g1423)) + ((g147) & (!g1388) & (!g1411) & (!g1423)) + ((g147) & (g1388) & (!g1411) & (g1423)) + ((g147) & (g1388) & (g1411) & (!g1423)) + ((g147) & (g1388) & (g1411) & (g1423)));
	assign g1461 = (((!g174) & (!g198) & (!g1390) & (g1391) & (g1410) & (!g1423)) + ((!g174) & (!g198) & (g1390) & (!g1391) & (!g1410) & (!g1423)) + ((!g174) & (!g198) & (g1390) & (!g1391) & (!g1410) & (g1423)) + ((!g174) & (!g198) & (g1390) & (!g1391) & (g1410) & (!g1423)) + ((!g174) & (!g198) & (g1390) & (!g1391) & (g1410) & (g1423)) + ((!g174) & (!g198) & (g1390) & (g1391) & (!g1410) & (!g1423)) + ((!g174) & (!g198) & (g1390) & (g1391) & (!g1410) & (g1423)) + ((!g174) & (!g198) & (g1390) & (g1391) & (g1410) & (g1423)) + ((!g174) & (g198) & (!g1390) & (!g1391) & (g1410) & (!g1423)) + ((!g174) & (g198) & (!g1390) & (g1391) & (!g1410) & (!g1423)) + ((!g174) & (g198) & (!g1390) & (g1391) & (g1410) & (!g1423)) + ((!g174) & (g198) & (g1390) & (!g1391) & (!g1410) & (!g1423)) + ((!g174) & (g198) & (g1390) & (!g1391) & (!g1410) & (g1423)) + ((!g174) & (g198) & (g1390) & (!g1391) & (g1410) & (g1423)) + ((!g174) & (g198) & (g1390) & (g1391) & (!g1410) & (g1423)) + ((!g174) & (g198) & (g1390) & (g1391) & (g1410) & (g1423)) + ((g174) & (!g198) & (!g1390) & (!g1391) & (!g1410) & (!g1423)) + ((g174) & (!g198) & (!g1390) & (!g1391) & (g1410) & (!g1423)) + ((g174) & (!g198) & (!g1390) & (g1391) & (!g1410) & (!g1423)) + ((g174) & (!g198) & (g1390) & (!g1391) & (!g1410) & (g1423)) + ((g174) & (!g198) & (g1390) & (!g1391) & (g1410) & (g1423)) + ((g174) & (!g198) & (g1390) & (g1391) & (!g1410) & (g1423)) + ((g174) & (!g198) & (g1390) & (g1391) & (g1410) & (!g1423)) + ((g174) & (!g198) & (g1390) & (g1391) & (g1410) & (g1423)) + ((g174) & (g198) & (!g1390) & (!g1391) & (!g1410) & (!g1423)) + ((g174) & (g198) & (g1390) & (!g1391) & (!g1410) & (g1423)) + ((g174) & (g198) & (g1390) & (!g1391) & (g1410) & (!g1423)) + ((g174) & (g198) & (g1390) & (!g1391) & (g1410) & (g1423)) + ((g174) & (g198) & (g1390) & (g1391) & (!g1410) & (!g1423)) + ((g174) & (g198) & (g1390) & (g1391) & (!g1410) & (g1423)) + ((g174) & (g198) & (g1390) & (g1391) & (g1410) & (!g1423)) + ((g174) & (g198) & (g1390) & (g1391) & (g1410) & (g1423)));
	assign g1462 = (((!g198) & (!g1391) & (g1410) & (!g1423)) + ((!g198) & (g1391) & (!g1410) & (!g1423)) + ((!g198) & (g1391) & (!g1410) & (g1423)) + ((!g198) & (g1391) & (g1410) & (g1423)) + ((g198) & (!g1391) & (!g1410) & (!g1423)) + ((g198) & (g1391) & (!g1410) & (g1423)) + ((g198) & (g1391) & (g1410) & (!g1423)) + ((g198) & (g1391) & (g1410) & (g1423)));
	assign g1463 = (((!g229) & (!g255) & (!g1393) & (g1394) & (g1409) & (!g1423)) + ((!g229) & (!g255) & (g1393) & (!g1394) & (!g1409) & (!g1423)) + ((!g229) & (!g255) & (g1393) & (!g1394) & (!g1409) & (g1423)) + ((!g229) & (!g255) & (g1393) & (!g1394) & (g1409) & (!g1423)) + ((!g229) & (!g255) & (g1393) & (!g1394) & (g1409) & (g1423)) + ((!g229) & (!g255) & (g1393) & (g1394) & (!g1409) & (!g1423)) + ((!g229) & (!g255) & (g1393) & (g1394) & (!g1409) & (g1423)) + ((!g229) & (!g255) & (g1393) & (g1394) & (g1409) & (g1423)) + ((!g229) & (g255) & (!g1393) & (!g1394) & (g1409) & (!g1423)) + ((!g229) & (g255) & (!g1393) & (g1394) & (!g1409) & (!g1423)) + ((!g229) & (g255) & (!g1393) & (g1394) & (g1409) & (!g1423)) + ((!g229) & (g255) & (g1393) & (!g1394) & (!g1409) & (!g1423)) + ((!g229) & (g255) & (g1393) & (!g1394) & (!g1409) & (g1423)) + ((!g229) & (g255) & (g1393) & (!g1394) & (g1409) & (g1423)) + ((!g229) & (g255) & (g1393) & (g1394) & (!g1409) & (g1423)) + ((!g229) & (g255) & (g1393) & (g1394) & (g1409) & (g1423)) + ((g229) & (!g255) & (!g1393) & (!g1394) & (!g1409) & (!g1423)) + ((g229) & (!g255) & (!g1393) & (!g1394) & (g1409) & (!g1423)) + ((g229) & (!g255) & (!g1393) & (g1394) & (!g1409) & (!g1423)) + ((g229) & (!g255) & (g1393) & (!g1394) & (!g1409) & (g1423)) + ((g229) & (!g255) & (g1393) & (!g1394) & (g1409) & (g1423)) + ((g229) & (!g255) & (g1393) & (g1394) & (!g1409) & (g1423)) + ((g229) & (!g255) & (g1393) & (g1394) & (g1409) & (!g1423)) + ((g229) & (!g255) & (g1393) & (g1394) & (g1409) & (g1423)) + ((g229) & (g255) & (!g1393) & (!g1394) & (!g1409) & (!g1423)) + ((g229) & (g255) & (g1393) & (!g1394) & (!g1409) & (g1423)) + ((g229) & (g255) & (g1393) & (!g1394) & (g1409) & (!g1423)) + ((g229) & (g255) & (g1393) & (!g1394) & (g1409) & (g1423)) + ((g229) & (g255) & (g1393) & (g1394) & (!g1409) & (!g1423)) + ((g229) & (g255) & (g1393) & (g1394) & (!g1409) & (g1423)) + ((g229) & (g255) & (g1393) & (g1394) & (g1409) & (!g1423)) + ((g229) & (g255) & (g1393) & (g1394) & (g1409) & (g1423)));
	assign g1464 = (((!g255) & (!g1394) & (g1409) & (!g1423)) + ((!g255) & (g1394) & (!g1409) & (!g1423)) + ((!g255) & (g1394) & (!g1409) & (g1423)) + ((!g255) & (g1394) & (g1409) & (g1423)) + ((g255) & (!g1394) & (!g1409) & (!g1423)) + ((g255) & (g1394) & (!g1409) & (g1423)) + ((g255) & (g1394) & (g1409) & (!g1423)) + ((g255) & (g1394) & (g1409) & (g1423)));
	assign g1465 = (((!g290) & (!g319) & (!g1396) & (g1397) & (g1408) & (!g1423)) + ((!g290) & (!g319) & (g1396) & (!g1397) & (!g1408) & (!g1423)) + ((!g290) & (!g319) & (g1396) & (!g1397) & (!g1408) & (g1423)) + ((!g290) & (!g319) & (g1396) & (!g1397) & (g1408) & (!g1423)) + ((!g290) & (!g319) & (g1396) & (!g1397) & (g1408) & (g1423)) + ((!g290) & (!g319) & (g1396) & (g1397) & (!g1408) & (!g1423)) + ((!g290) & (!g319) & (g1396) & (g1397) & (!g1408) & (g1423)) + ((!g290) & (!g319) & (g1396) & (g1397) & (g1408) & (g1423)) + ((!g290) & (g319) & (!g1396) & (!g1397) & (g1408) & (!g1423)) + ((!g290) & (g319) & (!g1396) & (g1397) & (!g1408) & (!g1423)) + ((!g290) & (g319) & (!g1396) & (g1397) & (g1408) & (!g1423)) + ((!g290) & (g319) & (g1396) & (!g1397) & (!g1408) & (!g1423)) + ((!g290) & (g319) & (g1396) & (!g1397) & (!g1408) & (g1423)) + ((!g290) & (g319) & (g1396) & (!g1397) & (g1408) & (g1423)) + ((!g290) & (g319) & (g1396) & (g1397) & (!g1408) & (g1423)) + ((!g290) & (g319) & (g1396) & (g1397) & (g1408) & (g1423)) + ((g290) & (!g319) & (!g1396) & (!g1397) & (!g1408) & (!g1423)) + ((g290) & (!g319) & (!g1396) & (!g1397) & (g1408) & (!g1423)) + ((g290) & (!g319) & (!g1396) & (g1397) & (!g1408) & (!g1423)) + ((g290) & (!g319) & (g1396) & (!g1397) & (!g1408) & (g1423)) + ((g290) & (!g319) & (g1396) & (!g1397) & (g1408) & (g1423)) + ((g290) & (!g319) & (g1396) & (g1397) & (!g1408) & (g1423)) + ((g290) & (!g319) & (g1396) & (g1397) & (g1408) & (!g1423)) + ((g290) & (!g319) & (g1396) & (g1397) & (g1408) & (g1423)) + ((g290) & (g319) & (!g1396) & (!g1397) & (!g1408) & (!g1423)) + ((g290) & (g319) & (g1396) & (!g1397) & (!g1408) & (g1423)) + ((g290) & (g319) & (g1396) & (!g1397) & (g1408) & (!g1423)) + ((g290) & (g319) & (g1396) & (!g1397) & (g1408) & (g1423)) + ((g290) & (g319) & (g1396) & (g1397) & (!g1408) & (!g1423)) + ((g290) & (g319) & (g1396) & (g1397) & (!g1408) & (g1423)) + ((g290) & (g319) & (g1396) & (g1397) & (g1408) & (!g1423)) + ((g290) & (g319) & (g1396) & (g1397) & (g1408) & (g1423)));
	assign g1466 = (((!g319) & (!g1397) & (g1408) & (!g1423)) + ((!g319) & (g1397) & (!g1408) & (!g1423)) + ((!g319) & (g1397) & (!g1408) & (g1423)) + ((!g319) & (g1397) & (g1408) & (g1423)) + ((g319) & (!g1397) & (!g1408) & (!g1423)) + ((g319) & (g1397) & (!g1408) & (g1423)) + ((g319) & (g1397) & (g1408) & (!g1423)) + ((g319) & (g1397) & (g1408) & (g1423)));
	assign g1467 = (((!g358) & (!g390) & (!g1399) & (g1400) & (g1407) & (!g1423)) + ((!g358) & (!g390) & (g1399) & (!g1400) & (!g1407) & (!g1423)) + ((!g358) & (!g390) & (g1399) & (!g1400) & (!g1407) & (g1423)) + ((!g358) & (!g390) & (g1399) & (!g1400) & (g1407) & (!g1423)) + ((!g358) & (!g390) & (g1399) & (!g1400) & (g1407) & (g1423)) + ((!g358) & (!g390) & (g1399) & (g1400) & (!g1407) & (!g1423)) + ((!g358) & (!g390) & (g1399) & (g1400) & (!g1407) & (g1423)) + ((!g358) & (!g390) & (g1399) & (g1400) & (g1407) & (g1423)) + ((!g358) & (g390) & (!g1399) & (!g1400) & (g1407) & (!g1423)) + ((!g358) & (g390) & (!g1399) & (g1400) & (!g1407) & (!g1423)) + ((!g358) & (g390) & (!g1399) & (g1400) & (g1407) & (!g1423)) + ((!g358) & (g390) & (g1399) & (!g1400) & (!g1407) & (!g1423)) + ((!g358) & (g390) & (g1399) & (!g1400) & (!g1407) & (g1423)) + ((!g358) & (g390) & (g1399) & (!g1400) & (g1407) & (g1423)) + ((!g358) & (g390) & (g1399) & (g1400) & (!g1407) & (g1423)) + ((!g358) & (g390) & (g1399) & (g1400) & (g1407) & (g1423)) + ((g358) & (!g390) & (!g1399) & (!g1400) & (!g1407) & (!g1423)) + ((g358) & (!g390) & (!g1399) & (!g1400) & (g1407) & (!g1423)) + ((g358) & (!g390) & (!g1399) & (g1400) & (!g1407) & (!g1423)) + ((g358) & (!g390) & (g1399) & (!g1400) & (!g1407) & (g1423)) + ((g358) & (!g390) & (g1399) & (!g1400) & (g1407) & (g1423)) + ((g358) & (!g390) & (g1399) & (g1400) & (!g1407) & (g1423)) + ((g358) & (!g390) & (g1399) & (g1400) & (g1407) & (!g1423)) + ((g358) & (!g390) & (g1399) & (g1400) & (g1407) & (g1423)) + ((g358) & (g390) & (!g1399) & (!g1400) & (!g1407) & (!g1423)) + ((g358) & (g390) & (g1399) & (!g1400) & (!g1407) & (g1423)) + ((g358) & (g390) & (g1399) & (!g1400) & (g1407) & (!g1423)) + ((g358) & (g390) & (g1399) & (!g1400) & (g1407) & (g1423)) + ((g358) & (g390) & (g1399) & (g1400) & (!g1407) & (!g1423)) + ((g358) & (g390) & (g1399) & (g1400) & (!g1407) & (g1423)) + ((g358) & (g390) & (g1399) & (g1400) & (g1407) & (!g1423)) + ((g358) & (g390) & (g1399) & (g1400) & (g1407) & (g1423)));
	assign g1468 = (((!g390) & (!g1400) & (g1407) & (!g1423)) + ((!g390) & (g1400) & (!g1407) & (!g1423)) + ((!g390) & (g1400) & (!g1407) & (g1423)) + ((!g390) & (g1400) & (g1407) & (g1423)) + ((g390) & (!g1400) & (!g1407) & (!g1423)) + ((g390) & (g1400) & (!g1407) & (g1423)) + ((g390) & (g1400) & (g1407) & (!g1423)) + ((g390) & (g1400) & (g1407) & (g1423)));
	assign g1469 = (((!g433) & (!g468) & (!g1402) & (g1403) & (g1406) & (!g1423)) + ((!g433) & (!g468) & (g1402) & (!g1403) & (!g1406) & (!g1423)) + ((!g433) & (!g468) & (g1402) & (!g1403) & (!g1406) & (g1423)) + ((!g433) & (!g468) & (g1402) & (!g1403) & (g1406) & (!g1423)) + ((!g433) & (!g468) & (g1402) & (!g1403) & (g1406) & (g1423)) + ((!g433) & (!g468) & (g1402) & (g1403) & (!g1406) & (!g1423)) + ((!g433) & (!g468) & (g1402) & (g1403) & (!g1406) & (g1423)) + ((!g433) & (!g468) & (g1402) & (g1403) & (g1406) & (g1423)) + ((!g433) & (g468) & (!g1402) & (!g1403) & (g1406) & (!g1423)) + ((!g433) & (g468) & (!g1402) & (g1403) & (!g1406) & (!g1423)) + ((!g433) & (g468) & (!g1402) & (g1403) & (g1406) & (!g1423)) + ((!g433) & (g468) & (g1402) & (!g1403) & (!g1406) & (!g1423)) + ((!g433) & (g468) & (g1402) & (!g1403) & (!g1406) & (g1423)) + ((!g433) & (g468) & (g1402) & (!g1403) & (g1406) & (g1423)) + ((!g433) & (g468) & (g1402) & (g1403) & (!g1406) & (g1423)) + ((!g433) & (g468) & (g1402) & (g1403) & (g1406) & (g1423)) + ((g433) & (!g468) & (!g1402) & (!g1403) & (!g1406) & (!g1423)) + ((g433) & (!g468) & (!g1402) & (!g1403) & (g1406) & (!g1423)) + ((g433) & (!g468) & (!g1402) & (g1403) & (!g1406) & (!g1423)) + ((g433) & (!g468) & (g1402) & (!g1403) & (!g1406) & (g1423)) + ((g433) & (!g468) & (g1402) & (!g1403) & (g1406) & (g1423)) + ((g433) & (!g468) & (g1402) & (g1403) & (!g1406) & (g1423)) + ((g433) & (!g468) & (g1402) & (g1403) & (g1406) & (!g1423)) + ((g433) & (!g468) & (g1402) & (g1403) & (g1406) & (g1423)) + ((g433) & (g468) & (!g1402) & (!g1403) & (!g1406) & (!g1423)) + ((g433) & (g468) & (g1402) & (!g1403) & (!g1406) & (g1423)) + ((g433) & (g468) & (g1402) & (!g1403) & (g1406) & (!g1423)) + ((g433) & (g468) & (g1402) & (!g1403) & (g1406) & (g1423)) + ((g433) & (g468) & (g1402) & (g1403) & (!g1406) & (!g1423)) + ((g433) & (g468) & (g1402) & (g1403) & (!g1406) & (g1423)) + ((g433) & (g468) & (g1402) & (g1403) & (g1406) & (!g1423)) + ((g433) & (g468) & (g1402) & (g1403) & (g1406) & (g1423)));
	assign g1470 = (((!g468) & (!g1403) & (g1406) & (!g1423)) + ((!g468) & (g1403) & (!g1406) & (!g1423)) + ((!g468) & (g1403) & (!g1406) & (g1423)) + ((!g468) & (g1403) & (g1406) & (g1423)) + ((g468) & (!g1403) & (!g1406) & (!g1423)) + ((g468) & (g1403) & (!g1406) & (g1423)) + ((g468) & (g1403) & (g1406) & (!g1423)) + ((g468) & (g1403) & (g1406) & (g1423)));
	assign g1471 = (((!g515) & (!g553) & (!g1405) & (g1345) & (g1371) & (!g1423)) + ((!g515) & (!g553) & (g1405) & (!g1345) & (!g1371) & (!g1423)) + ((!g515) & (!g553) & (g1405) & (!g1345) & (!g1371) & (g1423)) + ((!g515) & (!g553) & (g1405) & (!g1345) & (g1371) & (!g1423)) + ((!g515) & (!g553) & (g1405) & (!g1345) & (g1371) & (g1423)) + ((!g515) & (!g553) & (g1405) & (g1345) & (!g1371) & (!g1423)) + ((!g515) & (!g553) & (g1405) & (g1345) & (!g1371) & (g1423)) + ((!g515) & (!g553) & (g1405) & (g1345) & (g1371) & (g1423)) + ((!g515) & (g553) & (!g1405) & (!g1345) & (g1371) & (!g1423)) + ((!g515) & (g553) & (!g1405) & (g1345) & (!g1371) & (!g1423)) + ((!g515) & (g553) & (!g1405) & (g1345) & (g1371) & (!g1423)) + ((!g515) & (g553) & (g1405) & (!g1345) & (!g1371) & (!g1423)) + ((!g515) & (g553) & (g1405) & (!g1345) & (!g1371) & (g1423)) + ((!g515) & (g553) & (g1405) & (!g1345) & (g1371) & (g1423)) + ((!g515) & (g553) & (g1405) & (g1345) & (!g1371) & (g1423)) + ((!g515) & (g553) & (g1405) & (g1345) & (g1371) & (g1423)) + ((g515) & (!g553) & (!g1405) & (!g1345) & (!g1371) & (!g1423)) + ((g515) & (!g553) & (!g1405) & (!g1345) & (g1371) & (!g1423)) + ((g515) & (!g553) & (!g1405) & (g1345) & (!g1371) & (!g1423)) + ((g515) & (!g553) & (g1405) & (!g1345) & (!g1371) & (g1423)) + ((g515) & (!g553) & (g1405) & (!g1345) & (g1371) & (g1423)) + ((g515) & (!g553) & (g1405) & (g1345) & (!g1371) & (g1423)) + ((g515) & (!g553) & (g1405) & (g1345) & (g1371) & (!g1423)) + ((g515) & (!g553) & (g1405) & (g1345) & (g1371) & (g1423)) + ((g515) & (g553) & (!g1405) & (!g1345) & (!g1371) & (!g1423)) + ((g515) & (g553) & (g1405) & (!g1345) & (!g1371) & (g1423)) + ((g515) & (g553) & (g1405) & (!g1345) & (g1371) & (!g1423)) + ((g515) & (g553) & (g1405) & (!g1345) & (g1371) & (g1423)) + ((g515) & (g553) & (g1405) & (g1345) & (!g1371) & (!g1423)) + ((g515) & (g553) & (g1405) & (g1345) & (!g1371) & (g1423)) + ((g515) & (g553) & (g1405) & (g1345) & (g1371) & (!g1423)) + ((g515) & (g553) & (g1405) & (g1345) & (g1371) & (g1423)));
	assign g1472 = (((!g468) & (!g515) & (g1471) & (g1424) & (g1448)) + ((!g468) & (g515) & (g1471) & (!g1424) & (g1448)) + ((!g468) & (g515) & (g1471) & (g1424) & (!g1448)) + ((!g468) & (g515) & (g1471) & (g1424) & (g1448)) + ((g468) & (!g515) & (!g1471) & (g1424) & (g1448)) + ((g468) & (!g515) & (g1471) & (!g1424) & (!g1448)) + ((g468) & (!g515) & (g1471) & (!g1424) & (g1448)) + ((g468) & (!g515) & (g1471) & (g1424) & (!g1448)) + ((g468) & (!g515) & (g1471) & (g1424) & (g1448)) + ((g468) & (g515) & (!g1471) & (!g1424) & (g1448)) + ((g468) & (g515) & (!g1471) & (g1424) & (!g1448)) + ((g468) & (g515) & (!g1471) & (g1424) & (g1448)) + ((g468) & (g515) & (g1471) & (!g1424) & (!g1448)) + ((g468) & (g515) & (g1471) & (!g1424) & (g1448)) + ((g468) & (g515) & (g1471) & (g1424) & (!g1448)) + ((g468) & (g515) & (g1471) & (g1424) & (g1448)));
	assign g1473 = (((!g390) & (!g433) & (g1469) & (g1470) & (g1472)) + ((!g390) & (g433) & (g1469) & (!g1470) & (g1472)) + ((!g390) & (g433) & (g1469) & (g1470) & (!g1472)) + ((!g390) & (g433) & (g1469) & (g1470) & (g1472)) + ((g390) & (!g433) & (!g1469) & (g1470) & (g1472)) + ((g390) & (!g433) & (g1469) & (!g1470) & (!g1472)) + ((g390) & (!g433) & (g1469) & (!g1470) & (g1472)) + ((g390) & (!g433) & (g1469) & (g1470) & (!g1472)) + ((g390) & (!g433) & (g1469) & (g1470) & (g1472)) + ((g390) & (g433) & (!g1469) & (!g1470) & (g1472)) + ((g390) & (g433) & (!g1469) & (g1470) & (!g1472)) + ((g390) & (g433) & (!g1469) & (g1470) & (g1472)) + ((g390) & (g433) & (g1469) & (!g1470) & (!g1472)) + ((g390) & (g433) & (g1469) & (!g1470) & (g1472)) + ((g390) & (g433) & (g1469) & (g1470) & (!g1472)) + ((g390) & (g433) & (g1469) & (g1470) & (g1472)));
	assign g1474 = (((!g319) & (!g358) & (g1467) & (g1468) & (g1473)) + ((!g319) & (g358) & (g1467) & (!g1468) & (g1473)) + ((!g319) & (g358) & (g1467) & (g1468) & (!g1473)) + ((!g319) & (g358) & (g1467) & (g1468) & (g1473)) + ((g319) & (!g358) & (!g1467) & (g1468) & (g1473)) + ((g319) & (!g358) & (g1467) & (!g1468) & (!g1473)) + ((g319) & (!g358) & (g1467) & (!g1468) & (g1473)) + ((g319) & (!g358) & (g1467) & (g1468) & (!g1473)) + ((g319) & (!g358) & (g1467) & (g1468) & (g1473)) + ((g319) & (g358) & (!g1467) & (!g1468) & (g1473)) + ((g319) & (g358) & (!g1467) & (g1468) & (!g1473)) + ((g319) & (g358) & (!g1467) & (g1468) & (g1473)) + ((g319) & (g358) & (g1467) & (!g1468) & (!g1473)) + ((g319) & (g358) & (g1467) & (!g1468) & (g1473)) + ((g319) & (g358) & (g1467) & (g1468) & (!g1473)) + ((g319) & (g358) & (g1467) & (g1468) & (g1473)));
	assign g1475 = (((!g255) & (!g290) & (g1465) & (g1466) & (g1474)) + ((!g255) & (g290) & (g1465) & (!g1466) & (g1474)) + ((!g255) & (g290) & (g1465) & (g1466) & (!g1474)) + ((!g255) & (g290) & (g1465) & (g1466) & (g1474)) + ((g255) & (!g290) & (!g1465) & (g1466) & (g1474)) + ((g255) & (!g290) & (g1465) & (!g1466) & (!g1474)) + ((g255) & (!g290) & (g1465) & (!g1466) & (g1474)) + ((g255) & (!g290) & (g1465) & (g1466) & (!g1474)) + ((g255) & (!g290) & (g1465) & (g1466) & (g1474)) + ((g255) & (g290) & (!g1465) & (!g1466) & (g1474)) + ((g255) & (g290) & (!g1465) & (g1466) & (!g1474)) + ((g255) & (g290) & (!g1465) & (g1466) & (g1474)) + ((g255) & (g290) & (g1465) & (!g1466) & (!g1474)) + ((g255) & (g290) & (g1465) & (!g1466) & (g1474)) + ((g255) & (g290) & (g1465) & (g1466) & (!g1474)) + ((g255) & (g290) & (g1465) & (g1466) & (g1474)));
	assign g1476 = (((!g198) & (!g229) & (g1463) & (g1464) & (g1475)) + ((!g198) & (g229) & (g1463) & (!g1464) & (g1475)) + ((!g198) & (g229) & (g1463) & (g1464) & (!g1475)) + ((!g198) & (g229) & (g1463) & (g1464) & (g1475)) + ((g198) & (!g229) & (!g1463) & (g1464) & (g1475)) + ((g198) & (!g229) & (g1463) & (!g1464) & (!g1475)) + ((g198) & (!g229) & (g1463) & (!g1464) & (g1475)) + ((g198) & (!g229) & (g1463) & (g1464) & (!g1475)) + ((g198) & (!g229) & (g1463) & (g1464) & (g1475)) + ((g198) & (g229) & (!g1463) & (!g1464) & (g1475)) + ((g198) & (g229) & (!g1463) & (g1464) & (!g1475)) + ((g198) & (g229) & (!g1463) & (g1464) & (g1475)) + ((g198) & (g229) & (g1463) & (!g1464) & (!g1475)) + ((g198) & (g229) & (g1463) & (!g1464) & (g1475)) + ((g198) & (g229) & (g1463) & (g1464) & (!g1475)) + ((g198) & (g229) & (g1463) & (g1464) & (g1475)));
	assign g1477 = (((!g147) & (!g174) & (g1461) & (g1462) & (g1476)) + ((!g147) & (g174) & (g1461) & (!g1462) & (g1476)) + ((!g147) & (g174) & (g1461) & (g1462) & (!g1476)) + ((!g147) & (g174) & (g1461) & (g1462) & (g1476)) + ((g147) & (!g174) & (!g1461) & (g1462) & (g1476)) + ((g147) & (!g174) & (g1461) & (!g1462) & (!g1476)) + ((g147) & (!g174) & (g1461) & (!g1462) & (g1476)) + ((g147) & (!g174) & (g1461) & (g1462) & (!g1476)) + ((g147) & (!g174) & (g1461) & (g1462) & (g1476)) + ((g147) & (g174) & (!g1461) & (!g1462) & (g1476)) + ((g147) & (g174) & (!g1461) & (g1462) & (!g1476)) + ((g147) & (g174) & (!g1461) & (g1462) & (g1476)) + ((g147) & (g174) & (g1461) & (!g1462) & (!g1476)) + ((g147) & (g174) & (g1461) & (!g1462) & (g1476)) + ((g147) & (g174) & (g1461) & (g1462) & (!g1476)) + ((g147) & (g174) & (g1461) & (g1462) & (g1476)));
	assign g1478 = (((!g104) & (!g127) & (g1459) & (g1460) & (g1477)) + ((!g104) & (g127) & (g1459) & (!g1460) & (g1477)) + ((!g104) & (g127) & (g1459) & (g1460) & (!g1477)) + ((!g104) & (g127) & (g1459) & (g1460) & (g1477)) + ((g104) & (!g127) & (!g1459) & (g1460) & (g1477)) + ((g104) & (!g127) & (g1459) & (!g1460) & (!g1477)) + ((g104) & (!g127) & (g1459) & (!g1460) & (g1477)) + ((g104) & (!g127) & (g1459) & (g1460) & (!g1477)) + ((g104) & (!g127) & (g1459) & (g1460) & (g1477)) + ((g104) & (g127) & (!g1459) & (!g1460) & (g1477)) + ((g104) & (g127) & (!g1459) & (g1460) & (!g1477)) + ((g104) & (g127) & (!g1459) & (g1460) & (g1477)) + ((g104) & (g127) & (g1459) & (!g1460) & (!g1477)) + ((g104) & (g127) & (g1459) & (!g1460) & (g1477)) + ((g104) & (g127) & (g1459) & (g1460) & (!g1477)) + ((g104) & (g127) & (g1459) & (g1460) & (g1477)));
	assign g1479 = (((!g68) & (!g87) & (g1457) & (g1458) & (g1478)) + ((!g68) & (g87) & (g1457) & (!g1458) & (g1478)) + ((!g68) & (g87) & (g1457) & (g1458) & (!g1478)) + ((!g68) & (g87) & (g1457) & (g1458) & (g1478)) + ((g68) & (!g87) & (!g1457) & (g1458) & (g1478)) + ((g68) & (!g87) & (g1457) & (!g1458) & (!g1478)) + ((g68) & (!g87) & (g1457) & (!g1458) & (g1478)) + ((g68) & (!g87) & (g1457) & (g1458) & (!g1478)) + ((g68) & (!g87) & (g1457) & (g1458) & (g1478)) + ((g68) & (g87) & (!g1457) & (!g1458) & (g1478)) + ((g68) & (g87) & (!g1457) & (g1458) & (!g1478)) + ((g68) & (g87) & (!g1457) & (g1458) & (g1478)) + ((g68) & (g87) & (g1457) & (!g1458) & (!g1478)) + ((g68) & (g87) & (g1457) & (!g1458) & (g1478)) + ((g68) & (g87) & (g1457) & (g1458) & (!g1478)) + ((g68) & (g87) & (g1457) & (g1458) & (g1478)));
	assign g1480 = (((!g39) & (!g54) & (g1455) & (g1456) & (g1479)) + ((!g39) & (g54) & (g1455) & (!g1456) & (g1479)) + ((!g39) & (g54) & (g1455) & (g1456) & (!g1479)) + ((!g39) & (g54) & (g1455) & (g1456) & (g1479)) + ((g39) & (!g54) & (!g1455) & (g1456) & (g1479)) + ((g39) & (!g54) & (g1455) & (!g1456) & (!g1479)) + ((g39) & (!g54) & (g1455) & (!g1456) & (g1479)) + ((g39) & (!g54) & (g1455) & (g1456) & (!g1479)) + ((g39) & (!g54) & (g1455) & (g1456) & (g1479)) + ((g39) & (g54) & (!g1455) & (!g1456) & (g1479)) + ((g39) & (g54) & (!g1455) & (g1456) & (!g1479)) + ((g39) & (g54) & (!g1455) & (g1456) & (g1479)) + ((g39) & (g54) & (g1455) & (!g1456) & (!g1479)) + ((g39) & (g54) & (g1455) & (!g1456) & (g1479)) + ((g39) & (g54) & (g1455) & (g1456) & (!g1479)) + ((g39) & (g54) & (g1455) & (g1456) & (g1479)));
	assign g1481 = (((!g18) & (!g27) & (g1453) & (g1454) & (g1480)) + ((!g18) & (g27) & (g1453) & (!g1454) & (g1480)) + ((!g18) & (g27) & (g1453) & (g1454) & (!g1480)) + ((!g18) & (g27) & (g1453) & (g1454) & (g1480)) + ((g18) & (!g27) & (!g1453) & (g1454) & (g1480)) + ((g18) & (!g27) & (g1453) & (!g1454) & (!g1480)) + ((g18) & (!g27) & (g1453) & (!g1454) & (g1480)) + ((g18) & (!g27) & (g1453) & (g1454) & (!g1480)) + ((g18) & (!g27) & (g1453) & (g1454) & (g1480)) + ((g18) & (g27) & (!g1453) & (!g1454) & (g1480)) + ((g18) & (g27) & (!g1453) & (g1454) & (!g1480)) + ((g18) & (g27) & (!g1453) & (g1454) & (g1480)) + ((g18) & (g27) & (g1453) & (!g1454) & (!g1480)) + ((g18) & (g27) & (g1453) & (!g1454) & (g1480)) + ((g18) & (g27) & (g1453) & (g1454) & (!g1480)) + ((g18) & (g27) & (g1453) & (g1454) & (g1480)));
	assign g1482 = (((!g2) & (!g8) & (g1451) & (g1452) & (g1481)) + ((!g2) & (g8) & (g1451) & (!g1452) & (g1481)) + ((!g2) & (g8) & (g1451) & (g1452) & (!g1481)) + ((!g2) & (g8) & (g1451) & (g1452) & (g1481)) + ((g2) & (!g8) & (!g1451) & (g1452) & (g1481)) + ((g2) & (!g8) & (g1451) & (!g1452) & (!g1481)) + ((g2) & (!g8) & (g1451) & (!g1452) & (g1481)) + ((g2) & (!g8) & (g1451) & (g1452) & (!g1481)) + ((g2) & (!g8) & (g1451) & (g1452) & (g1481)) + ((g2) & (g8) & (!g1451) & (!g1452) & (g1481)) + ((g2) & (g8) & (!g1451) & (g1452) & (!g1481)) + ((g2) & (g8) & (!g1451) & (g1452) & (g1481)) + ((g2) & (g8) & (g1451) & (!g1452) & (!g1481)) + ((g2) & (g8) & (g1451) & (!g1452) & (g1481)) + ((g2) & (g8) & (g1451) & (g1452) & (!g1481)) + ((g2) & (g8) & (g1451) & (g1452) & (g1481)));
	assign g1483 = (((!g2) & (!g1373) & (g1416) & (!g1423)) + ((!g2) & (g1373) & (!g1416) & (!g1423)) + ((!g2) & (g1373) & (!g1416) & (g1423)) + ((!g2) & (g1373) & (g1416) & (g1423)) + ((g2) & (!g1373) & (!g1416) & (!g1423)) + ((g2) & (g1373) & (!g1416) & (g1423)) + ((g2) & (g1373) & (g1416) & (!g1423)) + ((g2) & (g1373) & (g1416) & (g1423)));
	assign g1484 = (((!g1) & (!g1372) & (!g1419) & (!g1421) & (g1422)) + ((!g1) & (!g1372) & (!g1419) & (g1421) & (!g1422)) + ((!g1) & (!g1372) & (!g1419) & (g1421) & (g1422)) + ((!g1) & (g1372) & (g1419) & (!g1421) & (!g1422)) + ((!g1) & (g1372) & (g1419) & (!g1421) & (g1422)) + ((!g1) & (g1372) & (g1419) & (g1421) & (!g1422)) + ((!g1) & (g1372) & (g1419) & (g1421) & (g1422)) + ((g1) & (!g1372) & (!g1419) & (!g1421) & (g1422)) + ((g1) & (!g1372) & (!g1419) & (g1421) & (g1422)) + ((g1) & (g1372) & (g1419) & (!g1421) & (!g1422)) + ((g1) & (g1372) & (g1419) & (!g1421) & (g1422)) + ((g1) & (g1372) & (g1419) & (g1421) & (!g1422)) + ((g1) & (g1372) & (g1419) & (g1421) & (g1422)));
	assign g1485 = (((!g4) & (!g1) & (!g1450) & (!g1482) & (!g1483) & (!g1484)) + ((!g4) & (g1) & (!g1450) & (!g1482) & (!g1483) & (!g1484)) + ((!g4) & (g1) & (!g1450) & (!g1482) & (!g1483) & (g1484)) + ((!g4) & (g1) & (!g1450) & (!g1482) & (g1483) & (!g1484)) + ((!g4) & (g1) & (!g1450) & (!g1482) & (g1483) & (g1484)) + ((!g4) & (g1) & (!g1450) & (g1482) & (!g1483) & (!g1484)) + ((!g4) & (g1) & (!g1450) & (g1482) & (!g1483) & (g1484)) + ((!g4) & (g1) & (!g1450) & (g1482) & (g1483) & (!g1484)) + ((!g4) & (g1) & (!g1450) & (g1482) & (g1483) & (g1484)) + ((!g4) & (g1) & (g1450) & (!g1482) & (!g1483) & (!g1484)) + ((!g4) & (g1) & (g1450) & (!g1482) & (!g1483) & (g1484)) + ((g4) & (!g1) & (!g1450) & (!g1482) & (!g1483) & (!g1484)) + ((g4) & (!g1) & (!g1450) & (!g1482) & (g1483) & (!g1484)) + ((g4) & (!g1) & (!g1450) & (g1482) & (!g1483) & (!g1484)) + ((g4) & (g1) & (!g1450) & (!g1482) & (!g1483) & (!g1484)) + ((g4) & (g1) & (!g1450) & (!g1482) & (!g1483) & (g1484)) + ((g4) & (g1) & (!g1450) & (!g1482) & (g1483) & (!g1484)) + ((g4) & (g1) & (!g1450) & (!g1482) & (g1483) & (g1484)) + ((g4) & (g1) & (!g1450) & (g1482) & (!g1483) & (!g1484)) + ((g4) & (g1) & (!g1450) & (g1482) & (!g1483) & (g1484)) + ((g4) & (g1) & (!g1450) & (g1482) & (g1483) & (!g1484)) + ((g4) & (g1) & (!g1450) & (g1482) & (g1483) & (g1484)) + ((g4) & (g1) & (g1450) & (!g1482) & (!g1483) & (!g1484)) + ((g4) & (g1) & (g1450) & (!g1482) & (!g1483) & (g1484)) + ((g4) & (g1) & (g1450) & (!g1482) & (g1483) & (!g1484)) + ((g4) & (g1) & (g1450) & (!g1482) & (g1483) & (g1484)) + ((g4) & (g1) & (g1450) & (g1482) & (!g1483) & (!g1484)) + ((g4) & (g1) & (g1450) & (g1482) & (!g1483) & (g1484)));
	assign g1486 = (((!g515) & (!g1424) & (g1448) & (!g1449) & (!g1485)) + ((!g515) & (!g1424) & (g1448) & (g1449) & (!g1485)) + ((!g515) & (!g1424) & (g1448) & (g1449) & (g1485)) + ((!g515) & (g1424) & (!g1448) & (!g1449) & (!g1485)) + ((!g515) & (g1424) & (!g1448) & (!g1449) & (g1485)) + ((!g515) & (g1424) & (!g1448) & (g1449) & (!g1485)) + ((!g515) & (g1424) & (!g1448) & (g1449) & (g1485)) + ((!g515) & (g1424) & (g1448) & (!g1449) & (g1485)) + ((g515) & (!g1424) & (!g1448) & (!g1449) & (!g1485)) + ((g515) & (!g1424) & (!g1448) & (g1449) & (!g1485)) + ((g515) & (!g1424) & (!g1448) & (g1449) & (g1485)) + ((g515) & (g1424) & (!g1448) & (!g1449) & (g1485)) + ((g515) & (g1424) & (g1448) & (!g1449) & (!g1485)) + ((g515) & (g1424) & (g1448) & (!g1449) & (g1485)) + ((g515) & (g1424) & (g1448) & (g1449) & (!g1485)) + ((g515) & (g1424) & (g1448) & (g1449) & (g1485)));
	assign g1487 = (((!g553) & (!g604) & (g1426) & (g1447)) + ((!g553) & (g604) & (!g1426) & (g1447)) + ((!g553) & (g604) & (g1426) & (!g1447)) + ((!g553) & (g604) & (g1426) & (g1447)) + ((g553) & (!g604) & (!g1426) & (!g1447)) + ((g553) & (!g604) & (!g1426) & (g1447)) + ((g553) & (!g604) & (g1426) & (!g1447)) + ((g553) & (g604) & (!g1426) & (!g1447)));
	assign g1488 = (((!g1425) & (!g1449) & (!g1485) & (g1487)) + ((!g1425) & (g1449) & (!g1485) & (g1487)) + ((!g1425) & (g1449) & (g1485) & (g1487)) + ((g1425) & (!g1449) & (!g1485) & (!g1487)) + ((g1425) & (!g1449) & (g1485) & (!g1487)) + ((g1425) & (!g1449) & (g1485) & (g1487)) + ((g1425) & (g1449) & (!g1485) & (!g1487)) + ((g1425) & (g1449) & (g1485) & (!g1487)));
	assign g1489 = (((!g604) & (!g1426) & (g1447) & (!g1449) & (!g1485)) + ((!g604) & (!g1426) & (g1447) & (g1449) & (!g1485)) + ((!g604) & (!g1426) & (g1447) & (g1449) & (g1485)) + ((!g604) & (g1426) & (!g1447) & (!g1449) & (!g1485)) + ((!g604) & (g1426) & (!g1447) & (!g1449) & (g1485)) + ((!g604) & (g1426) & (!g1447) & (g1449) & (!g1485)) + ((!g604) & (g1426) & (!g1447) & (g1449) & (g1485)) + ((!g604) & (g1426) & (g1447) & (!g1449) & (g1485)) + ((g604) & (!g1426) & (!g1447) & (!g1449) & (!g1485)) + ((g604) & (!g1426) & (!g1447) & (g1449) & (!g1485)) + ((g604) & (!g1426) & (!g1447) & (g1449) & (g1485)) + ((g604) & (g1426) & (!g1447) & (!g1449) & (g1485)) + ((g604) & (g1426) & (g1447) & (!g1449) & (!g1485)) + ((g604) & (g1426) & (g1447) & (!g1449) & (g1485)) + ((g604) & (g1426) & (g1447) & (g1449) & (!g1485)) + ((g604) & (g1426) & (g1447) & (g1449) & (g1485)));
	assign g1490 = (((!g645) & (!g700) & (g1428) & (g1446)) + ((!g645) & (g700) & (!g1428) & (g1446)) + ((!g645) & (g700) & (g1428) & (!g1446)) + ((!g645) & (g700) & (g1428) & (g1446)) + ((g645) & (!g700) & (!g1428) & (!g1446)) + ((g645) & (!g700) & (!g1428) & (g1446)) + ((g645) & (!g700) & (g1428) & (!g1446)) + ((g645) & (g700) & (!g1428) & (!g1446)));
	assign g1491 = (((!g1427) & (!g1449) & (!g1485) & (g1490)) + ((!g1427) & (g1449) & (!g1485) & (g1490)) + ((!g1427) & (g1449) & (g1485) & (g1490)) + ((g1427) & (!g1449) & (!g1485) & (!g1490)) + ((g1427) & (!g1449) & (g1485) & (!g1490)) + ((g1427) & (!g1449) & (g1485) & (g1490)) + ((g1427) & (g1449) & (!g1485) & (!g1490)) + ((g1427) & (g1449) & (g1485) & (!g1490)));
	assign g1492 = (((!g700) & (!g1428) & (g1446) & (!g1449) & (!g1485)) + ((!g700) & (!g1428) & (g1446) & (g1449) & (!g1485)) + ((!g700) & (!g1428) & (g1446) & (g1449) & (g1485)) + ((!g700) & (g1428) & (!g1446) & (!g1449) & (!g1485)) + ((!g700) & (g1428) & (!g1446) & (!g1449) & (g1485)) + ((!g700) & (g1428) & (!g1446) & (g1449) & (!g1485)) + ((!g700) & (g1428) & (!g1446) & (g1449) & (g1485)) + ((!g700) & (g1428) & (g1446) & (!g1449) & (g1485)) + ((g700) & (!g1428) & (!g1446) & (!g1449) & (!g1485)) + ((g700) & (!g1428) & (!g1446) & (g1449) & (!g1485)) + ((g700) & (!g1428) & (!g1446) & (g1449) & (g1485)) + ((g700) & (g1428) & (!g1446) & (!g1449) & (g1485)) + ((g700) & (g1428) & (g1446) & (!g1449) & (!g1485)) + ((g700) & (g1428) & (g1446) & (!g1449) & (g1485)) + ((g700) & (g1428) & (g1446) & (g1449) & (!g1485)) + ((g700) & (g1428) & (g1446) & (g1449) & (g1485)));
	assign g1493 = (((!g744) & (!g803) & (g1430) & (g1445)) + ((!g744) & (g803) & (!g1430) & (g1445)) + ((!g744) & (g803) & (g1430) & (!g1445)) + ((!g744) & (g803) & (g1430) & (g1445)) + ((g744) & (!g803) & (!g1430) & (!g1445)) + ((g744) & (!g803) & (!g1430) & (g1445)) + ((g744) & (!g803) & (g1430) & (!g1445)) + ((g744) & (g803) & (!g1430) & (!g1445)));
	assign g1494 = (((!g1429) & (!g1449) & (!g1485) & (g1493)) + ((!g1429) & (g1449) & (!g1485) & (g1493)) + ((!g1429) & (g1449) & (g1485) & (g1493)) + ((g1429) & (!g1449) & (!g1485) & (!g1493)) + ((g1429) & (!g1449) & (g1485) & (!g1493)) + ((g1429) & (!g1449) & (g1485) & (g1493)) + ((g1429) & (g1449) & (!g1485) & (!g1493)) + ((g1429) & (g1449) & (g1485) & (!g1493)));
	assign g1495 = (((!g803) & (!g1430) & (g1445) & (!g1449) & (!g1485)) + ((!g803) & (!g1430) & (g1445) & (g1449) & (!g1485)) + ((!g803) & (!g1430) & (g1445) & (g1449) & (g1485)) + ((!g803) & (g1430) & (!g1445) & (!g1449) & (!g1485)) + ((!g803) & (g1430) & (!g1445) & (!g1449) & (g1485)) + ((!g803) & (g1430) & (!g1445) & (g1449) & (!g1485)) + ((!g803) & (g1430) & (!g1445) & (g1449) & (g1485)) + ((!g803) & (g1430) & (g1445) & (!g1449) & (g1485)) + ((g803) & (!g1430) & (!g1445) & (!g1449) & (!g1485)) + ((g803) & (!g1430) & (!g1445) & (g1449) & (!g1485)) + ((g803) & (!g1430) & (!g1445) & (g1449) & (g1485)) + ((g803) & (g1430) & (!g1445) & (!g1449) & (g1485)) + ((g803) & (g1430) & (g1445) & (!g1449) & (!g1485)) + ((g803) & (g1430) & (g1445) & (!g1449) & (g1485)) + ((g803) & (g1430) & (g1445) & (g1449) & (!g1485)) + ((g803) & (g1430) & (g1445) & (g1449) & (g1485)));
	assign g1496 = (((!g851) & (!g914) & (g1432) & (g1444)) + ((!g851) & (g914) & (!g1432) & (g1444)) + ((!g851) & (g914) & (g1432) & (!g1444)) + ((!g851) & (g914) & (g1432) & (g1444)) + ((g851) & (!g914) & (!g1432) & (!g1444)) + ((g851) & (!g914) & (!g1432) & (g1444)) + ((g851) & (!g914) & (g1432) & (!g1444)) + ((g851) & (g914) & (!g1432) & (!g1444)));
	assign g1497 = (((!g1431) & (!g1449) & (!g1485) & (g1496)) + ((!g1431) & (g1449) & (!g1485) & (g1496)) + ((!g1431) & (g1449) & (g1485) & (g1496)) + ((g1431) & (!g1449) & (!g1485) & (!g1496)) + ((g1431) & (!g1449) & (g1485) & (!g1496)) + ((g1431) & (!g1449) & (g1485) & (g1496)) + ((g1431) & (g1449) & (!g1485) & (!g1496)) + ((g1431) & (g1449) & (g1485) & (!g1496)));
	assign g1498 = (((!g914) & (!g1432) & (g1444) & (!g1449) & (!g1485)) + ((!g914) & (!g1432) & (g1444) & (g1449) & (!g1485)) + ((!g914) & (!g1432) & (g1444) & (g1449) & (g1485)) + ((!g914) & (g1432) & (!g1444) & (!g1449) & (!g1485)) + ((!g914) & (g1432) & (!g1444) & (!g1449) & (g1485)) + ((!g914) & (g1432) & (!g1444) & (g1449) & (!g1485)) + ((!g914) & (g1432) & (!g1444) & (g1449) & (g1485)) + ((!g914) & (g1432) & (g1444) & (!g1449) & (g1485)) + ((g914) & (!g1432) & (!g1444) & (!g1449) & (!g1485)) + ((g914) & (!g1432) & (!g1444) & (g1449) & (!g1485)) + ((g914) & (!g1432) & (!g1444) & (g1449) & (g1485)) + ((g914) & (g1432) & (!g1444) & (!g1449) & (g1485)) + ((g914) & (g1432) & (g1444) & (!g1449) & (!g1485)) + ((g914) & (g1432) & (g1444) & (!g1449) & (g1485)) + ((g914) & (g1432) & (g1444) & (g1449) & (!g1485)) + ((g914) & (g1432) & (g1444) & (g1449) & (g1485)));
	assign g1499 = (((!g1032) & (!g1030) & (g1434) & (g1443)) + ((!g1032) & (g1030) & (!g1434) & (g1443)) + ((!g1032) & (g1030) & (g1434) & (!g1443)) + ((!g1032) & (g1030) & (g1434) & (g1443)) + ((g1032) & (!g1030) & (!g1434) & (!g1443)) + ((g1032) & (!g1030) & (!g1434) & (g1443)) + ((g1032) & (!g1030) & (g1434) & (!g1443)) + ((g1032) & (g1030) & (!g1434) & (!g1443)));
	assign g1500 = (((!g1433) & (!g1449) & (!g1485) & (g1499)) + ((!g1433) & (g1449) & (!g1485) & (g1499)) + ((!g1433) & (g1449) & (g1485) & (g1499)) + ((g1433) & (!g1449) & (!g1485) & (!g1499)) + ((g1433) & (!g1449) & (g1485) & (!g1499)) + ((g1433) & (!g1449) & (g1485) & (g1499)) + ((g1433) & (g1449) & (!g1485) & (!g1499)) + ((g1433) & (g1449) & (g1485) & (!g1499)));
	assign g1501 = (((!g1030) & (!g1434) & (g1443) & (!g1449) & (!g1485)) + ((!g1030) & (!g1434) & (g1443) & (g1449) & (!g1485)) + ((!g1030) & (!g1434) & (g1443) & (g1449) & (g1485)) + ((!g1030) & (g1434) & (!g1443) & (!g1449) & (!g1485)) + ((!g1030) & (g1434) & (!g1443) & (!g1449) & (g1485)) + ((!g1030) & (g1434) & (!g1443) & (g1449) & (!g1485)) + ((!g1030) & (g1434) & (!g1443) & (g1449) & (g1485)) + ((!g1030) & (g1434) & (g1443) & (!g1449) & (g1485)) + ((g1030) & (!g1434) & (!g1443) & (!g1449) & (!g1485)) + ((g1030) & (!g1434) & (!g1443) & (g1449) & (!g1485)) + ((g1030) & (!g1434) & (!g1443) & (g1449) & (g1485)) + ((g1030) & (g1434) & (!g1443) & (!g1449) & (g1485)) + ((g1030) & (g1434) & (g1443) & (!g1449) & (!g1485)) + ((g1030) & (g1434) & (g1443) & (!g1449) & (g1485)) + ((g1030) & (g1434) & (g1443) & (g1449) & (!g1485)) + ((g1030) & (g1434) & (g1443) & (g1449) & (g1485)));
	assign g1502 = (((!g1160) & (!g1154) & (g1436) & (g1442)) + ((!g1160) & (g1154) & (!g1436) & (g1442)) + ((!g1160) & (g1154) & (g1436) & (!g1442)) + ((!g1160) & (g1154) & (g1436) & (g1442)) + ((g1160) & (!g1154) & (!g1436) & (!g1442)) + ((g1160) & (!g1154) & (!g1436) & (g1442)) + ((g1160) & (!g1154) & (g1436) & (!g1442)) + ((g1160) & (g1154) & (!g1436) & (!g1442)));
	assign g1503 = (((!g1435) & (!g1449) & (!g1485) & (g1502)) + ((!g1435) & (g1449) & (!g1485) & (g1502)) + ((!g1435) & (g1449) & (g1485) & (g1502)) + ((g1435) & (!g1449) & (!g1485) & (!g1502)) + ((g1435) & (!g1449) & (g1485) & (!g1502)) + ((g1435) & (!g1449) & (g1485) & (g1502)) + ((g1435) & (g1449) & (!g1485) & (!g1502)) + ((g1435) & (g1449) & (g1485) & (!g1502)));
	assign g1504 = (((!g1154) & (!g1436) & (g1442) & (!g1449) & (!g1485)) + ((!g1154) & (!g1436) & (g1442) & (g1449) & (!g1485)) + ((!g1154) & (!g1436) & (g1442) & (g1449) & (g1485)) + ((!g1154) & (g1436) & (!g1442) & (!g1449) & (!g1485)) + ((!g1154) & (g1436) & (!g1442) & (!g1449) & (g1485)) + ((!g1154) & (g1436) & (!g1442) & (g1449) & (!g1485)) + ((!g1154) & (g1436) & (!g1442) & (g1449) & (g1485)) + ((!g1154) & (g1436) & (g1442) & (!g1449) & (g1485)) + ((g1154) & (!g1436) & (!g1442) & (!g1449) & (!g1485)) + ((g1154) & (!g1436) & (!g1442) & (g1449) & (!g1485)) + ((g1154) & (!g1436) & (!g1442) & (g1449) & (g1485)) + ((g1154) & (g1436) & (!g1442) & (!g1449) & (g1485)) + ((g1154) & (g1436) & (g1442) & (!g1449) & (!g1485)) + ((g1154) & (g1436) & (g1442) & (!g1449) & (g1485)) + ((g1154) & (g1436) & (g1442) & (g1449) & (!g1485)) + ((g1154) & (g1436) & (g1442) & (g1449) & (g1485)));
	assign g1505 = (((!g1295) & (!g1285) & (g1439) & (g1441)) + ((!g1295) & (g1285) & (!g1439) & (g1441)) + ((!g1295) & (g1285) & (g1439) & (!g1441)) + ((!g1295) & (g1285) & (g1439) & (g1441)) + ((g1295) & (!g1285) & (!g1439) & (!g1441)) + ((g1295) & (!g1285) & (!g1439) & (g1441)) + ((g1295) & (!g1285) & (g1439) & (!g1441)) + ((g1295) & (g1285) & (!g1439) & (!g1441)));
	assign g1506 = (((!g1438) & (!g1449) & (!g1485) & (g1505)) + ((!g1438) & (g1449) & (!g1485) & (g1505)) + ((!g1438) & (g1449) & (g1485) & (g1505)) + ((g1438) & (!g1449) & (!g1485) & (!g1505)) + ((g1438) & (!g1449) & (g1485) & (!g1505)) + ((g1438) & (!g1449) & (g1485) & (g1505)) + ((g1438) & (g1449) & (!g1485) & (!g1505)) + ((g1438) & (g1449) & (g1485) & (!g1505)));
	assign g1507 = (((!g1285) & (!g1439) & (g1441) & (!g1449) & (!g1485)) + ((!g1285) & (!g1439) & (g1441) & (g1449) & (!g1485)) + ((!g1285) & (!g1439) & (g1441) & (g1449) & (g1485)) + ((!g1285) & (g1439) & (!g1441) & (!g1449) & (!g1485)) + ((!g1285) & (g1439) & (!g1441) & (!g1449) & (g1485)) + ((!g1285) & (g1439) & (!g1441) & (g1449) & (!g1485)) + ((!g1285) & (g1439) & (!g1441) & (g1449) & (g1485)) + ((!g1285) & (g1439) & (g1441) & (!g1449) & (g1485)) + ((g1285) & (!g1439) & (!g1441) & (!g1449) & (!g1485)) + ((g1285) & (!g1439) & (!g1441) & (g1449) & (!g1485)) + ((g1285) & (!g1439) & (!g1441) & (g1449) & (g1485)) + ((g1285) & (g1439) & (!g1441) & (!g1449) & (g1485)) + ((g1285) & (g1439) & (g1441) & (!g1449) & (!g1485)) + ((g1285) & (g1439) & (g1441) & (!g1449) & (g1485)) + ((g1285) & (g1439) & (g1441) & (g1449) & (!g1485)) + ((g1285) & (g1439) & (g1441) & (g1449) & (g1485)));
	assign g1508 = (((!g1437) & (!ax48x) & (!g1423) & (g1440)) + ((!g1437) & (!ax48x) & (g1423) & (g1440)) + ((!g1437) & (ax48x) & (!g1423) & (!g1440)) + ((!g1437) & (ax48x) & (!g1423) & (g1440)) + ((g1437) & (!ax48x) & (!g1423) & (!g1440)) + ((g1437) & (!ax48x) & (g1423) & (!g1440)) + ((g1437) & (ax48x) & (g1423) & (!g1440)) + ((g1437) & (ax48x) & (g1423) & (g1440)));
	assign g1509 = (((!ax48x) & (!ax49x) & (!g1423) & (!g1449) & (!g1485) & (g1508)) + ((!ax48x) & (!ax49x) & (!g1423) & (!g1449) & (g1485) & (!g1508)) + ((!ax48x) & (!ax49x) & (!g1423) & (!g1449) & (g1485) & (g1508)) + ((!ax48x) & (!ax49x) & (!g1423) & (g1449) & (!g1485) & (g1508)) + ((!ax48x) & (!ax49x) & (!g1423) & (g1449) & (g1485) & (g1508)) + ((!ax48x) & (!ax49x) & (g1423) & (!g1449) & (!g1485) & (!g1508)) + ((!ax48x) & (!ax49x) & (g1423) & (g1449) & (!g1485) & (!g1508)) + ((!ax48x) & (!ax49x) & (g1423) & (g1449) & (g1485) & (!g1508)) + ((!ax48x) & (ax49x) & (!g1423) & (!g1449) & (!g1485) & (!g1508)) + ((!ax48x) & (ax49x) & (!g1423) & (g1449) & (!g1485) & (!g1508)) + ((!ax48x) & (ax49x) & (!g1423) & (g1449) & (g1485) & (!g1508)) + ((!ax48x) & (ax49x) & (g1423) & (!g1449) & (!g1485) & (g1508)) + ((!ax48x) & (ax49x) & (g1423) & (!g1449) & (g1485) & (!g1508)) + ((!ax48x) & (ax49x) & (g1423) & (!g1449) & (g1485) & (g1508)) + ((!ax48x) & (ax49x) & (g1423) & (g1449) & (!g1485) & (g1508)) + ((!ax48x) & (ax49x) & (g1423) & (g1449) & (g1485) & (g1508)) + ((ax48x) & (!ax49x) & (!g1423) & (!g1449) & (!g1485) & (!g1508)) + ((ax48x) & (!ax49x) & (!g1423) & (g1449) & (!g1485) & (!g1508)) + ((ax48x) & (!ax49x) & (!g1423) & (g1449) & (g1485) & (!g1508)) + ((ax48x) & (!ax49x) & (g1423) & (!g1449) & (!g1485) & (!g1508)) + ((ax48x) & (!ax49x) & (g1423) & (g1449) & (!g1485) & (!g1508)) + ((ax48x) & (!ax49x) & (g1423) & (g1449) & (g1485) & (!g1508)) + ((ax48x) & (ax49x) & (!g1423) & (!g1449) & (!g1485) & (g1508)) + ((ax48x) & (ax49x) & (!g1423) & (!g1449) & (g1485) & (!g1508)) + ((ax48x) & (ax49x) & (!g1423) & (!g1449) & (g1485) & (g1508)) + ((ax48x) & (ax49x) & (!g1423) & (g1449) & (!g1485) & (g1508)) + ((ax48x) & (ax49x) & (!g1423) & (g1449) & (g1485) & (g1508)) + ((ax48x) & (ax49x) & (g1423) & (!g1449) & (!g1485) & (g1508)) + ((ax48x) & (ax49x) & (g1423) & (!g1449) & (g1485) & (!g1508)) + ((ax48x) & (ax49x) & (g1423) & (!g1449) & (g1485) & (g1508)) + ((ax48x) & (ax49x) & (g1423) & (g1449) & (!g1485) & (g1508)) + ((ax48x) & (ax49x) & (g1423) & (g1449) & (g1485) & (g1508)));
	assign g1510 = (((!ax48x) & (!g1423) & (!g1440) & (!g1449) & (g1485)) + ((!ax48x) & (!g1423) & (g1440) & (!g1449) & (!g1485)) + ((!ax48x) & (!g1423) & (g1440) & (!g1449) & (g1485)) + ((!ax48x) & (!g1423) & (g1440) & (g1449) & (!g1485)) + ((!ax48x) & (!g1423) & (g1440) & (g1449) & (g1485)) + ((!ax48x) & (g1423) & (g1440) & (!g1449) & (!g1485)) + ((!ax48x) & (g1423) & (g1440) & (g1449) & (!g1485)) + ((!ax48x) & (g1423) & (g1440) & (g1449) & (g1485)) + ((ax48x) & (!g1423) & (!g1440) & (!g1449) & (!g1485)) + ((ax48x) & (!g1423) & (!g1440) & (g1449) & (!g1485)) + ((ax48x) & (!g1423) & (!g1440) & (g1449) & (g1485)) + ((ax48x) & (g1423) & (!g1440) & (!g1449) & (!g1485)) + ((ax48x) & (g1423) & (!g1440) & (!g1449) & (g1485)) + ((ax48x) & (g1423) & (!g1440) & (g1449) & (!g1485)) + ((ax48x) & (g1423) & (!g1440) & (g1449) & (g1485)) + ((ax48x) & (g1423) & (g1440) & (!g1449) & (g1485)));
	assign g1511 = (((!ax44x) & (!ax45x)));
	assign g1512 = (((!g1423) & (!ax46x) & (!ax47x) & (!g1449) & (!g1485) & (!g1511)) + ((!g1423) & (!ax46x) & (!ax47x) & (g1449) & (!g1485) & (!g1511)) + ((!g1423) & (!ax46x) & (!ax47x) & (g1449) & (g1485) & (!g1511)) + ((!g1423) & (!ax46x) & (ax47x) & (!g1449) & (g1485) & (!g1511)) + ((!g1423) & (ax46x) & (ax47x) & (!g1449) & (g1485) & (!g1511)) + ((!g1423) & (ax46x) & (ax47x) & (!g1449) & (g1485) & (g1511)) + ((g1423) & (!ax46x) & (!ax47x) & (!g1449) & (!g1485) & (!g1511)) + ((g1423) & (!ax46x) & (!ax47x) & (!g1449) & (!g1485) & (g1511)) + ((g1423) & (!ax46x) & (!ax47x) & (!g1449) & (g1485) & (!g1511)) + ((g1423) & (!ax46x) & (!ax47x) & (g1449) & (!g1485) & (!g1511)) + ((g1423) & (!ax46x) & (!ax47x) & (g1449) & (!g1485) & (g1511)) + ((g1423) & (!ax46x) & (!ax47x) & (g1449) & (g1485) & (!g1511)) + ((g1423) & (!ax46x) & (!ax47x) & (g1449) & (g1485) & (g1511)) + ((g1423) & (!ax46x) & (ax47x) & (!g1449) & (!g1485) & (!g1511)) + ((g1423) & (!ax46x) & (ax47x) & (!g1449) & (g1485) & (!g1511)) + ((g1423) & (!ax46x) & (ax47x) & (!g1449) & (g1485) & (g1511)) + ((g1423) & (!ax46x) & (ax47x) & (g1449) & (!g1485) & (!g1511)) + ((g1423) & (!ax46x) & (ax47x) & (g1449) & (g1485) & (!g1511)) + ((g1423) & (ax46x) & (!ax47x) & (!g1449) & (g1485) & (!g1511)) + ((g1423) & (ax46x) & (!ax47x) & (!g1449) & (g1485) & (g1511)) + ((g1423) & (ax46x) & (ax47x) & (!g1449) & (!g1485) & (!g1511)) + ((g1423) & (ax46x) & (ax47x) & (!g1449) & (!g1485) & (g1511)) + ((g1423) & (ax46x) & (ax47x) & (!g1449) & (g1485) & (!g1511)) + ((g1423) & (ax46x) & (ax47x) & (!g1449) & (g1485) & (g1511)) + ((g1423) & (ax46x) & (ax47x) & (g1449) & (!g1485) & (!g1511)) + ((g1423) & (ax46x) & (ax47x) & (g1449) & (!g1485) & (g1511)) + ((g1423) & (ax46x) & (ax47x) & (g1449) & (g1485) & (!g1511)) + ((g1423) & (ax46x) & (ax47x) & (g1449) & (g1485) & (g1511)));
	assign g1513 = (((!g1285) & (!g1437) & (g1509) & (g1510) & (g1512)) + ((!g1285) & (g1437) & (g1509) & (!g1510) & (g1512)) + ((!g1285) & (g1437) & (g1509) & (g1510) & (!g1512)) + ((!g1285) & (g1437) & (g1509) & (g1510) & (g1512)) + ((g1285) & (!g1437) & (!g1509) & (g1510) & (g1512)) + ((g1285) & (!g1437) & (g1509) & (!g1510) & (!g1512)) + ((g1285) & (!g1437) & (g1509) & (!g1510) & (g1512)) + ((g1285) & (!g1437) & (g1509) & (g1510) & (!g1512)) + ((g1285) & (!g1437) & (g1509) & (g1510) & (g1512)) + ((g1285) & (g1437) & (!g1509) & (!g1510) & (g1512)) + ((g1285) & (g1437) & (!g1509) & (g1510) & (!g1512)) + ((g1285) & (g1437) & (!g1509) & (g1510) & (g1512)) + ((g1285) & (g1437) & (g1509) & (!g1510) & (!g1512)) + ((g1285) & (g1437) & (g1509) & (!g1510) & (g1512)) + ((g1285) & (g1437) & (g1509) & (g1510) & (!g1512)) + ((g1285) & (g1437) & (g1509) & (g1510) & (g1512)));
	assign g1514 = (((!g1154) & (!g1295) & (g1506) & (g1507) & (g1513)) + ((!g1154) & (g1295) & (g1506) & (!g1507) & (g1513)) + ((!g1154) & (g1295) & (g1506) & (g1507) & (!g1513)) + ((!g1154) & (g1295) & (g1506) & (g1507) & (g1513)) + ((g1154) & (!g1295) & (!g1506) & (g1507) & (g1513)) + ((g1154) & (!g1295) & (g1506) & (!g1507) & (!g1513)) + ((g1154) & (!g1295) & (g1506) & (!g1507) & (g1513)) + ((g1154) & (!g1295) & (g1506) & (g1507) & (!g1513)) + ((g1154) & (!g1295) & (g1506) & (g1507) & (g1513)) + ((g1154) & (g1295) & (!g1506) & (!g1507) & (g1513)) + ((g1154) & (g1295) & (!g1506) & (g1507) & (!g1513)) + ((g1154) & (g1295) & (!g1506) & (g1507) & (g1513)) + ((g1154) & (g1295) & (g1506) & (!g1507) & (!g1513)) + ((g1154) & (g1295) & (g1506) & (!g1507) & (g1513)) + ((g1154) & (g1295) & (g1506) & (g1507) & (!g1513)) + ((g1154) & (g1295) & (g1506) & (g1507) & (g1513)));
	assign g1515 = (((!g1030) & (!g1160) & (g1503) & (g1504) & (g1514)) + ((!g1030) & (g1160) & (g1503) & (!g1504) & (g1514)) + ((!g1030) & (g1160) & (g1503) & (g1504) & (!g1514)) + ((!g1030) & (g1160) & (g1503) & (g1504) & (g1514)) + ((g1030) & (!g1160) & (!g1503) & (g1504) & (g1514)) + ((g1030) & (!g1160) & (g1503) & (!g1504) & (!g1514)) + ((g1030) & (!g1160) & (g1503) & (!g1504) & (g1514)) + ((g1030) & (!g1160) & (g1503) & (g1504) & (!g1514)) + ((g1030) & (!g1160) & (g1503) & (g1504) & (g1514)) + ((g1030) & (g1160) & (!g1503) & (!g1504) & (g1514)) + ((g1030) & (g1160) & (!g1503) & (g1504) & (!g1514)) + ((g1030) & (g1160) & (!g1503) & (g1504) & (g1514)) + ((g1030) & (g1160) & (g1503) & (!g1504) & (!g1514)) + ((g1030) & (g1160) & (g1503) & (!g1504) & (g1514)) + ((g1030) & (g1160) & (g1503) & (g1504) & (!g1514)) + ((g1030) & (g1160) & (g1503) & (g1504) & (g1514)));
	assign g1516 = (((!g914) & (!g1032) & (g1500) & (g1501) & (g1515)) + ((!g914) & (g1032) & (g1500) & (!g1501) & (g1515)) + ((!g914) & (g1032) & (g1500) & (g1501) & (!g1515)) + ((!g914) & (g1032) & (g1500) & (g1501) & (g1515)) + ((g914) & (!g1032) & (!g1500) & (g1501) & (g1515)) + ((g914) & (!g1032) & (g1500) & (!g1501) & (!g1515)) + ((g914) & (!g1032) & (g1500) & (!g1501) & (g1515)) + ((g914) & (!g1032) & (g1500) & (g1501) & (!g1515)) + ((g914) & (!g1032) & (g1500) & (g1501) & (g1515)) + ((g914) & (g1032) & (!g1500) & (!g1501) & (g1515)) + ((g914) & (g1032) & (!g1500) & (g1501) & (!g1515)) + ((g914) & (g1032) & (!g1500) & (g1501) & (g1515)) + ((g914) & (g1032) & (g1500) & (!g1501) & (!g1515)) + ((g914) & (g1032) & (g1500) & (!g1501) & (g1515)) + ((g914) & (g1032) & (g1500) & (g1501) & (!g1515)) + ((g914) & (g1032) & (g1500) & (g1501) & (g1515)));
	assign g1517 = (((!g803) & (!g851) & (g1497) & (g1498) & (g1516)) + ((!g803) & (g851) & (g1497) & (!g1498) & (g1516)) + ((!g803) & (g851) & (g1497) & (g1498) & (!g1516)) + ((!g803) & (g851) & (g1497) & (g1498) & (g1516)) + ((g803) & (!g851) & (!g1497) & (g1498) & (g1516)) + ((g803) & (!g851) & (g1497) & (!g1498) & (!g1516)) + ((g803) & (!g851) & (g1497) & (!g1498) & (g1516)) + ((g803) & (!g851) & (g1497) & (g1498) & (!g1516)) + ((g803) & (!g851) & (g1497) & (g1498) & (g1516)) + ((g803) & (g851) & (!g1497) & (!g1498) & (g1516)) + ((g803) & (g851) & (!g1497) & (g1498) & (!g1516)) + ((g803) & (g851) & (!g1497) & (g1498) & (g1516)) + ((g803) & (g851) & (g1497) & (!g1498) & (!g1516)) + ((g803) & (g851) & (g1497) & (!g1498) & (g1516)) + ((g803) & (g851) & (g1497) & (g1498) & (!g1516)) + ((g803) & (g851) & (g1497) & (g1498) & (g1516)));
	assign g1518 = (((!g700) & (!g744) & (g1494) & (g1495) & (g1517)) + ((!g700) & (g744) & (g1494) & (!g1495) & (g1517)) + ((!g700) & (g744) & (g1494) & (g1495) & (!g1517)) + ((!g700) & (g744) & (g1494) & (g1495) & (g1517)) + ((g700) & (!g744) & (!g1494) & (g1495) & (g1517)) + ((g700) & (!g744) & (g1494) & (!g1495) & (!g1517)) + ((g700) & (!g744) & (g1494) & (!g1495) & (g1517)) + ((g700) & (!g744) & (g1494) & (g1495) & (!g1517)) + ((g700) & (!g744) & (g1494) & (g1495) & (g1517)) + ((g700) & (g744) & (!g1494) & (!g1495) & (g1517)) + ((g700) & (g744) & (!g1494) & (g1495) & (!g1517)) + ((g700) & (g744) & (!g1494) & (g1495) & (g1517)) + ((g700) & (g744) & (g1494) & (!g1495) & (!g1517)) + ((g700) & (g744) & (g1494) & (!g1495) & (g1517)) + ((g700) & (g744) & (g1494) & (g1495) & (!g1517)) + ((g700) & (g744) & (g1494) & (g1495) & (g1517)));
	assign g1519 = (((!g604) & (!g645) & (g1491) & (g1492) & (g1518)) + ((!g604) & (g645) & (g1491) & (!g1492) & (g1518)) + ((!g604) & (g645) & (g1491) & (g1492) & (!g1518)) + ((!g604) & (g645) & (g1491) & (g1492) & (g1518)) + ((g604) & (!g645) & (!g1491) & (g1492) & (g1518)) + ((g604) & (!g645) & (g1491) & (!g1492) & (!g1518)) + ((g604) & (!g645) & (g1491) & (!g1492) & (g1518)) + ((g604) & (!g645) & (g1491) & (g1492) & (!g1518)) + ((g604) & (!g645) & (g1491) & (g1492) & (g1518)) + ((g604) & (g645) & (!g1491) & (!g1492) & (g1518)) + ((g604) & (g645) & (!g1491) & (g1492) & (!g1518)) + ((g604) & (g645) & (!g1491) & (g1492) & (g1518)) + ((g604) & (g645) & (g1491) & (!g1492) & (!g1518)) + ((g604) & (g645) & (g1491) & (!g1492) & (g1518)) + ((g604) & (g645) & (g1491) & (g1492) & (!g1518)) + ((g604) & (g645) & (g1491) & (g1492) & (g1518)));
	assign g1520 = (((!g515) & (!g553) & (g1488) & (g1489) & (g1519)) + ((!g515) & (g553) & (g1488) & (!g1489) & (g1519)) + ((!g515) & (g553) & (g1488) & (g1489) & (!g1519)) + ((!g515) & (g553) & (g1488) & (g1489) & (g1519)) + ((g515) & (!g553) & (!g1488) & (g1489) & (g1519)) + ((g515) & (!g553) & (g1488) & (!g1489) & (!g1519)) + ((g515) & (!g553) & (g1488) & (!g1489) & (g1519)) + ((g515) & (!g553) & (g1488) & (g1489) & (!g1519)) + ((g515) & (!g553) & (g1488) & (g1489) & (g1519)) + ((g515) & (g553) & (!g1488) & (!g1489) & (g1519)) + ((g515) & (g553) & (!g1488) & (g1489) & (!g1519)) + ((g515) & (g553) & (!g1488) & (g1489) & (g1519)) + ((g515) & (g553) & (g1488) & (!g1489) & (!g1519)) + ((g515) & (g553) & (g1488) & (!g1489) & (g1519)) + ((g515) & (g553) & (g1488) & (g1489) & (!g1519)) + ((g515) & (g553) & (g1488) & (g1489) & (g1519)));
	assign g1521 = (((!g4) & (!g1482) & (!g1483) & (!g1449) & (!g1485)) + ((!g4) & (!g1482) & (!g1483) & (g1449) & (!g1485)) + ((!g4) & (!g1482) & (!g1483) & (g1449) & (g1485)) + ((!g4) & (!g1482) & (g1483) & (!g1449) & (g1485)) + ((!g4) & (g1482) & (g1483) & (!g1449) & (!g1485)) + ((!g4) & (g1482) & (g1483) & (!g1449) & (g1485)) + ((!g4) & (g1482) & (g1483) & (g1449) & (!g1485)) + ((!g4) & (g1482) & (g1483) & (g1449) & (g1485)) + ((g4) & (!g1482) & (g1483) & (!g1449) & (!g1485)) + ((g4) & (!g1482) & (g1483) & (!g1449) & (g1485)) + ((g4) & (!g1482) & (g1483) & (g1449) & (!g1485)) + ((g4) & (!g1482) & (g1483) & (g1449) & (g1485)) + ((g4) & (g1482) & (!g1483) & (!g1449) & (!g1485)) + ((g4) & (g1482) & (!g1483) & (g1449) & (!g1485)) + ((g4) & (g1482) & (!g1483) & (g1449) & (g1485)) + ((g4) & (g1482) & (g1483) & (!g1449) & (g1485)));
	assign g1522 = (((!g8) & (!g1452) & (g1481) & (!g1449) & (!g1485)) + ((!g8) & (!g1452) & (g1481) & (g1449) & (!g1485)) + ((!g8) & (!g1452) & (g1481) & (g1449) & (g1485)) + ((!g8) & (g1452) & (!g1481) & (!g1449) & (!g1485)) + ((!g8) & (g1452) & (!g1481) & (!g1449) & (g1485)) + ((!g8) & (g1452) & (!g1481) & (g1449) & (!g1485)) + ((!g8) & (g1452) & (!g1481) & (g1449) & (g1485)) + ((!g8) & (g1452) & (g1481) & (!g1449) & (g1485)) + ((g8) & (!g1452) & (!g1481) & (!g1449) & (!g1485)) + ((g8) & (!g1452) & (!g1481) & (g1449) & (!g1485)) + ((g8) & (!g1452) & (!g1481) & (g1449) & (g1485)) + ((g8) & (g1452) & (!g1481) & (!g1449) & (g1485)) + ((g8) & (g1452) & (g1481) & (!g1449) & (!g1485)) + ((g8) & (g1452) & (g1481) & (!g1449) & (g1485)) + ((g8) & (g1452) & (g1481) & (g1449) & (!g1485)) + ((g8) & (g1452) & (g1481) & (g1449) & (g1485)));
	assign g1523 = (((!g18) & (!g27) & (g1454) & (g1480)) + ((!g18) & (g27) & (!g1454) & (g1480)) + ((!g18) & (g27) & (g1454) & (!g1480)) + ((!g18) & (g27) & (g1454) & (g1480)) + ((g18) & (!g27) & (!g1454) & (!g1480)) + ((g18) & (!g27) & (!g1454) & (g1480)) + ((g18) & (!g27) & (g1454) & (!g1480)) + ((g18) & (g27) & (!g1454) & (!g1480)));
	assign g1524 = (((!g1453) & (!g1449) & (!g1485) & (g1523)) + ((!g1453) & (g1449) & (!g1485) & (g1523)) + ((!g1453) & (g1449) & (g1485) & (g1523)) + ((g1453) & (!g1449) & (!g1485) & (!g1523)) + ((g1453) & (!g1449) & (g1485) & (!g1523)) + ((g1453) & (!g1449) & (g1485) & (g1523)) + ((g1453) & (g1449) & (!g1485) & (!g1523)) + ((g1453) & (g1449) & (g1485) & (!g1523)));
	assign g1525 = (((!g27) & (!g1454) & (g1480) & (!g1449) & (!g1485)) + ((!g27) & (!g1454) & (g1480) & (g1449) & (!g1485)) + ((!g27) & (!g1454) & (g1480) & (g1449) & (g1485)) + ((!g27) & (g1454) & (!g1480) & (!g1449) & (!g1485)) + ((!g27) & (g1454) & (!g1480) & (!g1449) & (g1485)) + ((!g27) & (g1454) & (!g1480) & (g1449) & (!g1485)) + ((!g27) & (g1454) & (!g1480) & (g1449) & (g1485)) + ((!g27) & (g1454) & (g1480) & (!g1449) & (g1485)) + ((g27) & (!g1454) & (!g1480) & (!g1449) & (!g1485)) + ((g27) & (!g1454) & (!g1480) & (g1449) & (!g1485)) + ((g27) & (!g1454) & (!g1480) & (g1449) & (g1485)) + ((g27) & (g1454) & (!g1480) & (!g1449) & (g1485)) + ((g27) & (g1454) & (g1480) & (!g1449) & (!g1485)) + ((g27) & (g1454) & (g1480) & (!g1449) & (g1485)) + ((g27) & (g1454) & (g1480) & (g1449) & (!g1485)) + ((g27) & (g1454) & (g1480) & (g1449) & (g1485)));
	assign g1526 = (((!g39) & (!g54) & (g1456) & (g1479)) + ((!g39) & (g54) & (!g1456) & (g1479)) + ((!g39) & (g54) & (g1456) & (!g1479)) + ((!g39) & (g54) & (g1456) & (g1479)) + ((g39) & (!g54) & (!g1456) & (!g1479)) + ((g39) & (!g54) & (!g1456) & (g1479)) + ((g39) & (!g54) & (g1456) & (!g1479)) + ((g39) & (g54) & (!g1456) & (!g1479)));
	assign g1527 = (((!g1455) & (!g1449) & (!g1485) & (g1526)) + ((!g1455) & (g1449) & (!g1485) & (g1526)) + ((!g1455) & (g1449) & (g1485) & (g1526)) + ((g1455) & (!g1449) & (!g1485) & (!g1526)) + ((g1455) & (!g1449) & (g1485) & (!g1526)) + ((g1455) & (!g1449) & (g1485) & (g1526)) + ((g1455) & (g1449) & (!g1485) & (!g1526)) + ((g1455) & (g1449) & (g1485) & (!g1526)));
	assign g1528 = (((!g54) & (!g1456) & (g1479) & (!g1449) & (!g1485)) + ((!g54) & (!g1456) & (g1479) & (g1449) & (!g1485)) + ((!g54) & (!g1456) & (g1479) & (g1449) & (g1485)) + ((!g54) & (g1456) & (!g1479) & (!g1449) & (!g1485)) + ((!g54) & (g1456) & (!g1479) & (!g1449) & (g1485)) + ((!g54) & (g1456) & (!g1479) & (g1449) & (!g1485)) + ((!g54) & (g1456) & (!g1479) & (g1449) & (g1485)) + ((!g54) & (g1456) & (g1479) & (!g1449) & (g1485)) + ((g54) & (!g1456) & (!g1479) & (!g1449) & (!g1485)) + ((g54) & (!g1456) & (!g1479) & (g1449) & (!g1485)) + ((g54) & (!g1456) & (!g1479) & (g1449) & (g1485)) + ((g54) & (g1456) & (!g1479) & (!g1449) & (g1485)) + ((g54) & (g1456) & (g1479) & (!g1449) & (!g1485)) + ((g54) & (g1456) & (g1479) & (!g1449) & (g1485)) + ((g54) & (g1456) & (g1479) & (g1449) & (!g1485)) + ((g54) & (g1456) & (g1479) & (g1449) & (g1485)));
	assign g1529 = (((!g68) & (!g87) & (g1458) & (g1478)) + ((!g68) & (g87) & (!g1458) & (g1478)) + ((!g68) & (g87) & (g1458) & (!g1478)) + ((!g68) & (g87) & (g1458) & (g1478)) + ((g68) & (!g87) & (!g1458) & (!g1478)) + ((g68) & (!g87) & (!g1458) & (g1478)) + ((g68) & (!g87) & (g1458) & (!g1478)) + ((g68) & (g87) & (!g1458) & (!g1478)));
	assign g1530 = (((!g1457) & (!g1449) & (!g1485) & (g1529)) + ((!g1457) & (g1449) & (!g1485) & (g1529)) + ((!g1457) & (g1449) & (g1485) & (g1529)) + ((g1457) & (!g1449) & (!g1485) & (!g1529)) + ((g1457) & (!g1449) & (g1485) & (!g1529)) + ((g1457) & (!g1449) & (g1485) & (g1529)) + ((g1457) & (g1449) & (!g1485) & (!g1529)) + ((g1457) & (g1449) & (g1485) & (!g1529)));
	assign g1531 = (((!g87) & (!g1458) & (g1478) & (!g1449) & (!g1485)) + ((!g87) & (!g1458) & (g1478) & (g1449) & (!g1485)) + ((!g87) & (!g1458) & (g1478) & (g1449) & (g1485)) + ((!g87) & (g1458) & (!g1478) & (!g1449) & (!g1485)) + ((!g87) & (g1458) & (!g1478) & (!g1449) & (g1485)) + ((!g87) & (g1458) & (!g1478) & (g1449) & (!g1485)) + ((!g87) & (g1458) & (!g1478) & (g1449) & (g1485)) + ((!g87) & (g1458) & (g1478) & (!g1449) & (g1485)) + ((g87) & (!g1458) & (!g1478) & (!g1449) & (!g1485)) + ((g87) & (!g1458) & (!g1478) & (g1449) & (!g1485)) + ((g87) & (!g1458) & (!g1478) & (g1449) & (g1485)) + ((g87) & (g1458) & (!g1478) & (!g1449) & (g1485)) + ((g87) & (g1458) & (g1478) & (!g1449) & (!g1485)) + ((g87) & (g1458) & (g1478) & (!g1449) & (g1485)) + ((g87) & (g1458) & (g1478) & (g1449) & (!g1485)) + ((g87) & (g1458) & (g1478) & (g1449) & (g1485)));
	assign g1532 = (((!g104) & (!g127) & (g1460) & (g1477)) + ((!g104) & (g127) & (!g1460) & (g1477)) + ((!g104) & (g127) & (g1460) & (!g1477)) + ((!g104) & (g127) & (g1460) & (g1477)) + ((g104) & (!g127) & (!g1460) & (!g1477)) + ((g104) & (!g127) & (!g1460) & (g1477)) + ((g104) & (!g127) & (g1460) & (!g1477)) + ((g104) & (g127) & (!g1460) & (!g1477)));
	assign g1533 = (((!g1459) & (!g1449) & (!g1485) & (g1532)) + ((!g1459) & (g1449) & (!g1485) & (g1532)) + ((!g1459) & (g1449) & (g1485) & (g1532)) + ((g1459) & (!g1449) & (!g1485) & (!g1532)) + ((g1459) & (!g1449) & (g1485) & (!g1532)) + ((g1459) & (!g1449) & (g1485) & (g1532)) + ((g1459) & (g1449) & (!g1485) & (!g1532)) + ((g1459) & (g1449) & (g1485) & (!g1532)));
	assign g1534 = (((!g127) & (!g1460) & (g1477) & (!g1449) & (!g1485)) + ((!g127) & (!g1460) & (g1477) & (g1449) & (!g1485)) + ((!g127) & (!g1460) & (g1477) & (g1449) & (g1485)) + ((!g127) & (g1460) & (!g1477) & (!g1449) & (!g1485)) + ((!g127) & (g1460) & (!g1477) & (!g1449) & (g1485)) + ((!g127) & (g1460) & (!g1477) & (g1449) & (!g1485)) + ((!g127) & (g1460) & (!g1477) & (g1449) & (g1485)) + ((!g127) & (g1460) & (g1477) & (!g1449) & (g1485)) + ((g127) & (!g1460) & (!g1477) & (!g1449) & (!g1485)) + ((g127) & (!g1460) & (!g1477) & (g1449) & (!g1485)) + ((g127) & (!g1460) & (!g1477) & (g1449) & (g1485)) + ((g127) & (g1460) & (!g1477) & (!g1449) & (g1485)) + ((g127) & (g1460) & (g1477) & (!g1449) & (!g1485)) + ((g127) & (g1460) & (g1477) & (!g1449) & (g1485)) + ((g127) & (g1460) & (g1477) & (g1449) & (!g1485)) + ((g127) & (g1460) & (g1477) & (g1449) & (g1485)));
	assign g1535 = (((!g147) & (!g174) & (g1462) & (g1476)) + ((!g147) & (g174) & (!g1462) & (g1476)) + ((!g147) & (g174) & (g1462) & (!g1476)) + ((!g147) & (g174) & (g1462) & (g1476)) + ((g147) & (!g174) & (!g1462) & (!g1476)) + ((g147) & (!g174) & (!g1462) & (g1476)) + ((g147) & (!g174) & (g1462) & (!g1476)) + ((g147) & (g174) & (!g1462) & (!g1476)));
	assign g1536 = (((!g1461) & (!g1449) & (!g1485) & (g1535)) + ((!g1461) & (g1449) & (!g1485) & (g1535)) + ((!g1461) & (g1449) & (g1485) & (g1535)) + ((g1461) & (!g1449) & (!g1485) & (!g1535)) + ((g1461) & (!g1449) & (g1485) & (!g1535)) + ((g1461) & (!g1449) & (g1485) & (g1535)) + ((g1461) & (g1449) & (!g1485) & (!g1535)) + ((g1461) & (g1449) & (g1485) & (!g1535)));
	assign g1537 = (((!g174) & (!g1462) & (g1476) & (!g1449) & (!g1485)) + ((!g174) & (!g1462) & (g1476) & (g1449) & (!g1485)) + ((!g174) & (!g1462) & (g1476) & (g1449) & (g1485)) + ((!g174) & (g1462) & (!g1476) & (!g1449) & (!g1485)) + ((!g174) & (g1462) & (!g1476) & (!g1449) & (g1485)) + ((!g174) & (g1462) & (!g1476) & (g1449) & (!g1485)) + ((!g174) & (g1462) & (!g1476) & (g1449) & (g1485)) + ((!g174) & (g1462) & (g1476) & (!g1449) & (g1485)) + ((g174) & (!g1462) & (!g1476) & (!g1449) & (!g1485)) + ((g174) & (!g1462) & (!g1476) & (g1449) & (!g1485)) + ((g174) & (!g1462) & (!g1476) & (g1449) & (g1485)) + ((g174) & (g1462) & (!g1476) & (!g1449) & (g1485)) + ((g174) & (g1462) & (g1476) & (!g1449) & (!g1485)) + ((g174) & (g1462) & (g1476) & (!g1449) & (g1485)) + ((g174) & (g1462) & (g1476) & (g1449) & (!g1485)) + ((g174) & (g1462) & (g1476) & (g1449) & (g1485)));
	assign g1538 = (((!g198) & (!g229) & (g1464) & (g1475)) + ((!g198) & (g229) & (!g1464) & (g1475)) + ((!g198) & (g229) & (g1464) & (!g1475)) + ((!g198) & (g229) & (g1464) & (g1475)) + ((g198) & (!g229) & (!g1464) & (!g1475)) + ((g198) & (!g229) & (!g1464) & (g1475)) + ((g198) & (!g229) & (g1464) & (!g1475)) + ((g198) & (g229) & (!g1464) & (!g1475)));
	assign g1539 = (((!g1463) & (!g1449) & (!g1485) & (g1538)) + ((!g1463) & (g1449) & (!g1485) & (g1538)) + ((!g1463) & (g1449) & (g1485) & (g1538)) + ((g1463) & (!g1449) & (!g1485) & (!g1538)) + ((g1463) & (!g1449) & (g1485) & (!g1538)) + ((g1463) & (!g1449) & (g1485) & (g1538)) + ((g1463) & (g1449) & (!g1485) & (!g1538)) + ((g1463) & (g1449) & (g1485) & (!g1538)));
	assign g1540 = (((!g229) & (!g1464) & (g1475) & (!g1449) & (!g1485)) + ((!g229) & (!g1464) & (g1475) & (g1449) & (!g1485)) + ((!g229) & (!g1464) & (g1475) & (g1449) & (g1485)) + ((!g229) & (g1464) & (!g1475) & (!g1449) & (!g1485)) + ((!g229) & (g1464) & (!g1475) & (!g1449) & (g1485)) + ((!g229) & (g1464) & (!g1475) & (g1449) & (!g1485)) + ((!g229) & (g1464) & (!g1475) & (g1449) & (g1485)) + ((!g229) & (g1464) & (g1475) & (!g1449) & (g1485)) + ((g229) & (!g1464) & (!g1475) & (!g1449) & (!g1485)) + ((g229) & (!g1464) & (!g1475) & (g1449) & (!g1485)) + ((g229) & (!g1464) & (!g1475) & (g1449) & (g1485)) + ((g229) & (g1464) & (!g1475) & (!g1449) & (g1485)) + ((g229) & (g1464) & (g1475) & (!g1449) & (!g1485)) + ((g229) & (g1464) & (g1475) & (!g1449) & (g1485)) + ((g229) & (g1464) & (g1475) & (g1449) & (!g1485)) + ((g229) & (g1464) & (g1475) & (g1449) & (g1485)));
	assign g1541 = (((!g255) & (!g290) & (g1466) & (g1474)) + ((!g255) & (g290) & (!g1466) & (g1474)) + ((!g255) & (g290) & (g1466) & (!g1474)) + ((!g255) & (g290) & (g1466) & (g1474)) + ((g255) & (!g290) & (!g1466) & (!g1474)) + ((g255) & (!g290) & (!g1466) & (g1474)) + ((g255) & (!g290) & (g1466) & (!g1474)) + ((g255) & (g290) & (!g1466) & (!g1474)));
	assign g1542 = (((!g1465) & (!g1449) & (!g1485) & (g1541)) + ((!g1465) & (g1449) & (!g1485) & (g1541)) + ((!g1465) & (g1449) & (g1485) & (g1541)) + ((g1465) & (!g1449) & (!g1485) & (!g1541)) + ((g1465) & (!g1449) & (g1485) & (!g1541)) + ((g1465) & (!g1449) & (g1485) & (g1541)) + ((g1465) & (g1449) & (!g1485) & (!g1541)) + ((g1465) & (g1449) & (g1485) & (!g1541)));
	assign g1543 = (((!g290) & (!g1466) & (g1474) & (!g1449) & (!g1485)) + ((!g290) & (!g1466) & (g1474) & (g1449) & (!g1485)) + ((!g290) & (!g1466) & (g1474) & (g1449) & (g1485)) + ((!g290) & (g1466) & (!g1474) & (!g1449) & (!g1485)) + ((!g290) & (g1466) & (!g1474) & (!g1449) & (g1485)) + ((!g290) & (g1466) & (!g1474) & (g1449) & (!g1485)) + ((!g290) & (g1466) & (!g1474) & (g1449) & (g1485)) + ((!g290) & (g1466) & (g1474) & (!g1449) & (g1485)) + ((g290) & (!g1466) & (!g1474) & (!g1449) & (!g1485)) + ((g290) & (!g1466) & (!g1474) & (g1449) & (!g1485)) + ((g290) & (!g1466) & (!g1474) & (g1449) & (g1485)) + ((g290) & (g1466) & (!g1474) & (!g1449) & (g1485)) + ((g290) & (g1466) & (g1474) & (!g1449) & (!g1485)) + ((g290) & (g1466) & (g1474) & (!g1449) & (g1485)) + ((g290) & (g1466) & (g1474) & (g1449) & (!g1485)) + ((g290) & (g1466) & (g1474) & (g1449) & (g1485)));
	assign g1544 = (((!g319) & (!g358) & (g1468) & (g1473)) + ((!g319) & (g358) & (!g1468) & (g1473)) + ((!g319) & (g358) & (g1468) & (!g1473)) + ((!g319) & (g358) & (g1468) & (g1473)) + ((g319) & (!g358) & (!g1468) & (!g1473)) + ((g319) & (!g358) & (!g1468) & (g1473)) + ((g319) & (!g358) & (g1468) & (!g1473)) + ((g319) & (g358) & (!g1468) & (!g1473)));
	assign g1545 = (((!g1467) & (!g1449) & (!g1485) & (g1544)) + ((!g1467) & (g1449) & (!g1485) & (g1544)) + ((!g1467) & (g1449) & (g1485) & (g1544)) + ((g1467) & (!g1449) & (!g1485) & (!g1544)) + ((g1467) & (!g1449) & (g1485) & (!g1544)) + ((g1467) & (!g1449) & (g1485) & (g1544)) + ((g1467) & (g1449) & (!g1485) & (!g1544)) + ((g1467) & (g1449) & (g1485) & (!g1544)));
	assign g1546 = (((!g358) & (!g1468) & (g1473) & (!g1449) & (!g1485)) + ((!g358) & (!g1468) & (g1473) & (g1449) & (!g1485)) + ((!g358) & (!g1468) & (g1473) & (g1449) & (g1485)) + ((!g358) & (g1468) & (!g1473) & (!g1449) & (!g1485)) + ((!g358) & (g1468) & (!g1473) & (!g1449) & (g1485)) + ((!g358) & (g1468) & (!g1473) & (g1449) & (!g1485)) + ((!g358) & (g1468) & (!g1473) & (g1449) & (g1485)) + ((!g358) & (g1468) & (g1473) & (!g1449) & (g1485)) + ((g358) & (!g1468) & (!g1473) & (!g1449) & (!g1485)) + ((g358) & (!g1468) & (!g1473) & (g1449) & (!g1485)) + ((g358) & (!g1468) & (!g1473) & (g1449) & (g1485)) + ((g358) & (g1468) & (!g1473) & (!g1449) & (g1485)) + ((g358) & (g1468) & (g1473) & (!g1449) & (!g1485)) + ((g358) & (g1468) & (g1473) & (!g1449) & (g1485)) + ((g358) & (g1468) & (g1473) & (g1449) & (!g1485)) + ((g358) & (g1468) & (g1473) & (g1449) & (g1485)));
	assign g1547 = (((!g390) & (!g433) & (g1470) & (g1472)) + ((!g390) & (g433) & (!g1470) & (g1472)) + ((!g390) & (g433) & (g1470) & (!g1472)) + ((!g390) & (g433) & (g1470) & (g1472)) + ((g390) & (!g433) & (!g1470) & (!g1472)) + ((g390) & (!g433) & (!g1470) & (g1472)) + ((g390) & (!g433) & (g1470) & (!g1472)) + ((g390) & (g433) & (!g1470) & (!g1472)));
	assign g1548 = (((!g1469) & (!g1449) & (!g1485) & (g1547)) + ((!g1469) & (g1449) & (!g1485) & (g1547)) + ((!g1469) & (g1449) & (g1485) & (g1547)) + ((g1469) & (!g1449) & (!g1485) & (!g1547)) + ((g1469) & (!g1449) & (g1485) & (!g1547)) + ((g1469) & (!g1449) & (g1485) & (g1547)) + ((g1469) & (g1449) & (!g1485) & (!g1547)) + ((g1469) & (g1449) & (g1485) & (!g1547)));
	assign g1549 = (((!g433) & (!g1470) & (g1472) & (!g1449) & (!g1485)) + ((!g433) & (!g1470) & (g1472) & (g1449) & (!g1485)) + ((!g433) & (!g1470) & (g1472) & (g1449) & (g1485)) + ((!g433) & (g1470) & (!g1472) & (!g1449) & (!g1485)) + ((!g433) & (g1470) & (!g1472) & (!g1449) & (g1485)) + ((!g433) & (g1470) & (!g1472) & (g1449) & (!g1485)) + ((!g433) & (g1470) & (!g1472) & (g1449) & (g1485)) + ((!g433) & (g1470) & (g1472) & (!g1449) & (g1485)) + ((g433) & (!g1470) & (!g1472) & (!g1449) & (!g1485)) + ((g433) & (!g1470) & (!g1472) & (g1449) & (!g1485)) + ((g433) & (!g1470) & (!g1472) & (g1449) & (g1485)) + ((g433) & (g1470) & (!g1472) & (!g1449) & (g1485)) + ((g433) & (g1470) & (g1472) & (!g1449) & (!g1485)) + ((g433) & (g1470) & (g1472) & (!g1449) & (g1485)) + ((g433) & (g1470) & (g1472) & (g1449) & (!g1485)) + ((g433) & (g1470) & (g1472) & (g1449) & (g1485)));
	assign g1550 = (((!g468) & (!g515) & (g1424) & (g1448)) + ((!g468) & (g515) & (!g1424) & (g1448)) + ((!g468) & (g515) & (g1424) & (!g1448)) + ((!g468) & (g515) & (g1424) & (g1448)) + ((g468) & (!g515) & (!g1424) & (!g1448)) + ((g468) & (!g515) & (!g1424) & (g1448)) + ((g468) & (!g515) & (g1424) & (!g1448)) + ((g468) & (g515) & (!g1424) & (!g1448)));
	assign g1551 = (((!g1471) & (!g1449) & (!g1485) & (g1550)) + ((!g1471) & (g1449) & (!g1485) & (g1550)) + ((!g1471) & (g1449) & (g1485) & (g1550)) + ((g1471) & (!g1449) & (!g1485) & (!g1550)) + ((g1471) & (!g1449) & (g1485) & (!g1550)) + ((g1471) & (!g1449) & (g1485) & (g1550)) + ((g1471) & (g1449) & (!g1485) & (!g1550)) + ((g1471) & (g1449) & (g1485) & (!g1550)));
	assign g1552 = (((!g433) & (!g468) & (g1551) & (g1486) & (g1520)) + ((!g433) & (g468) & (g1551) & (!g1486) & (g1520)) + ((!g433) & (g468) & (g1551) & (g1486) & (!g1520)) + ((!g433) & (g468) & (g1551) & (g1486) & (g1520)) + ((g433) & (!g468) & (!g1551) & (g1486) & (g1520)) + ((g433) & (!g468) & (g1551) & (!g1486) & (!g1520)) + ((g433) & (!g468) & (g1551) & (!g1486) & (g1520)) + ((g433) & (!g468) & (g1551) & (g1486) & (!g1520)) + ((g433) & (!g468) & (g1551) & (g1486) & (g1520)) + ((g433) & (g468) & (!g1551) & (!g1486) & (g1520)) + ((g433) & (g468) & (!g1551) & (g1486) & (!g1520)) + ((g433) & (g468) & (!g1551) & (g1486) & (g1520)) + ((g433) & (g468) & (g1551) & (!g1486) & (!g1520)) + ((g433) & (g468) & (g1551) & (!g1486) & (g1520)) + ((g433) & (g468) & (g1551) & (g1486) & (!g1520)) + ((g433) & (g468) & (g1551) & (g1486) & (g1520)));
	assign g1553 = (((!g358) & (!g390) & (g1548) & (g1549) & (g1552)) + ((!g358) & (g390) & (g1548) & (!g1549) & (g1552)) + ((!g358) & (g390) & (g1548) & (g1549) & (!g1552)) + ((!g358) & (g390) & (g1548) & (g1549) & (g1552)) + ((g358) & (!g390) & (!g1548) & (g1549) & (g1552)) + ((g358) & (!g390) & (g1548) & (!g1549) & (!g1552)) + ((g358) & (!g390) & (g1548) & (!g1549) & (g1552)) + ((g358) & (!g390) & (g1548) & (g1549) & (!g1552)) + ((g358) & (!g390) & (g1548) & (g1549) & (g1552)) + ((g358) & (g390) & (!g1548) & (!g1549) & (g1552)) + ((g358) & (g390) & (!g1548) & (g1549) & (!g1552)) + ((g358) & (g390) & (!g1548) & (g1549) & (g1552)) + ((g358) & (g390) & (g1548) & (!g1549) & (!g1552)) + ((g358) & (g390) & (g1548) & (!g1549) & (g1552)) + ((g358) & (g390) & (g1548) & (g1549) & (!g1552)) + ((g358) & (g390) & (g1548) & (g1549) & (g1552)));
	assign g1554 = (((!g290) & (!g319) & (g1545) & (g1546) & (g1553)) + ((!g290) & (g319) & (g1545) & (!g1546) & (g1553)) + ((!g290) & (g319) & (g1545) & (g1546) & (!g1553)) + ((!g290) & (g319) & (g1545) & (g1546) & (g1553)) + ((g290) & (!g319) & (!g1545) & (g1546) & (g1553)) + ((g290) & (!g319) & (g1545) & (!g1546) & (!g1553)) + ((g290) & (!g319) & (g1545) & (!g1546) & (g1553)) + ((g290) & (!g319) & (g1545) & (g1546) & (!g1553)) + ((g290) & (!g319) & (g1545) & (g1546) & (g1553)) + ((g290) & (g319) & (!g1545) & (!g1546) & (g1553)) + ((g290) & (g319) & (!g1545) & (g1546) & (!g1553)) + ((g290) & (g319) & (!g1545) & (g1546) & (g1553)) + ((g290) & (g319) & (g1545) & (!g1546) & (!g1553)) + ((g290) & (g319) & (g1545) & (!g1546) & (g1553)) + ((g290) & (g319) & (g1545) & (g1546) & (!g1553)) + ((g290) & (g319) & (g1545) & (g1546) & (g1553)));
	assign g1555 = (((!g229) & (!g255) & (g1542) & (g1543) & (g1554)) + ((!g229) & (g255) & (g1542) & (!g1543) & (g1554)) + ((!g229) & (g255) & (g1542) & (g1543) & (!g1554)) + ((!g229) & (g255) & (g1542) & (g1543) & (g1554)) + ((g229) & (!g255) & (!g1542) & (g1543) & (g1554)) + ((g229) & (!g255) & (g1542) & (!g1543) & (!g1554)) + ((g229) & (!g255) & (g1542) & (!g1543) & (g1554)) + ((g229) & (!g255) & (g1542) & (g1543) & (!g1554)) + ((g229) & (!g255) & (g1542) & (g1543) & (g1554)) + ((g229) & (g255) & (!g1542) & (!g1543) & (g1554)) + ((g229) & (g255) & (!g1542) & (g1543) & (!g1554)) + ((g229) & (g255) & (!g1542) & (g1543) & (g1554)) + ((g229) & (g255) & (g1542) & (!g1543) & (!g1554)) + ((g229) & (g255) & (g1542) & (!g1543) & (g1554)) + ((g229) & (g255) & (g1542) & (g1543) & (!g1554)) + ((g229) & (g255) & (g1542) & (g1543) & (g1554)));
	assign g1556 = (((!g174) & (!g198) & (g1539) & (g1540) & (g1555)) + ((!g174) & (g198) & (g1539) & (!g1540) & (g1555)) + ((!g174) & (g198) & (g1539) & (g1540) & (!g1555)) + ((!g174) & (g198) & (g1539) & (g1540) & (g1555)) + ((g174) & (!g198) & (!g1539) & (g1540) & (g1555)) + ((g174) & (!g198) & (g1539) & (!g1540) & (!g1555)) + ((g174) & (!g198) & (g1539) & (!g1540) & (g1555)) + ((g174) & (!g198) & (g1539) & (g1540) & (!g1555)) + ((g174) & (!g198) & (g1539) & (g1540) & (g1555)) + ((g174) & (g198) & (!g1539) & (!g1540) & (g1555)) + ((g174) & (g198) & (!g1539) & (g1540) & (!g1555)) + ((g174) & (g198) & (!g1539) & (g1540) & (g1555)) + ((g174) & (g198) & (g1539) & (!g1540) & (!g1555)) + ((g174) & (g198) & (g1539) & (!g1540) & (g1555)) + ((g174) & (g198) & (g1539) & (g1540) & (!g1555)) + ((g174) & (g198) & (g1539) & (g1540) & (g1555)));
	assign g1557 = (((!g127) & (!g147) & (g1536) & (g1537) & (g1556)) + ((!g127) & (g147) & (g1536) & (!g1537) & (g1556)) + ((!g127) & (g147) & (g1536) & (g1537) & (!g1556)) + ((!g127) & (g147) & (g1536) & (g1537) & (g1556)) + ((g127) & (!g147) & (!g1536) & (g1537) & (g1556)) + ((g127) & (!g147) & (g1536) & (!g1537) & (!g1556)) + ((g127) & (!g147) & (g1536) & (!g1537) & (g1556)) + ((g127) & (!g147) & (g1536) & (g1537) & (!g1556)) + ((g127) & (!g147) & (g1536) & (g1537) & (g1556)) + ((g127) & (g147) & (!g1536) & (!g1537) & (g1556)) + ((g127) & (g147) & (!g1536) & (g1537) & (!g1556)) + ((g127) & (g147) & (!g1536) & (g1537) & (g1556)) + ((g127) & (g147) & (g1536) & (!g1537) & (!g1556)) + ((g127) & (g147) & (g1536) & (!g1537) & (g1556)) + ((g127) & (g147) & (g1536) & (g1537) & (!g1556)) + ((g127) & (g147) & (g1536) & (g1537) & (g1556)));
	assign g1558 = (((!g87) & (!g104) & (g1533) & (g1534) & (g1557)) + ((!g87) & (g104) & (g1533) & (!g1534) & (g1557)) + ((!g87) & (g104) & (g1533) & (g1534) & (!g1557)) + ((!g87) & (g104) & (g1533) & (g1534) & (g1557)) + ((g87) & (!g104) & (!g1533) & (g1534) & (g1557)) + ((g87) & (!g104) & (g1533) & (!g1534) & (!g1557)) + ((g87) & (!g104) & (g1533) & (!g1534) & (g1557)) + ((g87) & (!g104) & (g1533) & (g1534) & (!g1557)) + ((g87) & (!g104) & (g1533) & (g1534) & (g1557)) + ((g87) & (g104) & (!g1533) & (!g1534) & (g1557)) + ((g87) & (g104) & (!g1533) & (g1534) & (!g1557)) + ((g87) & (g104) & (!g1533) & (g1534) & (g1557)) + ((g87) & (g104) & (g1533) & (!g1534) & (!g1557)) + ((g87) & (g104) & (g1533) & (!g1534) & (g1557)) + ((g87) & (g104) & (g1533) & (g1534) & (!g1557)) + ((g87) & (g104) & (g1533) & (g1534) & (g1557)));
	assign g1559 = (((!g54) & (!g68) & (g1530) & (g1531) & (g1558)) + ((!g54) & (g68) & (g1530) & (!g1531) & (g1558)) + ((!g54) & (g68) & (g1530) & (g1531) & (!g1558)) + ((!g54) & (g68) & (g1530) & (g1531) & (g1558)) + ((g54) & (!g68) & (!g1530) & (g1531) & (g1558)) + ((g54) & (!g68) & (g1530) & (!g1531) & (!g1558)) + ((g54) & (!g68) & (g1530) & (!g1531) & (g1558)) + ((g54) & (!g68) & (g1530) & (g1531) & (!g1558)) + ((g54) & (!g68) & (g1530) & (g1531) & (g1558)) + ((g54) & (g68) & (!g1530) & (!g1531) & (g1558)) + ((g54) & (g68) & (!g1530) & (g1531) & (!g1558)) + ((g54) & (g68) & (!g1530) & (g1531) & (g1558)) + ((g54) & (g68) & (g1530) & (!g1531) & (!g1558)) + ((g54) & (g68) & (g1530) & (!g1531) & (g1558)) + ((g54) & (g68) & (g1530) & (g1531) & (!g1558)) + ((g54) & (g68) & (g1530) & (g1531) & (g1558)));
	assign g1560 = (((!g27) & (!g39) & (g1527) & (g1528) & (g1559)) + ((!g27) & (g39) & (g1527) & (!g1528) & (g1559)) + ((!g27) & (g39) & (g1527) & (g1528) & (!g1559)) + ((!g27) & (g39) & (g1527) & (g1528) & (g1559)) + ((g27) & (!g39) & (!g1527) & (g1528) & (g1559)) + ((g27) & (!g39) & (g1527) & (!g1528) & (!g1559)) + ((g27) & (!g39) & (g1527) & (!g1528) & (g1559)) + ((g27) & (!g39) & (g1527) & (g1528) & (!g1559)) + ((g27) & (!g39) & (g1527) & (g1528) & (g1559)) + ((g27) & (g39) & (!g1527) & (!g1528) & (g1559)) + ((g27) & (g39) & (!g1527) & (g1528) & (!g1559)) + ((g27) & (g39) & (!g1527) & (g1528) & (g1559)) + ((g27) & (g39) & (g1527) & (!g1528) & (!g1559)) + ((g27) & (g39) & (g1527) & (!g1528) & (g1559)) + ((g27) & (g39) & (g1527) & (g1528) & (!g1559)) + ((g27) & (g39) & (g1527) & (g1528) & (g1559)));
	assign g1561 = (((!g8) & (!g18) & (g1524) & (g1525) & (g1560)) + ((!g8) & (g18) & (g1524) & (!g1525) & (g1560)) + ((!g8) & (g18) & (g1524) & (g1525) & (!g1560)) + ((!g8) & (g18) & (g1524) & (g1525) & (g1560)) + ((g8) & (!g18) & (!g1524) & (g1525) & (g1560)) + ((g8) & (!g18) & (g1524) & (!g1525) & (!g1560)) + ((g8) & (!g18) & (g1524) & (!g1525) & (g1560)) + ((g8) & (!g18) & (g1524) & (g1525) & (!g1560)) + ((g8) & (!g18) & (g1524) & (g1525) & (g1560)) + ((g8) & (g18) & (!g1524) & (!g1525) & (g1560)) + ((g8) & (g18) & (!g1524) & (g1525) & (!g1560)) + ((g8) & (g18) & (!g1524) & (g1525) & (g1560)) + ((g8) & (g18) & (g1524) & (!g1525) & (!g1560)) + ((g8) & (g18) & (g1524) & (!g1525) & (g1560)) + ((g8) & (g18) & (g1524) & (g1525) & (!g1560)) + ((g8) & (g18) & (g1524) & (g1525) & (g1560)));
	assign g1562 = (((!g2) & (!g8) & (g1452) & (g1481)) + ((!g2) & (g8) & (!g1452) & (g1481)) + ((!g2) & (g8) & (g1452) & (!g1481)) + ((!g2) & (g8) & (g1452) & (g1481)) + ((g2) & (!g8) & (!g1452) & (!g1481)) + ((g2) & (!g8) & (!g1452) & (g1481)) + ((g2) & (!g8) & (g1452) & (!g1481)) + ((g2) & (g8) & (!g1452) & (!g1481)));
	assign g1563 = (((!g1451) & (!g1449) & (!g1485) & (g1562)) + ((!g1451) & (g1449) & (!g1485) & (g1562)) + ((!g1451) & (g1449) & (g1485) & (g1562)) + ((g1451) & (!g1449) & (!g1485) & (!g1562)) + ((g1451) & (!g1449) & (g1485) & (!g1562)) + ((g1451) & (!g1449) & (g1485) & (g1562)) + ((g1451) & (g1449) & (!g1485) & (!g1562)) + ((g1451) & (g1449) & (g1485) & (!g1562)));
	assign g1564 = (((!g4) & (!g2) & (!g1522) & (!g1561) & (g1563)) + ((!g4) & (!g2) & (!g1522) & (g1561) & (g1563)) + ((!g4) & (!g2) & (g1522) & (!g1561) & (g1563)) + ((!g4) & (!g2) & (g1522) & (g1561) & (!g1563)) + ((!g4) & (!g2) & (g1522) & (g1561) & (g1563)) + ((!g4) & (g2) & (!g1522) & (!g1561) & (g1563)) + ((!g4) & (g2) & (!g1522) & (g1561) & (!g1563)) + ((!g4) & (g2) & (!g1522) & (g1561) & (g1563)) + ((!g4) & (g2) & (g1522) & (!g1561) & (!g1563)) + ((!g4) & (g2) & (g1522) & (!g1561) & (g1563)) + ((!g4) & (g2) & (g1522) & (g1561) & (!g1563)) + ((!g4) & (g2) & (g1522) & (g1561) & (g1563)) + ((g4) & (!g2) & (g1522) & (g1561) & (g1563)) + ((g4) & (g2) & (!g1522) & (g1561) & (g1563)) + ((g4) & (g2) & (g1522) & (!g1561) & (g1563)) + ((g4) & (g2) & (g1522) & (g1561) & (g1563)));
	assign g1565 = (((!g4) & (!g1482) & (g1483)) + ((!g4) & (g1482) & (!g1483)) + ((!g4) & (g1482) & (g1483)) + ((g4) & (g1482) & (g1483)));
	assign g1566 = (((!g1450) & (!g1565) & (!g1449) & (!g1485)) + ((!g1450) & (!g1565) & (g1449) & (!g1485)) + ((!g1450) & (!g1565) & (g1449) & (g1485)) + ((g1450) & (g1565) & (!g1449) & (!g1485)) + ((g1450) & (g1565) & (!g1449) & (g1485)) + ((g1450) & (g1565) & (g1449) & (!g1485)) + ((g1450) & (g1565) & (g1449) & (g1485)));
	assign g1567 = (((!g1) & (g1450) & (!g1565) & (!g1449) & (g1485)) + ((!g1) & (g1450) & (g1565) & (!g1449) & (g1485)) + ((g1) & (!g1450) & (g1565) & (g1449) & (!g1485)) + ((g1) & (!g1450) & (g1565) & (g1449) & (g1485)) + ((g1) & (g1450) & (!g1565) & (!g1449) & (!g1485)) + ((g1) & (g1450) & (!g1565) & (!g1449) & (g1485)) + ((g1) & (g1450) & (!g1565) & (g1449) & (!g1485)) + ((g1) & (g1450) & (!g1565) & (g1449) & (g1485)) + ((g1) & (g1450) & (g1565) & (!g1449) & (g1485)));
	assign g1568 = (((!g1) & (!g1521) & (!g1564) & (!g1566) & (!g1567)) + ((g1) & (!g1521) & (!g1564) & (!g1566) & (!g1567)) + ((g1) & (!g1521) & (!g1564) & (g1566) & (!g1567)) + ((g1) & (!g1521) & (g1564) & (!g1566) & (!g1567)) + ((g1) & (!g1521) & (g1564) & (g1566) & (!g1567)) + ((g1) & (g1521) & (!g1564) & (!g1566) & (!g1567)) + ((g1) & (g1521) & (!g1564) & (g1566) & (!g1567)));
	assign g1569 = (((!g468) & (!g1486) & (g1520) & (!g1568)) + ((!g468) & (g1486) & (!g1520) & (!g1568)) + ((!g468) & (g1486) & (!g1520) & (g1568)) + ((!g468) & (g1486) & (g1520) & (g1568)) + ((g468) & (!g1486) & (!g1520) & (!g1568)) + ((g468) & (g1486) & (!g1520) & (g1568)) + ((g468) & (g1486) & (g1520) & (!g1568)) + ((g468) & (g1486) & (g1520) & (g1568)));
	assign g1570 = (((!g515) & (!g553) & (!g1488) & (g1489) & (g1519) & (!g1568)) + ((!g515) & (!g553) & (g1488) & (!g1489) & (!g1519) & (!g1568)) + ((!g515) & (!g553) & (g1488) & (!g1489) & (!g1519) & (g1568)) + ((!g515) & (!g553) & (g1488) & (!g1489) & (g1519) & (!g1568)) + ((!g515) & (!g553) & (g1488) & (!g1489) & (g1519) & (g1568)) + ((!g515) & (!g553) & (g1488) & (g1489) & (!g1519) & (!g1568)) + ((!g515) & (!g553) & (g1488) & (g1489) & (!g1519) & (g1568)) + ((!g515) & (!g553) & (g1488) & (g1489) & (g1519) & (g1568)) + ((!g515) & (g553) & (!g1488) & (!g1489) & (g1519) & (!g1568)) + ((!g515) & (g553) & (!g1488) & (g1489) & (!g1519) & (!g1568)) + ((!g515) & (g553) & (!g1488) & (g1489) & (g1519) & (!g1568)) + ((!g515) & (g553) & (g1488) & (!g1489) & (!g1519) & (!g1568)) + ((!g515) & (g553) & (g1488) & (!g1489) & (!g1519) & (g1568)) + ((!g515) & (g553) & (g1488) & (!g1489) & (g1519) & (g1568)) + ((!g515) & (g553) & (g1488) & (g1489) & (!g1519) & (g1568)) + ((!g515) & (g553) & (g1488) & (g1489) & (g1519) & (g1568)) + ((g515) & (!g553) & (!g1488) & (!g1489) & (!g1519) & (!g1568)) + ((g515) & (!g553) & (!g1488) & (!g1489) & (g1519) & (!g1568)) + ((g515) & (!g553) & (!g1488) & (g1489) & (!g1519) & (!g1568)) + ((g515) & (!g553) & (g1488) & (!g1489) & (!g1519) & (g1568)) + ((g515) & (!g553) & (g1488) & (!g1489) & (g1519) & (g1568)) + ((g515) & (!g553) & (g1488) & (g1489) & (!g1519) & (g1568)) + ((g515) & (!g553) & (g1488) & (g1489) & (g1519) & (!g1568)) + ((g515) & (!g553) & (g1488) & (g1489) & (g1519) & (g1568)) + ((g515) & (g553) & (!g1488) & (!g1489) & (!g1519) & (!g1568)) + ((g515) & (g553) & (g1488) & (!g1489) & (!g1519) & (g1568)) + ((g515) & (g553) & (g1488) & (!g1489) & (g1519) & (!g1568)) + ((g515) & (g553) & (g1488) & (!g1489) & (g1519) & (g1568)) + ((g515) & (g553) & (g1488) & (g1489) & (!g1519) & (!g1568)) + ((g515) & (g553) & (g1488) & (g1489) & (!g1519) & (g1568)) + ((g515) & (g553) & (g1488) & (g1489) & (g1519) & (!g1568)) + ((g515) & (g553) & (g1488) & (g1489) & (g1519) & (g1568)));
	assign g1571 = (((!g553) & (!g1489) & (g1519) & (!g1568)) + ((!g553) & (g1489) & (!g1519) & (!g1568)) + ((!g553) & (g1489) & (!g1519) & (g1568)) + ((!g553) & (g1489) & (g1519) & (g1568)) + ((g553) & (!g1489) & (!g1519) & (!g1568)) + ((g553) & (g1489) & (!g1519) & (g1568)) + ((g553) & (g1489) & (g1519) & (!g1568)) + ((g553) & (g1489) & (g1519) & (g1568)));
	assign g1572 = (((!g604) & (!g645) & (!g1491) & (g1492) & (g1518) & (!g1568)) + ((!g604) & (!g645) & (g1491) & (!g1492) & (!g1518) & (!g1568)) + ((!g604) & (!g645) & (g1491) & (!g1492) & (!g1518) & (g1568)) + ((!g604) & (!g645) & (g1491) & (!g1492) & (g1518) & (!g1568)) + ((!g604) & (!g645) & (g1491) & (!g1492) & (g1518) & (g1568)) + ((!g604) & (!g645) & (g1491) & (g1492) & (!g1518) & (!g1568)) + ((!g604) & (!g645) & (g1491) & (g1492) & (!g1518) & (g1568)) + ((!g604) & (!g645) & (g1491) & (g1492) & (g1518) & (g1568)) + ((!g604) & (g645) & (!g1491) & (!g1492) & (g1518) & (!g1568)) + ((!g604) & (g645) & (!g1491) & (g1492) & (!g1518) & (!g1568)) + ((!g604) & (g645) & (!g1491) & (g1492) & (g1518) & (!g1568)) + ((!g604) & (g645) & (g1491) & (!g1492) & (!g1518) & (!g1568)) + ((!g604) & (g645) & (g1491) & (!g1492) & (!g1518) & (g1568)) + ((!g604) & (g645) & (g1491) & (!g1492) & (g1518) & (g1568)) + ((!g604) & (g645) & (g1491) & (g1492) & (!g1518) & (g1568)) + ((!g604) & (g645) & (g1491) & (g1492) & (g1518) & (g1568)) + ((g604) & (!g645) & (!g1491) & (!g1492) & (!g1518) & (!g1568)) + ((g604) & (!g645) & (!g1491) & (!g1492) & (g1518) & (!g1568)) + ((g604) & (!g645) & (!g1491) & (g1492) & (!g1518) & (!g1568)) + ((g604) & (!g645) & (g1491) & (!g1492) & (!g1518) & (g1568)) + ((g604) & (!g645) & (g1491) & (!g1492) & (g1518) & (g1568)) + ((g604) & (!g645) & (g1491) & (g1492) & (!g1518) & (g1568)) + ((g604) & (!g645) & (g1491) & (g1492) & (g1518) & (!g1568)) + ((g604) & (!g645) & (g1491) & (g1492) & (g1518) & (g1568)) + ((g604) & (g645) & (!g1491) & (!g1492) & (!g1518) & (!g1568)) + ((g604) & (g645) & (g1491) & (!g1492) & (!g1518) & (g1568)) + ((g604) & (g645) & (g1491) & (!g1492) & (g1518) & (!g1568)) + ((g604) & (g645) & (g1491) & (!g1492) & (g1518) & (g1568)) + ((g604) & (g645) & (g1491) & (g1492) & (!g1518) & (!g1568)) + ((g604) & (g645) & (g1491) & (g1492) & (!g1518) & (g1568)) + ((g604) & (g645) & (g1491) & (g1492) & (g1518) & (!g1568)) + ((g604) & (g645) & (g1491) & (g1492) & (g1518) & (g1568)));
	assign g1573 = (((!g645) & (!g1492) & (g1518) & (!g1568)) + ((!g645) & (g1492) & (!g1518) & (!g1568)) + ((!g645) & (g1492) & (!g1518) & (g1568)) + ((!g645) & (g1492) & (g1518) & (g1568)) + ((g645) & (!g1492) & (!g1518) & (!g1568)) + ((g645) & (g1492) & (!g1518) & (g1568)) + ((g645) & (g1492) & (g1518) & (!g1568)) + ((g645) & (g1492) & (g1518) & (g1568)));
	assign g1574 = (((!g700) & (!g744) & (!g1494) & (g1495) & (g1517) & (!g1568)) + ((!g700) & (!g744) & (g1494) & (!g1495) & (!g1517) & (!g1568)) + ((!g700) & (!g744) & (g1494) & (!g1495) & (!g1517) & (g1568)) + ((!g700) & (!g744) & (g1494) & (!g1495) & (g1517) & (!g1568)) + ((!g700) & (!g744) & (g1494) & (!g1495) & (g1517) & (g1568)) + ((!g700) & (!g744) & (g1494) & (g1495) & (!g1517) & (!g1568)) + ((!g700) & (!g744) & (g1494) & (g1495) & (!g1517) & (g1568)) + ((!g700) & (!g744) & (g1494) & (g1495) & (g1517) & (g1568)) + ((!g700) & (g744) & (!g1494) & (!g1495) & (g1517) & (!g1568)) + ((!g700) & (g744) & (!g1494) & (g1495) & (!g1517) & (!g1568)) + ((!g700) & (g744) & (!g1494) & (g1495) & (g1517) & (!g1568)) + ((!g700) & (g744) & (g1494) & (!g1495) & (!g1517) & (!g1568)) + ((!g700) & (g744) & (g1494) & (!g1495) & (!g1517) & (g1568)) + ((!g700) & (g744) & (g1494) & (!g1495) & (g1517) & (g1568)) + ((!g700) & (g744) & (g1494) & (g1495) & (!g1517) & (g1568)) + ((!g700) & (g744) & (g1494) & (g1495) & (g1517) & (g1568)) + ((g700) & (!g744) & (!g1494) & (!g1495) & (!g1517) & (!g1568)) + ((g700) & (!g744) & (!g1494) & (!g1495) & (g1517) & (!g1568)) + ((g700) & (!g744) & (!g1494) & (g1495) & (!g1517) & (!g1568)) + ((g700) & (!g744) & (g1494) & (!g1495) & (!g1517) & (g1568)) + ((g700) & (!g744) & (g1494) & (!g1495) & (g1517) & (g1568)) + ((g700) & (!g744) & (g1494) & (g1495) & (!g1517) & (g1568)) + ((g700) & (!g744) & (g1494) & (g1495) & (g1517) & (!g1568)) + ((g700) & (!g744) & (g1494) & (g1495) & (g1517) & (g1568)) + ((g700) & (g744) & (!g1494) & (!g1495) & (!g1517) & (!g1568)) + ((g700) & (g744) & (g1494) & (!g1495) & (!g1517) & (g1568)) + ((g700) & (g744) & (g1494) & (!g1495) & (g1517) & (!g1568)) + ((g700) & (g744) & (g1494) & (!g1495) & (g1517) & (g1568)) + ((g700) & (g744) & (g1494) & (g1495) & (!g1517) & (!g1568)) + ((g700) & (g744) & (g1494) & (g1495) & (!g1517) & (g1568)) + ((g700) & (g744) & (g1494) & (g1495) & (g1517) & (!g1568)) + ((g700) & (g744) & (g1494) & (g1495) & (g1517) & (g1568)));
	assign g1575 = (((!g744) & (!g1495) & (g1517) & (!g1568)) + ((!g744) & (g1495) & (!g1517) & (!g1568)) + ((!g744) & (g1495) & (!g1517) & (g1568)) + ((!g744) & (g1495) & (g1517) & (g1568)) + ((g744) & (!g1495) & (!g1517) & (!g1568)) + ((g744) & (g1495) & (!g1517) & (g1568)) + ((g744) & (g1495) & (g1517) & (!g1568)) + ((g744) & (g1495) & (g1517) & (g1568)));
	assign g1576 = (((!g803) & (!g851) & (!g1497) & (g1498) & (g1516) & (!g1568)) + ((!g803) & (!g851) & (g1497) & (!g1498) & (!g1516) & (!g1568)) + ((!g803) & (!g851) & (g1497) & (!g1498) & (!g1516) & (g1568)) + ((!g803) & (!g851) & (g1497) & (!g1498) & (g1516) & (!g1568)) + ((!g803) & (!g851) & (g1497) & (!g1498) & (g1516) & (g1568)) + ((!g803) & (!g851) & (g1497) & (g1498) & (!g1516) & (!g1568)) + ((!g803) & (!g851) & (g1497) & (g1498) & (!g1516) & (g1568)) + ((!g803) & (!g851) & (g1497) & (g1498) & (g1516) & (g1568)) + ((!g803) & (g851) & (!g1497) & (!g1498) & (g1516) & (!g1568)) + ((!g803) & (g851) & (!g1497) & (g1498) & (!g1516) & (!g1568)) + ((!g803) & (g851) & (!g1497) & (g1498) & (g1516) & (!g1568)) + ((!g803) & (g851) & (g1497) & (!g1498) & (!g1516) & (!g1568)) + ((!g803) & (g851) & (g1497) & (!g1498) & (!g1516) & (g1568)) + ((!g803) & (g851) & (g1497) & (!g1498) & (g1516) & (g1568)) + ((!g803) & (g851) & (g1497) & (g1498) & (!g1516) & (g1568)) + ((!g803) & (g851) & (g1497) & (g1498) & (g1516) & (g1568)) + ((g803) & (!g851) & (!g1497) & (!g1498) & (!g1516) & (!g1568)) + ((g803) & (!g851) & (!g1497) & (!g1498) & (g1516) & (!g1568)) + ((g803) & (!g851) & (!g1497) & (g1498) & (!g1516) & (!g1568)) + ((g803) & (!g851) & (g1497) & (!g1498) & (!g1516) & (g1568)) + ((g803) & (!g851) & (g1497) & (!g1498) & (g1516) & (g1568)) + ((g803) & (!g851) & (g1497) & (g1498) & (!g1516) & (g1568)) + ((g803) & (!g851) & (g1497) & (g1498) & (g1516) & (!g1568)) + ((g803) & (!g851) & (g1497) & (g1498) & (g1516) & (g1568)) + ((g803) & (g851) & (!g1497) & (!g1498) & (!g1516) & (!g1568)) + ((g803) & (g851) & (g1497) & (!g1498) & (!g1516) & (g1568)) + ((g803) & (g851) & (g1497) & (!g1498) & (g1516) & (!g1568)) + ((g803) & (g851) & (g1497) & (!g1498) & (g1516) & (g1568)) + ((g803) & (g851) & (g1497) & (g1498) & (!g1516) & (!g1568)) + ((g803) & (g851) & (g1497) & (g1498) & (!g1516) & (g1568)) + ((g803) & (g851) & (g1497) & (g1498) & (g1516) & (!g1568)) + ((g803) & (g851) & (g1497) & (g1498) & (g1516) & (g1568)));
	assign g1577 = (((!g851) & (!g1498) & (g1516) & (!g1568)) + ((!g851) & (g1498) & (!g1516) & (!g1568)) + ((!g851) & (g1498) & (!g1516) & (g1568)) + ((!g851) & (g1498) & (g1516) & (g1568)) + ((g851) & (!g1498) & (!g1516) & (!g1568)) + ((g851) & (g1498) & (!g1516) & (g1568)) + ((g851) & (g1498) & (g1516) & (!g1568)) + ((g851) & (g1498) & (g1516) & (g1568)));
	assign g1578 = (((!g914) & (!g1032) & (!g1500) & (g1501) & (g1515) & (!g1568)) + ((!g914) & (!g1032) & (g1500) & (!g1501) & (!g1515) & (!g1568)) + ((!g914) & (!g1032) & (g1500) & (!g1501) & (!g1515) & (g1568)) + ((!g914) & (!g1032) & (g1500) & (!g1501) & (g1515) & (!g1568)) + ((!g914) & (!g1032) & (g1500) & (!g1501) & (g1515) & (g1568)) + ((!g914) & (!g1032) & (g1500) & (g1501) & (!g1515) & (!g1568)) + ((!g914) & (!g1032) & (g1500) & (g1501) & (!g1515) & (g1568)) + ((!g914) & (!g1032) & (g1500) & (g1501) & (g1515) & (g1568)) + ((!g914) & (g1032) & (!g1500) & (!g1501) & (g1515) & (!g1568)) + ((!g914) & (g1032) & (!g1500) & (g1501) & (!g1515) & (!g1568)) + ((!g914) & (g1032) & (!g1500) & (g1501) & (g1515) & (!g1568)) + ((!g914) & (g1032) & (g1500) & (!g1501) & (!g1515) & (!g1568)) + ((!g914) & (g1032) & (g1500) & (!g1501) & (!g1515) & (g1568)) + ((!g914) & (g1032) & (g1500) & (!g1501) & (g1515) & (g1568)) + ((!g914) & (g1032) & (g1500) & (g1501) & (!g1515) & (g1568)) + ((!g914) & (g1032) & (g1500) & (g1501) & (g1515) & (g1568)) + ((g914) & (!g1032) & (!g1500) & (!g1501) & (!g1515) & (!g1568)) + ((g914) & (!g1032) & (!g1500) & (!g1501) & (g1515) & (!g1568)) + ((g914) & (!g1032) & (!g1500) & (g1501) & (!g1515) & (!g1568)) + ((g914) & (!g1032) & (g1500) & (!g1501) & (!g1515) & (g1568)) + ((g914) & (!g1032) & (g1500) & (!g1501) & (g1515) & (g1568)) + ((g914) & (!g1032) & (g1500) & (g1501) & (!g1515) & (g1568)) + ((g914) & (!g1032) & (g1500) & (g1501) & (g1515) & (!g1568)) + ((g914) & (!g1032) & (g1500) & (g1501) & (g1515) & (g1568)) + ((g914) & (g1032) & (!g1500) & (!g1501) & (!g1515) & (!g1568)) + ((g914) & (g1032) & (g1500) & (!g1501) & (!g1515) & (g1568)) + ((g914) & (g1032) & (g1500) & (!g1501) & (g1515) & (!g1568)) + ((g914) & (g1032) & (g1500) & (!g1501) & (g1515) & (g1568)) + ((g914) & (g1032) & (g1500) & (g1501) & (!g1515) & (!g1568)) + ((g914) & (g1032) & (g1500) & (g1501) & (!g1515) & (g1568)) + ((g914) & (g1032) & (g1500) & (g1501) & (g1515) & (!g1568)) + ((g914) & (g1032) & (g1500) & (g1501) & (g1515) & (g1568)));
	assign g1579 = (((!g1032) & (!g1501) & (g1515) & (!g1568)) + ((!g1032) & (g1501) & (!g1515) & (!g1568)) + ((!g1032) & (g1501) & (!g1515) & (g1568)) + ((!g1032) & (g1501) & (g1515) & (g1568)) + ((g1032) & (!g1501) & (!g1515) & (!g1568)) + ((g1032) & (g1501) & (!g1515) & (g1568)) + ((g1032) & (g1501) & (g1515) & (!g1568)) + ((g1032) & (g1501) & (g1515) & (g1568)));
	assign g1580 = (((!g1030) & (!g1160) & (!g1503) & (g1504) & (g1514) & (!g1568)) + ((!g1030) & (!g1160) & (g1503) & (!g1504) & (!g1514) & (!g1568)) + ((!g1030) & (!g1160) & (g1503) & (!g1504) & (!g1514) & (g1568)) + ((!g1030) & (!g1160) & (g1503) & (!g1504) & (g1514) & (!g1568)) + ((!g1030) & (!g1160) & (g1503) & (!g1504) & (g1514) & (g1568)) + ((!g1030) & (!g1160) & (g1503) & (g1504) & (!g1514) & (!g1568)) + ((!g1030) & (!g1160) & (g1503) & (g1504) & (!g1514) & (g1568)) + ((!g1030) & (!g1160) & (g1503) & (g1504) & (g1514) & (g1568)) + ((!g1030) & (g1160) & (!g1503) & (!g1504) & (g1514) & (!g1568)) + ((!g1030) & (g1160) & (!g1503) & (g1504) & (!g1514) & (!g1568)) + ((!g1030) & (g1160) & (!g1503) & (g1504) & (g1514) & (!g1568)) + ((!g1030) & (g1160) & (g1503) & (!g1504) & (!g1514) & (!g1568)) + ((!g1030) & (g1160) & (g1503) & (!g1504) & (!g1514) & (g1568)) + ((!g1030) & (g1160) & (g1503) & (!g1504) & (g1514) & (g1568)) + ((!g1030) & (g1160) & (g1503) & (g1504) & (!g1514) & (g1568)) + ((!g1030) & (g1160) & (g1503) & (g1504) & (g1514) & (g1568)) + ((g1030) & (!g1160) & (!g1503) & (!g1504) & (!g1514) & (!g1568)) + ((g1030) & (!g1160) & (!g1503) & (!g1504) & (g1514) & (!g1568)) + ((g1030) & (!g1160) & (!g1503) & (g1504) & (!g1514) & (!g1568)) + ((g1030) & (!g1160) & (g1503) & (!g1504) & (!g1514) & (g1568)) + ((g1030) & (!g1160) & (g1503) & (!g1504) & (g1514) & (g1568)) + ((g1030) & (!g1160) & (g1503) & (g1504) & (!g1514) & (g1568)) + ((g1030) & (!g1160) & (g1503) & (g1504) & (g1514) & (!g1568)) + ((g1030) & (!g1160) & (g1503) & (g1504) & (g1514) & (g1568)) + ((g1030) & (g1160) & (!g1503) & (!g1504) & (!g1514) & (!g1568)) + ((g1030) & (g1160) & (g1503) & (!g1504) & (!g1514) & (g1568)) + ((g1030) & (g1160) & (g1503) & (!g1504) & (g1514) & (!g1568)) + ((g1030) & (g1160) & (g1503) & (!g1504) & (g1514) & (g1568)) + ((g1030) & (g1160) & (g1503) & (g1504) & (!g1514) & (!g1568)) + ((g1030) & (g1160) & (g1503) & (g1504) & (!g1514) & (g1568)) + ((g1030) & (g1160) & (g1503) & (g1504) & (g1514) & (!g1568)) + ((g1030) & (g1160) & (g1503) & (g1504) & (g1514) & (g1568)));
	assign g1581 = (((!g1160) & (!g1504) & (g1514) & (!g1568)) + ((!g1160) & (g1504) & (!g1514) & (!g1568)) + ((!g1160) & (g1504) & (!g1514) & (g1568)) + ((!g1160) & (g1504) & (g1514) & (g1568)) + ((g1160) & (!g1504) & (!g1514) & (!g1568)) + ((g1160) & (g1504) & (!g1514) & (g1568)) + ((g1160) & (g1504) & (g1514) & (!g1568)) + ((g1160) & (g1504) & (g1514) & (g1568)));
	assign g1582 = (((!g1154) & (!g1295) & (!g1506) & (g1507) & (g1513) & (!g1568)) + ((!g1154) & (!g1295) & (g1506) & (!g1507) & (!g1513) & (!g1568)) + ((!g1154) & (!g1295) & (g1506) & (!g1507) & (!g1513) & (g1568)) + ((!g1154) & (!g1295) & (g1506) & (!g1507) & (g1513) & (!g1568)) + ((!g1154) & (!g1295) & (g1506) & (!g1507) & (g1513) & (g1568)) + ((!g1154) & (!g1295) & (g1506) & (g1507) & (!g1513) & (!g1568)) + ((!g1154) & (!g1295) & (g1506) & (g1507) & (!g1513) & (g1568)) + ((!g1154) & (!g1295) & (g1506) & (g1507) & (g1513) & (g1568)) + ((!g1154) & (g1295) & (!g1506) & (!g1507) & (g1513) & (!g1568)) + ((!g1154) & (g1295) & (!g1506) & (g1507) & (!g1513) & (!g1568)) + ((!g1154) & (g1295) & (!g1506) & (g1507) & (g1513) & (!g1568)) + ((!g1154) & (g1295) & (g1506) & (!g1507) & (!g1513) & (!g1568)) + ((!g1154) & (g1295) & (g1506) & (!g1507) & (!g1513) & (g1568)) + ((!g1154) & (g1295) & (g1506) & (!g1507) & (g1513) & (g1568)) + ((!g1154) & (g1295) & (g1506) & (g1507) & (!g1513) & (g1568)) + ((!g1154) & (g1295) & (g1506) & (g1507) & (g1513) & (g1568)) + ((g1154) & (!g1295) & (!g1506) & (!g1507) & (!g1513) & (!g1568)) + ((g1154) & (!g1295) & (!g1506) & (!g1507) & (g1513) & (!g1568)) + ((g1154) & (!g1295) & (!g1506) & (g1507) & (!g1513) & (!g1568)) + ((g1154) & (!g1295) & (g1506) & (!g1507) & (!g1513) & (g1568)) + ((g1154) & (!g1295) & (g1506) & (!g1507) & (g1513) & (g1568)) + ((g1154) & (!g1295) & (g1506) & (g1507) & (!g1513) & (g1568)) + ((g1154) & (!g1295) & (g1506) & (g1507) & (g1513) & (!g1568)) + ((g1154) & (!g1295) & (g1506) & (g1507) & (g1513) & (g1568)) + ((g1154) & (g1295) & (!g1506) & (!g1507) & (!g1513) & (!g1568)) + ((g1154) & (g1295) & (g1506) & (!g1507) & (!g1513) & (g1568)) + ((g1154) & (g1295) & (g1506) & (!g1507) & (g1513) & (!g1568)) + ((g1154) & (g1295) & (g1506) & (!g1507) & (g1513) & (g1568)) + ((g1154) & (g1295) & (g1506) & (g1507) & (!g1513) & (!g1568)) + ((g1154) & (g1295) & (g1506) & (g1507) & (!g1513) & (g1568)) + ((g1154) & (g1295) & (g1506) & (g1507) & (g1513) & (!g1568)) + ((g1154) & (g1295) & (g1506) & (g1507) & (g1513) & (g1568)));
	assign g1583 = (((!g1295) & (!g1507) & (g1513) & (!g1568)) + ((!g1295) & (g1507) & (!g1513) & (!g1568)) + ((!g1295) & (g1507) & (!g1513) & (g1568)) + ((!g1295) & (g1507) & (g1513) & (g1568)) + ((g1295) & (!g1507) & (!g1513) & (!g1568)) + ((g1295) & (g1507) & (!g1513) & (g1568)) + ((g1295) & (g1507) & (g1513) & (!g1568)) + ((g1295) & (g1507) & (g1513) & (g1568)));
	assign g1584 = (((!g1285) & (!g1437) & (!g1509) & (g1510) & (g1512) & (!g1568)) + ((!g1285) & (!g1437) & (g1509) & (!g1510) & (!g1512) & (!g1568)) + ((!g1285) & (!g1437) & (g1509) & (!g1510) & (!g1512) & (g1568)) + ((!g1285) & (!g1437) & (g1509) & (!g1510) & (g1512) & (!g1568)) + ((!g1285) & (!g1437) & (g1509) & (!g1510) & (g1512) & (g1568)) + ((!g1285) & (!g1437) & (g1509) & (g1510) & (!g1512) & (!g1568)) + ((!g1285) & (!g1437) & (g1509) & (g1510) & (!g1512) & (g1568)) + ((!g1285) & (!g1437) & (g1509) & (g1510) & (g1512) & (g1568)) + ((!g1285) & (g1437) & (!g1509) & (!g1510) & (g1512) & (!g1568)) + ((!g1285) & (g1437) & (!g1509) & (g1510) & (!g1512) & (!g1568)) + ((!g1285) & (g1437) & (!g1509) & (g1510) & (g1512) & (!g1568)) + ((!g1285) & (g1437) & (g1509) & (!g1510) & (!g1512) & (!g1568)) + ((!g1285) & (g1437) & (g1509) & (!g1510) & (!g1512) & (g1568)) + ((!g1285) & (g1437) & (g1509) & (!g1510) & (g1512) & (g1568)) + ((!g1285) & (g1437) & (g1509) & (g1510) & (!g1512) & (g1568)) + ((!g1285) & (g1437) & (g1509) & (g1510) & (g1512) & (g1568)) + ((g1285) & (!g1437) & (!g1509) & (!g1510) & (!g1512) & (!g1568)) + ((g1285) & (!g1437) & (!g1509) & (!g1510) & (g1512) & (!g1568)) + ((g1285) & (!g1437) & (!g1509) & (g1510) & (!g1512) & (!g1568)) + ((g1285) & (!g1437) & (g1509) & (!g1510) & (!g1512) & (g1568)) + ((g1285) & (!g1437) & (g1509) & (!g1510) & (g1512) & (g1568)) + ((g1285) & (!g1437) & (g1509) & (g1510) & (!g1512) & (g1568)) + ((g1285) & (!g1437) & (g1509) & (g1510) & (g1512) & (!g1568)) + ((g1285) & (!g1437) & (g1509) & (g1510) & (g1512) & (g1568)) + ((g1285) & (g1437) & (!g1509) & (!g1510) & (!g1512) & (!g1568)) + ((g1285) & (g1437) & (g1509) & (!g1510) & (!g1512) & (g1568)) + ((g1285) & (g1437) & (g1509) & (!g1510) & (g1512) & (!g1568)) + ((g1285) & (g1437) & (g1509) & (!g1510) & (g1512) & (g1568)) + ((g1285) & (g1437) & (g1509) & (g1510) & (!g1512) & (!g1568)) + ((g1285) & (g1437) & (g1509) & (g1510) & (!g1512) & (g1568)) + ((g1285) & (g1437) & (g1509) & (g1510) & (g1512) & (!g1568)) + ((g1285) & (g1437) & (g1509) & (g1510) & (g1512) & (g1568)));
	assign g1585 = (((!g1437) & (!g1510) & (g1512) & (!g1568)) + ((!g1437) & (g1510) & (!g1512) & (!g1568)) + ((!g1437) & (g1510) & (!g1512) & (g1568)) + ((!g1437) & (g1510) & (g1512) & (g1568)) + ((g1437) & (!g1510) & (!g1512) & (!g1568)) + ((g1437) & (g1510) & (!g1512) & (g1568)) + ((g1437) & (g1510) & (g1512) & (!g1568)) + ((g1437) & (g1510) & (g1512) & (g1568)));
	assign g1586 = (((!g1449) & (g1485)));
	assign g1587 = (((!g1423) & (!ax46x) & (!ax47x) & (!g1586) & (!g1511) & (g1568)) + ((!g1423) & (!ax46x) & (!ax47x) & (!g1586) & (g1511) & (!g1568)) + ((!g1423) & (!ax46x) & (!ax47x) & (!g1586) & (g1511) & (g1568)) + ((!g1423) & (!ax46x) & (!ax47x) & (g1586) & (!g1511) & (!g1568)) + ((!g1423) & (!ax46x) & (ax47x) & (!g1586) & (!g1511) & (!g1568)) + ((!g1423) & (!ax46x) & (ax47x) & (g1586) & (!g1511) & (g1568)) + ((!g1423) & (!ax46x) & (ax47x) & (g1586) & (g1511) & (!g1568)) + ((!g1423) & (!ax46x) & (ax47x) & (g1586) & (g1511) & (g1568)) + ((!g1423) & (ax46x) & (!ax47x) & (g1586) & (!g1511) & (!g1568)) + ((!g1423) & (ax46x) & (!ax47x) & (g1586) & (g1511) & (!g1568)) + ((!g1423) & (ax46x) & (ax47x) & (!g1586) & (!g1511) & (!g1568)) + ((!g1423) & (ax46x) & (ax47x) & (!g1586) & (!g1511) & (g1568)) + ((!g1423) & (ax46x) & (ax47x) & (!g1586) & (g1511) & (!g1568)) + ((!g1423) & (ax46x) & (ax47x) & (!g1586) & (g1511) & (g1568)) + ((!g1423) & (ax46x) & (ax47x) & (g1586) & (!g1511) & (g1568)) + ((!g1423) & (ax46x) & (ax47x) & (g1586) & (g1511) & (g1568)) + ((g1423) & (!ax46x) & (!ax47x) & (!g1586) & (!g1511) & (!g1568)) + ((g1423) & (!ax46x) & (!ax47x) & (!g1586) & (!g1511) & (g1568)) + ((g1423) & (!ax46x) & (!ax47x) & (!g1586) & (g1511) & (g1568)) + ((g1423) & (!ax46x) & (!ax47x) & (g1586) & (g1511) & (!g1568)) + ((g1423) & (!ax46x) & (ax47x) & (!g1586) & (g1511) & (!g1568)) + ((g1423) & (!ax46x) & (ax47x) & (g1586) & (!g1511) & (!g1568)) + ((g1423) & (!ax46x) & (ax47x) & (g1586) & (!g1511) & (g1568)) + ((g1423) & (!ax46x) & (ax47x) & (g1586) & (g1511) & (g1568)) + ((g1423) & (ax46x) & (!ax47x) & (!g1586) & (!g1511) & (!g1568)) + ((g1423) & (ax46x) & (!ax47x) & (!g1586) & (g1511) & (!g1568)) + ((g1423) & (ax46x) & (ax47x) & (!g1586) & (!g1511) & (g1568)) + ((g1423) & (ax46x) & (ax47x) & (!g1586) & (g1511) & (g1568)) + ((g1423) & (ax46x) & (ax47x) & (g1586) & (!g1511) & (!g1568)) + ((g1423) & (ax46x) & (ax47x) & (g1586) & (!g1511) & (g1568)) + ((g1423) & (ax46x) & (ax47x) & (g1586) & (g1511) & (!g1568)) + ((g1423) & (ax46x) & (ax47x) & (g1586) & (g1511) & (g1568)));
	assign g1588 = (((!ax46x) & (!g1586) & (!g1511) & (g1568)) + ((!ax46x) & (!g1586) & (g1511) & (!g1568)) + ((!ax46x) & (!g1586) & (g1511) & (g1568)) + ((!ax46x) & (g1586) & (g1511) & (!g1568)) + ((ax46x) & (!g1586) & (!g1511) & (!g1568)) + ((ax46x) & (g1586) & (!g1511) & (!g1568)) + ((ax46x) & (g1586) & (!g1511) & (g1568)) + ((ax46x) & (g1586) & (g1511) & (g1568)));
	assign g1589 = (((!ax42x) & (!ax43x)));
	assign g1590 = (((!g1586) & (!ax44x) & (!ax45x) & (!g1568) & (!g1589)) + ((!g1586) & (!ax44x) & (ax45x) & (g1568) & (!g1589)) + ((!g1586) & (ax44x) & (ax45x) & (g1568) & (!g1589)) + ((!g1586) & (ax44x) & (ax45x) & (g1568) & (g1589)) + ((g1586) & (!ax44x) & (!ax45x) & (!g1568) & (!g1589)) + ((g1586) & (!ax44x) & (!ax45x) & (!g1568) & (g1589)) + ((g1586) & (!ax44x) & (!ax45x) & (g1568) & (!g1589)) + ((g1586) & (!ax44x) & (ax45x) & (!g1568) & (!g1589)) + ((g1586) & (!ax44x) & (ax45x) & (g1568) & (!g1589)) + ((g1586) & (!ax44x) & (ax45x) & (g1568) & (g1589)) + ((g1586) & (ax44x) & (!ax45x) & (g1568) & (!g1589)) + ((g1586) & (ax44x) & (!ax45x) & (g1568) & (g1589)) + ((g1586) & (ax44x) & (ax45x) & (!g1568) & (!g1589)) + ((g1586) & (ax44x) & (ax45x) & (!g1568) & (g1589)) + ((g1586) & (ax44x) & (ax45x) & (g1568) & (!g1589)) + ((g1586) & (ax44x) & (ax45x) & (g1568) & (g1589)));
	assign g1591 = (((!g1437) & (!g1423) & (g1587) & (g1588) & (g1590)) + ((!g1437) & (g1423) & (g1587) & (!g1588) & (g1590)) + ((!g1437) & (g1423) & (g1587) & (g1588) & (!g1590)) + ((!g1437) & (g1423) & (g1587) & (g1588) & (g1590)) + ((g1437) & (!g1423) & (!g1587) & (g1588) & (g1590)) + ((g1437) & (!g1423) & (g1587) & (!g1588) & (!g1590)) + ((g1437) & (!g1423) & (g1587) & (!g1588) & (g1590)) + ((g1437) & (!g1423) & (g1587) & (g1588) & (!g1590)) + ((g1437) & (!g1423) & (g1587) & (g1588) & (g1590)) + ((g1437) & (g1423) & (!g1587) & (!g1588) & (g1590)) + ((g1437) & (g1423) & (!g1587) & (g1588) & (!g1590)) + ((g1437) & (g1423) & (!g1587) & (g1588) & (g1590)) + ((g1437) & (g1423) & (g1587) & (!g1588) & (!g1590)) + ((g1437) & (g1423) & (g1587) & (!g1588) & (g1590)) + ((g1437) & (g1423) & (g1587) & (g1588) & (!g1590)) + ((g1437) & (g1423) & (g1587) & (g1588) & (g1590)));
	assign g1592 = (((!g1295) & (!g1285) & (g1584) & (g1585) & (g1591)) + ((!g1295) & (g1285) & (g1584) & (!g1585) & (g1591)) + ((!g1295) & (g1285) & (g1584) & (g1585) & (!g1591)) + ((!g1295) & (g1285) & (g1584) & (g1585) & (g1591)) + ((g1295) & (!g1285) & (!g1584) & (g1585) & (g1591)) + ((g1295) & (!g1285) & (g1584) & (!g1585) & (!g1591)) + ((g1295) & (!g1285) & (g1584) & (!g1585) & (g1591)) + ((g1295) & (!g1285) & (g1584) & (g1585) & (!g1591)) + ((g1295) & (!g1285) & (g1584) & (g1585) & (g1591)) + ((g1295) & (g1285) & (!g1584) & (!g1585) & (g1591)) + ((g1295) & (g1285) & (!g1584) & (g1585) & (!g1591)) + ((g1295) & (g1285) & (!g1584) & (g1585) & (g1591)) + ((g1295) & (g1285) & (g1584) & (!g1585) & (!g1591)) + ((g1295) & (g1285) & (g1584) & (!g1585) & (g1591)) + ((g1295) & (g1285) & (g1584) & (g1585) & (!g1591)) + ((g1295) & (g1285) & (g1584) & (g1585) & (g1591)));
	assign g1593 = (((!g1160) & (!g1154) & (g1582) & (g1583) & (g1592)) + ((!g1160) & (g1154) & (g1582) & (!g1583) & (g1592)) + ((!g1160) & (g1154) & (g1582) & (g1583) & (!g1592)) + ((!g1160) & (g1154) & (g1582) & (g1583) & (g1592)) + ((g1160) & (!g1154) & (!g1582) & (g1583) & (g1592)) + ((g1160) & (!g1154) & (g1582) & (!g1583) & (!g1592)) + ((g1160) & (!g1154) & (g1582) & (!g1583) & (g1592)) + ((g1160) & (!g1154) & (g1582) & (g1583) & (!g1592)) + ((g1160) & (!g1154) & (g1582) & (g1583) & (g1592)) + ((g1160) & (g1154) & (!g1582) & (!g1583) & (g1592)) + ((g1160) & (g1154) & (!g1582) & (g1583) & (!g1592)) + ((g1160) & (g1154) & (!g1582) & (g1583) & (g1592)) + ((g1160) & (g1154) & (g1582) & (!g1583) & (!g1592)) + ((g1160) & (g1154) & (g1582) & (!g1583) & (g1592)) + ((g1160) & (g1154) & (g1582) & (g1583) & (!g1592)) + ((g1160) & (g1154) & (g1582) & (g1583) & (g1592)));
	assign g1594 = (((!g1032) & (!g1030) & (g1580) & (g1581) & (g1593)) + ((!g1032) & (g1030) & (g1580) & (!g1581) & (g1593)) + ((!g1032) & (g1030) & (g1580) & (g1581) & (!g1593)) + ((!g1032) & (g1030) & (g1580) & (g1581) & (g1593)) + ((g1032) & (!g1030) & (!g1580) & (g1581) & (g1593)) + ((g1032) & (!g1030) & (g1580) & (!g1581) & (!g1593)) + ((g1032) & (!g1030) & (g1580) & (!g1581) & (g1593)) + ((g1032) & (!g1030) & (g1580) & (g1581) & (!g1593)) + ((g1032) & (!g1030) & (g1580) & (g1581) & (g1593)) + ((g1032) & (g1030) & (!g1580) & (!g1581) & (g1593)) + ((g1032) & (g1030) & (!g1580) & (g1581) & (!g1593)) + ((g1032) & (g1030) & (!g1580) & (g1581) & (g1593)) + ((g1032) & (g1030) & (g1580) & (!g1581) & (!g1593)) + ((g1032) & (g1030) & (g1580) & (!g1581) & (g1593)) + ((g1032) & (g1030) & (g1580) & (g1581) & (!g1593)) + ((g1032) & (g1030) & (g1580) & (g1581) & (g1593)));
	assign g1595 = (((!g851) & (!g914) & (g1578) & (g1579) & (g1594)) + ((!g851) & (g914) & (g1578) & (!g1579) & (g1594)) + ((!g851) & (g914) & (g1578) & (g1579) & (!g1594)) + ((!g851) & (g914) & (g1578) & (g1579) & (g1594)) + ((g851) & (!g914) & (!g1578) & (g1579) & (g1594)) + ((g851) & (!g914) & (g1578) & (!g1579) & (!g1594)) + ((g851) & (!g914) & (g1578) & (!g1579) & (g1594)) + ((g851) & (!g914) & (g1578) & (g1579) & (!g1594)) + ((g851) & (!g914) & (g1578) & (g1579) & (g1594)) + ((g851) & (g914) & (!g1578) & (!g1579) & (g1594)) + ((g851) & (g914) & (!g1578) & (g1579) & (!g1594)) + ((g851) & (g914) & (!g1578) & (g1579) & (g1594)) + ((g851) & (g914) & (g1578) & (!g1579) & (!g1594)) + ((g851) & (g914) & (g1578) & (!g1579) & (g1594)) + ((g851) & (g914) & (g1578) & (g1579) & (!g1594)) + ((g851) & (g914) & (g1578) & (g1579) & (g1594)));
	assign g1596 = (((!g744) & (!g803) & (g1576) & (g1577) & (g1595)) + ((!g744) & (g803) & (g1576) & (!g1577) & (g1595)) + ((!g744) & (g803) & (g1576) & (g1577) & (!g1595)) + ((!g744) & (g803) & (g1576) & (g1577) & (g1595)) + ((g744) & (!g803) & (!g1576) & (g1577) & (g1595)) + ((g744) & (!g803) & (g1576) & (!g1577) & (!g1595)) + ((g744) & (!g803) & (g1576) & (!g1577) & (g1595)) + ((g744) & (!g803) & (g1576) & (g1577) & (!g1595)) + ((g744) & (!g803) & (g1576) & (g1577) & (g1595)) + ((g744) & (g803) & (!g1576) & (!g1577) & (g1595)) + ((g744) & (g803) & (!g1576) & (g1577) & (!g1595)) + ((g744) & (g803) & (!g1576) & (g1577) & (g1595)) + ((g744) & (g803) & (g1576) & (!g1577) & (!g1595)) + ((g744) & (g803) & (g1576) & (!g1577) & (g1595)) + ((g744) & (g803) & (g1576) & (g1577) & (!g1595)) + ((g744) & (g803) & (g1576) & (g1577) & (g1595)));
	assign g1597 = (((!g645) & (!g700) & (g1574) & (g1575) & (g1596)) + ((!g645) & (g700) & (g1574) & (!g1575) & (g1596)) + ((!g645) & (g700) & (g1574) & (g1575) & (!g1596)) + ((!g645) & (g700) & (g1574) & (g1575) & (g1596)) + ((g645) & (!g700) & (!g1574) & (g1575) & (g1596)) + ((g645) & (!g700) & (g1574) & (!g1575) & (!g1596)) + ((g645) & (!g700) & (g1574) & (!g1575) & (g1596)) + ((g645) & (!g700) & (g1574) & (g1575) & (!g1596)) + ((g645) & (!g700) & (g1574) & (g1575) & (g1596)) + ((g645) & (g700) & (!g1574) & (!g1575) & (g1596)) + ((g645) & (g700) & (!g1574) & (g1575) & (!g1596)) + ((g645) & (g700) & (!g1574) & (g1575) & (g1596)) + ((g645) & (g700) & (g1574) & (!g1575) & (!g1596)) + ((g645) & (g700) & (g1574) & (!g1575) & (g1596)) + ((g645) & (g700) & (g1574) & (g1575) & (!g1596)) + ((g645) & (g700) & (g1574) & (g1575) & (g1596)));
	assign g1598 = (((!g553) & (!g604) & (g1572) & (g1573) & (g1597)) + ((!g553) & (g604) & (g1572) & (!g1573) & (g1597)) + ((!g553) & (g604) & (g1572) & (g1573) & (!g1597)) + ((!g553) & (g604) & (g1572) & (g1573) & (g1597)) + ((g553) & (!g604) & (!g1572) & (g1573) & (g1597)) + ((g553) & (!g604) & (g1572) & (!g1573) & (!g1597)) + ((g553) & (!g604) & (g1572) & (!g1573) & (g1597)) + ((g553) & (!g604) & (g1572) & (g1573) & (!g1597)) + ((g553) & (!g604) & (g1572) & (g1573) & (g1597)) + ((g553) & (g604) & (!g1572) & (!g1573) & (g1597)) + ((g553) & (g604) & (!g1572) & (g1573) & (!g1597)) + ((g553) & (g604) & (!g1572) & (g1573) & (g1597)) + ((g553) & (g604) & (g1572) & (!g1573) & (!g1597)) + ((g553) & (g604) & (g1572) & (!g1573) & (g1597)) + ((g553) & (g604) & (g1572) & (g1573) & (!g1597)) + ((g553) & (g604) & (g1572) & (g1573) & (g1597)));
	assign g1599 = (((!g468) & (!g515) & (g1570) & (g1571) & (g1598)) + ((!g468) & (g515) & (g1570) & (!g1571) & (g1598)) + ((!g468) & (g515) & (g1570) & (g1571) & (!g1598)) + ((!g468) & (g515) & (g1570) & (g1571) & (g1598)) + ((g468) & (!g515) & (!g1570) & (g1571) & (g1598)) + ((g468) & (!g515) & (g1570) & (!g1571) & (!g1598)) + ((g468) & (!g515) & (g1570) & (!g1571) & (g1598)) + ((g468) & (!g515) & (g1570) & (g1571) & (!g1598)) + ((g468) & (!g515) & (g1570) & (g1571) & (g1598)) + ((g468) & (g515) & (!g1570) & (!g1571) & (g1598)) + ((g468) & (g515) & (!g1570) & (g1571) & (!g1598)) + ((g468) & (g515) & (!g1570) & (g1571) & (g1598)) + ((g468) & (g515) & (g1570) & (!g1571) & (!g1598)) + ((g468) & (g515) & (g1570) & (!g1571) & (g1598)) + ((g468) & (g515) & (g1570) & (g1571) & (!g1598)) + ((g468) & (g515) & (g1570) & (g1571) & (g1598)));
	assign g1600 = (((g1) & (!g1521) & (g1564) & (g1567)) + ((g1) & (g1521) & (!g1564) & (!g1567)) + ((g1) & (g1521) & (!g1564) & (g1567)));
	assign g1601 = (((!g4) & (!g2) & (!g1522) & (!g1561) & (!g1563) & (!g1568)) + ((!g4) & (!g2) & (!g1522) & (!g1561) & (g1563) & (g1568)) + ((!g4) & (!g2) & (!g1522) & (g1561) & (!g1563) & (!g1568)) + ((!g4) & (!g2) & (!g1522) & (g1561) & (g1563) & (g1568)) + ((!g4) & (!g2) & (g1522) & (!g1561) & (!g1563) & (!g1568)) + ((!g4) & (!g2) & (g1522) & (!g1561) & (g1563) & (g1568)) + ((!g4) & (!g2) & (g1522) & (g1561) & (g1563) & (!g1568)) + ((!g4) & (!g2) & (g1522) & (g1561) & (g1563) & (g1568)) + ((!g4) & (g2) & (!g1522) & (!g1561) & (!g1563) & (!g1568)) + ((!g4) & (g2) & (!g1522) & (!g1561) & (g1563) & (g1568)) + ((!g4) & (g2) & (!g1522) & (g1561) & (g1563) & (!g1568)) + ((!g4) & (g2) & (!g1522) & (g1561) & (g1563) & (g1568)) + ((!g4) & (g2) & (g1522) & (!g1561) & (g1563) & (!g1568)) + ((!g4) & (g2) & (g1522) & (!g1561) & (g1563) & (g1568)) + ((!g4) & (g2) & (g1522) & (g1561) & (g1563) & (!g1568)) + ((!g4) & (g2) & (g1522) & (g1561) & (g1563) & (g1568)) + ((g4) & (!g2) & (!g1522) & (!g1561) & (g1563) & (!g1568)) + ((g4) & (!g2) & (!g1522) & (!g1561) & (g1563) & (g1568)) + ((g4) & (!g2) & (!g1522) & (g1561) & (g1563) & (!g1568)) + ((g4) & (!g2) & (!g1522) & (g1561) & (g1563) & (g1568)) + ((g4) & (!g2) & (g1522) & (!g1561) & (g1563) & (!g1568)) + ((g4) & (!g2) & (g1522) & (!g1561) & (g1563) & (g1568)) + ((g4) & (!g2) & (g1522) & (g1561) & (!g1563) & (!g1568)) + ((g4) & (!g2) & (g1522) & (g1561) & (g1563) & (g1568)) + ((g4) & (g2) & (!g1522) & (!g1561) & (g1563) & (!g1568)) + ((g4) & (g2) & (!g1522) & (!g1561) & (g1563) & (g1568)) + ((g4) & (g2) & (!g1522) & (g1561) & (!g1563) & (!g1568)) + ((g4) & (g2) & (!g1522) & (g1561) & (g1563) & (g1568)) + ((g4) & (g2) & (g1522) & (!g1561) & (!g1563) & (!g1568)) + ((g4) & (g2) & (g1522) & (!g1561) & (g1563) & (g1568)) + ((g4) & (g2) & (g1522) & (g1561) & (!g1563) & (!g1568)) + ((g4) & (g2) & (g1522) & (g1561) & (g1563) & (g1568)));
	assign g1602 = (((!g8) & (!g18) & (!g1524) & (g1525) & (g1560) & (!g1568)) + ((!g8) & (!g18) & (g1524) & (!g1525) & (!g1560) & (!g1568)) + ((!g8) & (!g18) & (g1524) & (!g1525) & (!g1560) & (g1568)) + ((!g8) & (!g18) & (g1524) & (!g1525) & (g1560) & (!g1568)) + ((!g8) & (!g18) & (g1524) & (!g1525) & (g1560) & (g1568)) + ((!g8) & (!g18) & (g1524) & (g1525) & (!g1560) & (!g1568)) + ((!g8) & (!g18) & (g1524) & (g1525) & (!g1560) & (g1568)) + ((!g8) & (!g18) & (g1524) & (g1525) & (g1560) & (g1568)) + ((!g8) & (g18) & (!g1524) & (!g1525) & (g1560) & (!g1568)) + ((!g8) & (g18) & (!g1524) & (g1525) & (!g1560) & (!g1568)) + ((!g8) & (g18) & (!g1524) & (g1525) & (g1560) & (!g1568)) + ((!g8) & (g18) & (g1524) & (!g1525) & (!g1560) & (!g1568)) + ((!g8) & (g18) & (g1524) & (!g1525) & (!g1560) & (g1568)) + ((!g8) & (g18) & (g1524) & (!g1525) & (g1560) & (g1568)) + ((!g8) & (g18) & (g1524) & (g1525) & (!g1560) & (g1568)) + ((!g8) & (g18) & (g1524) & (g1525) & (g1560) & (g1568)) + ((g8) & (!g18) & (!g1524) & (!g1525) & (!g1560) & (!g1568)) + ((g8) & (!g18) & (!g1524) & (!g1525) & (g1560) & (!g1568)) + ((g8) & (!g18) & (!g1524) & (g1525) & (!g1560) & (!g1568)) + ((g8) & (!g18) & (g1524) & (!g1525) & (!g1560) & (g1568)) + ((g8) & (!g18) & (g1524) & (!g1525) & (g1560) & (g1568)) + ((g8) & (!g18) & (g1524) & (g1525) & (!g1560) & (g1568)) + ((g8) & (!g18) & (g1524) & (g1525) & (g1560) & (!g1568)) + ((g8) & (!g18) & (g1524) & (g1525) & (g1560) & (g1568)) + ((g8) & (g18) & (!g1524) & (!g1525) & (!g1560) & (!g1568)) + ((g8) & (g18) & (g1524) & (!g1525) & (!g1560) & (g1568)) + ((g8) & (g18) & (g1524) & (!g1525) & (g1560) & (!g1568)) + ((g8) & (g18) & (g1524) & (!g1525) & (g1560) & (g1568)) + ((g8) & (g18) & (g1524) & (g1525) & (!g1560) & (!g1568)) + ((g8) & (g18) & (g1524) & (g1525) & (!g1560) & (g1568)) + ((g8) & (g18) & (g1524) & (g1525) & (g1560) & (!g1568)) + ((g8) & (g18) & (g1524) & (g1525) & (g1560) & (g1568)));
	assign g1603 = (((!g18) & (!g1525) & (g1560) & (!g1568)) + ((!g18) & (g1525) & (!g1560) & (!g1568)) + ((!g18) & (g1525) & (!g1560) & (g1568)) + ((!g18) & (g1525) & (g1560) & (g1568)) + ((g18) & (!g1525) & (!g1560) & (!g1568)) + ((g18) & (g1525) & (!g1560) & (g1568)) + ((g18) & (g1525) & (g1560) & (!g1568)) + ((g18) & (g1525) & (g1560) & (g1568)));
	assign g1604 = (((!g27) & (!g39) & (!g1527) & (g1528) & (g1559) & (!g1568)) + ((!g27) & (!g39) & (g1527) & (!g1528) & (!g1559) & (!g1568)) + ((!g27) & (!g39) & (g1527) & (!g1528) & (!g1559) & (g1568)) + ((!g27) & (!g39) & (g1527) & (!g1528) & (g1559) & (!g1568)) + ((!g27) & (!g39) & (g1527) & (!g1528) & (g1559) & (g1568)) + ((!g27) & (!g39) & (g1527) & (g1528) & (!g1559) & (!g1568)) + ((!g27) & (!g39) & (g1527) & (g1528) & (!g1559) & (g1568)) + ((!g27) & (!g39) & (g1527) & (g1528) & (g1559) & (g1568)) + ((!g27) & (g39) & (!g1527) & (!g1528) & (g1559) & (!g1568)) + ((!g27) & (g39) & (!g1527) & (g1528) & (!g1559) & (!g1568)) + ((!g27) & (g39) & (!g1527) & (g1528) & (g1559) & (!g1568)) + ((!g27) & (g39) & (g1527) & (!g1528) & (!g1559) & (!g1568)) + ((!g27) & (g39) & (g1527) & (!g1528) & (!g1559) & (g1568)) + ((!g27) & (g39) & (g1527) & (!g1528) & (g1559) & (g1568)) + ((!g27) & (g39) & (g1527) & (g1528) & (!g1559) & (g1568)) + ((!g27) & (g39) & (g1527) & (g1528) & (g1559) & (g1568)) + ((g27) & (!g39) & (!g1527) & (!g1528) & (!g1559) & (!g1568)) + ((g27) & (!g39) & (!g1527) & (!g1528) & (g1559) & (!g1568)) + ((g27) & (!g39) & (!g1527) & (g1528) & (!g1559) & (!g1568)) + ((g27) & (!g39) & (g1527) & (!g1528) & (!g1559) & (g1568)) + ((g27) & (!g39) & (g1527) & (!g1528) & (g1559) & (g1568)) + ((g27) & (!g39) & (g1527) & (g1528) & (!g1559) & (g1568)) + ((g27) & (!g39) & (g1527) & (g1528) & (g1559) & (!g1568)) + ((g27) & (!g39) & (g1527) & (g1528) & (g1559) & (g1568)) + ((g27) & (g39) & (!g1527) & (!g1528) & (!g1559) & (!g1568)) + ((g27) & (g39) & (g1527) & (!g1528) & (!g1559) & (g1568)) + ((g27) & (g39) & (g1527) & (!g1528) & (g1559) & (!g1568)) + ((g27) & (g39) & (g1527) & (!g1528) & (g1559) & (g1568)) + ((g27) & (g39) & (g1527) & (g1528) & (!g1559) & (!g1568)) + ((g27) & (g39) & (g1527) & (g1528) & (!g1559) & (g1568)) + ((g27) & (g39) & (g1527) & (g1528) & (g1559) & (!g1568)) + ((g27) & (g39) & (g1527) & (g1528) & (g1559) & (g1568)));
	assign g1605 = (((!g39) & (!g1528) & (g1559) & (!g1568)) + ((!g39) & (g1528) & (!g1559) & (!g1568)) + ((!g39) & (g1528) & (!g1559) & (g1568)) + ((!g39) & (g1528) & (g1559) & (g1568)) + ((g39) & (!g1528) & (!g1559) & (!g1568)) + ((g39) & (g1528) & (!g1559) & (g1568)) + ((g39) & (g1528) & (g1559) & (!g1568)) + ((g39) & (g1528) & (g1559) & (g1568)));
	assign g1606 = (((!g54) & (!g68) & (!g1530) & (g1531) & (g1558) & (!g1568)) + ((!g54) & (!g68) & (g1530) & (!g1531) & (!g1558) & (!g1568)) + ((!g54) & (!g68) & (g1530) & (!g1531) & (!g1558) & (g1568)) + ((!g54) & (!g68) & (g1530) & (!g1531) & (g1558) & (!g1568)) + ((!g54) & (!g68) & (g1530) & (!g1531) & (g1558) & (g1568)) + ((!g54) & (!g68) & (g1530) & (g1531) & (!g1558) & (!g1568)) + ((!g54) & (!g68) & (g1530) & (g1531) & (!g1558) & (g1568)) + ((!g54) & (!g68) & (g1530) & (g1531) & (g1558) & (g1568)) + ((!g54) & (g68) & (!g1530) & (!g1531) & (g1558) & (!g1568)) + ((!g54) & (g68) & (!g1530) & (g1531) & (!g1558) & (!g1568)) + ((!g54) & (g68) & (!g1530) & (g1531) & (g1558) & (!g1568)) + ((!g54) & (g68) & (g1530) & (!g1531) & (!g1558) & (!g1568)) + ((!g54) & (g68) & (g1530) & (!g1531) & (!g1558) & (g1568)) + ((!g54) & (g68) & (g1530) & (!g1531) & (g1558) & (g1568)) + ((!g54) & (g68) & (g1530) & (g1531) & (!g1558) & (g1568)) + ((!g54) & (g68) & (g1530) & (g1531) & (g1558) & (g1568)) + ((g54) & (!g68) & (!g1530) & (!g1531) & (!g1558) & (!g1568)) + ((g54) & (!g68) & (!g1530) & (!g1531) & (g1558) & (!g1568)) + ((g54) & (!g68) & (!g1530) & (g1531) & (!g1558) & (!g1568)) + ((g54) & (!g68) & (g1530) & (!g1531) & (!g1558) & (g1568)) + ((g54) & (!g68) & (g1530) & (!g1531) & (g1558) & (g1568)) + ((g54) & (!g68) & (g1530) & (g1531) & (!g1558) & (g1568)) + ((g54) & (!g68) & (g1530) & (g1531) & (g1558) & (!g1568)) + ((g54) & (!g68) & (g1530) & (g1531) & (g1558) & (g1568)) + ((g54) & (g68) & (!g1530) & (!g1531) & (!g1558) & (!g1568)) + ((g54) & (g68) & (g1530) & (!g1531) & (!g1558) & (g1568)) + ((g54) & (g68) & (g1530) & (!g1531) & (g1558) & (!g1568)) + ((g54) & (g68) & (g1530) & (!g1531) & (g1558) & (g1568)) + ((g54) & (g68) & (g1530) & (g1531) & (!g1558) & (!g1568)) + ((g54) & (g68) & (g1530) & (g1531) & (!g1558) & (g1568)) + ((g54) & (g68) & (g1530) & (g1531) & (g1558) & (!g1568)) + ((g54) & (g68) & (g1530) & (g1531) & (g1558) & (g1568)));
	assign g1607 = (((!g68) & (!g1531) & (g1558) & (!g1568)) + ((!g68) & (g1531) & (!g1558) & (!g1568)) + ((!g68) & (g1531) & (!g1558) & (g1568)) + ((!g68) & (g1531) & (g1558) & (g1568)) + ((g68) & (!g1531) & (!g1558) & (!g1568)) + ((g68) & (g1531) & (!g1558) & (g1568)) + ((g68) & (g1531) & (g1558) & (!g1568)) + ((g68) & (g1531) & (g1558) & (g1568)));
	assign g1608 = (((!g87) & (!g104) & (!g1533) & (g1534) & (g1557) & (!g1568)) + ((!g87) & (!g104) & (g1533) & (!g1534) & (!g1557) & (!g1568)) + ((!g87) & (!g104) & (g1533) & (!g1534) & (!g1557) & (g1568)) + ((!g87) & (!g104) & (g1533) & (!g1534) & (g1557) & (!g1568)) + ((!g87) & (!g104) & (g1533) & (!g1534) & (g1557) & (g1568)) + ((!g87) & (!g104) & (g1533) & (g1534) & (!g1557) & (!g1568)) + ((!g87) & (!g104) & (g1533) & (g1534) & (!g1557) & (g1568)) + ((!g87) & (!g104) & (g1533) & (g1534) & (g1557) & (g1568)) + ((!g87) & (g104) & (!g1533) & (!g1534) & (g1557) & (!g1568)) + ((!g87) & (g104) & (!g1533) & (g1534) & (!g1557) & (!g1568)) + ((!g87) & (g104) & (!g1533) & (g1534) & (g1557) & (!g1568)) + ((!g87) & (g104) & (g1533) & (!g1534) & (!g1557) & (!g1568)) + ((!g87) & (g104) & (g1533) & (!g1534) & (!g1557) & (g1568)) + ((!g87) & (g104) & (g1533) & (!g1534) & (g1557) & (g1568)) + ((!g87) & (g104) & (g1533) & (g1534) & (!g1557) & (g1568)) + ((!g87) & (g104) & (g1533) & (g1534) & (g1557) & (g1568)) + ((g87) & (!g104) & (!g1533) & (!g1534) & (!g1557) & (!g1568)) + ((g87) & (!g104) & (!g1533) & (!g1534) & (g1557) & (!g1568)) + ((g87) & (!g104) & (!g1533) & (g1534) & (!g1557) & (!g1568)) + ((g87) & (!g104) & (g1533) & (!g1534) & (!g1557) & (g1568)) + ((g87) & (!g104) & (g1533) & (!g1534) & (g1557) & (g1568)) + ((g87) & (!g104) & (g1533) & (g1534) & (!g1557) & (g1568)) + ((g87) & (!g104) & (g1533) & (g1534) & (g1557) & (!g1568)) + ((g87) & (!g104) & (g1533) & (g1534) & (g1557) & (g1568)) + ((g87) & (g104) & (!g1533) & (!g1534) & (!g1557) & (!g1568)) + ((g87) & (g104) & (g1533) & (!g1534) & (!g1557) & (g1568)) + ((g87) & (g104) & (g1533) & (!g1534) & (g1557) & (!g1568)) + ((g87) & (g104) & (g1533) & (!g1534) & (g1557) & (g1568)) + ((g87) & (g104) & (g1533) & (g1534) & (!g1557) & (!g1568)) + ((g87) & (g104) & (g1533) & (g1534) & (!g1557) & (g1568)) + ((g87) & (g104) & (g1533) & (g1534) & (g1557) & (!g1568)) + ((g87) & (g104) & (g1533) & (g1534) & (g1557) & (g1568)));
	assign g1609 = (((!g104) & (!g1534) & (g1557) & (!g1568)) + ((!g104) & (g1534) & (!g1557) & (!g1568)) + ((!g104) & (g1534) & (!g1557) & (g1568)) + ((!g104) & (g1534) & (g1557) & (g1568)) + ((g104) & (!g1534) & (!g1557) & (!g1568)) + ((g104) & (g1534) & (!g1557) & (g1568)) + ((g104) & (g1534) & (g1557) & (!g1568)) + ((g104) & (g1534) & (g1557) & (g1568)));
	assign g1610 = (((!g127) & (!g147) & (!g1536) & (g1537) & (g1556) & (!g1568)) + ((!g127) & (!g147) & (g1536) & (!g1537) & (!g1556) & (!g1568)) + ((!g127) & (!g147) & (g1536) & (!g1537) & (!g1556) & (g1568)) + ((!g127) & (!g147) & (g1536) & (!g1537) & (g1556) & (!g1568)) + ((!g127) & (!g147) & (g1536) & (!g1537) & (g1556) & (g1568)) + ((!g127) & (!g147) & (g1536) & (g1537) & (!g1556) & (!g1568)) + ((!g127) & (!g147) & (g1536) & (g1537) & (!g1556) & (g1568)) + ((!g127) & (!g147) & (g1536) & (g1537) & (g1556) & (g1568)) + ((!g127) & (g147) & (!g1536) & (!g1537) & (g1556) & (!g1568)) + ((!g127) & (g147) & (!g1536) & (g1537) & (!g1556) & (!g1568)) + ((!g127) & (g147) & (!g1536) & (g1537) & (g1556) & (!g1568)) + ((!g127) & (g147) & (g1536) & (!g1537) & (!g1556) & (!g1568)) + ((!g127) & (g147) & (g1536) & (!g1537) & (!g1556) & (g1568)) + ((!g127) & (g147) & (g1536) & (!g1537) & (g1556) & (g1568)) + ((!g127) & (g147) & (g1536) & (g1537) & (!g1556) & (g1568)) + ((!g127) & (g147) & (g1536) & (g1537) & (g1556) & (g1568)) + ((g127) & (!g147) & (!g1536) & (!g1537) & (!g1556) & (!g1568)) + ((g127) & (!g147) & (!g1536) & (!g1537) & (g1556) & (!g1568)) + ((g127) & (!g147) & (!g1536) & (g1537) & (!g1556) & (!g1568)) + ((g127) & (!g147) & (g1536) & (!g1537) & (!g1556) & (g1568)) + ((g127) & (!g147) & (g1536) & (!g1537) & (g1556) & (g1568)) + ((g127) & (!g147) & (g1536) & (g1537) & (!g1556) & (g1568)) + ((g127) & (!g147) & (g1536) & (g1537) & (g1556) & (!g1568)) + ((g127) & (!g147) & (g1536) & (g1537) & (g1556) & (g1568)) + ((g127) & (g147) & (!g1536) & (!g1537) & (!g1556) & (!g1568)) + ((g127) & (g147) & (g1536) & (!g1537) & (!g1556) & (g1568)) + ((g127) & (g147) & (g1536) & (!g1537) & (g1556) & (!g1568)) + ((g127) & (g147) & (g1536) & (!g1537) & (g1556) & (g1568)) + ((g127) & (g147) & (g1536) & (g1537) & (!g1556) & (!g1568)) + ((g127) & (g147) & (g1536) & (g1537) & (!g1556) & (g1568)) + ((g127) & (g147) & (g1536) & (g1537) & (g1556) & (!g1568)) + ((g127) & (g147) & (g1536) & (g1537) & (g1556) & (g1568)));
	assign g1611 = (((!g147) & (!g1537) & (g1556) & (!g1568)) + ((!g147) & (g1537) & (!g1556) & (!g1568)) + ((!g147) & (g1537) & (!g1556) & (g1568)) + ((!g147) & (g1537) & (g1556) & (g1568)) + ((g147) & (!g1537) & (!g1556) & (!g1568)) + ((g147) & (g1537) & (!g1556) & (g1568)) + ((g147) & (g1537) & (g1556) & (!g1568)) + ((g147) & (g1537) & (g1556) & (g1568)));
	assign g1612 = (((!g174) & (!g198) & (!g1539) & (g1540) & (g1555) & (!g1568)) + ((!g174) & (!g198) & (g1539) & (!g1540) & (!g1555) & (!g1568)) + ((!g174) & (!g198) & (g1539) & (!g1540) & (!g1555) & (g1568)) + ((!g174) & (!g198) & (g1539) & (!g1540) & (g1555) & (!g1568)) + ((!g174) & (!g198) & (g1539) & (!g1540) & (g1555) & (g1568)) + ((!g174) & (!g198) & (g1539) & (g1540) & (!g1555) & (!g1568)) + ((!g174) & (!g198) & (g1539) & (g1540) & (!g1555) & (g1568)) + ((!g174) & (!g198) & (g1539) & (g1540) & (g1555) & (g1568)) + ((!g174) & (g198) & (!g1539) & (!g1540) & (g1555) & (!g1568)) + ((!g174) & (g198) & (!g1539) & (g1540) & (!g1555) & (!g1568)) + ((!g174) & (g198) & (!g1539) & (g1540) & (g1555) & (!g1568)) + ((!g174) & (g198) & (g1539) & (!g1540) & (!g1555) & (!g1568)) + ((!g174) & (g198) & (g1539) & (!g1540) & (!g1555) & (g1568)) + ((!g174) & (g198) & (g1539) & (!g1540) & (g1555) & (g1568)) + ((!g174) & (g198) & (g1539) & (g1540) & (!g1555) & (g1568)) + ((!g174) & (g198) & (g1539) & (g1540) & (g1555) & (g1568)) + ((g174) & (!g198) & (!g1539) & (!g1540) & (!g1555) & (!g1568)) + ((g174) & (!g198) & (!g1539) & (!g1540) & (g1555) & (!g1568)) + ((g174) & (!g198) & (!g1539) & (g1540) & (!g1555) & (!g1568)) + ((g174) & (!g198) & (g1539) & (!g1540) & (!g1555) & (g1568)) + ((g174) & (!g198) & (g1539) & (!g1540) & (g1555) & (g1568)) + ((g174) & (!g198) & (g1539) & (g1540) & (!g1555) & (g1568)) + ((g174) & (!g198) & (g1539) & (g1540) & (g1555) & (!g1568)) + ((g174) & (!g198) & (g1539) & (g1540) & (g1555) & (g1568)) + ((g174) & (g198) & (!g1539) & (!g1540) & (!g1555) & (!g1568)) + ((g174) & (g198) & (g1539) & (!g1540) & (!g1555) & (g1568)) + ((g174) & (g198) & (g1539) & (!g1540) & (g1555) & (!g1568)) + ((g174) & (g198) & (g1539) & (!g1540) & (g1555) & (g1568)) + ((g174) & (g198) & (g1539) & (g1540) & (!g1555) & (!g1568)) + ((g174) & (g198) & (g1539) & (g1540) & (!g1555) & (g1568)) + ((g174) & (g198) & (g1539) & (g1540) & (g1555) & (!g1568)) + ((g174) & (g198) & (g1539) & (g1540) & (g1555) & (g1568)));
	assign g1613 = (((!g198) & (!g1540) & (g1555) & (!g1568)) + ((!g198) & (g1540) & (!g1555) & (!g1568)) + ((!g198) & (g1540) & (!g1555) & (g1568)) + ((!g198) & (g1540) & (g1555) & (g1568)) + ((g198) & (!g1540) & (!g1555) & (!g1568)) + ((g198) & (g1540) & (!g1555) & (g1568)) + ((g198) & (g1540) & (g1555) & (!g1568)) + ((g198) & (g1540) & (g1555) & (g1568)));
	assign g1614 = (((!g229) & (!g255) & (!g1542) & (g1543) & (g1554) & (!g1568)) + ((!g229) & (!g255) & (g1542) & (!g1543) & (!g1554) & (!g1568)) + ((!g229) & (!g255) & (g1542) & (!g1543) & (!g1554) & (g1568)) + ((!g229) & (!g255) & (g1542) & (!g1543) & (g1554) & (!g1568)) + ((!g229) & (!g255) & (g1542) & (!g1543) & (g1554) & (g1568)) + ((!g229) & (!g255) & (g1542) & (g1543) & (!g1554) & (!g1568)) + ((!g229) & (!g255) & (g1542) & (g1543) & (!g1554) & (g1568)) + ((!g229) & (!g255) & (g1542) & (g1543) & (g1554) & (g1568)) + ((!g229) & (g255) & (!g1542) & (!g1543) & (g1554) & (!g1568)) + ((!g229) & (g255) & (!g1542) & (g1543) & (!g1554) & (!g1568)) + ((!g229) & (g255) & (!g1542) & (g1543) & (g1554) & (!g1568)) + ((!g229) & (g255) & (g1542) & (!g1543) & (!g1554) & (!g1568)) + ((!g229) & (g255) & (g1542) & (!g1543) & (!g1554) & (g1568)) + ((!g229) & (g255) & (g1542) & (!g1543) & (g1554) & (g1568)) + ((!g229) & (g255) & (g1542) & (g1543) & (!g1554) & (g1568)) + ((!g229) & (g255) & (g1542) & (g1543) & (g1554) & (g1568)) + ((g229) & (!g255) & (!g1542) & (!g1543) & (!g1554) & (!g1568)) + ((g229) & (!g255) & (!g1542) & (!g1543) & (g1554) & (!g1568)) + ((g229) & (!g255) & (!g1542) & (g1543) & (!g1554) & (!g1568)) + ((g229) & (!g255) & (g1542) & (!g1543) & (!g1554) & (g1568)) + ((g229) & (!g255) & (g1542) & (!g1543) & (g1554) & (g1568)) + ((g229) & (!g255) & (g1542) & (g1543) & (!g1554) & (g1568)) + ((g229) & (!g255) & (g1542) & (g1543) & (g1554) & (!g1568)) + ((g229) & (!g255) & (g1542) & (g1543) & (g1554) & (g1568)) + ((g229) & (g255) & (!g1542) & (!g1543) & (!g1554) & (!g1568)) + ((g229) & (g255) & (g1542) & (!g1543) & (!g1554) & (g1568)) + ((g229) & (g255) & (g1542) & (!g1543) & (g1554) & (!g1568)) + ((g229) & (g255) & (g1542) & (!g1543) & (g1554) & (g1568)) + ((g229) & (g255) & (g1542) & (g1543) & (!g1554) & (!g1568)) + ((g229) & (g255) & (g1542) & (g1543) & (!g1554) & (g1568)) + ((g229) & (g255) & (g1542) & (g1543) & (g1554) & (!g1568)) + ((g229) & (g255) & (g1542) & (g1543) & (g1554) & (g1568)));
	assign g1615 = (((!g255) & (!g1543) & (g1554) & (!g1568)) + ((!g255) & (g1543) & (!g1554) & (!g1568)) + ((!g255) & (g1543) & (!g1554) & (g1568)) + ((!g255) & (g1543) & (g1554) & (g1568)) + ((g255) & (!g1543) & (!g1554) & (!g1568)) + ((g255) & (g1543) & (!g1554) & (g1568)) + ((g255) & (g1543) & (g1554) & (!g1568)) + ((g255) & (g1543) & (g1554) & (g1568)));
	assign g1616 = (((!g290) & (!g319) & (!g1545) & (g1546) & (g1553) & (!g1568)) + ((!g290) & (!g319) & (g1545) & (!g1546) & (!g1553) & (!g1568)) + ((!g290) & (!g319) & (g1545) & (!g1546) & (!g1553) & (g1568)) + ((!g290) & (!g319) & (g1545) & (!g1546) & (g1553) & (!g1568)) + ((!g290) & (!g319) & (g1545) & (!g1546) & (g1553) & (g1568)) + ((!g290) & (!g319) & (g1545) & (g1546) & (!g1553) & (!g1568)) + ((!g290) & (!g319) & (g1545) & (g1546) & (!g1553) & (g1568)) + ((!g290) & (!g319) & (g1545) & (g1546) & (g1553) & (g1568)) + ((!g290) & (g319) & (!g1545) & (!g1546) & (g1553) & (!g1568)) + ((!g290) & (g319) & (!g1545) & (g1546) & (!g1553) & (!g1568)) + ((!g290) & (g319) & (!g1545) & (g1546) & (g1553) & (!g1568)) + ((!g290) & (g319) & (g1545) & (!g1546) & (!g1553) & (!g1568)) + ((!g290) & (g319) & (g1545) & (!g1546) & (!g1553) & (g1568)) + ((!g290) & (g319) & (g1545) & (!g1546) & (g1553) & (g1568)) + ((!g290) & (g319) & (g1545) & (g1546) & (!g1553) & (g1568)) + ((!g290) & (g319) & (g1545) & (g1546) & (g1553) & (g1568)) + ((g290) & (!g319) & (!g1545) & (!g1546) & (!g1553) & (!g1568)) + ((g290) & (!g319) & (!g1545) & (!g1546) & (g1553) & (!g1568)) + ((g290) & (!g319) & (!g1545) & (g1546) & (!g1553) & (!g1568)) + ((g290) & (!g319) & (g1545) & (!g1546) & (!g1553) & (g1568)) + ((g290) & (!g319) & (g1545) & (!g1546) & (g1553) & (g1568)) + ((g290) & (!g319) & (g1545) & (g1546) & (!g1553) & (g1568)) + ((g290) & (!g319) & (g1545) & (g1546) & (g1553) & (!g1568)) + ((g290) & (!g319) & (g1545) & (g1546) & (g1553) & (g1568)) + ((g290) & (g319) & (!g1545) & (!g1546) & (!g1553) & (!g1568)) + ((g290) & (g319) & (g1545) & (!g1546) & (!g1553) & (g1568)) + ((g290) & (g319) & (g1545) & (!g1546) & (g1553) & (!g1568)) + ((g290) & (g319) & (g1545) & (!g1546) & (g1553) & (g1568)) + ((g290) & (g319) & (g1545) & (g1546) & (!g1553) & (!g1568)) + ((g290) & (g319) & (g1545) & (g1546) & (!g1553) & (g1568)) + ((g290) & (g319) & (g1545) & (g1546) & (g1553) & (!g1568)) + ((g290) & (g319) & (g1545) & (g1546) & (g1553) & (g1568)));
	assign g1617 = (((!g319) & (!g1546) & (g1553) & (!g1568)) + ((!g319) & (g1546) & (!g1553) & (!g1568)) + ((!g319) & (g1546) & (!g1553) & (g1568)) + ((!g319) & (g1546) & (g1553) & (g1568)) + ((g319) & (!g1546) & (!g1553) & (!g1568)) + ((g319) & (g1546) & (!g1553) & (g1568)) + ((g319) & (g1546) & (g1553) & (!g1568)) + ((g319) & (g1546) & (g1553) & (g1568)));
	assign g1618 = (((!g358) & (!g390) & (!g1548) & (g1549) & (g1552) & (!g1568)) + ((!g358) & (!g390) & (g1548) & (!g1549) & (!g1552) & (!g1568)) + ((!g358) & (!g390) & (g1548) & (!g1549) & (!g1552) & (g1568)) + ((!g358) & (!g390) & (g1548) & (!g1549) & (g1552) & (!g1568)) + ((!g358) & (!g390) & (g1548) & (!g1549) & (g1552) & (g1568)) + ((!g358) & (!g390) & (g1548) & (g1549) & (!g1552) & (!g1568)) + ((!g358) & (!g390) & (g1548) & (g1549) & (!g1552) & (g1568)) + ((!g358) & (!g390) & (g1548) & (g1549) & (g1552) & (g1568)) + ((!g358) & (g390) & (!g1548) & (!g1549) & (g1552) & (!g1568)) + ((!g358) & (g390) & (!g1548) & (g1549) & (!g1552) & (!g1568)) + ((!g358) & (g390) & (!g1548) & (g1549) & (g1552) & (!g1568)) + ((!g358) & (g390) & (g1548) & (!g1549) & (!g1552) & (!g1568)) + ((!g358) & (g390) & (g1548) & (!g1549) & (!g1552) & (g1568)) + ((!g358) & (g390) & (g1548) & (!g1549) & (g1552) & (g1568)) + ((!g358) & (g390) & (g1548) & (g1549) & (!g1552) & (g1568)) + ((!g358) & (g390) & (g1548) & (g1549) & (g1552) & (g1568)) + ((g358) & (!g390) & (!g1548) & (!g1549) & (!g1552) & (!g1568)) + ((g358) & (!g390) & (!g1548) & (!g1549) & (g1552) & (!g1568)) + ((g358) & (!g390) & (!g1548) & (g1549) & (!g1552) & (!g1568)) + ((g358) & (!g390) & (g1548) & (!g1549) & (!g1552) & (g1568)) + ((g358) & (!g390) & (g1548) & (!g1549) & (g1552) & (g1568)) + ((g358) & (!g390) & (g1548) & (g1549) & (!g1552) & (g1568)) + ((g358) & (!g390) & (g1548) & (g1549) & (g1552) & (!g1568)) + ((g358) & (!g390) & (g1548) & (g1549) & (g1552) & (g1568)) + ((g358) & (g390) & (!g1548) & (!g1549) & (!g1552) & (!g1568)) + ((g358) & (g390) & (g1548) & (!g1549) & (!g1552) & (g1568)) + ((g358) & (g390) & (g1548) & (!g1549) & (g1552) & (!g1568)) + ((g358) & (g390) & (g1548) & (!g1549) & (g1552) & (g1568)) + ((g358) & (g390) & (g1548) & (g1549) & (!g1552) & (!g1568)) + ((g358) & (g390) & (g1548) & (g1549) & (!g1552) & (g1568)) + ((g358) & (g390) & (g1548) & (g1549) & (g1552) & (!g1568)) + ((g358) & (g390) & (g1548) & (g1549) & (g1552) & (g1568)));
	assign g1619 = (((!g390) & (!g1549) & (g1552) & (!g1568)) + ((!g390) & (g1549) & (!g1552) & (!g1568)) + ((!g390) & (g1549) & (!g1552) & (g1568)) + ((!g390) & (g1549) & (g1552) & (g1568)) + ((g390) & (!g1549) & (!g1552) & (!g1568)) + ((g390) & (g1549) & (!g1552) & (g1568)) + ((g390) & (g1549) & (g1552) & (!g1568)) + ((g390) & (g1549) & (g1552) & (g1568)));
	assign g1620 = (((!g433) & (!g468) & (!g1551) & (g1486) & (g1520) & (!g1568)) + ((!g433) & (!g468) & (g1551) & (!g1486) & (!g1520) & (!g1568)) + ((!g433) & (!g468) & (g1551) & (!g1486) & (!g1520) & (g1568)) + ((!g433) & (!g468) & (g1551) & (!g1486) & (g1520) & (!g1568)) + ((!g433) & (!g468) & (g1551) & (!g1486) & (g1520) & (g1568)) + ((!g433) & (!g468) & (g1551) & (g1486) & (!g1520) & (!g1568)) + ((!g433) & (!g468) & (g1551) & (g1486) & (!g1520) & (g1568)) + ((!g433) & (!g468) & (g1551) & (g1486) & (g1520) & (g1568)) + ((!g433) & (g468) & (!g1551) & (!g1486) & (g1520) & (!g1568)) + ((!g433) & (g468) & (!g1551) & (g1486) & (!g1520) & (!g1568)) + ((!g433) & (g468) & (!g1551) & (g1486) & (g1520) & (!g1568)) + ((!g433) & (g468) & (g1551) & (!g1486) & (!g1520) & (!g1568)) + ((!g433) & (g468) & (g1551) & (!g1486) & (!g1520) & (g1568)) + ((!g433) & (g468) & (g1551) & (!g1486) & (g1520) & (g1568)) + ((!g433) & (g468) & (g1551) & (g1486) & (!g1520) & (g1568)) + ((!g433) & (g468) & (g1551) & (g1486) & (g1520) & (g1568)) + ((g433) & (!g468) & (!g1551) & (!g1486) & (!g1520) & (!g1568)) + ((g433) & (!g468) & (!g1551) & (!g1486) & (g1520) & (!g1568)) + ((g433) & (!g468) & (!g1551) & (g1486) & (!g1520) & (!g1568)) + ((g433) & (!g468) & (g1551) & (!g1486) & (!g1520) & (g1568)) + ((g433) & (!g468) & (g1551) & (!g1486) & (g1520) & (g1568)) + ((g433) & (!g468) & (g1551) & (g1486) & (!g1520) & (g1568)) + ((g433) & (!g468) & (g1551) & (g1486) & (g1520) & (!g1568)) + ((g433) & (!g468) & (g1551) & (g1486) & (g1520) & (g1568)) + ((g433) & (g468) & (!g1551) & (!g1486) & (!g1520) & (!g1568)) + ((g433) & (g468) & (g1551) & (!g1486) & (!g1520) & (g1568)) + ((g433) & (g468) & (g1551) & (!g1486) & (g1520) & (!g1568)) + ((g433) & (g468) & (g1551) & (!g1486) & (g1520) & (g1568)) + ((g433) & (g468) & (g1551) & (g1486) & (!g1520) & (!g1568)) + ((g433) & (g468) & (g1551) & (g1486) & (!g1520) & (g1568)) + ((g433) & (g468) & (g1551) & (g1486) & (g1520) & (!g1568)) + ((g433) & (g468) & (g1551) & (g1486) & (g1520) & (g1568)));
	assign g1621 = (((!g390) & (!g433) & (g1620) & (g1569) & (g1599)) + ((!g390) & (g433) & (g1620) & (!g1569) & (g1599)) + ((!g390) & (g433) & (g1620) & (g1569) & (!g1599)) + ((!g390) & (g433) & (g1620) & (g1569) & (g1599)) + ((g390) & (!g433) & (!g1620) & (g1569) & (g1599)) + ((g390) & (!g433) & (g1620) & (!g1569) & (!g1599)) + ((g390) & (!g433) & (g1620) & (!g1569) & (g1599)) + ((g390) & (!g433) & (g1620) & (g1569) & (!g1599)) + ((g390) & (!g433) & (g1620) & (g1569) & (g1599)) + ((g390) & (g433) & (!g1620) & (!g1569) & (g1599)) + ((g390) & (g433) & (!g1620) & (g1569) & (!g1599)) + ((g390) & (g433) & (!g1620) & (g1569) & (g1599)) + ((g390) & (g433) & (g1620) & (!g1569) & (!g1599)) + ((g390) & (g433) & (g1620) & (!g1569) & (g1599)) + ((g390) & (g433) & (g1620) & (g1569) & (!g1599)) + ((g390) & (g433) & (g1620) & (g1569) & (g1599)));
	assign g1622 = (((!g319) & (!g358) & (g1618) & (g1619) & (g1621)) + ((!g319) & (g358) & (g1618) & (!g1619) & (g1621)) + ((!g319) & (g358) & (g1618) & (g1619) & (!g1621)) + ((!g319) & (g358) & (g1618) & (g1619) & (g1621)) + ((g319) & (!g358) & (!g1618) & (g1619) & (g1621)) + ((g319) & (!g358) & (g1618) & (!g1619) & (!g1621)) + ((g319) & (!g358) & (g1618) & (!g1619) & (g1621)) + ((g319) & (!g358) & (g1618) & (g1619) & (!g1621)) + ((g319) & (!g358) & (g1618) & (g1619) & (g1621)) + ((g319) & (g358) & (!g1618) & (!g1619) & (g1621)) + ((g319) & (g358) & (!g1618) & (g1619) & (!g1621)) + ((g319) & (g358) & (!g1618) & (g1619) & (g1621)) + ((g319) & (g358) & (g1618) & (!g1619) & (!g1621)) + ((g319) & (g358) & (g1618) & (!g1619) & (g1621)) + ((g319) & (g358) & (g1618) & (g1619) & (!g1621)) + ((g319) & (g358) & (g1618) & (g1619) & (g1621)));
	assign g1623 = (((!g255) & (!g290) & (g1616) & (g1617) & (g1622)) + ((!g255) & (g290) & (g1616) & (!g1617) & (g1622)) + ((!g255) & (g290) & (g1616) & (g1617) & (!g1622)) + ((!g255) & (g290) & (g1616) & (g1617) & (g1622)) + ((g255) & (!g290) & (!g1616) & (g1617) & (g1622)) + ((g255) & (!g290) & (g1616) & (!g1617) & (!g1622)) + ((g255) & (!g290) & (g1616) & (!g1617) & (g1622)) + ((g255) & (!g290) & (g1616) & (g1617) & (!g1622)) + ((g255) & (!g290) & (g1616) & (g1617) & (g1622)) + ((g255) & (g290) & (!g1616) & (!g1617) & (g1622)) + ((g255) & (g290) & (!g1616) & (g1617) & (!g1622)) + ((g255) & (g290) & (!g1616) & (g1617) & (g1622)) + ((g255) & (g290) & (g1616) & (!g1617) & (!g1622)) + ((g255) & (g290) & (g1616) & (!g1617) & (g1622)) + ((g255) & (g290) & (g1616) & (g1617) & (!g1622)) + ((g255) & (g290) & (g1616) & (g1617) & (g1622)));
	assign g1624 = (((!g198) & (!g229) & (g1614) & (g1615) & (g1623)) + ((!g198) & (g229) & (g1614) & (!g1615) & (g1623)) + ((!g198) & (g229) & (g1614) & (g1615) & (!g1623)) + ((!g198) & (g229) & (g1614) & (g1615) & (g1623)) + ((g198) & (!g229) & (!g1614) & (g1615) & (g1623)) + ((g198) & (!g229) & (g1614) & (!g1615) & (!g1623)) + ((g198) & (!g229) & (g1614) & (!g1615) & (g1623)) + ((g198) & (!g229) & (g1614) & (g1615) & (!g1623)) + ((g198) & (!g229) & (g1614) & (g1615) & (g1623)) + ((g198) & (g229) & (!g1614) & (!g1615) & (g1623)) + ((g198) & (g229) & (!g1614) & (g1615) & (!g1623)) + ((g198) & (g229) & (!g1614) & (g1615) & (g1623)) + ((g198) & (g229) & (g1614) & (!g1615) & (!g1623)) + ((g198) & (g229) & (g1614) & (!g1615) & (g1623)) + ((g198) & (g229) & (g1614) & (g1615) & (!g1623)) + ((g198) & (g229) & (g1614) & (g1615) & (g1623)));
	assign g1625 = (((!g147) & (!g174) & (g1612) & (g1613) & (g1624)) + ((!g147) & (g174) & (g1612) & (!g1613) & (g1624)) + ((!g147) & (g174) & (g1612) & (g1613) & (!g1624)) + ((!g147) & (g174) & (g1612) & (g1613) & (g1624)) + ((g147) & (!g174) & (!g1612) & (g1613) & (g1624)) + ((g147) & (!g174) & (g1612) & (!g1613) & (!g1624)) + ((g147) & (!g174) & (g1612) & (!g1613) & (g1624)) + ((g147) & (!g174) & (g1612) & (g1613) & (!g1624)) + ((g147) & (!g174) & (g1612) & (g1613) & (g1624)) + ((g147) & (g174) & (!g1612) & (!g1613) & (g1624)) + ((g147) & (g174) & (!g1612) & (g1613) & (!g1624)) + ((g147) & (g174) & (!g1612) & (g1613) & (g1624)) + ((g147) & (g174) & (g1612) & (!g1613) & (!g1624)) + ((g147) & (g174) & (g1612) & (!g1613) & (g1624)) + ((g147) & (g174) & (g1612) & (g1613) & (!g1624)) + ((g147) & (g174) & (g1612) & (g1613) & (g1624)));
	assign g1626 = (((!g104) & (!g127) & (g1610) & (g1611) & (g1625)) + ((!g104) & (g127) & (g1610) & (!g1611) & (g1625)) + ((!g104) & (g127) & (g1610) & (g1611) & (!g1625)) + ((!g104) & (g127) & (g1610) & (g1611) & (g1625)) + ((g104) & (!g127) & (!g1610) & (g1611) & (g1625)) + ((g104) & (!g127) & (g1610) & (!g1611) & (!g1625)) + ((g104) & (!g127) & (g1610) & (!g1611) & (g1625)) + ((g104) & (!g127) & (g1610) & (g1611) & (!g1625)) + ((g104) & (!g127) & (g1610) & (g1611) & (g1625)) + ((g104) & (g127) & (!g1610) & (!g1611) & (g1625)) + ((g104) & (g127) & (!g1610) & (g1611) & (!g1625)) + ((g104) & (g127) & (!g1610) & (g1611) & (g1625)) + ((g104) & (g127) & (g1610) & (!g1611) & (!g1625)) + ((g104) & (g127) & (g1610) & (!g1611) & (g1625)) + ((g104) & (g127) & (g1610) & (g1611) & (!g1625)) + ((g104) & (g127) & (g1610) & (g1611) & (g1625)));
	assign g1627 = (((!g68) & (!g87) & (g1608) & (g1609) & (g1626)) + ((!g68) & (g87) & (g1608) & (!g1609) & (g1626)) + ((!g68) & (g87) & (g1608) & (g1609) & (!g1626)) + ((!g68) & (g87) & (g1608) & (g1609) & (g1626)) + ((g68) & (!g87) & (!g1608) & (g1609) & (g1626)) + ((g68) & (!g87) & (g1608) & (!g1609) & (!g1626)) + ((g68) & (!g87) & (g1608) & (!g1609) & (g1626)) + ((g68) & (!g87) & (g1608) & (g1609) & (!g1626)) + ((g68) & (!g87) & (g1608) & (g1609) & (g1626)) + ((g68) & (g87) & (!g1608) & (!g1609) & (g1626)) + ((g68) & (g87) & (!g1608) & (g1609) & (!g1626)) + ((g68) & (g87) & (!g1608) & (g1609) & (g1626)) + ((g68) & (g87) & (g1608) & (!g1609) & (!g1626)) + ((g68) & (g87) & (g1608) & (!g1609) & (g1626)) + ((g68) & (g87) & (g1608) & (g1609) & (!g1626)) + ((g68) & (g87) & (g1608) & (g1609) & (g1626)));
	assign g1628 = (((!g39) & (!g54) & (g1606) & (g1607) & (g1627)) + ((!g39) & (g54) & (g1606) & (!g1607) & (g1627)) + ((!g39) & (g54) & (g1606) & (g1607) & (!g1627)) + ((!g39) & (g54) & (g1606) & (g1607) & (g1627)) + ((g39) & (!g54) & (!g1606) & (g1607) & (g1627)) + ((g39) & (!g54) & (g1606) & (!g1607) & (!g1627)) + ((g39) & (!g54) & (g1606) & (!g1607) & (g1627)) + ((g39) & (!g54) & (g1606) & (g1607) & (!g1627)) + ((g39) & (!g54) & (g1606) & (g1607) & (g1627)) + ((g39) & (g54) & (!g1606) & (!g1607) & (g1627)) + ((g39) & (g54) & (!g1606) & (g1607) & (!g1627)) + ((g39) & (g54) & (!g1606) & (g1607) & (g1627)) + ((g39) & (g54) & (g1606) & (!g1607) & (!g1627)) + ((g39) & (g54) & (g1606) & (!g1607) & (g1627)) + ((g39) & (g54) & (g1606) & (g1607) & (!g1627)) + ((g39) & (g54) & (g1606) & (g1607) & (g1627)));
	assign g1629 = (((!g18) & (!g27) & (g1604) & (g1605) & (g1628)) + ((!g18) & (g27) & (g1604) & (!g1605) & (g1628)) + ((!g18) & (g27) & (g1604) & (g1605) & (!g1628)) + ((!g18) & (g27) & (g1604) & (g1605) & (g1628)) + ((g18) & (!g27) & (!g1604) & (g1605) & (g1628)) + ((g18) & (!g27) & (g1604) & (!g1605) & (!g1628)) + ((g18) & (!g27) & (g1604) & (!g1605) & (g1628)) + ((g18) & (!g27) & (g1604) & (g1605) & (!g1628)) + ((g18) & (!g27) & (g1604) & (g1605) & (g1628)) + ((g18) & (g27) & (!g1604) & (!g1605) & (g1628)) + ((g18) & (g27) & (!g1604) & (g1605) & (!g1628)) + ((g18) & (g27) & (!g1604) & (g1605) & (g1628)) + ((g18) & (g27) & (g1604) & (!g1605) & (!g1628)) + ((g18) & (g27) & (g1604) & (!g1605) & (g1628)) + ((g18) & (g27) & (g1604) & (g1605) & (!g1628)) + ((g18) & (g27) & (g1604) & (g1605) & (g1628)));
	assign g1630 = (((!g2) & (!g8) & (g1602) & (g1603) & (g1629)) + ((!g2) & (g8) & (g1602) & (!g1603) & (g1629)) + ((!g2) & (g8) & (g1602) & (g1603) & (!g1629)) + ((!g2) & (g8) & (g1602) & (g1603) & (g1629)) + ((g2) & (!g8) & (!g1602) & (g1603) & (g1629)) + ((g2) & (!g8) & (g1602) & (!g1603) & (!g1629)) + ((g2) & (!g8) & (g1602) & (!g1603) & (g1629)) + ((g2) & (!g8) & (g1602) & (g1603) & (!g1629)) + ((g2) & (!g8) & (g1602) & (g1603) & (g1629)) + ((g2) & (g8) & (!g1602) & (!g1603) & (g1629)) + ((g2) & (g8) & (!g1602) & (g1603) & (!g1629)) + ((g2) & (g8) & (!g1602) & (g1603) & (g1629)) + ((g2) & (g8) & (g1602) & (!g1603) & (!g1629)) + ((g2) & (g8) & (g1602) & (!g1603) & (g1629)) + ((g2) & (g8) & (g1602) & (g1603) & (!g1629)) + ((g2) & (g8) & (g1602) & (g1603) & (g1629)));
	assign g1631 = (((!g2) & (!g1522) & (g1561) & (!g1568)) + ((!g2) & (g1522) & (!g1561) & (!g1568)) + ((!g2) & (g1522) & (!g1561) & (g1568)) + ((!g2) & (g1522) & (g1561) & (g1568)) + ((g2) & (!g1522) & (!g1561) & (!g1568)) + ((g2) & (g1522) & (!g1561) & (g1568)) + ((g2) & (g1522) & (g1561) & (!g1568)) + ((g2) & (g1522) & (g1561) & (g1568)));
	assign g1632 = (((!g1) & (!g1521) & (!g1564) & (!g1566) & (g1567)) + ((!g1) & (!g1521) & (!g1564) & (g1566) & (!g1567)) + ((!g1) & (!g1521) & (!g1564) & (g1566) & (g1567)) + ((!g1) & (g1521) & (g1564) & (!g1566) & (!g1567)) + ((!g1) & (g1521) & (g1564) & (!g1566) & (g1567)) + ((!g1) & (g1521) & (g1564) & (g1566) & (!g1567)) + ((!g1) & (g1521) & (g1564) & (g1566) & (g1567)) + ((g1) & (!g1521) & (!g1564) & (!g1566) & (g1567)) + ((g1) & (!g1521) & (!g1564) & (g1566) & (g1567)) + ((g1) & (g1521) & (g1564) & (!g1566) & (!g1567)) + ((g1) & (g1521) & (g1564) & (!g1566) & (g1567)) + ((g1) & (g1521) & (g1564) & (g1566) & (!g1567)) + ((g1) & (g1521) & (g1564) & (g1566) & (g1567)));
	assign g1633 = (((!g4) & (!g1) & (!g1601) & (!g1630) & (!g1631) & (!g1632)) + ((!g4) & (g1) & (!g1601) & (!g1630) & (!g1631) & (!g1632)) + ((!g4) & (g1) & (!g1601) & (!g1630) & (!g1631) & (g1632)) + ((!g4) & (g1) & (!g1601) & (!g1630) & (g1631) & (!g1632)) + ((!g4) & (g1) & (!g1601) & (!g1630) & (g1631) & (g1632)) + ((!g4) & (g1) & (!g1601) & (g1630) & (!g1631) & (!g1632)) + ((!g4) & (g1) & (!g1601) & (g1630) & (!g1631) & (g1632)) + ((!g4) & (g1) & (!g1601) & (g1630) & (g1631) & (!g1632)) + ((!g4) & (g1) & (!g1601) & (g1630) & (g1631) & (g1632)) + ((!g4) & (g1) & (g1601) & (!g1630) & (!g1631) & (!g1632)) + ((!g4) & (g1) & (g1601) & (!g1630) & (!g1631) & (g1632)) + ((g4) & (!g1) & (!g1601) & (!g1630) & (!g1631) & (!g1632)) + ((g4) & (!g1) & (!g1601) & (!g1630) & (g1631) & (!g1632)) + ((g4) & (!g1) & (!g1601) & (g1630) & (!g1631) & (!g1632)) + ((g4) & (g1) & (!g1601) & (!g1630) & (!g1631) & (!g1632)) + ((g4) & (g1) & (!g1601) & (!g1630) & (!g1631) & (g1632)) + ((g4) & (g1) & (!g1601) & (!g1630) & (g1631) & (!g1632)) + ((g4) & (g1) & (!g1601) & (!g1630) & (g1631) & (g1632)) + ((g4) & (g1) & (!g1601) & (g1630) & (!g1631) & (!g1632)) + ((g4) & (g1) & (!g1601) & (g1630) & (!g1631) & (g1632)) + ((g4) & (g1) & (!g1601) & (g1630) & (g1631) & (!g1632)) + ((g4) & (g1) & (!g1601) & (g1630) & (g1631) & (g1632)) + ((g4) & (g1) & (g1601) & (!g1630) & (!g1631) & (!g1632)) + ((g4) & (g1) & (g1601) & (!g1630) & (!g1631) & (g1632)) + ((g4) & (g1) & (g1601) & (!g1630) & (g1631) & (!g1632)) + ((g4) & (g1) & (g1601) & (!g1630) & (g1631) & (g1632)) + ((g4) & (g1) & (g1601) & (g1630) & (!g1631) & (!g1632)) + ((g4) & (g1) & (g1601) & (g1630) & (!g1631) & (g1632)));
	assign g1634 = (((!g433) & (!g1569) & (g1599) & (!g1600) & (!g1633)) + ((!g433) & (!g1569) & (g1599) & (g1600) & (!g1633)) + ((!g433) & (!g1569) & (g1599) & (g1600) & (g1633)) + ((!g433) & (g1569) & (!g1599) & (!g1600) & (!g1633)) + ((!g433) & (g1569) & (!g1599) & (!g1600) & (g1633)) + ((!g433) & (g1569) & (!g1599) & (g1600) & (!g1633)) + ((!g433) & (g1569) & (!g1599) & (g1600) & (g1633)) + ((!g433) & (g1569) & (g1599) & (!g1600) & (g1633)) + ((g433) & (!g1569) & (!g1599) & (!g1600) & (!g1633)) + ((g433) & (!g1569) & (!g1599) & (g1600) & (!g1633)) + ((g433) & (!g1569) & (!g1599) & (g1600) & (g1633)) + ((g433) & (g1569) & (!g1599) & (!g1600) & (g1633)) + ((g433) & (g1569) & (g1599) & (!g1600) & (!g1633)) + ((g433) & (g1569) & (g1599) & (!g1600) & (g1633)) + ((g433) & (g1569) & (g1599) & (g1600) & (!g1633)) + ((g433) & (g1569) & (g1599) & (g1600) & (g1633)));
	assign g1635 = (((!g468) & (!g515) & (g1571) & (g1598)) + ((!g468) & (g515) & (!g1571) & (g1598)) + ((!g468) & (g515) & (g1571) & (!g1598)) + ((!g468) & (g515) & (g1571) & (g1598)) + ((g468) & (!g515) & (!g1571) & (!g1598)) + ((g468) & (!g515) & (!g1571) & (g1598)) + ((g468) & (!g515) & (g1571) & (!g1598)) + ((g468) & (g515) & (!g1571) & (!g1598)));
	assign g1636 = (((!g1570) & (!g1600) & (!g1633) & (g1635)) + ((!g1570) & (g1600) & (!g1633) & (g1635)) + ((!g1570) & (g1600) & (g1633) & (g1635)) + ((g1570) & (!g1600) & (!g1633) & (!g1635)) + ((g1570) & (!g1600) & (g1633) & (!g1635)) + ((g1570) & (!g1600) & (g1633) & (g1635)) + ((g1570) & (g1600) & (!g1633) & (!g1635)) + ((g1570) & (g1600) & (g1633) & (!g1635)));
	assign g1637 = (((!g515) & (!g1571) & (g1598) & (!g1600) & (!g1633)) + ((!g515) & (!g1571) & (g1598) & (g1600) & (!g1633)) + ((!g515) & (!g1571) & (g1598) & (g1600) & (g1633)) + ((!g515) & (g1571) & (!g1598) & (!g1600) & (!g1633)) + ((!g515) & (g1571) & (!g1598) & (!g1600) & (g1633)) + ((!g515) & (g1571) & (!g1598) & (g1600) & (!g1633)) + ((!g515) & (g1571) & (!g1598) & (g1600) & (g1633)) + ((!g515) & (g1571) & (g1598) & (!g1600) & (g1633)) + ((g515) & (!g1571) & (!g1598) & (!g1600) & (!g1633)) + ((g515) & (!g1571) & (!g1598) & (g1600) & (!g1633)) + ((g515) & (!g1571) & (!g1598) & (g1600) & (g1633)) + ((g515) & (g1571) & (!g1598) & (!g1600) & (g1633)) + ((g515) & (g1571) & (g1598) & (!g1600) & (!g1633)) + ((g515) & (g1571) & (g1598) & (!g1600) & (g1633)) + ((g515) & (g1571) & (g1598) & (g1600) & (!g1633)) + ((g515) & (g1571) & (g1598) & (g1600) & (g1633)));
	assign g1638 = (((!g553) & (!g604) & (g1573) & (g1597)) + ((!g553) & (g604) & (!g1573) & (g1597)) + ((!g553) & (g604) & (g1573) & (!g1597)) + ((!g553) & (g604) & (g1573) & (g1597)) + ((g553) & (!g604) & (!g1573) & (!g1597)) + ((g553) & (!g604) & (!g1573) & (g1597)) + ((g553) & (!g604) & (g1573) & (!g1597)) + ((g553) & (g604) & (!g1573) & (!g1597)));
	assign g1639 = (((!g1572) & (!g1600) & (!g1633) & (g1638)) + ((!g1572) & (g1600) & (!g1633) & (g1638)) + ((!g1572) & (g1600) & (g1633) & (g1638)) + ((g1572) & (!g1600) & (!g1633) & (!g1638)) + ((g1572) & (!g1600) & (g1633) & (!g1638)) + ((g1572) & (!g1600) & (g1633) & (g1638)) + ((g1572) & (g1600) & (!g1633) & (!g1638)) + ((g1572) & (g1600) & (g1633) & (!g1638)));
	assign g1640 = (((!g604) & (!g1573) & (g1597) & (!g1600) & (!g1633)) + ((!g604) & (!g1573) & (g1597) & (g1600) & (!g1633)) + ((!g604) & (!g1573) & (g1597) & (g1600) & (g1633)) + ((!g604) & (g1573) & (!g1597) & (!g1600) & (!g1633)) + ((!g604) & (g1573) & (!g1597) & (!g1600) & (g1633)) + ((!g604) & (g1573) & (!g1597) & (g1600) & (!g1633)) + ((!g604) & (g1573) & (!g1597) & (g1600) & (g1633)) + ((!g604) & (g1573) & (g1597) & (!g1600) & (g1633)) + ((g604) & (!g1573) & (!g1597) & (!g1600) & (!g1633)) + ((g604) & (!g1573) & (!g1597) & (g1600) & (!g1633)) + ((g604) & (!g1573) & (!g1597) & (g1600) & (g1633)) + ((g604) & (g1573) & (!g1597) & (!g1600) & (g1633)) + ((g604) & (g1573) & (g1597) & (!g1600) & (!g1633)) + ((g604) & (g1573) & (g1597) & (!g1600) & (g1633)) + ((g604) & (g1573) & (g1597) & (g1600) & (!g1633)) + ((g604) & (g1573) & (g1597) & (g1600) & (g1633)));
	assign g1641 = (((!g645) & (!g700) & (g1575) & (g1596)) + ((!g645) & (g700) & (!g1575) & (g1596)) + ((!g645) & (g700) & (g1575) & (!g1596)) + ((!g645) & (g700) & (g1575) & (g1596)) + ((g645) & (!g700) & (!g1575) & (!g1596)) + ((g645) & (!g700) & (!g1575) & (g1596)) + ((g645) & (!g700) & (g1575) & (!g1596)) + ((g645) & (g700) & (!g1575) & (!g1596)));
	assign g1642 = (((!g1574) & (!g1600) & (!g1633) & (g1641)) + ((!g1574) & (g1600) & (!g1633) & (g1641)) + ((!g1574) & (g1600) & (g1633) & (g1641)) + ((g1574) & (!g1600) & (!g1633) & (!g1641)) + ((g1574) & (!g1600) & (g1633) & (!g1641)) + ((g1574) & (!g1600) & (g1633) & (g1641)) + ((g1574) & (g1600) & (!g1633) & (!g1641)) + ((g1574) & (g1600) & (g1633) & (!g1641)));
	assign g1643 = (((!g700) & (!g1575) & (g1596) & (!g1600) & (!g1633)) + ((!g700) & (!g1575) & (g1596) & (g1600) & (!g1633)) + ((!g700) & (!g1575) & (g1596) & (g1600) & (g1633)) + ((!g700) & (g1575) & (!g1596) & (!g1600) & (!g1633)) + ((!g700) & (g1575) & (!g1596) & (!g1600) & (g1633)) + ((!g700) & (g1575) & (!g1596) & (g1600) & (!g1633)) + ((!g700) & (g1575) & (!g1596) & (g1600) & (g1633)) + ((!g700) & (g1575) & (g1596) & (!g1600) & (g1633)) + ((g700) & (!g1575) & (!g1596) & (!g1600) & (!g1633)) + ((g700) & (!g1575) & (!g1596) & (g1600) & (!g1633)) + ((g700) & (!g1575) & (!g1596) & (g1600) & (g1633)) + ((g700) & (g1575) & (!g1596) & (!g1600) & (g1633)) + ((g700) & (g1575) & (g1596) & (!g1600) & (!g1633)) + ((g700) & (g1575) & (g1596) & (!g1600) & (g1633)) + ((g700) & (g1575) & (g1596) & (g1600) & (!g1633)) + ((g700) & (g1575) & (g1596) & (g1600) & (g1633)));
	assign g1644 = (((!g744) & (!g803) & (g1577) & (g1595)) + ((!g744) & (g803) & (!g1577) & (g1595)) + ((!g744) & (g803) & (g1577) & (!g1595)) + ((!g744) & (g803) & (g1577) & (g1595)) + ((g744) & (!g803) & (!g1577) & (!g1595)) + ((g744) & (!g803) & (!g1577) & (g1595)) + ((g744) & (!g803) & (g1577) & (!g1595)) + ((g744) & (g803) & (!g1577) & (!g1595)));
	assign g1645 = (((!g1576) & (!g1600) & (!g1633) & (g1644)) + ((!g1576) & (g1600) & (!g1633) & (g1644)) + ((!g1576) & (g1600) & (g1633) & (g1644)) + ((g1576) & (!g1600) & (!g1633) & (!g1644)) + ((g1576) & (!g1600) & (g1633) & (!g1644)) + ((g1576) & (!g1600) & (g1633) & (g1644)) + ((g1576) & (g1600) & (!g1633) & (!g1644)) + ((g1576) & (g1600) & (g1633) & (!g1644)));
	assign g1646 = (((!g803) & (!g1577) & (g1595) & (!g1600) & (!g1633)) + ((!g803) & (!g1577) & (g1595) & (g1600) & (!g1633)) + ((!g803) & (!g1577) & (g1595) & (g1600) & (g1633)) + ((!g803) & (g1577) & (!g1595) & (!g1600) & (!g1633)) + ((!g803) & (g1577) & (!g1595) & (!g1600) & (g1633)) + ((!g803) & (g1577) & (!g1595) & (g1600) & (!g1633)) + ((!g803) & (g1577) & (!g1595) & (g1600) & (g1633)) + ((!g803) & (g1577) & (g1595) & (!g1600) & (g1633)) + ((g803) & (!g1577) & (!g1595) & (!g1600) & (!g1633)) + ((g803) & (!g1577) & (!g1595) & (g1600) & (!g1633)) + ((g803) & (!g1577) & (!g1595) & (g1600) & (g1633)) + ((g803) & (g1577) & (!g1595) & (!g1600) & (g1633)) + ((g803) & (g1577) & (g1595) & (!g1600) & (!g1633)) + ((g803) & (g1577) & (g1595) & (!g1600) & (g1633)) + ((g803) & (g1577) & (g1595) & (g1600) & (!g1633)) + ((g803) & (g1577) & (g1595) & (g1600) & (g1633)));
	assign g1647 = (((!g851) & (!g914) & (g1579) & (g1594)) + ((!g851) & (g914) & (!g1579) & (g1594)) + ((!g851) & (g914) & (g1579) & (!g1594)) + ((!g851) & (g914) & (g1579) & (g1594)) + ((g851) & (!g914) & (!g1579) & (!g1594)) + ((g851) & (!g914) & (!g1579) & (g1594)) + ((g851) & (!g914) & (g1579) & (!g1594)) + ((g851) & (g914) & (!g1579) & (!g1594)));
	assign g1648 = (((!g1578) & (!g1600) & (!g1633) & (g1647)) + ((!g1578) & (g1600) & (!g1633) & (g1647)) + ((!g1578) & (g1600) & (g1633) & (g1647)) + ((g1578) & (!g1600) & (!g1633) & (!g1647)) + ((g1578) & (!g1600) & (g1633) & (!g1647)) + ((g1578) & (!g1600) & (g1633) & (g1647)) + ((g1578) & (g1600) & (!g1633) & (!g1647)) + ((g1578) & (g1600) & (g1633) & (!g1647)));
	assign g1649 = (((!g914) & (!g1579) & (g1594) & (!g1600) & (!g1633)) + ((!g914) & (!g1579) & (g1594) & (g1600) & (!g1633)) + ((!g914) & (!g1579) & (g1594) & (g1600) & (g1633)) + ((!g914) & (g1579) & (!g1594) & (!g1600) & (!g1633)) + ((!g914) & (g1579) & (!g1594) & (!g1600) & (g1633)) + ((!g914) & (g1579) & (!g1594) & (g1600) & (!g1633)) + ((!g914) & (g1579) & (!g1594) & (g1600) & (g1633)) + ((!g914) & (g1579) & (g1594) & (!g1600) & (g1633)) + ((g914) & (!g1579) & (!g1594) & (!g1600) & (!g1633)) + ((g914) & (!g1579) & (!g1594) & (g1600) & (!g1633)) + ((g914) & (!g1579) & (!g1594) & (g1600) & (g1633)) + ((g914) & (g1579) & (!g1594) & (!g1600) & (g1633)) + ((g914) & (g1579) & (g1594) & (!g1600) & (!g1633)) + ((g914) & (g1579) & (g1594) & (!g1600) & (g1633)) + ((g914) & (g1579) & (g1594) & (g1600) & (!g1633)) + ((g914) & (g1579) & (g1594) & (g1600) & (g1633)));
	assign g1650 = (((!g1032) & (!g1030) & (g1581) & (g1593)) + ((!g1032) & (g1030) & (!g1581) & (g1593)) + ((!g1032) & (g1030) & (g1581) & (!g1593)) + ((!g1032) & (g1030) & (g1581) & (g1593)) + ((g1032) & (!g1030) & (!g1581) & (!g1593)) + ((g1032) & (!g1030) & (!g1581) & (g1593)) + ((g1032) & (!g1030) & (g1581) & (!g1593)) + ((g1032) & (g1030) & (!g1581) & (!g1593)));
	assign g1651 = (((!g1580) & (!g1600) & (!g1633) & (g1650)) + ((!g1580) & (g1600) & (!g1633) & (g1650)) + ((!g1580) & (g1600) & (g1633) & (g1650)) + ((g1580) & (!g1600) & (!g1633) & (!g1650)) + ((g1580) & (!g1600) & (g1633) & (!g1650)) + ((g1580) & (!g1600) & (g1633) & (g1650)) + ((g1580) & (g1600) & (!g1633) & (!g1650)) + ((g1580) & (g1600) & (g1633) & (!g1650)));
	assign g1652 = (((!g1030) & (!g1581) & (g1593) & (!g1600) & (!g1633)) + ((!g1030) & (!g1581) & (g1593) & (g1600) & (!g1633)) + ((!g1030) & (!g1581) & (g1593) & (g1600) & (g1633)) + ((!g1030) & (g1581) & (!g1593) & (!g1600) & (!g1633)) + ((!g1030) & (g1581) & (!g1593) & (!g1600) & (g1633)) + ((!g1030) & (g1581) & (!g1593) & (g1600) & (!g1633)) + ((!g1030) & (g1581) & (!g1593) & (g1600) & (g1633)) + ((!g1030) & (g1581) & (g1593) & (!g1600) & (g1633)) + ((g1030) & (!g1581) & (!g1593) & (!g1600) & (!g1633)) + ((g1030) & (!g1581) & (!g1593) & (g1600) & (!g1633)) + ((g1030) & (!g1581) & (!g1593) & (g1600) & (g1633)) + ((g1030) & (g1581) & (!g1593) & (!g1600) & (g1633)) + ((g1030) & (g1581) & (g1593) & (!g1600) & (!g1633)) + ((g1030) & (g1581) & (g1593) & (!g1600) & (g1633)) + ((g1030) & (g1581) & (g1593) & (g1600) & (!g1633)) + ((g1030) & (g1581) & (g1593) & (g1600) & (g1633)));
	assign g1653 = (((!g1160) & (!g1154) & (g1583) & (g1592)) + ((!g1160) & (g1154) & (!g1583) & (g1592)) + ((!g1160) & (g1154) & (g1583) & (!g1592)) + ((!g1160) & (g1154) & (g1583) & (g1592)) + ((g1160) & (!g1154) & (!g1583) & (!g1592)) + ((g1160) & (!g1154) & (!g1583) & (g1592)) + ((g1160) & (!g1154) & (g1583) & (!g1592)) + ((g1160) & (g1154) & (!g1583) & (!g1592)));
	assign g1654 = (((!g1582) & (!g1600) & (!g1633) & (g1653)) + ((!g1582) & (g1600) & (!g1633) & (g1653)) + ((!g1582) & (g1600) & (g1633) & (g1653)) + ((g1582) & (!g1600) & (!g1633) & (!g1653)) + ((g1582) & (!g1600) & (g1633) & (!g1653)) + ((g1582) & (!g1600) & (g1633) & (g1653)) + ((g1582) & (g1600) & (!g1633) & (!g1653)) + ((g1582) & (g1600) & (g1633) & (!g1653)));
	assign g1655 = (((!g1154) & (!g1583) & (g1592) & (!g1600) & (!g1633)) + ((!g1154) & (!g1583) & (g1592) & (g1600) & (!g1633)) + ((!g1154) & (!g1583) & (g1592) & (g1600) & (g1633)) + ((!g1154) & (g1583) & (!g1592) & (!g1600) & (!g1633)) + ((!g1154) & (g1583) & (!g1592) & (!g1600) & (g1633)) + ((!g1154) & (g1583) & (!g1592) & (g1600) & (!g1633)) + ((!g1154) & (g1583) & (!g1592) & (g1600) & (g1633)) + ((!g1154) & (g1583) & (g1592) & (!g1600) & (g1633)) + ((g1154) & (!g1583) & (!g1592) & (!g1600) & (!g1633)) + ((g1154) & (!g1583) & (!g1592) & (g1600) & (!g1633)) + ((g1154) & (!g1583) & (!g1592) & (g1600) & (g1633)) + ((g1154) & (g1583) & (!g1592) & (!g1600) & (g1633)) + ((g1154) & (g1583) & (g1592) & (!g1600) & (!g1633)) + ((g1154) & (g1583) & (g1592) & (!g1600) & (g1633)) + ((g1154) & (g1583) & (g1592) & (g1600) & (!g1633)) + ((g1154) & (g1583) & (g1592) & (g1600) & (g1633)));
	assign g1656 = (((!g1295) & (!g1285) & (g1585) & (g1591)) + ((!g1295) & (g1285) & (!g1585) & (g1591)) + ((!g1295) & (g1285) & (g1585) & (!g1591)) + ((!g1295) & (g1285) & (g1585) & (g1591)) + ((g1295) & (!g1285) & (!g1585) & (!g1591)) + ((g1295) & (!g1285) & (!g1585) & (g1591)) + ((g1295) & (!g1285) & (g1585) & (!g1591)) + ((g1295) & (g1285) & (!g1585) & (!g1591)));
	assign g1657 = (((!g1584) & (!g1600) & (!g1633) & (g1656)) + ((!g1584) & (g1600) & (!g1633) & (g1656)) + ((!g1584) & (g1600) & (g1633) & (g1656)) + ((g1584) & (!g1600) & (!g1633) & (!g1656)) + ((g1584) & (!g1600) & (g1633) & (!g1656)) + ((g1584) & (!g1600) & (g1633) & (g1656)) + ((g1584) & (g1600) & (!g1633) & (!g1656)) + ((g1584) & (g1600) & (g1633) & (!g1656)));
	assign g1658 = (((!g1285) & (!g1585) & (g1591) & (!g1600) & (!g1633)) + ((!g1285) & (!g1585) & (g1591) & (g1600) & (!g1633)) + ((!g1285) & (!g1585) & (g1591) & (g1600) & (g1633)) + ((!g1285) & (g1585) & (!g1591) & (!g1600) & (!g1633)) + ((!g1285) & (g1585) & (!g1591) & (!g1600) & (g1633)) + ((!g1285) & (g1585) & (!g1591) & (g1600) & (!g1633)) + ((!g1285) & (g1585) & (!g1591) & (g1600) & (g1633)) + ((!g1285) & (g1585) & (g1591) & (!g1600) & (g1633)) + ((g1285) & (!g1585) & (!g1591) & (!g1600) & (!g1633)) + ((g1285) & (!g1585) & (!g1591) & (g1600) & (!g1633)) + ((g1285) & (!g1585) & (!g1591) & (g1600) & (g1633)) + ((g1285) & (g1585) & (!g1591) & (!g1600) & (g1633)) + ((g1285) & (g1585) & (g1591) & (!g1600) & (!g1633)) + ((g1285) & (g1585) & (g1591) & (!g1600) & (g1633)) + ((g1285) & (g1585) & (g1591) & (g1600) & (!g1633)) + ((g1285) & (g1585) & (g1591) & (g1600) & (g1633)));
	assign g1659 = (((!g1437) & (!g1423) & (g1588) & (g1590)) + ((!g1437) & (g1423) & (!g1588) & (g1590)) + ((!g1437) & (g1423) & (g1588) & (!g1590)) + ((!g1437) & (g1423) & (g1588) & (g1590)) + ((g1437) & (!g1423) & (!g1588) & (!g1590)) + ((g1437) & (!g1423) & (!g1588) & (g1590)) + ((g1437) & (!g1423) & (g1588) & (!g1590)) + ((g1437) & (g1423) & (!g1588) & (!g1590)));
	assign g1660 = (((!g1587) & (!g1600) & (!g1633) & (g1659)) + ((!g1587) & (g1600) & (!g1633) & (g1659)) + ((!g1587) & (g1600) & (g1633) & (g1659)) + ((g1587) & (!g1600) & (!g1633) & (!g1659)) + ((g1587) & (!g1600) & (g1633) & (!g1659)) + ((g1587) & (!g1600) & (g1633) & (g1659)) + ((g1587) & (g1600) & (!g1633) & (!g1659)) + ((g1587) & (g1600) & (g1633) & (!g1659)));
	assign g1661 = (((!g1423) & (!g1588) & (g1590) & (!g1600) & (!g1633)) + ((!g1423) & (!g1588) & (g1590) & (g1600) & (!g1633)) + ((!g1423) & (!g1588) & (g1590) & (g1600) & (g1633)) + ((!g1423) & (g1588) & (!g1590) & (!g1600) & (!g1633)) + ((!g1423) & (g1588) & (!g1590) & (!g1600) & (g1633)) + ((!g1423) & (g1588) & (!g1590) & (g1600) & (!g1633)) + ((!g1423) & (g1588) & (!g1590) & (g1600) & (g1633)) + ((!g1423) & (g1588) & (g1590) & (!g1600) & (g1633)) + ((g1423) & (!g1588) & (!g1590) & (!g1600) & (!g1633)) + ((g1423) & (!g1588) & (!g1590) & (g1600) & (!g1633)) + ((g1423) & (!g1588) & (!g1590) & (g1600) & (g1633)) + ((g1423) & (g1588) & (!g1590) & (!g1600) & (g1633)) + ((g1423) & (g1588) & (g1590) & (!g1600) & (!g1633)) + ((g1423) & (g1588) & (g1590) & (!g1600) & (g1633)) + ((g1423) & (g1588) & (g1590) & (g1600) & (!g1633)) + ((g1423) & (g1588) & (g1590) & (g1600) & (g1633)));
	assign g1662 = (((!g1586) & (!ax44x) & (!g1568) & (g1589)) + ((!g1586) & (!ax44x) & (g1568) & (g1589)) + ((!g1586) & (ax44x) & (!g1568) & (!g1589)) + ((!g1586) & (ax44x) & (!g1568) & (g1589)) + ((g1586) & (!ax44x) & (!g1568) & (!g1589)) + ((g1586) & (!ax44x) & (g1568) & (!g1589)) + ((g1586) & (ax44x) & (g1568) & (!g1589)) + ((g1586) & (ax44x) & (g1568) & (g1589)));
	assign g1663 = (((!ax44x) & (!ax45x) & (!g1568) & (!g1600) & (!g1633) & (g1662)) + ((!ax44x) & (!ax45x) & (!g1568) & (!g1600) & (g1633) & (!g1662)) + ((!ax44x) & (!ax45x) & (!g1568) & (!g1600) & (g1633) & (g1662)) + ((!ax44x) & (!ax45x) & (!g1568) & (g1600) & (!g1633) & (g1662)) + ((!ax44x) & (!ax45x) & (!g1568) & (g1600) & (g1633) & (g1662)) + ((!ax44x) & (!ax45x) & (g1568) & (!g1600) & (!g1633) & (!g1662)) + ((!ax44x) & (!ax45x) & (g1568) & (g1600) & (!g1633) & (!g1662)) + ((!ax44x) & (!ax45x) & (g1568) & (g1600) & (g1633) & (!g1662)) + ((!ax44x) & (ax45x) & (!g1568) & (!g1600) & (!g1633) & (!g1662)) + ((!ax44x) & (ax45x) & (!g1568) & (g1600) & (!g1633) & (!g1662)) + ((!ax44x) & (ax45x) & (!g1568) & (g1600) & (g1633) & (!g1662)) + ((!ax44x) & (ax45x) & (g1568) & (!g1600) & (!g1633) & (g1662)) + ((!ax44x) & (ax45x) & (g1568) & (!g1600) & (g1633) & (!g1662)) + ((!ax44x) & (ax45x) & (g1568) & (!g1600) & (g1633) & (g1662)) + ((!ax44x) & (ax45x) & (g1568) & (g1600) & (!g1633) & (g1662)) + ((!ax44x) & (ax45x) & (g1568) & (g1600) & (g1633) & (g1662)) + ((ax44x) & (!ax45x) & (!g1568) & (!g1600) & (!g1633) & (!g1662)) + ((ax44x) & (!ax45x) & (!g1568) & (g1600) & (!g1633) & (!g1662)) + ((ax44x) & (!ax45x) & (!g1568) & (g1600) & (g1633) & (!g1662)) + ((ax44x) & (!ax45x) & (g1568) & (!g1600) & (!g1633) & (!g1662)) + ((ax44x) & (!ax45x) & (g1568) & (g1600) & (!g1633) & (!g1662)) + ((ax44x) & (!ax45x) & (g1568) & (g1600) & (g1633) & (!g1662)) + ((ax44x) & (ax45x) & (!g1568) & (!g1600) & (!g1633) & (g1662)) + ((ax44x) & (ax45x) & (!g1568) & (!g1600) & (g1633) & (!g1662)) + ((ax44x) & (ax45x) & (!g1568) & (!g1600) & (g1633) & (g1662)) + ((ax44x) & (ax45x) & (!g1568) & (g1600) & (!g1633) & (g1662)) + ((ax44x) & (ax45x) & (!g1568) & (g1600) & (g1633) & (g1662)) + ((ax44x) & (ax45x) & (g1568) & (!g1600) & (!g1633) & (g1662)) + ((ax44x) & (ax45x) & (g1568) & (!g1600) & (g1633) & (!g1662)) + ((ax44x) & (ax45x) & (g1568) & (!g1600) & (g1633) & (g1662)) + ((ax44x) & (ax45x) & (g1568) & (g1600) & (!g1633) & (g1662)) + ((ax44x) & (ax45x) & (g1568) & (g1600) & (g1633) & (g1662)));
	assign g1664 = (((!ax44x) & (!g1568) & (!g1589) & (!g1600) & (g1633)) + ((!ax44x) & (!g1568) & (g1589) & (!g1600) & (!g1633)) + ((!ax44x) & (!g1568) & (g1589) & (!g1600) & (g1633)) + ((!ax44x) & (!g1568) & (g1589) & (g1600) & (!g1633)) + ((!ax44x) & (!g1568) & (g1589) & (g1600) & (g1633)) + ((!ax44x) & (g1568) & (g1589) & (!g1600) & (!g1633)) + ((!ax44x) & (g1568) & (g1589) & (g1600) & (!g1633)) + ((!ax44x) & (g1568) & (g1589) & (g1600) & (g1633)) + ((ax44x) & (!g1568) & (!g1589) & (!g1600) & (!g1633)) + ((ax44x) & (!g1568) & (!g1589) & (g1600) & (!g1633)) + ((ax44x) & (!g1568) & (!g1589) & (g1600) & (g1633)) + ((ax44x) & (g1568) & (!g1589) & (!g1600) & (!g1633)) + ((ax44x) & (g1568) & (!g1589) & (!g1600) & (g1633)) + ((ax44x) & (g1568) & (!g1589) & (g1600) & (!g1633)) + ((ax44x) & (g1568) & (!g1589) & (g1600) & (g1633)) + ((ax44x) & (g1568) & (g1589) & (!g1600) & (g1633)));
	assign g1665 = (((!ax40x) & (!ax41x)));
	assign g1666 = (((!g1568) & (!ax42x) & (!ax43x) & (!g1600) & (!g1633) & (!g1665)) + ((!g1568) & (!ax42x) & (!ax43x) & (g1600) & (!g1633) & (!g1665)) + ((!g1568) & (!ax42x) & (!ax43x) & (g1600) & (g1633) & (!g1665)) + ((!g1568) & (!ax42x) & (ax43x) & (!g1600) & (g1633) & (!g1665)) + ((!g1568) & (ax42x) & (ax43x) & (!g1600) & (g1633) & (!g1665)) + ((!g1568) & (ax42x) & (ax43x) & (!g1600) & (g1633) & (g1665)) + ((g1568) & (!ax42x) & (!ax43x) & (!g1600) & (!g1633) & (!g1665)) + ((g1568) & (!ax42x) & (!ax43x) & (!g1600) & (!g1633) & (g1665)) + ((g1568) & (!ax42x) & (!ax43x) & (!g1600) & (g1633) & (!g1665)) + ((g1568) & (!ax42x) & (!ax43x) & (g1600) & (!g1633) & (!g1665)) + ((g1568) & (!ax42x) & (!ax43x) & (g1600) & (!g1633) & (g1665)) + ((g1568) & (!ax42x) & (!ax43x) & (g1600) & (g1633) & (!g1665)) + ((g1568) & (!ax42x) & (!ax43x) & (g1600) & (g1633) & (g1665)) + ((g1568) & (!ax42x) & (ax43x) & (!g1600) & (!g1633) & (!g1665)) + ((g1568) & (!ax42x) & (ax43x) & (!g1600) & (g1633) & (!g1665)) + ((g1568) & (!ax42x) & (ax43x) & (!g1600) & (g1633) & (g1665)) + ((g1568) & (!ax42x) & (ax43x) & (g1600) & (!g1633) & (!g1665)) + ((g1568) & (!ax42x) & (ax43x) & (g1600) & (g1633) & (!g1665)) + ((g1568) & (ax42x) & (!ax43x) & (!g1600) & (g1633) & (!g1665)) + ((g1568) & (ax42x) & (!ax43x) & (!g1600) & (g1633) & (g1665)) + ((g1568) & (ax42x) & (ax43x) & (!g1600) & (!g1633) & (!g1665)) + ((g1568) & (ax42x) & (ax43x) & (!g1600) & (!g1633) & (g1665)) + ((g1568) & (ax42x) & (ax43x) & (!g1600) & (g1633) & (!g1665)) + ((g1568) & (ax42x) & (ax43x) & (!g1600) & (g1633) & (g1665)) + ((g1568) & (ax42x) & (ax43x) & (g1600) & (!g1633) & (!g1665)) + ((g1568) & (ax42x) & (ax43x) & (g1600) & (!g1633) & (g1665)) + ((g1568) & (ax42x) & (ax43x) & (g1600) & (g1633) & (!g1665)) + ((g1568) & (ax42x) & (ax43x) & (g1600) & (g1633) & (g1665)));
	assign g1667 = (((!g1423) & (!g1586) & (g1663) & (g1664) & (g1666)) + ((!g1423) & (g1586) & (g1663) & (!g1664) & (g1666)) + ((!g1423) & (g1586) & (g1663) & (g1664) & (!g1666)) + ((!g1423) & (g1586) & (g1663) & (g1664) & (g1666)) + ((g1423) & (!g1586) & (!g1663) & (g1664) & (g1666)) + ((g1423) & (!g1586) & (g1663) & (!g1664) & (!g1666)) + ((g1423) & (!g1586) & (g1663) & (!g1664) & (g1666)) + ((g1423) & (!g1586) & (g1663) & (g1664) & (!g1666)) + ((g1423) & (!g1586) & (g1663) & (g1664) & (g1666)) + ((g1423) & (g1586) & (!g1663) & (!g1664) & (g1666)) + ((g1423) & (g1586) & (!g1663) & (g1664) & (!g1666)) + ((g1423) & (g1586) & (!g1663) & (g1664) & (g1666)) + ((g1423) & (g1586) & (g1663) & (!g1664) & (!g1666)) + ((g1423) & (g1586) & (g1663) & (!g1664) & (g1666)) + ((g1423) & (g1586) & (g1663) & (g1664) & (!g1666)) + ((g1423) & (g1586) & (g1663) & (g1664) & (g1666)));
	assign g1668 = (((!g1285) & (!g1437) & (g1660) & (g1661) & (g1667)) + ((!g1285) & (g1437) & (g1660) & (!g1661) & (g1667)) + ((!g1285) & (g1437) & (g1660) & (g1661) & (!g1667)) + ((!g1285) & (g1437) & (g1660) & (g1661) & (g1667)) + ((g1285) & (!g1437) & (!g1660) & (g1661) & (g1667)) + ((g1285) & (!g1437) & (g1660) & (!g1661) & (!g1667)) + ((g1285) & (!g1437) & (g1660) & (!g1661) & (g1667)) + ((g1285) & (!g1437) & (g1660) & (g1661) & (!g1667)) + ((g1285) & (!g1437) & (g1660) & (g1661) & (g1667)) + ((g1285) & (g1437) & (!g1660) & (!g1661) & (g1667)) + ((g1285) & (g1437) & (!g1660) & (g1661) & (!g1667)) + ((g1285) & (g1437) & (!g1660) & (g1661) & (g1667)) + ((g1285) & (g1437) & (g1660) & (!g1661) & (!g1667)) + ((g1285) & (g1437) & (g1660) & (!g1661) & (g1667)) + ((g1285) & (g1437) & (g1660) & (g1661) & (!g1667)) + ((g1285) & (g1437) & (g1660) & (g1661) & (g1667)));
	assign g1669 = (((!g1154) & (!g1295) & (g1657) & (g1658) & (g1668)) + ((!g1154) & (g1295) & (g1657) & (!g1658) & (g1668)) + ((!g1154) & (g1295) & (g1657) & (g1658) & (!g1668)) + ((!g1154) & (g1295) & (g1657) & (g1658) & (g1668)) + ((g1154) & (!g1295) & (!g1657) & (g1658) & (g1668)) + ((g1154) & (!g1295) & (g1657) & (!g1658) & (!g1668)) + ((g1154) & (!g1295) & (g1657) & (!g1658) & (g1668)) + ((g1154) & (!g1295) & (g1657) & (g1658) & (!g1668)) + ((g1154) & (!g1295) & (g1657) & (g1658) & (g1668)) + ((g1154) & (g1295) & (!g1657) & (!g1658) & (g1668)) + ((g1154) & (g1295) & (!g1657) & (g1658) & (!g1668)) + ((g1154) & (g1295) & (!g1657) & (g1658) & (g1668)) + ((g1154) & (g1295) & (g1657) & (!g1658) & (!g1668)) + ((g1154) & (g1295) & (g1657) & (!g1658) & (g1668)) + ((g1154) & (g1295) & (g1657) & (g1658) & (!g1668)) + ((g1154) & (g1295) & (g1657) & (g1658) & (g1668)));
	assign g1670 = (((!g1030) & (!g1160) & (g1654) & (g1655) & (g1669)) + ((!g1030) & (g1160) & (g1654) & (!g1655) & (g1669)) + ((!g1030) & (g1160) & (g1654) & (g1655) & (!g1669)) + ((!g1030) & (g1160) & (g1654) & (g1655) & (g1669)) + ((g1030) & (!g1160) & (!g1654) & (g1655) & (g1669)) + ((g1030) & (!g1160) & (g1654) & (!g1655) & (!g1669)) + ((g1030) & (!g1160) & (g1654) & (!g1655) & (g1669)) + ((g1030) & (!g1160) & (g1654) & (g1655) & (!g1669)) + ((g1030) & (!g1160) & (g1654) & (g1655) & (g1669)) + ((g1030) & (g1160) & (!g1654) & (!g1655) & (g1669)) + ((g1030) & (g1160) & (!g1654) & (g1655) & (!g1669)) + ((g1030) & (g1160) & (!g1654) & (g1655) & (g1669)) + ((g1030) & (g1160) & (g1654) & (!g1655) & (!g1669)) + ((g1030) & (g1160) & (g1654) & (!g1655) & (g1669)) + ((g1030) & (g1160) & (g1654) & (g1655) & (!g1669)) + ((g1030) & (g1160) & (g1654) & (g1655) & (g1669)));
	assign g1671 = (((!g914) & (!g1032) & (g1651) & (g1652) & (g1670)) + ((!g914) & (g1032) & (g1651) & (!g1652) & (g1670)) + ((!g914) & (g1032) & (g1651) & (g1652) & (!g1670)) + ((!g914) & (g1032) & (g1651) & (g1652) & (g1670)) + ((g914) & (!g1032) & (!g1651) & (g1652) & (g1670)) + ((g914) & (!g1032) & (g1651) & (!g1652) & (!g1670)) + ((g914) & (!g1032) & (g1651) & (!g1652) & (g1670)) + ((g914) & (!g1032) & (g1651) & (g1652) & (!g1670)) + ((g914) & (!g1032) & (g1651) & (g1652) & (g1670)) + ((g914) & (g1032) & (!g1651) & (!g1652) & (g1670)) + ((g914) & (g1032) & (!g1651) & (g1652) & (!g1670)) + ((g914) & (g1032) & (!g1651) & (g1652) & (g1670)) + ((g914) & (g1032) & (g1651) & (!g1652) & (!g1670)) + ((g914) & (g1032) & (g1651) & (!g1652) & (g1670)) + ((g914) & (g1032) & (g1651) & (g1652) & (!g1670)) + ((g914) & (g1032) & (g1651) & (g1652) & (g1670)));
	assign g1672 = (((!g803) & (!g851) & (g1648) & (g1649) & (g1671)) + ((!g803) & (g851) & (g1648) & (!g1649) & (g1671)) + ((!g803) & (g851) & (g1648) & (g1649) & (!g1671)) + ((!g803) & (g851) & (g1648) & (g1649) & (g1671)) + ((g803) & (!g851) & (!g1648) & (g1649) & (g1671)) + ((g803) & (!g851) & (g1648) & (!g1649) & (!g1671)) + ((g803) & (!g851) & (g1648) & (!g1649) & (g1671)) + ((g803) & (!g851) & (g1648) & (g1649) & (!g1671)) + ((g803) & (!g851) & (g1648) & (g1649) & (g1671)) + ((g803) & (g851) & (!g1648) & (!g1649) & (g1671)) + ((g803) & (g851) & (!g1648) & (g1649) & (!g1671)) + ((g803) & (g851) & (!g1648) & (g1649) & (g1671)) + ((g803) & (g851) & (g1648) & (!g1649) & (!g1671)) + ((g803) & (g851) & (g1648) & (!g1649) & (g1671)) + ((g803) & (g851) & (g1648) & (g1649) & (!g1671)) + ((g803) & (g851) & (g1648) & (g1649) & (g1671)));
	assign g1673 = (((!g700) & (!g744) & (g1645) & (g1646) & (g1672)) + ((!g700) & (g744) & (g1645) & (!g1646) & (g1672)) + ((!g700) & (g744) & (g1645) & (g1646) & (!g1672)) + ((!g700) & (g744) & (g1645) & (g1646) & (g1672)) + ((g700) & (!g744) & (!g1645) & (g1646) & (g1672)) + ((g700) & (!g744) & (g1645) & (!g1646) & (!g1672)) + ((g700) & (!g744) & (g1645) & (!g1646) & (g1672)) + ((g700) & (!g744) & (g1645) & (g1646) & (!g1672)) + ((g700) & (!g744) & (g1645) & (g1646) & (g1672)) + ((g700) & (g744) & (!g1645) & (!g1646) & (g1672)) + ((g700) & (g744) & (!g1645) & (g1646) & (!g1672)) + ((g700) & (g744) & (!g1645) & (g1646) & (g1672)) + ((g700) & (g744) & (g1645) & (!g1646) & (!g1672)) + ((g700) & (g744) & (g1645) & (!g1646) & (g1672)) + ((g700) & (g744) & (g1645) & (g1646) & (!g1672)) + ((g700) & (g744) & (g1645) & (g1646) & (g1672)));
	assign g1674 = (((!g604) & (!g645) & (g1642) & (g1643) & (g1673)) + ((!g604) & (g645) & (g1642) & (!g1643) & (g1673)) + ((!g604) & (g645) & (g1642) & (g1643) & (!g1673)) + ((!g604) & (g645) & (g1642) & (g1643) & (g1673)) + ((g604) & (!g645) & (!g1642) & (g1643) & (g1673)) + ((g604) & (!g645) & (g1642) & (!g1643) & (!g1673)) + ((g604) & (!g645) & (g1642) & (!g1643) & (g1673)) + ((g604) & (!g645) & (g1642) & (g1643) & (!g1673)) + ((g604) & (!g645) & (g1642) & (g1643) & (g1673)) + ((g604) & (g645) & (!g1642) & (!g1643) & (g1673)) + ((g604) & (g645) & (!g1642) & (g1643) & (!g1673)) + ((g604) & (g645) & (!g1642) & (g1643) & (g1673)) + ((g604) & (g645) & (g1642) & (!g1643) & (!g1673)) + ((g604) & (g645) & (g1642) & (!g1643) & (g1673)) + ((g604) & (g645) & (g1642) & (g1643) & (!g1673)) + ((g604) & (g645) & (g1642) & (g1643) & (g1673)));
	assign g1675 = (((!g515) & (!g553) & (g1639) & (g1640) & (g1674)) + ((!g515) & (g553) & (g1639) & (!g1640) & (g1674)) + ((!g515) & (g553) & (g1639) & (g1640) & (!g1674)) + ((!g515) & (g553) & (g1639) & (g1640) & (g1674)) + ((g515) & (!g553) & (!g1639) & (g1640) & (g1674)) + ((g515) & (!g553) & (g1639) & (!g1640) & (!g1674)) + ((g515) & (!g553) & (g1639) & (!g1640) & (g1674)) + ((g515) & (!g553) & (g1639) & (g1640) & (!g1674)) + ((g515) & (!g553) & (g1639) & (g1640) & (g1674)) + ((g515) & (g553) & (!g1639) & (!g1640) & (g1674)) + ((g515) & (g553) & (!g1639) & (g1640) & (!g1674)) + ((g515) & (g553) & (!g1639) & (g1640) & (g1674)) + ((g515) & (g553) & (g1639) & (!g1640) & (!g1674)) + ((g515) & (g553) & (g1639) & (!g1640) & (g1674)) + ((g515) & (g553) & (g1639) & (g1640) & (!g1674)) + ((g515) & (g553) & (g1639) & (g1640) & (g1674)));
	assign g1676 = (((!g433) & (!g468) & (g1636) & (g1637) & (g1675)) + ((!g433) & (g468) & (g1636) & (!g1637) & (g1675)) + ((!g433) & (g468) & (g1636) & (g1637) & (!g1675)) + ((!g433) & (g468) & (g1636) & (g1637) & (g1675)) + ((g433) & (!g468) & (!g1636) & (g1637) & (g1675)) + ((g433) & (!g468) & (g1636) & (!g1637) & (!g1675)) + ((g433) & (!g468) & (g1636) & (!g1637) & (g1675)) + ((g433) & (!g468) & (g1636) & (g1637) & (!g1675)) + ((g433) & (!g468) & (g1636) & (g1637) & (g1675)) + ((g433) & (g468) & (!g1636) & (!g1637) & (g1675)) + ((g433) & (g468) & (!g1636) & (g1637) & (!g1675)) + ((g433) & (g468) & (!g1636) & (g1637) & (g1675)) + ((g433) & (g468) & (g1636) & (!g1637) & (!g1675)) + ((g433) & (g468) & (g1636) & (!g1637) & (g1675)) + ((g433) & (g468) & (g1636) & (g1637) & (!g1675)) + ((g433) & (g468) & (g1636) & (g1637) & (g1675)));
	assign g1677 = (((!g4) & (!g1630) & (!g1631) & (!g1600) & (!g1633)) + ((!g4) & (!g1630) & (!g1631) & (g1600) & (!g1633)) + ((!g4) & (!g1630) & (!g1631) & (g1600) & (g1633)) + ((!g4) & (!g1630) & (g1631) & (!g1600) & (g1633)) + ((!g4) & (g1630) & (g1631) & (!g1600) & (!g1633)) + ((!g4) & (g1630) & (g1631) & (!g1600) & (g1633)) + ((!g4) & (g1630) & (g1631) & (g1600) & (!g1633)) + ((!g4) & (g1630) & (g1631) & (g1600) & (g1633)) + ((g4) & (!g1630) & (g1631) & (!g1600) & (!g1633)) + ((g4) & (!g1630) & (g1631) & (!g1600) & (g1633)) + ((g4) & (!g1630) & (g1631) & (g1600) & (!g1633)) + ((g4) & (!g1630) & (g1631) & (g1600) & (g1633)) + ((g4) & (g1630) & (!g1631) & (!g1600) & (!g1633)) + ((g4) & (g1630) & (!g1631) & (g1600) & (!g1633)) + ((g4) & (g1630) & (!g1631) & (g1600) & (g1633)) + ((g4) & (g1630) & (g1631) & (!g1600) & (g1633)));
	assign g1678 = (((!g8) & (!g1603) & (g1629) & (!g1600) & (!g1633)) + ((!g8) & (!g1603) & (g1629) & (g1600) & (!g1633)) + ((!g8) & (!g1603) & (g1629) & (g1600) & (g1633)) + ((!g8) & (g1603) & (!g1629) & (!g1600) & (!g1633)) + ((!g8) & (g1603) & (!g1629) & (!g1600) & (g1633)) + ((!g8) & (g1603) & (!g1629) & (g1600) & (!g1633)) + ((!g8) & (g1603) & (!g1629) & (g1600) & (g1633)) + ((!g8) & (g1603) & (g1629) & (!g1600) & (g1633)) + ((g8) & (!g1603) & (!g1629) & (!g1600) & (!g1633)) + ((g8) & (!g1603) & (!g1629) & (g1600) & (!g1633)) + ((g8) & (!g1603) & (!g1629) & (g1600) & (g1633)) + ((g8) & (g1603) & (!g1629) & (!g1600) & (g1633)) + ((g8) & (g1603) & (g1629) & (!g1600) & (!g1633)) + ((g8) & (g1603) & (g1629) & (!g1600) & (g1633)) + ((g8) & (g1603) & (g1629) & (g1600) & (!g1633)) + ((g8) & (g1603) & (g1629) & (g1600) & (g1633)));
	assign g1679 = (((!g18) & (!g27) & (g1605) & (g1628)) + ((!g18) & (g27) & (!g1605) & (g1628)) + ((!g18) & (g27) & (g1605) & (!g1628)) + ((!g18) & (g27) & (g1605) & (g1628)) + ((g18) & (!g27) & (!g1605) & (!g1628)) + ((g18) & (!g27) & (!g1605) & (g1628)) + ((g18) & (!g27) & (g1605) & (!g1628)) + ((g18) & (g27) & (!g1605) & (!g1628)));
	assign g1680 = (((!g1604) & (!g1600) & (!g1633) & (g1679)) + ((!g1604) & (g1600) & (!g1633) & (g1679)) + ((!g1604) & (g1600) & (g1633) & (g1679)) + ((g1604) & (!g1600) & (!g1633) & (!g1679)) + ((g1604) & (!g1600) & (g1633) & (!g1679)) + ((g1604) & (!g1600) & (g1633) & (g1679)) + ((g1604) & (g1600) & (!g1633) & (!g1679)) + ((g1604) & (g1600) & (g1633) & (!g1679)));
	assign g1681 = (((!g27) & (!g1605) & (g1628) & (!g1600) & (!g1633)) + ((!g27) & (!g1605) & (g1628) & (g1600) & (!g1633)) + ((!g27) & (!g1605) & (g1628) & (g1600) & (g1633)) + ((!g27) & (g1605) & (!g1628) & (!g1600) & (!g1633)) + ((!g27) & (g1605) & (!g1628) & (!g1600) & (g1633)) + ((!g27) & (g1605) & (!g1628) & (g1600) & (!g1633)) + ((!g27) & (g1605) & (!g1628) & (g1600) & (g1633)) + ((!g27) & (g1605) & (g1628) & (!g1600) & (g1633)) + ((g27) & (!g1605) & (!g1628) & (!g1600) & (!g1633)) + ((g27) & (!g1605) & (!g1628) & (g1600) & (!g1633)) + ((g27) & (!g1605) & (!g1628) & (g1600) & (g1633)) + ((g27) & (g1605) & (!g1628) & (!g1600) & (g1633)) + ((g27) & (g1605) & (g1628) & (!g1600) & (!g1633)) + ((g27) & (g1605) & (g1628) & (!g1600) & (g1633)) + ((g27) & (g1605) & (g1628) & (g1600) & (!g1633)) + ((g27) & (g1605) & (g1628) & (g1600) & (g1633)));
	assign g1682 = (((!g39) & (!g54) & (g1607) & (g1627)) + ((!g39) & (g54) & (!g1607) & (g1627)) + ((!g39) & (g54) & (g1607) & (!g1627)) + ((!g39) & (g54) & (g1607) & (g1627)) + ((g39) & (!g54) & (!g1607) & (!g1627)) + ((g39) & (!g54) & (!g1607) & (g1627)) + ((g39) & (!g54) & (g1607) & (!g1627)) + ((g39) & (g54) & (!g1607) & (!g1627)));
	assign g1683 = (((!g1606) & (!g1600) & (!g1633) & (g1682)) + ((!g1606) & (g1600) & (!g1633) & (g1682)) + ((!g1606) & (g1600) & (g1633) & (g1682)) + ((g1606) & (!g1600) & (!g1633) & (!g1682)) + ((g1606) & (!g1600) & (g1633) & (!g1682)) + ((g1606) & (!g1600) & (g1633) & (g1682)) + ((g1606) & (g1600) & (!g1633) & (!g1682)) + ((g1606) & (g1600) & (g1633) & (!g1682)));
	assign g1684 = (((!g54) & (!g1607) & (g1627) & (!g1600) & (!g1633)) + ((!g54) & (!g1607) & (g1627) & (g1600) & (!g1633)) + ((!g54) & (!g1607) & (g1627) & (g1600) & (g1633)) + ((!g54) & (g1607) & (!g1627) & (!g1600) & (!g1633)) + ((!g54) & (g1607) & (!g1627) & (!g1600) & (g1633)) + ((!g54) & (g1607) & (!g1627) & (g1600) & (!g1633)) + ((!g54) & (g1607) & (!g1627) & (g1600) & (g1633)) + ((!g54) & (g1607) & (g1627) & (!g1600) & (g1633)) + ((g54) & (!g1607) & (!g1627) & (!g1600) & (!g1633)) + ((g54) & (!g1607) & (!g1627) & (g1600) & (!g1633)) + ((g54) & (!g1607) & (!g1627) & (g1600) & (g1633)) + ((g54) & (g1607) & (!g1627) & (!g1600) & (g1633)) + ((g54) & (g1607) & (g1627) & (!g1600) & (!g1633)) + ((g54) & (g1607) & (g1627) & (!g1600) & (g1633)) + ((g54) & (g1607) & (g1627) & (g1600) & (!g1633)) + ((g54) & (g1607) & (g1627) & (g1600) & (g1633)));
	assign g1685 = (((!g68) & (!g87) & (g1609) & (g1626)) + ((!g68) & (g87) & (!g1609) & (g1626)) + ((!g68) & (g87) & (g1609) & (!g1626)) + ((!g68) & (g87) & (g1609) & (g1626)) + ((g68) & (!g87) & (!g1609) & (!g1626)) + ((g68) & (!g87) & (!g1609) & (g1626)) + ((g68) & (!g87) & (g1609) & (!g1626)) + ((g68) & (g87) & (!g1609) & (!g1626)));
	assign g1686 = (((!g1608) & (!g1600) & (!g1633) & (g1685)) + ((!g1608) & (g1600) & (!g1633) & (g1685)) + ((!g1608) & (g1600) & (g1633) & (g1685)) + ((g1608) & (!g1600) & (!g1633) & (!g1685)) + ((g1608) & (!g1600) & (g1633) & (!g1685)) + ((g1608) & (!g1600) & (g1633) & (g1685)) + ((g1608) & (g1600) & (!g1633) & (!g1685)) + ((g1608) & (g1600) & (g1633) & (!g1685)));
	assign g1687 = (((!g87) & (!g1609) & (g1626) & (!g1600) & (!g1633)) + ((!g87) & (!g1609) & (g1626) & (g1600) & (!g1633)) + ((!g87) & (!g1609) & (g1626) & (g1600) & (g1633)) + ((!g87) & (g1609) & (!g1626) & (!g1600) & (!g1633)) + ((!g87) & (g1609) & (!g1626) & (!g1600) & (g1633)) + ((!g87) & (g1609) & (!g1626) & (g1600) & (!g1633)) + ((!g87) & (g1609) & (!g1626) & (g1600) & (g1633)) + ((!g87) & (g1609) & (g1626) & (!g1600) & (g1633)) + ((g87) & (!g1609) & (!g1626) & (!g1600) & (!g1633)) + ((g87) & (!g1609) & (!g1626) & (g1600) & (!g1633)) + ((g87) & (!g1609) & (!g1626) & (g1600) & (g1633)) + ((g87) & (g1609) & (!g1626) & (!g1600) & (g1633)) + ((g87) & (g1609) & (g1626) & (!g1600) & (!g1633)) + ((g87) & (g1609) & (g1626) & (!g1600) & (g1633)) + ((g87) & (g1609) & (g1626) & (g1600) & (!g1633)) + ((g87) & (g1609) & (g1626) & (g1600) & (g1633)));
	assign g1688 = (((!g104) & (!g127) & (g1611) & (g1625)) + ((!g104) & (g127) & (!g1611) & (g1625)) + ((!g104) & (g127) & (g1611) & (!g1625)) + ((!g104) & (g127) & (g1611) & (g1625)) + ((g104) & (!g127) & (!g1611) & (!g1625)) + ((g104) & (!g127) & (!g1611) & (g1625)) + ((g104) & (!g127) & (g1611) & (!g1625)) + ((g104) & (g127) & (!g1611) & (!g1625)));
	assign g1689 = (((!g1610) & (!g1600) & (!g1633) & (g1688)) + ((!g1610) & (g1600) & (!g1633) & (g1688)) + ((!g1610) & (g1600) & (g1633) & (g1688)) + ((g1610) & (!g1600) & (!g1633) & (!g1688)) + ((g1610) & (!g1600) & (g1633) & (!g1688)) + ((g1610) & (!g1600) & (g1633) & (g1688)) + ((g1610) & (g1600) & (!g1633) & (!g1688)) + ((g1610) & (g1600) & (g1633) & (!g1688)));
	assign g1690 = (((!g127) & (!g1611) & (g1625) & (!g1600) & (!g1633)) + ((!g127) & (!g1611) & (g1625) & (g1600) & (!g1633)) + ((!g127) & (!g1611) & (g1625) & (g1600) & (g1633)) + ((!g127) & (g1611) & (!g1625) & (!g1600) & (!g1633)) + ((!g127) & (g1611) & (!g1625) & (!g1600) & (g1633)) + ((!g127) & (g1611) & (!g1625) & (g1600) & (!g1633)) + ((!g127) & (g1611) & (!g1625) & (g1600) & (g1633)) + ((!g127) & (g1611) & (g1625) & (!g1600) & (g1633)) + ((g127) & (!g1611) & (!g1625) & (!g1600) & (!g1633)) + ((g127) & (!g1611) & (!g1625) & (g1600) & (!g1633)) + ((g127) & (!g1611) & (!g1625) & (g1600) & (g1633)) + ((g127) & (g1611) & (!g1625) & (!g1600) & (g1633)) + ((g127) & (g1611) & (g1625) & (!g1600) & (!g1633)) + ((g127) & (g1611) & (g1625) & (!g1600) & (g1633)) + ((g127) & (g1611) & (g1625) & (g1600) & (!g1633)) + ((g127) & (g1611) & (g1625) & (g1600) & (g1633)));
	assign g1691 = (((!g147) & (!g174) & (g1613) & (g1624)) + ((!g147) & (g174) & (!g1613) & (g1624)) + ((!g147) & (g174) & (g1613) & (!g1624)) + ((!g147) & (g174) & (g1613) & (g1624)) + ((g147) & (!g174) & (!g1613) & (!g1624)) + ((g147) & (!g174) & (!g1613) & (g1624)) + ((g147) & (!g174) & (g1613) & (!g1624)) + ((g147) & (g174) & (!g1613) & (!g1624)));
	assign g1692 = (((!g1612) & (!g1600) & (!g1633) & (g1691)) + ((!g1612) & (g1600) & (!g1633) & (g1691)) + ((!g1612) & (g1600) & (g1633) & (g1691)) + ((g1612) & (!g1600) & (!g1633) & (!g1691)) + ((g1612) & (!g1600) & (g1633) & (!g1691)) + ((g1612) & (!g1600) & (g1633) & (g1691)) + ((g1612) & (g1600) & (!g1633) & (!g1691)) + ((g1612) & (g1600) & (g1633) & (!g1691)));
	assign g1693 = (((!g174) & (!g1613) & (g1624) & (!g1600) & (!g1633)) + ((!g174) & (!g1613) & (g1624) & (g1600) & (!g1633)) + ((!g174) & (!g1613) & (g1624) & (g1600) & (g1633)) + ((!g174) & (g1613) & (!g1624) & (!g1600) & (!g1633)) + ((!g174) & (g1613) & (!g1624) & (!g1600) & (g1633)) + ((!g174) & (g1613) & (!g1624) & (g1600) & (!g1633)) + ((!g174) & (g1613) & (!g1624) & (g1600) & (g1633)) + ((!g174) & (g1613) & (g1624) & (!g1600) & (g1633)) + ((g174) & (!g1613) & (!g1624) & (!g1600) & (!g1633)) + ((g174) & (!g1613) & (!g1624) & (g1600) & (!g1633)) + ((g174) & (!g1613) & (!g1624) & (g1600) & (g1633)) + ((g174) & (g1613) & (!g1624) & (!g1600) & (g1633)) + ((g174) & (g1613) & (g1624) & (!g1600) & (!g1633)) + ((g174) & (g1613) & (g1624) & (!g1600) & (g1633)) + ((g174) & (g1613) & (g1624) & (g1600) & (!g1633)) + ((g174) & (g1613) & (g1624) & (g1600) & (g1633)));
	assign g1694 = (((!g198) & (!g229) & (g1615) & (g1623)) + ((!g198) & (g229) & (!g1615) & (g1623)) + ((!g198) & (g229) & (g1615) & (!g1623)) + ((!g198) & (g229) & (g1615) & (g1623)) + ((g198) & (!g229) & (!g1615) & (!g1623)) + ((g198) & (!g229) & (!g1615) & (g1623)) + ((g198) & (!g229) & (g1615) & (!g1623)) + ((g198) & (g229) & (!g1615) & (!g1623)));
	assign g1695 = (((!g1614) & (!g1600) & (!g1633) & (g1694)) + ((!g1614) & (g1600) & (!g1633) & (g1694)) + ((!g1614) & (g1600) & (g1633) & (g1694)) + ((g1614) & (!g1600) & (!g1633) & (!g1694)) + ((g1614) & (!g1600) & (g1633) & (!g1694)) + ((g1614) & (!g1600) & (g1633) & (g1694)) + ((g1614) & (g1600) & (!g1633) & (!g1694)) + ((g1614) & (g1600) & (g1633) & (!g1694)));
	assign g1696 = (((!g229) & (!g1615) & (g1623) & (!g1600) & (!g1633)) + ((!g229) & (!g1615) & (g1623) & (g1600) & (!g1633)) + ((!g229) & (!g1615) & (g1623) & (g1600) & (g1633)) + ((!g229) & (g1615) & (!g1623) & (!g1600) & (!g1633)) + ((!g229) & (g1615) & (!g1623) & (!g1600) & (g1633)) + ((!g229) & (g1615) & (!g1623) & (g1600) & (!g1633)) + ((!g229) & (g1615) & (!g1623) & (g1600) & (g1633)) + ((!g229) & (g1615) & (g1623) & (!g1600) & (g1633)) + ((g229) & (!g1615) & (!g1623) & (!g1600) & (!g1633)) + ((g229) & (!g1615) & (!g1623) & (g1600) & (!g1633)) + ((g229) & (!g1615) & (!g1623) & (g1600) & (g1633)) + ((g229) & (g1615) & (!g1623) & (!g1600) & (g1633)) + ((g229) & (g1615) & (g1623) & (!g1600) & (!g1633)) + ((g229) & (g1615) & (g1623) & (!g1600) & (g1633)) + ((g229) & (g1615) & (g1623) & (g1600) & (!g1633)) + ((g229) & (g1615) & (g1623) & (g1600) & (g1633)));
	assign g1697 = (((!g255) & (!g290) & (g1617) & (g1622)) + ((!g255) & (g290) & (!g1617) & (g1622)) + ((!g255) & (g290) & (g1617) & (!g1622)) + ((!g255) & (g290) & (g1617) & (g1622)) + ((g255) & (!g290) & (!g1617) & (!g1622)) + ((g255) & (!g290) & (!g1617) & (g1622)) + ((g255) & (!g290) & (g1617) & (!g1622)) + ((g255) & (g290) & (!g1617) & (!g1622)));
	assign g1698 = (((!g1616) & (!g1600) & (!g1633) & (g1697)) + ((!g1616) & (g1600) & (!g1633) & (g1697)) + ((!g1616) & (g1600) & (g1633) & (g1697)) + ((g1616) & (!g1600) & (!g1633) & (!g1697)) + ((g1616) & (!g1600) & (g1633) & (!g1697)) + ((g1616) & (!g1600) & (g1633) & (g1697)) + ((g1616) & (g1600) & (!g1633) & (!g1697)) + ((g1616) & (g1600) & (g1633) & (!g1697)));
	assign g1699 = (((!g290) & (!g1617) & (g1622) & (!g1600) & (!g1633)) + ((!g290) & (!g1617) & (g1622) & (g1600) & (!g1633)) + ((!g290) & (!g1617) & (g1622) & (g1600) & (g1633)) + ((!g290) & (g1617) & (!g1622) & (!g1600) & (!g1633)) + ((!g290) & (g1617) & (!g1622) & (!g1600) & (g1633)) + ((!g290) & (g1617) & (!g1622) & (g1600) & (!g1633)) + ((!g290) & (g1617) & (!g1622) & (g1600) & (g1633)) + ((!g290) & (g1617) & (g1622) & (!g1600) & (g1633)) + ((g290) & (!g1617) & (!g1622) & (!g1600) & (!g1633)) + ((g290) & (!g1617) & (!g1622) & (g1600) & (!g1633)) + ((g290) & (!g1617) & (!g1622) & (g1600) & (g1633)) + ((g290) & (g1617) & (!g1622) & (!g1600) & (g1633)) + ((g290) & (g1617) & (g1622) & (!g1600) & (!g1633)) + ((g290) & (g1617) & (g1622) & (!g1600) & (g1633)) + ((g290) & (g1617) & (g1622) & (g1600) & (!g1633)) + ((g290) & (g1617) & (g1622) & (g1600) & (g1633)));
	assign g1700 = (((!g319) & (!g358) & (g1619) & (g1621)) + ((!g319) & (g358) & (!g1619) & (g1621)) + ((!g319) & (g358) & (g1619) & (!g1621)) + ((!g319) & (g358) & (g1619) & (g1621)) + ((g319) & (!g358) & (!g1619) & (!g1621)) + ((g319) & (!g358) & (!g1619) & (g1621)) + ((g319) & (!g358) & (g1619) & (!g1621)) + ((g319) & (g358) & (!g1619) & (!g1621)));
	assign g1701 = (((!g1618) & (!g1600) & (!g1633) & (g1700)) + ((!g1618) & (g1600) & (!g1633) & (g1700)) + ((!g1618) & (g1600) & (g1633) & (g1700)) + ((g1618) & (!g1600) & (!g1633) & (!g1700)) + ((g1618) & (!g1600) & (g1633) & (!g1700)) + ((g1618) & (!g1600) & (g1633) & (g1700)) + ((g1618) & (g1600) & (!g1633) & (!g1700)) + ((g1618) & (g1600) & (g1633) & (!g1700)));
	assign g1702 = (((!g358) & (!g1619) & (g1621) & (!g1600) & (!g1633)) + ((!g358) & (!g1619) & (g1621) & (g1600) & (!g1633)) + ((!g358) & (!g1619) & (g1621) & (g1600) & (g1633)) + ((!g358) & (g1619) & (!g1621) & (!g1600) & (!g1633)) + ((!g358) & (g1619) & (!g1621) & (!g1600) & (g1633)) + ((!g358) & (g1619) & (!g1621) & (g1600) & (!g1633)) + ((!g358) & (g1619) & (!g1621) & (g1600) & (g1633)) + ((!g358) & (g1619) & (g1621) & (!g1600) & (g1633)) + ((g358) & (!g1619) & (!g1621) & (!g1600) & (!g1633)) + ((g358) & (!g1619) & (!g1621) & (g1600) & (!g1633)) + ((g358) & (!g1619) & (!g1621) & (g1600) & (g1633)) + ((g358) & (g1619) & (!g1621) & (!g1600) & (g1633)) + ((g358) & (g1619) & (g1621) & (!g1600) & (!g1633)) + ((g358) & (g1619) & (g1621) & (!g1600) & (g1633)) + ((g358) & (g1619) & (g1621) & (g1600) & (!g1633)) + ((g358) & (g1619) & (g1621) & (g1600) & (g1633)));
	assign g1703 = (((!g390) & (!g433) & (g1569) & (g1599)) + ((!g390) & (g433) & (!g1569) & (g1599)) + ((!g390) & (g433) & (g1569) & (!g1599)) + ((!g390) & (g433) & (g1569) & (g1599)) + ((g390) & (!g433) & (!g1569) & (!g1599)) + ((g390) & (!g433) & (!g1569) & (g1599)) + ((g390) & (!g433) & (g1569) & (!g1599)) + ((g390) & (g433) & (!g1569) & (!g1599)));
	assign g1704 = (((!g1620) & (!g1600) & (!g1633) & (g1703)) + ((!g1620) & (g1600) & (!g1633) & (g1703)) + ((!g1620) & (g1600) & (g1633) & (g1703)) + ((g1620) & (!g1600) & (!g1633) & (!g1703)) + ((g1620) & (!g1600) & (g1633) & (!g1703)) + ((g1620) & (!g1600) & (g1633) & (g1703)) + ((g1620) & (g1600) & (!g1633) & (!g1703)) + ((g1620) & (g1600) & (g1633) & (!g1703)));
	assign g1705 = (((!g358) & (!g390) & (g1704) & (g1634) & (g1676)) + ((!g358) & (g390) & (g1704) & (!g1634) & (g1676)) + ((!g358) & (g390) & (g1704) & (g1634) & (!g1676)) + ((!g358) & (g390) & (g1704) & (g1634) & (g1676)) + ((g358) & (!g390) & (!g1704) & (g1634) & (g1676)) + ((g358) & (!g390) & (g1704) & (!g1634) & (!g1676)) + ((g358) & (!g390) & (g1704) & (!g1634) & (g1676)) + ((g358) & (!g390) & (g1704) & (g1634) & (!g1676)) + ((g358) & (!g390) & (g1704) & (g1634) & (g1676)) + ((g358) & (g390) & (!g1704) & (!g1634) & (g1676)) + ((g358) & (g390) & (!g1704) & (g1634) & (!g1676)) + ((g358) & (g390) & (!g1704) & (g1634) & (g1676)) + ((g358) & (g390) & (g1704) & (!g1634) & (!g1676)) + ((g358) & (g390) & (g1704) & (!g1634) & (g1676)) + ((g358) & (g390) & (g1704) & (g1634) & (!g1676)) + ((g358) & (g390) & (g1704) & (g1634) & (g1676)));
	assign g1706 = (((!g290) & (!g319) & (g1701) & (g1702) & (g1705)) + ((!g290) & (g319) & (g1701) & (!g1702) & (g1705)) + ((!g290) & (g319) & (g1701) & (g1702) & (!g1705)) + ((!g290) & (g319) & (g1701) & (g1702) & (g1705)) + ((g290) & (!g319) & (!g1701) & (g1702) & (g1705)) + ((g290) & (!g319) & (g1701) & (!g1702) & (!g1705)) + ((g290) & (!g319) & (g1701) & (!g1702) & (g1705)) + ((g290) & (!g319) & (g1701) & (g1702) & (!g1705)) + ((g290) & (!g319) & (g1701) & (g1702) & (g1705)) + ((g290) & (g319) & (!g1701) & (!g1702) & (g1705)) + ((g290) & (g319) & (!g1701) & (g1702) & (!g1705)) + ((g290) & (g319) & (!g1701) & (g1702) & (g1705)) + ((g290) & (g319) & (g1701) & (!g1702) & (!g1705)) + ((g290) & (g319) & (g1701) & (!g1702) & (g1705)) + ((g290) & (g319) & (g1701) & (g1702) & (!g1705)) + ((g290) & (g319) & (g1701) & (g1702) & (g1705)));
	assign g1707 = (((!g229) & (!g255) & (g1698) & (g1699) & (g1706)) + ((!g229) & (g255) & (g1698) & (!g1699) & (g1706)) + ((!g229) & (g255) & (g1698) & (g1699) & (!g1706)) + ((!g229) & (g255) & (g1698) & (g1699) & (g1706)) + ((g229) & (!g255) & (!g1698) & (g1699) & (g1706)) + ((g229) & (!g255) & (g1698) & (!g1699) & (!g1706)) + ((g229) & (!g255) & (g1698) & (!g1699) & (g1706)) + ((g229) & (!g255) & (g1698) & (g1699) & (!g1706)) + ((g229) & (!g255) & (g1698) & (g1699) & (g1706)) + ((g229) & (g255) & (!g1698) & (!g1699) & (g1706)) + ((g229) & (g255) & (!g1698) & (g1699) & (!g1706)) + ((g229) & (g255) & (!g1698) & (g1699) & (g1706)) + ((g229) & (g255) & (g1698) & (!g1699) & (!g1706)) + ((g229) & (g255) & (g1698) & (!g1699) & (g1706)) + ((g229) & (g255) & (g1698) & (g1699) & (!g1706)) + ((g229) & (g255) & (g1698) & (g1699) & (g1706)));
	assign g1708 = (((!g174) & (!g198) & (g1695) & (g1696) & (g1707)) + ((!g174) & (g198) & (g1695) & (!g1696) & (g1707)) + ((!g174) & (g198) & (g1695) & (g1696) & (!g1707)) + ((!g174) & (g198) & (g1695) & (g1696) & (g1707)) + ((g174) & (!g198) & (!g1695) & (g1696) & (g1707)) + ((g174) & (!g198) & (g1695) & (!g1696) & (!g1707)) + ((g174) & (!g198) & (g1695) & (!g1696) & (g1707)) + ((g174) & (!g198) & (g1695) & (g1696) & (!g1707)) + ((g174) & (!g198) & (g1695) & (g1696) & (g1707)) + ((g174) & (g198) & (!g1695) & (!g1696) & (g1707)) + ((g174) & (g198) & (!g1695) & (g1696) & (!g1707)) + ((g174) & (g198) & (!g1695) & (g1696) & (g1707)) + ((g174) & (g198) & (g1695) & (!g1696) & (!g1707)) + ((g174) & (g198) & (g1695) & (!g1696) & (g1707)) + ((g174) & (g198) & (g1695) & (g1696) & (!g1707)) + ((g174) & (g198) & (g1695) & (g1696) & (g1707)));
	assign g1709 = (((!g127) & (!g147) & (g1692) & (g1693) & (g1708)) + ((!g127) & (g147) & (g1692) & (!g1693) & (g1708)) + ((!g127) & (g147) & (g1692) & (g1693) & (!g1708)) + ((!g127) & (g147) & (g1692) & (g1693) & (g1708)) + ((g127) & (!g147) & (!g1692) & (g1693) & (g1708)) + ((g127) & (!g147) & (g1692) & (!g1693) & (!g1708)) + ((g127) & (!g147) & (g1692) & (!g1693) & (g1708)) + ((g127) & (!g147) & (g1692) & (g1693) & (!g1708)) + ((g127) & (!g147) & (g1692) & (g1693) & (g1708)) + ((g127) & (g147) & (!g1692) & (!g1693) & (g1708)) + ((g127) & (g147) & (!g1692) & (g1693) & (!g1708)) + ((g127) & (g147) & (!g1692) & (g1693) & (g1708)) + ((g127) & (g147) & (g1692) & (!g1693) & (!g1708)) + ((g127) & (g147) & (g1692) & (!g1693) & (g1708)) + ((g127) & (g147) & (g1692) & (g1693) & (!g1708)) + ((g127) & (g147) & (g1692) & (g1693) & (g1708)));
	assign g1710 = (((!g87) & (!g104) & (g1689) & (g1690) & (g1709)) + ((!g87) & (g104) & (g1689) & (!g1690) & (g1709)) + ((!g87) & (g104) & (g1689) & (g1690) & (!g1709)) + ((!g87) & (g104) & (g1689) & (g1690) & (g1709)) + ((g87) & (!g104) & (!g1689) & (g1690) & (g1709)) + ((g87) & (!g104) & (g1689) & (!g1690) & (!g1709)) + ((g87) & (!g104) & (g1689) & (!g1690) & (g1709)) + ((g87) & (!g104) & (g1689) & (g1690) & (!g1709)) + ((g87) & (!g104) & (g1689) & (g1690) & (g1709)) + ((g87) & (g104) & (!g1689) & (!g1690) & (g1709)) + ((g87) & (g104) & (!g1689) & (g1690) & (!g1709)) + ((g87) & (g104) & (!g1689) & (g1690) & (g1709)) + ((g87) & (g104) & (g1689) & (!g1690) & (!g1709)) + ((g87) & (g104) & (g1689) & (!g1690) & (g1709)) + ((g87) & (g104) & (g1689) & (g1690) & (!g1709)) + ((g87) & (g104) & (g1689) & (g1690) & (g1709)));
	assign g1711 = (((!g54) & (!g68) & (g1686) & (g1687) & (g1710)) + ((!g54) & (g68) & (g1686) & (!g1687) & (g1710)) + ((!g54) & (g68) & (g1686) & (g1687) & (!g1710)) + ((!g54) & (g68) & (g1686) & (g1687) & (g1710)) + ((g54) & (!g68) & (!g1686) & (g1687) & (g1710)) + ((g54) & (!g68) & (g1686) & (!g1687) & (!g1710)) + ((g54) & (!g68) & (g1686) & (!g1687) & (g1710)) + ((g54) & (!g68) & (g1686) & (g1687) & (!g1710)) + ((g54) & (!g68) & (g1686) & (g1687) & (g1710)) + ((g54) & (g68) & (!g1686) & (!g1687) & (g1710)) + ((g54) & (g68) & (!g1686) & (g1687) & (!g1710)) + ((g54) & (g68) & (!g1686) & (g1687) & (g1710)) + ((g54) & (g68) & (g1686) & (!g1687) & (!g1710)) + ((g54) & (g68) & (g1686) & (!g1687) & (g1710)) + ((g54) & (g68) & (g1686) & (g1687) & (!g1710)) + ((g54) & (g68) & (g1686) & (g1687) & (g1710)));
	assign g1712 = (((!g27) & (!g39) & (g1683) & (g1684) & (g1711)) + ((!g27) & (g39) & (g1683) & (!g1684) & (g1711)) + ((!g27) & (g39) & (g1683) & (g1684) & (!g1711)) + ((!g27) & (g39) & (g1683) & (g1684) & (g1711)) + ((g27) & (!g39) & (!g1683) & (g1684) & (g1711)) + ((g27) & (!g39) & (g1683) & (!g1684) & (!g1711)) + ((g27) & (!g39) & (g1683) & (!g1684) & (g1711)) + ((g27) & (!g39) & (g1683) & (g1684) & (!g1711)) + ((g27) & (!g39) & (g1683) & (g1684) & (g1711)) + ((g27) & (g39) & (!g1683) & (!g1684) & (g1711)) + ((g27) & (g39) & (!g1683) & (g1684) & (!g1711)) + ((g27) & (g39) & (!g1683) & (g1684) & (g1711)) + ((g27) & (g39) & (g1683) & (!g1684) & (!g1711)) + ((g27) & (g39) & (g1683) & (!g1684) & (g1711)) + ((g27) & (g39) & (g1683) & (g1684) & (!g1711)) + ((g27) & (g39) & (g1683) & (g1684) & (g1711)));
	assign g1713 = (((!g8) & (!g18) & (g1680) & (g1681) & (g1712)) + ((!g8) & (g18) & (g1680) & (!g1681) & (g1712)) + ((!g8) & (g18) & (g1680) & (g1681) & (!g1712)) + ((!g8) & (g18) & (g1680) & (g1681) & (g1712)) + ((g8) & (!g18) & (!g1680) & (g1681) & (g1712)) + ((g8) & (!g18) & (g1680) & (!g1681) & (!g1712)) + ((g8) & (!g18) & (g1680) & (!g1681) & (g1712)) + ((g8) & (!g18) & (g1680) & (g1681) & (!g1712)) + ((g8) & (!g18) & (g1680) & (g1681) & (g1712)) + ((g8) & (g18) & (!g1680) & (!g1681) & (g1712)) + ((g8) & (g18) & (!g1680) & (g1681) & (!g1712)) + ((g8) & (g18) & (!g1680) & (g1681) & (g1712)) + ((g8) & (g18) & (g1680) & (!g1681) & (!g1712)) + ((g8) & (g18) & (g1680) & (!g1681) & (g1712)) + ((g8) & (g18) & (g1680) & (g1681) & (!g1712)) + ((g8) & (g18) & (g1680) & (g1681) & (g1712)));
	assign g1714 = (((!g2) & (!g8) & (g1603) & (g1629)) + ((!g2) & (g8) & (!g1603) & (g1629)) + ((!g2) & (g8) & (g1603) & (!g1629)) + ((!g2) & (g8) & (g1603) & (g1629)) + ((g2) & (!g8) & (!g1603) & (!g1629)) + ((g2) & (!g8) & (!g1603) & (g1629)) + ((g2) & (!g8) & (g1603) & (!g1629)) + ((g2) & (g8) & (!g1603) & (!g1629)));
	assign g1715 = (((!g1602) & (!g1600) & (!g1633) & (g1714)) + ((!g1602) & (g1600) & (!g1633) & (g1714)) + ((!g1602) & (g1600) & (g1633) & (g1714)) + ((g1602) & (!g1600) & (!g1633) & (!g1714)) + ((g1602) & (!g1600) & (g1633) & (!g1714)) + ((g1602) & (!g1600) & (g1633) & (g1714)) + ((g1602) & (g1600) & (!g1633) & (!g1714)) + ((g1602) & (g1600) & (g1633) & (!g1714)));
	assign g1716 = (((!g4) & (!g2) & (!g1678) & (!g1713) & (g1715)) + ((!g4) & (!g2) & (!g1678) & (g1713) & (g1715)) + ((!g4) & (!g2) & (g1678) & (!g1713) & (g1715)) + ((!g4) & (!g2) & (g1678) & (g1713) & (!g1715)) + ((!g4) & (!g2) & (g1678) & (g1713) & (g1715)) + ((!g4) & (g2) & (!g1678) & (!g1713) & (g1715)) + ((!g4) & (g2) & (!g1678) & (g1713) & (!g1715)) + ((!g4) & (g2) & (!g1678) & (g1713) & (g1715)) + ((!g4) & (g2) & (g1678) & (!g1713) & (!g1715)) + ((!g4) & (g2) & (g1678) & (!g1713) & (g1715)) + ((!g4) & (g2) & (g1678) & (g1713) & (!g1715)) + ((!g4) & (g2) & (g1678) & (g1713) & (g1715)) + ((g4) & (!g2) & (g1678) & (g1713) & (g1715)) + ((g4) & (g2) & (!g1678) & (g1713) & (g1715)) + ((g4) & (g2) & (g1678) & (!g1713) & (g1715)) + ((g4) & (g2) & (g1678) & (g1713) & (g1715)));
	assign g1717 = (((!g4) & (!g1630) & (g1631)) + ((!g4) & (g1630) & (!g1631)) + ((!g4) & (g1630) & (g1631)) + ((g4) & (g1630) & (g1631)));
	assign g1718 = (((!g1601) & (!g1717) & (!g1600) & (!g1633)) + ((!g1601) & (!g1717) & (g1600) & (!g1633)) + ((!g1601) & (!g1717) & (g1600) & (g1633)) + ((g1601) & (g1717) & (!g1600) & (!g1633)) + ((g1601) & (g1717) & (!g1600) & (g1633)) + ((g1601) & (g1717) & (g1600) & (!g1633)) + ((g1601) & (g1717) & (g1600) & (g1633)));
	assign g1719 = (((!g1) & (g1601) & (!g1717) & (!g1600) & (g1633)) + ((!g1) & (g1601) & (g1717) & (!g1600) & (g1633)) + ((g1) & (!g1601) & (g1717) & (g1600) & (!g1633)) + ((g1) & (!g1601) & (g1717) & (g1600) & (g1633)) + ((g1) & (g1601) & (!g1717) & (!g1600) & (!g1633)) + ((g1) & (g1601) & (!g1717) & (!g1600) & (g1633)) + ((g1) & (g1601) & (!g1717) & (g1600) & (!g1633)) + ((g1) & (g1601) & (!g1717) & (g1600) & (g1633)) + ((g1) & (g1601) & (g1717) & (!g1600) & (g1633)));
	assign g1720 = (((!g1) & (!g1677) & (!g1716) & (!g1718) & (!g1719)) + ((g1) & (!g1677) & (!g1716) & (!g1718) & (!g1719)) + ((g1) & (!g1677) & (!g1716) & (g1718) & (!g1719)) + ((g1) & (!g1677) & (g1716) & (!g1718) & (!g1719)) + ((g1) & (!g1677) & (g1716) & (g1718) & (!g1719)) + ((g1) & (g1677) & (!g1716) & (!g1718) & (!g1719)) + ((g1) & (g1677) & (!g1716) & (g1718) & (!g1719)));
	assign g1721 = (((!g390) & (!g1634) & (g1676) & (!g1720)) + ((!g390) & (g1634) & (!g1676) & (!g1720)) + ((!g390) & (g1634) & (!g1676) & (g1720)) + ((!g390) & (g1634) & (g1676) & (g1720)) + ((g390) & (!g1634) & (!g1676) & (!g1720)) + ((g390) & (g1634) & (!g1676) & (g1720)) + ((g390) & (g1634) & (g1676) & (!g1720)) + ((g390) & (g1634) & (g1676) & (g1720)));
	assign g1722 = (((!g433) & (!g468) & (!g1636) & (g1637) & (g1675) & (!g1720)) + ((!g433) & (!g468) & (g1636) & (!g1637) & (!g1675) & (!g1720)) + ((!g433) & (!g468) & (g1636) & (!g1637) & (!g1675) & (g1720)) + ((!g433) & (!g468) & (g1636) & (!g1637) & (g1675) & (!g1720)) + ((!g433) & (!g468) & (g1636) & (!g1637) & (g1675) & (g1720)) + ((!g433) & (!g468) & (g1636) & (g1637) & (!g1675) & (!g1720)) + ((!g433) & (!g468) & (g1636) & (g1637) & (!g1675) & (g1720)) + ((!g433) & (!g468) & (g1636) & (g1637) & (g1675) & (g1720)) + ((!g433) & (g468) & (!g1636) & (!g1637) & (g1675) & (!g1720)) + ((!g433) & (g468) & (!g1636) & (g1637) & (!g1675) & (!g1720)) + ((!g433) & (g468) & (!g1636) & (g1637) & (g1675) & (!g1720)) + ((!g433) & (g468) & (g1636) & (!g1637) & (!g1675) & (!g1720)) + ((!g433) & (g468) & (g1636) & (!g1637) & (!g1675) & (g1720)) + ((!g433) & (g468) & (g1636) & (!g1637) & (g1675) & (g1720)) + ((!g433) & (g468) & (g1636) & (g1637) & (!g1675) & (g1720)) + ((!g433) & (g468) & (g1636) & (g1637) & (g1675) & (g1720)) + ((g433) & (!g468) & (!g1636) & (!g1637) & (!g1675) & (!g1720)) + ((g433) & (!g468) & (!g1636) & (!g1637) & (g1675) & (!g1720)) + ((g433) & (!g468) & (!g1636) & (g1637) & (!g1675) & (!g1720)) + ((g433) & (!g468) & (g1636) & (!g1637) & (!g1675) & (g1720)) + ((g433) & (!g468) & (g1636) & (!g1637) & (g1675) & (g1720)) + ((g433) & (!g468) & (g1636) & (g1637) & (!g1675) & (g1720)) + ((g433) & (!g468) & (g1636) & (g1637) & (g1675) & (!g1720)) + ((g433) & (!g468) & (g1636) & (g1637) & (g1675) & (g1720)) + ((g433) & (g468) & (!g1636) & (!g1637) & (!g1675) & (!g1720)) + ((g433) & (g468) & (g1636) & (!g1637) & (!g1675) & (g1720)) + ((g433) & (g468) & (g1636) & (!g1637) & (g1675) & (!g1720)) + ((g433) & (g468) & (g1636) & (!g1637) & (g1675) & (g1720)) + ((g433) & (g468) & (g1636) & (g1637) & (!g1675) & (!g1720)) + ((g433) & (g468) & (g1636) & (g1637) & (!g1675) & (g1720)) + ((g433) & (g468) & (g1636) & (g1637) & (g1675) & (!g1720)) + ((g433) & (g468) & (g1636) & (g1637) & (g1675) & (g1720)));
	assign g1723 = (((!g468) & (!g1637) & (g1675) & (!g1720)) + ((!g468) & (g1637) & (!g1675) & (!g1720)) + ((!g468) & (g1637) & (!g1675) & (g1720)) + ((!g468) & (g1637) & (g1675) & (g1720)) + ((g468) & (!g1637) & (!g1675) & (!g1720)) + ((g468) & (g1637) & (!g1675) & (g1720)) + ((g468) & (g1637) & (g1675) & (!g1720)) + ((g468) & (g1637) & (g1675) & (g1720)));
	assign g1724 = (((!g515) & (!g553) & (!g1639) & (g1640) & (g1674) & (!g1720)) + ((!g515) & (!g553) & (g1639) & (!g1640) & (!g1674) & (!g1720)) + ((!g515) & (!g553) & (g1639) & (!g1640) & (!g1674) & (g1720)) + ((!g515) & (!g553) & (g1639) & (!g1640) & (g1674) & (!g1720)) + ((!g515) & (!g553) & (g1639) & (!g1640) & (g1674) & (g1720)) + ((!g515) & (!g553) & (g1639) & (g1640) & (!g1674) & (!g1720)) + ((!g515) & (!g553) & (g1639) & (g1640) & (!g1674) & (g1720)) + ((!g515) & (!g553) & (g1639) & (g1640) & (g1674) & (g1720)) + ((!g515) & (g553) & (!g1639) & (!g1640) & (g1674) & (!g1720)) + ((!g515) & (g553) & (!g1639) & (g1640) & (!g1674) & (!g1720)) + ((!g515) & (g553) & (!g1639) & (g1640) & (g1674) & (!g1720)) + ((!g515) & (g553) & (g1639) & (!g1640) & (!g1674) & (!g1720)) + ((!g515) & (g553) & (g1639) & (!g1640) & (!g1674) & (g1720)) + ((!g515) & (g553) & (g1639) & (!g1640) & (g1674) & (g1720)) + ((!g515) & (g553) & (g1639) & (g1640) & (!g1674) & (g1720)) + ((!g515) & (g553) & (g1639) & (g1640) & (g1674) & (g1720)) + ((g515) & (!g553) & (!g1639) & (!g1640) & (!g1674) & (!g1720)) + ((g515) & (!g553) & (!g1639) & (!g1640) & (g1674) & (!g1720)) + ((g515) & (!g553) & (!g1639) & (g1640) & (!g1674) & (!g1720)) + ((g515) & (!g553) & (g1639) & (!g1640) & (!g1674) & (g1720)) + ((g515) & (!g553) & (g1639) & (!g1640) & (g1674) & (g1720)) + ((g515) & (!g553) & (g1639) & (g1640) & (!g1674) & (g1720)) + ((g515) & (!g553) & (g1639) & (g1640) & (g1674) & (!g1720)) + ((g515) & (!g553) & (g1639) & (g1640) & (g1674) & (g1720)) + ((g515) & (g553) & (!g1639) & (!g1640) & (!g1674) & (!g1720)) + ((g515) & (g553) & (g1639) & (!g1640) & (!g1674) & (g1720)) + ((g515) & (g553) & (g1639) & (!g1640) & (g1674) & (!g1720)) + ((g515) & (g553) & (g1639) & (!g1640) & (g1674) & (g1720)) + ((g515) & (g553) & (g1639) & (g1640) & (!g1674) & (!g1720)) + ((g515) & (g553) & (g1639) & (g1640) & (!g1674) & (g1720)) + ((g515) & (g553) & (g1639) & (g1640) & (g1674) & (!g1720)) + ((g515) & (g553) & (g1639) & (g1640) & (g1674) & (g1720)));
	assign g1725 = (((!g553) & (!g1640) & (g1674) & (!g1720)) + ((!g553) & (g1640) & (!g1674) & (!g1720)) + ((!g553) & (g1640) & (!g1674) & (g1720)) + ((!g553) & (g1640) & (g1674) & (g1720)) + ((g553) & (!g1640) & (!g1674) & (!g1720)) + ((g553) & (g1640) & (!g1674) & (g1720)) + ((g553) & (g1640) & (g1674) & (!g1720)) + ((g553) & (g1640) & (g1674) & (g1720)));
	assign g1726 = (((!g604) & (!g645) & (!g1642) & (g1643) & (g1673) & (!g1720)) + ((!g604) & (!g645) & (g1642) & (!g1643) & (!g1673) & (!g1720)) + ((!g604) & (!g645) & (g1642) & (!g1643) & (!g1673) & (g1720)) + ((!g604) & (!g645) & (g1642) & (!g1643) & (g1673) & (!g1720)) + ((!g604) & (!g645) & (g1642) & (!g1643) & (g1673) & (g1720)) + ((!g604) & (!g645) & (g1642) & (g1643) & (!g1673) & (!g1720)) + ((!g604) & (!g645) & (g1642) & (g1643) & (!g1673) & (g1720)) + ((!g604) & (!g645) & (g1642) & (g1643) & (g1673) & (g1720)) + ((!g604) & (g645) & (!g1642) & (!g1643) & (g1673) & (!g1720)) + ((!g604) & (g645) & (!g1642) & (g1643) & (!g1673) & (!g1720)) + ((!g604) & (g645) & (!g1642) & (g1643) & (g1673) & (!g1720)) + ((!g604) & (g645) & (g1642) & (!g1643) & (!g1673) & (!g1720)) + ((!g604) & (g645) & (g1642) & (!g1643) & (!g1673) & (g1720)) + ((!g604) & (g645) & (g1642) & (!g1643) & (g1673) & (g1720)) + ((!g604) & (g645) & (g1642) & (g1643) & (!g1673) & (g1720)) + ((!g604) & (g645) & (g1642) & (g1643) & (g1673) & (g1720)) + ((g604) & (!g645) & (!g1642) & (!g1643) & (!g1673) & (!g1720)) + ((g604) & (!g645) & (!g1642) & (!g1643) & (g1673) & (!g1720)) + ((g604) & (!g645) & (!g1642) & (g1643) & (!g1673) & (!g1720)) + ((g604) & (!g645) & (g1642) & (!g1643) & (!g1673) & (g1720)) + ((g604) & (!g645) & (g1642) & (!g1643) & (g1673) & (g1720)) + ((g604) & (!g645) & (g1642) & (g1643) & (!g1673) & (g1720)) + ((g604) & (!g645) & (g1642) & (g1643) & (g1673) & (!g1720)) + ((g604) & (!g645) & (g1642) & (g1643) & (g1673) & (g1720)) + ((g604) & (g645) & (!g1642) & (!g1643) & (!g1673) & (!g1720)) + ((g604) & (g645) & (g1642) & (!g1643) & (!g1673) & (g1720)) + ((g604) & (g645) & (g1642) & (!g1643) & (g1673) & (!g1720)) + ((g604) & (g645) & (g1642) & (!g1643) & (g1673) & (g1720)) + ((g604) & (g645) & (g1642) & (g1643) & (!g1673) & (!g1720)) + ((g604) & (g645) & (g1642) & (g1643) & (!g1673) & (g1720)) + ((g604) & (g645) & (g1642) & (g1643) & (g1673) & (!g1720)) + ((g604) & (g645) & (g1642) & (g1643) & (g1673) & (g1720)));
	assign g1727 = (((!g645) & (!g1643) & (g1673) & (!g1720)) + ((!g645) & (g1643) & (!g1673) & (!g1720)) + ((!g645) & (g1643) & (!g1673) & (g1720)) + ((!g645) & (g1643) & (g1673) & (g1720)) + ((g645) & (!g1643) & (!g1673) & (!g1720)) + ((g645) & (g1643) & (!g1673) & (g1720)) + ((g645) & (g1643) & (g1673) & (!g1720)) + ((g645) & (g1643) & (g1673) & (g1720)));
	assign g1728 = (((!g700) & (!g744) & (!g1645) & (g1646) & (g1672) & (!g1720)) + ((!g700) & (!g744) & (g1645) & (!g1646) & (!g1672) & (!g1720)) + ((!g700) & (!g744) & (g1645) & (!g1646) & (!g1672) & (g1720)) + ((!g700) & (!g744) & (g1645) & (!g1646) & (g1672) & (!g1720)) + ((!g700) & (!g744) & (g1645) & (!g1646) & (g1672) & (g1720)) + ((!g700) & (!g744) & (g1645) & (g1646) & (!g1672) & (!g1720)) + ((!g700) & (!g744) & (g1645) & (g1646) & (!g1672) & (g1720)) + ((!g700) & (!g744) & (g1645) & (g1646) & (g1672) & (g1720)) + ((!g700) & (g744) & (!g1645) & (!g1646) & (g1672) & (!g1720)) + ((!g700) & (g744) & (!g1645) & (g1646) & (!g1672) & (!g1720)) + ((!g700) & (g744) & (!g1645) & (g1646) & (g1672) & (!g1720)) + ((!g700) & (g744) & (g1645) & (!g1646) & (!g1672) & (!g1720)) + ((!g700) & (g744) & (g1645) & (!g1646) & (!g1672) & (g1720)) + ((!g700) & (g744) & (g1645) & (!g1646) & (g1672) & (g1720)) + ((!g700) & (g744) & (g1645) & (g1646) & (!g1672) & (g1720)) + ((!g700) & (g744) & (g1645) & (g1646) & (g1672) & (g1720)) + ((g700) & (!g744) & (!g1645) & (!g1646) & (!g1672) & (!g1720)) + ((g700) & (!g744) & (!g1645) & (!g1646) & (g1672) & (!g1720)) + ((g700) & (!g744) & (!g1645) & (g1646) & (!g1672) & (!g1720)) + ((g700) & (!g744) & (g1645) & (!g1646) & (!g1672) & (g1720)) + ((g700) & (!g744) & (g1645) & (!g1646) & (g1672) & (g1720)) + ((g700) & (!g744) & (g1645) & (g1646) & (!g1672) & (g1720)) + ((g700) & (!g744) & (g1645) & (g1646) & (g1672) & (!g1720)) + ((g700) & (!g744) & (g1645) & (g1646) & (g1672) & (g1720)) + ((g700) & (g744) & (!g1645) & (!g1646) & (!g1672) & (!g1720)) + ((g700) & (g744) & (g1645) & (!g1646) & (!g1672) & (g1720)) + ((g700) & (g744) & (g1645) & (!g1646) & (g1672) & (!g1720)) + ((g700) & (g744) & (g1645) & (!g1646) & (g1672) & (g1720)) + ((g700) & (g744) & (g1645) & (g1646) & (!g1672) & (!g1720)) + ((g700) & (g744) & (g1645) & (g1646) & (!g1672) & (g1720)) + ((g700) & (g744) & (g1645) & (g1646) & (g1672) & (!g1720)) + ((g700) & (g744) & (g1645) & (g1646) & (g1672) & (g1720)));
	assign g1729 = (((!g744) & (!g1646) & (g1672) & (!g1720)) + ((!g744) & (g1646) & (!g1672) & (!g1720)) + ((!g744) & (g1646) & (!g1672) & (g1720)) + ((!g744) & (g1646) & (g1672) & (g1720)) + ((g744) & (!g1646) & (!g1672) & (!g1720)) + ((g744) & (g1646) & (!g1672) & (g1720)) + ((g744) & (g1646) & (g1672) & (!g1720)) + ((g744) & (g1646) & (g1672) & (g1720)));
	assign g1730 = (((!g803) & (!g851) & (!g1648) & (g1649) & (g1671) & (!g1720)) + ((!g803) & (!g851) & (g1648) & (!g1649) & (!g1671) & (!g1720)) + ((!g803) & (!g851) & (g1648) & (!g1649) & (!g1671) & (g1720)) + ((!g803) & (!g851) & (g1648) & (!g1649) & (g1671) & (!g1720)) + ((!g803) & (!g851) & (g1648) & (!g1649) & (g1671) & (g1720)) + ((!g803) & (!g851) & (g1648) & (g1649) & (!g1671) & (!g1720)) + ((!g803) & (!g851) & (g1648) & (g1649) & (!g1671) & (g1720)) + ((!g803) & (!g851) & (g1648) & (g1649) & (g1671) & (g1720)) + ((!g803) & (g851) & (!g1648) & (!g1649) & (g1671) & (!g1720)) + ((!g803) & (g851) & (!g1648) & (g1649) & (!g1671) & (!g1720)) + ((!g803) & (g851) & (!g1648) & (g1649) & (g1671) & (!g1720)) + ((!g803) & (g851) & (g1648) & (!g1649) & (!g1671) & (!g1720)) + ((!g803) & (g851) & (g1648) & (!g1649) & (!g1671) & (g1720)) + ((!g803) & (g851) & (g1648) & (!g1649) & (g1671) & (g1720)) + ((!g803) & (g851) & (g1648) & (g1649) & (!g1671) & (g1720)) + ((!g803) & (g851) & (g1648) & (g1649) & (g1671) & (g1720)) + ((g803) & (!g851) & (!g1648) & (!g1649) & (!g1671) & (!g1720)) + ((g803) & (!g851) & (!g1648) & (!g1649) & (g1671) & (!g1720)) + ((g803) & (!g851) & (!g1648) & (g1649) & (!g1671) & (!g1720)) + ((g803) & (!g851) & (g1648) & (!g1649) & (!g1671) & (g1720)) + ((g803) & (!g851) & (g1648) & (!g1649) & (g1671) & (g1720)) + ((g803) & (!g851) & (g1648) & (g1649) & (!g1671) & (g1720)) + ((g803) & (!g851) & (g1648) & (g1649) & (g1671) & (!g1720)) + ((g803) & (!g851) & (g1648) & (g1649) & (g1671) & (g1720)) + ((g803) & (g851) & (!g1648) & (!g1649) & (!g1671) & (!g1720)) + ((g803) & (g851) & (g1648) & (!g1649) & (!g1671) & (g1720)) + ((g803) & (g851) & (g1648) & (!g1649) & (g1671) & (!g1720)) + ((g803) & (g851) & (g1648) & (!g1649) & (g1671) & (g1720)) + ((g803) & (g851) & (g1648) & (g1649) & (!g1671) & (!g1720)) + ((g803) & (g851) & (g1648) & (g1649) & (!g1671) & (g1720)) + ((g803) & (g851) & (g1648) & (g1649) & (g1671) & (!g1720)) + ((g803) & (g851) & (g1648) & (g1649) & (g1671) & (g1720)));
	assign g1731 = (((!g851) & (!g1649) & (g1671) & (!g1720)) + ((!g851) & (g1649) & (!g1671) & (!g1720)) + ((!g851) & (g1649) & (!g1671) & (g1720)) + ((!g851) & (g1649) & (g1671) & (g1720)) + ((g851) & (!g1649) & (!g1671) & (!g1720)) + ((g851) & (g1649) & (!g1671) & (g1720)) + ((g851) & (g1649) & (g1671) & (!g1720)) + ((g851) & (g1649) & (g1671) & (g1720)));
	assign g1732 = (((!g914) & (!g1032) & (!g1651) & (g1652) & (g1670) & (!g1720)) + ((!g914) & (!g1032) & (g1651) & (!g1652) & (!g1670) & (!g1720)) + ((!g914) & (!g1032) & (g1651) & (!g1652) & (!g1670) & (g1720)) + ((!g914) & (!g1032) & (g1651) & (!g1652) & (g1670) & (!g1720)) + ((!g914) & (!g1032) & (g1651) & (!g1652) & (g1670) & (g1720)) + ((!g914) & (!g1032) & (g1651) & (g1652) & (!g1670) & (!g1720)) + ((!g914) & (!g1032) & (g1651) & (g1652) & (!g1670) & (g1720)) + ((!g914) & (!g1032) & (g1651) & (g1652) & (g1670) & (g1720)) + ((!g914) & (g1032) & (!g1651) & (!g1652) & (g1670) & (!g1720)) + ((!g914) & (g1032) & (!g1651) & (g1652) & (!g1670) & (!g1720)) + ((!g914) & (g1032) & (!g1651) & (g1652) & (g1670) & (!g1720)) + ((!g914) & (g1032) & (g1651) & (!g1652) & (!g1670) & (!g1720)) + ((!g914) & (g1032) & (g1651) & (!g1652) & (!g1670) & (g1720)) + ((!g914) & (g1032) & (g1651) & (!g1652) & (g1670) & (g1720)) + ((!g914) & (g1032) & (g1651) & (g1652) & (!g1670) & (g1720)) + ((!g914) & (g1032) & (g1651) & (g1652) & (g1670) & (g1720)) + ((g914) & (!g1032) & (!g1651) & (!g1652) & (!g1670) & (!g1720)) + ((g914) & (!g1032) & (!g1651) & (!g1652) & (g1670) & (!g1720)) + ((g914) & (!g1032) & (!g1651) & (g1652) & (!g1670) & (!g1720)) + ((g914) & (!g1032) & (g1651) & (!g1652) & (!g1670) & (g1720)) + ((g914) & (!g1032) & (g1651) & (!g1652) & (g1670) & (g1720)) + ((g914) & (!g1032) & (g1651) & (g1652) & (!g1670) & (g1720)) + ((g914) & (!g1032) & (g1651) & (g1652) & (g1670) & (!g1720)) + ((g914) & (!g1032) & (g1651) & (g1652) & (g1670) & (g1720)) + ((g914) & (g1032) & (!g1651) & (!g1652) & (!g1670) & (!g1720)) + ((g914) & (g1032) & (g1651) & (!g1652) & (!g1670) & (g1720)) + ((g914) & (g1032) & (g1651) & (!g1652) & (g1670) & (!g1720)) + ((g914) & (g1032) & (g1651) & (!g1652) & (g1670) & (g1720)) + ((g914) & (g1032) & (g1651) & (g1652) & (!g1670) & (!g1720)) + ((g914) & (g1032) & (g1651) & (g1652) & (!g1670) & (g1720)) + ((g914) & (g1032) & (g1651) & (g1652) & (g1670) & (!g1720)) + ((g914) & (g1032) & (g1651) & (g1652) & (g1670) & (g1720)));
	assign g1733 = (((!g1032) & (!g1652) & (g1670) & (!g1720)) + ((!g1032) & (g1652) & (!g1670) & (!g1720)) + ((!g1032) & (g1652) & (!g1670) & (g1720)) + ((!g1032) & (g1652) & (g1670) & (g1720)) + ((g1032) & (!g1652) & (!g1670) & (!g1720)) + ((g1032) & (g1652) & (!g1670) & (g1720)) + ((g1032) & (g1652) & (g1670) & (!g1720)) + ((g1032) & (g1652) & (g1670) & (g1720)));
	assign g1734 = (((!g1030) & (!g1160) & (!g1654) & (g1655) & (g1669) & (!g1720)) + ((!g1030) & (!g1160) & (g1654) & (!g1655) & (!g1669) & (!g1720)) + ((!g1030) & (!g1160) & (g1654) & (!g1655) & (!g1669) & (g1720)) + ((!g1030) & (!g1160) & (g1654) & (!g1655) & (g1669) & (!g1720)) + ((!g1030) & (!g1160) & (g1654) & (!g1655) & (g1669) & (g1720)) + ((!g1030) & (!g1160) & (g1654) & (g1655) & (!g1669) & (!g1720)) + ((!g1030) & (!g1160) & (g1654) & (g1655) & (!g1669) & (g1720)) + ((!g1030) & (!g1160) & (g1654) & (g1655) & (g1669) & (g1720)) + ((!g1030) & (g1160) & (!g1654) & (!g1655) & (g1669) & (!g1720)) + ((!g1030) & (g1160) & (!g1654) & (g1655) & (!g1669) & (!g1720)) + ((!g1030) & (g1160) & (!g1654) & (g1655) & (g1669) & (!g1720)) + ((!g1030) & (g1160) & (g1654) & (!g1655) & (!g1669) & (!g1720)) + ((!g1030) & (g1160) & (g1654) & (!g1655) & (!g1669) & (g1720)) + ((!g1030) & (g1160) & (g1654) & (!g1655) & (g1669) & (g1720)) + ((!g1030) & (g1160) & (g1654) & (g1655) & (!g1669) & (g1720)) + ((!g1030) & (g1160) & (g1654) & (g1655) & (g1669) & (g1720)) + ((g1030) & (!g1160) & (!g1654) & (!g1655) & (!g1669) & (!g1720)) + ((g1030) & (!g1160) & (!g1654) & (!g1655) & (g1669) & (!g1720)) + ((g1030) & (!g1160) & (!g1654) & (g1655) & (!g1669) & (!g1720)) + ((g1030) & (!g1160) & (g1654) & (!g1655) & (!g1669) & (g1720)) + ((g1030) & (!g1160) & (g1654) & (!g1655) & (g1669) & (g1720)) + ((g1030) & (!g1160) & (g1654) & (g1655) & (!g1669) & (g1720)) + ((g1030) & (!g1160) & (g1654) & (g1655) & (g1669) & (!g1720)) + ((g1030) & (!g1160) & (g1654) & (g1655) & (g1669) & (g1720)) + ((g1030) & (g1160) & (!g1654) & (!g1655) & (!g1669) & (!g1720)) + ((g1030) & (g1160) & (g1654) & (!g1655) & (!g1669) & (g1720)) + ((g1030) & (g1160) & (g1654) & (!g1655) & (g1669) & (!g1720)) + ((g1030) & (g1160) & (g1654) & (!g1655) & (g1669) & (g1720)) + ((g1030) & (g1160) & (g1654) & (g1655) & (!g1669) & (!g1720)) + ((g1030) & (g1160) & (g1654) & (g1655) & (!g1669) & (g1720)) + ((g1030) & (g1160) & (g1654) & (g1655) & (g1669) & (!g1720)) + ((g1030) & (g1160) & (g1654) & (g1655) & (g1669) & (g1720)));
	assign g1735 = (((!g1160) & (!g1655) & (g1669) & (!g1720)) + ((!g1160) & (g1655) & (!g1669) & (!g1720)) + ((!g1160) & (g1655) & (!g1669) & (g1720)) + ((!g1160) & (g1655) & (g1669) & (g1720)) + ((g1160) & (!g1655) & (!g1669) & (!g1720)) + ((g1160) & (g1655) & (!g1669) & (g1720)) + ((g1160) & (g1655) & (g1669) & (!g1720)) + ((g1160) & (g1655) & (g1669) & (g1720)));
	assign g1736 = (((!g1154) & (!g1295) & (!g1657) & (g1658) & (g1668) & (!g1720)) + ((!g1154) & (!g1295) & (g1657) & (!g1658) & (!g1668) & (!g1720)) + ((!g1154) & (!g1295) & (g1657) & (!g1658) & (!g1668) & (g1720)) + ((!g1154) & (!g1295) & (g1657) & (!g1658) & (g1668) & (!g1720)) + ((!g1154) & (!g1295) & (g1657) & (!g1658) & (g1668) & (g1720)) + ((!g1154) & (!g1295) & (g1657) & (g1658) & (!g1668) & (!g1720)) + ((!g1154) & (!g1295) & (g1657) & (g1658) & (!g1668) & (g1720)) + ((!g1154) & (!g1295) & (g1657) & (g1658) & (g1668) & (g1720)) + ((!g1154) & (g1295) & (!g1657) & (!g1658) & (g1668) & (!g1720)) + ((!g1154) & (g1295) & (!g1657) & (g1658) & (!g1668) & (!g1720)) + ((!g1154) & (g1295) & (!g1657) & (g1658) & (g1668) & (!g1720)) + ((!g1154) & (g1295) & (g1657) & (!g1658) & (!g1668) & (!g1720)) + ((!g1154) & (g1295) & (g1657) & (!g1658) & (!g1668) & (g1720)) + ((!g1154) & (g1295) & (g1657) & (!g1658) & (g1668) & (g1720)) + ((!g1154) & (g1295) & (g1657) & (g1658) & (!g1668) & (g1720)) + ((!g1154) & (g1295) & (g1657) & (g1658) & (g1668) & (g1720)) + ((g1154) & (!g1295) & (!g1657) & (!g1658) & (!g1668) & (!g1720)) + ((g1154) & (!g1295) & (!g1657) & (!g1658) & (g1668) & (!g1720)) + ((g1154) & (!g1295) & (!g1657) & (g1658) & (!g1668) & (!g1720)) + ((g1154) & (!g1295) & (g1657) & (!g1658) & (!g1668) & (g1720)) + ((g1154) & (!g1295) & (g1657) & (!g1658) & (g1668) & (g1720)) + ((g1154) & (!g1295) & (g1657) & (g1658) & (!g1668) & (g1720)) + ((g1154) & (!g1295) & (g1657) & (g1658) & (g1668) & (!g1720)) + ((g1154) & (!g1295) & (g1657) & (g1658) & (g1668) & (g1720)) + ((g1154) & (g1295) & (!g1657) & (!g1658) & (!g1668) & (!g1720)) + ((g1154) & (g1295) & (g1657) & (!g1658) & (!g1668) & (g1720)) + ((g1154) & (g1295) & (g1657) & (!g1658) & (g1668) & (!g1720)) + ((g1154) & (g1295) & (g1657) & (!g1658) & (g1668) & (g1720)) + ((g1154) & (g1295) & (g1657) & (g1658) & (!g1668) & (!g1720)) + ((g1154) & (g1295) & (g1657) & (g1658) & (!g1668) & (g1720)) + ((g1154) & (g1295) & (g1657) & (g1658) & (g1668) & (!g1720)) + ((g1154) & (g1295) & (g1657) & (g1658) & (g1668) & (g1720)));
	assign g1737 = (((!g1295) & (!g1658) & (g1668) & (!g1720)) + ((!g1295) & (g1658) & (!g1668) & (!g1720)) + ((!g1295) & (g1658) & (!g1668) & (g1720)) + ((!g1295) & (g1658) & (g1668) & (g1720)) + ((g1295) & (!g1658) & (!g1668) & (!g1720)) + ((g1295) & (g1658) & (!g1668) & (g1720)) + ((g1295) & (g1658) & (g1668) & (!g1720)) + ((g1295) & (g1658) & (g1668) & (g1720)));
	assign g1738 = (((!g1285) & (!g1437) & (!g1660) & (g1661) & (g1667) & (!g1720)) + ((!g1285) & (!g1437) & (g1660) & (!g1661) & (!g1667) & (!g1720)) + ((!g1285) & (!g1437) & (g1660) & (!g1661) & (!g1667) & (g1720)) + ((!g1285) & (!g1437) & (g1660) & (!g1661) & (g1667) & (!g1720)) + ((!g1285) & (!g1437) & (g1660) & (!g1661) & (g1667) & (g1720)) + ((!g1285) & (!g1437) & (g1660) & (g1661) & (!g1667) & (!g1720)) + ((!g1285) & (!g1437) & (g1660) & (g1661) & (!g1667) & (g1720)) + ((!g1285) & (!g1437) & (g1660) & (g1661) & (g1667) & (g1720)) + ((!g1285) & (g1437) & (!g1660) & (!g1661) & (g1667) & (!g1720)) + ((!g1285) & (g1437) & (!g1660) & (g1661) & (!g1667) & (!g1720)) + ((!g1285) & (g1437) & (!g1660) & (g1661) & (g1667) & (!g1720)) + ((!g1285) & (g1437) & (g1660) & (!g1661) & (!g1667) & (!g1720)) + ((!g1285) & (g1437) & (g1660) & (!g1661) & (!g1667) & (g1720)) + ((!g1285) & (g1437) & (g1660) & (!g1661) & (g1667) & (g1720)) + ((!g1285) & (g1437) & (g1660) & (g1661) & (!g1667) & (g1720)) + ((!g1285) & (g1437) & (g1660) & (g1661) & (g1667) & (g1720)) + ((g1285) & (!g1437) & (!g1660) & (!g1661) & (!g1667) & (!g1720)) + ((g1285) & (!g1437) & (!g1660) & (!g1661) & (g1667) & (!g1720)) + ((g1285) & (!g1437) & (!g1660) & (g1661) & (!g1667) & (!g1720)) + ((g1285) & (!g1437) & (g1660) & (!g1661) & (!g1667) & (g1720)) + ((g1285) & (!g1437) & (g1660) & (!g1661) & (g1667) & (g1720)) + ((g1285) & (!g1437) & (g1660) & (g1661) & (!g1667) & (g1720)) + ((g1285) & (!g1437) & (g1660) & (g1661) & (g1667) & (!g1720)) + ((g1285) & (!g1437) & (g1660) & (g1661) & (g1667) & (g1720)) + ((g1285) & (g1437) & (!g1660) & (!g1661) & (!g1667) & (!g1720)) + ((g1285) & (g1437) & (g1660) & (!g1661) & (!g1667) & (g1720)) + ((g1285) & (g1437) & (g1660) & (!g1661) & (g1667) & (!g1720)) + ((g1285) & (g1437) & (g1660) & (!g1661) & (g1667) & (g1720)) + ((g1285) & (g1437) & (g1660) & (g1661) & (!g1667) & (!g1720)) + ((g1285) & (g1437) & (g1660) & (g1661) & (!g1667) & (g1720)) + ((g1285) & (g1437) & (g1660) & (g1661) & (g1667) & (!g1720)) + ((g1285) & (g1437) & (g1660) & (g1661) & (g1667) & (g1720)));
	assign g1739 = (((!g1437) & (!g1661) & (g1667) & (!g1720)) + ((!g1437) & (g1661) & (!g1667) & (!g1720)) + ((!g1437) & (g1661) & (!g1667) & (g1720)) + ((!g1437) & (g1661) & (g1667) & (g1720)) + ((g1437) & (!g1661) & (!g1667) & (!g1720)) + ((g1437) & (g1661) & (!g1667) & (g1720)) + ((g1437) & (g1661) & (g1667) & (!g1720)) + ((g1437) & (g1661) & (g1667) & (g1720)));
	assign g1740 = (((!g1423) & (!g1586) & (!g1663) & (g1664) & (g1666) & (!g1720)) + ((!g1423) & (!g1586) & (g1663) & (!g1664) & (!g1666) & (!g1720)) + ((!g1423) & (!g1586) & (g1663) & (!g1664) & (!g1666) & (g1720)) + ((!g1423) & (!g1586) & (g1663) & (!g1664) & (g1666) & (!g1720)) + ((!g1423) & (!g1586) & (g1663) & (!g1664) & (g1666) & (g1720)) + ((!g1423) & (!g1586) & (g1663) & (g1664) & (!g1666) & (!g1720)) + ((!g1423) & (!g1586) & (g1663) & (g1664) & (!g1666) & (g1720)) + ((!g1423) & (!g1586) & (g1663) & (g1664) & (g1666) & (g1720)) + ((!g1423) & (g1586) & (!g1663) & (!g1664) & (g1666) & (!g1720)) + ((!g1423) & (g1586) & (!g1663) & (g1664) & (!g1666) & (!g1720)) + ((!g1423) & (g1586) & (!g1663) & (g1664) & (g1666) & (!g1720)) + ((!g1423) & (g1586) & (g1663) & (!g1664) & (!g1666) & (!g1720)) + ((!g1423) & (g1586) & (g1663) & (!g1664) & (!g1666) & (g1720)) + ((!g1423) & (g1586) & (g1663) & (!g1664) & (g1666) & (g1720)) + ((!g1423) & (g1586) & (g1663) & (g1664) & (!g1666) & (g1720)) + ((!g1423) & (g1586) & (g1663) & (g1664) & (g1666) & (g1720)) + ((g1423) & (!g1586) & (!g1663) & (!g1664) & (!g1666) & (!g1720)) + ((g1423) & (!g1586) & (!g1663) & (!g1664) & (g1666) & (!g1720)) + ((g1423) & (!g1586) & (!g1663) & (g1664) & (!g1666) & (!g1720)) + ((g1423) & (!g1586) & (g1663) & (!g1664) & (!g1666) & (g1720)) + ((g1423) & (!g1586) & (g1663) & (!g1664) & (g1666) & (g1720)) + ((g1423) & (!g1586) & (g1663) & (g1664) & (!g1666) & (g1720)) + ((g1423) & (!g1586) & (g1663) & (g1664) & (g1666) & (!g1720)) + ((g1423) & (!g1586) & (g1663) & (g1664) & (g1666) & (g1720)) + ((g1423) & (g1586) & (!g1663) & (!g1664) & (!g1666) & (!g1720)) + ((g1423) & (g1586) & (g1663) & (!g1664) & (!g1666) & (g1720)) + ((g1423) & (g1586) & (g1663) & (!g1664) & (g1666) & (!g1720)) + ((g1423) & (g1586) & (g1663) & (!g1664) & (g1666) & (g1720)) + ((g1423) & (g1586) & (g1663) & (g1664) & (!g1666) & (!g1720)) + ((g1423) & (g1586) & (g1663) & (g1664) & (!g1666) & (g1720)) + ((g1423) & (g1586) & (g1663) & (g1664) & (g1666) & (!g1720)) + ((g1423) & (g1586) & (g1663) & (g1664) & (g1666) & (g1720)));
	assign g1741 = (((!g1586) & (!g1664) & (g1666) & (!g1720)) + ((!g1586) & (g1664) & (!g1666) & (!g1720)) + ((!g1586) & (g1664) & (!g1666) & (g1720)) + ((!g1586) & (g1664) & (g1666) & (g1720)) + ((g1586) & (!g1664) & (!g1666) & (!g1720)) + ((g1586) & (g1664) & (!g1666) & (g1720)) + ((g1586) & (g1664) & (g1666) & (!g1720)) + ((g1586) & (g1664) & (g1666) & (g1720)));
	assign g1742 = (((!g1600) & (g1633)));
	assign g1743 = (((!g1568) & (!ax42x) & (!ax43x) & (!g1742) & (!g1665) & (g1720)) + ((!g1568) & (!ax42x) & (!ax43x) & (!g1742) & (g1665) & (!g1720)) + ((!g1568) & (!ax42x) & (!ax43x) & (!g1742) & (g1665) & (g1720)) + ((!g1568) & (!ax42x) & (!ax43x) & (g1742) & (!g1665) & (!g1720)) + ((!g1568) & (!ax42x) & (ax43x) & (!g1742) & (!g1665) & (!g1720)) + ((!g1568) & (!ax42x) & (ax43x) & (g1742) & (!g1665) & (g1720)) + ((!g1568) & (!ax42x) & (ax43x) & (g1742) & (g1665) & (!g1720)) + ((!g1568) & (!ax42x) & (ax43x) & (g1742) & (g1665) & (g1720)) + ((!g1568) & (ax42x) & (!ax43x) & (g1742) & (!g1665) & (!g1720)) + ((!g1568) & (ax42x) & (!ax43x) & (g1742) & (g1665) & (!g1720)) + ((!g1568) & (ax42x) & (ax43x) & (!g1742) & (!g1665) & (!g1720)) + ((!g1568) & (ax42x) & (ax43x) & (!g1742) & (!g1665) & (g1720)) + ((!g1568) & (ax42x) & (ax43x) & (!g1742) & (g1665) & (!g1720)) + ((!g1568) & (ax42x) & (ax43x) & (!g1742) & (g1665) & (g1720)) + ((!g1568) & (ax42x) & (ax43x) & (g1742) & (!g1665) & (g1720)) + ((!g1568) & (ax42x) & (ax43x) & (g1742) & (g1665) & (g1720)) + ((g1568) & (!ax42x) & (!ax43x) & (!g1742) & (!g1665) & (!g1720)) + ((g1568) & (!ax42x) & (!ax43x) & (!g1742) & (!g1665) & (g1720)) + ((g1568) & (!ax42x) & (!ax43x) & (!g1742) & (g1665) & (g1720)) + ((g1568) & (!ax42x) & (!ax43x) & (g1742) & (g1665) & (!g1720)) + ((g1568) & (!ax42x) & (ax43x) & (!g1742) & (g1665) & (!g1720)) + ((g1568) & (!ax42x) & (ax43x) & (g1742) & (!g1665) & (!g1720)) + ((g1568) & (!ax42x) & (ax43x) & (g1742) & (!g1665) & (g1720)) + ((g1568) & (!ax42x) & (ax43x) & (g1742) & (g1665) & (g1720)) + ((g1568) & (ax42x) & (!ax43x) & (!g1742) & (!g1665) & (!g1720)) + ((g1568) & (ax42x) & (!ax43x) & (!g1742) & (g1665) & (!g1720)) + ((g1568) & (ax42x) & (ax43x) & (!g1742) & (!g1665) & (g1720)) + ((g1568) & (ax42x) & (ax43x) & (!g1742) & (g1665) & (g1720)) + ((g1568) & (ax42x) & (ax43x) & (g1742) & (!g1665) & (!g1720)) + ((g1568) & (ax42x) & (ax43x) & (g1742) & (!g1665) & (g1720)) + ((g1568) & (ax42x) & (ax43x) & (g1742) & (g1665) & (!g1720)) + ((g1568) & (ax42x) & (ax43x) & (g1742) & (g1665) & (g1720)));
	assign g1744 = (((!ax42x) & (!g1742) & (!g1665) & (g1720)) + ((!ax42x) & (!g1742) & (g1665) & (!g1720)) + ((!ax42x) & (!g1742) & (g1665) & (g1720)) + ((!ax42x) & (g1742) & (g1665) & (!g1720)) + ((ax42x) & (!g1742) & (!g1665) & (!g1720)) + ((ax42x) & (g1742) & (!g1665) & (!g1720)) + ((ax42x) & (g1742) & (!g1665) & (g1720)) + ((ax42x) & (g1742) & (g1665) & (g1720)));
	assign g1745 = (((!ax38x) & (!ax39x)));
	assign g1746 = (((!g1742) & (!ax40x) & (!ax41x) & (!g1720) & (!g1745)) + ((!g1742) & (!ax40x) & (ax41x) & (g1720) & (!g1745)) + ((!g1742) & (ax40x) & (ax41x) & (g1720) & (!g1745)) + ((!g1742) & (ax40x) & (ax41x) & (g1720) & (g1745)) + ((g1742) & (!ax40x) & (!ax41x) & (!g1720) & (!g1745)) + ((g1742) & (!ax40x) & (!ax41x) & (!g1720) & (g1745)) + ((g1742) & (!ax40x) & (!ax41x) & (g1720) & (!g1745)) + ((g1742) & (!ax40x) & (ax41x) & (!g1720) & (!g1745)) + ((g1742) & (!ax40x) & (ax41x) & (g1720) & (!g1745)) + ((g1742) & (!ax40x) & (ax41x) & (g1720) & (g1745)) + ((g1742) & (ax40x) & (!ax41x) & (g1720) & (!g1745)) + ((g1742) & (ax40x) & (!ax41x) & (g1720) & (g1745)) + ((g1742) & (ax40x) & (ax41x) & (!g1720) & (!g1745)) + ((g1742) & (ax40x) & (ax41x) & (!g1720) & (g1745)) + ((g1742) & (ax40x) & (ax41x) & (g1720) & (!g1745)) + ((g1742) & (ax40x) & (ax41x) & (g1720) & (g1745)));
	assign g1747 = (((!g1586) & (!g1568) & (g1743) & (g1744) & (g1746)) + ((!g1586) & (g1568) & (g1743) & (!g1744) & (g1746)) + ((!g1586) & (g1568) & (g1743) & (g1744) & (!g1746)) + ((!g1586) & (g1568) & (g1743) & (g1744) & (g1746)) + ((g1586) & (!g1568) & (!g1743) & (g1744) & (g1746)) + ((g1586) & (!g1568) & (g1743) & (!g1744) & (!g1746)) + ((g1586) & (!g1568) & (g1743) & (!g1744) & (g1746)) + ((g1586) & (!g1568) & (g1743) & (g1744) & (!g1746)) + ((g1586) & (!g1568) & (g1743) & (g1744) & (g1746)) + ((g1586) & (g1568) & (!g1743) & (!g1744) & (g1746)) + ((g1586) & (g1568) & (!g1743) & (g1744) & (!g1746)) + ((g1586) & (g1568) & (!g1743) & (g1744) & (g1746)) + ((g1586) & (g1568) & (g1743) & (!g1744) & (!g1746)) + ((g1586) & (g1568) & (g1743) & (!g1744) & (g1746)) + ((g1586) & (g1568) & (g1743) & (g1744) & (!g1746)) + ((g1586) & (g1568) & (g1743) & (g1744) & (g1746)));
	assign g1748 = (((!g1437) & (!g1423) & (g1740) & (g1741) & (g1747)) + ((!g1437) & (g1423) & (g1740) & (!g1741) & (g1747)) + ((!g1437) & (g1423) & (g1740) & (g1741) & (!g1747)) + ((!g1437) & (g1423) & (g1740) & (g1741) & (g1747)) + ((g1437) & (!g1423) & (!g1740) & (g1741) & (g1747)) + ((g1437) & (!g1423) & (g1740) & (!g1741) & (!g1747)) + ((g1437) & (!g1423) & (g1740) & (!g1741) & (g1747)) + ((g1437) & (!g1423) & (g1740) & (g1741) & (!g1747)) + ((g1437) & (!g1423) & (g1740) & (g1741) & (g1747)) + ((g1437) & (g1423) & (!g1740) & (!g1741) & (g1747)) + ((g1437) & (g1423) & (!g1740) & (g1741) & (!g1747)) + ((g1437) & (g1423) & (!g1740) & (g1741) & (g1747)) + ((g1437) & (g1423) & (g1740) & (!g1741) & (!g1747)) + ((g1437) & (g1423) & (g1740) & (!g1741) & (g1747)) + ((g1437) & (g1423) & (g1740) & (g1741) & (!g1747)) + ((g1437) & (g1423) & (g1740) & (g1741) & (g1747)));
	assign g1749 = (((!g1295) & (!g1285) & (g1738) & (g1739) & (g1748)) + ((!g1295) & (g1285) & (g1738) & (!g1739) & (g1748)) + ((!g1295) & (g1285) & (g1738) & (g1739) & (!g1748)) + ((!g1295) & (g1285) & (g1738) & (g1739) & (g1748)) + ((g1295) & (!g1285) & (!g1738) & (g1739) & (g1748)) + ((g1295) & (!g1285) & (g1738) & (!g1739) & (!g1748)) + ((g1295) & (!g1285) & (g1738) & (!g1739) & (g1748)) + ((g1295) & (!g1285) & (g1738) & (g1739) & (!g1748)) + ((g1295) & (!g1285) & (g1738) & (g1739) & (g1748)) + ((g1295) & (g1285) & (!g1738) & (!g1739) & (g1748)) + ((g1295) & (g1285) & (!g1738) & (g1739) & (!g1748)) + ((g1295) & (g1285) & (!g1738) & (g1739) & (g1748)) + ((g1295) & (g1285) & (g1738) & (!g1739) & (!g1748)) + ((g1295) & (g1285) & (g1738) & (!g1739) & (g1748)) + ((g1295) & (g1285) & (g1738) & (g1739) & (!g1748)) + ((g1295) & (g1285) & (g1738) & (g1739) & (g1748)));
	assign g1750 = (((!g1160) & (!g1154) & (g1736) & (g1737) & (g1749)) + ((!g1160) & (g1154) & (g1736) & (!g1737) & (g1749)) + ((!g1160) & (g1154) & (g1736) & (g1737) & (!g1749)) + ((!g1160) & (g1154) & (g1736) & (g1737) & (g1749)) + ((g1160) & (!g1154) & (!g1736) & (g1737) & (g1749)) + ((g1160) & (!g1154) & (g1736) & (!g1737) & (!g1749)) + ((g1160) & (!g1154) & (g1736) & (!g1737) & (g1749)) + ((g1160) & (!g1154) & (g1736) & (g1737) & (!g1749)) + ((g1160) & (!g1154) & (g1736) & (g1737) & (g1749)) + ((g1160) & (g1154) & (!g1736) & (!g1737) & (g1749)) + ((g1160) & (g1154) & (!g1736) & (g1737) & (!g1749)) + ((g1160) & (g1154) & (!g1736) & (g1737) & (g1749)) + ((g1160) & (g1154) & (g1736) & (!g1737) & (!g1749)) + ((g1160) & (g1154) & (g1736) & (!g1737) & (g1749)) + ((g1160) & (g1154) & (g1736) & (g1737) & (!g1749)) + ((g1160) & (g1154) & (g1736) & (g1737) & (g1749)));
	assign g1751 = (((!g1032) & (!g1030) & (g1734) & (g1735) & (g1750)) + ((!g1032) & (g1030) & (g1734) & (!g1735) & (g1750)) + ((!g1032) & (g1030) & (g1734) & (g1735) & (!g1750)) + ((!g1032) & (g1030) & (g1734) & (g1735) & (g1750)) + ((g1032) & (!g1030) & (!g1734) & (g1735) & (g1750)) + ((g1032) & (!g1030) & (g1734) & (!g1735) & (!g1750)) + ((g1032) & (!g1030) & (g1734) & (!g1735) & (g1750)) + ((g1032) & (!g1030) & (g1734) & (g1735) & (!g1750)) + ((g1032) & (!g1030) & (g1734) & (g1735) & (g1750)) + ((g1032) & (g1030) & (!g1734) & (!g1735) & (g1750)) + ((g1032) & (g1030) & (!g1734) & (g1735) & (!g1750)) + ((g1032) & (g1030) & (!g1734) & (g1735) & (g1750)) + ((g1032) & (g1030) & (g1734) & (!g1735) & (!g1750)) + ((g1032) & (g1030) & (g1734) & (!g1735) & (g1750)) + ((g1032) & (g1030) & (g1734) & (g1735) & (!g1750)) + ((g1032) & (g1030) & (g1734) & (g1735) & (g1750)));
	assign g1752 = (((!g851) & (!g914) & (g1732) & (g1733) & (g1751)) + ((!g851) & (g914) & (g1732) & (!g1733) & (g1751)) + ((!g851) & (g914) & (g1732) & (g1733) & (!g1751)) + ((!g851) & (g914) & (g1732) & (g1733) & (g1751)) + ((g851) & (!g914) & (!g1732) & (g1733) & (g1751)) + ((g851) & (!g914) & (g1732) & (!g1733) & (!g1751)) + ((g851) & (!g914) & (g1732) & (!g1733) & (g1751)) + ((g851) & (!g914) & (g1732) & (g1733) & (!g1751)) + ((g851) & (!g914) & (g1732) & (g1733) & (g1751)) + ((g851) & (g914) & (!g1732) & (!g1733) & (g1751)) + ((g851) & (g914) & (!g1732) & (g1733) & (!g1751)) + ((g851) & (g914) & (!g1732) & (g1733) & (g1751)) + ((g851) & (g914) & (g1732) & (!g1733) & (!g1751)) + ((g851) & (g914) & (g1732) & (!g1733) & (g1751)) + ((g851) & (g914) & (g1732) & (g1733) & (!g1751)) + ((g851) & (g914) & (g1732) & (g1733) & (g1751)));
	assign g1753 = (((!g744) & (!g803) & (g1730) & (g1731) & (g1752)) + ((!g744) & (g803) & (g1730) & (!g1731) & (g1752)) + ((!g744) & (g803) & (g1730) & (g1731) & (!g1752)) + ((!g744) & (g803) & (g1730) & (g1731) & (g1752)) + ((g744) & (!g803) & (!g1730) & (g1731) & (g1752)) + ((g744) & (!g803) & (g1730) & (!g1731) & (!g1752)) + ((g744) & (!g803) & (g1730) & (!g1731) & (g1752)) + ((g744) & (!g803) & (g1730) & (g1731) & (!g1752)) + ((g744) & (!g803) & (g1730) & (g1731) & (g1752)) + ((g744) & (g803) & (!g1730) & (!g1731) & (g1752)) + ((g744) & (g803) & (!g1730) & (g1731) & (!g1752)) + ((g744) & (g803) & (!g1730) & (g1731) & (g1752)) + ((g744) & (g803) & (g1730) & (!g1731) & (!g1752)) + ((g744) & (g803) & (g1730) & (!g1731) & (g1752)) + ((g744) & (g803) & (g1730) & (g1731) & (!g1752)) + ((g744) & (g803) & (g1730) & (g1731) & (g1752)));
	assign g1754 = (((!g645) & (!g700) & (g1728) & (g1729) & (g1753)) + ((!g645) & (g700) & (g1728) & (!g1729) & (g1753)) + ((!g645) & (g700) & (g1728) & (g1729) & (!g1753)) + ((!g645) & (g700) & (g1728) & (g1729) & (g1753)) + ((g645) & (!g700) & (!g1728) & (g1729) & (g1753)) + ((g645) & (!g700) & (g1728) & (!g1729) & (!g1753)) + ((g645) & (!g700) & (g1728) & (!g1729) & (g1753)) + ((g645) & (!g700) & (g1728) & (g1729) & (!g1753)) + ((g645) & (!g700) & (g1728) & (g1729) & (g1753)) + ((g645) & (g700) & (!g1728) & (!g1729) & (g1753)) + ((g645) & (g700) & (!g1728) & (g1729) & (!g1753)) + ((g645) & (g700) & (!g1728) & (g1729) & (g1753)) + ((g645) & (g700) & (g1728) & (!g1729) & (!g1753)) + ((g645) & (g700) & (g1728) & (!g1729) & (g1753)) + ((g645) & (g700) & (g1728) & (g1729) & (!g1753)) + ((g645) & (g700) & (g1728) & (g1729) & (g1753)));
	assign g1755 = (((!g553) & (!g604) & (g1726) & (g1727) & (g1754)) + ((!g553) & (g604) & (g1726) & (!g1727) & (g1754)) + ((!g553) & (g604) & (g1726) & (g1727) & (!g1754)) + ((!g553) & (g604) & (g1726) & (g1727) & (g1754)) + ((g553) & (!g604) & (!g1726) & (g1727) & (g1754)) + ((g553) & (!g604) & (g1726) & (!g1727) & (!g1754)) + ((g553) & (!g604) & (g1726) & (!g1727) & (g1754)) + ((g553) & (!g604) & (g1726) & (g1727) & (!g1754)) + ((g553) & (!g604) & (g1726) & (g1727) & (g1754)) + ((g553) & (g604) & (!g1726) & (!g1727) & (g1754)) + ((g553) & (g604) & (!g1726) & (g1727) & (!g1754)) + ((g553) & (g604) & (!g1726) & (g1727) & (g1754)) + ((g553) & (g604) & (g1726) & (!g1727) & (!g1754)) + ((g553) & (g604) & (g1726) & (!g1727) & (g1754)) + ((g553) & (g604) & (g1726) & (g1727) & (!g1754)) + ((g553) & (g604) & (g1726) & (g1727) & (g1754)));
	assign g1756 = (((!g468) & (!g515) & (g1724) & (g1725) & (g1755)) + ((!g468) & (g515) & (g1724) & (!g1725) & (g1755)) + ((!g468) & (g515) & (g1724) & (g1725) & (!g1755)) + ((!g468) & (g515) & (g1724) & (g1725) & (g1755)) + ((g468) & (!g515) & (!g1724) & (g1725) & (g1755)) + ((g468) & (!g515) & (g1724) & (!g1725) & (!g1755)) + ((g468) & (!g515) & (g1724) & (!g1725) & (g1755)) + ((g468) & (!g515) & (g1724) & (g1725) & (!g1755)) + ((g468) & (!g515) & (g1724) & (g1725) & (g1755)) + ((g468) & (g515) & (!g1724) & (!g1725) & (g1755)) + ((g468) & (g515) & (!g1724) & (g1725) & (!g1755)) + ((g468) & (g515) & (!g1724) & (g1725) & (g1755)) + ((g468) & (g515) & (g1724) & (!g1725) & (!g1755)) + ((g468) & (g515) & (g1724) & (!g1725) & (g1755)) + ((g468) & (g515) & (g1724) & (g1725) & (!g1755)) + ((g468) & (g515) & (g1724) & (g1725) & (g1755)));
	assign g1757 = (((!g390) & (!g433) & (g1722) & (g1723) & (g1756)) + ((!g390) & (g433) & (g1722) & (!g1723) & (g1756)) + ((!g390) & (g433) & (g1722) & (g1723) & (!g1756)) + ((!g390) & (g433) & (g1722) & (g1723) & (g1756)) + ((g390) & (!g433) & (!g1722) & (g1723) & (g1756)) + ((g390) & (!g433) & (g1722) & (!g1723) & (!g1756)) + ((g390) & (!g433) & (g1722) & (!g1723) & (g1756)) + ((g390) & (!g433) & (g1722) & (g1723) & (!g1756)) + ((g390) & (!g433) & (g1722) & (g1723) & (g1756)) + ((g390) & (g433) & (!g1722) & (!g1723) & (g1756)) + ((g390) & (g433) & (!g1722) & (g1723) & (!g1756)) + ((g390) & (g433) & (!g1722) & (g1723) & (g1756)) + ((g390) & (g433) & (g1722) & (!g1723) & (!g1756)) + ((g390) & (g433) & (g1722) & (!g1723) & (g1756)) + ((g390) & (g433) & (g1722) & (g1723) & (!g1756)) + ((g390) & (g433) & (g1722) & (g1723) & (g1756)));
	assign g1758 = (((g1) & (!g1677) & (g1716) & (g1719)) + ((g1) & (g1677) & (!g1716) & (!g1719)) + ((g1) & (g1677) & (!g1716) & (g1719)));
	assign g1759 = (((!g4) & (!g2) & (!g1678) & (!g1713) & (!g1715) & (!g1720)) + ((!g4) & (!g2) & (!g1678) & (!g1713) & (g1715) & (g1720)) + ((!g4) & (!g2) & (!g1678) & (g1713) & (!g1715) & (!g1720)) + ((!g4) & (!g2) & (!g1678) & (g1713) & (g1715) & (g1720)) + ((!g4) & (!g2) & (g1678) & (!g1713) & (!g1715) & (!g1720)) + ((!g4) & (!g2) & (g1678) & (!g1713) & (g1715) & (g1720)) + ((!g4) & (!g2) & (g1678) & (g1713) & (g1715) & (!g1720)) + ((!g4) & (!g2) & (g1678) & (g1713) & (g1715) & (g1720)) + ((!g4) & (g2) & (!g1678) & (!g1713) & (!g1715) & (!g1720)) + ((!g4) & (g2) & (!g1678) & (!g1713) & (g1715) & (g1720)) + ((!g4) & (g2) & (!g1678) & (g1713) & (g1715) & (!g1720)) + ((!g4) & (g2) & (!g1678) & (g1713) & (g1715) & (g1720)) + ((!g4) & (g2) & (g1678) & (!g1713) & (g1715) & (!g1720)) + ((!g4) & (g2) & (g1678) & (!g1713) & (g1715) & (g1720)) + ((!g4) & (g2) & (g1678) & (g1713) & (g1715) & (!g1720)) + ((!g4) & (g2) & (g1678) & (g1713) & (g1715) & (g1720)) + ((g4) & (!g2) & (!g1678) & (!g1713) & (g1715) & (!g1720)) + ((g4) & (!g2) & (!g1678) & (!g1713) & (g1715) & (g1720)) + ((g4) & (!g2) & (!g1678) & (g1713) & (g1715) & (!g1720)) + ((g4) & (!g2) & (!g1678) & (g1713) & (g1715) & (g1720)) + ((g4) & (!g2) & (g1678) & (!g1713) & (g1715) & (!g1720)) + ((g4) & (!g2) & (g1678) & (!g1713) & (g1715) & (g1720)) + ((g4) & (!g2) & (g1678) & (g1713) & (!g1715) & (!g1720)) + ((g4) & (!g2) & (g1678) & (g1713) & (g1715) & (g1720)) + ((g4) & (g2) & (!g1678) & (!g1713) & (g1715) & (!g1720)) + ((g4) & (g2) & (!g1678) & (!g1713) & (g1715) & (g1720)) + ((g4) & (g2) & (!g1678) & (g1713) & (!g1715) & (!g1720)) + ((g4) & (g2) & (!g1678) & (g1713) & (g1715) & (g1720)) + ((g4) & (g2) & (g1678) & (!g1713) & (!g1715) & (!g1720)) + ((g4) & (g2) & (g1678) & (!g1713) & (g1715) & (g1720)) + ((g4) & (g2) & (g1678) & (g1713) & (!g1715) & (!g1720)) + ((g4) & (g2) & (g1678) & (g1713) & (g1715) & (g1720)));
	assign g1760 = (((!g8) & (!g18) & (!g1680) & (g1681) & (g1712) & (!g1720)) + ((!g8) & (!g18) & (g1680) & (!g1681) & (!g1712) & (!g1720)) + ((!g8) & (!g18) & (g1680) & (!g1681) & (!g1712) & (g1720)) + ((!g8) & (!g18) & (g1680) & (!g1681) & (g1712) & (!g1720)) + ((!g8) & (!g18) & (g1680) & (!g1681) & (g1712) & (g1720)) + ((!g8) & (!g18) & (g1680) & (g1681) & (!g1712) & (!g1720)) + ((!g8) & (!g18) & (g1680) & (g1681) & (!g1712) & (g1720)) + ((!g8) & (!g18) & (g1680) & (g1681) & (g1712) & (g1720)) + ((!g8) & (g18) & (!g1680) & (!g1681) & (g1712) & (!g1720)) + ((!g8) & (g18) & (!g1680) & (g1681) & (!g1712) & (!g1720)) + ((!g8) & (g18) & (!g1680) & (g1681) & (g1712) & (!g1720)) + ((!g8) & (g18) & (g1680) & (!g1681) & (!g1712) & (!g1720)) + ((!g8) & (g18) & (g1680) & (!g1681) & (!g1712) & (g1720)) + ((!g8) & (g18) & (g1680) & (!g1681) & (g1712) & (g1720)) + ((!g8) & (g18) & (g1680) & (g1681) & (!g1712) & (g1720)) + ((!g8) & (g18) & (g1680) & (g1681) & (g1712) & (g1720)) + ((g8) & (!g18) & (!g1680) & (!g1681) & (!g1712) & (!g1720)) + ((g8) & (!g18) & (!g1680) & (!g1681) & (g1712) & (!g1720)) + ((g8) & (!g18) & (!g1680) & (g1681) & (!g1712) & (!g1720)) + ((g8) & (!g18) & (g1680) & (!g1681) & (!g1712) & (g1720)) + ((g8) & (!g18) & (g1680) & (!g1681) & (g1712) & (g1720)) + ((g8) & (!g18) & (g1680) & (g1681) & (!g1712) & (g1720)) + ((g8) & (!g18) & (g1680) & (g1681) & (g1712) & (!g1720)) + ((g8) & (!g18) & (g1680) & (g1681) & (g1712) & (g1720)) + ((g8) & (g18) & (!g1680) & (!g1681) & (!g1712) & (!g1720)) + ((g8) & (g18) & (g1680) & (!g1681) & (!g1712) & (g1720)) + ((g8) & (g18) & (g1680) & (!g1681) & (g1712) & (!g1720)) + ((g8) & (g18) & (g1680) & (!g1681) & (g1712) & (g1720)) + ((g8) & (g18) & (g1680) & (g1681) & (!g1712) & (!g1720)) + ((g8) & (g18) & (g1680) & (g1681) & (!g1712) & (g1720)) + ((g8) & (g18) & (g1680) & (g1681) & (g1712) & (!g1720)) + ((g8) & (g18) & (g1680) & (g1681) & (g1712) & (g1720)));
	assign g1761 = (((!g18) & (!g1681) & (g1712) & (!g1720)) + ((!g18) & (g1681) & (!g1712) & (!g1720)) + ((!g18) & (g1681) & (!g1712) & (g1720)) + ((!g18) & (g1681) & (g1712) & (g1720)) + ((g18) & (!g1681) & (!g1712) & (!g1720)) + ((g18) & (g1681) & (!g1712) & (g1720)) + ((g18) & (g1681) & (g1712) & (!g1720)) + ((g18) & (g1681) & (g1712) & (g1720)));
	assign g1762 = (((!g27) & (!g39) & (!g1683) & (g1684) & (g1711) & (!g1720)) + ((!g27) & (!g39) & (g1683) & (!g1684) & (!g1711) & (!g1720)) + ((!g27) & (!g39) & (g1683) & (!g1684) & (!g1711) & (g1720)) + ((!g27) & (!g39) & (g1683) & (!g1684) & (g1711) & (!g1720)) + ((!g27) & (!g39) & (g1683) & (!g1684) & (g1711) & (g1720)) + ((!g27) & (!g39) & (g1683) & (g1684) & (!g1711) & (!g1720)) + ((!g27) & (!g39) & (g1683) & (g1684) & (!g1711) & (g1720)) + ((!g27) & (!g39) & (g1683) & (g1684) & (g1711) & (g1720)) + ((!g27) & (g39) & (!g1683) & (!g1684) & (g1711) & (!g1720)) + ((!g27) & (g39) & (!g1683) & (g1684) & (!g1711) & (!g1720)) + ((!g27) & (g39) & (!g1683) & (g1684) & (g1711) & (!g1720)) + ((!g27) & (g39) & (g1683) & (!g1684) & (!g1711) & (!g1720)) + ((!g27) & (g39) & (g1683) & (!g1684) & (!g1711) & (g1720)) + ((!g27) & (g39) & (g1683) & (!g1684) & (g1711) & (g1720)) + ((!g27) & (g39) & (g1683) & (g1684) & (!g1711) & (g1720)) + ((!g27) & (g39) & (g1683) & (g1684) & (g1711) & (g1720)) + ((g27) & (!g39) & (!g1683) & (!g1684) & (!g1711) & (!g1720)) + ((g27) & (!g39) & (!g1683) & (!g1684) & (g1711) & (!g1720)) + ((g27) & (!g39) & (!g1683) & (g1684) & (!g1711) & (!g1720)) + ((g27) & (!g39) & (g1683) & (!g1684) & (!g1711) & (g1720)) + ((g27) & (!g39) & (g1683) & (!g1684) & (g1711) & (g1720)) + ((g27) & (!g39) & (g1683) & (g1684) & (!g1711) & (g1720)) + ((g27) & (!g39) & (g1683) & (g1684) & (g1711) & (!g1720)) + ((g27) & (!g39) & (g1683) & (g1684) & (g1711) & (g1720)) + ((g27) & (g39) & (!g1683) & (!g1684) & (!g1711) & (!g1720)) + ((g27) & (g39) & (g1683) & (!g1684) & (!g1711) & (g1720)) + ((g27) & (g39) & (g1683) & (!g1684) & (g1711) & (!g1720)) + ((g27) & (g39) & (g1683) & (!g1684) & (g1711) & (g1720)) + ((g27) & (g39) & (g1683) & (g1684) & (!g1711) & (!g1720)) + ((g27) & (g39) & (g1683) & (g1684) & (!g1711) & (g1720)) + ((g27) & (g39) & (g1683) & (g1684) & (g1711) & (!g1720)) + ((g27) & (g39) & (g1683) & (g1684) & (g1711) & (g1720)));
	assign g1763 = (((!g39) & (!g1684) & (g1711) & (!g1720)) + ((!g39) & (g1684) & (!g1711) & (!g1720)) + ((!g39) & (g1684) & (!g1711) & (g1720)) + ((!g39) & (g1684) & (g1711) & (g1720)) + ((g39) & (!g1684) & (!g1711) & (!g1720)) + ((g39) & (g1684) & (!g1711) & (g1720)) + ((g39) & (g1684) & (g1711) & (!g1720)) + ((g39) & (g1684) & (g1711) & (g1720)));
	assign g1764 = (((!g54) & (!g68) & (!g1686) & (g1687) & (g1710) & (!g1720)) + ((!g54) & (!g68) & (g1686) & (!g1687) & (!g1710) & (!g1720)) + ((!g54) & (!g68) & (g1686) & (!g1687) & (!g1710) & (g1720)) + ((!g54) & (!g68) & (g1686) & (!g1687) & (g1710) & (!g1720)) + ((!g54) & (!g68) & (g1686) & (!g1687) & (g1710) & (g1720)) + ((!g54) & (!g68) & (g1686) & (g1687) & (!g1710) & (!g1720)) + ((!g54) & (!g68) & (g1686) & (g1687) & (!g1710) & (g1720)) + ((!g54) & (!g68) & (g1686) & (g1687) & (g1710) & (g1720)) + ((!g54) & (g68) & (!g1686) & (!g1687) & (g1710) & (!g1720)) + ((!g54) & (g68) & (!g1686) & (g1687) & (!g1710) & (!g1720)) + ((!g54) & (g68) & (!g1686) & (g1687) & (g1710) & (!g1720)) + ((!g54) & (g68) & (g1686) & (!g1687) & (!g1710) & (!g1720)) + ((!g54) & (g68) & (g1686) & (!g1687) & (!g1710) & (g1720)) + ((!g54) & (g68) & (g1686) & (!g1687) & (g1710) & (g1720)) + ((!g54) & (g68) & (g1686) & (g1687) & (!g1710) & (g1720)) + ((!g54) & (g68) & (g1686) & (g1687) & (g1710) & (g1720)) + ((g54) & (!g68) & (!g1686) & (!g1687) & (!g1710) & (!g1720)) + ((g54) & (!g68) & (!g1686) & (!g1687) & (g1710) & (!g1720)) + ((g54) & (!g68) & (!g1686) & (g1687) & (!g1710) & (!g1720)) + ((g54) & (!g68) & (g1686) & (!g1687) & (!g1710) & (g1720)) + ((g54) & (!g68) & (g1686) & (!g1687) & (g1710) & (g1720)) + ((g54) & (!g68) & (g1686) & (g1687) & (!g1710) & (g1720)) + ((g54) & (!g68) & (g1686) & (g1687) & (g1710) & (!g1720)) + ((g54) & (!g68) & (g1686) & (g1687) & (g1710) & (g1720)) + ((g54) & (g68) & (!g1686) & (!g1687) & (!g1710) & (!g1720)) + ((g54) & (g68) & (g1686) & (!g1687) & (!g1710) & (g1720)) + ((g54) & (g68) & (g1686) & (!g1687) & (g1710) & (!g1720)) + ((g54) & (g68) & (g1686) & (!g1687) & (g1710) & (g1720)) + ((g54) & (g68) & (g1686) & (g1687) & (!g1710) & (!g1720)) + ((g54) & (g68) & (g1686) & (g1687) & (!g1710) & (g1720)) + ((g54) & (g68) & (g1686) & (g1687) & (g1710) & (!g1720)) + ((g54) & (g68) & (g1686) & (g1687) & (g1710) & (g1720)));
	assign g1765 = (((!g68) & (!g1687) & (g1710) & (!g1720)) + ((!g68) & (g1687) & (!g1710) & (!g1720)) + ((!g68) & (g1687) & (!g1710) & (g1720)) + ((!g68) & (g1687) & (g1710) & (g1720)) + ((g68) & (!g1687) & (!g1710) & (!g1720)) + ((g68) & (g1687) & (!g1710) & (g1720)) + ((g68) & (g1687) & (g1710) & (!g1720)) + ((g68) & (g1687) & (g1710) & (g1720)));
	assign g1766 = (((!g87) & (!g104) & (!g1689) & (g1690) & (g1709) & (!g1720)) + ((!g87) & (!g104) & (g1689) & (!g1690) & (!g1709) & (!g1720)) + ((!g87) & (!g104) & (g1689) & (!g1690) & (!g1709) & (g1720)) + ((!g87) & (!g104) & (g1689) & (!g1690) & (g1709) & (!g1720)) + ((!g87) & (!g104) & (g1689) & (!g1690) & (g1709) & (g1720)) + ((!g87) & (!g104) & (g1689) & (g1690) & (!g1709) & (!g1720)) + ((!g87) & (!g104) & (g1689) & (g1690) & (!g1709) & (g1720)) + ((!g87) & (!g104) & (g1689) & (g1690) & (g1709) & (g1720)) + ((!g87) & (g104) & (!g1689) & (!g1690) & (g1709) & (!g1720)) + ((!g87) & (g104) & (!g1689) & (g1690) & (!g1709) & (!g1720)) + ((!g87) & (g104) & (!g1689) & (g1690) & (g1709) & (!g1720)) + ((!g87) & (g104) & (g1689) & (!g1690) & (!g1709) & (!g1720)) + ((!g87) & (g104) & (g1689) & (!g1690) & (!g1709) & (g1720)) + ((!g87) & (g104) & (g1689) & (!g1690) & (g1709) & (g1720)) + ((!g87) & (g104) & (g1689) & (g1690) & (!g1709) & (g1720)) + ((!g87) & (g104) & (g1689) & (g1690) & (g1709) & (g1720)) + ((g87) & (!g104) & (!g1689) & (!g1690) & (!g1709) & (!g1720)) + ((g87) & (!g104) & (!g1689) & (!g1690) & (g1709) & (!g1720)) + ((g87) & (!g104) & (!g1689) & (g1690) & (!g1709) & (!g1720)) + ((g87) & (!g104) & (g1689) & (!g1690) & (!g1709) & (g1720)) + ((g87) & (!g104) & (g1689) & (!g1690) & (g1709) & (g1720)) + ((g87) & (!g104) & (g1689) & (g1690) & (!g1709) & (g1720)) + ((g87) & (!g104) & (g1689) & (g1690) & (g1709) & (!g1720)) + ((g87) & (!g104) & (g1689) & (g1690) & (g1709) & (g1720)) + ((g87) & (g104) & (!g1689) & (!g1690) & (!g1709) & (!g1720)) + ((g87) & (g104) & (g1689) & (!g1690) & (!g1709) & (g1720)) + ((g87) & (g104) & (g1689) & (!g1690) & (g1709) & (!g1720)) + ((g87) & (g104) & (g1689) & (!g1690) & (g1709) & (g1720)) + ((g87) & (g104) & (g1689) & (g1690) & (!g1709) & (!g1720)) + ((g87) & (g104) & (g1689) & (g1690) & (!g1709) & (g1720)) + ((g87) & (g104) & (g1689) & (g1690) & (g1709) & (!g1720)) + ((g87) & (g104) & (g1689) & (g1690) & (g1709) & (g1720)));
	assign g1767 = (((!g104) & (!g1690) & (g1709) & (!g1720)) + ((!g104) & (g1690) & (!g1709) & (!g1720)) + ((!g104) & (g1690) & (!g1709) & (g1720)) + ((!g104) & (g1690) & (g1709) & (g1720)) + ((g104) & (!g1690) & (!g1709) & (!g1720)) + ((g104) & (g1690) & (!g1709) & (g1720)) + ((g104) & (g1690) & (g1709) & (!g1720)) + ((g104) & (g1690) & (g1709) & (g1720)));
	assign g1768 = (((!g127) & (!g147) & (!g1692) & (g1693) & (g1708) & (!g1720)) + ((!g127) & (!g147) & (g1692) & (!g1693) & (!g1708) & (!g1720)) + ((!g127) & (!g147) & (g1692) & (!g1693) & (!g1708) & (g1720)) + ((!g127) & (!g147) & (g1692) & (!g1693) & (g1708) & (!g1720)) + ((!g127) & (!g147) & (g1692) & (!g1693) & (g1708) & (g1720)) + ((!g127) & (!g147) & (g1692) & (g1693) & (!g1708) & (!g1720)) + ((!g127) & (!g147) & (g1692) & (g1693) & (!g1708) & (g1720)) + ((!g127) & (!g147) & (g1692) & (g1693) & (g1708) & (g1720)) + ((!g127) & (g147) & (!g1692) & (!g1693) & (g1708) & (!g1720)) + ((!g127) & (g147) & (!g1692) & (g1693) & (!g1708) & (!g1720)) + ((!g127) & (g147) & (!g1692) & (g1693) & (g1708) & (!g1720)) + ((!g127) & (g147) & (g1692) & (!g1693) & (!g1708) & (!g1720)) + ((!g127) & (g147) & (g1692) & (!g1693) & (!g1708) & (g1720)) + ((!g127) & (g147) & (g1692) & (!g1693) & (g1708) & (g1720)) + ((!g127) & (g147) & (g1692) & (g1693) & (!g1708) & (g1720)) + ((!g127) & (g147) & (g1692) & (g1693) & (g1708) & (g1720)) + ((g127) & (!g147) & (!g1692) & (!g1693) & (!g1708) & (!g1720)) + ((g127) & (!g147) & (!g1692) & (!g1693) & (g1708) & (!g1720)) + ((g127) & (!g147) & (!g1692) & (g1693) & (!g1708) & (!g1720)) + ((g127) & (!g147) & (g1692) & (!g1693) & (!g1708) & (g1720)) + ((g127) & (!g147) & (g1692) & (!g1693) & (g1708) & (g1720)) + ((g127) & (!g147) & (g1692) & (g1693) & (!g1708) & (g1720)) + ((g127) & (!g147) & (g1692) & (g1693) & (g1708) & (!g1720)) + ((g127) & (!g147) & (g1692) & (g1693) & (g1708) & (g1720)) + ((g127) & (g147) & (!g1692) & (!g1693) & (!g1708) & (!g1720)) + ((g127) & (g147) & (g1692) & (!g1693) & (!g1708) & (g1720)) + ((g127) & (g147) & (g1692) & (!g1693) & (g1708) & (!g1720)) + ((g127) & (g147) & (g1692) & (!g1693) & (g1708) & (g1720)) + ((g127) & (g147) & (g1692) & (g1693) & (!g1708) & (!g1720)) + ((g127) & (g147) & (g1692) & (g1693) & (!g1708) & (g1720)) + ((g127) & (g147) & (g1692) & (g1693) & (g1708) & (!g1720)) + ((g127) & (g147) & (g1692) & (g1693) & (g1708) & (g1720)));
	assign g1769 = (((!g147) & (!g1693) & (g1708) & (!g1720)) + ((!g147) & (g1693) & (!g1708) & (!g1720)) + ((!g147) & (g1693) & (!g1708) & (g1720)) + ((!g147) & (g1693) & (g1708) & (g1720)) + ((g147) & (!g1693) & (!g1708) & (!g1720)) + ((g147) & (g1693) & (!g1708) & (g1720)) + ((g147) & (g1693) & (g1708) & (!g1720)) + ((g147) & (g1693) & (g1708) & (g1720)));
	assign g1770 = (((!g174) & (!g198) & (!g1695) & (g1696) & (g1707) & (!g1720)) + ((!g174) & (!g198) & (g1695) & (!g1696) & (!g1707) & (!g1720)) + ((!g174) & (!g198) & (g1695) & (!g1696) & (!g1707) & (g1720)) + ((!g174) & (!g198) & (g1695) & (!g1696) & (g1707) & (!g1720)) + ((!g174) & (!g198) & (g1695) & (!g1696) & (g1707) & (g1720)) + ((!g174) & (!g198) & (g1695) & (g1696) & (!g1707) & (!g1720)) + ((!g174) & (!g198) & (g1695) & (g1696) & (!g1707) & (g1720)) + ((!g174) & (!g198) & (g1695) & (g1696) & (g1707) & (g1720)) + ((!g174) & (g198) & (!g1695) & (!g1696) & (g1707) & (!g1720)) + ((!g174) & (g198) & (!g1695) & (g1696) & (!g1707) & (!g1720)) + ((!g174) & (g198) & (!g1695) & (g1696) & (g1707) & (!g1720)) + ((!g174) & (g198) & (g1695) & (!g1696) & (!g1707) & (!g1720)) + ((!g174) & (g198) & (g1695) & (!g1696) & (!g1707) & (g1720)) + ((!g174) & (g198) & (g1695) & (!g1696) & (g1707) & (g1720)) + ((!g174) & (g198) & (g1695) & (g1696) & (!g1707) & (g1720)) + ((!g174) & (g198) & (g1695) & (g1696) & (g1707) & (g1720)) + ((g174) & (!g198) & (!g1695) & (!g1696) & (!g1707) & (!g1720)) + ((g174) & (!g198) & (!g1695) & (!g1696) & (g1707) & (!g1720)) + ((g174) & (!g198) & (!g1695) & (g1696) & (!g1707) & (!g1720)) + ((g174) & (!g198) & (g1695) & (!g1696) & (!g1707) & (g1720)) + ((g174) & (!g198) & (g1695) & (!g1696) & (g1707) & (g1720)) + ((g174) & (!g198) & (g1695) & (g1696) & (!g1707) & (g1720)) + ((g174) & (!g198) & (g1695) & (g1696) & (g1707) & (!g1720)) + ((g174) & (!g198) & (g1695) & (g1696) & (g1707) & (g1720)) + ((g174) & (g198) & (!g1695) & (!g1696) & (!g1707) & (!g1720)) + ((g174) & (g198) & (g1695) & (!g1696) & (!g1707) & (g1720)) + ((g174) & (g198) & (g1695) & (!g1696) & (g1707) & (!g1720)) + ((g174) & (g198) & (g1695) & (!g1696) & (g1707) & (g1720)) + ((g174) & (g198) & (g1695) & (g1696) & (!g1707) & (!g1720)) + ((g174) & (g198) & (g1695) & (g1696) & (!g1707) & (g1720)) + ((g174) & (g198) & (g1695) & (g1696) & (g1707) & (!g1720)) + ((g174) & (g198) & (g1695) & (g1696) & (g1707) & (g1720)));
	assign g1771 = (((!g198) & (!g1696) & (g1707) & (!g1720)) + ((!g198) & (g1696) & (!g1707) & (!g1720)) + ((!g198) & (g1696) & (!g1707) & (g1720)) + ((!g198) & (g1696) & (g1707) & (g1720)) + ((g198) & (!g1696) & (!g1707) & (!g1720)) + ((g198) & (g1696) & (!g1707) & (g1720)) + ((g198) & (g1696) & (g1707) & (!g1720)) + ((g198) & (g1696) & (g1707) & (g1720)));
	assign g1772 = (((!g229) & (!g255) & (!g1698) & (g1699) & (g1706) & (!g1720)) + ((!g229) & (!g255) & (g1698) & (!g1699) & (!g1706) & (!g1720)) + ((!g229) & (!g255) & (g1698) & (!g1699) & (!g1706) & (g1720)) + ((!g229) & (!g255) & (g1698) & (!g1699) & (g1706) & (!g1720)) + ((!g229) & (!g255) & (g1698) & (!g1699) & (g1706) & (g1720)) + ((!g229) & (!g255) & (g1698) & (g1699) & (!g1706) & (!g1720)) + ((!g229) & (!g255) & (g1698) & (g1699) & (!g1706) & (g1720)) + ((!g229) & (!g255) & (g1698) & (g1699) & (g1706) & (g1720)) + ((!g229) & (g255) & (!g1698) & (!g1699) & (g1706) & (!g1720)) + ((!g229) & (g255) & (!g1698) & (g1699) & (!g1706) & (!g1720)) + ((!g229) & (g255) & (!g1698) & (g1699) & (g1706) & (!g1720)) + ((!g229) & (g255) & (g1698) & (!g1699) & (!g1706) & (!g1720)) + ((!g229) & (g255) & (g1698) & (!g1699) & (!g1706) & (g1720)) + ((!g229) & (g255) & (g1698) & (!g1699) & (g1706) & (g1720)) + ((!g229) & (g255) & (g1698) & (g1699) & (!g1706) & (g1720)) + ((!g229) & (g255) & (g1698) & (g1699) & (g1706) & (g1720)) + ((g229) & (!g255) & (!g1698) & (!g1699) & (!g1706) & (!g1720)) + ((g229) & (!g255) & (!g1698) & (!g1699) & (g1706) & (!g1720)) + ((g229) & (!g255) & (!g1698) & (g1699) & (!g1706) & (!g1720)) + ((g229) & (!g255) & (g1698) & (!g1699) & (!g1706) & (g1720)) + ((g229) & (!g255) & (g1698) & (!g1699) & (g1706) & (g1720)) + ((g229) & (!g255) & (g1698) & (g1699) & (!g1706) & (g1720)) + ((g229) & (!g255) & (g1698) & (g1699) & (g1706) & (!g1720)) + ((g229) & (!g255) & (g1698) & (g1699) & (g1706) & (g1720)) + ((g229) & (g255) & (!g1698) & (!g1699) & (!g1706) & (!g1720)) + ((g229) & (g255) & (g1698) & (!g1699) & (!g1706) & (g1720)) + ((g229) & (g255) & (g1698) & (!g1699) & (g1706) & (!g1720)) + ((g229) & (g255) & (g1698) & (!g1699) & (g1706) & (g1720)) + ((g229) & (g255) & (g1698) & (g1699) & (!g1706) & (!g1720)) + ((g229) & (g255) & (g1698) & (g1699) & (!g1706) & (g1720)) + ((g229) & (g255) & (g1698) & (g1699) & (g1706) & (!g1720)) + ((g229) & (g255) & (g1698) & (g1699) & (g1706) & (g1720)));
	assign g1773 = (((!g255) & (!g1699) & (g1706) & (!g1720)) + ((!g255) & (g1699) & (!g1706) & (!g1720)) + ((!g255) & (g1699) & (!g1706) & (g1720)) + ((!g255) & (g1699) & (g1706) & (g1720)) + ((g255) & (!g1699) & (!g1706) & (!g1720)) + ((g255) & (g1699) & (!g1706) & (g1720)) + ((g255) & (g1699) & (g1706) & (!g1720)) + ((g255) & (g1699) & (g1706) & (g1720)));
	assign g1774 = (((!g290) & (!g319) & (!g1701) & (g1702) & (g1705) & (!g1720)) + ((!g290) & (!g319) & (g1701) & (!g1702) & (!g1705) & (!g1720)) + ((!g290) & (!g319) & (g1701) & (!g1702) & (!g1705) & (g1720)) + ((!g290) & (!g319) & (g1701) & (!g1702) & (g1705) & (!g1720)) + ((!g290) & (!g319) & (g1701) & (!g1702) & (g1705) & (g1720)) + ((!g290) & (!g319) & (g1701) & (g1702) & (!g1705) & (!g1720)) + ((!g290) & (!g319) & (g1701) & (g1702) & (!g1705) & (g1720)) + ((!g290) & (!g319) & (g1701) & (g1702) & (g1705) & (g1720)) + ((!g290) & (g319) & (!g1701) & (!g1702) & (g1705) & (!g1720)) + ((!g290) & (g319) & (!g1701) & (g1702) & (!g1705) & (!g1720)) + ((!g290) & (g319) & (!g1701) & (g1702) & (g1705) & (!g1720)) + ((!g290) & (g319) & (g1701) & (!g1702) & (!g1705) & (!g1720)) + ((!g290) & (g319) & (g1701) & (!g1702) & (!g1705) & (g1720)) + ((!g290) & (g319) & (g1701) & (!g1702) & (g1705) & (g1720)) + ((!g290) & (g319) & (g1701) & (g1702) & (!g1705) & (g1720)) + ((!g290) & (g319) & (g1701) & (g1702) & (g1705) & (g1720)) + ((g290) & (!g319) & (!g1701) & (!g1702) & (!g1705) & (!g1720)) + ((g290) & (!g319) & (!g1701) & (!g1702) & (g1705) & (!g1720)) + ((g290) & (!g319) & (!g1701) & (g1702) & (!g1705) & (!g1720)) + ((g290) & (!g319) & (g1701) & (!g1702) & (!g1705) & (g1720)) + ((g290) & (!g319) & (g1701) & (!g1702) & (g1705) & (g1720)) + ((g290) & (!g319) & (g1701) & (g1702) & (!g1705) & (g1720)) + ((g290) & (!g319) & (g1701) & (g1702) & (g1705) & (!g1720)) + ((g290) & (!g319) & (g1701) & (g1702) & (g1705) & (g1720)) + ((g290) & (g319) & (!g1701) & (!g1702) & (!g1705) & (!g1720)) + ((g290) & (g319) & (g1701) & (!g1702) & (!g1705) & (g1720)) + ((g290) & (g319) & (g1701) & (!g1702) & (g1705) & (!g1720)) + ((g290) & (g319) & (g1701) & (!g1702) & (g1705) & (g1720)) + ((g290) & (g319) & (g1701) & (g1702) & (!g1705) & (!g1720)) + ((g290) & (g319) & (g1701) & (g1702) & (!g1705) & (g1720)) + ((g290) & (g319) & (g1701) & (g1702) & (g1705) & (!g1720)) + ((g290) & (g319) & (g1701) & (g1702) & (g1705) & (g1720)));
	assign g1775 = (((!g319) & (!g1702) & (g1705) & (!g1720)) + ((!g319) & (g1702) & (!g1705) & (!g1720)) + ((!g319) & (g1702) & (!g1705) & (g1720)) + ((!g319) & (g1702) & (g1705) & (g1720)) + ((g319) & (!g1702) & (!g1705) & (!g1720)) + ((g319) & (g1702) & (!g1705) & (g1720)) + ((g319) & (g1702) & (g1705) & (!g1720)) + ((g319) & (g1702) & (g1705) & (g1720)));
	assign g1776 = (((!g358) & (!g390) & (!g1704) & (g1634) & (g1676) & (!g1720)) + ((!g358) & (!g390) & (g1704) & (!g1634) & (!g1676) & (!g1720)) + ((!g358) & (!g390) & (g1704) & (!g1634) & (!g1676) & (g1720)) + ((!g358) & (!g390) & (g1704) & (!g1634) & (g1676) & (!g1720)) + ((!g358) & (!g390) & (g1704) & (!g1634) & (g1676) & (g1720)) + ((!g358) & (!g390) & (g1704) & (g1634) & (!g1676) & (!g1720)) + ((!g358) & (!g390) & (g1704) & (g1634) & (!g1676) & (g1720)) + ((!g358) & (!g390) & (g1704) & (g1634) & (g1676) & (g1720)) + ((!g358) & (g390) & (!g1704) & (!g1634) & (g1676) & (!g1720)) + ((!g358) & (g390) & (!g1704) & (g1634) & (!g1676) & (!g1720)) + ((!g358) & (g390) & (!g1704) & (g1634) & (g1676) & (!g1720)) + ((!g358) & (g390) & (g1704) & (!g1634) & (!g1676) & (!g1720)) + ((!g358) & (g390) & (g1704) & (!g1634) & (!g1676) & (g1720)) + ((!g358) & (g390) & (g1704) & (!g1634) & (g1676) & (g1720)) + ((!g358) & (g390) & (g1704) & (g1634) & (!g1676) & (g1720)) + ((!g358) & (g390) & (g1704) & (g1634) & (g1676) & (g1720)) + ((g358) & (!g390) & (!g1704) & (!g1634) & (!g1676) & (!g1720)) + ((g358) & (!g390) & (!g1704) & (!g1634) & (g1676) & (!g1720)) + ((g358) & (!g390) & (!g1704) & (g1634) & (!g1676) & (!g1720)) + ((g358) & (!g390) & (g1704) & (!g1634) & (!g1676) & (g1720)) + ((g358) & (!g390) & (g1704) & (!g1634) & (g1676) & (g1720)) + ((g358) & (!g390) & (g1704) & (g1634) & (!g1676) & (g1720)) + ((g358) & (!g390) & (g1704) & (g1634) & (g1676) & (!g1720)) + ((g358) & (!g390) & (g1704) & (g1634) & (g1676) & (g1720)) + ((g358) & (g390) & (!g1704) & (!g1634) & (!g1676) & (!g1720)) + ((g358) & (g390) & (g1704) & (!g1634) & (!g1676) & (g1720)) + ((g358) & (g390) & (g1704) & (!g1634) & (g1676) & (!g1720)) + ((g358) & (g390) & (g1704) & (!g1634) & (g1676) & (g1720)) + ((g358) & (g390) & (g1704) & (g1634) & (!g1676) & (!g1720)) + ((g358) & (g390) & (g1704) & (g1634) & (!g1676) & (g1720)) + ((g358) & (g390) & (g1704) & (g1634) & (g1676) & (!g1720)) + ((g358) & (g390) & (g1704) & (g1634) & (g1676) & (g1720)));
	assign g1777 = (((!g319) & (!g358) & (g1776) & (g1721) & (g1757)) + ((!g319) & (g358) & (g1776) & (!g1721) & (g1757)) + ((!g319) & (g358) & (g1776) & (g1721) & (!g1757)) + ((!g319) & (g358) & (g1776) & (g1721) & (g1757)) + ((g319) & (!g358) & (!g1776) & (g1721) & (g1757)) + ((g319) & (!g358) & (g1776) & (!g1721) & (!g1757)) + ((g319) & (!g358) & (g1776) & (!g1721) & (g1757)) + ((g319) & (!g358) & (g1776) & (g1721) & (!g1757)) + ((g319) & (!g358) & (g1776) & (g1721) & (g1757)) + ((g319) & (g358) & (!g1776) & (!g1721) & (g1757)) + ((g319) & (g358) & (!g1776) & (g1721) & (!g1757)) + ((g319) & (g358) & (!g1776) & (g1721) & (g1757)) + ((g319) & (g358) & (g1776) & (!g1721) & (!g1757)) + ((g319) & (g358) & (g1776) & (!g1721) & (g1757)) + ((g319) & (g358) & (g1776) & (g1721) & (!g1757)) + ((g319) & (g358) & (g1776) & (g1721) & (g1757)));
	assign g1778 = (((!g255) & (!g290) & (g1774) & (g1775) & (g1777)) + ((!g255) & (g290) & (g1774) & (!g1775) & (g1777)) + ((!g255) & (g290) & (g1774) & (g1775) & (!g1777)) + ((!g255) & (g290) & (g1774) & (g1775) & (g1777)) + ((g255) & (!g290) & (!g1774) & (g1775) & (g1777)) + ((g255) & (!g290) & (g1774) & (!g1775) & (!g1777)) + ((g255) & (!g290) & (g1774) & (!g1775) & (g1777)) + ((g255) & (!g290) & (g1774) & (g1775) & (!g1777)) + ((g255) & (!g290) & (g1774) & (g1775) & (g1777)) + ((g255) & (g290) & (!g1774) & (!g1775) & (g1777)) + ((g255) & (g290) & (!g1774) & (g1775) & (!g1777)) + ((g255) & (g290) & (!g1774) & (g1775) & (g1777)) + ((g255) & (g290) & (g1774) & (!g1775) & (!g1777)) + ((g255) & (g290) & (g1774) & (!g1775) & (g1777)) + ((g255) & (g290) & (g1774) & (g1775) & (!g1777)) + ((g255) & (g290) & (g1774) & (g1775) & (g1777)));
	assign g1779 = (((!g198) & (!g229) & (g1772) & (g1773) & (g1778)) + ((!g198) & (g229) & (g1772) & (!g1773) & (g1778)) + ((!g198) & (g229) & (g1772) & (g1773) & (!g1778)) + ((!g198) & (g229) & (g1772) & (g1773) & (g1778)) + ((g198) & (!g229) & (!g1772) & (g1773) & (g1778)) + ((g198) & (!g229) & (g1772) & (!g1773) & (!g1778)) + ((g198) & (!g229) & (g1772) & (!g1773) & (g1778)) + ((g198) & (!g229) & (g1772) & (g1773) & (!g1778)) + ((g198) & (!g229) & (g1772) & (g1773) & (g1778)) + ((g198) & (g229) & (!g1772) & (!g1773) & (g1778)) + ((g198) & (g229) & (!g1772) & (g1773) & (!g1778)) + ((g198) & (g229) & (!g1772) & (g1773) & (g1778)) + ((g198) & (g229) & (g1772) & (!g1773) & (!g1778)) + ((g198) & (g229) & (g1772) & (!g1773) & (g1778)) + ((g198) & (g229) & (g1772) & (g1773) & (!g1778)) + ((g198) & (g229) & (g1772) & (g1773) & (g1778)));
	assign g1780 = (((!g147) & (!g174) & (g1770) & (g1771) & (g1779)) + ((!g147) & (g174) & (g1770) & (!g1771) & (g1779)) + ((!g147) & (g174) & (g1770) & (g1771) & (!g1779)) + ((!g147) & (g174) & (g1770) & (g1771) & (g1779)) + ((g147) & (!g174) & (!g1770) & (g1771) & (g1779)) + ((g147) & (!g174) & (g1770) & (!g1771) & (!g1779)) + ((g147) & (!g174) & (g1770) & (!g1771) & (g1779)) + ((g147) & (!g174) & (g1770) & (g1771) & (!g1779)) + ((g147) & (!g174) & (g1770) & (g1771) & (g1779)) + ((g147) & (g174) & (!g1770) & (!g1771) & (g1779)) + ((g147) & (g174) & (!g1770) & (g1771) & (!g1779)) + ((g147) & (g174) & (!g1770) & (g1771) & (g1779)) + ((g147) & (g174) & (g1770) & (!g1771) & (!g1779)) + ((g147) & (g174) & (g1770) & (!g1771) & (g1779)) + ((g147) & (g174) & (g1770) & (g1771) & (!g1779)) + ((g147) & (g174) & (g1770) & (g1771) & (g1779)));
	assign g1781 = (((!g104) & (!g127) & (g1768) & (g1769) & (g1780)) + ((!g104) & (g127) & (g1768) & (!g1769) & (g1780)) + ((!g104) & (g127) & (g1768) & (g1769) & (!g1780)) + ((!g104) & (g127) & (g1768) & (g1769) & (g1780)) + ((g104) & (!g127) & (!g1768) & (g1769) & (g1780)) + ((g104) & (!g127) & (g1768) & (!g1769) & (!g1780)) + ((g104) & (!g127) & (g1768) & (!g1769) & (g1780)) + ((g104) & (!g127) & (g1768) & (g1769) & (!g1780)) + ((g104) & (!g127) & (g1768) & (g1769) & (g1780)) + ((g104) & (g127) & (!g1768) & (!g1769) & (g1780)) + ((g104) & (g127) & (!g1768) & (g1769) & (!g1780)) + ((g104) & (g127) & (!g1768) & (g1769) & (g1780)) + ((g104) & (g127) & (g1768) & (!g1769) & (!g1780)) + ((g104) & (g127) & (g1768) & (!g1769) & (g1780)) + ((g104) & (g127) & (g1768) & (g1769) & (!g1780)) + ((g104) & (g127) & (g1768) & (g1769) & (g1780)));
	assign g1782 = (((!g68) & (!g87) & (g1766) & (g1767) & (g1781)) + ((!g68) & (g87) & (g1766) & (!g1767) & (g1781)) + ((!g68) & (g87) & (g1766) & (g1767) & (!g1781)) + ((!g68) & (g87) & (g1766) & (g1767) & (g1781)) + ((g68) & (!g87) & (!g1766) & (g1767) & (g1781)) + ((g68) & (!g87) & (g1766) & (!g1767) & (!g1781)) + ((g68) & (!g87) & (g1766) & (!g1767) & (g1781)) + ((g68) & (!g87) & (g1766) & (g1767) & (!g1781)) + ((g68) & (!g87) & (g1766) & (g1767) & (g1781)) + ((g68) & (g87) & (!g1766) & (!g1767) & (g1781)) + ((g68) & (g87) & (!g1766) & (g1767) & (!g1781)) + ((g68) & (g87) & (!g1766) & (g1767) & (g1781)) + ((g68) & (g87) & (g1766) & (!g1767) & (!g1781)) + ((g68) & (g87) & (g1766) & (!g1767) & (g1781)) + ((g68) & (g87) & (g1766) & (g1767) & (!g1781)) + ((g68) & (g87) & (g1766) & (g1767) & (g1781)));
	assign g1783 = (((!g39) & (!g54) & (g1764) & (g1765) & (g1782)) + ((!g39) & (g54) & (g1764) & (!g1765) & (g1782)) + ((!g39) & (g54) & (g1764) & (g1765) & (!g1782)) + ((!g39) & (g54) & (g1764) & (g1765) & (g1782)) + ((g39) & (!g54) & (!g1764) & (g1765) & (g1782)) + ((g39) & (!g54) & (g1764) & (!g1765) & (!g1782)) + ((g39) & (!g54) & (g1764) & (!g1765) & (g1782)) + ((g39) & (!g54) & (g1764) & (g1765) & (!g1782)) + ((g39) & (!g54) & (g1764) & (g1765) & (g1782)) + ((g39) & (g54) & (!g1764) & (!g1765) & (g1782)) + ((g39) & (g54) & (!g1764) & (g1765) & (!g1782)) + ((g39) & (g54) & (!g1764) & (g1765) & (g1782)) + ((g39) & (g54) & (g1764) & (!g1765) & (!g1782)) + ((g39) & (g54) & (g1764) & (!g1765) & (g1782)) + ((g39) & (g54) & (g1764) & (g1765) & (!g1782)) + ((g39) & (g54) & (g1764) & (g1765) & (g1782)));
	assign g1784 = (((!g18) & (!g27) & (g1762) & (g1763) & (g1783)) + ((!g18) & (g27) & (g1762) & (!g1763) & (g1783)) + ((!g18) & (g27) & (g1762) & (g1763) & (!g1783)) + ((!g18) & (g27) & (g1762) & (g1763) & (g1783)) + ((g18) & (!g27) & (!g1762) & (g1763) & (g1783)) + ((g18) & (!g27) & (g1762) & (!g1763) & (!g1783)) + ((g18) & (!g27) & (g1762) & (!g1763) & (g1783)) + ((g18) & (!g27) & (g1762) & (g1763) & (!g1783)) + ((g18) & (!g27) & (g1762) & (g1763) & (g1783)) + ((g18) & (g27) & (!g1762) & (!g1763) & (g1783)) + ((g18) & (g27) & (!g1762) & (g1763) & (!g1783)) + ((g18) & (g27) & (!g1762) & (g1763) & (g1783)) + ((g18) & (g27) & (g1762) & (!g1763) & (!g1783)) + ((g18) & (g27) & (g1762) & (!g1763) & (g1783)) + ((g18) & (g27) & (g1762) & (g1763) & (!g1783)) + ((g18) & (g27) & (g1762) & (g1763) & (g1783)));
	assign g1785 = (((!g2) & (!g8) & (g1760) & (g1761) & (g1784)) + ((!g2) & (g8) & (g1760) & (!g1761) & (g1784)) + ((!g2) & (g8) & (g1760) & (g1761) & (!g1784)) + ((!g2) & (g8) & (g1760) & (g1761) & (g1784)) + ((g2) & (!g8) & (!g1760) & (g1761) & (g1784)) + ((g2) & (!g8) & (g1760) & (!g1761) & (!g1784)) + ((g2) & (!g8) & (g1760) & (!g1761) & (g1784)) + ((g2) & (!g8) & (g1760) & (g1761) & (!g1784)) + ((g2) & (!g8) & (g1760) & (g1761) & (g1784)) + ((g2) & (g8) & (!g1760) & (!g1761) & (g1784)) + ((g2) & (g8) & (!g1760) & (g1761) & (!g1784)) + ((g2) & (g8) & (!g1760) & (g1761) & (g1784)) + ((g2) & (g8) & (g1760) & (!g1761) & (!g1784)) + ((g2) & (g8) & (g1760) & (!g1761) & (g1784)) + ((g2) & (g8) & (g1760) & (g1761) & (!g1784)) + ((g2) & (g8) & (g1760) & (g1761) & (g1784)));
	assign g1786 = (((!g2) & (!g1678) & (g1713) & (!g1720)) + ((!g2) & (g1678) & (!g1713) & (!g1720)) + ((!g2) & (g1678) & (!g1713) & (g1720)) + ((!g2) & (g1678) & (g1713) & (g1720)) + ((g2) & (!g1678) & (!g1713) & (!g1720)) + ((g2) & (g1678) & (!g1713) & (g1720)) + ((g2) & (g1678) & (g1713) & (!g1720)) + ((g2) & (g1678) & (g1713) & (g1720)));
	assign g1787 = (((!g1) & (!g1677) & (!g1716) & (!g1718) & (g1719)) + ((!g1) & (!g1677) & (!g1716) & (g1718) & (!g1719)) + ((!g1) & (!g1677) & (!g1716) & (g1718) & (g1719)) + ((!g1) & (g1677) & (g1716) & (!g1718) & (!g1719)) + ((!g1) & (g1677) & (g1716) & (!g1718) & (g1719)) + ((!g1) & (g1677) & (g1716) & (g1718) & (!g1719)) + ((!g1) & (g1677) & (g1716) & (g1718) & (g1719)) + ((g1) & (!g1677) & (!g1716) & (!g1718) & (g1719)) + ((g1) & (!g1677) & (!g1716) & (g1718) & (g1719)) + ((g1) & (g1677) & (g1716) & (!g1718) & (!g1719)) + ((g1) & (g1677) & (g1716) & (!g1718) & (g1719)) + ((g1) & (g1677) & (g1716) & (g1718) & (!g1719)) + ((g1) & (g1677) & (g1716) & (g1718) & (g1719)));
	assign g1788 = (((!g4) & (!g1) & (!g1759) & (!g1785) & (!g1786) & (!g1787)) + ((!g4) & (g1) & (!g1759) & (!g1785) & (!g1786) & (!g1787)) + ((!g4) & (g1) & (!g1759) & (!g1785) & (!g1786) & (g1787)) + ((!g4) & (g1) & (!g1759) & (!g1785) & (g1786) & (!g1787)) + ((!g4) & (g1) & (!g1759) & (!g1785) & (g1786) & (g1787)) + ((!g4) & (g1) & (!g1759) & (g1785) & (!g1786) & (!g1787)) + ((!g4) & (g1) & (!g1759) & (g1785) & (!g1786) & (g1787)) + ((!g4) & (g1) & (!g1759) & (g1785) & (g1786) & (!g1787)) + ((!g4) & (g1) & (!g1759) & (g1785) & (g1786) & (g1787)) + ((!g4) & (g1) & (g1759) & (!g1785) & (!g1786) & (!g1787)) + ((!g4) & (g1) & (g1759) & (!g1785) & (!g1786) & (g1787)) + ((g4) & (!g1) & (!g1759) & (!g1785) & (!g1786) & (!g1787)) + ((g4) & (!g1) & (!g1759) & (!g1785) & (g1786) & (!g1787)) + ((g4) & (!g1) & (!g1759) & (g1785) & (!g1786) & (!g1787)) + ((g4) & (g1) & (!g1759) & (!g1785) & (!g1786) & (!g1787)) + ((g4) & (g1) & (!g1759) & (!g1785) & (!g1786) & (g1787)) + ((g4) & (g1) & (!g1759) & (!g1785) & (g1786) & (!g1787)) + ((g4) & (g1) & (!g1759) & (!g1785) & (g1786) & (g1787)) + ((g4) & (g1) & (!g1759) & (g1785) & (!g1786) & (!g1787)) + ((g4) & (g1) & (!g1759) & (g1785) & (!g1786) & (g1787)) + ((g4) & (g1) & (!g1759) & (g1785) & (g1786) & (!g1787)) + ((g4) & (g1) & (!g1759) & (g1785) & (g1786) & (g1787)) + ((g4) & (g1) & (g1759) & (!g1785) & (!g1786) & (!g1787)) + ((g4) & (g1) & (g1759) & (!g1785) & (!g1786) & (g1787)) + ((g4) & (g1) & (g1759) & (!g1785) & (g1786) & (!g1787)) + ((g4) & (g1) & (g1759) & (!g1785) & (g1786) & (g1787)) + ((g4) & (g1) & (g1759) & (g1785) & (!g1786) & (!g1787)) + ((g4) & (g1) & (g1759) & (g1785) & (!g1786) & (g1787)));
	assign g1789 = (((!g358) & (!g1721) & (g1757) & (!g1758) & (!g1788)) + ((!g358) & (!g1721) & (g1757) & (g1758) & (!g1788)) + ((!g358) & (!g1721) & (g1757) & (g1758) & (g1788)) + ((!g358) & (g1721) & (!g1757) & (!g1758) & (!g1788)) + ((!g358) & (g1721) & (!g1757) & (!g1758) & (g1788)) + ((!g358) & (g1721) & (!g1757) & (g1758) & (!g1788)) + ((!g358) & (g1721) & (!g1757) & (g1758) & (g1788)) + ((!g358) & (g1721) & (g1757) & (!g1758) & (g1788)) + ((g358) & (!g1721) & (!g1757) & (!g1758) & (!g1788)) + ((g358) & (!g1721) & (!g1757) & (g1758) & (!g1788)) + ((g358) & (!g1721) & (!g1757) & (g1758) & (g1788)) + ((g358) & (g1721) & (!g1757) & (!g1758) & (g1788)) + ((g358) & (g1721) & (g1757) & (!g1758) & (!g1788)) + ((g358) & (g1721) & (g1757) & (!g1758) & (g1788)) + ((g358) & (g1721) & (g1757) & (g1758) & (!g1788)) + ((g358) & (g1721) & (g1757) & (g1758) & (g1788)));
	assign g1790 = (((!g390) & (!g433) & (g1723) & (g1756)) + ((!g390) & (g433) & (!g1723) & (g1756)) + ((!g390) & (g433) & (g1723) & (!g1756)) + ((!g390) & (g433) & (g1723) & (g1756)) + ((g390) & (!g433) & (!g1723) & (!g1756)) + ((g390) & (!g433) & (!g1723) & (g1756)) + ((g390) & (!g433) & (g1723) & (!g1756)) + ((g390) & (g433) & (!g1723) & (!g1756)));
	assign g1791 = (((!g1722) & (!g1758) & (!g1788) & (g1790)) + ((!g1722) & (g1758) & (!g1788) & (g1790)) + ((!g1722) & (g1758) & (g1788) & (g1790)) + ((g1722) & (!g1758) & (!g1788) & (!g1790)) + ((g1722) & (!g1758) & (g1788) & (!g1790)) + ((g1722) & (!g1758) & (g1788) & (g1790)) + ((g1722) & (g1758) & (!g1788) & (!g1790)) + ((g1722) & (g1758) & (g1788) & (!g1790)));
	assign g1792 = (((!g433) & (!g1723) & (g1756) & (!g1758) & (!g1788)) + ((!g433) & (!g1723) & (g1756) & (g1758) & (!g1788)) + ((!g433) & (!g1723) & (g1756) & (g1758) & (g1788)) + ((!g433) & (g1723) & (!g1756) & (!g1758) & (!g1788)) + ((!g433) & (g1723) & (!g1756) & (!g1758) & (g1788)) + ((!g433) & (g1723) & (!g1756) & (g1758) & (!g1788)) + ((!g433) & (g1723) & (!g1756) & (g1758) & (g1788)) + ((!g433) & (g1723) & (g1756) & (!g1758) & (g1788)) + ((g433) & (!g1723) & (!g1756) & (!g1758) & (!g1788)) + ((g433) & (!g1723) & (!g1756) & (g1758) & (!g1788)) + ((g433) & (!g1723) & (!g1756) & (g1758) & (g1788)) + ((g433) & (g1723) & (!g1756) & (!g1758) & (g1788)) + ((g433) & (g1723) & (g1756) & (!g1758) & (!g1788)) + ((g433) & (g1723) & (g1756) & (!g1758) & (g1788)) + ((g433) & (g1723) & (g1756) & (g1758) & (!g1788)) + ((g433) & (g1723) & (g1756) & (g1758) & (g1788)));
	assign g1793 = (((!g468) & (!g515) & (g1725) & (g1755)) + ((!g468) & (g515) & (!g1725) & (g1755)) + ((!g468) & (g515) & (g1725) & (!g1755)) + ((!g468) & (g515) & (g1725) & (g1755)) + ((g468) & (!g515) & (!g1725) & (!g1755)) + ((g468) & (!g515) & (!g1725) & (g1755)) + ((g468) & (!g515) & (g1725) & (!g1755)) + ((g468) & (g515) & (!g1725) & (!g1755)));
	assign g1794 = (((!g1724) & (!g1758) & (!g1788) & (g1793)) + ((!g1724) & (g1758) & (!g1788) & (g1793)) + ((!g1724) & (g1758) & (g1788) & (g1793)) + ((g1724) & (!g1758) & (!g1788) & (!g1793)) + ((g1724) & (!g1758) & (g1788) & (!g1793)) + ((g1724) & (!g1758) & (g1788) & (g1793)) + ((g1724) & (g1758) & (!g1788) & (!g1793)) + ((g1724) & (g1758) & (g1788) & (!g1793)));
	assign g1795 = (((!g515) & (!g1725) & (g1755) & (!g1758) & (!g1788)) + ((!g515) & (!g1725) & (g1755) & (g1758) & (!g1788)) + ((!g515) & (!g1725) & (g1755) & (g1758) & (g1788)) + ((!g515) & (g1725) & (!g1755) & (!g1758) & (!g1788)) + ((!g515) & (g1725) & (!g1755) & (!g1758) & (g1788)) + ((!g515) & (g1725) & (!g1755) & (g1758) & (!g1788)) + ((!g515) & (g1725) & (!g1755) & (g1758) & (g1788)) + ((!g515) & (g1725) & (g1755) & (!g1758) & (g1788)) + ((g515) & (!g1725) & (!g1755) & (!g1758) & (!g1788)) + ((g515) & (!g1725) & (!g1755) & (g1758) & (!g1788)) + ((g515) & (!g1725) & (!g1755) & (g1758) & (g1788)) + ((g515) & (g1725) & (!g1755) & (!g1758) & (g1788)) + ((g515) & (g1725) & (g1755) & (!g1758) & (!g1788)) + ((g515) & (g1725) & (g1755) & (!g1758) & (g1788)) + ((g515) & (g1725) & (g1755) & (g1758) & (!g1788)) + ((g515) & (g1725) & (g1755) & (g1758) & (g1788)));
	assign g1796 = (((!g553) & (!g604) & (g1727) & (g1754)) + ((!g553) & (g604) & (!g1727) & (g1754)) + ((!g553) & (g604) & (g1727) & (!g1754)) + ((!g553) & (g604) & (g1727) & (g1754)) + ((g553) & (!g604) & (!g1727) & (!g1754)) + ((g553) & (!g604) & (!g1727) & (g1754)) + ((g553) & (!g604) & (g1727) & (!g1754)) + ((g553) & (g604) & (!g1727) & (!g1754)));
	assign g1797 = (((!g1726) & (!g1758) & (!g1788) & (g1796)) + ((!g1726) & (g1758) & (!g1788) & (g1796)) + ((!g1726) & (g1758) & (g1788) & (g1796)) + ((g1726) & (!g1758) & (!g1788) & (!g1796)) + ((g1726) & (!g1758) & (g1788) & (!g1796)) + ((g1726) & (!g1758) & (g1788) & (g1796)) + ((g1726) & (g1758) & (!g1788) & (!g1796)) + ((g1726) & (g1758) & (g1788) & (!g1796)));
	assign g1798 = (((!g604) & (!g1727) & (g1754) & (!g1758) & (!g1788)) + ((!g604) & (!g1727) & (g1754) & (g1758) & (!g1788)) + ((!g604) & (!g1727) & (g1754) & (g1758) & (g1788)) + ((!g604) & (g1727) & (!g1754) & (!g1758) & (!g1788)) + ((!g604) & (g1727) & (!g1754) & (!g1758) & (g1788)) + ((!g604) & (g1727) & (!g1754) & (g1758) & (!g1788)) + ((!g604) & (g1727) & (!g1754) & (g1758) & (g1788)) + ((!g604) & (g1727) & (g1754) & (!g1758) & (g1788)) + ((g604) & (!g1727) & (!g1754) & (!g1758) & (!g1788)) + ((g604) & (!g1727) & (!g1754) & (g1758) & (!g1788)) + ((g604) & (!g1727) & (!g1754) & (g1758) & (g1788)) + ((g604) & (g1727) & (!g1754) & (!g1758) & (g1788)) + ((g604) & (g1727) & (g1754) & (!g1758) & (!g1788)) + ((g604) & (g1727) & (g1754) & (!g1758) & (g1788)) + ((g604) & (g1727) & (g1754) & (g1758) & (!g1788)) + ((g604) & (g1727) & (g1754) & (g1758) & (g1788)));
	assign g1799 = (((!g645) & (!g700) & (g1729) & (g1753)) + ((!g645) & (g700) & (!g1729) & (g1753)) + ((!g645) & (g700) & (g1729) & (!g1753)) + ((!g645) & (g700) & (g1729) & (g1753)) + ((g645) & (!g700) & (!g1729) & (!g1753)) + ((g645) & (!g700) & (!g1729) & (g1753)) + ((g645) & (!g700) & (g1729) & (!g1753)) + ((g645) & (g700) & (!g1729) & (!g1753)));
	assign g1800 = (((!g1728) & (!g1758) & (!g1788) & (g1799)) + ((!g1728) & (g1758) & (!g1788) & (g1799)) + ((!g1728) & (g1758) & (g1788) & (g1799)) + ((g1728) & (!g1758) & (!g1788) & (!g1799)) + ((g1728) & (!g1758) & (g1788) & (!g1799)) + ((g1728) & (!g1758) & (g1788) & (g1799)) + ((g1728) & (g1758) & (!g1788) & (!g1799)) + ((g1728) & (g1758) & (g1788) & (!g1799)));
	assign g1801 = (((!g700) & (!g1729) & (g1753) & (!g1758) & (!g1788)) + ((!g700) & (!g1729) & (g1753) & (g1758) & (!g1788)) + ((!g700) & (!g1729) & (g1753) & (g1758) & (g1788)) + ((!g700) & (g1729) & (!g1753) & (!g1758) & (!g1788)) + ((!g700) & (g1729) & (!g1753) & (!g1758) & (g1788)) + ((!g700) & (g1729) & (!g1753) & (g1758) & (!g1788)) + ((!g700) & (g1729) & (!g1753) & (g1758) & (g1788)) + ((!g700) & (g1729) & (g1753) & (!g1758) & (g1788)) + ((g700) & (!g1729) & (!g1753) & (!g1758) & (!g1788)) + ((g700) & (!g1729) & (!g1753) & (g1758) & (!g1788)) + ((g700) & (!g1729) & (!g1753) & (g1758) & (g1788)) + ((g700) & (g1729) & (!g1753) & (!g1758) & (g1788)) + ((g700) & (g1729) & (g1753) & (!g1758) & (!g1788)) + ((g700) & (g1729) & (g1753) & (!g1758) & (g1788)) + ((g700) & (g1729) & (g1753) & (g1758) & (!g1788)) + ((g700) & (g1729) & (g1753) & (g1758) & (g1788)));
	assign g1802 = (((!g744) & (!g803) & (g1731) & (g1752)) + ((!g744) & (g803) & (!g1731) & (g1752)) + ((!g744) & (g803) & (g1731) & (!g1752)) + ((!g744) & (g803) & (g1731) & (g1752)) + ((g744) & (!g803) & (!g1731) & (!g1752)) + ((g744) & (!g803) & (!g1731) & (g1752)) + ((g744) & (!g803) & (g1731) & (!g1752)) + ((g744) & (g803) & (!g1731) & (!g1752)));
	assign g1803 = (((!g1730) & (!g1758) & (!g1788) & (g1802)) + ((!g1730) & (g1758) & (!g1788) & (g1802)) + ((!g1730) & (g1758) & (g1788) & (g1802)) + ((g1730) & (!g1758) & (!g1788) & (!g1802)) + ((g1730) & (!g1758) & (g1788) & (!g1802)) + ((g1730) & (!g1758) & (g1788) & (g1802)) + ((g1730) & (g1758) & (!g1788) & (!g1802)) + ((g1730) & (g1758) & (g1788) & (!g1802)));
	assign g1804 = (((!g803) & (!g1731) & (g1752) & (!g1758) & (!g1788)) + ((!g803) & (!g1731) & (g1752) & (g1758) & (!g1788)) + ((!g803) & (!g1731) & (g1752) & (g1758) & (g1788)) + ((!g803) & (g1731) & (!g1752) & (!g1758) & (!g1788)) + ((!g803) & (g1731) & (!g1752) & (!g1758) & (g1788)) + ((!g803) & (g1731) & (!g1752) & (g1758) & (!g1788)) + ((!g803) & (g1731) & (!g1752) & (g1758) & (g1788)) + ((!g803) & (g1731) & (g1752) & (!g1758) & (g1788)) + ((g803) & (!g1731) & (!g1752) & (!g1758) & (!g1788)) + ((g803) & (!g1731) & (!g1752) & (g1758) & (!g1788)) + ((g803) & (!g1731) & (!g1752) & (g1758) & (g1788)) + ((g803) & (g1731) & (!g1752) & (!g1758) & (g1788)) + ((g803) & (g1731) & (g1752) & (!g1758) & (!g1788)) + ((g803) & (g1731) & (g1752) & (!g1758) & (g1788)) + ((g803) & (g1731) & (g1752) & (g1758) & (!g1788)) + ((g803) & (g1731) & (g1752) & (g1758) & (g1788)));
	assign g1805 = (((!g851) & (!g914) & (g1733) & (g1751)) + ((!g851) & (g914) & (!g1733) & (g1751)) + ((!g851) & (g914) & (g1733) & (!g1751)) + ((!g851) & (g914) & (g1733) & (g1751)) + ((g851) & (!g914) & (!g1733) & (!g1751)) + ((g851) & (!g914) & (!g1733) & (g1751)) + ((g851) & (!g914) & (g1733) & (!g1751)) + ((g851) & (g914) & (!g1733) & (!g1751)));
	assign g1806 = (((!g1732) & (!g1758) & (!g1788) & (g1805)) + ((!g1732) & (g1758) & (!g1788) & (g1805)) + ((!g1732) & (g1758) & (g1788) & (g1805)) + ((g1732) & (!g1758) & (!g1788) & (!g1805)) + ((g1732) & (!g1758) & (g1788) & (!g1805)) + ((g1732) & (!g1758) & (g1788) & (g1805)) + ((g1732) & (g1758) & (!g1788) & (!g1805)) + ((g1732) & (g1758) & (g1788) & (!g1805)));
	assign g1807 = (((!g914) & (!g1733) & (g1751) & (!g1758) & (!g1788)) + ((!g914) & (!g1733) & (g1751) & (g1758) & (!g1788)) + ((!g914) & (!g1733) & (g1751) & (g1758) & (g1788)) + ((!g914) & (g1733) & (!g1751) & (!g1758) & (!g1788)) + ((!g914) & (g1733) & (!g1751) & (!g1758) & (g1788)) + ((!g914) & (g1733) & (!g1751) & (g1758) & (!g1788)) + ((!g914) & (g1733) & (!g1751) & (g1758) & (g1788)) + ((!g914) & (g1733) & (g1751) & (!g1758) & (g1788)) + ((g914) & (!g1733) & (!g1751) & (!g1758) & (!g1788)) + ((g914) & (!g1733) & (!g1751) & (g1758) & (!g1788)) + ((g914) & (!g1733) & (!g1751) & (g1758) & (g1788)) + ((g914) & (g1733) & (!g1751) & (!g1758) & (g1788)) + ((g914) & (g1733) & (g1751) & (!g1758) & (!g1788)) + ((g914) & (g1733) & (g1751) & (!g1758) & (g1788)) + ((g914) & (g1733) & (g1751) & (g1758) & (!g1788)) + ((g914) & (g1733) & (g1751) & (g1758) & (g1788)));
	assign g1808 = (((!g1032) & (!g1030) & (g1735) & (g1750)) + ((!g1032) & (g1030) & (!g1735) & (g1750)) + ((!g1032) & (g1030) & (g1735) & (!g1750)) + ((!g1032) & (g1030) & (g1735) & (g1750)) + ((g1032) & (!g1030) & (!g1735) & (!g1750)) + ((g1032) & (!g1030) & (!g1735) & (g1750)) + ((g1032) & (!g1030) & (g1735) & (!g1750)) + ((g1032) & (g1030) & (!g1735) & (!g1750)));
	assign g1809 = (((!g1734) & (!g1758) & (!g1788) & (g1808)) + ((!g1734) & (g1758) & (!g1788) & (g1808)) + ((!g1734) & (g1758) & (g1788) & (g1808)) + ((g1734) & (!g1758) & (!g1788) & (!g1808)) + ((g1734) & (!g1758) & (g1788) & (!g1808)) + ((g1734) & (!g1758) & (g1788) & (g1808)) + ((g1734) & (g1758) & (!g1788) & (!g1808)) + ((g1734) & (g1758) & (g1788) & (!g1808)));
	assign g1810 = (((!g1030) & (!g1735) & (g1750) & (!g1758) & (!g1788)) + ((!g1030) & (!g1735) & (g1750) & (g1758) & (!g1788)) + ((!g1030) & (!g1735) & (g1750) & (g1758) & (g1788)) + ((!g1030) & (g1735) & (!g1750) & (!g1758) & (!g1788)) + ((!g1030) & (g1735) & (!g1750) & (!g1758) & (g1788)) + ((!g1030) & (g1735) & (!g1750) & (g1758) & (!g1788)) + ((!g1030) & (g1735) & (!g1750) & (g1758) & (g1788)) + ((!g1030) & (g1735) & (g1750) & (!g1758) & (g1788)) + ((g1030) & (!g1735) & (!g1750) & (!g1758) & (!g1788)) + ((g1030) & (!g1735) & (!g1750) & (g1758) & (!g1788)) + ((g1030) & (!g1735) & (!g1750) & (g1758) & (g1788)) + ((g1030) & (g1735) & (!g1750) & (!g1758) & (g1788)) + ((g1030) & (g1735) & (g1750) & (!g1758) & (!g1788)) + ((g1030) & (g1735) & (g1750) & (!g1758) & (g1788)) + ((g1030) & (g1735) & (g1750) & (g1758) & (!g1788)) + ((g1030) & (g1735) & (g1750) & (g1758) & (g1788)));
	assign g1811 = (((!g1160) & (!g1154) & (g1737) & (g1749)) + ((!g1160) & (g1154) & (!g1737) & (g1749)) + ((!g1160) & (g1154) & (g1737) & (!g1749)) + ((!g1160) & (g1154) & (g1737) & (g1749)) + ((g1160) & (!g1154) & (!g1737) & (!g1749)) + ((g1160) & (!g1154) & (!g1737) & (g1749)) + ((g1160) & (!g1154) & (g1737) & (!g1749)) + ((g1160) & (g1154) & (!g1737) & (!g1749)));
	assign g1812 = (((!g1736) & (!g1758) & (!g1788) & (g1811)) + ((!g1736) & (g1758) & (!g1788) & (g1811)) + ((!g1736) & (g1758) & (g1788) & (g1811)) + ((g1736) & (!g1758) & (!g1788) & (!g1811)) + ((g1736) & (!g1758) & (g1788) & (!g1811)) + ((g1736) & (!g1758) & (g1788) & (g1811)) + ((g1736) & (g1758) & (!g1788) & (!g1811)) + ((g1736) & (g1758) & (g1788) & (!g1811)));
	assign g1813 = (((!g1154) & (!g1737) & (g1749) & (!g1758) & (!g1788)) + ((!g1154) & (!g1737) & (g1749) & (g1758) & (!g1788)) + ((!g1154) & (!g1737) & (g1749) & (g1758) & (g1788)) + ((!g1154) & (g1737) & (!g1749) & (!g1758) & (!g1788)) + ((!g1154) & (g1737) & (!g1749) & (!g1758) & (g1788)) + ((!g1154) & (g1737) & (!g1749) & (g1758) & (!g1788)) + ((!g1154) & (g1737) & (!g1749) & (g1758) & (g1788)) + ((!g1154) & (g1737) & (g1749) & (!g1758) & (g1788)) + ((g1154) & (!g1737) & (!g1749) & (!g1758) & (!g1788)) + ((g1154) & (!g1737) & (!g1749) & (g1758) & (!g1788)) + ((g1154) & (!g1737) & (!g1749) & (g1758) & (g1788)) + ((g1154) & (g1737) & (!g1749) & (!g1758) & (g1788)) + ((g1154) & (g1737) & (g1749) & (!g1758) & (!g1788)) + ((g1154) & (g1737) & (g1749) & (!g1758) & (g1788)) + ((g1154) & (g1737) & (g1749) & (g1758) & (!g1788)) + ((g1154) & (g1737) & (g1749) & (g1758) & (g1788)));
	assign g1814 = (((!g1295) & (!g1285) & (g1739) & (g1748)) + ((!g1295) & (g1285) & (!g1739) & (g1748)) + ((!g1295) & (g1285) & (g1739) & (!g1748)) + ((!g1295) & (g1285) & (g1739) & (g1748)) + ((g1295) & (!g1285) & (!g1739) & (!g1748)) + ((g1295) & (!g1285) & (!g1739) & (g1748)) + ((g1295) & (!g1285) & (g1739) & (!g1748)) + ((g1295) & (g1285) & (!g1739) & (!g1748)));
	assign g1815 = (((!g1738) & (!g1758) & (!g1788) & (g1814)) + ((!g1738) & (g1758) & (!g1788) & (g1814)) + ((!g1738) & (g1758) & (g1788) & (g1814)) + ((g1738) & (!g1758) & (!g1788) & (!g1814)) + ((g1738) & (!g1758) & (g1788) & (!g1814)) + ((g1738) & (!g1758) & (g1788) & (g1814)) + ((g1738) & (g1758) & (!g1788) & (!g1814)) + ((g1738) & (g1758) & (g1788) & (!g1814)));
	assign g1816 = (((!g1285) & (!g1739) & (g1748) & (!g1758) & (!g1788)) + ((!g1285) & (!g1739) & (g1748) & (g1758) & (!g1788)) + ((!g1285) & (!g1739) & (g1748) & (g1758) & (g1788)) + ((!g1285) & (g1739) & (!g1748) & (!g1758) & (!g1788)) + ((!g1285) & (g1739) & (!g1748) & (!g1758) & (g1788)) + ((!g1285) & (g1739) & (!g1748) & (g1758) & (!g1788)) + ((!g1285) & (g1739) & (!g1748) & (g1758) & (g1788)) + ((!g1285) & (g1739) & (g1748) & (!g1758) & (g1788)) + ((g1285) & (!g1739) & (!g1748) & (!g1758) & (!g1788)) + ((g1285) & (!g1739) & (!g1748) & (g1758) & (!g1788)) + ((g1285) & (!g1739) & (!g1748) & (g1758) & (g1788)) + ((g1285) & (g1739) & (!g1748) & (!g1758) & (g1788)) + ((g1285) & (g1739) & (g1748) & (!g1758) & (!g1788)) + ((g1285) & (g1739) & (g1748) & (!g1758) & (g1788)) + ((g1285) & (g1739) & (g1748) & (g1758) & (!g1788)) + ((g1285) & (g1739) & (g1748) & (g1758) & (g1788)));
	assign g1817 = (((!g1437) & (!g1423) & (g1741) & (g1747)) + ((!g1437) & (g1423) & (!g1741) & (g1747)) + ((!g1437) & (g1423) & (g1741) & (!g1747)) + ((!g1437) & (g1423) & (g1741) & (g1747)) + ((g1437) & (!g1423) & (!g1741) & (!g1747)) + ((g1437) & (!g1423) & (!g1741) & (g1747)) + ((g1437) & (!g1423) & (g1741) & (!g1747)) + ((g1437) & (g1423) & (!g1741) & (!g1747)));
	assign g1818 = (((!g1740) & (!g1758) & (!g1788) & (g1817)) + ((!g1740) & (g1758) & (!g1788) & (g1817)) + ((!g1740) & (g1758) & (g1788) & (g1817)) + ((g1740) & (!g1758) & (!g1788) & (!g1817)) + ((g1740) & (!g1758) & (g1788) & (!g1817)) + ((g1740) & (!g1758) & (g1788) & (g1817)) + ((g1740) & (g1758) & (!g1788) & (!g1817)) + ((g1740) & (g1758) & (g1788) & (!g1817)));
	assign g1819 = (((!g1423) & (!g1741) & (g1747) & (!g1758) & (!g1788)) + ((!g1423) & (!g1741) & (g1747) & (g1758) & (!g1788)) + ((!g1423) & (!g1741) & (g1747) & (g1758) & (g1788)) + ((!g1423) & (g1741) & (!g1747) & (!g1758) & (!g1788)) + ((!g1423) & (g1741) & (!g1747) & (!g1758) & (g1788)) + ((!g1423) & (g1741) & (!g1747) & (g1758) & (!g1788)) + ((!g1423) & (g1741) & (!g1747) & (g1758) & (g1788)) + ((!g1423) & (g1741) & (g1747) & (!g1758) & (g1788)) + ((g1423) & (!g1741) & (!g1747) & (!g1758) & (!g1788)) + ((g1423) & (!g1741) & (!g1747) & (g1758) & (!g1788)) + ((g1423) & (!g1741) & (!g1747) & (g1758) & (g1788)) + ((g1423) & (g1741) & (!g1747) & (!g1758) & (g1788)) + ((g1423) & (g1741) & (g1747) & (!g1758) & (!g1788)) + ((g1423) & (g1741) & (g1747) & (!g1758) & (g1788)) + ((g1423) & (g1741) & (g1747) & (g1758) & (!g1788)) + ((g1423) & (g1741) & (g1747) & (g1758) & (g1788)));
	assign g1820 = (((!g1586) & (!g1568) & (g1744) & (g1746)) + ((!g1586) & (g1568) & (!g1744) & (g1746)) + ((!g1586) & (g1568) & (g1744) & (!g1746)) + ((!g1586) & (g1568) & (g1744) & (g1746)) + ((g1586) & (!g1568) & (!g1744) & (!g1746)) + ((g1586) & (!g1568) & (!g1744) & (g1746)) + ((g1586) & (!g1568) & (g1744) & (!g1746)) + ((g1586) & (g1568) & (!g1744) & (!g1746)));
	assign g1821 = (((!g1743) & (!g1758) & (!g1788) & (g1820)) + ((!g1743) & (g1758) & (!g1788) & (g1820)) + ((!g1743) & (g1758) & (g1788) & (g1820)) + ((g1743) & (!g1758) & (!g1788) & (!g1820)) + ((g1743) & (!g1758) & (g1788) & (!g1820)) + ((g1743) & (!g1758) & (g1788) & (g1820)) + ((g1743) & (g1758) & (!g1788) & (!g1820)) + ((g1743) & (g1758) & (g1788) & (!g1820)));
	assign g1822 = (((!g1568) & (!g1744) & (g1746) & (!g1758) & (!g1788)) + ((!g1568) & (!g1744) & (g1746) & (g1758) & (!g1788)) + ((!g1568) & (!g1744) & (g1746) & (g1758) & (g1788)) + ((!g1568) & (g1744) & (!g1746) & (!g1758) & (!g1788)) + ((!g1568) & (g1744) & (!g1746) & (!g1758) & (g1788)) + ((!g1568) & (g1744) & (!g1746) & (g1758) & (!g1788)) + ((!g1568) & (g1744) & (!g1746) & (g1758) & (g1788)) + ((!g1568) & (g1744) & (g1746) & (!g1758) & (g1788)) + ((g1568) & (!g1744) & (!g1746) & (!g1758) & (!g1788)) + ((g1568) & (!g1744) & (!g1746) & (g1758) & (!g1788)) + ((g1568) & (!g1744) & (!g1746) & (g1758) & (g1788)) + ((g1568) & (g1744) & (!g1746) & (!g1758) & (g1788)) + ((g1568) & (g1744) & (g1746) & (!g1758) & (!g1788)) + ((g1568) & (g1744) & (g1746) & (!g1758) & (g1788)) + ((g1568) & (g1744) & (g1746) & (g1758) & (!g1788)) + ((g1568) & (g1744) & (g1746) & (g1758) & (g1788)));
	assign g1823 = (((!g1742) & (!ax40x) & (!g1720) & (g1745)) + ((!g1742) & (!ax40x) & (g1720) & (g1745)) + ((!g1742) & (ax40x) & (!g1720) & (!g1745)) + ((!g1742) & (ax40x) & (!g1720) & (g1745)) + ((g1742) & (!ax40x) & (!g1720) & (!g1745)) + ((g1742) & (!ax40x) & (g1720) & (!g1745)) + ((g1742) & (ax40x) & (g1720) & (!g1745)) + ((g1742) & (ax40x) & (g1720) & (g1745)));
	assign g1824 = (((!ax40x) & (!ax41x) & (!g1720) & (!g1758) & (!g1788) & (g1823)) + ((!ax40x) & (!ax41x) & (!g1720) & (!g1758) & (g1788) & (!g1823)) + ((!ax40x) & (!ax41x) & (!g1720) & (!g1758) & (g1788) & (g1823)) + ((!ax40x) & (!ax41x) & (!g1720) & (g1758) & (!g1788) & (g1823)) + ((!ax40x) & (!ax41x) & (!g1720) & (g1758) & (g1788) & (g1823)) + ((!ax40x) & (!ax41x) & (g1720) & (!g1758) & (!g1788) & (!g1823)) + ((!ax40x) & (!ax41x) & (g1720) & (g1758) & (!g1788) & (!g1823)) + ((!ax40x) & (!ax41x) & (g1720) & (g1758) & (g1788) & (!g1823)) + ((!ax40x) & (ax41x) & (!g1720) & (!g1758) & (!g1788) & (!g1823)) + ((!ax40x) & (ax41x) & (!g1720) & (g1758) & (!g1788) & (!g1823)) + ((!ax40x) & (ax41x) & (!g1720) & (g1758) & (g1788) & (!g1823)) + ((!ax40x) & (ax41x) & (g1720) & (!g1758) & (!g1788) & (g1823)) + ((!ax40x) & (ax41x) & (g1720) & (!g1758) & (g1788) & (!g1823)) + ((!ax40x) & (ax41x) & (g1720) & (!g1758) & (g1788) & (g1823)) + ((!ax40x) & (ax41x) & (g1720) & (g1758) & (!g1788) & (g1823)) + ((!ax40x) & (ax41x) & (g1720) & (g1758) & (g1788) & (g1823)) + ((ax40x) & (!ax41x) & (!g1720) & (!g1758) & (!g1788) & (!g1823)) + ((ax40x) & (!ax41x) & (!g1720) & (g1758) & (!g1788) & (!g1823)) + ((ax40x) & (!ax41x) & (!g1720) & (g1758) & (g1788) & (!g1823)) + ((ax40x) & (!ax41x) & (g1720) & (!g1758) & (!g1788) & (!g1823)) + ((ax40x) & (!ax41x) & (g1720) & (g1758) & (!g1788) & (!g1823)) + ((ax40x) & (!ax41x) & (g1720) & (g1758) & (g1788) & (!g1823)) + ((ax40x) & (ax41x) & (!g1720) & (!g1758) & (!g1788) & (g1823)) + ((ax40x) & (ax41x) & (!g1720) & (!g1758) & (g1788) & (!g1823)) + ((ax40x) & (ax41x) & (!g1720) & (!g1758) & (g1788) & (g1823)) + ((ax40x) & (ax41x) & (!g1720) & (g1758) & (!g1788) & (g1823)) + ((ax40x) & (ax41x) & (!g1720) & (g1758) & (g1788) & (g1823)) + ((ax40x) & (ax41x) & (g1720) & (!g1758) & (!g1788) & (g1823)) + ((ax40x) & (ax41x) & (g1720) & (!g1758) & (g1788) & (!g1823)) + ((ax40x) & (ax41x) & (g1720) & (!g1758) & (g1788) & (g1823)) + ((ax40x) & (ax41x) & (g1720) & (g1758) & (!g1788) & (g1823)) + ((ax40x) & (ax41x) & (g1720) & (g1758) & (g1788) & (g1823)));
	assign g1825 = (((!ax40x) & (!g1720) & (!g1745) & (!g1758) & (g1788)) + ((!ax40x) & (!g1720) & (g1745) & (!g1758) & (!g1788)) + ((!ax40x) & (!g1720) & (g1745) & (!g1758) & (g1788)) + ((!ax40x) & (!g1720) & (g1745) & (g1758) & (!g1788)) + ((!ax40x) & (!g1720) & (g1745) & (g1758) & (g1788)) + ((!ax40x) & (g1720) & (g1745) & (!g1758) & (!g1788)) + ((!ax40x) & (g1720) & (g1745) & (g1758) & (!g1788)) + ((!ax40x) & (g1720) & (g1745) & (g1758) & (g1788)) + ((ax40x) & (!g1720) & (!g1745) & (!g1758) & (!g1788)) + ((ax40x) & (!g1720) & (!g1745) & (g1758) & (!g1788)) + ((ax40x) & (!g1720) & (!g1745) & (g1758) & (g1788)) + ((ax40x) & (g1720) & (!g1745) & (!g1758) & (!g1788)) + ((ax40x) & (g1720) & (!g1745) & (!g1758) & (g1788)) + ((ax40x) & (g1720) & (!g1745) & (g1758) & (!g1788)) + ((ax40x) & (g1720) & (!g1745) & (g1758) & (g1788)) + ((ax40x) & (g1720) & (g1745) & (!g1758) & (g1788)));
	assign g1826 = (((!ax36x) & (!ax37x)));
	assign g1827 = (((!g1720) & (!ax38x) & (!ax39x) & (!g1758) & (!g1788) & (!g1826)) + ((!g1720) & (!ax38x) & (!ax39x) & (g1758) & (!g1788) & (!g1826)) + ((!g1720) & (!ax38x) & (!ax39x) & (g1758) & (g1788) & (!g1826)) + ((!g1720) & (!ax38x) & (ax39x) & (!g1758) & (g1788) & (!g1826)) + ((!g1720) & (ax38x) & (ax39x) & (!g1758) & (g1788) & (!g1826)) + ((!g1720) & (ax38x) & (ax39x) & (!g1758) & (g1788) & (g1826)) + ((g1720) & (!ax38x) & (!ax39x) & (!g1758) & (!g1788) & (!g1826)) + ((g1720) & (!ax38x) & (!ax39x) & (!g1758) & (!g1788) & (g1826)) + ((g1720) & (!ax38x) & (!ax39x) & (!g1758) & (g1788) & (!g1826)) + ((g1720) & (!ax38x) & (!ax39x) & (g1758) & (!g1788) & (!g1826)) + ((g1720) & (!ax38x) & (!ax39x) & (g1758) & (!g1788) & (g1826)) + ((g1720) & (!ax38x) & (!ax39x) & (g1758) & (g1788) & (!g1826)) + ((g1720) & (!ax38x) & (!ax39x) & (g1758) & (g1788) & (g1826)) + ((g1720) & (!ax38x) & (ax39x) & (!g1758) & (!g1788) & (!g1826)) + ((g1720) & (!ax38x) & (ax39x) & (!g1758) & (g1788) & (!g1826)) + ((g1720) & (!ax38x) & (ax39x) & (!g1758) & (g1788) & (g1826)) + ((g1720) & (!ax38x) & (ax39x) & (g1758) & (!g1788) & (!g1826)) + ((g1720) & (!ax38x) & (ax39x) & (g1758) & (g1788) & (!g1826)) + ((g1720) & (ax38x) & (!ax39x) & (!g1758) & (g1788) & (!g1826)) + ((g1720) & (ax38x) & (!ax39x) & (!g1758) & (g1788) & (g1826)) + ((g1720) & (ax38x) & (ax39x) & (!g1758) & (!g1788) & (!g1826)) + ((g1720) & (ax38x) & (ax39x) & (!g1758) & (!g1788) & (g1826)) + ((g1720) & (ax38x) & (ax39x) & (!g1758) & (g1788) & (!g1826)) + ((g1720) & (ax38x) & (ax39x) & (!g1758) & (g1788) & (g1826)) + ((g1720) & (ax38x) & (ax39x) & (g1758) & (!g1788) & (!g1826)) + ((g1720) & (ax38x) & (ax39x) & (g1758) & (!g1788) & (g1826)) + ((g1720) & (ax38x) & (ax39x) & (g1758) & (g1788) & (!g1826)) + ((g1720) & (ax38x) & (ax39x) & (g1758) & (g1788) & (g1826)));
	assign g1828 = (((!g1568) & (!g1742) & (g1824) & (g1825) & (g1827)) + ((!g1568) & (g1742) & (g1824) & (!g1825) & (g1827)) + ((!g1568) & (g1742) & (g1824) & (g1825) & (!g1827)) + ((!g1568) & (g1742) & (g1824) & (g1825) & (g1827)) + ((g1568) & (!g1742) & (!g1824) & (g1825) & (g1827)) + ((g1568) & (!g1742) & (g1824) & (!g1825) & (!g1827)) + ((g1568) & (!g1742) & (g1824) & (!g1825) & (g1827)) + ((g1568) & (!g1742) & (g1824) & (g1825) & (!g1827)) + ((g1568) & (!g1742) & (g1824) & (g1825) & (g1827)) + ((g1568) & (g1742) & (!g1824) & (!g1825) & (g1827)) + ((g1568) & (g1742) & (!g1824) & (g1825) & (!g1827)) + ((g1568) & (g1742) & (!g1824) & (g1825) & (g1827)) + ((g1568) & (g1742) & (g1824) & (!g1825) & (!g1827)) + ((g1568) & (g1742) & (g1824) & (!g1825) & (g1827)) + ((g1568) & (g1742) & (g1824) & (g1825) & (!g1827)) + ((g1568) & (g1742) & (g1824) & (g1825) & (g1827)));
	assign g1829 = (((!g1423) & (!g1586) & (g1821) & (g1822) & (g1828)) + ((!g1423) & (g1586) & (g1821) & (!g1822) & (g1828)) + ((!g1423) & (g1586) & (g1821) & (g1822) & (!g1828)) + ((!g1423) & (g1586) & (g1821) & (g1822) & (g1828)) + ((g1423) & (!g1586) & (!g1821) & (g1822) & (g1828)) + ((g1423) & (!g1586) & (g1821) & (!g1822) & (!g1828)) + ((g1423) & (!g1586) & (g1821) & (!g1822) & (g1828)) + ((g1423) & (!g1586) & (g1821) & (g1822) & (!g1828)) + ((g1423) & (!g1586) & (g1821) & (g1822) & (g1828)) + ((g1423) & (g1586) & (!g1821) & (!g1822) & (g1828)) + ((g1423) & (g1586) & (!g1821) & (g1822) & (!g1828)) + ((g1423) & (g1586) & (!g1821) & (g1822) & (g1828)) + ((g1423) & (g1586) & (g1821) & (!g1822) & (!g1828)) + ((g1423) & (g1586) & (g1821) & (!g1822) & (g1828)) + ((g1423) & (g1586) & (g1821) & (g1822) & (!g1828)) + ((g1423) & (g1586) & (g1821) & (g1822) & (g1828)));
	assign g1830 = (((!g1285) & (!g1437) & (g1818) & (g1819) & (g1829)) + ((!g1285) & (g1437) & (g1818) & (!g1819) & (g1829)) + ((!g1285) & (g1437) & (g1818) & (g1819) & (!g1829)) + ((!g1285) & (g1437) & (g1818) & (g1819) & (g1829)) + ((g1285) & (!g1437) & (!g1818) & (g1819) & (g1829)) + ((g1285) & (!g1437) & (g1818) & (!g1819) & (!g1829)) + ((g1285) & (!g1437) & (g1818) & (!g1819) & (g1829)) + ((g1285) & (!g1437) & (g1818) & (g1819) & (!g1829)) + ((g1285) & (!g1437) & (g1818) & (g1819) & (g1829)) + ((g1285) & (g1437) & (!g1818) & (!g1819) & (g1829)) + ((g1285) & (g1437) & (!g1818) & (g1819) & (!g1829)) + ((g1285) & (g1437) & (!g1818) & (g1819) & (g1829)) + ((g1285) & (g1437) & (g1818) & (!g1819) & (!g1829)) + ((g1285) & (g1437) & (g1818) & (!g1819) & (g1829)) + ((g1285) & (g1437) & (g1818) & (g1819) & (!g1829)) + ((g1285) & (g1437) & (g1818) & (g1819) & (g1829)));
	assign g1831 = (((!g1154) & (!g1295) & (g1815) & (g1816) & (g1830)) + ((!g1154) & (g1295) & (g1815) & (!g1816) & (g1830)) + ((!g1154) & (g1295) & (g1815) & (g1816) & (!g1830)) + ((!g1154) & (g1295) & (g1815) & (g1816) & (g1830)) + ((g1154) & (!g1295) & (!g1815) & (g1816) & (g1830)) + ((g1154) & (!g1295) & (g1815) & (!g1816) & (!g1830)) + ((g1154) & (!g1295) & (g1815) & (!g1816) & (g1830)) + ((g1154) & (!g1295) & (g1815) & (g1816) & (!g1830)) + ((g1154) & (!g1295) & (g1815) & (g1816) & (g1830)) + ((g1154) & (g1295) & (!g1815) & (!g1816) & (g1830)) + ((g1154) & (g1295) & (!g1815) & (g1816) & (!g1830)) + ((g1154) & (g1295) & (!g1815) & (g1816) & (g1830)) + ((g1154) & (g1295) & (g1815) & (!g1816) & (!g1830)) + ((g1154) & (g1295) & (g1815) & (!g1816) & (g1830)) + ((g1154) & (g1295) & (g1815) & (g1816) & (!g1830)) + ((g1154) & (g1295) & (g1815) & (g1816) & (g1830)));
	assign g1832 = (((!g1030) & (!g1160) & (g1812) & (g1813) & (g1831)) + ((!g1030) & (g1160) & (g1812) & (!g1813) & (g1831)) + ((!g1030) & (g1160) & (g1812) & (g1813) & (!g1831)) + ((!g1030) & (g1160) & (g1812) & (g1813) & (g1831)) + ((g1030) & (!g1160) & (!g1812) & (g1813) & (g1831)) + ((g1030) & (!g1160) & (g1812) & (!g1813) & (!g1831)) + ((g1030) & (!g1160) & (g1812) & (!g1813) & (g1831)) + ((g1030) & (!g1160) & (g1812) & (g1813) & (!g1831)) + ((g1030) & (!g1160) & (g1812) & (g1813) & (g1831)) + ((g1030) & (g1160) & (!g1812) & (!g1813) & (g1831)) + ((g1030) & (g1160) & (!g1812) & (g1813) & (!g1831)) + ((g1030) & (g1160) & (!g1812) & (g1813) & (g1831)) + ((g1030) & (g1160) & (g1812) & (!g1813) & (!g1831)) + ((g1030) & (g1160) & (g1812) & (!g1813) & (g1831)) + ((g1030) & (g1160) & (g1812) & (g1813) & (!g1831)) + ((g1030) & (g1160) & (g1812) & (g1813) & (g1831)));
	assign g1833 = (((!g914) & (!g1032) & (g1809) & (g1810) & (g1832)) + ((!g914) & (g1032) & (g1809) & (!g1810) & (g1832)) + ((!g914) & (g1032) & (g1809) & (g1810) & (!g1832)) + ((!g914) & (g1032) & (g1809) & (g1810) & (g1832)) + ((g914) & (!g1032) & (!g1809) & (g1810) & (g1832)) + ((g914) & (!g1032) & (g1809) & (!g1810) & (!g1832)) + ((g914) & (!g1032) & (g1809) & (!g1810) & (g1832)) + ((g914) & (!g1032) & (g1809) & (g1810) & (!g1832)) + ((g914) & (!g1032) & (g1809) & (g1810) & (g1832)) + ((g914) & (g1032) & (!g1809) & (!g1810) & (g1832)) + ((g914) & (g1032) & (!g1809) & (g1810) & (!g1832)) + ((g914) & (g1032) & (!g1809) & (g1810) & (g1832)) + ((g914) & (g1032) & (g1809) & (!g1810) & (!g1832)) + ((g914) & (g1032) & (g1809) & (!g1810) & (g1832)) + ((g914) & (g1032) & (g1809) & (g1810) & (!g1832)) + ((g914) & (g1032) & (g1809) & (g1810) & (g1832)));
	assign g1834 = (((!g803) & (!g851) & (g1806) & (g1807) & (g1833)) + ((!g803) & (g851) & (g1806) & (!g1807) & (g1833)) + ((!g803) & (g851) & (g1806) & (g1807) & (!g1833)) + ((!g803) & (g851) & (g1806) & (g1807) & (g1833)) + ((g803) & (!g851) & (!g1806) & (g1807) & (g1833)) + ((g803) & (!g851) & (g1806) & (!g1807) & (!g1833)) + ((g803) & (!g851) & (g1806) & (!g1807) & (g1833)) + ((g803) & (!g851) & (g1806) & (g1807) & (!g1833)) + ((g803) & (!g851) & (g1806) & (g1807) & (g1833)) + ((g803) & (g851) & (!g1806) & (!g1807) & (g1833)) + ((g803) & (g851) & (!g1806) & (g1807) & (!g1833)) + ((g803) & (g851) & (!g1806) & (g1807) & (g1833)) + ((g803) & (g851) & (g1806) & (!g1807) & (!g1833)) + ((g803) & (g851) & (g1806) & (!g1807) & (g1833)) + ((g803) & (g851) & (g1806) & (g1807) & (!g1833)) + ((g803) & (g851) & (g1806) & (g1807) & (g1833)));
	assign g1835 = (((!g700) & (!g744) & (g1803) & (g1804) & (g1834)) + ((!g700) & (g744) & (g1803) & (!g1804) & (g1834)) + ((!g700) & (g744) & (g1803) & (g1804) & (!g1834)) + ((!g700) & (g744) & (g1803) & (g1804) & (g1834)) + ((g700) & (!g744) & (!g1803) & (g1804) & (g1834)) + ((g700) & (!g744) & (g1803) & (!g1804) & (!g1834)) + ((g700) & (!g744) & (g1803) & (!g1804) & (g1834)) + ((g700) & (!g744) & (g1803) & (g1804) & (!g1834)) + ((g700) & (!g744) & (g1803) & (g1804) & (g1834)) + ((g700) & (g744) & (!g1803) & (!g1804) & (g1834)) + ((g700) & (g744) & (!g1803) & (g1804) & (!g1834)) + ((g700) & (g744) & (!g1803) & (g1804) & (g1834)) + ((g700) & (g744) & (g1803) & (!g1804) & (!g1834)) + ((g700) & (g744) & (g1803) & (!g1804) & (g1834)) + ((g700) & (g744) & (g1803) & (g1804) & (!g1834)) + ((g700) & (g744) & (g1803) & (g1804) & (g1834)));
	assign g1836 = (((!g604) & (!g645) & (g1800) & (g1801) & (g1835)) + ((!g604) & (g645) & (g1800) & (!g1801) & (g1835)) + ((!g604) & (g645) & (g1800) & (g1801) & (!g1835)) + ((!g604) & (g645) & (g1800) & (g1801) & (g1835)) + ((g604) & (!g645) & (!g1800) & (g1801) & (g1835)) + ((g604) & (!g645) & (g1800) & (!g1801) & (!g1835)) + ((g604) & (!g645) & (g1800) & (!g1801) & (g1835)) + ((g604) & (!g645) & (g1800) & (g1801) & (!g1835)) + ((g604) & (!g645) & (g1800) & (g1801) & (g1835)) + ((g604) & (g645) & (!g1800) & (!g1801) & (g1835)) + ((g604) & (g645) & (!g1800) & (g1801) & (!g1835)) + ((g604) & (g645) & (!g1800) & (g1801) & (g1835)) + ((g604) & (g645) & (g1800) & (!g1801) & (!g1835)) + ((g604) & (g645) & (g1800) & (!g1801) & (g1835)) + ((g604) & (g645) & (g1800) & (g1801) & (!g1835)) + ((g604) & (g645) & (g1800) & (g1801) & (g1835)));
	assign g1837 = (((!g515) & (!g553) & (g1797) & (g1798) & (g1836)) + ((!g515) & (g553) & (g1797) & (!g1798) & (g1836)) + ((!g515) & (g553) & (g1797) & (g1798) & (!g1836)) + ((!g515) & (g553) & (g1797) & (g1798) & (g1836)) + ((g515) & (!g553) & (!g1797) & (g1798) & (g1836)) + ((g515) & (!g553) & (g1797) & (!g1798) & (!g1836)) + ((g515) & (!g553) & (g1797) & (!g1798) & (g1836)) + ((g515) & (!g553) & (g1797) & (g1798) & (!g1836)) + ((g515) & (!g553) & (g1797) & (g1798) & (g1836)) + ((g515) & (g553) & (!g1797) & (!g1798) & (g1836)) + ((g515) & (g553) & (!g1797) & (g1798) & (!g1836)) + ((g515) & (g553) & (!g1797) & (g1798) & (g1836)) + ((g515) & (g553) & (g1797) & (!g1798) & (!g1836)) + ((g515) & (g553) & (g1797) & (!g1798) & (g1836)) + ((g515) & (g553) & (g1797) & (g1798) & (!g1836)) + ((g515) & (g553) & (g1797) & (g1798) & (g1836)));
	assign g1838 = (((!g433) & (!g468) & (g1794) & (g1795) & (g1837)) + ((!g433) & (g468) & (g1794) & (!g1795) & (g1837)) + ((!g433) & (g468) & (g1794) & (g1795) & (!g1837)) + ((!g433) & (g468) & (g1794) & (g1795) & (g1837)) + ((g433) & (!g468) & (!g1794) & (g1795) & (g1837)) + ((g433) & (!g468) & (g1794) & (!g1795) & (!g1837)) + ((g433) & (!g468) & (g1794) & (!g1795) & (g1837)) + ((g433) & (!g468) & (g1794) & (g1795) & (!g1837)) + ((g433) & (!g468) & (g1794) & (g1795) & (g1837)) + ((g433) & (g468) & (!g1794) & (!g1795) & (g1837)) + ((g433) & (g468) & (!g1794) & (g1795) & (!g1837)) + ((g433) & (g468) & (!g1794) & (g1795) & (g1837)) + ((g433) & (g468) & (g1794) & (!g1795) & (!g1837)) + ((g433) & (g468) & (g1794) & (!g1795) & (g1837)) + ((g433) & (g468) & (g1794) & (g1795) & (!g1837)) + ((g433) & (g468) & (g1794) & (g1795) & (g1837)));
	assign g1839 = (((!g358) & (!g390) & (g1791) & (g1792) & (g1838)) + ((!g358) & (g390) & (g1791) & (!g1792) & (g1838)) + ((!g358) & (g390) & (g1791) & (g1792) & (!g1838)) + ((!g358) & (g390) & (g1791) & (g1792) & (g1838)) + ((g358) & (!g390) & (!g1791) & (g1792) & (g1838)) + ((g358) & (!g390) & (g1791) & (!g1792) & (!g1838)) + ((g358) & (!g390) & (g1791) & (!g1792) & (g1838)) + ((g358) & (!g390) & (g1791) & (g1792) & (!g1838)) + ((g358) & (!g390) & (g1791) & (g1792) & (g1838)) + ((g358) & (g390) & (!g1791) & (!g1792) & (g1838)) + ((g358) & (g390) & (!g1791) & (g1792) & (!g1838)) + ((g358) & (g390) & (!g1791) & (g1792) & (g1838)) + ((g358) & (g390) & (g1791) & (!g1792) & (!g1838)) + ((g358) & (g390) & (g1791) & (!g1792) & (g1838)) + ((g358) & (g390) & (g1791) & (g1792) & (!g1838)) + ((g358) & (g390) & (g1791) & (g1792) & (g1838)));
	assign g1840 = (((!g4) & (!g1785) & (!g1786) & (!g1758) & (!g1788)) + ((!g4) & (!g1785) & (!g1786) & (g1758) & (!g1788)) + ((!g4) & (!g1785) & (!g1786) & (g1758) & (g1788)) + ((!g4) & (!g1785) & (g1786) & (!g1758) & (g1788)) + ((!g4) & (g1785) & (g1786) & (!g1758) & (!g1788)) + ((!g4) & (g1785) & (g1786) & (!g1758) & (g1788)) + ((!g4) & (g1785) & (g1786) & (g1758) & (!g1788)) + ((!g4) & (g1785) & (g1786) & (g1758) & (g1788)) + ((g4) & (!g1785) & (g1786) & (!g1758) & (!g1788)) + ((g4) & (!g1785) & (g1786) & (!g1758) & (g1788)) + ((g4) & (!g1785) & (g1786) & (g1758) & (!g1788)) + ((g4) & (!g1785) & (g1786) & (g1758) & (g1788)) + ((g4) & (g1785) & (!g1786) & (!g1758) & (!g1788)) + ((g4) & (g1785) & (!g1786) & (g1758) & (!g1788)) + ((g4) & (g1785) & (!g1786) & (g1758) & (g1788)) + ((g4) & (g1785) & (g1786) & (!g1758) & (g1788)));
	assign g1841 = (((!g8) & (!g1761) & (g1784) & (!g1758) & (!g1788)) + ((!g8) & (!g1761) & (g1784) & (g1758) & (!g1788)) + ((!g8) & (!g1761) & (g1784) & (g1758) & (g1788)) + ((!g8) & (g1761) & (!g1784) & (!g1758) & (!g1788)) + ((!g8) & (g1761) & (!g1784) & (!g1758) & (g1788)) + ((!g8) & (g1761) & (!g1784) & (g1758) & (!g1788)) + ((!g8) & (g1761) & (!g1784) & (g1758) & (g1788)) + ((!g8) & (g1761) & (g1784) & (!g1758) & (g1788)) + ((g8) & (!g1761) & (!g1784) & (!g1758) & (!g1788)) + ((g8) & (!g1761) & (!g1784) & (g1758) & (!g1788)) + ((g8) & (!g1761) & (!g1784) & (g1758) & (g1788)) + ((g8) & (g1761) & (!g1784) & (!g1758) & (g1788)) + ((g8) & (g1761) & (g1784) & (!g1758) & (!g1788)) + ((g8) & (g1761) & (g1784) & (!g1758) & (g1788)) + ((g8) & (g1761) & (g1784) & (g1758) & (!g1788)) + ((g8) & (g1761) & (g1784) & (g1758) & (g1788)));
	assign g1842 = (((!g18) & (!g27) & (g1763) & (g1783)) + ((!g18) & (g27) & (!g1763) & (g1783)) + ((!g18) & (g27) & (g1763) & (!g1783)) + ((!g18) & (g27) & (g1763) & (g1783)) + ((g18) & (!g27) & (!g1763) & (!g1783)) + ((g18) & (!g27) & (!g1763) & (g1783)) + ((g18) & (!g27) & (g1763) & (!g1783)) + ((g18) & (g27) & (!g1763) & (!g1783)));
	assign g1843 = (((!g1762) & (!g1758) & (!g1788) & (g1842)) + ((!g1762) & (g1758) & (!g1788) & (g1842)) + ((!g1762) & (g1758) & (g1788) & (g1842)) + ((g1762) & (!g1758) & (!g1788) & (!g1842)) + ((g1762) & (!g1758) & (g1788) & (!g1842)) + ((g1762) & (!g1758) & (g1788) & (g1842)) + ((g1762) & (g1758) & (!g1788) & (!g1842)) + ((g1762) & (g1758) & (g1788) & (!g1842)));
	assign g1844 = (((!g27) & (!g1763) & (g1783) & (!g1758) & (!g1788)) + ((!g27) & (!g1763) & (g1783) & (g1758) & (!g1788)) + ((!g27) & (!g1763) & (g1783) & (g1758) & (g1788)) + ((!g27) & (g1763) & (!g1783) & (!g1758) & (!g1788)) + ((!g27) & (g1763) & (!g1783) & (!g1758) & (g1788)) + ((!g27) & (g1763) & (!g1783) & (g1758) & (!g1788)) + ((!g27) & (g1763) & (!g1783) & (g1758) & (g1788)) + ((!g27) & (g1763) & (g1783) & (!g1758) & (g1788)) + ((g27) & (!g1763) & (!g1783) & (!g1758) & (!g1788)) + ((g27) & (!g1763) & (!g1783) & (g1758) & (!g1788)) + ((g27) & (!g1763) & (!g1783) & (g1758) & (g1788)) + ((g27) & (g1763) & (!g1783) & (!g1758) & (g1788)) + ((g27) & (g1763) & (g1783) & (!g1758) & (!g1788)) + ((g27) & (g1763) & (g1783) & (!g1758) & (g1788)) + ((g27) & (g1763) & (g1783) & (g1758) & (!g1788)) + ((g27) & (g1763) & (g1783) & (g1758) & (g1788)));
	assign g1845 = (((!g39) & (!g54) & (g1765) & (g1782)) + ((!g39) & (g54) & (!g1765) & (g1782)) + ((!g39) & (g54) & (g1765) & (!g1782)) + ((!g39) & (g54) & (g1765) & (g1782)) + ((g39) & (!g54) & (!g1765) & (!g1782)) + ((g39) & (!g54) & (!g1765) & (g1782)) + ((g39) & (!g54) & (g1765) & (!g1782)) + ((g39) & (g54) & (!g1765) & (!g1782)));
	assign g1846 = (((!g1764) & (!g1758) & (!g1788) & (g1845)) + ((!g1764) & (g1758) & (!g1788) & (g1845)) + ((!g1764) & (g1758) & (g1788) & (g1845)) + ((g1764) & (!g1758) & (!g1788) & (!g1845)) + ((g1764) & (!g1758) & (g1788) & (!g1845)) + ((g1764) & (!g1758) & (g1788) & (g1845)) + ((g1764) & (g1758) & (!g1788) & (!g1845)) + ((g1764) & (g1758) & (g1788) & (!g1845)));
	assign g1847 = (((!g54) & (!g1765) & (g1782) & (!g1758) & (!g1788)) + ((!g54) & (!g1765) & (g1782) & (g1758) & (!g1788)) + ((!g54) & (!g1765) & (g1782) & (g1758) & (g1788)) + ((!g54) & (g1765) & (!g1782) & (!g1758) & (!g1788)) + ((!g54) & (g1765) & (!g1782) & (!g1758) & (g1788)) + ((!g54) & (g1765) & (!g1782) & (g1758) & (!g1788)) + ((!g54) & (g1765) & (!g1782) & (g1758) & (g1788)) + ((!g54) & (g1765) & (g1782) & (!g1758) & (g1788)) + ((g54) & (!g1765) & (!g1782) & (!g1758) & (!g1788)) + ((g54) & (!g1765) & (!g1782) & (g1758) & (!g1788)) + ((g54) & (!g1765) & (!g1782) & (g1758) & (g1788)) + ((g54) & (g1765) & (!g1782) & (!g1758) & (g1788)) + ((g54) & (g1765) & (g1782) & (!g1758) & (!g1788)) + ((g54) & (g1765) & (g1782) & (!g1758) & (g1788)) + ((g54) & (g1765) & (g1782) & (g1758) & (!g1788)) + ((g54) & (g1765) & (g1782) & (g1758) & (g1788)));
	assign g1848 = (((!g68) & (!g87) & (g1767) & (g1781)) + ((!g68) & (g87) & (!g1767) & (g1781)) + ((!g68) & (g87) & (g1767) & (!g1781)) + ((!g68) & (g87) & (g1767) & (g1781)) + ((g68) & (!g87) & (!g1767) & (!g1781)) + ((g68) & (!g87) & (!g1767) & (g1781)) + ((g68) & (!g87) & (g1767) & (!g1781)) + ((g68) & (g87) & (!g1767) & (!g1781)));
	assign g1849 = (((!g1766) & (!g1758) & (!g1788) & (g1848)) + ((!g1766) & (g1758) & (!g1788) & (g1848)) + ((!g1766) & (g1758) & (g1788) & (g1848)) + ((g1766) & (!g1758) & (!g1788) & (!g1848)) + ((g1766) & (!g1758) & (g1788) & (!g1848)) + ((g1766) & (!g1758) & (g1788) & (g1848)) + ((g1766) & (g1758) & (!g1788) & (!g1848)) + ((g1766) & (g1758) & (g1788) & (!g1848)));
	assign g1850 = (((!g87) & (!g1767) & (g1781) & (!g1758) & (!g1788)) + ((!g87) & (!g1767) & (g1781) & (g1758) & (!g1788)) + ((!g87) & (!g1767) & (g1781) & (g1758) & (g1788)) + ((!g87) & (g1767) & (!g1781) & (!g1758) & (!g1788)) + ((!g87) & (g1767) & (!g1781) & (!g1758) & (g1788)) + ((!g87) & (g1767) & (!g1781) & (g1758) & (!g1788)) + ((!g87) & (g1767) & (!g1781) & (g1758) & (g1788)) + ((!g87) & (g1767) & (g1781) & (!g1758) & (g1788)) + ((g87) & (!g1767) & (!g1781) & (!g1758) & (!g1788)) + ((g87) & (!g1767) & (!g1781) & (g1758) & (!g1788)) + ((g87) & (!g1767) & (!g1781) & (g1758) & (g1788)) + ((g87) & (g1767) & (!g1781) & (!g1758) & (g1788)) + ((g87) & (g1767) & (g1781) & (!g1758) & (!g1788)) + ((g87) & (g1767) & (g1781) & (!g1758) & (g1788)) + ((g87) & (g1767) & (g1781) & (g1758) & (!g1788)) + ((g87) & (g1767) & (g1781) & (g1758) & (g1788)));
	assign g1851 = (((!g104) & (!g127) & (g1769) & (g1780)) + ((!g104) & (g127) & (!g1769) & (g1780)) + ((!g104) & (g127) & (g1769) & (!g1780)) + ((!g104) & (g127) & (g1769) & (g1780)) + ((g104) & (!g127) & (!g1769) & (!g1780)) + ((g104) & (!g127) & (!g1769) & (g1780)) + ((g104) & (!g127) & (g1769) & (!g1780)) + ((g104) & (g127) & (!g1769) & (!g1780)));
	assign g1852 = (((!g1768) & (!g1758) & (!g1788) & (g1851)) + ((!g1768) & (g1758) & (!g1788) & (g1851)) + ((!g1768) & (g1758) & (g1788) & (g1851)) + ((g1768) & (!g1758) & (!g1788) & (!g1851)) + ((g1768) & (!g1758) & (g1788) & (!g1851)) + ((g1768) & (!g1758) & (g1788) & (g1851)) + ((g1768) & (g1758) & (!g1788) & (!g1851)) + ((g1768) & (g1758) & (g1788) & (!g1851)));
	assign g1853 = (((!g127) & (!g1769) & (g1780) & (!g1758) & (!g1788)) + ((!g127) & (!g1769) & (g1780) & (g1758) & (!g1788)) + ((!g127) & (!g1769) & (g1780) & (g1758) & (g1788)) + ((!g127) & (g1769) & (!g1780) & (!g1758) & (!g1788)) + ((!g127) & (g1769) & (!g1780) & (!g1758) & (g1788)) + ((!g127) & (g1769) & (!g1780) & (g1758) & (!g1788)) + ((!g127) & (g1769) & (!g1780) & (g1758) & (g1788)) + ((!g127) & (g1769) & (g1780) & (!g1758) & (g1788)) + ((g127) & (!g1769) & (!g1780) & (!g1758) & (!g1788)) + ((g127) & (!g1769) & (!g1780) & (g1758) & (!g1788)) + ((g127) & (!g1769) & (!g1780) & (g1758) & (g1788)) + ((g127) & (g1769) & (!g1780) & (!g1758) & (g1788)) + ((g127) & (g1769) & (g1780) & (!g1758) & (!g1788)) + ((g127) & (g1769) & (g1780) & (!g1758) & (g1788)) + ((g127) & (g1769) & (g1780) & (g1758) & (!g1788)) + ((g127) & (g1769) & (g1780) & (g1758) & (g1788)));
	assign g1854 = (((!g147) & (!g174) & (g1771) & (g1779)) + ((!g147) & (g174) & (!g1771) & (g1779)) + ((!g147) & (g174) & (g1771) & (!g1779)) + ((!g147) & (g174) & (g1771) & (g1779)) + ((g147) & (!g174) & (!g1771) & (!g1779)) + ((g147) & (!g174) & (!g1771) & (g1779)) + ((g147) & (!g174) & (g1771) & (!g1779)) + ((g147) & (g174) & (!g1771) & (!g1779)));
	assign g1855 = (((!g1770) & (!g1758) & (!g1788) & (g1854)) + ((!g1770) & (g1758) & (!g1788) & (g1854)) + ((!g1770) & (g1758) & (g1788) & (g1854)) + ((g1770) & (!g1758) & (!g1788) & (!g1854)) + ((g1770) & (!g1758) & (g1788) & (!g1854)) + ((g1770) & (!g1758) & (g1788) & (g1854)) + ((g1770) & (g1758) & (!g1788) & (!g1854)) + ((g1770) & (g1758) & (g1788) & (!g1854)));
	assign g1856 = (((!g174) & (!g1771) & (g1779) & (!g1758) & (!g1788)) + ((!g174) & (!g1771) & (g1779) & (g1758) & (!g1788)) + ((!g174) & (!g1771) & (g1779) & (g1758) & (g1788)) + ((!g174) & (g1771) & (!g1779) & (!g1758) & (!g1788)) + ((!g174) & (g1771) & (!g1779) & (!g1758) & (g1788)) + ((!g174) & (g1771) & (!g1779) & (g1758) & (!g1788)) + ((!g174) & (g1771) & (!g1779) & (g1758) & (g1788)) + ((!g174) & (g1771) & (g1779) & (!g1758) & (g1788)) + ((g174) & (!g1771) & (!g1779) & (!g1758) & (!g1788)) + ((g174) & (!g1771) & (!g1779) & (g1758) & (!g1788)) + ((g174) & (!g1771) & (!g1779) & (g1758) & (g1788)) + ((g174) & (g1771) & (!g1779) & (!g1758) & (g1788)) + ((g174) & (g1771) & (g1779) & (!g1758) & (!g1788)) + ((g174) & (g1771) & (g1779) & (!g1758) & (g1788)) + ((g174) & (g1771) & (g1779) & (g1758) & (!g1788)) + ((g174) & (g1771) & (g1779) & (g1758) & (g1788)));
	assign g1857 = (((!g198) & (!g229) & (g1773) & (g1778)) + ((!g198) & (g229) & (!g1773) & (g1778)) + ((!g198) & (g229) & (g1773) & (!g1778)) + ((!g198) & (g229) & (g1773) & (g1778)) + ((g198) & (!g229) & (!g1773) & (!g1778)) + ((g198) & (!g229) & (!g1773) & (g1778)) + ((g198) & (!g229) & (g1773) & (!g1778)) + ((g198) & (g229) & (!g1773) & (!g1778)));
	assign g1858 = (((!g1772) & (!g1758) & (!g1788) & (g1857)) + ((!g1772) & (g1758) & (!g1788) & (g1857)) + ((!g1772) & (g1758) & (g1788) & (g1857)) + ((g1772) & (!g1758) & (!g1788) & (!g1857)) + ((g1772) & (!g1758) & (g1788) & (!g1857)) + ((g1772) & (!g1758) & (g1788) & (g1857)) + ((g1772) & (g1758) & (!g1788) & (!g1857)) + ((g1772) & (g1758) & (g1788) & (!g1857)));
	assign g1859 = (((!g229) & (!g1773) & (g1778) & (!g1758) & (!g1788)) + ((!g229) & (!g1773) & (g1778) & (g1758) & (!g1788)) + ((!g229) & (!g1773) & (g1778) & (g1758) & (g1788)) + ((!g229) & (g1773) & (!g1778) & (!g1758) & (!g1788)) + ((!g229) & (g1773) & (!g1778) & (!g1758) & (g1788)) + ((!g229) & (g1773) & (!g1778) & (g1758) & (!g1788)) + ((!g229) & (g1773) & (!g1778) & (g1758) & (g1788)) + ((!g229) & (g1773) & (g1778) & (!g1758) & (g1788)) + ((g229) & (!g1773) & (!g1778) & (!g1758) & (!g1788)) + ((g229) & (!g1773) & (!g1778) & (g1758) & (!g1788)) + ((g229) & (!g1773) & (!g1778) & (g1758) & (g1788)) + ((g229) & (g1773) & (!g1778) & (!g1758) & (g1788)) + ((g229) & (g1773) & (g1778) & (!g1758) & (!g1788)) + ((g229) & (g1773) & (g1778) & (!g1758) & (g1788)) + ((g229) & (g1773) & (g1778) & (g1758) & (!g1788)) + ((g229) & (g1773) & (g1778) & (g1758) & (g1788)));
	assign g1860 = (((!g255) & (!g290) & (g1775) & (g1777)) + ((!g255) & (g290) & (!g1775) & (g1777)) + ((!g255) & (g290) & (g1775) & (!g1777)) + ((!g255) & (g290) & (g1775) & (g1777)) + ((g255) & (!g290) & (!g1775) & (!g1777)) + ((g255) & (!g290) & (!g1775) & (g1777)) + ((g255) & (!g290) & (g1775) & (!g1777)) + ((g255) & (g290) & (!g1775) & (!g1777)));
	assign g1861 = (((!g1774) & (!g1758) & (!g1788) & (g1860)) + ((!g1774) & (g1758) & (!g1788) & (g1860)) + ((!g1774) & (g1758) & (g1788) & (g1860)) + ((g1774) & (!g1758) & (!g1788) & (!g1860)) + ((g1774) & (!g1758) & (g1788) & (!g1860)) + ((g1774) & (!g1758) & (g1788) & (g1860)) + ((g1774) & (g1758) & (!g1788) & (!g1860)) + ((g1774) & (g1758) & (g1788) & (!g1860)));
	assign g1862 = (((!g290) & (!g1775) & (g1777) & (!g1758) & (!g1788)) + ((!g290) & (!g1775) & (g1777) & (g1758) & (!g1788)) + ((!g290) & (!g1775) & (g1777) & (g1758) & (g1788)) + ((!g290) & (g1775) & (!g1777) & (!g1758) & (!g1788)) + ((!g290) & (g1775) & (!g1777) & (!g1758) & (g1788)) + ((!g290) & (g1775) & (!g1777) & (g1758) & (!g1788)) + ((!g290) & (g1775) & (!g1777) & (g1758) & (g1788)) + ((!g290) & (g1775) & (g1777) & (!g1758) & (g1788)) + ((g290) & (!g1775) & (!g1777) & (!g1758) & (!g1788)) + ((g290) & (!g1775) & (!g1777) & (g1758) & (!g1788)) + ((g290) & (!g1775) & (!g1777) & (g1758) & (g1788)) + ((g290) & (g1775) & (!g1777) & (!g1758) & (g1788)) + ((g290) & (g1775) & (g1777) & (!g1758) & (!g1788)) + ((g290) & (g1775) & (g1777) & (!g1758) & (g1788)) + ((g290) & (g1775) & (g1777) & (g1758) & (!g1788)) + ((g290) & (g1775) & (g1777) & (g1758) & (g1788)));
	assign g1863 = (((!g319) & (!g358) & (g1721) & (g1757)) + ((!g319) & (g358) & (!g1721) & (g1757)) + ((!g319) & (g358) & (g1721) & (!g1757)) + ((!g319) & (g358) & (g1721) & (g1757)) + ((g319) & (!g358) & (!g1721) & (!g1757)) + ((g319) & (!g358) & (!g1721) & (g1757)) + ((g319) & (!g358) & (g1721) & (!g1757)) + ((g319) & (g358) & (!g1721) & (!g1757)));
	assign g1864 = (((!g1776) & (!g1758) & (!g1788) & (g1863)) + ((!g1776) & (g1758) & (!g1788) & (g1863)) + ((!g1776) & (g1758) & (g1788) & (g1863)) + ((g1776) & (!g1758) & (!g1788) & (!g1863)) + ((g1776) & (!g1758) & (g1788) & (!g1863)) + ((g1776) & (!g1758) & (g1788) & (g1863)) + ((g1776) & (g1758) & (!g1788) & (!g1863)) + ((g1776) & (g1758) & (g1788) & (!g1863)));
	assign g1865 = (((!g290) & (!g319) & (g1864) & (g1789) & (g1839)) + ((!g290) & (g319) & (g1864) & (!g1789) & (g1839)) + ((!g290) & (g319) & (g1864) & (g1789) & (!g1839)) + ((!g290) & (g319) & (g1864) & (g1789) & (g1839)) + ((g290) & (!g319) & (!g1864) & (g1789) & (g1839)) + ((g290) & (!g319) & (g1864) & (!g1789) & (!g1839)) + ((g290) & (!g319) & (g1864) & (!g1789) & (g1839)) + ((g290) & (!g319) & (g1864) & (g1789) & (!g1839)) + ((g290) & (!g319) & (g1864) & (g1789) & (g1839)) + ((g290) & (g319) & (!g1864) & (!g1789) & (g1839)) + ((g290) & (g319) & (!g1864) & (g1789) & (!g1839)) + ((g290) & (g319) & (!g1864) & (g1789) & (g1839)) + ((g290) & (g319) & (g1864) & (!g1789) & (!g1839)) + ((g290) & (g319) & (g1864) & (!g1789) & (g1839)) + ((g290) & (g319) & (g1864) & (g1789) & (!g1839)) + ((g290) & (g319) & (g1864) & (g1789) & (g1839)));
	assign g1866 = (((!g229) & (!g255) & (g1861) & (g1862) & (g1865)) + ((!g229) & (g255) & (g1861) & (!g1862) & (g1865)) + ((!g229) & (g255) & (g1861) & (g1862) & (!g1865)) + ((!g229) & (g255) & (g1861) & (g1862) & (g1865)) + ((g229) & (!g255) & (!g1861) & (g1862) & (g1865)) + ((g229) & (!g255) & (g1861) & (!g1862) & (!g1865)) + ((g229) & (!g255) & (g1861) & (!g1862) & (g1865)) + ((g229) & (!g255) & (g1861) & (g1862) & (!g1865)) + ((g229) & (!g255) & (g1861) & (g1862) & (g1865)) + ((g229) & (g255) & (!g1861) & (!g1862) & (g1865)) + ((g229) & (g255) & (!g1861) & (g1862) & (!g1865)) + ((g229) & (g255) & (!g1861) & (g1862) & (g1865)) + ((g229) & (g255) & (g1861) & (!g1862) & (!g1865)) + ((g229) & (g255) & (g1861) & (!g1862) & (g1865)) + ((g229) & (g255) & (g1861) & (g1862) & (!g1865)) + ((g229) & (g255) & (g1861) & (g1862) & (g1865)));
	assign g1867 = (((!g174) & (!g198) & (g1858) & (g1859) & (g1866)) + ((!g174) & (g198) & (g1858) & (!g1859) & (g1866)) + ((!g174) & (g198) & (g1858) & (g1859) & (!g1866)) + ((!g174) & (g198) & (g1858) & (g1859) & (g1866)) + ((g174) & (!g198) & (!g1858) & (g1859) & (g1866)) + ((g174) & (!g198) & (g1858) & (!g1859) & (!g1866)) + ((g174) & (!g198) & (g1858) & (!g1859) & (g1866)) + ((g174) & (!g198) & (g1858) & (g1859) & (!g1866)) + ((g174) & (!g198) & (g1858) & (g1859) & (g1866)) + ((g174) & (g198) & (!g1858) & (!g1859) & (g1866)) + ((g174) & (g198) & (!g1858) & (g1859) & (!g1866)) + ((g174) & (g198) & (!g1858) & (g1859) & (g1866)) + ((g174) & (g198) & (g1858) & (!g1859) & (!g1866)) + ((g174) & (g198) & (g1858) & (!g1859) & (g1866)) + ((g174) & (g198) & (g1858) & (g1859) & (!g1866)) + ((g174) & (g198) & (g1858) & (g1859) & (g1866)));
	assign g1868 = (((!g127) & (!g147) & (g1855) & (g1856) & (g1867)) + ((!g127) & (g147) & (g1855) & (!g1856) & (g1867)) + ((!g127) & (g147) & (g1855) & (g1856) & (!g1867)) + ((!g127) & (g147) & (g1855) & (g1856) & (g1867)) + ((g127) & (!g147) & (!g1855) & (g1856) & (g1867)) + ((g127) & (!g147) & (g1855) & (!g1856) & (!g1867)) + ((g127) & (!g147) & (g1855) & (!g1856) & (g1867)) + ((g127) & (!g147) & (g1855) & (g1856) & (!g1867)) + ((g127) & (!g147) & (g1855) & (g1856) & (g1867)) + ((g127) & (g147) & (!g1855) & (!g1856) & (g1867)) + ((g127) & (g147) & (!g1855) & (g1856) & (!g1867)) + ((g127) & (g147) & (!g1855) & (g1856) & (g1867)) + ((g127) & (g147) & (g1855) & (!g1856) & (!g1867)) + ((g127) & (g147) & (g1855) & (!g1856) & (g1867)) + ((g127) & (g147) & (g1855) & (g1856) & (!g1867)) + ((g127) & (g147) & (g1855) & (g1856) & (g1867)));
	assign g1869 = (((!g87) & (!g104) & (g1852) & (g1853) & (g1868)) + ((!g87) & (g104) & (g1852) & (!g1853) & (g1868)) + ((!g87) & (g104) & (g1852) & (g1853) & (!g1868)) + ((!g87) & (g104) & (g1852) & (g1853) & (g1868)) + ((g87) & (!g104) & (!g1852) & (g1853) & (g1868)) + ((g87) & (!g104) & (g1852) & (!g1853) & (!g1868)) + ((g87) & (!g104) & (g1852) & (!g1853) & (g1868)) + ((g87) & (!g104) & (g1852) & (g1853) & (!g1868)) + ((g87) & (!g104) & (g1852) & (g1853) & (g1868)) + ((g87) & (g104) & (!g1852) & (!g1853) & (g1868)) + ((g87) & (g104) & (!g1852) & (g1853) & (!g1868)) + ((g87) & (g104) & (!g1852) & (g1853) & (g1868)) + ((g87) & (g104) & (g1852) & (!g1853) & (!g1868)) + ((g87) & (g104) & (g1852) & (!g1853) & (g1868)) + ((g87) & (g104) & (g1852) & (g1853) & (!g1868)) + ((g87) & (g104) & (g1852) & (g1853) & (g1868)));
	assign g1870 = (((!g54) & (!g68) & (g1849) & (g1850) & (g1869)) + ((!g54) & (g68) & (g1849) & (!g1850) & (g1869)) + ((!g54) & (g68) & (g1849) & (g1850) & (!g1869)) + ((!g54) & (g68) & (g1849) & (g1850) & (g1869)) + ((g54) & (!g68) & (!g1849) & (g1850) & (g1869)) + ((g54) & (!g68) & (g1849) & (!g1850) & (!g1869)) + ((g54) & (!g68) & (g1849) & (!g1850) & (g1869)) + ((g54) & (!g68) & (g1849) & (g1850) & (!g1869)) + ((g54) & (!g68) & (g1849) & (g1850) & (g1869)) + ((g54) & (g68) & (!g1849) & (!g1850) & (g1869)) + ((g54) & (g68) & (!g1849) & (g1850) & (!g1869)) + ((g54) & (g68) & (!g1849) & (g1850) & (g1869)) + ((g54) & (g68) & (g1849) & (!g1850) & (!g1869)) + ((g54) & (g68) & (g1849) & (!g1850) & (g1869)) + ((g54) & (g68) & (g1849) & (g1850) & (!g1869)) + ((g54) & (g68) & (g1849) & (g1850) & (g1869)));
	assign g1871 = (((!g27) & (!g39) & (g1846) & (g1847) & (g1870)) + ((!g27) & (g39) & (g1846) & (!g1847) & (g1870)) + ((!g27) & (g39) & (g1846) & (g1847) & (!g1870)) + ((!g27) & (g39) & (g1846) & (g1847) & (g1870)) + ((g27) & (!g39) & (!g1846) & (g1847) & (g1870)) + ((g27) & (!g39) & (g1846) & (!g1847) & (!g1870)) + ((g27) & (!g39) & (g1846) & (!g1847) & (g1870)) + ((g27) & (!g39) & (g1846) & (g1847) & (!g1870)) + ((g27) & (!g39) & (g1846) & (g1847) & (g1870)) + ((g27) & (g39) & (!g1846) & (!g1847) & (g1870)) + ((g27) & (g39) & (!g1846) & (g1847) & (!g1870)) + ((g27) & (g39) & (!g1846) & (g1847) & (g1870)) + ((g27) & (g39) & (g1846) & (!g1847) & (!g1870)) + ((g27) & (g39) & (g1846) & (!g1847) & (g1870)) + ((g27) & (g39) & (g1846) & (g1847) & (!g1870)) + ((g27) & (g39) & (g1846) & (g1847) & (g1870)));
	assign g1872 = (((!g8) & (!g18) & (g1843) & (g1844) & (g1871)) + ((!g8) & (g18) & (g1843) & (!g1844) & (g1871)) + ((!g8) & (g18) & (g1843) & (g1844) & (!g1871)) + ((!g8) & (g18) & (g1843) & (g1844) & (g1871)) + ((g8) & (!g18) & (!g1843) & (g1844) & (g1871)) + ((g8) & (!g18) & (g1843) & (!g1844) & (!g1871)) + ((g8) & (!g18) & (g1843) & (!g1844) & (g1871)) + ((g8) & (!g18) & (g1843) & (g1844) & (!g1871)) + ((g8) & (!g18) & (g1843) & (g1844) & (g1871)) + ((g8) & (g18) & (!g1843) & (!g1844) & (g1871)) + ((g8) & (g18) & (!g1843) & (g1844) & (!g1871)) + ((g8) & (g18) & (!g1843) & (g1844) & (g1871)) + ((g8) & (g18) & (g1843) & (!g1844) & (!g1871)) + ((g8) & (g18) & (g1843) & (!g1844) & (g1871)) + ((g8) & (g18) & (g1843) & (g1844) & (!g1871)) + ((g8) & (g18) & (g1843) & (g1844) & (g1871)));
	assign g1873 = (((!g2) & (!g8) & (g1761) & (g1784)) + ((!g2) & (g8) & (!g1761) & (g1784)) + ((!g2) & (g8) & (g1761) & (!g1784)) + ((!g2) & (g8) & (g1761) & (g1784)) + ((g2) & (!g8) & (!g1761) & (!g1784)) + ((g2) & (!g8) & (!g1761) & (g1784)) + ((g2) & (!g8) & (g1761) & (!g1784)) + ((g2) & (g8) & (!g1761) & (!g1784)));
	assign g1874 = (((!g1760) & (!g1758) & (!g1788) & (g1873)) + ((!g1760) & (g1758) & (!g1788) & (g1873)) + ((!g1760) & (g1758) & (g1788) & (g1873)) + ((g1760) & (!g1758) & (!g1788) & (!g1873)) + ((g1760) & (!g1758) & (g1788) & (!g1873)) + ((g1760) & (!g1758) & (g1788) & (g1873)) + ((g1760) & (g1758) & (!g1788) & (!g1873)) + ((g1760) & (g1758) & (g1788) & (!g1873)));
	assign g1875 = (((!g4) & (!g2) & (!g1841) & (!g1872) & (g1874)) + ((!g4) & (!g2) & (!g1841) & (g1872) & (g1874)) + ((!g4) & (!g2) & (g1841) & (!g1872) & (g1874)) + ((!g4) & (!g2) & (g1841) & (g1872) & (!g1874)) + ((!g4) & (!g2) & (g1841) & (g1872) & (g1874)) + ((!g4) & (g2) & (!g1841) & (!g1872) & (g1874)) + ((!g4) & (g2) & (!g1841) & (g1872) & (!g1874)) + ((!g4) & (g2) & (!g1841) & (g1872) & (g1874)) + ((!g4) & (g2) & (g1841) & (!g1872) & (!g1874)) + ((!g4) & (g2) & (g1841) & (!g1872) & (g1874)) + ((!g4) & (g2) & (g1841) & (g1872) & (!g1874)) + ((!g4) & (g2) & (g1841) & (g1872) & (g1874)) + ((g4) & (!g2) & (g1841) & (g1872) & (g1874)) + ((g4) & (g2) & (!g1841) & (g1872) & (g1874)) + ((g4) & (g2) & (g1841) & (!g1872) & (g1874)) + ((g4) & (g2) & (g1841) & (g1872) & (g1874)));
	assign g1876 = (((!g4) & (!g1785) & (g1786)) + ((!g4) & (g1785) & (!g1786)) + ((!g4) & (g1785) & (g1786)) + ((g4) & (g1785) & (g1786)));
	assign g1877 = (((!g1759) & (!g1876) & (!g1758) & (!g1788)) + ((!g1759) & (!g1876) & (g1758) & (!g1788)) + ((!g1759) & (!g1876) & (g1758) & (g1788)) + ((g1759) & (g1876) & (!g1758) & (!g1788)) + ((g1759) & (g1876) & (!g1758) & (g1788)) + ((g1759) & (g1876) & (g1758) & (!g1788)) + ((g1759) & (g1876) & (g1758) & (g1788)));
	assign g1878 = (((!g1) & (g1759) & (!g1876) & (!g1758) & (g1788)) + ((!g1) & (g1759) & (g1876) & (!g1758) & (g1788)) + ((g1) & (!g1759) & (g1876) & (g1758) & (!g1788)) + ((g1) & (!g1759) & (g1876) & (g1758) & (g1788)) + ((g1) & (g1759) & (!g1876) & (!g1758) & (!g1788)) + ((g1) & (g1759) & (!g1876) & (!g1758) & (g1788)) + ((g1) & (g1759) & (!g1876) & (g1758) & (!g1788)) + ((g1) & (g1759) & (!g1876) & (g1758) & (g1788)) + ((g1) & (g1759) & (g1876) & (!g1758) & (g1788)));
	assign g1879 = (((!g1) & (!g1840) & (!g1875) & (!g1877) & (!g1878)) + ((g1) & (!g1840) & (!g1875) & (!g1877) & (!g1878)) + ((g1) & (!g1840) & (!g1875) & (g1877) & (!g1878)) + ((g1) & (!g1840) & (g1875) & (!g1877) & (!g1878)) + ((g1) & (!g1840) & (g1875) & (g1877) & (!g1878)) + ((g1) & (g1840) & (!g1875) & (!g1877) & (!g1878)) + ((g1) & (g1840) & (!g1875) & (g1877) & (!g1878)));
	assign g1880 = (((!g319) & (!g1789) & (g1839) & (!g1879)) + ((!g319) & (g1789) & (!g1839) & (!g1879)) + ((!g319) & (g1789) & (!g1839) & (g1879)) + ((!g319) & (g1789) & (g1839) & (g1879)) + ((g319) & (!g1789) & (!g1839) & (!g1879)) + ((g319) & (g1789) & (!g1839) & (g1879)) + ((g319) & (g1789) & (g1839) & (!g1879)) + ((g319) & (g1789) & (g1839) & (g1879)));
	assign g1881 = (((!g358) & (!g390) & (!g1791) & (g1792) & (g1838) & (!g1879)) + ((!g358) & (!g390) & (g1791) & (!g1792) & (!g1838) & (!g1879)) + ((!g358) & (!g390) & (g1791) & (!g1792) & (!g1838) & (g1879)) + ((!g358) & (!g390) & (g1791) & (!g1792) & (g1838) & (!g1879)) + ((!g358) & (!g390) & (g1791) & (!g1792) & (g1838) & (g1879)) + ((!g358) & (!g390) & (g1791) & (g1792) & (!g1838) & (!g1879)) + ((!g358) & (!g390) & (g1791) & (g1792) & (!g1838) & (g1879)) + ((!g358) & (!g390) & (g1791) & (g1792) & (g1838) & (g1879)) + ((!g358) & (g390) & (!g1791) & (!g1792) & (g1838) & (!g1879)) + ((!g358) & (g390) & (!g1791) & (g1792) & (!g1838) & (!g1879)) + ((!g358) & (g390) & (!g1791) & (g1792) & (g1838) & (!g1879)) + ((!g358) & (g390) & (g1791) & (!g1792) & (!g1838) & (!g1879)) + ((!g358) & (g390) & (g1791) & (!g1792) & (!g1838) & (g1879)) + ((!g358) & (g390) & (g1791) & (!g1792) & (g1838) & (g1879)) + ((!g358) & (g390) & (g1791) & (g1792) & (!g1838) & (g1879)) + ((!g358) & (g390) & (g1791) & (g1792) & (g1838) & (g1879)) + ((g358) & (!g390) & (!g1791) & (!g1792) & (!g1838) & (!g1879)) + ((g358) & (!g390) & (!g1791) & (!g1792) & (g1838) & (!g1879)) + ((g358) & (!g390) & (!g1791) & (g1792) & (!g1838) & (!g1879)) + ((g358) & (!g390) & (g1791) & (!g1792) & (!g1838) & (g1879)) + ((g358) & (!g390) & (g1791) & (!g1792) & (g1838) & (g1879)) + ((g358) & (!g390) & (g1791) & (g1792) & (!g1838) & (g1879)) + ((g358) & (!g390) & (g1791) & (g1792) & (g1838) & (!g1879)) + ((g358) & (!g390) & (g1791) & (g1792) & (g1838) & (g1879)) + ((g358) & (g390) & (!g1791) & (!g1792) & (!g1838) & (!g1879)) + ((g358) & (g390) & (g1791) & (!g1792) & (!g1838) & (g1879)) + ((g358) & (g390) & (g1791) & (!g1792) & (g1838) & (!g1879)) + ((g358) & (g390) & (g1791) & (!g1792) & (g1838) & (g1879)) + ((g358) & (g390) & (g1791) & (g1792) & (!g1838) & (!g1879)) + ((g358) & (g390) & (g1791) & (g1792) & (!g1838) & (g1879)) + ((g358) & (g390) & (g1791) & (g1792) & (g1838) & (!g1879)) + ((g358) & (g390) & (g1791) & (g1792) & (g1838) & (g1879)));
	assign g1882 = (((!g390) & (!g1792) & (g1838) & (!g1879)) + ((!g390) & (g1792) & (!g1838) & (!g1879)) + ((!g390) & (g1792) & (!g1838) & (g1879)) + ((!g390) & (g1792) & (g1838) & (g1879)) + ((g390) & (!g1792) & (!g1838) & (!g1879)) + ((g390) & (g1792) & (!g1838) & (g1879)) + ((g390) & (g1792) & (g1838) & (!g1879)) + ((g390) & (g1792) & (g1838) & (g1879)));
	assign g1883 = (((!g433) & (!g468) & (!g1794) & (g1795) & (g1837) & (!g1879)) + ((!g433) & (!g468) & (g1794) & (!g1795) & (!g1837) & (!g1879)) + ((!g433) & (!g468) & (g1794) & (!g1795) & (!g1837) & (g1879)) + ((!g433) & (!g468) & (g1794) & (!g1795) & (g1837) & (!g1879)) + ((!g433) & (!g468) & (g1794) & (!g1795) & (g1837) & (g1879)) + ((!g433) & (!g468) & (g1794) & (g1795) & (!g1837) & (!g1879)) + ((!g433) & (!g468) & (g1794) & (g1795) & (!g1837) & (g1879)) + ((!g433) & (!g468) & (g1794) & (g1795) & (g1837) & (g1879)) + ((!g433) & (g468) & (!g1794) & (!g1795) & (g1837) & (!g1879)) + ((!g433) & (g468) & (!g1794) & (g1795) & (!g1837) & (!g1879)) + ((!g433) & (g468) & (!g1794) & (g1795) & (g1837) & (!g1879)) + ((!g433) & (g468) & (g1794) & (!g1795) & (!g1837) & (!g1879)) + ((!g433) & (g468) & (g1794) & (!g1795) & (!g1837) & (g1879)) + ((!g433) & (g468) & (g1794) & (!g1795) & (g1837) & (g1879)) + ((!g433) & (g468) & (g1794) & (g1795) & (!g1837) & (g1879)) + ((!g433) & (g468) & (g1794) & (g1795) & (g1837) & (g1879)) + ((g433) & (!g468) & (!g1794) & (!g1795) & (!g1837) & (!g1879)) + ((g433) & (!g468) & (!g1794) & (!g1795) & (g1837) & (!g1879)) + ((g433) & (!g468) & (!g1794) & (g1795) & (!g1837) & (!g1879)) + ((g433) & (!g468) & (g1794) & (!g1795) & (!g1837) & (g1879)) + ((g433) & (!g468) & (g1794) & (!g1795) & (g1837) & (g1879)) + ((g433) & (!g468) & (g1794) & (g1795) & (!g1837) & (g1879)) + ((g433) & (!g468) & (g1794) & (g1795) & (g1837) & (!g1879)) + ((g433) & (!g468) & (g1794) & (g1795) & (g1837) & (g1879)) + ((g433) & (g468) & (!g1794) & (!g1795) & (!g1837) & (!g1879)) + ((g433) & (g468) & (g1794) & (!g1795) & (!g1837) & (g1879)) + ((g433) & (g468) & (g1794) & (!g1795) & (g1837) & (!g1879)) + ((g433) & (g468) & (g1794) & (!g1795) & (g1837) & (g1879)) + ((g433) & (g468) & (g1794) & (g1795) & (!g1837) & (!g1879)) + ((g433) & (g468) & (g1794) & (g1795) & (!g1837) & (g1879)) + ((g433) & (g468) & (g1794) & (g1795) & (g1837) & (!g1879)) + ((g433) & (g468) & (g1794) & (g1795) & (g1837) & (g1879)));
	assign g1884 = (((!g468) & (!g1795) & (g1837) & (!g1879)) + ((!g468) & (g1795) & (!g1837) & (!g1879)) + ((!g468) & (g1795) & (!g1837) & (g1879)) + ((!g468) & (g1795) & (g1837) & (g1879)) + ((g468) & (!g1795) & (!g1837) & (!g1879)) + ((g468) & (g1795) & (!g1837) & (g1879)) + ((g468) & (g1795) & (g1837) & (!g1879)) + ((g468) & (g1795) & (g1837) & (g1879)));
	assign g1885 = (((!g515) & (!g553) & (!g1797) & (g1798) & (g1836) & (!g1879)) + ((!g515) & (!g553) & (g1797) & (!g1798) & (!g1836) & (!g1879)) + ((!g515) & (!g553) & (g1797) & (!g1798) & (!g1836) & (g1879)) + ((!g515) & (!g553) & (g1797) & (!g1798) & (g1836) & (!g1879)) + ((!g515) & (!g553) & (g1797) & (!g1798) & (g1836) & (g1879)) + ((!g515) & (!g553) & (g1797) & (g1798) & (!g1836) & (!g1879)) + ((!g515) & (!g553) & (g1797) & (g1798) & (!g1836) & (g1879)) + ((!g515) & (!g553) & (g1797) & (g1798) & (g1836) & (g1879)) + ((!g515) & (g553) & (!g1797) & (!g1798) & (g1836) & (!g1879)) + ((!g515) & (g553) & (!g1797) & (g1798) & (!g1836) & (!g1879)) + ((!g515) & (g553) & (!g1797) & (g1798) & (g1836) & (!g1879)) + ((!g515) & (g553) & (g1797) & (!g1798) & (!g1836) & (!g1879)) + ((!g515) & (g553) & (g1797) & (!g1798) & (!g1836) & (g1879)) + ((!g515) & (g553) & (g1797) & (!g1798) & (g1836) & (g1879)) + ((!g515) & (g553) & (g1797) & (g1798) & (!g1836) & (g1879)) + ((!g515) & (g553) & (g1797) & (g1798) & (g1836) & (g1879)) + ((g515) & (!g553) & (!g1797) & (!g1798) & (!g1836) & (!g1879)) + ((g515) & (!g553) & (!g1797) & (!g1798) & (g1836) & (!g1879)) + ((g515) & (!g553) & (!g1797) & (g1798) & (!g1836) & (!g1879)) + ((g515) & (!g553) & (g1797) & (!g1798) & (!g1836) & (g1879)) + ((g515) & (!g553) & (g1797) & (!g1798) & (g1836) & (g1879)) + ((g515) & (!g553) & (g1797) & (g1798) & (!g1836) & (g1879)) + ((g515) & (!g553) & (g1797) & (g1798) & (g1836) & (!g1879)) + ((g515) & (!g553) & (g1797) & (g1798) & (g1836) & (g1879)) + ((g515) & (g553) & (!g1797) & (!g1798) & (!g1836) & (!g1879)) + ((g515) & (g553) & (g1797) & (!g1798) & (!g1836) & (g1879)) + ((g515) & (g553) & (g1797) & (!g1798) & (g1836) & (!g1879)) + ((g515) & (g553) & (g1797) & (!g1798) & (g1836) & (g1879)) + ((g515) & (g553) & (g1797) & (g1798) & (!g1836) & (!g1879)) + ((g515) & (g553) & (g1797) & (g1798) & (!g1836) & (g1879)) + ((g515) & (g553) & (g1797) & (g1798) & (g1836) & (!g1879)) + ((g515) & (g553) & (g1797) & (g1798) & (g1836) & (g1879)));
	assign g1886 = (((!g553) & (!g1798) & (g1836) & (!g1879)) + ((!g553) & (g1798) & (!g1836) & (!g1879)) + ((!g553) & (g1798) & (!g1836) & (g1879)) + ((!g553) & (g1798) & (g1836) & (g1879)) + ((g553) & (!g1798) & (!g1836) & (!g1879)) + ((g553) & (g1798) & (!g1836) & (g1879)) + ((g553) & (g1798) & (g1836) & (!g1879)) + ((g553) & (g1798) & (g1836) & (g1879)));
	assign g1887 = (((!g604) & (!g645) & (!g1800) & (g1801) & (g1835) & (!g1879)) + ((!g604) & (!g645) & (g1800) & (!g1801) & (!g1835) & (!g1879)) + ((!g604) & (!g645) & (g1800) & (!g1801) & (!g1835) & (g1879)) + ((!g604) & (!g645) & (g1800) & (!g1801) & (g1835) & (!g1879)) + ((!g604) & (!g645) & (g1800) & (!g1801) & (g1835) & (g1879)) + ((!g604) & (!g645) & (g1800) & (g1801) & (!g1835) & (!g1879)) + ((!g604) & (!g645) & (g1800) & (g1801) & (!g1835) & (g1879)) + ((!g604) & (!g645) & (g1800) & (g1801) & (g1835) & (g1879)) + ((!g604) & (g645) & (!g1800) & (!g1801) & (g1835) & (!g1879)) + ((!g604) & (g645) & (!g1800) & (g1801) & (!g1835) & (!g1879)) + ((!g604) & (g645) & (!g1800) & (g1801) & (g1835) & (!g1879)) + ((!g604) & (g645) & (g1800) & (!g1801) & (!g1835) & (!g1879)) + ((!g604) & (g645) & (g1800) & (!g1801) & (!g1835) & (g1879)) + ((!g604) & (g645) & (g1800) & (!g1801) & (g1835) & (g1879)) + ((!g604) & (g645) & (g1800) & (g1801) & (!g1835) & (g1879)) + ((!g604) & (g645) & (g1800) & (g1801) & (g1835) & (g1879)) + ((g604) & (!g645) & (!g1800) & (!g1801) & (!g1835) & (!g1879)) + ((g604) & (!g645) & (!g1800) & (!g1801) & (g1835) & (!g1879)) + ((g604) & (!g645) & (!g1800) & (g1801) & (!g1835) & (!g1879)) + ((g604) & (!g645) & (g1800) & (!g1801) & (!g1835) & (g1879)) + ((g604) & (!g645) & (g1800) & (!g1801) & (g1835) & (g1879)) + ((g604) & (!g645) & (g1800) & (g1801) & (!g1835) & (g1879)) + ((g604) & (!g645) & (g1800) & (g1801) & (g1835) & (!g1879)) + ((g604) & (!g645) & (g1800) & (g1801) & (g1835) & (g1879)) + ((g604) & (g645) & (!g1800) & (!g1801) & (!g1835) & (!g1879)) + ((g604) & (g645) & (g1800) & (!g1801) & (!g1835) & (g1879)) + ((g604) & (g645) & (g1800) & (!g1801) & (g1835) & (!g1879)) + ((g604) & (g645) & (g1800) & (!g1801) & (g1835) & (g1879)) + ((g604) & (g645) & (g1800) & (g1801) & (!g1835) & (!g1879)) + ((g604) & (g645) & (g1800) & (g1801) & (!g1835) & (g1879)) + ((g604) & (g645) & (g1800) & (g1801) & (g1835) & (!g1879)) + ((g604) & (g645) & (g1800) & (g1801) & (g1835) & (g1879)));
	assign g1888 = (((!g645) & (!g1801) & (g1835) & (!g1879)) + ((!g645) & (g1801) & (!g1835) & (!g1879)) + ((!g645) & (g1801) & (!g1835) & (g1879)) + ((!g645) & (g1801) & (g1835) & (g1879)) + ((g645) & (!g1801) & (!g1835) & (!g1879)) + ((g645) & (g1801) & (!g1835) & (g1879)) + ((g645) & (g1801) & (g1835) & (!g1879)) + ((g645) & (g1801) & (g1835) & (g1879)));
	assign g1889 = (((!g700) & (!g744) & (!g1803) & (g1804) & (g1834) & (!g1879)) + ((!g700) & (!g744) & (g1803) & (!g1804) & (!g1834) & (!g1879)) + ((!g700) & (!g744) & (g1803) & (!g1804) & (!g1834) & (g1879)) + ((!g700) & (!g744) & (g1803) & (!g1804) & (g1834) & (!g1879)) + ((!g700) & (!g744) & (g1803) & (!g1804) & (g1834) & (g1879)) + ((!g700) & (!g744) & (g1803) & (g1804) & (!g1834) & (!g1879)) + ((!g700) & (!g744) & (g1803) & (g1804) & (!g1834) & (g1879)) + ((!g700) & (!g744) & (g1803) & (g1804) & (g1834) & (g1879)) + ((!g700) & (g744) & (!g1803) & (!g1804) & (g1834) & (!g1879)) + ((!g700) & (g744) & (!g1803) & (g1804) & (!g1834) & (!g1879)) + ((!g700) & (g744) & (!g1803) & (g1804) & (g1834) & (!g1879)) + ((!g700) & (g744) & (g1803) & (!g1804) & (!g1834) & (!g1879)) + ((!g700) & (g744) & (g1803) & (!g1804) & (!g1834) & (g1879)) + ((!g700) & (g744) & (g1803) & (!g1804) & (g1834) & (g1879)) + ((!g700) & (g744) & (g1803) & (g1804) & (!g1834) & (g1879)) + ((!g700) & (g744) & (g1803) & (g1804) & (g1834) & (g1879)) + ((g700) & (!g744) & (!g1803) & (!g1804) & (!g1834) & (!g1879)) + ((g700) & (!g744) & (!g1803) & (!g1804) & (g1834) & (!g1879)) + ((g700) & (!g744) & (!g1803) & (g1804) & (!g1834) & (!g1879)) + ((g700) & (!g744) & (g1803) & (!g1804) & (!g1834) & (g1879)) + ((g700) & (!g744) & (g1803) & (!g1804) & (g1834) & (g1879)) + ((g700) & (!g744) & (g1803) & (g1804) & (!g1834) & (g1879)) + ((g700) & (!g744) & (g1803) & (g1804) & (g1834) & (!g1879)) + ((g700) & (!g744) & (g1803) & (g1804) & (g1834) & (g1879)) + ((g700) & (g744) & (!g1803) & (!g1804) & (!g1834) & (!g1879)) + ((g700) & (g744) & (g1803) & (!g1804) & (!g1834) & (g1879)) + ((g700) & (g744) & (g1803) & (!g1804) & (g1834) & (!g1879)) + ((g700) & (g744) & (g1803) & (!g1804) & (g1834) & (g1879)) + ((g700) & (g744) & (g1803) & (g1804) & (!g1834) & (!g1879)) + ((g700) & (g744) & (g1803) & (g1804) & (!g1834) & (g1879)) + ((g700) & (g744) & (g1803) & (g1804) & (g1834) & (!g1879)) + ((g700) & (g744) & (g1803) & (g1804) & (g1834) & (g1879)));
	assign g1890 = (((!g744) & (!g1804) & (g1834) & (!g1879)) + ((!g744) & (g1804) & (!g1834) & (!g1879)) + ((!g744) & (g1804) & (!g1834) & (g1879)) + ((!g744) & (g1804) & (g1834) & (g1879)) + ((g744) & (!g1804) & (!g1834) & (!g1879)) + ((g744) & (g1804) & (!g1834) & (g1879)) + ((g744) & (g1804) & (g1834) & (!g1879)) + ((g744) & (g1804) & (g1834) & (g1879)));
	assign g1891 = (((!g803) & (!g851) & (!g1806) & (g1807) & (g1833) & (!g1879)) + ((!g803) & (!g851) & (g1806) & (!g1807) & (!g1833) & (!g1879)) + ((!g803) & (!g851) & (g1806) & (!g1807) & (!g1833) & (g1879)) + ((!g803) & (!g851) & (g1806) & (!g1807) & (g1833) & (!g1879)) + ((!g803) & (!g851) & (g1806) & (!g1807) & (g1833) & (g1879)) + ((!g803) & (!g851) & (g1806) & (g1807) & (!g1833) & (!g1879)) + ((!g803) & (!g851) & (g1806) & (g1807) & (!g1833) & (g1879)) + ((!g803) & (!g851) & (g1806) & (g1807) & (g1833) & (g1879)) + ((!g803) & (g851) & (!g1806) & (!g1807) & (g1833) & (!g1879)) + ((!g803) & (g851) & (!g1806) & (g1807) & (!g1833) & (!g1879)) + ((!g803) & (g851) & (!g1806) & (g1807) & (g1833) & (!g1879)) + ((!g803) & (g851) & (g1806) & (!g1807) & (!g1833) & (!g1879)) + ((!g803) & (g851) & (g1806) & (!g1807) & (!g1833) & (g1879)) + ((!g803) & (g851) & (g1806) & (!g1807) & (g1833) & (g1879)) + ((!g803) & (g851) & (g1806) & (g1807) & (!g1833) & (g1879)) + ((!g803) & (g851) & (g1806) & (g1807) & (g1833) & (g1879)) + ((g803) & (!g851) & (!g1806) & (!g1807) & (!g1833) & (!g1879)) + ((g803) & (!g851) & (!g1806) & (!g1807) & (g1833) & (!g1879)) + ((g803) & (!g851) & (!g1806) & (g1807) & (!g1833) & (!g1879)) + ((g803) & (!g851) & (g1806) & (!g1807) & (!g1833) & (g1879)) + ((g803) & (!g851) & (g1806) & (!g1807) & (g1833) & (g1879)) + ((g803) & (!g851) & (g1806) & (g1807) & (!g1833) & (g1879)) + ((g803) & (!g851) & (g1806) & (g1807) & (g1833) & (!g1879)) + ((g803) & (!g851) & (g1806) & (g1807) & (g1833) & (g1879)) + ((g803) & (g851) & (!g1806) & (!g1807) & (!g1833) & (!g1879)) + ((g803) & (g851) & (g1806) & (!g1807) & (!g1833) & (g1879)) + ((g803) & (g851) & (g1806) & (!g1807) & (g1833) & (!g1879)) + ((g803) & (g851) & (g1806) & (!g1807) & (g1833) & (g1879)) + ((g803) & (g851) & (g1806) & (g1807) & (!g1833) & (!g1879)) + ((g803) & (g851) & (g1806) & (g1807) & (!g1833) & (g1879)) + ((g803) & (g851) & (g1806) & (g1807) & (g1833) & (!g1879)) + ((g803) & (g851) & (g1806) & (g1807) & (g1833) & (g1879)));
	assign g1892 = (((!g851) & (!g1807) & (g1833) & (!g1879)) + ((!g851) & (g1807) & (!g1833) & (!g1879)) + ((!g851) & (g1807) & (!g1833) & (g1879)) + ((!g851) & (g1807) & (g1833) & (g1879)) + ((g851) & (!g1807) & (!g1833) & (!g1879)) + ((g851) & (g1807) & (!g1833) & (g1879)) + ((g851) & (g1807) & (g1833) & (!g1879)) + ((g851) & (g1807) & (g1833) & (g1879)));
	assign g1893 = (((!g914) & (!g1032) & (!g1809) & (g1810) & (g1832) & (!g1879)) + ((!g914) & (!g1032) & (g1809) & (!g1810) & (!g1832) & (!g1879)) + ((!g914) & (!g1032) & (g1809) & (!g1810) & (!g1832) & (g1879)) + ((!g914) & (!g1032) & (g1809) & (!g1810) & (g1832) & (!g1879)) + ((!g914) & (!g1032) & (g1809) & (!g1810) & (g1832) & (g1879)) + ((!g914) & (!g1032) & (g1809) & (g1810) & (!g1832) & (!g1879)) + ((!g914) & (!g1032) & (g1809) & (g1810) & (!g1832) & (g1879)) + ((!g914) & (!g1032) & (g1809) & (g1810) & (g1832) & (g1879)) + ((!g914) & (g1032) & (!g1809) & (!g1810) & (g1832) & (!g1879)) + ((!g914) & (g1032) & (!g1809) & (g1810) & (!g1832) & (!g1879)) + ((!g914) & (g1032) & (!g1809) & (g1810) & (g1832) & (!g1879)) + ((!g914) & (g1032) & (g1809) & (!g1810) & (!g1832) & (!g1879)) + ((!g914) & (g1032) & (g1809) & (!g1810) & (!g1832) & (g1879)) + ((!g914) & (g1032) & (g1809) & (!g1810) & (g1832) & (g1879)) + ((!g914) & (g1032) & (g1809) & (g1810) & (!g1832) & (g1879)) + ((!g914) & (g1032) & (g1809) & (g1810) & (g1832) & (g1879)) + ((g914) & (!g1032) & (!g1809) & (!g1810) & (!g1832) & (!g1879)) + ((g914) & (!g1032) & (!g1809) & (!g1810) & (g1832) & (!g1879)) + ((g914) & (!g1032) & (!g1809) & (g1810) & (!g1832) & (!g1879)) + ((g914) & (!g1032) & (g1809) & (!g1810) & (!g1832) & (g1879)) + ((g914) & (!g1032) & (g1809) & (!g1810) & (g1832) & (g1879)) + ((g914) & (!g1032) & (g1809) & (g1810) & (!g1832) & (g1879)) + ((g914) & (!g1032) & (g1809) & (g1810) & (g1832) & (!g1879)) + ((g914) & (!g1032) & (g1809) & (g1810) & (g1832) & (g1879)) + ((g914) & (g1032) & (!g1809) & (!g1810) & (!g1832) & (!g1879)) + ((g914) & (g1032) & (g1809) & (!g1810) & (!g1832) & (g1879)) + ((g914) & (g1032) & (g1809) & (!g1810) & (g1832) & (!g1879)) + ((g914) & (g1032) & (g1809) & (!g1810) & (g1832) & (g1879)) + ((g914) & (g1032) & (g1809) & (g1810) & (!g1832) & (!g1879)) + ((g914) & (g1032) & (g1809) & (g1810) & (!g1832) & (g1879)) + ((g914) & (g1032) & (g1809) & (g1810) & (g1832) & (!g1879)) + ((g914) & (g1032) & (g1809) & (g1810) & (g1832) & (g1879)));
	assign g1894 = (((!g1032) & (!g1810) & (g1832) & (!g1879)) + ((!g1032) & (g1810) & (!g1832) & (!g1879)) + ((!g1032) & (g1810) & (!g1832) & (g1879)) + ((!g1032) & (g1810) & (g1832) & (g1879)) + ((g1032) & (!g1810) & (!g1832) & (!g1879)) + ((g1032) & (g1810) & (!g1832) & (g1879)) + ((g1032) & (g1810) & (g1832) & (!g1879)) + ((g1032) & (g1810) & (g1832) & (g1879)));
	assign g1895 = (((!g1030) & (!g1160) & (!g1812) & (g1813) & (g1831) & (!g1879)) + ((!g1030) & (!g1160) & (g1812) & (!g1813) & (!g1831) & (!g1879)) + ((!g1030) & (!g1160) & (g1812) & (!g1813) & (!g1831) & (g1879)) + ((!g1030) & (!g1160) & (g1812) & (!g1813) & (g1831) & (!g1879)) + ((!g1030) & (!g1160) & (g1812) & (!g1813) & (g1831) & (g1879)) + ((!g1030) & (!g1160) & (g1812) & (g1813) & (!g1831) & (!g1879)) + ((!g1030) & (!g1160) & (g1812) & (g1813) & (!g1831) & (g1879)) + ((!g1030) & (!g1160) & (g1812) & (g1813) & (g1831) & (g1879)) + ((!g1030) & (g1160) & (!g1812) & (!g1813) & (g1831) & (!g1879)) + ((!g1030) & (g1160) & (!g1812) & (g1813) & (!g1831) & (!g1879)) + ((!g1030) & (g1160) & (!g1812) & (g1813) & (g1831) & (!g1879)) + ((!g1030) & (g1160) & (g1812) & (!g1813) & (!g1831) & (!g1879)) + ((!g1030) & (g1160) & (g1812) & (!g1813) & (!g1831) & (g1879)) + ((!g1030) & (g1160) & (g1812) & (!g1813) & (g1831) & (g1879)) + ((!g1030) & (g1160) & (g1812) & (g1813) & (!g1831) & (g1879)) + ((!g1030) & (g1160) & (g1812) & (g1813) & (g1831) & (g1879)) + ((g1030) & (!g1160) & (!g1812) & (!g1813) & (!g1831) & (!g1879)) + ((g1030) & (!g1160) & (!g1812) & (!g1813) & (g1831) & (!g1879)) + ((g1030) & (!g1160) & (!g1812) & (g1813) & (!g1831) & (!g1879)) + ((g1030) & (!g1160) & (g1812) & (!g1813) & (!g1831) & (g1879)) + ((g1030) & (!g1160) & (g1812) & (!g1813) & (g1831) & (g1879)) + ((g1030) & (!g1160) & (g1812) & (g1813) & (!g1831) & (g1879)) + ((g1030) & (!g1160) & (g1812) & (g1813) & (g1831) & (!g1879)) + ((g1030) & (!g1160) & (g1812) & (g1813) & (g1831) & (g1879)) + ((g1030) & (g1160) & (!g1812) & (!g1813) & (!g1831) & (!g1879)) + ((g1030) & (g1160) & (g1812) & (!g1813) & (!g1831) & (g1879)) + ((g1030) & (g1160) & (g1812) & (!g1813) & (g1831) & (!g1879)) + ((g1030) & (g1160) & (g1812) & (!g1813) & (g1831) & (g1879)) + ((g1030) & (g1160) & (g1812) & (g1813) & (!g1831) & (!g1879)) + ((g1030) & (g1160) & (g1812) & (g1813) & (!g1831) & (g1879)) + ((g1030) & (g1160) & (g1812) & (g1813) & (g1831) & (!g1879)) + ((g1030) & (g1160) & (g1812) & (g1813) & (g1831) & (g1879)));
	assign g1896 = (((!g1160) & (!g1813) & (g1831) & (!g1879)) + ((!g1160) & (g1813) & (!g1831) & (!g1879)) + ((!g1160) & (g1813) & (!g1831) & (g1879)) + ((!g1160) & (g1813) & (g1831) & (g1879)) + ((g1160) & (!g1813) & (!g1831) & (!g1879)) + ((g1160) & (g1813) & (!g1831) & (g1879)) + ((g1160) & (g1813) & (g1831) & (!g1879)) + ((g1160) & (g1813) & (g1831) & (g1879)));
	assign g1897 = (((!g1154) & (!g1295) & (!g1815) & (g1816) & (g1830) & (!g1879)) + ((!g1154) & (!g1295) & (g1815) & (!g1816) & (!g1830) & (!g1879)) + ((!g1154) & (!g1295) & (g1815) & (!g1816) & (!g1830) & (g1879)) + ((!g1154) & (!g1295) & (g1815) & (!g1816) & (g1830) & (!g1879)) + ((!g1154) & (!g1295) & (g1815) & (!g1816) & (g1830) & (g1879)) + ((!g1154) & (!g1295) & (g1815) & (g1816) & (!g1830) & (!g1879)) + ((!g1154) & (!g1295) & (g1815) & (g1816) & (!g1830) & (g1879)) + ((!g1154) & (!g1295) & (g1815) & (g1816) & (g1830) & (g1879)) + ((!g1154) & (g1295) & (!g1815) & (!g1816) & (g1830) & (!g1879)) + ((!g1154) & (g1295) & (!g1815) & (g1816) & (!g1830) & (!g1879)) + ((!g1154) & (g1295) & (!g1815) & (g1816) & (g1830) & (!g1879)) + ((!g1154) & (g1295) & (g1815) & (!g1816) & (!g1830) & (!g1879)) + ((!g1154) & (g1295) & (g1815) & (!g1816) & (!g1830) & (g1879)) + ((!g1154) & (g1295) & (g1815) & (!g1816) & (g1830) & (g1879)) + ((!g1154) & (g1295) & (g1815) & (g1816) & (!g1830) & (g1879)) + ((!g1154) & (g1295) & (g1815) & (g1816) & (g1830) & (g1879)) + ((g1154) & (!g1295) & (!g1815) & (!g1816) & (!g1830) & (!g1879)) + ((g1154) & (!g1295) & (!g1815) & (!g1816) & (g1830) & (!g1879)) + ((g1154) & (!g1295) & (!g1815) & (g1816) & (!g1830) & (!g1879)) + ((g1154) & (!g1295) & (g1815) & (!g1816) & (!g1830) & (g1879)) + ((g1154) & (!g1295) & (g1815) & (!g1816) & (g1830) & (g1879)) + ((g1154) & (!g1295) & (g1815) & (g1816) & (!g1830) & (g1879)) + ((g1154) & (!g1295) & (g1815) & (g1816) & (g1830) & (!g1879)) + ((g1154) & (!g1295) & (g1815) & (g1816) & (g1830) & (g1879)) + ((g1154) & (g1295) & (!g1815) & (!g1816) & (!g1830) & (!g1879)) + ((g1154) & (g1295) & (g1815) & (!g1816) & (!g1830) & (g1879)) + ((g1154) & (g1295) & (g1815) & (!g1816) & (g1830) & (!g1879)) + ((g1154) & (g1295) & (g1815) & (!g1816) & (g1830) & (g1879)) + ((g1154) & (g1295) & (g1815) & (g1816) & (!g1830) & (!g1879)) + ((g1154) & (g1295) & (g1815) & (g1816) & (!g1830) & (g1879)) + ((g1154) & (g1295) & (g1815) & (g1816) & (g1830) & (!g1879)) + ((g1154) & (g1295) & (g1815) & (g1816) & (g1830) & (g1879)));
	assign g1898 = (((!g1295) & (!g1816) & (g1830) & (!g1879)) + ((!g1295) & (g1816) & (!g1830) & (!g1879)) + ((!g1295) & (g1816) & (!g1830) & (g1879)) + ((!g1295) & (g1816) & (g1830) & (g1879)) + ((g1295) & (!g1816) & (!g1830) & (!g1879)) + ((g1295) & (g1816) & (!g1830) & (g1879)) + ((g1295) & (g1816) & (g1830) & (!g1879)) + ((g1295) & (g1816) & (g1830) & (g1879)));
	assign g1899 = (((!g1285) & (!g1437) & (!g1818) & (g1819) & (g1829) & (!g1879)) + ((!g1285) & (!g1437) & (g1818) & (!g1819) & (!g1829) & (!g1879)) + ((!g1285) & (!g1437) & (g1818) & (!g1819) & (!g1829) & (g1879)) + ((!g1285) & (!g1437) & (g1818) & (!g1819) & (g1829) & (!g1879)) + ((!g1285) & (!g1437) & (g1818) & (!g1819) & (g1829) & (g1879)) + ((!g1285) & (!g1437) & (g1818) & (g1819) & (!g1829) & (!g1879)) + ((!g1285) & (!g1437) & (g1818) & (g1819) & (!g1829) & (g1879)) + ((!g1285) & (!g1437) & (g1818) & (g1819) & (g1829) & (g1879)) + ((!g1285) & (g1437) & (!g1818) & (!g1819) & (g1829) & (!g1879)) + ((!g1285) & (g1437) & (!g1818) & (g1819) & (!g1829) & (!g1879)) + ((!g1285) & (g1437) & (!g1818) & (g1819) & (g1829) & (!g1879)) + ((!g1285) & (g1437) & (g1818) & (!g1819) & (!g1829) & (!g1879)) + ((!g1285) & (g1437) & (g1818) & (!g1819) & (!g1829) & (g1879)) + ((!g1285) & (g1437) & (g1818) & (!g1819) & (g1829) & (g1879)) + ((!g1285) & (g1437) & (g1818) & (g1819) & (!g1829) & (g1879)) + ((!g1285) & (g1437) & (g1818) & (g1819) & (g1829) & (g1879)) + ((g1285) & (!g1437) & (!g1818) & (!g1819) & (!g1829) & (!g1879)) + ((g1285) & (!g1437) & (!g1818) & (!g1819) & (g1829) & (!g1879)) + ((g1285) & (!g1437) & (!g1818) & (g1819) & (!g1829) & (!g1879)) + ((g1285) & (!g1437) & (g1818) & (!g1819) & (!g1829) & (g1879)) + ((g1285) & (!g1437) & (g1818) & (!g1819) & (g1829) & (g1879)) + ((g1285) & (!g1437) & (g1818) & (g1819) & (!g1829) & (g1879)) + ((g1285) & (!g1437) & (g1818) & (g1819) & (g1829) & (!g1879)) + ((g1285) & (!g1437) & (g1818) & (g1819) & (g1829) & (g1879)) + ((g1285) & (g1437) & (!g1818) & (!g1819) & (!g1829) & (!g1879)) + ((g1285) & (g1437) & (g1818) & (!g1819) & (!g1829) & (g1879)) + ((g1285) & (g1437) & (g1818) & (!g1819) & (g1829) & (!g1879)) + ((g1285) & (g1437) & (g1818) & (!g1819) & (g1829) & (g1879)) + ((g1285) & (g1437) & (g1818) & (g1819) & (!g1829) & (!g1879)) + ((g1285) & (g1437) & (g1818) & (g1819) & (!g1829) & (g1879)) + ((g1285) & (g1437) & (g1818) & (g1819) & (g1829) & (!g1879)) + ((g1285) & (g1437) & (g1818) & (g1819) & (g1829) & (g1879)));
	assign g1900 = (((!g1437) & (!g1819) & (g1829) & (!g1879)) + ((!g1437) & (g1819) & (!g1829) & (!g1879)) + ((!g1437) & (g1819) & (!g1829) & (g1879)) + ((!g1437) & (g1819) & (g1829) & (g1879)) + ((g1437) & (!g1819) & (!g1829) & (!g1879)) + ((g1437) & (g1819) & (!g1829) & (g1879)) + ((g1437) & (g1819) & (g1829) & (!g1879)) + ((g1437) & (g1819) & (g1829) & (g1879)));
	assign g1901 = (((!g1423) & (!g1586) & (!g1821) & (g1822) & (g1828) & (!g1879)) + ((!g1423) & (!g1586) & (g1821) & (!g1822) & (!g1828) & (!g1879)) + ((!g1423) & (!g1586) & (g1821) & (!g1822) & (!g1828) & (g1879)) + ((!g1423) & (!g1586) & (g1821) & (!g1822) & (g1828) & (!g1879)) + ((!g1423) & (!g1586) & (g1821) & (!g1822) & (g1828) & (g1879)) + ((!g1423) & (!g1586) & (g1821) & (g1822) & (!g1828) & (!g1879)) + ((!g1423) & (!g1586) & (g1821) & (g1822) & (!g1828) & (g1879)) + ((!g1423) & (!g1586) & (g1821) & (g1822) & (g1828) & (g1879)) + ((!g1423) & (g1586) & (!g1821) & (!g1822) & (g1828) & (!g1879)) + ((!g1423) & (g1586) & (!g1821) & (g1822) & (!g1828) & (!g1879)) + ((!g1423) & (g1586) & (!g1821) & (g1822) & (g1828) & (!g1879)) + ((!g1423) & (g1586) & (g1821) & (!g1822) & (!g1828) & (!g1879)) + ((!g1423) & (g1586) & (g1821) & (!g1822) & (!g1828) & (g1879)) + ((!g1423) & (g1586) & (g1821) & (!g1822) & (g1828) & (g1879)) + ((!g1423) & (g1586) & (g1821) & (g1822) & (!g1828) & (g1879)) + ((!g1423) & (g1586) & (g1821) & (g1822) & (g1828) & (g1879)) + ((g1423) & (!g1586) & (!g1821) & (!g1822) & (!g1828) & (!g1879)) + ((g1423) & (!g1586) & (!g1821) & (!g1822) & (g1828) & (!g1879)) + ((g1423) & (!g1586) & (!g1821) & (g1822) & (!g1828) & (!g1879)) + ((g1423) & (!g1586) & (g1821) & (!g1822) & (!g1828) & (g1879)) + ((g1423) & (!g1586) & (g1821) & (!g1822) & (g1828) & (g1879)) + ((g1423) & (!g1586) & (g1821) & (g1822) & (!g1828) & (g1879)) + ((g1423) & (!g1586) & (g1821) & (g1822) & (g1828) & (!g1879)) + ((g1423) & (!g1586) & (g1821) & (g1822) & (g1828) & (g1879)) + ((g1423) & (g1586) & (!g1821) & (!g1822) & (!g1828) & (!g1879)) + ((g1423) & (g1586) & (g1821) & (!g1822) & (!g1828) & (g1879)) + ((g1423) & (g1586) & (g1821) & (!g1822) & (g1828) & (!g1879)) + ((g1423) & (g1586) & (g1821) & (!g1822) & (g1828) & (g1879)) + ((g1423) & (g1586) & (g1821) & (g1822) & (!g1828) & (!g1879)) + ((g1423) & (g1586) & (g1821) & (g1822) & (!g1828) & (g1879)) + ((g1423) & (g1586) & (g1821) & (g1822) & (g1828) & (!g1879)) + ((g1423) & (g1586) & (g1821) & (g1822) & (g1828) & (g1879)));
	assign g1902 = (((!g1586) & (!g1822) & (g1828) & (!g1879)) + ((!g1586) & (g1822) & (!g1828) & (!g1879)) + ((!g1586) & (g1822) & (!g1828) & (g1879)) + ((!g1586) & (g1822) & (g1828) & (g1879)) + ((g1586) & (!g1822) & (!g1828) & (!g1879)) + ((g1586) & (g1822) & (!g1828) & (g1879)) + ((g1586) & (g1822) & (g1828) & (!g1879)) + ((g1586) & (g1822) & (g1828) & (g1879)));
	assign g1903 = (((!g1568) & (!g1742) & (!g1824) & (g1825) & (g1827) & (!g1879)) + ((!g1568) & (!g1742) & (g1824) & (!g1825) & (!g1827) & (!g1879)) + ((!g1568) & (!g1742) & (g1824) & (!g1825) & (!g1827) & (g1879)) + ((!g1568) & (!g1742) & (g1824) & (!g1825) & (g1827) & (!g1879)) + ((!g1568) & (!g1742) & (g1824) & (!g1825) & (g1827) & (g1879)) + ((!g1568) & (!g1742) & (g1824) & (g1825) & (!g1827) & (!g1879)) + ((!g1568) & (!g1742) & (g1824) & (g1825) & (!g1827) & (g1879)) + ((!g1568) & (!g1742) & (g1824) & (g1825) & (g1827) & (g1879)) + ((!g1568) & (g1742) & (!g1824) & (!g1825) & (g1827) & (!g1879)) + ((!g1568) & (g1742) & (!g1824) & (g1825) & (!g1827) & (!g1879)) + ((!g1568) & (g1742) & (!g1824) & (g1825) & (g1827) & (!g1879)) + ((!g1568) & (g1742) & (g1824) & (!g1825) & (!g1827) & (!g1879)) + ((!g1568) & (g1742) & (g1824) & (!g1825) & (!g1827) & (g1879)) + ((!g1568) & (g1742) & (g1824) & (!g1825) & (g1827) & (g1879)) + ((!g1568) & (g1742) & (g1824) & (g1825) & (!g1827) & (g1879)) + ((!g1568) & (g1742) & (g1824) & (g1825) & (g1827) & (g1879)) + ((g1568) & (!g1742) & (!g1824) & (!g1825) & (!g1827) & (!g1879)) + ((g1568) & (!g1742) & (!g1824) & (!g1825) & (g1827) & (!g1879)) + ((g1568) & (!g1742) & (!g1824) & (g1825) & (!g1827) & (!g1879)) + ((g1568) & (!g1742) & (g1824) & (!g1825) & (!g1827) & (g1879)) + ((g1568) & (!g1742) & (g1824) & (!g1825) & (g1827) & (g1879)) + ((g1568) & (!g1742) & (g1824) & (g1825) & (!g1827) & (g1879)) + ((g1568) & (!g1742) & (g1824) & (g1825) & (g1827) & (!g1879)) + ((g1568) & (!g1742) & (g1824) & (g1825) & (g1827) & (g1879)) + ((g1568) & (g1742) & (!g1824) & (!g1825) & (!g1827) & (!g1879)) + ((g1568) & (g1742) & (g1824) & (!g1825) & (!g1827) & (g1879)) + ((g1568) & (g1742) & (g1824) & (!g1825) & (g1827) & (!g1879)) + ((g1568) & (g1742) & (g1824) & (!g1825) & (g1827) & (g1879)) + ((g1568) & (g1742) & (g1824) & (g1825) & (!g1827) & (!g1879)) + ((g1568) & (g1742) & (g1824) & (g1825) & (!g1827) & (g1879)) + ((g1568) & (g1742) & (g1824) & (g1825) & (g1827) & (!g1879)) + ((g1568) & (g1742) & (g1824) & (g1825) & (g1827) & (g1879)));
	assign g1904 = (((!g1742) & (!g1825) & (g1827) & (!g1879)) + ((!g1742) & (g1825) & (!g1827) & (!g1879)) + ((!g1742) & (g1825) & (!g1827) & (g1879)) + ((!g1742) & (g1825) & (g1827) & (g1879)) + ((g1742) & (!g1825) & (!g1827) & (!g1879)) + ((g1742) & (g1825) & (!g1827) & (g1879)) + ((g1742) & (g1825) & (g1827) & (!g1879)) + ((g1742) & (g1825) & (g1827) & (g1879)));
	assign g1905 = (((!g1758) & (g1788)));
	assign g1906 = (((!g1720) & (!ax38x) & (!ax39x) & (!g1905) & (!g1826) & (g1879)) + ((!g1720) & (!ax38x) & (!ax39x) & (!g1905) & (g1826) & (!g1879)) + ((!g1720) & (!ax38x) & (!ax39x) & (!g1905) & (g1826) & (g1879)) + ((!g1720) & (!ax38x) & (!ax39x) & (g1905) & (!g1826) & (!g1879)) + ((!g1720) & (!ax38x) & (ax39x) & (!g1905) & (!g1826) & (!g1879)) + ((!g1720) & (!ax38x) & (ax39x) & (g1905) & (!g1826) & (g1879)) + ((!g1720) & (!ax38x) & (ax39x) & (g1905) & (g1826) & (!g1879)) + ((!g1720) & (!ax38x) & (ax39x) & (g1905) & (g1826) & (g1879)) + ((!g1720) & (ax38x) & (!ax39x) & (g1905) & (!g1826) & (!g1879)) + ((!g1720) & (ax38x) & (!ax39x) & (g1905) & (g1826) & (!g1879)) + ((!g1720) & (ax38x) & (ax39x) & (!g1905) & (!g1826) & (!g1879)) + ((!g1720) & (ax38x) & (ax39x) & (!g1905) & (!g1826) & (g1879)) + ((!g1720) & (ax38x) & (ax39x) & (!g1905) & (g1826) & (!g1879)) + ((!g1720) & (ax38x) & (ax39x) & (!g1905) & (g1826) & (g1879)) + ((!g1720) & (ax38x) & (ax39x) & (g1905) & (!g1826) & (g1879)) + ((!g1720) & (ax38x) & (ax39x) & (g1905) & (g1826) & (g1879)) + ((g1720) & (!ax38x) & (!ax39x) & (!g1905) & (!g1826) & (!g1879)) + ((g1720) & (!ax38x) & (!ax39x) & (!g1905) & (!g1826) & (g1879)) + ((g1720) & (!ax38x) & (!ax39x) & (!g1905) & (g1826) & (g1879)) + ((g1720) & (!ax38x) & (!ax39x) & (g1905) & (g1826) & (!g1879)) + ((g1720) & (!ax38x) & (ax39x) & (!g1905) & (g1826) & (!g1879)) + ((g1720) & (!ax38x) & (ax39x) & (g1905) & (!g1826) & (!g1879)) + ((g1720) & (!ax38x) & (ax39x) & (g1905) & (!g1826) & (g1879)) + ((g1720) & (!ax38x) & (ax39x) & (g1905) & (g1826) & (g1879)) + ((g1720) & (ax38x) & (!ax39x) & (!g1905) & (!g1826) & (!g1879)) + ((g1720) & (ax38x) & (!ax39x) & (!g1905) & (g1826) & (!g1879)) + ((g1720) & (ax38x) & (ax39x) & (!g1905) & (!g1826) & (g1879)) + ((g1720) & (ax38x) & (ax39x) & (!g1905) & (g1826) & (g1879)) + ((g1720) & (ax38x) & (ax39x) & (g1905) & (!g1826) & (!g1879)) + ((g1720) & (ax38x) & (ax39x) & (g1905) & (!g1826) & (g1879)) + ((g1720) & (ax38x) & (ax39x) & (g1905) & (g1826) & (!g1879)) + ((g1720) & (ax38x) & (ax39x) & (g1905) & (g1826) & (g1879)));
	assign g1907 = (((!ax38x) & (!g1905) & (!g1826) & (g1879)) + ((!ax38x) & (!g1905) & (g1826) & (!g1879)) + ((!ax38x) & (!g1905) & (g1826) & (g1879)) + ((!ax38x) & (g1905) & (g1826) & (!g1879)) + ((ax38x) & (!g1905) & (!g1826) & (!g1879)) + ((ax38x) & (g1905) & (!g1826) & (!g1879)) + ((ax38x) & (g1905) & (!g1826) & (g1879)) + ((ax38x) & (g1905) & (g1826) & (g1879)));
	assign g1908 = (((!ax34x) & (!ax35x)));
	assign g1909 = (((!g1905) & (!ax36x) & (!ax37x) & (!g1879) & (!g1908)) + ((!g1905) & (!ax36x) & (ax37x) & (g1879) & (!g1908)) + ((!g1905) & (ax36x) & (ax37x) & (g1879) & (!g1908)) + ((!g1905) & (ax36x) & (ax37x) & (g1879) & (g1908)) + ((g1905) & (!ax36x) & (!ax37x) & (!g1879) & (!g1908)) + ((g1905) & (!ax36x) & (!ax37x) & (!g1879) & (g1908)) + ((g1905) & (!ax36x) & (!ax37x) & (g1879) & (!g1908)) + ((g1905) & (!ax36x) & (ax37x) & (!g1879) & (!g1908)) + ((g1905) & (!ax36x) & (ax37x) & (g1879) & (!g1908)) + ((g1905) & (!ax36x) & (ax37x) & (g1879) & (g1908)) + ((g1905) & (ax36x) & (!ax37x) & (g1879) & (!g1908)) + ((g1905) & (ax36x) & (!ax37x) & (g1879) & (g1908)) + ((g1905) & (ax36x) & (ax37x) & (!g1879) & (!g1908)) + ((g1905) & (ax36x) & (ax37x) & (!g1879) & (g1908)) + ((g1905) & (ax36x) & (ax37x) & (g1879) & (!g1908)) + ((g1905) & (ax36x) & (ax37x) & (g1879) & (g1908)));
	assign g1910 = (((!g1742) & (!g1720) & (g1906) & (g1907) & (g1909)) + ((!g1742) & (g1720) & (g1906) & (!g1907) & (g1909)) + ((!g1742) & (g1720) & (g1906) & (g1907) & (!g1909)) + ((!g1742) & (g1720) & (g1906) & (g1907) & (g1909)) + ((g1742) & (!g1720) & (!g1906) & (g1907) & (g1909)) + ((g1742) & (!g1720) & (g1906) & (!g1907) & (!g1909)) + ((g1742) & (!g1720) & (g1906) & (!g1907) & (g1909)) + ((g1742) & (!g1720) & (g1906) & (g1907) & (!g1909)) + ((g1742) & (!g1720) & (g1906) & (g1907) & (g1909)) + ((g1742) & (g1720) & (!g1906) & (!g1907) & (g1909)) + ((g1742) & (g1720) & (!g1906) & (g1907) & (!g1909)) + ((g1742) & (g1720) & (!g1906) & (g1907) & (g1909)) + ((g1742) & (g1720) & (g1906) & (!g1907) & (!g1909)) + ((g1742) & (g1720) & (g1906) & (!g1907) & (g1909)) + ((g1742) & (g1720) & (g1906) & (g1907) & (!g1909)) + ((g1742) & (g1720) & (g1906) & (g1907) & (g1909)));
	assign g1911 = (((!g1586) & (!g1568) & (g1903) & (g1904) & (g1910)) + ((!g1586) & (g1568) & (g1903) & (!g1904) & (g1910)) + ((!g1586) & (g1568) & (g1903) & (g1904) & (!g1910)) + ((!g1586) & (g1568) & (g1903) & (g1904) & (g1910)) + ((g1586) & (!g1568) & (!g1903) & (g1904) & (g1910)) + ((g1586) & (!g1568) & (g1903) & (!g1904) & (!g1910)) + ((g1586) & (!g1568) & (g1903) & (!g1904) & (g1910)) + ((g1586) & (!g1568) & (g1903) & (g1904) & (!g1910)) + ((g1586) & (!g1568) & (g1903) & (g1904) & (g1910)) + ((g1586) & (g1568) & (!g1903) & (!g1904) & (g1910)) + ((g1586) & (g1568) & (!g1903) & (g1904) & (!g1910)) + ((g1586) & (g1568) & (!g1903) & (g1904) & (g1910)) + ((g1586) & (g1568) & (g1903) & (!g1904) & (!g1910)) + ((g1586) & (g1568) & (g1903) & (!g1904) & (g1910)) + ((g1586) & (g1568) & (g1903) & (g1904) & (!g1910)) + ((g1586) & (g1568) & (g1903) & (g1904) & (g1910)));
	assign g1912 = (((!g1437) & (!g1423) & (g1901) & (g1902) & (g1911)) + ((!g1437) & (g1423) & (g1901) & (!g1902) & (g1911)) + ((!g1437) & (g1423) & (g1901) & (g1902) & (!g1911)) + ((!g1437) & (g1423) & (g1901) & (g1902) & (g1911)) + ((g1437) & (!g1423) & (!g1901) & (g1902) & (g1911)) + ((g1437) & (!g1423) & (g1901) & (!g1902) & (!g1911)) + ((g1437) & (!g1423) & (g1901) & (!g1902) & (g1911)) + ((g1437) & (!g1423) & (g1901) & (g1902) & (!g1911)) + ((g1437) & (!g1423) & (g1901) & (g1902) & (g1911)) + ((g1437) & (g1423) & (!g1901) & (!g1902) & (g1911)) + ((g1437) & (g1423) & (!g1901) & (g1902) & (!g1911)) + ((g1437) & (g1423) & (!g1901) & (g1902) & (g1911)) + ((g1437) & (g1423) & (g1901) & (!g1902) & (!g1911)) + ((g1437) & (g1423) & (g1901) & (!g1902) & (g1911)) + ((g1437) & (g1423) & (g1901) & (g1902) & (!g1911)) + ((g1437) & (g1423) & (g1901) & (g1902) & (g1911)));
	assign g1913 = (((!g1295) & (!g1285) & (g1899) & (g1900) & (g1912)) + ((!g1295) & (g1285) & (g1899) & (!g1900) & (g1912)) + ((!g1295) & (g1285) & (g1899) & (g1900) & (!g1912)) + ((!g1295) & (g1285) & (g1899) & (g1900) & (g1912)) + ((g1295) & (!g1285) & (!g1899) & (g1900) & (g1912)) + ((g1295) & (!g1285) & (g1899) & (!g1900) & (!g1912)) + ((g1295) & (!g1285) & (g1899) & (!g1900) & (g1912)) + ((g1295) & (!g1285) & (g1899) & (g1900) & (!g1912)) + ((g1295) & (!g1285) & (g1899) & (g1900) & (g1912)) + ((g1295) & (g1285) & (!g1899) & (!g1900) & (g1912)) + ((g1295) & (g1285) & (!g1899) & (g1900) & (!g1912)) + ((g1295) & (g1285) & (!g1899) & (g1900) & (g1912)) + ((g1295) & (g1285) & (g1899) & (!g1900) & (!g1912)) + ((g1295) & (g1285) & (g1899) & (!g1900) & (g1912)) + ((g1295) & (g1285) & (g1899) & (g1900) & (!g1912)) + ((g1295) & (g1285) & (g1899) & (g1900) & (g1912)));
	assign g1914 = (((!g1160) & (!g1154) & (g1897) & (g1898) & (g1913)) + ((!g1160) & (g1154) & (g1897) & (!g1898) & (g1913)) + ((!g1160) & (g1154) & (g1897) & (g1898) & (!g1913)) + ((!g1160) & (g1154) & (g1897) & (g1898) & (g1913)) + ((g1160) & (!g1154) & (!g1897) & (g1898) & (g1913)) + ((g1160) & (!g1154) & (g1897) & (!g1898) & (!g1913)) + ((g1160) & (!g1154) & (g1897) & (!g1898) & (g1913)) + ((g1160) & (!g1154) & (g1897) & (g1898) & (!g1913)) + ((g1160) & (!g1154) & (g1897) & (g1898) & (g1913)) + ((g1160) & (g1154) & (!g1897) & (!g1898) & (g1913)) + ((g1160) & (g1154) & (!g1897) & (g1898) & (!g1913)) + ((g1160) & (g1154) & (!g1897) & (g1898) & (g1913)) + ((g1160) & (g1154) & (g1897) & (!g1898) & (!g1913)) + ((g1160) & (g1154) & (g1897) & (!g1898) & (g1913)) + ((g1160) & (g1154) & (g1897) & (g1898) & (!g1913)) + ((g1160) & (g1154) & (g1897) & (g1898) & (g1913)));
	assign g1915 = (((!g1032) & (!g1030) & (g1895) & (g1896) & (g1914)) + ((!g1032) & (g1030) & (g1895) & (!g1896) & (g1914)) + ((!g1032) & (g1030) & (g1895) & (g1896) & (!g1914)) + ((!g1032) & (g1030) & (g1895) & (g1896) & (g1914)) + ((g1032) & (!g1030) & (!g1895) & (g1896) & (g1914)) + ((g1032) & (!g1030) & (g1895) & (!g1896) & (!g1914)) + ((g1032) & (!g1030) & (g1895) & (!g1896) & (g1914)) + ((g1032) & (!g1030) & (g1895) & (g1896) & (!g1914)) + ((g1032) & (!g1030) & (g1895) & (g1896) & (g1914)) + ((g1032) & (g1030) & (!g1895) & (!g1896) & (g1914)) + ((g1032) & (g1030) & (!g1895) & (g1896) & (!g1914)) + ((g1032) & (g1030) & (!g1895) & (g1896) & (g1914)) + ((g1032) & (g1030) & (g1895) & (!g1896) & (!g1914)) + ((g1032) & (g1030) & (g1895) & (!g1896) & (g1914)) + ((g1032) & (g1030) & (g1895) & (g1896) & (!g1914)) + ((g1032) & (g1030) & (g1895) & (g1896) & (g1914)));
	assign g1916 = (((!g851) & (!g914) & (g1893) & (g1894) & (g1915)) + ((!g851) & (g914) & (g1893) & (!g1894) & (g1915)) + ((!g851) & (g914) & (g1893) & (g1894) & (!g1915)) + ((!g851) & (g914) & (g1893) & (g1894) & (g1915)) + ((g851) & (!g914) & (!g1893) & (g1894) & (g1915)) + ((g851) & (!g914) & (g1893) & (!g1894) & (!g1915)) + ((g851) & (!g914) & (g1893) & (!g1894) & (g1915)) + ((g851) & (!g914) & (g1893) & (g1894) & (!g1915)) + ((g851) & (!g914) & (g1893) & (g1894) & (g1915)) + ((g851) & (g914) & (!g1893) & (!g1894) & (g1915)) + ((g851) & (g914) & (!g1893) & (g1894) & (!g1915)) + ((g851) & (g914) & (!g1893) & (g1894) & (g1915)) + ((g851) & (g914) & (g1893) & (!g1894) & (!g1915)) + ((g851) & (g914) & (g1893) & (!g1894) & (g1915)) + ((g851) & (g914) & (g1893) & (g1894) & (!g1915)) + ((g851) & (g914) & (g1893) & (g1894) & (g1915)));
	assign g1917 = (((!g744) & (!g803) & (g1891) & (g1892) & (g1916)) + ((!g744) & (g803) & (g1891) & (!g1892) & (g1916)) + ((!g744) & (g803) & (g1891) & (g1892) & (!g1916)) + ((!g744) & (g803) & (g1891) & (g1892) & (g1916)) + ((g744) & (!g803) & (!g1891) & (g1892) & (g1916)) + ((g744) & (!g803) & (g1891) & (!g1892) & (!g1916)) + ((g744) & (!g803) & (g1891) & (!g1892) & (g1916)) + ((g744) & (!g803) & (g1891) & (g1892) & (!g1916)) + ((g744) & (!g803) & (g1891) & (g1892) & (g1916)) + ((g744) & (g803) & (!g1891) & (!g1892) & (g1916)) + ((g744) & (g803) & (!g1891) & (g1892) & (!g1916)) + ((g744) & (g803) & (!g1891) & (g1892) & (g1916)) + ((g744) & (g803) & (g1891) & (!g1892) & (!g1916)) + ((g744) & (g803) & (g1891) & (!g1892) & (g1916)) + ((g744) & (g803) & (g1891) & (g1892) & (!g1916)) + ((g744) & (g803) & (g1891) & (g1892) & (g1916)));
	assign g1918 = (((!g645) & (!g700) & (g1889) & (g1890) & (g1917)) + ((!g645) & (g700) & (g1889) & (!g1890) & (g1917)) + ((!g645) & (g700) & (g1889) & (g1890) & (!g1917)) + ((!g645) & (g700) & (g1889) & (g1890) & (g1917)) + ((g645) & (!g700) & (!g1889) & (g1890) & (g1917)) + ((g645) & (!g700) & (g1889) & (!g1890) & (!g1917)) + ((g645) & (!g700) & (g1889) & (!g1890) & (g1917)) + ((g645) & (!g700) & (g1889) & (g1890) & (!g1917)) + ((g645) & (!g700) & (g1889) & (g1890) & (g1917)) + ((g645) & (g700) & (!g1889) & (!g1890) & (g1917)) + ((g645) & (g700) & (!g1889) & (g1890) & (!g1917)) + ((g645) & (g700) & (!g1889) & (g1890) & (g1917)) + ((g645) & (g700) & (g1889) & (!g1890) & (!g1917)) + ((g645) & (g700) & (g1889) & (!g1890) & (g1917)) + ((g645) & (g700) & (g1889) & (g1890) & (!g1917)) + ((g645) & (g700) & (g1889) & (g1890) & (g1917)));
	assign g1919 = (((!g553) & (!g604) & (g1887) & (g1888) & (g1918)) + ((!g553) & (g604) & (g1887) & (!g1888) & (g1918)) + ((!g553) & (g604) & (g1887) & (g1888) & (!g1918)) + ((!g553) & (g604) & (g1887) & (g1888) & (g1918)) + ((g553) & (!g604) & (!g1887) & (g1888) & (g1918)) + ((g553) & (!g604) & (g1887) & (!g1888) & (!g1918)) + ((g553) & (!g604) & (g1887) & (!g1888) & (g1918)) + ((g553) & (!g604) & (g1887) & (g1888) & (!g1918)) + ((g553) & (!g604) & (g1887) & (g1888) & (g1918)) + ((g553) & (g604) & (!g1887) & (!g1888) & (g1918)) + ((g553) & (g604) & (!g1887) & (g1888) & (!g1918)) + ((g553) & (g604) & (!g1887) & (g1888) & (g1918)) + ((g553) & (g604) & (g1887) & (!g1888) & (!g1918)) + ((g553) & (g604) & (g1887) & (!g1888) & (g1918)) + ((g553) & (g604) & (g1887) & (g1888) & (!g1918)) + ((g553) & (g604) & (g1887) & (g1888) & (g1918)));
	assign g1920 = (((!g468) & (!g515) & (g1885) & (g1886) & (g1919)) + ((!g468) & (g515) & (g1885) & (!g1886) & (g1919)) + ((!g468) & (g515) & (g1885) & (g1886) & (!g1919)) + ((!g468) & (g515) & (g1885) & (g1886) & (g1919)) + ((g468) & (!g515) & (!g1885) & (g1886) & (g1919)) + ((g468) & (!g515) & (g1885) & (!g1886) & (!g1919)) + ((g468) & (!g515) & (g1885) & (!g1886) & (g1919)) + ((g468) & (!g515) & (g1885) & (g1886) & (!g1919)) + ((g468) & (!g515) & (g1885) & (g1886) & (g1919)) + ((g468) & (g515) & (!g1885) & (!g1886) & (g1919)) + ((g468) & (g515) & (!g1885) & (g1886) & (!g1919)) + ((g468) & (g515) & (!g1885) & (g1886) & (g1919)) + ((g468) & (g515) & (g1885) & (!g1886) & (!g1919)) + ((g468) & (g515) & (g1885) & (!g1886) & (g1919)) + ((g468) & (g515) & (g1885) & (g1886) & (!g1919)) + ((g468) & (g515) & (g1885) & (g1886) & (g1919)));
	assign g1921 = (((!g390) & (!g433) & (g1883) & (g1884) & (g1920)) + ((!g390) & (g433) & (g1883) & (!g1884) & (g1920)) + ((!g390) & (g433) & (g1883) & (g1884) & (!g1920)) + ((!g390) & (g433) & (g1883) & (g1884) & (g1920)) + ((g390) & (!g433) & (!g1883) & (g1884) & (g1920)) + ((g390) & (!g433) & (g1883) & (!g1884) & (!g1920)) + ((g390) & (!g433) & (g1883) & (!g1884) & (g1920)) + ((g390) & (!g433) & (g1883) & (g1884) & (!g1920)) + ((g390) & (!g433) & (g1883) & (g1884) & (g1920)) + ((g390) & (g433) & (!g1883) & (!g1884) & (g1920)) + ((g390) & (g433) & (!g1883) & (g1884) & (!g1920)) + ((g390) & (g433) & (!g1883) & (g1884) & (g1920)) + ((g390) & (g433) & (g1883) & (!g1884) & (!g1920)) + ((g390) & (g433) & (g1883) & (!g1884) & (g1920)) + ((g390) & (g433) & (g1883) & (g1884) & (!g1920)) + ((g390) & (g433) & (g1883) & (g1884) & (g1920)));
	assign g1922 = (((!g319) & (!g358) & (g1881) & (g1882) & (g1921)) + ((!g319) & (g358) & (g1881) & (!g1882) & (g1921)) + ((!g319) & (g358) & (g1881) & (g1882) & (!g1921)) + ((!g319) & (g358) & (g1881) & (g1882) & (g1921)) + ((g319) & (!g358) & (!g1881) & (g1882) & (g1921)) + ((g319) & (!g358) & (g1881) & (!g1882) & (!g1921)) + ((g319) & (!g358) & (g1881) & (!g1882) & (g1921)) + ((g319) & (!g358) & (g1881) & (g1882) & (!g1921)) + ((g319) & (!g358) & (g1881) & (g1882) & (g1921)) + ((g319) & (g358) & (!g1881) & (!g1882) & (g1921)) + ((g319) & (g358) & (!g1881) & (g1882) & (!g1921)) + ((g319) & (g358) & (!g1881) & (g1882) & (g1921)) + ((g319) & (g358) & (g1881) & (!g1882) & (!g1921)) + ((g319) & (g358) & (g1881) & (!g1882) & (g1921)) + ((g319) & (g358) & (g1881) & (g1882) & (!g1921)) + ((g319) & (g358) & (g1881) & (g1882) & (g1921)));
	assign g1923 = (((g1) & (!g1840) & (g1875) & (g1878)) + ((g1) & (g1840) & (!g1875) & (!g1878)) + ((g1) & (g1840) & (!g1875) & (g1878)));
	assign g1924 = (((!g4) & (!g2) & (!g1841) & (!g1872) & (!g1874) & (!g1879)) + ((!g4) & (!g2) & (!g1841) & (!g1872) & (g1874) & (g1879)) + ((!g4) & (!g2) & (!g1841) & (g1872) & (!g1874) & (!g1879)) + ((!g4) & (!g2) & (!g1841) & (g1872) & (g1874) & (g1879)) + ((!g4) & (!g2) & (g1841) & (!g1872) & (!g1874) & (!g1879)) + ((!g4) & (!g2) & (g1841) & (!g1872) & (g1874) & (g1879)) + ((!g4) & (!g2) & (g1841) & (g1872) & (g1874) & (!g1879)) + ((!g4) & (!g2) & (g1841) & (g1872) & (g1874) & (g1879)) + ((!g4) & (g2) & (!g1841) & (!g1872) & (!g1874) & (!g1879)) + ((!g4) & (g2) & (!g1841) & (!g1872) & (g1874) & (g1879)) + ((!g4) & (g2) & (!g1841) & (g1872) & (g1874) & (!g1879)) + ((!g4) & (g2) & (!g1841) & (g1872) & (g1874) & (g1879)) + ((!g4) & (g2) & (g1841) & (!g1872) & (g1874) & (!g1879)) + ((!g4) & (g2) & (g1841) & (!g1872) & (g1874) & (g1879)) + ((!g4) & (g2) & (g1841) & (g1872) & (g1874) & (!g1879)) + ((!g4) & (g2) & (g1841) & (g1872) & (g1874) & (g1879)) + ((g4) & (!g2) & (!g1841) & (!g1872) & (g1874) & (!g1879)) + ((g4) & (!g2) & (!g1841) & (!g1872) & (g1874) & (g1879)) + ((g4) & (!g2) & (!g1841) & (g1872) & (g1874) & (!g1879)) + ((g4) & (!g2) & (!g1841) & (g1872) & (g1874) & (g1879)) + ((g4) & (!g2) & (g1841) & (!g1872) & (g1874) & (!g1879)) + ((g4) & (!g2) & (g1841) & (!g1872) & (g1874) & (g1879)) + ((g4) & (!g2) & (g1841) & (g1872) & (!g1874) & (!g1879)) + ((g4) & (!g2) & (g1841) & (g1872) & (g1874) & (g1879)) + ((g4) & (g2) & (!g1841) & (!g1872) & (g1874) & (!g1879)) + ((g4) & (g2) & (!g1841) & (!g1872) & (g1874) & (g1879)) + ((g4) & (g2) & (!g1841) & (g1872) & (!g1874) & (!g1879)) + ((g4) & (g2) & (!g1841) & (g1872) & (g1874) & (g1879)) + ((g4) & (g2) & (g1841) & (!g1872) & (!g1874) & (!g1879)) + ((g4) & (g2) & (g1841) & (!g1872) & (g1874) & (g1879)) + ((g4) & (g2) & (g1841) & (g1872) & (!g1874) & (!g1879)) + ((g4) & (g2) & (g1841) & (g1872) & (g1874) & (g1879)));
	assign g1925 = (((!g8) & (!g18) & (!g1843) & (g1844) & (g1871) & (!g1879)) + ((!g8) & (!g18) & (g1843) & (!g1844) & (!g1871) & (!g1879)) + ((!g8) & (!g18) & (g1843) & (!g1844) & (!g1871) & (g1879)) + ((!g8) & (!g18) & (g1843) & (!g1844) & (g1871) & (!g1879)) + ((!g8) & (!g18) & (g1843) & (!g1844) & (g1871) & (g1879)) + ((!g8) & (!g18) & (g1843) & (g1844) & (!g1871) & (!g1879)) + ((!g8) & (!g18) & (g1843) & (g1844) & (!g1871) & (g1879)) + ((!g8) & (!g18) & (g1843) & (g1844) & (g1871) & (g1879)) + ((!g8) & (g18) & (!g1843) & (!g1844) & (g1871) & (!g1879)) + ((!g8) & (g18) & (!g1843) & (g1844) & (!g1871) & (!g1879)) + ((!g8) & (g18) & (!g1843) & (g1844) & (g1871) & (!g1879)) + ((!g8) & (g18) & (g1843) & (!g1844) & (!g1871) & (!g1879)) + ((!g8) & (g18) & (g1843) & (!g1844) & (!g1871) & (g1879)) + ((!g8) & (g18) & (g1843) & (!g1844) & (g1871) & (g1879)) + ((!g8) & (g18) & (g1843) & (g1844) & (!g1871) & (g1879)) + ((!g8) & (g18) & (g1843) & (g1844) & (g1871) & (g1879)) + ((g8) & (!g18) & (!g1843) & (!g1844) & (!g1871) & (!g1879)) + ((g8) & (!g18) & (!g1843) & (!g1844) & (g1871) & (!g1879)) + ((g8) & (!g18) & (!g1843) & (g1844) & (!g1871) & (!g1879)) + ((g8) & (!g18) & (g1843) & (!g1844) & (!g1871) & (g1879)) + ((g8) & (!g18) & (g1843) & (!g1844) & (g1871) & (g1879)) + ((g8) & (!g18) & (g1843) & (g1844) & (!g1871) & (g1879)) + ((g8) & (!g18) & (g1843) & (g1844) & (g1871) & (!g1879)) + ((g8) & (!g18) & (g1843) & (g1844) & (g1871) & (g1879)) + ((g8) & (g18) & (!g1843) & (!g1844) & (!g1871) & (!g1879)) + ((g8) & (g18) & (g1843) & (!g1844) & (!g1871) & (g1879)) + ((g8) & (g18) & (g1843) & (!g1844) & (g1871) & (!g1879)) + ((g8) & (g18) & (g1843) & (!g1844) & (g1871) & (g1879)) + ((g8) & (g18) & (g1843) & (g1844) & (!g1871) & (!g1879)) + ((g8) & (g18) & (g1843) & (g1844) & (!g1871) & (g1879)) + ((g8) & (g18) & (g1843) & (g1844) & (g1871) & (!g1879)) + ((g8) & (g18) & (g1843) & (g1844) & (g1871) & (g1879)));
	assign g1926 = (((!g18) & (!g1844) & (g1871) & (!g1879)) + ((!g18) & (g1844) & (!g1871) & (!g1879)) + ((!g18) & (g1844) & (!g1871) & (g1879)) + ((!g18) & (g1844) & (g1871) & (g1879)) + ((g18) & (!g1844) & (!g1871) & (!g1879)) + ((g18) & (g1844) & (!g1871) & (g1879)) + ((g18) & (g1844) & (g1871) & (!g1879)) + ((g18) & (g1844) & (g1871) & (g1879)));
	assign g1927 = (((!g27) & (!g39) & (!g1846) & (g1847) & (g1870) & (!g1879)) + ((!g27) & (!g39) & (g1846) & (!g1847) & (!g1870) & (!g1879)) + ((!g27) & (!g39) & (g1846) & (!g1847) & (!g1870) & (g1879)) + ((!g27) & (!g39) & (g1846) & (!g1847) & (g1870) & (!g1879)) + ((!g27) & (!g39) & (g1846) & (!g1847) & (g1870) & (g1879)) + ((!g27) & (!g39) & (g1846) & (g1847) & (!g1870) & (!g1879)) + ((!g27) & (!g39) & (g1846) & (g1847) & (!g1870) & (g1879)) + ((!g27) & (!g39) & (g1846) & (g1847) & (g1870) & (g1879)) + ((!g27) & (g39) & (!g1846) & (!g1847) & (g1870) & (!g1879)) + ((!g27) & (g39) & (!g1846) & (g1847) & (!g1870) & (!g1879)) + ((!g27) & (g39) & (!g1846) & (g1847) & (g1870) & (!g1879)) + ((!g27) & (g39) & (g1846) & (!g1847) & (!g1870) & (!g1879)) + ((!g27) & (g39) & (g1846) & (!g1847) & (!g1870) & (g1879)) + ((!g27) & (g39) & (g1846) & (!g1847) & (g1870) & (g1879)) + ((!g27) & (g39) & (g1846) & (g1847) & (!g1870) & (g1879)) + ((!g27) & (g39) & (g1846) & (g1847) & (g1870) & (g1879)) + ((g27) & (!g39) & (!g1846) & (!g1847) & (!g1870) & (!g1879)) + ((g27) & (!g39) & (!g1846) & (!g1847) & (g1870) & (!g1879)) + ((g27) & (!g39) & (!g1846) & (g1847) & (!g1870) & (!g1879)) + ((g27) & (!g39) & (g1846) & (!g1847) & (!g1870) & (g1879)) + ((g27) & (!g39) & (g1846) & (!g1847) & (g1870) & (g1879)) + ((g27) & (!g39) & (g1846) & (g1847) & (!g1870) & (g1879)) + ((g27) & (!g39) & (g1846) & (g1847) & (g1870) & (!g1879)) + ((g27) & (!g39) & (g1846) & (g1847) & (g1870) & (g1879)) + ((g27) & (g39) & (!g1846) & (!g1847) & (!g1870) & (!g1879)) + ((g27) & (g39) & (g1846) & (!g1847) & (!g1870) & (g1879)) + ((g27) & (g39) & (g1846) & (!g1847) & (g1870) & (!g1879)) + ((g27) & (g39) & (g1846) & (!g1847) & (g1870) & (g1879)) + ((g27) & (g39) & (g1846) & (g1847) & (!g1870) & (!g1879)) + ((g27) & (g39) & (g1846) & (g1847) & (!g1870) & (g1879)) + ((g27) & (g39) & (g1846) & (g1847) & (g1870) & (!g1879)) + ((g27) & (g39) & (g1846) & (g1847) & (g1870) & (g1879)));
	assign g1928 = (((!g39) & (!g1847) & (g1870) & (!g1879)) + ((!g39) & (g1847) & (!g1870) & (!g1879)) + ((!g39) & (g1847) & (!g1870) & (g1879)) + ((!g39) & (g1847) & (g1870) & (g1879)) + ((g39) & (!g1847) & (!g1870) & (!g1879)) + ((g39) & (g1847) & (!g1870) & (g1879)) + ((g39) & (g1847) & (g1870) & (!g1879)) + ((g39) & (g1847) & (g1870) & (g1879)));
	assign g1929 = (((!g54) & (!g68) & (!g1849) & (g1850) & (g1869) & (!g1879)) + ((!g54) & (!g68) & (g1849) & (!g1850) & (!g1869) & (!g1879)) + ((!g54) & (!g68) & (g1849) & (!g1850) & (!g1869) & (g1879)) + ((!g54) & (!g68) & (g1849) & (!g1850) & (g1869) & (!g1879)) + ((!g54) & (!g68) & (g1849) & (!g1850) & (g1869) & (g1879)) + ((!g54) & (!g68) & (g1849) & (g1850) & (!g1869) & (!g1879)) + ((!g54) & (!g68) & (g1849) & (g1850) & (!g1869) & (g1879)) + ((!g54) & (!g68) & (g1849) & (g1850) & (g1869) & (g1879)) + ((!g54) & (g68) & (!g1849) & (!g1850) & (g1869) & (!g1879)) + ((!g54) & (g68) & (!g1849) & (g1850) & (!g1869) & (!g1879)) + ((!g54) & (g68) & (!g1849) & (g1850) & (g1869) & (!g1879)) + ((!g54) & (g68) & (g1849) & (!g1850) & (!g1869) & (!g1879)) + ((!g54) & (g68) & (g1849) & (!g1850) & (!g1869) & (g1879)) + ((!g54) & (g68) & (g1849) & (!g1850) & (g1869) & (g1879)) + ((!g54) & (g68) & (g1849) & (g1850) & (!g1869) & (g1879)) + ((!g54) & (g68) & (g1849) & (g1850) & (g1869) & (g1879)) + ((g54) & (!g68) & (!g1849) & (!g1850) & (!g1869) & (!g1879)) + ((g54) & (!g68) & (!g1849) & (!g1850) & (g1869) & (!g1879)) + ((g54) & (!g68) & (!g1849) & (g1850) & (!g1869) & (!g1879)) + ((g54) & (!g68) & (g1849) & (!g1850) & (!g1869) & (g1879)) + ((g54) & (!g68) & (g1849) & (!g1850) & (g1869) & (g1879)) + ((g54) & (!g68) & (g1849) & (g1850) & (!g1869) & (g1879)) + ((g54) & (!g68) & (g1849) & (g1850) & (g1869) & (!g1879)) + ((g54) & (!g68) & (g1849) & (g1850) & (g1869) & (g1879)) + ((g54) & (g68) & (!g1849) & (!g1850) & (!g1869) & (!g1879)) + ((g54) & (g68) & (g1849) & (!g1850) & (!g1869) & (g1879)) + ((g54) & (g68) & (g1849) & (!g1850) & (g1869) & (!g1879)) + ((g54) & (g68) & (g1849) & (!g1850) & (g1869) & (g1879)) + ((g54) & (g68) & (g1849) & (g1850) & (!g1869) & (!g1879)) + ((g54) & (g68) & (g1849) & (g1850) & (!g1869) & (g1879)) + ((g54) & (g68) & (g1849) & (g1850) & (g1869) & (!g1879)) + ((g54) & (g68) & (g1849) & (g1850) & (g1869) & (g1879)));
	assign g1930 = (((!g68) & (!g1850) & (g1869) & (!g1879)) + ((!g68) & (g1850) & (!g1869) & (!g1879)) + ((!g68) & (g1850) & (!g1869) & (g1879)) + ((!g68) & (g1850) & (g1869) & (g1879)) + ((g68) & (!g1850) & (!g1869) & (!g1879)) + ((g68) & (g1850) & (!g1869) & (g1879)) + ((g68) & (g1850) & (g1869) & (!g1879)) + ((g68) & (g1850) & (g1869) & (g1879)));
	assign g1931 = (((!g87) & (!g104) & (!g1852) & (g1853) & (g1868) & (!g1879)) + ((!g87) & (!g104) & (g1852) & (!g1853) & (!g1868) & (!g1879)) + ((!g87) & (!g104) & (g1852) & (!g1853) & (!g1868) & (g1879)) + ((!g87) & (!g104) & (g1852) & (!g1853) & (g1868) & (!g1879)) + ((!g87) & (!g104) & (g1852) & (!g1853) & (g1868) & (g1879)) + ((!g87) & (!g104) & (g1852) & (g1853) & (!g1868) & (!g1879)) + ((!g87) & (!g104) & (g1852) & (g1853) & (!g1868) & (g1879)) + ((!g87) & (!g104) & (g1852) & (g1853) & (g1868) & (g1879)) + ((!g87) & (g104) & (!g1852) & (!g1853) & (g1868) & (!g1879)) + ((!g87) & (g104) & (!g1852) & (g1853) & (!g1868) & (!g1879)) + ((!g87) & (g104) & (!g1852) & (g1853) & (g1868) & (!g1879)) + ((!g87) & (g104) & (g1852) & (!g1853) & (!g1868) & (!g1879)) + ((!g87) & (g104) & (g1852) & (!g1853) & (!g1868) & (g1879)) + ((!g87) & (g104) & (g1852) & (!g1853) & (g1868) & (g1879)) + ((!g87) & (g104) & (g1852) & (g1853) & (!g1868) & (g1879)) + ((!g87) & (g104) & (g1852) & (g1853) & (g1868) & (g1879)) + ((g87) & (!g104) & (!g1852) & (!g1853) & (!g1868) & (!g1879)) + ((g87) & (!g104) & (!g1852) & (!g1853) & (g1868) & (!g1879)) + ((g87) & (!g104) & (!g1852) & (g1853) & (!g1868) & (!g1879)) + ((g87) & (!g104) & (g1852) & (!g1853) & (!g1868) & (g1879)) + ((g87) & (!g104) & (g1852) & (!g1853) & (g1868) & (g1879)) + ((g87) & (!g104) & (g1852) & (g1853) & (!g1868) & (g1879)) + ((g87) & (!g104) & (g1852) & (g1853) & (g1868) & (!g1879)) + ((g87) & (!g104) & (g1852) & (g1853) & (g1868) & (g1879)) + ((g87) & (g104) & (!g1852) & (!g1853) & (!g1868) & (!g1879)) + ((g87) & (g104) & (g1852) & (!g1853) & (!g1868) & (g1879)) + ((g87) & (g104) & (g1852) & (!g1853) & (g1868) & (!g1879)) + ((g87) & (g104) & (g1852) & (!g1853) & (g1868) & (g1879)) + ((g87) & (g104) & (g1852) & (g1853) & (!g1868) & (!g1879)) + ((g87) & (g104) & (g1852) & (g1853) & (!g1868) & (g1879)) + ((g87) & (g104) & (g1852) & (g1853) & (g1868) & (!g1879)) + ((g87) & (g104) & (g1852) & (g1853) & (g1868) & (g1879)));
	assign g1932 = (((!g104) & (!g1853) & (g1868) & (!g1879)) + ((!g104) & (g1853) & (!g1868) & (!g1879)) + ((!g104) & (g1853) & (!g1868) & (g1879)) + ((!g104) & (g1853) & (g1868) & (g1879)) + ((g104) & (!g1853) & (!g1868) & (!g1879)) + ((g104) & (g1853) & (!g1868) & (g1879)) + ((g104) & (g1853) & (g1868) & (!g1879)) + ((g104) & (g1853) & (g1868) & (g1879)));
	assign g1933 = (((!g127) & (!g147) & (!g1855) & (g1856) & (g1867) & (!g1879)) + ((!g127) & (!g147) & (g1855) & (!g1856) & (!g1867) & (!g1879)) + ((!g127) & (!g147) & (g1855) & (!g1856) & (!g1867) & (g1879)) + ((!g127) & (!g147) & (g1855) & (!g1856) & (g1867) & (!g1879)) + ((!g127) & (!g147) & (g1855) & (!g1856) & (g1867) & (g1879)) + ((!g127) & (!g147) & (g1855) & (g1856) & (!g1867) & (!g1879)) + ((!g127) & (!g147) & (g1855) & (g1856) & (!g1867) & (g1879)) + ((!g127) & (!g147) & (g1855) & (g1856) & (g1867) & (g1879)) + ((!g127) & (g147) & (!g1855) & (!g1856) & (g1867) & (!g1879)) + ((!g127) & (g147) & (!g1855) & (g1856) & (!g1867) & (!g1879)) + ((!g127) & (g147) & (!g1855) & (g1856) & (g1867) & (!g1879)) + ((!g127) & (g147) & (g1855) & (!g1856) & (!g1867) & (!g1879)) + ((!g127) & (g147) & (g1855) & (!g1856) & (!g1867) & (g1879)) + ((!g127) & (g147) & (g1855) & (!g1856) & (g1867) & (g1879)) + ((!g127) & (g147) & (g1855) & (g1856) & (!g1867) & (g1879)) + ((!g127) & (g147) & (g1855) & (g1856) & (g1867) & (g1879)) + ((g127) & (!g147) & (!g1855) & (!g1856) & (!g1867) & (!g1879)) + ((g127) & (!g147) & (!g1855) & (!g1856) & (g1867) & (!g1879)) + ((g127) & (!g147) & (!g1855) & (g1856) & (!g1867) & (!g1879)) + ((g127) & (!g147) & (g1855) & (!g1856) & (!g1867) & (g1879)) + ((g127) & (!g147) & (g1855) & (!g1856) & (g1867) & (g1879)) + ((g127) & (!g147) & (g1855) & (g1856) & (!g1867) & (g1879)) + ((g127) & (!g147) & (g1855) & (g1856) & (g1867) & (!g1879)) + ((g127) & (!g147) & (g1855) & (g1856) & (g1867) & (g1879)) + ((g127) & (g147) & (!g1855) & (!g1856) & (!g1867) & (!g1879)) + ((g127) & (g147) & (g1855) & (!g1856) & (!g1867) & (g1879)) + ((g127) & (g147) & (g1855) & (!g1856) & (g1867) & (!g1879)) + ((g127) & (g147) & (g1855) & (!g1856) & (g1867) & (g1879)) + ((g127) & (g147) & (g1855) & (g1856) & (!g1867) & (!g1879)) + ((g127) & (g147) & (g1855) & (g1856) & (!g1867) & (g1879)) + ((g127) & (g147) & (g1855) & (g1856) & (g1867) & (!g1879)) + ((g127) & (g147) & (g1855) & (g1856) & (g1867) & (g1879)));
	assign g1934 = (((!g147) & (!g1856) & (g1867) & (!g1879)) + ((!g147) & (g1856) & (!g1867) & (!g1879)) + ((!g147) & (g1856) & (!g1867) & (g1879)) + ((!g147) & (g1856) & (g1867) & (g1879)) + ((g147) & (!g1856) & (!g1867) & (!g1879)) + ((g147) & (g1856) & (!g1867) & (g1879)) + ((g147) & (g1856) & (g1867) & (!g1879)) + ((g147) & (g1856) & (g1867) & (g1879)));
	assign g1935 = (((!g174) & (!g198) & (!g1858) & (g1859) & (g1866) & (!g1879)) + ((!g174) & (!g198) & (g1858) & (!g1859) & (!g1866) & (!g1879)) + ((!g174) & (!g198) & (g1858) & (!g1859) & (!g1866) & (g1879)) + ((!g174) & (!g198) & (g1858) & (!g1859) & (g1866) & (!g1879)) + ((!g174) & (!g198) & (g1858) & (!g1859) & (g1866) & (g1879)) + ((!g174) & (!g198) & (g1858) & (g1859) & (!g1866) & (!g1879)) + ((!g174) & (!g198) & (g1858) & (g1859) & (!g1866) & (g1879)) + ((!g174) & (!g198) & (g1858) & (g1859) & (g1866) & (g1879)) + ((!g174) & (g198) & (!g1858) & (!g1859) & (g1866) & (!g1879)) + ((!g174) & (g198) & (!g1858) & (g1859) & (!g1866) & (!g1879)) + ((!g174) & (g198) & (!g1858) & (g1859) & (g1866) & (!g1879)) + ((!g174) & (g198) & (g1858) & (!g1859) & (!g1866) & (!g1879)) + ((!g174) & (g198) & (g1858) & (!g1859) & (!g1866) & (g1879)) + ((!g174) & (g198) & (g1858) & (!g1859) & (g1866) & (g1879)) + ((!g174) & (g198) & (g1858) & (g1859) & (!g1866) & (g1879)) + ((!g174) & (g198) & (g1858) & (g1859) & (g1866) & (g1879)) + ((g174) & (!g198) & (!g1858) & (!g1859) & (!g1866) & (!g1879)) + ((g174) & (!g198) & (!g1858) & (!g1859) & (g1866) & (!g1879)) + ((g174) & (!g198) & (!g1858) & (g1859) & (!g1866) & (!g1879)) + ((g174) & (!g198) & (g1858) & (!g1859) & (!g1866) & (g1879)) + ((g174) & (!g198) & (g1858) & (!g1859) & (g1866) & (g1879)) + ((g174) & (!g198) & (g1858) & (g1859) & (!g1866) & (g1879)) + ((g174) & (!g198) & (g1858) & (g1859) & (g1866) & (!g1879)) + ((g174) & (!g198) & (g1858) & (g1859) & (g1866) & (g1879)) + ((g174) & (g198) & (!g1858) & (!g1859) & (!g1866) & (!g1879)) + ((g174) & (g198) & (g1858) & (!g1859) & (!g1866) & (g1879)) + ((g174) & (g198) & (g1858) & (!g1859) & (g1866) & (!g1879)) + ((g174) & (g198) & (g1858) & (!g1859) & (g1866) & (g1879)) + ((g174) & (g198) & (g1858) & (g1859) & (!g1866) & (!g1879)) + ((g174) & (g198) & (g1858) & (g1859) & (!g1866) & (g1879)) + ((g174) & (g198) & (g1858) & (g1859) & (g1866) & (!g1879)) + ((g174) & (g198) & (g1858) & (g1859) & (g1866) & (g1879)));
	assign g1936 = (((!g198) & (!g1859) & (g1866) & (!g1879)) + ((!g198) & (g1859) & (!g1866) & (!g1879)) + ((!g198) & (g1859) & (!g1866) & (g1879)) + ((!g198) & (g1859) & (g1866) & (g1879)) + ((g198) & (!g1859) & (!g1866) & (!g1879)) + ((g198) & (g1859) & (!g1866) & (g1879)) + ((g198) & (g1859) & (g1866) & (!g1879)) + ((g198) & (g1859) & (g1866) & (g1879)));
	assign g1937 = (((!g229) & (!g255) & (!g1861) & (g1862) & (g1865) & (!g1879)) + ((!g229) & (!g255) & (g1861) & (!g1862) & (!g1865) & (!g1879)) + ((!g229) & (!g255) & (g1861) & (!g1862) & (!g1865) & (g1879)) + ((!g229) & (!g255) & (g1861) & (!g1862) & (g1865) & (!g1879)) + ((!g229) & (!g255) & (g1861) & (!g1862) & (g1865) & (g1879)) + ((!g229) & (!g255) & (g1861) & (g1862) & (!g1865) & (!g1879)) + ((!g229) & (!g255) & (g1861) & (g1862) & (!g1865) & (g1879)) + ((!g229) & (!g255) & (g1861) & (g1862) & (g1865) & (g1879)) + ((!g229) & (g255) & (!g1861) & (!g1862) & (g1865) & (!g1879)) + ((!g229) & (g255) & (!g1861) & (g1862) & (!g1865) & (!g1879)) + ((!g229) & (g255) & (!g1861) & (g1862) & (g1865) & (!g1879)) + ((!g229) & (g255) & (g1861) & (!g1862) & (!g1865) & (!g1879)) + ((!g229) & (g255) & (g1861) & (!g1862) & (!g1865) & (g1879)) + ((!g229) & (g255) & (g1861) & (!g1862) & (g1865) & (g1879)) + ((!g229) & (g255) & (g1861) & (g1862) & (!g1865) & (g1879)) + ((!g229) & (g255) & (g1861) & (g1862) & (g1865) & (g1879)) + ((g229) & (!g255) & (!g1861) & (!g1862) & (!g1865) & (!g1879)) + ((g229) & (!g255) & (!g1861) & (!g1862) & (g1865) & (!g1879)) + ((g229) & (!g255) & (!g1861) & (g1862) & (!g1865) & (!g1879)) + ((g229) & (!g255) & (g1861) & (!g1862) & (!g1865) & (g1879)) + ((g229) & (!g255) & (g1861) & (!g1862) & (g1865) & (g1879)) + ((g229) & (!g255) & (g1861) & (g1862) & (!g1865) & (g1879)) + ((g229) & (!g255) & (g1861) & (g1862) & (g1865) & (!g1879)) + ((g229) & (!g255) & (g1861) & (g1862) & (g1865) & (g1879)) + ((g229) & (g255) & (!g1861) & (!g1862) & (!g1865) & (!g1879)) + ((g229) & (g255) & (g1861) & (!g1862) & (!g1865) & (g1879)) + ((g229) & (g255) & (g1861) & (!g1862) & (g1865) & (!g1879)) + ((g229) & (g255) & (g1861) & (!g1862) & (g1865) & (g1879)) + ((g229) & (g255) & (g1861) & (g1862) & (!g1865) & (!g1879)) + ((g229) & (g255) & (g1861) & (g1862) & (!g1865) & (g1879)) + ((g229) & (g255) & (g1861) & (g1862) & (g1865) & (!g1879)) + ((g229) & (g255) & (g1861) & (g1862) & (g1865) & (g1879)));
	assign g1938 = (((!g255) & (!g1862) & (g1865) & (!g1879)) + ((!g255) & (g1862) & (!g1865) & (!g1879)) + ((!g255) & (g1862) & (!g1865) & (g1879)) + ((!g255) & (g1862) & (g1865) & (g1879)) + ((g255) & (!g1862) & (!g1865) & (!g1879)) + ((g255) & (g1862) & (!g1865) & (g1879)) + ((g255) & (g1862) & (g1865) & (!g1879)) + ((g255) & (g1862) & (g1865) & (g1879)));
	assign g1939 = (((!g290) & (!g319) & (!g1864) & (g1789) & (g1839) & (!g1879)) + ((!g290) & (!g319) & (g1864) & (!g1789) & (!g1839) & (!g1879)) + ((!g290) & (!g319) & (g1864) & (!g1789) & (!g1839) & (g1879)) + ((!g290) & (!g319) & (g1864) & (!g1789) & (g1839) & (!g1879)) + ((!g290) & (!g319) & (g1864) & (!g1789) & (g1839) & (g1879)) + ((!g290) & (!g319) & (g1864) & (g1789) & (!g1839) & (!g1879)) + ((!g290) & (!g319) & (g1864) & (g1789) & (!g1839) & (g1879)) + ((!g290) & (!g319) & (g1864) & (g1789) & (g1839) & (g1879)) + ((!g290) & (g319) & (!g1864) & (!g1789) & (g1839) & (!g1879)) + ((!g290) & (g319) & (!g1864) & (g1789) & (!g1839) & (!g1879)) + ((!g290) & (g319) & (!g1864) & (g1789) & (g1839) & (!g1879)) + ((!g290) & (g319) & (g1864) & (!g1789) & (!g1839) & (!g1879)) + ((!g290) & (g319) & (g1864) & (!g1789) & (!g1839) & (g1879)) + ((!g290) & (g319) & (g1864) & (!g1789) & (g1839) & (g1879)) + ((!g290) & (g319) & (g1864) & (g1789) & (!g1839) & (g1879)) + ((!g290) & (g319) & (g1864) & (g1789) & (g1839) & (g1879)) + ((g290) & (!g319) & (!g1864) & (!g1789) & (!g1839) & (!g1879)) + ((g290) & (!g319) & (!g1864) & (!g1789) & (g1839) & (!g1879)) + ((g290) & (!g319) & (!g1864) & (g1789) & (!g1839) & (!g1879)) + ((g290) & (!g319) & (g1864) & (!g1789) & (!g1839) & (g1879)) + ((g290) & (!g319) & (g1864) & (!g1789) & (g1839) & (g1879)) + ((g290) & (!g319) & (g1864) & (g1789) & (!g1839) & (g1879)) + ((g290) & (!g319) & (g1864) & (g1789) & (g1839) & (!g1879)) + ((g290) & (!g319) & (g1864) & (g1789) & (g1839) & (g1879)) + ((g290) & (g319) & (!g1864) & (!g1789) & (!g1839) & (!g1879)) + ((g290) & (g319) & (g1864) & (!g1789) & (!g1839) & (g1879)) + ((g290) & (g319) & (g1864) & (!g1789) & (g1839) & (!g1879)) + ((g290) & (g319) & (g1864) & (!g1789) & (g1839) & (g1879)) + ((g290) & (g319) & (g1864) & (g1789) & (!g1839) & (!g1879)) + ((g290) & (g319) & (g1864) & (g1789) & (!g1839) & (g1879)) + ((g290) & (g319) & (g1864) & (g1789) & (g1839) & (!g1879)) + ((g290) & (g319) & (g1864) & (g1789) & (g1839) & (g1879)));
	assign g1940 = (((!g255) & (!g290) & (g1939) & (g1880) & (g1922)) + ((!g255) & (g290) & (g1939) & (!g1880) & (g1922)) + ((!g255) & (g290) & (g1939) & (g1880) & (!g1922)) + ((!g255) & (g290) & (g1939) & (g1880) & (g1922)) + ((g255) & (!g290) & (!g1939) & (g1880) & (g1922)) + ((g255) & (!g290) & (g1939) & (!g1880) & (!g1922)) + ((g255) & (!g290) & (g1939) & (!g1880) & (g1922)) + ((g255) & (!g290) & (g1939) & (g1880) & (!g1922)) + ((g255) & (!g290) & (g1939) & (g1880) & (g1922)) + ((g255) & (g290) & (!g1939) & (!g1880) & (g1922)) + ((g255) & (g290) & (!g1939) & (g1880) & (!g1922)) + ((g255) & (g290) & (!g1939) & (g1880) & (g1922)) + ((g255) & (g290) & (g1939) & (!g1880) & (!g1922)) + ((g255) & (g290) & (g1939) & (!g1880) & (g1922)) + ((g255) & (g290) & (g1939) & (g1880) & (!g1922)) + ((g255) & (g290) & (g1939) & (g1880) & (g1922)));
	assign g1941 = (((!g198) & (!g229) & (g1937) & (g1938) & (g1940)) + ((!g198) & (g229) & (g1937) & (!g1938) & (g1940)) + ((!g198) & (g229) & (g1937) & (g1938) & (!g1940)) + ((!g198) & (g229) & (g1937) & (g1938) & (g1940)) + ((g198) & (!g229) & (!g1937) & (g1938) & (g1940)) + ((g198) & (!g229) & (g1937) & (!g1938) & (!g1940)) + ((g198) & (!g229) & (g1937) & (!g1938) & (g1940)) + ((g198) & (!g229) & (g1937) & (g1938) & (!g1940)) + ((g198) & (!g229) & (g1937) & (g1938) & (g1940)) + ((g198) & (g229) & (!g1937) & (!g1938) & (g1940)) + ((g198) & (g229) & (!g1937) & (g1938) & (!g1940)) + ((g198) & (g229) & (!g1937) & (g1938) & (g1940)) + ((g198) & (g229) & (g1937) & (!g1938) & (!g1940)) + ((g198) & (g229) & (g1937) & (!g1938) & (g1940)) + ((g198) & (g229) & (g1937) & (g1938) & (!g1940)) + ((g198) & (g229) & (g1937) & (g1938) & (g1940)));
	assign g1942 = (((!g147) & (!g174) & (g1935) & (g1936) & (g1941)) + ((!g147) & (g174) & (g1935) & (!g1936) & (g1941)) + ((!g147) & (g174) & (g1935) & (g1936) & (!g1941)) + ((!g147) & (g174) & (g1935) & (g1936) & (g1941)) + ((g147) & (!g174) & (!g1935) & (g1936) & (g1941)) + ((g147) & (!g174) & (g1935) & (!g1936) & (!g1941)) + ((g147) & (!g174) & (g1935) & (!g1936) & (g1941)) + ((g147) & (!g174) & (g1935) & (g1936) & (!g1941)) + ((g147) & (!g174) & (g1935) & (g1936) & (g1941)) + ((g147) & (g174) & (!g1935) & (!g1936) & (g1941)) + ((g147) & (g174) & (!g1935) & (g1936) & (!g1941)) + ((g147) & (g174) & (!g1935) & (g1936) & (g1941)) + ((g147) & (g174) & (g1935) & (!g1936) & (!g1941)) + ((g147) & (g174) & (g1935) & (!g1936) & (g1941)) + ((g147) & (g174) & (g1935) & (g1936) & (!g1941)) + ((g147) & (g174) & (g1935) & (g1936) & (g1941)));
	assign g1943 = (((!g104) & (!g127) & (g1933) & (g1934) & (g1942)) + ((!g104) & (g127) & (g1933) & (!g1934) & (g1942)) + ((!g104) & (g127) & (g1933) & (g1934) & (!g1942)) + ((!g104) & (g127) & (g1933) & (g1934) & (g1942)) + ((g104) & (!g127) & (!g1933) & (g1934) & (g1942)) + ((g104) & (!g127) & (g1933) & (!g1934) & (!g1942)) + ((g104) & (!g127) & (g1933) & (!g1934) & (g1942)) + ((g104) & (!g127) & (g1933) & (g1934) & (!g1942)) + ((g104) & (!g127) & (g1933) & (g1934) & (g1942)) + ((g104) & (g127) & (!g1933) & (!g1934) & (g1942)) + ((g104) & (g127) & (!g1933) & (g1934) & (!g1942)) + ((g104) & (g127) & (!g1933) & (g1934) & (g1942)) + ((g104) & (g127) & (g1933) & (!g1934) & (!g1942)) + ((g104) & (g127) & (g1933) & (!g1934) & (g1942)) + ((g104) & (g127) & (g1933) & (g1934) & (!g1942)) + ((g104) & (g127) & (g1933) & (g1934) & (g1942)));
	assign g1944 = (((!g68) & (!g87) & (g1931) & (g1932) & (g1943)) + ((!g68) & (g87) & (g1931) & (!g1932) & (g1943)) + ((!g68) & (g87) & (g1931) & (g1932) & (!g1943)) + ((!g68) & (g87) & (g1931) & (g1932) & (g1943)) + ((g68) & (!g87) & (!g1931) & (g1932) & (g1943)) + ((g68) & (!g87) & (g1931) & (!g1932) & (!g1943)) + ((g68) & (!g87) & (g1931) & (!g1932) & (g1943)) + ((g68) & (!g87) & (g1931) & (g1932) & (!g1943)) + ((g68) & (!g87) & (g1931) & (g1932) & (g1943)) + ((g68) & (g87) & (!g1931) & (!g1932) & (g1943)) + ((g68) & (g87) & (!g1931) & (g1932) & (!g1943)) + ((g68) & (g87) & (!g1931) & (g1932) & (g1943)) + ((g68) & (g87) & (g1931) & (!g1932) & (!g1943)) + ((g68) & (g87) & (g1931) & (!g1932) & (g1943)) + ((g68) & (g87) & (g1931) & (g1932) & (!g1943)) + ((g68) & (g87) & (g1931) & (g1932) & (g1943)));
	assign g1945 = (((!g39) & (!g54) & (g1929) & (g1930) & (g1944)) + ((!g39) & (g54) & (g1929) & (!g1930) & (g1944)) + ((!g39) & (g54) & (g1929) & (g1930) & (!g1944)) + ((!g39) & (g54) & (g1929) & (g1930) & (g1944)) + ((g39) & (!g54) & (!g1929) & (g1930) & (g1944)) + ((g39) & (!g54) & (g1929) & (!g1930) & (!g1944)) + ((g39) & (!g54) & (g1929) & (!g1930) & (g1944)) + ((g39) & (!g54) & (g1929) & (g1930) & (!g1944)) + ((g39) & (!g54) & (g1929) & (g1930) & (g1944)) + ((g39) & (g54) & (!g1929) & (!g1930) & (g1944)) + ((g39) & (g54) & (!g1929) & (g1930) & (!g1944)) + ((g39) & (g54) & (!g1929) & (g1930) & (g1944)) + ((g39) & (g54) & (g1929) & (!g1930) & (!g1944)) + ((g39) & (g54) & (g1929) & (!g1930) & (g1944)) + ((g39) & (g54) & (g1929) & (g1930) & (!g1944)) + ((g39) & (g54) & (g1929) & (g1930) & (g1944)));
	assign g1946 = (((!g18) & (!g27) & (g1927) & (g1928) & (g1945)) + ((!g18) & (g27) & (g1927) & (!g1928) & (g1945)) + ((!g18) & (g27) & (g1927) & (g1928) & (!g1945)) + ((!g18) & (g27) & (g1927) & (g1928) & (g1945)) + ((g18) & (!g27) & (!g1927) & (g1928) & (g1945)) + ((g18) & (!g27) & (g1927) & (!g1928) & (!g1945)) + ((g18) & (!g27) & (g1927) & (!g1928) & (g1945)) + ((g18) & (!g27) & (g1927) & (g1928) & (!g1945)) + ((g18) & (!g27) & (g1927) & (g1928) & (g1945)) + ((g18) & (g27) & (!g1927) & (!g1928) & (g1945)) + ((g18) & (g27) & (!g1927) & (g1928) & (!g1945)) + ((g18) & (g27) & (!g1927) & (g1928) & (g1945)) + ((g18) & (g27) & (g1927) & (!g1928) & (!g1945)) + ((g18) & (g27) & (g1927) & (!g1928) & (g1945)) + ((g18) & (g27) & (g1927) & (g1928) & (!g1945)) + ((g18) & (g27) & (g1927) & (g1928) & (g1945)));
	assign g1947 = (((!g2) & (!g8) & (g1925) & (g1926) & (g1946)) + ((!g2) & (g8) & (g1925) & (!g1926) & (g1946)) + ((!g2) & (g8) & (g1925) & (g1926) & (!g1946)) + ((!g2) & (g8) & (g1925) & (g1926) & (g1946)) + ((g2) & (!g8) & (!g1925) & (g1926) & (g1946)) + ((g2) & (!g8) & (g1925) & (!g1926) & (!g1946)) + ((g2) & (!g8) & (g1925) & (!g1926) & (g1946)) + ((g2) & (!g8) & (g1925) & (g1926) & (!g1946)) + ((g2) & (!g8) & (g1925) & (g1926) & (g1946)) + ((g2) & (g8) & (!g1925) & (!g1926) & (g1946)) + ((g2) & (g8) & (!g1925) & (g1926) & (!g1946)) + ((g2) & (g8) & (!g1925) & (g1926) & (g1946)) + ((g2) & (g8) & (g1925) & (!g1926) & (!g1946)) + ((g2) & (g8) & (g1925) & (!g1926) & (g1946)) + ((g2) & (g8) & (g1925) & (g1926) & (!g1946)) + ((g2) & (g8) & (g1925) & (g1926) & (g1946)));
	assign g1948 = (((!g2) & (!g1841) & (g1872) & (!g1879)) + ((!g2) & (g1841) & (!g1872) & (!g1879)) + ((!g2) & (g1841) & (!g1872) & (g1879)) + ((!g2) & (g1841) & (g1872) & (g1879)) + ((g2) & (!g1841) & (!g1872) & (!g1879)) + ((g2) & (g1841) & (!g1872) & (g1879)) + ((g2) & (g1841) & (g1872) & (!g1879)) + ((g2) & (g1841) & (g1872) & (g1879)));
	assign g1949 = (((!g1) & (!g1840) & (!g1875) & (!g1877) & (g1878)) + ((!g1) & (!g1840) & (!g1875) & (g1877) & (!g1878)) + ((!g1) & (!g1840) & (!g1875) & (g1877) & (g1878)) + ((!g1) & (g1840) & (g1875) & (!g1877) & (!g1878)) + ((!g1) & (g1840) & (g1875) & (!g1877) & (g1878)) + ((!g1) & (g1840) & (g1875) & (g1877) & (!g1878)) + ((!g1) & (g1840) & (g1875) & (g1877) & (g1878)) + ((g1) & (!g1840) & (!g1875) & (!g1877) & (g1878)) + ((g1) & (!g1840) & (!g1875) & (g1877) & (g1878)) + ((g1) & (g1840) & (g1875) & (!g1877) & (!g1878)) + ((g1) & (g1840) & (g1875) & (!g1877) & (g1878)) + ((g1) & (g1840) & (g1875) & (g1877) & (!g1878)) + ((g1) & (g1840) & (g1875) & (g1877) & (g1878)));
	assign g1950 = (((!g4) & (!g1) & (!g1924) & (!g1947) & (!g1948) & (!g1949)) + ((!g4) & (g1) & (!g1924) & (!g1947) & (!g1948) & (!g1949)) + ((!g4) & (g1) & (!g1924) & (!g1947) & (!g1948) & (g1949)) + ((!g4) & (g1) & (!g1924) & (!g1947) & (g1948) & (!g1949)) + ((!g4) & (g1) & (!g1924) & (!g1947) & (g1948) & (g1949)) + ((!g4) & (g1) & (!g1924) & (g1947) & (!g1948) & (!g1949)) + ((!g4) & (g1) & (!g1924) & (g1947) & (!g1948) & (g1949)) + ((!g4) & (g1) & (!g1924) & (g1947) & (g1948) & (!g1949)) + ((!g4) & (g1) & (!g1924) & (g1947) & (g1948) & (g1949)) + ((!g4) & (g1) & (g1924) & (!g1947) & (!g1948) & (!g1949)) + ((!g4) & (g1) & (g1924) & (!g1947) & (!g1948) & (g1949)) + ((g4) & (!g1) & (!g1924) & (!g1947) & (!g1948) & (!g1949)) + ((g4) & (!g1) & (!g1924) & (!g1947) & (g1948) & (!g1949)) + ((g4) & (!g1) & (!g1924) & (g1947) & (!g1948) & (!g1949)) + ((g4) & (g1) & (!g1924) & (!g1947) & (!g1948) & (!g1949)) + ((g4) & (g1) & (!g1924) & (!g1947) & (!g1948) & (g1949)) + ((g4) & (g1) & (!g1924) & (!g1947) & (g1948) & (!g1949)) + ((g4) & (g1) & (!g1924) & (!g1947) & (g1948) & (g1949)) + ((g4) & (g1) & (!g1924) & (g1947) & (!g1948) & (!g1949)) + ((g4) & (g1) & (!g1924) & (g1947) & (!g1948) & (g1949)) + ((g4) & (g1) & (!g1924) & (g1947) & (g1948) & (!g1949)) + ((g4) & (g1) & (!g1924) & (g1947) & (g1948) & (g1949)) + ((g4) & (g1) & (g1924) & (!g1947) & (!g1948) & (!g1949)) + ((g4) & (g1) & (g1924) & (!g1947) & (!g1948) & (g1949)) + ((g4) & (g1) & (g1924) & (!g1947) & (g1948) & (!g1949)) + ((g4) & (g1) & (g1924) & (!g1947) & (g1948) & (g1949)) + ((g4) & (g1) & (g1924) & (g1947) & (!g1948) & (!g1949)) + ((g4) & (g1) & (g1924) & (g1947) & (!g1948) & (g1949)));
	assign g1951 = (((!g290) & (!g1880) & (g1922) & (!g1923) & (!g1950)) + ((!g290) & (!g1880) & (g1922) & (g1923) & (!g1950)) + ((!g290) & (!g1880) & (g1922) & (g1923) & (g1950)) + ((!g290) & (g1880) & (!g1922) & (!g1923) & (!g1950)) + ((!g290) & (g1880) & (!g1922) & (!g1923) & (g1950)) + ((!g290) & (g1880) & (!g1922) & (g1923) & (!g1950)) + ((!g290) & (g1880) & (!g1922) & (g1923) & (g1950)) + ((!g290) & (g1880) & (g1922) & (!g1923) & (g1950)) + ((g290) & (!g1880) & (!g1922) & (!g1923) & (!g1950)) + ((g290) & (!g1880) & (!g1922) & (g1923) & (!g1950)) + ((g290) & (!g1880) & (!g1922) & (g1923) & (g1950)) + ((g290) & (g1880) & (!g1922) & (!g1923) & (g1950)) + ((g290) & (g1880) & (g1922) & (!g1923) & (!g1950)) + ((g290) & (g1880) & (g1922) & (!g1923) & (g1950)) + ((g290) & (g1880) & (g1922) & (g1923) & (!g1950)) + ((g290) & (g1880) & (g1922) & (g1923) & (g1950)));
	assign g1952 = (((!g319) & (!g358) & (g1882) & (g1921)) + ((!g319) & (g358) & (!g1882) & (g1921)) + ((!g319) & (g358) & (g1882) & (!g1921)) + ((!g319) & (g358) & (g1882) & (g1921)) + ((g319) & (!g358) & (!g1882) & (!g1921)) + ((g319) & (!g358) & (!g1882) & (g1921)) + ((g319) & (!g358) & (g1882) & (!g1921)) + ((g319) & (g358) & (!g1882) & (!g1921)));
	assign g1953 = (((!g1881) & (!g1923) & (!g1950) & (g1952)) + ((!g1881) & (g1923) & (!g1950) & (g1952)) + ((!g1881) & (g1923) & (g1950) & (g1952)) + ((g1881) & (!g1923) & (!g1950) & (!g1952)) + ((g1881) & (!g1923) & (g1950) & (!g1952)) + ((g1881) & (!g1923) & (g1950) & (g1952)) + ((g1881) & (g1923) & (!g1950) & (!g1952)) + ((g1881) & (g1923) & (g1950) & (!g1952)));
	assign g1954 = (((!g358) & (!g1882) & (g1921) & (!g1923) & (!g1950)) + ((!g358) & (!g1882) & (g1921) & (g1923) & (!g1950)) + ((!g358) & (!g1882) & (g1921) & (g1923) & (g1950)) + ((!g358) & (g1882) & (!g1921) & (!g1923) & (!g1950)) + ((!g358) & (g1882) & (!g1921) & (!g1923) & (g1950)) + ((!g358) & (g1882) & (!g1921) & (g1923) & (!g1950)) + ((!g358) & (g1882) & (!g1921) & (g1923) & (g1950)) + ((!g358) & (g1882) & (g1921) & (!g1923) & (g1950)) + ((g358) & (!g1882) & (!g1921) & (!g1923) & (!g1950)) + ((g358) & (!g1882) & (!g1921) & (g1923) & (!g1950)) + ((g358) & (!g1882) & (!g1921) & (g1923) & (g1950)) + ((g358) & (g1882) & (!g1921) & (!g1923) & (g1950)) + ((g358) & (g1882) & (g1921) & (!g1923) & (!g1950)) + ((g358) & (g1882) & (g1921) & (!g1923) & (g1950)) + ((g358) & (g1882) & (g1921) & (g1923) & (!g1950)) + ((g358) & (g1882) & (g1921) & (g1923) & (g1950)));
	assign g1955 = (((!g390) & (!g433) & (g1884) & (g1920)) + ((!g390) & (g433) & (!g1884) & (g1920)) + ((!g390) & (g433) & (g1884) & (!g1920)) + ((!g390) & (g433) & (g1884) & (g1920)) + ((g390) & (!g433) & (!g1884) & (!g1920)) + ((g390) & (!g433) & (!g1884) & (g1920)) + ((g390) & (!g433) & (g1884) & (!g1920)) + ((g390) & (g433) & (!g1884) & (!g1920)));
	assign g1956 = (((!g1883) & (!g1923) & (!g1950) & (g1955)) + ((!g1883) & (g1923) & (!g1950) & (g1955)) + ((!g1883) & (g1923) & (g1950) & (g1955)) + ((g1883) & (!g1923) & (!g1950) & (!g1955)) + ((g1883) & (!g1923) & (g1950) & (!g1955)) + ((g1883) & (!g1923) & (g1950) & (g1955)) + ((g1883) & (g1923) & (!g1950) & (!g1955)) + ((g1883) & (g1923) & (g1950) & (!g1955)));
	assign g1957 = (((!g433) & (!g1884) & (g1920) & (!g1923) & (!g1950)) + ((!g433) & (!g1884) & (g1920) & (g1923) & (!g1950)) + ((!g433) & (!g1884) & (g1920) & (g1923) & (g1950)) + ((!g433) & (g1884) & (!g1920) & (!g1923) & (!g1950)) + ((!g433) & (g1884) & (!g1920) & (!g1923) & (g1950)) + ((!g433) & (g1884) & (!g1920) & (g1923) & (!g1950)) + ((!g433) & (g1884) & (!g1920) & (g1923) & (g1950)) + ((!g433) & (g1884) & (g1920) & (!g1923) & (g1950)) + ((g433) & (!g1884) & (!g1920) & (!g1923) & (!g1950)) + ((g433) & (!g1884) & (!g1920) & (g1923) & (!g1950)) + ((g433) & (!g1884) & (!g1920) & (g1923) & (g1950)) + ((g433) & (g1884) & (!g1920) & (!g1923) & (g1950)) + ((g433) & (g1884) & (g1920) & (!g1923) & (!g1950)) + ((g433) & (g1884) & (g1920) & (!g1923) & (g1950)) + ((g433) & (g1884) & (g1920) & (g1923) & (!g1950)) + ((g433) & (g1884) & (g1920) & (g1923) & (g1950)));
	assign g1958 = (((!g468) & (!g515) & (g1886) & (g1919)) + ((!g468) & (g515) & (!g1886) & (g1919)) + ((!g468) & (g515) & (g1886) & (!g1919)) + ((!g468) & (g515) & (g1886) & (g1919)) + ((g468) & (!g515) & (!g1886) & (!g1919)) + ((g468) & (!g515) & (!g1886) & (g1919)) + ((g468) & (!g515) & (g1886) & (!g1919)) + ((g468) & (g515) & (!g1886) & (!g1919)));
	assign g1959 = (((!g1885) & (!g1923) & (!g1950) & (g1958)) + ((!g1885) & (g1923) & (!g1950) & (g1958)) + ((!g1885) & (g1923) & (g1950) & (g1958)) + ((g1885) & (!g1923) & (!g1950) & (!g1958)) + ((g1885) & (!g1923) & (g1950) & (!g1958)) + ((g1885) & (!g1923) & (g1950) & (g1958)) + ((g1885) & (g1923) & (!g1950) & (!g1958)) + ((g1885) & (g1923) & (g1950) & (!g1958)));
	assign g1960 = (((!g515) & (!g1886) & (g1919) & (!g1923) & (!g1950)) + ((!g515) & (!g1886) & (g1919) & (g1923) & (!g1950)) + ((!g515) & (!g1886) & (g1919) & (g1923) & (g1950)) + ((!g515) & (g1886) & (!g1919) & (!g1923) & (!g1950)) + ((!g515) & (g1886) & (!g1919) & (!g1923) & (g1950)) + ((!g515) & (g1886) & (!g1919) & (g1923) & (!g1950)) + ((!g515) & (g1886) & (!g1919) & (g1923) & (g1950)) + ((!g515) & (g1886) & (g1919) & (!g1923) & (g1950)) + ((g515) & (!g1886) & (!g1919) & (!g1923) & (!g1950)) + ((g515) & (!g1886) & (!g1919) & (g1923) & (!g1950)) + ((g515) & (!g1886) & (!g1919) & (g1923) & (g1950)) + ((g515) & (g1886) & (!g1919) & (!g1923) & (g1950)) + ((g515) & (g1886) & (g1919) & (!g1923) & (!g1950)) + ((g515) & (g1886) & (g1919) & (!g1923) & (g1950)) + ((g515) & (g1886) & (g1919) & (g1923) & (!g1950)) + ((g515) & (g1886) & (g1919) & (g1923) & (g1950)));
	assign g1961 = (((!g553) & (!g604) & (g1888) & (g1918)) + ((!g553) & (g604) & (!g1888) & (g1918)) + ((!g553) & (g604) & (g1888) & (!g1918)) + ((!g553) & (g604) & (g1888) & (g1918)) + ((g553) & (!g604) & (!g1888) & (!g1918)) + ((g553) & (!g604) & (!g1888) & (g1918)) + ((g553) & (!g604) & (g1888) & (!g1918)) + ((g553) & (g604) & (!g1888) & (!g1918)));
	assign g1962 = (((!g1887) & (!g1923) & (!g1950) & (g1961)) + ((!g1887) & (g1923) & (!g1950) & (g1961)) + ((!g1887) & (g1923) & (g1950) & (g1961)) + ((g1887) & (!g1923) & (!g1950) & (!g1961)) + ((g1887) & (!g1923) & (g1950) & (!g1961)) + ((g1887) & (!g1923) & (g1950) & (g1961)) + ((g1887) & (g1923) & (!g1950) & (!g1961)) + ((g1887) & (g1923) & (g1950) & (!g1961)));
	assign g1963 = (((!g604) & (!g1888) & (g1918) & (!g1923) & (!g1950)) + ((!g604) & (!g1888) & (g1918) & (g1923) & (!g1950)) + ((!g604) & (!g1888) & (g1918) & (g1923) & (g1950)) + ((!g604) & (g1888) & (!g1918) & (!g1923) & (!g1950)) + ((!g604) & (g1888) & (!g1918) & (!g1923) & (g1950)) + ((!g604) & (g1888) & (!g1918) & (g1923) & (!g1950)) + ((!g604) & (g1888) & (!g1918) & (g1923) & (g1950)) + ((!g604) & (g1888) & (g1918) & (!g1923) & (g1950)) + ((g604) & (!g1888) & (!g1918) & (!g1923) & (!g1950)) + ((g604) & (!g1888) & (!g1918) & (g1923) & (!g1950)) + ((g604) & (!g1888) & (!g1918) & (g1923) & (g1950)) + ((g604) & (g1888) & (!g1918) & (!g1923) & (g1950)) + ((g604) & (g1888) & (g1918) & (!g1923) & (!g1950)) + ((g604) & (g1888) & (g1918) & (!g1923) & (g1950)) + ((g604) & (g1888) & (g1918) & (g1923) & (!g1950)) + ((g604) & (g1888) & (g1918) & (g1923) & (g1950)));
	assign g1964 = (((!g645) & (!g700) & (g1890) & (g1917)) + ((!g645) & (g700) & (!g1890) & (g1917)) + ((!g645) & (g700) & (g1890) & (!g1917)) + ((!g645) & (g700) & (g1890) & (g1917)) + ((g645) & (!g700) & (!g1890) & (!g1917)) + ((g645) & (!g700) & (!g1890) & (g1917)) + ((g645) & (!g700) & (g1890) & (!g1917)) + ((g645) & (g700) & (!g1890) & (!g1917)));
	assign g1965 = (((!g1889) & (!g1923) & (!g1950) & (g1964)) + ((!g1889) & (g1923) & (!g1950) & (g1964)) + ((!g1889) & (g1923) & (g1950) & (g1964)) + ((g1889) & (!g1923) & (!g1950) & (!g1964)) + ((g1889) & (!g1923) & (g1950) & (!g1964)) + ((g1889) & (!g1923) & (g1950) & (g1964)) + ((g1889) & (g1923) & (!g1950) & (!g1964)) + ((g1889) & (g1923) & (g1950) & (!g1964)));
	assign g1966 = (((!g700) & (!g1890) & (g1917) & (!g1923) & (!g1950)) + ((!g700) & (!g1890) & (g1917) & (g1923) & (!g1950)) + ((!g700) & (!g1890) & (g1917) & (g1923) & (g1950)) + ((!g700) & (g1890) & (!g1917) & (!g1923) & (!g1950)) + ((!g700) & (g1890) & (!g1917) & (!g1923) & (g1950)) + ((!g700) & (g1890) & (!g1917) & (g1923) & (!g1950)) + ((!g700) & (g1890) & (!g1917) & (g1923) & (g1950)) + ((!g700) & (g1890) & (g1917) & (!g1923) & (g1950)) + ((g700) & (!g1890) & (!g1917) & (!g1923) & (!g1950)) + ((g700) & (!g1890) & (!g1917) & (g1923) & (!g1950)) + ((g700) & (!g1890) & (!g1917) & (g1923) & (g1950)) + ((g700) & (g1890) & (!g1917) & (!g1923) & (g1950)) + ((g700) & (g1890) & (g1917) & (!g1923) & (!g1950)) + ((g700) & (g1890) & (g1917) & (!g1923) & (g1950)) + ((g700) & (g1890) & (g1917) & (g1923) & (!g1950)) + ((g700) & (g1890) & (g1917) & (g1923) & (g1950)));
	assign g1967 = (((!g744) & (!g803) & (g1892) & (g1916)) + ((!g744) & (g803) & (!g1892) & (g1916)) + ((!g744) & (g803) & (g1892) & (!g1916)) + ((!g744) & (g803) & (g1892) & (g1916)) + ((g744) & (!g803) & (!g1892) & (!g1916)) + ((g744) & (!g803) & (!g1892) & (g1916)) + ((g744) & (!g803) & (g1892) & (!g1916)) + ((g744) & (g803) & (!g1892) & (!g1916)));
	assign g1968 = (((!g1891) & (!g1923) & (!g1950) & (g1967)) + ((!g1891) & (g1923) & (!g1950) & (g1967)) + ((!g1891) & (g1923) & (g1950) & (g1967)) + ((g1891) & (!g1923) & (!g1950) & (!g1967)) + ((g1891) & (!g1923) & (g1950) & (!g1967)) + ((g1891) & (!g1923) & (g1950) & (g1967)) + ((g1891) & (g1923) & (!g1950) & (!g1967)) + ((g1891) & (g1923) & (g1950) & (!g1967)));
	assign g1969 = (((!g803) & (!g1892) & (g1916) & (!g1923) & (!g1950)) + ((!g803) & (!g1892) & (g1916) & (g1923) & (!g1950)) + ((!g803) & (!g1892) & (g1916) & (g1923) & (g1950)) + ((!g803) & (g1892) & (!g1916) & (!g1923) & (!g1950)) + ((!g803) & (g1892) & (!g1916) & (!g1923) & (g1950)) + ((!g803) & (g1892) & (!g1916) & (g1923) & (!g1950)) + ((!g803) & (g1892) & (!g1916) & (g1923) & (g1950)) + ((!g803) & (g1892) & (g1916) & (!g1923) & (g1950)) + ((g803) & (!g1892) & (!g1916) & (!g1923) & (!g1950)) + ((g803) & (!g1892) & (!g1916) & (g1923) & (!g1950)) + ((g803) & (!g1892) & (!g1916) & (g1923) & (g1950)) + ((g803) & (g1892) & (!g1916) & (!g1923) & (g1950)) + ((g803) & (g1892) & (g1916) & (!g1923) & (!g1950)) + ((g803) & (g1892) & (g1916) & (!g1923) & (g1950)) + ((g803) & (g1892) & (g1916) & (g1923) & (!g1950)) + ((g803) & (g1892) & (g1916) & (g1923) & (g1950)));
	assign g1970 = (((!g851) & (!g914) & (g1894) & (g1915)) + ((!g851) & (g914) & (!g1894) & (g1915)) + ((!g851) & (g914) & (g1894) & (!g1915)) + ((!g851) & (g914) & (g1894) & (g1915)) + ((g851) & (!g914) & (!g1894) & (!g1915)) + ((g851) & (!g914) & (!g1894) & (g1915)) + ((g851) & (!g914) & (g1894) & (!g1915)) + ((g851) & (g914) & (!g1894) & (!g1915)));
	assign g1971 = (((!g1893) & (!g1923) & (!g1950) & (g1970)) + ((!g1893) & (g1923) & (!g1950) & (g1970)) + ((!g1893) & (g1923) & (g1950) & (g1970)) + ((g1893) & (!g1923) & (!g1950) & (!g1970)) + ((g1893) & (!g1923) & (g1950) & (!g1970)) + ((g1893) & (!g1923) & (g1950) & (g1970)) + ((g1893) & (g1923) & (!g1950) & (!g1970)) + ((g1893) & (g1923) & (g1950) & (!g1970)));
	assign g1972 = (((!g914) & (!g1894) & (g1915) & (!g1923) & (!g1950)) + ((!g914) & (!g1894) & (g1915) & (g1923) & (!g1950)) + ((!g914) & (!g1894) & (g1915) & (g1923) & (g1950)) + ((!g914) & (g1894) & (!g1915) & (!g1923) & (!g1950)) + ((!g914) & (g1894) & (!g1915) & (!g1923) & (g1950)) + ((!g914) & (g1894) & (!g1915) & (g1923) & (!g1950)) + ((!g914) & (g1894) & (!g1915) & (g1923) & (g1950)) + ((!g914) & (g1894) & (g1915) & (!g1923) & (g1950)) + ((g914) & (!g1894) & (!g1915) & (!g1923) & (!g1950)) + ((g914) & (!g1894) & (!g1915) & (g1923) & (!g1950)) + ((g914) & (!g1894) & (!g1915) & (g1923) & (g1950)) + ((g914) & (g1894) & (!g1915) & (!g1923) & (g1950)) + ((g914) & (g1894) & (g1915) & (!g1923) & (!g1950)) + ((g914) & (g1894) & (g1915) & (!g1923) & (g1950)) + ((g914) & (g1894) & (g1915) & (g1923) & (!g1950)) + ((g914) & (g1894) & (g1915) & (g1923) & (g1950)));
	assign g1973 = (((!g1032) & (!g1030) & (g1896) & (g1914)) + ((!g1032) & (g1030) & (!g1896) & (g1914)) + ((!g1032) & (g1030) & (g1896) & (!g1914)) + ((!g1032) & (g1030) & (g1896) & (g1914)) + ((g1032) & (!g1030) & (!g1896) & (!g1914)) + ((g1032) & (!g1030) & (!g1896) & (g1914)) + ((g1032) & (!g1030) & (g1896) & (!g1914)) + ((g1032) & (g1030) & (!g1896) & (!g1914)));
	assign g1974 = (((!g1895) & (!g1923) & (!g1950) & (g1973)) + ((!g1895) & (g1923) & (!g1950) & (g1973)) + ((!g1895) & (g1923) & (g1950) & (g1973)) + ((g1895) & (!g1923) & (!g1950) & (!g1973)) + ((g1895) & (!g1923) & (g1950) & (!g1973)) + ((g1895) & (!g1923) & (g1950) & (g1973)) + ((g1895) & (g1923) & (!g1950) & (!g1973)) + ((g1895) & (g1923) & (g1950) & (!g1973)));
	assign g1975 = (((!g1030) & (!g1896) & (g1914) & (!g1923) & (!g1950)) + ((!g1030) & (!g1896) & (g1914) & (g1923) & (!g1950)) + ((!g1030) & (!g1896) & (g1914) & (g1923) & (g1950)) + ((!g1030) & (g1896) & (!g1914) & (!g1923) & (!g1950)) + ((!g1030) & (g1896) & (!g1914) & (!g1923) & (g1950)) + ((!g1030) & (g1896) & (!g1914) & (g1923) & (!g1950)) + ((!g1030) & (g1896) & (!g1914) & (g1923) & (g1950)) + ((!g1030) & (g1896) & (g1914) & (!g1923) & (g1950)) + ((g1030) & (!g1896) & (!g1914) & (!g1923) & (!g1950)) + ((g1030) & (!g1896) & (!g1914) & (g1923) & (!g1950)) + ((g1030) & (!g1896) & (!g1914) & (g1923) & (g1950)) + ((g1030) & (g1896) & (!g1914) & (!g1923) & (g1950)) + ((g1030) & (g1896) & (g1914) & (!g1923) & (!g1950)) + ((g1030) & (g1896) & (g1914) & (!g1923) & (g1950)) + ((g1030) & (g1896) & (g1914) & (g1923) & (!g1950)) + ((g1030) & (g1896) & (g1914) & (g1923) & (g1950)));
	assign g1976 = (((!g1160) & (!g1154) & (g1898) & (g1913)) + ((!g1160) & (g1154) & (!g1898) & (g1913)) + ((!g1160) & (g1154) & (g1898) & (!g1913)) + ((!g1160) & (g1154) & (g1898) & (g1913)) + ((g1160) & (!g1154) & (!g1898) & (!g1913)) + ((g1160) & (!g1154) & (!g1898) & (g1913)) + ((g1160) & (!g1154) & (g1898) & (!g1913)) + ((g1160) & (g1154) & (!g1898) & (!g1913)));
	assign g1977 = (((!g1897) & (!g1923) & (!g1950) & (g1976)) + ((!g1897) & (g1923) & (!g1950) & (g1976)) + ((!g1897) & (g1923) & (g1950) & (g1976)) + ((g1897) & (!g1923) & (!g1950) & (!g1976)) + ((g1897) & (!g1923) & (g1950) & (!g1976)) + ((g1897) & (!g1923) & (g1950) & (g1976)) + ((g1897) & (g1923) & (!g1950) & (!g1976)) + ((g1897) & (g1923) & (g1950) & (!g1976)));
	assign g1978 = (((!g1154) & (!g1898) & (g1913) & (!g1923) & (!g1950)) + ((!g1154) & (!g1898) & (g1913) & (g1923) & (!g1950)) + ((!g1154) & (!g1898) & (g1913) & (g1923) & (g1950)) + ((!g1154) & (g1898) & (!g1913) & (!g1923) & (!g1950)) + ((!g1154) & (g1898) & (!g1913) & (!g1923) & (g1950)) + ((!g1154) & (g1898) & (!g1913) & (g1923) & (!g1950)) + ((!g1154) & (g1898) & (!g1913) & (g1923) & (g1950)) + ((!g1154) & (g1898) & (g1913) & (!g1923) & (g1950)) + ((g1154) & (!g1898) & (!g1913) & (!g1923) & (!g1950)) + ((g1154) & (!g1898) & (!g1913) & (g1923) & (!g1950)) + ((g1154) & (!g1898) & (!g1913) & (g1923) & (g1950)) + ((g1154) & (g1898) & (!g1913) & (!g1923) & (g1950)) + ((g1154) & (g1898) & (g1913) & (!g1923) & (!g1950)) + ((g1154) & (g1898) & (g1913) & (!g1923) & (g1950)) + ((g1154) & (g1898) & (g1913) & (g1923) & (!g1950)) + ((g1154) & (g1898) & (g1913) & (g1923) & (g1950)));
	assign g1979 = (((!g1295) & (!g1285) & (g1900) & (g1912)) + ((!g1295) & (g1285) & (!g1900) & (g1912)) + ((!g1295) & (g1285) & (g1900) & (!g1912)) + ((!g1295) & (g1285) & (g1900) & (g1912)) + ((g1295) & (!g1285) & (!g1900) & (!g1912)) + ((g1295) & (!g1285) & (!g1900) & (g1912)) + ((g1295) & (!g1285) & (g1900) & (!g1912)) + ((g1295) & (g1285) & (!g1900) & (!g1912)));
	assign g1980 = (((!g1899) & (!g1923) & (!g1950) & (g1979)) + ((!g1899) & (g1923) & (!g1950) & (g1979)) + ((!g1899) & (g1923) & (g1950) & (g1979)) + ((g1899) & (!g1923) & (!g1950) & (!g1979)) + ((g1899) & (!g1923) & (g1950) & (!g1979)) + ((g1899) & (!g1923) & (g1950) & (g1979)) + ((g1899) & (g1923) & (!g1950) & (!g1979)) + ((g1899) & (g1923) & (g1950) & (!g1979)));
	assign g1981 = (((!g1285) & (!g1900) & (g1912) & (!g1923) & (!g1950)) + ((!g1285) & (!g1900) & (g1912) & (g1923) & (!g1950)) + ((!g1285) & (!g1900) & (g1912) & (g1923) & (g1950)) + ((!g1285) & (g1900) & (!g1912) & (!g1923) & (!g1950)) + ((!g1285) & (g1900) & (!g1912) & (!g1923) & (g1950)) + ((!g1285) & (g1900) & (!g1912) & (g1923) & (!g1950)) + ((!g1285) & (g1900) & (!g1912) & (g1923) & (g1950)) + ((!g1285) & (g1900) & (g1912) & (!g1923) & (g1950)) + ((g1285) & (!g1900) & (!g1912) & (!g1923) & (!g1950)) + ((g1285) & (!g1900) & (!g1912) & (g1923) & (!g1950)) + ((g1285) & (!g1900) & (!g1912) & (g1923) & (g1950)) + ((g1285) & (g1900) & (!g1912) & (!g1923) & (g1950)) + ((g1285) & (g1900) & (g1912) & (!g1923) & (!g1950)) + ((g1285) & (g1900) & (g1912) & (!g1923) & (g1950)) + ((g1285) & (g1900) & (g1912) & (g1923) & (!g1950)) + ((g1285) & (g1900) & (g1912) & (g1923) & (g1950)));
	assign g1982 = (((!g1437) & (!g1423) & (g1902) & (g1911)) + ((!g1437) & (g1423) & (!g1902) & (g1911)) + ((!g1437) & (g1423) & (g1902) & (!g1911)) + ((!g1437) & (g1423) & (g1902) & (g1911)) + ((g1437) & (!g1423) & (!g1902) & (!g1911)) + ((g1437) & (!g1423) & (!g1902) & (g1911)) + ((g1437) & (!g1423) & (g1902) & (!g1911)) + ((g1437) & (g1423) & (!g1902) & (!g1911)));
	assign g1983 = (((!g1901) & (!g1923) & (!g1950) & (g1982)) + ((!g1901) & (g1923) & (!g1950) & (g1982)) + ((!g1901) & (g1923) & (g1950) & (g1982)) + ((g1901) & (!g1923) & (!g1950) & (!g1982)) + ((g1901) & (!g1923) & (g1950) & (!g1982)) + ((g1901) & (!g1923) & (g1950) & (g1982)) + ((g1901) & (g1923) & (!g1950) & (!g1982)) + ((g1901) & (g1923) & (g1950) & (!g1982)));
	assign g1984 = (((!g1423) & (!g1902) & (g1911) & (!g1923) & (!g1950)) + ((!g1423) & (!g1902) & (g1911) & (g1923) & (!g1950)) + ((!g1423) & (!g1902) & (g1911) & (g1923) & (g1950)) + ((!g1423) & (g1902) & (!g1911) & (!g1923) & (!g1950)) + ((!g1423) & (g1902) & (!g1911) & (!g1923) & (g1950)) + ((!g1423) & (g1902) & (!g1911) & (g1923) & (!g1950)) + ((!g1423) & (g1902) & (!g1911) & (g1923) & (g1950)) + ((!g1423) & (g1902) & (g1911) & (!g1923) & (g1950)) + ((g1423) & (!g1902) & (!g1911) & (!g1923) & (!g1950)) + ((g1423) & (!g1902) & (!g1911) & (g1923) & (!g1950)) + ((g1423) & (!g1902) & (!g1911) & (g1923) & (g1950)) + ((g1423) & (g1902) & (!g1911) & (!g1923) & (g1950)) + ((g1423) & (g1902) & (g1911) & (!g1923) & (!g1950)) + ((g1423) & (g1902) & (g1911) & (!g1923) & (g1950)) + ((g1423) & (g1902) & (g1911) & (g1923) & (!g1950)) + ((g1423) & (g1902) & (g1911) & (g1923) & (g1950)));
	assign g1985 = (((!g1586) & (!g1568) & (g1904) & (g1910)) + ((!g1586) & (g1568) & (!g1904) & (g1910)) + ((!g1586) & (g1568) & (g1904) & (!g1910)) + ((!g1586) & (g1568) & (g1904) & (g1910)) + ((g1586) & (!g1568) & (!g1904) & (!g1910)) + ((g1586) & (!g1568) & (!g1904) & (g1910)) + ((g1586) & (!g1568) & (g1904) & (!g1910)) + ((g1586) & (g1568) & (!g1904) & (!g1910)));
	assign g1986 = (((!g1903) & (!g1923) & (!g1950) & (g1985)) + ((!g1903) & (g1923) & (!g1950) & (g1985)) + ((!g1903) & (g1923) & (g1950) & (g1985)) + ((g1903) & (!g1923) & (!g1950) & (!g1985)) + ((g1903) & (!g1923) & (g1950) & (!g1985)) + ((g1903) & (!g1923) & (g1950) & (g1985)) + ((g1903) & (g1923) & (!g1950) & (!g1985)) + ((g1903) & (g1923) & (g1950) & (!g1985)));
	assign g1987 = (((!g1568) & (!g1904) & (g1910) & (!g1923) & (!g1950)) + ((!g1568) & (!g1904) & (g1910) & (g1923) & (!g1950)) + ((!g1568) & (!g1904) & (g1910) & (g1923) & (g1950)) + ((!g1568) & (g1904) & (!g1910) & (!g1923) & (!g1950)) + ((!g1568) & (g1904) & (!g1910) & (!g1923) & (g1950)) + ((!g1568) & (g1904) & (!g1910) & (g1923) & (!g1950)) + ((!g1568) & (g1904) & (!g1910) & (g1923) & (g1950)) + ((!g1568) & (g1904) & (g1910) & (!g1923) & (g1950)) + ((g1568) & (!g1904) & (!g1910) & (!g1923) & (!g1950)) + ((g1568) & (!g1904) & (!g1910) & (g1923) & (!g1950)) + ((g1568) & (!g1904) & (!g1910) & (g1923) & (g1950)) + ((g1568) & (g1904) & (!g1910) & (!g1923) & (g1950)) + ((g1568) & (g1904) & (g1910) & (!g1923) & (!g1950)) + ((g1568) & (g1904) & (g1910) & (!g1923) & (g1950)) + ((g1568) & (g1904) & (g1910) & (g1923) & (!g1950)) + ((g1568) & (g1904) & (g1910) & (g1923) & (g1950)));
	assign g1988 = (((!g1742) & (!g1720) & (g1907) & (g1909)) + ((!g1742) & (g1720) & (!g1907) & (g1909)) + ((!g1742) & (g1720) & (g1907) & (!g1909)) + ((!g1742) & (g1720) & (g1907) & (g1909)) + ((g1742) & (!g1720) & (!g1907) & (!g1909)) + ((g1742) & (!g1720) & (!g1907) & (g1909)) + ((g1742) & (!g1720) & (g1907) & (!g1909)) + ((g1742) & (g1720) & (!g1907) & (!g1909)));
	assign g1989 = (((!g1906) & (!g1923) & (!g1950) & (g1988)) + ((!g1906) & (g1923) & (!g1950) & (g1988)) + ((!g1906) & (g1923) & (g1950) & (g1988)) + ((g1906) & (!g1923) & (!g1950) & (!g1988)) + ((g1906) & (!g1923) & (g1950) & (!g1988)) + ((g1906) & (!g1923) & (g1950) & (g1988)) + ((g1906) & (g1923) & (!g1950) & (!g1988)) + ((g1906) & (g1923) & (g1950) & (!g1988)));
	assign g1990 = (((!g1720) & (!g1907) & (g1909) & (!g1923) & (!g1950)) + ((!g1720) & (!g1907) & (g1909) & (g1923) & (!g1950)) + ((!g1720) & (!g1907) & (g1909) & (g1923) & (g1950)) + ((!g1720) & (g1907) & (!g1909) & (!g1923) & (!g1950)) + ((!g1720) & (g1907) & (!g1909) & (!g1923) & (g1950)) + ((!g1720) & (g1907) & (!g1909) & (g1923) & (!g1950)) + ((!g1720) & (g1907) & (!g1909) & (g1923) & (g1950)) + ((!g1720) & (g1907) & (g1909) & (!g1923) & (g1950)) + ((g1720) & (!g1907) & (!g1909) & (!g1923) & (!g1950)) + ((g1720) & (!g1907) & (!g1909) & (g1923) & (!g1950)) + ((g1720) & (!g1907) & (!g1909) & (g1923) & (g1950)) + ((g1720) & (g1907) & (!g1909) & (!g1923) & (g1950)) + ((g1720) & (g1907) & (g1909) & (!g1923) & (!g1950)) + ((g1720) & (g1907) & (g1909) & (!g1923) & (g1950)) + ((g1720) & (g1907) & (g1909) & (g1923) & (!g1950)) + ((g1720) & (g1907) & (g1909) & (g1923) & (g1950)));
	assign g1991 = (((!g1905) & (!ax36x) & (!g1879) & (g1908)) + ((!g1905) & (!ax36x) & (g1879) & (g1908)) + ((!g1905) & (ax36x) & (!g1879) & (!g1908)) + ((!g1905) & (ax36x) & (!g1879) & (g1908)) + ((g1905) & (!ax36x) & (!g1879) & (!g1908)) + ((g1905) & (!ax36x) & (g1879) & (!g1908)) + ((g1905) & (ax36x) & (g1879) & (!g1908)) + ((g1905) & (ax36x) & (g1879) & (g1908)));
	assign g1992 = (((!ax36x) & (!ax37x) & (!g1879) & (!g1923) & (!g1950) & (g1991)) + ((!ax36x) & (!ax37x) & (!g1879) & (!g1923) & (g1950) & (!g1991)) + ((!ax36x) & (!ax37x) & (!g1879) & (!g1923) & (g1950) & (g1991)) + ((!ax36x) & (!ax37x) & (!g1879) & (g1923) & (!g1950) & (g1991)) + ((!ax36x) & (!ax37x) & (!g1879) & (g1923) & (g1950) & (g1991)) + ((!ax36x) & (!ax37x) & (g1879) & (!g1923) & (!g1950) & (!g1991)) + ((!ax36x) & (!ax37x) & (g1879) & (g1923) & (!g1950) & (!g1991)) + ((!ax36x) & (!ax37x) & (g1879) & (g1923) & (g1950) & (!g1991)) + ((!ax36x) & (ax37x) & (!g1879) & (!g1923) & (!g1950) & (!g1991)) + ((!ax36x) & (ax37x) & (!g1879) & (g1923) & (!g1950) & (!g1991)) + ((!ax36x) & (ax37x) & (!g1879) & (g1923) & (g1950) & (!g1991)) + ((!ax36x) & (ax37x) & (g1879) & (!g1923) & (!g1950) & (g1991)) + ((!ax36x) & (ax37x) & (g1879) & (!g1923) & (g1950) & (!g1991)) + ((!ax36x) & (ax37x) & (g1879) & (!g1923) & (g1950) & (g1991)) + ((!ax36x) & (ax37x) & (g1879) & (g1923) & (!g1950) & (g1991)) + ((!ax36x) & (ax37x) & (g1879) & (g1923) & (g1950) & (g1991)) + ((ax36x) & (!ax37x) & (!g1879) & (!g1923) & (!g1950) & (!g1991)) + ((ax36x) & (!ax37x) & (!g1879) & (g1923) & (!g1950) & (!g1991)) + ((ax36x) & (!ax37x) & (!g1879) & (g1923) & (g1950) & (!g1991)) + ((ax36x) & (!ax37x) & (g1879) & (!g1923) & (!g1950) & (!g1991)) + ((ax36x) & (!ax37x) & (g1879) & (g1923) & (!g1950) & (!g1991)) + ((ax36x) & (!ax37x) & (g1879) & (g1923) & (g1950) & (!g1991)) + ((ax36x) & (ax37x) & (!g1879) & (!g1923) & (!g1950) & (g1991)) + ((ax36x) & (ax37x) & (!g1879) & (!g1923) & (g1950) & (!g1991)) + ((ax36x) & (ax37x) & (!g1879) & (!g1923) & (g1950) & (g1991)) + ((ax36x) & (ax37x) & (!g1879) & (g1923) & (!g1950) & (g1991)) + ((ax36x) & (ax37x) & (!g1879) & (g1923) & (g1950) & (g1991)) + ((ax36x) & (ax37x) & (g1879) & (!g1923) & (!g1950) & (g1991)) + ((ax36x) & (ax37x) & (g1879) & (!g1923) & (g1950) & (!g1991)) + ((ax36x) & (ax37x) & (g1879) & (!g1923) & (g1950) & (g1991)) + ((ax36x) & (ax37x) & (g1879) & (g1923) & (!g1950) & (g1991)) + ((ax36x) & (ax37x) & (g1879) & (g1923) & (g1950) & (g1991)));
	assign g1993 = (((!ax36x) & (!g1879) & (!g1908) & (!g1923) & (g1950)) + ((!ax36x) & (!g1879) & (g1908) & (!g1923) & (!g1950)) + ((!ax36x) & (!g1879) & (g1908) & (!g1923) & (g1950)) + ((!ax36x) & (!g1879) & (g1908) & (g1923) & (!g1950)) + ((!ax36x) & (!g1879) & (g1908) & (g1923) & (g1950)) + ((!ax36x) & (g1879) & (g1908) & (!g1923) & (!g1950)) + ((!ax36x) & (g1879) & (g1908) & (g1923) & (!g1950)) + ((!ax36x) & (g1879) & (g1908) & (g1923) & (g1950)) + ((ax36x) & (!g1879) & (!g1908) & (!g1923) & (!g1950)) + ((ax36x) & (!g1879) & (!g1908) & (g1923) & (!g1950)) + ((ax36x) & (!g1879) & (!g1908) & (g1923) & (g1950)) + ((ax36x) & (g1879) & (!g1908) & (!g1923) & (!g1950)) + ((ax36x) & (g1879) & (!g1908) & (!g1923) & (g1950)) + ((ax36x) & (g1879) & (!g1908) & (g1923) & (!g1950)) + ((ax36x) & (g1879) & (!g1908) & (g1923) & (g1950)) + ((ax36x) & (g1879) & (g1908) & (!g1923) & (g1950)));
	assign g1994 = (((!ax32x) & (!ax33x)));
	assign g1995 = (((!g1879) & (!ax34x) & (!ax35x) & (!g1923) & (!g1950) & (!g1994)) + ((!g1879) & (!ax34x) & (!ax35x) & (g1923) & (!g1950) & (!g1994)) + ((!g1879) & (!ax34x) & (!ax35x) & (g1923) & (g1950) & (!g1994)) + ((!g1879) & (!ax34x) & (ax35x) & (!g1923) & (g1950) & (!g1994)) + ((!g1879) & (ax34x) & (ax35x) & (!g1923) & (g1950) & (!g1994)) + ((!g1879) & (ax34x) & (ax35x) & (!g1923) & (g1950) & (g1994)) + ((g1879) & (!ax34x) & (!ax35x) & (!g1923) & (!g1950) & (!g1994)) + ((g1879) & (!ax34x) & (!ax35x) & (!g1923) & (!g1950) & (g1994)) + ((g1879) & (!ax34x) & (!ax35x) & (!g1923) & (g1950) & (!g1994)) + ((g1879) & (!ax34x) & (!ax35x) & (g1923) & (!g1950) & (!g1994)) + ((g1879) & (!ax34x) & (!ax35x) & (g1923) & (!g1950) & (g1994)) + ((g1879) & (!ax34x) & (!ax35x) & (g1923) & (g1950) & (!g1994)) + ((g1879) & (!ax34x) & (!ax35x) & (g1923) & (g1950) & (g1994)) + ((g1879) & (!ax34x) & (ax35x) & (!g1923) & (!g1950) & (!g1994)) + ((g1879) & (!ax34x) & (ax35x) & (!g1923) & (g1950) & (!g1994)) + ((g1879) & (!ax34x) & (ax35x) & (!g1923) & (g1950) & (g1994)) + ((g1879) & (!ax34x) & (ax35x) & (g1923) & (!g1950) & (!g1994)) + ((g1879) & (!ax34x) & (ax35x) & (g1923) & (g1950) & (!g1994)) + ((g1879) & (ax34x) & (!ax35x) & (!g1923) & (g1950) & (!g1994)) + ((g1879) & (ax34x) & (!ax35x) & (!g1923) & (g1950) & (g1994)) + ((g1879) & (ax34x) & (ax35x) & (!g1923) & (!g1950) & (!g1994)) + ((g1879) & (ax34x) & (ax35x) & (!g1923) & (!g1950) & (g1994)) + ((g1879) & (ax34x) & (ax35x) & (!g1923) & (g1950) & (!g1994)) + ((g1879) & (ax34x) & (ax35x) & (!g1923) & (g1950) & (g1994)) + ((g1879) & (ax34x) & (ax35x) & (g1923) & (!g1950) & (!g1994)) + ((g1879) & (ax34x) & (ax35x) & (g1923) & (!g1950) & (g1994)) + ((g1879) & (ax34x) & (ax35x) & (g1923) & (g1950) & (!g1994)) + ((g1879) & (ax34x) & (ax35x) & (g1923) & (g1950) & (g1994)));
	assign g1996 = (((!g1720) & (!g1905) & (g1992) & (g1993) & (g1995)) + ((!g1720) & (g1905) & (g1992) & (!g1993) & (g1995)) + ((!g1720) & (g1905) & (g1992) & (g1993) & (!g1995)) + ((!g1720) & (g1905) & (g1992) & (g1993) & (g1995)) + ((g1720) & (!g1905) & (!g1992) & (g1993) & (g1995)) + ((g1720) & (!g1905) & (g1992) & (!g1993) & (!g1995)) + ((g1720) & (!g1905) & (g1992) & (!g1993) & (g1995)) + ((g1720) & (!g1905) & (g1992) & (g1993) & (!g1995)) + ((g1720) & (!g1905) & (g1992) & (g1993) & (g1995)) + ((g1720) & (g1905) & (!g1992) & (!g1993) & (g1995)) + ((g1720) & (g1905) & (!g1992) & (g1993) & (!g1995)) + ((g1720) & (g1905) & (!g1992) & (g1993) & (g1995)) + ((g1720) & (g1905) & (g1992) & (!g1993) & (!g1995)) + ((g1720) & (g1905) & (g1992) & (!g1993) & (g1995)) + ((g1720) & (g1905) & (g1992) & (g1993) & (!g1995)) + ((g1720) & (g1905) & (g1992) & (g1993) & (g1995)));
	assign g1997 = (((!g1568) & (!g1742) & (g1989) & (g1990) & (g1996)) + ((!g1568) & (g1742) & (g1989) & (!g1990) & (g1996)) + ((!g1568) & (g1742) & (g1989) & (g1990) & (!g1996)) + ((!g1568) & (g1742) & (g1989) & (g1990) & (g1996)) + ((g1568) & (!g1742) & (!g1989) & (g1990) & (g1996)) + ((g1568) & (!g1742) & (g1989) & (!g1990) & (!g1996)) + ((g1568) & (!g1742) & (g1989) & (!g1990) & (g1996)) + ((g1568) & (!g1742) & (g1989) & (g1990) & (!g1996)) + ((g1568) & (!g1742) & (g1989) & (g1990) & (g1996)) + ((g1568) & (g1742) & (!g1989) & (!g1990) & (g1996)) + ((g1568) & (g1742) & (!g1989) & (g1990) & (!g1996)) + ((g1568) & (g1742) & (!g1989) & (g1990) & (g1996)) + ((g1568) & (g1742) & (g1989) & (!g1990) & (!g1996)) + ((g1568) & (g1742) & (g1989) & (!g1990) & (g1996)) + ((g1568) & (g1742) & (g1989) & (g1990) & (!g1996)) + ((g1568) & (g1742) & (g1989) & (g1990) & (g1996)));
	assign g1998 = (((!g1423) & (!g1586) & (g1986) & (g1987) & (g1997)) + ((!g1423) & (g1586) & (g1986) & (!g1987) & (g1997)) + ((!g1423) & (g1586) & (g1986) & (g1987) & (!g1997)) + ((!g1423) & (g1586) & (g1986) & (g1987) & (g1997)) + ((g1423) & (!g1586) & (!g1986) & (g1987) & (g1997)) + ((g1423) & (!g1586) & (g1986) & (!g1987) & (!g1997)) + ((g1423) & (!g1586) & (g1986) & (!g1987) & (g1997)) + ((g1423) & (!g1586) & (g1986) & (g1987) & (!g1997)) + ((g1423) & (!g1586) & (g1986) & (g1987) & (g1997)) + ((g1423) & (g1586) & (!g1986) & (!g1987) & (g1997)) + ((g1423) & (g1586) & (!g1986) & (g1987) & (!g1997)) + ((g1423) & (g1586) & (!g1986) & (g1987) & (g1997)) + ((g1423) & (g1586) & (g1986) & (!g1987) & (!g1997)) + ((g1423) & (g1586) & (g1986) & (!g1987) & (g1997)) + ((g1423) & (g1586) & (g1986) & (g1987) & (!g1997)) + ((g1423) & (g1586) & (g1986) & (g1987) & (g1997)));
	assign g1999 = (((!g1285) & (!g1437) & (g1983) & (g1984) & (g1998)) + ((!g1285) & (g1437) & (g1983) & (!g1984) & (g1998)) + ((!g1285) & (g1437) & (g1983) & (g1984) & (!g1998)) + ((!g1285) & (g1437) & (g1983) & (g1984) & (g1998)) + ((g1285) & (!g1437) & (!g1983) & (g1984) & (g1998)) + ((g1285) & (!g1437) & (g1983) & (!g1984) & (!g1998)) + ((g1285) & (!g1437) & (g1983) & (!g1984) & (g1998)) + ((g1285) & (!g1437) & (g1983) & (g1984) & (!g1998)) + ((g1285) & (!g1437) & (g1983) & (g1984) & (g1998)) + ((g1285) & (g1437) & (!g1983) & (!g1984) & (g1998)) + ((g1285) & (g1437) & (!g1983) & (g1984) & (!g1998)) + ((g1285) & (g1437) & (!g1983) & (g1984) & (g1998)) + ((g1285) & (g1437) & (g1983) & (!g1984) & (!g1998)) + ((g1285) & (g1437) & (g1983) & (!g1984) & (g1998)) + ((g1285) & (g1437) & (g1983) & (g1984) & (!g1998)) + ((g1285) & (g1437) & (g1983) & (g1984) & (g1998)));
	assign g2000 = (((!g1154) & (!g1295) & (g1980) & (g1981) & (g1999)) + ((!g1154) & (g1295) & (g1980) & (!g1981) & (g1999)) + ((!g1154) & (g1295) & (g1980) & (g1981) & (!g1999)) + ((!g1154) & (g1295) & (g1980) & (g1981) & (g1999)) + ((g1154) & (!g1295) & (!g1980) & (g1981) & (g1999)) + ((g1154) & (!g1295) & (g1980) & (!g1981) & (!g1999)) + ((g1154) & (!g1295) & (g1980) & (!g1981) & (g1999)) + ((g1154) & (!g1295) & (g1980) & (g1981) & (!g1999)) + ((g1154) & (!g1295) & (g1980) & (g1981) & (g1999)) + ((g1154) & (g1295) & (!g1980) & (!g1981) & (g1999)) + ((g1154) & (g1295) & (!g1980) & (g1981) & (!g1999)) + ((g1154) & (g1295) & (!g1980) & (g1981) & (g1999)) + ((g1154) & (g1295) & (g1980) & (!g1981) & (!g1999)) + ((g1154) & (g1295) & (g1980) & (!g1981) & (g1999)) + ((g1154) & (g1295) & (g1980) & (g1981) & (!g1999)) + ((g1154) & (g1295) & (g1980) & (g1981) & (g1999)));
	assign g2001 = (((!g1030) & (!g1160) & (g1977) & (g1978) & (g2000)) + ((!g1030) & (g1160) & (g1977) & (!g1978) & (g2000)) + ((!g1030) & (g1160) & (g1977) & (g1978) & (!g2000)) + ((!g1030) & (g1160) & (g1977) & (g1978) & (g2000)) + ((g1030) & (!g1160) & (!g1977) & (g1978) & (g2000)) + ((g1030) & (!g1160) & (g1977) & (!g1978) & (!g2000)) + ((g1030) & (!g1160) & (g1977) & (!g1978) & (g2000)) + ((g1030) & (!g1160) & (g1977) & (g1978) & (!g2000)) + ((g1030) & (!g1160) & (g1977) & (g1978) & (g2000)) + ((g1030) & (g1160) & (!g1977) & (!g1978) & (g2000)) + ((g1030) & (g1160) & (!g1977) & (g1978) & (!g2000)) + ((g1030) & (g1160) & (!g1977) & (g1978) & (g2000)) + ((g1030) & (g1160) & (g1977) & (!g1978) & (!g2000)) + ((g1030) & (g1160) & (g1977) & (!g1978) & (g2000)) + ((g1030) & (g1160) & (g1977) & (g1978) & (!g2000)) + ((g1030) & (g1160) & (g1977) & (g1978) & (g2000)));
	assign g2002 = (((!g914) & (!g1032) & (g1974) & (g1975) & (g2001)) + ((!g914) & (g1032) & (g1974) & (!g1975) & (g2001)) + ((!g914) & (g1032) & (g1974) & (g1975) & (!g2001)) + ((!g914) & (g1032) & (g1974) & (g1975) & (g2001)) + ((g914) & (!g1032) & (!g1974) & (g1975) & (g2001)) + ((g914) & (!g1032) & (g1974) & (!g1975) & (!g2001)) + ((g914) & (!g1032) & (g1974) & (!g1975) & (g2001)) + ((g914) & (!g1032) & (g1974) & (g1975) & (!g2001)) + ((g914) & (!g1032) & (g1974) & (g1975) & (g2001)) + ((g914) & (g1032) & (!g1974) & (!g1975) & (g2001)) + ((g914) & (g1032) & (!g1974) & (g1975) & (!g2001)) + ((g914) & (g1032) & (!g1974) & (g1975) & (g2001)) + ((g914) & (g1032) & (g1974) & (!g1975) & (!g2001)) + ((g914) & (g1032) & (g1974) & (!g1975) & (g2001)) + ((g914) & (g1032) & (g1974) & (g1975) & (!g2001)) + ((g914) & (g1032) & (g1974) & (g1975) & (g2001)));
	assign g2003 = (((!g803) & (!g851) & (g1971) & (g1972) & (g2002)) + ((!g803) & (g851) & (g1971) & (!g1972) & (g2002)) + ((!g803) & (g851) & (g1971) & (g1972) & (!g2002)) + ((!g803) & (g851) & (g1971) & (g1972) & (g2002)) + ((g803) & (!g851) & (!g1971) & (g1972) & (g2002)) + ((g803) & (!g851) & (g1971) & (!g1972) & (!g2002)) + ((g803) & (!g851) & (g1971) & (!g1972) & (g2002)) + ((g803) & (!g851) & (g1971) & (g1972) & (!g2002)) + ((g803) & (!g851) & (g1971) & (g1972) & (g2002)) + ((g803) & (g851) & (!g1971) & (!g1972) & (g2002)) + ((g803) & (g851) & (!g1971) & (g1972) & (!g2002)) + ((g803) & (g851) & (!g1971) & (g1972) & (g2002)) + ((g803) & (g851) & (g1971) & (!g1972) & (!g2002)) + ((g803) & (g851) & (g1971) & (!g1972) & (g2002)) + ((g803) & (g851) & (g1971) & (g1972) & (!g2002)) + ((g803) & (g851) & (g1971) & (g1972) & (g2002)));
	assign g2004 = (((!g700) & (!g744) & (g1968) & (g1969) & (g2003)) + ((!g700) & (g744) & (g1968) & (!g1969) & (g2003)) + ((!g700) & (g744) & (g1968) & (g1969) & (!g2003)) + ((!g700) & (g744) & (g1968) & (g1969) & (g2003)) + ((g700) & (!g744) & (!g1968) & (g1969) & (g2003)) + ((g700) & (!g744) & (g1968) & (!g1969) & (!g2003)) + ((g700) & (!g744) & (g1968) & (!g1969) & (g2003)) + ((g700) & (!g744) & (g1968) & (g1969) & (!g2003)) + ((g700) & (!g744) & (g1968) & (g1969) & (g2003)) + ((g700) & (g744) & (!g1968) & (!g1969) & (g2003)) + ((g700) & (g744) & (!g1968) & (g1969) & (!g2003)) + ((g700) & (g744) & (!g1968) & (g1969) & (g2003)) + ((g700) & (g744) & (g1968) & (!g1969) & (!g2003)) + ((g700) & (g744) & (g1968) & (!g1969) & (g2003)) + ((g700) & (g744) & (g1968) & (g1969) & (!g2003)) + ((g700) & (g744) & (g1968) & (g1969) & (g2003)));
	assign g2005 = (((!g604) & (!g645) & (g1965) & (g1966) & (g2004)) + ((!g604) & (g645) & (g1965) & (!g1966) & (g2004)) + ((!g604) & (g645) & (g1965) & (g1966) & (!g2004)) + ((!g604) & (g645) & (g1965) & (g1966) & (g2004)) + ((g604) & (!g645) & (!g1965) & (g1966) & (g2004)) + ((g604) & (!g645) & (g1965) & (!g1966) & (!g2004)) + ((g604) & (!g645) & (g1965) & (!g1966) & (g2004)) + ((g604) & (!g645) & (g1965) & (g1966) & (!g2004)) + ((g604) & (!g645) & (g1965) & (g1966) & (g2004)) + ((g604) & (g645) & (!g1965) & (!g1966) & (g2004)) + ((g604) & (g645) & (!g1965) & (g1966) & (!g2004)) + ((g604) & (g645) & (!g1965) & (g1966) & (g2004)) + ((g604) & (g645) & (g1965) & (!g1966) & (!g2004)) + ((g604) & (g645) & (g1965) & (!g1966) & (g2004)) + ((g604) & (g645) & (g1965) & (g1966) & (!g2004)) + ((g604) & (g645) & (g1965) & (g1966) & (g2004)));
	assign g2006 = (((!g515) & (!g553) & (g1962) & (g1963) & (g2005)) + ((!g515) & (g553) & (g1962) & (!g1963) & (g2005)) + ((!g515) & (g553) & (g1962) & (g1963) & (!g2005)) + ((!g515) & (g553) & (g1962) & (g1963) & (g2005)) + ((g515) & (!g553) & (!g1962) & (g1963) & (g2005)) + ((g515) & (!g553) & (g1962) & (!g1963) & (!g2005)) + ((g515) & (!g553) & (g1962) & (!g1963) & (g2005)) + ((g515) & (!g553) & (g1962) & (g1963) & (!g2005)) + ((g515) & (!g553) & (g1962) & (g1963) & (g2005)) + ((g515) & (g553) & (!g1962) & (!g1963) & (g2005)) + ((g515) & (g553) & (!g1962) & (g1963) & (!g2005)) + ((g515) & (g553) & (!g1962) & (g1963) & (g2005)) + ((g515) & (g553) & (g1962) & (!g1963) & (!g2005)) + ((g515) & (g553) & (g1962) & (!g1963) & (g2005)) + ((g515) & (g553) & (g1962) & (g1963) & (!g2005)) + ((g515) & (g553) & (g1962) & (g1963) & (g2005)));
	assign g2007 = (((!g433) & (!g468) & (g1959) & (g1960) & (g2006)) + ((!g433) & (g468) & (g1959) & (!g1960) & (g2006)) + ((!g433) & (g468) & (g1959) & (g1960) & (!g2006)) + ((!g433) & (g468) & (g1959) & (g1960) & (g2006)) + ((g433) & (!g468) & (!g1959) & (g1960) & (g2006)) + ((g433) & (!g468) & (g1959) & (!g1960) & (!g2006)) + ((g433) & (!g468) & (g1959) & (!g1960) & (g2006)) + ((g433) & (!g468) & (g1959) & (g1960) & (!g2006)) + ((g433) & (!g468) & (g1959) & (g1960) & (g2006)) + ((g433) & (g468) & (!g1959) & (!g1960) & (g2006)) + ((g433) & (g468) & (!g1959) & (g1960) & (!g2006)) + ((g433) & (g468) & (!g1959) & (g1960) & (g2006)) + ((g433) & (g468) & (g1959) & (!g1960) & (!g2006)) + ((g433) & (g468) & (g1959) & (!g1960) & (g2006)) + ((g433) & (g468) & (g1959) & (g1960) & (!g2006)) + ((g433) & (g468) & (g1959) & (g1960) & (g2006)));
	assign g2008 = (((!g358) & (!g390) & (g1956) & (g1957) & (g2007)) + ((!g358) & (g390) & (g1956) & (!g1957) & (g2007)) + ((!g358) & (g390) & (g1956) & (g1957) & (!g2007)) + ((!g358) & (g390) & (g1956) & (g1957) & (g2007)) + ((g358) & (!g390) & (!g1956) & (g1957) & (g2007)) + ((g358) & (!g390) & (g1956) & (!g1957) & (!g2007)) + ((g358) & (!g390) & (g1956) & (!g1957) & (g2007)) + ((g358) & (!g390) & (g1956) & (g1957) & (!g2007)) + ((g358) & (!g390) & (g1956) & (g1957) & (g2007)) + ((g358) & (g390) & (!g1956) & (!g1957) & (g2007)) + ((g358) & (g390) & (!g1956) & (g1957) & (!g2007)) + ((g358) & (g390) & (!g1956) & (g1957) & (g2007)) + ((g358) & (g390) & (g1956) & (!g1957) & (!g2007)) + ((g358) & (g390) & (g1956) & (!g1957) & (g2007)) + ((g358) & (g390) & (g1956) & (g1957) & (!g2007)) + ((g358) & (g390) & (g1956) & (g1957) & (g2007)));
	assign g2009 = (((!g290) & (!g319) & (g1953) & (g1954) & (g2008)) + ((!g290) & (g319) & (g1953) & (!g1954) & (g2008)) + ((!g290) & (g319) & (g1953) & (g1954) & (!g2008)) + ((!g290) & (g319) & (g1953) & (g1954) & (g2008)) + ((g290) & (!g319) & (!g1953) & (g1954) & (g2008)) + ((g290) & (!g319) & (g1953) & (!g1954) & (!g2008)) + ((g290) & (!g319) & (g1953) & (!g1954) & (g2008)) + ((g290) & (!g319) & (g1953) & (g1954) & (!g2008)) + ((g290) & (!g319) & (g1953) & (g1954) & (g2008)) + ((g290) & (g319) & (!g1953) & (!g1954) & (g2008)) + ((g290) & (g319) & (!g1953) & (g1954) & (!g2008)) + ((g290) & (g319) & (!g1953) & (g1954) & (g2008)) + ((g290) & (g319) & (g1953) & (!g1954) & (!g2008)) + ((g290) & (g319) & (g1953) & (!g1954) & (g2008)) + ((g290) & (g319) & (g1953) & (g1954) & (!g2008)) + ((g290) & (g319) & (g1953) & (g1954) & (g2008)));
	assign g2010 = (((!g4) & (!g1947) & (!g1948) & (!g1923) & (!g1950)) + ((!g4) & (!g1947) & (!g1948) & (g1923) & (!g1950)) + ((!g4) & (!g1947) & (!g1948) & (g1923) & (g1950)) + ((!g4) & (!g1947) & (g1948) & (!g1923) & (g1950)) + ((!g4) & (g1947) & (g1948) & (!g1923) & (!g1950)) + ((!g4) & (g1947) & (g1948) & (!g1923) & (g1950)) + ((!g4) & (g1947) & (g1948) & (g1923) & (!g1950)) + ((!g4) & (g1947) & (g1948) & (g1923) & (g1950)) + ((g4) & (!g1947) & (g1948) & (!g1923) & (!g1950)) + ((g4) & (!g1947) & (g1948) & (!g1923) & (g1950)) + ((g4) & (!g1947) & (g1948) & (g1923) & (!g1950)) + ((g4) & (!g1947) & (g1948) & (g1923) & (g1950)) + ((g4) & (g1947) & (!g1948) & (!g1923) & (!g1950)) + ((g4) & (g1947) & (!g1948) & (g1923) & (!g1950)) + ((g4) & (g1947) & (!g1948) & (g1923) & (g1950)) + ((g4) & (g1947) & (g1948) & (!g1923) & (g1950)));
	assign g2011 = (((!g8) & (!g1926) & (g1946) & (!g1923) & (!g1950)) + ((!g8) & (!g1926) & (g1946) & (g1923) & (!g1950)) + ((!g8) & (!g1926) & (g1946) & (g1923) & (g1950)) + ((!g8) & (g1926) & (!g1946) & (!g1923) & (!g1950)) + ((!g8) & (g1926) & (!g1946) & (!g1923) & (g1950)) + ((!g8) & (g1926) & (!g1946) & (g1923) & (!g1950)) + ((!g8) & (g1926) & (!g1946) & (g1923) & (g1950)) + ((!g8) & (g1926) & (g1946) & (!g1923) & (g1950)) + ((g8) & (!g1926) & (!g1946) & (!g1923) & (!g1950)) + ((g8) & (!g1926) & (!g1946) & (g1923) & (!g1950)) + ((g8) & (!g1926) & (!g1946) & (g1923) & (g1950)) + ((g8) & (g1926) & (!g1946) & (!g1923) & (g1950)) + ((g8) & (g1926) & (g1946) & (!g1923) & (!g1950)) + ((g8) & (g1926) & (g1946) & (!g1923) & (g1950)) + ((g8) & (g1926) & (g1946) & (g1923) & (!g1950)) + ((g8) & (g1926) & (g1946) & (g1923) & (g1950)));
	assign g2012 = (((!g18) & (!g27) & (g1928) & (g1945)) + ((!g18) & (g27) & (!g1928) & (g1945)) + ((!g18) & (g27) & (g1928) & (!g1945)) + ((!g18) & (g27) & (g1928) & (g1945)) + ((g18) & (!g27) & (!g1928) & (!g1945)) + ((g18) & (!g27) & (!g1928) & (g1945)) + ((g18) & (!g27) & (g1928) & (!g1945)) + ((g18) & (g27) & (!g1928) & (!g1945)));
	assign g2013 = (((!g1927) & (!g1923) & (!g1950) & (g2012)) + ((!g1927) & (g1923) & (!g1950) & (g2012)) + ((!g1927) & (g1923) & (g1950) & (g2012)) + ((g1927) & (!g1923) & (!g1950) & (!g2012)) + ((g1927) & (!g1923) & (g1950) & (!g2012)) + ((g1927) & (!g1923) & (g1950) & (g2012)) + ((g1927) & (g1923) & (!g1950) & (!g2012)) + ((g1927) & (g1923) & (g1950) & (!g2012)));
	assign g2014 = (((!g27) & (!g1928) & (g1945) & (!g1923) & (!g1950)) + ((!g27) & (!g1928) & (g1945) & (g1923) & (!g1950)) + ((!g27) & (!g1928) & (g1945) & (g1923) & (g1950)) + ((!g27) & (g1928) & (!g1945) & (!g1923) & (!g1950)) + ((!g27) & (g1928) & (!g1945) & (!g1923) & (g1950)) + ((!g27) & (g1928) & (!g1945) & (g1923) & (!g1950)) + ((!g27) & (g1928) & (!g1945) & (g1923) & (g1950)) + ((!g27) & (g1928) & (g1945) & (!g1923) & (g1950)) + ((g27) & (!g1928) & (!g1945) & (!g1923) & (!g1950)) + ((g27) & (!g1928) & (!g1945) & (g1923) & (!g1950)) + ((g27) & (!g1928) & (!g1945) & (g1923) & (g1950)) + ((g27) & (g1928) & (!g1945) & (!g1923) & (g1950)) + ((g27) & (g1928) & (g1945) & (!g1923) & (!g1950)) + ((g27) & (g1928) & (g1945) & (!g1923) & (g1950)) + ((g27) & (g1928) & (g1945) & (g1923) & (!g1950)) + ((g27) & (g1928) & (g1945) & (g1923) & (g1950)));
	assign g2015 = (((!g39) & (!g54) & (g1930) & (g1944)) + ((!g39) & (g54) & (!g1930) & (g1944)) + ((!g39) & (g54) & (g1930) & (!g1944)) + ((!g39) & (g54) & (g1930) & (g1944)) + ((g39) & (!g54) & (!g1930) & (!g1944)) + ((g39) & (!g54) & (!g1930) & (g1944)) + ((g39) & (!g54) & (g1930) & (!g1944)) + ((g39) & (g54) & (!g1930) & (!g1944)));
	assign g2016 = (((!g1929) & (!g1923) & (!g1950) & (g2015)) + ((!g1929) & (g1923) & (!g1950) & (g2015)) + ((!g1929) & (g1923) & (g1950) & (g2015)) + ((g1929) & (!g1923) & (!g1950) & (!g2015)) + ((g1929) & (!g1923) & (g1950) & (!g2015)) + ((g1929) & (!g1923) & (g1950) & (g2015)) + ((g1929) & (g1923) & (!g1950) & (!g2015)) + ((g1929) & (g1923) & (g1950) & (!g2015)));
	assign g2017 = (((!g54) & (!g1930) & (g1944) & (!g1923) & (!g1950)) + ((!g54) & (!g1930) & (g1944) & (g1923) & (!g1950)) + ((!g54) & (!g1930) & (g1944) & (g1923) & (g1950)) + ((!g54) & (g1930) & (!g1944) & (!g1923) & (!g1950)) + ((!g54) & (g1930) & (!g1944) & (!g1923) & (g1950)) + ((!g54) & (g1930) & (!g1944) & (g1923) & (!g1950)) + ((!g54) & (g1930) & (!g1944) & (g1923) & (g1950)) + ((!g54) & (g1930) & (g1944) & (!g1923) & (g1950)) + ((g54) & (!g1930) & (!g1944) & (!g1923) & (!g1950)) + ((g54) & (!g1930) & (!g1944) & (g1923) & (!g1950)) + ((g54) & (!g1930) & (!g1944) & (g1923) & (g1950)) + ((g54) & (g1930) & (!g1944) & (!g1923) & (g1950)) + ((g54) & (g1930) & (g1944) & (!g1923) & (!g1950)) + ((g54) & (g1930) & (g1944) & (!g1923) & (g1950)) + ((g54) & (g1930) & (g1944) & (g1923) & (!g1950)) + ((g54) & (g1930) & (g1944) & (g1923) & (g1950)));
	assign g2018 = (((!g68) & (!g87) & (g1932) & (g1943)) + ((!g68) & (g87) & (!g1932) & (g1943)) + ((!g68) & (g87) & (g1932) & (!g1943)) + ((!g68) & (g87) & (g1932) & (g1943)) + ((g68) & (!g87) & (!g1932) & (!g1943)) + ((g68) & (!g87) & (!g1932) & (g1943)) + ((g68) & (!g87) & (g1932) & (!g1943)) + ((g68) & (g87) & (!g1932) & (!g1943)));
	assign g2019 = (((!g1931) & (!g1923) & (!g1950) & (g2018)) + ((!g1931) & (g1923) & (!g1950) & (g2018)) + ((!g1931) & (g1923) & (g1950) & (g2018)) + ((g1931) & (!g1923) & (!g1950) & (!g2018)) + ((g1931) & (!g1923) & (g1950) & (!g2018)) + ((g1931) & (!g1923) & (g1950) & (g2018)) + ((g1931) & (g1923) & (!g1950) & (!g2018)) + ((g1931) & (g1923) & (g1950) & (!g2018)));
	assign g2020 = (((!g87) & (!g1932) & (g1943) & (!g1923) & (!g1950)) + ((!g87) & (!g1932) & (g1943) & (g1923) & (!g1950)) + ((!g87) & (!g1932) & (g1943) & (g1923) & (g1950)) + ((!g87) & (g1932) & (!g1943) & (!g1923) & (!g1950)) + ((!g87) & (g1932) & (!g1943) & (!g1923) & (g1950)) + ((!g87) & (g1932) & (!g1943) & (g1923) & (!g1950)) + ((!g87) & (g1932) & (!g1943) & (g1923) & (g1950)) + ((!g87) & (g1932) & (g1943) & (!g1923) & (g1950)) + ((g87) & (!g1932) & (!g1943) & (!g1923) & (!g1950)) + ((g87) & (!g1932) & (!g1943) & (g1923) & (!g1950)) + ((g87) & (!g1932) & (!g1943) & (g1923) & (g1950)) + ((g87) & (g1932) & (!g1943) & (!g1923) & (g1950)) + ((g87) & (g1932) & (g1943) & (!g1923) & (!g1950)) + ((g87) & (g1932) & (g1943) & (!g1923) & (g1950)) + ((g87) & (g1932) & (g1943) & (g1923) & (!g1950)) + ((g87) & (g1932) & (g1943) & (g1923) & (g1950)));
	assign g2021 = (((!g104) & (!g127) & (g1934) & (g1942)) + ((!g104) & (g127) & (!g1934) & (g1942)) + ((!g104) & (g127) & (g1934) & (!g1942)) + ((!g104) & (g127) & (g1934) & (g1942)) + ((g104) & (!g127) & (!g1934) & (!g1942)) + ((g104) & (!g127) & (!g1934) & (g1942)) + ((g104) & (!g127) & (g1934) & (!g1942)) + ((g104) & (g127) & (!g1934) & (!g1942)));
	assign g2022 = (((!g1933) & (!g1923) & (!g1950) & (g2021)) + ((!g1933) & (g1923) & (!g1950) & (g2021)) + ((!g1933) & (g1923) & (g1950) & (g2021)) + ((g1933) & (!g1923) & (!g1950) & (!g2021)) + ((g1933) & (!g1923) & (g1950) & (!g2021)) + ((g1933) & (!g1923) & (g1950) & (g2021)) + ((g1933) & (g1923) & (!g1950) & (!g2021)) + ((g1933) & (g1923) & (g1950) & (!g2021)));
	assign g2023 = (((!g127) & (!g1934) & (g1942) & (!g1923) & (!g1950)) + ((!g127) & (!g1934) & (g1942) & (g1923) & (!g1950)) + ((!g127) & (!g1934) & (g1942) & (g1923) & (g1950)) + ((!g127) & (g1934) & (!g1942) & (!g1923) & (!g1950)) + ((!g127) & (g1934) & (!g1942) & (!g1923) & (g1950)) + ((!g127) & (g1934) & (!g1942) & (g1923) & (!g1950)) + ((!g127) & (g1934) & (!g1942) & (g1923) & (g1950)) + ((!g127) & (g1934) & (g1942) & (!g1923) & (g1950)) + ((g127) & (!g1934) & (!g1942) & (!g1923) & (!g1950)) + ((g127) & (!g1934) & (!g1942) & (g1923) & (!g1950)) + ((g127) & (!g1934) & (!g1942) & (g1923) & (g1950)) + ((g127) & (g1934) & (!g1942) & (!g1923) & (g1950)) + ((g127) & (g1934) & (g1942) & (!g1923) & (!g1950)) + ((g127) & (g1934) & (g1942) & (!g1923) & (g1950)) + ((g127) & (g1934) & (g1942) & (g1923) & (!g1950)) + ((g127) & (g1934) & (g1942) & (g1923) & (g1950)));
	assign g2024 = (((!g147) & (!g174) & (g1936) & (g1941)) + ((!g147) & (g174) & (!g1936) & (g1941)) + ((!g147) & (g174) & (g1936) & (!g1941)) + ((!g147) & (g174) & (g1936) & (g1941)) + ((g147) & (!g174) & (!g1936) & (!g1941)) + ((g147) & (!g174) & (!g1936) & (g1941)) + ((g147) & (!g174) & (g1936) & (!g1941)) + ((g147) & (g174) & (!g1936) & (!g1941)));
	assign g2025 = (((!g1935) & (!g1923) & (!g1950) & (g2024)) + ((!g1935) & (g1923) & (!g1950) & (g2024)) + ((!g1935) & (g1923) & (g1950) & (g2024)) + ((g1935) & (!g1923) & (!g1950) & (!g2024)) + ((g1935) & (!g1923) & (g1950) & (!g2024)) + ((g1935) & (!g1923) & (g1950) & (g2024)) + ((g1935) & (g1923) & (!g1950) & (!g2024)) + ((g1935) & (g1923) & (g1950) & (!g2024)));
	assign g2026 = (((!g174) & (!g1936) & (g1941) & (!g1923) & (!g1950)) + ((!g174) & (!g1936) & (g1941) & (g1923) & (!g1950)) + ((!g174) & (!g1936) & (g1941) & (g1923) & (g1950)) + ((!g174) & (g1936) & (!g1941) & (!g1923) & (!g1950)) + ((!g174) & (g1936) & (!g1941) & (!g1923) & (g1950)) + ((!g174) & (g1936) & (!g1941) & (g1923) & (!g1950)) + ((!g174) & (g1936) & (!g1941) & (g1923) & (g1950)) + ((!g174) & (g1936) & (g1941) & (!g1923) & (g1950)) + ((g174) & (!g1936) & (!g1941) & (!g1923) & (!g1950)) + ((g174) & (!g1936) & (!g1941) & (g1923) & (!g1950)) + ((g174) & (!g1936) & (!g1941) & (g1923) & (g1950)) + ((g174) & (g1936) & (!g1941) & (!g1923) & (g1950)) + ((g174) & (g1936) & (g1941) & (!g1923) & (!g1950)) + ((g174) & (g1936) & (g1941) & (!g1923) & (g1950)) + ((g174) & (g1936) & (g1941) & (g1923) & (!g1950)) + ((g174) & (g1936) & (g1941) & (g1923) & (g1950)));
	assign g2027 = (((!g198) & (!g229) & (g1938) & (g1940)) + ((!g198) & (g229) & (!g1938) & (g1940)) + ((!g198) & (g229) & (g1938) & (!g1940)) + ((!g198) & (g229) & (g1938) & (g1940)) + ((g198) & (!g229) & (!g1938) & (!g1940)) + ((g198) & (!g229) & (!g1938) & (g1940)) + ((g198) & (!g229) & (g1938) & (!g1940)) + ((g198) & (g229) & (!g1938) & (!g1940)));
	assign g2028 = (((!g1937) & (!g1923) & (!g1950) & (g2027)) + ((!g1937) & (g1923) & (!g1950) & (g2027)) + ((!g1937) & (g1923) & (g1950) & (g2027)) + ((g1937) & (!g1923) & (!g1950) & (!g2027)) + ((g1937) & (!g1923) & (g1950) & (!g2027)) + ((g1937) & (!g1923) & (g1950) & (g2027)) + ((g1937) & (g1923) & (!g1950) & (!g2027)) + ((g1937) & (g1923) & (g1950) & (!g2027)));
	assign g2029 = (((!g229) & (!g1938) & (g1940) & (!g1923) & (!g1950)) + ((!g229) & (!g1938) & (g1940) & (g1923) & (!g1950)) + ((!g229) & (!g1938) & (g1940) & (g1923) & (g1950)) + ((!g229) & (g1938) & (!g1940) & (!g1923) & (!g1950)) + ((!g229) & (g1938) & (!g1940) & (!g1923) & (g1950)) + ((!g229) & (g1938) & (!g1940) & (g1923) & (!g1950)) + ((!g229) & (g1938) & (!g1940) & (g1923) & (g1950)) + ((!g229) & (g1938) & (g1940) & (!g1923) & (g1950)) + ((g229) & (!g1938) & (!g1940) & (!g1923) & (!g1950)) + ((g229) & (!g1938) & (!g1940) & (g1923) & (!g1950)) + ((g229) & (!g1938) & (!g1940) & (g1923) & (g1950)) + ((g229) & (g1938) & (!g1940) & (!g1923) & (g1950)) + ((g229) & (g1938) & (g1940) & (!g1923) & (!g1950)) + ((g229) & (g1938) & (g1940) & (!g1923) & (g1950)) + ((g229) & (g1938) & (g1940) & (g1923) & (!g1950)) + ((g229) & (g1938) & (g1940) & (g1923) & (g1950)));
	assign g2030 = (((!g255) & (!g290) & (g1880) & (g1922)) + ((!g255) & (g290) & (!g1880) & (g1922)) + ((!g255) & (g290) & (g1880) & (!g1922)) + ((!g255) & (g290) & (g1880) & (g1922)) + ((g255) & (!g290) & (!g1880) & (!g1922)) + ((g255) & (!g290) & (!g1880) & (g1922)) + ((g255) & (!g290) & (g1880) & (!g1922)) + ((g255) & (g290) & (!g1880) & (!g1922)));
	assign g2031 = (((!g1939) & (!g1923) & (!g1950) & (g2030)) + ((!g1939) & (g1923) & (!g1950) & (g2030)) + ((!g1939) & (g1923) & (g1950) & (g2030)) + ((g1939) & (!g1923) & (!g1950) & (!g2030)) + ((g1939) & (!g1923) & (g1950) & (!g2030)) + ((g1939) & (!g1923) & (g1950) & (g2030)) + ((g1939) & (g1923) & (!g1950) & (!g2030)) + ((g1939) & (g1923) & (g1950) & (!g2030)));
	assign g2032 = (((!g229) & (!g255) & (g2031) & (g1951) & (g2009)) + ((!g229) & (g255) & (g2031) & (!g1951) & (g2009)) + ((!g229) & (g255) & (g2031) & (g1951) & (!g2009)) + ((!g229) & (g255) & (g2031) & (g1951) & (g2009)) + ((g229) & (!g255) & (!g2031) & (g1951) & (g2009)) + ((g229) & (!g255) & (g2031) & (!g1951) & (!g2009)) + ((g229) & (!g255) & (g2031) & (!g1951) & (g2009)) + ((g229) & (!g255) & (g2031) & (g1951) & (!g2009)) + ((g229) & (!g255) & (g2031) & (g1951) & (g2009)) + ((g229) & (g255) & (!g2031) & (!g1951) & (g2009)) + ((g229) & (g255) & (!g2031) & (g1951) & (!g2009)) + ((g229) & (g255) & (!g2031) & (g1951) & (g2009)) + ((g229) & (g255) & (g2031) & (!g1951) & (!g2009)) + ((g229) & (g255) & (g2031) & (!g1951) & (g2009)) + ((g229) & (g255) & (g2031) & (g1951) & (!g2009)) + ((g229) & (g255) & (g2031) & (g1951) & (g2009)));
	assign g2033 = (((!g174) & (!g198) & (g2028) & (g2029) & (g2032)) + ((!g174) & (g198) & (g2028) & (!g2029) & (g2032)) + ((!g174) & (g198) & (g2028) & (g2029) & (!g2032)) + ((!g174) & (g198) & (g2028) & (g2029) & (g2032)) + ((g174) & (!g198) & (!g2028) & (g2029) & (g2032)) + ((g174) & (!g198) & (g2028) & (!g2029) & (!g2032)) + ((g174) & (!g198) & (g2028) & (!g2029) & (g2032)) + ((g174) & (!g198) & (g2028) & (g2029) & (!g2032)) + ((g174) & (!g198) & (g2028) & (g2029) & (g2032)) + ((g174) & (g198) & (!g2028) & (!g2029) & (g2032)) + ((g174) & (g198) & (!g2028) & (g2029) & (!g2032)) + ((g174) & (g198) & (!g2028) & (g2029) & (g2032)) + ((g174) & (g198) & (g2028) & (!g2029) & (!g2032)) + ((g174) & (g198) & (g2028) & (!g2029) & (g2032)) + ((g174) & (g198) & (g2028) & (g2029) & (!g2032)) + ((g174) & (g198) & (g2028) & (g2029) & (g2032)));
	assign g2034 = (((!g127) & (!g147) & (g2025) & (g2026) & (g2033)) + ((!g127) & (g147) & (g2025) & (!g2026) & (g2033)) + ((!g127) & (g147) & (g2025) & (g2026) & (!g2033)) + ((!g127) & (g147) & (g2025) & (g2026) & (g2033)) + ((g127) & (!g147) & (!g2025) & (g2026) & (g2033)) + ((g127) & (!g147) & (g2025) & (!g2026) & (!g2033)) + ((g127) & (!g147) & (g2025) & (!g2026) & (g2033)) + ((g127) & (!g147) & (g2025) & (g2026) & (!g2033)) + ((g127) & (!g147) & (g2025) & (g2026) & (g2033)) + ((g127) & (g147) & (!g2025) & (!g2026) & (g2033)) + ((g127) & (g147) & (!g2025) & (g2026) & (!g2033)) + ((g127) & (g147) & (!g2025) & (g2026) & (g2033)) + ((g127) & (g147) & (g2025) & (!g2026) & (!g2033)) + ((g127) & (g147) & (g2025) & (!g2026) & (g2033)) + ((g127) & (g147) & (g2025) & (g2026) & (!g2033)) + ((g127) & (g147) & (g2025) & (g2026) & (g2033)));
	assign g2035 = (((!g87) & (!g104) & (g2022) & (g2023) & (g2034)) + ((!g87) & (g104) & (g2022) & (!g2023) & (g2034)) + ((!g87) & (g104) & (g2022) & (g2023) & (!g2034)) + ((!g87) & (g104) & (g2022) & (g2023) & (g2034)) + ((g87) & (!g104) & (!g2022) & (g2023) & (g2034)) + ((g87) & (!g104) & (g2022) & (!g2023) & (!g2034)) + ((g87) & (!g104) & (g2022) & (!g2023) & (g2034)) + ((g87) & (!g104) & (g2022) & (g2023) & (!g2034)) + ((g87) & (!g104) & (g2022) & (g2023) & (g2034)) + ((g87) & (g104) & (!g2022) & (!g2023) & (g2034)) + ((g87) & (g104) & (!g2022) & (g2023) & (!g2034)) + ((g87) & (g104) & (!g2022) & (g2023) & (g2034)) + ((g87) & (g104) & (g2022) & (!g2023) & (!g2034)) + ((g87) & (g104) & (g2022) & (!g2023) & (g2034)) + ((g87) & (g104) & (g2022) & (g2023) & (!g2034)) + ((g87) & (g104) & (g2022) & (g2023) & (g2034)));
	assign g2036 = (((!g54) & (!g68) & (g2019) & (g2020) & (g2035)) + ((!g54) & (g68) & (g2019) & (!g2020) & (g2035)) + ((!g54) & (g68) & (g2019) & (g2020) & (!g2035)) + ((!g54) & (g68) & (g2019) & (g2020) & (g2035)) + ((g54) & (!g68) & (!g2019) & (g2020) & (g2035)) + ((g54) & (!g68) & (g2019) & (!g2020) & (!g2035)) + ((g54) & (!g68) & (g2019) & (!g2020) & (g2035)) + ((g54) & (!g68) & (g2019) & (g2020) & (!g2035)) + ((g54) & (!g68) & (g2019) & (g2020) & (g2035)) + ((g54) & (g68) & (!g2019) & (!g2020) & (g2035)) + ((g54) & (g68) & (!g2019) & (g2020) & (!g2035)) + ((g54) & (g68) & (!g2019) & (g2020) & (g2035)) + ((g54) & (g68) & (g2019) & (!g2020) & (!g2035)) + ((g54) & (g68) & (g2019) & (!g2020) & (g2035)) + ((g54) & (g68) & (g2019) & (g2020) & (!g2035)) + ((g54) & (g68) & (g2019) & (g2020) & (g2035)));
	assign g2037 = (((!g27) & (!g39) & (g2016) & (g2017) & (g2036)) + ((!g27) & (g39) & (g2016) & (!g2017) & (g2036)) + ((!g27) & (g39) & (g2016) & (g2017) & (!g2036)) + ((!g27) & (g39) & (g2016) & (g2017) & (g2036)) + ((g27) & (!g39) & (!g2016) & (g2017) & (g2036)) + ((g27) & (!g39) & (g2016) & (!g2017) & (!g2036)) + ((g27) & (!g39) & (g2016) & (!g2017) & (g2036)) + ((g27) & (!g39) & (g2016) & (g2017) & (!g2036)) + ((g27) & (!g39) & (g2016) & (g2017) & (g2036)) + ((g27) & (g39) & (!g2016) & (!g2017) & (g2036)) + ((g27) & (g39) & (!g2016) & (g2017) & (!g2036)) + ((g27) & (g39) & (!g2016) & (g2017) & (g2036)) + ((g27) & (g39) & (g2016) & (!g2017) & (!g2036)) + ((g27) & (g39) & (g2016) & (!g2017) & (g2036)) + ((g27) & (g39) & (g2016) & (g2017) & (!g2036)) + ((g27) & (g39) & (g2016) & (g2017) & (g2036)));
	assign g2038 = (((!g8) & (!g18) & (g2013) & (g2014) & (g2037)) + ((!g8) & (g18) & (g2013) & (!g2014) & (g2037)) + ((!g8) & (g18) & (g2013) & (g2014) & (!g2037)) + ((!g8) & (g18) & (g2013) & (g2014) & (g2037)) + ((g8) & (!g18) & (!g2013) & (g2014) & (g2037)) + ((g8) & (!g18) & (g2013) & (!g2014) & (!g2037)) + ((g8) & (!g18) & (g2013) & (!g2014) & (g2037)) + ((g8) & (!g18) & (g2013) & (g2014) & (!g2037)) + ((g8) & (!g18) & (g2013) & (g2014) & (g2037)) + ((g8) & (g18) & (!g2013) & (!g2014) & (g2037)) + ((g8) & (g18) & (!g2013) & (g2014) & (!g2037)) + ((g8) & (g18) & (!g2013) & (g2014) & (g2037)) + ((g8) & (g18) & (g2013) & (!g2014) & (!g2037)) + ((g8) & (g18) & (g2013) & (!g2014) & (g2037)) + ((g8) & (g18) & (g2013) & (g2014) & (!g2037)) + ((g8) & (g18) & (g2013) & (g2014) & (g2037)));
	assign g2039 = (((!g2) & (!g8) & (g1926) & (g1946)) + ((!g2) & (g8) & (!g1926) & (g1946)) + ((!g2) & (g8) & (g1926) & (!g1946)) + ((!g2) & (g8) & (g1926) & (g1946)) + ((g2) & (!g8) & (!g1926) & (!g1946)) + ((g2) & (!g8) & (!g1926) & (g1946)) + ((g2) & (!g8) & (g1926) & (!g1946)) + ((g2) & (g8) & (!g1926) & (!g1946)));
	assign g2040 = (((!g1925) & (!g1923) & (!g1950) & (g2039)) + ((!g1925) & (g1923) & (!g1950) & (g2039)) + ((!g1925) & (g1923) & (g1950) & (g2039)) + ((g1925) & (!g1923) & (!g1950) & (!g2039)) + ((g1925) & (!g1923) & (g1950) & (!g2039)) + ((g1925) & (!g1923) & (g1950) & (g2039)) + ((g1925) & (g1923) & (!g1950) & (!g2039)) + ((g1925) & (g1923) & (g1950) & (!g2039)));
	assign g2041 = (((!g4) & (!g2) & (!g2011) & (!g2038) & (g2040)) + ((!g4) & (!g2) & (!g2011) & (g2038) & (g2040)) + ((!g4) & (!g2) & (g2011) & (!g2038) & (g2040)) + ((!g4) & (!g2) & (g2011) & (g2038) & (!g2040)) + ((!g4) & (!g2) & (g2011) & (g2038) & (g2040)) + ((!g4) & (g2) & (!g2011) & (!g2038) & (g2040)) + ((!g4) & (g2) & (!g2011) & (g2038) & (!g2040)) + ((!g4) & (g2) & (!g2011) & (g2038) & (g2040)) + ((!g4) & (g2) & (g2011) & (!g2038) & (!g2040)) + ((!g4) & (g2) & (g2011) & (!g2038) & (g2040)) + ((!g4) & (g2) & (g2011) & (g2038) & (!g2040)) + ((!g4) & (g2) & (g2011) & (g2038) & (g2040)) + ((g4) & (!g2) & (g2011) & (g2038) & (g2040)) + ((g4) & (g2) & (!g2011) & (g2038) & (g2040)) + ((g4) & (g2) & (g2011) & (!g2038) & (g2040)) + ((g4) & (g2) & (g2011) & (g2038) & (g2040)));
	assign g2042 = (((!g4) & (!g1947) & (g1948)) + ((!g4) & (g1947) & (!g1948)) + ((!g4) & (g1947) & (g1948)) + ((g4) & (g1947) & (g1948)));
	assign g2043 = (((!g1924) & (!g2042) & (!g1923) & (!g1950)) + ((!g1924) & (!g2042) & (g1923) & (!g1950)) + ((!g1924) & (!g2042) & (g1923) & (g1950)) + ((g1924) & (g2042) & (!g1923) & (!g1950)) + ((g1924) & (g2042) & (!g1923) & (g1950)) + ((g1924) & (g2042) & (g1923) & (!g1950)) + ((g1924) & (g2042) & (g1923) & (g1950)));
	assign g2044 = (((!g1) & (g1924) & (!g2042) & (!g1923) & (g1950)) + ((!g1) & (g1924) & (g2042) & (!g1923) & (g1950)) + ((g1) & (!g1924) & (g2042) & (g1923) & (!g1950)) + ((g1) & (!g1924) & (g2042) & (g1923) & (g1950)) + ((g1) & (g1924) & (!g2042) & (!g1923) & (!g1950)) + ((g1) & (g1924) & (!g2042) & (!g1923) & (g1950)) + ((g1) & (g1924) & (!g2042) & (g1923) & (!g1950)) + ((g1) & (g1924) & (!g2042) & (g1923) & (g1950)) + ((g1) & (g1924) & (g2042) & (!g1923) & (g1950)));
	assign g2045 = (((!g1) & (!g2010) & (!g2041) & (!g2043) & (!g2044)) + ((g1) & (!g2010) & (!g2041) & (!g2043) & (!g2044)) + ((g1) & (!g2010) & (!g2041) & (g2043) & (!g2044)) + ((g1) & (!g2010) & (g2041) & (!g2043) & (!g2044)) + ((g1) & (!g2010) & (g2041) & (g2043) & (!g2044)) + ((g1) & (g2010) & (!g2041) & (!g2043) & (!g2044)) + ((g1) & (g2010) & (!g2041) & (g2043) & (!g2044)));
	assign g2046 = (((!g255) & (!g1951) & (g2009) & (!g2045)) + ((!g255) & (g1951) & (!g2009) & (!g2045)) + ((!g255) & (g1951) & (!g2009) & (g2045)) + ((!g255) & (g1951) & (g2009) & (g2045)) + ((g255) & (!g1951) & (!g2009) & (!g2045)) + ((g255) & (g1951) & (!g2009) & (g2045)) + ((g255) & (g1951) & (g2009) & (!g2045)) + ((g255) & (g1951) & (g2009) & (g2045)));
	assign g2047 = (((!g290) & (!g319) & (!g1953) & (g1954) & (g2008) & (!g2045)) + ((!g290) & (!g319) & (g1953) & (!g1954) & (!g2008) & (!g2045)) + ((!g290) & (!g319) & (g1953) & (!g1954) & (!g2008) & (g2045)) + ((!g290) & (!g319) & (g1953) & (!g1954) & (g2008) & (!g2045)) + ((!g290) & (!g319) & (g1953) & (!g1954) & (g2008) & (g2045)) + ((!g290) & (!g319) & (g1953) & (g1954) & (!g2008) & (!g2045)) + ((!g290) & (!g319) & (g1953) & (g1954) & (!g2008) & (g2045)) + ((!g290) & (!g319) & (g1953) & (g1954) & (g2008) & (g2045)) + ((!g290) & (g319) & (!g1953) & (!g1954) & (g2008) & (!g2045)) + ((!g290) & (g319) & (!g1953) & (g1954) & (!g2008) & (!g2045)) + ((!g290) & (g319) & (!g1953) & (g1954) & (g2008) & (!g2045)) + ((!g290) & (g319) & (g1953) & (!g1954) & (!g2008) & (!g2045)) + ((!g290) & (g319) & (g1953) & (!g1954) & (!g2008) & (g2045)) + ((!g290) & (g319) & (g1953) & (!g1954) & (g2008) & (g2045)) + ((!g290) & (g319) & (g1953) & (g1954) & (!g2008) & (g2045)) + ((!g290) & (g319) & (g1953) & (g1954) & (g2008) & (g2045)) + ((g290) & (!g319) & (!g1953) & (!g1954) & (!g2008) & (!g2045)) + ((g290) & (!g319) & (!g1953) & (!g1954) & (g2008) & (!g2045)) + ((g290) & (!g319) & (!g1953) & (g1954) & (!g2008) & (!g2045)) + ((g290) & (!g319) & (g1953) & (!g1954) & (!g2008) & (g2045)) + ((g290) & (!g319) & (g1953) & (!g1954) & (g2008) & (g2045)) + ((g290) & (!g319) & (g1953) & (g1954) & (!g2008) & (g2045)) + ((g290) & (!g319) & (g1953) & (g1954) & (g2008) & (!g2045)) + ((g290) & (!g319) & (g1953) & (g1954) & (g2008) & (g2045)) + ((g290) & (g319) & (!g1953) & (!g1954) & (!g2008) & (!g2045)) + ((g290) & (g319) & (g1953) & (!g1954) & (!g2008) & (g2045)) + ((g290) & (g319) & (g1953) & (!g1954) & (g2008) & (!g2045)) + ((g290) & (g319) & (g1953) & (!g1954) & (g2008) & (g2045)) + ((g290) & (g319) & (g1953) & (g1954) & (!g2008) & (!g2045)) + ((g290) & (g319) & (g1953) & (g1954) & (!g2008) & (g2045)) + ((g290) & (g319) & (g1953) & (g1954) & (g2008) & (!g2045)) + ((g290) & (g319) & (g1953) & (g1954) & (g2008) & (g2045)));
	assign g2048 = (((!g319) & (!g1954) & (g2008) & (!g2045)) + ((!g319) & (g1954) & (!g2008) & (!g2045)) + ((!g319) & (g1954) & (!g2008) & (g2045)) + ((!g319) & (g1954) & (g2008) & (g2045)) + ((g319) & (!g1954) & (!g2008) & (!g2045)) + ((g319) & (g1954) & (!g2008) & (g2045)) + ((g319) & (g1954) & (g2008) & (!g2045)) + ((g319) & (g1954) & (g2008) & (g2045)));
	assign g2049 = (((!g358) & (!g390) & (!g1956) & (g1957) & (g2007) & (!g2045)) + ((!g358) & (!g390) & (g1956) & (!g1957) & (!g2007) & (!g2045)) + ((!g358) & (!g390) & (g1956) & (!g1957) & (!g2007) & (g2045)) + ((!g358) & (!g390) & (g1956) & (!g1957) & (g2007) & (!g2045)) + ((!g358) & (!g390) & (g1956) & (!g1957) & (g2007) & (g2045)) + ((!g358) & (!g390) & (g1956) & (g1957) & (!g2007) & (!g2045)) + ((!g358) & (!g390) & (g1956) & (g1957) & (!g2007) & (g2045)) + ((!g358) & (!g390) & (g1956) & (g1957) & (g2007) & (g2045)) + ((!g358) & (g390) & (!g1956) & (!g1957) & (g2007) & (!g2045)) + ((!g358) & (g390) & (!g1956) & (g1957) & (!g2007) & (!g2045)) + ((!g358) & (g390) & (!g1956) & (g1957) & (g2007) & (!g2045)) + ((!g358) & (g390) & (g1956) & (!g1957) & (!g2007) & (!g2045)) + ((!g358) & (g390) & (g1956) & (!g1957) & (!g2007) & (g2045)) + ((!g358) & (g390) & (g1956) & (!g1957) & (g2007) & (g2045)) + ((!g358) & (g390) & (g1956) & (g1957) & (!g2007) & (g2045)) + ((!g358) & (g390) & (g1956) & (g1957) & (g2007) & (g2045)) + ((g358) & (!g390) & (!g1956) & (!g1957) & (!g2007) & (!g2045)) + ((g358) & (!g390) & (!g1956) & (!g1957) & (g2007) & (!g2045)) + ((g358) & (!g390) & (!g1956) & (g1957) & (!g2007) & (!g2045)) + ((g358) & (!g390) & (g1956) & (!g1957) & (!g2007) & (g2045)) + ((g358) & (!g390) & (g1956) & (!g1957) & (g2007) & (g2045)) + ((g358) & (!g390) & (g1956) & (g1957) & (!g2007) & (g2045)) + ((g358) & (!g390) & (g1956) & (g1957) & (g2007) & (!g2045)) + ((g358) & (!g390) & (g1956) & (g1957) & (g2007) & (g2045)) + ((g358) & (g390) & (!g1956) & (!g1957) & (!g2007) & (!g2045)) + ((g358) & (g390) & (g1956) & (!g1957) & (!g2007) & (g2045)) + ((g358) & (g390) & (g1956) & (!g1957) & (g2007) & (!g2045)) + ((g358) & (g390) & (g1956) & (!g1957) & (g2007) & (g2045)) + ((g358) & (g390) & (g1956) & (g1957) & (!g2007) & (!g2045)) + ((g358) & (g390) & (g1956) & (g1957) & (!g2007) & (g2045)) + ((g358) & (g390) & (g1956) & (g1957) & (g2007) & (!g2045)) + ((g358) & (g390) & (g1956) & (g1957) & (g2007) & (g2045)));
	assign g2050 = (((!g390) & (!g1957) & (g2007) & (!g2045)) + ((!g390) & (g1957) & (!g2007) & (!g2045)) + ((!g390) & (g1957) & (!g2007) & (g2045)) + ((!g390) & (g1957) & (g2007) & (g2045)) + ((g390) & (!g1957) & (!g2007) & (!g2045)) + ((g390) & (g1957) & (!g2007) & (g2045)) + ((g390) & (g1957) & (g2007) & (!g2045)) + ((g390) & (g1957) & (g2007) & (g2045)));
	assign g2051 = (((!g433) & (!g468) & (!g1959) & (g1960) & (g2006) & (!g2045)) + ((!g433) & (!g468) & (g1959) & (!g1960) & (!g2006) & (!g2045)) + ((!g433) & (!g468) & (g1959) & (!g1960) & (!g2006) & (g2045)) + ((!g433) & (!g468) & (g1959) & (!g1960) & (g2006) & (!g2045)) + ((!g433) & (!g468) & (g1959) & (!g1960) & (g2006) & (g2045)) + ((!g433) & (!g468) & (g1959) & (g1960) & (!g2006) & (!g2045)) + ((!g433) & (!g468) & (g1959) & (g1960) & (!g2006) & (g2045)) + ((!g433) & (!g468) & (g1959) & (g1960) & (g2006) & (g2045)) + ((!g433) & (g468) & (!g1959) & (!g1960) & (g2006) & (!g2045)) + ((!g433) & (g468) & (!g1959) & (g1960) & (!g2006) & (!g2045)) + ((!g433) & (g468) & (!g1959) & (g1960) & (g2006) & (!g2045)) + ((!g433) & (g468) & (g1959) & (!g1960) & (!g2006) & (!g2045)) + ((!g433) & (g468) & (g1959) & (!g1960) & (!g2006) & (g2045)) + ((!g433) & (g468) & (g1959) & (!g1960) & (g2006) & (g2045)) + ((!g433) & (g468) & (g1959) & (g1960) & (!g2006) & (g2045)) + ((!g433) & (g468) & (g1959) & (g1960) & (g2006) & (g2045)) + ((g433) & (!g468) & (!g1959) & (!g1960) & (!g2006) & (!g2045)) + ((g433) & (!g468) & (!g1959) & (!g1960) & (g2006) & (!g2045)) + ((g433) & (!g468) & (!g1959) & (g1960) & (!g2006) & (!g2045)) + ((g433) & (!g468) & (g1959) & (!g1960) & (!g2006) & (g2045)) + ((g433) & (!g468) & (g1959) & (!g1960) & (g2006) & (g2045)) + ((g433) & (!g468) & (g1959) & (g1960) & (!g2006) & (g2045)) + ((g433) & (!g468) & (g1959) & (g1960) & (g2006) & (!g2045)) + ((g433) & (!g468) & (g1959) & (g1960) & (g2006) & (g2045)) + ((g433) & (g468) & (!g1959) & (!g1960) & (!g2006) & (!g2045)) + ((g433) & (g468) & (g1959) & (!g1960) & (!g2006) & (g2045)) + ((g433) & (g468) & (g1959) & (!g1960) & (g2006) & (!g2045)) + ((g433) & (g468) & (g1959) & (!g1960) & (g2006) & (g2045)) + ((g433) & (g468) & (g1959) & (g1960) & (!g2006) & (!g2045)) + ((g433) & (g468) & (g1959) & (g1960) & (!g2006) & (g2045)) + ((g433) & (g468) & (g1959) & (g1960) & (g2006) & (!g2045)) + ((g433) & (g468) & (g1959) & (g1960) & (g2006) & (g2045)));
	assign g2052 = (((!g468) & (!g1960) & (g2006) & (!g2045)) + ((!g468) & (g1960) & (!g2006) & (!g2045)) + ((!g468) & (g1960) & (!g2006) & (g2045)) + ((!g468) & (g1960) & (g2006) & (g2045)) + ((g468) & (!g1960) & (!g2006) & (!g2045)) + ((g468) & (g1960) & (!g2006) & (g2045)) + ((g468) & (g1960) & (g2006) & (!g2045)) + ((g468) & (g1960) & (g2006) & (g2045)));
	assign g2053 = (((!g515) & (!g553) & (!g1962) & (g1963) & (g2005) & (!g2045)) + ((!g515) & (!g553) & (g1962) & (!g1963) & (!g2005) & (!g2045)) + ((!g515) & (!g553) & (g1962) & (!g1963) & (!g2005) & (g2045)) + ((!g515) & (!g553) & (g1962) & (!g1963) & (g2005) & (!g2045)) + ((!g515) & (!g553) & (g1962) & (!g1963) & (g2005) & (g2045)) + ((!g515) & (!g553) & (g1962) & (g1963) & (!g2005) & (!g2045)) + ((!g515) & (!g553) & (g1962) & (g1963) & (!g2005) & (g2045)) + ((!g515) & (!g553) & (g1962) & (g1963) & (g2005) & (g2045)) + ((!g515) & (g553) & (!g1962) & (!g1963) & (g2005) & (!g2045)) + ((!g515) & (g553) & (!g1962) & (g1963) & (!g2005) & (!g2045)) + ((!g515) & (g553) & (!g1962) & (g1963) & (g2005) & (!g2045)) + ((!g515) & (g553) & (g1962) & (!g1963) & (!g2005) & (!g2045)) + ((!g515) & (g553) & (g1962) & (!g1963) & (!g2005) & (g2045)) + ((!g515) & (g553) & (g1962) & (!g1963) & (g2005) & (g2045)) + ((!g515) & (g553) & (g1962) & (g1963) & (!g2005) & (g2045)) + ((!g515) & (g553) & (g1962) & (g1963) & (g2005) & (g2045)) + ((g515) & (!g553) & (!g1962) & (!g1963) & (!g2005) & (!g2045)) + ((g515) & (!g553) & (!g1962) & (!g1963) & (g2005) & (!g2045)) + ((g515) & (!g553) & (!g1962) & (g1963) & (!g2005) & (!g2045)) + ((g515) & (!g553) & (g1962) & (!g1963) & (!g2005) & (g2045)) + ((g515) & (!g553) & (g1962) & (!g1963) & (g2005) & (g2045)) + ((g515) & (!g553) & (g1962) & (g1963) & (!g2005) & (g2045)) + ((g515) & (!g553) & (g1962) & (g1963) & (g2005) & (!g2045)) + ((g515) & (!g553) & (g1962) & (g1963) & (g2005) & (g2045)) + ((g515) & (g553) & (!g1962) & (!g1963) & (!g2005) & (!g2045)) + ((g515) & (g553) & (g1962) & (!g1963) & (!g2005) & (g2045)) + ((g515) & (g553) & (g1962) & (!g1963) & (g2005) & (!g2045)) + ((g515) & (g553) & (g1962) & (!g1963) & (g2005) & (g2045)) + ((g515) & (g553) & (g1962) & (g1963) & (!g2005) & (!g2045)) + ((g515) & (g553) & (g1962) & (g1963) & (!g2005) & (g2045)) + ((g515) & (g553) & (g1962) & (g1963) & (g2005) & (!g2045)) + ((g515) & (g553) & (g1962) & (g1963) & (g2005) & (g2045)));
	assign g2054 = (((!g553) & (!g1963) & (g2005) & (!g2045)) + ((!g553) & (g1963) & (!g2005) & (!g2045)) + ((!g553) & (g1963) & (!g2005) & (g2045)) + ((!g553) & (g1963) & (g2005) & (g2045)) + ((g553) & (!g1963) & (!g2005) & (!g2045)) + ((g553) & (g1963) & (!g2005) & (g2045)) + ((g553) & (g1963) & (g2005) & (!g2045)) + ((g553) & (g1963) & (g2005) & (g2045)));
	assign g2055 = (((!g604) & (!g645) & (!g1965) & (g1966) & (g2004) & (!g2045)) + ((!g604) & (!g645) & (g1965) & (!g1966) & (!g2004) & (!g2045)) + ((!g604) & (!g645) & (g1965) & (!g1966) & (!g2004) & (g2045)) + ((!g604) & (!g645) & (g1965) & (!g1966) & (g2004) & (!g2045)) + ((!g604) & (!g645) & (g1965) & (!g1966) & (g2004) & (g2045)) + ((!g604) & (!g645) & (g1965) & (g1966) & (!g2004) & (!g2045)) + ((!g604) & (!g645) & (g1965) & (g1966) & (!g2004) & (g2045)) + ((!g604) & (!g645) & (g1965) & (g1966) & (g2004) & (g2045)) + ((!g604) & (g645) & (!g1965) & (!g1966) & (g2004) & (!g2045)) + ((!g604) & (g645) & (!g1965) & (g1966) & (!g2004) & (!g2045)) + ((!g604) & (g645) & (!g1965) & (g1966) & (g2004) & (!g2045)) + ((!g604) & (g645) & (g1965) & (!g1966) & (!g2004) & (!g2045)) + ((!g604) & (g645) & (g1965) & (!g1966) & (!g2004) & (g2045)) + ((!g604) & (g645) & (g1965) & (!g1966) & (g2004) & (g2045)) + ((!g604) & (g645) & (g1965) & (g1966) & (!g2004) & (g2045)) + ((!g604) & (g645) & (g1965) & (g1966) & (g2004) & (g2045)) + ((g604) & (!g645) & (!g1965) & (!g1966) & (!g2004) & (!g2045)) + ((g604) & (!g645) & (!g1965) & (!g1966) & (g2004) & (!g2045)) + ((g604) & (!g645) & (!g1965) & (g1966) & (!g2004) & (!g2045)) + ((g604) & (!g645) & (g1965) & (!g1966) & (!g2004) & (g2045)) + ((g604) & (!g645) & (g1965) & (!g1966) & (g2004) & (g2045)) + ((g604) & (!g645) & (g1965) & (g1966) & (!g2004) & (g2045)) + ((g604) & (!g645) & (g1965) & (g1966) & (g2004) & (!g2045)) + ((g604) & (!g645) & (g1965) & (g1966) & (g2004) & (g2045)) + ((g604) & (g645) & (!g1965) & (!g1966) & (!g2004) & (!g2045)) + ((g604) & (g645) & (g1965) & (!g1966) & (!g2004) & (g2045)) + ((g604) & (g645) & (g1965) & (!g1966) & (g2004) & (!g2045)) + ((g604) & (g645) & (g1965) & (!g1966) & (g2004) & (g2045)) + ((g604) & (g645) & (g1965) & (g1966) & (!g2004) & (!g2045)) + ((g604) & (g645) & (g1965) & (g1966) & (!g2004) & (g2045)) + ((g604) & (g645) & (g1965) & (g1966) & (g2004) & (!g2045)) + ((g604) & (g645) & (g1965) & (g1966) & (g2004) & (g2045)));
	assign g2056 = (((!g645) & (!g1966) & (g2004) & (!g2045)) + ((!g645) & (g1966) & (!g2004) & (!g2045)) + ((!g645) & (g1966) & (!g2004) & (g2045)) + ((!g645) & (g1966) & (g2004) & (g2045)) + ((g645) & (!g1966) & (!g2004) & (!g2045)) + ((g645) & (g1966) & (!g2004) & (g2045)) + ((g645) & (g1966) & (g2004) & (!g2045)) + ((g645) & (g1966) & (g2004) & (g2045)));
	assign g2057 = (((!g700) & (!g744) & (!g1968) & (g1969) & (g2003) & (!g2045)) + ((!g700) & (!g744) & (g1968) & (!g1969) & (!g2003) & (!g2045)) + ((!g700) & (!g744) & (g1968) & (!g1969) & (!g2003) & (g2045)) + ((!g700) & (!g744) & (g1968) & (!g1969) & (g2003) & (!g2045)) + ((!g700) & (!g744) & (g1968) & (!g1969) & (g2003) & (g2045)) + ((!g700) & (!g744) & (g1968) & (g1969) & (!g2003) & (!g2045)) + ((!g700) & (!g744) & (g1968) & (g1969) & (!g2003) & (g2045)) + ((!g700) & (!g744) & (g1968) & (g1969) & (g2003) & (g2045)) + ((!g700) & (g744) & (!g1968) & (!g1969) & (g2003) & (!g2045)) + ((!g700) & (g744) & (!g1968) & (g1969) & (!g2003) & (!g2045)) + ((!g700) & (g744) & (!g1968) & (g1969) & (g2003) & (!g2045)) + ((!g700) & (g744) & (g1968) & (!g1969) & (!g2003) & (!g2045)) + ((!g700) & (g744) & (g1968) & (!g1969) & (!g2003) & (g2045)) + ((!g700) & (g744) & (g1968) & (!g1969) & (g2003) & (g2045)) + ((!g700) & (g744) & (g1968) & (g1969) & (!g2003) & (g2045)) + ((!g700) & (g744) & (g1968) & (g1969) & (g2003) & (g2045)) + ((g700) & (!g744) & (!g1968) & (!g1969) & (!g2003) & (!g2045)) + ((g700) & (!g744) & (!g1968) & (!g1969) & (g2003) & (!g2045)) + ((g700) & (!g744) & (!g1968) & (g1969) & (!g2003) & (!g2045)) + ((g700) & (!g744) & (g1968) & (!g1969) & (!g2003) & (g2045)) + ((g700) & (!g744) & (g1968) & (!g1969) & (g2003) & (g2045)) + ((g700) & (!g744) & (g1968) & (g1969) & (!g2003) & (g2045)) + ((g700) & (!g744) & (g1968) & (g1969) & (g2003) & (!g2045)) + ((g700) & (!g744) & (g1968) & (g1969) & (g2003) & (g2045)) + ((g700) & (g744) & (!g1968) & (!g1969) & (!g2003) & (!g2045)) + ((g700) & (g744) & (g1968) & (!g1969) & (!g2003) & (g2045)) + ((g700) & (g744) & (g1968) & (!g1969) & (g2003) & (!g2045)) + ((g700) & (g744) & (g1968) & (!g1969) & (g2003) & (g2045)) + ((g700) & (g744) & (g1968) & (g1969) & (!g2003) & (!g2045)) + ((g700) & (g744) & (g1968) & (g1969) & (!g2003) & (g2045)) + ((g700) & (g744) & (g1968) & (g1969) & (g2003) & (!g2045)) + ((g700) & (g744) & (g1968) & (g1969) & (g2003) & (g2045)));
	assign g2058 = (((!g744) & (!g1969) & (g2003) & (!g2045)) + ((!g744) & (g1969) & (!g2003) & (!g2045)) + ((!g744) & (g1969) & (!g2003) & (g2045)) + ((!g744) & (g1969) & (g2003) & (g2045)) + ((g744) & (!g1969) & (!g2003) & (!g2045)) + ((g744) & (g1969) & (!g2003) & (g2045)) + ((g744) & (g1969) & (g2003) & (!g2045)) + ((g744) & (g1969) & (g2003) & (g2045)));
	assign g2059 = (((!g803) & (!g851) & (!g1971) & (g1972) & (g2002) & (!g2045)) + ((!g803) & (!g851) & (g1971) & (!g1972) & (!g2002) & (!g2045)) + ((!g803) & (!g851) & (g1971) & (!g1972) & (!g2002) & (g2045)) + ((!g803) & (!g851) & (g1971) & (!g1972) & (g2002) & (!g2045)) + ((!g803) & (!g851) & (g1971) & (!g1972) & (g2002) & (g2045)) + ((!g803) & (!g851) & (g1971) & (g1972) & (!g2002) & (!g2045)) + ((!g803) & (!g851) & (g1971) & (g1972) & (!g2002) & (g2045)) + ((!g803) & (!g851) & (g1971) & (g1972) & (g2002) & (g2045)) + ((!g803) & (g851) & (!g1971) & (!g1972) & (g2002) & (!g2045)) + ((!g803) & (g851) & (!g1971) & (g1972) & (!g2002) & (!g2045)) + ((!g803) & (g851) & (!g1971) & (g1972) & (g2002) & (!g2045)) + ((!g803) & (g851) & (g1971) & (!g1972) & (!g2002) & (!g2045)) + ((!g803) & (g851) & (g1971) & (!g1972) & (!g2002) & (g2045)) + ((!g803) & (g851) & (g1971) & (!g1972) & (g2002) & (g2045)) + ((!g803) & (g851) & (g1971) & (g1972) & (!g2002) & (g2045)) + ((!g803) & (g851) & (g1971) & (g1972) & (g2002) & (g2045)) + ((g803) & (!g851) & (!g1971) & (!g1972) & (!g2002) & (!g2045)) + ((g803) & (!g851) & (!g1971) & (!g1972) & (g2002) & (!g2045)) + ((g803) & (!g851) & (!g1971) & (g1972) & (!g2002) & (!g2045)) + ((g803) & (!g851) & (g1971) & (!g1972) & (!g2002) & (g2045)) + ((g803) & (!g851) & (g1971) & (!g1972) & (g2002) & (g2045)) + ((g803) & (!g851) & (g1971) & (g1972) & (!g2002) & (g2045)) + ((g803) & (!g851) & (g1971) & (g1972) & (g2002) & (!g2045)) + ((g803) & (!g851) & (g1971) & (g1972) & (g2002) & (g2045)) + ((g803) & (g851) & (!g1971) & (!g1972) & (!g2002) & (!g2045)) + ((g803) & (g851) & (g1971) & (!g1972) & (!g2002) & (g2045)) + ((g803) & (g851) & (g1971) & (!g1972) & (g2002) & (!g2045)) + ((g803) & (g851) & (g1971) & (!g1972) & (g2002) & (g2045)) + ((g803) & (g851) & (g1971) & (g1972) & (!g2002) & (!g2045)) + ((g803) & (g851) & (g1971) & (g1972) & (!g2002) & (g2045)) + ((g803) & (g851) & (g1971) & (g1972) & (g2002) & (!g2045)) + ((g803) & (g851) & (g1971) & (g1972) & (g2002) & (g2045)));
	assign g2060 = (((!g851) & (!g1972) & (g2002) & (!g2045)) + ((!g851) & (g1972) & (!g2002) & (!g2045)) + ((!g851) & (g1972) & (!g2002) & (g2045)) + ((!g851) & (g1972) & (g2002) & (g2045)) + ((g851) & (!g1972) & (!g2002) & (!g2045)) + ((g851) & (g1972) & (!g2002) & (g2045)) + ((g851) & (g1972) & (g2002) & (!g2045)) + ((g851) & (g1972) & (g2002) & (g2045)));
	assign g2061 = (((!g914) & (!g1032) & (!g1974) & (g1975) & (g2001) & (!g2045)) + ((!g914) & (!g1032) & (g1974) & (!g1975) & (!g2001) & (!g2045)) + ((!g914) & (!g1032) & (g1974) & (!g1975) & (!g2001) & (g2045)) + ((!g914) & (!g1032) & (g1974) & (!g1975) & (g2001) & (!g2045)) + ((!g914) & (!g1032) & (g1974) & (!g1975) & (g2001) & (g2045)) + ((!g914) & (!g1032) & (g1974) & (g1975) & (!g2001) & (!g2045)) + ((!g914) & (!g1032) & (g1974) & (g1975) & (!g2001) & (g2045)) + ((!g914) & (!g1032) & (g1974) & (g1975) & (g2001) & (g2045)) + ((!g914) & (g1032) & (!g1974) & (!g1975) & (g2001) & (!g2045)) + ((!g914) & (g1032) & (!g1974) & (g1975) & (!g2001) & (!g2045)) + ((!g914) & (g1032) & (!g1974) & (g1975) & (g2001) & (!g2045)) + ((!g914) & (g1032) & (g1974) & (!g1975) & (!g2001) & (!g2045)) + ((!g914) & (g1032) & (g1974) & (!g1975) & (!g2001) & (g2045)) + ((!g914) & (g1032) & (g1974) & (!g1975) & (g2001) & (g2045)) + ((!g914) & (g1032) & (g1974) & (g1975) & (!g2001) & (g2045)) + ((!g914) & (g1032) & (g1974) & (g1975) & (g2001) & (g2045)) + ((g914) & (!g1032) & (!g1974) & (!g1975) & (!g2001) & (!g2045)) + ((g914) & (!g1032) & (!g1974) & (!g1975) & (g2001) & (!g2045)) + ((g914) & (!g1032) & (!g1974) & (g1975) & (!g2001) & (!g2045)) + ((g914) & (!g1032) & (g1974) & (!g1975) & (!g2001) & (g2045)) + ((g914) & (!g1032) & (g1974) & (!g1975) & (g2001) & (g2045)) + ((g914) & (!g1032) & (g1974) & (g1975) & (!g2001) & (g2045)) + ((g914) & (!g1032) & (g1974) & (g1975) & (g2001) & (!g2045)) + ((g914) & (!g1032) & (g1974) & (g1975) & (g2001) & (g2045)) + ((g914) & (g1032) & (!g1974) & (!g1975) & (!g2001) & (!g2045)) + ((g914) & (g1032) & (g1974) & (!g1975) & (!g2001) & (g2045)) + ((g914) & (g1032) & (g1974) & (!g1975) & (g2001) & (!g2045)) + ((g914) & (g1032) & (g1974) & (!g1975) & (g2001) & (g2045)) + ((g914) & (g1032) & (g1974) & (g1975) & (!g2001) & (!g2045)) + ((g914) & (g1032) & (g1974) & (g1975) & (!g2001) & (g2045)) + ((g914) & (g1032) & (g1974) & (g1975) & (g2001) & (!g2045)) + ((g914) & (g1032) & (g1974) & (g1975) & (g2001) & (g2045)));
	assign g2062 = (((!g1032) & (!g1975) & (g2001) & (!g2045)) + ((!g1032) & (g1975) & (!g2001) & (!g2045)) + ((!g1032) & (g1975) & (!g2001) & (g2045)) + ((!g1032) & (g1975) & (g2001) & (g2045)) + ((g1032) & (!g1975) & (!g2001) & (!g2045)) + ((g1032) & (g1975) & (!g2001) & (g2045)) + ((g1032) & (g1975) & (g2001) & (!g2045)) + ((g1032) & (g1975) & (g2001) & (g2045)));
	assign g2063 = (((!g1030) & (!g1160) & (!g1977) & (g1978) & (g2000) & (!g2045)) + ((!g1030) & (!g1160) & (g1977) & (!g1978) & (!g2000) & (!g2045)) + ((!g1030) & (!g1160) & (g1977) & (!g1978) & (!g2000) & (g2045)) + ((!g1030) & (!g1160) & (g1977) & (!g1978) & (g2000) & (!g2045)) + ((!g1030) & (!g1160) & (g1977) & (!g1978) & (g2000) & (g2045)) + ((!g1030) & (!g1160) & (g1977) & (g1978) & (!g2000) & (!g2045)) + ((!g1030) & (!g1160) & (g1977) & (g1978) & (!g2000) & (g2045)) + ((!g1030) & (!g1160) & (g1977) & (g1978) & (g2000) & (g2045)) + ((!g1030) & (g1160) & (!g1977) & (!g1978) & (g2000) & (!g2045)) + ((!g1030) & (g1160) & (!g1977) & (g1978) & (!g2000) & (!g2045)) + ((!g1030) & (g1160) & (!g1977) & (g1978) & (g2000) & (!g2045)) + ((!g1030) & (g1160) & (g1977) & (!g1978) & (!g2000) & (!g2045)) + ((!g1030) & (g1160) & (g1977) & (!g1978) & (!g2000) & (g2045)) + ((!g1030) & (g1160) & (g1977) & (!g1978) & (g2000) & (g2045)) + ((!g1030) & (g1160) & (g1977) & (g1978) & (!g2000) & (g2045)) + ((!g1030) & (g1160) & (g1977) & (g1978) & (g2000) & (g2045)) + ((g1030) & (!g1160) & (!g1977) & (!g1978) & (!g2000) & (!g2045)) + ((g1030) & (!g1160) & (!g1977) & (!g1978) & (g2000) & (!g2045)) + ((g1030) & (!g1160) & (!g1977) & (g1978) & (!g2000) & (!g2045)) + ((g1030) & (!g1160) & (g1977) & (!g1978) & (!g2000) & (g2045)) + ((g1030) & (!g1160) & (g1977) & (!g1978) & (g2000) & (g2045)) + ((g1030) & (!g1160) & (g1977) & (g1978) & (!g2000) & (g2045)) + ((g1030) & (!g1160) & (g1977) & (g1978) & (g2000) & (!g2045)) + ((g1030) & (!g1160) & (g1977) & (g1978) & (g2000) & (g2045)) + ((g1030) & (g1160) & (!g1977) & (!g1978) & (!g2000) & (!g2045)) + ((g1030) & (g1160) & (g1977) & (!g1978) & (!g2000) & (g2045)) + ((g1030) & (g1160) & (g1977) & (!g1978) & (g2000) & (!g2045)) + ((g1030) & (g1160) & (g1977) & (!g1978) & (g2000) & (g2045)) + ((g1030) & (g1160) & (g1977) & (g1978) & (!g2000) & (!g2045)) + ((g1030) & (g1160) & (g1977) & (g1978) & (!g2000) & (g2045)) + ((g1030) & (g1160) & (g1977) & (g1978) & (g2000) & (!g2045)) + ((g1030) & (g1160) & (g1977) & (g1978) & (g2000) & (g2045)));
	assign g2064 = (((!g1160) & (!g1978) & (g2000) & (!g2045)) + ((!g1160) & (g1978) & (!g2000) & (!g2045)) + ((!g1160) & (g1978) & (!g2000) & (g2045)) + ((!g1160) & (g1978) & (g2000) & (g2045)) + ((g1160) & (!g1978) & (!g2000) & (!g2045)) + ((g1160) & (g1978) & (!g2000) & (g2045)) + ((g1160) & (g1978) & (g2000) & (!g2045)) + ((g1160) & (g1978) & (g2000) & (g2045)));
	assign g2065 = (((!g1154) & (!g1295) & (!g1980) & (g1981) & (g1999) & (!g2045)) + ((!g1154) & (!g1295) & (g1980) & (!g1981) & (!g1999) & (!g2045)) + ((!g1154) & (!g1295) & (g1980) & (!g1981) & (!g1999) & (g2045)) + ((!g1154) & (!g1295) & (g1980) & (!g1981) & (g1999) & (!g2045)) + ((!g1154) & (!g1295) & (g1980) & (!g1981) & (g1999) & (g2045)) + ((!g1154) & (!g1295) & (g1980) & (g1981) & (!g1999) & (!g2045)) + ((!g1154) & (!g1295) & (g1980) & (g1981) & (!g1999) & (g2045)) + ((!g1154) & (!g1295) & (g1980) & (g1981) & (g1999) & (g2045)) + ((!g1154) & (g1295) & (!g1980) & (!g1981) & (g1999) & (!g2045)) + ((!g1154) & (g1295) & (!g1980) & (g1981) & (!g1999) & (!g2045)) + ((!g1154) & (g1295) & (!g1980) & (g1981) & (g1999) & (!g2045)) + ((!g1154) & (g1295) & (g1980) & (!g1981) & (!g1999) & (!g2045)) + ((!g1154) & (g1295) & (g1980) & (!g1981) & (!g1999) & (g2045)) + ((!g1154) & (g1295) & (g1980) & (!g1981) & (g1999) & (g2045)) + ((!g1154) & (g1295) & (g1980) & (g1981) & (!g1999) & (g2045)) + ((!g1154) & (g1295) & (g1980) & (g1981) & (g1999) & (g2045)) + ((g1154) & (!g1295) & (!g1980) & (!g1981) & (!g1999) & (!g2045)) + ((g1154) & (!g1295) & (!g1980) & (!g1981) & (g1999) & (!g2045)) + ((g1154) & (!g1295) & (!g1980) & (g1981) & (!g1999) & (!g2045)) + ((g1154) & (!g1295) & (g1980) & (!g1981) & (!g1999) & (g2045)) + ((g1154) & (!g1295) & (g1980) & (!g1981) & (g1999) & (g2045)) + ((g1154) & (!g1295) & (g1980) & (g1981) & (!g1999) & (g2045)) + ((g1154) & (!g1295) & (g1980) & (g1981) & (g1999) & (!g2045)) + ((g1154) & (!g1295) & (g1980) & (g1981) & (g1999) & (g2045)) + ((g1154) & (g1295) & (!g1980) & (!g1981) & (!g1999) & (!g2045)) + ((g1154) & (g1295) & (g1980) & (!g1981) & (!g1999) & (g2045)) + ((g1154) & (g1295) & (g1980) & (!g1981) & (g1999) & (!g2045)) + ((g1154) & (g1295) & (g1980) & (!g1981) & (g1999) & (g2045)) + ((g1154) & (g1295) & (g1980) & (g1981) & (!g1999) & (!g2045)) + ((g1154) & (g1295) & (g1980) & (g1981) & (!g1999) & (g2045)) + ((g1154) & (g1295) & (g1980) & (g1981) & (g1999) & (!g2045)) + ((g1154) & (g1295) & (g1980) & (g1981) & (g1999) & (g2045)));
	assign g2066 = (((!g1295) & (!g1981) & (g1999) & (!g2045)) + ((!g1295) & (g1981) & (!g1999) & (!g2045)) + ((!g1295) & (g1981) & (!g1999) & (g2045)) + ((!g1295) & (g1981) & (g1999) & (g2045)) + ((g1295) & (!g1981) & (!g1999) & (!g2045)) + ((g1295) & (g1981) & (!g1999) & (g2045)) + ((g1295) & (g1981) & (g1999) & (!g2045)) + ((g1295) & (g1981) & (g1999) & (g2045)));
	assign g2067 = (((!g1285) & (!g1437) & (!g1983) & (g1984) & (g1998) & (!g2045)) + ((!g1285) & (!g1437) & (g1983) & (!g1984) & (!g1998) & (!g2045)) + ((!g1285) & (!g1437) & (g1983) & (!g1984) & (!g1998) & (g2045)) + ((!g1285) & (!g1437) & (g1983) & (!g1984) & (g1998) & (!g2045)) + ((!g1285) & (!g1437) & (g1983) & (!g1984) & (g1998) & (g2045)) + ((!g1285) & (!g1437) & (g1983) & (g1984) & (!g1998) & (!g2045)) + ((!g1285) & (!g1437) & (g1983) & (g1984) & (!g1998) & (g2045)) + ((!g1285) & (!g1437) & (g1983) & (g1984) & (g1998) & (g2045)) + ((!g1285) & (g1437) & (!g1983) & (!g1984) & (g1998) & (!g2045)) + ((!g1285) & (g1437) & (!g1983) & (g1984) & (!g1998) & (!g2045)) + ((!g1285) & (g1437) & (!g1983) & (g1984) & (g1998) & (!g2045)) + ((!g1285) & (g1437) & (g1983) & (!g1984) & (!g1998) & (!g2045)) + ((!g1285) & (g1437) & (g1983) & (!g1984) & (!g1998) & (g2045)) + ((!g1285) & (g1437) & (g1983) & (!g1984) & (g1998) & (g2045)) + ((!g1285) & (g1437) & (g1983) & (g1984) & (!g1998) & (g2045)) + ((!g1285) & (g1437) & (g1983) & (g1984) & (g1998) & (g2045)) + ((g1285) & (!g1437) & (!g1983) & (!g1984) & (!g1998) & (!g2045)) + ((g1285) & (!g1437) & (!g1983) & (!g1984) & (g1998) & (!g2045)) + ((g1285) & (!g1437) & (!g1983) & (g1984) & (!g1998) & (!g2045)) + ((g1285) & (!g1437) & (g1983) & (!g1984) & (!g1998) & (g2045)) + ((g1285) & (!g1437) & (g1983) & (!g1984) & (g1998) & (g2045)) + ((g1285) & (!g1437) & (g1983) & (g1984) & (!g1998) & (g2045)) + ((g1285) & (!g1437) & (g1983) & (g1984) & (g1998) & (!g2045)) + ((g1285) & (!g1437) & (g1983) & (g1984) & (g1998) & (g2045)) + ((g1285) & (g1437) & (!g1983) & (!g1984) & (!g1998) & (!g2045)) + ((g1285) & (g1437) & (g1983) & (!g1984) & (!g1998) & (g2045)) + ((g1285) & (g1437) & (g1983) & (!g1984) & (g1998) & (!g2045)) + ((g1285) & (g1437) & (g1983) & (!g1984) & (g1998) & (g2045)) + ((g1285) & (g1437) & (g1983) & (g1984) & (!g1998) & (!g2045)) + ((g1285) & (g1437) & (g1983) & (g1984) & (!g1998) & (g2045)) + ((g1285) & (g1437) & (g1983) & (g1984) & (g1998) & (!g2045)) + ((g1285) & (g1437) & (g1983) & (g1984) & (g1998) & (g2045)));
	assign g2068 = (((!g1437) & (!g1984) & (g1998) & (!g2045)) + ((!g1437) & (g1984) & (!g1998) & (!g2045)) + ((!g1437) & (g1984) & (!g1998) & (g2045)) + ((!g1437) & (g1984) & (g1998) & (g2045)) + ((g1437) & (!g1984) & (!g1998) & (!g2045)) + ((g1437) & (g1984) & (!g1998) & (g2045)) + ((g1437) & (g1984) & (g1998) & (!g2045)) + ((g1437) & (g1984) & (g1998) & (g2045)));
	assign g2069 = (((!g1423) & (!g1586) & (!g1986) & (g1987) & (g1997) & (!g2045)) + ((!g1423) & (!g1586) & (g1986) & (!g1987) & (!g1997) & (!g2045)) + ((!g1423) & (!g1586) & (g1986) & (!g1987) & (!g1997) & (g2045)) + ((!g1423) & (!g1586) & (g1986) & (!g1987) & (g1997) & (!g2045)) + ((!g1423) & (!g1586) & (g1986) & (!g1987) & (g1997) & (g2045)) + ((!g1423) & (!g1586) & (g1986) & (g1987) & (!g1997) & (!g2045)) + ((!g1423) & (!g1586) & (g1986) & (g1987) & (!g1997) & (g2045)) + ((!g1423) & (!g1586) & (g1986) & (g1987) & (g1997) & (g2045)) + ((!g1423) & (g1586) & (!g1986) & (!g1987) & (g1997) & (!g2045)) + ((!g1423) & (g1586) & (!g1986) & (g1987) & (!g1997) & (!g2045)) + ((!g1423) & (g1586) & (!g1986) & (g1987) & (g1997) & (!g2045)) + ((!g1423) & (g1586) & (g1986) & (!g1987) & (!g1997) & (!g2045)) + ((!g1423) & (g1586) & (g1986) & (!g1987) & (!g1997) & (g2045)) + ((!g1423) & (g1586) & (g1986) & (!g1987) & (g1997) & (g2045)) + ((!g1423) & (g1586) & (g1986) & (g1987) & (!g1997) & (g2045)) + ((!g1423) & (g1586) & (g1986) & (g1987) & (g1997) & (g2045)) + ((g1423) & (!g1586) & (!g1986) & (!g1987) & (!g1997) & (!g2045)) + ((g1423) & (!g1586) & (!g1986) & (!g1987) & (g1997) & (!g2045)) + ((g1423) & (!g1586) & (!g1986) & (g1987) & (!g1997) & (!g2045)) + ((g1423) & (!g1586) & (g1986) & (!g1987) & (!g1997) & (g2045)) + ((g1423) & (!g1586) & (g1986) & (!g1987) & (g1997) & (g2045)) + ((g1423) & (!g1586) & (g1986) & (g1987) & (!g1997) & (g2045)) + ((g1423) & (!g1586) & (g1986) & (g1987) & (g1997) & (!g2045)) + ((g1423) & (!g1586) & (g1986) & (g1987) & (g1997) & (g2045)) + ((g1423) & (g1586) & (!g1986) & (!g1987) & (!g1997) & (!g2045)) + ((g1423) & (g1586) & (g1986) & (!g1987) & (!g1997) & (g2045)) + ((g1423) & (g1586) & (g1986) & (!g1987) & (g1997) & (!g2045)) + ((g1423) & (g1586) & (g1986) & (!g1987) & (g1997) & (g2045)) + ((g1423) & (g1586) & (g1986) & (g1987) & (!g1997) & (!g2045)) + ((g1423) & (g1586) & (g1986) & (g1987) & (!g1997) & (g2045)) + ((g1423) & (g1586) & (g1986) & (g1987) & (g1997) & (!g2045)) + ((g1423) & (g1586) & (g1986) & (g1987) & (g1997) & (g2045)));
	assign g2070 = (((!g1586) & (!g1987) & (g1997) & (!g2045)) + ((!g1586) & (g1987) & (!g1997) & (!g2045)) + ((!g1586) & (g1987) & (!g1997) & (g2045)) + ((!g1586) & (g1987) & (g1997) & (g2045)) + ((g1586) & (!g1987) & (!g1997) & (!g2045)) + ((g1586) & (g1987) & (!g1997) & (g2045)) + ((g1586) & (g1987) & (g1997) & (!g2045)) + ((g1586) & (g1987) & (g1997) & (g2045)));
	assign g2071 = (((!g1568) & (!g1742) & (!g1989) & (g1990) & (g1996) & (!g2045)) + ((!g1568) & (!g1742) & (g1989) & (!g1990) & (!g1996) & (!g2045)) + ((!g1568) & (!g1742) & (g1989) & (!g1990) & (!g1996) & (g2045)) + ((!g1568) & (!g1742) & (g1989) & (!g1990) & (g1996) & (!g2045)) + ((!g1568) & (!g1742) & (g1989) & (!g1990) & (g1996) & (g2045)) + ((!g1568) & (!g1742) & (g1989) & (g1990) & (!g1996) & (!g2045)) + ((!g1568) & (!g1742) & (g1989) & (g1990) & (!g1996) & (g2045)) + ((!g1568) & (!g1742) & (g1989) & (g1990) & (g1996) & (g2045)) + ((!g1568) & (g1742) & (!g1989) & (!g1990) & (g1996) & (!g2045)) + ((!g1568) & (g1742) & (!g1989) & (g1990) & (!g1996) & (!g2045)) + ((!g1568) & (g1742) & (!g1989) & (g1990) & (g1996) & (!g2045)) + ((!g1568) & (g1742) & (g1989) & (!g1990) & (!g1996) & (!g2045)) + ((!g1568) & (g1742) & (g1989) & (!g1990) & (!g1996) & (g2045)) + ((!g1568) & (g1742) & (g1989) & (!g1990) & (g1996) & (g2045)) + ((!g1568) & (g1742) & (g1989) & (g1990) & (!g1996) & (g2045)) + ((!g1568) & (g1742) & (g1989) & (g1990) & (g1996) & (g2045)) + ((g1568) & (!g1742) & (!g1989) & (!g1990) & (!g1996) & (!g2045)) + ((g1568) & (!g1742) & (!g1989) & (!g1990) & (g1996) & (!g2045)) + ((g1568) & (!g1742) & (!g1989) & (g1990) & (!g1996) & (!g2045)) + ((g1568) & (!g1742) & (g1989) & (!g1990) & (!g1996) & (g2045)) + ((g1568) & (!g1742) & (g1989) & (!g1990) & (g1996) & (g2045)) + ((g1568) & (!g1742) & (g1989) & (g1990) & (!g1996) & (g2045)) + ((g1568) & (!g1742) & (g1989) & (g1990) & (g1996) & (!g2045)) + ((g1568) & (!g1742) & (g1989) & (g1990) & (g1996) & (g2045)) + ((g1568) & (g1742) & (!g1989) & (!g1990) & (!g1996) & (!g2045)) + ((g1568) & (g1742) & (g1989) & (!g1990) & (!g1996) & (g2045)) + ((g1568) & (g1742) & (g1989) & (!g1990) & (g1996) & (!g2045)) + ((g1568) & (g1742) & (g1989) & (!g1990) & (g1996) & (g2045)) + ((g1568) & (g1742) & (g1989) & (g1990) & (!g1996) & (!g2045)) + ((g1568) & (g1742) & (g1989) & (g1990) & (!g1996) & (g2045)) + ((g1568) & (g1742) & (g1989) & (g1990) & (g1996) & (!g2045)) + ((g1568) & (g1742) & (g1989) & (g1990) & (g1996) & (g2045)));
	assign g2072 = (((!g1742) & (!g1990) & (g1996) & (!g2045)) + ((!g1742) & (g1990) & (!g1996) & (!g2045)) + ((!g1742) & (g1990) & (!g1996) & (g2045)) + ((!g1742) & (g1990) & (g1996) & (g2045)) + ((g1742) & (!g1990) & (!g1996) & (!g2045)) + ((g1742) & (g1990) & (!g1996) & (g2045)) + ((g1742) & (g1990) & (g1996) & (!g2045)) + ((g1742) & (g1990) & (g1996) & (g2045)));
	assign g2073 = (((!g1720) & (!g1905) & (!g1992) & (g1993) & (g1995) & (!g2045)) + ((!g1720) & (!g1905) & (g1992) & (!g1993) & (!g1995) & (!g2045)) + ((!g1720) & (!g1905) & (g1992) & (!g1993) & (!g1995) & (g2045)) + ((!g1720) & (!g1905) & (g1992) & (!g1993) & (g1995) & (!g2045)) + ((!g1720) & (!g1905) & (g1992) & (!g1993) & (g1995) & (g2045)) + ((!g1720) & (!g1905) & (g1992) & (g1993) & (!g1995) & (!g2045)) + ((!g1720) & (!g1905) & (g1992) & (g1993) & (!g1995) & (g2045)) + ((!g1720) & (!g1905) & (g1992) & (g1993) & (g1995) & (g2045)) + ((!g1720) & (g1905) & (!g1992) & (!g1993) & (g1995) & (!g2045)) + ((!g1720) & (g1905) & (!g1992) & (g1993) & (!g1995) & (!g2045)) + ((!g1720) & (g1905) & (!g1992) & (g1993) & (g1995) & (!g2045)) + ((!g1720) & (g1905) & (g1992) & (!g1993) & (!g1995) & (!g2045)) + ((!g1720) & (g1905) & (g1992) & (!g1993) & (!g1995) & (g2045)) + ((!g1720) & (g1905) & (g1992) & (!g1993) & (g1995) & (g2045)) + ((!g1720) & (g1905) & (g1992) & (g1993) & (!g1995) & (g2045)) + ((!g1720) & (g1905) & (g1992) & (g1993) & (g1995) & (g2045)) + ((g1720) & (!g1905) & (!g1992) & (!g1993) & (!g1995) & (!g2045)) + ((g1720) & (!g1905) & (!g1992) & (!g1993) & (g1995) & (!g2045)) + ((g1720) & (!g1905) & (!g1992) & (g1993) & (!g1995) & (!g2045)) + ((g1720) & (!g1905) & (g1992) & (!g1993) & (!g1995) & (g2045)) + ((g1720) & (!g1905) & (g1992) & (!g1993) & (g1995) & (g2045)) + ((g1720) & (!g1905) & (g1992) & (g1993) & (!g1995) & (g2045)) + ((g1720) & (!g1905) & (g1992) & (g1993) & (g1995) & (!g2045)) + ((g1720) & (!g1905) & (g1992) & (g1993) & (g1995) & (g2045)) + ((g1720) & (g1905) & (!g1992) & (!g1993) & (!g1995) & (!g2045)) + ((g1720) & (g1905) & (g1992) & (!g1993) & (!g1995) & (g2045)) + ((g1720) & (g1905) & (g1992) & (!g1993) & (g1995) & (!g2045)) + ((g1720) & (g1905) & (g1992) & (!g1993) & (g1995) & (g2045)) + ((g1720) & (g1905) & (g1992) & (g1993) & (!g1995) & (!g2045)) + ((g1720) & (g1905) & (g1992) & (g1993) & (!g1995) & (g2045)) + ((g1720) & (g1905) & (g1992) & (g1993) & (g1995) & (!g2045)) + ((g1720) & (g1905) & (g1992) & (g1993) & (g1995) & (g2045)));
	assign g2074 = (((!g1905) & (!g1993) & (g1995) & (!g2045)) + ((!g1905) & (g1993) & (!g1995) & (!g2045)) + ((!g1905) & (g1993) & (!g1995) & (g2045)) + ((!g1905) & (g1993) & (g1995) & (g2045)) + ((g1905) & (!g1993) & (!g1995) & (!g2045)) + ((g1905) & (g1993) & (!g1995) & (g2045)) + ((g1905) & (g1993) & (g1995) & (!g2045)) + ((g1905) & (g1993) & (g1995) & (g2045)));
	assign g2075 = (((!g1923) & (g1950)));
	assign g2076 = (((!g1879) & (!ax34x) & (!ax35x) & (!g2075) & (!g1994) & (g2045)) + ((!g1879) & (!ax34x) & (!ax35x) & (!g2075) & (g1994) & (!g2045)) + ((!g1879) & (!ax34x) & (!ax35x) & (!g2075) & (g1994) & (g2045)) + ((!g1879) & (!ax34x) & (!ax35x) & (g2075) & (!g1994) & (!g2045)) + ((!g1879) & (!ax34x) & (ax35x) & (!g2075) & (!g1994) & (!g2045)) + ((!g1879) & (!ax34x) & (ax35x) & (g2075) & (!g1994) & (g2045)) + ((!g1879) & (!ax34x) & (ax35x) & (g2075) & (g1994) & (!g2045)) + ((!g1879) & (!ax34x) & (ax35x) & (g2075) & (g1994) & (g2045)) + ((!g1879) & (ax34x) & (!ax35x) & (g2075) & (!g1994) & (!g2045)) + ((!g1879) & (ax34x) & (!ax35x) & (g2075) & (g1994) & (!g2045)) + ((!g1879) & (ax34x) & (ax35x) & (!g2075) & (!g1994) & (!g2045)) + ((!g1879) & (ax34x) & (ax35x) & (!g2075) & (!g1994) & (g2045)) + ((!g1879) & (ax34x) & (ax35x) & (!g2075) & (g1994) & (!g2045)) + ((!g1879) & (ax34x) & (ax35x) & (!g2075) & (g1994) & (g2045)) + ((!g1879) & (ax34x) & (ax35x) & (g2075) & (!g1994) & (g2045)) + ((!g1879) & (ax34x) & (ax35x) & (g2075) & (g1994) & (g2045)) + ((g1879) & (!ax34x) & (!ax35x) & (!g2075) & (!g1994) & (!g2045)) + ((g1879) & (!ax34x) & (!ax35x) & (!g2075) & (!g1994) & (g2045)) + ((g1879) & (!ax34x) & (!ax35x) & (!g2075) & (g1994) & (g2045)) + ((g1879) & (!ax34x) & (!ax35x) & (g2075) & (g1994) & (!g2045)) + ((g1879) & (!ax34x) & (ax35x) & (!g2075) & (g1994) & (!g2045)) + ((g1879) & (!ax34x) & (ax35x) & (g2075) & (!g1994) & (!g2045)) + ((g1879) & (!ax34x) & (ax35x) & (g2075) & (!g1994) & (g2045)) + ((g1879) & (!ax34x) & (ax35x) & (g2075) & (g1994) & (g2045)) + ((g1879) & (ax34x) & (!ax35x) & (!g2075) & (!g1994) & (!g2045)) + ((g1879) & (ax34x) & (!ax35x) & (!g2075) & (g1994) & (!g2045)) + ((g1879) & (ax34x) & (ax35x) & (!g2075) & (!g1994) & (g2045)) + ((g1879) & (ax34x) & (ax35x) & (!g2075) & (g1994) & (g2045)) + ((g1879) & (ax34x) & (ax35x) & (g2075) & (!g1994) & (!g2045)) + ((g1879) & (ax34x) & (ax35x) & (g2075) & (!g1994) & (g2045)) + ((g1879) & (ax34x) & (ax35x) & (g2075) & (g1994) & (!g2045)) + ((g1879) & (ax34x) & (ax35x) & (g2075) & (g1994) & (g2045)));
	assign g2077 = (((!ax34x) & (!g2075) & (!g1994) & (g2045)) + ((!ax34x) & (!g2075) & (g1994) & (!g2045)) + ((!ax34x) & (!g2075) & (g1994) & (g2045)) + ((!ax34x) & (g2075) & (g1994) & (!g2045)) + ((ax34x) & (!g2075) & (!g1994) & (!g2045)) + ((ax34x) & (g2075) & (!g1994) & (!g2045)) + ((ax34x) & (g2075) & (!g1994) & (g2045)) + ((ax34x) & (g2075) & (g1994) & (g2045)));
	assign g2078 = (((!ax30x) & (!ax31x)));
	assign g2079 = (((!g2075) & (!ax32x) & (!ax33x) & (!g2045) & (!g2078)) + ((!g2075) & (!ax32x) & (ax33x) & (g2045) & (!g2078)) + ((!g2075) & (ax32x) & (ax33x) & (g2045) & (!g2078)) + ((!g2075) & (ax32x) & (ax33x) & (g2045) & (g2078)) + ((g2075) & (!ax32x) & (!ax33x) & (!g2045) & (!g2078)) + ((g2075) & (!ax32x) & (!ax33x) & (!g2045) & (g2078)) + ((g2075) & (!ax32x) & (!ax33x) & (g2045) & (!g2078)) + ((g2075) & (!ax32x) & (ax33x) & (!g2045) & (!g2078)) + ((g2075) & (!ax32x) & (ax33x) & (g2045) & (!g2078)) + ((g2075) & (!ax32x) & (ax33x) & (g2045) & (g2078)) + ((g2075) & (ax32x) & (!ax33x) & (g2045) & (!g2078)) + ((g2075) & (ax32x) & (!ax33x) & (g2045) & (g2078)) + ((g2075) & (ax32x) & (ax33x) & (!g2045) & (!g2078)) + ((g2075) & (ax32x) & (ax33x) & (!g2045) & (g2078)) + ((g2075) & (ax32x) & (ax33x) & (g2045) & (!g2078)) + ((g2075) & (ax32x) & (ax33x) & (g2045) & (g2078)));
	assign g2080 = (((!g1905) & (!g1879) & (g2076) & (g2077) & (g2079)) + ((!g1905) & (g1879) & (g2076) & (!g2077) & (g2079)) + ((!g1905) & (g1879) & (g2076) & (g2077) & (!g2079)) + ((!g1905) & (g1879) & (g2076) & (g2077) & (g2079)) + ((g1905) & (!g1879) & (!g2076) & (g2077) & (g2079)) + ((g1905) & (!g1879) & (g2076) & (!g2077) & (!g2079)) + ((g1905) & (!g1879) & (g2076) & (!g2077) & (g2079)) + ((g1905) & (!g1879) & (g2076) & (g2077) & (!g2079)) + ((g1905) & (!g1879) & (g2076) & (g2077) & (g2079)) + ((g1905) & (g1879) & (!g2076) & (!g2077) & (g2079)) + ((g1905) & (g1879) & (!g2076) & (g2077) & (!g2079)) + ((g1905) & (g1879) & (!g2076) & (g2077) & (g2079)) + ((g1905) & (g1879) & (g2076) & (!g2077) & (!g2079)) + ((g1905) & (g1879) & (g2076) & (!g2077) & (g2079)) + ((g1905) & (g1879) & (g2076) & (g2077) & (!g2079)) + ((g1905) & (g1879) & (g2076) & (g2077) & (g2079)));
	assign g2081 = (((!g1742) & (!g1720) & (g2073) & (g2074) & (g2080)) + ((!g1742) & (g1720) & (g2073) & (!g2074) & (g2080)) + ((!g1742) & (g1720) & (g2073) & (g2074) & (!g2080)) + ((!g1742) & (g1720) & (g2073) & (g2074) & (g2080)) + ((g1742) & (!g1720) & (!g2073) & (g2074) & (g2080)) + ((g1742) & (!g1720) & (g2073) & (!g2074) & (!g2080)) + ((g1742) & (!g1720) & (g2073) & (!g2074) & (g2080)) + ((g1742) & (!g1720) & (g2073) & (g2074) & (!g2080)) + ((g1742) & (!g1720) & (g2073) & (g2074) & (g2080)) + ((g1742) & (g1720) & (!g2073) & (!g2074) & (g2080)) + ((g1742) & (g1720) & (!g2073) & (g2074) & (!g2080)) + ((g1742) & (g1720) & (!g2073) & (g2074) & (g2080)) + ((g1742) & (g1720) & (g2073) & (!g2074) & (!g2080)) + ((g1742) & (g1720) & (g2073) & (!g2074) & (g2080)) + ((g1742) & (g1720) & (g2073) & (g2074) & (!g2080)) + ((g1742) & (g1720) & (g2073) & (g2074) & (g2080)));
	assign g2082 = (((!g1586) & (!g1568) & (g2071) & (g2072) & (g2081)) + ((!g1586) & (g1568) & (g2071) & (!g2072) & (g2081)) + ((!g1586) & (g1568) & (g2071) & (g2072) & (!g2081)) + ((!g1586) & (g1568) & (g2071) & (g2072) & (g2081)) + ((g1586) & (!g1568) & (!g2071) & (g2072) & (g2081)) + ((g1586) & (!g1568) & (g2071) & (!g2072) & (!g2081)) + ((g1586) & (!g1568) & (g2071) & (!g2072) & (g2081)) + ((g1586) & (!g1568) & (g2071) & (g2072) & (!g2081)) + ((g1586) & (!g1568) & (g2071) & (g2072) & (g2081)) + ((g1586) & (g1568) & (!g2071) & (!g2072) & (g2081)) + ((g1586) & (g1568) & (!g2071) & (g2072) & (!g2081)) + ((g1586) & (g1568) & (!g2071) & (g2072) & (g2081)) + ((g1586) & (g1568) & (g2071) & (!g2072) & (!g2081)) + ((g1586) & (g1568) & (g2071) & (!g2072) & (g2081)) + ((g1586) & (g1568) & (g2071) & (g2072) & (!g2081)) + ((g1586) & (g1568) & (g2071) & (g2072) & (g2081)));
	assign g2083 = (((!g1437) & (!g1423) & (g2069) & (g2070) & (g2082)) + ((!g1437) & (g1423) & (g2069) & (!g2070) & (g2082)) + ((!g1437) & (g1423) & (g2069) & (g2070) & (!g2082)) + ((!g1437) & (g1423) & (g2069) & (g2070) & (g2082)) + ((g1437) & (!g1423) & (!g2069) & (g2070) & (g2082)) + ((g1437) & (!g1423) & (g2069) & (!g2070) & (!g2082)) + ((g1437) & (!g1423) & (g2069) & (!g2070) & (g2082)) + ((g1437) & (!g1423) & (g2069) & (g2070) & (!g2082)) + ((g1437) & (!g1423) & (g2069) & (g2070) & (g2082)) + ((g1437) & (g1423) & (!g2069) & (!g2070) & (g2082)) + ((g1437) & (g1423) & (!g2069) & (g2070) & (!g2082)) + ((g1437) & (g1423) & (!g2069) & (g2070) & (g2082)) + ((g1437) & (g1423) & (g2069) & (!g2070) & (!g2082)) + ((g1437) & (g1423) & (g2069) & (!g2070) & (g2082)) + ((g1437) & (g1423) & (g2069) & (g2070) & (!g2082)) + ((g1437) & (g1423) & (g2069) & (g2070) & (g2082)));
	assign g2084 = (((!g1295) & (!g1285) & (g2067) & (g2068) & (g2083)) + ((!g1295) & (g1285) & (g2067) & (!g2068) & (g2083)) + ((!g1295) & (g1285) & (g2067) & (g2068) & (!g2083)) + ((!g1295) & (g1285) & (g2067) & (g2068) & (g2083)) + ((g1295) & (!g1285) & (!g2067) & (g2068) & (g2083)) + ((g1295) & (!g1285) & (g2067) & (!g2068) & (!g2083)) + ((g1295) & (!g1285) & (g2067) & (!g2068) & (g2083)) + ((g1295) & (!g1285) & (g2067) & (g2068) & (!g2083)) + ((g1295) & (!g1285) & (g2067) & (g2068) & (g2083)) + ((g1295) & (g1285) & (!g2067) & (!g2068) & (g2083)) + ((g1295) & (g1285) & (!g2067) & (g2068) & (!g2083)) + ((g1295) & (g1285) & (!g2067) & (g2068) & (g2083)) + ((g1295) & (g1285) & (g2067) & (!g2068) & (!g2083)) + ((g1295) & (g1285) & (g2067) & (!g2068) & (g2083)) + ((g1295) & (g1285) & (g2067) & (g2068) & (!g2083)) + ((g1295) & (g1285) & (g2067) & (g2068) & (g2083)));
	assign g2085 = (((!g1160) & (!g1154) & (g2065) & (g2066) & (g2084)) + ((!g1160) & (g1154) & (g2065) & (!g2066) & (g2084)) + ((!g1160) & (g1154) & (g2065) & (g2066) & (!g2084)) + ((!g1160) & (g1154) & (g2065) & (g2066) & (g2084)) + ((g1160) & (!g1154) & (!g2065) & (g2066) & (g2084)) + ((g1160) & (!g1154) & (g2065) & (!g2066) & (!g2084)) + ((g1160) & (!g1154) & (g2065) & (!g2066) & (g2084)) + ((g1160) & (!g1154) & (g2065) & (g2066) & (!g2084)) + ((g1160) & (!g1154) & (g2065) & (g2066) & (g2084)) + ((g1160) & (g1154) & (!g2065) & (!g2066) & (g2084)) + ((g1160) & (g1154) & (!g2065) & (g2066) & (!g2084)) + ((g1160) & (g1154) & (!g2065) & (g2066) & (g2084)) + ((g1160) & (g1154) & (g2065) & (!g2066) & (!g2084)) + ((g1160) & (g1154) & (g2065) & (!g2066) & (g2084)) + ((g1160) & (g1154) & (g2065) & (g2066) & (!g2084)) + ((g1160) & (g1154) & (g2065) & (g2066) & (g2084)));
	assign g2086 = (((!g1032) & (!g1030) & (g2063) & (g2064) & (g2085)) + ((!g1032) & (g1030) & (g2063) & (!g2064) & (g2085)) + ((!g1032) & (g1030) & (g2063) & (g2064) & (!g2085)) + ((!g1032) & (g1030) & (g2063) & (g2064) & (g2085)) + ((g1032) & (!g1030) & (!g2063) & (g2064) & (g2085)) + ((g1032) & (!g1030) & (g2063) & (!g2064) & (!g2085)) + ((g1032) & (!g1030) & (g2063) & (!g2064) & (g2085)) + ((g1032) & (!g1030) & (g2063) & (g2064) & (!g2085)) + ((g1032) & (!g1030) & (g2063) & (g2064) & (g2085)) + ((g1032) & (g1030) & (!g2063) & (!g2064) & (g2085)) + ((g1032) & (g1030) & (!g2063) & (g2064) & (!g2085)) + ((g1032) & (g1030) & (!g2063) & (g2064) & (g2085)) + ((g1032) & (g1030) & (g2063) & (!g2064) & (!g2085)) + ((g1032) & (g1030) & (g2063) & (!g2064) & (g2085)) + ((g1032) & (g1030) & (g2063) & (g2064) & (!g2085)) + ((g1032) & (g1030) & (g2063) & (g2064) & (g2085)));
	assign g2087 = (((!g851) & (!g914) & (g2061) & (g2062) & (g2086)) + ((!g851) & (g914) & (g2061) & (!g2062) & (g2086)) + ((!g851) & (g914) & (g2061) & (g2062) & (!g2086)) + ((!g851) & (g914) & (g2061) & (g2062) & (g2086)) + ((g851) & (!g914) & (!g2061) & (g2062) & (g2086)) + ((g851) & (!g914) & (g2061) & (!g2062) & (!g2086)) + ((g851) & (!g914) & (g2061) & (!g2062) & (g2086)) + ((g851) & (!g914) & (g2061) & (g2062) & (!g2086)) + ((g851) & (!g914) & (g2061) & (g2062) & (g2086)) + ((g851) & (g914) & (!g2061) & (!g2062) & (g2086)) + ((g851) & (g914) & (!g2061) & (g2062) & (!g2086)) + ((g851) & (g914) & (!g2061) & (g2062) & (g2086)) + ((g851) & (g914) & (g2061) & (!g2062) & (!g2086)) + ((g851) & (g914) & (g2061) & (!g2062) & (g2086)) + ((g851) & (g914) & (g2061) & (g2062) & (!g2086)) + ((g851) & (g914) & (g2061) & (g2062) & (g2086)));
	assign g2088 = (((!g744) & (!g803) & (g2059) & (g2060) & (g2087)) + ((!g744) & (g803) & (g2059) & (!g2060) & (g2087)) + ((!g744) & (g803) & (g2059) & (g2060) & (!g2087)) + ((!g744) & (g803) & (g2059) & (g2060) & (g2087)) + ((g744) & (!g803) & (!g2059) & (g2060) & (g2087)) + ((g744) & (!g803) & (g2059) & (!g2060) & (!g2087)) + ((g744) & (!g803) & (g2059) & (!g2060) & (g2087)) + ((g744) & (!g803) & (g2059) & (g2060) & (!g2087)) + ((g744) & (!g803) & (g2059) & (g2060) & (g2087)) + ((g744) & (g803) & (!g2059) & (!g2060) & (g2087)) + ((g744) & (g803) & (!g2059) & (g2060) & (!g2087)) + ((g744) & (g803) & (!g2059) & (g2060) & (g2087)) + ((g744) & (g803) & (g2059) & (!g2060) & (!g2087)) + ((g744) & (g803) & (g2059) & (!g2060) & (g2087)) + ((g744) & (g803) & (g2059) & (g2060) & (!g2087)) + ((g744) & (g803) & (g2059) & (g2060) & (g2087)));
	assign g2089 = (((!g645) & (!g700) & (g2057) & (g2058) & (g2088)) + ((!g645) & (g700) & (g2057) & (!g2058) & (g2088)) + ((!g645) & (g700) & (g2057) & (g2058) & (!g2088)) + ((!g645) & (g700) & (g2057) & (g2058) & (g2088)) + ((g645) & (!g700) & (!g2057) & (g2058) & (g2088)) + ((g645) & (!g700) & (g2057) & (!g2058) & (!g2088)) + ((g645) & (!g700) & (g2057) & (!g2058) & (g2088)) + ((g645) & (!g700) & (g2057) & (g2058) & (!g2088)) + ((g645) & (!g700) & (g2057) & (g2058) & (g2088)) + ((g645) & (g700) & (!g2057) & (!g2058) & (g2088)) + ((g645) & (g700) & (!g2057) & (g2058) & (!g2088)) + ((g645) & (g700) & (!g2057) & (g2058) & (g2088)) + ((g645) & (g700) & (g2057) & (!g2058) & (!g2088)) + ((g645) & (g700) & (g2057) & (!g2058) & (g2088)) + ((g645) & (g700) & (g2057) & (g2058) & (!g2088)) + ((g645) & (g700) & (g2057) & (g2058) & (g2088)));
	assign g2090 = (((!g553) & (!g604) & (g2055) & (g2056) & (g2089)) + ((!g553) & (g604) & (g2055) & (!g2056) & (g2089)) + ((!g553) & (g604) & (g2055) & (g2056) & (!g2089)) + ((!g553) & (g604) & (g2055) & (g2056) & (g2089)) + ((g553) & (!g604) & (!g2055) & (g2056) & (g2089)) + ((g553) & (!g604) & (g2055) & (!g2056) & (!g2089)) + ((g553) & (!g604) & (g2055) & (!g2056) & (g2089)) + ((g553) & (!g604) & (g2055) & (g2056) & (!g2089)) + ((g553) & (!g604) & (g2055) & (g2056) & (g2089)) + ((g553) & (g604) & (!g2055) & (!g2056) & (g2089)) + ((g553) & (g604) & (!g2055) & (g2056) & (!g2089)) + ((g553) & (g604) & (!g2055) & (g2056) & (g2089)) + ((g553) & (g604) & (g2055) & (!g2056) & (!g2089)) + ((g553) & (g604) & (g2055) & (!g2056) & (g2089)) + ((g553) & (g604) & (g2055) & (g2056) & (!g2089)) + ((g553) & (g604) & (g2055) & (g2056) & (g2089)));
	assign g2091 = (((!g468) & (!g515) & (g2053) & (g2054) & (g2090)) + ((!g468) & (g515) & (g2053) & (!g2054) & (g2090)) + ((!g468) & (g515) & (g2053) & (g2054) & (!g2090)) + ((!g468) & (g515) & (g2053) & (g2054) & (g2090)) + ((g468) & (!g515) & (!g2053) & (g2054) & (g2090)) + ((g468) & (!g515) & (g2053) & (!g2054) & (!g2090)) + ((g468) & (!g515) & (g2053) & (!g2054) & (g2090)) + ((g468) & (!g515) & (g2053) & (g2054) & (!g2090)) + ((g468) & (!g515) & (g2053) & (g2054) & (g2090)) + ((g468) & (g515) & (!g2053) & (!g2054) & (g2090)) + ((g468) & (g515) & (!g2053) & (g2054) & (!g2090)) + ((g468) & (g515) & (!g2053) & (g2054) & (g2090)) + ((g468) & (g515) & (g2053) & (!g2054) & (!g2090)) + ((g468) & (g515) & (g2053) & (!g2054) & (g2090)) + ((g468) & (g515) & (g2053) & (g2054) & (!g2090)) + ((g468) & (g515) & (g2053) & (g2054) & (g2090)));
	assign g2092 = (((!g390) & (!g433) & (g2051) & (g2052) & (g2091)) + ((!g390) & (g433) & (g2051) & (!g2052) & (g2091)) + ((!g390) & (g433) & (g2051) & (g2052) & (!g2091)) + ((!g390) & (g433) & (g2051) & (g2052) & (g2091)) + ((g390) & (!g433) & (!g2051) & (g2052) & (g2091)) + ((g390) & (!g433) & (g2051) & (!g2052) & (!g2091)) + ((g390) & (!g433) & (g2051) & (!g2052) & (g2091)) + ((g390) & (!g433) & (g2051) & (g2052) & (!g2091)) + ((g390) & (!g433) & (g2051) & (g2052) & (g2091)) + ((g390) & (g433) & (!g2051) & (!g2052) & (g2091)) + ((g390) & (g433) & (!g2051) & (g2052) & (!g2091)) + ((g390) & (g433) & (!g2051) & (g2052) & (g2091)) + ((g390) & (g433) & (g2051) & (!g2052) & (!g2091)) + ((g390) & (g433) & (g2051) & (!g2052) & (g2091)) + ((g390) & (g433) & (g2051) & (g2052) & (!g2091)) + ((g390) & (g433) & (g2051) & (g2052) & (g2091)));
	assign g2093 = (((!g319) & (!g358) & (g2049) & (g2050) & (g2092)) + ((!g319) & (g358) & (g2049) & (!g2050) & (g2092)) + ((!g319) & (g358) & (g2049) & (g2050) & (!g2092)) + ((!g319) & (g358) & (g2049) & (g2050) & (g2092)) + ((g319) & (!g358) & (!g2049) & (g2050) & (g2092)) + ((g319) & (!g358) & (g2049) & (!g2050) & (!g2092)) + ((g319) & (!g358) & (g2049) & (!g2050) & (g2092)) + ((g319) & (!g358) & (g2049) & (g2050) & (!g2092)) + ((g319) & (!g358) & (g2049) & (g2050) & (g2092)) + ((g319) & (g358) & (!g2049) & (!g2050) & (g2092)) + ((g319) & (g358) & (!g2049) & (g2050) & (!g2092)) + ((g319) & (g358) & (!g2049) & (g2050) & (g2092)) + ((g319) & (g358) & (g2049) & (!g2050) & (!g2092)) + ((g319) & (g358) & (g2049) & (!g2050) & (g2092)) + ((g319) & (g358) & (g2049) & (g2050) & (!g2092)) + ((g319) & (g358) & (g2049) & (g2050) & (g2092)));
	assign g2094 = (((!g255) & (!g290) & (g2047) & (g2048) & (g2093)) + ((!g255) & (g290) & (g2047) & (!g2048) & (g2093)) + ((!g255) & (g290) & (g2047) & (g2048) & (!g2093)) + ((!g255) & (g290) & (g2047) & (g2048) & (g2093)) + ((g255) & (!g290) & (!g2047) & (g2048) & (g2093)) + ((g255) & (!g290) & (g2047) & (!g2048) & (!g2093)) + ((g255) & (!g290) & (g2047) & (!g2048) & (g2093)) + ((g255) & (!g290) & (g2047) & (g2048) & (!g2093)) + ((g255) & (!g290) & (g2047) & (g2048) & (g2093)) + ((g255) & (g290) & (!g2047) & (!g2048) & (g2093)) + ((g255) & (g290) & (!g2047) & (g2048) & (!g2093)) + ((g255) & (g290) & (!g2047) & (g2048) & (g2093)) + ((g255) & (g290) & (g2047) & (!g2048) & (!g2093)) + ((g255) & (g290) & (g2047) & (!g2048) & (g2093)) + ((g255) & (g290) & (g2047) & (g2048) & (!g2093)) + ((g255) & (g290) & (g2047) & (g2048) & (g2093)));
	assign g2095 = (((g1) & (!g2010) & (g2041) & (g2044)) + ((g1) & (g2010) & (!g2041) & (!g2044)) + ((g1) & (g2010) & (!g2041) & (g2044)));
	assign g2096 = (((!g4) & (!g2) & (!g2011) & (!g2038) & (!g2040) & (!g2045)) + ((!g4) & (!g2) & (!g2011) & (!g2038) & (g2040) & (g2045)) + ((!g4) & (!g2) & (!g2011) & (g2038) & (!g2040) & (!g2045)) + ((!g4) & (!g2) & (!g2011) & (g2038) & (g2040) & (g2045)) + ((!g4) & (!g2) & (g2011) & (!g2038) & (!g2040) & (!g2045)) + ((!g4) & (!g2) & (g2011) & (!g2038) & (g2040) & (g2045)) + ((!g4) & (!g2) & (g2011) & (g2038) & (g2040) & (!g2045)) + ((!g4) & (!g2) & (g2011) & (g2038) & (g2040) & (g2045)) + ((!g4) & (g2) & (!g2011) & (!g2038) & (!g2040) & (!g2045)) + ((!g4) & (g2) & (!g2011) & (!g2038) & (g2040) & (g2045)) + ((!g4) & (g2) & (!g2011) & (g2038) & (g2040) & (!g2045)) + ((!g4) & (g2) & (!g2011) & (g2038) & (g2040) & (g2045)) + ((!g4) & (g2) & (g2011) & (!g2038) & (g2040) & (!g2045)) + ((!g4) & (g2) & (g2011) & (!g2038) & (g2040) & (g2045)) + ((!g4) & (g2) & (g2011) & (g2038) & (g2040) & (!g2045)) + ((!g4) & (g2) & (g2011) & (g2038) & (g2040) & (g2045)) + ((g4) & (!g2) & (!g2011) & (!g2038) & (g2040) & (!g2045)) + ((g4) & (!g2) & (!g2011) & (!g2038) & (g2040) & (g2045)) + ((g4) & (!g2) & (!g2011) & (g2038) & (g2040) & (!g2045)) + ((g4) & (!g2) & (!g2011) & (g2038) & (g2040) & (g2045)) + ((g4) & (!g2) & (g2011) & (!g2038) & (g2040) & (!g2045)) + ((g4) & (!g2) & (g2011) & (!g2038) & (g2040) & (g2045)) + ((g4) & (!g2) & (g2011) & (g2038) & (!g2040) & (!g2045)) + ((g4) & (!g2) & (g2011) & (g2038) & (g2040) & (g2045)) + ((g4) & (g2) & (!g2011) & (!g2038) & (g2040) & (!g2045)) + ((g4) & (g2) & (!g2011) & (!g2038) & (g2040) & (g2045)) + ((g4) & (g2) & (!g2011) & (g2038) & (!g2040) & (!g2045)) + ((g4) & (g2) & (!g2011) & (g2038) & (g2040) & (g2045)) + ((g4) & (g2) & (g2011) & (!g2038) & (!g2040) & (!g2045)) + ((g4) & (g2) & (g2011) & (!g2038) & (g2040) & (g2045)) + ((g4) & (g2) & (g2011) & (g2038) & (!g2040) & (!g2045)) + ((g4) & (g2) & (g2011) & (g2038) & (g2040) & (g2045)));
	assign g2097 = (((!g8) & (!g18) & (!g2013) & (g2014) & (g2037) & (!g2045)) + ((!g8) & (!g18) & (g2013) & (!g2014) & (!g2037) & (!g2045)) + ((!g8) & (!g18) & (g2013) & (!g2014) & (!g2037) & (g2045)) + ((!g8) & (!g18) & (g2013) & (!g2014) & (g2037) & (!g2045)) + ((!g8) & (!g18) & (g2013) & (!g2014) & (g2037) & (g2045)) + ((!g8) & (!g18) & (g2013) & (g2014) & (!g2037) & (!g2045)) + ((!g8) & (!g18) & (g2013) & (g2014) & (!g2037) & (g2045)) + ((!g8) & (!g18) & (g2013) & (g2014) & (g2037) & (g2045)) + ((!g8) & (g18) & (!g2013) & (!g2014) & (g2037) & (!g2045)) + ((!g8) & (g18) & (!g2013) & (g2014) & (!g2037) & (!g2045)) + ((!g8) & (g18) & (!g2013) & (g2014) & (g2037) & (!g2045)) + ((!g8) & (g18) & (g2013) & (!g2014) & (!g2037) & (!g2045)) + ((!g8) & (g18) & (g2013) & (!g2014) & (!g2037) & (g2045)) + ((!g8) & (g18) & (g2013) & (!g2014) & (g2037) & (g2045)) + ((!g8) & (g18) & (g2013) & (g2014) & (!g2037) & (g2045)) + ((!g8) & (g18) & (g2013) & (g2014) & (g2037) & (g2045)) + ((g8) & (!g18) & (!g2013) & (!g2014) & (!g2037) & (!g2045)) + ((g8) & (!g18) & (!g2013) & (!g2014) & (g2037) & (!g2045)) + ((g8) & (!g18) & (!g2013) & (g2014) & (!g2037) & (!g2045)) + ((g8) & (!g18) & (g2013) & (!g2014) & (!g2037) & (g2045)) + ((g8) & (!g18) & (g2013) & (!g2014) & (g2037) & (g2045)) + ((g8) & (!g18) & (g2013) & (g2014) & (!g2037) & (g2045)) + ((g8) & (!g18) & (g2013) & (g2014) & (g2037) & (!g2045)) + ((g8) & (!g18) & (g2013) & (g2014) & (g2037) & (g2045)) + ((g8) & (g18) & (!g2013) & (!g2014) & (!g2037) & (!g2045)) + ((g8) & (g18) & (g2013) & (!g2014) & (!g2037) & (g2045)) + ((g8) & (g18) & (g2013) & (!g2014) & (g2037) & (!g2045)) + ((g8) & (g18) & (g2013) & (!g2014) & (g2037) & (g2045)) + ((g8) & (g18) & (g2013) & (g2014) & (!g2037) & (!g2045)) + ((g8) & (g18) & (g2013) & (g2014) & (!g2037) & (g2045)) + ((g8) & (g18) & (g2013) & (g2014) & (g2037) & (!g2045)) + ((g8) & (g18) & (g2013) & (g2014) & (g2037) & (g2045)));
	assign g2098 = (((!g18) & (!g2014) & (g2037) & (!g2045)) + ((!g18) & (g2014) & (!g2037) & (!g2045)) + ((!g18) & (g2014) & (!g2037) & (g2045)) + ((!g18) & (g2014) & (g2037) & (g2045)) + ((g18) & (!g2014) & (!g2037) & (!g2045)) + ((g18) & (g2014) & (!g2037) & (g2045)) + ((g18) & (g2014) & (g2037) & (!g2045)) + ((g18) & (g2014) & (g2037) & (g2045)));
	assign g2099 = (((!g27) & (!g39) & (!g2016) & (g2017) & (g2036) & (!g2045)) + ((!g27) & (!g39) & (g2016) & (!g2017) & (!g2036) & (!g2045)) + ((!g27) & (!g39) & (g2016) & (!g2017) & (!g2036) & (g2045)) + ((!g27) & (!g39) & (g2016) & (!g2017) & (g2036) & (!g2045)) + ((!g27) & (!g39) & (g2016) & (!g2017) & (g2036) & (g2045)) + ((!g27) & (!g39) & (g2016) & (g2017) & (!g2036) & (!g2045)) + ((!g27) & (!g39) & (g2016) & (g2017) & (!g2036) & (g2045)) + ((!g27) & (!g39) & (g2016) & (g2017) & (g2036) & (g2045)) + ((!g27) & (g39) & (!g2016) & (!g2017) & (g2036) & (!g2045)) + ((!g27) & (g39) & (!g2016) & (g2017) & (!g2036) & (!g2045)) + ((!g27) & (g39) & (!g2016) & (g2017) & (g2036) & (!g2045)) + ((!g27) & (g39) & (g2016) & (!g2017) & (!g2036) & (!g2045)) + ((!g27) & (g39) & (g2016) & (!g2017) & (!g2036) & (g2045)) + ((!g27) & (g39) & (g2016) & (!g2017) & (g2036) & (g2045)) + ((!g27) & (g39) & (g2016) & (g2017) & (!g2036) & (g2045)) + ((!g27) & (g39) & (g2016) & (g2017) & (g2036) & (g2045)) + ((g27) & (!g39) & (!g2016) & (!g2017) & (!g2036) & (!g2045)) + ((g27) & (!g39) & (!g2016) & (!g2017) & (g2036) & (!g2045)) + ((g27) & (!g39) & (!g2016) & (g2017) & (!g2036) & (!g2045)) + ((g27) & (!g39) & (g2016) & (!g2017) & (!g2036) & (g2045)) + ((g27) & (!g39) & (g2016) & (!g2017) & (g2036) & (g2045)) + ((g27) & (!g39) & (g2016) & (g2017) & (!g2036) & (g2045)) + ((g27) & (!g39) & (g2016) & (g2017) & (g2036) & (!g2045)) + ((g27) & (!g39) & (g2016) & (g2017) & (g2036) & (g2045)) + ((g27) & (g39) & (!g2016) & (!g2017) & (!g2036) & (!g2045)) + ((g27) & (g39) & (g2016) & (!g2017) & (!g2036) & (g2045)) + ((g27) & (g39) & (g2016) & (!g2017) & (g2036) & (!g2045)) + ((g27) & (g39) & (g2016) & (!g2017) & (g2036) & (g2045)) + ((g27) & (g39) & (g2016) & (g2017) & (!g2036) & (!g2045)) + ((g27) & (g39) & (g2016) & (g2017) & (!g2036) & (g2045)) + ((g27) & (g39) & (g2016) & (g2017) & (g2036) & (!g2045)) + ((g27) & (g39) & (g2016) & (g2017) & (g2036) & (g2045)));
	assign g2100 = (((!g39) & (!g2017) & (g2036) & (!g2045)) + ((!g39) & (g2017) & (!g2036) & (!g2045)) + ((!g39) & (g2017) & (!g2036) & (g2045)) + ((!g39) & (g2017) & (g2036) & (g2045)) + ((g39) & (!g2017) & (!g2036) & (!g2045)) + ((g39) & (g2017) & (!g2036) & (g2045)) + ((g39) & (g2017) & (g2036) & (!g2045)) + ((g39) & (g2017) & (g2036) & (g2045)));
	assign g2101 = (((!g54) & (!g68) & (!g2019) & (g2020) & (g2035) & (!g2045)) + ((!g54) & (!g68) & (g2019) & (!g2020) & (!g2035) & (!g2045)) + ((!g54) & (!g68) & (g2019) & (!g2020) & (!g2035) & (g2045)) + ((!g54) & (!g68) & (g2019) & (!g2020) & (g2035) & (!g2045)) + ((!g54) & (!g68) & (g2019) & (!g2020) & (g2035) & (g2045)) + ((!g54) & (!g68) & (g2019) & (g2020) & (!g2035) & (!g2045)) + ((!g54) & (!g68) & (g2019) & (g2020) & (!g2035) & (g2045)) + ((!g54) & (!g68) & (g2019) & (g2020) & (g2035) & (g2045)) + ((!g54) & (g68) & (!g2019) & (!g2020) & (g2035) & (!g2045)) + ((!g54) & (g68) & (!g2019) & (g2020) & (!g2035) & (!g2045)) + ((!g54) & (g68) & (!g2019) & (g2020) & (g2035) & (!g2045)) + ((!g54) & (g68) & (g2019) & (!g2020) & (!g2035) & (!g2045)) + ((!g54) & (g68) & (g2019) & (!g2020) & (!g2035) & (g2045)) + ((!g54) & (g68) & (g2019) & (!g2020) & (g2035) & (g2045)) + ((!g54) & (g68) & (g2019) & (g2020) & (!g2035) & (g2045)) + ((!g54) & (g68) & (g2019) & (g2020) & (g2035) & (g2045)) + ((g54) & (!g68) & (!g2019) & (!g2020) & (!g2035) & (!g2045)) + ((g54) & (!g68) & (!g2019) & (!g2020) & (g2035) & (!g2045)) + ((g54) & (!g68) & (!g2019) & (g2020) & (!g2035) & (!g2045)) + ((g54) & (!g68) & (g2019) & (!g2020) & (!g2035) & (g2045)) + ((g54) & (!g68) & (g2019) & (!g2020) & (g2035) & (g2045)) + ((g54) & (!g68) & (g2019) & (g2020) & (!g2035) & (g2045)) + ((g54) & (!g68) & (g2019) & (g2020) & (g2035) & (!g2045)) + ((g54) & (!g68) & (g2019) & (g2020) & (g2035) & (g2045)) + ((g54) & (g68) & (!g2019) & (!g2020) & (!g2035) & (!g2045)) + ((g54) & (g68) & (g2019) & (!g2020) & (!g2035) & (g2045)) + ((g54) & (g68) & (g2019) & (!g2020) & (g2035) & (!g2045)) + ((g54) & (g68) & (g2019) & (!g2020) & (g2035) & (g2045)) + ((g54) & (g68) & (g2019) & (g2020) & (!g2035) & (!g2045)) + ((g54) & (g68) & (g2019) & (g2020) & (!g2035) & (g2045)) + ((g54) & (g68) & (g2019) & (g2020) & (g2035) & (!g2045)) + ((g54) & (g68) & (g2019) & (g2020) & (g2035) & (g2045)));
	assign g2102 = (((!g68) & (!g2020) & (g2035) & (!g2045)) + ((!g68) & (g2020) & (!g2035) & (!g2045)) + ((!g68) & (g2020) & (!g2035) & (g2045)) + ((!g68) & (g2020) & (g2035) & (g2045)) + ((g68) & (!g2020) & (!g2035) & (!g2045)) + ((g68) & (g2020) & (!g2035) & (g2045)) + ((g68) & (g2020) & (g2035) & (!g2045)) + ((g68) & (g2020) & (g2035) & (g2045)));
	assign g2103 = (((!g87) & (!g104) & (!g2022) & (g2023) & (g2034) & (!g2045)) + ((!g87) & (!g104) & (g2022) & (!g2023) & (!g2034) & (!g2045)) + ((!g87) & (!g104) & (g2022) & (!g2023) & (!g2034) & (g2045)) + ((!g87) & (!g104) & (g2022) & (!g2023) & (g2034) & (!g2045)) + ((!g87) & (!g104) & (g2022) & (!g2023) & (g2034) & (g2045)) + ((!g87) & (!g104) & (g2022) & (g2023) & (!g2034) & (!g2045)) + ((!g87) & (!g104) & (g2022) & (g2023) & (!g2034) & (g2045)) + ((!g87) & (!g104) & (g2022) & (g2023) & (g2034) & (g2045)) + ((!g87) & (g104) & (!g2022) & (!g2023) & (g2034) & (!g2045)) + ((!g87) & (g104) & (!g2022) & (g2023) & (!g2034) & (!g2045)) + ((!g87) & (g104) & (!g2022) & (g2023) & (g2034) & (!g2045)) + ((!g87) & (g104) & (g2022) & (!g2023) & (!g2034) & (!g2045)) + ((!g87) & (g104) & (g2022) & (!g2023) & (!g2034) & (g2045)) + ((!g87) & (g104) & (g2022) & (!g2023) & (g2034) & (g2045)) + ((!g87) & (g104) & (g2022) & (g2023) & (!g2034) & (g2045)) + ((!g87) & (g104) & (g2022) & (g2023) & (g2034) & (g2045)) + ((g87) & (!g104) & (!g2022) & (!g2023) & (!g2034) & (!g2045)) + ((g87) & (!g104) & (!g2022) & (!g2023) & (g2034) & (!g2045)) + ((g87) & (!g104) & (!g2022) & (g2023) & (!g2034) & (!g2045)) + ((g87) & (!g104) & (g2022) & (!g2023) & (!g2034) & (g2045)) + ((g87) & (!g104) & (g2022) & (!g2023) & (g2034) & (g2045)) + ((g87) & (!g104) & (g2022) & (g2023) & (!g2034) & (g2045)) + ((g87) & (!g104) & (g2022) & (g2023) & (g2034) & (!g2045)) + ((g87) & (!g104) & (g2022) & (g2023) & (g2034) & (g2045)) + ((g87) & (g104) & (!g2022) & (!g2023) & (!g2034) & (!g2045)) + ((g87) & (g104) & (g2022) & (!g2023) & (!g2034) & (g2045)) + ((g87) & (g104) & (g2022) & (!g2023) & (g2034) & (!g2045)) + ((g87) & (g104) & (g2022) & (!g2023) & (g2034) & (g2045)) + ((g87) & (g104) & (g2022) & (g2023) & (!g2034) & (!g2045)) + ((g87) & (g104) & (g2022) & (g2023) & (!g2034) & (g2045)) + ((g87) & (g104) & (g2022) & (g2023) & (g2034) & (!g2045)) + ((g87) & (g104) & (g2022) & (g2023) & (g2034) & (g2045)));
	assign g2104 = (((!g104) & (!g2023) & (g2034) & (!g2045)) + ((!g104) & (g2023) & (!g2034) & (!g2045)) + ((!g104) & (g2023) & (!g2034) & (g2045)) + ((!g104) & (g2023) & (g2034) & (g2045)) + ((g104) & (!g2023) & (!g2034) & (!g2045)) + ((g104) & (g2023) & (!g2034) & (g2045)) + ((g104) & (g2023) & (g2034) & (!g2045)) + ((g104) & (g2023) & (g2034) & (g2045)));
	assign g2105 = (((!g127) & (!g147) & (!g2025) & (g2026) & (g2033) & (!g2045)) + ((!g127) & (!g147) & (g2025) & (!g2026) & (!g2033) & (!g2045)) + ((!g127) & (!g147) & (g2025) & (!g2026) & (!g2033) & (g2045)) + ((!g127) & (!g147) & (g2025) & (!g2026) & (g2033) & (!g2045)) + ((!g127) & (!g147) & (g2025) & (!g2026) & (g2033) & (g2045)) + ((!g127) & (!g147) & (g2025) & (g2026) & (!g2033) & (!g2045)) + ((!g127) & (!g147) & (g2025) & (g2026) & (!g2033) & (g2045)) + ((!g127) & (!g147) & (g2025) & (g2026) & (g2033) & (g2045)) + ((!g127) & (g147) & (!g2025) & (!g2026) & (g2033) & (!g2045)) + ((!g127) & (g147) & (!g2025) & (g2026) & (!g2033) & (!g2045)) + ((!g127) & (g147) & (!g2025) & (g2026) & (g2033) & (!g2045)) + ((!g127) & (g147) & (g2025) & (!g2026) & (!g2033) & (!g2045)) + ((!g127) & (g147) & (g2025) & (!g2026) & (!g2033) & (g2045)) + ((!g127) & (g147) & (g2025) & (!g2026) & (g2033) & (g2045)) + ((!g127) & (g147) & (g2025) & (g2026) & (!g2033) & (g2045)) + ((!g127) & (g147) & (g2025) & (g2026) & (g2033) & (g2045)) + ((g127) & (!g147) & (!g2025) & (!g2026) & (!g2033) & (!g2045)) + ((g127) & (!g147) & (!g2025) & (!g2026) & (g2033) & (!g2045)) + ((g127) & (!g147) & (!g2025) & (g2026) & (!g2033) & (!g2045)) + ((g127) & (!g147) & (g2025) & (!g2026) & (!g2033) & (g2045)) + ((g127) & (!g147) & (g2025) & (!g2026) & (g2033) & (g2045)) + ((g127) & (!g147) & (g2025) & (g2026) & (!g2033) & (g2045)) + ((g127) & (!g147) & (g2025) & (g2026) & (g2033) & (!g2045)) + ((g127) & (!g147) & (g2025) & (g2026) & (g2033) & (g2045)) + ((g127) & (g147) & (!g2025) & (!g2026) & (!g2033) & (!g2045)) + ((g127) & (g147) & (g2025) & (!g2026) & (!g2033) & (g2045)) + ((g127) & (g147) & (g2025) & (!g2026) & (g2033) & (!g2045)) + ((g127) & (g147) & (g2025) & (!g2026) & (g2033) & (g2045)) + ((g127) & (g147) & (g2025) & (g2026) & (!g2033) & (!g2045)) + ((g127) & (g147) & (g2025) & (g2026) & (!g2033) & (g2045)) + ((g127) & (g147) & (g2025) & (g2026) & (g2033) & (!g2045)) + ((g127) & (g147) & (g2025) & (g2026) & (g2033) & (g2045)));
	assign g2106 = (((!g147) & (!g2026) & (g2033) & (!g2045)) + ((!g147) & (g2026) & (!g2033) & (!g2045)) + ((!g147) & (g2026) & (!g2033) & (g2045)) + ((!g147) & (g2026) & (g2033) & (g2045)) + ((g147) & (!g2026) & (!g2033) & (!g2045)) + ((g147) & (g2026) & (!g2033) & (g2045)) + ((g147) & (g2026) & (g2033) & (!g2045)) + ((g147) & (g2026) & (g2033) & (g2045)));
	assign g2107 = (((!g174) & (!g198) & (!g2028) & (g2029) & (g2032) & (!g2045)) + ((!g174) & (!g198) & (g2028) & (!g2029) & (!g2032) & (!g2045)) + ((!g174) & (!g198) & (g2028) & (!g2029) & (!g2032) & (g2045)) + ((!g174) & (!g198) & (g2028) & (!g2029) & (g2032) & (!g2045)) + ((!g174) & (!g198) & (g2028) & (!g2029) & (g2032) & (g2045)) + ((!g174) & (!g198) & (g2028) & (g2029) & (!g2032) & (!g2045)) + ((!g174) & (!g198) & (g2028) & (g2029) & (!g2032) & (g2045)) + ((!g174) & (!g198) & (g2028) & (g2029) & (g2032) & (g2045)) + ((!g174) & (g198) & (!g2028) & (!g2029) & (g2032) & (!g2045)) + ((!g174) & (g198) & (!g2028) & (g2029) & (!g2032) & (!g2045)) + ((!g174) & (g198) & (!g2028) & (g2029) & (g2032) & (!g2045)) + ((!g174) & (g198) & (g2028) & (!g2029) & (!g2032) & (!g2045)) + ((!g174) & (g198) & (g2028) & (!g2029) & (!g2032) & (g2045)) + ((!g174) & (g198) & (g2028) & (!g2029) & (g2032) & (g2045)) + ((!g174) & (g198) & (g2028) & (g2029) & (!g2032) & (g2045)) + ((!g174) & (g198) & (g2028) & (g2029) & (g2032) & (g2045)) + ((g174) & (!g198) & (!g2028) & (!g2029) & (!g2032) & (!g2045)) + ((g174) & (!g198) & (!g2028) & (!g2029) & (g2032) & (!g2045)) + ((g174) & (!g198) & (!g2028) & (g2029) & (!g2032) & (!g2045)) + ((g174) & (!g198) & (g2028) & (!g2029) & (!g2032) & (g2045)) + ((g174) & (!g198) & (g2028) & (!g2029) & (g2032) & (g2045)) + ((g174) & (!g198) & (g2028) & (g2029) & (!g2032) & (g2045)) + ((g174) & (!g198) & (g2028) & (g2029) & (g2032) & (!g2045)) + ((g174) & (!g198) & (g2028) & (g2029) & (g2032) & (g2045)) + ((g174) & (g198) & (!g2028) & (!g2029) & (!g2032) & (!g2045)) + ((g174) & (g198) & (g2028) & (!g2029) & (!g2032) & (g2045)) + ((g174) & (g198) & (g2028) & (!g2029) & (g2032) & (!g2045)) + ((g174) & (g198) & (g2028) & (!g2029) & (g2032) & (g2045)) + ((g174) & (g198) & (g2028) & (g2029) & (!g2032) & (!g2045)) + ((g174) & (g198) & (g2028) & (g2029) & (!g2032) & (g2045)) + ((g174) & (g198) & (g2028) & (g2029) & (g2032) & (!g2045)) + ((g174) & (g198) & (g2028) & (g2029) & (g2032) & (g2045)));
	assign g2108 = (((!g198) & (!g2029) & (g2032) & (!g2045)) + ((!g198) & (g2029) & (!g2032) & (!g2045)) + ((!g198) & (g2029) & (!g2032) & (g2045)) + ((!g198) & (g2029) & (g2032) & (g2045)) + ((g198) & (!g2029) & (!g2032) & (!g2045)) + ((g198) & (g2029) & (!g2032) & (g2045)) + ((g198) & (g2029) & (g2032) & (!g2045)) + ((g198) & (g2029) & (g2032) & (g2045)));
	assign g2109 = (((!g229) & (!g255) & (!g2031) & (g1951) & (g2009) & (!g2045)) + ((!g229) & (!g255) & (g2031) & (!g1951) & (!g2009) & (!g2045)) + ((!g229) & (!g255) & (g2031) & (!g1951) & (!g2009) & (g2045)) + ((!g229) & (!g255) & (g2031) & (!g1951) & (g2009) & (!g2045)) + ((!g229) & (!g255) & (g2031) & (!g1951) & (g2009) & (g2045)) + ((!g229) & (!g255) & (g2031) & (g1951) & (!g2009) & (!g2045)) + ((!g229) & (!g255) & (g2031) & (g1951) & (!g2009) & (g2045)) + ((!g229) & (!g255) & (g2031) & (g1951) & (g2009) & (g2045)) + ((!g229) & (g255) & (!g2031) & (!g1951) & (g2009) & (!g2045)) + ((!g229) & (g255) & (!g2031) & (g1951) & (!g2009) & (!g2045)) + ((!g229) & (g255) & (!g2031) & (g1951) & (g2009) & (!g2045)) + ((!g229) & (g255) & (g2031) & (!g1951) & (!g2009) & (!g2045)) + ((!g229) & (g255) & (g2031) & (!g1951) & (!g2009) & (g2045)) + ((!g229) & (g255) & (g2031) & (!g1951) & (g2009) & (g2045)) + ((!g229) & (g255) & (g2031) & (g1951) & (!g2009) & (g2045)) + ((!g229) & (g255) & (g2031) & (g1951) & (g2009) & (g2045)) + ((g229) & (!g255) & (!g2031) & (!g1951) & (!g2009) & (!g2045)) + ((g229) & (!g255) & (!g2031) & (!g1951) & (g2009) & (!g2045)) + ((g229) & (!g255) & (!g2031) & (g1951) & (!g2009) & (!g2045)) + ((g229) & (!g255) & (g2031) & (!g1951) & (!g2009) & (g2045)) + ((g229) & (!g255) & (g2031) & (!g1951) & (g2009) & (g2045)) + ((g229) & (!g255) & (g2031) & (g1951) & (!g2009) & (g2045)) + ((g229) & (!g255) & (g2031) & (g1951) & (g2009) & (!g2045)) + ((g229) & (!g255) & (g2031) & (g1951) & (g2009) & (g2045)) + ((g229) & (g255) & (!g2031) & (!g1951) & (!g2009) & (!g2045)) + ((g229) & (g255) & (g2031) & (!g1951) & (!g2009) & (g2045)) + ((g229) & (g255) & (g2031) & (!g1951) & (g2009) & (!g2045)) + ((g229) & (g255) & (g2031) & (!g1951) & (g2009) & (g2045)) + ((g229) & (g255) & (g2031) & (g1951) & (!g2009) & (!g2045)) + ((g229) & (g255) & (g2031) & (g1951) & (!g2009) & (g2045)) + ((g229) & (g255) & (g2031) & (g1951) & (g2009) & (!g2045)) + ((g229) & (g255) & (g2031) & (g1951) & (g2009) & (g2045)));
	assign g2110 = (((!g198) & (!g229) & (g2109) & (g2046) & (g2094)) + ((!g198) & (g229) & (g2109) & (!g2046) & (g2094)) + ((!g198) & (g229) & (g2109) & (g2046) & (!g2094)) + ((!g198) & (g229) & (g2109) & (g2046) & (g2094)) + ((g198) & (!g229) & (!g2109) & (g2046) & (g2094)) + ((g198) & (!g229) & (g2109) & (!g2046) & (!g2094)) + ((g198) & (!g229) & (g2109) & (!g2046) & (g2094)) + ((g198) & (!g229) & (g2109) & (g2046) & (!g2094)) + ((g198) & (!g229) & (g2109) & (g2046) & (g2094)) + ((g198) & (g229) & (!g2109) & (!g2046) & (g2094)) + ((g198) & (g229) & (!g2109) & (g2046) & (!g2094)) + ((g198) & (g229) & (!g2109) & (g2046) & (g2094)) + ((g198) & (g229) & (g2109) & (!g2046) & (!g2094)) + ((g198) & (g229) & (g2109) & (!g2046) & (g2094)) + ((g198) & (g229) & (g2109) & (g2046) & (!g2094)) + ((g198) & (g229) & (g2109) & (g2046) & (g2094)));
	assign g2111 = (((!g147) & (!g174) & (g2107) & (g2108) & (g2110)) + ((!g147) & (g174) & (g2107) & (!g2108) & (g2110)) + ((!g147) & (g174) & (g2107) & (g2108) & (!g2110)) + ((!g147) & (g174) & (g2107) & (g2108) & (g2110)) + ((g147) & (!g174) & (!g2107) & (g2108) & (g2110)) + ((g147) & (!g174) & (g2107) & (!g2108) & (!g2110)) + ((g147) & (!g174) & (g2107) & (!g2108) & (g2110)) + ((g147) & (!g174) & (g2107) & (g2108) & (!g2110)) + ((g147) & (!g174) & (g2107) & (g2108) & (g2110)) + ((g147) & (g174) & (!g2107) & (!g2108) & (g2110)) + ((g147) & (g174) & (!g2107) & (g2108) & (!g2110)) + ((g147) & (g174) & (!g2107) & (g2108) & (g2110)) + ((g147) & (g174) & (g2107) & (!g2108) & (!g2110)) + ((g147) & (g174) & (g2107) & (!g2108) & (g2110)) + ((g147) & (g174) & (g2107) & (g2108) & (!g2110)) + ((g147) & (g174) & (g2107) & (g2108) & (g2110)));
	assign g2112 = (((!g104) & (!g127) & (g2105) & (g2106) & (g2111)) + ((!g104) & (g127) & (g2105) & (!g2106) & (g2111)) + ((!g104) & (g127) & (g2105) & (g2106) & (!g2111)) + ((!g104) & (g127) & (g2105) & (g2106) & (g2111)) + ((g104) & (!g127) & (!g2105) & (g2106) & (g2111)) + ((g104) & (!g127) & (g2105) & (!g2106) & (!g2111)) + ((g104) & (!g127) & (g2105) & (!g2106) & (g2111)) + ((g104) & (!g127) & (g2105) & (g2106) & (!g2111)) + ((g104) & (!g127) & (g2105) & (g2106) & (g2111)) + ((g104) & (g127) & (!g2105) & (!g2106) & (g2111)) + ((g104) & (g127) & (!g2105) & (g2106) & (!g2111)) + ((g104) & (g127) & (!g2105) & (g2106) & (g2111)) + ((g104) & (g127) & (g2105) & (!g2106) & (!g2111)) + ((g104) & (g127) & (g2105) & (!g2106) & (g2111)) + ((g104) & (g127) & (g2105) & (g2106) & (!g2111)) + ((g104) & (g127) & (g2105) & (g2106) & (g2111)));
	assign g2113 = (((!g68) & (!g87) & (g2103) & (g2104) & (g2112)) + ((!g68) & (g87) & (g2103) & (!g2104) & (g2112)) + ((!g68) & (g87) & (g2103) & (g2104) & (!g2112)) + ((!g68) & (g87) & (g2103) & (g2104) & (g2112)) + ((g68) & (!g87) & (!g2103) & (g2104) & (g2112)) + ((g68) & (!g87) & (g2103) & (!g2104) & (!g2112)) + ((g68) & (!g87) & (g2103) & (!g2104) & (g2112)) + ((g68) & (!g87) & (g2103) & (g2104) & (!g2112)) + ((g68) & (!g87) & (g2103) & (g2104) & (g2112)) + ((g68) & (g87) & (!g2103) & (!g2104) & (g2112)) + ((g68) & (g87) & (!g2103) & (g2104) & (!g2112)) + ((g68) & (g87) & (!g2103) & (g2104) & (g2112)) + ((g68) & (g87) & (g2103) & (!g2104) & (!g2112)) + ((g68) & (g87) & (g2103) & (!g2104) & (g2112)) + ((g68) & (g87) & (g2103) & (g2104) & (!g2112)) + ((g68) & (g87) & (g2103) & (g2104) & (g2112)));
	assign g2114 = (((!g39) & (!g54) & (g2101) & (g2102) & (g2113)) + ((!g39) & (g54) & (g2101) & (!g2102) & (g2113)) + ((!g39) & (g54) & (g2101) & (g2102) & (!g2113)) + ((!g39) & (g54) & (g2101) & (g2102) & (g2113)) + ((g39) & (!g54) & (!g2101) & (g2102) & (g2113)) + ((g39) & (!g54) & (g2101) & (!g2102) & (!g2113)) + ((g39) & (!g54) & (g2101) & (!g2102) & (g2113)) + ((g39) & (!g54) & (g2101) & (g2102) & (!g2113)) + ((g39) & (!g54) & (g2101) & (g2102) & (g2113)) + ((g39) & (g54) & (!g2101) & (!g2102) & (g2113)) + ((g39) & (g54) & (!g2101) & (g2102) & (!g2113)) + ((g39) & (g54) & (!g2101) & (g2102) & (g2113)) + ((g39) & (g54) & (g2101) & (!g2102) & (!g2113)) + ((g39) & (g54) & (g2101) & (!g2102) & (g2113)) + ((g39) & (g54) & (g2101) & (g2102) & (!g2113)) + ((g39) & (g54) & (g2101) & (g2102) & (g2113)));
	assign g2115 = (((!g18) & (!g27) & (g2099) & (g2100) & (g2114)) + ((!g18) & (g27) & (g2099) & (!g2100) & (g2114)) + ((!g18) & (g27) & (g2099) & (g2100) & (!g2114)) + ((!g18) & (g27) & (g2099) & (g2100) & (g2114)) + ((g18) & (!g27) & (!g2099) & (g2100) & (g2114)) + ((g18) & (!g27) & (g2099) & (!g2100) & (!g2114)) + ((g18) & (!g27) & (g2099) & (!g2100) & (g2114)) + ((g18) & (!g27) & (g2099) & (g2100) & (!g2114)) + ((g18) & (!g27) & (g2099) & (g2100) & (g2114)) + ((g18) & (g27) & (!g2099) & (!g2100) & (g2114)) + ((g18) & (g27) & (!g2099) & (g2100) & (!g2114)) + ((g18) & (g27) & (!g2099) & (g2100) & (g2114)) + ((g18) & (g27) & (g2099) & (!g2100) & (!g2114)) + ((g18) & (g27) & (g2099) & (!g2100) & (g2114)) + ((g18) & (g27) & (g2099) & (g2100) & (!g2114)) + ((g18) & (g27) & (g2099) & (g2100) & (g2114)));
	assign g2116 = (((!g2) & (!g8) & (g2097) & (g2098) & (g2115)) + ((!g2) & (g8) & (g2097) & (!g2098) & (g2115)) + ((!g2) & (g8) & (g2097) & (g2098) & (!g2115)) + ((!g2) & (g8) & (g2097) & (g2098) & (g2115)) + ((g2) & (!g8) & (!g2097) & (g2098) & (g2115)) + ((g2) & (!g8) & (g2097) & (!g2098) & (!g2115)) + ((g2) & (!g8) & (g2097) & (!g2098) & (g2115)) + ((g2) & (!g8) & (g2097) & (g2098) & (!g2115)) + ((g2) & (!g8) & (g2097) & (g2098) & (g2115)) + ((g2) & (g8) & (!g2097) & (!g2098) & (g2115)) + ((g2) & (g8) & (!g2097) & (g2098) & (!g2115)) + ((g2) & (g8) & (!g2097) & (g2098) & (g2115)) + ((g2) & (g8) & (g2097) & (!g2098) & (!g2115)) + ((g2) & (g8) & (g2097) & (!g2098) & (g2115)) + ((g2) & (g8) & (g2097) & (g2098) & (!g2115)) + ((g2) & (g8) & (g2097) & (g2098) & (g2115)));
	assign g2117 = (((!g2) & (!g2011) & (g2038) & (!g2045)) + ((!g2) & (g2011) & (!g2038) & (!g2045)) + ((!g2) & (g2011) & (!g2038) & (g2045)) + ((!g2) & (g2011) & (g2038) & (g2045)) + ((g2) & (!g2011) & (!g2038) & (!g2045)) + ((g2) & (g2011) & (!g2038) & (g2045)) + ((g2) & (g2011) & (g2038) & (!g2045)) + ((g2) & (g2011) & (g2038) & (g2045)));
	assign g2118 = (((!g1) & (!g2010) & (!g2041) & (!g2043) & (g2044)) + ((!g1) & (!g2010) & (!g2041) & (g2043) & (!g2044)) + ((!g1) & (!g2010) & (!g2041) & (g2043) & (g2044)) + ((!g1) & (g2010) & (g2041) & (!g2043) & (!g2044)) + ((!g1) & (g2010) & (g2041) & (!g2043) & (g2044)) + ((!g1) & (g2010) & (g2041) & (g2043) & (!g2044)) + ((!g1) & (g2010) & (g2041) & (g2043) & (g2044)) + ((g1) & (!g2010) & (!g2041) & (!g2043) & (g2044)) + ((g1) & (!g2010) & (!g2041) & (g2043) & (g2044)) + ((g1) & (g2010) & (g2041) & (!g2043) & (!g2044)) + ((g1) & (g2010) & (g2041) & (!g2043) & (g2044)) + ((g1) & (g2010) & (g2041) & (g2043) & (!g2044)) + ((g1) & (g2010) & (g2041) & (g2043) & (g2044)));
	assign g2119 = (((!g4) & (!g1) & (!g2096) & (!g2116) & (!g2117) & (!g2118)) + ((!g4) & (g1) & (!g2096) & (!g2116) & (!g2117) & (!g2118)) + ((!g4) & (g1) & (!g2096) & (!g2116) & (!g2117) & (g2118)) + ((!g4) & (g1) & (!g2096) & (!g2116) & (g2117) & (!g2118)) + ((!g4) & (g1) & (!g2096) & (!g2116) & (g2117) & (g2118)) + ((!g4) & (g1) & (!g2096) & (g2116) & (!g2117) & (!g2118)) + ((!g4) & (g1) & (!g2096) & (g2116) & (!g2117) & (g2118)) + ((!g4) & (g1) & (!g2096) & (g2116) & (g2117) & (!g2118)) + ((!g4) & (g1) & (!g2096) & (g2116) & (g2117) & (g2118)) + ((!g4) & (g1) & (g2096) & (!g2116) & (!g2117) & (!g2118)) + ((!g4) & (g1) & (g2096) & (!g2116) & (!g2117) & (g2118)) + ((g4) & (!g1) & (!g2096) & (!g2116) & (!g2117) & (!g2118)) + ((g4) & (!g1) & (!g2096) & (!g2116) & (g2117) & (!g2118)) + ((g4) & (!g1) & (!g2096) & (g2116) & (!g2117) & (!g2118)) + ((g4) & (g1) & (!g2096) & (!g2116) & (!g2117) & (!g2118)) + ((g4) & (g1) & (!g2096) & (!g2116) & (!g2117) & (g2118)) + ((g4) & (g1) & (!g2096) & (!g2116) & (g2117) & (!g2118)) + ((g4) & (g1) & (!g2096) & (!g2116) & (g2117) & (g2118)) + ((g4) & (g1) & (!g2096) & (g2116) & (!g2117) & (!g2118)) + ((g4) & (g1) & (!g2096) & (g2116) & (!g2117) & (g2118)) + ((g4) & (g1) & (!g2096) & (g2116) & (g2117) & (!g2118)) + ((g4) & (g1) & (!g2096) & (g2116) & (g2117) & (g2118)) + ((g4) & (g1) & (g2096) & (!g2116) & (!g2117) & (!g2118)) + ((g4) & (g1) & (g2096) & (!g2116) & (!g2117) & (g2118)) + ((g4) & (g1) & (g2096) & (!g2116) & (g2117) & (!g2118)) + ((g4) & (g1) & (g2096) & (!g2116) & (g2117) & (g2118)) + ((g4) & (g1) & (g2096) & (g2116) & (!g2117) & (!g2118)) + ((g4) & (g1) & (g2096) & (g2116) & (!g2117) & (g2118)));
	assign g2120 = (((!g229) & (!g2046) & (g2094) & (!g2095) & (!g2119)) + ((!g229) & (!g2046) & (g2094) & (g2095) & (!g2119)) + ((!g229) & (!g2046) & (g2094) & (g2095) & (g2119)) + ((!g229) & (g2046) & (!g2094) & (!g2095) & (!g2119)) + ((!g229) & (g2046) & (!g2094) & (!g2095) & (g2119)) + ((!g229) & (g2046) & (!g2094) & (g2095) & (!g2119)) + ((!g229) & (g2046) & (!g2094) & (g2095) & (g2119)) + ((!g229) & (g2046) & (g2094) & (!g2095) & (g2119)) + ((g229) & (!g2046) & (!g2094) & (!g2095) & (!g2119)) + ((g229) & (!g2046) & (!g2094) & (g2095) & (!g2119)) + ((g229) & (!g2046) & (!g2094) & (g2095) & (g2119)) + ((g229) & (g2046) & (!g2094) & (!g2095) & (g2119)) + ((g229) & (g2046) & (g2094) & (!g2095) & (!g2119)) + ((g229) & (g2046) & (g2094) & (!g2095) & (g2119)) + ((g229) & (g2046) & (g2094) & (g2095) & (!g2119)) + ((g229) & (g2046) & (g2094) & (g2095) & (g2119)));
	assign g2121 = (((!g255) & (!g290) & (g2048) & (g2093)) + ((!g255) & (g290) & (!g2048) & (g2093)) + ((!g255) & (g290) & (g2048) & (!g2093)) + ((!g255) & (g290) & (g2048) & (g2093)) + ((g255) & (!g290) & (!g2048) & (!g2093)) + ((g255) & (!g290) & (!g2048) & (g2093)) + ((g255) & (!g290) & (g2048) & (!g2093)) + ((g255) & (g290) & (!g2048) & (!g2093)));
	assign g2122 = (((!g2047) & (!g2095) & (!g2119) & (g2121)) + ((!g2047) & (g2095) & (!g2119) & (g2121)) + ((!g2047) & (g2095) & (g2119) & (g2121)) + ((g2047) & (!g2095) & (!g2119) & (!g2121)) + ((g2047) & (!g2095) & (g2119) & (!g2121)) + ((g2047) & (!g2095) & (g2119) & (g2121)) + ((g2047) & (g2095) & (!g2119) & (!g2121)) + ((g2047) & (g2095) & (g2119) & (!g2121)));
	assign g2123 = (((!g290) & (!g2048) & (g2093) & (!g2095) & (!g2119)) + ((!g290) & (!g2048) & (g2093) & (g2095) & (!g2119)) + ((!g290) & (!g2048) & (g2093) & (g2095) & (g2119)) + ((!g290) & (g2048) & (!g2093) & (!g2095) & (!g2119)) + ((!g290) & (g2048) & (!g2093) & (!g2095) & (g2119)) + ((!g290) & (g2048) & (!g2093) & (g2095) & (!g2119)) + ((!g290) & (g2048) & (!g2093) & (g2095) & (g2119)) + ((!g290) & (g2048) & (g2093) & (!g2095) & (g2119)) + ((g290) & (!g2048) & (!g2093) & (!g2095) & (!g2119)) + ((g290) & (!g2048) & (!g2093) & (g2095) & (!g2119)) + ((g290) & (!g2048) & (!g2093) & (g2095) & (g2119)) + ((g290) & (g2048) & (!g2093) & (!g2095) & (g2119)) + ((g290) & (g2048) & (g2093) & (!g2095) & (!g2119)) + ((g290) & (g2048) & (g2093) & (!g2095) & (g2119)) + ((g290) & (g2048) & (g2093) & (g2095) & (!g2119)) + ((g290) & (g2048) & (g2093) & (g2095) & (g2119)));
	assign g2124 = (((!g319) & (!g358) & (g2050) & (g2092)) + ((!g319) & (g358) & (!g2050) & (g2092)) + ((!g319) & (g358) & (g2050) & (!g2092)) + ((!g319) & (g358) & (g2050) & (g2092)) + ((g319) & (!g358) & (!g2050) & (!g2092)) + ((g319) & (!g358) & (!g2050) & (g2092)) + ((g319) & (!g358) & (g2050) & (!g2092)) + ((g319) & (g358) & (!g2050) & (!g2092)));
	assign g2125 = (((!g2049) & (!g2095) & (!g2119) & (g2124)) + ((!g2049) & (g2095) & (!g2119) & (g2124)) + ((!g2049) & (g2095) & (g2119) & (g2124)) + ((g2049) & (!g2095) & (!g2119) & (!g2124)) + ((g2049) & (!g2095) & (g2119) & (!g2124)) + ((g2049) & (!g2095) & (g2119) & (g2124)) + ((g2049) & (g2095) & (!g2119) & (!g2124)) + ((g2049) & (g2095) & (g2119) & (!g2124)));
	assign g2126 = (((!g358) & (!g2050) & (g2092) & (!g2095) & (!g2119)) + ((!g358) & (!g2050) & (g2092) & (g2095) & (!g2119)) + ((!g358) & (!g2050) & (g2092) & (g2095) & (g2119)) + ((!g358) & (g2050) & (!g2092) & (!g2095) & (!g2119)) + ((!g358) & (g2050) & (!g2092) & (!g2095) & (g2119)) + ((!g358) & (g2050) & (!g2092) & (g2095) & (!g2119)) + ((!g358) & (g2050) & (!g2092) & (g2095) & (g2119)) + ((!g358) & (g2050) & (g2092) & (!g2095) & (g2119)) + ((g358) & (!g2050) & (!g2092) & (!g2095) & (!g2119)) + ((g358) & (!g2050) & (!g2092) & (g2095) & (!g2119)) + ((g358) & (!g2050) & (!g2092) & (g2095) & (g2119)) + ((g358) & (g2050) & (!g2092) & (!g2095) & (g2119)) + ((g358) & (g2050) & (g2092) & (!g2095) & (!g2119)) + ((g358) & (g2050) & (g2092) & (!g2095) & (g2119)) + ((g358) & (g2050) & (g2092) & (g2095) & (!g2119)) + ((g358) & (g2050) & (g2092) & (g2095) & (g2119)));
	assign g2127 = (((!g390) & (!g433) & (g2052) & (g2091)) + ((!g390) & (g433) & (!g2052) & (g2091)) + ((!g390) & (g433) & (g2052) & (!g2091)) + ((!g390) & (g433) & (g2052) & (g2091)) + ((g390) & (!g433) & (!g2052) & (!g2091)) + ((g390) & (!g433) & (!g2052) & (g2091)) + ((g390) & (!g433) & (g2052) & (!g2091)) + ((g390) & (g433) & (!g2052) & (!g2091)));
	assign g2128 = (((!g2051) & (!g2095) & (!g2119) & (g2127)) + ((!g2051) & (g2095) & (!g2119) & (g2127)) + ((!g2051) & (g2095) & (g2119) & (g2127)) + ((g2051) & (!g2095) & (!g2119) & (!g2127)) + ((g2051) & (!g2095) & (g2119) & (!g2127)) + ((g2051) & (!g2095) & (g2119) & (g2127)) + ((g2051) & (g2095) & (!g2119) & (!g2127)) + ((g2051) & (g2095) & (g2119) & (!g2127)));
	assign g2129 = (((!g433) & (!g2052) & (g2091) & (!g2095) & (!g2119)) + ((!g433) & (!g2052) & (g2091) & (g2095) & (!g2119)) + ((!g433) & (!g2052) & (g2091) & (g2095) & (g2119)) + ((!g433) & (g2052) & (!g2091) & (!g2095) & (!g2119)) + ((!g433) & (g2052) & (!g2091) & (!g2095) & (g2119)) + ((!g433) & (g2052) & (!g2091) & (g2095) & (!g2119)) + ((!g433) & (g2052) & (!g2091) & (g2095) & (g2119)) + ((!g433) & (g2052) & (g2091) & (!g2095) & (g2119)) + ((g433) & (!g2052) & (!g2091) & (!g2095) & (!g2119)) + ((g433) & (!g2052) & (!g2091) & (g2095) & (!g2119)) + ((g433) & (!g2052) & (!g2091) & (g2095) & (g2119)) + ((g433) & (g2052) & (!g2091) & (!g2095) & (g2119)) + ((g433) & (g2052) & (g2091) & (!g2095) & (!g2119)) + ((g433) & (g2052) & (g2091) & (!g2095) & (g2119)) + ((g433) & (g2052) & (g2091) & (g2095) & (!g2119)) + ((g433) & (g2052) & (g2091) & (g2095) & (g2119)));
	assign g2130 = (((!g468) & (!g515) & (g2054) & (g2090)) + ((!g468) & (g515) & (!g2054) & (g2090)) + ((!g468) & (g515) & (g2054) & (!g2090)) + ((!g468) & (g515) & (g2054) & (g2090)) + ((g468) & (!g515) & (!g2054) & (!g2090)) + ((g468) & (!g515) & (!g2054) & (g2090)) + ((g468) & (!g515) & (g2054) & (!g2090)) + ((g468) & (g515) & (!g2054) & (!g2090)));
	assign g2131 = (((!g2053) & (!g2095) & (!g2119) & (g2130)) + ((!g2053) & (g2095) & (!g2119) & (g2130)) + ((!g2053) & (g2095) & (g2119) & (g2130)) + ((g2053) & (!g2095) & (!g2119) & (!g2130)) + ((g2053) & (!g2095) & (g2119) & (!g2130)) + ((g2053) & (!g2095) & (g2119) & (g2130)) + ((g2053) & (g2095) & (!g2119) & (!g2130)) + ((g2053) & (g2095) & (g2119) & (!g2130)));
	assign g2132 = (((!g515) & (!g2054) & (g2090) & (!g2095) & (!g2119)) + ((!g515) & (!g2054) & (g2090) & (g2095) & (!g2119)) + ((!g515) & (!g2054) & (g2090) & (g2095) & (g2119)) + ((!g515) & (g2054) & (!g2090) & (!g2095) & (!g2119)) + ((!g515) & (g2054) & (!g2090) & (!g2095) & (g2119)) + ((!g515) & (g2054) & (!g2090) & (g2095) & (!g2119)) + ((!g515) & (g2054) & (!g2090) & (g2095) & (g2119)) + ((!g515) & (g2054) & (g2090) & (!g2095) & (g2119)) + ((g515) & (!g2054) & (!g2090) & (!g2095) & (!g2119)) + ((g515) & (!g2054) & (!g2090) & (g2095) & (!g2119)) + ((g515) & (!g2054) & (!g2090) & (g2095) & (g2119)) + ((g515) & (g2054) & (!g2090) & (!g2095) & (g2119)) + ((g515) & (g2054) & (g2090) & (!g2095) & (!g2119)) + ((g515) & (g2054) & (g2090) & (!g2095) & (g2119)) + ((g515) & (g2054) & (g2090) & (g2095) & (!g2119)) + ((g515) & (g2054) & (g2090) & (g2095) & (g2119)));
	assign g2133 = (((!g553) & (!g604) & (g2056) & (g2089)) + ((!g553) & (g604) & (!g2056) & (g2089)) + ((!g553) & (g604) & (g2056) & (!g2089)) + ((!g553) & (g604) & (g2056) & (g2089)) + ((g553) & (!g604) & (!g2056) & (!g2089)) + ((g553) & (!g604) & (!g2056) & (g2089)) + ((g553) & (!g604) & (g2056) & (!g2089)) + ((g553) & (g604) & (!g2056) & (!g2089)));
	assign g2134 = (((!g2055) & (!g2095) & (!g2119) & (g2133)) + ((!g2055) & (g2095) & (!g2119) & (g2133)) + ((!g2055) & (g2095) & (g2119) & (g2133)) + ((g2055) & (!g2095) & (!g2119) & (!g2133)) + ((g2055) & (!g2095) & (g2119) & (!g2133)) + ((g2055) & (!g2095) & (g2119) & (g2133)) + ((g2055) & (g2095) & (!g2119) & (!g2133)) + ((g2055) & (g2095) & (g2119) & (!g2133)));
	assign g2135 = (((!g604) & (!g2056) & (g2089) & (!g2095) & (!g2119)) + ((!g604) & (!g2056) & (g2089) & (g2095) & (!g2119)) + ((!g604) & (!g2056) & (g2089) & (g2095) & (g2119)) + ((!g604) & (g2056) & (!g2089) & (!g2095) & (!g2119)) + ((!g604) & (g2056) & (!g2089) & (!g2095) & (g2119)) + ((!g604) & (g2056) & (!g2089) & (g2095) & (!g2119)) + ((!g604) & (g2056) & (!g2089) & (g2095) & (g2119)) + ((!g604) & (g2056) & (g2089) & (!g2095) & (g2119)) + ((g604) & (!g2056) & (!g2089) & (!g2095) & (!g2119)) + ((g604) & (!g2056) & (!g2089) & (g2095) & (!g2119)) + ((g604) & (!g2056) & (!g2089) & (g2095) & (g2119)) + ((g604) & (g2056) & (!g2089) & (!g2095) & (g2119)) + ((g604) & (g2056) & (g2089) & (!g2095) & (!g2119)) + ((g604) & (g2056) & (g2089) & (!g2095) & (g2119)) + ((g604) & (g2056) & (g2089) & (g2095) & (!g2119)) + ((g604) & (g2056) & (g2089) & (g2095) & (g2119)));
	assign g2136 = (((!g645) & (!g700) & (g2058) & (g2088)) + ((!g645) & (g700) & (!g2058) & (g2088)) + ((!g645) & (g700) & (g2058) & (!g2088)) + ((!g645) & (g700) & (g2058) & (g2088)) + ((g645) & (!g700) & (!g2058) & (!g2088)) + ((g645) & (!g700) & (!g2058) & (g2088)) + ((g645) & (!g700) & (g2058) & (!g2088)) + ((g645) & (g700) & (!g2058) & (!g2088)));
	assign g2137 = (((!g2057) & (!g2095) & (!g2119) & (g2136)) + ((!g2057) & (g2095) & (!g2119) & (g2136)) + ((!g2057) & (g2095) & (g2119) & (g2136)) + ((g2057) & (!g2095) & (!g2119) & (!g2136)) + ((g2057) & (!g2095) & (g2119) & (!g2136)) + ((g2057) & (!g2095) & (g2119) & (g2136)) + ((g2057) & (g2095) & (!g2119) & (!g2136)) + ((g2057) & (g2095) & (g2119) & (!g2136)));
	assign g2138 = (((!g700) & (!g2058) & (g2088) & (!g2095) & (!g2119)) + ((!g700) & (!g2058) & (g2088) & (g2095) & (!g2119)) + ((!g700) & (!g2058) & (g2088) & (g2095) & (g2119)) + ((!g700) & (g2058) & (!g2088) & (!g2095) & (!g2119)) + ((!g700) & (g2058) & (!g2088) & (!g2095) & (g2119)) + ((!g700) & (g2058) & (!g2088) & (g2095) & (!g2119)) + ((!g700) & (g2058) & (!g2088) & (g2095) & (g2119)) + ((!g700) & (g2058) & (g2088) & (!g2095) & (g2119)) + ((g700) & (!g2058) & (!g2088) & (!g2095) & (!g2119)) + ((g700) & (!g2058) & (!g2088) & (g2095) & (!g2119)) + ((g700) & (!g2058) & (!g2088) & (g2095) & (g2119)) + ((g700) & (g2058) & (!g2088) & (!g2095) & (g2119)) + ((g700) & (g2058) & (g2088) & (!g2095) & (!g2119)) + ((g700) & (g2058) & (g2088) & (!g2095) & (g2119)) + ((g700) & (g2058) & (g2088) & (g2095) & (!g2119)) + ((g700) & (g2058) & (g2088) & (g2095) & (g2119)));
	assign g2139 = (((!g744) & (!g803) & (g2060) & (g2087)) + ((!g744) & (g803) & (!g2060) & (g2087)) + ((!g744) & (g803) & (g2060) & (!g2087)) + ((!g744) & (g803) & (g2060) & (g2087)) + ((g744) & (!g803) & (!g2060) & (!g2087)) + ((g744) & (!g803) & (!g2060) & (g2087)) + ((g744) & (!g803) & (g2060) & (!g2087)) + ((g744) & (g803) & (!g2060) & (!g2087)));
	assign g2140 = (((!g2059) & (!g2095) & (!g2119) & (g2139)) + ((!g2059) & (g2095) & (!g2119) & (g2139)) + ((!g2059) & (g2095) & (g2119) & (g2139)) + ((g2059) & (!g2095) & (!g2119) & (!g2139)) + ((g2059) & (!g2095) & (g2119) & (!g2139)) + ((g2059) & (!g2095) & (g2119) & (g2139)) + ((g2059) & (g2095) & (!g2119) & (!g2139)) + ((g2059) & (g2095) & (g2119) & (!g2139)));
	assign g2141 = (((!g803) & (!g2060) & (g2087) & (!g2095) & (!g2119)) + ((!g803) & (!g2060) & (g2087) & (g2095) & (!g2119)) + ((!g803) & (!g2060) & (g2087) & (g2095) & (g2119)) + ((!g803) & (g2060) & (!g2087) & (!g2095) & (!g2119)) + ((!g803) & (g2060) & (!g2087) & (!g2095) & (g2119)) + ((!g803) & (g2060) & (!g2087) & (g2095) & (!g2119)) + ((!g803) & (g2060) & (!g2087) & (g2095) & (g2119)) + ((!g803) & (g2060) & (g2087) & (!g2095) & (g2119)) + ((g803) & (!g2060) & (!g2087) & (!g2095) & (!g2119)) + ((g803) & (!g2060) & (!g2087) & (g2095) & (!g2119)) + ((g803) & (!g2060) & (!g2087) & (g2095) & (g2119)) + ((g803) & (g2060) & (!g2087) & (!g2095) & (g2119)) + ((g803) & (g2060) & (g2087) & (!g2095) & (!g2119)) + ((g803) & (g2060) & (g2087) & (!g2095) & (g2119)) + ((g803) & (g2060) & (g2087) & (g2095) & (!g2119)) + ((g803) & (g2060) & (g2087) & (g2095) & (g2119)));
	assign g2142 = (((!g851) & (!g914) & (g2062) & (g2086)) + ((!g851) & (g914) & (!g2062) & (g2086)) + ((!g851) & (g914) & (g2062) & (!g2086)) + ((!g851) & (g914) & (g2062) & (g2086)) + ((g851) & (!g914) & (!g2062) & (!g2086)) + ((g851) & (!g914) & (!g2062) & (g2086)) + ((g851) & (!g914) & (g2062) & (!g2086)) + ((g851) & (g914) & (!g2062) & (!g2086)));
	assign g2143 = (((!g2061) & (!g2095) & (!g2119) & (g2142)) + ((!g2061) & (g2095) & (!g2119) & (g2142)) + ((!g2061) & (g2095) & (g2119) & (g2142)) + ((g2061) & (!g2095) & (!g2119) & (!g2142)) + ((g2061) & (!g2095) & (g2119) & (!g2142)) + ((g2061) & (!g2095) & (g2119) & (g2142)) + ((g2061) & (g2095) & (!g2119) & (!g2142)) + ((g2061) & (g2095) & (g2119) & (!g2142)));
	assign g2144 = (((!g914) & (!g2062) & (g2086) & (!g2095) & (!g2119)) + ((!g914) & (!g2062) & (g2086) & (g2095) & (!g2119)) + ((!g914) & (!g2062) & (g2086) & (g2095) & (g2119)) + ((!g914) & (g2062) & (!g2086) & (!g2095) & (!g2119)) + ((!g914) & (g2062) & (!g2086) & (!g2095) & (g2119)) + ((!g914) & (g2062) & (!g2086) & (g2095) & (!g2119)) + ((!g914) & (g2062) & (!g2086) & (g2095) & (g2119)) + ((!g914) & (g2062) & (g2086) & (!g2095) & (g2119)) + ((g914) & (!g2062) & (!g2086) & (!g2095) & (!g2119)) + ((g914) & (!g2062) & (!g2086) & (g2095) & (!g2119)) + ((g914) & (!g2062) & (!g2086) & (g2095) & (g2119)) + ((g914) & (g2062) & (!g2086) & (!g2095) & (g2119)) + ((g914) & (g2062) & (g2086) & (!g2095) & (!g2119)) + ((g914) & (g2062) & (g2086) & (!g2095) & (g2119)) + ((g914) & (g2062) & (g2086) & (g2095) & (!g2119)) + ((g914) & (g2062) & (g2086) & (g2095) & (g2119)));
	assign g2145 = (((!g1032) & (!g1030) & (g2064) & (g2085)) + ((!g1032) & (g1030) & (!g2064) & (g2085)) + ((!g1032) & (g1030) & (g2064) & (!g2085)) + ((!g1032) & (g1030) & (g2064) & (g2085)) + ((g1032) & (!g1030) & (!g2064) & (!g2085)) + ((g1032) & (!g1030) & (!g2064) & (g2085)) + ((g1032) & (!g1030) & (g2064) & (!g2085)) + ((g1032) & (g1030) & (!g2064) & (!g2085)));
	assign g2146 = (((!g2063) & (!g2095) & (!g2119) & (g2145)) + ((!g2063) & (g2095) & (!g2119) & (g2145)) + ((!g2063) & (g2095) & (g2119) & (g2145)) + ((g2063) & (!g2095) & (!g2119) & (!g2145)) + ((g2063) & (!g2095) & (g2119) & (!g2145)) + ((g2063) & (!g2095) & (g2119) & (g2145)) + ((g2063) & (g2095) & (!g2119) & (!g2145)) + ((g2063) & (g2095) & (g2119) & (!g2145)));
	assign g2147 = (((!g1030) & (!g2064) & (g2085) & (!g2095) & (!g2119)) + ((!g1030) & (!g2064) & (g2085) & (g2095) & (!g2119)) + ((!g1030) & (!g2064) & (g2085) & (g2095) & (g2119)) + ((!g1030) & (g2064) & (!g2085) & (!g2095) & (!g2119)) + ((!g1030) & (g2064) & (!g2085) & (!g2095) & (g2119)) + ((!g1030) & (g2064) & (!g2085) & (g2095) & (!g2119)) + ((!g1030) & (g2064) & (!g2085) & (g2095) & (g2119)) + ((!g1030) & (g2064) & (g2085) & (!g2095) & (g2119)) + ((g1030) & (!g2064) & (!g2085) & (!g2095) & (!g2119)) + ((g1030) & (!g2064) & (!g2085) & (g2095) & (!g2119)) + ((g1030) & (!g2064) & (!g2085) & (g2095) & (g2119)) + ((g1030) & (g2064) & (!g2085) & (!g2095) & (g2119)) + ((g1030) & (g2064) & (g2085) & (!g2095) & (!g2119)) + ((g1030) & (g2064) & (g2085) & (!g2095) & (g2119)) + ((g1030) & (g2064) & (g2085) & (g2095) & (!g2119)) + ((g1030) & (g2064) & (g2085) & (g2095) & (g2119)));
	assign g2148 = (((!g1160) & (!g1154) & (g2066) & (g2084)) + ((!g1160) & (g1154) & (!g2066) & (g2084)) + ((!g1160) & (g1154) & (g2066) & (!g2084)) + ((!g1160) & (g1154) & (g2066) & (g2084)) + ((g1160) & (!g1154) & (!g2066) & (!g2084)) + ((g1160) & (!g1154) & (!g2066) & (g2084)) + ((g1160) & (!g1154) & (g2066) & (!g2084)) + ((g1160) & (g1154) & (!g2066) & (!g2084)));
	assign g2149 = (((!g2065) & (!g2095) & (!g2119) & (g2148)) + ((!g2065) & (g2095) & (!g2119) & (g2148)) + ((!g2065) & (g2095) & (g2119) & (g2148)) + ((g2065) & (!g2095) & (!g2119) & (!g2148)) + ((g2065) & (!g2095) & (g2119) & (!g2148)) + ((g2065) & (!g2095) & (g2119) & (g2148)) + ((g2065) & (g2095) & (!g2119) & (!g2148)) + ((g2065) & (g2095) & (g2119) & (!g2148)));
	assign g2150 = (((!g1154) & (!g2066) & (g2084) & (!g2095) & (!g2119)) + ((!g1154) & (!g2066) & (g2084) & (g2095) & (!g2119)) + ((!g1154) & (!g2066) & (g2084) & (g2095) & (g2119)) + ((!g1154) & (g2066) & (!g2084) & (!g2095) & (!g2119)) + ((!g1154) & (g2066) & (!g2084) & (!g2095) & (g2119)) + ((!g1154) & (g2066) & (!g2084) & (g2095) & (!g2119)) + ((!g1154) & (g2066) & (!g2084) & (g2095) & (g2119)) + ((!g1154) & (g2066) & (g2084) & (!g2095) & (g2119)) + ((g1154) & (!g2066) & (!g2084) & (!g2095) & (!g2119)) + ((g1154) & (!g2066) & (!g2084) & (g2095) & (!g2119)) + ((g1154) & (!g2066) & (!g2084) & (g2095) & (g2119)) + ((g1154) & (g2066) & (!g2084) & (!g2095) & (g2119)) + ((g1154) & (g2066) & (g2084) & (!g2095) & (!g2119)) + ((g1154) & (g2066) & (g2084) & (!g2095) & (g2119)) + ((g1154) & (g2066) & (g2084) & (g2095) & (!g2119)) + ((g1154) & (g2066) & (g2084) & (g2095) & (g2119)));
	assign g2151 = (((!g1295) & (!g1285) & (g2068) & (g2083)) + ((!g1295) & (g1285) & (!g2068) & (g2083)) + ((!g1295) & (g1285) & (g2068) & (!g2083)) + ((!g1295) & (g1285) & (g2068) & (g2083)) + ((g1295) & (!g1285) & (!g2068) & (!g2083)) + ((g1295) & (!g1285) & (!g2068) & (g2083)) + ((g1295) & (!g1285) & (g2068) & (!g2083)) + ((g1295) & (g1285) & (!g2068) & (!g2083)));
	assign g2152 = (((!g2067) & (!g2095) & (!g2119) & (g2151)) + ((!g2067) & (g2095) & (!g2119) & (g2151)) + ((!g2067) & (g2095) & (g2119) & (g2151)) + ((g2067) & (!g2095) & (!g2119) & (!g2151)) + ((g2067) & (!g2095) & (g2119) & (!g2151)) + ((g2067) & (!g2095) & (g2119) & (g2151)) + ((g2067) & (g2095) & (!g2119) & (!g2151)) + ((g2067) & (g2095) & (g2119) & (!g2151)));
	assign g2153 = (((!g1285) & (!g2068) & (g2083) & (!g2095) & (!g2119)) + ((!g1285) & (!g2068) & (g2083) & (g2095) & (!g2119)) + ((!g1285) & (!g2068) & (g2083) & (g2095) & (g2119)) + ((!g1285) & (g2068) & (!g2083) & (!g2095) & (!g2119)) + ((!g1285) & (g2068) & (!g2083) & (!g2095) & (g2119)) + ((!g1285) & (g2068) & (!g2083) & (g2095) & (!g2119)) + ((!g1285) & (g2068) & (!g2083) & (g2095) & (g2119)) + ((!g1285) & (g2068) & (g2083) & (!g2095) & (g2119)) + ((g1285) & (!g2068) & (!g2083) & (!g2095) & (!g2119)) + ((g1285) & (!g2068) & (!g2083) & (g2095) & (!g2119)) + ((g1285) & (!g2068) & (!g2083) & (g2095) & (g2119)) + ((g1285) & (g2068) & (!g2083) & (!g2095) & (g2119)) + ((g1285) & (g2068) & (g2083) & (!g2095) & (!g2119)) + ((g1285) & (g2068) & (g2083) & (!g2095) & (g2119)) + ((g1285) & (g2068) & (g2083) & (g2095) & (!g2119)) + ((g1285) & (g2068) & (g2083) & (g2095) & (g2119)));
	assign g2154 = (((!g1437) & (!g1423) & (g2070) & (g2082)) + ((!g1437) & (g1423) & (!g2070) & (g2082)) + ((!g1437) & (g1423) & (g2070) & (!g2082)) + ((!g1437) & (g1423) & (g2070) & (g2082)) + ((g1437) & (!g1423) & (!g2070) & (!g2082)) + ((g1437) & (!g1423) & (!g2070) & (g2082)) + ((g1437) & (!g1423) & (g2070) & (!g2082)) + ((g1437) & (g1423) & (!g2070) & (!g2082)));
	assign g2155 = (((!g2069) & (!g2095) & (!g2119) & (g2154)) + ((!g2069) & (g2095) & (!g2119) & (g2154)) + ((!g2069) & (g2095) & (g2119) & (g2154)) + ((g2069) & (!g2095) & (!g2119) & (!g2154)) + ((g2069) & (!g2095) & (g2119) & (!g2154)) + ((g2069) & (!g2095) & (g2119) & (g2154)) + ((g2069) & (g2095) & (!g2119) & (!g2154)) + ((g2069) & (g2095) & (g2119) & (!g2154)));
	assign g2156 = (((!g1423) & (!g2070) & (g2082) & (!g2095) & (!g2119)) + ((!g1423) & (!g2070) & (g2082) & (g2095) & (!g2119)) + ((!g1423) & (!g2070) & (g2082) & (g2095) & (g2119)) + ((!g1423) & (g2070) & (!g2082) & (!g2095) & (!g2119)) + ((!g1423) & (g2070) & (!g2082) & (!g2095) & (g2119)) + ((!g1423) & (g2070) & (!g2082) & (g2095) & (!g2119)) + ((!g1423) & (g2070) & (!g2082) & (g2095) & (g2119)) + ((!g1423) & (g2070) & (g2082) & (!g2095) & (g2119)) + ((g1423) & (!g2070) & (!g2082) & (!g2095) & (!g2119)) + ((g1423) & (!g2070) & (!g2082) & (g2095) & (!g2119)) + ((g1423) & (!g2070) & (!g2082) & (g2095) & (g2119)) + ((g1423) & (g2070) & (!g2082) & (!g2095) & (g2119)) + ((g1423) & (g2070) & (g2082) & (!g2095) & (!g2119)) + ((g1423) & (g2070) & (g2082) & (!g2095) & (g2119)) + ((g1423) & (g2070) & (g2082) & (g2095) & (!g2119)) + ((g1423) & (g2070) & (g2082) & (g2095) & (g2119)));
	assign g2157 = (((!g1586) & (!g1568) & (g2072) & (g2081)) + ((!g1586) & (g1568) & (!g2072) & (g2081)) + ((!g1586) & (g1568) & (g2072) & (!g2081)) + ((!g1586) & (g1568) & (g2072) & (g2081)) + ((g1586) & (!g1568) & (!g2072) & (!g2081)) + ((g1586) & (!g1568) & (!g2072) & (g2081)) + ((g1586) & (!g1568) & (g2072) & (!g2081)) + ((g1586) & (g1568) & (!g2072) & (!g2081)));
	assign g2158 = (((!g2071) & (!g2095) & (!g2119) & (g2157)) + ((!g2071) & (g2095) & (!g2119) & (g2157)) + ((!g2071) & (g2095) & (g2119) & (g2157)) + ((g2071) & (!g2095) & (!g2119) & (!g2157)) + ((g2071) & (!g2095) & (g2119) & (!g2157)) + ((g2071) & (!g2095) & (g2119) & (g2157)) + ((g2071) & (g2095) & (!g2119) & (!g2157)) + ((g2071) & (g2095) & (g2119) & (!g2157)));
	assign g2159 = (((!g1568) & (!g2072) & (g2081) & (!g2095) & (!g2119)) + ((!g1568) & (!g2072) & (g2081) & (g2095) & (!g2119)) + ((!g1568) & (!g2072) & (g2081) & (g2095) & (g2119)) + ((!g1568) & (g2072) & (!g2081) & (!g2095) & (!g2119)) + ((!g1568) & (g2072) & (!g2081) & (!g2095) & (g2119)) + ((!g1568) & (g2072) & (!g2081) & (g2095) & (!g2119)) + ((!g1568) & (g2072) & (!g2081) & (g2095) & (g2119)) + ((!g1568) & (g2072) & (g2081) & (!g2095) & (g2119)) + ((g1568) & (!g2072) & (!g2081) & (!g2095) & (!g2119)) + ((g1568) & (!g2072) & (!g2081) & (g2095) & (!g2119)) + ((g1568) & (!g2072) & (!g2081) & (g2095) & (g2119)) + ((g1568) & (g2072) & (!g2081) & (!g2095) & (g2119)) + ((g1568) & (g2072) & (g2081) & (!g2095) & (!g2119)) + ((g1568) & (g2072) & (g2081) & (!g2095) & (g2119)) + ((g1568) & (g2072) & (g2081) & (g2095) & (!g2119)) + ((g1568) & (g2072) & (g2081) & (g2095) & (g2119)));
	assign g2160 = (((!g1742) & (!g1720) & (g2074) & (g2080)) + ((!g1742) & (g1720) & (!g2074) & (g2080)) + ((!g1742) & (g1720) & (g2074) & (!g2080)) + ((!g1742) & (g1720) & (g2074) & (g2080)) + ((g1742) & (!g1720) & (!g2074) & (!g2080)) + ((g1742) & (!g1720) & (!g2074) & (g2080)) + ((g1742) & (!g1720) & (g2074) & (!g2080)) + ((g1742) & (g1720) & (!g2074) & (!g2080)));
	assign g2161 = (((!g2073) & (!g2095) & (!g2119) & (g2160)) + ((!g2073) & (g2095) & (!g2119) & (g2160)) + ((!g2073) & (g2095) & (g2119) & (g2160)) + ((g2073) & (!g2095) & (!g2119) & (!g2160)) + ((g2073) & (!g2095) & (g2119) & (!g2160)) + ((g2073) & (!g2095) & (g2119) & (g2160)) + ((g2073) & (g2095) & (!g2119) & (!g2160)) + ((g2073) & (g2095) & (g2119) & (!g2160)));
	assign g2162 = (((!g1720) & (!g2074) & (g2080) & (!g2095) & (!g2119)) + ((!g1720) & (!g2074) & (g2080) & (g2095) & (!g2119)) + ((!g1720) & (!g2074) & (g2080) & (g2095) & (g2119)) + ((!g1720) & (g2074) & (!g2080) & (!g2095) & (!g2119)) + ((!g1720) & (g2074) & (!g2080) & (!g2095) & (g2119)) + ((!g1720) & (g2074) & (!g2080) & (g2095) & (!g2119)) + ((!g1720) & (g2074) & (!g2080) & (g2095) & (g2119)) + ((!g1720) & (g2074) & (g2080) & (!g2095) & (g2119)) + ((g1720) & (!g2074) & (!g2080) & (!g2095) & (!g2119)) + ((g1720) & (!g2074) & (!g2080) & (g2095) & (!g2119)) + ((g1720) & (!g2074) & (!g2080) & (g2095) & (g2119)) + ((g1720) & (g2074) & (!g2080) & (!g2095) & (g2119)) + ((g1720) & (g2074) & (g2080) & (!g2095) & (!g2119)) + ((g1720) & (g2074) & (g2080) & (!g2095) & (g2119)) + ((g1720) & (g2074) & (g2080) & (g2095) & (!g2119)) + ((g1720) & (g2074) & (g2080) & (g2095) & (g2119)));
	assign g2163 = (((!g1905) & (!g1879) & (g2077) & (g2079)) + ((!g1905) & (g1879) & (!g2077) & (g2079)) + ((!g1905) & (g1879) & (g2077) & (!g2079)) + ((!g1905) & (g1879) & (g2077) & (g2079)) + ((g1905) & (!g1879) & (!g2077) & (!g2079)) + ((g1905) & (!g1879) & (!g2077) & (g2079)) + ((g1905) & (!g1879) & (g2077) & (!g2079)) + ((g1905) & (g1879) & (!g2077) & (!g2079)));
	assign g2164 = (((!g2076) & (!g2095) & (!g2119) & (g2163)) + ((!g2076) & (g2095) & (!g2119) & (g2163)) + ((!g2076) & (g2095) & (g2119) & (g2163)) + ((g2076) & (!g2095) & (!g2119) & (!g2163)) + ((g2076) & (!g2095) & (g2119) & (!g2163)) + ((g2076) & (!g2095) & (g2119) & (g2163)) + ((g2076) & (g2095) & (!g2119) & (!g2163)) + ((g2076) & (g2095) & (g2119) & (!g2163)));
	assign g2165 = (((!g1879) & (!g2077) & (g2079) & (!g2095) & (!g2119)) + ((!g1879) & (!g2077) & (g2079) & (g2095) & (!g2119)) + ((!g1879) & (!g2077) & (g2079) & (g2095) & (g2119)) + ((!g1879) & (g2077) & (!g2079) & (!g2095) & (!g2119)) + ((!g1879) & (g2077) & (!g2079) & (!g2095) & (g2119)) + ((!g1879) & (g2077) & (!g2079) & (g2095) & (!g2119)) + ((!g1879) & (g2077) & (!g2079) & (g2095) & (g2119)) + ((!g1879) & (g2077) & (g2079) & (!g2095) & (g2119)) + ((g1879) & (!g2077) & (!g2079) & (!g2095) & (!g2119)) + ((g1879) & (!g2077) & (!g2079) & (g2095) & (!g2119)) + ((g1879) & (!g2077) & (!g2079) & (g2095) & (g2119)) + ((g1879) & (g2077) & (!g2079) & (!g2095) & (g2119)) + ((g1879) & (g2077) & (g2079) & (!g2095) & (!g2119)) + ((g1879) & (g2077) & (g2079) & (!g2095) & (g2119)) + ((g1879) & (g2077) & (g2079) & (g2095) & (!g2119)) + ((g1879) & (g2077) & (g2079) & (g2095) & (g2119)));
	assign g2166 = (((!g2075) & (!ax32x) & (!g2045) & (g2078)) + ((!g2075) & (!ax32x) & (g2045) & (g2078)) + ((!g2075) & (ax32x) & (!g2045) & (!g2078)) + ((!g2075) & (ax32x) & (!g2045) & (g2078)) + ((g2075) & (!ax32x) & (!g2045) & (!g2078)) + ((g2075) & (!ax32x) & (g2045) & (!g2078)) + ((g2075) & (ax32x) & (g2045) & (!g2078)) + ((g2075) & (ax32x) & (g2045) & (g2078)));
	assign g2167 = (((!ax32x) & (!ax33x) & (!g2045) & (!g2095) & (!g2119) & (g2166)) + ((!ax32x) & (!ax33x) & (!g2045) & (!g2095) & (g2119) & (!g2166)) + ((!ax32x) & (!ax33x) & (!g2045) & (!g2095) & (g2119) & (g2166)) + ((!ax32x) & (!ax33x) & (!g2045) & (g2095) & (!g2119) & (g2166)) + ((!ax32x) & (!ax33x) & (!g2045) & (g2095) & (g2119) & (g2166)) + ((!ax32x) & (!ax33x) & (g2045) & (!g2095) & (!g2119) & (!g2166)) + ((!ax32x) & (!ax33x) & (g2045) & (g2095) & (!g2119) & (!g2166)) + ((!ax32x) & (!ax33x) & (g2045) & (g2095) & (g2119) & (!g2166)) + ((!ax32x) & (ax33x) & (!g2045) & (!g2095) & (!g2119) & (!g2166)) + ((!ax32x) & (ax33x) & (!g2045) & (g2095) & (!g2119) & (!g2166)) + ((!ax32x) & (ax33x) & (!g2045) & (g2095) & (g2119) & (!g2166)) + ((!ax32x) & (ax33x) & (g2045) & (!g2095) & (!g2119) & (g2166)) + ((!ax32x) & (ax33x) & (g2045) & (!g2095) & (g2119) & (!g2166)) + ((!ax32x) & (ax33x) & (g2045) & (!g2095) & (g2119) & (g2166)) + ((!ax32x) & (ax33x) & (g2045) & (g2095) & (!g2119) & (g2166)) + ((!ax32x) & (ax33x) & (g2045) & (g2095) & (g2119) & (g2166)) + ((ax32x) & (!ax33x) & (!g2045) & (!g2095) & (!g2119) & (!g2166)) + ((ax32x) & (!ax33x) & (!g2045) & (g2095) & (!g2119) & (!g2166)) + ((ax32x) & (!ax33x) & (!g2045) & (g2095) & (g2119) & (!g2166)) + ((ax32x) & (!ax33x) & (g2045) & (!g2095) & (!g2119) & (!g2166)) + ((ax32x) & (!ax33x) & (g2045) & (g2095) & (!g2119) & (!g2166)) + ((ax32x) & (!ax33x) & (g2045) & (g2095) & (g2119) & (!g2166)) + ((ax32x) & (ax33x) & (!g2045) & (!g2095) & (!g2119) & (g2166)) + ((ax32x) & (ax33x) & (!g2045) & (!g2095) & (g2119) & (!g2166)) + ((ax32x) & (ax33x) & (!g2045) & (!g2095) & (g2119) & (g2166)) + ((ax32x) & (ax33x) & (!g2045) & (g2095) & (!g2119) & (g2166)) + ((ax32x) & (ax33x) & (!g2045) & (g2095) & (g2119) & (g2166)) + ((ax32x) & (ax33x) & (g2045) & (!g2095) & (!g2119) & (g2166)) + ((ax32x) & (ax33x) & (g2045) & (!g2095) & (g2119) & (!g2166)) + ((ax32x) & (ax33x) & (g2045) & (!g2095) & (g2119) & (g2166)) + ((ax32x) & (ax33x) & (g2045) & (g2095) & (!g2119) & (g2166)) + ((ax32x) & (ax33x) & (g2045) & (g2095) & (g2119) & (g2166)));
	assign g2168 = (((!ax32x) & (!g2045) & (!g2078) & (!g2095) & (g2119)) + ((!ax32x) & (!g2045) & (g2078) & (!g2095) & (!g2119)) + ((!ax32x) & (!g2045) & (g2078) & (!g2095) & (g2119)) + ((!ax32x) & (!g2045) & (g2078) & (g2095) & (!g2119)) + ((!ax32x) & (!g2045) & (g2078) & (g2095) & (g2119)) + ((!ax32x) & (g2045) & (g2078) & (!g2095) & (!g2119)) + ((!ax32x) & (g2045) & (g2078) & (g2095) & (!g2119)) + ((!ax32x) & (g2045) & (g2078) & (g2095) & (g2119)) + ((ax32x) & (!g2045) & (!g2078) & (!g2095) & (!g2119)) + ((ax32x) & (!g2045) & (!g2078) & (g2095) & (!g2119)) + ((ax32x) & (!g2045) & (!g2078) & (g2095) & (g2119)) + ((ax32x) & (g2045) & (!g2078) & (!g2095) & (!g2119)) + ((ax32x) & (g2045) & (!g2078) & (!g2095) & (g2119)) + ((ax32x) & (g2045) & (!g2078) & (g2095) & (!g2119)) + ((ax32x) & (g2045) & (!g2078) & (g2095) & (g2119)) + ((ax32x) & (g2045) & (g2078) & (!g2095) & (g2119)));
	assign g2169 = (((!ax28x) & (!ax29x)));
	assign g2170 = (((!g2045) & (!ax30x) & (!ax31x) & (!g2095) & (!g2119) & (!g2169)) + ((!g2045) & (!ax30x) & (!ax31x) & (g2095) & (!g2119) & (!g2169)) + ((!g2045) & (!ax30x) & (!ax31x) & (g2095) & (g2119) & (!g2169)) + ((!g2045) & (!ax30x) & (ax31x) & (!g2095) & (g2119) & (!g2169)) + ((!g2045) & (ax30x) & (ax31x) & (!g2095) & (g2119) & (!g2169)) + ((!g2045) & (ax30x) & (ax31x) & (!g2095) & (g2119) & (g2169)) + ((g2045) & (!ax30x) & (!ax31x) & (!g2095) & (!g2119) & (!g2169)) + ((g2045) & (!ax30x) & (!ax31x) & (!g2095) & (!g2119) & (g2169)) + ((g2045) & (!ax30x) & (!ax31x) & (!g2095) & (g2119) & (!g2169)) + ((g2045) & (!ax30x) & (!ax31x) & (g2095) & (!g2119) & (!g2169)) + ((g2045) & (!ax30x) & (!ax31x) & (g2095) & (!g2119) & (g2169)) + ((g2045) & (!ax30x) & (!ax31x) & (g2095) & (g2119) & (!g2169)) + ((g2045) & (!ax30x) & (!ax31x) & (g2095) & (g2119) & (g2169)) + ((g2045) & (!ax30x) & (ax31x) & (!g2095) & (!g2119) & (!g2169)) + ((g2045) & (!ax30x) & (ax31x) & (!g2095) & (g2119) & (!g2169)) + ((g2045) & (!ax30x) & (ax31x) & (!g2095) & (g2119) & (g2169)) + ((g2045) & (!ax30x) & (ax31x) & (g2095) & (!g2119) & (!g2169)) + ((g2045) & (!ax30x) & (ax31x) & (g2095) & (g2119) & (!g2169)) + ((g2045) & (ax30x) & (!ax31x) & (!g2095) & (g2119) & (!g2169)) + ((g2045) & (ax30x) & (!ax31x) & (!g2095) & (g2119) & (g2169)) + ((g2045) & (ax30x) & (ax31x) & (!g2095) & (!g2119) & (!g2169)) + ((g2045) & (ax30x) & (ax31x) & (!g2095) & (!g2119) & (g2169)) + ((g2045) & (ax30x) & (ax31x) & (!g2095) & (g2119) & (!g2169)) + ((g2045) & (ax30x) & (ax31x) & (!g2095) & (g2119) & (g2169)) + ((g2045) & (ax30x) & (ax31x) & (g2095) & (!g2119) & (!g2169)) + ((g2045) & (ax30x) & (ax31x) & (g2095) & (!g2119) & (g2169)) + ((g2045) & (ax30x) & (ax31x) & (g2095) & (g2119) & (!g2169)) + ((g2045) & (ax30x) & (ax31x) & (g2095) & (g2119) & (g2169)));
	assign g2171 = (((!g1879) & (!g2075) & (g2167) & (g2168) & (g2170)) + ((!g1879) & (g2075) & (g2167) & (!g2168) & (g2170)) + ((!g1879) & (g2075) & (g2167) & (g2168) & (!g2170)) + ((!g1879) & (g2075) & (g2167) & (g2168) & (g2170)) + ((g1879) & (!g2075) & (!g2167) & (g2168) & (g2170)) + ((g1879) & (!g2075) & (g2167) & (!g2168) & (!g2170)) + ((g1879) & (!g2075) & (g2167) & (!g2168) & (g2170)) + ((g1879) & (!g2075) & (g2167) & (g2168) & (!g2170)) + ((g1879) & (!g2075) & (g2167) & (g2168) & (g2170)) + ((g1879) & (g2075) & (!g2167) & (!g2168) & (g2170)) + ((g1879) & (g2075) & (!g2167) & (g2168) & (!g2170)) + ((g1879) & (g2075) & (!g2167) & (g2168) & (g2170)) + ((g1879) & (g2075) & (g2167) & (!g2168) & (!g2170)) + ((g1879) & (g2075) & (g2167) & (!g2168) & (g2170)) + ((g1879) & (g2075) & (g2167) & (g2168) & (!g2170)) + ((g1879) & (g2075) & (g2167) & (g2168) & (g2170)));
	assign g2172 = (((!g1720) & (!g1905) & (g2164) & (g2165) & (g2171)) + ((!g1720) & (g1905) & (g2164) & (!g2165) & (g2171)) + ((!g1720) & (g1905) & (g2164) & (g2165) & (!g2171)) + ((!g1720) & (g1905) & (g2164) & (g2165) & (g2171)) + ((g1720) & (!g1905) & (!g2164) & (g2165) & (g2171)) + ((g1720) & (!g1905) & (g2164) & (!g2165) & (!g2171)) + ((g1720) & (!g1905) & (g2164) & (!g2165) & (g2171)) + ((g1720) & (!g1905) & (g2164) & (g2165) & (!g2171)) + ((g1720) & (!g1905) & (g2164) & (g2165) & (g2171)) + ((g1720) & (g1905) & (!g2164) & (!g2165) & (g2171)) + ((g1720) & (g1905) & (!g2164) & (g2165) & (!g2171)) + ((g1720) & (g1905) & (!g2164) & (g2165) & (g2171)) + ((g1720) & (g1905) & (g2164) & (!g2165) & (!g2171)) + ((g1720) & (g1905) & (g2164) & (!g2165) & (g2171)) + ((g1720) & (g1905) & (g2164) & (g2165) & (!g2171)) + ((g1720) & (g1905) & (g2164) & (g2165) & (g2171)));
	assign g2173 = (((!g1568) & (!g1742) & (g2161) & (g2162) & (g2172)) + ((!g1568) & (g1742) & (g2161) & (!g2162) & (g2172)) + ((!g1568) & (g1742) & (g2161) & (g2162) & (!g2172)) + ((!g1568) & (g1742) & (g2161) & (g2162) & (g2172)) + ((g1568) & (!g1742) & (!g2161) & (g2162) & (g2172)) + ((g1568) & (!g1742) & (g2161) & (!g2162) & (!g2172)) + ((g1568) & (!g1742) & (g2161) & (!g2162) & (g2172)) + ((g1568) & (!g1742) & (g2161) & (g2162) & (!g2172)) + ((g1568) & (!g1742) & (g2161) & (g2162) & (g2172)) + ((g1568) & (g1742) & (!g2161) & (!g2162) & (g2172)) + ((g1568) & (g1742) & (!g2161) & (g2162) & (!g2172)) + ((g1568) & (g1742) & (!g2161) & (g2162) & (g2172)) + ((g1568) & (g1742) & (g2161) & (!g2162) & (!g2172)) + ((g1568) & (g1742) & (g2161) & (!g2162) & (g2172)) + ((g1568) & (g1742) & (g2161) & (g2162) & (!g2172)) + ((g1568) & (g1742) & (g2161) & (g2162) & (g2172)));
	assign g2174 = (((!g1423) & (!g1586) & (g2158) & (g2159) & (g2173)) + ((!g1423) & (g1586) & (g2158) & (!g2159) & (g2173)) + ((!g1423) & (g1586) & (g2158) & (g2159) & (!g2173)) + ((!g1423) & (g1586) & (g2158) & (g2159) & (g2173)) + ((g1423) & (!g1586) & (!g2158) & (g2159) & (g2173)) + ((g1423) & (!g1586) & (g2158) & (!g2159) & (!g2173)) + ((g1423) & (!g1586) & (g2158) & (!g2159) & (g2173)) + ((g1423) & (!g1586) & (g2158) & (g2159) & (!g2173)) + ((g1423) & (!g1586) & (g2158) & (g2159) & (g2173)) + ((g1423) & (g1586) & (!g2158) & (!g2159) & (g2173)) + ((g1423) & (g1586) & (!g2158) & (g2159) & (!g2173)) + ((g1423) & (g1586) & (!g2158) & (g2159) & (g2173)) + ((g1423) & (g1586) & (g2158) & (!g2159) & (!g2173)) + ((g1423) & (g1586) & (g2158) & (!g2159) & (g2173)) + ((g1423) & (g1586) & (g2158) & (g2159) & (!g2173)) + ((g1423) & (g1586) & (g2158) & (g2159) & (g2173)));
	assign g2175 = (((!g1285) & (!g1437) & (g2155) & (g2156) & (g2174)) + ((!g1285) & (g1437) & (g2155) & (!g2156) & (g2174)) + ((!g1285) & (g1437) & (g2155) & (g2156) & (!g2174)) + ((!g1285) & (g1437) & (g2155) & (g2156) & (g2174)) + ((g1285) & (!g1437) & (!g2155) & (g2156) & (g2174)) + ((g1285) & (!g1437) & (g2155) & (!g2156) & (!g2174)) + ((g1285) & (!g1437) & (g2155) & (!g2156) & (g2174)) + ((g1285) & (!g1437) & (g2155) & (g2156) & (!g2174)) + ((g1285) & (!g1437) & (g2155) & (g2156) & (g2174)) + ((g1285) & (g1437) & (!g2155) & (!g2156) & (g2174)) + ((g1285) & (g1437) & (!g2155) & (g2156) & (!g2174)) + ((g1285) & (g1437) & (!g2155) & (g2156) & (g2174)) + ((g1285) & (g1437) & (g2155) & (!g2156) & (!g2174)) + ((g1285) & (g1437) & (g2155) & (!g2156) & (g2174)) + ((g1285) & (g1437) & (g2155) & (g2156) & (!g2174)) + ((g1285) & (g1437) & (g2155) & (g2156) & (g2174)));
	assign g2176 = (((!g1154) & (!g1295) & (g2152) & (g2153) & (g2175)) + ((!g1154) & (g1295) & (g2152) & (!g2153) & (g2175)) + ((!g1154) & (g1295) & (g2152) & (g2153) & (!g2175)) + ((!g1154) & (g1295) & (g2152) & (g2153) & (g2175)) + ((g1154) & (!g1295) & (!g2152) & (g2153) & (g2175)) + ((g1154) & (!g1295) & (g2152) & (!g2153) & (!g2175)) + ((g1154) & (!g1295) & (g2152) & (!g2153) & (g2175)) + ((g1154) & (!g1295) & (g2152) & (g2153) & (!g2175)) + ((g1154) & (!g1295) & (g2152) & (g2153) & (g2175)) + ((g1154) & (g1295) & (!g2152) & (!g2153) & (g2175)) + ((g1154) & (g1295) & (!g2152) & (g2153) & (!g2175)) + ((g1154) & (g1295) & (!g2152) & (g2153) & (g2175)) + ((g1154) & (g1295) & (g2152) & (!g2153) & (!g2175)) + ((g1154) & (g1295) & (g2152) & (!g2153) & (g2175)) + ((g1154) & (g1295) & (g2152) & (g2153) & (!g2175)) + ((g1154) & (g1295) & (g2152) & (g2153) & (g2175)));
	assign g2177 = (((!g1030) & (!g1160) & (g2149) & (g2150) & (g2176)) + ((!g1030) & (g1160) & (g2149) & (!g2150) & (g2176)) + ((!g1030) & (g1160) & (g2149) & (g2150) & (!g2176)) + ((!g1030) & (g1160) & (g2149) & (g2150) & (g2176)) + ((g1030) & (!g1160) & (!g2149) & (g2150) & (g2176)) + ((g1030) & (!g1160) & (g2149) & (!g2150) & (!g2176)) + ((g1030) & (!g1160) & (g2149) & (!g2150) & (g2176)) + ((g1030) & (!g1160) & (g2149) & (g2150) & (!g2176)) + ((g1030) & (!g1160) & (g2149) & (g2150) & (g2176)) + ((g1030) & (g1160) & (!g2149) & (!g2150) & (g2176)) + ((g1030) & (g1160) & (!g2149) & (g2150) & (!g2176)) + ((g1030) & (g1160) & (!g2149) & (g2150) & (g2176)) + ((g1030) & (g1160) & (g2149) & (!g2150) & (!g2176)) + ((g1030) & (g1160) & (g2149) & (!g2150) & (g2176)) + ((g1030) & (g1160) & (g2149) & (g2150) & (!g2176)) + ((g1030) & (g1160) & (g2149) & (g2150) & (g2176)));
	assign g2178 = (((!g914) & (!g1032) & (g2146) & (g2147) & (g2177)) + ((!g914) & (g1032) & (g2146) & (!g2147) & (g2177)) + ((!g914) & (g1032) & (g2146) & (g2147) & (!g2177)) + ((!g914) & (g1032) & (g2146) & (g2147) & (g2177)) + ((g914) & (!g1032) & (!g2146) & (g2147) & (g2177)) + ((g914) & (!g1032) & (g2146) & (!g2147) & (!g2177)) + ((g914) & (!g1032) & (g2146) & (!g2147) & (g2177)) + ((g914) & (!g1032) & (g2146) & (g2147) & (!g2177)) + ((g914) & (!g1032) & (g2146) & (g2147) & (g2177)) + ((g914) & (g1032) & (!g2146) & (!g2147) & (g2177)) + ((g914) & (g1032) & (!g2146) & (g2147) & (!g2177)) + ((g914) & (g1032) & (!g2146) & (g2147) & (g2177)) + ((g914) & (g1032) & (g2146) & (!g2147) & (!g2177)) + ((g914) & (g1032) & (g2146) & (!g2147) & (g2177)) + ((g914) & (g1032) & (g2146) & (g2147) & (!g2177)) + ((g914) & (g1032) & (g2146) & (g2147) & (g2177)));
	assign g2179 = (((!g803) & (!g851) & (g2143) & (g2144) & (g2178)) + ((!g803) & (g851) & (g2143) & (!g2144) & (g2178)) + ((!g803) & (g851) & (g2143) & (g2144) & (!g2178)) + ((!g803) & (g851) & (g2143) & (g2144) & (g2178)) + ((g803) & (!g851) & (!g2143) & (g2144) & (g2178)) + ((g803) & (!g851) & (g2143) & (!g2144) & (!g2178)) + ((g803) & (!g851) & (g2143) & (!g2144) & (g2178)) + ((g803) & (!g851) & (g2143) & (g2144) & (!g2178)) + ((g803) & (!g851) & (g2143) & (g2144) & (g2178)) + ((g803) & (g851) & (!g2143) & (!g2144) & (g2178)) + ((g803) & (g851) & (!g2143) & (g2144) & (!g2178)) + ((g803) & (g851) & (!g2143) & (g2144) & (g2178)) + ((g803) & (g851) & (g2143) & (!g2144) & (!g2178)) + ((g803) & (g851) & (g2143) & (!g2144) & (g2178)) + ((g803) & (g851) & (g2143) & (g2144) & (!g2178)) + ((g803) & (g851) & (g2143) & (g2144) & (g2178)));
	assign g2180 = (((!g700) & (!g744) & (g2140) & (g2141) & (g2179)) + ((!g700) & (g744) & (g2140) & (!g2141) & (g2179)) + ((!g700) & (g744) & (g2140) & (g2141) & (!g2179)) + ((!g700) & (g744) & (g2140) & (g2141) & (g2179)) + ((g700) & (!g744) & (!g2140) & (g2141) & (g2179)) + ((g700) & (!g744) & (g2140) & (!g2141) & (!g2179)) + ((g700) & (!g744) & (g2140) & (!g2141) & (g2179)) + ((g700) & (!g744) & (g2140) & (g2141) & (!g2179)) + ((g700) & (!g744) & (g2140) & (g2141) & (g2179)) + ((g700) & (g744) & (!g2140) & (!g2141) & (g2179)) + ((g700) & (g744) & (!g2140) & (g2141) & (!g2179)) + ((g700) & (g744) & (!g2140) & (g2141) & (g2179)) + ((g700) & (g744) & (g2140) & (!g2141) & (!g2179)) + ((g700) & (g744) & (g2140) & (!g2141) & (g2179)) + ((g700) & (g744) & (g2140) & (g2141) & (!g2179)) + ((g700) & (g744) & (g2140) & (g2141) & (g2179)));
	assign g2181 = (((!g604) & (!g645) & (g2137) & (g2138) & (g2180)) + ((!g604) & (g645) & (g2137) & (!g2138) & (g2180)) + ((!g604) & (g645) & (g2137) & (g2138) & (!g2180)) + ((!g604) & (g645) & (g2137) & (g2138) & (g2180)) + ((g604) & (!g645) & (!g2137) & (g2138) & (g2180)) + ((g604) & (!g645) & (g2137) & (!g2138) & (!g2180)) + ((g604) & (!g645) & (g2137) & (!g2138) & (g2180)) + ((g604) & (!g645) & (g2137) & (g2138) & (!g2180)) + ((g604) & (!g645) & (g2137) & (g2138) & (g2180)) + ((g604) & (g645) & (!g2137) & (!g2138) & (g2180)) + ((g604) & (g645) & (!g2137) & (g2138) & (!g2180)) + ((g604) & (g645) & (!g2137) & (g2138) & (g2180)) + ((g604) & (g645) & (g2137) & (!g2138) & (!g2180)) + ((g604) & (g645) & (g2137) & (!g2138) & (g2180)) + ((g604) & (g645) & (g2137) & (g2138) & (!g2180)) + ((g604) & (g645) & (g2137) & (g2138) & (g2180)));
	assign g2182 = (((!g515) & (!g553) & (g2134) & (g2135) & (g2181)) + ((!g515) & (g553) & (g2134) & (!g2135) & (g2181)) + ((!g515) & (g553) & (g2134) & (g2135) & (!g2181)) + ((!g515) & (g553) & (g2134) & (g2135) & (g2181)) + ((g515) & (!g553) & (!g2134) & (g2135) & (g2181)) + ((g515) & (!g553) & (g2134) & (!g2135) & (!g2181)) + ((g515) & (!g553) & (g2134) & (!g2135) & (g2181)) + ((g515) & (!g553) & (g2134) & (g2135) & (!g2181)) + ((g515) & (!g553) & (g2134) & (g2135) & (g2181)) + ((g515) & (g553) & (!g2134) & (!g2135) & (g2181)) + ((g515) & (g553) & (!g2134) & (g2135) & (!g2181)) + ((g515) & (g553) & (!g2134) & (g2135) & (g2181)) + ((g515) & (g553) & (g2134) & (!g2135) & (!g2181)) + ((g515) & (g553) & (g2134) & (!g2135) & (g2181)) + ((g515) & (g553) & (g2134) & (g2135) & (!g2181)) + ((g515) & (g553) & (g2134) & (g2135) & (g2181)));
	assign g2183 = (((!g433) & (!g468) & (g2131) & (g2132) & (g2182)) + ((!g433) & (g468) & (g2131) & (!g2132) & (g2182)) + ((!g433) & (g468) & (g2131) & (g2132) & (!g2182)) + ((!g433) & (g468) & (g2131) & (g2132) & (g2182)) + ((g433) & (!g468) & (!g2131) & (g2132) & (g2182)) + ((g433) & (!g468) & (g2131) & (!g2132) & (!g2182)) + ((g433) & (!g468) & (g2131) & (!g2132) & (g2182)) + ((g433) & (!g468) & (g2131) & (g2132) & (!g2182)) + ((g433) & (!g468) & (g2131) & (g2132) & (g2182)) + ((g433) & (g468) & (!g2131) & (!g2132) & (g2182)) + ((g433) & (g468) & (!g2131) & (g2132) & (!g2182)) + ((g433) & (g468) & (!g2131) & (g2132) & (g2182)) + ((g433) & (g468) & (g2131) & (!g2132) & (!g2182)) + ((g433) & (g468) & (g2131) & (!g2132) & (g2182)) + ((g433) & (g468) & (g2131) & (g2132) & (!g2182)) + ((g433) & (g468) & (g2131) & (g2132) & (g2182)));
	assign g2184 = (((!g358) & (!g390) & (g2128) & (g2129) & (g2183)) + ((!g358) & (g390) & (g2128) & (!g2129) & (g2183)) + ((!g358) & (g390) & (g2128) & (g2129) & (!g2183)) + ((!g358) & (g390) & (g2128) & (g2129) & (g2183)) + ((g358) & (!g390) & (!g2128) & (g2129) & (g2183)) + ((g358) & (!g390) & (g2128) & (!g2129) & (!g2183)) + ((g358) & (!g390) & (g2128) & (!g2129) & (g2183)) + ((g358) & (!g390) & (g2128) & (g2129) & (!g2183)) + ((g358) & (!g390) & (g2128) & (g2129) & (g2183)) + ((g358) & (g390) & (!g2128) & (!g2129) & (g2183)) + ((g358) & (g390) & (!g2128) & (g2129) & (!g2183)) + ((g358) & (g390) & (!g2128) & (g2129) & (g2183)) + ((g358) & (g390) & (g2128) & (!g2129) & (!g2183)) + ((g358) & (g390) & (g2128) & (!g2129) & (g2183)) + ((g358) & (g390) & (g2128) & (g2129) & (!g2183)) + ((g358) & (g390) & (g2128) & (g2129) & (g2183)));
	assign g2185 = (((!g290) & (!g319) & (g2125) & (g2126) & (g2184)) + ((!g290) & (g319) & (g2125) & (!g2126) & (g2184)) + ((!g290) & (g319) & (g2125) & (g2126) & (!g2184)) + ((!g290) & (g319) & (g2125) & (g2126) & (g2184)) + ((g290) & (!g319) & (!g2125) & (g2126) & (g2184)) + ((g290) & (!g319) & (g2125) & (!g2126) & (!g2184)) + ((g290) & (!g319) & (g2125) & (!g2126) & (g2184)) + ((g290) & (!g319) & (g2125) & (g2126) & (!g2184)) + ((g290) & (!g319) & (g2125) & (g2126) & (g2184)) + ((g290) & (g319) & (!g2125) & (!g2126) & (g2184)) + ((g290) & (g319) & (!g2125) & (g2126) & (!g2184)) + ((g290) & (g319) & (!g2125) & (g2126) & (g2184)) + ((g290) & (g319) & (g2125) & (!g2126) & (!g2184)) + ((g290) & (g319) & (g2125) & (!g2126) & (g2184)) + ((g290) & (g319) & (g2125) & (g2126) & (!g2184)) + ((g290) & (g319) & (g2125) & (g2126) & (g2184)));
	assign g2186 = (((!g229) & (!g255) & (g2122) & (g2123) & (g2185)) + ((!g229) & (g255) & (g2122) & (!g2123) & (g2185)) + ((!g229) & (g255) & (g2122) & (g2123) & (!g2185)) + ((!g229) & (g255) & (g2122) & (g2123) & (g2185)) + ((g229) & (!g255) & (!g2122) & (g2123) & (g2185)) + ((g229) & (!g255) & (g2122) & (!g2123) & (!g2185)) + ((g229) & (!g255) & (g2122) & (!g2123) & (g2185)) + ((g229) & (!g255) & (g2122) & (g2123) & (!g2185)) + ((g229) & (!g255) & (g2122) & (g2123) & (g2185)) + ((g229) & (g255) & (!g2122) & (!g2123) & (g2185)) + ((g229) & (g255) & (!g2122) & (g2123) & (!g2185)) + ((g229) & (g255) & (!g2122) & (g2123) & (g2185)) + ((g229) & (g255) & (g2122) & (!g2123) & (!g2185)) + ((g229) & (g255) & (g2122) & (!g2123) & (g2185)) + ((g229) & (g255) & (g2122) & (g2123) & (!g2185)) + ((g229) & (g255) & (g2122) & (g2123) & (g2185)));
	assign g2187 = (((!g4) & (!g2116) & (!g2117) & (!g2095) & (!g2119)) + ((!g4) & (!g2116) & (!g2117) & (g2095) & (!g2119)) + ((!g4) & (!g2116) & (!g2117) & (g2095) & (g2119)) + ((!g4) & (!g2116) & (g2117) & (!g2095) & (g2119)) + ((!g4) & (g2116) & (g2117) & (!g2095) & (!g2119)) + ((!g4) & (g2116) & (g2117) & (!g2095) & (g2119)) + ((!g4) & (g2116) & (g2117) & (g2095) & (!g2119)) + ((!g4) & (g2116) & (g2117) & (g2095) & (g2119)) + ((g4) & (!g2116) & (g2117) & (!g2095) & (!g2119)) + ((g4) & (!g2116) & (g2117) & (!g2095) & (g2119)) + ((g4) & (!g2116) & (g2117) & (g2095) & (!g2119)) + ((g4) & (!g2116) & (g2117) & (g2095) & (g2119)) + ((g4) & (g2116) & (!g2117) & (!g2095) & (!g2119)) + ((g4) & (g2116) & (!g2117) & (g2095) & (!g2119)) + ((g4) & (g2116) & (!g2117) & (g2095) & (g2119)) + ((g4) & (g2116) & (g2117) & (!g2095) & (g2119)));
	assign g2188 = (((!g8) & (!g2098) & (g2115) & (!g2095) & (!g2119)) + ((!g8) & (!g2098) & (g2115) & (g2095) & (!g2119)) + ((!g8) & (!g2098) & (g2115) & (g2095) & (g2119)) + ((!g8) & (g2098) & (!g2115) & (!g2095) & (!g2119)) + ((!g8) & (g2098) & (!g2115) & (!g2095) & (g2119)) + ((!g8) & (g2098) & (!g2115) & (g2095) & (!g2119)) + ((!g8) & (g2098) & (!g2115) & (g2095) & (g2119)) + ((!g8) & (g2098) & (g2115) & (!g2095) & (g2119)) + ((g8) & (!g2098) & (!g2115) & (!g2095) & (!g2119)) + ((g8) & (!g2098) & (!g2115) & (g2095) & (!g2119)) + ((g8) & (!g2098) & (!g2115) & (g2095) & (g2119)) + ((g8) & (g2098) & (!g2115) & (!g2095) & (g2119)) + ((g8) & (g2098) & (g2115) & (!g2095) & (!g2119)) + ((g8) & (g2098) & (g2115) & (!g2095) & (g2119)) + ((g8) & (g2098) & (g2115) & (g2095) & (!g2119)) + ((g8) & (g2098) & (g2115) & (g2095) & (g2119)));
	assign g2189 = (((!g18) & (!g27) & (g2100) & (g2114)) + ((!g18) & (g27) & (!g2100) & (g2114)) + ((!g18) & (g27) & (g2100) & (!g2114)) + ((!g18) & (g27) & (g2100) & (g2114)) + ((g18) & (!g27) & (!g2100) & (!g2114)) + ((g18) & (!g27) & (!g2100) & (g2114)) + ((g18) & (!g27) & (g2100) & (!g2114)) + ((g18) & (g27) & (!g2100) & (!g2114)));
	assign g2190 = (((!g2099) & (!g2095) & (!g2119) & (g2189)) + ((!g2099) & (g2095) & (!g2119) & (g2189)) + ((!g2099) & (g2095) & (g2119) & (g2189)) + ((g2099) & (!g2095) & (!g2119) & (!g2189)) + ((g2099) & (!g2095) & (g2119) & (!g2189)) + ((g2099) & (!g2095) & (g2119) & (g2189)) + ((g2099) & (g2095) & (!g2119) & (!g2189)) + ((g2099) & (g2095) & (g2119) & (!g2189)));
	assign g2191 = (((!g27) & (!g2100) & (g2114) & (!g2095) & (!g2119)) + ((!g27) & (!g2100) & (g2114) & (g2095) & (!g2119)) + ((!g27) & (!g2100) & (g2114) & (g2095) & (g2119)) + ((!g27) & (g2100) & (!g2114) & (!g2095) & (!g2119)) + ((!g27) & (g2100) & (!g2114) & (!g2095) & (g2119)) + ((!g27) & (g2100) & (!g2114) & (g2095) & (!g2119)) + ((!g27) & (g2100) & (!g2114) & (g2095) & (g2119)) + ((!g27) & (g2100) & (g2114) & (!g2095) & (g2119)) + ((g27) & (!g2100) & (!g2114) & (!g2095) & (!g2119)) + ((g27) & (!g2100) & (!g2114) & (g2095) & (!g2119)) + ((g27) & (!g2100) & (!g2114) & (g2095) & (g2119)) + ((g27) & (g2100) & (!g2114) & (!g2095) & (g2119)) + ((g27) & (g2100) & (g2114) & (!g2095) & (!g2119)) + ((g27) & (g2100) & (g2114) & (!g2095) & (g2119)) + ((g27) & (g2100) & (g2114) & (g2095) & (!g2119)) + ((g27) & (g2100) & (g2114) & (g2095) & (g2119)));
	assign g2192 = (((!g39) & (!g54) & (g2102) & (g2113)) + ((!g39) & (g54) & (!g2102) & (g2113)) + ((!g39) & (g54) & (g2102) & (!g2113)) + ((!g39) & (g54) & (g2102) & (g2113)) + ((g39) & (!g54) & (!g2102) & (!g2113)) + ((g39) & (!g54) & (!g2102) & (g2113)) + ((g39) & (!g54) & (g2102) & (!g2113)) + ((g39) & (g54) & (!g2102) & (!g2113)));
	assign g2193 = (((!g2101) & (!g2095) & (!g2119) & (g2192)) + ((!g2101) & (g2095) & (!g2119) & (g2192)) + ((!g2101) & (g2095) & (g2119) & (g2192)) + ((g2101) & (!g2095) & (!g2119) & (!g2192)) + ((g2101) & (!g2095) & (g2119) & (!g2192)) + ((g2101) & (!g2095) & (g2119) & (g2192)) + ((g2101) & (g2095) & (!g2119) & (!g2192)) + ((g2101) & (g2095) & (g2119) & (!g2192)));
	assign g2194 = (((!g54) & (!g2102) & (g2113) & (!g2095) & (!g2119)) + ((!g54) & (!g2102) & (g2113) & (g2095) & (!g2119)) + ((!g54) & (!g2102) & (g2113) & (g2095) & (g2119)) + ((!g54) & (g2102) & (!g2113) & (!g2095) & (!g2119)) + ((!g54) & (g2102) & (!g2113) & (!g2095) & (g2119)) + ((!g54) & (g2102) & (!g2113) & (g2095) & (!g2119)) + ((!g54) & (g2102) & (!g2113) & (g2095) & (g2119)) + ((!g54) & (g2102) & (g2113) & (!g2095) & (g2119)) + ((g54) & (!g2102) & (!g2113) & (!g2095) & (!g2119)) + ((g54) & (!g2102) & (!g2113) & (g2095) & (!g2119)) + ((g54) & (!g2102) & (!g2113) & (g2095) & (g2119)) + ((g54) & (g2102) & (!g2113) & (!g2095) & (g2119)) + ((g54) & (g2102) & (g2113) & (!g2095) & (!g2119)) + ((g54) & (g2102) & (g2113) & (!g2095) & (g2119)) + ((g54) & (g2102) & (g2113) & (g2095) & (!g2119)) + ((g54) & (g2102) & (g2113) & (g2095) & (g2119)));
	assign g2195 = (((!g68) & (!g87) & (g2104) & (g2112)) + ((!g68) & (g87) & (!g2104) & (g2112)) + ((!g68) & (g87) & (g2104) & (!g2112)) + ((!g68) & (g87) & (g2104) & (g2112)) + ((g68) & (!g87) & (!g2104) & (!g2112)) + ((g68) & (!g87) & (!g2104) & (g2112)) + ((g68) & (!g87) & (g2104) & (!g2112)) + ((g68) & (g87) & (!g2104) & (!g2112)));
	assign g2196 = (((!g2103) & (!g2095) & (!g2119) & (g2195)) + ((!g2103) & (g2095) & (!g2119) & (g2195)) + ((!g2103) & (g2095) & (g2119) & (g2195)) + ((g2103) & (!g2095) & (!g2119) & (!g2195)) + ((g2103) & (!g2095) & (g2119) & (!g2195)) + ((g2103) & (!g2095) & (g2119) & (g2195)) + ((g2103) & (g2095) & (!g2119) & (!g2195)) + ((g2103) & (g2095) & (g2119) & (!g2195)));
	assign g2197 = (((!g87) & (!g2104) & (g2112) & (!g2095) & (!g2119)) + ((!g87) & (!g2104) & (g2112) & (g2095) & (!g2119)) + ((!g87) & (!g2104) & (g2112) & (g2095) & (g2119)) + ((!g87) & (g2104) & (!g2112) & (!g2095) & (!g2119)) + ((!g87) & (g2104) & (!g2112) & (!g2095) & (g2119)) + ((!g87) & (g2104) & (!g2112) & (g2095) & (!g2119)) + ((!g87) & (g2104) & (!g2112) & (g2095) & (g2119)) + ((!g87) & (g2104) & (g2112) & (!g2095) & (g2119)) + ((g87) & (!g2104) & (!g2112) & (!g2095) & (!g2119)) + ((g87) & (!g2104) & (!g2112) & (g2095) & (!g2119)) + ((g87) & (!g2104) & (!g2112) & (g2095) & (g2119)) + ((g87) & (g2104) & (!g2112) & (!g2095) & (g2119)) + ((g87) & (g2104) & (g2112) & (!g2095) & (!g2119)) + ((g87) & (g2104) & (g2112) & (!g2095) & (g2119)) + ((g87) & (g2104) & (g2112) & (g2095) & (!g2119)) + ((g87) & (g2104) & (g2112) & (g2095) & (g2119)));
	assign g2198 = (((!g104) & (!g127) & (g2106) & (g2111)) + ((!g104) & (g127) & (!g2106) & (g2111)) + ((!g104) & (g127) & (g2106) & (!g2111)) + ((!g104) & (g127) & (g2106) & (g2111)) + ((g104) & (!g127) & (!g2106) & (!g2111)) + ((g104) & (!g127) & (!g2106) & (g2111)) + ((g104) & (!g127) & (g2106) & (!g2111)) + ((g104) & (g127) & (!g2106) & (!g2111)));
	assign g2199 = (((!g2105) & (!g2095) & (!g2119) & (g2198)) + ((!g2105) & (g2095) & (!g2119) & (g2198)) + ((!g2105) & (g2095) & (g2119) & (g2198)) + ((g2105) & (!g2095) & (!g2119) & (!g2198)) + ((g2105) & (!g2095) & (g2119) & (!g2198)) + ((g2105) & (!g2095) & (g2119) & (g2198)) + ((g2105) & (g2095) & (!g2119) & (!g2198)) + ((g2105) & (g2095) & (g2119) & (!g2198)));
	assign g2200 = (((!g127) & (!g2106) & (g2111) & (!g2095) & (!g2119)) + ((!g127) & (!g2106) & (g2111) & (g2095) & (!g2119)) + ((!g127) & (!g2106) & (g2111) & (g2095) & (g2119)) + ((!g127) & (g2106) & (!g2111) & (!g2095) & (!g2119)) + ((!g127) & (g2106) & (!g2111) & (!g2095) & (g2119)) + ((!g127) & (g2106) & (!g2111) & (g2095) & (!g2119)) + ((!g127) & (g2106) & (!g2111) & (g2095) & (g2119)) + ((!g127) & (g2106) & (g2111) & (!g2095) & (g2119)) + ((g127) & (!g2106) & (!g2111) & (!g2095) & (!g2119)) + ((g127) & (!g2106) & (!g2111) & (g2095) & (!g2119)) + ((g127) & (!g2106) & (!g2111) & (g2095) & (g2119)) + ((g127) & (g2106) & (!g2111) & (!g2095) & (g2119)) + ((g127) & (g2106) & (g2111) & (!g2095) & (!g2119)) + ((g127) & (g2106) & (g2111) & (!g2095) & (g2119)) + ((g127) & (g2106) & (g2111) & (g2095) & (!g2119)) + ((g127) & (g2106) & (g2111) & (g2095) & (g2119)));
	assign g2201 = (((!g147) & (!g174) & (g2108) & (g2110)) + ((!g147) & (g174) & (!g2108) & (g2110)) + ((!g147) & (g174) & (g2108) & (!g2110)) + ((!g147) & (g174) & (g2108) & (g2110)) + ((g147) & (!g174) & (!g2108) & (!g2110)) + ((g147) & (!g174) & (!g2108) & (g2110)) + ((g147) & (!g174) & (g2108) & (!g2110)) + ((g147) & (g174) & (!g2108) & (!g2110)));
	assign g2202 = (((!g2107) & (!g2095) & (!g2119) & (g2201)) + ((!g2107) & (g2095) & (!g2119) & (g2201)) + ((!g2107) & (g2095) & (g2119) & (g2201)) + ((g2107) & (!g2095) & (!g2119) & (!g2201)) + ((g2107) & (!g2095) & (g2119) & (!g2201)) + ((g2107) & (!g2095) & (g2119) & (g2201)) + ((g2107) & (g2095) & (!g2119) & (!g2201)) + ((g2107) & (g2095) & (g2119) & (!g2201)));
	assign g2203 = (((!g174) & (!g2108) & (g2110) & (!g2095) & (!g2119)) + ((!g174) & (!g2108) & (g2110) & (g2095) & (!g2119)) + ((!g174) & (!g2108) & (g2110) & (g2095) & (g2119)) + ((!g174) & (g2108) & (!g2110) & (!g2095) & (!g2119)) + ((!g174) & (g2108) & (!g2110) & (!g2095) & (g2119)) + ((!g174) & (g2108) & (!g2110) & (g2095) & (!g2119)) + ((!g174) & (g2108) & (!g2110) & (g2095) & (g2119)) + ((!g174) & (g2108) & (g2110) & (!g2095) & (g2119)) + ((g174) & (!g2108) & (!g2110) & (!g2095) & (!g2119)) + ((g174) & (!g2108) & (!g2110) & (g2095) & (!g2119)) + ((g174) & (!g2108) & (!g2110) & (g2095) & (g2119)) + ((g174) & (g2108) & (!g2110) & (!g2095) & (g2119)) + ((g174) & (g2108) & (g2110) & (!g2095) & (!g2119)) + ((g174) & (g2108) & (g2110) & (!g2095) & (g2119)) + ((g174) & (g2108) & (g2110) & (g2095) & (!g2119)) + ((g174) & (g2108) & (g2110) & (g2095) & (g2119)));
	assign g2204 = (((!g198) & (!g229) & (g2046) & (g2094)) + ((!g198) & (g229) & (!g2046) & (g2094)) + ((!g198) & (g229) & (g2046) & (!g2094)) + ((!g198) & (g229) & (g2046) & (g2094)) + ((g198) & (!g229) & (!g2046) & (!g2094)) + ((g198) & (!g229) & (!g2046) & (g2094)) + ((g198) & (!g229) & (g2046) & (!g2094)) + ((g198) & (g229) & (!g2046) & (!g2094)));
	assign g2205 = (((!g2109) & (!g2095) & (!g2119) & (g2204)) + ((!g2109) & (g2095) & (!g2119) & (g2204)) + ((!g2109) & (g2095) & (g2119) & (g2204)) + ((g2109) & (!g2095) & (!g2119) & (!g2204)) + ((g2109) & (!g2095) & (g2119) & (!g2204)) + ((g2109) & (!g2095) & (g2119) & (g2204)) + ((g2109) & (g2095) & (!g2119) & (!g2204)) + ((g2109) & (g2095) & (g2119) & (!g2204)));
	assign g2206 = (((!g174) & (!g198) & (g2205) & (g2120) & (g2186)) + ((!g174) & (g198) & (g2205) & (!g2120) & (g2186)) + ((!g174) & (g198) & (g2205) & (g2120) & (!g2186)) + ((!g174) & (g198) & (g2205) & (g2120) & (g2186)) + ((g174) & (!g198) & (!g2205) & (g2120) & (g2186)) + ((g174) & (!g198) & (g2205) & (!g2120) & (!g2186)) + ((g174) & (!g198) & (g2205) & (!g2120) & (g2186)) + ((g174) & (!g198) & (g2205) & (g2120) & (!g2186)) + ((g174) & (!g198) & (g2205) & (g2120) & (g2186)) + ((g174) & (g198) & (!g2205) & (!g2120) & (g2186)) + ((g174) & (g198) & (!g2205) & (g2120) & (!g2186)) + ((g174) & (g198) & (!g2205) & (g2120) & (g2186)) + ((g174) & (g198) & (g2205) & (!g2120) & (!g2186)) + ((g174) & (g198) & (g2205) & (!g2120) & (g2186)) + ((g174) & (g198) & (g2205) & (g2120) & (!g2186)) + ((g174) & (g198) & (g2205) & (g2120) & (g2186)));
	assign g2207 = (((!g127) & (!g147) & (g2202) & (g2203) & (g2206)) + ((!g127) & (g147) & (g2202) & (!g2203) & (g2206)) + ((!g127) & (g147) & (g2202) & (g2203) & (!g2206)) + ((!g127) & (g147) & (g2202) & (g2203) & (g2206)) + ((g127) & (!g147) & (!g2202) & (g2203) & (g2206)) + ((g127) & (!g147) & (g2202) & (!g2203) & (!g2206)) + ((g127) & (!g147) & (g2202) & (!g2203) & (g2206)) + ((g127) & (!g147) & (g2202) & (g2203) & (!g2206)) + ((g127) & (!g147) & (g2202) & (g2203) & (g2206)) + ((g127) & (g147) & (!g2202) & (!g2203) & (g2206)) + ((g127) & (g147) & (!g2202) & (g2203) & (!g2206)) + ((g127) & (g147) & (!g2202) & (g2203) & (g2206)) + ((g127) & (g147) & (g2202) & (!g2203) & (!g2206)) + ((g127) & (g147) & (g2202) & (!g2203) & (g2206)) + ((g127) & (g147) & (g2202) & (g2203) & (!g2206)) + ((g127) & (g147) & (g2202) & (g2203) & (g2206)));
	assign g2208 = (((!g87) & (!g104) & (g2199) & (g2200) & (g2207)) + ((!g87) & (g104) & (g2199) & (!g2200) & (g2207)) + ((!g87) & (g104) & (g2199) & (g2200) & (!g2207)) + ((!g87) & (g104) & (g2199) & (g2200) & (g2207)) + ((g87) & (!g104) & (!g2199) & (g2200) & (g2207)) + ((g87) & (!g104) & (g2199) & (!g2200) & (!g2207)) + ((g87) & (!g104) & (g2199) & (!g2200) & (g2207)) + ((g87) & (!g104) & (g2199) & (g2200) & (!g2207)) + ((g87) & (!g104) & (g2199) & (g2200) & (g2207)) + ((g87) & (g104) & (!g2199) & (!g2200) & (g2207)) + ((g87) & (g104) & (!g2199) & (g2200) & (!g2207)) + ((g87) & (g104) & (!g2199) & (g2200) & (g2207)) + ((g87) & (g104) & (g2199) & (!g2200) & (!g2207)) + ((g87) & (g104) & (g2199) & (!g2200) & (g2207)) + ((g87) & (g104) & (g2199) & (g2200) & (!g2207)) + ((g87) & (g104) & (g2199) & (g2200) & (g2207)));
	assign g2209 = (((!g54) & (!g68) & (g2196) & (g2197) & (g2208)) + ((!g54) & (g68) & (g2196) & (!g2197) & (g2208)) + ((!g54) & (g68) & (g2196) & (g2197) & (!g2208)) + ((!g54) & (g68) & (g2196) & (g2197) & (g2208)) + ((g54) & (!g68) & (!g2196) & (g2197) & (g2208)) + ((g54) & (!g68) & (g2196) & (!g2197) & (!g2208)) + ((g54) & (!g68) & (g2196) & (!g2197) & (g2208)) + ((g54) & (!g68) & (g2196) & (g2197) & (!g2208)) + ((g54) & (!g68) & (g2196) & (g2197) & (g2208)) + ((g54) & (g68) & (!g2196) & (!g2197) & (g2208)) + ((g54) & (g68) & (!g2196) & (g2197) & (!g2208)) + ((g54) & (g68) & (!g2196) & (g2197) & (g2208)) + ((g54) & (g68) & (g2196) & (!g2197) & (!g2208)) + ((g54) & (g68) & (g2196) & (!g2197) & (g2208)) + ((g54) & (g68) & (g2196) & (g2197) & (!g2208)) + ((g54) & (g68) & (g2196) & (g2197) & (g2208)));
	assign g2210 = (((!g27) & (!g39) & (g2193) & (g2194) & (g2209)) + ((!g27) & (g39) & (g2193) & (!g2194) & (g2209)) + ((!g27) & (g39) & (g2193) & (g2194) & (!g2209)) + ((!g27) & (g39) & (g2193) & (g2194) & (g2209)) + ((g27) & (!g39) & (!g2193) & (g2194) & (g2209)) + ((g27) & (!g39) & (g2193) & (!g2194) & (!g2209)) + ((g27) & (!g39) & (g2193) & (!g2194) & (g2209)) + ((g27) & (!g39) & (g2193) & (g2194) & (!g2209)) + ((g27) & (!g39) & (g2193) & (g2194) & (g2209)) + ((g27) & (g39) & (!g2193) & (!g2194) & (g2209)) + ((g27) & (g39) & (!g2193) & (g2194) & (!g2209)) + ((g27) & (g39) & (!g2193) & (g2194) & (g2209)) + ((g27) & (g39) & (g2193) & (!g2194) & (!g2209)) + ((g27) & (g39) & (g2193) & (!g2194) & (g2209)) + ((g27) & (g39) & (g2193) & (g2194) & (!g2209)) + ((g27) & (g39) & (g2193) & (g2194) & (g2209)));
	assign g2211 = (((!g8) & (!g18) & (g2190) & (g2191) & (g2210)) + ((!g8) & (g18) & (g2190) & (!g2191) & (g2210)) + ((!g8) & (g18) & (g2190) & (g2191) & (!g2210)) + ((!g8) & (g18) & (g2190) & (g2191) & (g2210)) + ((g8) & (!g18) & (!g2190) & (g2191) & (g2210)) + ((g8) & (!g18) & (g2190) & (!g2191) & (!g2210)) + ((g8) & (!g18) & (g2190) & (!g2191) & (g2210)) + ((g8) & (!g18) & (g2190) & (g2191) & (!g2210)) + ((g8) & (!g18) & (g2190) & (g2191) & (g2210)) + ((g8) & (g18) & (!g2190) & (!g2191) & (g2210)) + ((g8) & (g18) & (!g2190) & (g2191) & (!g2210)) + ((g8) & (g18) & (!g2190) & (g2191) & (g2210)) + ((g8) & (g18) & (g2190) & (!g2191) & (!g2210)) + ((g8) & (g18) & (g2190) & (!g2191) & (g2210)) + ((g8) & (g18) & (g2190) & (g2191) & (!g2210)) + ((g8) & (g18) & (g2190) & (g2191) & (g2210)));
	assign g2212 = (((!g2) & (!g8) & (g2098) & (g2115)) + ((!g2) & (g8) & (!g2098) & (g2115)) + ((!g2) & (g8) & (g2098) & (!g2115)) + ((!g2) & (g8) & (g2098) & (g2115)) + ((g2) & (!g8) & (!g2098) & (!g2115)) + ((g2) & (!g8) & (!g2098) & (g2115)) + ((g2) & (!g8) & (g2098) & (!g2115)) + ((g2) & (g8) & (!g2098) & (!g2115)));
	assign g2213 = (((!g2097) & (!g2095) & (!g2119) & (g2212)) + ((!g2097) & (g2095) & (!g2119) & (g2212)) + ((!g2097) & (g2095) & (g2119) & (g2212)) + ((g2097) & (!g2095) & (!g2119) & (!g2212)) + ((g2097) & (!g2095) & (g2119) & (!g2212)) + ((g2097) & (!g2095) & (g2119) & (g2212)) + ((g2097) & (g2095) & (!g2119) & (!g2212)) + ((g2097) & (g2095) & (g2119) & (!g2212)));
	assign g2214 = (((!g4) & (!g2) & (!g2188) & (!g2211) & (g2213)) + ((!g4) & (!g2) & (!g2188) & (g2211) & (g2213)) + ((!g4) & (!g2) & (g2188) & (!g2211) & (g2213)) + ((!g4) & (!g2) & (g2188) & (g2211) & (!g2213)) + ((!g4) & (!g2) & (g2188) & (g2211) & (g2213)) + ((!g4) & (g2) & (!g2188) & (!g2211) & (g2213)) + ((!g4) & (g2) & (!g2188) & (g2211) & (!g2213)) + ((!g4) & (g2) & (!g2188) & (g2211) & (g2213)) + ((!g4) & (g2) & (g2188) & (!g2211) & (!g2213)) + ((!g4) & (g2) & (g2188) & (!g2211) & (g2213)) + ((!g4) & (g2) & (g2188) & (g2211) & (!g2213)) + ((!g4) & (g2) & (g2188) & (g2211) & (g2213)) + ((g4) & (!g2) & (g2188) & (g2211) & (g2213)) + ((g4) & (g2) & (!g2188) & (g2211) & (g2213)) + ((g4) & (g2) & (g2188) & (!g2211) & (g2213)) + ((g4) & (g2) & (g2188) & (g2211) & (g2213)));
	assign g2215 = (((!g4) & (!g2116) & (g2117)) + ((!g4) & (g2116) & (!g2117)) + ((!g4) & (g2116) & (g2117)) + ((g4) & (g2116) & (g2117)));
	assign g2216 = (((!g2096) & (!g2215) & (!g2095) & (!g2119)) + ((!g2096) & (!g2215) & (g2095) & (!g2119)) + ((!g2096) & (!g2215) & (g2095) & (g2119)) + ((g2096) & (g2215) & (!g2095) & (!g2119)) + ((g2096) & (g2215) & (!g2095) & (g2119)) + ((g2096) & (g2215) & (g2095) & (!g2119)) + ((g2096) & (g2215) & (g2095) & (g2119)));
	assign g2217 = (((!g1) & (g2096) & (!g2215) & (!g2095) & (g2119)) + ((!g1) & (g2096) & (g2215) & (!g2095) & (g2119)) + ((g1) & (!g2096) & (g2215) & (g2095) & (!g2119)) + ((g1) & (!g2096) & (g2215) & (g2095) & (g2119)) + ((g1) & (g2096) & (!g2215) & (!g2095) & (!g2119)) + ((g1) & (g2096) & (!g2215) & (!g2095) & (g2119)) + ((g1) & (g2096) & (!g2215) & (g2095) & (!g2119)) + ((g1) & (g2096) & (!g2215) & (g2095) & (g2119)) + ((g1) & (g2096) & (g2215) & (!g2095) & (g2119)));
	assign g2218 = (((!g1) & (!g2187) & (!g2214) & (!g2216) & (!g2217)) + ((g1) & (!g2187) & (!g2214) & (!g2216) & (!g2217)) + ((g1) & (!g2187) & (!g2214) & (g2216) & (!g2217)) + ((g1) & (!g2187) & (g2214) & (!g2216) & (!g2217)) + ((g1) & (!g2187) & (g2214) & (g2216) & (!g2217)) + ((g1) & (g2187) & (!g2214) & (!g2216) & (!g2217)) + ((g1) & (g2187) & (!g2214) & (g2216) & (!g2217)));
	assign g2219 = (((!g198) & (!g2120) & (g2186) & (!g2218)) + ((!g198) & (g2120) & (!g2186) & (!g2218)) + ((!g198) & (g2120) & (!g2186) & (g2218)) + ((!g198) & (g2120) & (g2186) & (g2218)) + ((g198) & (!g2120) & (!g2186) & (!g2218)) + ((g198) & (g2120) & (!g2186) & (g2218)) + ((g198) & (g2120) & (g2186) & (!g2218)) + ((g198) & (g2120) & (g2186) & (g2218)));
	assign g2220 = (((!g229) & (!g255) & (!g2122) & (g2123) & (g2185) & (!g2218)) + ((!g229) & (!g255) & (g2122) & (!g2123) & (!g2185) & (!g2218)) + ((!g229) & (!g255) & (g2122) & (!g2123) & (!g2185) & (g2218)) + ((!g229) & (!g255) & (g2122) & (!g2123) & (g2185) & (!g2218)) + ((!g229) & (!g255) & (g2122) & (!g2123) & (g2185) & (g2218)) + ((!g229) & (!g255) & (g2122) & (g2123) & (!g2185) & (!g2218)) + ((!g229) & (!g255) & (g2122) & (g2123) & (!g2185) & (g2218)) + ((!g229) & (!g255) & (g2122) & (g2123) & (g2185) & (g2218)) + ((!g229) & (g255) & (!g2122) & (!g2123) & (g2185) & (!g2218)) + ((!g229) & (g255) & (!g2122) & (g2123) & (!g2185) & (!g2218)) + ((!g229) & (g255) & (!g2122) & (g2123) & (g2185) & (!g2218)) + ((!g229) & (g255) & (g2122) & (!g2123) & (!g2185) & (!g2218)) + ((!g229) & (g255) & (g2122) & (!g2123) & (!g2185) & (g2218)) + ((!g229) & (g255) & (g2122) & (!g2123) & (g2185) & (g2218)) + ((!g229) & (g255) & (g2122) & (g2123) & (!g2185) & (g2218)) + ((!g229) & (g255) & (g2122) & (g2123) & (g2185) & (g2218)) + ((g229) & (!g255) & (!g2122) & (!g2123) & (!g2185) & (!g2218)) + ((g229) & (!g255) & (!g2122) & (!g2123) & (g2185) & (!g2218)) + ((g229) & (!g255) & (!g2122) & (g2123) & (!g2185) & (!g2218)) + ((g229) & (!g255) & (g2122) & (!g2123) & (!g2185) & (g2218)) + ((g229) & (!g255) & (g2122) & (!g2123) & (g2185) & (g2218)) + ((g229) & (!g255) & (g2122) & (g2123) & (!g2185) & (g2218)) + ((g229) & (!g255) & (g2122) & (g2123) & (g2185) & (!g2218)) + ((g229) & (!g255) & (g2122) & (g2123) & (g2185) & (g2218)) + ((g229) & (g255) & (!g2122) & (!g2123) & (!g2185) & (!g2218)) + ((g229) & (g255) & (g2122) & (!g2123) & (!g2185) & (g2218)) + ((g229) & (g255) & (g2122) & (!g2123) & (g2185) & (!g2218)) + ((g229) & (g255) & (g2122) & (!g2123) & (g2185) & (g2218)) + ((g229) & (g255) & (g2122) & (g2123) & (!g2185) & (!g2218)) + ((g229) & (g255) & (g2122) & (g2123) & (!g2185) & (g2218)) + ((g229) & (g255) & (g2122) & (g2123) & (g2185) & (!g2218)) + ((g229) & (g255) & (g2122) & (g2123) & (g2185) & (g2218)));
	assign g2221 = (((!g255) & (!g2123) & (g2185) & (!g2218)) + ((!g255) & (g2123) & (!g2185) & (!g2218)) + ((!g255) & (g2123) & (!g2185) & (g2218)) + ((!g255) & (g2123) & (g2185) & (g2218)) + ((g255) & (!g2123) & (!g2185) & (!g2218)) + ((g255) & (g2123) & (!g2185) & (g2218)) + ((g255) & (g2123) & (g2185) & (!g2218)) + ((g255) & (g2123) & (g2185) & (g2218)));
	assign g2222 = (((!g290) & (!g319) & (!g2125) & (g2126) & (g2184) & (!g2218)) + ((!g290) & (!g319) & (g2125) & (!g2126) & (!g2184) & (!g2218)) + ((!g290) & (!g319) & (g2125) & (!g2126) & (!g2184) & (g2218)) + ((!g290) & (!g319) & (g2125) & (!g2126) & (g2184) & (!g2218)) + ((!g290) & (!g319) & (g2125) & (!g2126) & (g2184) & (g2218)) + ((!g290) & (!g319) & (g2125) & (g2126) & (!g2184) & (!g2218)) + ((!g290) & (!g319) & (g2125) & (g2126) & (!g2184) & (g2218)) + ((!g290) & (!g319) & (g2125) & (g2126) & (g2184) & (g2218)) + ((!g290) & (g319) & (!g2125) & (!g2126) & (g2184) & (!g2218)) + ((!g290) & (g319) & (!g2125) & (g2126) & (!g2184) & (!g2218)) + ((!g290) & (g319) & (!g2125) & (g2126) & (g2184) & (!g2218)) + ((!g290) & (g319) & (g2125) & (!g2126) & (!g2184) & (!g2218)) + ((!g290) & (g319) & (g2125) & (!g2126) & (!g2184) & (g2218)) + ((!g290) & (g319) & (g2125) & (!g2126) & (g2184) & (g2218)) + ((!g290) & (g319) & (g2125) & (g2126) & (!g2184) & (g2218)) + ((!g290) & (g319) & (g2125) & (g2126) & (g2184) & (g2218)) + ((g290) & (!g319) & (!g2125) & (!g2126) & (!g2184) & (!g2218)) + ((g290) & (!g319) & (!g2125) & (!g2126) & (g2184) & (!g2218)) + ((g290) & (!g319) & (!g2125) & (g2126) & (!g2184) & (!g2218)) + ((g290) & (!g319) & (g2125) & (!g2126) & (!g2184) & (g2218)) + ((g290) & (!g319) & (g2125) & (!g2126) & (g2184) & (g2218)) + ((g290) & (!g319) & (g2125) & (g2126) & (!g2184) & (g2218)) + ((g290) & (!g319) & (g2125) & (g2126) & (g2184) & (!g2218)) + ((g290) & (!g319) & (g2125) & (g2126) & (g2184) & (g2218)) + ((g290) & (g319) & (!g2125) & (!g2126) & (!g2184) & (!g2218)) + ((g290) & (g319) & (g2125) & (!g2126) & (!g2184) & (g2218)) + ((g290) & (g319) & (g2125) & (!g2126) & (g2184) & (!g2218)) + ((g290) & (g319) & (g2125) & (!g2126) & (g2184) & (g2218)) + ((g290) & (g319) & (g2125) & (g2126) & (!g2184) & (!g2218)) + ((g290) & (g319) & (g2125) & (g2126) & (!g2184) & (g2218)) + ((g290) & (g319) & (g2125) & (g2126) & (g2184) & (!g2218)) + ((g290) & (g319) & (g2125) & (g2126) & (g2184) & (g2218)));
	assign g2223 = (((!g319) & (!g2126) & (g2184) & (!g2218)) + ((!g319) & (g2126) & (!g2184) & (!g2218)) + ((!g319) & (g2126) & (!g2184) & (g2218)) + ((!g319) & (g2126) & (g2184) & (g2218)) + ((g319) & (!g2126) & (!g2184) & (!g2218)) + ((g319) & (g2126) & (!g2184) & (g2218)) + ((g319) & (g2126) & (g2184) & (!g2218)) + ((g319) & (g2126) & (g2184) & (g2218)));
	assign g2224 = (((!g358) & (!g390) & (!g2128) & (g2129) & (g2183) & (!g2218)) + ((!g358) & (!g390) & (g2128) & (!g2129) & (!g2183) & (!g2218)) + ((!g358) & (!g390) & (g2128) & (!g2129) & (!g2183) & (g2218)) + ((!g358) & (!g390) & (g2128) & (!g2129) & (g2183) & (!g2218)) + ((!g358) & (!g390) & (g2128) & (!g2129) & (g2183) & (g2218)) + ((!g358) & (!g390) & (g2128) & (g2129) & (!g2183) & (!g2218)) + ((!g358) & (!g390) & (g2128) & (g2129) & (!g2183) & (g2218)) + ((!g358) & (!g390) & (g2128) & (g2129) & (g2183) & (g2218)) + ((!g358) & (g390) & (!g2128) & (!g2129) & (g2183) & (!g2218)) + ((!g358) & (g390) & (!g2128) & (g2129) & (!g2183) & (!g2218)) + ((!g358) & (g390) & (!g2128) & (g2129) & (g2183) & (!g2218)) + ((!g358) & (g390) & (g2128) & (!g2129) & (!g2183) & (!g2218)) + ((!g358) & (g390) & (g2128) & (!g2129) & (!g2183) & (g2218)) + ((!g358) & (g390) & (g2128) & (!g2129) & (g2183) & (g2218)) + ((!g358) & (g390) & (g2128) & (g2129) & (!g2183) & (g2218)) + ((!g358) & (g390) & (g2128) & (g2129) & (g2183) & (g2218)) + ((g358) & (!g390) & (!g2128) & (!g2129) & (!g2183) & (!g2218)) + ((g358) & (!g390) & (!g2128) & (!g2129) & (g2183) & (!g2218)) + ((g358) & (!g390) & (!g2128) & (g2129) & (!g2183) & (!g2218)) + ((g358) & (!g390) & (g2128) & (!g2129) & (!g2183) & (g2218)) + ((g358) & (!g390) & (g2128) & (!g2129) & (g2183) & (g2218)) + ((g358) & (!g390) & (g2128) & (g2129) & (!g2183) & (g2218)) + ((g358) & (!g390) & (g2128) & (g2129) & (g2183) & (!g2218)) + ((g358) & (!g390) & (g2128) & (g2129) & (g2183) & (g2218)) + ((g358) & (g390) & (!g2128) & (!g2129) & (!g2183) & (!g2218)) + ((g358) & (g390) & (g2128) & (!g2129) & (!g2183) & (g2218)) + ((g358) & (g390) & (g2128) & (!g2129) & (g2183) & (!g2218)) + ((g358) & (g390) & (g2128) & (!g2129) & (g2183) & (g2218)) + ((g358) & (g390) & (g2128) & (g2129) & (!g2183) & (!g2218)) + ((g358) & (g390) & (g2128) & (g2129) & (!g2183) & (g2218)) + ((g358) & (g390) & (g2128) & (g2129) & (g2183) & (!g2218)) + ((g358) & (g390) & (g2128) & (g2129) & (g2183) & (g2218)));
	assign g2225 = (((!g390) & (!g2129) & (g2183) & (!g2218)) + ((!g390) & (g2129) & (!g2183) & (!g2218)) + ((!g390) & (g2129) & (!g2183) & (g2218)) + ((!g390) & (g2129) & (g2183) & (g2218)) + ((g390) & (!g2129) & (!g2183) & (!g2218)) + ((g390) & (g2129) & (!g2183) & (g2218)) + ((g390) & (g2129) & (g2183) & (!g2218)) + ((g390) & (g2129) & (g2183) & (g2218)));
	assign g2226 = (((!g433) & (!g468) & (!g2131) & (g2132) & (g2182) & (!g2218)) + ((!g433) & (!g468) & (g2131) & (!g2132) & (!g2182) & (!g2218)) + ((!g433) & (!g468) & (g2131) & (!g2132) & (!g2182) & (g2218)) + ((!g433) & (!g468) & (g2131) & (!g2132) & (g2182) & (!g2218)) + ((!g433) & (!g468) & (g2131) & (!g2132) & (g2182) & (g2218)) + ((!g433) & (!g468) & (g2131) & (g2132) & (!g2182) & (!g2218)) + ((!g433) & (!g468) & (g2131) & (g2132) & (!g2182) & (g2218)) + ((!g433) & (!g468) & (g2131) & (g2132) & (g2182) & (g2218)) + ((!g433) & (g468) & (!g2131) & (!g2132) & (g2182) & (!g2218)) + ((!g433) & (g468) & (!g2131) & (g2132) & (!g2182) & (!g2218)) + ((!g433) & (g468) & (!g2131) & (g2132) & (g2182) & (!g2218)) + ((!g433) & (g468) & (g2131) & (!g2132) & (!g2182) & (!g2218)) + ((!g433) & (g468) & (g2131) & (!g2132) & (!g2182) & (g2218)) + ((!g433) & (g468) & (g2131) & (!g2132) & (g2182) & (g2218)) + ((!g433) & (g468) & (g2131) & (g2132) & (!g2182) & (g2218)) + ((!g433) & (g468) & (g2131) & (g2132) & (g2182) & (g2218)) + ((g433) & (!g468) & (!g2131) & (!g2132) & (!g2182) & (!g2218)) + ((g433) & (!g468) & (!g2131) & (!g2132) & (g2182) & (!g2218)) + ((g433) & (!g468) & (!g2131) & (g2132) & (!g2182) & (!g2218)) + ((g433) & (!g468) & (g2131) & (!g2132) & (!g2182) & (g2218)) + ((g433) & (!g468) & (g2131) & (!g2132) & (g2182) & (g2218)) + ((g433) & (!g468) & (g2131) & (g2132) & (!g2182) & (g2218)) + ((g433) & (!g468) & (g2131) & (g2132) & (g2182) & (!g2218)) + ((g433) & (!g468) & (g2131) & (g2132) & (g2182) & (g2218)) + ((g433) & (g468) & (!g2131) & (!g2132) & (!g2182) & (!g2218)) + ((g433) & (g468) & (g2131) & (!g2132) & (!g2182) & (g2218)) + ((g433) & (g468) & (g2131) & (!g2132) & (g2182) & (!g2218)) + ((g433) & (g468) & (g2131) & (!g2132) & (g2182) & (g2218)) + ((g433) & (g468) & (g2131) & (g2132) & (!g2182) & (!g2218)) + ((g433) & (g468) & (g2131) & (g2132) & (!g2182) & (g2218)) + ((g433) & (g468) & (g2131) & (g2132) & (g2182) & (!g2218)) + ((g433) & (g468) & (g2131) & (g2132) & (g2182) & (g2218)));
	assign g2227 = (((!g468) & (!g2132) & (g2182) & (!g2218)) + ((!g468) & (g2132) & (!g2182) & (!g2218)) + ((!g468) & (g2132) & (!g2182) & (g2218)) + ((!g468) & (g2132) & (g2182) & (g2218)) + ((g468) & (!g2132) & (!g2182) & (!g2218)) + ((g468) & (g2132) & (!g2182) & (g2218)) + ((g468) & (g2132) & (g2182) & (!g2218)) + ((g468) & (g2132) & (g2182) & (g2218)));
	assign g2228 = (((!g515) & (!g553) & (!g2134) & (g2135) & (g2181) & (!g2218)) + ((!g515) & (!g553) & (g2134) & (!g2135) & (!g2181) & (!g2218)) + ((!g515) & (!g553) & (g2134) & (!g2135) & (!g2181) & (g2218)) + ((!g515) & (!g553) & (g2134) & (!g2135) & (g2181) & (!g2218)) + ((!g515) & (!g553) & (g2134) & (!g2135) & (g2181) & (g2218)) + ((!g515) & (!g553) & (g2134) & (g2135) & (!g2181) & (!g2218)) + ((!g515) & (!g553) & (g2134) & (g2135) & (!g2181) & (g2218)) + ((!g515) & (!g553) & (g2134) & (g2135) & (g2181) & (g2218)) + ((!g515) & (g553) & (!g2134) & (!g2135) & (g2181) & (!g2218)) + ((!g515) & (g553) & (!g2134) & (g2135) & (!g2181) & (!g2218)) + ((!g515) & (g553) & (!g2134) & (g2135) & (g2181) & (!g2218)) + ((!g515) & (g553) & (g2134) & (!g2135) & (!g2181) & (!g2218)) + ((!g515) & (g553) & (g2134) & (!g2135) & (!g2181) & (g2218)) + ((!g515) & (g553) & (g2134) & (!g2135) & (g2181) & (g2218)) + ((!g515) & (g553) & (g2134) & (g2135) & (!g2181) & (g2218)) + ((!g515) & (g553) & (g2134) & (g2135) & (g2181) & (g2218)) + ((g515) & (!g553) & (!g2134) & (!g2135) & (!g2181) & (!g2218)) + ((g515) & (!g553) & (!g2134) & (!g2135) & (g2181) & (!g2218)) + ((g515) & (!g553) & (!g2134) & (g2135) & (!g2181) & (!g2218)) + ((g515) & (!g553) & (g2134) & (!g2135) & (!g2181) & (g2218)) + ((g515) & (!g553) & (g2134) & (!g2135) & (g2181) & (g2218)) + ((g515) & (!g553) & (g2134) & (g2135) & (!g2181) & (g2218)) + ((g515) & (!g553) & (g2134) & (g2135) & (g2181) & (!g2218)) + ((g515) & (!g553) & (g2134) & (g2135) & (g2181) & (g2218)) + ((g515) & (g553) & (!g2134) & (!g2135) & (!g2181) & (!g2218)) + ((g515) & (g553) & (g2134) & (!g2135) & (!g2181) & (g2218)) + ((g515) & (g553) & (g2134) & (!g2135) & (g2181) & (!g2218)) + ((g515) & (g553) & (g2134) & (!g2135) & (g2181) & (g2218)) + ((g515) & (g553) & (g2134) & (g2135) & (!g2181) & (!g2218)) + ((g515) & (g553) & (g2134) & (g2135) & (!g2181) & (g2218)) + ((g515) & (g553) & (g2134) & (g2135) & (g2181) & (!g2218)) + ((g515) & (g553) & (g2134) & (g2135) & (g2181) & (g2218)));
	assign g2229 = (((!g553) & (!g2135) & (g2181) & (!g2218)) + ((!g553) & (g2135) & (!g2181) & (!g2218)) + ((!g553) & (g2135) & (!g2181) & (g2218)) + ((!g553) & (g2135) & (g2181) & (g2218)) + ((g553) & (!g2135) & (!g2181) & (!g2218)) + ((g553) & (g2135) & (!g2181) & (g2218)) + ((g553) & (g2135) & (g2181) & (!g2218)) + ((g553) & (g2135) & (g2181) & (g2218)));
	assign g2230 = (((!g604) & (!g645) & (!g2137) & (g2138) & (g2180) & (!g2218)) + ((!g604) & (!g645) & (g2137) & (!g2138) & (!g2180) & (!g2218)) + ((!g604) & (!g645) & (g2137) & (!g2138) & (!g2180) & (g2218)) + ((!g604) & (!g645) & (g2137) & (!g2138) & (g2180) & (!g2218)) + ((!g604) & (!g645) & (g2137) & (!g2138) & (g2180) & (g2218)) + ((!g604) & (!g645) & (g2137) & (g2138) & (!g2180) & (!g2218)) + ((!g604) & (!g645) & (g2137) & (g2138) & (!g2180) & (g2218)) + ((!g604) & (!g645) & (g2137) & (g2138) & (g2180) & (g2218)) + ((!g604) & (g645) & (!g2137) & (!g2138) & (g2180) & (!g2218)) + ((!g604) & (g645) & (!g2137) & (g2138) & (!g2180) & (!g2218)) + ((!g604) & (g645) & (!g2137) & (g2138) & (g2180) & (!g2218)) + ((!g604) & (g645) & (g2137) & (!g2138) & (!g2180) & (!g2218)) + ((!g604) & (g645) & (g2137) & (!g2138) & (!g2180) & (g2218)) + ((!g604) & (g645) & (g2137) & (!g2138) & (g2180) & (g2218)) + ((!g604) & (g645) & (g2137) & (g2138) & (!g2180) & (g2218)) + ((!g604) & (g645) & (g2137) & (g2138) & (g2180) & (g2218)) + ((g604) & (!g645) & (!g2137) & (!g2138) & (!g2180) & (!g2218)) + ((g604) & (!g645) & (!g2137) & (!g2138) & (g2180) & (!g2218)) + ((g604) & (!g645) & (!g2137) & (g2138) & (!g2180) & (!g2218)) + ((g604) & (!g645) & (g2137) & (!g2138) & (!g2180) & (g2218)) + ((g604) & (!g645) & (g2137) & (!g2138) & (g2180) & (g2218)) + ((g604) & (!g645) & (g2137) & (g2138) & (!g2180) & (g2218)) + ((g604) & (!g645) & (g2137) & (g2138) & (g2180) & (!g2218)) + ((g604) & (!g645) & (g2137) & (g2138) & (g2180) & (g2218)) + ((g604) & (g645) & (!g2137) & (!g2138) & (!g2180) & (!g2218)) + ((g604) & (g645) & (g2137) & (!g2138) & (!g2180) & (g2218)) + ((g604) & (g645) & (g2137) & (!g2138) & (g2180) & (!g2218)) + ((g604) & (g645) & (g2137) & (!g2138) & (g2180) & (g2218)) + ((g604) & (g645) & (g2137) & (g2138) & (!g2180) & (!g2218)) + ((g604) & (g645) & (g2137) & (g2138) & (!g2180) & (g2218)) + ((g604) & (g645) & (g2137) & (g2138) & (g2180) & (!g2218)) + ((g604) & (g645) & (g2137) & (g2138) & (g2180) & (g2218)));
	assign g2231 = (((!g645) & (!g2138) & (g2180) & (!g2218)) + ((!g645) & (g2138) & (!g2180) & (!g2218)) + ((!g645) & (g2138) & (!g2180) & (g2218)) + ((!g645) & (g2138) & (g2180) & (g2218)) + ((g645) & (!g2138) & (!g2180) & (!g2218)) + ((g645) & (g2138) & (!g2180) & (g2218)) + ((g645) & (g2138) & (g2180) & (!g2218)) + ((g645) & (g2138) & (g2180) & (g2218)));
	assign g2232 = (((!g700) & (!g744) & (!g2140) & (g2141) & (g2179) & (!g2218)) + ((!g700) & (!g744) & (g2140) & (!g2141) & (!g2179) & (!g2218)) + ((!g700) & (!g744) & (g2140) & (!g2141) & (!g2179) & (g2218)) + ((!g700) & (!g744) & (g2140) & (!g2141) & (g2179) & (!g2218)) + ((!g700) & (!g744) & (g2140) & (!g2141) & (g2179) & (g2218)) + ((!g700) & (!g744) & (g2140) & (g2141) & (!g2179) & (!g2218)) + ((!g700) & (!g744) & (g2140) & (g2141) & (!g2179) & (g2218)) + ((!g700) & (!g744) & (g2140) & (g2141) & (g2179) & (g2218)) + ((!g700) & (g744) & (!g2140) & (!g2141) & (g2179) & (!g2218)) + ((!g700) & (g744) & (!g2140) & (g2141) & (!g2179) & (!g2218)) + ((!g700) & (g744) & (!g2140) & (g2141) & (g2179) & (!g2218)) + ((!g700) & (g744) & (g2140) & (!g2141) & (!g2179) & (!g2218)) + ((!g700) & (g744) & (g2140) & (!g2141) & (!g2179) & (g2218)) + ((!g700) & (g744) & (g2140) & (!g2141) & (g2179) & (g2218)) + ((!g700) & (g744) & (g2140) & (g2141) & (!g2179) & (g2218)) + ((!g700) & (g744) & (g2140) & (g2141) & (g2179) & (g2218)) + ((g700) & (!g744) & (!g2140) & (!g2141) & (!g2179) & (!g2218)) + ((g700) & (!g744) & (!g2140) & (!g2141) & (g2179) & (!g2218)) + ((g700) & (!g744) & (!g2140) & (g2141) & (!g2179) & (!g2218)) + ((g700) & (!g744) & (g2140) & (!g2141) & (!g2179) & (g2218)) + ((g700) & (!g744) & (g2140) & (!g2141) & (g2179) & (g2218)) + ((g700) & (!g744) & (g2140) & (g2141) & (!g2179) & (g2218)) + ((g700) & (!g744) & (g2140) & (g2141) & (g2179) & (!g2218)) + ((g700) & (!g744) & (g2140) & (g2141) & (g2179) & (g2218)) + ((g700) & (g744) & (!g2140) & (!g2141) & (!g2179) & (!g2218)) + ((g700) & (g744) & (g2140) & (!g2141) & (!g2179) & (g2218)) + ((g700) & (g744) & (g2140) & (!g2141) & (g2179) & (!g2218)) + ((g700) & (g744) & (g2140) & (!g2141) & (g2179) & (g2218)) + ((g700) & (g744) & (g2140) & (g2141) & (!g2179) & (!g2218)) + ((g700) & (g744) & (g2140) & (g2141) & (!g2179) & (g2218)) + ((g700) & (g744) & (g2140) & (g2141) & (g2179) & (!g2218)) + ((g700) & (g744) & (g2140) & (g2141) & (g2179) & (g2218)));
	assign g2233 = (((!g744) & (!g2141) & (g2179) & (!g2218)) + ((!g744) & (g2141) & (!g2179) & (!g2218)) + ((!g744) & (g2141) & (!g2179) & (g2218)) + ((!g744) & (g2141) & (g2179) & (g2218)) + ((g744) & (!g2141) & (!g2179) & (!g2218)) + ((g744) & (g2141) & (!g2179) & (g2218)) + ((g744) & (g2141) & (g2179) & (!g2218)) + ((g744) & (g2141) & (g2179) & (g2218)));
	assign g2234 = (((!g803) & (!g851) & (!g2143) & (g2144) & (g2178) & (!g2218)) + ((!g803) & (!g851) & (g2143) & (!g2144) & (!g2178) & (!g2218)) + ((!g803) & (!g851) & (g2143) & (!g2144) & (!g2178) & (g2218)) + ((!g803) & (!g851) & (g2143) & (!g2144) & (g2178) & (!g2218)) + ((!g803) & (!g851) & (g2143) & (!g2144) & (g2178) & (g2218)) + ((!g803) & (!g851) & (g2143) & (g2144) & (!g2178) & (!g2218)) + ((!g803) & (!g851) & (g2143) & (g2144) & (!g2178) & (g2218)) + ((!g803) & (!g851) & (g2143) & (g2144) & (g2178) & (g2218)) + ((!g803) & (g851) & (!g2143) & (!g2144) & (g2178) & (!g2218)) + ((!g803) & (g851) & (!g2143) & (g2144) & (!g2178) & (!g2218)) + ((!g803) & (g851) & (!g2143) & (g2144) & (g2178) & (!g2218)) + ((!g803) & (g851) & (g2143) & (!g2144) & (!g2178) & (!g2218)) + ((!g803) & (g851) & (g2143) & (!g2144) & (!g2178) & (g2218)) + ((!g803) & (g851) & (g2143) & (!g2144) & (g2178) & (g2218)) + ((!g803) & (g851) & (g2143) & (g2144) & (!g2178) & (g2218)) + ((!g803) & (g851) & (g2143) & (g2144) & (g2178) & (g2218)) + ((g803) & (!g851) & (!g2143) & (!g2144) & (!g2178) & (!g2218)) + ((g803) & (!g851) & (!g2143) & (!g2144) & (g2178) & (!g2218)) + ((g803) & (!g851) & (!g2143) & (g2144) & (!g2178) & (!g2218)) + ((g803) & (!g851) & (g2143) & (!g2144) & (!g2178) & (g2218)) + ((g803) & (!g851) & (g2143) & (!g2144) & (g2178) & (g2218)) + ((g803) & (!g851) & (g2143) & (g2144) & (!g2178) & (g2218)) + ((g803) & (!g851) & (g2143) & (g2144) & (g2178) & (!g2218)) + ((g803) & (!g851) & (g2143) & (g2144) & (g2178) & (g2218)) + ((g803) & (g851) & (!g2143) & (!g2144) & (!g2178) & (!g2218)) + ((g803) & (g851) & (g2143) & (!g2144) & (!g2178) & (g2218)) + ((g803) & (g851) & (g2143) & (!g2144) & (g2178) & (!g2218)) + ((g803) & (g851) & (g2143) & (!g2144) & (g2178) & (g2218)) + ((g803) & (g851) & (g2143) & (g2144) & (!g2178) & (!g2218)) + ((g803) & (g851) & (g2143) & (g2144) & (!g2178) & (g2218)) + ((g803) & (g851) & (g2143) & (g2144) & (g2178) & (!g2218)) + ((g803) & (g851) & (g2143) & (g2144) & (g2178) & (g2218)));
	assign g2235 = (((!g851) & (!g2144) & (g2178) & (!g2218)) + ((!g851) & (g2144) & (!g2178) & (!g2218)) + ((!g851) & (g2144) & (!g2178) & (g2218)) + ((!g851) & (g2144) & (g2178) & (g2218)) + ((g851) & (!g2144) & (!g2178) & (!g2218)) + ((g851) & (g2144) & (!g2178) & (g2218)) + ((g851) & (g2144) & (g2178) & (!g2218)) + ((g851) & (g2144) & (g2178) & (g2218)));
	assign g2236 = (((!g914) & (!g1032) & (!g2146) & (g2147) & (g2177) & (!g2218)) + ((!g914) & (!g1032) & (g2146) & (!g2147) & (!g2177) & (!g2218)) + ((!g914) & (!g1032) & (g2146) & (!g2147) & (!g2177) & (g2218)) + ((!g914) & (!g1032) & (g2146) & (!g2147) & (g2177) & (!g2218)) + ((!g914) & (!g1032) & (g2146) & (!g2147) & (g2177) & (g2218)) + ((!g914) & (!g1032) & (g2146) & (g2147) & (!g2177) & (!g2218)) + ((!g914) & (!g1032) & (g2146) & (g2147) & (!g2177) & (g2218)) + ((!g914) & (!g1032) & (g2146) & (g2147) & (g2177) & (g2218)) + ((!g914) & (g1032) & (!g2146) & (!g2147) & (g2177) & (!g2218)) + ((!g914) & (g1032) & (!g2146) & (g2147) & (!g2177) & (!g2218)) + ((!g914) & (g1032) & (!g2146) & (g2147) & (g2177) & (!g2218)) + ((!g914) & (g1032) & (g2146) & (!g2147) & (!g2177) & (!g2218)) + ((!g914) & (g1032) & (g2146) & (!g2147) & (!g2177) & (g2218)) + ((!g914) & (g1032) & (g2146) & (!g2147) & (g2177) & (g2218)) + ((!g914) & (g1032) & (g2146) & (g2147) & (!g2177) & (g2218)) + ((!g914) & (g1032) & (g2146) & (g2147) & (g2177) & (g2218)) + ((g914) & (!g1032) & (!g2146) & (!g2147) & (!g2177) & (!g2218)) + ((g914) & (!g1032) & (!g2146) & (!g2147) & (g2177) & (!g2218)) + ((g914) & (!g1032) & (!g2146) & (g2147) & (!g2177) & (!g2218)) + ((g914) & (!g1032) & (g2146) & (!g2147) & (!g2177) & (g2218)) + ((g914) & (!g1032) & (g2146) & (!g2147) & (g2177) & (g2218)) + ((g914) & (!g1032) & (g2146) & (g2147) & (!g2177) & (g2218)) + ((g914) & (!g1032) & (g2146) & (g2147) & (g2177) & (!g2218)) + ((g914) & (!g1032) & (g2146) & (g2147) & (g2177) & (g2218)) + ((g914) & (g1032) & (!g2146) & (!g2147) & (!g2177) & (!g2218)) + ((g914) & (g1032) & (g2146) & (!g2147) & (!g2177) & (g2218)) + ((g914) & (g1032) & (g2146) & (!g2147) & (g2177) & (!g2218)) + ((g914) & (g1032) & (g2146) & (!g2147) & (g2177) & (g2218)) + ((g914) & (g1032) & (g2146) & (g2147) & (!g2177) & (!g2218)) + ((g914) & (g1032) & (g2146) & (g2147) & (!g2177) & (g2218)) + ((g914) & (g1032) & (g2146) & (g2147) & (g2177) & (!g2218)) + ((g914) & (g1032) & (g2146) & (g2147) & (g2177) & (g2218)));
	assign g2237 = (((!g1032) & (!g2147) & (g2177) & (!g2218)) + ((!g1032) & (g2147) & (!g2177) & (!g2218)) + ((!g1032) & (g2147) & (!g2177) & (g2218)) + ((!g1032) & (g2147) & (g2177) & (g2218)) + ((g1032) & (!g2147) & (!g2177) & (!g2218)) + ((g1032) & (g2147) & (!g2177) & (g2218)) + ((g1032) & (g2147) & (g2177) & (!g2218)) + ((g1032) & (g2147) & (g2177) & (g2218)));
	assign g2238 = (((!g1030) & (!g1160) & (!g2149) & (g2150) & (g2176) & (!g2218)) + ((!g1030) & (!g1160) & (g2149) & (!g2150) & (!g2176) & (!g2218)) + ((!g1030) & (!g1160) & (g2149) & (!g2150) & (!g2176) & (g2218)) + ((!g1030) & (!g1160) & (g2149) & (!g2150) & (g2176) & (!g2218)) + ((!g1030) & (!g1160) & (g2149) & (!g2150) & (g2176) & (g2218)) + ((!g1030) & (!g1160) & (g2149) & (g2150) & (!g2176) & (!g2218)) + ((!g1030) & (!g1160) & (g2149) & (g2150) & (!g2176) & (g2218)) + ((!g1030) & (!g1160) & (g2149) & (g2150) & (g2176) & (g2218)) + ((!g1030) & (g1160) & (!g2149) & (!g2150) & (g2176) & (!g2218)) + ((!g1030) & (g1160) & (!g2149) & (g2150) & (!g2176) & (!g2218)) + ((!g1030) & (g1160) & (!g2149) & (g2150) & (g2176) & (!g2218)) + ((!g1030) & (g1160) & (g2149) & (!g2150) & (!g2176) & (!g2218)) + ((!g1030) & (g1160) & (g2149) & (!g2150) & (!g2176) & (g2218)) + ((!g1030) & (g1160) & (g2149) & (!g2150) & (g2176) & (g2218)) + ((!g1030) & (g1160) & (g2149) & (g2150) & (!g2176) & (g2218)) + ((!g1030) & (g1160) & (g2149) & (g2150) & (g2176) & (g2218)) + ((g1030) & (!g1160) & (!g2149) & (!g2150) & (!g2176) & (!g2218)) + ((g1030) & (!g1160) & (!g2149) & (!g2150) & (g2176) & (!g2218)) + ((g1030) & (!g1160) & (!g2149) & (g2150) & (!g2176) & (!g2218)) + ((g1030) & (!g1160) & (g2149) & (!g2150) & (!g2176) & (g2218)) + ((g1030) & (!g1160) & (g2149) & (!g2150) & (g2176) & (g2218)) + ((g1030) & (!g1160) & (g2149) & (g2150) & (!g2176) & (g2218)) + ((g1030) & (!g1160) & (g2149) & (g2150) & (g2176) & (!g2218)) + ((g1030) & (!g1160) & (g2149) & (g2150) & (g2176) & (g2218)) + ((g1030) & (g1160) & (!g2149) & (!g2150) & (!g2176) & (!g2218)) + ((g1030) & (g1160) & (g2149) & (!g2150) & (!g2176) & (g2218)) + ((g1030) & (g1160) & (g2149) & (!g2150) & (g2176) & (!g2218)) + ((g1030) & (g1160) & (g2149) & (!g2150) & (g2176) & (g2218)) + ((g1030) & (g1160) & (g2149) & (g2150) & (!g2176) & (!g2218)) + ((g1030) & (g1160) & (g2149) & (g2150) & (!g2176) & (g2218)) + ((g1030) & (g1160) & (g2149) & (g2150) & (g2176) & (!g2218)) + ((g1030) & (g1160) & (g2149) & (g2150) & (g2176) & (g2218)));
	assign g2239 = (((!g1160) & (!g2150) & (g2176) & (!g2218)) + ((!g1160) & (g2150) & (!g2176) & (!g2218)) + ((!g1160) & (g2150) & (!g2176) & (g2218)) + ((!g1160) & (g2150) & (g2176) & (g2218)) + ((g1160) & (!g2150) & (!g2176) & (!g2218)) + ((g1160) & (g2150) & (!g2176) & (g2218)) + ((g1160) & (g2150) & (g2176) & (!g2218)) + ((g1160) & (g2150) & (g2176) & (g2218)));
	assign g2240 = (((!g1154) & (!g1295) & (!g2152) & (g2153) & (g2175) & (!g2218)) + ((!g1154) & (!g1295) & (g2152) & (!g2153) & (!g2175) & (!g2218)) + ((!g1154) & (!g1295) & (g2152) & (!g2153) & (!g2175) & (g2218)) + ((!g1154) & (!g1295) & (g2152) & (!g2153) & (g2175) & (!g2218)) + ((!g1154) & (!g1295) & (g2152) & (!g2153) & (g2175) & (g2218)) + ((!g1154) & (!g1295) & (g2152) & (g2153) & (!g2175) & (!g2218)) + ((!g1154) & (!g1295) & (g2152) & (g2153) & (!g2175) & (g2218)) + ((!g1154) & (!g1295) & (g2152) & (g2153) & (g2175) & (g2218)) + ((!g1154) & (g1295) & (!g2152) & (!g2153) & (g2175) & (!g2218)) + ((!g1154) & (g1295) & (!g2152) & (g2153) & (!g2175) & (!g2218)) + ((!g1154) & (g1295) & (!g2152) & (g2153) & (g2175) & (!g2218)) + ((!g1154) & (g1295) & (g2152) & (!g2153) & (!g2175) & (!g2218)) + ((!g1154) & (g1295) & (g2152) & (!g2153) & (!g2175) & (g2218)) + ((!g1154) & (g1295) & (g2152) & (!g2153) & (g2175) & (g2218)) + ((!g1154) & (g1295) & (g2152) & (g2153) & (!g2175) & (g2218)) + ((!g1154) & (g1295) & (g2152) & (g2153) & (g2175) & (g2218)) + ((g1154) & (!g1295) & (!g2152) & (!g2153) & (!g2175) & (!g2218)) + ((g1154) & (!g1295) & (!g2152) & (!g2153) & (g2175) & (!g2218)) + ((g1154) & (!g1295) & (!g2152) & (g2153) & (!g2175) & (!g2218)) + ((g1154) & (!g1295) & (g2152) & (!g2153) & (!g2175) & (g2218)) + ((g1154) & (!g1295) & (g2152) & (!g2153) & (g2175) & (g2218)) + ((g1154) & (!g1295) & (g2152) & (g2153) & (!g2175) & (g2218)) + ((g1154) & (!g1295) & (g2152) & (g2153) & (g2175) & (!g2218)) + ((g1154) & (!g1295) & (g2152) & (g2153) & (g2175) & (g2218)) + ((g1154) & (g1295) & (!g2152) & (!g2153) & (!g2175) & (!g2218)) + ((g1154) & (g1295) & (g2152) & (!g2153) & (!g2175) & (g2218)) + ((g1154) & (g1295) & (g2152) & (!g2153) & (g2175) & (!g2218)) + ((g1154) & (g1295) & (g2152) & (!g2153) & (g2175) & (g2218)) + ((g1154) & (g1295) & (g2152) & (g2153) & (!g2175) & (!g2218)) + ((g1154) & (g1295) & (g2152) & (g2153) & (!g2175) & (g2218)) + ((g1154) & (g1295) & (g2152) & (g2153) & (g2175) & (!g2218)) + ((g1154) & (g1295) & (g2152) & (g2153) & (g2175) & (g2218)));
	assign g2241 = (((!g1295) & (!g2153) & (g2175) & (!g2218)) + ((!g1295) & (g2153) & (!g2175) & (!g2218)) + ((!g1295) & (g2153) & (!g2175) & (g2218)) + ((!g1295) & (g2153) & (g2175) & (g2218)) + ((g1295) & (!g2153) & (!g2175) & (!g2218)) + ((g1295) & (g2153) & (!g2175) & (g2218)) + ((g1295) & (g2153) & (g2175) & (!g2218)) + ((g1295) & (g2153) & (g2175) & (g2218)));
	assign g2242 = (((!g1285) & (!g1437) & (!g2155) & (g2156) & (g2174) & (!g2218)) + ((!g1285) & (!g1437) & (g2155) & (!g2156) & (!g2174) & (!g2218)) + ((!g1285) & (!g1437) & (g2155) & (!g2156) & (!g2174) & (g2218)) + ((!g1285) & (!g1437) & (g2155) & (!g2156) & (g2174) & (!g2218)) + ((!g1285) & (!g1437) & (g2155) & (!g2156) & (g2174) & (g2218)) + ((!g1285) & (!g1437) & (g2155) & (g2156) & (!g2174) & (!g2218)) + ((!g1285) & (!g1437) & (g2155) & (g2156) & (!g2174) & (g2218)) + ((!g1285) & (!g1437) & (g2155) & (g2156) & (g2174) & (g2218)) + ((!g1285) & (g1437) & (!g2155) & (!g2156) & (g2174) & (!g2218)) + ((!g1285) & (g1437) & (!g2155) & (g2156) & (!g2174) & (!g2218)) + ((!g1285) & (g1437) & (!g2155) & (g2156) & (g2174) & (!g2218)) + ((!g1285) & (g1437) & (g2155) & (!g2156) & (!g2174) & (!g2218)) + ((!g1285) & (g1437) & (g2155) & (!g2156) & (!g2174) & (g2218)) + ((!g1285) & (g1437) & (g2155) & (!g2156) & (g2174) & (g2218)) + ((!g1285) & (g1437) & (g2155) & (g2156) & (!g2174) & (g2218)) + ((!g1285) & (g1437) & (g2155) & (g2156) & (g2174) & (g2218)) + ((g1285) & (!g1437) & (!g2155) & (!g2156) & (!g2174) & (!g2218)) + ((g1285) & (!g1437) & (!g2155) & (!g2156) & (g2174) & (!g2218)) + ((g1285) & (!g1437) & (!g2155) & (g2156) & (!g2174) & (!g2218)) + ((g1285) & (!g1437) & (g2155) & (!g2156) & (!g2174) & (g2218)) + ((g1285) & (!g1437) & (g2155) & (!g2156) & (g2174) & (g2218)) + ((g1285) & (!g1437) & (g2155) & (g2156) & (!g2174) & (g2218)) + ((g1285) & (!g1437) & (g2155) & (g2156) & (g2174) & (!g2218)) + ((g1285) & (!g1437) & (g2155) & (g2156) & (g2174) & (g2218)) + ((g1285) & (g1437) & (!g2155) & (!g2156) & (!g2174) & (!g2218)) + ((g1285) & (g1437) & (g2155) & (!g2156) & (!g2174) & (g2218)) + ((g1285) & (g1437) & (g2155) & (!g2156) & (g2174) & (!g2218)) + ((g1285) & (g1437) & (g2155) & (!g2156) & (g2174) & (g2218)) + ((g1285) & (g1437) & (g2155) & (g2156) & (!g2174) & (!g2218)) + ((g1285) & (g1437) & (g2155) & (g2156) & (!g2174) & (g2218)) + ((g1285) & (g1437) & (g2155) & (g2156) & (g2174) & (!g2218)) + ((g1285) & (g1437) & (g2155) & (g2156) & (g2174) & (g2218)));
	assign g2243 = (((!g1437) & (!g2156) & (g2174) & (!g2218)) + ((!g1437) & (g2156) & (!g2174) & (!g2218)) + ((!g1437) & (g2156) & (!g2174) & (g2218)) + ((!g1437) & (g2156) & (g2174) & (g2218)) + ((g1437) & (!g2156) & (!g2174) & (!g2218)) + ((g1437) & (g2156) & (!g2174) & (g2218)) + ((g1437) & (g2156) & (g2174) & (!g2218)) + ((g1437) & (g2156) & (g2174) & (g2218)));
	assign g2244 = (((!g1423) & (!g1586) & (!g2158) & (g2159) & (g2173) & (!g2218)) + ((!g1423) & (!g1586) & (g2158) & (!g2159) & (!g2173) & (!g2218)) + ((!g1423) & (!g1586) & (g2158) & (!g2159) & (!g2173) & (g2218)) + ((!g1423) & (!g1586) & (g2158) & (!g2159) & (g2173) & (!g2218)) + ((!g1423) & (!g1586) & (g2158) & (!g2159) & (g2173) & (g2218)) + ((!g1423) & (!g1586) & (g2158) & (g2159) & (!g2173) & (!g2218)) + ((!g1423) & (!g1586) & (g2158) & (g2159) & (!g2173) & (g2218)) + ((!g1423) & (!g1586) & (g2158) & (g2159) & (g2173) & (g2218)) + ((!g1423) & (g1586) & (!g2158) & (!g2159) & (g2173) & (!g2218)) + ((!g1423) & (g1586) & (!g2158) & (g2159) & (!g2173) & (!g2218)) + ((!g1423) & (g1586) & (!g2158) & (g2159) & (g2173) & (!g2218)) + ((!g1423) & (g1586) & (g2158) & (!g2159) & (!g2173) & (!g2218)) + ((!g1423) & (g1586) & (g2158) & (!g2159) & (!g2173) & (g2218)) + ((!g1423) & (g1586) & (g2158) & (!g2159) & (g2173) & (g2218)) + ((!g1423) & (g1586) & (g2158) & (g2159) & (!g2173) & (g2218)) + ((!g1423) & (g1586) & (g2158) & (g2159) & (g2173) & (g2218)) + ((g1423) & (!g1586) & (!g2158) & (!g2159) & (!g2173) & (!g2218)) + ((g1423) & (!g1586) & (!g2158) & (!g2159) & (g2173) & (!g2218)) + ((g1423) & (!g1586) & (!g2158) & (g2159) & (!g2173) & (!g2218)) + ((g1423) & (!g1586) & (g2158) & (!g2159) & (!g2173) & (g2218)) + ((g1423) & (!g1586) & (g2158) & (!g2159) & (g2173) & (g2218)) + ((g1423) & (!g1586) & (g2158) & (g2159) & (!g2173) & (g2218)) + ((g1423) & (!g1586) & (g2158) & (g2159) & (g2173) & (!g2218)) + ((g1423) & (!g1586) & (g2158) & (g2159) & (g2173) & (g2218)) + ((g1423) & (g1586) & (!g2158) & (!g2159) & (!g2173) & (!g2218)) + ((g1423) & (g1586) & (g2158) & (!g2159) & (!g2173) & (g2218)) + ((g1423) & (g1586) & (g2158) & (!g2159) & (g2173) & (!g2218)) + ((g1423) & (g1586) & (g2158) & (!g2159) & (g2173) & (g2218)) + ((g1423) & (g1586) & (g2158) & (g2159) & (!g2173) & (!g2218)) + ((g1423) & (g1586) & (g2158) & (g2159) & (!g2173) & (g2218)) + ((g1423) & (g1586) & (g2158) & (g2159) & (g2173) & (!g2218)) + ((g1423) & (g1586) & (g2158) & (g2159) & (g2173) & (g2218)));
	assign g2245 = (((!g1586) & (!g2159) & (g2173) & (!g2218)) + ((!g1586) & (g2159) & (!g2173) & (!g2218)) + ((!g1586) & (g2159) & (!g2173) & (g2218)) + ((!g1586) & (g2159) & (g2173) & (g2218)) + ((g1586) & (!g2159) & (!g2173) & (!g2218)) + ((g1586) & (g2159) & (!g2173) & (g2218)) + ((g1586) & (g2159) & (g2173) & (!g2218)) + ((g1586) & (g2159) & (g2173) & (g2218)));
	assign g2246 = (((!g1568) & (!g1742) & (!g2161) & (g2162) & (g2172) & (!g2218)) + ((!g1568) & (!g1742) & (g2161) & (!g2162) & (!g2172) & (!g2218)) + ((!g1568) & (!g1742) & (g2161) & (!g2162) & (!g2172) & (g2218)) + ((!g1568) & (!g1742) & (g2161) & (!g2162) & (g2172) & (!g2218)) + ((!g1568) & (!g1742) & (g2161) & (!g2162) & (g2172) & (g2218)) + ((!g1568) & (!g1742) & (g2161) & (g2162) & (!g2172) & (!g2218)) + ((!g1568) & (!g1742) & (g2161) & (g2162) & (!g2172) & (g2218)) + ((!g1568) & (!g1742) & (g2161) & (g2162) & (g2172) & (g2218)) + ((!g1568) & (g1742) & (!g2161) & (!g2162) & (g2172) & (!g2218)) + ((!g1568) & (g1742) & (!g2161) & (g2162) & (!g2172) & (!g2218)) + ((!g1568) & (g1742) & (!g2161) & (g2162) & (g2172) & (!g2218)) + ((!g1568) & (g1742) & (g2161) & (!g2162) & (!g2172) & (!g2218)) + ((!g1568) & (g1742) & (g2161) & (!g2162) & (!g2172) & (g2218)) + ((!g1568) & (g1742) & (g2161) & (!g2162) & (g2172) & (g2218)) + ((!g1568) & (g1742) & (g2161) & (g2162) & (!g2172) & (g2218)) + ((!g1568) & (g1742) & (g2161) & (g2162) & (g2172) & (g2218)) + ((g1568) & (!g1742) & (!g2161) & (!g2162) & (!g2172) & (!g2218)) + ((g1568) & (!g1742) & (!g2161) & (!g2162) & (g2172) & (!g2218)) + ((g1568) & (!g1742) & (!g2161) & (g2162) & (!g2172) & (!g2218)) + ((g1568) & (!g1742) & (g2161) & (!g2162) & (!g2172) & (g2218)) + ((g1568) & (!g1742) & (g2161) & (!g2162) & (g2172) & (g2218)) + ((g1568) & (!g1742) & (g2161) & (g2162) & (!g2172) & (g2218)) + ((g1568) & (!g1742) & (g2161) & (g2162) & (g2172) & (!g2218)) + ((g1568) & (!g1742) & (g2161) & (g2162) & (g2172) & (g2218)) + ((g1568) & (g1742) & (!g2161) & (!g2162) & (!g2172) & (!g2218)) + ((g1568) & (g1742) & (g2161) & (!g2162) & (!g2172) & (g2218)) + ((g1568) & (g1742) & (g2161) & (!g2162) & (g2172) & (!g2218)) + ((g1568) & (g1742) & (g2161) & (!g2162) & (g2172) & (g2218)) + ((g1568) & (g1742) & (g2161) & (g2162) & (!g2172) & (!g2218)) + ((g1568) & (g1742) & (g2161) & (g2162) & (!g2172) & (g2218)) + ((g1568) & (g1742) & (g2161) & (g2162) & (g2172) & (!g2218)) + ((g1568) & (g1742) & (g2161) & (g2162) & (g2172) & (g2218)));
	assign g2247 = (((!g1742) & (!g2162) & (g2172) & (!g2218)) + ((!g1742) & (g2162) & (!g2172) & (!g2218)) + ((!g1742) & (g2162) & (!g2172) & (g2218)) + ((!g1742) & (g2162) & (g2172) & (g2218)) + ((g1742) & (!g2162) & (!g2172) & (!g2218)) + ((g1742) & (g2162) & (!g2172) & (g2218)) + ((g1742) & (g2162) & (g2172) & (!g2218)) + ((g1742) & (g2162) & (g2172) & (g2218)));
	assign g2248 = (((!g1720) & (!g1905) & (!g2164) & (g2165) & (g2171) & (!g2218)) + ((!g1720) & (!g1905) & (g2164) & (!g2165) & (!g2171) & (!g2218)) + ((!g1720) & (!g1905) & (g2164) & (!g2165) & (!g2171) & (g2218)) + ((!g1720) & (!g1905) & (g2164) & (!g2165) & (g2171) & (!g2218)) + ((!g1720) & (!g1905) & (g2164) & (!g2165) & (g2171) & (g2218)) + ((!g1720) & (!g1905) & (g2164) & (g2165) & (!g2171) & (!g2218)) + ((!g1720) & (!g1905) & (g2164) & (g2165) & (!g2171) & (g2218)) + ((!g1720) & (!g1905) & (g2164) & (g2165) & (g2171) & (g2218)) + ((!g1720) & (g1905) & (!g2164) & (!g2165) & (g2171) & (!g2218)) + ((!g1720) & (g1905) & (!g2164) & (g2165) & (!g2171) & (!g2218)) + ((!g1720) & (g1905) & (!g2164) & (g2165) & (g2171) & (!g2218)) + ((!g1720) & (g1905) & (g2164) & (!g2165) & (!g2171) & (!g2218)) + ((!g1720) & (g1905) & (g2164) & (!g2165) & (!g2171) & (g2218)) + ((!g1720) & (g1905) & (g2164) & (!g2165) & (g2171) & (g2218)) + ((!g1720) & (g1905) & (g2164) & (g2165) & (!g2171) & (g2218)) + ((!g1720) & (g1905) & (g2164) & (g2165) & (g2171) & (g2218)) + ((g1720) & (!g1905) & (!g2164) & (!g2165) & (!g2171) & (!g2218)) + ((g1720) & (!g1905) & (!g2164) & (!g2165) & (g2171) & (!g2218)) + ((g1720) & (!g1905) & (!g2164) & (g2165) & (!g2171) & (!g2218)) + ((g1720) & (!g1905) & (g2164) & (!g2165) & (!g2171) & (g2218)) + ((g1720) & (!g1905) & (g2164) & (!g2165) & (g2171) & (g2218)) + ((g1720) & (!g1905) & (g2164) & (g2165) & (!g2171) & (g2218)) + ((g1720) & (!g1905) & (g2164) & (g2165) & (g2171) & (!g2218)) + ((g1720) & (!g1905) & (g2164) & (g2165) & (g2171) & (g2218)) + ((g1720) & (g1905) & (!g2164) & (!g2165) & (!g2171) & (!g2218)) + ((g1720) & (g1905) & (g2164) & (!g2165) & (!g2171) & (g2218)) + ((g1720) & (g1905) & (g2164) & (!g2165) & (g2171) & (!g2218)) + ((g1720) & (g1905) & (g2164) & (!g2165) & (g2171) & (g2218)) + ((g1720) & (g1905) & (g2164) & (g2165) & (!g2171) & (!g2218)) + ((g1720) & (g1905) & (g2164) & (g2165) & (!g2171) & (g2218)) + ((g1720) & (g1905) & (g2164) & (g2165) & (g2171) & (!g2218)) + ((g1720) & (g1905) & (g2164) & (g2165) & (g2171) & (g2218)));
	assign g2249 = (((!g1905) & (!g2165) & (g2171) & (!g2218)) + ((!g1905) & (g2165) & (!g2171) & (!g2218)) + ((!g1905) & (g2165) & (!g2171) & (g2218)) + ((!g1905) & (g2165) & (g2171) & (g2218)) + ((g1905) & (!g2165) & (!g2171) & (!g2218)) + ((g1905) & (g2165) & (!g2171) & (g2218)) + ((g1905) & (g2165) & (g2171) & (!g2218)) + ((g1905) & (g2165) & (g2171) & (g2218)));
	assign g2250 = (((!g1879) & (!g2075) & (!g2167) & (g2168) & (g2170) & (!g2218)) + ((!g1879) & (!g2075) & (g2167) & (!g2168) & (!g2170) & (!g2218)) + ((!g1879) & (!g2075) & (g2167) & (!g2168) & (!g2170) & (g2218)) + ((!g1879) & (!g2075) & (g2167) & (!g2168) & (g2170) & (!g2218)) + ((!g1879) & (!g2075) & (g2167) & (!g2168) & (g2170) & (g2218)) + ((!g1879) & (!g2075) & (g2167) & (g2168) & (!g2170) & (!g2218)) + ((!g1879) & (!g2075) & (g2167) & (g2168) & (!g2170) & (g2218)) + ((!g1879) & (!g2075) & (g2167) & (g2168) & (g2170) & (g2218)) + ((!g1879) & (g2075) & (!g2167) & (!g2168) & (g2170) & (!g2218)) + ((!g1879) & (g2075) & (!g2167) & (g2168) & (!g2170) & (!g2218)) + ((!g1879) & (g2075) & (!g2167) & (g2168) & (g2170) & (!g2218)) + ((!g1879) & (g2075) & (g2167) & (!g2168) & (!g2170) & (!g2218)) + ((!g1879) & (g2075) & (g2167) & (!g2168) & (!g2170) & (g2218)) + ((!g1879) & (g2075) & (g2167) & (!g2168) & (g2170) & (g2218)) + ((!g1879) & (g2075) & (g2167) & (g2168) & (!g2170) & (g2218)) + ((!g1879) & (g2075) & (g2167) & (g2168) & (g2170) & (g2218)) + ((g1879) & (!g2075) & (!g2167) & (!g2168) & (!g2170) & (!g2218)) + ((g1879) & (!g2075) & (!g2167) & (!g2168) & (g2170) & (!g2218)) + ((g1879) & (!g2075) & (!g2167) & (g2168) & (!g2170) & (!g2218)) + ((g1879) & (!g2075) & (g2167) & (!g2168) & (!g2170) & (g2218)) + ((g1879) & (!g2075) & (g2167) & (!g2168) & (g2170) & (g2218)) + ((g1879) & (!g2075) & (g2167) & (g2168) & (!g2170) & (g2218)) + ((g1879) & (!g2075) & (g2167) & (g2168) & (g2170) & (!g2218)) + ((g1879) & (!g2075) & (g2167) & (g2168) & (g2170) & (g2218)) + ((g1879) & (g2075) & (!g2167) & (!g2168) & (!g2170) & (!g2218)) + ((g1879) & (g2075) & (g2167) & (!g2168) & (!g2170) & (g2218)) + ((g1879) & (g2075) & (g2167) & (!g2168) & (g2170) & (!g2218)) + ((g1879) & (g2075) & (g2167) & (!g2168) & (g2170) & (g2218)) + ((g1879) & (g2075) & (g2167) & (g2168) & (!g2170) & (!g2218)) + ((g1879) & (g2075) & (g2167) & (g2168) & (!g2170) & (g2218)) + ((g1879) & (g2075) & (g2167) & (g2168) & (g2170) & (!g2218)) + ((g1879) & (g2075) & (g2167) & (g2168) & (g2170) & (g2218)));
	assign g2251 = (((!g2075) & (!g2168) & (g2170) & (!g2218)) + ((!g2075) & (g2168) & (!g2170) & (!g2218)) + ((!g2075) & (g2168) & (!g2170) & (g2218)) + ((!g2075) & (g2168) & (g2170) & (g2218)) + ((g2075) & (!g2168) & (!g2170) & (!g2218)) + ((g2075) & (g2168) & (!g2170) & (g2218)) + ((g2075) & (g2168) & (g2170) & (!g2218)) + ((g2075) & (g2168) & (g2170) & (g2218)));
	assign g2252 = (((!g2095) & (g2119)));
	assign g2253 = (((!g2045) & (!ax30x) & (!ax31x) & (!g2252) & (!g2169) & (g2218)) + ((!g2045) & (!ax30x) & (!ax31x) & (!g2252) & (g2169) & (!g2218)) + ((!g2045) & (!ax30x) & (!ax31x) & (!g2252) & (g2169) & (g2218)) + ((!g2045) & (!ax30x) & (!ax31x) & (g2252) & (!g2169) & (!g2218)) + ((!g2045) & (!ax30x) & (ax31x) & (!g2252) & (!g2169) & (!g2218)) + ((!g2045) & (!ax30x) & (ax31x) & (g2252) & (!g2169) & (g2218)) + ((!g2045) & (!ax30x) & (ax31x) & (g2252) & (g2169) & (!g2218)) + ((!g2045) & (!ax30x) & (ax31x) & (g2252) & (g2169) & (g2218)) + ((!g2045) & (ax30x) & (!ax31x) & (g2252) & (!g2169) & (!g2218)) + ((!g2045) & (ax30x) & (!ax31x) & (g2252) & (g2169) & (!g2218)) + ((!g2045) & (ax30x) & (ax31x) & (!g2252) & (!g2169) & (!g2218)) + ((!g2045) & (ax30x) & (ax31x) & (!g2252) & (!g2169) & (g2218)) + ((!g2045) & (ax30x) & (ax31x) & (!g2252) & (g2169) & (!g2218)) + ((!g2045) & (ax30x) & (ax31x) & (!g2252) & (g2169) & (g2218)) + ((!g2045) & (ax30x) & (ax31x) & (g2252) & (!g2169) & (g2218)) + ((!g2045) & (ax30x) & (ax31x) & (g2252) & (g2169) & (g2218)) + ((g2045) & (!ax30x) & (!ax31x) & (!g2252) & (!g2169) & (!g2218)) + ((g2045) & (!ax30x) & (!ax31x) & (!g2252) & (!g2169) & (g2218)) + ((g2045) & (!ax30x) & (!ax31x) & (!g2252) & (g2169) & (g2218)) + ((g2045) & (!ax30x) & (!ax31x) & (g2252) & (g2169) & (!g2218)) + ((g2045) & (!ax30x) & (ax31x) & (!g2252) & (g2169) & (!g2218)) + ((g2045) & (!ax30x) & (ax31x) & (g2252) & (!g2169) & (!g2218)) + ((g2045) & (!ax30x) & (ax31x) & (g2252) & (!g2169) & (g2218)) + ((g2045) & (!ax30x) & (ax31x) & (g2252) & (g2169) & (g2218)) + ((g2045) & (ax30x) & (!ax31x) & (!g2252) & (!g2169) & (!g2218)) + ((g2045) & (ax30x) & (!ax31x) & (!g2252) & (g2169) & (!g2218)) + ((g2045) & (ax30x) & (ax31x) & (!g2252) & (!g2169) & (g2218)) + ((g2045) & (ax30x) & (ax31x) & (!g2252) & (g2169) & (g2218)) + ((g2045) & (ax30x) & (ax31x) & (g2252) & (!g2169) & (!g2218)) + ((g2045) & (ax30x) & (ax31x) & (g2252) & (!g2169) & (g2218)) + ((g2045) & (ax30x) & (ax31x) & (g2252) & (g2169) & (!g2218)) + ((g2045) & (ax30x) & (ax31x) & (g2252) & (g2169) & (g2218)));
	assign g2254 = (((!ax30x) & (!g2252) & (!g2169) & (g2218)) + ((!ax30x) & (!g2252) & (g2169) & (!g2218)) + ((!ax30x) & (!g2252) & (g2169) & (g2218)) + ((!ax30x) & (g2252) & (g2169) & (!g2218)) + ((ax30x) & (!g2252) & (!g2169) & (!g2218)) + ((ax30x) & (g2252) & (!g2169) & (!g2218)) + ((ax30x) & (g2252) & (!g2169) & (g2218)) + ((ax30x) & (g2252) & (g2169) & (g2218)));
	assign g2255 = (((!ax26x) & (!ax27x)));
	assign g2256 = (((!g2252) & (!ax28x) & (!ax29x) & (!g2218) & (!g2255)) + ((!g2252) & (!ax28x) & (ax29x) & (g2218) & (!g2255)) + ((!g2252) & (ax28x) & (ax29x) & (g2218) & (!g2255)) + ((!g2252) & (ax28x) & (ax29x) & (g2218) & (g2255)) + ((g2252) & (!ax28x) & (!ax29x) & (!g2218) & (!g2255)) + ((g2252) & (!ax28x) & (!ax29x) & (!g2218) & (g2255)) + ((g2252) & (!ax28x) & (!ax29x) & (g2218) & (!g2255)) + ((g2252) & (!ax28x) & (ax29x) & (!g2218) & (!g2255)) + ((g2252) & (!ax28x) & (ax29x) & (g2218) & (!g2255)) + ((g2252) & (!ax28x) & (ax29x) & (g2218) & (g2255)) + ((g2252) & (ax28x) & (!ax29x) & (g2218) & (!g2255)) + ((g2252) & (ax28x) & (!ax29x) & (g2218) & (g2255)) + ((g2252) & (ax28x) & (ax29x) & (!g2218) & (!g2255)) + ((g2252) & (ax28x) & (ax29x) & (!g2218) & (g2255)) + ((g2252) & (ax28x) & (ax29x) & (g2218) & (!g2255)) + ((g2252) & (ax28x) & (ax29x) & (g2218) & (g2255)));
	assign g2257 = (((!g2075) & (!g2045) & (g2253) & (g2254) & (g2256)) + ((!g2075) & (g2045) & (g2253) & (!g2254) & (g2256)) + ((!g2075) & (g2045) & (g2253) & (g2254) & (!g2256)) + ((!g2075) & (g2045) & (g2253) & (g2254) & (g2256)) + ((g2075) & (!g2045) & (!g2253) & (g2254) & (g2256)) + ((g2075) & (!g2045) & (g2253) & (!g2254) & (!g2256)) + ((g2075) & (!g2045) & (g2253) & (!g2254) & (g2256)) + ((g2075) & (!g2045) & (g2253) & (g2254) & (!g2256)) + ((g2075) & (!g2045) & (g2253) & (g2254) & (g2256)) + ((g2075) & (g2045) & (!g2253) & (!g2254) & (g2256)) + ((g2075) & (g2045) & (!g2253) & (g2254) & (!g2256)) + ((g2075) & (g2045) & (!g2253) & (g2254) & (g2256)) + ((g2075) & (g2045) & (g2253) & (!g2254) & (!g2256)) + ((g2075) & (g2045) & (g2253) & (!g2254) & (g2256)) + ((g2075) & (g2045) & (g2253) & (g2254) & (!g2256)) + ((g2075) & (g2045) & (g2253) & (g2254) & (g2256)));
	assign g2258 = (((!g1905) & (!g1879) & (g2250) & (g2251) & (g2257)) + ((!g1905) & (g1879) & (g2250) & (!g2251) & (g2257)) + ((!g1905) & (g1879) & (g2250) & (g2251) & (!g2257)) + ((!g1905) & (g1879) & (g2250) & (g2251) & (g2257)) + ((g1905) & (!g1879) & (!g2250) & (g2251) & (g2257)) + ((g1905) & (!g1879) & (g2250) & (!g2251) & (!g2257)) + ((g1905) & (!g1879) & (g2250) & (!g2251) & (g2257)) + ((g1905) & (!g1879) & (g2250) & (g2251) & (!g2257)) + ((g1905) & (!g1879) & (g2250) & (g2251) & (g2257)) + ((g1905) & (g1879) & (!g2250) & (!g2251) & (g2257)) + ((g1905) & (g1879) & (!g2250) & (g2251) & (!g2257)) + ((g1905) & (g1879) & (!g2250) & (g2251) & (g2257)) + ((g1905) & (g1879) & (g2250) & (!g2251) & (!g2257)) + ((g1905) & (g1879) & (g2250) & (!g2251) & (g2257)) + ((g1905) & (g1879) & (g2250) & (g2251) & (!g2257)) + ((g1905) & (g1879) & (g2250) & (g2251) & (g2257)));
	assign g2259 = (((!g1742) & (!g1720) & (g2248) & (g2249) & (g2258)) + ((!g1742) & (g1720) & (g2248) & (!g2249) & (g2258)) + ((!g1742) & (g1720) & (g2248) & (g2249) & (!g2258)) + ((!g1742) & (g1720) & (g2248) & (g2249) & (g2258)) + ((g1742) & (!g1720) & (!g2248) & (g2249) & (g2258)) + ((g1742) & (!g1720) & (g2248) & (!g2249) & (!g2258)) + ((g1742) & (!g1720) & (g2248) & (!g2249) & (g2258)) + ((g1742) & (!g1720) & (g2248) & (g2249) & (!g2258)) + ((g1742) & (!g1720) & (g2248) & (g2249) & (g2258)) + ((g1742) & (g1720) & (!g2248) & (!g2249) & (g2258)) + ((g1742) & (g1720) & (!g2248) & (g2249) & (!g2258)) + ((g1742) & (g1720) & (!g2248) & (g2249) & (g2258)) + ((g1742) & (g1720) & (g2248) & (!g2249) & (!g2258)) + ((g1742) & (g1720) & (g2248) & (!g2249) & (g2258)) + ((g1742) & (g1720) & (g2248) & (g2249) & (!g2258)) + ((g1742) & (g1720) & (g2248) & (g2249) & (g2258)));
	assign g2260 = (((!g1586) & (!g1568) & (g2246) & (g2247) & (g2259)) + ((!g1586) & (g1568) & (g2246) & (!g2247) & (g2259)) + ((!g1586) & (g1568) & (g2246) & (g2247) & (!g2259)) + ((!g1586) & (g1568) & (g2246) & (g2247) & (g2259)) + ((g1586) & (!g1568) & (!g2246) & (g2247) & (g2259)) + ((g1586) & (!g1568) & (g2246) & (!g2247) & (!g2259)) + ((g1586) & (!g1568) & (g2246) & (!g2247) & (g2259)) + ((g1586) & (!g1568) & (g2246) & (g2247) & (!g2259)) + ((g1586) & (!g1568) & (g2246) & (g2247) & (g2259)) + ((g1586) & (g1568) & (!g2246) & (!g2247) & (g2259)) + ((g1586) & (g1568) & (!g2246) & (g2247) & (!g2259)) + ((g1586) & (g1568) & (!g2246) & (g2247) & (g2259)) + ((g1586) & (g1568) & (g2246) & (!g2247) & (!g2259)) + ((g1586) & (g1568) & (g2246) & (!g2247) & (g2259)) + ((g1586) & (g1568) & (g2246) & (g2247) & (!g2259)) + ((g1586) & (g1568) & (g2246) & (g2247) & (g2259)));
	assign g2261 = (((!g1437) & (!g1423) & (g2244) & (g2245) & (g2260)) + ((!g1437) & (g1423) & (g2244) & (!g2245) & (g2260)) + ((!g1437) & (g1423) & (g2244) & (g2245) & (!g2260)) + ((!g1437) & (g1423) & (g2244) & (g2245) & (g2260)) + ((g1437) & (!g1423) & (!g2244) & (g2245) & (g2260)) + ((g1437) & (!g1423) & (g2244) & (!g2245) & (!g2260)) + ((g1437) & (!g1423) & (g2244) & (!g2245) & (g2260)) + ((g1437) & (!g1423) & (g2244) & (g2245) & (!g2260)) + ((g1437) & (!g1423) & (g2244) & (g2245) & (g2260)) + ((g1437) & (g1423) & (!g2244) & (!g2245) & (g2260)) + ((g1437) & (g1423) & (!g2244) & (g2245) & (!g2260)) + ((g1437) & (g1423) & (!g2244) & (g2245) & (g2260)) + ((g1437) & (g1423) & (g2244) & (!g2245) & (!g2260)) + ((g1437) & (g1423) & (g2244) & (!g2245) & (g2260)) + ((g1437) & (g1423) & (g2244) & (g2245) & (!g2260)) + ((g1437) & (g1423) & (g2244) & (g2245) & (g2260)));
	assign g2262 = (((!g1295) & (!g1285) & (g2242) & (g2243) & (g2261)) + ((!g1295) & (g1285) & (g2242) & (!g2243) & (g2261)) + ((!g1295) & (g1285) & (g2242) & (g2243) & (!g2261)) + ((!g1295) & (g1285) & (g2242) & (g2243) & (g2261)) + ((g1295) & (!g1285) & (!g2242) & (g2243) & (g2261)) + ((g1295) & (!g1285) & (g2242) & (!g2243) & (!g2261)) + ((g1295) & (!g1285) & (g2242) & (!g2243) & (g2261)) + ((g1295) & (!g1285) & (g2242) & (g2243) & (!g2261)) + ((g1295) & (!g1285) & (g2242) & (g2243) & (g2261)) + ((g1295) & (g1285) & (!g2242) & (!g2243) & (g2261)) + ((g1295) & (g1285) & (!g2242) & (g2243) & (!g2261)) + ((g1295) & (g1285) & (!g2242) & (g2243) & (g2261)) + ((g1295) & (g1285) & (g2242) & (!g2243) & (!g2261)) + ((g1295) & (g1285) & (g2242) & (!g2243) & (g2261)) + ((g1295) & (g1285) & (g2242) & (g2243) & (!g2261)) + ((g1295) & (g1285) & (g2242) & (g2243) & (g2261)));
	assign g2263 = (((!g1160) & (!g1154) & (g2240) & (g2241) & (g2262)) + ((!g1160) & (g1154) & (g2240) & (!g2241) & (g2262)) + ((!g1160) & (g1154) & (g2240) & (g2241) & (!g2262)) + ((!g1160) & (g1154) & (g2240) & (g2241) & (g2262)) + ((g1160) & (!g1154) & (!g2240) & (g2241) & (g2262)) + ((g1160) & (!g1154) & (g2240) & (!g2241) & (!g2262)) + ((g1160) & (!g1154) & (g2240) & (!g2241) & (g2262)) + ((g1160) & (!g1154) & (g2240) & (g2241) & (!g2262)) + ((g1160) & (!g1154) & (g2240) & (g2241) & (g2262)) + ((g1160) & (g1154) & (!g2240) & (!g2241) & (g2262)) + ((g1160) & (g1154) & (!g2240) & (g2241) & (!g2262)) + ((g1160) & (g1154) & (!g2240) & (g2241) & (g2262)) + ((g1160) & (g1154) & (g2240) & (!g2241) & (!g2262)) + ((g1160) & (g1154) & (g2240) & (!g2241) & (g2262)) + ((g1160) & (g1154) & (g2240) & (g2241) & (!g2262)) + ((g1160) & (g1154) & (g2240) & (g2241) & (g2262)));
	assign g2264 = (((!g1032) & (!g1030) & (g2238) & (g2239) & (g2263)) + ((!g1032) & (g1030) & (g2238) & (!g2239) & (g2263)) + ((!g1032) & (g1030) & (g2238) & (g2239) & (!g2263)) + ((!g1032) & (g1030) & (g2238) & (g2239) & (g2263)) + ((g1032) & (!g1030) & (!g2238) & (g2239) & (g2263)) + ((g1032) & (!g1030) & (g2238) & (!g2239) & (!g2263)) + ((g1032) & (!g1030) & (g2238) & (!g2239) & (g2263)) + ((g1032) & (!g1030) & (g2238) & (g2239) & (!g2263)) + ((g1032) & (!g1030) & (g2238) & (g2239) & (g2263)) + ((g1032) & (g1030) & (!g2238) & (!g2239) & (g2263)) + ((g1032) & (g1030) & (!g2238) & (g2239) & (!g2263)) + ((g1032) & (g1030) & (!g2238) & (g2239) & (g2263)) + ((g1032) & (g1030) & (g2238) & (!g2239) & (!g2263)) + ((g1032) & (g1030) & (g2238) & (!g2239) & (g2263)) + ((g1032) & (g1030) & (g2238) & (g2239) & (!g2263)) + ((g1032) & (g1030) & (g2238) & (g2239) & (g2263)));
	assign g2265 = (((!g851) & (!g914) & (g2236) & (g2237) & (g2264)) + ((!g851) & (g914) & (g2236) & (!g2237) & (g2264)) + ((!g851) & (g914) & (g2236) & (g2237) & (!g2264)) + ((!g851) & (g914) & (g2236) & (g2237) & (g2264)) + ((g851) & (!g914) & (!g2236) & (g2237) & (g2264)) + ((g851) & (!g914) & (g2236) & (!g2237) & (!g2264)) + ((g851) & (!g914) & (g2236) & (!g2237) & (g2264)) + ((g851) & (!g914) & (g2236) & (g2237) & (!g2264)) + ((g851) & (!g914) & (g2236) & (g2237) & (g2264)) + ((g851) & (g914) & (!g2236) & (!g2237) & (g2264)) + ((g851) & (g914) & (!g2236) & (g2237) & (!g2264)) + ((g851) & (g914) & (!g2236) & (g2237) & (g2264)) + ((g851) & (g914) & (g2236) & (!g2237) & (!g2264)) + ((g851) & (g914) & (g2236) & (!g2237) & (g2264)) + ((g851) & (g914) & (g2236) & (g2237) & (!g2264)) + ((g851) & (g914) & (g2236) & (g2237) & (g2264)));
	assign g2266 = (((!g744) & (!g803) & (g2234) & (g2235) & (g2265)) + ((!g744) & (g803) & (g2234) & (!g2235) & (g2265)) + ((!g744) & (g803) & (g2234) & (g2235) & (!g2265)) + ((!g744) & (g803) & (g2234) & (g2235) & (g2265)) + ((g744) & (!g803) & (!g2234) & (g2235) & (g2265)) + ((g744) & (!g803) & (g2234) & (!g2235) & (!g2265)) + ((g744) & (!g803) & (g2234) & (!g2235) & (g2265)) + ((g744) & (!g803) & (g2234) & (g2235) & (!g2265)) + ((g744) & (!g803) & (g2234) & (g2235) & (g2265)) + ((g744) & (g803) & (!g2234) & (!g2235) & (g2265)) + ((g744) & (g803) & (!g2234) & (g2235) & (!g2265)) + ((g744) & (g803) & (!g2234) & (g2235) & (g2265)) + ((g744) & (g803) & (g2234) & (!g2235) & (!g2265)) + ((g744) & (g803) & (g2234) & (!g2235) & (g2265)) + ((g744) & (g803) & (g2234) & (g2235) & (!g2265)) + ((g744) & (g803) & (g2234) & (g2235) & (g2265)));
	assign g2267 = (((!g645) & (!g700) & (g2232) & (g2233) & (g2266)) + ((!g645) & (g700) & (g2232) & (!g2233) & (g2266)) + ((!g645) & (g700) & (g2232) & (g2233) & (!g2266)) + ((!g645) & (g700) & (g2232) & (g2233) & (g2266)) + ((g645) & (!g700) & (!g2232) & (g2233) & (g2266)) + ((g645) & (!g700) & (g2232) & (!g2233) & (!g2266)) + ((g645) & (!g700) & (g2232) & (!g2233) & (g2266)) + ((g645) & (!g700) & (g2232) & (g2233) & (!g2266)) + ((g645) & (!g700) & (g2232) & (g2233) & (g2266)) + ((g645) & (g700) & (!g2232) & (!g2233) & (g2266)) + ((g645) & (g700) & (!g2232) & (g2233) & (!g2266)) + ((g645) & (g700) & (!g2232) & (g2233) & (g2266)) + ((g645) & (g700) & (g2232) & (!g2233) & (!g2266)) + ((g645) & (g700) & (g2232) & (!g2233) & (g2266)) + ((g645) & (g700) & (g2232) & (g2233) & (!g2266)) + ((g645) & (g700) & (g2232) & (g2233) & (g2266)));
	assign g2268 = (((!g553) & (!g604) & (g2230) & (g2231) & (g2267)) + ((!g553) & (g604) & (g2230) & (!g2231) & (g2267)) + ((!g553) & (g604) & (g2230) & (g2231) & (!g2267)) + ((!g553) & (g604) & (g2230) & (g2231) & (g2267)) + ((g553) & (!g604) & (!g2230) & (g2231) & (g2267)) + ((g553) & (!g604) & (g2230) & (!g2231) & (!g2267)) + ((g553) & (!g604) & (g2230) & (!g2231) & (g2267)) + ((g553) & (!g604) & (g2230) & (g2231) & (!g2267)) + ((g553) & (!g604) & (g2230) & (g2231) & (g2267)) + ((g553) & (g604) & (!g2230) & (!g2231) & (g2267)) + ((g553) & (g604) & (!g2230) & (g2231) & (!g2267)) + ((g553) & (g604) & (!g2230) & (g2231) & (g2267)) + ((g553) & (g604) & (g2230) & (!g2231) & (!g2267)) + ((g553) & (g604) & (g2230) & (!g2231) & (g2267)) + ((g553) & (g604) & (g2230) & (g2231) & (!g2267)) + ((g553) & (g604) & (g2230) & (g2231) & (g2267)));
	assign g2269 = (((!g468) & (!g515) & (g2228) & (g2229) & (g2268)) + ((!g468) & (g515) & (g2228) & (!g2229) & (g2268)) + ((!g468) & (g515) & (g2228) & (g2229) & (!g2268)) + ((!g468) & (g515) & (g2228) & (g2229) & (g2268)) + ((g468) & (!g515) & (!g2228) & (g2229) & (g2268)) + ((g468) & (!g515) & (g2228) & (!g2229) & (!g2268)) + ((g468) & (!g515) & (g2228) & (!g2229) & (g2268)) + ((g468) & (!g515) & (g2228) & (g2229) & (!g2268)) + ((g468) & (!g515) & (g2228) & (g2229) & (g2268)) + ((g468) & (g515) & (!g2228) & (!g2229) & (g2268)) + ((g468) & (g515) & (!g2228) & (g2229) & (!g2268)) + ((g468) & (g515) & (!g2228) & (g2229) & (g2268)) + ((g468) & (g515) & (g2228) & (!g2229) & (!g2268)) + ((g468) & (g515) & (g2228) & (!g2229) & (g2268)) + ((g468) & (g515) & (g2228) & (g2229) & (!g2268)) + ((g468) & (g515) & (g2228) & (g2229) & (g2268)));
	assign g2270 = (((!g390) & (!g433) & (g2226) & (g2227) & (g2269)) + ((!g390) & (g433) & (g2226) & (!g2227) & (g2269)) + ((!g390) & (g433) & (g2226) & (g2227) & (!g2269)) + ((!g390) & (g433) & (g2226) & (g2227) & (g2269)) + ((g390) & (!g433) & (!g2226) & (g2227) & (g2269)) + ((g390) & (!g433) & (g2226) & (!g2227) & (!g2269)) + ((g390) & (!g433) & (g2226) & (!g2227) & (g2269)) + ((g390) & (!g433) & (g2226) & (g2227) & (!g2269)) + ((g390) & (!g433) & (g2226) & (g2227) & (g2269)) + ((g390) & (g433) & (!g2226) & (!g2227) & (g2269)) + ((g390) & (g433) & (!g2226) & (g2227) & (!g2269)) + ((g390) & (g433) & (!g2226) & (g2227) & (g2269)) + ((g390) & (g433) & (g2226) & (!g2227) & (!g2269)) + ((g390) & (g433) & (g2226) & (!g2227) & (g2269)) + ((g390) & (g433) & (g2226) & (g2227) & (!g2269)) + ((g390) & (g433) & (g2226) & (g2227) & (g2269)));
	assign g2271 = (((!g319) & (!g358) & (g2224) & (g2225) & (g2270)) + ((!g319) & (g358) & (g2224) & (!g2225) & (g2270)) + ((!g319) & (g358) & (g2224) & (g2225) & (!g2270)) + ((!g319) & (g358) & (g2224) & (g2225) & (g2270)) + ((g319) & (!g358) & (!g2224) & (g2225) & (g2270)) + ((g319) & (!g358) & (g2224) & (!g2225) & (!g2270)) + ((g319) & (!g358) & (g2224) & (!g2225) & (g2270)) + ((g319) & (!g358) & (g2224) & (g2225) & (!g2270)) + ((g319) & (!g358) & (g2224) & (g2225) & (g2270)) + ((g319) & (g358) & (!g2224) & (!g2225) & (g2270)) + ((g319) & (g358) & (!g2224) & (g2225) & (!g2270)) + ((g319) & (g358) & (!g2224) & (g2225) & (g2270)) + ((g319) & (g358) & (g2224) & (!g2225) & (!g2270)) + ((g319) & (g358) & (g2224) & (!g2225) & (g2270)) + ((g319) & (g358) & (g2224) & (g2225) & (!g2270)) + ((g319) & (g358) & (g2224) & (g2225) & (g2270)));
	assign g2272 = (((!g255) & (!g290) & (g2222) & (g2223) & (g2271)) + ((!g255) & (g290) & (g2222) & (!g2223) & (g2271)) + ((!g255) & (g290) & (g2222) & (g2223) & (!g2271)) + ((!g255) & (g290) & (g2222) & (g2223) & (g2271)) + ((g255) & (!g290) & (!g2222) & (g2223) & (g2271)) + ((g255) & (!g290) & (g2222) & (!g2223) & (!g2271)) + ((g255) & (!g290) & (g2222) & (!g2223) & (g2271)) + ((g255) & (!g290) & (g2222) & (g2223) & (!g2271)) + ((g255) & (!g290) & (g2222) & (g2223) & (g2271)) + ((g255) & (g290) & (!g2222) & (!g2223) & (g2271)) + ((g255) & (g290) & (!g2222) & (g2223) & (!g2271)) + ((g255) & (g290) & (!g2222) & (g2223) & (g2271)) + ((g255) & (g290) & (g2222) & (!g2223) & (!g2271)) + ((g255) & (g290) & (g2222) & (!g2223) & (g2271)) + ((g255) & (g290) & (g2222) & (g2223) & (!g2271)) + ((g255) & (g290) & (g2222) & (g2223) & (g2271)));
	assign g2273 = (((!g198) & (!g229) & (g2220) & (g2221) & (g2272)) + ((!g198) & (g229) & (g2220) & (!g2221) & (g2272)) + ((!g198) & (g229) & (g2220) & (g2221) & (!g2272)) + ((!g198) & (g229) & (g2220) & (g2221) & (g2272)) + ((g198) & (!g229) & (!g2220) & (g2221) & (g2272)) + ((g198) & (!g229) & (g2220) & (!g2221) & (!g2272)) + ((g198) & (!g229) & (g2220) & (!g2221) & (g2272)) + ((g198) & (!g229) & (g2220) & (g2221) & (!g2272)) + ((g198) & (!g229) & (g2220) & (g2221) & (g2272)) + ((g198) & (g229) & (!g2220) & (!g2221) & (g2272)) + ((g198) & (g229) & (!g2220) & (g2221) & (!g2272)) + ((g198) & (g229) & (!g2220) & (g2221) & (g2272)) + ((g198) & (g229) & (g2220) & (!g2221) & (!g2272)) + ((g198) & (g229) & (g2220) & (!g2221) & (g2272)) + ((g198) & (g229) & (g2220) & (g2221) & (!g2272)) + ((g198) & (g229) & (g2220) & (g2221) & (g2272)));
	assign g2274 = (((g1) & (!g2187) & (g2214) & (g2217)) + ((g1) & (g2187) & (!g2214) & (!g2217)) + ((g1) & (g2187) & (!g2214) & (g2217)));
	assign g2275 = (((!g4) & (!g2) & (!g2188) & (!g2211) & (!g2213) & (!g2218)) + ((!g4) & (!g2) & (!g2188) & (!g2211) & (g2213) & (g2218)) + ((!g4) & (!g2) & (!g2188) & (g2211) & (!g2213) & (!g2218)) + ((!g4) & (!g2) & (!g2188) & (g2211) & (g2213) & (g2218)) + ((!g4) & (!g2) & (g2188) & (!g2211) & (!g2213) & (!g2218)) + ((!g4) & (!g2) & (g2188) & (!g2211) & (g2213) & (g2218)) + ((!g4) & (!g2) & (g2188) & (g2211) & (g2213) & (!g2218)) + ((!g4) & (!g2) & (g2188) & (g2211) & (g2213) & (g2218)) + ((!g4) & (g2) & (!g2188) & (!g2211) & (!g2213) & (!g2218)) + ((!g4) & (g2) & (!g2188) & (!g2211) & (g2213) & (g2218)) + ((!g4) & (g2) & (!g2188) & (g2211) & (g2213) & (!g2218)) + ((!g4) & (g2) & (!g2188) & (g2211) & (g2213) & (g2218)) + ((!g4) & (g2) & (g2188) & (!g2211) & (g2213) & (!g2218)) + ((!g4) & (g2) & (g2188) & (!g2211) & (g2213) & (g2218)) + ((!g4) & (g2) & (g2188) & (g2211) & (g2213) & (!g2218)) + ((!g4) & (g2) & (g2188) & (g2211) & (g2213) & (g2218)) + ((g4) & (!g2) & (!g2188) & (!g2211) & (g2213) & (!g2218)) + ((g4) & (!g2) & (!g2188) & (!g2211) & (g2213) & (g2218)) + ((g4) & (!g2) & (!g2188) & (g2211) & (g2213) & (!g2218)) + ((g4) & (!g2) & (!g2188) & (g2211) & (g2213) & (g2218)) + ((g4) & (!g2) & (g2188) & (!g2211) & (g2213) & (!g2218)) + ((g4) & (!g2) & (g2188) & (!g2211) & (g2213) & (g2218)) + ((g4) & (!g2) & (g2188) & (g2211) & (!g2213) & (!g2218)) + ((g4) & (!g2) & (g2188) & (g2211) & (g2213) & (g2218)) + ((g4) & (g2) & (!g2188) & (!g2211) & (g2213) & (!g2218)) + ((g4) & (g2) & (!g2188) & (!g2211) & (g2213) & (g2218)) + ((g4) & (g2) & (!g2188) & (g2211) & (!g2213) & (!g2218)) + ((g4) & (g2) & (!g2188) & (g2211) & (g2213) & (g2218)) + ((g4) & (g2) & (g2188) & (!g2211) & (!g2213) & (!g2218)) + ((g4) & (g2) & (g2188) & (!g2211) & (g2213) & (g2218)) + ((g4) & (g2) & (g2188) & (g2211) & (!g2213) & (!g2218)) + ((g4) & (g2) & (g2188) & (g2211) & (g2213) & (g2218)));
	assign g2276 = (((!g8) & (!g18) & (!g2190) & (g2191) & (g2210) & (!g2218)) + ((!g8) & (!g18) & (g2190) & (!g2191) & (!g2210) & (!g2218)) + ((!g8) & (!g18) & (g2190) & (!g2191) & (!g2210) & (g2218)) + ((!g8) & (!g18) & (g2190) & (!g2191) & (g2210) & (!g2218)) + ((!g8) & (!g18) & (g2190) & (!g2191) & (g2210) & (g2218)) + ((!g8) & (!g18) & (g2190) & (g2191) & (!g2210) & (!g2218)) + ((!g8) & (!g18) & (g2190) & (g2191) & (!g2210) & (g2218)) + ((!g8) & (!g18) & (g2190) & (g2191) & (g2210) & (g2218)) + ((!g8) & (g18) & (!g2190) & (!g2191) & (g2210) & (!g2218)) + ((!g8) & (g18) & (!g2190) & (g2191) & (!g2210) & (!g2218)) + ((!g8) & (g18) & (!g2190) & (g2191) & (g2210) & (!g2218)) + ((!g8) & (g18) & (g2190) & (!g2191) & (!g2210) & (!g2218)) + ((!g8) & (g18) & (g2190) & (!g2191) & (!g2210) & (g2218)) + ((!g8) & (g18) & (g2190) & (!g2191) & (g2210) & (g2218)) + ((!g8) & (g18) & (g2190) & (g2191) & (!g2210) & (g2218)) + ((!g8) & (g18) & (g2190) & (g2191) & (g2210) & (g2218)) + ((g8) & (!g18) & (!g2190) & (!g2191) & (!g2210) & (!g2218)) + ((g8) & (!g18) & (!g2190) & (!g2191) & (g2210) & (!g2218)) + ((g8) & (!g18) & (!g2190) & (g2191) & (!g2210) & (!g2218)) + ((g8) & (!g18) & (g2190) & (!g2191) & (!g2210) & (g2218)) + ((g8) & (!g18) & (g2190) & (!g2191) & (g2210) & (g2218)) + ((g8) & (!g18) & (g2190) & (g2191) & (!g2210) & (g2218)) + ((g8) & (!g18) & (g2190) & (g2191) & (g2210) & (!g2218)) + ((g8) & (!g18) & (g2190) & (g2191) & (g2210) & (g2218)) + ((g8) & (g18) & (!g2190) & (!g2191) & (!g2210) & (!g2218)) + ((g8) & (g18) & (g2190) & (!g2191) & (!g2210) & (g2218)) + ((g8) & (g18) & (g2190) & (!g2191) & (g2210) & (!g2218)) + ((g8) & (g18) & (g2190) & (!g2191) & (g2210) & (g2218)) + ((g8) & (g18) & (g2190) & (g2191) & (!g2210) & (!g2218)) + ((g8) & (g18) & (g2190) & (g2191) & (!g2210) & (g2218)) + ((g8) & (g18) & (g2190) & (g2191) & (g2210) & (!g2218)) + ((g8) & (g18) & (g2190) & (g2191) & (g2210) & (g2218)));
	assign g2277 = (((!g18) & (!g2191) & (g2210) & (!g2218)) + ((!g18) & (g2191) & (!g2210) & (!g2218)) + ((!g18) & (g2191) & (!g2210) & (g2218)) + ((!g18) & (g2191) & (g2210) & (g2218)) + ((g18) & (!g2191) & (!g2210) & (!g2218)) + ((g18) & (g2191) & (!g2210) & (g2218)) + ((g18) & (g2191) & (g2210) & (!g2218)) + ((g18) & (g2191) & (g2210) & (g2218)));
	assign g2278 = (((!g27) & (!g39) & (!g2193) & (g2194) & (g2209) & (!g2218)) + ((!g27) & (!g39) & (g2193) & (!g2194) & (!g2209) & (!g2218)) + ((!g27) & (!g39) & (g2193) & (!g2194) & (!g2209) & (g2218)) + ((!g27) & (!g39) & (g2193) & (!g2194) & (g2209) & (!g2218)) + ((!g27) & (!g39) & (g2193) & (!g2194) & (g2209) & (g2218)) + ((!g27) & (!g39) & (g2193) & (g2194) & (!g2209) & (!g2218)) + ((!g27) & (!g39) & (g2193) & (g2194) & (!g2209) & (g2218)) + ((!g27) & (!g39) & (g2193) & (g2194) & (g2209) & (g2218)) + ((!g27) & (g39) & (!g2193) & (!g2194) & (g2209) & (!g2218)) + ((!g27) & (g39) & (!g2193) & (g2194) & (!g2209) & (!g2218)) + ((!g27) & (g39) & (!g2193) & (g2194) & (g2209) & (!g2218)) + ((!g27) & (g39) & (g2193) & (!g2194) & (!g2209) & (!g2218)) + ((!g27) & (g39) & (g2193) & (!g2194) & (!g2209) & (g2218)) + ((!g27) & (g39) & (g2193) & (!g2194) & (g2209) & (g2218)) + ((!g27) & (g39) & (g2193) & (g2194) & (!g2209) & (g2218)) + ((!g27) & (g39) & (g2193) & (g2194) & (g2209) & (g2218)) + ((g27) & (!g39) & (!g2193) & (!g2194) & (!g2209) & (!g2218)) + ((g27) & (!g39) & (!g2193) & (!g2194) & (g2209) & (!g2218)) + ((g27) & (!g39) & (!g2193) & (g2194) & (!g2209) & (!g2218)) + ((g27) & (!g39) & (g2193) & (!g2194) & (!g2209) & (g2218)) + ((g27) & (!g39) & (g2193) & (!g2194) & (g2209) & (g2218)) + ((g27) & (!g39) & (g2193) & (g2194) & (!g2209) & (g2218)) + ((g27) & (!g39) & (g2193) & (g2194) & (g2209) & (!g2218)) + ((g27) & (!g39) & (g2193) & (g2194) & (g2209) & (g2218)) + ((g27) & (g39) & (!g2193) & (!g2194) & (!g2209) & (!g2218)) + ((g27) & (g39) & (g2193) & (!g2194) & (!g2209) & (g2218)) + ((g27) & (g39) & (g2193) & (!g2194) & (g2209) & (!g2218)) + ((g27) & (g39) & (g2193) & (!g2194) & (g2209) & (g2218)) + ((g27) & (g39) & (g2193) & (g2194) & (!g2209) & (!g2218)) + ((g27) & (g39) & (g2193) & (g2194) & (!g2209) & (g2218)) + ((g27) & (g39) & (g2193) & (g2194) & (g2209) & (!g2218)) + ((g27) & (g39) & (g2193) & (g2194) & (g2209) & (g2218)));
	assign g2279 = (((!g39) & (!g2194) & (g2209) & (!g2218)) + ((!g39) & (g2194) & (!g2209) & (!g2218)) + ((!g39) & (g2194) & (!g2209) & (g2218)) + ((!g39) & (g2194) & (g2209) & (g2218)) + ((g39) & (!g2194) & (!g2209) & (!g2218)) + ((g39) & (g2194) & (!g2209) & (g2218)) + ((g39) & (g2194) & (g2209) & (!g2218)) + ((g39) & (g2194) & (g2209) & (g2218)));
	assign g2280 = (((!g54) & (!g68) & (!g2196) & (g2197) & (g2208) & (!g2218)) + ((!g54) & (!g68) & (g2196) & (!g2197) & (!g2208) & (!g2218)) + ((!g54) & (!g68) & (g2196) & (!g2197) & (!g2208) & (g2218)) + ((!g54) & (!g68) & (g2196) & (!g2197) & (g2208) & (!g2218)) + ((!g54) & (!g68) & (g2196) & (!g2197) & (g2208) & (g2218)) + ((!g54) & (!g68) & (g2196) & (g2197) & (!g2208) & (!g2218)) + ((!g54) & (!g68) & (g2196) & (g2197) & (!g2208) & (g2218)) + ((!g54) & (!g68) & (g2196) & (g2197) & (g2208) & (g2218)) + ((!g54) & (g68) & (!g2196) & (!g2197) & (g2208) & (!g2218)) + ((!g54) & (g68) & (!g2196) & (g2197) & (!g2208) & (!g2218)) + ((!g54) & (g68) & (!g2196) & (g2197) & (g2208) & (!g2218)) + ((!g54) & (g68) & (g2196) & (!g2197) & (!g2208) & (!g2218)) + ((!g54) & (g68) & (g2196) & (!g2197) & (!g2208) & (g2218)) + ((!g54) & (g68) & (g2196) & (!g2197) & (g2208) & (g2218)) + ((!g54) & (g68) & (g2196) & (g2197) & (!g2208) & (g2218)) + ((!g54) & (g68) & (g2196) & (g2197) & (g2208) & (g2218)) + ((g54) & (!g68) & (!g2196) & (!g2197) & (!g2208) & (!g2218)) + ((g54) & (!g68) & (!g2196) & (!g2197) & (g2208) & (!g2218)) + ((g54) & (!g68) & (!g2196) & (g2197) & (!g2208) & (!g2218)) + ((g54) & (!g68) & (g2196) & (!g2197) & (!g2208) & (g2218)) + ((g54) & (!g68) & (g2196) & (!g2197) & (g2208) & (g2218)) + ((g54) & (!g68) & (g2196) & (g2197) & (!g2208) & (g2218)) + ((g54) & (!g68) & (g2196) & (g2197) & (g2208) & (!g2218)) + ((g54) & (!g68) & (g2196) & (g2197) & (g2208) & (g2218)) + ((g54) & (g68) & (!g2196) & (!g2197) & (!g2208) & (!g2218)) + ((g54) & (g68) & (g2196) & (!g2197) & (!g2208) & (g2218)) + ((g54) & (g68) & (g2196) & (!g2197) & (g2208) & (!g2218)) + ((g54) & (g68) & (g2196) & (!g2197) & (g2208) & (g2218)) + ((g54) & (g68) & (g2196) & (g2197) & (!g2208) & (!g2218)) + ((g54) & (g68) & (g2196) & (g2197) & (!g2208) & (g2218)) + ((g54) & (g68) & (g2196) & (g2197) & (g2208) & (!g2218)) + ((g54) & (g68) & (g2196) & (g2197) & (g2208) & (g2218)));
	assign g2281 = (((!g68) & (!g2197) & (g2208) & (!g2218)) + ((!g68) & (g2197) & (!g2208) & (!g2218)) + ((!g68) & (g2197) & (!g2208) & (g2218)) + ((!g68) & (g2197) & (g2208) & (g2218)) + ((g68) & (!g2197) & (!g2208) & (!g2218)) + ((g68) & (g2197) & (!g2208) & (g2218)) + ((g68) & (g2197) & (g2208) & (!g2218)) + ((g68) & (g2197) & (g2208) & (g2218)));
	assign g2282 = (((!g87) & (!g104) & (!g2199) & (g2200) & (g2207) & (!g2218)) + ((!g87) & (!g104) & (g2199) & (!g2200) & (!g2207) & (!g2218)) + ((!g87) & (!g104) & (g2199) & (!g2200) & (!g2207) & (g2218)) + ((!g87) & (!g104) & (g2199) & (!g2200) & (g2207) & (!g2218)) + ((!g87) & (!g104) & (g2199) & (!g2200) & (g2207) & (g2218)) + ((!g87) & (!g104) & (g2199) & (g2200) & (!g2207) & (!g2218)) + ((!g87) & (!g104) & (g2199) & (g2200) & (!g2207) & (g2218)) + ((!g87) & (!g104) & (g2199) & (g2200) & (g2207) & (g2218)) + ((!g87) & (g104) & (!g2199) & (!g2200) & (g2207) & (!g2218)) + ((!g87) & (g104) & (!g2199) & (g2200) & (!g2207) & (!g2218)) + ((!g87) & (g104) & (!g2199) & (g2200) & (g2207) & (!g2218)) + ((!g87) & (g104) & (g2199) & (!g2200) & (!g2207) & (!g2218)) + ((!g87) & (g104) & (g2199) & (!g2200) & (!g2207) & (g2218)) + ((!g87) & (g104) & (g2199) & (!g2200) & (g2207) & (g2218)) + ((!g87) & (g104) & (g2199) & (g2200) & (!g2207) & (g2218)) + ((!g87) & (g104) & (g2199) & (g2200) & (g2207) & (g2218)) + ((g87) & (!g104) & (!g2199) & (!g2200) & (!g2207) & (!g2218)) + ((g87) & (!g104) & (!g2199) & (!g2200) & (g2207) & (!g2218)) + ((g87) & (!g104) & (!g2199) & (g2200) & (!g2207) & (!g2218)) + ((g87) & (!g104) & (g2199) & (!g2200) & (!g2207) & (g2218)) + ((g87) & (!g104) & (g2199) & (!g2200) & (g2207) & (g2218)) + ((g87) & (!g104) & (g2199) & (g2200) & (!g2207) & (g2218)) + ((g87) & (!g104) & (g2199) & (g2200) & (g2207) & (!g2218)) + ((g87) & (!g104) & (g2199) & (g2200) & (g2207) & (g2218)) + ((g87) & (g104) & (!g2199) & (!g2200) & (!g2207) & (!g2218)) + ((g87) & (g104) & (g2199) & (!g2200) & (!g2207) & (g2218)) + ((g87) & (g104) & (g2199) & (!g2200) & (g2207) & (!g2218)) + ((g87) & (g104) & (g2199) & (!g2200) & (g2207) & (g2218)) + ((g87) & (g104) & (g2199) & (g2200) & (!g2207) & (!g2218)) + ((g87) & (g104) & (g2199) & (g2200) & (!g2207) & (g2218)) + ((g87) & (g104) & (g2199) & (g2200) & (g2207) & (!g2218)) + ((g87) & (g104) & (g2199) & (g2200) & (g2207) & (g2218)));
	assign g2283 = (((!g104) & (!g2200) & (g2207) & (!g2218)) + ((!g104) & (g2200) & (!g2207) & (!g2218)) + ((!g104) & (g2200) & (!g2207) & (g2218)) + ((!g104) & (g2200) & (g2207) & (g2218)) + ((g104) & (!g2200) & (!g2207) & (!g2218)) + ((g104) & (g2200) & (!g2207) & (g2218)) + ((g104) & (g2200) & (g2207) & (!g2218)) + ((g104) & (g2200) & (g2207) & (g2218)));
	assign g2284 = (((!g127) & (!g147) & (!g2202) & (g2203) & (g2206) & (!g2218)) + ((!g127) & (!g147) & (g2202) & (!g2203) & (!g2206) & (!g2218)) + ((!g127) & (!g147) & (g2202) & (!g2203) & (!g2206) & (g2218)) + ((!g127) & (!g147) & (g2202) & (!g2203) & (g2206) & (!g2218)) + ((!g127) & (!g147) & (g2202) & (!g2203) & (g2206) & (g2218)) + ((!g127) & (!g147) & (g2202) & (g2203) & (!g2206) & (!g2218)) + ((!g127) & (!g147) & (g2202) & (g2203) & (!g2206) & (g2218)) + ((!g127) & (!g147) & (g2202) & (g2203) & (g2206) & (g2218)) + ((!g127) & (g147) & (!g2202) & (!g2203) & (g2206) & (!g2218)) + ((!g127) & (g147) & (!g2202) & (g2203) & (!g2206) & (!g2218)) + ((!g127) & (g147) & (!g2202) & (g2203) & (g2206) & (!g2218)) + ((!g127) & (g147) & (g2202) & (!g2203) & (!g2206) & (!g2218)) + ((!g127) & (g147) & (g2202) & (!g2203) & (!g2206) & (g2218)) + ((!g127) & (g147) & (g2202) & (!g2203) & (g2206) & (g2218)) + ((!g127) & (g147) & (g2202) & (g2203) & (!g2206) & (g2218)) + ((!g127) & (g147) & (g2202) & (g2203) & (g2206) & (g2218)) + ((g127) & (!g147) & (!g2202) & (!g2203) & (!g2206) & (!g2218)) + ((g127) & (!g147) & (!g2202) & (!g2203) & (g2206) & (!g2218)) + ((g127) & (!g147) & (!g2202) & (g2203) & (!g2206) & (!g2218)) + ((g127) & (!g147) & (g2202) & (!g2203) & (!g2206) & (g2218)) + ((g127) & (!g147) & (g2202) & (!g2203) & (g2206) & (g2218)) + ((g127) & (!g147) & (g2202) & (g2203) & (!g2206) & (g2218)) + ((g127) & (!g147) & (g2202) & (g2203) & (g2206) & (!g2218)) + ((g127) & (!g147) & (g2202) & (g2203) & (g2206) & (g2218)) + ((g127) & (g147) & (!g2202) & (!g2203) & (!g2206) & (!g2218)) + ((g127) & (g147) & (g2202) & (!g2203) & (!g2206) & (g2218)) + ((g127) & (g147) & (g2202) & (!g2203) & (g2206) & (!g2218)) + ((g127) & (g147) & (g2202) & (!g2203) & (g2206) & (g2218)) + ((g127) & (g147) & (g2202) & (g2203) & (!g2206) & (!g2218)) + ((g127) & (g147) & (g2202) & (g2203) & (!g2206) & (g2218)) + ((g127) & (g147) & (g2202) & (g2203) & (g2206) & (!g2218)) + ((g127) & (g147) & (g2202) & (g2203) & (g2206) & (g2218)));
	assign g2285 = (((!g147) & (!g2203) & (g2206) & (!g2218)) + ((!g147) & (g2203) & (!g2206) & (!g2218)) + ((!g147) & (g2203) & (!g2206) & (g2218)) + ((!g147) & (g2203) & (g2206) & (g2218)) + ((g147) & (!g2203) & (!g2206) & (!g2218)) + ((g147) & (g2203) & (!g2206) & (g2218)) + ((g147) & (g2203) & (g2206) & (!g2218)) + ((g147) & (g2203) & (g2206) & (g2218)));
	assign g2286 = (((!g174) & (!g198) & (!g2205) & (g2120) & (g2186) & (!g2218)) + ((!g174) & (!g198) & (g2205) & (!g2120) & (!g2186) & (!g2218)) + ((!g174) & (!g198) & (g2205) & (!g2120) & (!g2186) & (g2218)) + ((!g174) & (!g198) & (g2205) & (!g2120) & (g2186) & (!g2218)) + ((!g174) & (!g198) & (g2205) & (!g2120) & (g2186) & (g2218)) + ((!g174) & (!g198) & (g2205) & (g2120) & (!g2186) & (!g2218)) + ((!g174) & (!g198) & (g2205) & (g2120) & (!g2186) & (g2218)) + ((!g174) & (!g198) & (g2205) & (g2120) & (g2186) & (g2218)) + ((!g174) & (g198) & (!g2205) & (!g2120) & (g2186) & (!g2218)) + ((!g174) & (g198) & (!g2205) & (g2120) & (!g2186) & (!g2218)) + ((!g174) & (g198) & (!g2205) & (g2120) & (g2186) & (!g2218)) + ((!g174) & (g198) & (g2205) & (!g2120) & (!g2186) & (!g2218)) + ((!g174) & (g198) & (g2205) & (!g2120) & (!g2186) & (g2218)) + ((!g174) & (g198) & (g2205) & (!g2120) & (g2186) & (g2218)) + ((!g174) & (g198) & (g2205) & (g2120) & (!g2186) & (g2218)) + ((!g174) & (g198) & (g2205) & (g2120) & (g2186) & (g2218)) + ((g174) & (!g198) & (!g2205) & (!g2120) & (!g2186) & (!g2218)) + ((g174) & (!g198) & (!g2205) & (!g2120) & (g2186) & (!g2218)) + ((g174) & (!g198) & (!g2205) & (g2120) & (!g2186) & (!g2218)) + ((g174) & (!g198) & (g2205) & (!g2120) & (!g2186) & (g2218)) + ((g174) & (!g198) & (g2205) & (!g2120) & (g2186) & (g2218)) + ((g174) & (!g198) & (g2205) & (g2120) & (!g2186) & (g2218)) + ((g174) & (!g198) & (g2205) & (g2120) & (g2186) & (!g2218)) + ((g174) & (!g198) & (g2205) & (g2120) & (g2186) & (g2218)) + ((g174) & (g198) & (!g2205) & (!g2120) & (!g2186) & (!g2218)) + ((g174) & (g198) & (g2205) & (!g2120) & (!g2186) & (g2218)) + ((g174) & (g198) & (g2205) & (!g2120) & (g2186) & (!g2218)) + ((g174) & (g198) & (g2205) & (!g2120) & (g2186) & (g2218)) + ((g174) & (g198) & (g2205) & (g2120) & (!g2186) & (!g2218)) + ((g174) & (g198) & (g2205) & (g2120) & (!g2186) & (g2218)) + ((g174) & (g198) & (g2205) & (g2120) & (g2186) & (!g2218)) + ((g174) & (g198) & (g2205) & (g2120) & (g2186) & (g2218)));
	assign g2287 = (((!g147) & (!g174) & (g2286) & (g2219) & (g2273)) + ((!g147) & (g174) & (g2286) & (!g2219) & (g2273)) + ((!g147) & (g174) & (g2286) & (g2219) & (!g2273)) + ((!g147) & (g174) & (g2286) & (g2219) & (g2273)) + ((g147) & (!g174) & (!g2286) & (g2219) & (g2273)) + ((g147) & (!g174) & (g2286) & (!g2219) & (!g2273)) + ((g147) & (!g174) & (g2286) & (!g2219) & (g2273)) + ((g147) & (!g174) & (g2286) & (g2219) & (!g2273)) + ((g147) & (!g174) & (g2286) & (g2219) & (g2273)) + ((g147) & (g174) & (!g2286) & (!g2219) & (g2273)) + ((g147) & (g174) & (!g2286) & (g2219) & (!g2273)) + ((g147) & (g174) & (!g2286) & (g2219) & (g2273)) + ((g147) & (g174) & (g2286) & (!g2219) & (!g2273)) + ((g147) & (g174) & (g2286) & (!g2219) & (g2273)) + ((g147) & (g174) & (g2286) & (g2219) & (!g2273)) + ((g147) & (g174) & (g2286) & (g2219) & (g2273)));
	assign g2288 = (((!g104) & (!g127) & (g2284) & (g2285) & (g2287)) + ((!g104) & (g127) & (g2284) & (!g2285) & (g2287)) + ((!g104) & (g127) & (g2284) & (g2285) & (!g2287)) + ((!g104) & (g127) & (g2284) & (g2285) & (g2287)) + ((g104) & (!g127) & (!g2284) & (g2285) & (g2287)) + ((g104) & (!g127) & (g2284) & (!g2285) & (!g2287)) + ((g104) & (!g127) & (g2284) & (!g2285) & (g2287)) + ((g104) & (!g127) & (g2284) & (g2285) & (!g2287)) + ((g104) & (!g127) & (g2284) & (g2285) & (g2287)) + ((g104) & (g127) & (!g2284) & (!g2285) & (g2287)) + ((g104) & (g127) & (!g2284) & (g2285) & (!g2287)) + ((g104) & (g127) & (!g2284) & (g2285) & (g2287)) + ((g104) & (g127) & (g2284) & (!g2285) & (!g2287)) + ((g104) & (g127) & (g2284) & (!g2285) & (g2287)) + ((g104) & (g127) & (g2284) & (g2285) & (!g2287)) + ((g104) & (g127) & (g2284) & (g2285) & (g2287)));
	assign g2289 = (((!g68) & (!g87) & (g2282) & (g2283) & (g2288)) + ((!g68) & (g87) & (g2282) & (!g2283) & (g2288)) + ((!g68) & (g87) & (g2282) & (g2283) & (!g2288)) + ((!g68) & (g87) & (g2282) & (g2283) & (g2288)) + ((g68) & (!g87) & (!g2282) & (g2283) & (g2288)) + ((g68) & (!g87) & (g2282) & (!g2283) & (!g2288)) + ((g68) & (!g87) & (g2282) & (!g2283) & (g2288)) + ((g68) & (!g87) & (g2282) & (g2283) & (!g2288)) + ((g68) & (!g87) & (g2282) & (g2283) & (g2288)) + ((g68) & (g87) & (!g2282) & (!g2283) & (g2288)) + ((g68) & (g87) & (!g2282) & (g2283) & (!g2288)) + ((g68) & (g87) & (!g2282) & (g2283) & (g2288)) + ((g68) & (g87) & (g2282) & (!g2283) & (!g2288)) + ((g68) & (g87) & (g2282) & (!g2283) & (g2288)) + ((g68) & (g87) & (g2282) & (g2283) & (!g2288)) + ((g68) & (g87) & (g2282) & (g2283) & (g2288)));
	assign g2290 = (((!g39) & (!g54) & (g2280) & (g2281) & (g2289)) + ((!g39) & (g54) & (g2280) & (!g2281) & (g2289)) + ((!g39) & (g54) & (g2280) & (g2281) & (!g2289)) + ((!g39) & (g54) & (g2280) & (g2281) & (g2289)) + ((g39) & (!g54) & (!g2280) & (g2281) & (g2289)) + ((g39) & (!g54) & (g2280) & (!g2281) & (!g2289)) + ((g39) & (!g54) & (g2280) & (!g2281) & (g2289)) + ((g39) & (!g54) & (g2280) & (g2281) & (!g2289)) + ((g39) & (!g54) & (g2280) & (g2281) & (g2289)) + ((g39) & (g54) & (!g2280) & (!g2281) & (g2289)) + ((g39) & (g54) & (!g2280) & (g2281) & (!g2289)) + ((g39) & (g54) & (!g2280) & (g2281) & (g2289)) + ((g39) & (g54) & (g2280) & (!g2281) & (!g2289)) + ((g39) & (g54) & (g2280) & (!g2281) & (g2289)) + ((g39) & (g54) & (g2280) & (g2281) & (!g2289)) + ((g39) & (g54) & (g2280) & (g2281) & (g2289)));
	assign g2291 = (((!g18) & (!g27) & (g2278) & (g2279) & (g2290)) + ((!g18) & (g27) & (g2278) & (!g2279) & (g2290)) + ((!g18) & (g27) & (g2278) & (g2279) & (!g2290)) + ((!g18) & (g27) & (g2278) & (g2279) & (g2290)) + ((g18) & (!g27) & (!g2278) & (g2279) & (g2290)) + ((g18) & (!g27) & (g2278) & (!g2279) & (!g2290)) + ((g18) & (!g27) & (g2278) & (!g2279) & (g2290)) + ((g18) & (!g27) & (g2278) & (g2279) & (!g2290)) + ((g18) & (!g27) & (g2278) & (g2279) & (g2290)) + ((g18) & (g27) & (!g2278) & (!g2279) & (g2290)) + ((g18) & (g27) & (!g2278) & (g2279) & (!g2290)) + ((g18) & (g27) & (!g2278) & (g2279) & (g2290)) + ((g18) & (g27) & (g2278) & (!g2279) & (!g2290)) + ((g18) & (g27) & (g2278) & (!g2279) & (g2290)) + ((g18) & (g27) & (g2278) & (g2279) & (!g2290)) + ((g18) & (g27) & (g2278) & (g2279) & (g2290)));
	assign g2292 = (((!g2) & (!g8) & (g2276) & (g2277) & (g2291)) + ((!g2) & (g8) & (g2276) & (!g2277) & (g2291)) + ((!g2) & (g8) & (g2276) & (g2277) & (!g2291)) + ((!g2) & (g8) & (g2276) & (g2277) & (g2291)) + ((g2) & (!g8) & (!g2276) & (g2277) & (g2291)) + ((g2) & (!g8) & (g2276) & (!g2277) & (!g2291)) + ((g2) & (!g8) & (g2276) & (!g2277) & (g2291)) + ((g2) & (!g8) & (g2276) & (g2277) & (!g2291)) + ((g2) & (!g8) & (g2276) & (g2277) & (g2291)) + ((g2) & (g8) & (!g2276) & (!g2277) & (g2291)) + ((g2) & (g8) & (!g2276) & (g2277) & (!g2291)) + ((g2) & (g8) & (!g2276) & (g2277) & (g2291)) + ((g2) & (g8) & (g2276) & (!g2277) & (!g2291)) + ((g2) & (g8) & (g2276) & (!g2277) & (g2291)) + ((g2) & (g8) & (g2276) & (g2277) & (!g2291)) + ((g2) & (g8) & (g2276) & (g2277) & (g2291)));
	assign g2293 = (((!g2) & (!g2188) & (g2211) & (!g2218)) + ((!g2) & (g2188) & (!g2211) & (!g2218)) + ((!g2) & (g2188) & (!g2211) & (g2218)) + ((!g2) & (g2188) & (g2211) & (g2218)) + ((g2) & (!g2188) & (!g2211) & (!g2218)) + ((g2) & (g2188) & (!g2211) & (g2218)) + ((g2) & (g2188) & (g2211) & (!g2218)) + ((g2) & (g2188) & (g2211) & (g2218)));
	assign g2294 = (((!g1) & (!g2187) & (!g2214) & (!g2216) & (g2217)) + ((!g1) & (!g2187) & (!g2214) & (g2216) & (!g2217)) + ((!g1) & (!g2187) & (!g2214) & (g2216) & (g2217)) + ((!g1) & (g2187) & (g2214) & (!g2216) & (!g2217)) + ((!g1) & (g2187) & (g2214) & (!g2216) & (g2217)) + ((!g1) & (g2187) & (g2214) & (g2216) & (!g2217)) + ((!g1) & (g2187) & (g2214) & (g2216) & (g2217)) + ((g1) & (!g2187) & (!g2214) & (!g2216) & (g2217)) + ((g1) & (!g2187) & (!g2214) & (g2216) & (g2217)) + ((g1) & (g2187) & (g2214) & (!g2216) & (!g2217)) + ((g1) & (g2187) & (g2214) & (!g2216) & (g2217)) + ((g1) & (g2187) & (g2214) & (g2216) & (!g2217)) + ((g1) & (g2187) & (g2214) & (g2216) & (g2217)));
	assign g2295 = (((!g4) & (!g1) & (!g2275) & (!g2292) & (!g2293) & (!g2294)) + ((!g4) & (g1) & (!g2275) & (!g2292) & (!g2293) & (!g2294)) + ((!g4) & (g1) & (!g2275) & (!g2292) & (!g2293) & (g2294)) + ((!g4) & (g1) & (!g2275) & (!g2292) & (g2293) & (!g2294)) + ((!g4) & (g1) & (!g2275) & (!g2292) & (g2293) & (g2294)) + ((!g4) & (g1) & (!g2275) & (g2292) & (!g2293) & (!g2294)) + ((!g4) & (g1) & (!g2275) & (g2292) & (!g2293) & (g2294)) + ((!g4) & (g1) & (!g2275) & (g2292) & (g2293) & (!g2294)) + ((!g4) & (g1) & (!g2275) & (g2292) & (g2293) & (g2294)) + ((!g4) & (g1) & (g2275) & (!g2292) & (!g2293) & (!g2294)) + ((!g4) & (g1) & (g2275) & (!g2292) & (!g2293) & (g2294)) + ((g4) & (!g1) & (!g2275) & (!g2292) & (!g2293) & (!g2294)) + ((g4) & (!g1) & (!g2275) & (!g2292) & (g2293) & (!g2294)) + ((g4) & (!g1) & (!g2275) & (g2292) & (!g2293) & (!g2294)) + ((g4) & (g1) & (!g2275) & (!g2292) & (!g2293) & (!g2294)) + ((g4) & (g1) & (!g2275) & (!g2292) & (!g2293) & (g2294)) + ((g4) & (g1) & (!g2275) & (!g2292) & (g2293) & (!g2294)) + ((g4) & (g1) & (!g2275) & (!g2292) & (g2293) & (g2294)) + ((g4) & (g1) & (!g2275) & (g2292) & (!g2293) & (!g2294)) + ((g4) & (g1) & (!g2275) & (g2292) & (!g2293) & (g2294)) + ((g4) & (g1) & (!g2275) & (g2292) & (g2293) & (!g2294)) + ((g4) & (g1) & (!g2275) & (g2292) & (g2293) & (g2294)) + ((g4) & (g1) & (g2275) & (!g2292) & (!g2293) & (!g2294)) + ((g4) & (g1) & (g2275) & (!g2292) & (!g2293) & (g2294)) + ((g4) & (g1) & (g2275) & (!g2292) & (g2293) & (!g2294)) + ((g4) & (g1) & (g2275) & (!g2292) & (g2293) & (g2294)) + ((g4) & (g1) & (g2275) & (g2292) & (!g2293) & (!g2294)) + ((g4) & (g1) & (g2275) & (g2292) & (!g2293) & (g2294)));
	assign g2296 = (((!g174) & (!g2219) & (g2273) & (!g2274) & (!g2295)) + ((!g174) & (!g2219) & (g2273) & (g2274) & (!g2295)) + ((!g174) & (!g2219) & (g2273) & (g2274) & (g2295)) + ((!g174) & (g2219) & (!g2273) & (!g2274) & (!g2295)) + ((!g174) & (g2219) & (!g2273) & (!g2274) & (g2295)) + ((!g174) & (g2219) & (!g2273) & (g2274) & (!g2295)) + ((!g174) & (g2219) & (!g2273) & (g2274) & (g2295)) + ((!g174) & (g2219) & (g2273) & (!g2274) & (g2295)) + ((g174) & (!g2219) & (!g2273) & (!g2274) & (!g2295)) + ((g174) & (!g2219) & (!g2273) & (g2274) & (!g2295)) + ((g174) & (!g2219) & (!g2273) & (g2274) & (g2295)) + ((g174) & (g2219) & (!g2273) & (!g2274) & (g2295)) + ((g174) & (g2219) & (g2273) & (!g2274) & (!g2295)) + ((g174) & (g2219) & (g2273) & (!g2274) & (g2295)) + ((g174) & (g2219) & (g2273) & (g2274) & (!g2295)) + ((g174) & (g2219) & (g2273) & (g2274) & (g2295)));
	assign g2297 = (((!g198) & (!g229) & (g2221) & (g2272)) + ((!g198) & (g229) & (!g2221) & (g2272)) + ((!g198) & (g229) & (g2221) & (!g2272)) + ((!g198) & (g229) & (g2221) & (g2272)) + ((g198) & (!g229) & (!g2221) & (!g2272)) + ((g198) & (!g229) & (!g2221) & (g2272)) + ((g198) & (!g229) & (g2221) & (!g2272)) + ((g198) & (g229) & (!g2221) & (!g2272)));
	assign g2298 = (((!g2220) & (!g2274) & (!g2295) & (g2297)) + ((!g2220) & (g2274) & (!g2295) & (g2297)) + ((!g2220) & (g2274) & (g2295) & (g2297)) + ((g2220) & (!g2274) & (!g2295) & (!g2297)) + ((g2220) & (!g2274) & (g2295) & (!g2297)) + ((g2220) & (!g2274) & (g2295) & (g2297)) + ((g2220) & (g2274) & (!g2295) & (!g2297)) + ((g2220) & (g2274) & (g2295) & (!g2297)));
	assign g2299 = (((!g229) & (!g2221) & (g2272) & (!g2274) & (!g2295)) + ((!g229) & (!g2221) & (g2272) & (g2274) & (!g2295)) + ((!g229) & (!g2221) & (g2272) & (g2274) & (g2295)) + ((!g229) & (g2221) & (!g2272) & (!g2274) & (!g2295)) + ((!g229) & (g2221) & (!g2272) & (!g2274) & (g2295)) + ((!g229) & (g2221) & (!g2272) & (g2274) & (!g2295)) + ((!g229) & (g2221) & (!g2272) & (g2274) & (g2295)) + ((!g229) & (g2221) & (g2272) & (!g2274) & (g2295)) + ((g229) & (!g2221) & (!g2272) & (!g2274) & (!g2295)) + ((g229) & (!g2221) & (!g2272) & (g2274) & (!g2295)) + ((g229) & (!g2221) & (!g2272) & (g2274) & (g2295)) + ((g229) & (g2221) & (!g2272) & (!g2274) & (g2295)) + ((g229) & (g2221) & (g2272) & (!g2274) & (!g2295)) + ((g229) & (g2221) & (g2272) & (!g2274) & (g2295)) + ((g229) & (g2221) & (g2272) & (g2274) & (!g2295)) + ((g229) & (g2221) & (g2272) & (g2274) & (g2295)));
	assign g2300 = (((!g255) & (!g290) & (g2223) & (g2271)) + ((!g255) & (g290) & (!g2223) & (g2271)) + ((!g255) & (g290) & (g2223) & (!g2271)) + ((!g255) & (g290) & (g2223) & (g2271)) + ((g255) & (!g290) & (!g2223) & (!g2271)) + ((g255) & (!g290) & (!g2223) & (g2271)) + ((g255) & (!g290) & (g2223) & (!g2271)) + ((g255) & (g290) & (!g2223) & (!g2271)));
	assign g2301 = (((!g2222) & (!g2274) & (!g2295) & (g2300)) + ((!g2222) & (g2274) & (!g2295) & (g2300)) + ((!g2222) & (g2274) & (g2295) & (g2300)) + ((g2222) & (!g2274) & (!g2295) & (!g2300)) + ((g2222) & (!g2274) & (g2295) & (!g2300)) + ((g2222) & (!g2274) & (g2295) & (g2300)) + ((g2222) & (g2274) & (!g2295) & (!g2300)) + ((g2222) & (g2274) & (g2295) & (!g2300)));
	assign g2302 = (((!g290) & (!g2223) & (g2271) & (!g2274) & (!g2295)) + ((!g290) & (!g2223) & (g2271) & (g2274) & (!g2295)) + ((!g290) & (!g2223) & (g2271) & (g2274) & (g2295)) + ((!g290) & (g2223) & (!g2271) & (!g2274) & (!g2295)) + ((!g290) & (g2223) & (!g2271) & (!g2274) & (g2295)) + ((!g290) & (g2223) & (!g2271) & (g2274) & (!g2295)) + ((!g290) & (g2223) & (!g2271) & (g2274) & (g2295)) + ((!g290) & (g2223) & (g2271) & (!g2274) & (g2295)) + ((g290) & (!g2223) & (!g2271) & (!g2274) & (!g2295)) + ((g290) & (!g2223) & (!g2271) & (g2274) & (!g2295)) + ((g290) & (!g2223) & (!g2271) & (g2274) & (g2295)) + ((g290) & (g2223) & (!g2271) & (!g2274) & (g2295)) + ((g290) & (g2223) & (g2271) & (!g2274) & (!g2295)) + ((g290) & (g2223) & (g2271) & (!g2274) & (g2295)) + ((g290) & (g2223) & (g2271) & (g2274) & (!g2295)) + ((g290) & (g2223) & (g2271) & (g2274) & (g2295)));
	assign g2303 = (((!g319) & (!g358) & (g2225) & (g2270)) + ((!g319) & (g358) & (!g2225) & (g2270)) + ((!g319) & (g358) & (g2225) & (!g2270)) + ((!g319) & (g358) & (g2225) & (g2270)) + ((g319) & (!g358) & (!g2225) & (!g2270)) + ((g319) & (!g358) & (!g2225) & (g2270)) + ((g319) & (!g358) & (g2225) & (!g2270)) + ((g319) & (g358) & (!g2225) & (!g2270)));
	assign g2304 = (((!g2224) & (!g2274) & (!g2295) & (g2303)) + ((!g2224) & (g2274) & (!g2295) & (g2303)) + ((!g2224) & (g2274) & (g2295) & (g2303)) + ((g2224) & (!g2274) & (!g2295) & (!g2303)) + ((g2224) & (!g2274) & (g2295) & (!g2303)) + ((g2224) & (!g2274) & (g2295) & (g2303)) + ((g2224) & (g2274) & (!g2295) & (!g2303)) + ((g2224) & (g2274) & (g2295) & (!g2303)));
	assign g2305 = (((!g358) & (!g2225) & (g2270) & (!g2274) & (!g2295)) + ((!g358) & (!g2225) & (g2270) & (g2274) & (!g2295)) + ((!g358) & (!g2225) & (g2270) & (g2274) & (g2295)) + ((!g358) & (g2225) & (!g2270) & (!g2274) & (!g2295)) + ((!g358) & (g2225) & (!g2270) & (!g2274) & (g2295)) + ((!g358) & (g2225) & (!g2270) & (g2274) & (!g2295)) + ((!g358) & (g2225) & (!g2270) & (g2274) & (g2295)) + ((!g358) & (g2225) & (g2270) & (!g2274) & (g2295)) + ((g358) & (!g2225) & (!g2270) & (!g2274) & (!g2295)) + ((g358) & (!g2225) & (!g2270) & (g2274) & (!g2295)) + ((g358) & (!g2225) & (!g2270) & (g2274) & (g2295)) + ((g358) & (g2225) & (!g2270) & (!g2274) & (g2295)) + ((g358) & (g2225) & (g2270) & (!g2274) & (!g2295)) + ((g358) & (g2225) & (g2270) & (!g2274) & (g2295)) + ((g358) & (g2225) & (g2270) & (g2274) & (!g2295)) + ((g358) & (g2225) & (g2270) & (g2274) & (g2295)));
	assign g2306 = (((!g390) & (!g433) & (g2227) & (g2269)) + ((!g390) & (g433) & (!g2227) & (g2269)) + ((!g390) & (g433) & (g2227) & (!g2269)) + ((!g390) & (g433) & (g2227) & (g2269)) + ((g390) & (!g433) & (!g2227) & (!g2269)) + ((g390) & (!g433) & (!g2227) & (g2269)) + ((g390) & (!g433) & (g2227) & (!g2269)) + ((g390) & (g433) & (!g2227) & (!g2269)));
	assign g2307 = (((!g2226) & (!g2274) & (!g2295) & (g2306)) + ((!g2226) & (g2274) & (!g2295) & (g2306)) + ((!g2226) & (g2274) & (g2295) & (g2306)) + ((g2226) & (!g2274) & (!g2295) & (!g2306)) + ((g2226) & (!g2274) & (g2295) & (!g2306)) + ((g2226) & (!g2274) & (g2295) & (g2306)) + ((g2226) & (g2274) & (!g2295) & (!g2306)) + ((g2226) & (g2274) & (g2295) & (!g2306)));
	assign g2308 = (((!g433) & (!g2227) & (g2269) & (!g2274) & (!g2295)) + ((!g433) & (!g2227) & (g2269) & (g2274) & (!g2295)) + ((!g433) & (!g2227) & (g2269) & (g2274) & (g2295)) + ((!g433) & (g2227) & (!g2269) & (!g2274) & (!g2295)) + ((!g433) & (g2227) & (!g2269) & (!g2274) & (g2295)) + ((!g433) & (g2227) & (!g2269) & (g2274) & (!g2295)) + ((!g433) & (g2227) & (!g2269) & (g2274) & (g2295)) + ((!g433) & (g2227) & (g2269) & (!g2274) & (g2295)) + ((g433) & (!g2227) & (!g2269) & (!g2274) & (!g2295)) + ((g433) & (!g2227) & (!g2269) & (g2274) & (!g2295)) + ((g433) & (!g2227) & (!g2269) & (g2274) & (g2295)) + ((g433) & (g2227) & (!g2269) & (!g2274) & (g2295)) + ((g433) & (g2227) & (g2269) & (!g2274) & (!g2295)) + ((g433) & (g2227) & (g2269) & (!g2274) & (g2295)) + ((g433) & (g2227) & (g2269) & (g2274) & (!g2295)) + ((g433) & (g2227) & (g2269) & (g2274) & (g2295)));
	assign g2309 = (((!g468) & (!g515) & (g2229) & (g2268)) + ((!g468) & (g515) & (!g2229) & (g2268)) + ((!g468) & (g515) & (g2229) & (!g2268)) + ((!g468) & (g515) & (g2229) & (g2268)) + ((g468) & (!g515) & (!g2229) & (!g2268)) + ((g468) & (!g515) & (!g2229) & (g2268)) + ((g468) & (!g515) & (g2229) & (!g2268)) + ((g468) & (g515) & (!g2229) & (!g2268)));
	assign g2310 = (((!g2228) & (!g2274) & (!g2295) & (g2309)) + ((!g2228) & (g2274) & (!g2295) & (g2309)) + ((!g2228) & (g2274) & (g2295) & (g2309)) + ((g2228) & (!g2274) & (!g2295) & (!g2309)) + ((g2228) & (!g2274) & (g2295) & (!g2309)) + ((g2228) & (!g2274) & (g2295) & (g2309)) + ((g2228) & (g2274) & (!g2295) & (!g2309)) + ((g2228) & (g2274) & (g2295) & (!g2309)));
	assign g2311 = (((!g515) & (!g2229) & (g2268) & (!g2274) & (!g2295)) + ((!g515) & (!g2229) & (g2268) & (g2274) & (!g2295)) + ((!g515) & (!g2229) & (g2268) & (g2274) & (g2295)) + ((!g515) & (g2229) & (!g2268) & (!g2274) & (!g2295)) + ((!g515) & (g2229) & (!g2268) & (!g2274) & (g2295)) + ((!g515) & (g2229) & (!g2268) & (g2274) & (!g2295)) + ((!g515) & (g2229) & (!g2268) & (g2274) & (g2295)) + ((!g515) & (g2229) & (g2268) & (!g2274) & (g2295)) + ((g515) & (!g2229) & (!g2268) & (!g2274) & (!g2295)) + ((g515) & (!g2229) & (!g2268) & (g2274) & (!g2295)) + ((g515) & (!g2229) & (!g2268) & (g2274) & (g2295)) + ((g515) & (g2229) & (!g2268) & (!g2274) & (g2295)) + ((g515) & (g2229) & (g2268) & (!g2274) & (!g2295)) + ((g515) & (g2229) & (g2268) & (!g2274) & (g2295)) + ((g515) & (g2229) & (g2268) & (g2274) & (!g2295)) + ((g515) & (g2229) & (g2268) & (g2274) & (g2295)));
	assign g2312 = (((!g553) & (!g604) & (g2231) & (g2267)) + ((!g553) & (g604) & (!g2231) & (g2267)) + ((!g553) & (g604) & (g2231) & (!g2267)) + ((!g553) & (g604) & (g2231) & (g2267)) + ((g553) & (!g604) & (!g2231) & (!g2267)) + ((g553) & (!g604) & (!g2231) & (g2267)) + ((g553) & (!g604) & (g2231) & (!g2267)) + ((g553) & (g604) & (!g2231) & (!g2267)));
	assign g2313 = (((!g2230) & (!g2274) & (!g2295) & (g2312)) + ((!g2230) & (g2274) & (!g2295) & (g2312)) + ((!g2230) & (g2274) & (g2295) & (g2312)) + ((g2230) & (!g2274) & (!g2295) & (!g2312)) + ((g2230) & (!g2274) & (g2295) & (!g2312)) + ((g2230) & (!g2274) & (g2295) & (g2312)) + ((g2230) & (g2274) & (!g2295) & (!g2312)) + ((g2230) & (g2274) & (g2295) & (!g2312)));
	assign g2314 = (((!g604) & (!g2231) & (g2267) & (!g2274) & (!g2295)) + ((!g604) & (!g2231) & (g2267) & (g2274) & (!g2295)) + ((!g604) & (!g2231) & (g2267) & (g2274) & (g2295)) + ((!g604) & (g2231) & (!g2267) & (!g2274) & (!g2295)) + ((!g604) & (g2231) & (!g2267) & (!g2274) & (g2295)) + ((!g604) & (g2231) & (!g2267) & (g2274) & (!g2295)) + ((!g604) & (g2231) & (!g2267) & (g2274) & (g2295)) + ((!g604) & (g2231) & (g2267) & (!g2274) & (g2295)) + ((g604) & (!g2231) & (!g2267) & (!g2274) & (!g2295)) + ((g604) & (!g2231) & (!g2267) & (g2274) & (!g2295)) + ((g604) & (!g2231) & (!g2267) & (g2274) & (g2295)) + ((g604) & (g2231) & (!g2267) & (!g2274) & (g2295)) + ((g604) & (g2231) & (g2267) & (!g2274) & (!g2295)) + ((g604) & (g2231) & (g2267) & (!g2274) & (g2295)) + ((g604) & (g2231) & (g2267) & (g2274) & (!g2295)) + ((g604) & (g2231) & (g2267) & (g2274) & (g2295)));
	assign g2315 = (((!g645) & (!g700) & (g2233) & (g2266)) + ((!g645) & (g700) & (!g2233) & (g2266)) + ((!g645) & (g700) & (g2233) & (!g2266)) + ((!g645) & (g700) & (g2233) & (g2266)) + ((g645) & (!g700) & (!g2233) & (!g2266)) + ((g645) & (!g700) & (!g2233) & (g2266)) + ((g645) & (!g700) & (g2233) & (!g2266)) + ((g645) & (g700) & (!g2233) & (!g2266)));
	assign g2316 = (((!g2232) & (!g2274) & (!g2295) & (g2315)) + ((!g2232) & (g2274) & (!g2295) & (g2315)) + ((!g2232) & (g2274) & (g2295) & (g2315)) + ((g2232) & (!g2274) & (!g2295) & (!g2315)) + ((g2232) & (!g2274) & (g2295) & (!g2315)) + ((g2232) & (!g2274) & (g2295) & (g2315)) + ((g2232) & (g2274) & (!g2295) & (!g2315)) + ((g2232) & (g2274) & (g2295) & (!g2315)));
	assign g2317 = (((!g700) & (!g2233) & (g2266) & (!g2274) & (!g2295)) + ((!g700) & (!g2233) & (g2266) & (g2274) & (!g2295)) + ((!g700) & (!g2233) & (g2266) & (g2274) & (g2295)) + ((!g700) & (g2233) & (!g2266) & (!g2274) & (!g2295)) + ((!g700) & (g2233) & (!g2266) & (!g2274) & (g2295)) + ((!g700) & (g2233) & (!g2266) & (g2274) & (!g2295)) + ((!g700) & (g2233) & (!g2266) & (g2274) & (g2295)) + ((!g700) & (g2233) & (g2266) & (!g2274) & (g2295)) + ((g700) & (!g2233) & (!g2266) & (!g2274) & (!g2295)) + ((g700) & (!g2233) & (!g2266) & (g2274) & (!g2295)) + ((g700) & (!g2233) & (!g2266) & (g2274) & (g2295)) + ((g700) & (g2233) & (!g2266) & (!g2274) & (g2295)) + ((g700) & (g2233) & (g2266) & (!g2274) & (!g2295)) + ((g700) & (g2233) & (g2266) & (!g2274) & (g2295)) + ((g700) & (g2233) & (g2266) & (g2274) & (!g2295)) + ((g700) & (g2233) & (g2266) & (g2274) & (g2295)));
	assign g2318 = (((!g744) & (!g803) & (g2235) & (g2265)) + ((!g744) & (g803) & (!g2235) & (g2265)) + ((!g744) & (g803) & (g2235) & (!g2265)) + ((!g744) & (g803) & (g2235) & (g2265)) + ((g744) & (!g803) & (!g2235) & (!g2265)) + ((g744) & (!g803) & (!g2235) & (g2265)) + ((g744) & (!g803) & (g2235) & (!g2265)) + ((g744) & (g803) & (!g2235) & (!g2265)));
	assign g2319 = (((!g2234) & (!g2274) & (!g2295) & (g2318)) + ((!g2234) & (g2274) & (!g2295) & (g2318)) + ((!g2234) & (g2274) & (g2295) & (g2318)) + ((g2234) & (!g2274) & (!g2295) & (!g2318)) + ((g2234) & (!g2274) & (g2295) & (!g2318)) + ((g2234) & (!g2274) & (g2295) & (g2318)) + ((g2234) & (g2274) & (!g2295) & (!g2318)) + ((g2234) & (g2274) & (g2295) & (!g2318)));
	assign g2320 = (((!g803) & (!g2235) & (g2265) & (!g2274) & (!g2295)) + ((!g803) & (!g2235) & (g2265) & (g2274) & (!g2295)) + ((!g803) & (!g2235) & (g2265) & (g2274) & (g2295)) + ((!g803) & (g2235) & (!g2265) & (!g2274) & (!g2295)) + ((!g803) & (g2235) & (!g2265) & (!g2274) & (g2295)) + ((!g803) & (g2235) & (!g2265) & (g2274) & (!g2295)) + ((!g803) & (g2235) & (!g2265) & (g2274) & (g2295)) + ((!g803) & (g2235) & (g2265) & (!g2274) & (g2295)) + ((g803) & (!g2235) & (!g2265) & (!g2274) & (!g2295)) + ((g803) & (!g2235) & (!g2265) & (g2274) & (!g2295)) + ((g803) & (!g2235) & (!g2265) & (g2274) & (g2295)) + ((g803) & (g2235) & (!g2265) & (!g2274) & (g2295)) + ((g803) & (g2235) & (g2265) & (!g2274) & (!g2295)) + ((g803) & (g2235) & (g2265) & (!g2274) & (g2295)) + ((g803) & (g2235) & (g2265) & (g2274) & (!g2295)) + ((g803) & (g2235) & (g2265) & (g2274) & (g2295)));
	assign g2321 = (((!g851) & (!g914) & (g2237) & (g2264)) + ((!g851) & (g914) & (!g2237) & (g2264)) + ((!g851) & (g914) & (g2237) & (!g2264)) + ((!g851) & (g914) & (g2237) & (g2264)) + ((g851) & (!g914) & (!g2237) & (!g2264)) + ((g851) & (!g914) & (!g2237) & (g2264)) + ((g851) & (!g914) & (g2237) & (!g2264)) + ((g851) & (g914) & (!g2237) & (!g2264)));
	assign g2322 = (((!g2236) & (!g2274) & (!g2295) & (g2321)) + ((!g2236) & (g2274) & (!g2295) & (g2321)) + ((!g2236) & (g2274) & (g2295) & (g2321)) + ((g2236) & (!g2274) & (!g2295) & (!g2321)) + ((g2236) & (!g2274) & (g2295) & (!g2321)) + ((g2236) & (!g2274) & (g2295) & (g2321)) + ((g2236) & (g2274) & (!g2295) & (!g2321)) + ((g2236) & (g2274) & (g2295) & (!g2321)));
	assign g2323 = (((!g914) & (!g2237) & (g2264) & (!g2274) & (!g2295)) + ((!g914) & (!g2237) & (g2264) & (g2274) & (!g2295)) + ((!g914) & (!g2237) & (g2264) & (g2274) & (g2295)) + ((!g914) & (g2237) & (!g2264) & (!g2274) & (!g2295)) + ((!g914) & (g2237) & (!g2264) & (!g2274) & (g2295)) + ((!g914) & (g2237) & (!g2264) & (g2274) & (!g2295)) + ((!g914) & (g2237) & (!g2264) & (g2274) & (g2295)) + ((!g914) & (g2237) & (g2264) & (!g2274) & (g2295)) + ((g914) & (!g2237) & (!g2264) & (!g2274) & (!g2295)) + ((g914) & (!g2237) & (!g2264) & (g2274) & (!g2295)) + ((g914) & (!g2237) & (!g2264) & (g2274) & (g2295)) + ((g914) & (g2237) & (!g2264) & (!g2274) & (g2295)) + ((g914) & (g2237) & (g2264) & (!g2274) & (!g2295)) + ((g914) & (g2237) & (g2264) & (!g2274) & (g2295)) + ((g914) & (g2237) & (g2264) & (g2274) & (!g2295)) + ((g914) & (g2237) & (g2264) & (g2274) & (g2295)));
	assign g2324 = (((!g1032) & (!g1030) & (g2239) & (g2263)) + ((!g1032) & (g1030) & (!g2239) & (g2263)) + ((!g1032) & (g1030) & (g2239) & (!g2263)) + ((!g1032) & (g1030) & (g2239) & (g2263)) + ((g1032) & (!g1030) & (!g2239) & (!g2263)) + ((g1032) & (!g1030) & (!g2239) & (g2263)) + ((g1032) & (!g1030) & (g2239) & (!g2263)) + ((g1032) & (g1030) & (!g2239) & (!g2263)));
	assign g2325 = (((!g2238) & (!g2274) & (!g2295) & (g2324)) + ((!g2238) & (g2274) & (!g2295) & (g2324)) + ((!g2238) & (g2274) & (g2295) & (g2324)) + ((g2238) & (!g2274) & (!g2295) & (!g2324)) + ((g2238) & (!g2274) & (g2295) & (!g2324)) + ((g2238) & (!g2274) & (g2295) & (g2324)) + ((g2238) & (g2274) & (!g2295) & (!g2324)) + ((g2238) & (g2274) & (g2295) & (!g2324)));
	assign g2326 = (((!g1030) & (!g2239) & (g2263) & (!g2274) & (!g2295)) + ((!g1030) & (!g2239) & (g2263) & (g2274) & (!g2295)) + ((!g1030) & (!g2239) & (g2263) & (g2274) & (g2295)) + ((!g1030) & (g2239) & (!g2263) & (!g2274) & (!g2295)) + ((!g1030) & (g2239) & (!g2263) & (!g2274) & (g2295)) + ((!g1030) & (g2239) & (!g2263) & (g2274) & (!g2295)) + ((!g1030) & (g2239) & (!g2263) & (g2274) & (g2295)) + ((!g1030) & (g2239) & (g2263) & (!g2274) & (g2295)) + ((g1030) & (!g2239) & (!g2263) & (!g2274) & (!g2295)) + ((g1030) & (!g2239) & (!g2263) & (g2274) & (!g2295)) + ((g1030) & (!g2239) & (!g2263) & (g2274) & (g2295)) + ((g1030) & (g2239) & (!g2263) & (!g2274) & (g2295)) + ((g1030) & (g2239) & (g2263) & (!g2274) & (!g2295)) + ((g1030) & (g2239) & (g2263) & (!g2274) & (g2295)) + ((g1030) & (g2239) & (g2263) & (g2274) & (!g2295)) + ((g1030) & (g2239) & (g2263) & (g2274) & (g2295)));
	assign g2327 = (((!g1160) & (!g1154) & (g2241) & (g2262)) + ((!g1160) & (g1154) & (!g2241) & (g2262)) + ((!g1160) & (g1154) & (g2241) & (!g2262)) + ((!g1160) & (g1154) & (g2241) & (g2262)) + ((g1160) & (!g1154) & (!g2241) & (!g2262)) + ((g1160) & (!g1154) & (!g2241) & (g2262)) + ((g1160) & (!g1154) & (g2241) & (!g2262)) + ((g1160) & (g1154) & (!g2241) & (!g2262)));
	assign g2328 = (((!g2240) & (!g2274) & (!g2295) & (g2327)) + ((!g2240) & (g2274) & (!g2295) & (g2327)) + ((!g2240) & (g2274) & (g2295) & (g2327)) + ((g2240) & (!g2274) & (!g2295) & (!g2327)) + ((g2240) & (!g2274) & (g2295) & (!g2327)) + ((g2240) & (!g2274) & (g2295) & (g2327)) + ((g2240) & (g2274) & (!g2295) & (!g2327)) + ((g2240) & (g2274) & (g2295) & (!g2327)));
	assign g2329 = (((!g1154) & (!g2241) & (g2262) & (!g2274) & (!g2295)) + ((!g1154) & (!g2241) & (g2262) & (g2274) & (!g2295)) + ((!g1154) & (!g2241) & (g2262) & (g2274) & (g2295)) + ((!g1154) & (g2241) & (!g2262) & (!g2274) & (!g2295)) + ((!g1154) & (g2241) & (!g2262) & (!g2274) & (g2295)) + ((!g1154) & (g2241) & (!g2262) & (g2274) & (!g2295)) + ((!g1154) & (g2241) & (!g2262) & (g2274) & (g2295)) + ((!g1154) & (g2241) & (g2262) & (!g2274) & (g2295)) + ((g1154) & (!g2241) & (!g2262) & (!g2274) & (!g2295)) + ((g1154) & (!g2241) & (!g2262) & (g2274) & (!g2295)) + ((g1154) & (!g2241) & (!g2262) & (g2274) & (g2295)) + ((g1154) & (g2241) & (!g2262) & (!g2274) & (g2295)) + ((g1154) & (g2241) & (g2262) & (!g2274) & (!g2295)) + ((g1154) & (g2241) & (g2262) & (!g2274) & (g2295)) + ((g1154) & (g2241) & (g2262) & (g2274) & (!g2295)) + ((g1154) & (g2241) & (g2262) & (g2274) & (g2295)));
	assign g2330 = (((!g1295) & (!g1285) & (g2243) & (g2261)) + ((!g1295) & (g1285) & (!g2243) & (g2261)) + ((!g1295) & (g1285) & (g2243) & (!g2261)) + ((!g1295) & (g1285) & (g2243) & (g2261)) + ((g1295) & (!g1285) & (!g2243) & (!g2261)) + ((g1295) & (!g1285) & (!g2243) & (g2261)) + ((g1295) & (!g1285) & (g2243) & (!g2261)) + ((g1295) & (g1285) & (!g2243) & (!g2261)));
	assign g2331 = (((!g2242) & (!g2274) & (!g2295) & (g2330)) + ((!g2242) & (g2274) & (!g2295) & (g2330)) + ((!g2242) & (g2274) & (g2295) & (g2330)) + ((g2242) & (!g2274) & (!g2295) & (!g2330)) + ((g2242) & (!g2274) & (g2295) & (!g2330)) + ((g2242) & (!g2274) & (g2295) & (g2330)) + ((g2242) & (g2274) & (!g2295) & (!g2330)) + ((g2242) & (g2274) & (g2295) & (!g2330)));
	assign g2332 = (((!g1285) & (!g2243) & (g2261) & (!g2274) & (!g2295)) + ((!g1285) & (!g2243) & (g2261) & (g2274) & (!g2295)) + ((!g1285) & (!g2243) & (g2261) & (g2274) & (g2295)) + ((!g1285) & (g2243) & (!g2261) & (!g2274) & (!g2295)) + ((!g1285) & (g2243) & (!g2261) & (!g2274) & (g2295)) + ((!g1285) & (g2243) & (!g2261) & (g2274) & (!g2295)) + ((!g1285) & (g2243) & (!g2261) & (g2274) & (g2295)) + ((!g1285) & (g2243) & (g2261) & (!g2274) & (g2295)) + ((g1285) & (!g2243) & (!g2261) & (!g2274) & (!g2295)) + ((g1285) & (!g2243) & (!g2261) & (g2274) & (!g2295)) + ((g1285) & (!g2243) & (!g2261) & (g2274) & (g2295)) + ((g1285) & (g2243) & (!g2261) & (!g2274) & (g2295)) + ((g1285) & (g2243) & (g2261) & (!g2274) & (!g2295)) + ((g1285) & (g2243) & (g2261) & (!g2274) & (g2295)) + ((g1285) & (g2243) & (g2261) & (g2274) & (!g2295)) + ((g1285) & (g2243) & (g2261) & (g2274) & (g2295)));
	assign g2333 = (((!g1437) & (!g1423) & (g2245) & (g2260)) + ((!g1437) & (g1423) & (!g2245) & (g2260)) + ((!g1437) & (g1423) & (g2245) & (!g2260)) + ((!g1437) & (g1423) & (g2245) & (g2260)) + ((g1437) & (!g1423) & (!g2245) & (!g2260)) + ((g1437) & (!g1423) & (!g2245) & (g2260)) + ((g1437) & (!g1423) & (g2245) & (!g2260)) + ((g1437) & (g1423) & (!g2245) & (!g2260)));
	assign g2334 = (((!g2244) & (!g2274) & (!g2295) & (g2333)) + ((!g2244) & (g2274) & (!g2295) & (g2333)) + ((!g2244) & (g2274) & (g2295) & (g2333)) + ((g2244) & (!g2274) & (!g2295) & (!g2333)) + ((g2244) & (!g2274) & (g2295) & (!g2333)) + ((g2244) & (!g2274) & (g2295) & (g2333)) + ((g2244) & (g2274) & (!g2295) & (!g2333)) + ((g2244) & (g2274) & (g2295) & (!g2333)));
	assign g2335 = (((!g1423) & (!g2245) & (g2260) & (!g2274) & (!g2295)) + ((!g1423) & (!g2245) & (g2260) & (g2274) & (!g2295)) + ((!g1423) & (!g2245) & (g2260) & (g2274) & (g2295)) + ((!g1423) & (g2245) & (!g2260) & (!g2274) & (!g2295)) + ((!g1423) & (g2245) & (!g2260) & (!g2274) & (g2295)) + ((!g1423) & (g2245) & (!g2260) & (g2274) & (!g2295)) + ((!g1423) & (g2245) & (!g2260) & (g2274) & (g2295)) + ((!g1423) & (g2245) & (g2260) & (!g2274) & (g2295)) + ((g1423) & (!g2245) & (!g2260) & (!g2274) & (!g2295)) + ((g1423) & (!g2245) & (!g2260) & (g2274) & (!g2295)) + ((g1423) & (!g2245) & (!g2260) & (g2274) & (g2295)) + ((g1423) & (g2245) & (!g2260) & (!g2274) & (g2295)) + ((g1423) & (g2245) & (g2260) & (!g2274) & (!g2295)) + ((g1423) & (g2245) & (g2260) & (!g2274) & (g2295)) + ((g1423) & (g2245) & (g2260) & (g2274) & (!g2295)) + ((g1423) & (g2245) & (g2260) & (g2274) & (g2295)));
	assign g2336 = (((!g1586) & (!g1568) & (g2247) & (g2259)) + ((!g1586) & (g1568) & (!g2247) & (g2259)) + ((!g1586) & (g1568) & (g2247) & (!g2259)) + ((!g1586) & (g1568) & (g2247) & (g2259)) + ((g1586) & (!g1568) & (!g2247) & (!g2259)) + ((g1586) & (!g1568) & (!g2247) & (g2259)) + ((g1586) & (!g1568) & (g2247) & (!g2259)) + ((g1586) & (g1568) & (!g2247) & (!g2259)));
	assign g2337 = (((!g2246) & (!g2274) & (!g2295) & (g2336)) + ((!g2246) & (g2274) & (!g2295) & (g2336)) + ((!g2246) & (g2274) & (g2295) & (g2336)) + ((g2246) & (!g2274) & (!g2295) & (!g2336)) + ((g2246) & (!g2274) & (g2295) & (!g2336)) + ((g2246) & (!g2274) & (g2295) & (g2336)) + ((g2246) & (g2274) & (!g2295) & (!g2336)) + ((g2246) & (g2274) & (g2295) & (!g2336)));
	assign g2338 = (((!g1568) & (!g2247) & (g2259) & (!g2274) & (!g2295)) + ((!g1568) & (!g2247) & (g2259) & (g2274) & (!g2295)) + ((!g1568) & (!g2247) & (g2259) & (g2274) & (g2295)) + ((!g1568) & (g2247) & (!g2259) & (!g2274) & (!g2295)) + ((!g1568) & (g2247) & (!g2259) & (!g2274) & (g2295)) + ((!g1568) & (g2247) & (!g2259) & (g2274) & (!g2295)) + ((!g1568) & (g2247) & (!g2259) & (g2274) & (g2295)) + ((!g1568) & (g2247) & (g2259) & (!g2274) & (g2295)) + ((g1568) & (!g2247) & (!g2259) & (!g2274) & (!g2295)) + ((g1568) & (!g2247) & (!g2259) & (g2274) & (!g2295)) + ((g1568) & (!g2247) & (!g2259) & (g2274) & (g2295)) + ((g1568) & (g2247) & (!g2259) & (!g2274) & (g2295)) + ((g1568) & (g2247) & (g2259) & (!g2274) & (!g2295)) + ((g1568) & (g2247) & (g2259) & (!g2274) & (g2295)) + ((g1568) & (g2247) & (g2259) & (g2274) & (!g2295)) + ((g1568) & (g2247) & (g2259) & (g2274) & (g2295)));
	assign g2339 = (((!g1742) & (!g1720) & (g2249) & (g2258)) + ((!g1742) & (g1720) & (!g2249) & (g2258)) + ((!g1742) & (g1720) & (g2249) & (!g2258)) + ((!g1742) & (g1720) & (g2249) & (g2258)) + ((g1742) & (!g1720) & (!g2249) & (!g2258)) + ((g1742) & (!g1720) & (!g2249) & (g2258)) + ((g1742) & (!g1720) & (g2249) & (!g2258)) + ((g1742) & (g1720) & (!g2249) & (!g2258)));
	assign g2340 = (((!g2248) & (!g2274) & (!g2295) & (g2339)) + ((!g2248) & (g2274) & (!g2295) & (g2339)) + ((!g2248) & (g2274) & (g2295) & (g2339)) + ((g2248) & (!g2274) & (!g2295) & (!g2339)) + ((g2248) & (!g2274) & (g2295) & (!g2339)) + ((g2248) & (!g2274) & (g2295) & (g2339)) + ((g2248) & (g2274) & (!g2295) & (!g2339)) + ((g2248) & (g2274) & (g2295) & (!g2339)));
	assign g2341 = (((!g1720) & (!g2249) & (g2258) & (!g2274) & (!g2295)) + ((!g1720) & (!g2249) & (g2258) & (g2274) & (!g2295)) + ((!g1720) & (!g2249) & (g2258) & (g2274) & (g2295)) + ((!g1720) & (g2249) & (!g2258) & (!g2274) & (!g2295)) + ((!g1720) & (g2249) & (!g2258) & (!g2274) & (g2295)) + ((!g1720) & (g2249) & (!g2258) & (g2274) & (!g2295)) + ((!g1720) & (g2249) & (!g2258) & (g2274) & (g2295)) + ((!g1720) & (g2249) & (g2258) & (!g2274) & (g2295)) + ((g1720) & (!g2249) & (!g2258) & (!g2274) & (!g2295)) + ((g1720) & (!g2249) & (!g2258) & (g2274) & (!g2295)) + ((g1720) & (!g2249) & (!g2258) & (g2274) & (g2295)) + ((g1720) & (g2249) & (!g2258) & (!g2274) & (g2295)) + ((g1720) & (g2249) & (g2258) & (!g2274) & (!g2295)) + ((g1720) & (g2249) & (g2258) & (!g2274) & (g2295)) + ((g1720) & (g2249) & (g2258) & (g2274) & (!g2295)) + ((g1720) & (g2249) & (g2258) & (g2274) & (g2295)));
	assign g2342 = (((!g1905) & (!g1879) & (g2251) & (g2257)) + ((!g1905) & (g1879) & (!g2251) & (g2257)) + ((!g1905) & (g1879) & (g2251) & (!g2257)) + ((!g1905) & (g1879) & (g2251) & (g2257)) + ((g1905) & (!g1879) & (!g2251) & (!g2257)) + ((g1905) & (!g1879) & (!g2251) & (g2257)) + ((g1905) & (!g1879) & (g2251) & (!g2257)) + ((g1905) & (g1879) & (!g2251) & (!g2257)));
	assign g2343 = (((!g2250) & (!g2274) & (!g2295) & (g2342)) + ((!g2250) & (g2274) & (!g2295) & (g2342)) + ((!g2250) & (g2274) & (g2295) & (g2342)) + ((g2250) & (!g2274) & (!g2295) & (!g2342)) + ((g2250) & (!g2274) & (g2295) & (!g2342)) + ((g2250) & (!g2274) & (g2295) & (g2342)) + ((g2250) & (g2274) & (!g2295) & (!g2342)) + ((g2250) & (g2274) & (g2295) & (!g2342)));
	assign g2344 = (((!g1879) & (!g2251) & (g2257) & (!g2274) & (!g2295)) + ((!g1879) & (!g2251) & (g2257) & (g2274) & (!g2295)) + ((!g1879) & (!g2251) & (g2257) & (g2274) & (g2295)) + ((!g1879) & (g2251) & (!g2257) & (!g2274) & (!g2295)) + ((!g1879) & (g2251) & (!g2257) & (!g2274) & (g2295)) + ((!g1879) & (g2251) & (!g2257) & (g2274) & (!g2295)) + ((!g1879) & (g2251) & (!g2257) & (g2274) & (g2295)) + ((!g1879) & (g2251) & (g2257) & (!g2274) & (g2295)) + ((g1879) & (!g2251) & (!g2257) & (!g2274) & (!g2295)) + ((g1879) & (!g2251) & (!g2257) & (g2274) & (!g2295)) + ((g1879) & (!g2251) & (!g2257) & (g2274) & (g2295)) + ((g1879) & (g2251) & (!g2257) & (!g2274) & (g2295)) + ((g1879) & (g2251) & (g2257) & (!g2274) & (!g2295)) + ((g1879) & (g2251) & (g2257) & (!g2274) & (g2295)) + ((g1879) & (g2251) & (g2257) & (g2274) & (!g2295)) + ((g1879) & (g2251) & (g2257) & (g2274) & (g2295)));
	assign g2345 = (((!g2075) & (!g2045) & (g2254) & (g2256)) + ((!g2075) & (g2045) & (!g2254) & (g2256)) + ((!g2075) & (g2045) & (g2254) & (!g2256)) + ((!g2075) & (g2045) & (g2254) & (g2256)) + ((g2075) & (!g2045) & (!g2254) & (!g2256)) + ((g2075) & (!g2045) & (!g2254) & (g2256)) + ((g2075) & (!g2045) & (g2254) & (!g2256)) + ((g2075) & (g2045) & (!g2254) & (!g2256)));
	assign g2346 = (((!g2253) & (!g2274) & (!g2295) & (g2345)) + ((!g2253) & (g2274) & (!g2295) & (g2345)) + ((!g2253) & (g2274) & (g2295) & (g2345)) + ((g2253) & (!g2274) & (!g2295) & (!g2345)) + ((g2253) & (!g2274) & (g2295) & (!g2345)) + ((g2253) & (!g2274) & (g2295) & (g2345)) + ((g2253) & (g2274) & (!g2295) & (!g2345)) + ((g2253) & (g2274) & (g2295) & (!g2345)));
	assign g2347 = (((!g2045) & (!g2254) & (g2256) & (!g2274) & (!g2295)) + ((!g2045) & (!g2254) & (g2256) & (g2274) & (!g2295)) + ((!g2045) & (!g2254) & (g2256) & (g2274) & (g2295)) + ((!g2045) & (g2254) & (!g2256) & (!g2274) & (!g2295)) + ((!g2045) & (g2254) & (!g2256) & (!g2274) & (g2295)) + ((!g2045) & (g2254) & (!g2256) & (g2274) & (!g2295)) + ((!g2045) & (g2254) & (!g2256) & (g2274) & (g2295)) + ((!g2045) & (g2254) & (g2256) & (!g2274) & (g2295)) + ((g2045) & (!g2254) & (!g2256) & (!g2274) & (!g2295)) + ((g2045) & (!g2254) & (!g2256) & (g2274) & (!g2295)) + ((g2045) & (!g2254) & (!g2256) & (g2274) & (g2295)) + ((g2045) & (g2254) & (!g2256) & (!g2274) & (g2295)) + ((g2045) & (g2254) & (g2256) & (!g2274) & (!g2295)) + ((g2045) & (g2254) & (g2256) & (!g2274) & (g2295)) + ((g2045) & (g2254) & (g2256) & (g2274) & (!g2295)) + ((g2045) & (g2254) & (g2256) & (g2274) & (g2295)));
	assign g2348 = (((!g2252) & (!ax28x) & (!g2218) & (g2255)) + ((!g2252) & (!ax28x) & (g2218) & (g2255)) + ((!g2252) & (ax28x) & (!g2218) & (!g2255)) + ((!g2252) & (ax28x) & (!g2218) & (g2255)) + ((g2252) & (!ax28x) & (!g2218) & (!g2255)) + ((g2252) & (!ax28x) & (g2218) & (!g2255)) + ((g2252) & (ax28x) & (g2218) & (!g2255)) + ((g2252) & (ax28x) & (g2218) & (g2255)));
	assign g2349 = (((!ax28x) & (!ax29x) & (!g2218) & (!g2274) & (!g2295) & (g2348)) + ((!ax28x) & (!ax29x) & (!g2218) & (!g2274) & (g2295) & (!g2348)) + ((!ax28x) & (!ax29x) & (!g2218) & (!g2274) & (g2295) & (g2348)) + ((!ax28x) & (!ax29x) & (!g2218) & (g2274) & (!g2295) & (g2348)) + ((!ax28x) & (!ax29x) & (!g2218) & (g2274) & (g2295) & (g2348)) + ((!ax28x) & (!ax29x) & (g2218) & (!g2274) & (!g2295) & (!g2348)) + ((!ax28x) & (!ax29x) & (g2218) & (g2274) & (!g2295) & (!g2348)) + ((!ax28x) & (!ax29x) & (g2218) & (g2274) & (g2295) & (!g2348)) + ((!ax28x) & (ax29x) & (!g2218) & (!g2274) & (!g2295) & (!g2348)) + ((!ax28x) & (ax29x) & (!g2218) & (g2274) & (!g2295) & (!g2348)) + ((!ax28x) & (ax29x) & (!g2218) & (g2274) & (g2295) & (!g2348)) + ((!ax28x) & (ax29x) & (g2218) & (!g2274) & (!g2295) & (g2348)) + ((!ax28x) & (ax29x) & (g2218) & (!g2274) & (g2295) & (!g2348)) + ((!ax28x) & (ax29x) & (g2218) & (!g2274) & (g2295) & (g2348)) + ((!ax28x) & (ax29x) & (g2218) & (g2274) & (!g2295) & (g2348)) + ((!ax28x) & (ax29x) & (g2218) & (g2274) & (g2295) & (g2348)) + ((ax28x) & (!ax29x) & (!g2218) & (!g2274) & (!g2295) & (!g2348)) + ((ax28x) & (!ax29x) & (!g2218) & (g2274) & (!g2295) & (!g2348)) + ((ax28x) & (!ax29x) & (!g2218) & (g2274) & (g2295) & (!g2348)) + ((ax28x) & (!ax29x) & (g2218) & (!g2274) & (!g2295) & (!g2348)) + ((ax28x) & (!ax29x) & (g2218) & (g2274) & (!g2295) & (!g2348)) + ((ax28x) & (!ax29x) & (g2218) & (g2274) & (g2295) & (!g2348)) + ((ax28x) & (ax29x) & (!g2218) & (!g2274) & (!g2295) & (g2348)) + ((ax28x) & (ax29x) & (!g2218) & (!g2274) & (g2295) & (!g2348)) + ((ax28x) & (ax29x) & (!g2218) & (!g2274) & (g2295) & (g2348)) + ((ax28x) & (ax29x) & (!g2218) & (g2274) & (!g2295) & (g2348)) + ((ax28x) & (ax29x) & (!g2218) & (g2274) & (g2295) & (g2348)) + ((ax28x) & (ax29x) & (g2218) & (!g2274) & (!g2295) & (g2348)) + ((ax28x) & (ax29x) & (g2218) & (!g2274) & (g2295) & (!g2348)) + ((ax28x) & (ax29x) & (g2218) & (!g2274) & (g2295) & (g2348)) + ((ax28x) & (ax29x) & (g2218) & (g2274) & (!g2295) & (g2348)) + ((ax28x) & (ax29x) & (g2218) & (g2274) & (g2295) & (g2348)));
	assign g2350 = (((!ax28x) & (!g2218) & (!g2255) & (!g2274) & (g2295)) + ((!ax28x) & (!g2218) & (g2255) & (!g2274) & (!g2295)) + ((!ax28x) & (!g2218) & (g2255) & (!g2274) & (g2295)) + ((!ax28x) & (!g2218) & (g2255) & (g2274) & (!g2295)) + ((!ax28x) & (!g2218) & (g2255) & (g2274) & (g2295)) + ((!ax28x) & (g2218) & (g2255) & (!g2274) & (!g2295)) + ((!ax28x) & (g2218) & (g2255) & (g2274) & (!g2295)) + ((!ax28x) & (g2218) & (g2255) & (g2274) & (g2295)) + ((ax28x) & (!g2218) & (!g2255) & (!g2274) & (!g2295)) + ((ax28x) & (!g2218) & (!g2255) & (g2274) & (!g2295)) + ((ax28x) & (!g2218) & (!g2255) & (g2274) & (g2295)) + ((ax28x) & (g2218) & (!g2255) & (!g2274) & (!g2295)) + ((ax28x) & (g2218) & (!g2255) & (!g2274) & (g2295)) + ((ax28x) & (g2218) & (!g2255) & (g2274) & (!g2295)) + ((ax28x) & (g2218) & (!g2255) & (g2274) & (g2295)) + ((ax28x) & (g2218) & (g2255) & (!g2274) & (g2295)));
	assign g2351 = (((!ax24x) & (!ax25x)));
	assign g2352 = (((!g2218) & (!ax26x) & (!ax27x) & (!g2274) & (!g2295) & (!g2351)) + ((!g2218) & (!ax26x) & (!ax27x) & (g2274) & (!g2295) & (!g2351)) + ((!g2218) & (!ax26x) & (!ax27x) & (g2274) & (g2295) & (!g2351)) + ((!g2218) & (!ax26x) & (ax27x) & (!g2274) & (g2295) & (!g2351)) + ((!g2218) & (ax26x) & (ax27x) & (!g2274) & (g2295) & (!g2351)) + ((!g2218) & (ax26x) & (ax27x) & (!g2274) & (g2295) & (g2351)) + ((g2218) & (!ax26x) & (!ax27x) & (!g2274) & (!g2295) & (!g2351)) + ((g2218) & (!ax26x) & (!ax27x) & (!g2274) & (!g2295) & (g2351)) + ((g2218) & (!ax26x) & (!ax27x) & (!g2274) & (g2295) & (!g2351)) + ((g2218) & (!ax26x) & (!ax27x) & (g2274) & (!g2295) & (!g2351)) + ((g2218) & (!ax26x) & (!ax27x) & (g2274) & (!g2295) & (g2351)) + ((g2218) & (!ax26x) & (!ax27x) & (g2274) & (g2295) & (!g2351)) + ((g2218) & (!ax26x) & (!ax27x) & (g2274) & (g2295) & (g2351)) + ((g2218) & (!ax26x) & (ax27x) & (!g2274) & (!g2295) & (!g2351)) + ((g2218) & (!ax26x) & (ax27x) & (!g2274) & (g2295) & (!g2351)) + ((g2218) & (!ax26x) & (ax27x) & (!g2274) & (g2295) & (g2351)) + ((g2218) & (!ax26x) & (ax27x) & (g2274) & (!g2295) & (!g2351)) + ((g2218) & (!ax26x) & (ax27x) & (g2274) & (g2295) & (!g2351)) + ((g2218) & (ax26x) & (!ax27x) & (!g2274) & (g2295) & (!g2351)) + ((g2218) & (ax26x) & (!ax27x) & (!g2274) & (g2295) & (g2351)) + ((g2218) & (ax26x) & (ax27x) & (!g2274) & (!g2295) & (!g2351)) + ((g2218) & (ax26x) & (ax27x) & (!g2274) & (!g2295) & (g2351)) + ((g2218) & (ax26x) & (ax27x) & (!g2274) & (g2295) & (!g2351)) + ((g2218) & (ax26x) & (ax27x) & (!g2274) & (g2295) & (g2351)) + ((g2218) & (ax26x) & (ax27x) & (g2274) & (!g2295) & (!g2351)) + ((g2218) & (ax26x) & (ax27x) & (g2274) & (!g2295) & (g2351)) + ((g2218) & (ax26x) & (ax27x) & (g2274) & (g2295) & (!g2351)) + ((g2218) & (ax26x) & (ax27x) & (g2274) & (g2295) & (g2351)));
	assign g2353 = (((!g2045) & (!g2252) & (g2349) & (g2350) & (g2352)) + ((!g2045) & (g2252) & (g2349) & (!g2350) & (g2352)) + ((!g2045) & (g2252) & (g2349) & (g2350) & (!g2352)) + ((!g2045) & (g2252) & (g2349) & (g2350) & (g2352)) + ((g2045) & (!g2252) & (!g2349) & (g2350) & (g2352)) + ((g2045) & (!g2252) & (g2349) & (!g2350) & (!g2352)) + ((g2045) & (!g2252) & (g2349) & (!g2350) & (g2352)) + ((g2045) & (!g2252) & (g2349) & (g2350) & (!g2352)) + ((g2045) & (!g2252) & (g2349) & (g2350) & (g2352)) + ((g2045) & (g2252) & (!g2349) & (!g2350) & (g2352)) + ((g2045) & (g2252) & (!g2349) & (g2350) & (!g2352)) + ((g2045) & (g2252) & (!g2349) & (g2350) & (g2352)) + ((g2045) & (g2252) & (g2349) & (!g2350) & (!g2352)) + ((g2045) & (g2252) & (g2349) & (!g2350) & (g2352)) + ((g2045) & (g2252) & (g2349) & (g2350) & (!g2352)) + ((g2045) & (g2252) & (g2349) & (g2350) & (g2352)));
	assign g2354 = (((!g1879) & (!g2075) & (g2346) & (g2347) & (g2353)) + ((!g1879) & (g2075) & (g2346) & (!g2347) & (g2353)) + ((!g1879) & (g2075) & (g2346) & (g2347) & (!g2353)) + ((!g1879) & (g2075) & (g2346) & (g2347) & (g2353)) + ((g1879) & (!g2075) & (!g2346) & (g2347) & (g2353)) + ((g1879) & (!g2075) & (g2346) & (!g2347) & (!g2353)) + ((g1879) & (!g2075) & (g2346) & (!g2347) & (g2353)) + ((g1879) & (!g2075) & (g2346) & (g2347) & (!g2353)) + ((g1879) & (!g2075) & (g2346) & (g2347) & (g2353)) + ((g1879) & (g2075) & (!g2346) & (!g2347) & (g2353)) + ((g1879) & (g2075) & (!g2346) & (g2347) & (!g2353)) + ((g1879) & (g2075) & (!g2346) & (g2347) & (g2353)) + ((g1879) & (g2075) & (g2346) & (!g2347) & (!g2353)) + ((g1879) & (g2075) & (g2346) & (!g2347) & (g2353)) + ((g1879) & (g2075) & (g2346) & (g2347) & (!g2353)) + ((g1879) & (g2075) & (g2346) & (g2347) & (g2353)));
	assign g2355 = (((!g1720) & (!g1905) & (g2343) & (g2344) & (g2354)) + ((!g1720) & (g1905) & (g2343) & (!g2344) & (g2354)) + ((!g1720) & (g1905) & (g2343) & (g2344) & (!g2354)) + ((!g1720) & (g1905) & (g2343) & (g2344) & (g2354)) + ((g1720) & (!g1905) & (!g2343) & (g2344) & (g2354)) + ((g1720) & (!g1905) & (g2343) & (!g2344) & (!g2354)) + ((g1720) & (!g1905) & (g2343) & (!g2344) & (g2354)) + ((g1720) & (!g1905) & (g2343) & (g2344) & (!g2354)) + ((g1720) & (!g1905) & (g2343) & (g2344) & (g2354)) + ((g1720) & (g1905) & (!g2343) & (!g2344) & (g2354)) + ((g1720) & (g1905) & (!g2343) & (g2344) & (!g2354)) + ((g1720) & (g1905) & (!g2343) & (g2344) & (g2354)) + ((g1720) & (g1905) & (g2343) & (!g2344) & (!g2354)) + ((g1720) & (g1905) & (g2343) & (!g2344) & (g2354)) + ((g1720) & (g1905) & (g2343) & (g2344) & (!g2354)) + ((g1720) & (g1905) & (g2343) & (g2344) & (g2354)));
	assign g2356 = (((!g1568) & (!g1742) & (g2340) & (g2341) & (g2355)) + ((!g1568) & (g1742) & (g2340) & (!g2341) & (g2355)) + ((!g1568) & (g1742) & (g2340) & (g2341) & (!g2355)) + ((!g1568) & (g1742) & (g2340) & (g2341) & (g2355)) + ((g1568) & (!g1742) & (!g2340) & (g2341) & (g2355)) + ((g1568) & (!g1742) & (g2340) & (!g2341) & (!g2355)) + ((g1568) & (!g1742) & (g2340) & (!g2341) & (g2355)) + ((g1568) & (!g1742) & (g2340) & (g2341) & (!g2355)) + ((g1568) & (!g1742) & (g2340) & (g2341) & (g2355)) + ((g1568) & (g1742) & (!g2340) & (!g2341) & (g2355)) + ((g1568) & (g1742) & (!g2340) & (g2341) & (!g2355)) + ((g1568) & (g1742) & (!g2340) & (g2341) & (g2355)) + ((g1568) & (g1742) & (g2340) & (!g2341) & (!g2355)) + ((g1568) & (g1742) & (g2340) & (!g2341) & (g2355)) + ((g1568) & (g1742) & (g2340) & (g2341) & (!g2355)) + ((g1568) & (g1742) & (g2340) & (g2341) & (g2355)));
	assign g2357 = (((!g1423) & (!g1586) & (g2337) & (g2338) & (g2356)) + ((!g1423) & (g1586) & (g2337) & (!g2338) & (g2356)) + ((!g1423) & (g1586) & (g2337) & (g2338) & (!g2356)) + ((!g1423) & (g1586) & (g2337) & (g2338) & (g2356)) + ((g1423) & (!g1586) & (!g2337) & (g2338) & (g2356)) + ((g1423) & (!g1586) & (g2337) & (!g2338) & (!g2356)) + ((g1423) & (!g1586) & (g2337) & (!g2338) & (g2356)) + ((g1423) & (!g1586) & (g2337) & (g2338) & (!g2356)) + ((g1423) & (!g1586) & (g2337) & (g2338) & (g2356)) + ((g1423) & (g1586) & (!g2337) & (!g2338) & (g2356)) + ((g1423) & (g1586) & (!g2337) & (g2338) & (!g2356)) + ((g1423) & (g1586) & (!g2337) & (g2338) & (g2356)) + ((g1423) & (g1586) & (g2337) & (!g2338) & (!g2356)) + ((g1423) & (g1586) & (g2337) & (!g2338) & (g2356)) + ((g1423) & (g1586) & (g2337) & (g2338) & (!g2356)) + ((g1423) & (g1586) & (g2337) & (g2338) & (g2356)));
	assign g2358 = (((!g1285) & (!g1437) & (g2334) & (g2335) & (g2357)) + ((!g1285) & (g1437) & (g2334) & (!g2335) & (g2357)) + ((!g1285) & (g1437) & (g2334) & (g2335) & (!g2357)) + ((!g1285) & (g1437) & (g2334) & (g2335) & (g2357)) + ((g1285) & (!g1437) & (!g2334) & (g2335) & (g2357)) + ((g1285) & (!g1437) & (g2334) & (!g2335) & (!g2357)) + ((g1285) & (!g1437) & (g2334) & (!g2335) & (g2357)) + ((g1285) & (!g1437) & (g2334) & (g2335) & (!g2357)) + ((g1285) & (!g1437) & (g2334) & (g2335) & (g2357)) + ((g1285) & (g1437) & (!g2334) & (!g2335) & (g2357)) + ((g1285) & (g1437) & (!g2334) & (g2335) & (!g2357)) + ((g1285) & (g1437) & (!g2334) & (g2335) & (g2357)) + ((g1285) & (g1437) & (g2334) & (!g2335) & (!g2357)) + ((g1285) & (g1437) & (g2334) & (!g2335) & (g2357)) + ((g1285) & (g1437) & (g2334) & (g2335) & (!g2357)) + ((g1285) & (g1437) & (g2334) & (g2335) & (g2357)));
	assign g2359 = (((!g1154) & (!g1295) & (g2331) & (g2332) & (g2358)) + ((!g1154) & (g1295) & (g2331) & (!g2332) & (g2358)) + ((!g1154) & (g1295) & (g2331) & (g2332) & (!g2358)) + ((!g1154) & (g1295) & (g2331) & (g2332) & (g2358)) + ((g1154) & (!g1295) & (!g2331) & (g2332) & (g2358)) + ((g1154) & (!g1295) & (g2331) & (!g2332) & (!g2358)) + ((g1154) & (!g1295) & (g2331) & (!g2332) & (g2358)) + ((g1154) & (!g1295) & (g2331) & (g2332) & (!g2358)) + ((g1154) & (!g1295) & (g2331) & (g2332) & (g2358)) + ((g1154) & (g1295) & (!g2331) & (!g2332) & (g2358)) + ((g1154) & (g1295) & (!g2331) & (g2332) & (!g2358)) + ((g1154) & (g1295) & (!g2331) & (g2332) & (g2358)) + ((g1154) & (g1295) & (g2331) & (!g2332) & (!g2358)) + ((g1154) & (g1295) & (g2331) & (!g2332) & (g2358)) + ((g1154) & (g1295) & (g2331) & (g2332) & (!g2358)) + ((g1154) & (g1295) & (g2331) & (g2332) & (g2358)));
	assign g2360 = (((!g1030) & (!g1160) & (g2328) & (g2329) & (g2359)) + ((!g1030) & (g1160) & (g2328) & (!g2329) & (g2359)) + ((!g1030) & (g1160) & (g2328) & (g2329) & (!g2359)) + ((!g1030) & (g1160) & (g2328) & (g2329) & (g2359)) + ((g1030) & (!g1160) & (!g2328) & (g2329) & (g2359)) + ((g1030) & (!g1160) & (g2328) & (!g2329) & (!g2359)) + ((g1030) & (!g1160) & (g2328) & (!g2329) & (g2359)) + ((g1030) & (!g1160) & (g2328) & (g2329) & (!g2359)) + ((g1030) & (!g1160) & (g2328) & (g2329) & (g2359)) + ((g1030) & (g1160) & (!g2328) & (!g2329) & (g2359)) + ((g1030) & (g1160) & (!g2328) & (g2329) & (!g2359)) + ((g1030) & (g1160) & (!g2328) & (g2329) & (g2359)) + ((g1030) & (g1160) & (g2328) & (!g2329) & (!g2359)) + ((g1030) & (g1160) & (g2328) & (!g2329) & (g2359)) + ((g1030) & (g1160) & (g2328) & (g2329) & (!g2359)) + ((g1030) & (g1160) & (g2328) & (g2329) & (g2359)));
	assign g2361 = (((!g914) & (!g1032) & (g2325) & (g2326) & (g2360)) + ((!g914) & (g1032) & (g2325) & (!g2326) & (g2360)) + ((!g914) & (g1032) & (g2325) & (g2326) & (!g2360)) + ((!g914) & (g1032) & (g2325) & (g2326) & (g2360)) + ((g914) & (!g1032) & (!g2325) & (g2326) & (g2360)) + ((g914) & (!g1032) & (g2325) & (!g2326) & (!g2360)) + ((g914) & (!g1032) & (g2325) & (!g2326) & (g2360)) + ((g914) & (!g1032) & (g2325) & (g2326) & (!g2360)) + ((g914) & (!g1032) & (g2325) & (g2326) & (g2360)) + ((g914) & (g1032) & (!g2325) & (!g2326) & (g2360)) + ((g914) & (g1032) & (!g2325) & (g2326) & (!g2360)) + ((g914) & (g1032) & (!g2325) & (g2326) & (g2360)) + ((g914) & (g1032) & (g2325) & (!g2326) & (!g2360)) + ((g914) & (g1032) & (g2325) & (!g2326) & (g2360)) + ((g914) & (g1032) & (g2325) & (g2326) & (!g2360)) + ((g914) & (g1032) & (g2325) & (g2326) & (g2360)));
	assign g2362 = (((!g803) & (!g851) & (g2322) & (g2323) & (g2361)) + ((!g803) & (g851) & (g2322) & (!g2323) & (g2361)) + ((!g803) & (g851) & (g2322) & (g2323) & (!g2361)) + ((!g803) & (g851) & (g2322) & (g2323) & (g2361)) + ((g803) & (!g851) & (!g2322) & (g2323) & (g2361)) + ((g803) & (!g851) & (g2322) & (!g2323) & (!g2361)) + ((g803) & (!g851) & (g2322) & (!g2323) & (g2361)) + ((g803) & (!g851) & (g2322) & (g2323) & (!g2361)) + ((g803) & (!g851) & (g2322) & (g2323) & (g2361)) + ((g803) & (g851) & (!g2322) & (!g2323) & (g2361)) + ((g803) & (g851) & (!g2322) & (g2323) & (!g2361)) + ((g803) & (g851) & (!g2322) & (g2323) & (g2361)) + ((g803) & (g851) & (g2322) & (!g2323) & (!g2361)) + ((g803) & (g851) & (g2322) & (!g2323) & (g2361)) + ((g803) & (g851) & (g2322) & (g2323) & (!g2361)) + ((g803) & (g851) & (g2322) & (g2323) & (g2361)));
	assign g2363 = (((!g700) & (!g744) & (g2319) & (g2320) & (g2362)) + ((!g700) & (g744) & (g2319) & (!g2320) & (g2362)) + ((!g700) & (g744) & (g2319) & (g2320) & (!g2362)) + ((!g700) & (g744) & (g2319) & (g2320) & (g2362)) + ((g700) & (!g744) & (!g2319) & (g2320) & (g2362)) + ((g700) & (!g744) & (g2319) & (!g2320) & (!g2362)) + ((g700) & (!g744) & (g2319) & (!g2320) & (g2362)) + ((g700) & (!g744) & (g2319) & (g2320) & (!g2362)) + ((g700) & (!g744) & (g2319) & (g2320) & (g2362)) + ((g700) & (g744) & (!g2319) & (!g2320) & (g2362)) + ((g700) & (g744) & (!g2319) & (g2320) & (!g2362)) + ((g700) & (g744) & (!g2319) & (g2320) & (g2362)) + ((g700) & (g744) & (g2319) & (!g2320) & (!g2362)) + ((g700) & (g744) & (g2319) & (!g2320) & (g2362)) + ((g700) & (g744) & (g2319) & (g2320) & (!g2362)) + ((g700) & (g744) & (g2319) & (g2320) & (g2362)));
	assign g2364 = (((!g604) & (!g645) & (g2316) & (g2317) & (g2363)) + ((!g604) & (g645) & (g2316) & (!g2317) & (g2363)) + ((!g604) & (g645) & (g2316) & (g2317) & (!g2363)) + ((!g604) & (g645) & (g2316) & (g2317) & (g2363)) + ((g604) & (!g645) & (!g2316) & (g2317) & (g2363)) + ((g604) & (!g645) & (g2316) & (!g2317) & (!g2363)) + ((g604) & (!g645) & (g2316) & (!g2317) & (g2363)) + ((g604) & (!g645) & (g2316) & (g2317) & (!g2363)) + ((g604) & (!g645) & (g2316) & (g2317) & (g2363)) + ((g604) & (g645) & (!g2316) & (!g2317) & (g2363)) + ((g604) & (g645) & (!g2316) & (g2317) & (!g2363)) + ((g604) & (g645) & (!g2316) & (g2317) & (g2363)) + ((g604) & (g645) & (g2316) & (!g2317) & (!g2363)) + ((g604) & (g645) & (g2316) & (!g2317) & (g2363)) + ((g604) & (g645) & (g2316) & (g2317) & (!g2363)) + ((g604) & (g645) & (g2316) & (g2317) & (g2363)));
	assign g2365 = (((!g515) & (!g553) & (g2313) & (g2314) & (g2364)) + ((!g515) & (g553) & (g2313) & (!g2314) & (g2364)) + ((!g515) & (g553) & (g2313) & (g2314) & (!g2364)) + ((!g515) & (g553) & (g2313) & (g2314) & (g2364)) + ((g515) & (!g553) & (!g2313) & (g2314) & (g2364)) + ((g515) & (!g553) & (g2313) & (!g2314) & (!g2364)) + ((g515) & (!g553) & (g2313) & (!g2314) & (g2364)) + ((g515) & (!g553) & (g2313) & (g2314) & (!g2364)) + ((g515) & (!g553) & (g2313) & (g2314) & (g2364)) + ((g515) & (g553) & (!g2313) & (!g2314) & (g2364)) + ((g515) & (g553) & (!g2313) & (g2314) & (!g2364)) + ((g515) & (g553) & (!g2313) & (g2314) & (g2364)) + ((g515) & (g553) & (g2313) & (!g2314) & (!g2364)) + ((g515) & (g553) & (g2313) & (!g2314) & (g2364)) + ((g515) & (g553) & (g2313) & (g2314) & (!g2364)) + ((g515) & (g553) & (g2313) & (g2314) & (g2364)));
	assign g2366 = (((!g433) & (!g468) & (g2310) & (g2311) & (g2365)) + ((!g433) & (g468) & (g2310) & (!g2311) & (g2365)) + ((!g433) & (g468) & (g2310) & (g2311) & (!g2365)) + ((!g433) & (g468) & (g2310) & (g2311) & (g2365)) + ((g433) & (!g468) & (!g2310) & (g2311) & (g2365)) + ((g433) & (!g468) & (g2310) & (!g2311) & (!g2365)) + ((g433) & (!g468) & (g2310) & (!g2311) & (g2365)) + ((g433) & (!g468) & (g2310) & (g2311) & (!g2365)) + ((g433) & (!g468) & (g2310) & (g2311) & (g2365)) + ((g433) & (g468) & (!g2310) & (!g2311) & (g2365)) + ((g433) & (g468) & (!g2310) & (g2311) & (!g2365)) + ((g433) & (g468) & (!g2310) & (g2311) & (g2365)) + ((g433) & (g468) & (g2310) & (!g2311) & (!g2365)) + ((g433) & (g468) & (g2310) & (!g2311) & (g2365)) + ((g433) & (g468) & (g2310) & (g2311) & (!g2365)) + ((g433) & (g468) & (g2310) & (g2311) & (g2365)));
	assign g2367 = (((!g358) & (!g390) & (g2307) & (g2308) & (g2366)) + ((!g358) & (g390) & (g2307) & (!g2308) & (g2366)) + ((!g358) & (g390) & (g2307) & (g2308) & (!g2366)) + ((!g358) & (g390) & (g2307) & (g2308) & (g2366)) + ((g358) & (!g390) & (!g2307) & (g2308) & (g2366)) + ((g358) & (!g390) & (g2307) & (!g2308) & (!g2366)) + ((g358) & (!g390) & (g2307) & (!g2308) & (g2366)) + ((g358) & (!g390) & (g2307) & (g2308) & (!g2366)) + ((g358) & (!g390) & (g2307) & (g2308) & (g2366)) + ((g358) & (g390) & (!g2307) & (!g2308) & (g2366)) + ((g358) & (g390) & (!g2307) & (g2308) & (!g2366)) + ((g358) & (g390) & (!g2307) & (g2308) & (g2366)) + ((g358) & (g390) & (g2307) & (!g2308) & (!g2366)) + ((g358) & (g390) & (g2307) & (!g2308) & (g2366)) + ((g358) & (g390) & (g2307) & (g2308) & (!g2366)) + ((g358) & (g390) & (g2307) & (g2308) & (g2366)));
	assign g2368 = (((!g290) & (!g319) & (g2304) & (g2305) & (g2367)) + ((!g290) & (g319) & (g2304) & (!g2305) & (g2367)) + ((!g290) & (g319) & (g2304) & (g2305) & (!g2367)) + ((!g290) & (g319) & (g2304) & (g2305) & (g2367)) + ((g290) & (!g319) & (!g2304) & (g2305) & (g2367)) + ((g290) & (!g319) & (g2304) & (!g2305) & (!g2367)) + ((g290) & (!g319) & (g2304) & (!g2305) & (g2367)) + ((g290) & (!g319) & (g2304) & (g2305) & (!g2367)) + ((g290) & (!g319) & (g2304) & (g2305) & (g2367)) + ((g290) & (g319) & (!g2304) & (!g2305) & (g2367)) + ((g290) & (g319) & (!g2304) & (g2305) & (!g2367)) + ((g290) & (g319) & (!g2304) & (g2305) & (g2367)) + ((g290) & (g319) & (g2304) & (!g2305) & (!g2367)) + ((g290) & (g319) & (g2304) & (!g2305) & (g2367)) + ((g290) & (g319) & (g2304) & (g2305) & (!g2367)) + ((g290) & (g319) & (g2304) & (g2305) & (g2367)));
	assign g2369 = (((!g229) & (!g255) & (g2301) & (g2302) & (g2368)) + ((!g229) & (g255) & (g2301) & (!g2302) & (g2368)) + ((!g229) & (g255) & (g2301) & (g2302) & (!g2368)) + ((!g229) & (g255) & (g2301) & (g2302) & (g2368)) + ((g229) & (!g255) & (!g2301) & (g2302) & (g2368)) + ((g229) & (!g255) & (g2301) & (!g2302) & (!g2368)) + ((g229) & (!g255) & (g2301) & (!g2302) & (g2368)) + ((g229) & (!g255) & (g2301) & (g2302) & (!g2368)) + ((g229) & (!g255) & (g2301) & (g2302) & (g2368)) + ((g229) & (g255) & (!g2301) & (!g2302) & (g2368)) + ((g229) & (g255) & (!g2301) & (g2302) & (!g2368)) + ((g229) & (g255) & (!g2301) & (g2302) & (g2368)) + ((g229) & (g255) & (g2301) & (!g2302) & (!g2368)) + ((g229) & (g255) & (g2301) & (!g2302) & (g2368)) + ((g229) & (g255) & (g2301) & (g2302) & (!g2368)) + ((g229) & (g255) & (g2301) & (g2302) & (g2368)));
	assign g2370 = (((!g174) & (!g198) & (g2298) & (g2299) & (g2369)) + ((!g174) & (g198) & (g2298) & (!g2299) & (g2369)) + ((!g174) & (g198) & (g2298) & (g2299) & (!g2369)) + ((!g174) & (g198) & (g2298) & (g2299) & (g2369)) + ((g174) & (!g198) & (!g2298) & (g2299) & (g2369)) + ((g174) & (!g198) & (g2298) & (!g2299) & (!g2369)) + ((g174) & (!g198) & (g2298) & (!g2299) & (g2369)) + ((g174) & (!g198) & (g2298) & (g2299) & (!g2369)) + ((g174) & (!g198) & (g2298) & (g2299) & (g2369)) + ((g174) & (g198) & (!g2298) & (!g2299) & (g2369)) + ((g174) & (g198) & (!g2298) & (g2299) & (!g2369)) + ((g174) & (g198) & (!g2298) & (g2299) & (g2369)) + ((g174) & (g198) & (g2298) & (!g2299) & (!g2369)) + ((g174) & (g198) & (g2298) & (!g2299) & (g2369)) + ((g174) & (g198) & (g2298) & (g2299) & (!g2369)) + ((g174) & (g198) & (g2298) & (g2299) & (g2369)));
	assign g2371 = (((!g4) & (!g2292) & (!g2293) & (!g2274) & (!g2295)) + ((!g4) & (!g2292) & (!g2293) & (g2274) & (!g2295)) + ((!g4) & (!g2292) & (!g2293) & (g2274) & (g2295)) + ((!g4) & (!g2292) & (g2293) & (!g2274) & (g2295)) + ((!g4) & (g2292) & (g2293) & (!g2274) & (!g2295)) + ((!g4) & (g2292) & (g2293) & (!g2274) & (g2295)) + ((!g4) & (g2292) & (g2293) & (g2274) & (!g2295)) + ((!g4) & (g2292) & (g2293) & (g2274) & (g2295)) + ((g4) & (!g2292) & (g2293) & (!g2274) & (!g2295)) + ((g4) & (!g2292) & (g2293) & (!g2274) & (g2295)) + ((g4) & (!g2292) & (g2293) & (g2274) & (!g2295)) + ((g4) & (!g2292) & (g2293) & (g2274) & (g2295)) + ((g4) & (g2292) & (!g2293) & (!g2274) & (!g2295)) + ((g4) & (g2292) & (!g2293) & (g2274) & (!g2295)) + ((g4) & (g2292) & (!g2293) & (g2274) & (g2295)) + ((g4) & (g2292) & (g2293) & (!g2274) & (g2295)));
	assign g2372 = (((!g8) & (!g2277) & (g2291) & (!g2274) & (!g2295)) + ((!g8) & (!g2277) & (g2291) & (g2274) & (!g2295)) + ((!g8) & (!g2277) & (g2291) & (g2274) & (g2295)) + ((!g8) & (g2277) & (!g2291) & (!g2274) & (!g2295)) + ((!g8) & (g2277) & (!g2291) & (!g2274) & (g2295)) + ((!g8) & (g2277) & (!g2291) & (g2274) & (!g2295)) + ((!g8) & (g2277) & (!g2291) & (g2274) & (g2295)) + ((!g8) & (g2277) & (g2291) & (!g2274) & (g2295)) + ((g8) & (!g2277) & (!g2291) & (!g2274) & (!g2295)) + ((g8) & (!g2277) & (!g2291) & (g2274) & (!g2295)) + ((g8) & (!g2277) & (!g2291) & (g2274) & (g2295)) + ((g8) & (g2277) & (!g2291) & (!g2274) & (g2295)) + ((g8) & (g2277) & (g2291) & (!g2274) & (!g2295)) + ((g8) & (g2277) & (g2291) & (!g2274) & (g2295)) + ((g8) & (g2277) & (g2291) & (g2274) & (!g2295)) + ((g8) & (g2277) & (g2291) & (g2274) & (g2295)));
	assign g2373 = (((!g18) & (!g27) & (g2279) & (g2290)) + ((!g18) & (g27) & (!g2279) & (g2290)) + ((!g18) & (g27) & (g2279) & (!g2290)) + ((!g18) & (g27) & (g2279) & (g2290)) + ((g18) & (!g27) & (!g2279) & (!g2290)) + ((g18) & (!g27) & (!g2279) & (g2290)) + ((g18) & (!g27) & (g2279) & (!g2290)) + ((g18) & (g27) & (!g2279) & (!g2290)));
	assign g2374 = (((!g2278) & (!g2274) & (!g2295) & (g2373)) + ((!g2278) & (g2274) & (!g2295) & (g2373)) + ((!g2278) & (g2274) & (g2295) & (g2373)) + ((g2278) & (!g2274) & (!g2295) & (!g2373)) + ((g2278) & (!g2274) & (g2295) & (!g2373)) + ((g2278) & (!g2274) & (g2295) & (g2373)) + ((g2278) & (g2274) & (!g2295) & (!g2373)) + ((g2278) & (g2274) & (g2295) & (!g2373)));
	assign g2375 = (((!g27) & (!g2279) & (g2290) & (!g2274) & (!g2295)) + ((!g27) & (!g2279) & (g2290) & (g2274) & (!g2295)) + ((!g27) & (!g2279) & (g2290) & (g2274) & (g2295)) + ((!g27) & (g2279) & (!g2290) & (!g2274) & (!g2295)) + ((!g27) & (g2279) & (!g2290) & (!g2274) & (g2295)) + ((!g27) & (g2279) & (!g2290) & (g2274) & (!g2295)) + ((!g27) & (g2279) & (!g2290) & (g2274) & (g2295)) + ((!g27) & (g2279) & (g2290) & (!g2274) & (g2295)) + ((g27) & (!g2279) & (!g2290) & (!g2274) & (!g2295)) + ((g27) & (!g2279) & (!g2290) & (g2274) & (!g2295)) + ((g27) & (!g2279) & (!g2290) & (g2274) & (g2295)) + ((g27) & (g2279) & (!g2290) & (!g2274) & (g2295)) + ((g27) & (g2279) & (g2290) & (!g2274) & (!g2295)) + ((g27) & (g2279) & (g2290) & (!g2274) & (g2295)) + ((g27) & (g2279) & (g2290) & (g2274) & (!g2295)) + ((g27) & (g2279) & (g2290) & (g2274) & (g2295)));
	assign g2376 = (((!g39) & (!g54) & (g2281) & (g2289)) + ((!g39) & (g54) & (!g2281) & (g2289)) + ((!g39) & (g54) & (g2281) & (!g2289)) + ((!g39) & (g54) & (g2281) & (g2289)) + ((g39) & (!g54) & (!g2281) & (!g2289)) + ((g39) & (!g54) & (!g2281) & (g2289)) + ((g39) & (!g54) & (g2281) & (!g2289)) + ((g39) & (g54) & (!g2281) & (!g2289)));
	assign g2377 = (((!g2280) & (!g2274) & (!g2295) & (g2376)) + ((!g2280) & (g2274) & (!g2295) & (g2376)) + ((!g2280) & (g2274) & (g2295) & (g2376)) + ((g2280) & (!g2274) & (!g2295) & (!g2376)) + ((g2280) & (!g2274) & (g2295) & (!g2376)) + ((g2280) & (!g2274) & (g2295) & (g2376)) + ((g2280) & (g2274) & (!g2295) & (!g2376)) + ((g2280) & (g2274) & (g2295) & (!g2376)));
	assign g2378 = (((!g54) & (!g2281) & (g2289) & (!g2274) & (!g2295)) + ((!g54) & (!g2281) & (g2289) & (g2274) & (!g2295)) + ((!g54) & (!g2281) & (g2289) & (g2274) & (g2295)) + ((!g54) & (g2281) & (!g2289) & (!g2274) & (!g2295)) + ((!g54) & (g2281) & (!g2289) & (!g2274) & (g2295)) + ((!g54) & (g2281) & (!g2289) & (g2274) & (!g2295)) + ((!g54) & (g2281) & (!g2289) & (g2274) & (g2295)) + ((!g54) & (g2281) & (g2289) & (!g2274) & (g2295)) + ((g54) & (!g2281) & (!g2289) & (!g2274) & (!g2295)) + ((g54) & (!g2281) & (!g2289) & (g2274) & (!g2295)) + ((g54) & (!g2281) & (!g2289) & (g2274) & (g2295)) + ((g54) & (g2281) & (!g2289) & (!g2274) & (g2295)) + ((g54) & (g2281) & (g2289) & (!g2274) & (!g2295)) + ((g54) & (g2281) & (g2289) & (!g2274) & (g2295)) + ((g54) & (g2281) & (g2289) & (g2274) & (!g2295)) + ((g54) & (g2281) & (g2289) & (g2274) & (g2295)));
	assign g2379 = (((!g68) & (!g87) & (g2283) & (g2288)) + ((!g68) & (g87) & (!g2283) & (g2288)) + ((!g68) & (g87) & (g2283) & (!g2288)) + ((!g68) & (g87) & (g2283) & (g2288)) + ((g68) & (!g87) & (!g2283) & (!g2288)) + ((g68) & (!g87) & (!g2283) & (g2288)) + ((g68) & (!g87) & (g2283) & (!g2288)) + ((g68) & (g87) & (!g2283) & (!g2288)));
	assign g2380 = (((!g2282) & (!g2274) & (!g2295) & (g2379)) + ((!g2282) & (g2274) & (!g2295) & (g2379)) + ((!g2282) & (g2274) & (g2295) & (g2379)) + ((g2282) & (!g2274) & (!g2295) & (!g2379)) + ((g2282) & (!g2274) & (g2295) & (!g2379)) + ((g2282) & (!g2274) & (g2295) & (g2379)) + ((g2282) & (g2274) & (!g2295) & (!g2379)) + ((g2282) & (g2274) & (g2295) & (!g2379)));
	assign g2381 = (((!g87) & (!g2283) & (g2288) & (!g2274) & (!g2295)) + ((!g87) & (!g2283) & (g2288) & (g2274) & (!g2295)) + ((!g87) & (!g2283) & (g2288) & (g2274) & (g2295)) + ((!g87) & (g2283) & (!g2288) & (!g2274) & (!g2295)) + ((!g87) & (g2283) & (!g2288) & (!g2274) & (g2295)) + ((!g87) & (g2283) & (!g2288) & (g2274) & (!g2295)) + ((!g87) & (g2283) & (!g2288) & (g2274) & (g2295)) + ((!g87) & (g2283) & (g2288) & (!g2274) & (g2295)) + ((g87) & (!g2283) & (!g2288) & (!g2274) & (!g2295)) + ((g87) & (!g2283) & (!g2288) & (g2274) & (!g2295)) + ((g87) & (!g2283) & (!g2288) & (g2274) & (g2295)) + ((g87) & (g2283) & (!g2288) & (!g2274) & (g2295)) + ((g87) & (g2283) & (g2288) & (!g2274) & (!g2295)) + ((g87) & (g2283) & (g2288) & (!g2274) & (g2295)) + ((g87) & (g2283) & (g2288) & (g2274) & (!g2295)) + ((g87) & (g2283) & (g2288) & (g2274) & (g2295)));
	assign g2382 = (((!g104) & (!g127) & (g2285) & (g2287)) + ((!g104) & (g127) & (!g2285) & (g2287)) + ((!g104) & (g127) & (g2285) & (!g2287)) + ((!g104) & (g127) & (g2285) & (g2287)) + ((g104) & (!g127) & (!g2285) & (!g2287)) + ((g104) & (!g127) & (!g2285) & (g2287)) + ((g104) & (!g127) & (g2285) & (!g2287)) + ((g104) & (g127) & (!g2285) & (!g2287)));
	assign g2383 = (((!g2284) & (!g2274) & (!g2295) & (g2382)) + ((!g2284) & (g2274) & (!g2295) & (g2382)) + ((!g2284) & (g2274) & (g2295) & (g2382)) + ((g2284) & (!g2274) & (!g2295) & (!g2382)) + ((g2284) & (!g2274) & (g2295) & (!g2382)) + ((g2284) & (!g2274) & (g2295) & (g2382)) + ((g2284) & (g2274) & (!g2295) & (!g2382)) + ((g2284) & (g2274) & (g2295) & (!g2382)));
	assign g2384 = (((!g127) & (!g2285) & (g2287) & (!g2274) & (!g2295)) + ((!g127) & (!g2285) & (g2287) & (g2274) & (!g2295)) + ((!g127) & (!g2285) & (g2287) & (g2274) & (g2295)) + ((!g127) & (g2285) & (!g2287) & (!g2274) & (!g2295)) + ((!g127) & (g2285) & (!g2287) & (!g2274) & (g2295)) + ((!g127) & (g2285) & (!g2287) & (g2274) & (!g2295)) + ((!g127) & (g2285) & (!g2287) & (g2274) & (g2295)) + ((!g127) & (g2285) & (g2287) & (!g2274) & (g2295)) + ((g127) & (!g2285) & (!g2287) & (!g2274) & (!g2295)) + ((g127) & (!g2285) & (!g2287) & (g2274) & (!g2295)) + ((g127) & (!g2285) & (!g2287) & (g2274) & (g2295)) + ((g127) & (g2285) & (!g2287) & (!g2274) & (g2295)) + ((g127) & (g2285) & (g2287) & (!g2274) & (!g2295)) + ((g127) & (g2285) & (g2287) & (!g2274) & (g2295)) + ((g127) & (g2285) & (g2287) & (g2274) & (!g2295)) + ((g127) & (g2285) & (g2287) & (g2274) & (g2295)));
	assign g2385 = (((!g147) & (!g174) & (g2219) & (g2273)) + ((!g147) & (g174) & (!g2219) & (g2273)) + ((!g147) & (g174) & (g2219) & (!g2273)) + ((!g147) & (g174) & (g2219) & (g2273)) + ((g147) & (!g174) & (!g2219) & (!g2273)) + ((g147) & (!g174) & (!g2219) & (g2273)) + ((g147) & (!g174) & (g2219) & (!g2273)) + ((g147) & (g174) & (!g2219) & (!g2273)));
	assign g2386 = (((!g2286) & (!g2274) & (!g2295) & (g2385)) + ((!g2286) & (g2274) & (!g2295) & (g2385)) + ((!g2286) & (g2274) & (g2295) & (g2385)) + ((g2286) & (!g2274) & (!g2295) & (!g2385)) + ((g2286) & (!g2274) & (g2295) & (!g2385)) + ((g2286) & (!g2274) & (g2295) & (g2385)) + ((g2286) & (g2274) & (!g2295) & (!g2385)) + ((g2286) & (g2274) & (g2295) & (!g2385)));
	assign g2387 = (((!g127) & (!g147) & (g2386) & (g2296) & (g2370)) + ((!g127) & (g147) & (g2386) & (!g2296) & (g2370)) + ((!g127) & (g147) & (g2386) & (g2296) & (!g2370)) + ((!g127) & (g147) & (g2386) & (g2296) & (g2370)) + ((g127) & (!g147) & (!g2386) & (g2296) & (g2370)) + ((g127) & (!g147) & (g2386) & (!g2296) & (!g2370)) + ((g127) & (!g147) & (g2386) & (!g2296) & (g2370)) + ((g127) & (!g147) & (g2386) & (g2296) & (!g2370)) + ((g127) & (!g147) & (g2386) & (g2296) & (g2370)) + ((g127) & (g147) & (!g2386) & (!g2296) & (g2370)) + ((g127) & (g147) & (!g2386) & (g2296) & (!g2370)) + ((g127) & (g147) & (!g2386) & (g2296) & (g2370)) + ((g127) & (g147) & (g2386) & (!g2296) & (!g2370)) + ((g127) & (g147) & (g2386) & (!g2296) & (g2370)) + ((g127) & (g147) & (g2386) & (g2296) & (!g2370)) + ((g127) & (g147) & (g2386) & (g2296) & (g2370)));
	assign g2388 = (((!g87) & (!g104) & (g2383) & (g2384) & (g2387)) + ((!g87) & (g104) & (g2383) & (!g2384) & (g2387)) + ((!g87) & (g104) & (g2383) & (g2384) & (!g2387)) + ((!g87) & (g104) & (g2383) & (g2384) & (g2387)) + ((g87) & (!g104) & (!g2383) & (g2384) & (g2387)) + ((g87) & (!g104) & (g2383) & (!g2384) & (!g2387)) + ((g87) & (!g104) & (g2383) & (!g2384) & (g2387)) + ((g87) & (!g104) & (g2383) & (g2384) & (!g2387)) + ((g87) & (!g104) & (g2383) & (g2384) & (g2387)) + ((g87) & (g104) & (!g2383) & (!g2384) & (g2387)) + ((g87) & (g104) & (!g2383) & (g2384) & (!g2387)) + ((g87) & (g104) & (!g2383) & (g2384) & (g2387)) + ((g87) & (g104) & (g2383) & (!g2384) & (!g2387)) + ((g87) & (g104) & (g2383) & (!g2384) & (g2387)) + ((g87) & (g104) & (g2383) & (g2384) & (!g2387)) + ((g87) & (g104) & (g2383) & (g2384) & (g2387)));
	assign g2389 = (((!g54) & (!g68) & (g2380) & (g2381) & (g2388)) + ((!g54) & (g68) & (g2380) & (!g2381) & (g2388)) + ((!g54) & (g68) & (g2380) & (g2381) & (!g2388)) + ((!g54) & (g68) & (g2380) & (g2381) & (g2388)) + ((g54) & (!g68) & (!g2380) & (g2381) & (g2388)) + ((g54) & (!g68) & (g2380) & (!g2381) & (!g2388)) + ((g54) & (!g68) & (g2380) & (!g2381) & (g2388)) + ((g54) & (!g68) & (g2380) & (g2381) & (!g2388)) + ((g54) & (!g68) & (g2380) & (g2381) & (g2388)) + ((g54) & (g68) & (!g2380) & (!g2381) & (g2388)) + ((g54) & (g68) & (!g2380) & (g2381) & (!g2388)) + ((g54) & (g68) & (!g2380) & (g2381) & (g2388)) + ((g54) & (g68) & (g2380) & (!g2381) & (!g2388)) + ((g54) & (g68) & (g2380) & (!g2381) & (g2388)) + ((g54) & (g68) & (g2380) & (g2381) & (!g2388)) + ((g54) & (g68) & (g2380) & (g2381) & (g2388)));
	assign g2390 = (((!g27) & (!g39) & (g2377) & (g2378) & (g2389)) + ((!g27) & (g39) & (g2377) & (!g2378) & (g2389)) + ((!g27) & (g39) & (g2377) & (g2378) & (!g2389)) + ((!g27) & (g39) & (g2377) & (g2378) & (g2389)) + ((g27) & (!g39) & (!g2377) & (g2378) & (g2389)) + ((g27) & (!g39) & (g2377) & (!g2378) & (!g2389)) + ((g27) & (!g39) & (g2377) & (!g2378) & (g2389)) + ((g27) & (!g39) & (g2377) & (g2378) & (!g2389)) + ((g27) & (!g39) & (g2377) & (g2378) & (g2389)) + ((g27) & (g39) & (!g2377) & (!g2378) & (g2389)) + ((g27) & (g39) & (!g2377) & (g2378) & (!g2389)) + ((g27) & (g39) & (!g2377) & (g2378) & (g2389)) + ((g27) & (g39) & (g2377) & (!g2378) & (!g2389)) + ((g27) & (g39) & (g2377) & (!g2378) & (g2389)) + ((g27) & (g39) & (g2377) & (g2378) & (!g2389)) + ((g27) & (g39) & (g2377) & (g2378) & (g2389)));
	assign g2391 = (((!g8) & (!g18) & (g2374) & (g2375) & (g2390)) + ((!g8) & (g18) & (g2374) & (!g2375) & (g2390)) + ((!g8) & (g18) & (g2374) & (g2375) & (!g2390)) + ((!g8) & (g18) & (g2374) & (g2375) & (g2390)) + ((g8) & (!g18) & (!g2374) & (g2375) & (g2390)) + ((g8) & (!g18) & (g2374) & (!g2375) & (!g2390)) + ((g8) & (!g18) & (g2374) & (!g2375) & (g2390)) + ((g8) & (!g18) & (g2374) & (g2375) & (!g2390)) + ((g8) & (!g18) & (g2374) & (g2375) & (g2390)) + ((g8) & (g18) & (!g2374) & (!g2375) & (g2390)) + ((g8) & (g18) & (!g2374) & (g2375) & (!g2390)) + ((g8) & (g18) & (!g2374) & (g2375) & (g2390)) + ((g8) & (g18) & (g2374) & (!g2375) & (!g2390)) + ((g8) & (g18) & (g2374) & (!g2375) & (g2390)) + ((g8) & (g18) & (g2374) & (g2375) & (!g2390)) + ((g8) & (g18) & (g2374) & (g2375) & (g2390)));
	assign g2392 = (((!g2) & (!g8) & (g2277) & (g2291)) + ((!g2) & (g8) & (!g2277) & (g2291)) + ((!g2) & (g8) & (g2277) & (!g2291)) + ((!g2) & (g8) & (g2277) & (g2291)) + ((g2) & (!g8) & (!g2277) & (!g2291)) + ((g2) & (!g8) & (!g2277) & (g2291)) + ((g2) & (!g8) & (g2277) & (!g2291)) + ((g2) & (g8) & (!g2277) & (!g2291)));
	assign g2393 = (((!g2276) & (!g2274) & (!g2295) & (g2392)) + ((!g2276) & (g2274) & (!g2295) & (g2392)) + ((!g2276) & (g2274) & (g2295) & (g2392)) + ((g2276) & (!g2274) & (!g2295) & (!g2392)) + ((g2276) & (!g2274) & (g2295) & (!g2392)) + ((g2276) & (!g2274) & (g2295) & (g2392)) + ((g2276) & (g2274) & (!g2295) & (!g2392)) + ((g2276) & (g2274) & (g2295) & (!g2392)));
	assign g2394 = (((!g4) & (!g2) & (!g2372) & (!g2391) & (g2393)) + ((!g4) & (!g2) & (!g2372) & (g2391) & (g2393)) + ((!g4) & (!g2) & (g2372) & (!g2391) & (g2393)) + ((!g4) & (!g2) & (g2372) & (g2391) & (!g2393)) + ((!g4) & (!g2) & (g2372) & (g2391) & (g2393)) + ((!g4) & (g2) & (!g2372) & (!g2391) & (g2393)) + ((!g4) & (g2) & (!g2372) & (g2391) & (!g2393)) + ((!g4) & (g2) & (!g2372) & (g2391) & (g2393)) + ((!g4) & (g2) & (g2372) & (!g2391) & (!g2393)) + ((!g4) & (g2) & (g2372) & (!g2391) & (g2393)) + ((!g4) & (g2) & (g2372) & (g2391) & (!g2393)) + ((!g4) & (g2) & (g2372) & (g2391) & (g2393)) + ((g4) & (!g2) & (g2372) & (g2391) & (g2393)) + ((g4) & (g2) & (!g2372) & (g2391) & (g2393)) + ((g4) & (g2) & (g2372) & (!g2391) & (g2393)) + ((g4) & (g2) & (g2372) & (g2391) & (g2393)));
	assign g2395 = (((!g4) & (!g2292) & (g2293)) + ((!g4) & (g2292) & (!g2293)) + ((!g4) & (g2292) & (g2293)) + ((g4) & (g2292) & (g2293)));
	assign g2396 = (((!g2275) & (!g2395) & (!g2274) & (!g2295)) + ((!g2275) & (!g2395) & (g2274) & (!g2295)) + ((!g2275) & (!g2395) & (g2274) & (g2295)) + ((g2275) & (g2395) & (!g2274) & (!g2295)) + ((g2275) & (g2395) & (!g2274) & (g2295)) + ((g2275) & (g2395) & (g2274) & (!g2295)) + ((g2275) & (g2395) & (g2274) & (g2295)));
	assign g2397 = (((!g1) & (g2275) & (!g2395) & (!g2274) & (g2295)) + ((!g1) & (g2275) & (g2395) & (!g2274) & (g2295)) + ((g1) & (!g2275) & (g2395) & (g2274) & (!g2295)) + ((g1) & (!g2275) & (g2395) & (g2274) & (g2295)) + ((g1) & (g2275) & (!g2395) & (!g2274) & (!g2295)) + ((g1) & (g2275) & (!g2395) & (!g2274) & (g2295)) + ((g1) & (g2275) & (!g2395) & (g2274) & (!g2295)) + ((g1) & (g2275) & (!g2395) & (g2274) & (g2295)) + ((g1) & (g2275) & (g2395) & (!g2274) & (g2295)));
	assign g2398 = (((!g1) & (!g2371) & (!g2394) & (!g2396) & (!g2397)) + ((g1) & (!g2371) & (!g2394) & (!g2396) & (!g2397)) + ((g1) & (!g2371) & (!g2394) & (g2396) & (!g2397)) + ((g1) & (!g2371) & (g2394) & (!g2396) & (!g2397)) + ((g1) & (!g2371) & (g2394) & (g2396) & (!g2397)) + ((g1) & (g2371) & (!g2394) & (!g2396) & (!g2397)) + ((g1) & (g2371) & (!g2394) & (g2396) & (!g2397)));
	assign g2399 = (((!g147) & (!g2296) & (g2370) & (!g2398)) + ((!g147) & (g2296) & (!g2370) & (!g2398)) + ((!g147) & (g2296) & (!g2370) & (g2398)) + ((!g147) & (g2296) & (g2370) & (g2398)) + ((g147) & (!g2296) & (!g2370) & (!g2398)) + ((g147) & (g2296) & (!g2370) & (g2398)) + ((g147) & (g2296) & (g2370) & (!g2398)) + ((g147) & (g2296) & (g2370) & (g2398)));
	assign g2400 = (((!g174) & (!g198) & (!g2298) & (g2299) & (g2369) & (!g2398)) + ((!g174) & (!g198) & (g2298) & (!g2299) & (!g2369) & (!g2398)) + ((!g174) & (!g198) & (g2298) & (!g2299) & (!g2369) & (g2398)) + ((!g174) & (!g198) & (g2298) & (!g2299) & (g2369) & (!g2398)) + ((!g174) & (!g198) & (g2298) & (!g2299) & (g2369) & (g2398)) + ((!g174) & (!g198) & (g2298) & (g2299) & (!g2369) & (!g2398)) + ((!g174) & (!g198) & (g2298) & (g2299) & (!g2369) & (g2398)) + ((!g174) & (!g198) & (g2298) & (g2299) & (g2369) & (g2398)) + ((!g174) & (g198) & (!g2298) & (!g2299) & (g2369) & (!g2398)) + ((!g174) & (g198) & (!g2298) & (g2299) & (!g2369) & (!g2398)) + ((!g174) & (g198) & (!g2298) & (g2299) & (g2369) & (!g2398)) + ((!g174) & (g198) & (g2298) & (!g2299) & (!g2369) & (!g2398)) + ((!g174) & (g198) & (g2298) & (!g2299) & (!g2369) & (g2398)) + ((!g174) & (g198) & (g2298) & (!g2299) & (g2369) & (g2398)) + ((!g174) & (g198) & (g2298) & (g2299) & (!g2369) & (g2398)) + ((!g174) & (g198) & (g2298) & (g2299) & (g2369) & (g2398)) + ((g174) & (!g198) & (!g2298) & (!g2299) & (!g2369) & (!g2398)) + ((g174) & (!g198) & (!g2298) & (!g2299) & (g2369) & (!g2398)) + ((g174) & (!g198) & (!g2298) & (g2299) & (!g2369) & (!g2398)) + ((g174) & (!g198) & (g2298) & (!g2299) & (!g2369) & (g2398)) + ((g174) & (!g198) & (g2298) & (!g2299) & (g2369) & (g2398)) + ((g174) & (!g198) & (g2298) & (g2299) & (!g2369) & (g2398)) + ((g174) & (!g198) & (g2298) & (g2299) & (g2369) & (!g2398)) + ((g174) & (!g198) & (g2298) & (g2299) & (g2369) & (g2398)) + ((g174) & (g198) & (!g2298) & (!g2299) & (!g2369) & (!g2398)) + ((g174) & (g198) & (g2298) & (!g2299) & (!g2369) & (g2398)) + ((g174) & (g198) & (g2298) & (!g2299) & (g2369) & (!g2398)) + ((g174) & (g198) & (g2298) & (!g2299) & (g2369) & (g2398)) + ((g174) & (g198) & (g2298) & (g2299) & (!g2369) & (!g2398)) + ((g174) & (g198) & (g2298) & (g2299) & (!g2369) & (g2398)) + ((g174) & (g198) & (g2298) & (g2299) & (g2369) & (!g2398)) + ((g174) & (g198) & (g2298) & (g2299) & (g2369) & (g2398)));
	assign g2401 = (((!g198) & (!g2299) & (g2369) & (!g2398)) + ((!g198) & (g2299) & (!g2369) & (!g2398)) + ((!g198) & (g2299) & (!g2369) & (g2398)) + ((!g198) & (g2299) & (g2369) & (g2398)) + ((g198) & (!g2299) & (!g2369) & (!g2398)) + ((g198) & (g2299) & (!g2369) & (g2398)) + ((g198) & (g2299) & (g2369) & (!g2398)) + ((g198) & (g2299) & (g2369) & (g2398)));
	assign g2402 = (((!g229) & (!g255) & (!g2301) & (g2302) & (g2368) & (!g2398)) + ((!g229) & (!g255) & (g2301) & (!g2302) & (!g2368) & (!g2398)) + ((!g229) & (!g255) & (g2301) & (!g2302) & (!g2368) & (g2398)) + ((!g229) & (!g255) & (g2301) & (!g2302) & (g2368) & (!g2398)) + ((!g229) & (!g255) & (g2301) & (!g2302) & (g2368) & (g2398)) + ((!g229) & (!g255) & (g2301) & (g2302) & (!g2368) & (!g2398)) + ((!g229) & (!g255) & (g2301) & (g2302) & (!g2368) & (g2398)) + ((!g229) & (!g255) & (g2301) & (g2302) & (g2368) & (g2398)) + ((!g229) & (g255) & (!g2301) & (!g2302) & (g2368) & (!g2398)) + ((!g229) & (g255) & (!g2301) & (g2302) & (!g2368) & (!g2398)) + ((!g229) & (g255) & (!g2301) & (g2302) & (g2368) & (!g2398)) + ((!g229) & (g255) & (g2301) & (!g2302) & (!g2368) & (!g2398)) + ((!g229) & (g255) & (g2301) & (!g2302) & (!g2368) & (g2398)) + ((!g229) & (g255) & (g2301) & (!g2302) & (g2368) & (g2398)) + ((!g229) & (g255) & (g2301) & (g2302) & (!g2368) & (g2398)) + ((!g229) & (g255) & (g2301) & (g2302) & (g2368) & (g2398)) + ((g229) & (!g255) & (!g2301) & (!g2302) & (!g2368) & (!g2398)) + ((g229) & (!g255) & (!g2301) & (!g2302) & (g2368) & (!g2398)) + ((g229) & (!g255) & (!g2301) & (g2302) & (!g2368) & (!g2398)) + ((g229) & (!g255) & (g2301) & (!g2302) & (!g2368) & (g2398)) + ((g229) & (!g255) & (g2301) & (!g2302) & (g2368) & (g2398)) + ((g229) & (!g255) & (g2301) & (g2302) & (!g2368) & (g2398)) + ((g229) & (!g255) & (g2301) & (g2302) & (g2368) & (!g2398)) + ((g229) & (!g255) & (g2301) & (g2302) & (g2368) & (g2398)) + ((g229) & (g255) & (!g2301) & (!g2302) & (!g2368) & (!g2398)) + ((g229) & (g255) & (g2301) & (!g2302) & (!g2368) & (g2398)) + ((g229) & (g255) & (g2301) & (!g2302) & (g2368) & (!g2398)) + ((g229) & (g255) & (g2301) & (!g2302) & (g2368) & (g2398)) + ((g229) & (g255) & (g2301) & (g2302) & (!g2368) & (!g2398)) + ((g229) & (g255) & (g2301) & (g2302) & (!g2368) & (g2398)) + ((g229) & (g255) & (g2301) & (g2302) & (g2368) & (!g2398)) + ((g229) & (g255) & (g2301) & (g2302) & (g2368) & (g2398)));
	assign g2403 = (((!g255) & (!g2302) & (g2368) & (!g2398)) + ((!g255) & (g2302) & (!g2368) & (!g2398)) + ((!g255) & (g2302) & (!g2368) & (g2398)) + ((!g255) & (g2302) & (g2368) & (g2398)) + ((g255) & (!g2302) & (!g2368) & (!g2398)) + ((g255) & (g2302) & (!g2368) & (g2398)) + ((g255) & (g2302) & (g2368) & (!g2398)) + ((g255) & (g2302) & (g2368) & (g2398)));
	assign g2404 = (((!g290) & (!g319) & (!g2304) & (g2305) & (g2367) & (!g2398)) + ((!g290) & (!g319) & (g2304) & (!g2305) & (!g2367) & (!g2398)) + ((!g290) & (!g319) & (g2304) & (!g2305) & (!g2367) & (g2398)) + ((!g290) & (!g319) & (g2304) & (!g2305) & (g2367) & (!g2398)) + ((!g290) & (!g319) & (g2304) & (!g2305) & (g2367) & (g2398)) + ((!g290) & (!g319) & (g2304) & (g2305) & (!g2367) & (!g2398)) + ((!g290) & (!g319) & (g2304) & (g2305) & (!g2367) & (g2398)) + ((!g290) & (!g319) & (g2304) & (g2305) & (g2367) & (g2398)) + ((!g290) & (g319) & (!g2304) & (!g2305) & (g2367) & (!g2398)) + ((!g290) & (g319) & (!g2304) & (g2305) & (!g2367) & (!g2398)) + ((!g290) & (g319) & (!g2304) & (g2305) & (g2367) & (!g2398)) + ((!g290) & (g319) & (g2304) & (!g2305) & (!g2367) & (!g2398)) + ((!g290) & (g319) & (g2304) & (!g2305) & (!g2367) & (g2398)) + ((!g290) & (g319) & (g2304) & (!g2305) & (g2367) & (g2398)) + ((!g290) & (g319) & (g2304) & (g2305) & (!g2367) & (g2398)) + ((!g290) & (g319) & (g2304) & (g2305) & (g2367) & (g2398)) + ((g290) & (!g319) & (!g2304) & (!g2305) & (!g2367) & (!g2398)) + ((g290) & (!g319) & (!g2304) & (!g2305) & (g2367) & (!g2398)) + ((g290) & (!g319) & (!g2304) & (g2305) & (!g2367) & (!g2398)) + ((g290) & (!g319) & (g2304) & (!g2305) & (!g2367) & (g2398)) + ((g290) & (!g319) & (g2304) & (!g2305) & (g2367) & (g2398)) + ((g290) & (!g319) & (g2304) & (g2305) & (!g2367) & (g2398)) + ((g290) & (!g319) & (g2304) & (g2305) & (g2367) & (!g2398)) + ((g290) & (!g319) & (g2304) & (g2305) & (g2367) & (g2398)) + ((g290) & (g319) & (!g2304) & (!g2305) & (!g2367) & (!g2398)) + ((g290) & (g319) & (g2304) & (!g2305) & (!g2367) & (g2398)) + ((g290) & (g319) & (g2304) & (!g2305) & (g2367) & (!g2398)) + ((g290) & (g319) & (g2304) & (!g2305) & (g2367) & (g2398)) + ((g290) & (g319) & (g2304) & (g2305) & (!g2367) & (!g2398)) + ((g290) & (g319) & (g2304) & (g2305) & (!g2367) & (g2398)) + ((g290) & (g319) & (g2304) & (g2305) & (g2367) & (!g2398)) + ((g290) & (g319) & (g2304) & (g2305) & (g2367) & (g2398)));
	assign g2405 = (((!g319) & (!g2305) & (g2367) & (!g2398)) + ((!g319) & (g2305) & (!g2367) & (!g2398)) + ((!g319) & (g2305) & (!g2367) & (g2398)) + ((!g319) & (g2305) & (g2367) & (g2398)) + ((g319) & (!g2305) & (!g2367) & (!g2398)) + ((g319) & (g2305) & (!g2367) & (g2398)) + ((g319) & (g2305) & (g2367) & (!g2398)) + ((g319) & (g2305) & (g2367) & (g2398)));
	assign g2406 = (((!g358) & (!g390) & (!g2307) & (g2308) & (g2366) & (!g2398)) + ((!g358) & (!g390) & (g2307) & (!g2308) & (!g2366) & (!g2398)) + ((!g358) & (!g390) & (g2307) & (!g2308) & (!g2366) & (g2398)) + ((!g358) & (!g390) & (g2307) & (!g2308) & (g2366) & (!g2398)) + ((!g358) & (!g390) & (g2307) & (!g2308) & (g2366) & (g2398)) + ((!g358) & (!g390) & (g2307) & (g2308) & (!g2366) & (!g2398)) + ((!g358) & (!g390) & (g2307) & (g2308) & (!g2366) & (g2398)) + ((!g358) & (!g390) & (g2307) & (g2308) & (g2366) & (g2398)) + ((!g358) & (g390) & (!g2307) & (!g2308) & (g2366) & (!g2398)) + ((!g358) & (g390) & (!g2307) & (g2308) & (!g2366) & (!g2398)) + ((!g358) & (g390) & (!g2307) & (g2308) & (g2366) & (!g2398)) + ((!g358) & (g390) & (g2307) & (!g2308) & (!g2366) & (!g2398)) + ((!g358) & (g390) & (g2307) & (!g2308) & (!g2366) & (g2398)) + ((!g358) & (g390) & (g2307) & (!g2308) & (g2366) & (g2398)) + ((!g358) & (g390) & (g2307) & (g2308) & (!g2366) & (g2398)) + ((!g358) & (g390) & (g2307) & (g2308) & (g2366) & (g2398)) + ((g358) & (!g390) & (!g2307) & (!g2308) & (!g2366) & (!g2398)) + ((g358) & (!g390) & (!g2307) & (!g2308) & (g2366) & (!g2398)) + ((g358) & (!g390) & (!g2307) & (g2308) & (!g2366) & (!g2398)) + ((g358) & (!g390) & (g2307) & (!g2308) & (!g2366) & (g2398)) + ((g358) & (!g390) & (g2307) & (!g2308) & (g2366) & (g2398)) + ((g358) & (!g390) & (g2307) & (g2308) & (!g2366) & (g2398)) + ((g358) & (!g390) & (g2307) & (g2308) & (g2366) & (!g2398)) + ((g358) & (!g390) & (g2307) & (g2308) & (g2366) & (g2398)) + ((g358) & (g390) & (!g2307) & (!g2308) & (!g2366) & (!g2398)) + ((g358) & (g390) & (g2307) & (!g2308) & (!g2366) & (g2398)) + ((g358) & (g390) & (g2307) & (!g2308) & (g2366) & (!g2398)) + ((g358) & (g390) & (g2307) & (!g2308) & (g2366) & (g2398)) + ((g358) & (g390) & (g2307) & (g2308) & (!g2366) & (!g2398)) + ((g358) & (g390) & (g2307) & (g2308) & (!g2366) & (g2398)) + ((g358) & (g390) & (g2307) & (g2308) & (g2366) & (!g2398)) + ((g358) & (g390) & (g2307) & (g2308) & (g2366) & (g2398)));
	assign g2407 = (((!g390) & (!g2308) & (g2366) & (!g2398)) + ((!g390) & (g2308) & (!g2366) & (!g2398)) + ((!g390) & (g2308) & (!g2366) & (g2398)) + ((!g390) & (g2308) & (g2366) & (g2398)) + ((g390) & (!g2308) & (!g2366) & (!g2398)) + ((g390) & (g2308) & (!g2366) & (g2398)) + ((g390) & (g2308) & (g2366) & (!g2398)) + ((g390) & (g2308) & (g2366) & (g2398)));
	assign g2408 = (((!g433) & (!g468) & (!g2310) & (g2311) & (g2365) & (!g2398)) + ((!g433) & (!g468) & (g2310) & (!g2311) & (!g2365) & (!g2398)) + ((!g433) & (!g468) & (g2310) & (!g2311) & (!g2365) & (g2398)) + ((!g433) & (!g468) & (g2310) & (!g2311) & (g2365) & (!g2398)) + ((!g433) & (!g468) & (g2310) & (!g2311) & (g2365) & (g2398)) + ((!g433) & (!g468) & (g2310) & (g2311) & (!g2365) & (!g2398)) + ((!g433) & (!g468) & (g2310) & (g2311) & (!g2365) & (g2398)) + ((!g433) & (!g468) & (g2310) & (g2311) & (g2365) & (g2398)) + ((!g433) & (g468) & (!g2310) & (!g2311) & (g2365) & (!g2398)) + ((!g433) & (g468) & (!g2310) & (g2311) & (!g2365) & (!g2398)) + ((!g433) & (g468) & (!g2310) & (g2311) & (g2365) & (!g2398)) + ((!g433) & (g468) & (g2310) & (!g2311) & (!g2365) & (!g2398)) + ((!g433) & (g468) & (g2310) & (!g2311) & (!g2365) & (g2398)) + ((!g433) & (g468) & (g2310) & (!g2311) & (g2365) & (g2398)) + ((!g433) & (g468) & (g2310) & (g2311) & (!g2365) & (g2398)) + ((!g433) & (g468) & (g2310) & (g2311) & (g2365) & (g2398)) + ((g433) & (!g468) & (!g2310) & (!g2311) & (!g2365) & (!g2398)) + ((g433) & (!g468) & (!g2310) & (!g2311) & (g2365) & (!g2398)) + ((g433) & (!g468) & (!g2310) & (g2311) & (!g2365) & (!g2398)) + ((g433) & (!g468) & (g2310) & (!g2311) & (!g2365) & (g2398)) + ((g433) & (!g468) & (g2310) & (!g2311) & (g2365) & (g2398)) + ((g433) & (!g468) & (g2310) & (g2311) & (!g2365) & (g2398)) + ((g433) & (!g468) & (g2310) & (g2311) & (g2365) & (!g2398)) + ((g433) & (!g468) & (g2310) & (g2311) & (g2365) & (g2398)) + ((g433) & (g468) & (!g2310) & (!g2311) & (!g2365) & (!g2398)) + ((g433) & (g468) & (g2310) & (!g2311) & (!g2365) & (g2398)) + ((g433) & (g468) & (g2310) & (!g2311) & (g2365) & (!g2398)) + ((g433) & (g468) & (g2310) & (!g2311) & (g2365) & (g2398)) + ((g433) & (g468) & (g2310) & (g2311) & (!g2365) & (!g2398)) + ((g433) & (g468) & (g2310) & (g2311) & (!g2365) & (g2398)) + ((g433) & (g468) & (g2310) & (g2311) & (g2365) & (!g2398)) + ((g433) & (g468) & (g2310) & (g2311) & (g2365) & (g2398)));
	assign g2409 = (((!g468) & (!g2311) & (g2365) & (!g2398)) + ((!g468) & (g2311) & (!g2365) & (!g2398)) + ((!g468) & (g2311) & (!g2365) & (g2398)) + ((!g468) & (g2311) & (g2365) & (g2398)) + ((g468) & (!g2311) & (!g2365) & (!g2398)) + ((g468) & (g2311) & (!g2365) & (g2398)) + ((g468) & (g2311) & (g2365) & (!g2398)) + ((g468) & (g2311) & (g2365) & (g2398)));
	assign g2410 = (((!g515) & (!g553) & (!g2313) & (g2314) & (g2364) & (!g2398)) + ((!g515) & (!g553) & (g2313) & (!g2314) & (!g2364) & (!g2398)) + ((!g515) & (!g553) & (g2313) & (!g2314) & (!g2364) & (g2398)) + ((!g515) & (!g553) & (g2313) & (!g2314) & (g2364) & (!g2398)) + ((!g515) & (!g553) & (g2313) & (!g2314) & (g2364) & (g2398)) + ((!g515) & (!g553) & (g2313) & (g2314) & (!g2364) & (!g2398)) + ((!g515) & (!g553) & (g2313) & (g2314) & (!g2364) & (g2398)) + ((!g515) & (!g553) & (g2313) & (g2314) & (g2364) & (g2398)) + ((!g515) & (g553) & (!g2313) & (!g2314) & (g2364) & (!g2398)) + ((!g515) & (g553) & (!g2313) & (g2314) & (!g2364) & (!g2398)) + ((!g515) & (g553) & (!g2313) & (g2314) & (g2364) & (!g2398)) + ((!g515) & (g553) & (g2313) & (!g2314) & (!g2364) & (!g2398)) + ((!g515) & (g553) & (g2313) & (!g2314) & (!g2364) & (g2398)) + ((!g515) & (g553) & (g2313) & (!g2314) & (g2364) & (g2398)) + ((!g515) & (g553) & (g2313) & (g2314) & (!g2364) & (g2398)) + ((!g515) & (g553) & (g2313) & (g2314) & (g2364) & (g2398)) + ((g515) & (!g553) & (!g2313) & (!g2314) & (!g2364) & (!g2398)) + ((g515) & (!g553) & (!g2313) & (!g2314) & (g2364) & (!g2398)) + ((g515) & (!g553) & (!g2313) & (g2314) & (!g2364) & (!g2398)) + ((g515) & (!g553) & (g2313) & (!g2314) & (!g2364) & (g2398)) + ((g515) & (!g553) & (g2313) & (!g2314) & (g2364) & (g2398)) + ((g515) & (!g553) & (g2313) & (g2314) & (!g2364) & (g2398)) + ((g515) & (!g553) & (g2313) & (g2314) & (g2364) & (!g2398)) + ((g515) & (!g553) & (g2313) & (g2314) & (g2364) & (g2398)) + ((g515) & (g553) & (!g2313) & (!g2314) & (!g2364) & (!g2398)) + ((g515) & (g553) & (g2313) & (!g2314) & (!g2364) & (g2398)) + ((g515) & (g553) & (g2313) & (!g2314) & (g2364) & (!g2398)) + ((g515) & (g553) & (g2313) & (!g2314) & (g2364) & (g2398)) + ((g515) & (g553) & (g2313) & (g2314) & (!g2364) & (!g2398)) + ((g515) & (g553) & (g2313) & (g2314) & (!g2364) & (g2398)) + ((g515) & (g553) & (g2313) & (g2314) & (g2364) & (!g2398)) + ((g515) & (g553) & (g2313) & (g2314) & (g2364) & (g2398)));
	assign g2411 = (((!g553) & (!g2314) & (g2364) & (!g2398)) + ((!g553) & (g2314) & (!g2364) & (!g2398)) + ((!g553) & (g2314) & (!g2364) & (g2398)) + ((!g553) & (g2314) & (g2364) & (g2398)) + ((g553) & (!g2314) & (!g2364) & (!g2398)) + ((g553) & (g2314) & (!g2364) & (g2398)) + ((g553) & (g2314) & (g2364) & (!g2398)) + ((g553) & (g2314) & (g2364) & (g2398)));
	assign g2412 = (((!g604) & (!g645) & (!g2316) & (g2317) & (g2363) & (!g2398)) + ((!g604) & (!g645) & (g2316) & (!g2317) & (!g2363) & (!g2398)) + ((!g604) & (!g645) & (g2316) & (!g2317) & (!g2363) & (g2398)) + ((!g604) & (!g645) & (g2316) & (!g2317) & (g2363) & (!g2398)) + ((!g604) & (!g645) & (g2316) & (!g2317) & (g2363) & (g2398)) + ((!g604) & (!g645) & (g2316) & (g2317) & (!g2363) & (!g2398)) + ((!g604) & (!g645) & (g2316) & (g2317) & (!g2363) & (g2398)) + ((!g604) & (!g645) & (g2316) & (g2317) & (g2363) & (g2398)) + ((!g604) & (g645) & (!g2316) & (!g2317) & (g2363) & (!g2398)) + ((!g604) & (g645) & (!g2316) & (g2317) & (!g2363) & (!g2398)) + ((!g604) & (g645) & (!g2316) & (g2317) & (g2363) & (!g2398)) + ((!g604) & (g645) & (g2316) & (!g2317) & (!g2363) & (!g2398)) + ((!g604) & (g645) & (g2316) & (!g2317) & (!g2363) & (g2398)) + ((!g604) & (g645) & (g2316) & (!g2317) & (g2363) & (g2398)) + ((!g604) & (g645) & (g2316) & (g2317) & (!g2363) & (g2398)) + ((!g604) & (g645) & (g2316) & (g2317) & (g2363) & (g2398)) + ((g604) & (!g645) & (!g2316) & (!g2317) & (!g2363) & (!g2398)) + ((g604) & (!g645) & (!g2316) & (!g2317) & (g2363) & (!g2398)) + ((g604) & (!g645) & (!g2316) & (g2317) & (!g2363) & (!g2398)) + ((g604) & (!g645) & (g2316) & (!g2317) & (!g2363) & (g2398)) + ((g604) & (!g645) & (g2316) & (!g2317) & (g2363) & (g2398)) + ((g604) & (!g645) & (g2316) & (g2317) & (!g2363) & (g2398)) + ((g604) & (!g645) & (g2316) & (g2317) & (g2363) & (!g2398)) + ((g604) & (!g645) & (g2316) & (g2317) & (g2363) & (g2398)) + ((g604) & (g645) & (!g2316) & (!g2317) & (!g2363) & (!g2398)) + ((g604) & (g645) & (g2316) & (!g2317) & (!g2363) & (g2398)) + ((g604) & (g645) & (g2316) & (!g2317) & (g2363) & (!g2398)) + ((g604) & (g645) & (g2316) & (!g2317) & (g2363) & (g2398)) + ((g604) & (g645) & (g2316) & (g2317) & (!g2363) & (!g2398)) + ((g604) & (g645) & (g2316) & (g2317) & (!g2363) & (g2398)) + ((g604) & (g645) & (g2316) & (g2317) & (g2363) & (!g2398)) + ((g604) & (g645) & (g2316) & (g2317) & (g2363) & (g2398)));
	assign g2413 = (((!g645) & (!g2317) & (g2363) & (!g2398)) + ((!g645) & (g2317) & (!g2363) & (!g2398)) + ((!g645) & (g2317) & (!g2363) & (g2398)) + ((!g645) & (g2317) & (g2363) & (g2398)) + ((g645) & (!g2317) & (!g2363) & (!g2398)) + ((g645) & (g2317) & (!g2363) & (g2398)) + ((g645) & (g2317) & (g2363) & (!g2398)) + ((g645) & (g2317) & (g2363) & (g2398)));
	assign g2414 = (((!g700) & (!g744) & (!g2319) & (g2320) & (g2362) & (!g2398)) + ((!g700) & (!g744) & (g2319) & (!g2320) & (!g2362) & (!g2398)) + ((!g700) & (!g744) & (g2319) & (!g2320) & (!g2362) & (g2398)) + ((!g700) & (!g744) & (g2319) & (!g2320) & (g2362) & (!g2398)) + ((!g700) & (!g744) & (g2319) & (!g2320) & (g2362) & (g2398)) + ((!g700) & (!g744) & (g2319) & (g2320) & (!g2362) & (!g2398)) + ((!g700) & (!g744) & (g2319) & (g2320) & (!g2362) & (g2398)) + ((!g700) & (!g744) & (g2319) & (g2320) & (g2362) & (g2398)) + ((!g700) & (g744) & (!g2319) & (!g2320) & (g2362) & (!g2398)) + ((!g700) & (g744) & (!g2319) & (g2320) & (!g2362) & (!g2398)) + ((!g700) & (g744) & (!g2319) & (g2320) & (g2362) & (!g2398)) + ((!g700) & (g744) & (g2319) & (!g2320) & (!g2362) & (!g2398)) + ((!g700) & (g744) & (g2319) & (!g2320) & (!g2362) & (g2398)) + ((!g700) & (g744) & (g2319) & (!g2320) & (g2362) & (g2398)) + ((!g700) & (g744) & (g2319) & (g2320) & (!g2362) & (g2398)) + ((!g700) & (g744) & (g2319) & (g2320) & (g2362) & (g2398)) + ((g700) & (!g744) & (!g2319) & (!g2320) & (!g2362) & (!g2398)) + ((g700) & (!g744) & (!g2319) & (!g2320) & (g2362) & (!g2398)) + ((g700) & (!g744) & (!g2319) & (g2320) & (!g2362) & (!g2398)) + ((g700) & (!g744) & (g2319) & (!g2320) & (!g2362) & (g2398)) + ((g700) & (!g744) & (g2319) & (!g2320) & (g2362) & (g2398)) + ((g700) & (!g744) & (g2319) & (g2320) & (!g2362) & (g2398)) + ((g700) & (!g744) & (g2319) & (g2320) & (g2362) & (!g2398)) + ((g700) & (!g744) & (g2319) & (g2320) & (g2362) & (g2398)) + ((g700) & (g744) & (!g2319) & (!g2320) & (!g2362) & (!g2398)) + ((g700) & (g744) & (g2319) & (!g2320) & (!g2362) & (g2398)) + ((g700) & (g744) & (g2319) & (!g2320) & (g2362) & (!g2398)) + ((g700) & (g744) & (g2319) & (!g2320) & (g2362) & (g2398)) + ((g700) & (g744) & (g2319) & (g2320) & (!g2362) & (!g2398)) + ((g700) & (g744) & (g2319) & (g2320) & (!g2362) & (g2398)) + ((g700) & (g744) & (g2319) & (g2320) & (g2362) & (!g2398)) + ((g700) & (g744) & (g2319) & (g2320) & (g2362) & (g2398)));
	assign g2415 = (((!g744) & (!g2320) & (g2362) & (!g2398)) + ((!g744) & (g2320) & (!g2362) & (!g2398)) + ((!g744) & (g2320) & (!g2362) & (g2398)) + ((!g744) & (g2320) & (g2362) & (g2398)) + ((g744) & (!g2320) & (!g2362) & (!g2398)) + ((g744) & (g2320) & (!g2362) & (g2398)) + ((g744) & (g2320) & (g2362) & (!g2398)) + ((g744) & (g2320) & (g2362) & (g2398)));
	assign g2416 = (((!g803) & (!g851) & (!g2322) & (g2323) & (g2361) & (!g2398)) + ((!g803) & (!g851) & (g2322) & (!g2323) & (!g2361) & (!g2398)) + ((!g803) & (!g851) & (g2322) & (!g2323) & (!g2361) & (g2398)) + ((!g803) & (!g851) & (g2322) & (!g2323) & (g2361) & (!g2398)) + ((!g803) & (!g851) & (g2322) & (!g2323) & (g2361) & (g2398)) + ((!g803) & (!g851) & (g2322) & (g2323) & (!g2361) & (!g2398)) + ((!g803) & (!g851) & (g2322) & (g2323) & (!g2361) & (g2398)) + ((!g803) & (!g851) & (g2322) & (g2323) & (g2361) & (g2398)) + ((!g803) & (g851) & (!g2322) & (!g2323) & (g2361) & (!g2398)) + ((!g803) & (g851) & (!g2322) & (g2323) & (!g2361) & (!g2398)) + ((!g803) & (g851) & (!g2322) & (g2323) & (g2361) & (!g2398)) + ((!g803) & (g851) & (g2322) & (!g2323) & (!g2361) & (!g2398)) + ((!g803) & (g851) & (g2322) & (!g2323) & (!g2361) & (g2398)) + ((!g803) & (g851) & (g2322) & (!g2323) & (g2361) & (g2398)) + ((!g803) & (g851) & (g2322) & (g2323) & (!g2361) & (g2398)) + ((!g803) & (g851) & (g2322) & (g2323) & (g2361) & (g2398)) + ((g803) & (!g851) & (!g2322) & (!g2323) & (!g2361) & (!g2398)) + ((g803) & (!g851) & (!g2322) & (!g2323) & (g2361) & (!g2398)) + ((g803) & (!g851) & (!g2322) & (g2323) & (!g2361) & (!g2398)) + ((g803) & (!g851) & (g2322) & (!g2323) & (!g2361) & (g2398)) + ((g803) & (!g851) & (g2322) & (!g2323) & (g2361) & (g2398)) + ((g803) & (!g851) & (g2322) & (g2323) & (!g2361) & (g2398)) + ((g803) & (!g851) & (g2322) & (g2323) & (g2361) & (!g2398)) + ((g803) & (!g851) & (g2322) & (g2323) & (g2361) & (g2398)) + ((g803) & (g851) & (!g2322) & (!g2323) & (!g2361) & (!g2398)) + ((g803) & (g851) & (g2322) & (!g2323) & (!g2361) & (g2398)) + ((g803) & (g851) & (g2322) & (!g2323) & (g2361) & (!g2398)) + ((g803) & (g851) & (g2322) & (!g2323) & (g2361) & (g2398)) + ((g803) & (g851) & (g2322) & (g2323) & (!g2361) & (!g2398)) + ((g803) & (g851) & (g2322) & (g2323) & (!g2361) & (g2398)) + ((g803) & (g851) & (g2322) & (g2323) & (g2361) & (!g2398)) + ((g803) & (g851) & (g2322) & (g2323) & (g2361) & (g2398)));
	assign g2417 = (((!g851) & (!g2323) & (g2361) & (!g2398)) + ((!g851) & (g2323) & (!g2361) & (!g2398)) + ((!g851) & (g2323) & (!g2361) & (g2398)) + ((!g851) & (g2323) & (g2361) & (g2398)) + ((g851) & (!g2323) & (!g2361) & (!g2398)) + ((g851) & (g2323) & (!g2361) & (g2398)) + ((g851) & (g2323) & (g2361) & (!g2398)) + ((g851) & (g2323) & (g2361) & (g2398)));
	assign g2418 = (((!g914) & (!g1032) & (!g2325) & (g2326) & (g2360) & (!g2398)) + ((!g914) & (!g1032) & (g2325) & (!g2326) & (!g2360) & (!g2398)) + ((!g914) & (!g1032) & (g2325) & (!g2326) & (!g2360) & (g2398)) + ((!g914) & (!g1032) & (g2325) & (!g2326) & (g2360) & (!g2398)) + ((!g914) & (!g1032) & (g2325) & (!g2326) & (g2360) & (g2398)) + ((!g914) & (!g1032) & (g2325) & (g2326) & (!g2360) & (!g2398)) + ((!g914) & (!g1032) & (g2325) & (g2326) & (!g2360) & (g2398)) + ((!g914) & (!g1032) & (g2325) & (g2326) & (g2360) & (g2398)) + ((!g914) & (g1032) & (!g2325) & (!g2326) & (g2360) & (!g2398)) + ((!g914) & (g1032) & (!g2325) & (g2326) & (!g2360) & (!g2398)) + ((!g914) & (g1032) & (!g2325) & (g2326) & (g2360) & (!g2398)) + ((!g914) & (g1032) & (g2325) & (!g2326) & (!g2360) & (!g2398)) + ((!g914) & (g1032) & (g2325) & (!g2326) & (!g2360) & (g2398)) + ((!g914) & (g1032) & (g2325) & (!g2326) & (g2360) & (g2398)) + ((!g914) & (g1032) & (g2325) & (g2326) & (!g2360) & (g2398)) + ((!g914) & (g1032) & (g2325) & (g2326) & (g2360) & (g2398)) + ((g914) & (!g1032) & (!g2325) & (!g2326) & (!g2360) & (!g2398)) + ((g914) & (!g1032) & (!g2325) & (!g2326) & (g2360) & (!g2398)) + ((g914) & (!g1032) & (!g2325) & (g2326) & (!g2360) & (!g2398)) + ((g914) & (!g1032) & (g2325) & (!g2326) & (!g2360) & (g2398)) + ((g914) & (!g1032) & (g2325) & (!g2326) & (g2360) & (g2398)) + ((g914) & (!g1032) & (g2325) & (g2326) & (!g2360) & (g2398)) + ((g914) & (!g1032) & (g2325) & (g2326) & (g2360) & (!g2398)) + ((g914) & (!g1032) & (g2325) & (g2326) & (g2360) & (g2398)) + ((g914) & (g1032) & (!g2325) & (!g2326) & (!g2360) & (!g2398)) + ((g914) & (g1032) & (g2325) & (!g2326) & (!g2360) & (g2398)) + ((g914) & (g1032) & (g2325) & (!g2326) & (g2360) & (!g2398)) + ((g914) & (g1032) & (g2325) & (!g2326) & (g2360) & (g2398)) + ((g914) & (g1032) & (g2325) & (g2326) & (!g2360) & (!g2398)) + ((g914) & (g1032) & (g2325) & (g2326) & (!g2360) & (g2398)) + ((g914) & (g1032) & (g2325) & (g2326) & (g2360) & (!g2398)) + ((g914) & (g1032) & (g2325) & (g2326) & (g2360) & (g2398)));
	assign g2419 = (((!g1032) & (!g2326) & (g2360) & (!g2398)) + ((!g1032) & (g2326) & (!g2360) & (!g2398)) + ((!g1032) & (g2326) & (!g2360) & (g2398)) + ((!g1032) & (g2326) & (g2360) & (g2398)) + ((g1032) & (!g2326) & (!g2360) & (!g2398)) + ((g1032) & (g2326) & (!g2360) & (g2398)) + ((g1032) & (g2326) & (g2360) & (!g2398)) + ((g1032) & (g2326) & (g2360) & (g2398)));
	assign g2420 = (((!g1030) & (!g1160) & (!g2328) & (g2329) & (g2359) & (!g2398)) + ((!g1030) & (!g1160) & (g2328) & (!g2329) & (!g2359) & (!g2398)) + ((!g1030) & (!g1160) & (g2328) & (!g2329) & (!g2359) & (g2398)) + ((!g1030) & (!g1160) & (g2328) & (!g2329) & (g2359) & (!g2398)) + ((!g1030) & (!g1160) & (g2328) & (!g2329) & (g2359) & (g2398)) + ((!g1030) & (!g1160) & (g2328) & (g2329) & (!g2359) & (!g2398)) + ((!g1030) & (!g1160) & (g2328) & (g2329) & (!g2359) & (g2398)) + ((!g1030) & (!g1160) & (g2328) & (g2329) & (g2359) & (g2398)) + ((!g1030) & (g1160) & (!g2328) & (!g2329) & (g2359) & (!g2398)) + ((!g1030) & (g1160) & (!g2328) & (g2329) & (!g2359) & (!g2398)) + ((!g1030) & (g1160) & (!g2328) & (g2329) & (g2359) & (!g2398)) + ((!g1030) & (g1160) & (g2328) & (!g2329) & (!g2359) & (!g2398)) + ((!g1030) & (g1160) & (g2328) & (!g2329) & (!g2359) & (g2398)) + ((!g1030) & (g1160) & (g2328) & (!g2329) & (g2359) & (g2398)) + ((!g1030) & (g1160) & (g2328) & (g2329) & (!g2359) & (g2398)) + ((!g1030) & (g1160) & (g2328) & (g2329) & (g2359) & (g2398)) + ((g1030) & (!g1160) & (!g2328) & (!g2329) & (!g2359) & (!g2398)) + ((g1030) & (!g1160) & (!g2328) & (!g2329) & (g2359) & (!g2398)) + ((g1030) & (!g1160) & (!g2328) & (g2329) & (!g2359) & (!g2398)) + ((g1030) & (!g1160) & (g2328) & (!g2329) & (!g2359) & (g2398)) + ((g1030) & (!g1160) & (g2328) & (!g2329) & (g2359) & (g2398)) + ((g1030) & (!g1160) & (g2328) & (g2329) & (!g2359) & (g2398)) + ((g1030) & (!g1160) & (g2328) & (g2329) & (g2359) & (!g2398)) + ((g1030) & (!g1160) & (g2328) & (g2329) & (g2359) & (g2398)) + ((g1030) & (g1160) & (!g2328) & (!g2329) & (!g2359) & (!g2398)) + ((g1030) & (g1160) & (g2328) & (!g2329) & (!g2359) & (g2398)) + ((g1030) & (g1160) & (g2328) & (!g2329) & (g2359) & (!g2398)) + ((g1030) & (g1160) & (g2328) & (!g2329) & (g2359) & (g2398)) + ((g1030) & (g1160) & (g2328) & (g2329) & (!g2359) & (!g2398)) + ((g1030) & (g1160) & (g2328) & (g2329) & (!g2359) & (g2398)) + ((g1030) & (g1160) & (g2328) & (g2329) & (g2359) & (!g2398)) + ((g1030) & (g1160) & (g2328) & (g2329) & (g2359) & (g2398)));
	assign g2421 = (((!g1160) & (!g2329) & (g2359) & (!g2398)) + ((!g1160) & (g2329) & (!g2359) & (!g2398)) + ((!g1160) & (g2329) & (!g2359) & (g2398)) + ((!g1160) & (g2329) & (g2359) & (g2398)) + ((g1160) & (!g2329) & (!g2359) & (!g2398)) + ((g1160) & (g2329) & (!g2359) & (g2398)) + ((g1160) & (g2329) & (g2359) & (!g2398)) + ((g1160) & (g2329) & (g2359) & (g2398)));
	assign g2422 = (((!g1154) & (!g1295) & (!g2331) & (g2332) & (g2358) & (!g2398)) + ((!g1154) & (!g1295) & (g2331) & (!g2332) & (!g2358) & (!g2398)) + ((!g1154) & (!g1295) & (g2331) & (!g2332) & (!g2358) & (g2398)) + ((!g1154) & (!g1295) & (g2331) & (!g2332) & (g2358) & (!g2398)) + ((!g1154) & (!g1295) & (g2331) & (!g2332) & (g2358) & (g2398)) + ((!g1154) & (!g1295) & (g2331) & (g2332) & (!g2358) & (!g2398)) + ((!g1154) & (!g1295) & (g2331) & (g2332) & (!g2358) & (g2398)) + ((!g1154) & (!g1295) & (g2331) & (g2332) & (g2358) & (g2398)) + ((!g1154) & (g1295) & (!g2331) & (!g2332) & (g2358) & (!g2398)) + ((!g1154) & (g1295) & (!g2331) & (g2332) & (!g2358) & (!g2398)) + ((!g1154) & (g1295) & (!g2331) & (g2332) & (g2358) & (!g2398)) + ((!g1154) & (g1295) & (g2331) & (!g2332) & (!g2358) & (!g2398)) + ((!g1154) & (g1295) & (g2331) & (!g2332) & (!g2358) & (g2398)) + ((!g1154) & (g1295) & (g2331) & (!g2332) & (g2358) & (g2398)) + ((!g1154) & (g1295) & (g2331) & (g2332) & (!g2358) & (g2398)) + ((!g1154) & (g1295) & (g2331) & (g2332) & (g2358) & (g2398)) + ((g1154) & (!g1295) & (!g2331) & (!g2332) & (!g2358) & (!g2398)) + ((g1154) & (!g1295) & (!g2331) & (!g2332) & (g2358) & (!g2398)) + ((g1154) & (!g1295) & (!g2331) & (g2332) & (!g2358) & (!g2398)) + ((g1154) & (!g1295) & (g2331) & (!g2332) & (!g2358) & (g2398)) + ((g1154) & (!g1295) & (g2331) & (!g2332) & (g2358) & (g2398)) + ((g1154) & (!g1295) & (g2331) & (g2332) & (!g2358) & (g2398)) + ((g1154) & (!g1295) & (g2331) & (g2332) & (g2358) & (!g2398)) + ((g1154) & (!g1295) & (g2331) & (g2332) & (g2358) & (g2398)) + ((g1154) & (g1295) & (!g2331) & (!g2332) & (!g2358) & (!g2398)) + ((g1154) & (g1295) & (g2331) & (!g2332) & (!g2358) & (g2398)) + ((g1154) & (g1295) & (g2331) & (!g2332) & (g2358) & (!g2398)) + ((g1154) & (g1295) & (g2331) & (!g2332) & (g2358) & (g2398)) + ((g1154) & (g1295) & (g2331) & (g2332) & (!g2358) & (!g2398)) + ((g1154) & (g1295) & (g2331) & (g2332) & (!g2358) & (g2398)) + ((g1154) & (g1295) & (g2331) & (g2332) & (g2358) & (!g2398)) + ((g1154) & (g1295) & (g2331) & (g2332) & (g2358) & (g2398)));
	assign g2423 = (((!g1295) & (!g2332) & (g2358) & (!g2398)) + ((!g1295) & (g2332) & (!g2358) & (!g2398)) + ((!g1295) & (g2332) & (!g2358) & (g2398)) + ((!g1295) & (g2332) & (g2358) & (g2398)) + ((g1295) & (!g2332) & (!g2358) & (!g2398)) + ((g1295) & (g2332) & (!g2358) & (g2398)) + ((g1295) & (g2332) & (g2358) & (!g2398)) + ((g1295) & (g2332) & (g2358) & (g2398)));
	assign g2424 = (((!g1285) & (!g1437) & (!g2334) & (g2335) & (g2357) & (!g2398)) + ((!g1285) & (!g1437) & (g2334) & (!g2335) & (!g2357) & (!g2398)) + ((!g1285) & (!g1437) & (g2334) & (!g2335) & (!g2357) & (g2398)) + ((!g1285) & (!g1437) & (g2334) & (!g2335) & (g2357) & (!g2398)) + ((!g1285) & (!g1437) & (g2334) & (!g2335) & (g2357) & (g2398)) + ((!g1285) & (!g1437) & (g2334) & (g2335) & (!g2357) & (!g2398)) + ((!g1285) & (!g1437) & (g2334) & (g2335) & (!g2357) & (g2398)) + ((!g1285) & (!g1437) & (g2334) & (g2335) & (g2357) & (g2398)) + ((!g1285) & (g1437) & (!g2334) & (!g2335) & (g2357) & (!g2398)) + ((!g1285) & (g1437) & (!g2334) & (g2335) & (!g2357) & (!g2398)) + ((!g1285) & (g1437) & (!g2334) & (g2335) & (g2357) & (!g2398)) + ((!g1285) & (g1437) & (g2334) & (!g2335) & (!g2357) & (!g2398)) + ((!g1285) & (g1437) & (g2334) & (!g2335) & (!g2357) & (g2398)) + ((!g1285) & (g1437) & (g2334) & (!g2335) & (g2357) & (g2398)) + ((!g1285) & (g1437) & (g2334) & (g2335) & (!g2357) & (g2398)) + ((!g1285) & (g1437) & (g2334) & (g2335) & (g2357) & (g2398)) + ((g1285) & (!g1437) & (!g2334) & (!g2335) & (!g2357) & (!g2398)) + ((g1285) & (!g1437) & (!g2334) & (!g2335) & (g2357) & (!g2398)) + ((g1285) & (!g1437) & (!g2334) & (g2335) & (!g2357) & (!g2398)) + ((g1285) & (!g1437) & (g2334) & (!g2335) & (!g2357) & (g2398)) + ((g1285) & (!g1437) & (g2334) & (!g2335) & (g2357) & (g2398)) + ((g1285) & (!g1437) & (g2334) & (g2335) & (!g2357) & (g2398)) + ((g1285) & (!g1437) & (g2334) & (g2335) & (g2357) & (!g2398)) + ((g1285) & (!g1437) & (g2334) & (g2335) & (g2357) & (g2398)) + ((g1285) & (g1437) & (!g2334) & (!g2335) & (!g2357) & (!g2398)) + ((g1285) & (g1437) & (g2334) & (!g2335) & (!g2357) & (g2398)) + ((g1285) & (g1437) & (g2334) & (!g2335) & (g2357) & (!g2398)) + ((g1285) & (g1437) & (g2334) & (!g2335) & (g2357) & (g2398)) + ((g1285) & (g1437) & (g2334) & (g2335) & (!g2357) & (!g2398)) + ((g1285) & (g1437) & (g2334) & (g2335) & (!g2357) & (g2398)) + ((g1285) & (g1437) & (g2334) & (g2335) & (g2357) & (!g2398)) + ((g1285) & (g1437) & (g2334) & (g2335) & (g2357) & (g2398)));
	assign g2425 = (((!g1437) & (!g2335) & (g2357) & (!g2398)) + ((!g1437) & (g2335) & (!g2357) & (!g2398)) + ((!g1437) & (g2335) & (!g2357) & (g2398)) + ((!g1437) & (g2335) & (g2357) & (g2398)) + ((g1437) & (!g2335) & (!g2357) & (!g2398)) + ((g1437) & (g2335) & (!g2357) & (g2398)) + ((g1437) & (g2335) & (g2357) & (!g2398)) + ((g1437) & (g2335) & (g2357) & (g2398)));
	assign g2426 = (((!g1423) & (!g1586) & (!g2337) & (g2338) & (g2356) & (!g2398)) + ((!g1423) & (!g1586) & (g2337) & (!g2338) & (!g2356) & (!g2398)) + ((!g1423) & (!g1586) & (g2337) & (!g2338) & (!g2356) & (g2398)) + ((!g1423) & (!g1586) & (g2337) & (!g2338) & (g2356) & (!g2398)) + ((!g1423) & (!g1586) & (g2337) & (!g2338) & (g2356) & (g2398)) + ((!g1423) & (!g1586) & (g2337) & (g2338) & (!g2356) & (!g2398)) + ((!g1423) & (!g1586) & (g2337) & (g2338) & (!g2356) & (g2398)) + ((!g1423) & (!g1586) & (g2337) & (g2338) & (g2356) & (g2398)) + ((!g1423) & (g1586) & (!g2337) & (!g2338) & (g2356) & (!g2398)) + ((!g1423) & (g1586) & (!g2337) & (g2338) & (!g2356) & (!g2398)) + ((!g1423) & (g1586) & (!g2337) & (g2338) & (g2356) & (!g2398)) + ((!g1423) & (g1586) & (g2337) & (!g2338) & (!g2356) & (!g2398)) + ((!g1423) & (g1586) & (g2337) & (!g2338) & (!g2356) & (g2398)) + ((!g1423) & (g1586) & (g2337) & (!g2338) & (g2356) & (g2398)) + ((!g1423) & (g1586) & (g2337) & (g2338) & (!g2356) & (g2398)) + ((!g1423) & (g1586) & (g2337) & (g2338) & (g2356) & (g2398)) + ((g1423) & (!g1586) & (!g2337) & (!g2338) & (!g2356) & (!g2398)) + ((g1423) & (!g1586) & (!g2337) & (!g2338) & (g2356) & (!g2398)) + ((g1423) & (!g1586) & (!g2337) & (g2338) & (!g2356) & (!g2398)) + ((g1423) & (!g1586) & (g2337) & (!g2338) & (!g2356) & (g2398)) + ((g1423) & (!g1586) & (g2337) & (!g2338) & (g2356) & (g2398)) + ((g1423) & (!g1586) & (g2337) & (g2338) & (!g2356) & (g2398)) + ((g1423) & (!g1586) & (g2337) & (g2338) & (g2356) & (!g2398)) + ((g1423) & (!g1586) & (g2337) & (g2338) & (g2356) & (g2398)) + ((g1423) & (g1586) & (!g2337) & (!g2338) & (!g2356) & (!g2398)) + ((g1423) & (g1586) & (g2337) & (!g2338) & (!g2356) & (g2398)) + ((g1423) & (g1586) & (g2337) & (!g2338) & (g2356) & (!g2398)) + ((g1423) & (g1586) & (g2337) & (!g2338) & (g2356) & (g2398)) + ((g1423) & (g1586) & (g2337) & (g2338) & (!g2356) & (!g2398)) + ((g1423) & (g1586) & (g2337) & (g2338) & (!g2356) & (g2398)) + ((g1423) & (g1586) & (g2337) & (g2338) & (g2356) & (!g2398)) + ((g1423) & (g1586) & (g2337) & (g2338) & (g2356) & (g2398)));
	assign g2427 = (((!g1586) & (!g2338) & (g2356) & (!g2398)) + ((!g1586) & (g2338) & (!g2356) & (!g2398)) + ((!g1586) & (g2338) & (!g2356) & (g2398)) + ((!g1586) & (g2338) & (g2356) & (g2398)) + ((g1586) & (!g2338) & (!g2356) & (!g2398)) + ((g1586) & (g2338) & (!g2356) & (g2398)) + ((g1586) & (g2338) & (g2356) & (!g2398)) + ((g1586) & (g2338) & (g2356) & (g2398)));
	assign g2428 = (((!g1568) & (!g1742) & (!g2340) & (g2341) & (g2355) & (!g2398)) + ((!g1568) & (!g1742) & (g2340) & (!g2341) & (!g2355) & (!g2398)) + ((!g1568) & (!g1742) & (g2340) & (!g2341) & (!g2355) & (g2398)) + ((!g1568) & (!g1742) & (g2340) & (!g2341) & (g2355) & (!g2398)) + ((!g1568) & (!g1742) & (g2340) & (!g2341) & (g2355) & (g2398)) + ((!g1568) & (!g1742) & (g2340) & (g2341) & (!g2355) & (!g2398)) + ((!g1568) & (!g1742) & (g2340) & (g2341) & (!g2355) & (g2398)) + ((!g1568) & (!g1742) & (g2340) & (g2341) & (g2355) & (g2398)) + ((!g1568) & (g1742) & (!g2340) & (!g2341) & (g2355) & (!g2398)) + ((!g1568) & (g1742) & (!g2340) & (g2341) & (!g2355) & (!g2398)) + ((!g1568) & (g1742) & (!g2340) & (g2341) & (g2355) & (!g2398)) + ((!g1568) & (g1742) & (g2340) & (!g2341) & (!g2355) & (!g2398)) + ((!g1568) & (g1742) & (g2340) & (!g2341) & (!g2355) & (g2398)) + ((!g1568) & (g1742) & (g2340) & (!g2341) & (g2355) & (g2398)) + ((!g1568) & (g1742) & (g2340) & (g2341) & (!g2355) & (g2398)) + ((!g1568) & (g1742) & (g2340) & (g2341) & (g2355) & (g2398)) + ((g1568) & (!g1742) & (!g2340) & (!g2341) & (!g2355) & (!g2398)) + ((g1568) & (!g1742) & (!g2340) & (!g2341) & (g2355) & (!g2398)) + ((g1568) & (!g1742) & (!g2340) & (g2341) & (!g2355) & (!g2398)) + ((g1568) & (!g1742) & (g2340) & (!g2341) & (!g2355) & (g2398)) + ((g1568) & (!g1742) & (g2340) & (!g2341) & (g2355) & (g2398)) + ((g1568) & (!g1742) & (g2340) & (g2341) & (!g2355) & (g2398)) + ((g1568) & (!g1742) & (g2340) & (g2341) & (g2355) & (!g2398)) + ((g1568) & (!g1742) & (g2340) & (g2341) & (g2355) & (g2398)) + ((g1568) & (g1742) & (!g2340) & (!g2341) & (!g2355) & (!g2398)) + ((g1568) & (g1742) & (g2340) & (!g2341) & (!g2355) & (g2398)) + ((g1568) & (g1742) & (g2340) & (!g2341) & (g2355) & (!g2398)) + ((g1568) & (g1742) & (g2340) & (!g2341) & (g2355) & (g2398)) + ((g1568) & (g1742) & (g2340) & (g2341) & (!g2355) & (!g2398)) + ((g1568) & (g1742) & (g2340) & (g2341) & (!g2355) & (g2398)) + ((g1568) & (g1742) & (g2340) & (g2341) & (g2355) & (!g2398)) + ((g1568) & (g1742) & (g2340) & (g2341) & (g2355) & (g2398)));
	assign g2429 = (((!g1742) & (!g2341) & (g2355) & (!g2398)) + ((!g1742) & (g2341) & (!g2355) & (!g2398)) + ((!g1742) & (g2341) & (!g2355) & (g2398)) + ((!g1742) & (g2341) & (g2355) & (g2398)) + ((g1742) & (!g2341) & (!g2355) & (!g2398)) + ((g1742) & (g2341) & (!g2355) & (g2398)) + ((g1742) & (g2341) & (g2355) & (!g2398)) + ((g1742) & (g2341) & (g2355) & (g2398)));
	assign g2430 = (((!g1720) & (!g1905) & (!g2343) & (g2344) & (g2354) & (!g2398)) + ((!g1720) & (!g1905) & (g2343) & (!g2344) & (!g2354) & (!g2398)) + ((!g1720) & (!g1905) & (g2343) & (!g2344) & (!g2354) & (g2398)) + ((!g1720) & (!g1905) & (g2343) & (!g2344) & (g2354) & (!g2398)) + ((!g1720) & (!g1905) & (g2343) & (!g2344) & (g2354) & (g2398)) + ((!g1720) & (!g1905) & (g2343) & (g2344) & (!g2354) & (!g2398)) + ((!g1720) & (!g1905) & (g2343) & (g2344) & (!g2354) & (g2398)) + ((!g1720) & (!g1905) & (g2343) & (g2344) & (g2354) & (g2398)) + ((!g1720) & (g1905) & (!g2343) & (!g2344) & (g2354) & (!g2398)) + ((!g1720) & (g1905) & (!g2343) & (g2344) & (!g2354) & (!g2398)) + ((!g1720) & (g1905) & (!g2343) & (g2344) & (g2354) & (!g2398)) + ((!g1720) & (g1905) & (g2343) & (!g2344) & (!g2354) & (!g2398)) + ((!g1720) & (g1905) & (g2343) & (!g2344) & (!g2354) & (g2398)) + ((!g1720) & (g1905) & (g2343) & (!g2344) & (g2354) & (g2398)) + ((!g1720) & (g1905) & (g2343) & (g2344) & (!g2354) & (g2398)) + ((!g1720) & (g1905) & (g2343) & (g2344) & (g2354) & (g2398)) + ((g1720) & (!g1905) & (!g2343) & (!g2344) & (!g2354) & (!g2398)) + ((g1720) & (!g1905) & (!g2343) & (!g2344) & (g2354) & (!g2398)) + ((g1720) & (!g1905) & (!g2343) & (g2344) & (!g2354) & (!g2398)) + ((g1720) & (!g1905) & (g2343) & (!g2344) & (!g2354) & (g2398)) + ((g1720) & (!g1905) & (g2343) & (!g2344) & (g2354) & (g2398)) + ((g1720) & (!g1905) & (g2343) & (g2344) & (!g2354) & (g2398)) + ((g1720) & (!g1905) & (g2343) & (g2344) & (g2354) & (!g2398)) + ((g1720) & (!g1905) & (g2343) & (g2344) & (g2354) & (g2398)) + ((g1720) & (g1905) & (!g2343) & (!g2344) & (!g2354) & (!g2398)) + ((g1720) & (g1905) & (g2343) & (!g2344) & (!g2354) & (g2398)) + ((g1720) & (g1905) & (g2343) & (!g2344) & (g2354) & (!g2398)) + ((g1720) & (g1905) & (g2343) & (!g2344) & (g2354) & (g2398)) + ((g1720) & (g1905) & (g2343) & (g2344) & (!g2354) & (!g2398)) + ((g1720) & (g1905) & (g2343) & (g2344) & (!g2354) & (g2398)) + ((g1720) & (g1905) & (g2343) & (g2344) & (g2354) & (!g2398)) + ((g1720) & (g1905) & (g2343) & (g2344) & (g2354) & (g2398)));
	assign g2431 = (((!g1905) & (!g2344) & (g2354) & (!g2398)) + ((!g1905) & (g2344) & (!g2354) & (!g2398)) + ((!g1905) & (g2344) & (!g2354) & (g2398)) + ((!g1905) & (g2344) & (g2354) & (g2398)) + ((g1905) & (!g2344) & (!g2354) & (!g2398)) + ((g1905) & (g2344) & (!g2354) & (g2398)) + ((g1905) & (g2344) & (g2354) & (!g2398)) + ((g1905) & (g2344) & (g2354) & (g2398)));
	assign g2432 = (((!g1879) & (!g2075) & (!g2346) & (g2347) & (g2353) & (!g2398)) + ((!g1879) & (!g2075) & (g2346) & (!g2347) & (!g2353) & (!g2398)) + ((!g1879) & (!g2075) & (g2346) & (!g2347) & (!g2353) & (g2398)) + ((!g1879) & (!g2075) & (g2346) & (!g2347) & (g2353) & (!g2398)) + ((!g1879) & (!g2075) & (g2346) & (!g2347) & (g2353) & (g2398)) + ((!g1879) & (!g2075) & (g2346) & (g2347) & (!g2353) & (!g2398)) + ((!g1879) & (!g2075) & (g2346) & (g2347) & (!g2353) & (g2398)) + ((!g1879) & (!g2075) & (g2346) & (g2347) & (g2353) & (g2398)) + ((!g1879) & (g2075) & (!g2346) & (!g2347) & (g2353) & (!g2398)) + ((!g1879) & (g2075) & (!g2346) & (g2347) & (!g2353) & (!g2398)) + ((!g1879) & (g2075) & (!g2346) & (g2347) & (g2353) & (!g2398)) + ((!g1879) & (g2075) & (g2346) & (!g2347) & (!g2353) & (!g2398)) + ((!g1879) & (g2075) & (g2346) & (!g2347) & (!g2353) & (g2398)) + ((!g1879) & (g2075) & (g2346) & (!g2347) & (g2353) & (g2398)) + ((!g1879) & (g2075) & (g2346) & (g2347) & (!g2353) & (g2398)) + ((!g1879) & (g2075) & (g2346) & (g2347) & (g2353) & (g2398)) + ((g1879) & (!g2075) & (!g2346) & (!g2347) & (!g2353) & (!g2398)) + ((g1879) & (!g2075) & (!g2346) & (!g2347) & (g2353) & (!g2398)) + ((g1879) & (!g2075) & (!g2346) & (g2347) & (!g2353) & (!g2398)) + ((g1879) & (!g2075) & (g2346) & (!g2347) & (!g2353) & (g2398)) + ((g1879) & (!g2075) & (g2346) & (!g2347) & (g2353) & (g2398)) + ((g1879) & (!g2075) & (g2346) & (g2347) & (!g2353) & (g2398)) + ((g1879) & (!g2075) & (g2346) & (g2347) & (g2353) & (!g2398)) + ((g1879) & (!g2075) & (g2346) & (g2347) & (g2353) & (g2398)) + ((g1879) & (g2075) & (!g2346) & (!g2347) & (!g2353) & (!g2398)) + ((g1879) & (g2075) & (g2346) & (!g2347) & (!g2353) & (g2398)) + ((g1879) & (g2075) & (g2346) & (!g2347) & (g2353) & (!g2398)) + ((g1879) & (g2075) & (g2346) & (!g2347) & (g2353) & (g2398)) + ((g1879) & (g2075) & (g2346) & (g2347) & (!g2353) & (!g2398)) + ((g1879) & (g2075) & (g2346) & (g2347) & (!g2353) & (g2398)) + ((g1879) & (g2075) & (g2346) & (g2347) & (g2353) & (!g2398)) + ((g1879) & (g2075) & (g2346) & (g2347) & (g2353) & (g2398)));
	assign g2433 = (((!g2075) & (!g2347) & (g2353) & (!g2398)) + ((!g2075) & (g2347) & (!g2353) & (!g2398)) + ((!g2075) & (g2347) & (!g2353) & (g2398)) + ((!g2075) & (g2347) & (g2353) & (g2398)) + ((g2075) & (!g2347) & (!g2353) & (!g2398)) + ((g2075) & (g2347) & (!g2353) & (g2398)) + ((g2075) & (g2347) & (g2353) & (!g2398)) + ((g2075) & (g2347) & (g2353) & (g2398)));
	assign g2434 = (((!g2045) & (!g2252) & (!g2349) & (g2350) & (g2352) & (!g2398)) + ((!g2045) & (!g2252) & (g2349) & (!g2350) & (!g2352) & (!g2398)) + ((!g2045) & (!g2252) & (g2349) & (!g2350) & (!g2352) & (g2398)) + ((!g2045) & (!g2252) & (g2349) & (!g2350) & (g2352) & (!g2398)) + ((!g2045) & (!g2252) & (g2349) & (!g2350) & (g2352) & (g2398)) + ((!g2045) & (!g2252) & (g2349) & (g2350) & (!g2352) & (!g2398)) + ((!g2045) & (!g2252) & (g2349) & (g2350) & (!g2352) & (g2398)) + ((!g2045) & (!g2252) & (g2349) & (g2350) & (g2352) & (g2398)) + ((!g2045) & (g2252) & (!g2349) & (!g2350) & (g2352) & (!g2398)) + ((!g2045) & (g2252) & (!g2349) & (g2350) & (!g2352) & (!g2398)) + ((!g2045) & (g2252) & (!g2349) & (g2350) & (g2352) & (!g2398)) + ((!g2045) & (g2252) & (g2349) & (!g2350) & (!g2352) & (!g2398)) + ((!g2045) & (g2252) & (g2349) & (!g2350) & (!g2352) & (g2398)) + ((!g2045) & (g2252) & (g2349) & (!g2350) & (g2352) & (g2398)) + ((!g2045) & (g2252) & (g2349) & (g2350) & (!g2352) & (g2398)) + ((!g2045) & (g2252) & (g2349) & (g2350) & (g2352) & (g2398)) + ((g2045) & (!g2252) & (!g2349) & (!g2350) & (!g2352) & (!g2398)) + ((g2045) & (!g2252) & (!g2349) & (!g2350) & (g2352) & (!g2398)) + ((g2045) & (!g2252) & (!g2349) & (g2350) & (!g2352) & (!g2398)) + ((g2045) & (!g2252) & (g2349) & (!g2350) & (!g2352) & (g2398)) + ((g2045) & (!g2252) & (g2349) & (!g2350) & (g2352) & (g2398)) + ((g2045) & (!g2252) & (g2349) & (g2350) & (!g2352) & (g2398)) + ((g2045) & (!g2252) & (g2349) & (g2350) & (g2352) & (!g2398)) + ((g2045) & (!g2252) & (g2349) & (g2350) & (g2352) & (g2398)) + ((g2045) & (g2252) & (!g2349) & (!g2350) & (!g2352) & (!g2398)) + ((g2045) & (g2252) & (g2349) & (!g2350) & (!g2352) & (g2398)) + ((g2045) & (g2252) & (g2349) & (!g2350) & (g2352) & (!g2398)) + ((g2045) & (g2252) & (g2349) & (!g2350) & (g2352) & (g2398)) + ((g2045) & (g2252) & (g2349) & (g2350) & (!g2352) & (!g2398)) + ((g2045) & (g2252) & (g2349) & (g2350) & (!g2352) & (g2398)) + ((g2045) & (g2252) & (g2349) & (g2350) & (g2352) & (!g2398)) + ((g2045) & (g2252) & (g2349) & (g2350) & (g2352) & (g2398)));
	assign g2435 = (((!g2252) & (!g2350) & (g2352) & (!g2398)) + ((!g2252) & (g2350) & (!g2352) & (!g2398)) + ((!g2252) & (g2350) & (!g2352) & (g2398)) + ((!g2252) & (g2350) & (g2352) & (g2398)) + ((g2252) & (!g2350) & (!g2352) & (!g2398)) + ((g2252) & (g2350) & (!g2352) & (g2398)) + ((g2252) & (g2350) & (g2352) & (!g2398)) + ((g2252) & (g2350) & (g2352) & (g2398)));
	assign g2436 = (((!g2274) & (g2295)));
	assign g2437 = (((!g2218) & (!ax26x) & (!ax27x) & (!g2436) & (!g2351) & (g2398)) + ((!g2218) & (!ax26x) & (!ax27x) & (!g2436) & (g2351) & (!g2398)) + ((!g2218) & (!ax26x) & (!ax27x) & (!g2436) & (g2351) & (g2398)) + ((!g2218) & (!ax26x) & (!ax27x) & (g2436) & (!g2351) & (!g2398)) + ((!g2218) & (!ax26x) & (ax27x) & (!g2436) & (!g2351) & (!g2398)) + ((!g2218) & (!ax26x) & (ax27x) & (g2436) & (!g2351) & (g2398)) + ((!g2218) & (!ax26x) & (ax27x) & (g2436) & (g2351) & (!g2398)) + ((!g2218) & (!ax26x) & (ax27x) & (g2436) & (g2351) & (g2398)) + ((!g2218) & (ax26x) & (!ax27x) & (g2436) & (!g2351) & (!g2398)) + ((!g2218) & (ax26x) & (!ax27x) & (g2436) & (g2351) & (!g2398)) + ((!g2218) & (ax26x) & (ax27x) & (!g2436) & (!g2351) & (!g2398)) + ((!g2218) & (ax26x) & (ax27x) & (!g2436) & (!g2351) & (g2398)) + ((!g2218) & (ax26x) & (ax27x) & (!g2436) & (g2351) & (!g2398)) + ((!g2218) & (ax26x) & (ax27x) & (!g2436) & (g2351) & (g2398)) + ((!g2218) & (ax26x) & (ax27x) & (g2436) & (!g2351) & (g2398)) + ((!g2218) & (ax26x) & (ax27x) & (g2436) & (g2351) & (g2398)) + ((g2218) & (!ax26x) & (!ax27x) & (!g2436) & (!g2351) & (!g2398)) + ((g2218) & (!ax26x) & (!ax27x) & (!g2436) & (!g2351) & (g2398)) + ((g2218) & (!ax26x) & (!ax27x) & (!g2436) & (g2351) & (g2398)) + ((g2218) & (!ax26x) & (!ax27x) & (g2436) & (g2351) & (!g2398)) + ((g2218) & (!ax26x) & (ax27x) & (!g2436) & (g2351) & (!g2398)) + ((g2218) & (!ax26x) & (ax27x) & (g2436) & (!g2351) & (!g2398)) + ((g2218) & (!ax26x) & (ax27x) & (g2436) & (!g2351) & (g2398)) + ((g2218) & (!ax26x) & (ax27x) & (g2436) & (g2351) & (g2398)) + ((g2218) & (ax26x) & (!ax27x) & (!g2436) & (!g2351) & (!g2398)) + ((g2218) & (ax26x) & (!ax27x) & (!g2436) & (g2351) & (!g2398)) + ((g2218) & (ax26x) & (ax27x) & (!g2436) & (!g2351) & (g2398)) + ((g2218) & (ax26x) & (ax27x) & (!g2436) & (g2351) & (g2398)) + ((g2218) & (ax26x) & (ax27x) & (g2436) & (!g2351) & (!g2398)) + ((g2218) & (ax26x) & (ax27x) & (g2436) & (!g2351) & (g2398)) + ((g2218) & (ax26x) & (ax27x) & (g2436) & (g2351) & (!g2398)) + ((g2218) & (ax26x) & (ax27x) & (g2436) & (g2351) & (g2398)));
	assign g2438 = (((!ax26x) & (!g2436) & (!g2351) & (g2398)) + ((!ax26x) & (!g2436) & (g2351) & (!g2398)) + ((!ax26x) & (!g2436) & (g2351) & (g2398)) + ((!ax26x) & (g2436) & (g2351) & (!g2398)) + ((ax26x) & (!g2436) & (!g2351) & (!g2398)) + ((ax26x) & (g2436) & (!g2351) & (!g2398)) + ((ax26x) & (g2436) & (!g2351) & (g2398)) + ((ax26x) & (g2436) & (g2351) & (g2398)));
	assign g2439 = (((!ax22x) & (!ax23x)));
	assign g2440 = (((!g2436) & (!ax24x) & (!ax25x) & (!g2398) & (!g2439)) + ((!g2436) & (!ax24x) & (ax25x) & (g2398) & (!g2439)) + ((!g2436) & (ax24x) & (ax25x) & (g2398) & (!g2439)) + ((!g2436) & (ax24x) & (ax25x) & (g2398) & (g2439)) + ((g2436) & (!ax24x) & (!ax25x) & (!g2398) & (!g2439)) + ((g2436) & (!ax24x) & (!ax25x) & (!g2398) & (g2439)) + ((g2436) & (!ax24x) & (!ax25x) & (g2398) & (!g2439)) + ((g2436) & (!ax24x) & (ax25x) & (!g2398) & (!g2439)) + ((g2436) & (!ax24x) & (ax25x) & (g2398) & (!g2439)) + ((g2436) & (!ax24x) & (ax25x) & (g2398) & (g2439)) + ((g2436) & (ax24x) & (!ax25x) & (g2398) & (!g2439)) + ((g2436) & (ax24x) & (!ax25x) & (g2398) & (g2439)) + ((g2436) & (ax24x) & (ax25x) & (!g2398) & (!g2439)) + ((g2436) & (ax24x) & (ax25x) & (!g2398) & (g2439)) + ((g2436) & (ax24x) & (ax25x) & (g2398) & (!g2439)) + ((g2436) & (ax24x) & (ax25x) & (g2398) & (g2439)));
	assign g2441 = (((!g2252) & (!g2218) & (g2437) & (g2438) & (g2440)) + ((!g2252) & (g2218) & (g2437) & (!g2438) & (g2440)) + ((!g2252) & (g2218) & (g2437) & (g2438) & (!g2440)) + ((!g2252) & (g2218) & (g2437) & (g2438) & (g2440)) + ((g2252) & (!g2218) & (!g2437) & (g2438) & (g2440)) + ((g2252) & (!g2218) & (g2437) & (!g2438) & (!g2440)) + ((g2252) & (!g2218) & (g2437) & (!g2438) & (g2440)) + ((g2252) & (!g2218) & (g2437) & (g2438) & (!g2440)) + ((g2252) & (!g2218) & (g2437) & (g2438) & (g2440)) + ((g2252) & (g2218) & (!g2437) & (!g2438) & (g2440)) + ((g2252) & (g2218) & (!g2437) & (g2438) & (!g2440)) + ((g2252) & (g2218) & (!g2437) & (g2438) & (g2440)) + ((g2252) & (g2218) & (g2437) & (!g2438) & (!g2440)) + ((g2252) & (g2218) & (g2437) & (!g2438) & (g2440)) + ((g2252) & (g2218) & (g2437) & (g2438) & (!g2440)) + ((g2252) & (g2218) & (g2437) & (g2438) & (g2440)));
	assign g2442 = (((!g2075) & (!g2045) & (g2434) & (g2435) & (g2441)) + ((!g2075) & (g2045) & (g2434) & (!g2435) & (g2441)) + ((!g2075) & (g2045) & (g2434) & (g2435) & (!g2441)) + ((!g2075) & (g2045) & (g2434) & (g2435) & (g2441)) + ((g2075) & (!g2045) & (!g2434) & (g2435) & (g2441)) + ((g2075) & (!g2045) & (g2434) & (!g2435) & (!g2441)) + ((g2075) & (!g2045) & (g2434) & (!g2435) & (g2441)) + ((g2075) & (!g2045) & (g2434) & (g2435) & (!g2441)) + ((g2075) & (!g2045) & (g2434) & (g2435) & (g2441)) + ((g2075) & (g2045) & (!g2434) & (!g2435) & (g2441)) + ((g2075) & (g2045) & (!g2434) & (g2435) & (!g2441)) + ((g2075) & (g2045) & (!g2434) & (g2435) & (g2441)) + ((g2075) & (g2045) & (g2434) & (!g2435) & (!g2441)) + ((g2075) & (g2045) & (g2434) & (!g2435) & (g2441)) + ((g2075) & (g2045) & (g2434) & (g2435) & (!g2441)) + ((g2075) & (g2045) & (g2434) & (g2435) & (g2441)));
	assign g2443 = (((!g1905) & (!g1879) & (g2432) & (g2433) & (g2442)) + ((!g1905) & (g1879) & (g2432) & (!g2433) & (g2442)) + ((!g1905) & (g1879) & (g2432) & (g2433) & (!g2442)) + ((!g1905) & (g1879) & (g2432) & (g2433) & (g2442)) + ((g1905) & (!g1879) & (!g2432) & (g2433) & (g2442)) + ((g1905) & (!g1879) & (g2432) & (!g2433) & (!g2442)) + ((g1905) & (!g1879) & (g2432) & (!g2433) & (g2442)) + ((g1905) & (!g1879) & (g2432) & (g2433) & (!g2442)) + ((g1905) & (!g1879) & (g2432) & (g2433) & (g2442)) + ((g1905) & (g1879) & (!g2432) & (!g2433) & (g2442)) + ((g1905) & (g1879) & (!g2432) & (g2433) & (!g2442)) + ((g1905) & (g1879) & (!g2432) & (g2433) & (g2442)) + ((g1905) & (g1879) & (g2432) & (!g2433) & (!g2442)) + ((g1905) & (g1879) & (g2432) & (!g2433) & (g2442)) + ((g1905) & (g1879) & (g2432) & (g2433) & (!g2442)) + ((g1905) & (g1879) & (g2432) & (g2433) & (g2442)));
	assign g2444 = (((!g1742) & (!g1720) & (g2430) & (g2431) & (g2443)) + ((!g1742) & (g1720) & (g2430) & (!g2431) & (g2443)) + ((!g1742) & (g1720) & (g2430) & (g2431) & (!g2443)) + ((!g1742) & (g1720) & (g2430) & (g2431) & (g2443)) + ((g1742) & (!g1720) & (!g2430) & (g2431) & (g2443)) + ((g1742) & (!g1720) & (g2430) & (!g2431) & (!g2443)) + ((g1742) & (!g1720) & (g2430) & (!g2431) & (g2443)) + ((g1742) & (!g1720) & (g2430) & (g2431) & (!g2443)) + ((g1742) & (!g1720) & (g2430) & (g2431) & (g2443)) + ((g1742) & (g1720) & (!g2430) & (!g2431) & (g2443)) + ((g1742) & (g1720) & (!g2430) & (g2431) & (!g2443)) + ((g1742) & (g1720) & (!g2430) & (g2431) & (g2443)) + ((g1742) & (g1720) & (g2430) & (!g2431) & (!g2443)) + ((g1742) & (g1720) & (g2430) & (!g2431) & (g2443)) + ((g1742) & (g1720) & (g2430) & (g2431) & (!g2443)) + ((g1742) & (g1720) & (g2430) & (g2431) & (g2443)));
	assign g2445 = (((!g1586) & (!g1568) & (g2428) & (g2429) & (g2444)) + ((!g1586) & (g1568) & (g2428) & (!g2429) & (g2444)) + ((!g1586) & (g1568) & (g2428) & (g2429) & (!g2444)) + ((!g1586) & (g1568) & (g2428) & (g2429) & (g2444)) + ((g1586) & (!g1568) & (!g2428) & (g2429) & (g2444)) + ((g1586) & (!g1568) & (g2428) & (!g2429) & (!g2444)) + ((g1586) & (!g1568) & (g2428) & (!g2429) & (g2444)) + ((g1586) & (!g1568) & (g2428) & (g2429) & (!g2444)) + ((g1586) & (!g1568) & (g2428) & (g2429) & (g2444)) + ((g1586) & (g1568) & (!g2428) & (!g2429) & (g2444)) + ((g1586) & (g1568) & (!g2428) & (g2429) & (!g2444)) + ((g1586) & (g1568) & (!g2428) & (g2429) & (g2444)) + ((g1586) & (g1568) & (g2428) & (!g2429) & (!g2444)) + ((g1586) & (g1568) & (g2428) & (!g2429) & (g2444)) + ((g1586) & (g1568) & (g2428) & (g2429) & (!g2444)) + ((g1586) & (g1568) & (g2428) & (g2429) & (g2444)));
	assign g2446 = (((!g1437) & (!g1423) & (g2426) & (g2427) & (g2445)) + ((!g1437) & (g1423) & (g2426) & (!g2427) & (g2445)) + ((!g1437) & (g1423) & (g2426) & (g2427) & (!g2445)) + ((!g1437) & (g1423) & (g2426) & (g2427) & (g2445)) + ((g1437) & (!g1423) & (!g2426) & (g2427) & (g2445)) + ((g1437) & (!g1423) & (g2426) & (!g2427) & (!g2445)) + ((g1437) & (!g1423) & (g2426) & (!g2427) & (g2445)) + ((g1437) & (!g1423) & (g2426) & (g2427) & (!g2445)) + ((g1437) & (!g1423) & (g2426) & (g2427) & (g2445)) + ((g1437) & (g1423) & (!g2426) & (!g2427) & (g2445)) + ((g1437) & (g1423) & (!g2426) & (g2427) & (!g2445)) + ((g1437) & (g1423) & (!g2426) & (g2427) & (g2445)) + ((g1437) & (g1423) & (g2426) & (!g2427) & (!g2445)) + ((g1437) & (g1423) & (g2426) & (!g2427) & (g2445)) + ((g1437) & (g1423) & (g2426) & (g2427) & (!g2445)) + ((g1437) & (g1423) & (g2426) & (g2427) & (g2445)));
	assign g2447 = (((!g1295) & (!g1285) & (g2424) & (g2425) & (g2446)) + ((!g1295) & (g1285) & (g2424) & (!g2425) & (g2446)) + ((!g1295) & (g1285) & (g2424) & (g2425) & (!g2446)) + ((!g1295) & (g1285) & (g2424) & (g2425) & (g2446)) + ((g1295) & (!g1285) & (!g2424) & (g2425) & (g2446)) + ((g1295) & (!g1285) & (g2424) & (!g2425) & (!g2446)) + ((g1295) & (!g1285) & (g2424) & (!g2425) & (g2446)) + ((g1295) & (!g1285) & (g2424) & (g2425) & (!g2446)) + ((g1295) & (!g1285) & (g2424) & (g2425) & (g2446)) + ((g1295) & (g1285) & (!g2424) & (!g2425) & (g2446)) + ((g1295) & (g1285) & (!g2424) & (g2425) & (!g2446)) + ((g1295) & (g1285) & (!g2424) & (g2425) & (g2446)) + ((g1295) & (g1285) & (g2424) & (!g2425) & (!g2446)) + ((g1295) & (g1285) & (g2424) & (!g2425) & (g2446)) + ((g1295) & (g1285) & (g2424) & (g2425) & (!g2446)) + ((g1295) & (g1285) & (g2424) & (g2425) & (g2446)));
	assign g2448 = (((!g1160) & (!g1154) & (g2422) & (g2423) & (g2447)) + ((!g1160) & (g1154) & (g2422) & (!g2423) & (g2447)) + ((!g1160) & (g1154) & (g2422) & (g2423) & (!g2447)) + ((!g1160) & (g1154) & (g2422) & (g2423) & (g2447)) + ((g1160) & (!g1154) & (!g2422) & (g2423) & (g2447)) + ((g1160) & (!g1154) & (g2422) & (!g2423) & (!g2447)) + ((g1160) & (!g1154) & (g2422) & (!g2423) & (g2447)) + ((g1160) & (!g1154) & (g2422) & (g2423) & (!g2447)) + ((g1160) & (!g1154) & (g2422) & (g2423) & (g2447)) + ((g1160) & (g1154) & (!g2422) & (!g2423) & (g2447)) + ((g1160) & (g1154) & (!g2422) & (g2423) & (!g2447)) + ((g1160) & (g1154) & (!g2422) & (g2423) & (g2447)) + ((g1160) & (g1154) & (g2422) & (!g2423) & (!g2447)) + ((g1160) & (g1154) & (g2422) & (!g2423) & (g2447)) + ((g1160) & (g1154) & (g2422) & (g2423) & (!g2447)) + ((g1160) & (g1154) & (g2422) & (g2423) & (g2447)));
	assign g2449 = (((!g1032) & (!g1030) & (g2420) & (g2421) & (g2448)) + ((!g1032) & (g1030) & (g2420) & (!g2421) & (g2448)) + ((!g1032) & (g1030) & (g2420) & (g2421) & (!g2448)) + ((!g1032) & (g1030) & (g2420) & (g2421) & (g2448)) + ((g1032) & (!g1030) & (!g2420) & (g2421) & (g2448)) + ((g1032) & (!g1030) & (g2420) & (!g2421) & (!g2448)) + ((g1032) & (!g1030) & (g2420) & (!g2421) & (g2448)) + ((g1032) & (!g1030) & (g2420) & (g2421) & (!g2448)) + ((g1032) & (!g1030) & (g2420) & (g2421) & (g2448)) + ((g1032) & (g1030) & (!g2420) & (!g2421) & (g2448)) + ((g1032) & (g1030) & (!g2420) & (g2421) & (!g2448)) + ((g1032) & (g1030) & (!g2420) & (g2421) & (g2448)) + ((g1032) & (g1030) & (g2420) & (!g2421) & (!g2448)) + ((g1032) & (g1030) & (g2420) & (!g2421) & (g2448)) + ((g1032) & (g1030) & (g2420) & (g2421) & (!g2448)) + ((g1032) & (g1030) & (g2420) & (g2421) & (g2448)));
	assign g2450 = (((!g851) & (!g914) & (g2418) & (g2419) & (g2449)) + ((!g851) & (g914) & (g2418) & (!g2419) & (g2449)) + ((!g851) & (g914) & (g2418) & (g2419) & (!g2449)) + ((!g851) & (g914) & (g2418) & (g2419) & (g2449)) + ((g851) & (!g914) & (!g2418) & (g2419) & (g2449)) + ((g851) & (!g914) & (g2418) & (!g2419) & (!g2449)) + ((g851) & (!g914) & (g2418) & (!g2419) & (g2449)) + ((g851) & (!g914) & (g2418) & (g2419) & (!g2449)) + ((g851) & (!g914) & (g2418) & (g2419) & (g2449)) + ((g851) & (g914) & (!g2418) & (!g2419) & (g2449)) + ((g851) & (g914) & (!g2418) & (g2419) & (!g2449)) + ((g851) & (g914) & (!g2418) & (g2419) & (g2449)) + ((g851) & (g914) & (g2418) & (!g2419) & (!g2449)) + ((g851) & (g914) & (g2418) & (!g2419) & (g2449)) + ((g851) & (g914) & (g2418) & (g2419) & (!g2449)) + ((g851) & (g914) & (g2418) & (g2419) & (g2449)));
	assign g2451 = (((!g744) & (!g803) & (g2416) & (g2417) & (g2450)) + ((!g744) & (g803) & (g2416) & (!g2417) & (g2450)) + ((!g744) & (g803) & (g2416) & (g2417) & (!g2450)) + ((!g744) & (g803) & (g2416) & (g2417) & (g2450)) + ((g744) & (!g803) & (!g2416) & (g2417) & (g2450)) + ((g744) & (!g803) & (g2416) & (!g2417) & (!g2450)) + ((g744) & (!g803) & (g2416) & (!g2417) & (g2450)) + ((g744) & (!g803) & (g2416) & (g2417) & (!g2450)) + ((g744) & (!g803) & (g2416) & (g2417) & (g2450)) + ((g744) & (g803) & (!g2416) & (!g2417) & (g2450)) + ((g744) & (g803) & (!g2416) & (g2417) & (!g2450)) + ((g744) & (g803) & (!g2416) & (g2417) & (g2450)) + ((g744) & (g803) & (g2416) & (!g2417) & (!g2450)) + ((g744) & (g803) & (g2416) & (!g2417) & (g2450)) + ((g744) & (g803) & (g2416) & (g2417) & (!g2450)) + ((g744) & (g803) & (g2416) & (g2417) & (g2450)));
	assign g2452 = (((!g645) & (!g700) & (g2414) & (g2415) & (g2451)) + ((!g645) & (g700) & (g2414) & (!g2415) & (g2451)) + ((!g645) & (g700) & (g2414) & (g2415) & (!g2451)) + ((!g645) & (g700) & (g2414) & (g2415) & (g2451)) + ((g645) & (!g700) & (!g2414) & (g2415) & (g2451)) + ((g645) & (!g700) & (g2414) & (!g2415) & (!g2451)) + ((g645) & (!g700) & (g2414) & (!g2415) & (g2451)) + ((g645) & (!g700) & (g2414) & (g2415) & (!g2451)) + ((g645) & (!g700) & (g2414) & (g2415) & (g2451)) + ((g645) & (g700) & (!g2414) & (!g2415) & (g2451)) + ((g645) & (g700) & (!g2414) & (g2415) & (!g2451)) + ((g645) & (g700) & (!g2414) & (g2415) & (g2451)) + ((g645) & (g700) & (g2414) & (!g2415) & (!g2451)) + ((g645) & (g700) & (g2414) & (!g2415) & (g2451)) + ((g645) & (g700) & (g2414) & (g2415) & (!g2451)) + ((g645) & (g700) & (g2414) & (g2415) & (g2451)));
	assign g2453 = (((!g553) & (!g604) & (g2412) & (g2413) & (g2452)) + ((!g553) & (g604) & (g2412) & (!g2413) & (g2452)) + ((!g553) & (g604) & (g2412) & (g2413) & (!g2452)) + ((!g553) & (g604) & (g2412) & (g2413) & (g2452)) + ((g553) & (!g604) & (!g2412) & (g2413) & (g2452)) + ((g553) & (!g604) & (g2412) & (!g2413) & (!g2452)) + ((g553) & (!g604) & (g2412) & (!g2413) & (g2452)) + ((g553) & (!g604) & (g2412) & (g2413) & (!g2452)) + ((g553) & (!g604) & (g2412) & (g2413) & (g2452)) + ((g553) & (g604) & (!g2412) & (!g2413) & (g2452)) + ((g553) & (g604) & (!g2412) & (g2413) & (!g2452)) + ((g553) & (g604) & (!g2412) & (g2413) & (g2452)) + ((g553) & (g604) & (g2412) & (!g2413) & (!g2452)) + ((g553) & (g604) & (g2412) & (!g2413) & (g2452)) + ((g553) & (g604) & (g2412) & (g2413) & (!g2452)) + ((g553) & (g604) & (g2412) & (g2413) & (g2452)));
	assign g2454 = (((!g468) & (!g515) & (g2410) & (g2411) & (g2453)) + ((!g468) & (g515) & (g2410) & (!g2411) & (g2453)) + ((!g468) & (g515) & (g2410) & (g2411) & (!g2453)) + ((!g468) & (g515) & (g2410) & (g2411) & (g2453)) + ((g468) & (!g515) & (!g2410) & (g2411) & (g2453)) + ((g468) & (!g515) & (g2410) & (!g2411) & (!g2453)) + ((g468) & (!g515) & (g2410) & (!g2411) & (g2453)) + ((g468) & (!g515) & (g2410) & (g2411) & (!g2453)) + ((g468) & (!g515) & (g2410) & (g2411) & (g2453)) + ((g468) & (g515) & (!g2410) & (!g2411) & (g2453)) + ((g468) & (g515) & (!g2410) & (g2411) & (!g2453)) + ((g468) & (g515) & (!g2410) & (g2411) & (g2453)) + ((g468) & (g515) & (g2410) & (!g2411) & (!g2453)) + ((g468) & (g515) & (g2410) & (!g2411) & (g2453)) + ((g468) & (g515) & (g2410) & (g2411) & (!g2453)) + ((g468) & (g515) & (g2410) & (g2411) & (g2453)));
	assign g2455 = (((!g390) & (!g433) & (g2408) & (g2409) & (g2454)) + ((!g390) & (g433) & (g2408) & (!g2409) & (g2454)) + ((!g390) & (g433) & (g2408) & (g2409) & (!g2454)) + ((!g390) & (g433) & (g2408) & (g2409) & (g2454)) + ((g390) & (!g433) & (!g2408) & (g2409) & (g2454)) + ((g390) & (!g433) & (g2408) & (!g2409) & (!g2454)) + ((g390) & (!g433) & (g2408) & (!g2409) & (g2454)) + ((g390) & (!g433) & (g2408) & (g2409) & (!g2454)) + ((g390) & (!g433) & (g2408) & (g2409) & (g2454)) + ((g390) & (g433) & (!g2408) & (!g2409) & (g2454)) + ((g390) & (g433) & (!g2408) & (g2409) & (!g2454)) + ((g390) & (g433) & (!g2408) & (g2409) & (g2454)) + ((g390) & (g433) & (g2408) & (!g2409) & (!g2454)) + ((g390) & (g433) & (g2408) & (!g2409) & (g2454)) + ((g390) & (g433) & (g2408) & (g2409) & (!g2454)) + ((g390) & (g433) & (g2408) & (g2409) & (g2454)));
	assign g2456 = (((!g319) & (!g358) & (g2406) & (g2407) & (g2455)) + ((!g319) & (g358) & (g2406) & (!g2407) & (g2455)) + ((!g319) & (g358) & (g2406) & (g2407) & (!g2455)) + ((!g319) & (g358) & (g2406) & (g2407) & (g2455)) + ((g319) & (!g358) & (!g2406) & (g2407) & (g2455)) + ((g319) & (!g358) & (g2406) & (!g2407) & (!g2455)) + ((g319) & (!g358) & (g2406) & (!g2407) & (g2455)) + ((g319) & (!g358) & (g2406) & (g2407) & (!g2455)) + ((g319) & (!g358) & (g2406) & (g2407) & (g2455)) + ((g319) & (g358) & (!g2406) & (!g2407) & (g2455)) + ((g319) & (g358) & (!g2406) & (g2407) & (!g2455)) + ((g319) & (g358) & (!g2406) & (g2407) & (g2455)) + ((g319) & (g358) & (g2406) & (!g2407) & (!g2455)) + ((g319) & (g358) & (g2406) & (!g2407) & (g2455)) + ((g319) & (g358) & (g2406) & (g2407) & (!g2455)) + ((g319) & (g358) & (g2406) & (g2407) & (g2455)));
	assign g2457 = (((!g255) & (!g290) & (g2404) & (g2405) & (g2456)) + ((!g255) & (g290) & (g2404) & (!g2405) & (g2456)) + ((!g255) & (g290) & (g2404) & (g2405) & (!g2456)) + ((!g255) & (g290) & (g2404) & (g2405) & (g2456)) + ((g255) & (!g290) & (!g2404) & (g2405) & (g2456)) + ((g255) & (!g290) & (g2404) & (!g2405) & (!g2456)) + ((g255) & (!g290) & (g2404) & (!g2405) & (g2456)) + ((g255) & (!g290) & (g2404) & (g2405) & (!g2456)) + ((g255) & (!g290) & (g2404) & (g2405) & (g2456)) + ((g255) & (g290) & (!g2404) & (!g2405) & (g2456)) + ((g255) & (g290) & (!g2404) & (g2405) & (!g2456)) + ((g255) & (g290) & (!g2404) & (g2405) & (g2456)) + ((g255) & (g290) & (g2404) & (!g2405) & (!g2456)) + ((g255) & (g290) & (g2404) & (!g2405) & (g2456)) + ((g255) & (g290) & (g2404) & (g2405) & (!g2456)) + ((g255) & (g290) & (g2404) & (g2405) & (g2456)));
	assign g2458 = (((!g198) & (!g229) & (g2402) & (g2403) & (g2457)) + ((!g198) & (g229) & (g2402) & (!g2403) & (g2457)) + ((!g198) & (g229) & (g2402) & (g2403) & (!g2457)) + ((!g198) & (g229) & (g2402) & (g2403) & (g2457)) + ((g198) & (!g229) & (!g2402) & (g2403) & (g2457)) + ((g198) & (!g229) & (g2402) & (!g2403) & (!g2457)) + ((g198) & (!g229) & (g2402) & (!g2403) & (g2457)) + ((g198) & (!g229) & (g2402) & (g2403) & (!g2457)) + ((g198) & (!g229) & (g2402) & (g2403) & (g2457)) + ((g198) & (g229) & (!g2402) & (!g2403) & (g2457)) + ((g198) & (g229) & (!g2402) & (g2403) & (!g2457)) + ((g198) & (g229) & (!g2402) & (g2403) & (g2457)) + ((g198) & (g229) & (g2402) & (!g2403) & (!g2457)) + ((g198) & (g229) & (g2402) & (!g2403) & (g2457)) + ((g198) & (g229) & (g2402) & (g2403) & (!g2457)) + ((g198) & (g229) & (g2402) & (g2403) & (g2457)));
	assign g2459 = (((!g147) & (!g174) & (g2400) & (g2401) & (g2458)) + ((!g147) & (g174) & (g2400) & (!g2401) & (g2458)) + ((!g147) & (g174) & (g2400) & (g2401) & (!g2458)) + ((!g147) & (g174) & (g2400) & (g2401) & (g2458)) + ((g147) & (!g174) & (!g2400) & (g2401) & (g2458)) + ((g147) & (!g174) & (g2400) & (!g2401) & (!g2458)) + ((g147) & (!g174) & (g2400) & (!g2401) & (g2458)) + ((g147) & (!g174) & (g2400) & (g2401) & (!g2458)) + ((g147) & (!g174) & (g2400) & (g2401) & (g2458)) + ((g147) & (g174) & (!g2400) & (!g2401) & (g2458)) + ((g147) & (g174) & (!g2400) & (g2401) & (!g2458)) + ((g147) & (g174) & (!g2400) & (g2401) & (g2458)) + ((g147) & (g174) & (g2400) & (!g2401) & (!g2458)) + ((g147) & (g174) & (g2400) & (!g2401) & (g2458)) + ((g147) & (g174) & (g2400) & (g2401) & (!g2458)) + ((g147) & (g174) & (g2400) & (g2401) & (g2458)));
	assign g2460 = (((g1) & (!g2371) & (g2394) & (g2397)) + ((g1) & (g2371) & (!g2394) & (!g2397)) + ((g1) & (g2371) & (!g2394) & (g2397)));
	assign g2461 = (((!g4) & (!g2) & (!g2372) & (!g2391) & (!g2393) & (!g2398)) + ((!g4) & (!g2) & (!g2372) & (!g2391) & (g2393) & (g2398)) + ((!g4) & (!g2) & (!g2372) & (g2391) & (!g2393) & (!g2398)) + ((!g4) & (!g2) & (!g2372) & (g2391) & (g2393) & (g2398)) + ((!g4) & (!g2) & (g2372) & (!g2391) & (!g2393) & (!g2398)) + ((!g4) & (!g2) & (g2372) & (!g2391) & (g2393) & (g2398)) + ((!g4) & (!g2) & (g2372) & (g2391) & (g2393) & (!g2398)) + ((!g4) & (!g2) & (g2372) & (g2391) & (g2393) & (g2398)) + ((!g4) & (g2) & (!g2372) & (!g2391) & (!g2393) & (!g2398)) + ((!g4) & (g2) & (!g2372) & (!g2391) & (g2393) & (g2398)) + ((!g4) & (g2) & (!g2372) & (g2391) & (g2393) & (!g2398)) + ((!g4) & (g2) & (!g2372) & (g2391) & (g2393) & (g2398)) + ((!g4) & (g2) & (g2372) & (!g2391) & (g2393) & (!g2398)) + ((!g4) & (g2) & (g2372) & (!g2391) & (g2393) & (g2398)) + ((!g4) & (g2) & (g2372) & (g2391) & (g2393) & (!g2398)) + ((!g4) & (g2) & (g2372) & (g2391) & (g2393) & (g2398)) + ((g4) & (!g2) & (!g2372) & (!g2391) & (g2393) & (!g2398)) + ((g4) & (!g2) & (!g2372) & (!g2391) & (g2393) & (g2398)) + ((g4) & (!g2) & (!g2372) & (g2391) & (g2393) & (!g2398)) + ((g4) & (!g2) & (!g2372) & (g2391) & (g2393) & (g2398)) + ((g4) & (!g2) & (g2372) & (!g2391) & (g2393) & (!g2398)) + ((g4) & (!g2) & (g2372) & (!g2391) & (g2393) & (g2398)) + ((g4) & (!g2) & (g2372) & (g2391) & (!g2393) & (!g2398)) + ((g4) & (!g2) & (g2372) & (g2391) & (g2393) & (g2398)) + ((g4) & (g2) & (!g2372) & (!g2391) & (g2393) & (!g2398)) + ((g4) & (g2) & (!g2372) & (!g2391) & (g2393) & (g2398)) + ((g4) & (g2) & (!g2372) & (g2391) & (!g2393) & (!g2398)) + ((g4) & (g2) & (!g2372) & (g2391) & (g2393) & (g2398)) + ((g4) & (g2) & (g2372) & (!g2391) & (!g2393) & (!g2398)) + ((g4) & (g2) & (g2372) & (!g2391) & (g2393) & (g2398)) + ((g4) & (g2) & (g2372) & (g2391) & (!g2393) & (!g2398)) + ((g4) & (g2) & (g2372) & (g2391) & (g2393) & (g2398)));
	assign g2462 = (((!g8) & (!g18) & (!g2374) & (g2375) & (g2390) & (!g2398)) + ((!g8) & (!g18) & (g2374) & (!g2375) & (!g2390) & (!g2398)) + ((!g8) & (!g18) & (g2374) & (!g2375) & (!g2390) & (g2398)) + ((!g8) & (!g18) & (g2374) & (!g2375) & (g2390) & (!g2398)) + ((!g8) & (!g18) & (g2374) & (!g2375) & (g2390) & (g2398)) + ((!g8) & (!g18) & (g2374) & (g2375) & (!g2390) & (!g2398)) + ((!g8) & (!g18) & (g2374) & (g2375) & (!g2390) & (g2398)) + ((!g8) & (!g18) & (g2374) & (g2375) & (g2390) & (g2398)) + ((!g8) & (g18) & (!g2374) & (!g2375) & (g2390) & (!g2398)) + ((!g8) & (g18) & (!g2374) & (g2375) & (!g2390) & (!g2398)) + ((!g8) & (g18) & (!g2374) & (g2375) & (g2390) & (!g2398)) + ((!g8) & (g18) & (g2374) & (!g2375) & (!g2390) & (!g2398)) + ((!g8) & (g18) & (g2374) & (!g2375) & (!g2390) & (g2398)) + ((!g8) & (g18) & (g2374) & (!g2375) & (g2390) & (g2398)) + ((!g8) & (g18) & (g2374) & (g2375) & (!g2390) & (g2398)) + ((!g8) & (g18) & (g2374) & (g2375) & (g2390) & (g2398)) + ((g8) & (!g18) & (!g2374) & (!g2375) & (!g2390) & (!g2398)) + ((g8) & (!g18) & (!g2374) & (!g2375) & (g2390) & (!g2398)) + ((g8) & (!g18) & (!g2374) & (g2375) & (!g2390) & (!g2398)) + ((g8) & (!g18) & (g2374) & (!g2375) & (!g2390) & (g2398)) + ((g8) & (!g18) & (g2374) & (!g2375) & (g2390) & (g2398)) + ((g8) & (!g18) & (g2374) & (g2375) & (!g2390) & (g2398)) + ((g8) & (!g18) & (g2374) & (g2375) & (g2390) & (!g2398)) + ((g8) & (!g18) & (g2374) & (g2375) & (g2390) & (g2398)) + ((g8) & (g18) & (!g2374) & (!g2375) & (!g2390) & (!g2398)) + ((g8) & (g18) & (g2374) & (!g2375) & (!g2390) & (g2398)) + ((g8) & (g18) & (g2374) & (!g2375) & (g2390) & (!g2398)) + ((g8) & (g18) & (g2374) & (!g2375) & (g2390) & (g2398)) + ((g8) & (g18) & (g2374) & (g2375) & (!g2390) & (!g2398)) + ((g8) & (g18) & (g2374) & (g2375) & (!g2390) & (g2398)) + ((g8) & (g18) & (g2374) & (g2375) & (g2390) & (!g2398)) + ((g8) & (g18) & (g2374) & (g2375) & (g2390) & (g2398)));
	assign g2463 = (((!g18) & (!g2375) & (g2390) & (!g2398)) + ((!g18) & (g2375) & (!g2390) & (!g2398)) + ((!g18) & (g2375) & (!g2390) & (g2398)) + ((!g18) & (g2375) & (g2390) & (g2398)) + ((g18) & (!g2375) & (!g2390) & (!g2398)) + ((g18) & (g2375) & (!g2390) & (g2398)) + ((g18) & (g2375) & (g2390) & (!g2398)) + ((g18) & (g2375) & (g2390) & (g2398)));
	assign g2464 = (((!g27) & (!g39) & (!g2377) & (g2378) & (g2389) & (!g2398)) + ((!g27) & (!g39) & (g2377) & (!g2378) & (!g2389) & (!g2398)) + ((!g27) & (!g39) & (g2377) & (!g2378) & (!g2389) & (g2398)) + ((!g27) & (!g39) & (g2377) & (!g2378) & (g2389) & (!g2398)) + ((!g27) & (!g39) & (g2377) & (!g2378) & (g2389) & (g2398)) + ((!g27) & (!g39) & (g2377) & (g2378) & (!g2389) & (!g2398)) + ((!g27) & (!g39) & (g2377) & (g2378) & (!g2389) & (g2398)) + ((!g27) & (!g39) & (g2377) & (g2378) & (g2389) & (g2398)) + ((!g27) & (g39) & (!g2377) & (!g2378) & (g2389) & (!g2398)) + ((!g27) & (g39) & (!g2377) & (g2378) & (!g2389) & (!g2398)) + ((!g27) & (g39) & (!g2377) & (g2378) & (g2389) & (!g2398)) + ((!g27) & (g39) & (g2377) & (!g2378) & (!g2389) & (!g2398)) + ((!g27) & (g39) & (g2377) & (!g2378) & (!g2389) & (g2398)) + ((!g27) & (g39) & (g2377) & (!g2378) & (g2389) & (g2398)) + ((!g27) & (g39) & (g2377) & (g2378) & (!g2389) & (g2398)) + ((!g27) & (g39) & (g2377) & (g2378) & (g2389) & (g2398)) + ((g27) & (!g39) & (!g2377) & (!g2378) & (!g2389) & (!g2398)) + ((g27) & (!g39) & (!g2377) & (!g2378) & (g2389) & (!g2398)) + ((g27) & (!g39) & (!g2377) & (g2378) & (!g2389) & (!g2398)) + ((g27) & (!g39) & (g2377) & (!g2378) & (!g2389) & (g2398)) + ((g27) & (!g39) & (g2377) & (!g2378) & (g2389) & (g2398)) + ((g27) & (!g39) & (g2377) & (g2378) & (!g2389) & (g2398)) + ((g27) & (!g39) & (g2377) & (g2378) & (g2389) & (!g2398)) + ((g27) & (!g39) & (g2377) & (g2378) & (g2389) & (g2398)) + ((g27) & (g39) & (!g2377) & (!g2378) & (!g2389) & (!g2398)) + ((g27) & (g39) & (g2377) & (!g2378) & (!g2389) & (g2398)) + ((g27) & (g39) & (g2377) & (!g2378) & (g2389) & (!g2398)) + ((g27) & (g39) & (g2377) & (!g2378) & (g2389) & (g2398)) + ((g27) & (g39) & (g2377) & (g2378) & (!g2389) & (!g2398)) + ((g27) & (g39) & (g2377) & (g2378) & (!g2389) & (g2398)) + ((g27) & (g39) & (g2377) & (g2378) & (g2389) & (!g2398)) + ((g27) & (g39) & (g2377) & (g2378) & (g2389) & (g2398)));
	assign g2465 = (((!g39) & (!g2378) & (g2389) & (!g2398)) + ((!g39) & (g2378) & (!g2389) & (!g2398)) + ((!g39) & (g2378) & (!g2389) & (g2398)) + ((!g39) & (g2378) & (g2389) & (g2398)) + ((g39) & (!g2378) & (!g2389) & (!g2398)) + ((g39) & (g2378) & (!g2389) & (g2398)) + ((g39) & (g2378) & (g2389) & (!g2398)) + ((g39) & (g2378) & (g2389) & (g2398)));
	assign g2466 = (((!g54) & (!g68) & (!g2380) & (g2381) & (g2388) & (!g2398)) + ((!g54) & (!g68) & (g2380) & (!g2381) & (!g2388) & (!g2398)) + ((!g54) & (!g68) & (g2380) & (!g2381) & (!g2388) & (g2398)) + ((!g54) & (!g68) & (g2380) & (!g2381) & (g2388) & (!g2398)) + ((!g54) & (!g68) & (g2380) & (!g2381) & (g2388) & (g2398)) + ((!g54) & (!g68) & (g2380) & (g2381) & (!g2388) & (!g2398)) + ((!g54) & (!g68) & (g2380) & (g2381) & (!g2388) & (g2398)) + ((!g54) & (!g68) & (g2380) & (g2381) & (g2388) & (g2398)) + ((!g54) & (g68) & (!g2380) & (!g2381) & (g2388) & (!g2398)) + ((!g54) & (g68) & (!g2380) & (g2381) & (!g2388) & (!g2398)) + ((!g54) & (g68) & (!g2380) & (g2381) & (g2388) & (!g2398)) + ((!g54) & (g68) & (g2380) & (!g2381) & (!g2388) & (!g2398)) + ((!g54) & (g68) & (g2380) & (!g2381) & (!g2388) & (g2398)) + ((!g54) & (g68) & (g2380) & (!g2381) & (g2388) & (g2398)) + ((!g54) & (g68) & (g2380) & (g2381) & (!g2388) & (g2398)) + ((!g54) & (g68) & (g2380) & (g2381) & (g2388) & (g2398)) + ((g54) & (!g68) & (!g2380) & (!g2381) & (!g2388) & (!g2398)) + ((g54) & (!g68) & (!g2380) & (!g2381) & (g2388) & (!g2398)) + ((g54) & (!g68) & (!g2380) & (g2381) & (!g2388) & (!g2398)) + ((g54) & (!g68) & (g2380) & (!g2381) & (!g2388) & (g2398)) + ((g54) & (!g68) & (g2380) & (!g2381) & (g2388) & (g2398)) + ((g54) & (!g68) & (g2380) & (g2381) & (!g2388) & (g2398)) + ((g54) & (!g68) & (g2380) & (g2381) & (g2388) & (!g2398)) + ((g54) & (!g68) & (g2380) & (g2381) & (g2388) & (g2398)) + ((g54) & (g68) & (!g2380) & (!g2381) & (!g2388) & (!g2398)) + ((g54) & (g68) & (g2380) & (!g2381) & (!g2388) & (g2398)) + ((g54) & (g68) & (g2380) & (!g2381) & (g2388) & (!g2398)) + ((g54) & (g68) & (g2380) & (!g2381) & (g2388) & (g2398)) + ((g54) & (g68) & (g2380) & (g2381) & (!g2388) & (!g2398)) + ((g54) & (g68) & (g2380) & (g2381) & (!g2388) & (g2398)) + ((g54) & (g68) & (g2380) & (g2381) & (g2388) & (!g2398)) + ((g54) & (g68) & (g2380) & (g2381) & (g2388) & (g2398)));
	assign g2467 = (((!g68) & (!g2381) & (g2388) & (!g2398)) + ((!g68) & (g2381) & (!g2388) & (!g2398)) + ((!g68) & (g2381) & (!g2388) & (g2398)) + ((!g68) & (g2381) & (g2388) & (g2398)) + ((g68) & (!g2381) & (!g2388) & (!g2398)) + ((g68) & (g2381) & (!g2388) & (g2398)) + ((g68) & (g2381) & (g2388) & (!g2398)) + ((g68) & (g2381) & (g2388) & (g2398)));
	assign g2468 = (((!g87) & (!g104) & (!g2383) & (g2384) & (g2387) & (!g2398)) + ((!g87) & (!g104) & (g2383) & (!g2384) & (!g2387) & (!g2398)) + ((!g87) & (!g104) & (g2383) & (!g2384) & (!g2387) & (g2398)) + ((!g87) & (!g104) & (g2383) & (!g2384) & (g2387) & (!g2398)) + ((!g87) & (!g104) & (g2383) & (!g2384) & (g2387) & (g2398)) + ((!g87) & (!g104) & (g2383) & (g2384) & (!g2387) & (!g2398)) + ((!g87) & (!g104) & (g2383) & (g2384) & (!g2387) & (g2398)) + ((!g87) & (!g104) & (g2383) & (g2384) & (g2387) & (g2398)) + ((!g87) & (g104) & (!g2383) & (!g2384) & (g2387) & (!g2398)) + ((!g87) & (g104) & (!g2383) & (g2384) & (!g2387) & (!g2398)) + ((!g87) & (g104) & (!g2383) & (g2384) & (g2387) & (!g2398)) + ((!g87) & (g104) & (g2383) & (!g2384) & (!g2387) & (!g2398)) + ((!g87) & (g104) & (g2383) & (!g2384) & (!g2387) & (g2398)) + ((!g87) & (g104) & (g2383) & (!g2384) & (g2387) & (g2398)) + ((!g87) & (g104) & (g2383) & (g2384) & (!g2387) & (g2398)) + ((!g87) & (g104) & (g2383) & (g2384) & (g2387) & (g2398)) + ((g87) & (!g104) & (!g2383) & (!g2384) & (!g2387) & (!g2398)) + ((g87) & (!g104) & (!g2383) & (!g2384) & (g2387) & (!g2398)) + ((g87) & (!g104) & (!g2383) & (g2384) & (!g2387) & (!g2398)) + ((g87) & (!g104) & (g2383) & (!g2384) & (!g2387) & (g2398)) + ((g87) & (!g104) & (g2383) & (!g2384) & (g2387) & (g2398)) + ((g87) & (!g104) & (g2383) & (g2384) & (!g2387) & (g2398)) + ((g87) & (!g104) & (g2383) & (g2384) & (g2387) & (!g2398)) + ((g87) & (!g104) & (g2383) & (g2384) & (g2387) & (g2398)) + ((g87) & (g104) & (!g2383) & (!g2384) & (!g2387) & (!g2398)) + ((g87) & (g104) & (g2383) & (!g2384) & (!g2387) & (g2398)) + ((g87) & (g104) & (g2383) & (!g2384) & (g2387) & (!g2398)) + ((g87) & (g104) & (g2383) & (!g2384) & (g2387) & (g2398)) + ((g87) & (g104) & (g2383) & (g2384) & (!g2387) & (!g2398)) + ((g87) & (g104) & (g2383) & (g2384) & (!g2387) & (g2398)) + ((g87) & (g104) & (g2383) & (g2384) & (g2387) & (!g2398)) + ((g87) & (g104) & (g2383) & (g2384) & (g2387) & (g2398)));
	assign g2469 = (((!g104) & (!g2384) & (g2387) & (!g2398)) + ((!g104) & (g2384) & (!g2387) & (!g2398)) + ((!g104) & (g2384) & (!g2387) & (g2398)) + ((!g104) & (g2384) & (g2387) & (g2398)) + ((g104) & (!g2384) & (!g2387) & (!g2398)) + ((g104) & (g2384) & (!g2387) & (g2398)) + ((g104) & (g2384) & (g2387) & (!g2398)) + ((g104) & (g2384) & (g2387) & (g2398)));
	assign g2470 = (((!g127) & (!g147) & (!g2386) & (g2296) & (g2370) & (!g2398)) + ((!g127) & (!g147) & (g2386) & (!g2296) & (!g2370) & (!g2398)) + ((!g127) & (!g147) & (g2386) & (!g2296) & (!g2370) & (g2398)) + ((!g127) & (!g147) & (g2386) & (!g2296) & (g2370) & (!g2398)) + ((!g127) & (!g147) & (g2386) & (!g2296) & (g2370) & (g2398)) + ((!g127) & (!g147) & (g2386) & (g2296) & (!g2370) & (!g2398)) + ((!g127) & (!g147) & (g2386) & (g2296) & (!g2370) & (g2398)) + ((!g127) & (!g147) & (g2386) & (g2296) & (g2370) & (g2398)) + ((!g127) & (g147) & (!g2386) & (!g2296) & (g2370) & (!g2398)) + ((!g127) & (g147) & (!g2386) & (g2296) & (!g2370) & (!g2398)) + ((!g127) & (g147) & (!g2386) & (g2296) & (g2370) & (!g2398)) + ((!g127) & (g147) & (g2386) & (!g2296) & (!g2370) & (!g2398)) + ((!g127) & (g147) & (g2386) & (!g2296) & (!g2370) & (g2398)) + ((!g127) & (g147) & (g2386) & (!g2296) & (g2370) & (g2398)) + ((!g127) & (g147) & (g2386) & (g2296) & (!g2370) & (g2398)) + ((!g127) & (g147) & (g2386) & (g2296) & (g2370) & (g2398)) + ((g127) & (!g147) & (!g2386) & (!g2296) & (!g2370) & (!g2398)) + ((g127) & (!g147) & (!g2386) & (!g2296) & (g2370) & (!g2398)) + ((g127) & (!g147) & (!g2386) & (g2296) & (!g2370) & (!g2398)) + ((g127) & (!g147) & (g2386) & (!g2296) & (!g2370) & (g2398)) + ((g127) & (!g147) & (g2386) & (!g2296) & (g2370) & (g2398)) + ((g127) & (!g147) & (g2386) & (g2296) & (!g2370) & (g2398)) + ((g127) & (!g147) & (g2386) & (g2296) & (g2370) & (!g2398)) + ((g127) & (!g147) & (g2386) & (g2296) & (g2370) & (g2398)) + ((g127) & (g147) & (!g2386) & (!g2296) & (!g2370) & (!g2398)) + ((g127) & (g147) & (g2386) & (!g2296) & (!g2370) & (g2398)) + ((g127) & (g147) & (g2386) & (!g2296) & (g2370) & (!g2398)) + ((g127) & (g147) & (g2386) & (!g2296) & (g2370) & (g2398)) + ((g127) & (g147) & (g2386) & (g2296) & (!g2370) & (!g2398)) + ((g127) & (g147) & (g2386) & (g2296) & (!g2370) & (g2398)) + ((g127) & (g147) & (g2386) & (g2296) & (g2370) & (!g2398)) + ((g127) & (g147) & (g2386) & (g2296) & (g2370) & (g2398)));
	assign g2471 = (((!g104) & (!g127) & (g2470) & (g2399) & (g2459)) + ((!g104) & (g127) & (g2470) & (!g2399) & (g2459)) + ((!g104) & (g127) & (g2470) & (g2399) & (!g2459)) + ((!g104) & (g127) & (g2470) & (g2399) & (g2459)) + ((g104) & (!g127) & (!g2470) & (g2399) & (g2459)) + ((g104) & (!g127) & (g2470) & (!g2399) & (!g2459)) + ((g104) & (!g127) & (g2470) & (!g2399) & (g2459)) + ((g104) & (!g127) & (g2470) & (g2399) & (!g2459)) + ((g104) & (!g127) & (g2470) & (g2399) & (g2459)) + ((g104) & (g127) & (!g2470) & (!g2399) & (g2459)) + ((g104) & (g127) & (!g2470) & (g2399) & (!g2459)) + ((g104) & (g127) & (!g2470) & (g2399) & (g2459)) + ((g104) & (g127) & (g2470) & (!g2399) & (!g2459)) + ((g104) & (g127) & (g2470) & (!g2399) & (g2459)) + ((g104) & (g127) & (g2470) & (g2399) & (!g2459)) + ((g104) & (g127) & (g2470) & (g2399) & (g2459)));
	assign g2472 = (((!g68) & (!g87) & (g2468) & (g2469) & (g2471)) + ((!g68) & (g87) & (g2468) & (!g2469) & (g2471)) + ((!g68) & (g87) & (g2468) & (g2469) & (!g2471)) + ((!g68) & (g87) & (g2468) & (g2469) & (g2471)) + ((g68) & (!g87) & (!g2468) & (g2469) & (g2471)) + ((g68) & (!g87) & (g2468) & (!g2469) & (!g2471)) + ((g68) & (!g87) & (g2468) & (!g2469) & (g2471)) + ((g68) & (!g87) & (g2468) & (g2469) & (!g2471)) + ((g68) & (!g87) & (g2468) & (g2469) & (g2471)) + ((g68) & (g87) & (!g2468) & (!g2469) & (g2471)) + ((g68) & (g87) & (!g2468) & (g2469) & (!g2471)) + ((g68) & (g87) & (!g2468) & (g2469) & (g2471)) + ((g68) & (g87) & (g2468) & (!g2469) & (!g2471)) + ((g68) & (g87) & (g2468) & (!g2469) & (g2471)) + ((g68) & (g87) & (g2468) & (g2469) & (!g2471)) + ((g68) & (g87) & (g2468) & (g2469) & (g2471)));
	assign g2473 = (((!g39) & (!g54) & (g2466) & (g2467) & (g2472)) + ((!g39) & (g54) & (g2466) & (!g2467) & (g2472)) + ((!g39) & (g54) & (g2466) & (g2467) & (!g2472)) + ((!g39) & (g54) & (g2466) & (g2467) & (g2472)) + ((g39) & (!g54) & (!g2466) & (g2467) & (g2472)) + ((g39) & (!g54) & (g2466) & (!g2467) & (!g2472)) + ((g39) & (!g54) & (g2466) & (!g2467) & (g2472)) + ((g39) & (!g54) & (g2466) & (g2467) & (!g2472)) + ((g39) & (!g54) & (g2466) & (g2467) & (g2472)) + ((g39) & (g54) & (!g2466) & (!g2467) & (g2472)) + ((g39) & (g54) & (!g2466) & (g2467) & (!g2472)) + ((g39) & (g54) & (!g2466) & (g2467) & (g2472)) + ((g39) & (g54) & (g2466) & (!g2467) & (!g2472)) + ((g39) & (g54) & (g2466) & (!g2467) & (g2472)) + ((g39) & (g54) & (g2466) & (g2467) & (!g2472)) + ((g39) & (g54) & (g2466) & (g2467) & (g2472)));
	assign g2474 = (((!g18) & (!g27) & (g2464) & (g2465) & (g2473)) + ((!g18) & (g27) & (g2464) & (!g2465) & (g2473)) + ((!g18) & (g27) & (g2464) & (g2465) & (!g2473)) + ((!g18) & (g27) & (g2464) & (g2465) & (g2473)) + ((g18) & (!g27) & (!g2464) & (g2465) & (g2473)) + ((g18) & (!g27) & (g2464) & (!g2465) & (!g2473)) + ((g18) & (!g27) & (g2464) & (!g2465) & (g2473)) + ((g18) & (!g27) & (g2464) & (g2465) & (!g2473)) + ((g18) & (!g27) & (g2464) & (g2465) & (g2473)) + ((g18) & (g27) & (!g2464) & (!g2465) & (g2473)) + ((g18) & (g27) & (!g2464) & (g2465) & (!g2473)) + ((g18) & (g27) & (!g2464) & (g2465) & (g2473)) + ((g18) & (g27) & (g2464) & (!g2465) & (!g2473)) + ((g18) & (g27) & (g2464) & (!g2465) & (g2473)) + ((g18) & (g27) & (g2464) & (g2465) & (!g2473)) + ((g18) & (g27) & (g2464) & (g2465) & (g2473)));
	assign g2475 = (((!g2) & (!g8) & (g2462) & (g2463) & (g2474)) + ((!g2) & (g8) & (g2462) & (!g2463) & (g2474)) + ((!g2) & (g8) & (g2462) & (g2463) & (!g2474)) + ((!g2) & (g8) & (g2462) & (g2463) & (g2474)) + ((g2) & (!g8) & (!g2462) & (g2463) & (g2474)) + ((g2) & (!g8) & (g2462) & (!g2463) & (!g2474)) + ((g2) & (!g8) & (g2462) & (!g2463) & (g2474)) + ((g2) & (!g8) & (g2462) & (g2463) & (!g2474)) + ((g2) & (!g8) & (g2462) & (g2463) & (g2474)) + ((g2) & (g8) & (!g2462) & (!g2463) & (g2474)) + ((g2) & (g8) & (!g2462) & (g2463) & (!g2474)) + ((g2) & (g8) & (!g2462) & (g2463) & (g2474)) + ((g2) & (g8) & (g2462) & (!g2463) & (!g2474)) + ((g2) & (g8) & (g2462) & (!g2463) & (g2474)) + ((g2) & (g8) & (g2462) & (g2463) & (!g2474)) + ((g2) & (g8) & (g2462) & (g2463) & (g2474)));
	assign g2476 = (((!g2) & (!g2372) & (g2391) & (!g2398)) + ((!g2) & (g2372) & (!g2391) & (!g2398)) + ((!g2) & (g2372) & (!g2391) & (g2398)) + ((!g2) & (g2372) & (g2391) & (g2398)) + ((g2) & (!g2372) & (!g2391) & (!g2398)) + ((g2) & (g2372) & (!g2391) & (g2398)) + ((g2) & (g2372) & (g2391) & (!g2398)) + ((g2) & (g2372) & (g2391) & (g2398)));
	assign g2477 = (((!g1) & (!g2371) & (!g2394) & (!g2396) & (g2397)) + ((!g1) & (!g2371) & (!g2394) & (g2396) & (!g2397)) + ((!g1) & (!g2371) & (!g2394) & (g2396) & (g2397)) + ((!g1) & (g2371) & (g2394) & (!g2396) & (!g2397)) + ((!g1) & (g2371) & (g2394) & (!g2396) & (g2397)) + ((!g1) & (g2371) & (g2394) & (g2396) & (!g2397)) + ((!g1) & (g2371) & (g2394) & (g2396) & (g2397)) + ((g1) & (!g2371) & (!g2394) & (!g2396) & (g2397)) + ((g1) & (!g2371) & (!g2394) & (g2396) & (g2397)) + ((g1) & (g2371) & (g2394) & (!g2396) & (!g2397)) + ((g1) & (g2371) & (g2394) & (!g2396) & (g2397)) + ((g1) & (g2371) & (g2394) & (g2396) & (!g2397)) + ((g1) & (g2371) & (g2394) & (g2396) & (g2397)));
	assign g2478 = (((!g4) & (!g1) & (!g2461) & (!g2475) & (!g2476) & (!g2477)) + ((!g4) & (g1) & (!g2461) & (!g2475) & (!g2476) & (!g2477)) + ((!g4) & (g1) & (!g2461) & (!g2475) & (!g2476) & (g2477)) + ((!g4) & (g1) & (!g2461) & (!g2475) & (g2476) & (!g2477)) + ((!g4) & (g1) & (!g2461) & (!g2475) & (g2476) & (g2477)) + ((!g4) & (g1) & (!g2461) & (g2475) & (!g2476) & (!g2477)) + ((!g4) & (g1) & (!g2461) & (g2475) & (!g2476) & (g2477)) + ((!g4) & (g1) & (!g2461) & (g2475) & (g2476) & (!g2477)) + ((!g4) & (g1) & (!g2461) & (g2475) & (g2476) & (g2477)) + ((!g4) & (g1) & (g2461) & (!g2475) & (!g2476) & (!g2477)) + ((!g4) & (g1) & (g2461) & (!g2475) & (!g2476) & (g2477)) + ((g4) & (!g1) & (!g2461) & (!g2475) & (!g2476) & (!g2477)) + ((g4) & (!g1) & (!g2461) & (!g2475) & (g2476) & (!g2477)) + ((g4) & (!g1) & (!g2461) & (g2475) & (!g2476) & (!g2477)) + ((g4) & (g1) & (!g2461) & (!g2475) & (!g2476) & (!g2477)) + ((g4) & (g1) & (!g2461) & (!g2475) & (!g2476) & (g2477)) + ((g4) & (g1) & (!g2461) & (!g2475) & (g2476) & (!g2477)) + ((g4) & (g1) & (!g2461) & (!g2475) & (g2476) & (g2477)) + ((g4) & (g1) & (!g2461) & (g2475) & (!g2476) & (!g2477)) + ((g4) & (g1) & (!g2461) & (g2475) & (!g2476) & (g2477)) + ((g4) & (g1) & (!g2461) & (g2475) & (g2476) & (!g2477)) + ((g4) & (g1) & (!g2461) & (g2475) & (g2476) & (g2477)) + ((g4) & (g1) & (g2461) & (!g2475) & (!g2476) & (!g2477)) + ((g4) & (g1) & (g2461) & (!g2475) & (!g2476) & (g2477)) + ((g4) & (g1) & (g2461) & (!g2475) & (g2476) & (!g2477)) + ((g4) & (g1) & (g2461) & (!g2475) & (g2476) & (g2477)) + ((g4) & (g1) & (g2461) & (g2475) & (!g2476) & (!g2477)) + ((g4) & (g1) & (g2461) & (g2475) & (!g2476) & (g2477)));
	assign g2479 = (((!g127) & (!g2399) & (g2459) & (!g2460) & (!g2478)) + ((!g127) & (!g2399) & (g2459) & (g2460) & (!g2478)) + ((!g127) & (!g2399) & (g2459) & (g2460) & (g2478)) + ((!g127) & (g2399) & (!g2459) & (!g2460) & (!g2478)) + ((!g127) & (g2399) & (!g2459) & (!g2460) & (g2478)) + ((!g127) & (g2399) & (!g2459) & (g2460) & (!g2478)) + ((!g127) & (g2399) & (!g2459) & (g2460) & (g2478)) + ((!g127) & (g2399) & (g2459) & (!g2460) & (g2478)) + ((g127) & (!g2399) & (!g2459) & (!g2460) & (!g2478)) + ((g127) & (!g2399) & (!g2459) & (g2460) & (!g2478)) + ((g127) & (!g2399) & (!g2459) & (g2460) & (g2478)) + ((g127) & (g2399) & (!g2459) & (!g2460) & (g2478)) + ((g127) & (g2399) & (g2459) & (!g2460) & (!g2478)) + ((g127) & (g2399) & (g2459) & (!g2460) & (g2478)) + ((g127) & (g2399) & (g2459) & (g2460) & (!g2478)) + ((g127) & (g2399) & (g2459) & (g2460) & (g2478)));
	assign g2480 = (((!g147) & (!g174) & (g2401) & (g2458)) + ((!g147) & (g174) & (!g2401) & (g2458)) + ((!g147) & (g174) & (g2401) & (!g2458)) + ((!g147) & (g174) & (g2401) & (g2458)) + ((g147) & (!g174) & (!g2401) & (!g2458)) + ((g147) & (!g174) & (!g2401) & (g2458)) + ((g147) & (!g174) & (g2401) & (!g2458)) + ((g147) & (g174) & (!g2401) & (!g2458)));
	assign g2481 = (((!g2400) & (!g2460) & (!g2478) & (g2480)) + ((!g2400) & (g2460) & (!g2478) & (g2480)) + ((!g2400) & (g2460) & (g2478) & (g2480)) + ((g2400) & (!g2460) & (!g2478) & (!g2480)) + ((g2400) & (!g2460) & (g2478) & (!g2480)) + ((g2400) & (!g2460) & (g2478) & (g2480)) + ((g2400) & (g2460) & (!g2478) & (!g2480)) + ((g2400) & (g2460) & (g2478) & (!g2480)));
	assign g2482 = (((!g174) & (!g2401) & (g2458) & (!g2460) & (!g2478)) + ((!g174) & (!g2401) & (g2458) & (g2460) & (!g2478)) + ((!g174) & (!g2401) & (g2458) & (g2460) & (g2478)) + ((!g174) & (g2401) & (!g2458) & (!g2460) & (!g2478)) + ((!g174) & (g2401) & (!g2458) & (!g2460) & (g2478)) + ((!g174) & (g2401) & (!g2458) & (g2460) & (!g2478)) + ((!g174) & (g2401) & (!g2458) & (g2460) & (g2478)) + ((!g174) & (g2401) & (g2458) & (!g2460) & (g2478)) + ((g174) & (!g2401) & (!g2458) & (!g2460) & (!g2478)) + ((g174) & (!g2401) & (!g2458) & (g2460) & (!g2478)) + ((g174) & (!g2401) & (!g2458) & (g2460) & (g2478)) + ((g174) & (g2401) & (!g2458) & (!g2460) & (g2478)) + ((g174) & (g2401) & (g2458) & (!g2460) & (!g2478)) + ((g174) & (g2401) & (g2458) & (!g2460) & (g2478)) + ((g174) & (g2401) & (g2458) & (g2460) & (!g2478)) + ((g174) & (g2401) & (g2458) & (g2460) & (g2478)));
	assign g2483 = (((!g198) & (!g229) & (g2403) & (g2457)) + ((!g198) & (g229) & (!g2403) & (g2457)) + ((!g198) & (g229) & (g2403) & (!g2457)) + ((!g198) & (g229) & (g2403) & (g2457)) + ((g198) & (!g229) & (!g2403) & (!g2457)) + ((g198) & (!g229) & (!g2403) & (g2457)) + ((g198) & (!g229) & (g2403) & (!g2457)) + ((g198) & (g229) & (!g2403) & (!g2457)));
	assign g2484 = (((!g2402) & (!g2460) & (!g2478) & (g2483)) + ((!g2402) & (g2460) & (!g2478) & (g2483)) + ((!g2402) & (g2460) & (g2478) & (g2483)) + ((g2402) & (!g2460) & (!g2478) & (!g2483)) + ((g2402) & (!g2460) & (g2478) & (!g2483)) + ((g2402) & (!g2460) & (g2478) & (g2483)) + ((g2402) & (g2460) & (!g2478) & (!g2483)) + ((g2402) & (g2460) & (g2478) & (!g2483)));
	assign g2485 = (((!g229) & (!g2403) & (g2457) & (!g2460) & (!g2478)) + ((!g229) & (!g2403) & (g2457) & (g2460) & (!g2478)) + ((!g229) & (!g2403) & (g2457) & (g2460) & (g2478)) + ((!g229) & (g2403) & (!g2457) & (!g2460) & (!g2478)) + ((!g229) & (g2403) & (!g2457) & (!g2460) & (g2478)) + ((!g229) & (g2403) & (!g2457) & (g2460) & (!g2478)) + ((!g229) & (g2403) & (!g2457) & (g2460) & (g2478)) + ((!g229) & (g2403) & (g2457) & (!g2460) & (g2478)) + ((g229) & (!g2403) & (!g2457) & (!g2460) & (!g2478)) + ((g229) & (!g2403) & (!g2457) & (g2460) & (!g2478)) + ((g229) & (!g2403) & (!g2457) & (g2460) & (g2478)) + ((g229) & (g2403) & (!g2457) & (!g2460) & (g2478)) + ((g229) & (g2403) & (g2457) & (!g2460) & (!g2478)) + ((g229) & (g2403) & (g2457) & (!g2460) & (g2478)) + ((g229) & (g2403) & (g2457) & (g2460) & (!g2478)) + ((g229) & (g2403) & (g2457) & (g2460) & (g2478)));
	assign g2486 = (((!g255) & (!g290) & (g2405) & (g2456)) + ((!g255) & (g290) & (!g2405) & (g2456)) + ((!g255) & (g290) & (g2405) & (!g2456)) + ((!g255) & (g290) & (g2405) & (g2456)) + ((g255) & (!g290) & (!g2405) & (!g2456)) + ((g255) & (!g290) & (!g2405) & (g2456)) + ((g255) & (!g290) & (g2405) & (!g2456)) + ((g255) & (g290) & (!g2405) & (!g2456)));
	assign g2487 = (((!g2404) & (!g2460) & (!g2478) & (g2486)) + ((!g2404) & (g2460) & (!g2478) & (g2486)) + ((!g2404) & (g2460) & (g2478) & (g2486)) + ((g2404) & (!g2460) & (!g2478) & (!g2486)) + ((g2404) & (!g2460) & (g2478) & (!g2486)) + ((g2404) & (!g2460) & (g2478) & (g2486)) + ((g2404) & (g2460) & (!g2478) & (!g2486)) + ((g2404) & (g2460) & (g2478) & (!g2486)));
	assign g2488 = (((!g290) & (!g2405) & (g2456) & (!g2460) & (!g2478)) + ((!g290) & (!g2405) & (g2456) & (g2460) & (!g2478)) + ((!g290) & (!g2405) & (g2456) & (g2460) & (g2478)) + ((!g290) & (g2405) & (!g2456) & (!g2460) & (!g2478)) + ((!g290) & (g2405) & (!g2456) & (!g2460) & (g2478)) + ((!g290) & (g2405) & (!g2456) & (g2460) & (!g2478)) + ((!g290) & (g2405) & (!g2456) & (g2460) & (g2478)) + ((!g290) & (g2405) & (g2456) & (!g2460) & (g2478)) + ((g290) & (!g2405) & (!g2456) & (!g2460) & (!g2478)) + ((g290) & (!g2405) & (!g2456) & (g2460) & (!g2478)) + ((g290) & (!g2405) & (!g2456) & (g2460) & (g2478)) + ((g290) & (g2405) & (!g2456) & (!g2460) & (g2478)) + ((g290) & (g2405) & (g2456) & (!g2460) & (!g2478)) + ((g290) & (g2405) & (g2456) & (!g2460) & (g2478)) + ((g290) & (g2405) & (g2456) & (g2460) & (!g2478)) + ((g290) & (g2405) & (g2456) & (g2460) & (g2478)));
	assign g2489 = (((!g319) & (!g358) & (g2407) & (g2455)) + ((!g319) & (g358) & (!g2407) & (g2455)) + ((!g319) & (g358) & (g2407) & (!g2455)) + ((!g319) & (g358) & (g2407) & (g2455)) + ((g319) & (!g358) & (!g2407) & (!g2455)) + ((g319) & (!g358) & (!g2407) & (g2455)) + ((g319) & (!g358) & (g2407) & (!g2455)) + ((g319) & (g358) & (!g2407) & (!g2455)));
	assign g2490 = (((!g2406) & (!g2460) & (!g2478) & (g2489)) + ((!g2406) & (g2460) & (!g2478) & (g2489)) + ((!g2406) & (g2460) & (g2478) & (g2489)) + ((g2406) & (!g2460) & (!g2478) & (!g2489)) + ((g2406) & (!g2460) & (g2478) & (!g2489)) + ((g2406) & (!g2460) & (g2478) & (g2489)) + ((g2406) & (g2460) & (!g2478) & (!g2489)) + ((g2406) & (g2460) & (g2478) & (!g2489)));
	assign g2491 = (((!g358) & (!g2407) & (g2455) & (!g2460) & (!g2478)) + ((!g358) & (!g2407) & (g2455) & (g2460) & (!g2478)) + ((!g358) & (!g2407) & (g2455) & (g2460) & (g2478)) + ((!g358) & (g2407) & (!g2455) & (!g2460) & (!g2478)) + ((!g358) & (g2407) & (!g2455) & (!g2460) & (g2478)) + ((!g358) & (g2407) & (!g2455) & (g2460) & (!g2478)) + ((!g358) & (g2407) & (!g2455) & (g2460) & (g2478)) + ((!g358) & (g2407) & (g2455) & (!g2460) & (g2478)) + ((g358) & (!g2407) & (!g2455) & (!g2460) & (!g2478)) + ((g358) & (!g2407) & (!g2455) & (g2460) & (!g2478)) + ((g358) & (!g2407) & (!g2455) & (g2460) & (g2478)) + ((g358) & (g2407) & (!g2455) & (!g2460) & (g2478)) + ((g358) & (g2407) & (g2455) & (!g2460) & (!g2478)) + ((g358) & (g2407) & (g2455) & (!g2460) & (g2478)) + ((g358) & (g2407) & (g2455) & (g2460) & (!g2478)) + ((g358) & (g2407) & (g2455) & (g2460) & (g2478)));
	assign g2492 = (((!g390) & (!g433) & (g2409) & (g2454)) + ((!g390) & (g433) & (!g2409) & (g2454)) + ((!g390) & (g433) & (g2409) & (!g2454)) + ((!g390) & (g433) & (g2409) & (g2454)) + ((g390) & (!g433) & (!g2409) & (!g2454)) + ((g390) & (!g433) & (!g2409) & (g2454)) + ((g390) & (!g433) & (g2409) & (!g2454)) + ((g390) & (g433) & (!g2409) & (!g2454)));
	assign g2493 = (((!g2408) & (!g2460) & (!g2478) & (g2492)) + ((!g2408) & (g2460) & (!g2478) & (g2492)) + ((!g2408) & (g2460) & (g2478) & (g2492)) + ((g2408) & (!g2460) & (!g2478) & (!g2492)) + ((g2408) & (!g2460) & (g2478) & (!g2492)) + ((g2408) & (!g2460) & (g2478) & (g2492)) + ((g2408) & (g2460) & (!g2478) & (!g2492)) + ((g2408) & (g2460) & (g2478) & (!g2492)));
	assign g2494 = (((!g433) & (!g2409) & (g2454) & (!g2460) & (!g2478)) + ((!g433) & (!g2409) & (g2454) & (g2460) & (!g2478)) + ((!g433) & (!g2409) & (g2454) & (g2460) & (g2478)) + ((!g433) & (g2409) & (!g2454) & (!g2460) & (!g2478)) + ((!g433) & (g2409) & (!g2454) & (!g2460) & (g2478)) + ((!g433) & (g2409) & (!g2454) & (g2460) & (!g2478)) + ((!g433) & (g2409) & (!g2454) & (g2460) & (g2478)) + ((!g433) & (g2409) & (g2454) & (!g2460) & (g2478)) + ((g433) & (!g2409) & (!g2454) & (!g2460) & (!g2478)) + ((g433) & (!g2409) & (!g2454) & (g2460) & (!g2478)) + ((g433) & (!g2409) & (!g2454) & (g2460) & (g2478)) + ((g433) & (g2409) & (!g2454) & (!g2460) & (g2478)) + ((g433) & (g2409) & (g2454) & (!g2460) & (!g2478)) + ((g433) & (g2409) & (g2454) & (!g2460) & (g2478)) + ((g433) & (g2409) & (g2454) & (g2460) & (!g2478)) + ((g433) & (g2409) & (g2454) & (g2460) & (g2478)));
	assign g2495 = (((!g468) & (!g515) & (g2411) & (g2453)) + ((!g468) & (g515) & (!g2411) & (g2453)) + ((!g468) & (g515) & (g2411) & (!g2453)) + ((!g468) & (g515) & (g2411) & (g2453)) + ((g468) & (!g515) & (!g2411) & (!g2453)) + ((g468) & (!g515) & (!g2411) & (g2453)) + ((g468) & (!g515) & (g2411) & (!g2453)) + ((g468) & (g515) & (!g2411) & (!g2453)));
	assign g2496 = (((!g2410) & (!g2460) & (!g2478) & (g2495)) + ((!g2410) & (g2460) & (!g2478) & (g2495)) + ((!g2410) & (g2460) & (g2478) & (g2495)) + ((g2410) & (!g2460) & (!g2478) & (!g2495)) + ((g2410) & (!g2460) & (g2478) & (!g2495)) + ((g2410) & (!g2460) & (g2478) & (g2495)) + ((g2410) & (g2460) & (!g2478) & (!g2495)) + ((g2410) & (g2460) & (g2478) & (!g2495)));
	assign g2497 = (((!g515) & (!g2411) & (g2453) & (!g2460) & (!g2478)) + ((!g515) & (!g2411) & (g2453) & (g2460) & (!g2478)) + ((!g515) & (!g2411) & (g2453) & (g2460) & (g2478)) + ((!g515) & (g2411) & (!g2453) & (!g2460) & (!g2478)) + ((!g515) & (g2411) & (!g2453) & (!g2460) & (g2478)) + ((!g515) & (g2411) & (!g2453) & (g2460) & (!g2478)) + ((!g515) & (g2411) & (!g2453) & (g2460) & (g2478)) + ((!g515) & (g2411) & (g2453) & (!g2460) & (g2478)) + ((g515) & (!g2411) & (!g2453) & (!g2460) & (!g2478)) + ((g515) & (!g2411) & (!g2453) & (g2460) & (!g2478)) + ((g515) & (!g2411) & (!g2453) & (g2460) & (g2478)) + ((g515) & (g2411) & (!g2453) & (!g2460) & (g2478)) + ((g515) & (g2411) & (g2453) & (!g2460) & (!g2478)) + ((g515) & (g2411) & (g2453) & (!g2460) & (g2478)) + ((g515) & (g2411) & (g2453) & (g2460) & (!g2478)) + ((g515) & (g2411) & (g2453) & (g2460) & (g2478)));
	assign g2498 = (((!g553) & (!g604) & (g2413) & (g2452)) + ((!g553) & (g604) & (!g2413) & (g2452)) + ((!g553) & (g604) & (g2413) & (!g2452)) + ((!g553) & (g604) & (g2413) & (g2452)) + ((g553) & (!g604) & (!g2413) & (!g2452)) + ((g553) & (!g604) & (!g2413) & (g2452)) + ((g553) & (!g604) & (g2413) & (!g2452)) + ((g553) & (g604) & (!g2413) & (!g2452)));
	assign g2499 = (((!g2412) & (!g2460) & (!g2478) & (g2498)) + ((!g2412) & (g2460) & (!g2478) & (g2498)) + ((!g2412) & (g2460) & (g2478) & (g2498)) + ((g2412) & (!g2460) & (!g2478) & (!g2498)) + ((g2412) & (!g2460) & (g2478) & (!g2498)) + ((g2412) & (!g2460) & (g2478) & (g2498)) + ((g2412) & (g2460) & (!g2478) & (!g2498)) + ((g2412) & (g2460) & (g2478) & (!g2498)));
	assign g2500 = (((!g604) & (!g2413) & (g2452) & (!g2460) & (!g2478)) + ((!g604) & (!g2413) & (g2452) & (g2460) & (!g2478)) + ((!g604) & (!g2413) & (g2452) & (g2460) & (g2478)) + ((!g604) & (g2413) & (!g2452) & (!g2460) & (!g2478)) + ((!g604) & (g2413) & (!g2452) & (!g2460) & (g2478)) + ((!g604) & (g2413) & (!g2452) & (g2460) & (!g2478)) + ((!g604) & (g2413) & (!g2452) & (g2460) & (g2478)) + ((!g604) & (g2413) & (g2452) & (!g2460) & (g2478)) + ((g604) & (!g2413) & (!g2452) & (!g2460) & (!g2478)) + ((g604) & (!g2413) & (!g2452) & (g2460) & (!g2478)) + ((g604) & (!g2413) & (!g2452) & (g2460) & (g2478)) + ((g604) & (g2413) & (!g2452) & (!g2460) & (g2478)) + ((g604) & (g2413) & (g2452) & (!g2460) & (!g2478)) + ((g604) & (g2413) & (g2452) & (!g2460) & (g2478)) + ((g604) & (g2413) & (g2452) & (g2460) & (!g2478)) + ((g604) & (g2413) & (g2452) & (g2460) & (g2478)));
	assign g2501 = (((!g645) & (!g700) & (g2415) & (g2451)) + ((!g645) & (g700) & (!g2415) & (g2451)) + ((!g645) & (g700) & (g2415) & (!g2451)) + ((!g645) & (g700) & (g2415) & (g2451)) + ((g645) & (!g700) & (!g2415) & (!g2451)) + ((g645) & (!g700) & (!g2415) & (g2451)) + ((g645) & (!g700) & (g2415) & (!g2451)) + ((g645) & (g700) & (!g2415) & (!g2451)));
	assign g2502 = (((!g2414) & (!g2460) & (!g2478) & (g2501)) + ((!g2414) & (g2460) & (!g2478) & (g2501)) + ((!g2414) & (g2460) & (g2478) & (g2501)) + ((g2414) & (!g2460) & (!g2478) & (!g2501)) + ((g2414) & (!g2460) & (g2478) & (!g2501)) + ((g2414) & (!g2460) & (g2478) & (g2501)) + ((g2414) & (g2460) & (!g2478) & (!g2501)) + ((g2414) & (g2460) & (g2478) & (!g2501)));
	assign g2503 = (((!g700) & (!g2415) & (g2451) & (!g2460) & (!g2478)) + ((!g700) & (!g2415) & (g2451) & (g2460) & (!g2478)) + ((!g700) & (!g2415) & (g2451) & (g2460) & (g2478)) + ((!g700) & (g2415) & (!g2451) & (!g2460) & (!g2478)) + ((!g700) & (g2415) & (!g2451) & (!g2460) & (g2478)) + ((!g700) & (g2415) & (!g2451) & (g2460) & (!g2478)) + ((!g700) & (g2415) & (!g2451) & (g2460) & (g2478)) + ((!g700) & (g2415) & (g2451) & (!g2460) & (g2478)) + ((g700) & (!g2415) & (!g2451) & (!g2460) & (!g2478)) + ((g700) & (!g2415) & (!g2451) & (g2460) & (!g2478)) + ((g700) & (!g2415) & (!g2451) & (g2460) & (g2478)) + ((g700) & (g2415) & (!g2451) & (!g2460) & (g2478)) + ((g700) & (g2415) & (g2451) & (!g2460) & (!g2478)) + ((g700) & (g2415) & (g2451) & (!g2460) & (g2478)) + ((g700) & (g2415) & (g2451) & (g2460) & (!g2478)) + ((g700) & (g2415) & (g2451) & (g2460) & (g2478)));
	assign g2504 = (((!g744) & (!g803) & (g2417) & (g2450)) + ((!g744) & (g803) & (!g2417) & (g2450)) + ((!g744) & (g803) & (g2417) & (!g2450)) + ((!g744) & (g803) & (g2417) & (g2450)) + ((g744) & (!g803) & (!g2417) & (!g2450)) + ((g744) & (!g803) & (!g2417) & (g2450)) + ((g744) & (!g803) & (g2417) & (!g2450)) + ((g744) & (g803) & (!g2417) & (!g2450)));
	assign g2505 = (((!g2416) & (!g2460) & (!g2478) & (g2504)) + ((!g2416) & (g2460) & (!g2478) & (g2504)) + ((!g2416) & (g2460) & (g2478) & (g2504)) + ((g2416) & (!g2460) & (!g2478) & (!g2504)) + ((g2416) & (!g2460) & (g2478) & (!g2504)) + ((g2416) & (!g2460) & (g2478) & (g2504)) + ((g2416) & (g2460) & (!g2478) & (!g2504)) + ((g2416) & (g2460) & (g2478) & (!g2504)));
	assign g2506 = (((!g803) & (!g2417) & (g2450) & (!g2460) & (!g2478)) + ((!g803) & (!g2417) & (g2450) & (g2460) & (!g2478)) + ((!g803) & (!g2417) & (g2450) & (g2460) & (g2478)) + ((!g803) & (g2417) & (!g2450) & (!g2460) & (!g2478)) + ((!g803) & (g2417) & (!g2450) & (!g2460) & (g2478)) + ((!g803) & (g2417) & (!g2450) & (g2460) & (!g2478)) + ((!g803) & (g2417) & (!g2450) & (g2460) & (g2478)) + ((!g803) & (g2417) & (g2450) & (!g2460) & (g2478)) + ((g803) & (!g2417) & (!g2450) & (!g2460) & (!g2478)) + ((g803) & (!g2417) & (!g2450) & (g2460) & (!g2478)) + ((g803) & (!g2417) & (!g2450) & (g2460) & (g2478)) + ((g803) & (g2417) & (!g2450) & (!g2460) & (g2478)) + ((g803) & (g2417) & (g2450) & (!g2460) & (!g2478)) + ((g803) & (g2417) & (g2450) & (!g2460) & (g2478)) + ((g803) & (g2417) & (g2450) & (g2460) & (!g2478)) + ((g803) & (g2417) & (g2450) & (g2460) & (g2478)));
	assign g2507 = (((!g851) & (!g914) & (g2419) & (g2449)) + ((!g851) & (g914) & (!g2419) & (g2449)) + ((!g851) & (g914) & (g2419) & (!g2449)) + ((!g851) & (g914) & (g2419) & (g2449)) + ((g851) & (!g914) & (!g2419) & (!g2449)) + ((g851) & (!g914) & (!g2419) & (g2449)) + ((g851) & (!g914) & (g2419) & (!g2449)) + ((g851) & (g914) & (!g2419) & (!g2449)));
	assign g2508 = (((!g2418) & (!g2460) & (!g2478) & (g2507)) + ((!g2418) & (g2460) & (!g2478) & (g2507)) + ((!g2418) & (g2460) & (g2478) & (g2507)) + ((g2418) & (!g2460) & (!g2478) & (!g2507)) + ((g2418) & (!g2460) & (g2478) & (!g2507)) + ((g2418) & (!g2460) & (g2478) & (g2507)) + ((g2418) & (g2460) & (!g2478) & (!g2507)) + ((g2418) & (g2460) & (g2478) & (!g2507)));
	assign g2509 = (((!g914) & (!g2419) & (g2449) & (!g2460) & (!g2478)) + ((!g914) & (!g2419) & (g2449) & (g2460) & (!g2478)) + ((!g914) & (!g2419) & (g2449) & (g2460) & (g2478)) + ((!g914) & (g2419) & (!g2449) & (!g2460) & (!g2478)) + ((!g914) & (g2419) & (!g2449) & (!g2460) & (g2478)) + ((!g914) & (g2419) & (!g2449) & (g2460) & (!g2478)) + ((!g914) & (g2419) & (!g2449) & (g2460) & (g2478)) + ((!g914) & (g2419) & (g2449) & (!g2460) & (g2478)) + ((g914) & (!g2419) & (!g2449) & (!g2460) & (!g2478)) + ((g914) & (!g2419) & (!g2449) & (g2460) & (!g2478)) + ((g914) & (!g2419) & (!g2449) & (g2460) & (g2478)) + ((g914) & (g2419) & (!g2449) & (!g2460) & (g2478)) + ((g914) & (g2419) & (g2449) & (!g2460) & (!g2478)) + ((g914) & (g2419) & (g2449) & (!g2460) & (g2478)) + ((g914) & (g2419) & (g2449) & (g2460) & (!g2478)) + ((g914) & (g2419) & (g2449) & (g2460) & (g2478)));
	assign g2510 = (((!g1032) & (!g1030) & (g2421) & (g2448)) + ((!g1032) & (g1030) & (!g2421) & (g2448)) + ((!g1032) & (g1030) & (g2421) & (!g2448)) + ((!g1032) & (g1030) & (g2421) & (g2448)) + ((g1032) & (!g1030) & (!g2421) & (!g2448)) + ((g1032) & (!g1030) & (!g2421) & (g2448)) + ((g1032) & (!g1030) & (g2421) & (!g2448)) + ((g1032) & (g1030) & (!g2421) & (!g2448)));
	assign g2511 = (((!g2420) & (!g2460) & (!g2478) & (g2510)) + ((!g2420) & (g2460) & (!g2478) & (g2510)) + ((!g2420) & (g2460) & (g2478) & (g2510)) + ((g2420) & (!g2460) & (!g2478) & (!g2510)) + ((g2420) & (!g2460) & (g2478) & (!g2510)) + ((g2420) & (!g2460) & (g2478) & (g2510)) + ((g2420) & (g2460) & (!g2478) & (!g2510)) + ((g2420) & (g2460) & (g2478) & (!g2510)));
	assign g2512 = (((!g1030) & (!g2421) & (g2448) & (!g2460) & (!g2478)) + ((!g1030) & (!g2421) & (g2448) & (g2460) & (!g2478)) + ((!g1030) & (!g2421) & (g2448) & (g2460) & (g2478)) + ((!g1030) & (g2421) & (!g2448) & (!g2460) & (!g2478)) + ((!g1030) & (g2421) & (!g2448) & (!g2460) & (g2478)) + ((!g1030) & (g2421) & (!g2448) & (g2460) & (!g2478)) + ((!g1030) & (g2421) & (!g2448) & (g2460) & (g2478)) + ((!g1030) & (g2421) & (g2448) & (!g2460) & (g2478)) + ((g1030) & (!g2421) & (!g2448) & (!g2460) & (!g2478)) + ((g1030) & (!g2421) & (!g2448) & (g2460) & (!g2478)) + ((g1030) & (!g2421) & (!g2448) & (g2460) & (g2478)) + ((g1030) & (g2421) & (!g2448) & (!g2460) & (g2478)) + ((g1030) & (g2421) & (g2448) & (!g2460) & (!g2478)) + ((g1030) & (g2421) & (g2448) & (!g2460) & (g2478)) + ((g1030) & (g2421) & (g2448) & (g2460) & (!g2478)) + ((g1030) & (g2421) & (g2448) & (g2460) & (g2478)));
	assign g2513 = (((!g1160) & (!g1154) & (g2423) & (g2447)) + ((!g1160) & (g1154) & (!g2423) & (g2447)) + ((!g1160) & (g1154) & (g2423) & (!g2447)) + ((!g1160) & (g1154) & (g2423) & (g2447)) + ((g1160) & (!g1154) & (!g2423) & (!g2447)) + ((g1160) & (!g1154) & (!g2423) & (g2447)) + ((g1160) & (!g1154) & (g2423) & (!g2447)) + ((g1160) & (g1154) & (!g2423) & (!g2447)));
	assign g2514 = (((!g2422) & (!g2460) & (!g2478) & (g2513)) + ((!g2422) & (g2460) & (!g2478) & (g2513)) + ((!g2422) & (g2460) & (g2478) & (g2513)) + ((g2422) & (!g2460) & (!g2478) & (!g2513)) + ((g2422) & (!g2460) & (g2478) & (!g2513)) + ((g2422) & (!g2460) & (g2478) & (g2513)) + ((g2422) & (g2460) & (!g2478) & (!g2513)) + ((g2422) & (g2460) & (g2478) & (!g2513)));
	assign g2515 = (((!g1154) & (!g2423) & (g2447) & (!g2460) & (!g2478)) + ((!g1154) & (!g2423) & (g2447) & (g2460) & (!g2478)) + ((!g1154) & (!g2423) & (g2447) & (g2460) & (g2478)) + ((!g1154) & (g2423) & (!g2447) & (!g2460) & (!g2478)) + ((!g1154) & (g2423) & (!g2447) & (!g2460) & (g2478)) + ((!g1154) & (g2423) & (!g2447) & (g2460) & (!g2478)) + ((!g1154) & (g2423) & (!g2447) & (g2460) & (g2478)) + ((!g1154) & (g2423) & (g2447) & (!g2460) & (g2478)) + ((g1154) & (!g2423) & (!g2447) & (!g2460) & (!g2478)) + ((g1154) & (!g2423) & (!g2447) & (g2460) & (!g2478)) + ((g1154) & (!g2423) & (!g2447) & (g2460) & (g2478)) + ((g1154) & (g2423) & (!g2447) & (!g2460) & (g2478)) + ((g1154) & (g2423) & (g2447) & (!g2460) & (!g2478)) + ((g1154) & (g2423) & (g2447) & (!g2460) & (g2478)) + ((g1154) & (g2423) & (g2447) & (g2460) & (!g2478)) + ((g1154) & (g2423) & (g2447) & (g2460) & (g2478)));
	assign g2516 = (((!g1295) & (!g1285) & (g2425) & (g2446)) + ((!g1295) & (g1285) & (!g2425) & (g2446)) + ((!g1295) & (g1285) & (g2425) & (!g2446)) + ((!g1295) & (g1285) & (g2425) & (g2446)) + ((g1295) & (!g1285) & (!g2425) & (!g2446)) + ((g1295) & (!g1285) & (!g2425) & (g2446)) + ((g1295) & (!g1285) & (g2425) & (!g2446)) + ((g1295) & (g1285) & (!g2425) & (!g2446)));
	assign g2517 = (((!g2424) & (!g2460) & (!g2478) & (g2516)) + ((!g2424) & (g2460) & (!g2478) & (g2516)) + ((!g2424) & (g2460) & (g2478) & (g2516)) + ((g2424) & (!g2460) & (!g2478) & (!g2516)) + ((g2424) & (!g2460) & (g2478) & (!g2516)) + ((g2424) & (!g2460) & (g2478) & (g2516)) + ((g2424) & (g2460) & (!g2478) & (!g2516)) + ((g2424) & (g2460) & (g2478) & (!g2516)));
	assign g2518 = (((!g1285) & (!g2425) & (g2446) & (!g2460) & (!g2478)) + ((!g1285) & (!g2425) & (g2446) & (g2460) & (!g2478)) + ((!g1285) & (!g2425) & (g2446) & (g2460) & (g2478)) + ((!g1285) & (g2425) & (!g2446) & (!g2460) & (!g2478)) + ((!g1285) & (g2425) & (!g2446) & (!g2460) & (g2478)) + ((!g1285) & (g2425) & (!g2446) & (g2460) & (!g2478)) + ((!g1285) & (g2425) & (!g2446) & (g2460) & (g2478)) + ((!g1285) & (g2425) & (g2446) & (!g2460) & (g2478)) + ((g1285) & (!g2425) & (!g2446) & (!g2460) & (!g2478)) + ((g1285) & (!g2425) & (!g2446) & (g2460) & (!g2478)) + ((g1285) & (!g2425) & (!g2446) & (g2460) & (g2478)) + ((g1285) & (g2425) & (!g2446) & (!g2460) & (g2478)) + ((g1285) & (g2425) & (g2446) & (!g2460) & (!g2478)) + ((g1285) & (g2425) & (g2446) & (!g2460) & (g2478)) + ((g1285) & (g2425) & (g2446) & (g2460) & (!g2478)) + ((g1285) & (g2425) & (g2446) & (g2460) & (g2478)));
	assign g2519 = (((!g1437) & (!g1423) & (g2427) & (g2445)) + ((!g1437) & (g1423) & (!g2427) & (g2445)) + ((!g1437) & (g1423) & (g2427) & (!g2445)) + ((!g1437) & (g1423) & (g2427) & (g2445)) + ((g1437) & (!g1423) & (!g2427) & (!g2445)) + ((g1437) & (!g1423) & (!g2427) & (g2445)) + ((g1437) & (!g1423) & (g2427) & (!g2445)) + ((g1437) & (g1423) & (!g2427) & (!g2445)));
	assign g2520 = (((!g2426) & (!g2460) & (!g2478) & (g2519)) + ((!g2426) & (g2460) & (!g2478) & (g2519)) + ((!g2426) & (g2460) & (g2478) & (g2519)) + ((g2426) & (!g2460) & (!g2478) & (!g2519)) + ((g2426) & (!g2460) & (g2478) & (!g2519)) + ((g2426) & (!g2460) & (g2478) & (g2519)) + ((g2426) & (g2460) & (!g2478) & (!g2519)) + ((g2426) & (g2460) & (g2478) & (!g2519)));
	assign g2521 = (((!g1423) & (!g2427) & (g2445) & (!g2460) & (!g2478)) + ((!g1423) & (!g2427) & (g2445) & (g2460) & (!g2478)) + ((!g1423) & (!g2427) & (g2445) & (g2460) & (g2478)) + ((!g1423) & (g2427) & (!g2445) & (!g2460) & (!g2478)) + ((!g1423) & (g2427) & (!g2445) & (!g2460) & (g2478)) + ((!g1423) & (g2427) & (!g2445) & (g2460) & (!g2478)) + ((!g1423) & (g2427) & (!g2445) & (g2460) & (g2478)) + ((!g1423) & (g2427) & (g2445) & (!g2460) & (g2478)) + ((g1423) & (!g2427) & (!g2445) & (!g2460) & (!g2478)) + ((g1423) & (!g2427) & (!g2445) & (g2460) & (!g2478)) + ((g1423) & (!g2427) & (!g2445) & (g2460) & (g2478)) + ((g1423) & (g2427) & (!g2445) & (!g2460) & (g2478)) + ((g1423) & (g2427) & (g2445) & (!g2460) & (!g2478)) + ((g1423) & (g2427) & (g2445) & (!g2460) & (g2478)) + ((g1423) & (g2427) & (g2445) & (g2460) & (!g2478)) + ((g1423) & (g2427) & (g2445) & (g2460) & (g2478)));
	assign g2522 = (((!g1586) & (!g1568) & (g2429) & (g2444)) + ((!g1586) & (g1568) & (!g2429) & (g2444)) + ((!g1586) & (g1568) & (g2429) & (!g2444)) + ((!g1586) & (g1568) & (g2429) & (g2444)) + ((g1586) & (!g1568) & (!g2429) & (!g2444)) + ((g1586) & (!g1568) & (!g2429) & (g2444)) + ((g1586) & (!g1568) & (g2429) & (!g2444)) + ((g1586) & (g1568) & (!g2429) & (!g2444)));
	assign g2523 = (((!g2428) & (!g2460) & (!g2478) & (g2522)) + ((!g2428) & (g2460) & (!g2478) & (g2522)) + ((!g2428) & (g2460) & (g2478) & (g2522)) + ((g2428) & (!g2460) & (!g2478) & (!g2522)) + ((g2428) & (!g2460) & (g2478) & (!g2522)) + ((g2428) & (!g2460) & (g2478) & (g2522)) + ((g2428) & (g2460) & (!g2478) & (!g2522)) + ((g2428) & (g2460) & (g2478) & (!g2522)));
	assign g2524 = (((!g1568) & (!g2429) & (g2444) & (!g2460) & (!g2478)) + ((!g1568) & (!g2429) & (g2444) & (g2460) & (!g2478)) + ((!g1568) & (!g2429) & (g2444) & (g2460) & (g2478)) + ((!g1568) & (g2429) & (!g2444) & (!g2460) & (!g2478)) + ((!g1568) & (g2429) & (!g2444) & (!g2460) & (g2478)) + ((!g1568) & (g2429) & (!g2444) & (g2460) & (!g2478)) + ((!g1568) & (g2429) & (!g2444) & (g2460) & (g2478)) + ((!g1568) & (g2429) & (g2444) & (!g2460) & (g2478)) + ((g1568) & (!g2429) & (!g2444) & (!g2460) & (!g2478)) + ((g1568) & (!g2429) & (!g2444) & (g2460) & (!g2478)) + ((g1568) & (!g2429) & (!g2444) & (g2460) & (g2478)) + ((g1568) & (g2429) & (!g2444) & (!g2460) & (g2478)) + ((g1568) & (g2429) & (g2444) & (!g2460) & (!g2478)) + ((g1568) & (g2429) & (g2444) & (!g2460) & (g2478)) + ((g1568) & (g2429) & (g2444) & (g2460) & (!g2478)) + ((g1568) & (g2429) & (g2444) & (g2460) & (g2478)));
	assign g2525 = (((!g1742) & (!g1720) & (g2431) & (g2443)) + ((!g1742) & (g1720) & (!g2431) & (g2443)) + ((!g1742) & (g1720) & (g2431) & (!g2443)) + ((!g1742) & (g1720) & (g2431) & (g2443)) + ((g1742) & (!g1720) & (!g2431) & (!g2443)) + ((g1742) & (!g1720) & (!g2431) & (g2443)) + ((g1742) & (!g1720) & (g2431) & (!g2443)) + ((g1742) & (g1720) & (!g2431) & (!g2443)));
	assign g2526 = (((!g2430) & (!g2460) & (!g2478) & (g2525)) + ((!g2430) & (g2460) & (!g2478) & (g2525)) + ((!g2430) & (g2460) & (g2478) & (g2525)) + ((g2430) & (!g2460) & (!g2478) & (!g2525)) + ((g2430) & (!g2460) & (g2478) & (!g2525)) + ((g2430) & (!g2460) & (g2478) & (g2525)) + ((g2430) & (g2460) & (!g2478) & (!g2525)) + ((g2430) & (g2460) & (g2478) & (!g2525)));
	assign g2527 = (((!g1720) & (!g2431) & (g2443) & (!g2460) & (!g2478)) + ((!g1720) & (!g2431) & (g2443) & (g2460) & (!g2478)) + ((!g1720) & (!g2431) & (g2443) & (g2460) & (g2478)) + ((!g1720) & (g2431) & (!g2443) & (!g2460) & (!g2478)) + ((!g1720) & (g2431) & (!g2443) & (!g2460) & (g2478)) + ((!g1720) & (g2431) & (!g2443) & (g2460) & (!g2478)) + ((!g1720) & (g2431) & (!g2443) & (g2460) & (g2478)) + ((!g1720) & (g2431) & (g2443) & (!g2460) & (g2478)) + ((g1720) & (!g2431) & (!g2443) & (!g2460) & (!g2478)) + ((g1720) & (!g2431) & (!g2443) & (g2460) & (!g2478)) + ((g1720) & (!g2431) & (!g2443) & (g2460) & (g2478)) + ((g1720) & (g2431) & (!g2443) & (!g2460) & (g2478)) + ((g1720) & (g2431) & (g2443) & (!g2460) & (!g2478)) + ((g1720) & (g2431) & (g2443) & (!g2460) & (g2478)) + ((g1720) & (g2431) & (g2443) & (g2460) & (!g2478)) + ((g1720) & (g2431) & (g2443) & (g2460) & (g2478)));
	assign g2528 = (((!g1905) & (!g1879) & (g2433) & (g2442)) + ((!g1905) & (g1879) & (!g2433) & (g2442)) + ((!g1905) & (g1879) & (g2433) & (!g2442)) + ((!g1905) & (g1879) & (g2433) & (g2442)) + ((g1905) & (!g1879) & (!g2433) & (!g2442)) + ((g1905) & (!g1879) & (!g2433) & (g2442)) + ((g1905) & (!g1879) & (g2433) & (!g2442)) + ((g1905) & (g1879) & (!g2433) & (!g2442)));
	assign g2529 = (((!g2432) & (!g2460) & (!g2478) & (g2528)) + ((!g2432) & (g2460) & (!g2478) & (g2528)) + ((!g2432) & (g2460) & (g2478) & (g2528)) + ((g2432) & (!g2460) & (!g2478) & (!g2528)) + ((g2432) & (!g2460) & (g2478) & (!g2528)) + ((g2432) & (!g2460) & (g2478) & (g2528)) + ((g2432) & (g2460) & (!g2478) & (!g2528)) + ((g2432) & (g2460) & (g2478) & (!g2528)));
	assign g2530 = (((!g1879) & (!g2433) & (g2442) & (!g2460) & (!g2478)) + ((!g1879) & (!g2433) & (g2442) & (g2460) & (!g2478)) + ((!g1879) & (!g2433) & (g2442) & (g2460) & (g2478)) + ((!g1879) & (g2433) & (!g2442) & (!g2460) & (!g2478)) + ((!g1879) & (g2433) & (!g2442) & (!g2460) & (g2478)) + ((!g1879) & (g2433) & (!g2442) & (g2460) & (!g2478)) + ((!g1879) & (g2433) & (!g2442) & (g2460) & (g2478)) + ((!g1879) & (g2433) & (g2442) & (!g2460) & (g2478)) + ((g1879) & (!g2433) & (!g2442) & (!g2460) & (!g2478)) + ((g1879) & (!g2433) & (!g2442) & (g2460) & (!g2478)) + ((g1879) & (!g2433) & (!g2442) & (g2460) & (g2478)) + ((g1879) & (g2433) & (!g2442) & (!g2460) & (g2478)) + ((g1879) & (g2433) & (g2442) & (!g2460) & (!g2478)) + ((g1879) & (g2433) & (g2442) & (!g2460) & (g2478)) + ((g1879) & (g2433) & (g2442) & (g2460) & (!g2478)) + ((g1879) & (g2433) & (g2442) & (g2460) & (g2478)));
	assign g2531 = (((!g2075) & (!g2045) & (g2435) & (g2441)) + ((!g2075) & (g2045) & (!g2435) & (g2441)) + ((!g2075) & (g2045) & (g2435) & (!g2441)) + ((!g2075) & (g2045) & (g2435) & (g2441)) + ((g2075) & (!g2045) & (!g2435) & (!g2441)) + ((g2075) & (!g2045) & (!g2435) & (g2441)) + ((g2075) & (!g2045) & (g2435) & (!g2441)) + ((g2075) & (g2045) & (!g2435) & (!g2441)));
	assign g2532 = (((!g2434) & (!g2460) & (!g2478) & (g2531)) + ((!g2434) & (g2460) & (!g2478) & (g2531)) + ((!g2434) & (g2460) & (g2478) & (g2531)) + ((g2434) & (!g2460) & (!g2478) & (!g2531)) + ((g2434) & (!g2460) & (g2478) & (!g2531)) + ((g2434) & (!g2460) & (g2478) & (g2531)) + ((g2434) & (g2460) & (!g2478) & (!g2531)) + ((g2434) & (g2460) & (g2478) & (!g2531)));
	assign g2533 = (((!g2045) & (!g2435) & (g2441) & (!g2460) & (!g2478)) + ((!g2045) & (!g2435) & (g2441) & (g2460) & (!g2478)) + ((!g2045) & (!g2435) & (g2441) & (g2460) & (g2478)) + ((!g2045) & (g2435) & (!g2441) & (!g2460) & (!g2478)) + ((!g2045) & (g2435) & (!g2441) & (!g2460) & (g2478)) + ((!g2045) & (g2435) & (!g2441) & (g2460) & (!g2478)) + ((!g2045) & (g2435) & (!g2441) & (g2460) & (g2478)) + ((!g2045) & (g2435) & (g2441) & (!g2460) & (g2478)) + ((g2045) & (!g2435) & (!g2441) & (!g2460) & (!g2478)) + ((g2045) & (!g2435) & (!g2441) & (g2460) & (!g2478)) + ((g2045) & (!g2435) & (!g2441) & (g2460) & (g2478)) + ((g2045) & (g2435) & (!g2441) & (!g2460) & (g2478)) + ((g2045) & (g2435) & (g2441) & (!g2460) & (!g2478)) + ((g2045) & (g2435) & (g2441) & (!g2460) & (g2478)) + ((g2045) & (g2435) & (g2441) & (g2460) & (!g2478)) + ((g2045) & (g2435) & (g2441) & (g2460) & (g2478)));
	assign g2534 = (((!g2252) & (!g2218) & (g2438) & (g2440)) + ((!g2252) & (g2218) & (!g2438) & (g2440)) + ((!g2252) & (g2218) & (g2438) & (!g2440)) + ((!g2252) & (g2218) & (g2438) & (g2440)) + ((g2252) & (!g2218) & (!g2438) & (!g2440)) + ((g2252) & (!g2218) & (!g2438) & (g2440)) + ((g2252) & (!g2218) & (g2438) & (!g2440)) + ((g2252) & (g2218) & (!g2438) & (!g2440)));
	assign g2535 = (((!g2437) & (!g2460) & (!g2478) & (g2534)) + ((!g2437) & (g2460) & (!g2478) & (g2534)) + ((!g2437) & (g2460) & (g2478) & (g2534)) + ((g2437) & (!g2460) & (!g2478) & (!g2534)) + ((g2437) & (!g2460) & (g2478) & (!g2534)) + ((g2437) & (!g2460) & (g2478) & (g2534)) + ((g2437) & (g2460) & (!g2478) & (!g2534)) + ((g2437) & (g2460) & (g2478) & (!g2534)));
	assign g2536 = (((!g2218) & (!g2438) & (g2440) & (!g2460) & (!g2478)) + ((!g2218) & (!g2438) & (g2440) & (g2460) & (!g2478)) + ((!g2218) & (!g2438) & (g2440) & (g2460) & (g2478)) + ((!g2218) & (g2438) & (!g2440) & (!g2460) & (!g2478)) + ((!g2218) & (g2438) & (!g2440) & (!g2460) & (g2478)) + ((!g2218) & (g2438) & (!g2440) & (g2460) & (!g2478)) + ((!g2218) & (g2438) & (!g2440) & (g2460) & (g2478)) + ((!g2218) & (g2438) & (g2440) & (!g2460) & (g2478)) + ((g2218) & (!g2438) & (!g2440) & (!g2460) & (!g2478)) + ((g2218) & (!g2438) & (!g2440) & (g2460) & (!g2478)) + ((g2218) & (!g2438) & (!g2440) & (g2460) & (g2478)) + ((g2218) & (g2438) & (!g2440) & (!g2460) & (g2478)) + ((g2218) & (g2438) & (g2440) & (!g2460) & (!g2478)) + ((g2218) & (g2438) & (g2440) & (!g2460) & (g2478)) + ((g2218) & (g2438) & (g2440) & (g2460) & (!g2478)) + ((g2218) & (g2438) & (g2440) & (g2460) & (g2478)));
	assign g2537 = (((!g2436) & (!ax24x) & (!g2398) & (g2439)) + ((!g2436) & (!ax24x) & (g2398) & (g2439)) + ((!g2436) & (ax24x) & (!g2398) & (!g2439)) + ((!g2436) & (ax24x) & (!g2398) & (g2439)) + ((g2436) & (!ax24x) & (!g2398) & (!g2439)) + ((g2436) & (!ax24x) & (g2398) & (!g2439)) + ((g2436) & (ax24x) & (g2398) & (!g2439)) + ((g2436) & (ax24x) & (g2398) & (g2439)));
	assign g2538 = (((!ax24x) & (!ax25x) & (!g2398) & (!g2460) & (!g2478) & (g2537)) + ((!ax24x) & (!ax25x) & (!g2398) & (!g2460) & (g2478) & (!g2537)) + ((!ax24x) & (!ax25x) & (!g2398) & (!g2460) & (g2478) & (g2537)) + ((!ax24x) & (!ax25x) & (!g2398) & (g2460) & (!g2478) & (g2537)) + ((!ax24x) & (!ax25x) & (!g2398) & (g2460) & (g2478) & (g2537)) + ((!ax24x) & (!ax25x) & (g2398) & (!g2460) & (!g2478) & (!g2537)) + ((!ax24x) & (!ax25x) & (g2398) & (g2460) & (!g2478) & (!g2537)) + ((!ax24x) & (!ax25x) & (g2398) & (g2460) & (g2478) & (!g2537)) + ((!ax24x) & (ax25x) & (!g2398) & (!g2460) & (!g2478) & (!g2537)) + ((!ax24x) & (ax25x) & (!g2398) & (g2460) & (!g2478) & (!g2537)) + ((!ax24x) & (ax25x) & (!g2398) & (g2460) & (g2478) & (!g2537)) + ((!ax24x) & (ax25x) & (g2398) & (!g2460) & (!g2478) & (g2537)) + ((!ax24x) & (ax25x) & (g2398) & (!g2460) & (g2478) & (!g2537)) + ((!ax24x) & (ax25x) & (g2398) & (!g2460) & (g2478) & (g2537)) + ((!ax24x) & (ax25x) & (g2398) & (g2460) & (!g2478) & (g2537)) + ((!ax24x) & (ax25x) & (g2398) & (g2460) & (g2478) & (g2537)) + ((ax24x) & (!ax25x) & (!g2398) & (!g2460) & (!g2478) & (!g2537)) + ((ax24x) & (!ax25x) & (!g2398) & (g2460) & (!g2478) & (!g2537)) + ((ax24x) & (!ax25x) & (!g2398) & (g2460) & (g2478) & (!g2537)) + ((ax24x) & (!ax25x) & (g2398) & (!g2460) & (!g2478) & (!g2537)) + ((ax24x) & (!ax25x) & (g2398) & (g2460) & (!g2478) & (!g2537)) + ((ax24x) & (!ax25x) & (g2398) & (g2460) & (g2478) & (!g2537)) + ((ax24x) & (ax25x) & (!g2398) & (!g2460) & (!g2478) & (g2537)) + ((ax24x) & (ax25x) & (!g2398) & (!g2460) & (g2478) & (!g2537)) + ((ax24x) & (ax25x) & (!g2398) & (!g2460) & (g2478) & (g2537)) + ((ax24x) & (ax25x) & (!g2398) & (g2460) & (!g2478) & (g2537)) + ((ax24x) & (ax25x) & (!g2398) & (g2460) & (g2478) & (g2537)) + ((ax24x) & (ax25x) & (g2398) & (!g2460) & (!g2478) & (g2537)) + ((ax24x) & (ax25x) & (g2398) & (!g2460) & (g2478) & (!g2537)) + ((ax24x) & (ax25x) & (g2398) & (!g2460) & (g2478) & (g2537)) + ((ax24x) & (ax25x) & (g2398) & (g2460) & (!g2478) & (g2537)) + ((ax24x) & (ax25x) & (g2398) & (g2460) & (g2478) & (g2537)));
	assign g2539 = (((!ax24x) & (!g2398) & (!g2439) & (!g2460) & (g2478)) + ((!ax24x) & (!g2398) & (g2439) & (!g2460) & (!g2478)) + ((!ax24x) & (!g2398) & (g2439) & (!g2460) & (g2478)) + ((!ax24x) & (!g2398) & (g2439) & (g2460) & (!g2478)) + ((!ax24x) & (!g2398) & (g2439) & (g2460) & (g2478)) + ((!ax24x) & (g2398) & (g2439) & (!g2460) & (!g2478)) + ((!ax24x) & (g2398) & (g2439) & (g2460) & (!g2478)) + ((!ax24x) & (g2398) & (g2439) & (g2460) & (g2478)) + ((ax24x) & (!g2398) & (!g2439) & (!g2460) & (!g2478)) + ((ax24x) & (!g2398) & (!g2439) & (g2460) & (!g2478)) + ((ax24x) & (!g2398) & (!g2439) & (g2460) & (g2478)) + ((ax24x) & (g2398) & (!g2439) & (!g2460) & (!g2478)) + ((ax24x) & (g2398) & (!g2439) & (!g2460) & (g2478)) + ((ax24x) & (g2398) & (!g2439) & (g2460) & (!g2478)) + ((ax24x) & (g2398) & (!g2439) & (g2460) & (g2478)) + ((ax24x) & (g2398) & (g2439) & (!g2460) & (g2478)));
	assign g2540 = (((!ax20x) & (!ax21x)));
	assign g2541 = (((!g2398) & (!ax22x) & (!ax23x) & (!g2460) & (!g2478) & (!g2540)) + ((!g2398) & (!ax22x) & (!ax23x) & (g2460) & (!g2478) & (!g2540)) + ((!g2398) & (!ax22x) & (!ax23x) & (g2460) & (g2478) & (!g2540)) + ((!g2398) & (!ax22x) & (ax23x) & (!g2460) & (g2478) & (!g2540)) + ((!g2398) & (ax22x) & (ax23x) & (!g2460) & (g2478) & (!g2540)) + ((!g2398) & (ax22x) & (ax23x) & (!g2460) & (g2478) & (g2540)) + ((g2398) & (!ax22x) & (!ax23x) & (!g2460) & (!g2478) & (!g2540)) + ((g2398) & (!ax22x) & (!ax23x) & (!g2460) & (!g2478) & (g2540)) + ((g2398) & (!ax22x) & (!ax23x) & (!g2460) & (g2478) & (!g2540)) + ((g2398) & (!ax22x) & (!ax23x) & (g2460) & (!g2478) & (!g2540)) + ((g2398) & (!ax22x) & (!ax23x) & (g2460) & (!g2478) & (g2540)) + ((g2398) & (!ax22x) & (!ax23x) & (g2460) & (g2478) & (!g2540)) + ((g2398) & (!ax22x) & (!ax23x) & (g2460) & (g2478) & (g2540)) + ((g2398) & (!ax22x) & (ax23x) & (!g2460) & (!g2478) & (!g2540)) + ((g2398) & (!ax22x) & (ax23x) & (!g2460) & (g2478) & (!g2540)) + ((g2398) & (!ax22x) & (ax23x) & (!g2460) & (g2478) & (g2540)) + ((g2398) & (!ax22x) & (ax23x) & (g2460) & (!g2478) & (!g2540)) + ((g2398) & (!ax22x) & (ax23x) & (g2460) & (g2478) & (!g2540)) + ((g2398) & (ax22x) & (!ax23x) & (!g2460) & (g2478) & (!g2540)) + ((g2398) & (ax22x) & (!ax23x) & (!g2460) & (g2478) & (g2540)) + ((g2398) & (ax22x) & (ax23x) & (!g2460) & (!g2478) & (!g2540)) + ((g2398) & (ax22x) & (ax23x) & (!g2460) & (!g2478) & (g2540)) + ((g2398) & (ax22x) & (ax23x) & (!g2460) & (g2478) & (!g2540)) + ((g2398) & (ax22x) & (ax23x) & (!g2460) & (g2478) & (g2540)) + ((g2398) & (ax22x) & (ax23x) & (g2460) & (!g2478) & (!g2540)) + ((g2398) & (ax22x) & (ax23x) & (g2460) & (!g2478) & (g2540)) + ((g2398) & (ax22x) & (ax23x) & (g2460) & (g2478) & (!g2540)) + ((g2398) & (ax22x) & (ax23x) & (g2460) & (g2478) & (g2540)));
	assign g2542 = (((!g2218) & (!g2436) & (g2538) & (g2539) & (g2541)) + ((!g2218) & (g2436) & (g2538) & (!g2539) & (g2541)) + ((!g2218) & (g2436) & (g2538) & (g2539) & (!g2541)) + ((!g2218) & (g2436) & (g2538) & (g2539) & (g2541)) + ((g2218) & (!g2436) & (!g2538) & (g2539) & (g2541)) + ((g2218) & (!g2436) & (g2538) & (!g2539) & (!g2541)) + ((g2218) & (!g2436) & (g2538) & (!g2539) & (g2541)) + ((g2218) & (!g2436) & (g2538) & (g2539) & (!g2541)) + ((g2218) & (!g2436) & (g2538) & (g2539) & (g2541)) + ((g2218) & (g2436) & (!g2538) & (!g2539) & (g2541)) + ((g2218) & (g2436) & (!g2538) & (g2539) & (!g2541)) + ((g2218) & (g2436) & (!g2538) & (g2539) & (g2541)) + ((g2218) & (g2436) & (g2538) & (!g2539) & (!g2541)) + ((g2218) & (g2436) & (g2538) & (!g2539) & (g2541)) + ((g2218) & (g2436) & (g2538) & (g2539) & (!g2541)) + ((g2218) & (g2436) & (g2538) & (g2539) & (g2541)));
	assign g2543 = (((!g2045) & (!g2252) & (g2535) & (g2536) & (g2542)) + ((!g2045) & (g2252) & (g2535) & (!g2536) & (g2542)) + ((!g2045) & (g2252) & (g2535) & (g2536) & (!g2542)) + ((!g2045) & (g2252) & (g2535) & (g2536) & (g2542)) + ((g2045) & (!g2252) & (!g2535) & (g2536) & (g2542)) + ((g2045) & (!g2252) & (g2535) & (!g2536) & (!g2542)) + ((g2045) & (!g2252) & (g2535) & (!g2536) & (g2542)) + ((g2045) & (!g2252) & (g2535) & (g2536) & (!g2542)) + ((g2045) & (!g2252) & (g2535) & (g2536) & (g2542)) + ((g2045) & (g2252) & (!g2535) & (!g2536) & (g2542)) + ((g2045) & (g2252) & (!g2535) & (g2536) & (!g2542)) + ((g2045) & (g2252) & (!g2535) & (g2536) & (g2542)) + ((g2045) & (g2252) & (g2535) & (!g2536) & (!g2542)) + ((g2045) & (g2252) & (g2535) & (!g2536) & (g2542)) + ((g2045) & (g2252) & (g2535) & (g2536) & (!g2542)) + ((g2045) & (g2252) & (g2535) & (g2536) & (g2542)));
	assign g2544 = (((!g1879) & (!g2075) & (g2532) & (g2533) & (g2543)) + ((!g1879) & (g2075) & (g2532) & (!g2533) & (g2543)) + ((!g1879) & (g2075) & (g2532) & (g2533) & (!g2543)) + ((!g1879) & (g2075) & (g2532) & (g2533) & (g2543)) + ((g1879) & (!g2075) & (!g2532) & (g2533) & (g2543)) + ((g1879) & (!g2075) & (g2532) & (!g2533) & (!g2543)) + ((g1879) & (!g2075) & (g2532) & (!g2533) & (g2543)) + ((g1879) & (!g2075) & (g2532) & (g2533) & (!g2543)) + ((g1879) & (!g2075) & (g2532) & (g2533) & (g2543)) + ((g1879) & (g2075) & (!g2532) & (!g2533) & (g2543)) + ((g1879) & (g2075) & (!g2532) & (g2533) & (!g2543)) + ((g1879) & (g2075) & (!g2532) & (g2533) & (g2543)) + ((g1879) & (g2075) & (g2532) & (!g2533) & (!g2543)) + ((g1879) & (g2075) & (g2532) & (!g2533) & (g2543)) + ((g1879) & (g2075) & (g2532) & (g2533) & (!g2543)) + ((g1879) & (g2075) & (g2532) & (g2533) & (g2543)));
	assign g2545 = (((!g1720) & (!g1905) & (g2529) & (g2530) & (g2544)) + ((!g1720) & (g1905) & (g2529) & (!g2530) & (g2544)) + ((!g1720) & (g1905) & (g2529) & (g2530) & (!g2544)) + ((!g1720) & (g1905) & (g2529) & (g2530) & (g2544)) + ((g1720) & (!g1905) & (!g2529) & (g2530) & (g2544)) + ((g1720) & (!g1905) & (g2529) & (!g2530) & (!g2544)) + ((g1720) & (!g1905) & (g2529) & (!g2530) & (g2544)) + ((g1720) & (!g1905) & (g2529) & (g2530) & (!g2544)) + ((g1720) & (!g1905) & (g2529) & (g2530) & (g2544)) + ((g1720) & (g1905) & (!g2529) & (!g2530) & (g2544)) + ((g1720) & (g1905) & (!g2529) & (g2530) & (!g2544)) + ((g1720) & (g1905) & (!g2529) & (g2530) & (g2544)) + ((g1720) & (g1905) & (g2529) & (!g2530) & (!g2544)) + ((g1720) & (g1905) & (g2529) & (!g2530) & (g2544)) + ((g1720) & (g1905) & (g2529) & (g2530) & (!g2544)) + ((g1720) & (g1905) & (g2529) & (g2530) & (g2544)));
	assign g2546 = (((!g1568) & (!g1742) & (g2526) & (g2527) & (g2545)) + ((!g1568) & (g1742) & (g2526) & (!g2527) & (g2545)) + ((!g1568) & (g1742) & (g2526) & (g2527) & (!g2545)) + ((!g1568) & (g1742) & (g2526) & (g2527) & (g2545)) + ((g1568) & (!g1742) & (!g2526) & (g2527) & (g2545)) + ((g1568) & (!g1742) & (g2526) & (!g2527) & (!g2545)) + ((g1568) & (!g1742) & (g2526) & (!g2527) & (g2545)) + ((g1568) & (!g1742) & (g2526) & (g2527) & (!g2545)) + ((g1568) & (!g1742) & (g2526) & (g2527) & (g2545)) + ((g1568) & (g1742) & (!g2526) & (!g2527) & (g2545)) + ((g1568) & (g1742) & (!g2526) & (g2527) & (!g2545)) + ((g1568) & (g1742) & (!g2526) & (g2527) & (g2545)) + ((g1568) & (g1742) & (g2526) & (!g2527) & (!g2545)) + ((g1568) & (g1742) & (g2526) & (!g2527) & (g2545)) + ((g1568) & (g1742) & (g2526) & (g2527) & (!g2545)) + ((g1568) & (g1742) & (g2526) & (g2527) & (g2545)));
	assign g2547 = (((!g1423) & (!g1586) & (g2523) & (g2524) & (g2546)) + ((!g1423) & (g1586) & (g2523) & (!g2524) & (g2546)) + ((!g1423) & (g1586) & (g2523) & (g2524) & (!g2546)) + ((!g1423) & (g1586) & (g2523) & (g2524) & (g2546)) + ((g1423) & (!g1586) & (!g2523) & (g2524) & (g2546)) + ((g1423) & (!g1586) & (g2523) & (!g2524) & (!g2546)) + ((g1423) & (!g1586) & (g2523) & (!g2524) & (g2546)) + ((g1423) & (!g1586) & (g2523) & (g2524) & (!g2546)) + ((g1423) & (!g1586) & (g2523) & (g2524) & (g2546)) + ((g1423) & (g1586) & (!g2523) & (!g2524) & (g2546)) + ((g1423) & (g1586) & (!g2523) & (g2524) & (!g2546)) + ((g1423) & (g1586) & (!g2523) & (g2524) & (g2546)) + ((g1423) & (g1586) & (g2523) & (!g2524) & (!g2546)) + ((g1423) & (g1586) & (g2523) & (!g2524) & (g2546)) + ((g1423) & (g1586) & (g2523) & (g2524) & (!g2546)) + ((g1423) & (g1586) & (g2523) & (g2524) & (g2546)));
	assign g2548 = (((!g1285) & (!g1437) & (g2520) & (g2521) & (g2547)) + ((!g1285) & (g1437) & (g2520) & (!g2521) & (g2547)) + ((!g1285) & (g1437) & (g2520) & (g2521) & (!g2547)) + ((!g1285) & (g1437) & (g2520) & (g2521) & (g2547)) + ((g1285) & (!g1437) & (!g2520) & (g2521) & (g2547)) + ((g1285) & (!g1437) & (g2520) & (!g2521) & (!g2547)) + ((g1285) & (!g1437) & (g2520) & (!g2521) & (g2547)) + ((g1285) & (!g1437) & (g2520) & (g2521) & (!g2547)) + ((g1285) & (!g1437) & (g2520) & (g2521) & (g2547)) + ((g1285) & (g1437) & (!g2520) & (!g2521) & (g2547)) + ((g1285) & (g1437) & (!g2520) & (g2521) & (!g2547)) + ((g1285) & (g1437) & (!g2520) & (g2521) & (g2547)) + ((g1285) & (g1437) & (g2520) & (!g2521) & (!g2547)) + ((g1285) & (g1437) & (g2520) & (!g2521) & (g2547)) + ((g1285) & (g1437) & (g2520) & (g2521) & (!g2547)) + ((g1285) & (g1437) & (g2520) & (g2521) & (g2547)));
	assign g2549 = (((!g1154) & (!g1295) & (g2517) & (g2518) & (g2548)) + ((!g1154) & (g1295) & (g2517) & (!g2518) & (g2548)) + ((!g1154) & (g1295) & (g2517) & (g2518) & (!g2548)) + ((!g1154) & (g1295) & (g2517) & (g2518) & (g2548)) + ((g1154) & (!g1295) & (!g2517) & (g2518) & (g2548)) + ((g1154) & (!g1295) & (g2517) & (!g2518) & (!g2548)) + ((g1154) & (!g1295) & (g2517) & (!g2518) & (g2548)) + ((g1154) & (!g1295) & (g2517) & (g2518) & (!g2548)) + ((g1154) & (!g1295) & (g2517) & (g2518) & (g2548)) + ((g1154) & (g1295) & (!g2517) & (!g2518) & (g2548)) + ((g1154) & (g1295) & (!g2517) & (g2518) & (!g2548)) + ((g1154) & (g1295) & (!g2517) & (g2518) & (g2548)) + ((g1154) & (g1295) & (g2517) & (!g2518) & (!g2548)) + ((g1154) & (g1295) & (g2517) & (!g2518) & (g2548)) + ((g1154) & (g1295) & (g2517) & (g2518) & (!g2548)) + ((g1154) & (g1295) & (g2517) & (g2518) & (g2548)));
	assign g2550 = (((!g1030) & (!g1160) & (g2514) & (g2515) & (g2549)) + ((!g1030) & (g1160) & (g2514) & (!g2515) & (g2549)) + ((!g1030) & (g1160) & (g2514) & (g2515) & (!g2549)) + ((!g1030) & (g1160) & (g2514) & (g2515) & (g2549)) + ((g1030) & (!g1160) & (!g2514) & (g2515) & (g2549)) + ((g1030) & (!g1160) & (g2514) & (!g2515) & (!g2549)) + ((g1030) & (!g1160) & (g2514) & (!g2515) & (g2549)) + ((g1030) & (!g1160) & (g2514) & (g2515) & (!g2549)) + ((g1030) & (!g1160) & (g2514) & (g2515) & (g2549)) + ((g1030) & (g1160) & (!g2514) & (!g2515) & (g2549)) + ((g1030) & (g1160) & (!g2514) & (g2515) & (!g2549)) + ((g1030) & (g1160) & (!g2514) & (g2515) & (g2549)) + ((g1030) & (g1160) & (g2514) & (!g2515) & (!g2549)) + ((g1030) & (g1160) & (g2514) & (!g2515) & (g2549)) + ((g1030) & (g1160) & (g2514) & (g2515) & (!g2549)) + ((g1030) & (g1160) & (g2514) & (g2515) & (g2549)));
	assign g2551 = (((!g914) & (!g1032) & (g2511) & (g2512) & (g2550)) + ((!g914) & (g1032) & (g2511) & (!g2512) & (g2550)) + ((!g914) & (g1032) & (g2511) & (g2512) & (!g2550)) + ((!g914) & (g1032) & (g2511) & (g2512) & (g2550)) + ((g914) & (!g1032) & (!g2511) & (g2512) & (g2550)) + ((g914) & (!g1032) & (g2511) & (!g2512) & (!g2550)) + ((g914) & (!g1032) & (g2511) & (!g2512) & (g2550)) + ((g914) & (!g1032) & (g2511) & (g2512) & (!g2550)) + ((g914) & (!g1032) & (g2511) & (g2512) & (g2550)) + ((g914) & (g1032) & (!g2511) & (!g2512) & (g2550)) + ((g914) & (g1032) & (!g2511) & (g2512) & (!g2550)) + ((g914) & (g1032) & (!g2511) & (g2512) & (g2550)) + ((g914) & (g1032) & (g2511) & (!g2512) & (!g2550)) + ((g914) & (g1032) & (g2511) & (!g2512) & (g2550)) + ((g914) & (g1032) & (g2511) & (g2512) & (!g2550)) + ((g914) & (g1032) & (g2511) & (g2512) & (g2550)));
	assign g2552 = (((!g803) & (!g851) & (g2508) & (g2509) & (g2551)) + ((!g803) & (g851) & (g2508) & (!g2509) & (g2551)) + ((!g803) & (g851) & (g2508) & (g2509) & (!g2551)) + ((!g803) & (g851) & (g2508) & (g2509) & (g2551)) + ((g803) & (!g851) & (!g2508) & (g2509) & (g2551)) + ((g803) & (!g851) & (g2508) & (!g2509) & (!g2551)) + ((g803) & (!g851) & (g2508) & (!g2509) & (g2551)) + ((g803) & (!g851) & (g2508) & (g2509) & (!g2551)) + ((g803) & (!g851) & (g2508) & (g2509) & (g2551)) + ((g803) & (g851) & (!g2508) & (!g2509) & (g2551)) + ((g803) & (g851) & (!g2508) & (g2509) & (!g2551)) + ((g803) & (g851) & (!g2508) & (g2509) & (g2551)) + ((g803) & (g851) & (g2508) & (!g2509) & (!g2551)) + ((g803) & (g851) & (g2508) & (!g2509) & (g2551)) + ((g803) & (g851) & (g2508) & (g2509) & (!g2551)) + ((g803) & (g851) & (g2508) & (g2509) & (g2551)));
	assign g2553 = (((!g700) & (!g744) & (g2505) & (g2506) & (g2552)) + ((!g700) & (g744) & (g2505) & (!g2506) & (g2552)) + ((!g700) & (g744) & (g2505) & (g2506) & (!g2552)) + ((!g700) & (g744) & (g2505) & (g2506) & (g2552)) + ((g700) & (!g744) & (!g2505) & (g2506) & (g2552)) + ((g700) & (!g744) & (g2505) & (!g2506) & (!g2552)) + ((g700) & (!g744) & (g2505) & (!g2506) & (g2552)) + ((g700) & (!g744) & (g2505) & (g2506) & (!g2552)) + ((g700) & (!g744) & (g2505) & (g2506) & (g2552)) + ((g700) & (g744) & (!g2505) & (!g2506) & (g2552)) + ((g700) & (g744) & (!g2505) & (g2506) & (!g2552)) + ((g700) & (g744) & (!g2505) & (g2506) & (g2552)) + ((g700) & (g744) & (g2505) & (!g2506) & (!g2552)) + ((g700) & (g744) & (g2505) & (!g2506) & (g2552)) + ((g700) & (g744) & (g2505) & (g2506) & (!g2552)) + ((g700) & (g744) & (g2505) & (g2506) & (g2552)));
	assign g2554 = (((!g604) & (!g645) & (g2502) & (g2503) & (g2553)) + ((!g604) & (g645) & (g2502) & (!g2503) & (g2553)) + ((!g604) & (g645) & (g2502) & (g2503) & (!g2553)) + ((!g604) & (g645) & (g2502) & (g2503) & (g2553)) + ((g604) & (!g645) & (!g2502) & (g2503) & (g2553)) + ((g604) & (!g645) & (g2502) & (!g2503) & (!g2553)) + ((g604) & (!g645) & (g2502) & (!g2503) & (g2553)) + ((g604) & (!g645) & (g2502) & (g2503) & (!g2553)) + ((g604) & (!g645) & (g2502) & (g2503) & (g2553)) + ((g604) & (g645) & (!g2502) & (!g2503) & (g2553)) + ((g604) & (g645) & (!g2502) & (g2503) & (!g2553)) + ((g604) & (g645) & (!g2502) & (g2503) & (g2553)) + ((g604) & (g645) & (g2502) & (!g2503) & (!g2553)) + ((g604) & (g645) & (g2502) & (!g2503) & (g2553)) + ((g604) & (g645) & (g2502) & (g2503) & (!g2553)) + ((g604) & (g645) & (g2502) & (g2503) & (g2553)));
	assign g2555 = (((!g515) & (!g553) & (g2499) & (g2500) & (g2554)) + ((!g515) & (g553) & (g2499) & (!g2500) & (g2554)) + ((!g515) & (g553) & (g2499) & (g2500) & (!g2554)) + ((!g515) & (g553) & (g2499) & (g2500) & (g2554)) + ((g515) & (!g553) & (!g2499) & (g2500) & (g2554)) + ((g515) & (!g553) & (g2499) & (!g2500) & (!g2554)) + ((g515) & (!g553) & (g2499) & (!g2500) & (g2554)) + ((g515) & (!g553) & (g2499) & (g2500) & (!g2554)) + ((g515) & (!g553) & (g2499) & (g2500) & (g2554)) + ((g515) & (g553) & (!g2499) & (!g2500) & (g2554)) + ((g515) & (g553) & (!g2499) & (g2500) & (!g2554)) + ((g515) & (g553) & (!g2499) & (g2500) & (g2554)) + ((g515) & (g553) & (g2499) & (!g2500) & (!g2554)) + ((g515) & (g553) & (g2499) & (!g2500) & (g2554)) + ((g515) & (g553) & (g2499) & (g2500) & (!g2554)) + ((g515) & (g553) & (g2499) & (g2500) & (g2554)));
	assign g2556 = (((!g433) & (!g468) & (g2496) & (g2497) & (g2555)) + ((!g433) & (g468) & (g2496) & (!g2497) & (g2555)) + ((!g433) & (g468) & (g2496) & (g2497) & (!g2555)) + ((!g433) & (g468) & (g2496) & (g2497) & (g2555)) + ((g433) & (!g468) & (!g2496) & (g2497) & (g2555)) + ((g433) & (!g468) & (g2496) & (!g2497) & (!g2555)) + ((g433) & (!g468) & (g2496) & (!g2497) & (g2555)) + ((g433) & (!g468) & (g2496) & (g2497) & (!g2555)) + ((g433) & (!g468) & (g2496) & (g2497) & (g2555)) + ((g433) & (g468) & (!g2496) & (!g2497) & (g2555)) + ((g433) & (g468) & (!g2496) & (g2497) & (!g2555)) + ((g433) & (g468) & (!g2496) & (g2497) & (g2555)) + ((g433) & (g468) & (g2496) & (!g2497) & (!g2555)) + ((g433) & (g468) & (g2496) & (!g2497) & (g2555)) + ((g433) & (g468) & (g2496) & (g2497) & (!g2555)) + ((g433) & (g468) & (g2496) & (g2497) & (g2555)));
	assign g2557 = (((!g358) & (!g390) & (g2493) & (g2494) & (g2556)) + ((!g358) & (g390) & (g2493) & (!g2494) & (g2556)) + ((!g358) & (g390) & (g2493) & (g2494) & (!g2556)) + ((!g358) & (g390) & (g2493) & (g2494) & (g2556)) + ((g358) & (!g390) & (!g2493) & (g2494) & (g2556)) + ((g358) & (!g390) & (g2493) & (!g2494) & (!g2556)) + ((g358) & (!g390) & (g2493) & (!g2494) & (g2556)) + ((g358) & (!g390) & (g2493) & (g2494) & (!g2556)) + ((g358) & (!g390) & (g2493) & (g2494) & (g2556)) + ((g358) & (g390) & (!g2493) & (!g2494) & (g2556)) + ((g358) & (g390) & (!g2493) & (g2494) & (!g2556)) + ((g358) & (g390) & (!g2493) & (g2494) & (g2556)) + ((g358) & (g390) & (g2493) & (!g2494) & (!g2556)) + ((g358) & (g390) & (g2493) & (!g2494) & (g2556)) + ((g358) & (g390) & (g2493) & (g2494) & (!g2556)) + ((g358) & (g390) & (g2493) & (g2494) & (g2556)));
	assign g2558 = (((!g290) & (!g319) & (g2490) & (g2491) & (g2557)) + ((!g290) & (g319) & (g2490) & (!g2491) & (g2557)) + ((!g290) & (g319) & (g2490) & (g2491) & (!g2557)) + ((!g290) & (g319) & (g2490) & (g2491) & (g2557)) + ((g290) & (!g319) & (!g2490) & (g2491) & (g2557)) + ((g290) & (!g319) & (g2490) & (!g2491) & (!g2557)) + ((g290) & (!g319) & (g2490) & (!g2491) & (g2557)) + ((g290) & (!g319) & (g2490) & (g2491) & (!g2557)) + ((g290) & (!g319) & (g2490) & (g2491) & (g2557)) + ((g290) & (g319) & (!g2490) & (!g2491) & (g2557)) + ((g290) & (g319) & (!g2490) & (g2491) & (!g2557)) + ((g290) & (g319) & (!g2490) & (g2491) & (g2557)) + ((g290) & (g319) & (g2490) & (!g2491) & (!g2557)) + ((g290) & (g319) & (g2490) & (!g2491) & (g2557)) + ((g290) & (g319) & (g2490) & (g2491) & (!g2557)) + ((g290) & (g319) & (g2490) & (g2491) & (g2557)));
	assign g2559 = (((!g229) & (!g255) & (g2487) & (g2488) & (g2558)) + ((!g229) & (g255) & (g2487) & (!g2488) & (g2558)) + ((!g229) & (g255) & (g2487) & (g2488) & (!g2558)) + ((!g229) & (g255) & (g2487) & (g2488) & (g2558)) + ((g229) & (!g255) & (!g2487) & (g2488) & (g2558)) + ((g229) & (!g255) & (g2487) & (!g2488) & (!g2558)) + ((g229) & (!g255) & (g2487) & (!g2488) & (g2558)) + ((g229) & (!g255) & (g2487) & (g2488) & (!g2558)) + ((g229) & (!g255) & (g2487) & (g2488) & (g2558)) + ((g229) & (g255) & (!g2487) & (!g2488) & (g2558)) + ((g229) & (g255) & (!g2487) & (g2488) & (!g2558)) + ((g229) & (g255) & (!g2487) & (g2488) & (g2558)) + ((g229) & (g255) & (g2487) & (!g2488) & (!g2558)) + ((g229) & (g255) & (g2487) & (!g2488) & (g2558)) + ((g229) & (g255) & (g2487) & (g2488) & (!g2558)) + ((g229) & (g255) & (g2487) & (g2488) & (g2558)));
	assign g2560 = (((!g174) & (!g198) & (g2484) & (g2485) & (g2559)) + ((!g174) & (g198) & (g2484) & (!g2485) & (g2559)) + ((!g174) & (g198) & (g2484) & (g2485) & (!g2559)) + ((!g174) & (g198) & (g2484) & (g2485) & (g2559)) + ((g174) & (!g198) & (!g2484) & (g2485) & (g2559)) + ((g174) & (!g198) & (g2484) & (!g2485) & (!g2559)) + ((g174) & (!g198) & (g2484) & (!g2485) & (g2559)) + ((g174) & (!g198) & (g2484) & (g2485) & (!g2559)) + ((g174) & (!g198) & (g2484) & (g2485) & (g2559)) + ((g174) & (g198) & (!g2484) & (!g2485) & (g2559)) + ((g174) & (g198) & (!g2484) & (g2485) & (!g2559)) + ((g174) & (g198) & (!g2484) & (g2485) & (g2559)) + ((g174) & (g198) & (g2484) & (!g2485) & (!g2559)) + ((g174) & (g198) & (g2484) & (!g2485) & (g2559)) + ((g174) & (g198) & (g2484) & (g2485) & (!g2559)) + ((g174) & (g198) & (g2484) & (g2485) & (g2559)));
	assign g2561 = (((!g127) & (!g147) & (g2481) & (g2482) & (g2560)) + ((!g127) & (g147) & (g2481) & (!g2482) & (g2560)) + ((!g127) & (g147) & (g2481) & (g2482) & (!g2560)) + ((!g127) & (g147) & (g2481) & (g2482) & (g2560)) + ((g127) & (!g147) & (!g2481) & (g2482) & (g2560)) + ((g127) & (!g147) & (g2481) & (!g2482) & (!g2560)) + ((g127) & (!g147) & (g2481) & (!g2482) & (g2560)) + ((g127) & (!g147) & (g2481) & (g2482) & (!g2560)) + ((g127) & (!g147) & (g2481) & (g2482) & (g2560)) + ((g127) & (g147) & (!g2481) & (!g2482) & (g2560)) + ((g127) & (g147) & (!g2481) & (g2482) & (!g2560)) + ((g127) & (g147) & (!g2481) & (g2482) & (g2560)) + ((g127) & (g147) & (g2481) & (!g2482) & (!g2560)) + ((g127) & (g147) & (g2481) & (!g2482) & (g2560)) + ((g127) & (g147) & (g2481) & (g2482) & (!g2560)) + ((g127) & (g147) & (g2481) & (g2482) & (g2560)));
	assign g2562 = (((!g4) & (!g2475) & (!g2476) & (!g2460) & (!g2478)) + ((!g4) & (!g2475) & (!g2476) & (g2460) & (!g2478)) + ((!g4) & (!g2475) & (!g2476) & (g2460) & (g2478)) + ((!g4) & (!g2475) & (g2476) & (!g2460) & (g2478)) + ((!g4) & (g2475) & (g2476) & (!g2460) & (!g2478)) + ((!g4) & (g2475) & (g2476) & (!g2460) & (g2478)) + ((!g4) & (g2475) & (g2476) & (g2460) & (!g2478)) + ((!g4) & (g2475) & (g2476) & (g2460) & (g2478)) + ((g4) & (!g2475) & (g2476) & (!g2460) & (!g2478)) + ((g4) & (!g2475) & (g2476) & (!g2460) & (g2478)) + ((g4) & (!g2475) & (g2476) & (g2460) & (!g2478)) + ((g4) & (!g2475) & (g2476) & (g2460) & (g2478)) + ((g4) & (g2475) & (!g2476) & (!g2460) & (!g2478)) + ((g4) & (g2475) & (!g2476) & (g2460) & (!g2478)) + ((g4) & (g2475) & (!g2476) & (g2460) & (g2478)) + ((g4) & (g2475) & (g2476) & (!g2460) & (g2478)));
	assign g2563 = (((!g8) & (!g2463) & (g2474) & (!g2460) & (!g2478)) + ((!g8) & (!g2463) & (g2474) & (g2460) & (!g2478)) + ((!g8) & (!g2463) & (g2474) & (g2460) & (g2478)) + ((!g8) & (g2463) & (!g2474) & (!g2460) & (!g2478)) + ((!g8) & (g2463) & (!g2474) & (!g2460) & (g2478)) + ((!g8) & (g2463) & (!g2474) & (g2460) & (!g2478)) + ((!g8) & (g2463) & (!g2474) & (g2460) & (g2478)) + ((!g8) & (g2463) & (g2474) & (!g2460) & (g2478)) + ((g8) & (!g2463) & (!g2474) & (!g2460) & (!g2478)) + ((g8) & (!g2463) & (!g2474) & (g2460) & (!g2478)) + ((g8) & (!g2463) & (!g2474) & (g2460) & (g2478)) + ((g8) & (g2463) & (!g2474) & (!g2460) & (g2478)) + ((g8) & (g2463) & (g2474) & (!g2460) & (!g2478)) + ((g8) & (g2463) & (g2474) & (!g2460) & (g2478)) + ((g8) & (g2463) & (g2474) & (g2460) & (!g2478)) + ((g8) & (g2463) & (g2474) & (g2460) & (g2478)));
	assign g2564 = (((!g18) & (!g27) & (g2465) & (g2473)) + ((!g18) & (g27) & (!g2465) & (g2473)) + ((!g18) & (g27) & (g2465) & (!g2473)) + ((!g18) & (g27) & (g2465) & (g2473)) + ((g18) & (!g27) & (!g2465) & (!g2473)) + ((g18) & (!g27) & (!g2465) & (g2473)) + ((g18) & (!g27) & (g2465) & (!g2473)) + ((g18) & (g27) & (!g2465) & (!g2473)));
	assign g2565 = (((!g2464) & (!g2460) & (!g2478) & (g2564)) + ((!g2464) & (g2460) & (!g2478) & (g2564)) + ((!g2464) & (g2460) & (g2478) & (g2564)) + ((g2464) & (!g2460) & (!g2478) & (!g2564)) + ((g2464) & (!g2460) & (g2478) & (!g2564)) + ((g2464) & (!g2460) & (g2478) & (g2564)) + ((g2464) & (g2460) & (!g2478) & (!g2564)) + ((g2464) & (g2460) & (g2478) & (!g2564)));
	assign g2566 = (((!g27) & (!g2465) & (g2473) & (!g2460) & (!g2478)) + ((!g27) & (!g2465) & (g2473) & (g2460) & (!g2478)) + ((!g27) & (!g2465) & (g2473) & (g2460) & (g2478)) + ((!g27) & (g2465) & (!g2473) & (!g2460) & (!g2478)) + ((!g27) & (g2465) & (!g2473) & (!g2460) & (g2478)) + ((!g27) & (g2465) & (!g2473) & (g2460) & (!g2478)) + ((!g27) & (g2465) & (!g2473) & (g2460) & (g2478)) + ((!g27) & (g2465) & (g2473) & (!g2460) & (g2478)) + ((g27) & (!g2465) & (!g2473) & (!g2460) & (!g2478)) + ((g27) & (!g2465) & (!g2473) & (g2460) & (!g2478)) + ((g27) & (!g2465) & (!g2473) & (g2460) & (g2478)) + ((g27) & (g2465) & (!g2473) & (!g2460) & (g2478)) + ((g27) & (g2465) & (g2473) & (!g2460) & (!g2478)) + ((g27) & (g2465) & (g2473) & (!g2460) & (g2478)) + ((g27) & (g2465) & (g2473) & (g2460) & (!g2478)) + ((g27) & (g2465) & (g2473) & (g2460) & (g2478)));
	assign g2567 = (((!g39) & (!g54) & (g2467) & (g2472)) + ((!g39) & (g54) & (!g2467) & (g2472)) + ((!g39) & (g54) & (g2467) & (!g2472)) + ((!g39) & (g54) & (g2467) & (g2472)) + ((g39) & (!g54) & (!g2467) & (!g2472)) + ((g39) & (!g54) & (!g2467) & (g2472)) + ((g39) & (!g54) & (g2467) & (!g2472)) + ((g39) & (g54) & (!g2467) & (!g2472)));
	assign g2568 = (((!g2466) & (!g2460) & (!g2478) & (g2567)) + ((!g2466) & (g2460) & (!g2478) & (g2567)) + ((!g2466) & (g2460) & (g2478) & (g2567)) + ((g2466) & (!g2460) & (!g2478) & (!g2567)) + ((g2466) & (!g2460) & (g2478) & (!g2567)) + ((g2466) & (!g2460) & (g2478) & (g2567)) + ((g2466) & (g2460) & (!g2478) & (!g2567)) + ((g2466) & (g2460) & (g2478) & (!g2567)));
	assign g2569 = (((!g54) & (!g2467) & (g2472) & (!g2460) & (!g2478)) + ((!g54) & (!g2467) & (g2472) & (g2460) & (!g2478)) + ((!g54) & (!g2467) & (g2472) & (g2460) & (g2478)) + ((!g54) & (g2467) & (!g2472) & (!g2460) & (!g2478)) + ((!g54) & (g2467) & (!g2472) & (!g2460) & (g2478)) + ((!g54) & (g2467) & (!g2472) & (g2460) & (!g2478)) + ((!g54) & (g2467) & (!g2472) & (g2460) & (g2478)) + ((!g54) & (g2467) & (g2472) & (!g2460) & (g2478)) + ((g54) & (!g2467) & (!g2472) & (!g2460) & (!g2478)) + ((g54) & (!g2467) & (!g2472) & (g2460) & (!g2478)) + ((g54) & (!g2467) & (!g2472) & (g2460) & (g2478)) + ((g54) & (g2467) & (!g2472) & (!g2460) & (g2478)) + ((g54) & (g2467) & (g2472) & (!g2460) & (!g2478)) + ((g54) & (g2467) & (g2472) & (!g2460) & (g2478)) + ((g54) & (g2467) & (g2472) & (g2460) & (!g2478)) + ((g54) & (g2467) & (g2472) & (g2460) & (g2478)));
	assign g2570 = (((!g68) & (!g87) & (g2469) & (g2471)) + ((!g68) & (g87) & (!g2469) & (g2471)) + ((!g68) & (g87) & (g2469) & (!g2471)) + ((!g68) & (g87) & (g2469) & (g2471)) + ((g68) & (!g87) & (!g2469) & (!g2471)) + ((g68) & (!g87) & (!g2469) & (g2471)) + ((g68) & (!g87) & (g2469) & (!g2471)) + ((g68) & (g87) & (!g2469) & (!g2471)));
	assign g2571 = (((!g2468) & (!g2460) & (!g2478) & (g2570)) + ((!g2468) & (g2460) & (!g2478) & (g2570)) + ((!g2468) & (g2460) & (g2478) & (g2570)) + ((g2468) & (!g2460) & (!g2478) & (!g2570)) + ((g2468) & (!g2460) & (g2478) & (!g2570)) + ((g2468) & (!g2460) & (g2478) & (g2570)) + ((g2468) & (g2460) & (!g2478) & (!g2570)) + ((g2468) & (g2460) & (g2478) & (!g2570)));
	assign g2572 = (((!g87) & (!g2469) & (g2471) & (!g2460) & (!g2478)) + ((!g87) & (!g2469) & (g2471) & (g2460) & (!g2478)) + ((!g87) & (!g2469) & (g2471) & (g2460) & (g2478)) + ((!g87) & (g2469) & (!g2471) & (!g2460) & (!g2478)) + ((!g87) & (g2469) & (!g2471) & (!g2460) & (g2478)) + ((!g87) & (g2469) & (!g2471) & (g2460) & (!g2478)) + ((!g87) & (g2469) & (!g2471) & (g2460) & (g2478)) + ((!g87) & (g2469) & (g2471) & (!g2460) & (g2478)) + ((g87) & (!g2469) & (!g2471) & (!g2460) & (!g2478)) + ((g87) & (!g2469) & (!g2471) & (g2460) & (!g2478)) + ((g87) & (!g2469) & (!g2471) & (g2460) & (g2478)) + ((g87) & (g2469) & (!g2471) & (!g2460) & (g2478)) + ((g87) & (g2469) & (g2471) & (!g2460) & (!g2478)) + ((g87) & (g2469) & (g2471) & (!g2460) & (g2478)) + ((g87) & (g2469) & (g2471) & (g2460) & (!g2478)) + ((g87) & (g2469) & (g2471) & (g2460) & (g2478)));
	assign g2573 = (((!g104) & (!g127) & (g2399) & (g2459)) + ((!g104) & (g127) & (!g2399) & (g2459)) + ((!g104) & (g127) & (g2399) & (!g2459)) + ((!g104) & (g127) & (g2399) & (g2459)) + ((g104) & (!g127) & (!g2399) & (!g2459)) + ((g104) & (!g127) & (!g2399) & (g2459)) + ((g104) & (!g127) & (g2399) & (!g2459)) + ((g104) & (g127) & (!g2399) & (!g2459)));
	assign g2574 = (((!g2470) & (!g2460) & (!g2478) & (g2573)) + ((!g2470) & (g2460) & (!g2478) & (g2573)) + ((!g2470) & (g2460) & (g2478) & (g2573)) + ((g2470) & (!g2460) & (!g2478) & (!g2573)) + ((g2470) & (!g2460) & (g2478) & (!g2573)) + ((g2470) & (!g2460) & (g2478) & (g2573)) + ((g2470) & (g2460) & (!g2478) & (!g2573)) + ((g2470) & (g2460) & (g2478) & (!g2573)));
	assign g2575 = (((!g87) & (!g104) & (g2574) & (g2479) & (g2561)) + ((!g87) & (g104) & (g2574) & (!g2479) & (g2561)) + ((!g87) & (g104) & (g2574) & (g2479) & (!g2561)) + ((!g87) & (g104) & (g2574) & (g2479) & (g2561)) + ((g87) & (!g104) & (!g2574) & (g2479) & (g2561)) + ((g87) & (!g104) & (g2574) & (!g2479) & (!g2561)) + ((g87) & (!g104) & (g2574) & (!g2479) & (g2561)) + ((g87) & (!g104) & (g2574) & (g2479) & (!g2561)) + ((g87) & (!g104) & (g2574) & (g2479) & (g2561)) + ((g87) & (g104) & (!g2574) & (!g2479) & (g2561)) + ((g87) & (g104) & (!g2574) & (g2479) & (!g2561)) + ((g87) & (g104) & (!g2574) & (g2479) & (g2561)) + ((g87) & (g104) & (g2574) & (!g2479) & (!g2561)) + ((g87) & (g104) & (g2574) & (!g2479) & (g2561)) + ((g87) & (g104) & (g2574) & (g2479) & (!g2561)) + ((g87) & (g104) & (g2574) & (g2479) & (g2561)));
	assign g2576 = (((!g54) & (!g68) & (g2571) & (g2572) & (g2575)) + ((!g54) & (g68) & (g2571) & (!g2572) & (g2575)) + ((!g54) & (g68) & (g2571) & (g2572) & (!g2575)) + ((!g54) & (g68) & (g2571) & (g2572) & (g2575)) + ((g54) & (!g68) & (!g2571) & (g2572) & (g2575)) + ((g54) & (!g68) & (g2571) & (!g2572) & (!g2575)) + ((g54) & (!g68) & (g2571) & (!g2572) & (g2575)) + ((g54) & (!g68) & (g2571) & (g2572) & (!g2575)) + ((g54) & (!g68) & (g2571) & (g2572) & (g2575)) + ((g54) & (g68) & (!g2571) & (!g2572) & (g2575)) + ((g54) & (g68) & (!g2571) & (g2572) & (!g2575)) + ((g54) & (g68) & (!g2571) & (g2572) & (g2575)) + ((g54) & (g68) & (g2571) & (!g2572) & (!g2575)) + ((g54) & (g68) & (g2571) & (!g2572) & (g2575)) + ((g54) & (g68) & (g2571) & (g2572) & (!g2575)) + ((g54) & (g68) & (g2571) & (g2572) & (g2575)));
	assign g2577 = (((!g27) & (!g39) & (g2568) & (g2569) & (g2576)) + ((!g27) & (g39) & (g2568) & (!g2569) & (g2576)) + ((!g27) & (g39) & (g2568) & (g2569) & (!g2576)) + ((!g27) & (g39) & (g2568) & (g2569) & (g2576)) + ((g27) & (!g39) & (!g2568) & (g2569) & (g2576)) + ((g27) & (!g39) & (g2568) & (!g2569) & (!g2576)) + ((g27) & (!g39) & (g2568) & (!g2569) & (g2576)) + ((g27) & (!g39) & (g2568) & (g2569) & (!g2576)) + ((g27) & (!g39) & (g2568) & (g2569) & (g2576)) + ((g27) & (g39) & (!g2568) & (!g2569) & (g2576)) + ((g27) & (g39) & (!g2568) & (g2569) & (!g2576)) + ((g27) & (g39) & (!g2568) & (g2569) & (g2576)) + ((g27) & (g39) & (g2568) & (!g2569) & (!g2576)) + ((g27) & (g39) & (g2568) & (!g2569) & (g2576)) + ((g27) & (g39) & (g2568) & (g2569) & (!g2576)) + ((g27) & (g39) & (g2568) & (g2569) & (g2576)));
	assign g2578 = (((!g8) & (!g18) & (g2565) & (g2566) & (g2577)) + ((!g8) & (g18) & (g2565) & (!g2566) & (g2577)) + ((!g8) & (g18) & (g2565) & (g2566) & (!g2577)) + ((!g8) & (g18) & (g2565) & (g2566) & (g2577)) + ((g8) & (!g18) & (!g2565) & (g2566) & (g2577)) + ((g8) & (!g18) & (g2565) & (!g2566) & (!g2577)) + ((g8) & (!g18) & (g2565) & (!g2566) & (g2577)) + ((g8) & (!g18) & (g2565) & (g2566) & (!g2577)) + ((g8) & (!g18) & (g2565) & (g2566) & (g2577)) + ((g8) & (g18) & (!g2565) & (!g2566) & (g2577)) + ((g8) & (g18) & (!g2565) & (g2566) & (!g2577)) + ((g8) & (g18) & (!g2565) & (g2566) & (g2577)) + ((g8) & (g18) & (g2565) & (!g2566) & (!g2577)) + ((g8) & (g18) & (g2565) & (!g2566) & (g2577)) + ((g8) & (g18) & (g2565) & (g2566) & (!g2577)) + ((g8) & (g18) & (g2565) & (g2566) & (g2577)));
	assign g2579 = (((!g2) & (!g8) & (g2463) & (g2474)) + ((!g2) & (g8) & (!g2463) & (g2474)) + ((!g2) & (g8) & (g2463) & (!g2474)) + ((!g2) & (g8) & (g2463) & (g2474)) + ((g2) & (!g8) & (!g2463) & (!g2474)) + ((g2) & (!g8) & (!g2463) & (g2474)) + ((g2) & (!g8) & (g2463) & (!g2474)) + ((g2) & (g8) & (!g2463) & (!g2474)));
	assign g2580 = (((!g2462) & (!g2460) & (!g2478) & (g2579)) + ((!g2462) & (g2460) & (!g2478) & (g2579)) + ((!g2462) & (g2460) & (g2478) & (g2579)) + ((g2462) & (!g2460) & (!g2478) & (!g2579)) + ((g2462) & (!g2460) & (g2478) & (!g2579)) + ((g2462) & (!g2460) & (g2478) & (g2579)) + ((g2462) & (g2460) & (!g2478) & (!g2579)) + ((g2462) & (g2460) & (g2478) & (!g2579)));
	assign g2581 = (((!g4) & (!g2) & (!g2563) & (!g2578) & (g2580)) + ((!g4) & (!g2) & (!g2563) & (g2578) & (g2580)) + ((!g4) & (!g2) & (g2563) & (!g2578) & (g2580)) + ((!g4) & (!g2) & (g2563) & (g2578) & (!g2580)) + ((!g4) & (!g2) & (g2563) & (g2578) & (g2580)) + ((!g4) & (g2) & (!g2563) & (!g2578) & (g2580)) + ((!g4) & (g2) & (!g2563) & (g2578) & (!g2580)) + ((!g4) & (g2) & (!g2563) & (g2578) & (g2580)) + ((!g4) & (g2) & (g2563) & (!g2578) & (!g2580)) + ((!g4) & (g2) & (g2563) & (!g2578) & (g2580)) + ((!g4) & (g2) & (g2563) & (g2578) & (!g2580)) + ((!g4) & (g2) & (g2563) & (g2578) & (g2580)) + ((g4) & (!g2) & (g2563) & (g2578) & (g2580)) + ((g4) & (g2) & (!g2563) & (g2578) & (g2580)) + ((g4) & (g2) & (g2563) & (!g2578) & (g2580)) + ((g4) & (g2) & (g2563) & (g2578) & (g2580)));
	assign g2582 = (((!g4) & (!g2475) & (g2476)) + ((!g4) & (g2475) & (!g2476)) + ((!g4) & (g2475) & (g2476)) + ((g4) & (g2475) & (g2476)));
	assign g2583 = (((!g2461) & (!g2582) & (!g2460) & (!g2478)) + ((!g2461) & (!g2582) & (g2460) & (!g2478)) + ((!g2461) & (!g2582) & (g2460) & (g2478)) + ((g2461) & (g2582) & (!g2460) & (!g2478)) + ((g2461) & (g2582) & (!g2460) & (g2478)) + ((g2461) & (g2582) & (g2460) & (!g2478)) + ((g2461) & (g2582) & (g2460) & (g2478)));
	assign g2584 = (((!g1) & (g2461) & (!g2582) & (!g2460) & (g2478)) + ((!g1) & (g2461) & (g2582) & (!g2460) & (g2478)) + ((g1) & (!g2461) & (g2582) & (g2460) & (!g2478)) + ((g1) & (!g2461) & (g2582) & (g2460) & (g2478)) + ((g1) & (g2461) & (!g2582) & (!g2460) & (!g2478)) + ((g1) & (g2461) & (!g2582) & (!g2460) & (g2478)) + ((g1) & (g2461) & (!g2582) & (g2460) & (!g2478)) + ((g1) & (g2461) & (!g2582) & (g2460) & (g2478)) + ((g1) & (g2461) & (g2582) & (!g2460) & (g2478)));
	assign g2585 = (((!g1) & (!g2562) & (!g2581) & (!g2583) & (!g2584)) + ((g1) & (!g2562) & (!g2581) & (!g2583) & (!g2584)) + ((g1) & (!g2562) & (!g2581) & (g2583) & (!g2584)) + ((g1) & (!g2562) & (g2581) & (!g2583) & (!g2584)) + ((g1) & (!g2562) & (g2581) & (g2583) & (!g2584)) + ((g1) & (g2562) & (!g2581) & (!g2583) & (!g2584)) + ((g1) & (g2562) & (!g2581) & (g2583) & (!g2584)));
	assign g2586 = (((!g104) & (!g2479) & (g2561) & (!g2585)) + ((!g104) & (g2479) & (!g2561) & (!g2585)) + ((!g104) & (g2479) & (!g2561) & (g2585)) + ((!g104) & (g2479) & (g2561) & (g2585)) + ((g104) & (!g2479) & (!g2561) & (!g2585)) + ((g104) & (g2479) & (!g2561) & (g2585)) + ((g104) & (g2479) & (g2561) & (!g2585)) + ((g104) & (g2479) & (g2561) & (g2585)));
	assign g2587 = (((!g127) & (!g147) & (!g2481) & (g2482) & (g2560) & (!g2585)) + ((!g127) & (!g147) & (g2481) & (!g2482) & (!g2560) & (!g2585)) + ((!g127) & (!g147) & (g2481) & (!g2482) & (!g2560) & (g2585)) + ((!g127) & (!g147) & (g2481) & (!g2482) & (g2560) & (!g2585)) + ((!g127) & (!g147) & (g2481) & (!g2482) & (g2560) & (g2585)) + ((!g127) & (!g147) & (g2481) & (g2482) & (!g2560) & (!g2585)) + ((!g127) & (!g147) & (g2481) & (g2482) & (!g2560) & (g2585)) + ((!g127) & (!g147) & (g2481) & (g2482) & (g2560) & (g2585)) + ((!g127) & (g147) & (!g2481) & (!g2482) & (g2560) & (!g2585)) + ((!g127) & (g147) & (!g2481) & (g2482) & (!g2560) & (!g2585)) + ((!g127) & (g147) & (!g2481) & (g2482) & (g2560) & (!g2585)) + ((!g127) & (g147) & (g2481) & (!g2482) & (!g2560) & (!g2585)) + ((!g127) & (g147) & (g2481) & (!g2482) & (!g2560) & (g2585)) + ((!g127) & (g147) & (g2481) & (!g2482) & (g2560) & (g2585)) + ((!g127) & (g147) & (g2481) & (g2482) & (!g2560) & (g2585)) + ((!g127) & (g147) & (g2481) & (g2482) & (g2560) & (g2585)) + ((g127) & (!g147) & (!g2481) & (!g2482) & (!g2560) & (!g2585)) + ((g127) & (!g147) & (!g2481) & (!g2482) & (g2560) & (!g2585)) + ((g127) & (!g147) & (!g2481) & (g2482) & (!g2560) & (!g2585)) + ((g127) & (!g147) & (g2481) & (!g2482) & (!g2560) & (g2585)) + ((g127) & (!g147) & (g2481) & (!g2482) & (g2560) & (g2585)) + ((g127) & (!g147) & (g2481) & (g2482) & (!g2560) & (g2585)) + ((g127) & (!g147) & (g2481) & (g2482) & (g2560) & (!g2585)) + ((g127) & (!g147) & (g2481) & (g2482) & (g2560) & (g2585)) + ((g127) & (g147) & (!g2481) & (!g2482) & (!g2560) & (!g2585)) + ((g127) & (g147) & (g2481) & (!g2482) & (!g2560) & (g2585)) + ((g127) & (g147) & (g2481) & (!g2482) & (g2560) & (!g2585)) + ((g127) & (g147) & (g2481) & (!g2482) & (g2560) & (g2585)) + ((g127) & (g147) & (g2481) & (g2482) & (!g2560) & (!g2585)) + ((g127) & (g147) & (g2481) & (g2482) & (!g2560) & (g2585)) + ((g127) & (g147) & (g2481) & (g2482) & (g2560) & (!g2585)) + ((g127) & (g147) & (g2481) & (g2482) & (g2560) & (g2585)));
	assign g2588 = (((!g147) & (!g2482) & (g2560) & (!g2585)) + ((!g147) & (g2482) & (!g2560) & (!g2585)) + ((!g147) & (g2482) & (!g2560) & (g2585)) + ((!g147) & (g2482) & (g2560) & (g2585)) + ((g147) & (!g2482) & (!g2560) & (!g2585)) + ((g147) & (g2482) & (!g2560) & (g2585)) + ((g147) & (g2482) & (g2560) & (!g2585)) + ((g147) & (g2482) & (g2560) & (g2585)));
	assign g2589 = (((!g174) & (!g198) & (!g2484) & (g2485) & (g2559) & (!g2585)) + ((!g174) & (!g198) & (g2484) & (!g2485) & (!g2559) & (!g2585)) + ((!g174) & (!g198) & (g2484) & (!g2485) & (!g2559) & (g2585)) + ((!g174) & (!g198) & (g2484) & (!g2485) & (g2559) & (!g2585)) + ((!g174) & (!g198) & (g2484) & (!g2485) & (g2559) & (g2585)) + ((!g174) & (!g198) & (g2484) & (g2485) & (!g2559) & (!g2585)) + ((!g174) & (!g198) & (g2484) & (g2485) & (!g2559) & (g2585)) + ((!g174) & (!g198) & (g2484) & (g2485) & (g2559) & (g2585)) + ((!g174) & (g198) & (!g2484) & (!g2485) & (g2559) & (!g2585)) + ((!g174) & (g198) & (!g2484) & (g2485) & (!g2559) & (!g2585)) + ((!g174) & (g198) & (!g2484) & (g2485) & (g2559) & (!g2585)) + ((!g174) & (g198) & (g2484) & (!g2485) & (!g2559) & (!g2585)) + ((!g174) & (g198) & (g2484) & (!g2485) & (!g2559) & (g2585)) + ((!g174) & (g198) & (g2484) & (!g2485) & (g2559) & (g2585)) + ((!g174) & (g198) & (g2484) & (g2485) & (!g2559) & (g2585)) + ((!g174) & (g198) & (g2484) & (g2485) & (g2559) & (g2585)) + ((g174) & (!g198) & (!g2484) & (!g2485) & (!g2559) & (!g2585)) + ((g174) & (!g198) & (!g2484) & (!g2485) & (g2559) & (!g2585)) + ((g174) & (!g198) & (!g2484) & (g2485) & (!g2559) & (!g2585)) + ((g174) & (!g198) & (g2484) & (!g2485) & (!g2559) & (g2585)) + ((g174) & (!g198) & (g2484) & (!g2485) & (g2559) & (g2585)) + ((g174) & (!g198) & (g2484) & (g2485) & (!g2559) & (g2585)) + ((g174) & (!g198) & (g2484) & (g2485) & (g2559) & (!g2585)) + ((g174) & (!g198) & (g2484) & (g2485) & (g2559) & (g2585)) + ((g174) & (g198) & (!g2484) & (!g2485) & (!g2559) & (!g2585)) + ((g174) & (g198) & (g2484) & (!g2485) & (!g2559) & (g2585)) + ((g174) & (g198) & (g2484) & (!g2485) & (g2559) & (!g2585)) + ((g174) & (g198) & (g2484) & (!g2485) & (g2559) & (g2585)) + ((g174) & (g198) & (g2484) & (g2485) & (!g2559) & (!g2585)) + ((g174) & (g198) & (g2484) & (g2485) & (!g2559) & (g2585)) + ((g174) & (g198) & (g2484) & (g2485) & (g2559) & (!g2585)) + ((g174) & (g198) & (g2484) & (g2485) & (g2559) & (g2585)));
	assign g2590 = (((!g198) & (!g2485) & (g2559) & (!g2585)) + ((!g198) & (g2485) & (!g2559) & (!g2585)) + ((!g198) & (g2485) & (!g2559) & (g2585)) + ((!g198) & (g2485) & (g2559) & (g2585)) + ((g198) & (!g2485) & (!g2559) & (!g2585)) + ((g198) & (g2485) & (!g2559) & (g2585)) + ((g198) & (g2485) & (g2559) & (!g2585)) + ((g198) & (g2485) & (g2559) & (g2585)));
	assign g2591 = (((!g229) & (!g255) & (!g2487) & (g2488) & (g2558) & (!g2585)) + ((!g229) & (!g255) & (g2487) & (!g2488) & (!g2558) & (!g2585)) + ((!g229) & (!g255) & (g2487) & (!g2488) & (!g2558) & (g2585)) + ((!g229) & (!g255) & (g2487) & (!g2488) & (g2558) & (!g2585)) + ((!g229) & (!g255) & (g2487) & (!g2488) & (g2558) & (g2585)) + ((!g229) & (!g255) & (g2487) & (g2488) & (!g2558) & (!g2585)) + ((!g229) & (!g255) & (g2487) & (g2488) & (!g2558) & (g2585)) + ((!g229) & (!g255) & (g2487) & (g2488) & (g2558) & (g2585)) + ((!g229) & (g255) & (!g2487) & (!g2488) & (g2558) & (!g2585)) + ((!g229) & (g255) & (!g2487) & (g2488) & (!g2558) & (!g2585)) + ((!g229) & (g255) & (!g2487) & (g2488) & (g2558) & (!g2585)) + ((!g229) & (g255) & (g2487) & (!g2488) & (!g2558) & (!g2585)) + ((!g229) & (g255) & (g2487) & (!g2488) & (!g2558) & (g2585)) + ((!g229) & (g255) & (g2487) & (!g2488) & (g2558) & (g2585)) + ((!g229) & (g255) & (g2487) & (g2488) & (!g2558) & (g2585)) + ((!g229) & (g255) & (g2487) & (g2488) & (g2558) & (g2585)) + ((g229) & (!g255) & (!g2487) & (!g2488) & (!g2558) & (!g2585)) + ((g229) & (!g255) & (!g2487) & (!g2488) & (g2558) & (!g2585)) + ((g229) & (!g255) & (!g2487) & (g2488) & (!g2558) & (!g2585)) + ((g229) & (!g255) & (g2487) & (!g2488) & (!g2558) & (g2585)) + ((g229) & (!g255) & (g2487) & (!g2488) & (g2558) & (g2585)) + ((g229) & (!g255) & (g2487) & (g2488) & (!g2558) & (g2585)) + ((g229) & (!g255) & (g2487) & (g2488) & (g2558) & (!g2585)) + ((g229) & (!g255) & (g2487) & (g2488) & (g2558) & (g2585)) + ((g229) & (g255) & (!g2487) & (!g2488) & (!g2558) & (!g2585)) + ((g229) & (g255) & (g2487) & (!g2488) & (!g2558) & (g2585)) + ((g229) & (g255) & (g2487) & (!g2488) & (g2558) & (!g2585)) + ((g229) & (g255) & (g2487) & (!g2488) & (g2558) & (g2585)) + ((g229) & (g255) & (g2487) & (g2488) & (!g2558) & (!g2585)) + ((g229) & (g255) & (g2487) & (g2488) & (!g2558) & (g2585)) + ((g229) & (g255) & (g2487) & (g2488) & (g2558) & (!g2585)) + ((g229) & (g255) & (g2487) & (g2488) & (g2558) & (g2585)));
	assign g2592 = (((!g255) & (!g2488) & (g2558) & (!g2585)) + ((!g255) & (g2488) & (!g2558) & (!g2585)) + ((!g255) & (g2488) & (!g2558) & (g2585)) + ((!g255) & (g2488) & (g2558) & (g2585)) + ((g255) & (!g2488) & (!g2558) & (!g2585)) + ((g255) & (g2488) & (!g2558) & (g2585)) + ((g255) & (g2488) & (g2558) & (!g2585)) + ((g255) & (g2488) & (g2558) & (g2585)));
	assign g2593 = (((!g290) & (!g319) & (!g2490) & (g2491) & (g2557) & (!g2585)) + ((!g290) & (!g319) & (g2490) & (!g2491) & (!g2557) & (!g2585)) + ((!g290) & (!g319) & (g2490) & (!g2491) & (!g2557) & (g2585)) + ((!g290) & (!g319) & (g2490) & (!g2491) & (g2557) & (!g2585)) + ((!g290) & (!g319) & (g2490) & (!g2491) & (g2557) & (g2585)) + ((!g290) & (!g319) & (g2490) & (g2491) & (!g2557) & (!g2585)) + ((!g290) & (!g319) & (g2490) & (g2491) & (!g2557) & (g2585)) + ((!g290) & (!g319) & (g2490) & (g2491) & (g2557) & (g2585)) + ((!g290) & (g319) & (!g2490) & (!g2491) & (g2557) & (!g2585)) + ((!g290) & (g319) & (!g2490) & (g2491) & (!g2557) & (!g2585)) + ((!g290) & (g319) & (!g2490) & (g2491) & (g2557) & (!g2585)) + ((!g290) & (g319) & (g2490) & (!g2491) & (!g2557) & (!g2585)) + ((!g290) & (g319) & (g2490) & (!g2491) & (!g2557) & (g2585)) + ((!g290) & (g319) & (g2490) & (!g2491) & (g2557) & (g2585)) + ((!g290) & (g319) & (g2490) & (g2491) & (!g2557) & (g2585)) + ((!g290) & (g319) & (g2490) & (g2491) & (g2557) & (g2585)) + ((g290) & (!g319) & (!g2490) & (!g2491) & (!g2557) & (!g2585)) + ((g290) & (!g319) & (!g2490) & (!g2491) & (g2557) & (!g2585)) + ((g290) & (!g319) & (!g2490) & (g2491) & (!g2557) & (!g2585)) + ((g290) & (!g319) & (g2490) & (!g2491) & (!g2557) & (g2585)) + ((g290) & (!g319) & (g2490) & (!g2491) & (g2557) & (g2585)) + ((g290) & (!g319) & (g2490) & (g2491) & (!g2557) & (g2585)) + ((g290) & (!g319) & (g2490) & (g2491) & (g2557) & (!g2585)) + ((g290) & (!g319) & (g2490) & (g2491) & (g2557) & (g2585)) + ((g290) & (g319) & (!g2490) & (!g2491) & (!g2557) & (!g2585)) + ((g290) & (g319) & (g2490) & (!g2491) & (!g2557) & (g2585)) + ((g290) & (g319) & (g2490) & (!g2491) & (g2557) & (!g2585)) + ((g290) & (g319) & (g2490) & (!g2491) & (g2557) & (g2585)) + ((g290) & (g319) & (g2490) & (g2491) & (!g2557) & (!g2585)) + ((g290) & (g319) & (g2490) & (g2491) & (!g2557) & (g2585)) + ((g290) & (g319) & (g2490) & (g2491) & (g2557) & (!g2585)) + ((g290) & (g319) & (g2490) & (g2491) & (g2557) & (g2585)));
	assign g2594 = (((!g319) & (!g2491) & (g2557) & (!g2585)) + ((!g319) & (g2491) & (!g2557) & (!g2585)) + ((!g319) & (g2491) & (!g2557) & (g2585)) + ((!g319) & (g2491) & (g2557) & (g2585)) + ((g319) & (!g2491) & (!g2557) & (!g2585)) + ((g319) & (g2491) & (!g2557) & (g2585)) + ((g319) & (g2491) & (g2557) & (!g2585)) + ((g319) & (g2491) & (g2557) & (g2585)));
	assign g2595 = (((!g358) & (!g390) & (!g2493) & (g2494) & (g2556) & (!g2585)) + ((!g358) & (!g390) & (g2493) & (!g2494) & (!g2556) & (!g2585)) + ((!g358) & (!g390) & (g2493) & (!g2494) & (!g2556) & (g2585)) + ((!g358) & (!g390) & (g2493) & (!g2494) & (g2556) & (!g2585)) + ((!g358) & (!g390) & (g2493) & (!g2494) & (g2556) & (g2585)) + ((!g358) & (!g390) & (g2493) & (g2494) & (!g2556) & (!g2585)) + ((!g358) & (!g390) & (g2493) & (g2494) & (!g2556) & (g2585)) + ((!g358) & (!g390) & (g2493) & (g2494) & (g2556) & (g2585)) + ((!g358) & (g390) & (!g2493) & (!g2494) & (g2556) & (!g2585)) + ((!g358) & (g390) & (!g2493) & (g2494) & (!g2556) & (!g2585)) + ((!g358) & (g390) & (!g2493) & (g2494) & (g2556) & (!g2585)) + ((!g358) & (g390) & (g2493) & (!g2494) & (!g2556) & (!g2585)) + ((!g358) & (g390) & (g2493) & (!g2494) & (!g2556) & (g2585)) + ((!g358) & (g390) & (g2493) & (!g2494) & (g2556) & (g2585)) + ((!g358) & (g390) & (g2493) & (g2494) & (!g2556) & (g2585)) + ((!g358) & (g390) & (g2493) & (g2494) & (g2556) & (g2585)) + ((g358) & (!g390) & (!g2493) & (!g2494) & (!g2556) & (!g2585)) + ((g358) & (!g390) & (!g2493) & (!g2494) & (g2556) & (!g2585)) + ((g358) & (!g390) & (!g2493) & (g2494) & (!g2556) & (!g2585)) + ((g358) & (!g390) & (g2493) & (!g2494) & (!g2556) & (g2585)) + ((g358) & (!g390) & (g2493) & (!g2494) & (g2556) & (g2585)) + ((g358) & (!g390) & (g2493) & (g2494) & (!g2556) & (g2585)) + ((g358) & (!g390) & (g2493) & (g2494) & (g2556) & (!g2585)) + ((g358) & (!g390) & (g2493) & (g2494) & (g2556) & (g2585)) + ((g358) & (g390) & (!g2493) & (!g2494) & (!g2556) & (!g2585)) + ((g358) & (g390) & (g2493) & (!g2494) & (!g2556) & (g2585)) + ((g358) & (g390) & (g2493) & (!g2494) & (g2556) & (!g2585)) + ((g358) & (g390) & (g2493) & (!g2494) & (g2556) & (g2585)) + ((g358) & (g390) & (g2493) & (g2494) & (!g2556) & (!g2585)) + ((g358) & (g390) & (g2493) & (g2494) & (!g2556) & (g2585)) + ((g358) & (g390) & (g2493) & (g2494) & (g2556) & (!g2585)) + ((g358) & (g390) & (g2493) & (g2494) & (g2556) & (g2585)));
	assign g2596 = (((!g390) & (!g2494) & (g2556) & (!g2585)) + ((!g390) & (g2494) & (!g2556) & (!g2585)) + ((!g390) & (g2494) & (!g2556) & (g2585)) + ((!g390) & (g2494) & (g2556) & (g2585)) + ((g390) & (!g2494) & (!g2556) & (!g2585)) + ((g390) & (g2494) & (!g2556) & (g2585)) + ((g390) & (g2494) & (g2556) & (!g2585)) + ((g390) & (g2494) & (g2556) & (g2585)));
	assign g2597 = (((!g433) & (!g468) & (!g2496) & (g2497) & (g2555) & (!g2585)) + ((!g433) & (!g468) & (g2496) & (!g2497) & (!g2555) & (!g2585)) + ((!g433) & (!g468) & (g2496) & (!g2497) & (!g2555) & (g2585)) + ((!g433) & (!g468) & (g2496) & (!g2497) & (g2555) & (!g2585)) + ((!g433) & (!g468) & (g2496) & (!g2497) & (g2555) & (g2585)) + ((!g433) & (!g468) & (g2496) & (g2497) & (!g2555) & (!g2585)) + ((!g433) & (!g468) & (g2496) & (g2497) & (!g2555) & (g2585)) + ((!g433) & (!g468) & (g2496) & (g2497) & (g2555) & (g2585)) + ((!g433) & (g468) & (!g2496) & (!g2497) & (g2555) & (!g2585)) + ((!g433) & (g468) & (!g2496) & (g2497) & (!g2555) & (!g2585)) + ((!g433) & (g468) & (!g2496) & (g2497) & (g2555) & (!g2585)) + ((!g433) & (g468) & (g2496) & (!g2497) & (!g2555) & (!g2585)) + ((!g433) & (g468) & (g2496) & (!g2497) & (!g2555) & (g2585)) + ((!g433) & (g468) & (g2496) & (!g2497) & (g2555) & (g2585)) + ((!g433) & (g468) & (g2496) & (g2497) & (!g2555) & (g2585)) + ((!g433) & (g468) & (g2496) & (g2497) & (g2555) & (g2585)) + ((g433) & (!g468) & (!g2496) & (!g2497) & (!g2555) & (!g2585)) + ((g433) & (!g468) & (!g2496) & (!g2497) & (g2555) & (!g2585)) + ((g433) & (!g468) & (!g2496) & (g2497) & (!g2555) & (!g2585)) + ((g433) & (!g468) & (g2496) & (!g2497) & (!g2555) & (g2585)) + ((g433) & (!g468) & (g2496) & (!g2497) & (g2555) & (g2585)) + ((g433) & (!g468) & (g2496) & (g2497) & (!g2555) & (g2585)) + ((g433) & (!g468) & (g2496) & (g2497) & (g2555) & (!g2585)) + ((g433) & (!g468) & (g2496) & (g2497) & (g2555) & (g2585)) + ((g433) & (g468) & (!g2496) & (!g2497) & (!g2555) & (!g2585)) + ((g433) & (g468) & (g2496) & (!g2497) & (!g2555) & (g2585)) + ((g433) & (g468) & (g2496) & (!g2497) & (g2555) & (!g2585)) + ((g433) & (g468) & (g2496) & (!g2497) & (g2555) & (g2585)) + ((g433) & (g468) & (g2496) & (g2497) & (!g2555) & (!g2585)) + ((g433) & (g468) & (g2496) & (g2497) & (!g2555) & (g2585)) + ((g433) & (g468) & (g2496) & (g2497) & (g2555) & (!g2585)) + ((g433) & (g468) & (g2496) & (g2497) & (g2555) & (g2585)));
	assign g2598 = (((!g468) & (!g2497) & (g2555) & (!g2585)) + ((!g468) & (g2497) & (!g2555) & (!g2585)) + ((!g468) & (g2497) & (!g2555) & (g2585)) + ((!g468) & (g2497) & (g2555) & (g2585)) + ((g468) & (!g2497) & (!g2555) & (!g2585)) + ((g468) & (g2497) & (!g2555) & (g2585)) + ((g468) & (g2497) & (g2555) & (!g2585)) + ((g468) & (g2497) & (g2555) & (g2585)));
	assign g2599 = (((!g515) & (!g553) & (!g2499) & (g2500) & (g2554) & (!g2585)) + ((!g515) & (!g553) & (g2499) & (!g2500) & (!g2554) & (!g2585)) + ((!g515) & (!g553) & (g2499) & (!g2500) & (!g2554) & (g2585)) + ((!g515) & (!g553) & (g2499) & (!g2500) & (g2554) & (!g2585)) + ((!g515) & (!g553) & (g2499) & (!g2500) & (g2554) & (g2585)) + ((!g515) & (!g553) & (g2499) & (g2500) & (!g2554) & (!g2585)) + ((!g515) & (!g553) & (g2499) & (g2500) & (!g2554) & (g2585)) + ((!g515) & (!g553) & (g2499) & (g2500) & (g2554) & (g2585)) + ((!g515) & (g553) & (!g2499) & (!g2500) & (g2554) & (!g2585)) + ((!g515) & (g553) & (!g2499) & (g2500) & (!g2554) & (!g2585)) + ((!g515) & (g553) & (!g2499) & (g2500) & (g2554) & (!g2585)) + ((!g515) & (g553) & (g2499) & (!g2500) & (!g2554) & (!g2585)) + ((!g515) & (g553) & (g2499) & (!g2500) & (!g2554) & (g2585)) + ((!g515) & (g553) & (g2499) & (!g2500) & (g2554) & (g2585)) + ((!g515) & (g553) & (g2499) & (g2500) & (!g2554) & (g2585)) + ((!g515) & (g553) & (g2499) & (g2500) & (g2554) & (g2585)) + ((g515) & (!g553) & (!g2499) & (!g2500) & (!g2554) & (!g2585)) + ((g515) & (!g553) & (!g2499) & (!g2500) & (g2554) & (!g2585)) + ((g515) & (!g553) & (!g2499) & (g2500) & (!g2554) & (!g2585)) + ((g515) & (!g553) & (g2499) & (!g2500) & (!g2554) & (g2585)) + ((g515) & (!g553) & (g2499) & (!g2500) & (g2554) & (g2585)) + ((g515) & (!g553) & (g2499) & (g2500) & (!g2554) & (g2585)) + ((g515) & (!g553) & (g2499) & (g2500) & (g2554) & (!g2585)) + ((g515) & (!g553) & (g2499) & (g2500) & (g2554) & (g2585)) + ((g515) & (g553) & (!g2499) & (!g2500) & (!g2554) & (!g2585)) + ((g515) & (g553) & (g2499) & (!g2500) & (!g2554) & (g2585)) + ((g515) & (g553) & (g2499) & (!g2500) & (g2554) & (!g2585)) + ((g515) & (g553) & (g2499) & (!g2500) & (g2554) & (g2585)) + ((g515) & (g553) & (g2499) & (g2500) & (!g2554) & (!g2585)) + ((g515) & (g553) & (g2499) & (g2500) & (!g2554) & (g2585)) + ((g515) & (g553) & (g2499) & (g2500) & (g2554) & (!g2585)) + ((g515) & (g553) & (g2499) & (g2500) & (g2554) & (g2585)));
	assign g2600 = (((!g553) & (!g2500) & (g2554) & (!g2585)) + ((!g553) & (g2500) & (!g2554) & (!g2585)) + ((!g553) & (g2500) & (!g2554) & (g2585)) + ((!g553) & (g2500) & (g2554) & (g2585)) + ((g553) & (!g2500) & (!g2554) & (!g2585)) + ((g553) & (g2500) & (!g2554) & (g2585)) + ((g553) & (g2500) & (g2554) & (!g2585)) + ((g553) & (g2500) & (g2554) & (g2585)));
	assign g2601 = (((!g604) & (!g645) & (!g2502) & (g2503) & (g2553) & (!g2585)) + ((!g604) & (!g645) & (g2502) & (!g2503) & (!g2553) & (!g2585)) + ((!g604) & (!g645) & (g2502) & (!g2503) & (!g2553) & (g2585)) + ((!g604) & (!g645) & (g2502) & (!g2503) & (g2553) & (!g2585)) + ((!g604) & (!g645) & (g2502) & (!g2503) & (g2553) & (g2585)) + ((!g604) & (!g645) & (g2502) & (g2503) & (!g2553) & (!g2585)) + ((!g604) & (!g645) & (g2502) & (g2503) & (!g2553) & (g2585)) + ((!g604) & (!g645) & (g2502) & (g2503) & (g2553) & (g2585)) + ((!g604) & (g645) & (!g2502) & (!g2503) & (g2553) & (!g2585)) + ((!g604) & (g645) & (!g2502) & (g2503) & (!g2553) & (!g2585)) + ((!g604) & (g645) & (!g2502) & (g2503) & (g2553) & (!g2585)) + ((!g604) & (g645) & (g2502) & (!g2503) & (!g2553) & (!g2585)) + ((!g604) & (g645) & (g2502) & (!g2503) & (!g2553) & (g2585)) + ((!g604) & (g645) & (g2502) & (!g2503) & (g2553) & (g2585)) + ((!g604) & (g645) & (g2502) & (g2503) & (!g2553) & (g2585)) + ((!g604) & (g645) & (g2502) & (g2503) & (g2553) & (g2585)) + ((g604) & (!g645) & (!g2502) & (!g2503) & (!g2553) & (!g2585)) + ((g604) & (!g645) & (!g2502) & (!g2503) & (g2553) & (!g2585)) + ((g604) & (!g645) & (!g2502) & (g2503) & (!g2553) & (!g2585)) + ((g604) & (!g645) & (g2502) & (!g2503) & (!g2553) & (g2585)) + ((g604) & (!g645) & (g2502) & (!g2503) & (g2553) & (g2585)) + ((g604) & (!g645) & (g2502) & (g2503) & (!g2553) & (g2585)) + ((g604) & (!g645) & (g2502) & (g2503) & (g2553) & (!g2585)) + ((g604) & (!g645) & (g2502) & (g2503) & (g2553) & (g2585)) + ((g604) & (g645) & (!g2502) & (!g2503) & (!g2553) & (!g2585)) + ((g604) & (g645) & (g2502) & (!g2503) & (!g2553) & (g2585)) + ((g604) & (g645) & (g2502) & (!g2503) & (g2553) & (!g2585)) + ((g604) & (g645) & (g2502) & (!g2503) & (g2553) & (g2585)) + ((g604) & (g645) & (g2502) & (g2503) & (!g2553) & (!g2585)) + ((g604) & (g645) & (g2502) & (g2503) & (!g2553) & (g2585)) + ((g604) & (g645) & (g2502) & (g2503) & (g2553) & (!g2585)) + ((g604) & (g645) & (g2502) & (g2503) & (g2553) & (g2585)));
	assign g2602 = (((!g645) & (!g2503) & (g2553) & (!g2585)) + ((!g645) & (g2503) & (!g2553) & (!g2585)) + ((!g645) & (g2503) & (!g2553) & (g2585)) + ((!g645) & (g2503) & (g2553) & (g2585)) + ((g645) & (!g2503) & (!g2553) & (!g2585)) + ((g645) & (g2503) & (!g2553) & (g2585)) + ((g645) & (g2503) & (g2553) & (!g2585)) + ((g645) & (g2503) & (g2553) & (g2585)));
	assign g2603 = (((!g700) & (!g744) & (!g2505) & (g2506) & (g2552) & (!g2585)) + ((!g700) & (!g744) & (g2505) & (!g2506) & (!g2552) & (!g2585)) + ((!g700) & (!g744) & (g2505) & (!g2506) & (!g2552) & (g2585)) + ((!g700) & (!g744) & (g2505) & (!g2506) & (g2552) & (!g2585)) + ((!g700) & (!g744) & (g2505) & (!g2506) & (g2552) & (g2585)) + ((!g700) & (!g744) & (g2505) & (g2506) & (!g2552) & (!g2585)) + ((!g700) & (!g744) & (g2505) & (g2506) & (!g2552) & (g2585)) + ((!g700) & (!g744) & (g2505) & (g2506) & (g2552) & (g2585)) + ((!g700) & (g744) & (!g2505) & (!g2506) & (g2552) & (!g2585)) + ((!g700) & (g744) & (!g2505) & (g2506) & (!g2552) & (!g2585)) + ((!g700) & (g744) & (!g2505) & (g2506) & (g2552) & (!g2585)) + ((!g700) & (g744) & (g2505) & (!g2506) & (!g2552) & (!g2585)) + ((!g700) & (g744) & (g2505) & (!g2506) & (!g2552) & (g2585)) + ((!g700) & (g744) & (g2505) & (!g2506) & (g2552) & (g2585)) + ((!g700) & (g744) & (g2505) & (g2506) & (!g2552) & (g2585)) + ((!g700) & (g744) & (g2505) & (g2506) & (g2552) & (g2585)) + ((g700) & (!g744) & (!g2505) & (!g2506) & (!g2552) & (!g2585)) + ((g700) & (!g744) & (!g2505) & (!g2506) & (g2552) & (!g2585)) + ((g700) & (!g744) & (!g2505) & (g2506) & (!g2552) & (!g2585)) + ((g700) & (!g744) & (g2505) & (!g2506) & (!g2552) & (g2585)) + ((g700) & (!g744) & (g2505) & (!g2506) & (g2552) & (g2585)) + ((g700) & (!g744) & (g2505) & (g2506) & (!g2552) & (g2585)) + ((g700) & (!g744) & (g2505) & (g2506) & (g2552) & (!g2585)) + ((g700) & (!g744) & (g2505) & (g2506) & (g2552) & (g2585)) + ((g700) & (g744) & (!g2505) & (!g2506) & (!g2552) & (!g2585)) + ((g700) & (g744) & (g2505) & (!g2506) & (!g2552) & (g2585)) + ((g700) & (g744) & (g2505) & (!g2506) & (g2552) & (!g2585)) + ((g700) & (g744) & (g2505) & (!g2506) & (g2552) & (g2585)) + ((g700) & (g744) & (g2505) & (g2506) & (!g2552) & (!g2585)) + ((g700) & (g744) & (g2505) & (g2506) & (!g2552) & (g2585)) + ((g700) & (g744) & (g2505) & (g2506) & (g2552) & (!g2585)) + ((g700) & (g744) & (g2505) & (g2506) & (g2552) & (g2585)));
	assign g2604 = (((!g744) & (!g2506) & (g2552) & (!g2585)) + ((!g744) & (g2506) & (!g2552) & (!g2585)) + ((!g744) & (g2506) & (!g2552) & (g2585)) + ((!g744) & (g2506) & (g2552) & (g2585)) + ((g744) & (!g2506) & (!g2552) & (!g2585)) + ((g744) & (g2506) & (!g2552) & (g2585)) + ((g744) & (g2506) & (g2552) & (!g2585)) + ((g744) & (g2506) & (g2552) & (g2585)));
	assign g2605 = (((!g803) & (!g851) & (!g2508) & (g2509) & (g2551) & (!g2585)) + ((!g803) & (!g851) & (g2508) & (!g2509) & (!g2551) & (!g2585)) + ((!g803) & (!g851) & (g2508) & (!g2509) & (!g2551) & (g2585)) + ((!g803) & (!g851) & (g2508) & (!g2509) & (g2551) & (!g2585)) + ((!g803) & (!g851) & (g2508) & (!g2509) & (g2551) & (g2585)) + ((!g803) & (!g851) & (g2508) & (g2509) & (!g2551) & (!g2585)) + ((!g803) & (!g851) & (g2508) & (g2509) & (!g2551) & (g2585)) + ((!g803) & (!g851) & (g2508) & (g2509) & (g2551) & (g2585)) + ((!g803) & (g851) & (!g2508) & (!g2509) & (g2551) & (!g2585)) + ((!g803) & (g851) & (!g2508) & (g2509) & (!g2551) & (!g2585)) + ((!g803) & (g851) & (!g2508) & (g2509) & (g2551) & (!g2585)) + ((!g803) & (g851) & (g2508) & (!g2509) & (!g2551) & (!g2585)) + ((!g803) & (g851) & (g2508) & (!g2509) & (!g2551) & (g2585)) + ((!g803) & (g851) & (g2508) & (!g2509) & (g2551) & (g2585)) + ((!g803) & (g851) & (g2508) & (g2509) & (!g2551) & (g2585)) + ((!g803) & (g851) & (g2508) & (g2509) & (g2551) & (g2585)) + ((g803) & (!g851) & (!g2508) & (!g2509) & (!g2551) & (!g2585)) + ((g803) & (!g851) & (!g2508) & (!g2509) & (g2551) & (!g2585)) + ((g803) & (!g851) & (!g2508) & (g2509) & (!g2551) & (!g2585)) + ((g803) & (!g851) & (g2508) & (!g2509) & (!g2551) & (g2585)) + ((g803) & (!g851) & (g2508) & (!g2509) & (g2551) & (g2585)) + ((g803) & (!g851) & (g2508) & (g2509) & (!g2551) & (g2585)) + ((g803) & (!g851) & (g2508) & (g2509) & (g2551) & (!g2585)) + ((g803) & (!g851) & (g2508) & (g2509) & (g2551) & (g2585)) + ((g803) & (g851) & (!g2508) & (!g2509) & (!g2551) & (!g2585)) + ((g803) & (g851) & (g2508) & (!g2509) & (!g2551) & (g2585)) + ((g803) & (g851) & (g2508) & (!g2509) & (g2551) & (!g2585)) + ((g803) & (g851) & (g2508) & (!g2509) & (g2551) & (g2585)) + ((g803) & (g851) & (g2508) & (g2509) & (!g2551) & (!g2585)) + ((g803) & (g851) & (g2508) & (g2509) & (!g2551) & (g2585)) + ((g803) & (g851) & (g2508) & (g2509) & (g2551) & (!g2585)) + ((g803) & (g851) & (g2508) & (g2509) & (g2551) & (g2585)));
	assign g2606 = (((!g851) & (!g2509) & (g2551) & (!g2585)) + ((!g851) & (g2509) & (!g2551) & (!g2585)) + ((!g851) & (g2509) & (!g2551) & (g2585)) + ((!g851) & (g2509) & (g2551) & (g2585)) + ((g851) & (!g2509) & (!g2551) & (!g2585)) + ((g851) & (g2509) & (!g2551) & (g2585)) + ((g851) & (g2509) & (g2551) & (!g2585)) + ((g851) & (g2509) & (g2551) & (g2585)));
	assign g2607 = (((!g914) & (!g1032) & (!g2511) & (g2512) & (g2550) & (!g2585)) + ((!g914) & (!g1032) & (g2511) & (!g2512) & (!g2550) & (!g2585)) + ((!g914) & (!g1032) & (g2511) & (!g2512) & (!g2550) & (g2585)) + ((!g914) & (!g1032) & (g2511) & (!g2512) & (g2550) & (!g2585)) + ((!g914) & (!g1032) & (g2511) & (!g2512) & (g2550) & (g2585)) + ((!g914) & (!g1032) & (g2511) & (g2512) & (!g2550) & (!g2585)) + ((!g914) & (!g1032) & (g2511) & (g2512) & (!g2550) & (g2585)) + ((!g914) & (!g1032) & (g2511) & (g2512) & (g2550) & (g2585)) + ((!g914) & (g1032) & (!g2511) & (!g2512) & (g2550) & (!g2585)) + ((!g914) & (g1032) & (!g2511) & (g2512) & (!g2550) & (!g2585)) + ((!g914) & (g1032) & (!g2511) & (g2512) & (g2550) & (!g2585)) + ((!g914) & (g1032) & (g2511) & (!g2512) & (!g2550) & (!g2585)) + ((!g914) & (g1032) & (g2511) & (!g2512) & (!g2550) & (g2585)) + ((!g914) & (g1032) & (g2511) & (!g2512) & (g2550) & (g2585)) + ((!g914) & (g1032) & (g2511) & (g2512) & (!g2550) & (g2585)) + ((!g914) & (g1032) & (g2511) & (g2512) & (g2550) & (g2585)) + ((g914) & (!g1032) & (!g2511) & (!g2512) & (!g2550) & (!g2585)) + ((g914) & (!g1032) & (!g2511) & (!g2512) & (g2550) & (!g2585)) + ((g914) & (!g1032) & (!g2511) & (g2512) & (!g2550) & (!g2585)) + ((g914) & (!g1032) & (g2511) & (!g2512) & (!g2550) & (g2585)) + ((g914) & (!g1032) & (g2511) & (!g2512) & (g2550) & (g2585)) + ((g914) & (!g1032) & (g2511) & (g2512) & (!g2550) & (g2585)) + ((g914) & (!g1032) & (g2511) & (g2512) & (g2550) & (!g2585)) + ((g914) & (!g1032) & (g2511) & (g2512) & (g2550) & (g2585)) + ((g914) & (g1032) & (!g2511) & (!g2512) & (!g2550) & (!g2585)) + ((g914) & (g1032) & (g2511) & (!g2512) & (!g2550) & (g2585)) + ((g914) & (g1032) & (g2511) & (!g2512) & (g2550) & (!g2585)) + ((g914) & (g1032) & (g2511) & (!g2512) & (g2550) & (g2585)) + ((g914) & (g1032) & (g2511) & (g2512) & (!g2550) & (!g2585)) + ((g914) & (g1032) & (g2511) & (g2512) & (!g2550) & (g2585)) + ((g914) & (g1032) & (g2511) & (g2512) & (g2550) & (!g2585)) + ((g914) & (g1032) & (g2511) & (g2512) & (g2550) & (g2585)));
	assign g2608 = (((!g1032) & (!g2512) & (g2550) & (!g2585)) + ((!g1032) & (g2512) & (!g2550) & (!g2585)) + ((!g1032) & (g2512) & (!g2550) & (g2585)) + ((!g1032) & (g2512) & (g2550) & (g2585)) + ((g1032) & (!g2512) & (!g2550) & (!g2585)) + ((g1032) & (g2512) & (!g2550) & (g2585)) + ((g1032) & (g2512) & (g2550) & (!g2585)) + ((g1032) & (g2512) & (g2550) & (g2585)));
	assign g2609 = (((!g1030) & (!g1160) & (!g2514) & (g2515) & (g2549) & (!g2585)) + ((!g1030) & (!g1160) & (g2514) & (!g2515) & (!g2549) & (!g2585)) + ((!g1030) & (!g1160) & (g2514) & (!g2515) & (!g2549) & (g2585)) + ((!g1030) & (!g1160) & (g2514) & (!g2515) & (g2549) & (!g2585)) + ((!g1030) & (!g1160) & (g2514) & (!g2515) & (g2549) & (g2585)) + ((!g1030) & (!g1160) & (g2514) & (g2515) & (!g2549) & (!g2585)) + ((!g1030) & (!g1160) & (g2514) & (g2515) & (!g2549) & (g2585)) + ((!g1030) & (!g1160) & (g2514) & (g2515) & (g2549) & (g2585)) + ((!g1030) & (g1160) & (!g2514) & (!g2515) & (g2549) & (!g2585)) + ((!g1030) & (g1160) & (!g2514) & (g2515) & (!g2549) & (!g2585)) + ((!g1030) & (g1160) & (!g2514) & (g2515) & (g2549) & (!g2585)) + ((!g1030) & (g1160) & (g2514) & (!g2515) & (!g2549) & (!g2585)) + ((!g1030) & (g1160) & (g2514) & (!g2515) & (!g2549) & (g2585)) + ((!g1030) & (g1160) & (g2514) & (!g2515) & (g2549) & (g2585)) + ((!g1030) & (g1160) & (g2514) & (g2515) & (!g2549) & (g2585)) + ((!g1030) & (g1160) & (g2514) & (g2515) & (g2549) & (g2585)) + ((g1030) & (!g1160) & (!g2514) & (!g2515) & (!g2549) & (!g2585)) + ((g1030) & (!g1160) & (!g2514) & (!g2515) & (g2549) & (!g2585)) + ((g1030) & (!g1160) & (!g2514) & (g2515) & (!g2549) & (!g2585)) + ((g1030) & (!g1160) & (g2514) & (!g2515) & (!g2549) & (g2585)) + ((g1030) & (!g1160) & (g2514) & (!g2515) & (g2549) & (g2585)) + ((g1030) & (!g1160) & (g2514) & (g2515) & (!g2549) & (g2585)) + ((g1030) & (!g1160) & (g2514) & (g2515) & (g2549) & (!g2585)) + ((g1030) & (!g1160) & (g2514) & (g2515) & (g2549) & (g2585)) + ((g1030) & (g1160) & (!g2514) & (!g2515) & (!g2549) & (!g2585)) + ((g1030) & (g1160) & (g2514) & (!g2515) & (!g2549) & (g2585)) + ((g1030) & (g1160) & (g2514) & (!g2515) & (g2549) & (!g2585)) + ((g1030) & (g1160) & (g2514) & (!g2515) & (g2549) & (g2585)) + ((g1030) & (g1160) & (g2514) & (g2515) & (!g2549) & (!g2585)) + ((g1030) & (g1160) & (g2514) & (g2515) & (!g2549) & (g2585)) + ((g1030) & (g1160) & (g2514) & (g2515) & (g2549) & (!g2585)) + ((g1030) & (g1160) & (g2514) & (g2515) & (g2549) & (g2585)));
	assign g2610 = (((!g1160) & (!g2515) & (g2549) & (!g2585)) + ((!g1160) & (g2515) & (!g2549) & (!g2585)) + ((!g1160) & (g2515) & (!g2549) & (g2585)) + ((!g1160) & (g2515) & (g2549) & (g2585)) + ((g1160) & (!g2515) & (!g2549) & (!g2585)) + ((g1160) & (g2515) & (!g2549) & (g2585)) + ((g1160) & (g2515) & (g2549) & (!g2585)) + ((g1160) & (g2515) & (g2549) & (g2585)));
	assign g2611 = (((!g1154) & (!g1295) & (!g2517) & (g2518) & (g2548) & (!g2585)) + ((!g1154) & (!g1295) & (g2517) & (!g2518) & (!g2548) & (!g2585)) + ((!g1154) & (!g1295) & (g2517) & (!g2518) & (!g2548) & (g2585)) + ((!g1154) & (!g1295) & (g2517) & (!g2518) & (g2548) & (!g2585)) + ((!g1154) & (!g1295) & (g2517) & (!g2518) & (g2548) & (g2585)) + ((!g1154) & (!g1295) & (g2517) & (g2518) & (!g2548) & (!g2585)) + ((!g1154) & (!g1295) & (g2517) & (g2518) & (!g2548) & (g2585)) + ((!g1154) & (!g1295) & (g2517) & (g2518) & (g2548) & (g2585)) + ((!g1154) & (g1295) & (!g2517) & (!g2518) & (g2548) & (!g2585)) + ((!g1154) & (g1295) & (!g2517) & (g2518) & (!g2548) & (!g2585)) + ((!g1154) & (g1295) & (!g2517) & (g2518) & (g2548) & (!g2585)) + ((!g1154) & (g1295) & (g2517) & (!g2518) & (!g2548) & (!g2585)) + ((!g1154) & (g1295) & (g2517) & (!g2518) & (!g2548) & (g2585)) + ((!g1154) & (g1295) & (g2517) & (!g2518) & (g2548) & (g2585)) + ((!g1154) & (g1295) & (g2517) & (g2518) & (!g2548) & (g2585)) + ((!g1154) & (g1295) & (g2517) & (g2518) & (g2548) & (g2585)) + ((g1154) & (!g1295) & (!g2517) & (!g2518) & (!g2548) & (!g2585)) + ((g1154) & (!g1295) & (!g2517) & (!g2518) & (g2548) & (!g2585)) + ((g1154) & (!g1295) & (!g2517) & (g2518) & (!g2548) & (!g2585)) + ((g1154) & (!g1295) & (g2517) & (!g2518) & (!g2548) & (g2585)) + ((g1154) & (!g1295) & (g2517) & (!g2518) & (g2548) & (g2585)) + ((g1154) & (!g1295) & (g2517) & (g2518) & (!g2548) & (g2585)) + ((g1154) & (!g1295) & (g2517) & (g2518) & (g2548) & (!g2585)) + ((g1154) & (!g1295) & (g2517) & (g2518) & (g2548) & (g2585)) + ((g1154) & (g1295) & (!g2517) & (!g2518) & (!g2548) & (!g2585)) + ((g1154) & (g1295) & (g2517) & (!g2518) & (!g2548) & (g2585)) + ((g1154) & (g1295) & (g2517) & (!g2518) & (g2548) & (!g2585)) + ((g1154) & (g1295) & (g2517) & (!g2518) & (g2548) & (g2585)) + ((g1154) & (g1295) & (g2517) & (g2518) & (!g2548) & (!g2585)) + ((g1154) & (g1295) & (g2517) & (g2518) & (!g2548) & (g2585)) + ((g1154) & (g1295) & (g2517) & (g2518) & (g2548) & (!g2585)) + ((g1154) & (g1295) & (g2517) & (g2518) & (g2548) & (g2585)));
	assign g2612 = (((!g1295) & (!g2518) & (g2548) & (!g2585)) + ((!g1295) & (g2518) & (!g2548) & (!g2585)) + ((!g1295) & (g2518) & (!g2548) & (g2585)) + ((!g1295) & (g2518) & (g2548) & (g2585)) + ((g1295) & (!g2518) & (!g2548) & (!g2585)) + ((g1295) & (g2518) & (!g2548) & (g2585)) + ((g1295) & (g2518) & (g2548) & (!g2585)) + ((g1295) & (g2518) & (g2548) & (g2585)));
	assign g2613 = (((!g1285) & (!g1437) & (!g2520) & (g2521) & (g2547) & (!g2585)) + ((!g1285) & (!g1437) & (g2520) & (!g2521) & (!g2547) & (!g2585)) + ((!g1285) & (!g1437) & (g2520) & (!g2521) & (!g2547) & (g2585)) + ((!g1285) & (!g1437) & (g2520) & (!g2521) & (g2547) & (!g2585)) + ((!g1285) & (!g1437) & (g2520) & (!g2521) & (g2547) & (g2585)) + ((!g1285) & (!g1437) & (g2520) & (g2521) & (!g2547) & (!g2585)) + ((!g1285) & (!g1437) & (g2520) & (g2521) & (!g2547) & (g2585)) + ((!g1285) & (!g1437) & (g2520) & (g2521) & (g2547) & (g2585)) + ((!g1285) & (g1437) & (!g2520) & (!g2521) & (g2547) & (!g2585)) + ((!g1285) & (g1437) & (!g2520) & (g2521) & (!g2547) & (!g2585)) + ((!g1285) & (g1437) & (!g2520) & (g2521) & (g2547) & (!g2585)) + ((!g1285) & (g1437) & (g2520) & (!g2521) & (!g2547) & (!g2585)) + ((!g1285) & (g1437) & (g2520) & (!g2521) & (!g2547) & (g2585)) + ((!g1285) & (g1437) & (g2520) & (!g2521) & (g2547) & (g2585)) + ((!g1285) & (g1437) & (g2520) & (g2521) & (!g2547) & (g2585)) + ((!g1285) & (g1437) & (g2520) & (g2521) & (g2547) & (g2585)) + ((g1285) & (!g1437) & (!g2520) & (!g2521) & (!g2547) & (!g2585)) + ((g1285) & (!g1437) & (!g2520) & (!g2521) & (g2547) & (!g2585)) + ((g1285) & (!g1437) & (!g2520) & (g2521) & (!g2547) & (!g2585)) + ((g1285) & (!g1437) & (g2520) & (!g2521) & (!g2547) & (g2585)) + ((g1285) & (!g1437) & (g2520) & (!g2521) & (g2547) & (g2585)) + ((g1285) & (!g1437) & (g2520) & (g2521) & (!g2547) & (g2585)) + ((g1285) & (!g1437) & (g2520) & (g2521) & (g2547) & (!g2585)) + ((g1285) & (!g1437) & (g2520) & (g2521) & (g2547) & (g2585)) + ((g1285) & (g1437) & (!g2520) & (!g2521) & (!g2547) & (!g2585)) + ((g1285) & (g1437) & (g2520) & (!g2521) & (!g2547) & (g2585)) + ((g1285) & (g1437) & (g2520) & (!g2521) & (g2547) & (!g2585)) + ((g1285) & (g1437) & (g2520) & (!g2521) & (g2547) & (g2585)) + ((g1285) & (g1437) & (g2520) & (g2521) & (!g2547) & (!g2585)) + ((g1285) & (g1437) & (g2520) & (g2521) & (!g2547) & (g2585)) + ((g1285) & (g1437) & (g2520) & (g2521) & (g2547) & (!g2585)) + ((g1285) & (g1437) & (g2520) & (g2521) & (g2547) & (g2585)));
	assign g2614 = (((!g1437) & (!g2521) & (g2547) & (!g2585)) + ((!g1437) & (g2521) & (!g2547) & (!g2585)) + ((!g1437) & (g2521) & (!g2547) & (g2585)) + ((!g1437) & (g2521) & (g2547) & (g2585)) + ((g1437) & (!g2521) & (!g2547) & (!g2585)) + ((g1437) & (g2521) & (!g2547) & (g2585)) + ((g1437) & (g2521) & (g2547) & (!g2585)) + ((g1437) & (g2521) & (g2547) & (g2585)));
	assign g2615 = (((!g1423) & (!g1586) & (!g2523) & (g2524) & (g2546) & (!g2585)) + ((!g1423) & (!g1586) & (g2523) & (!g2524) & (!g2546) & (!g2585)) + ((!g1423) & (!g1586) & (g2523) & (!g2524) & (!g2546) & (g2585)) + ((!g1423) & (!g1586) & (g2523) & (!g2524) & (g2546) & (!g2585)) + ((!g1423) & (!g1586) & (g2523) & (!g2524) & (g2546) & (g2585)) + ((!g1423) & (!g1586) & (g2523) & (g2524) & (!g2546) & (!g2585)) + ((!g1423) & (!g1586) & (g2523) & (g2524) & (!g2546) & (g2585)) + ((!g1423) & (!g1586) & (g2523) & (g2524) & (g2546) & (g2585)) + ((!g1423) & (g1586) & (!g2523) & (!g2524) & (g2546) & (!g2585)) + ((!g1423) & (g1586) & (!g2523) & (g2524) & (!g2546) & (!g2585)) + ((!g1423) & (g1586) & (!g2523) & (g2524) & (g2546) & (!g2585)) + ((!g1423) & (g1586) & (g2523) & (!g2524) & (!g2546) & (!g2585)) + ((!g1423) & (g1586) & (g2523) & (!g2524) & (!g2546) & (g2585)) + ((!g1423) & (g1586) & (g2523) & (!g2524) & (g2546) & (g2585)) + ((!g1423) & (g1586) & (g2523) & (g2524) & (!g2546) & (g2585)) + ((!g1423) & (g1586) & (g2523) & (g2524) & (g2546) & (g2585)) + ((g1423) & (!g1586) & (!g2523) & (!g2524) & (!g2546) & (!g2585)) + ((g1423) & (!g1586) & (!g2523) & (!g2524) & (g2546) & (!g2585)) + ((g1423) & (!g1586) & (!g2523) & (g2524) & (!g2546) & (!g2585)) + ((g1423) & (!g1586) & (g2523) & (!g2524) & (!g2546) & (g2585)) + ((g1423) & (!g1586) & (g2523) & (!g2524) & (g2546) & (g2585)) + ((g1423) & (!g1586) & (g2523) & (g2524) & (!g2546) & (g2585)) + ((g1423) & (!g1586) & (g2523) & (g2524) & (g2546) & (!g2585)) + ((g1423) & (!g1586) & (g2523) & (g2524) & (g2546) & (g2585)) + ((g1423) & (g1586) & (!g2523) & (!g2524) & (!g2546) & (!g2585)) + ((g1423) & (g1586) & (g2523) & (!g2524) & (!g2546) & (g2585)) + ((g1423) & (g1586) & (g2523) & (!g2524) & (g2546) & (!g2585)) + ((g1423) & (g1586) & (g2523) & (!g2524) & (g2546) & (g2585)) + ((g1423) & (g1586) & (g2523) & (g2524) & (!g2546) & (!g2585)) + ((g1423) & (g1586) & (g2523) & (g2524) & (!g2546) & (g2585)) + ((g1423) & (g1586) & (g2523) & (g2524) & (g2546) & (!g2585)) + ((g1423) & (g1586) & (g2523) & (g2524) & (g2546) & (g2585)));
	assign g2616 = (((!g1586) & (!g2524) & (g2546) & (!g2585)) + ((!g1586) & (g2524) & (!g2546) & (!g2585)) + ((!g1586) & (g2524) & (!g2546) & (g2585)) + ((!g1586) & (g2524) & (g2546) & (g2585)) + ((g1586) & (!g2524) & (!g2546) & (!g2585)) + ((g1586) & (g2524) & (!g2546) & (g2585)) + ((g1586) & (g2524) & (g2546) & (!g2585)) + ((g1586) & (g2524) & (g2546) & (g2585)));
	assign g2617 = (((!g1568) & (!g1742) & (!g2526) & (g2527) & (g2545) & (!g2585)) + ((!g1568) & (!g1742) & (g2526) & (!g2527) & (!g2545) & (!g2585)) + ((!g1568) & (!g1742) & (g2526) & (!g2527) & (!g2545) & (g2585)) + ((!g1568) & (!g1742) & (g2526) & (!g2527) & (g2545) & (!g2585)) + ((!g1568) & (!g1742) & (g2526) & (!g2527) & (g2545) & (g2585)) + ((!g1568) & (!g1742) & (g2526) & (g2527) & (!g2545) & (!g2585)) + ((!g1568) & (!g1742) & (g2526) & (g2527) & (!g2545) & (g2585)) + ((!g1568) & (!g1742) & (g2526) & (g2527) & (g2545) & (g2585)) + ((!g1568) & (g1742) & (!g2526) & (!g2527) & (g2545) & (!g2585)) + ((!g1568) & (g1742) & (!g2526) & (g2527) & (!g2545) & (!g2585)) + ((!g1568) & (g1742) & (!g2526) & (g2527) & (g2545) & (!g2585)) + ((!g1568) & (g1742) & (g2526) & (!g2527) & (!g2545) & (!g2585)) + ((!g1568) & (g1742) & (g2526) & (!g2527) & (!g2545) & (g2585)) + ((!g1568) & (g1742) & (g2526) & (!g2527) & (g2545) & (g2585)) + ((!g1568) & (g1742) & (g2526) & (g2527) & (!g2545) & (g2585)) + ((!g1568) & (g1742) & (g2526) & (g2527) & (g2545) & (g2585)) + ((g1568) & (!g1742) & (!g2526) & (!g2527) & (!g2545) & (!g2585)) + ((g1568) & (!g1742) & (!g2526) & (!g2527) & (g2545) & (!g2585)) + ((g1568) & (!g1742) & (!g2526) & (g2527) & (!g2545) & (!g2585)) + ((g1568) & (!g1742) & (g2526) & (!g2527) & (!g2545) & (g2585)) + ((g1568) & (!g1742) & (g2526) & (!g2527) & (g2545) & (g2585)) + ((g1568) & (!g1742) & (g2526) & (g2527) & (!g2545) & (g2585)) + ((g1568) & (!g1742) & (g2526) & (g2527) & (g2545) & (!g2585)) + ((g1568) & (!g1742) & (g2526) & (g2527) & (g2545) & (g2585)) + ((g1568) & (g1742) & (!g2526) & (!g2527) & (!g2545) & (!g2585)) + ((g1568) & (g1742) & (g2526) & (!g2527) & (!g2545) & (g2585)) + ((g1568) & (g1742) & (g2526) & (!g2527) & (g2545) & (!g2585)) + ((g1568) & (g1742) & (g2526) & (!g2527) & (g2545) & (g2585)) + ((g1568) & (g1742) & (g2526) & (g2527) & (!g2545) & (!g2585)) + ((g1568) & (g1742) & (g2526) & (g2527) & (!g2545) & (g2585)) + ((g1568) & (g1742) & (g2526) & (g2527) & (g2545) & (!g2585)) + ((g1568) & (g1742) & (g2526) & (g2527) & (g2545) & (g2585)));
	assign g2618 = (((!g1742) & (!g2527) & (g2545) & (!g2585)) + ((!g1742) & (g2527) & (!g2545) & (!g2585)) + ((!g1742) & (g2527) & (!g2545) & (g2585)) + ((!g1742) & (g2527) & (g2545) & (g2585)) + ((g1742) & (!g2527) & (!g2545) & (!g2585)) + ((g1742) & (g2527) & (!g2545) & (g2585)) + ((g1742) & (g2527) & (g2545) & (!g2585)) + ((g1742) & (g2527) & (g2545) & (g2585)));
	assign g2619 = (((!g1720) & (!g1905) & (!g2529) & (g2530) & (g2544) & (!g2585)) + ((!g1720) & (!g1905) & (g2529) & (!g2530) & (!g2544) & (!g2585)) + ((!g1720) & (!g1905) & (g2529) & (!g2530) & (!g2544) & (g2585)) + ((!g1720) & (!g1905) & (g2529) & (!g2530) & (g2544) & (!g2585)) + ((!g1720) & (!g1905) & (g2529) & (!g2530) & (g2544) & (g2585)) + ((!g1720) & (!g1905) & (g2529) & (g2530) & (!g2544) & (!g2585)) + ((!g1720) & (!g1905) & (g2529) & (g2530) & (!g2544) & (g2585)) + ((!g1720) & (!g1905) & (g2529) & (g2530) & (g2544) & (g2585)) + ((!g1720) & (g1905) & (!g2529) & (!g2530) & (g2544) & (!g2585)) + ((!g1720) & (g1905) & (!g2529) & (g2530) & (!g2544) & (!g2585)) + ((!g1720) & (g1905) & (!g2529) & (g2530) & (g2544) & (!g2585)) + ((!g1720) & (g1905) & (g2529) & (!g2530) & (!g2544) & (!g2585)) + ((!g1720) & (g1905) & (g2529) & (!g2530) & (!g2544) & (g2585)) + ((!g1720) & (g1905) & (g2529) & (!g2530) & (g2544) & (g2585)) + ((!g1720) & (g1905) & (g2529) & (g2530) & (!g2544) & (g2585)) + ((!g1720) & (g1905) & (g2529) & (g2530) & (g2544) & (g2585)) + ((g1720) & (!g1905) & (!g2529) & (!g2530) & (!g2544) & (!g2585)) + ((g1720) & (!g1905) & (!g2529) & (!g2530) & (g2544) & (!g2585)) + ((g1720) & (!g1905) & (!g2529) & (g2530) & (!g2544) & (!g2585)) + ((g1720) & (!g1905) & (g2529) & (!g2530) & (!g2544) & (g2585)) + ((g1720) & (!g1905) & (g2529) & (!g2530) & (g2544) & (g2585)) + ((g1720) & (!g1905) & (g2529) & (g2530) & (!g2544) & (g2585)) + ((g1720) & (!g1905) & (g2529) & (g2530) & (g2544) & (!g2585)) + ((g1720) & (!g1905) & (g2529) & (g2530) & (g2544) & (g2585)) + ((g1720) & (g1905) & (!g2529) & (!g2530) & (!g2544) & (!g2585)) + ((g1720) & (g1905) & (g2529) & (!g2530) & (!g2544) & (g2585)) + ((g1720) & (g1905) & (g2529) & (!g2530) & (g2544) & (!g2585)) + ((g1720) & (g1905) & (g2529) & (!g2530) & (g2544) & (g2585)) + ((g1720) & (g1905) & (g2529) & (g2530) & (!g2544) & (!g2585)) + ((g1720) & (g1905) & (g2529) & (g2530) & (!g2544) & (g2585)) + ((g1720) & (g1905) & (g2529) & (g2530) & (g2544) & (!g2585)) + ((g1720) & (g1905) & (g2529) & (g2530) & (g2544) & (g2585)));
	assign g2620 = (((!g1905) & (!g2530) & (g2544) & (!g2585)) + ((!g1905) & (g2530) & (!g2544) & (!g2585)) + ((!g1905) & (g2530) & (!g2544) & (g2585)) + ((!g1905) & (g2530) & (g2544) & (g2585)) + ((g1905) & (!g2530) & (!g2544) & (!g2585)) + ((g1905) & (g2530) & (!g2544) & (g2585)) + ((g1905) & (g2530) & (g2544) & (!g2585)) + ((g1905) & (g2530) & (g2544) & (g2585)));
	assign g2621 = (((!g1879) & (!g2075) & (!g2532) & (g2533) & (g2543) & (!g2585)) + ((!g1879) & (!g2075) & (g2532) & (!g2533) & (!g2543) & (!g2585)) + ((!g1879) & (!g2075) & (g2532) & (!g2533) & (!g2543) & (g2585)) + ((!g1879) & (!g2075) & (g2532) & (!g2533) & (g2543) & (!g2585)) + ((!g1879) & (!g2075) & (g2532) & (!g2533) & (g2543) & (g2585)) + ((!g1879) & (!g2075) & (g2532) & (g2533) & (!g2543) & (!g2585)) + ((!g1879) & (!g2075) & (g2532) & (g2533) & (!g2543) & (g2585)) + ((!g1879) & (!g2075) & (g2532) & (g2533) & (g2543) & (g2585)) + ((!g1879) & (g2075) & (!g2532) & (!g2533) & (g2543) & (!g2585)) + ((!g1879) & (g2075) & (!g2532) & (g2533) & (!g2543) & (!g2585)) + ((!g1879) & (g2075) & (!g2532) & (g2533) & (g2543) & (!g2585)) + ((!g1879) & (g2075) & (g2532) & (!g2533) & (!g2543) & (!g2585)) + ((!g1879) & (g2075) & (g2532) & (!g2533) & (!g2543) & (g2585)) + ((!g1879) & (g2075) & (g2532) & (!g2533) & (g2543) & (g2585)) + ((!g1879) & (g2075) & (g2532) & (g2533) & (!g2543) & (g2585)) + ((!g1879) & (g2075) & (g2532) & (g2533) & (g2543) & (g2585)) + ((g1879) & (!g2075) & (!g2532) & (!g2533) & (!g2543) & (!g2585)) + ((g1879) & (!g2075) & (!g2532) & (!g2533) & (g2543) & (!g2585)) + ((g1879) & (!g2075) & (!g2532) & (g2533) & (!g2543) & (!g2585)) + ((g1879) & (!g2075) & (g2532) & (!g2533) & (!g2543) & (g2585)) + ((g1879) & (!g2075) & (g2532) & (!g2533) & (g2543) & (g2585)) + ((g1879) & (!g2075) & (g2532) & (g2533) & (!g2543) & (g2585)) + ((g1879) & (!g2075) & (g2532) & (g2533) & (g2543) & (!g2585)) + ((g1879) & (!g2075) & (g2532) & (g2533) & (g2543) & (g2585)) + ((g1879) & (g2075) & (!g2532) & (!g2533) & (!g2543) & (!g2585)) + ((g1879) & (g2075) & (g2532) & (!g2533) & (!g2543) & (g2585)) + ((g1879) & (g2075) & (g2532) & (!g2533) & (g2543) & (!g2585)) + ((g1879) & (g2075) & (g2532) & (!g2533) & (g2543) & (g2585)) + ((g1879) & (g2075) & (g2532) & (g2533) & (!g2543) & (!g2585)) + ((g1879) & (g2075) & (g2532) & (g2533) & (!g2543) & (g2585)) + ((g1879) & (g2075) & (g2532) & (g2533) & (g2543) & (!g2585)) + ((g1879) & (g2075) & (g2532) & (g2533) & (g2543) & (g2585)));
	assign g2622 = (((!g2075) & (!g2533) & (g2543) & (!g2585)) + ((!g2075) & (g2533) & (!g2543) & (!g2585)) + ((!g2075) & (g2533) & (!g2543) & (g2585)) + ((!g2075) & (g2533) & (g2543) & (g2585)) + ((g2075) & (!g2533) & (!g2543) & (!g2585)) + ((g2075) & (g2533) & (!g2543) & (g2585)) + ((g2075) & (g2533) & (g2543) & (!g2585)) + ((g2075) & (g2533) & (g2543) & (g2585)));
	assign g2623 = (((!g2045) & (!g2252) & (!g2535) & (g2536) & (g2542) & (!g2585)) + ((!g2045) & (!g2252) & (g2535) & (!g2536) & (!g2542) & (!g2585)) + ((!g2045) & (!g2252) & (g2535) & (!g2536) & (!g2542) & (g2585)) + ((!g2045) & (!g2252) & (g2535) & (!g2536) & (g2542) & (!g2585)) + ((!g2045) & (!g2252) & (g2535) & (!g2536) & (g2542) & (g2585)) + ((!g2045) & (!g2252) & (g2535) & (g2536) & (!g2542) & (!g2585)) + ((!g2045) & (!g2252) & (g2535) & (g2536) & (!g2542) & (g2585)) + ((!g2045) & (!g2252) & (g2535) & (g2536) & (g2542) & (g2585)) + ((!g2045) & (g2252) & (!g2535) & (!g2536) & (g2542) & (!g2585)) + ((!g2045) & (g2252) & (!g2535) & (g2536) & (!g2542) & (!g2585)) + ((!g2045) & (g2252) & (!g2535) & (g2536) & (g2542) & (!g2585)) + ((!g2045) & (g2252) & (g2535) & (!g2536) & (!g2542) & (!g2585)) + ((!g2045) & (g2252) & (g2535) & (!g2536) & (!g2542) & (g2585)) + ((!g2045) & (g2252) & (g2535) & (!g2536) & (g2542) & (g2585)) + ((!g2045) & (g2252) & (g2535) & (g2536) & (!g2542) & (g2585)) + ((!g2045) & (g2252) & (g2535) & (g2536) & (g2542) & (g2585)) + ((g2045) & (!g2252) & (!g2535) & (!g2536) & (!g2542) & (!g2585)) + ((g2045) & (!g2252) & (!g2535) & (!g2536) & (g2542) & (!g2585)) + ((g2045) & (!g2252) & (!g2535) & (g2536) & (!g2542) & (!g2585)) + ((g2045) & (!g2252) & (g2535) & (!g2536) & (!g2542) & (g2585)) + ((g2045) & (!g2252) & (g2535) & (!g2536) & (g2542) & (g2585)) + ((g2045) & (!g2252) & (g2535) & (g2536) & (!g2542) & (g2585)) + ((g2045) & (!g2252) & (g2535) & (g2536) & (g2542) & (!g2585)) + ((g2045) & (!g2252) & (g2535) & (g2536) & (g2542) & (g2585)) + ((g2045) & (g2252) & (!g2535) & (!g2536) & (!g2542) & (!g2585)) + ((g2045) & (g2252) & (g2535) & (!g2536) & (!g2542) & (g2585)) + ((g2045) & (g2252) & (g2535) & (!g2536) & (g2542) & (!g2585)) + ((g2045) & (g2252) & (g2535) & (!g2536) & (g2542) & (g2585)) + ((g2045) & (g2252) & (g2535) & (g2536) & (!g2542) & (!g2585)) + ((g2045) & (g2252) & (g2535) & (g2536) & (!g2542) & (g2585)) + ((g2045) & (g2252) & (g2535) & (g2536) & (g2542) & (!g2585)) + ((g2045) & (g2252) & (g2535) & (g2536) & (g2542) & (g2585)));
	assign g2624 = (((!g2252) & (!g2536) & (g2542) & (!g2585)) + ((!g2252) & (g2536) & (!g2542) & (!g2585)) + ((!g2252) & (g2536) & (!g2542) & (g2585)) + ((!g2252) & (g2536) & (g2542) & (g2585)) + ((g2252) & (!g2536) & (!g2542) & (!g2585)) + ((g2252) & (g2536) & (!g2542) & (g2585)) + ((g2252) & (g2536) & (g2542) & (!g2585)) + ((g2252) & (g2536) & (g2542) & (g2585)));
	assign g2625 = (((!g2218) & (!g2436) & (!g2538) & (g2539) & (g2541) & (!g2585)) + ((!g2218) & (!g2436) & (g2538) & (!g2539) & (!g2541) & (!g2585)) + ((!g2218) & (!g2436) & (g2538) & (!g2539) & (!g2541) & (g2585)) + ((!g2218) & (!g2436) & (g2538) & (!g2539) & (g2541) & (!g2585)) + ((!g2218) & (!g2436) & (g2538) & (!g2539) & (g2541) & (g2585)) + ((!g2218) & (!g2436) & (g2538) & (g2539) & (!g2541) & (!g2585)) + ((!g2218) & (!g2436) & (g2538) & (g2539) & (!g2541) & (g2585)) + ((!g2218) & (!g2436) & (g2538) & (g2539) & (g2541) & (g2585)) + ((!g2218) & (g2436) & (!g2538) & (!g2539) & (g2541) & (!g2585)) + ((!g2218) & (g2436) & (!g2538) & (g2539) & (!g2541) & (!g2585)) + ((!g2218) & (g2436) & (!g2538) & (g2539) & (g2541) & (!g2585)) + ((!g2218) & (g2436) & (g2538) & (!g2539) & (!g2541) & (!g2585)) + ((!g2218) & (g2436) & (g2538) & (!g2539) & (!g2541) & (g2585)) + ((!g2218) & (g2436) & (g2538) & (!g2539) & (g2541) & (g2585)) + ((!g2218) & (g2436) & (g2538) & (g2539) & (!g2541) & (g2585)) + ((!g2218) & (g2436) & (g2538) & (g2539) & (g2541) & (g2585)) + ((g2218) & (!g2436) & (!g2538) & (!g2539) & (!g2541) & (!g2585)) + ((g2218) & (!g2436) & (!g2538) & (!g2539) & (g2541) & (!g2585)) + ((g2218) & (!g2436) & (!g2538) & (g2539) & (!g2541) & (!g2585)) + ((g2218) & (!g2436) & (g2538) & (!g2539) & (!g2541) & (g2585)) + ((g2218) & (!g2436) & (g2538) & (!g2539) & (g2541) & (g2585)) + ((g2218) & (!g2436) & (g2538) & (g2539) & (!g2541) & (g2585)) + ((g2218) & (!g2436) & (g2538) & (g2539) & (g2541) & (!g2585)) + ((g2218) & (!g2436) & (g2538) & (g2539) & (g2541) & (g2585)) + ((g2218) & (g2436) & (!g2538) & (!g2539) & (!g2541) & (!g2585)) + ((g2218) & (g2436) & (g2538) & (!g2539) & (!g2541) & (g2585)) + ((g2218) & (g2436) & (g2538) & (!g2539) & (g2541) & (!g2585)) + ((g2218) & (g2436) & (g2538) & (!g2539) & (g2541) & (g2585)) + ((g2218) & (g2436) & (g2538) & (g2539) & (!g2541) & (!g2585)) + ((g2218) & (g2436) & (g2538) & (g2539) & (!g2541) & (g2585)) + ((g2218) & (g2436) & (g2538) & (g2539) & (g2541) & (!g2585)) + ((g2218) & (g2436) & (g2538) & (g2539) & (g2541) & (g2585)));
	assign g2626 = (((!g2436) & (!g2539) & (g2541) & (!g2585)) + ((!g2436) & (g2539) & (!g2541) & (!g2585)) + ((!g2436) & (g2539) & (!g2541) & (g2585)) + ((!g2436) & (g2539) & (g2541) & (g2585)) + ((g2436) & (!g2539) & (!g2541) & (!g2585)) + ((g2436) & (g2539) & (!g2541) & (g2585)) + ((g2436) & (g2539) & (g2541) & (!g2585)) + ((g2436) & (g2539) & (g2541) & (g2585)));
	assign g2627 = (((!g2460) & (g2478)));
	assign g2628 = (((!g2398) & (!ax22x) & (!ax23x) & (!g2627) & (!g2540) & (g2585)) + ((!g2398) & (!ax22x) & (!ax23x) & (!g2627) & (g2540) & (!g2585)) + ((!g2398) & (!ax22x) & (!ax23x) & (!g2627) & (g2540) & (g2585)) + ((!g2398) & (!ax22x) & (!ax23x) & (g2627) & (!g2540) & (!g2585)) + ((!g2398) & (!ax22x) & (ax23x) & (!g2627) & (!g2540) & (!g2585)) + ((!g2398) & (!ax22x) & (ax23x) & (g2627) & (!g2540) & (g2585)) + ((!g2398) & (!ax22x) & (ax23x) & (g2627) & (g2540) & (!g2585)) + ((!g2398) & (!ax22x) & (ax23x) & (g2627) & (g2540) & (g2585)) + ((!g2398) & (ax22x) & (!ax23x) & (g2627) & (!g2540) & (!g2585)) + ((!g2398) & (ax22x) & (!ax23x) & (g2627) & (g2540) & (!g2585)) + ((!g2398) & (ax22x) & (ax23x) & (!g2627) & (!g2540) & (!g2585)) + ((!g2398) & (ax22x) & (ax23x) & (!g2627) & (!g2540) & (g2585)) + ((!g2398) & (ax22x) & (ax23x) & (!g2627) & (g2540) & (!g2585)) + ((!g2398) & (ax22x) & (ax23x) & (!g2627) & (g2540) & (g2585)) + ((!g2398) & (ax22x) & (ax23x) & (g2627) & (!g2540) & (g2585)) + ((!g2398) & (ax22x) & (ax23x) & (g2627) & (g2540) & (g2585)) + ((g2398) & (!ax22x) & (!ax23x) & (!g2627) & (!g2540) & (!g2585)) + ((g2398) & (!ax22x) & (!ax23x) & (!g2627) & (!g2540) & (g2585)) + ((g2398) & (!ax22x) & (!ax23x) & (!g2627) & (g2540) & (g2585)) + ((g2398) & (!ax22x) & (!ax23x) & (g2627) & (g2540) & (!g2585)) + ((g2398) & (!ax22x) & (ax23x) & (!g2627) & (g2540) & (!g2585)) + ((g2398) & (!ax22x) & (ax23x) & (g2627) & (!g2540) & (!g2585)) + ((g2398) & (!ax22x) & (ax23x) & (g2627) & (!g2540) & (g2585)) + ((g2398) & (!ax22x) & (ax23x) & (g2627) & (g2540) & (g2585)) + ((g2398) & (ax22x) & (!ax23x) & (!g2627) & (!g2540) & (!g2585)) + ((g2398) & (ax22x) & (!ax23x) & (!g2627) & (g2540) & (!g2585)) + ((g2398) & (ax22x) & (ax23x) & (!g2627) & (!g2540) & (g2585)) + ((g2398) & (ax22x) & (ax23x) & (!g2627) & (g2540) & (g2585)) + ((g2398) & (ax22x) & (ax23x) & (g2627) & (!g2540) & (!g2585)) + ((g2398) & (ax22x) & (ax23x) & (g2627) & (!g2540) & (g2585)) + ((g2398) & (ax22x) & (ax23x) & (g2627) & (g2540) & (!g2585)) + ((g2398) & (ax22x) & (ax23x) & (g2627) & (g2540) & (g2585)));
	assign g2629 = (((!ax22x) & (!g2627) & (!g2540) & (g2585)) + ((!ax22x) & (!g2627) & (g2540) & (!g2585)) + ((!ax22x) & (!g2627) & (g2540) & (g2585)) + ((!ax22x) & (g2627) & (g2540) & (!g2585)) + ((ax22x) & (!g2627) & (!g2540) & (!g2585)) + ((ax22x) & (g2627) & (!g2540) & (!g2585)) + ((ax22x) & (g2627) & (!g2540) & (g2585)) + ((ax22x) & (g2627) & (g2540) & (g2585)));
	assign g2630 = (((!ax18x) & (!ax19x)));
	assign g2631 = (((!g2627) & (!ax20x) & (!ax21x) & (!g2585) & (!g2630)) + ((!g2627) & (!ax20x) & (ax21x) & (g2585) & (!g2630)) + ((!g2627) & (ax20x) & (ax21x) & (g2585) & (!g2630)) + ((!g2627) & (ax20x) & (ax21x) & (g2585) & (g2630)) + ((g2627) & (!ax20x) & (!ax21x) & (!g2585) & (!g2630)) + ((g2627) & (!ax20x) & (!ax21x) & (!g2585) & (g2630)) + ((g2627) & (!ax20x) & (!ax21x) & (g2585) & (!g2630)) + ((g2627) & (!ax20x) & (ax21x) & (!g2585) & (!g2630)) + ((g2627) & (!ax20x) & (ax21x) & (g2585) & (!g2630)) + ((g2627) & (!ax20x) & (ax21x) & (g2585) & (g2630)) + ((g2627) & (ax20x) & (!ax21x) & (g2585) & (!g2630)) + ((g2627) & (ax20x) & (!ax21x) & (g2585) & (g2630)) + ((g2627) & (ax20x) & (ax21x) & (!g2585) & (!g2630)) + ((g2627) & (ax20x) & (ax21x) & (!g2585) & (g2630)) + ((g2627) & (ax20x) & (ax21x) & (g2585) & (!g2630)) + ((g2627) & (ax20x) & (ax21x) & (g2585) & (g2630)));
	assign g2632 = (((!g2436) & (!g2398) & (g2628) & (g2629) & (g2631)) + ((!g2436) & (g2398) & (g2628) & (!g2629) & (g2631)) + ((!g2436) & (g2398) & (g2628) & (g2629) & (!g2631)) + ((!g2436) & (g2398) & (g2628) & (g2629) & (g2631)) + ((g2436) & (!g2398) & (!g2628) & (g2629) & (g2631)) + ((g2436) & (!g2398) & (g2628) & (!g2629) & (!g2631)) + ((g2436) & (!g2398) & (g2628) & (!g2629) & (g2631)) + ((g2436) & (!g2398) & (g2628) & (g2629) & (!g2631)) + ((g2436) & (!g2398) & (g2628) & (g2629) & (g2631)) + ((g2436) & (g2398) & (!g2628) & (!g2629) & (g2631)) + ((g2436) & (g2398) & (!g2628) & (g2629) & (!g2631)) + ((g2436) & (g2398) & (!g2628) & (g2629) & (g2631)) + ((g2436) & (g2398) & (g2628) & (!g2629) & (!g2631)) + ((g2436) & (g2398) & (g2628) & (!g2629) & (g2631)) + ((g2436) & (g2398) & (g2628) & (g2629) & (!g2631)) + ((g2436) & (g2398) & (g2628) & (g2629) & (g2631)));
	assign g2633 = (((!g2252) & (!g2218) & (g2625) & (g2626) & (g2632)) + ((!g2252) & (g2218) & (g2625) & (!g2626) & (g2632)) + ((!g2252) & (g2218) & (g2625) & (g2626) & (!g2632)) + ((!g2252) & (g2218) & (g2625) & (g2626) & (g2632)) + ((g2252) & (!g2218) & (!g2625) & (g2626) & (g2632)) + ((g2252) & (!g2218) & (g2625) & (!g2626) & (!g2632)) + ((g2252) & (!g2218) & (g2625) & (!g2626) & (g2632)) + ((g2252) & (!g2218) & (g2625) & (g2626) & (!g2632)) + ((g2252) & (!g2218) & (g2625) & (g2626) & (g2632)) + ((g2252) & (g2218) & (!g2625) & (!g2626) & (g2632)) + ((g2252) & (g2218) & (!g2625) & (g2626) & (!g2632)) + ((g2252) & (g2218) & (!g2625) & (g2626) & (g2632)) + ((g2252) & (g2218) & (g2625) & (!g2626) & (!g2632)) + ((g2252) & (g2218) & (g2625) & (!g2626) & (g2632)) + ((g2252) & (g2218) & (g2625) & (g2626) & (!g2632)) + ((g2252) & (g2218) & (g2625) & (g2626) & (g2632)));
	assign g2634 = (((!g2075) & (!g2045) & (g2623) & (g2624) & (g2633)) + ((!g2075) & (g2045) & (g2623) & (!g2624) & (g2633)) + ((!g2075) & (g2045) & (g2623) & (g2624) & (!g2633)) + ((!g2075) & (g2045) & (g2623) & (g2624) & (g2633)) + ((g2075) & (!g2045) & (!g2623) & (g2624) & (g2633)) + ((g2075) & (!g2045) & (g2623) & (!g2624) & (!g2633)) + ((g2075) & (!g2045) & (g2623) & (!g2624) & (g2633)) + ((g2075) & (!g2045) & (g2623) & (g2624) & (!g2633)) + ((g2075) & (!g2045) & (g2623) & (g2624) & (g2633)) + ((g2075) & (g2045) & (!g2623) & (!g2624) & (g2633)) + ((g2075) & (g2045) & (!g2623) & (g2624) & (!g2633)) + ((g2075) & (g2045) & (!g2623) & (g2624) & (g2633)) + ((g2075) & (g2045) & (g2623) & (!g2624) & (!g2633)) + ((g2075) & (g2045) & (g2623) & (!g2624) & (g2633)) + ((g2075) & (g2045) & (g2623) & (g2624) & (!g2633)) + ((g2075) & (g2045) & (g2623) & (g2624) & (g2633)));
	assign g2635 = (((!g1905) & (!g1879) & (g2621) & (g2622) & (g2634)) + ((!g1905) & (g1879) & (g2621) & (!g2622) & (g2634)) + ((!g1905) & (g1879) & (g2621) & (g2622) & (!g2634)) + ((!g1905) & (g1879) & (g2621) & (g2622) & (g2634)) + ((g1905) & (!g1879) & (!g2621) & (g2622) & (g2634)) + ((g1905) & (!g1879) & (g2621) & (!g2622) & (!g2634)) + ((g1905) & (!g1879) & (g2621) & (!g2622) & (g2634)) + ((g1905) & (!g1879) & (g2621) & (g2622) & (!g2634)) + ((g1905) & (!g1879) & (g2621) & (g2622) & (g2634)) + ((g1905) & (g1879) & (!g2621) & (!g2622) & (g2634)) + ((g1905) & (g1879) & (!g2621) & (g2622) & (!g2634)) + ((g1905) & (g1879) & (!g2621) & (g2622) & (g2634)) + ((g1905) & (g1879) & (g2621) & (!g2622) & (!g2634)) + ((g1905) & (g1879) & (g2621) & (!g2622) & (g2634)) + ((g1905) & (g1879) & (g2621) & (g2622) & (!g2634)) + ((g1905) & (g1879) & (g2621) & (g2622) & (g2634)));
	assign g2636 = (((!g1742) & (!g1720) & (g2619) & (g2620) & (g2635)) + ((!g1742) & (g1720) & (g2619) & (!g2620) & (g2635)) + ((!g1742) & (g1720) & (g2619) & (g2620) & (!g2635)) + ((!g1742) & (g1720) & (g2619) & (g2620) & (g2635)) + ((g1742) & (!g1720) & (!g2619) & (g2620) & (g2635)) + ((g1742) & (!g1720) & (g2619) & (!g2620) & (!g2635)) + ((g1742) & (!g1720) & (g2619) & (!g2620) & (g2635)) + ((g1742) & (!g1720) & (g2619) & (g2620) & (!g2635)) + ((g1742) & (!g1720) & (g2619) & (g2620) & (g2635)) + ((g1742) & (g1720) & (!g2619) & (!g2620) & (g2635)) + ((g1742) & (g1720) & (!g2619) & (g2620) & (!g2635)) + ((g1742) & (g1720) & (!g2619) & (g2620) & (g2635)) + ((g1742) & (g1720) & (g2619) & (!g2620) & (!g2635)) + ((g1742) & (g1720) & (g2619) & (!g2620) & (g2635)) + ((g1742) & (g1720) & (g2619) & (g2620) & (!g2635)) + ((g1742) & (g1720) & (g2619) & (g2620) & (g2635)));
	assign g2637 = (((!g1586) & (!g1568) & (g2617) & (g2618) & (g2636)) + ((!g1586) & (g1568) & (g2617) & (!g2618) & (g2636)) + ((!g1586) & (g1568) & (g2617) & (g2618) & (!g2636)) + ((!g1586) & (g1568) & (g2617) & (g2618) & (g2636)) + ((g1586) & (!g1568) & (!g2617) & (g2618) & (g2636)) + ((g1586) & (!g1568) & (g2617) & (!g2618) & (!g2636)) + ((g1586) & (!g1568) & (g2617) & (!g2618) & (g2636)) + ((g1586) & (!g1568) & (g2617) & (g2618) & (!g2636)) + ((g1586) & (!g1568) & (g2617) & (g2618) & (g2636)) + ((g1586) & (g1568) & (!g2617) & (!g2618) & (g2636)) + ((g1586) & (g1568) & (!g2617) & (g2618) & (!g2636)) + ((g1586) & (g1568) & (!g2617) & (g2618) & (g2636)) + ((g1586) & (g1568) & (g2617) & (!g2618) & (!g2636)) + ((g1586) & (g1568) & (g2617) & (!g2618) & (g2636)) + ((g1586) & (g1568) & (g2617) & (g2618) & (!g2636)) + ((g1586) & (g1568) & (g2617) & (g2618) & (g2636)));
	assign g2638 = (((!g1437) & (!g1423) & (g2615) & (g2616) & (g2637)) + ((!g1437) & (g1423) & (g2615) & (!g2616) & (g2637)) + ((!g1437) & (g1423) & (g2615) & (g2616) & (!g2637)) + ((!g1437) & (g1423) & (g2615) & (g2616) & (g2637)) + ((g1437) & (!g1423) & (!g2615) & (g2616) & (g2637)) + ((g1437) & (!g1423) & (g2615) & (!g2616) & (!g2637)) + ((g1437) & (!g1423) & (g2615) & (!g2616) & (g2637)) + ((g1437) & (!g1423) & (g2615) & (g2616) & (!g2637)) + ((g1437) & (!g1423) & (g2615) & (g2616) & (g2637)) + ((g1437) & (g1423) & (!g2615) & (!g2616) & (g2637)) + ((g1437) & (g1423) & (!g2615) & (g2616) & (!g2637)) + ((g1437) & (g1423) & (!g2615) & (g2616) & (g2637)) + ((g1437) & (g1423) & (g2615) & (!g2616) & (!g2637)) + ((g1437) & (g1423) & (g2615) & (!g2616) & (g2637)) + ((g1437) & (g1423) & (g2615) & (g2616) & (!g2637)) + ((g1437) & (g1423) & (g2615) & (g2616) & (g2637)));
	assign g2639 = (((!g1295) & (!g1285) & (g2613) & (g2614) & (g2638)) + ((!g1295) & (g1285) & (g2613) & (!g2614) & (g2638)) + ((!g1295) & (g1285) & (g2613) & (g2614) & (!g2638)) + ((!g1295) & (g1285) & (g2613) & (g2614) & (g2638)) + ((g1295) & (!g1285) & (!g2613) & (g2614) & (g2638)) + ((g1295) & (!g1285) & (g2613) & (!g2614) & (!g2638)) + ((g1295) & (!g1285) & (g2613) & (!g2614) & (g2638)) + ((g1295) & (!g1285) & (g2613) & (g2614) & (!g2638)) + ((g1295) & (!g1285) & (g2613) & (g2614) & (g2638)) + ((g1295) & (g1285) & (!g2613) & (!g2614) & (g2638)) + ((g1295) & (g1285) & (!g2613) & (g2614) & (!g2638)) + ((g1295) & (g1285) & (!g2613) & (g2614) & (g2638)) + ((g1295) & (g1285) & (g2613) & (!g2614) & (!g2638)) + ((g1295) & (g1285) & (g2613) & (!g2614) & (g2638)) + ((g1295) & (g1285) & (g2613) & (g2614) & (!g2638)) + ((g1295) & (g1285) & (g2613) & (g2614) & (g2638)));
	assign g2640 = (((!g1160) & (!g1154) & (g2611) & (g2612) & (g2639)) + ((!g1160) & (g1154) & (g2611) & (!g2612) & (g2639)) + ((!g1160) & (g1154) & (g2611) & (g2612) & (!g2639)) + ((!g1160) & (g1154) & (g2611) & (g2612) & (g2639)) + ((g1160) & (!g1154) & (!g2611) & (g2612) & (g2639)) + ((g1160) & (!g1154) & (g2611) & (!g2612) & (!g2639)) + ((g1160) & (!g1154) & (g2611) & (!g2612) & (g2639)) + ((g1160) & (!g1154) & (g2611) & (g2612) & (!g2639)) + ((g1160) & (!g1154) & (g2611) & (g2612) & (g2639)) + ((g1160) & (g1154) & (!g2611) & (!g2612) & (g2639)) + ((g1160) & (g1154) & (!g2611) & (g2612) & (!g2639)) + ((g1160) & (g1154) & (!g2611) & (g2612) & (g2639)) + ((g1160) & (g1154) & (g2611) & (!g2612) & (!g2639)) + ((g1160) & (g1154) & (g2611) & (!g2612) & (g2639)) + ((g1160) & (g1154) & (g2611) & (g2612) & (!g2639)) + ((g1160) & (g1154) & (g2611) & (g2612) & (g2639)));
	assign g2641 = (((!g1032) & (!g1030) & (g2609) & (g2610) & (g2640)) + ((!g1032) & (g1030) & (g2609) & (!g2610) & (g2640)) + ((!g1032) & (g1030) & (g2609) & (g2610) & (!g2640)) + ((!g1032) & (g1030) & (g2609) & (g2610) & (g2640)) + ((g1032) & (!g1030) & (!g2609) & (g2610) & (g2640)) + ((g1032) & (!g1030) & (g2609) & (!g2610) & (!g2640)) + ((g1032) & (!g1030) & (g2609) & (!g2610) & (g2640)) + ((g1032) & (!g1030) & (g2609) & (g2610) & (!g2640)) + ((g1032) & (!g1030) & (g2609) & (g2610) & (g2640)) + ((g1032) & (g1030) & (!g2609) & (!g2610) & (g2640)) + ((g1032) & (g1030) & (!g2609) & (g2610) & (!g2640)) + ((g1032) & (g1030) & (!g2609) & (g2610) & (g2640)) + ((g1032) & (g1030) & (g2609) & (!g2610) & (!g2640)) + ((g1032) & (g1030) & (g2609) & (!g2610) & (g2640)) + ((g1032) & (g1030) & (g2609) & (g2610) & (!g2640)) + ((g1032) & (g1030) & (g2609) & (g2610) & (g2640)));
	assign g2642 = (((!g851) & (!g914) & (g2607) & (g2608) & (g2641)) + ((!g851) & (g914) & (g2607) & (!g2608) & (g2641)) + ((!g851) & (g914) & (g2607) & (g2608) & (!g2641)) + ((!g851) & (g914) & (g2607) & (g2608) & (g2641)) + ((g851) & (!g914) & (!g2607) & (g2608) & (g2641)) + ((g851) & (!g914) & (g2607) & (!g2608) & (!g2641)) + ((g851) & (!g914) & (g2607) & (!g2608) & (g2641)) + ((g851) & (!g914) & (g2607) & (g2608) & (!g2641)) + ((g851) & (!g914) & (g2607) & (g2608) & (g2641)) + ((g851) & (g914) & (!g2607) & (!g2608) & (g2641)) + ((g851) & (g914) & (!g2607) & (g2608) & (!g2641)) + ((g851) & (g914) & (!g2607) & (g2608) & (g2641)) + ((g851) & (g914) & (g2607) & (!g2608) & (!g2641)) + ((g851) & (g914) & (g2607) & (!g2608) & (g2641)) + ((g851) & (g914) & (g2607) & (g2608) & (!g2641)) + ((g851) & (g914) & (g2607) & (g2608) & (g2641)));
	assign g2643 = (((!g744) & (!g803) & (g2605) & (g2606) & (g2642)) + ((!g744) & (g803) & (g2605) & (!g2606) & (g2642)) + ((!g744) & (g803) & (g2605) & (g2606) & (!g2642)) + ((!g744) & (g803) & (g2605) & (g2606) & (g2642)) + ((g744) & (!g803) & (!g2605) & (g2606) & (g2642)) + ((g744) & (!g803) & (g2605) & (!g2606) & (!g2642)) + ((g744) & (!g803) & (g2605) & (!g2606) & (g2642)) + ((g744) & (!g803) & (g2605) & (g2606) & (!g2642)) + ((g744) & (!g803) & (g2605) & (g2606) & (g2642)) + ((g744) & (g803) & (!g2605) & (!g2606) & (g2642)) + ((g744) & (g803) & (!g2605) & (g2606) & (!g2642)) + ((g744) & (g803) & (!g2605) & (g2606) & (g2642)) + ((g744) & (g803) & (g2605) & (!g2606) & (!g2642)) + ((g744) & (g803) & (g2605) & (!g2606) & (g2642)) + ((g744) & (g803) & (g2605) & (g2606) & (!g2642)) + ((g744) & (g803) & (g2605) & (g2606) & (g2642)));
	assign g2644 = (((!g645) & (!g700) & (g2603) & (g2604) & (g2643)) + ((!g645) & (g700) & (g2603) & (!g2604) & (g2643)) + ((!g645) & (g700) & (g2603) & (g2604) & (!g2643)) + ((!g645) & (g700) & (g2603) & (g2604) & (g2643)) + ((g645) & (!g700) & (!g2603) & (g2604) & (g2643)) + ((g645) & (!g700) & (g2603) & (!g2604) & (!g2643)) + ((g645) & (!g700) & (g2603) & (!g2604) & (g2643)) + ((g645) & (!g700) & (g2603) & (g2604) & (!g2643)) + ((g645) & (!g700) & (g2603) & (g2604) & (g2643)) + ((g645) & (g700) & (!g2603) & (!g2604) & (g2643)) + ((g645) & (g700) & (!g2603) & (g2604) & (!g2643)) + ((g645) & (g700) & (!g2603) & (g2604) & (g2643)) + ((g645) & (g700) & (g2603) & (!g2604) & (!g2643)) + ((g645) & (g700) & (g2603) & (!g2604) & (g2643)) + ((g645) & (g700) & (g2603) & (g2604) & (!g2643)) + ((g645) & (g700) & (g2603) & (g2604) & (g2643)));
	assign g2645 = (((!g553) & (!g604) & (g2601) & (g2602) & (g2644)) + ((!g553) & (g604) & (g2601) & (!g2602) & (g2644)) + ((!g553) & (g604) & (g2601) & (g2602) & (!g2644)) + ((!g553) & (g604) & (g2601) & (g2602) & (g2644)) + ((g553) & (!g604) & (!g2601) & (g2602) & (g2644)) + ((g553) & (!g604) & (g2601) & (!g2602) & (!g2644)) + ((g553) & (!g604) & (g2601) & (!g2602) & (g2644)) + ((g553) & (!g604) & (g2601) & (g2602) & (!g2644)) + ((g553) & (!g604) & (g2601) & (g2602) & (g2644)) + ((g553) & (g604) & (!g2601) & (!g2602) & (g2644)) + ((g553) & (g604) & (!g2601) & (g2602) & (!g2644)) + ((g553) & (g604) & (!g2601) & (g2602) & (g2644)) + ((g553) & (g604) & (g2601) & (!g2602) & (!g2644)) + ((g553) & (g604) & (g2601) & (!g2602) & (g2644)) + ((g553) & (g604) & (g2601) & (g2602) & (!g2644)) + ((g553) & (g604) & (g2601) & (g2602) & (g2644)));
	assign g2646 = (((!g468) & (!g515) & (g2599) & (g2600) & (g2645)) + ((!g468) & (g515) & (g2599) & (!g2600) & (g2645)) + ((!g468) & (g515) & (g2599) & (g2600) & (!g2645)) + ((!g468) & (g515) & (g2599) & (g2600) & (g2645)) + ((g468) & (!g515) & (!g2599) & (g2600) & (g2645)) + ((g468) & (!g515) & (g2599) & (!g2600) & (!g2645)) + ((g468) & (!g515) & (g2599) & (!g2600) & (g2645)) + ((g468) & (!g515) & (g2599) & (g2600) & (!g2645)) + ((g468) & (!g515) & (g2599) & (g2600) & (g2645)) + ((g468) & (g515) & (!g2599) & (!g2600) & (g2645)) + ((g468) & (g515) & (!g2599) & (g2600) & (!g2645)) + ((g468) & (g515) & (!g2599) & (g2600) & (g2645)) + ((g468) & (g515) & (g2599) & (!g2600) & (!g2645)) + ((g468) & (g515) & (g2599) & (!g2600) & (g2645)) + ((g468) & (g515) & (g2599) & (g2600) & (!g2645)) + ((g468) & (g515) & (g2599) & (g2600) & (g2645)));
	assign g2647 = (((!g390) & (!g433) & (g2597) & (g2598) & (g2646)) + ((!g390) & (g433) & (g2597) & (!g2598) & (g2646)) + ((!g390) & (g433) & (g2597) & (g2598) & (!g2646)) + ((!g390) & (g433) & (g2597) & (g2598) & (g2646)) + ((g390) & (!g433) & (!g2597) & (g2598) & (g2646)) + ((g390) & (!g433) & (g2597) & (!g2598) & (!g2646)) + ((g390) & (!g433) & (g2597) & (!g2598) & (g2646)) + ((g390) & (!g433) & (g2597) & (g2598) & (!g2646)) + ((g390) & (!g433) & (g2597) & (g2598) & (g2646)) + ((g390) & (g433) & (!g2597) & (!g2598) & (g2646)) + ((g390) & (g433) & (!g2597) & (g2598) & (!g2646)) + ((g390) & (g433) & (!g2597) & (g2598) & (g2646)) + ((g390) & (g433) & (g2597) & (!g2598) & (!g2646)) + ((g390) & (g433) & (g2597) & (!g2598) & (g2646)) + ((g390) & (g433) & (g2597) & (g2598) & (!g2646)) + ((g390) & (g433) & (g2597) & (g2598) & (g2646)));
	assign g2648 = (((!g319) & (!g358) & (g2595) & (g2596) & (g2647)) + ((!g319) & (g358) & (g2595) & (!g2596) & (g2647)) + ((!g319) & (g358) & (g2595) & (g2596) & (!g2647)) + ((!g319) & (g358) & (g2595) & (g2596) & (g2647)) + ((g319) & (!g358) & (!g2595) & (g2596) & (g2647)) + ((g319) & (!g358) & (g2595) & (!g2596) & (!g2647)) + ((g319) & (!g358) & (g2595) & (!g2596) & (g2647)) + ((g319) & (!g358) & (g2595) & (g2596) & (!g2647)) + ((g319) & (!g358) & (g2595) & (g2596) & (g2647)) + ((g319) & (g358) & (!g2595) & (!g2596) & (g2647)) + ((g319) & (g358) & (!g2595) & (g2596) & (!g2647)) + ((g319) & (g358) & (!g2595) & (g2596) & (g2647)) + ((g319) & (g358) & (g2595) & (!g2596) & (!g2647)) + ((g319) & (g358) & (g2595) & (!g2596) & (g2647)) + ((g319) & (g358) & (g2595) & (g2596) & (!g2647)) + ((g319) & (g358) & (g2595) & (g2596) & (g2647)));
	assign g2649 = (((!g255) & (!g290) & (g2593) & (g2594) & (g2648)) + ((!g255) & (g290) & (g2593) & (!g2594) & (g2648)) + ((!g255) & (g290) & (g2593) & (g2594) & (!g2648)) + ((!g255) & (g290) & (g2593) & (g2594) & (g2648)) + ((g255) & (!g290) & (!g2593) & (g2594) & (g2648)) + ((g255) & (!g290) & (g2593) & (!g2594) & (!g2648)) + ((g255) & (!g290) & (g2593) & (!g2594) & (g2648)) + ((g255) & (!g290) & (g2593) & (g2594) & (!g2648)) + ((g255) & (!g290) & (g2593) & (g2594) & (g2648)) + ((g255) & (g290) & (!g2593) & (!g2594) & (g2648)) + ((g255) & (g290) & (!g2593) & (g2594) & (!g2648)) + ((g255) & (g290) & (!g2593) & (g2594) & (g2648)) + ((g255) & (g290) & (g2593) & (!g2594) & (!g2648)) + ((g255) & (g290) & (g2593) & (!g2594) & (g2648)) + ((g255) & (g290) & (g2593) & (g2594) & (!g2648)) + ((g255) & (g290) & (g2593) & (g2594) & (g2648)));
	assign g2650 = (((!g198) & (!g229) & (g2591) & (g2592) & (g2649)) + ((!g198) & (g229) & (g2591) & (!g2592) & (g2649)) + ((!g198) & (g229) & (g2591) & (g2592) & (!g2649)) + ((!g198) & (g229) & (g2591) & (g2592) & (g2649)) + ((g198) & (!g229) & (!g2591) & (g2592) & (g2649)) + ((g198) & (!g229) & (g2591) & (!g2592) & (!g2649)) + ((g198) & (!g229) & (g2591) & (!g2592) & (g2649)) + ((g198) & (!g229) & (g2591) & (g2592) & (!g2649)) + ((g198) & (!g229) & (g2591) & (g2592) & (g2649)) + ((g198) & (g229) & (!g2591) & (!g2592) & (g2649)) + ((g198) & (g229) & (!g2591) & (g2592) & (!g2649)) + ((g198) & (g229) & (!g2591) & (g2592) & (g2649)) + ((g198) & (g229) & (g2591) & (!g2592) & (!g2649)) + ((g198) & (g229) & (g2591) & (!g2592) & (g2649)) + ((g198) & (g229) & (g2591) & (g2592) & (!g2649)) + ((g198) & (g229) & (g2591) & (g2592) & (g2649)));
	assign g2651 = (((!g147) & (!g174) & (g2589) & (g2590) & (g2650)) + ((!g147) & (g174) & (g2589) & (!g2590) & (g2650)) + ((!g147) & (g174) & (g2589) & (g2590) & (!g2650)) + ((!g147) & (g174) & (g2589) & (g2590) & (g2650)) + ((g147) & (!g174) & (!g2589) & (g2590) & (g2650)) + ((g147) & (!g174) & (g2589) & (!g2590) & (!g2650)) + ((g147) & (!g174) & (g2589) & (!g2590) & (g2650)) + ((g147) & (!g174) & (g2589) & (g2590) & (!g2650)) + ((g147) & (!g174) & (g2589) & (g2590) & (g2650)) + ((g147) & (g174) & (!g2589) & (!g2590) & (g2650)) + ((g147) & (g174) & (!g2589) & (g2590) & (!g2650)) + ((g147) & (g174) & (!g2589) & (g2590) & (g2650)) + ((g147) & (g174) & (g2589) & (!g2590) & (!g2650)) + ((g147) & (g174) & (g2589) & (!g2590) & (g2650)) + ((g147) & (g174) & (g2589) & (g2590) & (!g2650)) + ((g147) & (g174) & (g2589) & (g2590) & (g2650)));
	assign g2652 = (((!g104) & (!g127) & (g2587) & (g2588) & (g2651)) + ((!g104) & (g127) & (g2587) & (!g2588) & (g2651)) + ((!g104) & (g127) & (g2587) & (g2588) & (!g2651)) + ((!g104) & (g127) & (g2587) & (g2588) & (g2651)) + ((g104) & (!g127) & (!g2587) & (g2588) & (g2651)) + ((g104) & (!g127) & (g2587) & (!g2588) & (!g2651)) + ((g104) & (!g127) & (g2587) & (!g2588) & (g2651)) + ((g104) & (!g127) & (g2587) & (g2588) & (!g2651)) + ((g104) & (!g127) & (g2587) & (g2588) & (g2651)) + ((g104) & (g127) & (!g2587) & (!g2588) & (g2651)) + ((g104) & (g127) & (!g2587) & (g2588) & (!g2651)) + ((g104) & (g127) & (!g2587) & (g2588) & (g2651)) + ((g104) & (g127) & (g2587) & (!g2588) & (!g2651)) + ((g104) & (g127) & (g2587) & (!g2588) & (g2651)) + ((g104) & (g127) & (g2587) & (g2588) & (!g2651)) + ((g104) & (g127) & (g2587) & (g2588) & (g2651)));
	assign g2653 = (((g1) & (!g2562) & (g2581) & (g2584)) + ((g1) & (g2562) & (!g2581) & (!g2584)) + ((g1) & (g2562) & (!g2581) & (g2584)));
	assign g2654 = (((!g4) & (!g2) & (!g2563) & (!g2578) & (!g2580) & (!g2585)) + ((!g4) & (!g2) & (!g2563) & (!g2578) & (g2580) & (g2585)) + ((!g4) & (!g2) & (!g2563) & (g2578) & (!g2580) & (!g2585)) + ((!g4) & (!g2) & (!g2563) & (g2578) & (g2580) & (g2585)) + ((!g4) & (!g2) & (g2563) & (!g2578) & (!g2580) & (!g2585)) + ((!g4) & (!g2) & (g2563) & (!g2578) & (g2580) & (g2585)) + ((!g4) & (!g2) & (g2563) & (g2578) & (g2580) & (!g2585)) + ((!g4) & (!g2) & (g2563) & (g2578) & (g2580) & (g2585)) + ((!g4) & (g2) & (!g2563) & (!g2578) & (!g2580) & (!g2585)) + ((!g4) & (g2) & (!g2563) & (!g2578) & (g2580) & (g2585)) + ((!g4) & (g2) & (!g2563) & (g2578) & (g2580) & (!g2585)) + ((!g4) & (g2) & (!g2563) & (g2578) & (g2580) & (g2585)) + ((!g4) & (g2) & (g2563) & (!g2578) & (g2580) & (!g2585)) + ((!g4) & (g2) & (g2563) & (!g2578) & (g2580) & (g2585)) + ((!g4) & (g2) & (g2563) & (g2578) & (g2580) & (!g2585)) + ((!g4) & (g2) & (g2563) & (g2578) & (g2580) & (g2585)) + ((g4) & (!g2) & (!g2563) & (!g2578) & (g2580) & (!g2585)) + ((g4) & (!g2) & (!g2563) & (!g2578) & (g2580) & (g2585)) + ((g4) & (!g2) & (!g2563) & (g2578) & (g2580) & (!g2585)) + ((g4) & (!g2) & (!g2563) & (g2578) & (g2580) & (g2585)) + ((g4) & (!g2) & (g2563) & (!g2578) & (g2580) & (!g2585)) + ((g4) & (!g2) & (g2563) & (!g2578) & (g2580) & (g2585)) + ((g4) & (!g2) & (g2563) & (g2578) & (!g2580) & (!g2585)) + ((g4) & (!g2) & (g2563) & (g2578) & (g2580) & (g2585)) + ((g4) & (g2) & (!g2563) & (!g2578) & (g2580) & (!g2585)) + ((g4) & (g2) & (!g2563) & (!g2578) & (g2580) & (g2585)) + ((g4) & (g2) & (!g2563) & (g2578) & (!g2580) & (!g2585)) + ((g4) & (g2) & (!g2563) & (g2578) & (g2580) & (g2585)) + ((g4) & (g2) & (g2563) & (!g2578) & (!g2580) & (!g2585)) + ((g4) & (g2) & (g2563) & (!g2578) & (g2580) & (g2585)) + ((g4) & (g2) & (g2563) & (g2578) & (!g2580) & (!g2585)) + ((g4) & (g2) & (g2563) & (g2578) & (g2580) & (g2585)));
	assign g2655 = (((!g8) & (!g18) & (!g2565) & (g2566) & (g2577) & (!g2585)) + ((!g8) & (!g18) & (g2565) & (!g2566) & (!g2577) & (!g2585)) + ((!g8) & (!g18) & (g2565) & (!g2566) & (!g2577) & (g2585)) + ((!g8) & (!g18) & (g2565) & (!g2566) & (g2577) & (!g2585)) + ((!g8) & (!g18) & (g2565) & (!g2566) & (g2577) & (g2585)) + ((!g8) & (!g18) & (g2565) & (g2566) & (!g2577) & (!g2585)) + ((!g8) & (!g18) & (g2565) & (g2566) & (!g2577) & (g2585)) + ((!g8) & (!g18) & (g2565) & (g2566) & (g2577) & (g2585)) + ((!g8) & (g18) & (!g2565) & (!g2566) & (g2577) & (!g2585)) + ((!g8) & (g18) & (!g2565) & (g2566) & (!g2577) & (!g2585)) + ((!g8) & (g18) & (!g2565) & (g2566) & (g2577) & (!g2585)) + ((!g8) & (g18) & (g2565) & (!g2566) & (!g2577) & (!g2585)) + ((!g8) & (g18) & (g2565) & (!g2566) & (!g2577) & (g2585)) + ((!g8) & (g18) & (g2565) & (!g2566) & (g2577) & (g2585)) + ((!g8) & (g18) & (g2565) & (g2566) & (!g2577) & (g2585)) + ((!g8) & (g18) & (g2565) & (g2566) & (g2577) & (g2585)) + ((g8) & (!g18) & (!g2565) & (!g2566) & (!g2577) & (!g2585)) + ((g8) & (!g18) & (!g2565) & (!g2566) & (g2577) & (!g2585)) + ((g8) & (!g18) & (!g2565) & (g2566) & (!g2577) & (!g2585)) + ((g8) & (!g18) & (g2565) & (!g2566) & (!g2577) & (g2585)) + ((g8) & (!g18) & (g2565) & (!g2566) & (g2577) & (g2585)) + ((g8) & (!g18) & (g2565) & (g2566) & (!g2577) & (g2585)) + ((g8) & (!g18) & (g2565) & (g2566) & (g2577) & (!g2585)) + ((g8) & (!g18) & (g2565) & (g2566) & (g2577) & (g2585)) + ((g8) & (g18) & (!g2565) & (!g2566) & (!g2577) & (!g2585)) + ((g8) & (g18) & (g2565) & (!g2566) & (!g2577) & (g2585)) + ((g8) & (g18) & (g2565) & (!g2566) & (g2577) & (!g2585)) + ((g8) & (g18) & (g2565) & (!g2566) & (g2577) & (g2585)) + ((g8) & (g18) & (g2565) & (g2566) & (!g2577) & (!g2585)) + ((g8) & (g18) & (g2565) & (g2566) & (!g2577) & (g2585)) + ((g8) & (g18) & (g2565) & (g2566) & (g2577) & (!g2585)) + ((g8) & (g18) & (g2565) & (g2566) & (g2577) & (g2585)));
	assign g2656 = (((!g18) & (!g2566) & (g2577) & (!g2585)) + ((!g18) & (g2566) & (!g2577) & (!g2585)) + ((!g18) & (g2566) & (!g2577) & (g2585)) + ((!g18) & (g2566) & (g2577) & (g2585)) + ((g18) & (!g2566) & (!g2577) & (!g2585)) + ((g18) & (g2566) & (!g2577) & (g2585)) + ((g18) & (g2566) & (g2577) & (!g2585)) + ((g18) & (g2566) & (g2577) & (g2585)));
	assign g2657 = (((!g27) & (!g39) & (!g2568) & (g2569) & (g2576) & (!g2585)) + ((!g27) & (!g39) & (g2568) & (!g2569) & (!g2576) & (!g2585)) + ((!g27) & (!g39) & (g2568) & (!g2569) & (!g2576) & (g2585)) + ((!g27) & (!g39) & (g2568) & (!g2569) & (g2576) & (!g2585)) + ((!g27) & (!g39) & (g2568) & (!g2569) & (g2576) & (g2585)) + ((!g27) & (!g39) & (g2568) & (g2569) & (!g2576) & (!g2585)) + ((!g27) & (!g39) & (g2568) & (g2569) & (!g2576) & (g2585)) + ((!g27) & (!g39) & (g2568) & (g2569) & (g2576) & (g2585)) + ((!g27) & (g39) & (!g2568) & (!g2569) & (g2576) & (!g2585)) + ((!g27) & (g39) & (!g2568) & (g2569) & (!g2576) & (!g2585)) + ((!g27) & (g39) & (!g2568) & (g2569) & (g2576) & (!g2585)) + ((!g27) & (g39) & (g2568) & (!g2569) & (!g2576) & (!g2585)) + ((!g27) & (g39) & (g2568) & (!g2569) & (!g2576) & (g2585)) + ((!g27) & (g39) & (g2568) & (!g2569) & (g2576) & (g2585)) + ((!g27) & (g39) & (g2568) & (g2569) & (!g2576) & (g2585)) + ((!g27) & (g39) & (g2568) & (g2569) & (g2576) & (g2585)) + ((g27) & (!g39) & (!g2568) & (!g2569) & (!g2576) & (!g2585)) + ((g27) & (!g39) & (!g2568) & (!g2569) & (g2576) & (!g2585)) + ((g27) & (!g39) & (!g2568) & (g2569) & (!g2576) & (!g2585)) + ((g27) & (!g39) & (g2568) & (!g2569) & (!g2576) & (g2585)) + ((g27) & (!g39) & (g2568) & (!g2569) & (g2576) & (g2585)) + ((g27) & (!g39) & (g2568) & (g2569) & (!g2576) & (g2585)) + ((g27) & (!g39) & (g2568) & (g2569) & (g2576) & (!g2585)) + ((g27) & (!g39) & (g2568) & (g2569) & (g2576) & (g2585)) + ((g27) & (g39) & (!g2568) & (!g2569) & (!g2576) & (!g2585)) + ((g27) & (g39) & (g2568) & (!g2569) & (!g2576) & (g2585)) + ((g27) & (g39) & (g2568) & (!g2569) & (g2576) & (!g2585)) + ((g27) & (g39) & (g2568) & (!g2569) & (g2576) & (g2585)) + ((g27) & (g39) & (g2568) & (g2569) & (!g2576) & (!g2585)) + ((g27) & (g39) & (g2568) & (g2569) & (!g2576) & (g2585)) + ((g27) & (g39) & (g2568) & (g2569) & (g2576) & (!g2585)) + ((g27) & (g39) & (g2568) & (g2569) & (g2576) & (g2585)));
	assign g2658 = (((!g39) & (!g2569) & (g2576) & (!g2585)) + ((!g39) & (g2569) & (!g2576) & (!g2585)) + ((!g39) & (g2569) & (!g2576) & (g2585)) + ((!g39) & (g2569) & (g2576) & (g2585)) + ((g39) & (!g2569) & (!g2576) & (!g2585)) + ((g39) & (g2569) & (!g2576) & (g2585)) + ((g39) & (g2569) & (g2576) & (!g2585)) + ((g39) & (g2569) & (g2576) & (g2585)));
	assign g2659 = (((!g54) & (!g68) & (!g2571) & (g2572) & (g2575) & (!g2585)) + ((!g54) & (!g68) & (g2571) & (!g2572) & (!g2575) & (!g2585)) + ((!g54) & (!g68) & (g2571) & (!g2572) & (!g2575) & (g2585)) + ((!g54) & (!g68) & (g2571) & (!g2572) & (g2575) & (!g2585)) + ((!g54) & (!g68) & (g2571) & (!g2572) & (g2575) & (g2585)) + ((!g54) & (!g68) & (g2571) & (g2572) & (!g2575) & (!g2585)) + ((!g54) & (!g68) & (g2571) & (g2572) & (!g2575) & (g2585)) + ((!g54) & (!g68) & (g2571) & (g2572) & (g2575) & (g2585)) + ((!g54) & (g68) & (!g2571) & (!g2572) & (g2575) & (!g2585)) + ((!g54) & (g68) & (!g2571) & (g2572) & (!g2575) & (!g2585)) + ((!g54) & (g68) & (!g2571) & (g2572) & (g2575) & (!g2585)) + ((!g54) & (g68) & (g2571) & (!g2572) & (!g2575) & (!g2585)) + ((!g54) & (g68) & (g2571) & (!g2572) & (!g2575) & (g2585)) + ((!g54) & (g68) & (g2571) & (!g2572) & (g2575) & (g2585)) + ((!g54) & (g68) & (g2571) & (g2572) & (!g2575) & (g2585)) + ((!g54) & (g68) & (g2571) & (g2572) & (g2575) & (g2585)) + ((g54) & (!g68) & (!g2571) & (!g2572) & (!g2575) & (!g2585)) + ((g54) & (!g68) & (!g2571) & (!g2572) & (g2575) & (!g2585)) + ((g54) & (!g68) & (!g2571) & (g2572) & (!g2575) & (!g2585)) + ((g54) & (!g68) & (g2571) & (!g2572) & (!g2575) & (g2585)) + ((g54) & (!g68) & (g2571) & (!g2572) & (g2575) & (g2585)) + ((g54) & (!g68) & (g2571) & (g2572) & (!g2575) & (g2585)) + ((g54) & (!g68) & (g2571) & (g2572) & (g2575) & (!g2585)) + ((g54) & (!g68) & (g2571) & (g2572) & (g2575) & (g2585)) + ((g54) & (g68) & (!g2571) & (!g2572) & (!g2575) & (!g2585)) + ((g54) & (g68) & (g2571) & (!g2572) & (!g2575) & (g2585)) + ((g54) & (g68) & (g2571) & (!g2572) & (g2575) & (!g2585)) + ((g54) & (g68) & (g2571) & (!g2572) & (g2575) & (g2585)) + ((g54) & (g68) & (g2571) & (g2572) & (!g2575) & (!g2585)) + ((g54) & (g68) & (g2571) & (g2572) & (!g2575) & (g2585)) + ((g54) & (g68) & (g2571) & (g2572) & (g2575) & (!g2585)) + ((g54) & (g68) & (g2571) & (g2572) & (g2575) & (g2585)));
	assign g2660 = (((!g68) & (!g2572) & (g2575) & (!g2585)) + ((!g68) & (g2572) & (!g2575) & (!g2585)) + ((!g68) & (g2572) & (!g2575) & (g2585)) + ((!g68) & (g2572) & (g2575) & (g2585)) + ((g68) & (!g2572) & (!g2575) & (!g2585)) + ((g68) & (g2572) & (!g2575) & (g2585)) + ((g68) & (g2572) & (g2575) & (!g2585)) + ((g68) & (g2572) & (g2575) & (g2585)));
	assign g2661 = (((!g87) & (!g104) & (!g2574) & (g2479) & (g2561) & (!g2585)) + ((!g87) & (!g104) & (g2574) & (!g2479) & (!g2561) & (!g2585)) + ((!g87) & (!g104) & (g2574) & (!g2479) & (!g2561) & (g2585)) + ((!g87) & (!g104) & (g2574) & (!g2479) & (g2561) & (!g2585)) + ((!g87) & (!g104) & (g2574) & (!g2479) & (g2561) & (g2585)) + ((!g87) & (!g104) & (g2574) & (g2479) & (!g2561) & (!g2585)) + ((!g87) & (!g104) & (g2574) & (g2479) & (!g2561) & (g2585)) + ((!g87) & (!g104) & (g2574) & (g2479) & (g2561) & (g2585)) + ((!g87) & (g104) & (!g2574) & (!g2479) & (g2561) & (!g2585)) + ((!g87) & (g104) & (!g2574) & (g2479) & (!g2561) & (!g2585)) + ((!g87) & (g104) & (!g2574) & (g2479) & (g2561) & (!g2585)) + ((!g87) & (g104) & (g2574) & (!g2479) & (!g2561) & (!g2585)) + ((!g87) & (g104) & (g2574) & (!g2479) & (!g2561) & (g2585)) + ((!g87) & (g104) & (g2574) & (!g2479) & (g2561) & (g2585)) + ((!g87) & (g104) & (g2574) & (g2479) & (!g2561) & (g2585)) + ((!g87) & (g104) & (g2574) & (g2479) & (g2561) & (g2585)) + ((g87) & (!g104) & (!g2574) & (!g2479) & (!g2561) & (!g2585)) + ((g87) & (!g104) & (!g2574) & (!g2479) & (g2561) & (!g2585)) + ((g87) & (!g104) & (!g2574) & (g2479) & (!g2561) & (!g2585)) + ((g87) & (!g104) & (g2574) & (!g2479) & (!g2561) & (g2585)) + ((g87) & (!g104) & (g2574) & (!g2479) & (g2561) & (g2585)) + ((g87) & (!g104) & (g2574) & (g2479) & (!g2561) & (g2585)) + ((g87) & (!g104) & (g2574) & (g2479) & (g2561) & (!g2585)) + ((g87) & (!g104) & (g2574) & (g2479) & (g2561) & (g2585)) + ((g87) & (g104) & (!g2574) & (!g2479) & (!g2561) & (!g2585)) + ((g87) & (g104) & (g2574) & (!g2479) & (!g2561) & (g2585)) + ((g87) & (g104) & (g2574) & (!g2479) & (g2561) & (!g2585)) + ((g87) & (g104) & (g2574) & (!g2479) & (g2561) & (g2585)) + ((g87) & (g104) & (g2574) & (g2479) & (!g2561) & (!g2585)) + ((g87) & (g104) & (g2574) & (g2479) & (!g2561) & (g2585)) + ((g87) & (g104) & (g2574) & (g2479) & (g2561) & (!g2585)) + ((g87) & (g104) & (g2574) & (g2479) & (g2561) & (g2585)));
	assign g2662 = (((!g68) & (!g87) & (g2661) & (g2586) & (g2652)) + ((!g68) & (g87) & (g2661) & (!g2586) & (g2652)) + ((!g68) & (g87) & (g2661) & (g2586) & (!g2652)) + ((!g68) & (g87) & (g2661) & (g2586) & (g2652)) + ((g68) & (!g87) & (!g2661) & (g2586) & (g2652)) + ((g68) & (!g87) & (g2661) & (!g2586) & (!g2652)) + ((g68) & (!g87) & (g2661) & (!g2586) & (g2652)) + ((g68) & (!g87) & (g2661) & (g2586) & (!g2652)) + ((g68) & (!g87) & (g2661) & (g2586) & (g2652)) + ((g68) & (g87) & (!g2661) & (!g2586) & (g2652)) + ((g68) & (g87) & (!g2661) & (g2586) & (!g2652)) + ((g68) & (g87) & (!g2661) & (g2586) & (g2652)) + ((g68) & (g87) & (g2661) & (!g2586) & (!g2652)) + ((g68) & (g87) & (g2661) & (!g2586) & (g2652)) + ((g68) & (g87) & (g2661) & (g2586) & (!g2652)) + ((g68) & (g87) & (g2661) & (g2586) & (g2652)));
	assign g2663 = (((!g39) & (!g54) & (g2659) & (g2660) & (g2662)) + ((!g39) & (g54) & (g2659) & (!g2660) & (g2662)) + ((!g39) & (g54) & (g2659) & (g2660) & (!g2662)) + ((!g39) & (g54) & (g2659) & (g2660) & (g2662)) + ((g39) & (!g54) & (!g2659) & (g2660) & (g2662)) + ((g39) & (!g54) & (g2659) & (!g2660) & (!g2662)) + ((g39) & (!g54) & (g2659) & (!g2660) & (g2662)) + ((g39) & (!g54) & (g2659) & (g2660) & (!g2662)) + ((g39) & (!g54) & (g2659) & (g2660) & (g2662)) + ((g39) & (g54) & (!g2659) & (!g2660) & (g2662)) + ((g39) & (g54) & (!g2659) & (g2660) & (!g2662)) + ((g39) & (g54) & (!g2659) & (g2660) & (g2662)) + ((g39) & (g54) & (g2659) & (!g2660) & (!g2662)) + ((g39) & (g54) & (g2659) & (!g2660) & (g2662)) + ((g39) & (g54) & (g2659) & (g2660) & (!g2662)) + ((g39) & (g54) & (g2659) & (g2660) & (g2662)));
	assign g2664 = (((!g18) & (!g27) & (g2657) & (g2658) & (g2663)) + ((!g18) & (g27) & (g2657) & (!g2658) & (g2663)) + ((!g18) & (g27) & (g2657) & (g2658) & (!g2663)) + ((!g18) & (g27) & (g2657) & (g2658) & (g2663)) + ((g18) & (!g27) & (!g2657) & (g2658) & (g2663)) + ((g18) & (!g27) & (g2657) & (!g2658) & (!g2663)) + ((g18) & (!g27) & (g2657) & (!g2658) & (g2663)) + ((g18) & (!g27) & (g2657) & (g2658) & (!g2663)) + ((g18) & (!g27) & (g2657) & (g2658) & (g2663)) + ((g18) & (g27) & (!g2657) & (!g2658) & (g2663)) + ((g18) & (g27) & (!g2657) & (g2658) & (!g2663)) + ((g18) & (g27) & (!g2657) & (g2658) & (g2663)) + ((g18) & (g27) & (g2657) & (!g2658) & (!g2663)) + ((g18) & (g27) & (g2657) & (!g2658) & (g2663)) + ((g18) & (g27) & (g2657) & (g2658) & (!g2663)) + ((g18) & (g27) & (g2657) & (g2658) & (g2663)));
	assign g2665 = (((!g2) & (!g8) & (g2655) & (g2656) & (g2664)) + ((!g2) & (g8) & (g2655) & (!g2656) & (g2664)) + ((!g2) & (g8) & (g2655) & (g2656) & (!g2664)) + ((!g2) & (g8) & (g2655) & (g2656) & (g2664)) + ((g2) & (!g8) & (!g2655) & (g2656) & (g2664)) + ((g2) & (!g8) & (g2655) & (!g2656) & (!g2664)) + ((g2) & (!g8) & (g2655) & (!g2656) & (g2664)) + ((g2) & (!g8) & (g2655) & (g2656) & (!g2664)) + ((g2) & (!g8) & (g2655) & (g2656) & (g2664)) + ((g2) & (g8) & (!g2655) & (!g2656) & (g2664)) + ((g2) & (g8) & (!g2655) & (g2656) & (!g2664)) + ((g2) & (g8) & (!g2655) & (g2656) & (g2664)) + ((g2) & (g8) & (g2655) & (!g2656) & (!g2664)) + ((g2) & (g8) & (g2655) & (!g2656) & (g2664)) + ((g2) & (g8) & (g2655) & (g2656) & (!g2664)) + ((g2) & (g8) & (g2655) & (g2656) & (g2664)));
	assign g2666 = (((!g2) & (!g2563) & (g2578) & (!g2585)) + ((!g2) & (g2563) & (!g2578) & (!g2585)) + ((!g2) & (g2563) & (!g2578) & (g2585)) + ((!g2) & (g2563) & (g2578) & (g2585)) + ((g2) & (!g2563) & (!g2578) & (!g2585)) + ((g2) & (g2563) & (!g2578) & (g2585)) + ((g2) & (g2563) & (g2578) & (!g2585)) + ((g2) & (g2563) & (g2578) & (g2585)));
	assign g2667 = (((!g1) & (!g2562) & (!g2581) & (!g2583) & (g2584)) + ((!g1) & (!g2562) & (!g2581) & (g2583) & (!g2584)) + ((!g1) & (!g2562) & (!g2581) & (g2583) & (g2584)) + ((!g1) & (g2562) & (g2581) & (!g2583) & (!g2584)) + ((!g1) & (g2562) & (g2581) & (!g2583) & (g2584)) + ((!g1) & (g2562) & (g2581) & (g2583) & (!g2584)) + ((!g1) & (g2562) & (g2581) & (g2583) & (g2584)) + ((g1) & (!g2562) & (!g2581) & (!g2583) & (g2584)) + ((g1) & (!g2562) & (!g2581) & (g2583) & (g2584)) + ((g1) & (g2562) & (g2581) & (!g2583) & (!g2584)) + ((g1) & (g2562) & (g2581) & (!g2583) & (g2584)) + ((g1) & (g2562) & (g2581) & (g2583) & (!g2584)) + ((g1) & (g2562) & (g2581) & (g2583) & (g2584)));
	assign g2668 = (((!g4) & (!g1) & (!g2654) & (!g2665) & (!g2666) & (!g2667)) + ((!g4) & (g1) & (!g2654) & (!g2665) & (!g2666) & (!g2667)) + ((!g4) & (g1) & (!g2654) & (!g2665) & (!g2666) & (g2667)) + ((!g4) & (g1) & (!g2654) & (!g2665) & (g2666) & (!g2667)) + ((!g4) & (g1) & (!g2654) & (!g2665) & (g2666) & (g2667)) + ((!g4) & (g1) & (!g2654) & (g2665) & (!g2666) & (!g2667)) + ((!g4) & (g1) & (!g2654) & (g2665) & (!g2666) & (g2667)) + ((!g4) & (g1) & (!g2654) & (g2665) & (g2666) & (!g2667)) + ((!g4) & (g1) & (!g2654) & (g2665) & (g2666) & (g2667)) + ((!g4) & (g1) & (g2654) & (!g2665) & (!g2666) & (!g2667)) + ((!g4) & (g1) & (g2654) & (!g2665) & (!g2666) & (g2667)) + ((g4) & (!g1) & (!g2654) & (!g2665) & (!g2666) & (!g2667)) + ((g4) & (!g1) & (!g2654) & (!g2665) & (g2666) & (!g2667)) + ((g4) & (!g1) & (!g2654) & (g2665) & (!g2666) & (!g2667)) + ((g4) & (g1) & (!g2654) & (!g2665) & (!g2666) & (!g2667)) + ((g4) & (g1) & (!g2654) & (!g2665) & (!g2666) & (g2667)) + ((g4) & (g1) & (!g2654) & (!g2665) & (g2666) & (!g2667)) + ((g4) & (g1) & (!g2654) & (!g2665) & (g2666) & (g2667)) + ((g4) & (g1) & (!g2654) & (g2665) & (!g2666) & (!g2667)) + ((g4) & (g1) & (!g2654) & (g2665) & (!g2666) & (g2667)) + ((g4) & (g1) & (!g2654) & (g2665) & (g2666) & (!g2667)) + ((g4) & (g1) & (!g2654) & (g2665) & (g2666) & (g2667)) + ((g4) & (g1) & (g2654) & (!g2665) & (!g2666) & (!g2667)) + ((g4) & (g1) & (g2654) & (!g2665) & (!g2666) & (g2667)) + ((g4) & (g1) & (g2654) & (!g2665) & (g2666) & (!g2667)) + ((g4) & (g1) & (g2654) & (!g2665) & (g2666) & (g2667)) + ((g4) & (g1) & (g2654) & (g2665) & (!g2666) & (!g2667)) + ((g4) & (g1) & (g2654) & (g2665) & (!g2666) & (g2667)));
	assign g2669 = (((!g87) & (!g2586) & (g2652) & (!g2653) & (!g2668)) + ((!g87) & (!g2586) & (g2652) & (g2653) & (!g2668)) + ((!g87) & (!g2586) & (g2652) & (g2653) & (g2668)) + ((!g87) & (g2586) & (!g2652) & (!g2653) & (!g2668)) + ((!g87) & (g2586) & (!g2652) & (!g2653) & (g2668)) + ((!g87) & (g2586) & (!g2652) & (g2653) & (!g2668)) + ((!g87) & (g2586) & (!g2652) & (g2653) & (g2668)) + ((!g87) & (g2586) & (g2652) & (!g2653) & (g2668)) + ((g87) & (!g2586) & (!g2652) & (!g2653) & (!g2668)) + ((g87) & (!g2586) & (!g2652) & (g2653) & (!g2668)) + ((g87) & (!g2586) & (!g2652) & (g2653) & (g2668)) + ((g87) & (g2586) & (!g2652) & (!g2653) & (g2668)) + ((g87) & (g2586) & (g2652) & (!g2653) & (!g2668)) + ((g87) & (g2586) & (g2652) & (!g2653) & (g2668)) + ((g87) & (g2586) & (g2652) & (g2653) & (!g2668)) + ((g87) & (g2586) & (g2652) & (g2653) & (g2668)));
	assign g2670 = (((!g104) & (!g127) & (g2588) & (g2651)) + ((!g104) & (g127) & (!g2588) & (g2651)) + ((!g104) & (g127) & (g2588) & (!g2651)) + ((!g104) & (g127) & (g2588) & (g2651)) + ((g104) & (!g127) & (!g2588) & (!g2651)) + ((g104) & (!g127) & (!g2588) & (g2651)) + ((g104) & (!g127) & (g2588) & (!g2651)) + ((g104) & (g127) & (!g2588) & (!g2651)));
	assign g2671 = (((!g2587) & (!g2653) & (!g2668) & (g2670)) + ((!g2587) & (g2653) & (!g2668) & (g2670)) + ((!g2587) & (g2653) & (g2668) & (g2670)) + ((g2587) & (!g2653) & (!g2668) & (!g2670)) + ((g2587) & (!g2653) & (g2668) & (!g2670)) + ((g2587) & (!g2653) & (g2668) & (g2670)) + ((g2587) & (g2653) & (!g2668) & (!g2670)) + ((g2587) & (g2653) & (g2668) & (!g2670)));
	assign g2672 = (((!g127) & (!g2588) & (g2651) & (!g2653) & (!g2668)) + ((!g127) & (!g2588) & (g2651) & (g2653) & (!g2668)) + ((!g127) & (!g2588) & (g2651) & (g2653) & (g2668)) + ((!g127) & (g2588) & (!g2651) & (!g2653) & (!g2668)) + ((!g127) & (g2588) & (!g2651) & (!g2653) & (g2668)) + ((!g127) & (g2588) & (!g2651) & (g2653) & (!g2668)) + ((!g127) & (g2588) & (!g2651) & (g2653) & (g2668)) + ((!g127) & (g2588) & (g2651) & (!g2653) & (g2668)) + ((g127) & (!g2588) & (!g2651) & (!g2653) & (!g2668)) + ((g127) & (!g2588) & (!g2651) & (g2653) & (!g2668)) + ((g127) & (!g2588) & (!g2651) & (g2653) & (g2668)) + ((g127) & (g2588) & (!g2651) & (!g2653) & (g2668)) + ((g127) & (g2588) & (g2651) & (!g2653) & (!g2668)) + ((g127) & (g2588) & (g2651) & (!g2653) & (g2668)) + ((g127) & (g2588) & (g2651) & (g2653) & (!g2668)) + ((g127) & (g2588) & (g2651) & (g2653) & (g2668)));
	assign g2673 = (((!g147) & (!g174) & (g2590) & (g2650)) + ((!g147) & (g174) & (!g2590) & (g2650)) + ((!g147) & (g174) & (g2590) & (!g2650)) + ((!g147) & (g174) & (g2590) & (g2650)) + ((g147) & (!g174) & (!g2590) & (!g2650)) + ((g147) & (!g174) & (!g2590) & (g2650)) + ((g147) & (!g174) & (g2590) & (!g2650)) + ((g147) & (g174) & (!g2590) & (!g2650)));
	assign g2674 = (((!g2589) & (!g2653) & (!g2668) & (g2673)) + ((!g2589) & (g2653) & (!g2668) & (g2673)) + ((!g2589) & (g2653) & (g2668) & (g2673)) + ((g2589) & (!g2653) & (!g2668) & (!g2673)) + ((g2589) & (!g2653) & (g2668) & (!g2673)) + ((g2589) & (!g2653) & (g2668) & (g2673)) + ((g2589) & (g2653) & (!g2668) & (!g2673)) + ((g2589) & (g2653) & (g2668) & (!g2673)));
	assign g2675 = (((!g174) & (!g2590) & (g2650) & (!g2653) & (!g2668)) + ((!g174) & (!g2590) & (g2650) & (g2653) & (!g2668)) + ((!g174) & (!g2590) & (g2650) & (g2653) & (g2668)) + ((!g174) & (g2590) & (!g2650) & (!g2653) & (!g2668)) + ((!g174) & (g2590) & (!g2650) & (!g2653) & (g2668)) + ((!g174) & (g2590) & (!g2650) & (g2653) & (!g2668)) + ((!g174) & (g2590) & (!g2650) & (g2653) & (g2668)) + ((!g174) & (g2590) & (g2650) & (!g2653) & (g2668)) + ((g174) & (!g2590) & (!g2650) & (!g2653) & (!g2668)) + ((g174) & (!g2590) & (!g2650) & (g2653) & (!g2668)) + ((g174) & (!g2590) & (!g2650) & (g2653) & (g2668)) + ((g174) & (g2590) & (!g2650) & (!g2653) & (g2668)) + ((g174) & (g2590) & (g2650) & (!g2653) & (!g2668)) + ((g174) & (g2590) & (g2650) & (!g2653) & (g2668)) + ((g174) & (g2590) & (g2650) & (g2653) & (!g2668)) + ((g174) & (g2590) & (g2650) & (g2653) & (g2668)));
	assign g2676 = (((!g198) & (!g229) & (g2592) & (g2649)) + ((!g198) & (g229) & (!g2592) & (g2649)) + ((!g198) & (g229) & (g2592) & (!g2649)) + ((!g198) & (g229) & (g2592) & (g2649)) + ((g198) & (!g229) & (!g2592) & (!g2649)) + ((g198) & (!g229) & (!g2592) & (g2649)) + ((g198) & (!g229) & (g2592) & (!g2649)) + ((g198) & (g229) & (!g2592) & (!g2649)));
	assign g2677 = (((!g2591) & (!g2653) & (!g2668) & (g2676)) + ((!g2591) & (g2653) & (!g2668) & (g2676)) + ((!g2591) & (g2653) & (g2668) & (g2676)) + ((g2591) & (!g2653) & (!g2668) & (!g2676)) + ((g2591) & (!g2653) & (g2668) & (!g2676)) + ((g2591) & (!g2653) & (g2668) & (g2676)) + ((g2591) & (g2653) & (!g2668) & (!g2676)) + ((g2591) & (g2653) & (g2668) & (!g2676)));
	assign g2678 = (((!g229) & (!g2592) & (g2649) & (!g2653) & (!g2668)) + ((!g229) & (!g2592) & (g2649) & (g2653) & (!g2668)) + ((!g229) & (!g2592) & (g2649) & (g2653) & (g2668)) + ((!g229) & (g2592) & (!g2649) & (!g2653) & (!g2668)) + ((!g229) & (g2592) & (!g2649) & (!g2653) & (g2668)) + ((!g229) & (g2592) & (!g2649) & (g2653) & (!g2668)) + ((!g229) & (g2592) & (!g2649) & (g2653) & (g2668)) + ((!g229) & (g2592) & (g2649) & (!g2653) & (g2668)) + ((g229) & (!g2592) & (!g2649) & (!g2653) & (!g2668)) + ((g229) & (!g2592) & (!g2649) & (g2653) & (!g2668)) + ((g229) & (!g2592) & (!g2649) & (g2653) & (g2668)) + ((g229) & (g2592) & (!g2649) & (!g2653) & (g2668)) + ((g229) & (g2592) & (g2649) & (!g2653) & (!g2668)) + ((g229) & (g2592) & (g2649) & (!g2653) & (g2668)) + ((g229) & (g2592) & (g2649) & (g2653) & (!g2668)) + ((g229) & (g2592) & (g2649) & (g2653) & (g2668)));
	assign g2679 = (((!g255) & (!g290) & (g2594) & (g2648)) + ((!g255) & (g290) & (!g2594) & (g2648)) + ((!g255) & (g290) & (g2594) & (!g2648)) + ((!g255) & (g290) & (g2594) & (g2648)) + ((g255) & (!g290) & (!g2594) & (!g2648)) + ((g255) & (!g290) & (!g2594) & (g2648)) + ((g255) & (!g290) & (g2594) & (!g2648)) + ((g255) & (g290) & (!g2594) & (!g2648)));
	assign g2680 = (((!g2593) & (!g2653) & (!g2668) & (g2679)) + ((!g2593) & (g2653) & (!g2668) & (g2679)) + ((!g2593) & (g2653) & (g2668) & (g2679)) + ((g2593) & (!g2653) & (!g2668) & (!g2679)) + ((g2593) & (!g2653) & (g2668) & (!g2679)) + ((g2593) & (!g2653) & (g2668) & (g2679)) + ((g2593) & (g2653) & (!g2668) & (!g2679)) + ((g2593) & (g2653) & (g2668) & (!g2679)));
	assign g2681 = (((!g290) & (!g2594) & (g2648) & (!g2653) & (!g2668)) + ((!g290) & (!g2594) & (g2648) & (g2653) & (!g2668)) + ((!g290) & (!g2594) & (g2648) & (g2653) & (g2668)) + ((!g290) & (g2594) & (!g2648) & (!g2653) & (!g2668)) + ((!g290) & (g2594) & (!g2648) & (!g2653) & (g2668)) + ((!g290) & (g2594) & (!g2648) & (g2653) & (!g2668)) + ((!g290) & (g2594) & (!g2648) & (g2653) & (g2668)) + ((!g290) & (g2594) & (g2648) & (!g2653) & (g2668)) + ((g290) & (!g2594) & (!g2648) & (!g2653) & (!g2668)) + ((g290) & (!g2594) & (!g2648) & (g2653) & (!g2668)) + ((g290) & (!g2594) & (!g2648) & (g2653) & (g2668)) + ((g290) & (g2594) & (!g2648) & (!g2653) & (g2668)) + ((g290) & (g2594) & (g2648) & (!g2653) & (!g2668)) + ((g290) & (g2594) & (g2648) & (!g2653) & (g2668)) + ((g290) & (g2594) & (g2648) & (g2653) & (!g2668)) + ((g290) & (g2594) & (g2648) & (g2653) & (g2668)));
	assign g2682 = (((!g319) & (!g358) & (g2596) & (g2647)) + ((!g319) & (g358) & (!g2596) & (g2647)) + ((!g319) & (g358) & (g2596) & (!g2647)) + ((!g319) & (g358) & (g2596) & (g2647)) + ((g319) & (!g358) & (!g2596) & (!g2647)) + ((g319) & (!g358) & (!g2596) & (g2647)) + ((g319) & (!g358) & (g2596) & (!g2647)) + ((g319) & (g358) & (!g2596) & (!g2647)));
	assign g2683 = (((!g2595) & (!g2653) & (!g2668) & (g2682)) + ((!g2595) & (g2653) & (!g2668) & (g2682)) + ((!g2595) & (g2653) & (g2668) & (g2682)) + ((g2595) & (!g2653) & (!g2668) & (!g2682)) + ((g2595) & (!g2653) & (g2668) & (!g2682)) + ((g2595) & (!g2653) & (g2668) & (g2682)) + ((g2595) & (g2653) & (!g2668) & (!g2682)) + ((g2595) & (g2653) & (g2668) & (!g2682)));
	assign g2684 = (((!g358) & (!g2596) & (g2647) & (!g2653) & (!g2668)) + ((!g358) & (!g2596) & (g2647) & (g2653) & (!g2668)) + ((!g358) & (!g2596) & (g2647) & (g2653) & (g2668)) + ((!g358) & (g2596) & (!g2647) & (!g2653) & (!g2668)) + ((!g358) & (g2596) & (!g2647) & (!g2653) & (g2668)) + ((!g358) & (g2596) & (!g2647) & (g2653) & (!g2668)) + ((!g358) & (g2596) & (!g2647) & (g2653) & (g2668)) + ((!g358) & (g2596) & (g2647) & (!g2653) & (g2668)) + ((g358) & (!g2596) & (!g2647) & (!g2653) & (!g2668)) + ((g358) & (!g2596) & (!g2647) & (g2653) & (!g2668)) + ((g358) & (!g2596) & (!g2647) & (g2653) & (g2668)) + ((g358) & (g2596) & (!g2647) & (!g2653) & (g2668)) + ((g358) & (g2596) & (g2647) & (!g2653) & (!g2668)) + ((g358) & (g2596) & (g2647) & (!g2653) & (g2668)) + ((g358) & (g2596) & (g2647) & (g2653) & (!g2668)) + ((g358) & (g2596) & (g2647) & (g2653) & (g2668)));
	assign g2685 = (((!g390) & (!g433) & (g2598) & (g2646)) + ((!g390) & (g433) & (!g2598) & (g2646)) + ((!g390) & (g433) & (g2598) & (!g2646)) + ((!g390) & (g433) & (g2598) & (g2646)) + ((g390) & (!g433) & (!g2598) & (!g2646)) + ((g390) & (!g433) & (!g2598) & (g2646)) + ((g390) & (!g433) & (g2598) & (!g2646)) + ((g390) & (g433) & (!g2598) & (!g2646)));
	assign g2686 = (((!g2597) & (!g2653) & (!g2668) & (g2685)) + ((!g2597) & (g2653) & (!g2668) & (g2685)) + ((!g2597) & (g2653) & (g2668) & (g2685)) + ((g2597) & (!g2653) & (!g2668) & (!g2685)) + ((g2597) & (!g2653) & (g2668) & (!g2685)) + ((g2597) & (!g2653) & (g2668) & (g2685)) + ((g2597) & (g2653) & (!g2668) & (!g2685)) + ((g2597) & (g2653) & (g2668) & (!g2685)));
	assign g2687 = (((!g433) & (!g2598) & (g2646) & (!g2653) & (!g2668)) + ((!g433) & (!g2598) & (g2646) & (g2653) & (!g2668)) + ((!g433) & (!g2598) & (g2646) & (g2653) & (g2668)) + ((!g433) & (g2598) & (!g2646) & (!g2653) & (!g2668)) + ((!g433) & (g2598) & (!g2646) & (!g2653) & (g2668)) + ((!g433) & (g2598) & (!g2646) & (g2653) & (!g2668)) + ((!g433) & (g2598) & (!g2646) & (g2653) & (g2668)) + ((!g433) & (g2598) & (g2646) & (!g2653) & (g2668)) + ((g433) & (!g2598) & (!g2646) & (!g2653) & (!g2668)) + ((g433) & (!g2598) & (!g2646) & (g2653) & (!g2668)) + ((g433) & (!g2598) & (!g2646) & (g2653) & (g2668)) + ((g433) & (g2598) & (!g2646) & (!g2653) & (g2668)) + ((g433) & (g2598) & (g2646) & (!g2653) & (!g2668)) + ((g433) & (g2598) & (g2646) & (!g2653) & (g2668)) + ((g433) & (g2598) & (g2646) & (g2653) & (!g2668)) + ((g433) & (g2598) & (g2646) & (g2653) & (g2668)));
	assign g2688 = (((!g468) & (!g515) & (g2600) & (g2645)) + ((!g468) & (g515) & (!g2600) & (g2645)) + ((!g468) & (g515) & (g2600) & (!g2645)) + ((!g468) & (g515) & (g2600) & (g2645)) + ((g468) & (!g515) & (!g2600) & (!g2645)) + ((g468) & (!g515) & (!g2600) & (g2645)) + ((g468) & (!g515) & (g2600) & (!g2645)) + ((g468) & (g515) & (!g2600) & (!g2645)));
	assign g2689 = (((!g2599) & (!g2653) & (!g2668) & (g2688)) + ((!g2599) & (g2653) & (!g2668) & (g2688)) + ((!g2599) & (g2653) & (g2668) & (g2688)) + ((g2599) & (!g2653) & (!g2668) & (!g2688)) + ((g2599) & (!g2653) & (g2668) & (!g2688)) + ((g2599) & (!g2653) & (g2668) & (g2688)) + ((g2599) & (g2653) & (!g2668) & (!g2688)) + ((g2599) & (g2653) & (g2668) & (!g2688)));
	assign g2690 = (((!g515) & (!g2600) & (g2645) & (!g2653) & (!g2668)) + ((!g515) & (!g2600) & (g2645) & (g2653) & (!g2668)) + ((!g515) & (!g2600) & (g2645) & (g2653) & (g2668)) + ((!g515) & (g2600) & (!g2645) & (!g2653) & (!g2668)) + ((!g515) & (g2600) & (!g2645) & (!g2653) & (g2668)) + ((!g515) & (g2600) & (!g2645) & (g2653) & (!g2668)) + ((!g515) & (g2600) & (!g2645) & (g2653) & (g2668)) + ((!g515) & (g2600) & (g2645) & (!g2653) & (g2668)) + ((g515) & (!g2600) & (!g2645) & (!g2653) & (!g2668)) + ((g515) & (!g2600) & (!g2645) & (g2653) & (!g2668)) + ((g515) & (!g2600) & (!g2645) & (g2653) & (g2668)) + ((g515) & (g2600) & (!g2645) & (!g2653) & (g2668)) + ((g515) & (g2600) & (g2645) & (!g2653) & (!g2668)) + ((g515) & (g2600) & (g2645) & (!g2653) & (g2668)) + ((g515) & (g2600) & (g2645) & (g2653) & (!g2668)) + ((g515) & (g2600) & (g2645) & (g2653) & (g2668)));
	assign g2691 = (((!g553) & (!g604) & (g2602) & (g2644)) + ((!g553) & (g604) & (!g2602) & (g2644)) + ((!g553) & (g604) & (g2602) & (!g2644)) + ((!g553) & (g604) & (g2602) & (g2644)) + ((g553) & (!g604) & (!g2602) & (!g2644)) + ((g553) & (!g604) & (!g2602) & (g2644)) + ((g553) & (!g604) & (g2602) & (!g2644)) + ((g553) & (g604) & (!g2602) & (!g2644)));
	assign g2692 = (((!g2601) & (!g2653) & (!g2668) & (g2691)) + ((!g2601) & (g2653) & (!g2668) & (g2691)) + ((!g2601) & (g2653) & (g2668) & (g2691)) + ((g2601) & (!g2653) & (!g2668) & (!g2691)) + ((g2601) & (!g2653) & (g2668) & (!g2691)) + ((g2601) & (!g2653) & (g2668) & (g2691)) + ((g2601) & (g2653) & (!g2668) & (!g2691)) + ((g2601) & (g2653) & (g2668) & (!g2691)));
	assign g2693 = (((!g604) & (!g2602) & (g2644) & (!g2653) & (!g2668)) + ((!g604) & (!g2602) & (g2644) & (g2653) & (!g2668)) + ((!g604) & (!g2602) & (g2644) & (g2653) & (g2668)) + ((!g604) & (g2602) & (!g2644) & (!g2653) & (!g2668)) + ((!g604) & (g2602) & (!g2644) & (!g2653) & (g2668)) + ((!g604) & (g2602) & (!g2644) & (g2653) & (!g2668)) + ((!g604) & (g2602) & (!g2644) & (g2653) & (g2668)) + ((!g604) & (g2602) & (g2644) & (!g2653) & (g2668)) + ((g604) & (!g2602) & (!g2644) & (!g2653) & (!g2668)) + ((g604) & (!g2602) & (!g2644) & (g2653) & (!g2668)) + ((g604) & (!g2602) & (!g2644) & (g2653) & (g2668)) + ((g604) & (g2602) & (!g2644) & (!g2653) & (g2668)) + ((g604) & (g2602) & (g2644) & (!g2653) & (!g2668)) + ((g604) & (g2602) & (g2644) & (!g2653) & (g2668)) + ((g604) & (g2602) & (g2644) & (g2653) & (!g2668)) + ((g604) & (g2602) & (g2644) & (g2653) & (g2668)));
	assign g2694 = (((!g645) & (!g700) & (g2604) & (g2643)) + ((!g645) & (g700) & (!g2604) & (g2643)) + ((!g645) & (g700) & (g2604) & (!g2643)) + ((!g645) & (g700) & (g2604) & (g2643)) + ((g645) & (!g700) & (!g2604) & (!g2643)) + ((g645) & (!g700) & (!g2604) & (g2643)) + ((g645) & (!g700) & (g2604) & (!g2643)) + ((g645) & (g700) & (!g2604) & (!g2643)));
	assign g2695 = (((!g2603) & (!g2653) & (!g2668) & (g2694)) + ((!g2603) & (g2653) & (!g2668) & (g2694)) + ((!g2603) & (g2653) & (g2668) & (g2694)) + ((g2603) & (!g2653) & (!g2668) & (!g2694)) + ((g2603) & (!g2653) & (g2668) & (!g2694)) + ((g2603) & (!g2653) & (g2668) & (g2694)) + ((g2603) & (g2653) & (!g2668) & (!g2694)) + ((g2603) & (g2653) & (g2668) & (!g2694)));
	assign g2696 = (((!g700) & (!g2604) & (g2643) & (!g2653) & (!g2668)) + ((!g700) & (!g2604) & (g2643) & (g2653) & (!g2668)) + ((!g700) & (!g2604) & (g2643) & (g2653) & (g2668)) + ((!g700) & (g2604) & (!g2643) & (!g2653) & (!g2668)) + ((!g700) & (g2604) & (!g2643) & (!g2653) & (g2668)) + ((!g700) & (g2604) & (!g2643) & (g2653) & (!g2668)) + ((!g700) & (g2604) & (!g2643) & (g2653) & (g2668)) + ((!g700) & (g2604) & (g2643) & (!g2653) & (g2668)) + ((g700) & (!g2604) & (!g2643) & (!g2653) & (!g2668)) + ((g700) & (!g2604) & (!g2643) & (g2653) & (!g2668)) + ((g700) & (!g2604) & (!g2643) & (g2653) & (g2668)) + ((g700) & (g2604) & (!g2643) & (!g2653) & (g2668)) + ((g700) & (g2604) & (g2643) & (!g2653) & (!g2668)) + ((g700) & (g2604) & (g2643) & (!g2653) & (g2668)) + ((g700) & (g2604) & (g2643) & (g2653) & (!g2668)) + ((g700) & (g2604) & (g2643) & (g2653) & (g2668)));
	assign g2697 = (((!g744) & (!g803) & (g2606) & (g2642)) + ((!g744) & (g803) & (!g2606) & (g2642)) + ((!g744) & (g803) & (g2606) & (!g2642)) + ((!g744) & (g803) & (g2606) & (g2642)) + ((g744) & (!g803) & (!g2606) & (!g2642)) + ((g744) & (!g803) & (!g2606) & (g2642)) + ((g744) & (!g803) & (g2606) & (!g2642)) + ((g744) & (g803) & (!g2606) & (!g2642)));
	assign g2698 = (((!g2605) & (!g2653) & (!g2668) & (g2697)) + ((!g2605) & (g2653) & (!g2668) & (g2697)) + ((!g2605) & (g2653) & (g2668) & (g2697)) + ((g2605) & (!g2653) & (!g2668) & (!g2697)) + ((g2605) & (!g2653) & (g2668) & (!g2697)) + ((g2605) & (!g2653) & (g2668) & (g2697)) + ((g2605) & (g2653) & (!g2668) & (!g2697)) + ((g2605) & (g2653) & (g2668) & (!g2697)));
	assign g2699 = (((!g803) & (!g2606) & (g2642) & (!g2653) & (!g2668)) + ((!g803) & (!g2606) & (g2642) & (g2653) & (!g2668)) + ((!g803) & (!g2606) & (g2642) & (g2653) & (g2668)) + ((!g803) & (g2606) & (!g2642) & (!g2653) & (!g2668)) + ((!g803) & (g2606) & (!g2642) & (!g2653) & (g2668)) + ((!g803) & (g2606) & (!g2642) & (g2653) & (!g2668)) + ((!g803) & (g2606) & (!g2642) & (g2653) & (g2668)) + ((!g803) & (g2606) & (g2642) & (!g2653) & (g2668)) + ((g803) & (!g2606) & (!g2642) & (!g2653) & (!g2668)) + ((g803) & (!g2606) & (!g2642) & (g2653) & (!g2668)) + ((g803) & (!g2606) & (!g2642) & (g2653) & (g2668)) + ((g803) & (g2606) & (!g2642) & (!g2653) & (g2668)) + ((g803) & (g2606) & (g2642) & (!g2653) & (!g2668)) + ((g803) & (g2606) & (g2642) & (!g2653) & (g2668)) + ((g803) & (g2606) & (g2642) & (g2653) & (!g2668)) + ((g803) & (g2606) & (g2642) & (g2653) & (g2668)));
	assign g2700 = (((!g851) & (!g914) & (g2608) & (g2641)) + ((!g851) & (g914) & (!g2608) & (g2641)) + ((!g851) & (g914) & (g2608) & (!g2641)) + ((!g851) & (g914) & (g2608) & (g2641)) + ((g851) & (!g914) & (!g2608) & (!g2641)) + ((g851) & (!g914) & (!g2608) & (g2641)) + ((g851) & (!g914) & (g2608) & (!g2641)) + ((g851) & (g914) & (!g2608) & (!g2641)));
	assign g2701 = (((!g2607) & (!g2653) & (!g2668) & (g2700)) + ((!g2607) & (g2653) & (!g2668) & (g2700)) + ((!g2607) & (g2653) & (g2668) & (g2700)) + ((g2607) & (!g2653) & (!g2668) & (!g2700)) + ((g2607) & (!g2653) & (g2668) & (!g2700)) + ((g2607) & (!g2653) & (g2668) & (g2700)) + ((g2607) & (g2653) & (!g2668) & (!g2700)) + ((g2607) & (g2653) & (g2668) & (!g2700)));
	assign g2702 = (((!g914) & (!g2608) & (g2641) & (!g2653) & (!g2668)) + ((!g914) & (!g2608) & (g2641) & (g2653) & (!g2668)) + ((!g914) & (!g2608) & (g2641) & (g2653) & (g2668)) + ((!g914) & (g2608) & (!g2641) & (!g2653) & (!g2668)) + ((!g914) & (g2608) & (!g2641) & (!g2653) & (g2668)) + ((!g914) & (g2608) & (!g2641) & (g2653) & (!g2668)) + ((!g914) & (g2608) & (!g2641) & (g2653) & (g2668)) + ((!g914) & (g2608) & (g2641) & (!g2653) & (g2668)) + ((g914) & (!g2608) & (!g2641) & (!g2653) & (!g2668)) + ((g914) & (!g2608) & (!g2641) & (g2653) & (!g2668)) + ((g914) & (!g2608) & (!g2641) & (g2653) & (g2668)) + ((g914) & (g2608) & (!g2641) & (!g2653) & (g2668)) + ((g914) & (g2608) & (g2641) & (!g2653) & (!g2668)) + ((g914) & (g2608) & (g2641) & (!g2653) & (g2668)) + ((g914) & (g2608) & (g2641) & (g2653) & (!g2668)) + ((g914) & (g2608) & (g2641) & (g2653) & (g2668)));
	assign g2703 = (((!g1032) & (!g1030) & (g2610) & (g2640)) + ((!g1032) & (g1030) & (!g2610) & (g2640)) + ((!g1032) & (g1030) & (g2610) & (!g2640)) + ((!g1032) & (g1030) & (g2610) & (g2640)) + ((g1032) & (!g1030) & (!g2610) & (!g2640)) + ((g1032) & (!g1030) & (!g2610) & (g2640)) + ((g1032) & (!g1030) & (g2610) & (!g2640)) + ((g1032) & (g1030) & (!g2610) & (!g2640)));
	assign g2704 = (((!g2609) & (!g2653) & (!g2668) & (g2703)) + ((!g2609) & (g2653) & (!g2668) & (g2703)) + ((!g2609) & (g2653) & (g2668) & (g2703)) + ((g2609) & (!g2653) & (!g2668) & (!g2703)) + ((g2609) & (!g2653) & (g2668) & (!g2703)) + ((g2609) & (!g2653) & (g2668) & (g2703)) + ((g2609) & (g2653) & (!g2668) & (!g2703)) + ((g2609) & (g2653) & (g2668) & (!g2703)));
	assign g2705 = (((!g1030) & (!g2610) & (g2640) & (!g2653) & (!g2668)) + ((!g1030) & (!g2610) & (g2640) & (g2653) & (!g2668)) + ((!g1030) & (!g2610) & (g2640) & (g2653) & (g2668)) + ((!g1030) & (g2610) & (!g2640) & (!g2653) & (!g2668)) + ((!g1030) & (g2610) & (!g2640) & (!g2653) & (g2668)) + ((!g1030) & (g2610) & (!g2640) & (g2653) & (!g2668)) + ((!g1030) & (g2610) & (!g2640) & (g2653) & (g2668)) + ((!g1030) & (g2610) & (g2640) & (!g2653) & (g2668)) + ((g1030) & (!g2610) & (!g2640) & (!g2653) & (!g2668)) + ((g1030) & (!g2610) & (!g2640) & (g2653) & (!g2668)) + ((g1030) & (!g2610) & (!g2640) & (g2653) & (g2668)) + ((g1030) & (g2610) & (!g2640) & (!g2653) & (g2668)) + ((g1030) & (g2610) & (g2640) & (!g2653) & (!g2668)) + ((g1030) & (g2610) & (g2640) & (!g2653) & (g2668)) + ((g1030) & (g2610) & (g2640) & (g2653) & (!g2668)) + ((g1030) & (g2610) & (g2640) & (g2653) & (g2668)));
	assign g2706 = (((!g1160) & (!g1154) & (g2612) & (g2639)) + ((!g1160) & (g1154) & (!g2612) & (g2639)) + ((!g1160) & (g1154) & (g2612) & (!g2639)) + ((!g1160) & (g1154) & (g2612) & (g2639)) + ((g1160) & (!g1154) & (!g2612) & (!g2639)) + ((g1160) & (!g1154) & (!g2612) & (g2639)) + ((g1160) & (!g1154) & (g2612) & (!g2639)) + ((g1160) & (g1154) & (!g2612) & (!g2639)));
	assign g2707 = (((!g2611) & (!g2653) & (!g2668) & (g2706)) + ((!g2611) & (g2653) & (!g2668) & (g2706)) + ((!g2611) & (g2653) & (g2668) & (g2706)) + ((g2611) & (!g2653) & (!g2668) & (!g2706)) + ((g2611) & (!g2653) & (g2668) & (!g2706)) + ((g2611) & (!g2653) & (g2668) & (g2706)) + ((g2611) & (g2653) & (!g2668) & (!g2706)) + ((g2611) & (g2653) & (g2668) & (!g2706)));
	assign g2708 = (((!g1154) & (!g2612) & (g2639) & (!g2653) & (!g2668)) + ((!g1154) & (!g2612) & (g2639) & (g2653) & (!g2668)) + ((!g1154) & (!g2612) & (g2639) & (g2653) & (g2668)) + ((!g1154) & (g2612) & (!g2639) & (!g2653) & (!g2668)) + ((!g1154) & (g2612) & (!g2639) & (!g2653) & (g2668)) + ((!g1154) & (g2612) & (!g2639) & (g2653) & (!g2668)) + ((!g1154) & (g2612) & (!g2639) & (g2653) & (g2668)) + ((!g1154) & (g2612) & (g2639) & (!g2653) & (g2668)) + ((g1154) & (!g2612) & (!g2639) & (!g2653) & (!g2668)) + ((g1154) & (!g2612) & (!g2639) & (g2653) & (!g2668)) + ((g1154) & (!g2612) & (!g2639) & (g2653) & (g2668)) + ((g1154) & (g2612) & (!g2639) & (!g2653) & (g2668)) + ((g1154) & (g2612) & (g2639) & (!g2653) & (!g2668)) + ((g1154) & (g2612) & (g2639) & (!g2653) & (g2668)) + ((g1154) & (g2612) & (g2639) & (g2653) & (!g2668)) + ((g1154) & (g2612) & (g2639) & (g2653) & (g2668)));
	assign g2709 = (((!g1295) & (!g1285) & (g2614) & (g2638)) + ((!g1295) & (g1285) & (!g2614) & (g2638)) + ((!g1295) & (g1285) & (g2614) & (!g2638)) + ((!g1295) & (g1285) & (g2614) & (g2638)) + ((g1295) & (!g1285) & (!g2614) & (!g2638)) + ((g1295) & (!g1285) & (!g2614) & (g2638)) + ((g1295) & (!g1285) & (g2614) & (!g2638)) + ((g1295) & (g1285) & (!g2614) & (!g2638)));
	assign g2710 = (((!g2613) & (!g2653) & (!g2668) & (g2709)) + ((!g2613) & (g2653) & (!g2668) & (g2709)) + ((!g2613) & (g2653) & (g2668) & (g2709)) + ((g2613) & (!g2653) & (!g2668) & (!g2709)) + ((g2613) & (!g2653) & (g2668) & (!g2709)) + ((g2613) & (!g2653) & (g2668) & (g2709)) + ((g2613) & (g2653) & (!g2668) & (!g2709)) + ((g2613) & (g2653) & (g2668) & (!g2709)));
	assign g2711 = (((!g1285) & (!g2614) & (g2638) & (!g2653) & (!g2668)) + ((!g1285) & (!g2614) & (g2638) & (g2653) & (!g2668)) + ((!g1285) & (!g2614) & (g2638) & (g2653) & (g2668)) + ((!g1285) & (g2614) & (!g2638) & (!g2653) & (!g2668)) + ((!g1285) & (g2614) & (!g2638) & (!g2653) & (g2668)) + ((!g1285) & (g2614) & (!g2638) & (g2653) & (!g2668)) + ((!g1285) & (g2614) & (!g2638) & (g2653) & (g2668)) + ((!g1285) & (g2614) & (g2638) & (!g2653) & (g2668)) + ((g1285) & (!g2614) & (!g2638) & (!g2653) & (!g2668)) + ((g1285) & (!g2614) & (!g2638) & (g2653) & (!g2668)) + ((g1285) & (!g2614) & (!g2638) & (g2653) & (g2668)) + ((g1285) & (g2614) & (!g2638) & (!g2653) & (g2668)) + ((g1285) & (g2614) & (g2638) & (!g2653) & (!g2668)) + ((g1285) & (g2614) & (g2638) & (!g2653) & (g2668)) + ((g1285) & (g2614) & (g2638) & (g2653) & (!g2668)) + ((g1285) & (g2614) & (g2638) & (g2653) & (g2668)));
	assign g2712 = (((!g1437) & (!g1423) & (g2616) & (g2637)) + ((!g1437) & (g1423) & (!g2616) & (g2637)) + ((!g1437) & (g1423) & (g2616) & (!g2637)) + ((!g1437) & (g1423) & (g2616) & (g2637)) + ((g1437) & (!g1423) & (!g2616) & (!g2637)) + ((g1437) & (!g1423) & (!g2616) & (g2637)) + ((g1437) & (!g1423) & (g2616) & (!g2637)) + ((g1437) & (g1423) & (!g2616) & (!g2637)));
	assign g2713 = (((!g2615) & (!g2653) & (!g2668) & (g2712)) + ((!g2615) & (g2653) & (!g2668) & (g2712)) + ((!g2615) & (g2653) & (g2668) & (g2712)) + ((g2615) & (!g2653) & (!g2668) & (!g2712)) + ((g2615) & (!g2653) & (g2668) & (!g2712)) + ((g2615) & (!g2653) & (g2668) & (g2712)) + ((g2615) & (g2653) & (!g2668) & (!g2712)) + ((g2615) & (g2653) & (g2668) & (!g2712)));
	assign g2714 = (((!g1423) & (!g2616) & (g2637) & (!g2653) & (!g2668)) + ((!g1423) & (!g2616) & (g2637) & (g2653) & (!g2668)) + ((!g1423) & (!g2616) & (g2637) & (g2653) & (g2668)) + ((!g1423) & (g2616) & (!g2637) & (!g2653) & (!g2668)) + ((!g1423) & (g2616) & (!g2637) & (!g2653) & (g2668)) + ((!g1423) & (g2616) & (!g2637) & (g2653) & (!g2668)) + ((!g1423) & (g2616) & (!g2637) & (g2653) & (g2668)) + ((!g1423) & (g2616) & (g2637) & (!g2653) & (g2668)) + ((g1423) & (!g2616) & (!g2637) & (!g2653) & (!g2668)) + ((g1423) & (!g2616) & (!g2637) & (g2653) & (!g2668)) + ((g1423) & (!g2616) & (!g2637) & (g2653) & (g2668)) + ((g1423) & (g2616) & (!g2637) & (!g2653) & (g2668)) + ((g1423) & (g2616) & (g2637) & (!g2653) & (!g2668)) + ((g1423) & (g2616) & (g2637) & (!g2653) & (g2668)) + ((g1423) & (g2616) & (g2637) & (g2653) & (!g2668)) + ((g1423) & (g2616) & (g2637) & (g2653) & (g2668)));
	assign g2715 = (((!g1586) & (!g1568) & (g2618) & (g2636)) + ((!g1586) & (g1568) & (!g2618) & (g2636)) + ((!g1586) & (g1568) & (g2618) & (!g2636)) + ((!g1586) & (g1568) & (g2618) & (g2636)) + ((g1586) & (!g1568) & (!g2618) & (!g2636)) + ((g1586) & (!g1568) & (!g2618) & (g2636)) + ((g1586) & (!g1568) & (g2618) & (!g2636)) + ((g1586) & (g1568) & (!g2618) & (!g2636)));
	assign g2716 = (((!g2617) & (!g2653) & (!g2668) & (g2715)) + ((!g2617) & (g2653) & (!g2668) & (g2715)) + ((!g2617) & (g2653) & (g2668) & (g2715)) + ((g2617) & (!g2653) & (!g2668) & (!g2715)) + ((g2617) & (!g2653) & (g2668) & (!g2715)) + ((g2617) & (!g2653) & (g2668) & (g2715)) + ((g2617) & (g2653) & (!g2668) & (!g2715)) + ((g2617) & (g2653) & (g2668) & (!g2715)));
	assign g2717 = (((!g1568) & (!g2618) & (g2636) & (!g2653) & (!g2668)) + ((!g1568) & (!g2618) & (g2636) & (g2653) & (!g2668)) + ((!g1568) & (!g2618) & (g2636) & (g2653) & (g2668)) + ((!g1568) & (g2618) & (!g2636) & (!g2653) & (!g2668)) + ((!g1568) & (g2618) & (!g2636) & (!g2653) & (g2668)) + ((!g1568) & (g2618) & (!g2636) & (g2653) & (!g2668)) + ((!g1568) & (g2618) & (!g2636) & (g2653) & (g2668)) + ((!g1568) & (g2618) & (g2636) & (!g2653) & (g2668)) + ((g1568) & (!g2618) & (!g2636) & (!g2653) & (!g2668)) + ((g1568) & (!g2618) & (!g2636) & (g2653) & (!g2668)) + ((g1568) & (!g2618) & (!g2636) & (g2653) & (g2668)) + ((g1568) & (g2618) & (!g2636) & (!g2653) & (g2668)) + ((g1568) & (g2618) & (g2636) & (!g2653) & (!g2668)) + ((g1568) & (g2618) & (g2636) & (!g2653) & (g2668)) + ((g1568) & (g2618) & (g2636) & (g2653) & (!g2668)) + ((g1568) & (g2618) & (g2636) & (g2653) & (g2668)));
	assign g2718 = (((!g1742) & (!g1720) & (g2620) & (g2635)) + ((!g1742) & (g1720) & (!g2620) & (g2635)) + ((!g1742) & (g1720) & (g2620) & (!g2635)) + ((!g1742) & (g1720) & (g2620) & (g2635)) + ((g1742) & (!g1720) & (!g2620) & (!g2635)) + ((g1742) & (!g1720) & (!g2620) & (g2635)) + ((g1742) & (!g1720) & (g2620) & (!g2635)) + ((g1742) & (g1720) & (!g2620) & (!g2635)));
	assign g2719 = (((!g2619) & (!g2653) & (!g2668) & (g2718)) + ((!g2619) & (g2653) & (!g2668) & (g2718)) + ((!g2619) & (g2653) & (g2668) & (g2718)) + ((g2619) & (!g2653) & (!g2668) & (!g2718)) + ((g2619) & (!g2653) & (g2668) & (!g2718)) + ((g2619) & (!g2653) & (g2668) & (g2718)) + ((g2619) & (g2653) & (!g2668) & (!g2718)) + ((g2619) & (g2653) & (g2668) & (!g2718)));
	assign g2720 = (((!g1720) & (!g2620) & (g2635) & (!g2653) & (!g2668)) + ((!g1720) & (!g2620) & (g2635) & (g2653) & (!g2668)) + ((!g1720) & (!g2620) & (g2635) & (g2653) & (g2668)) + ((!g1720) & (g2620) & (!g2635) & (!g2653) & (!g2668)) + ((!g1720) & (g2620) & (!g2635) & (!g2653) & (g2668)) + ((!g1720) & (g2620) & (!g2635) & (g2653) & (!g2668)) + ((!g1720) & (g2620) & (!g2635) & (g2653) & (g2668)) + ((!g1720) & (g2620) & (g2635) & (!g2653) & (g2668)) + ((g1720) & (!g2620) & (!g2635) & (!g2653) & (!g2668)) + ((g1720) & (!g2620) & (!g2635) & (g2653) & (!g2668)) + ((g1720) & (!g2620) & (!g2635) & (g2653) & (g2668)) + ((g1720) & (g2620) & (!g2635) & (!g2653) & (g2668)) + ((g1720) & (g2620) & (g2635) & (!g2653) & (!g2668)) + ((g1720) & (g2620) & (g2635) & (!g2653) & (g2668)) + ((g1720) & (g2620) & (g2635) & (g2653) & (!g2668)) + ((g1720) & (g2620) & (g2635) & (g2653) & (g2668)));
	assign g2721 = (((!g1905) & (!g1879) & (g2622) & (g2634)) + ((!g1905) & (g1879) & (!g2622) & (g2634)) + ((!g1905) & (g1879) & (g2622) & (!g2634)) + ((!g1905) & (g1879) & (g2622) & (g2634)) + ((g1905) & (!g1879) & (!g2622) & (!g2634)) + ((g1905) & (!g1879) & (!g2622) & (g2634)) + ((g1905) & (!g1879) & (g2622) & (!g2634)) + ((g1905) & (g1879) & (!g2622) & (!g2634)));
	assign g2722 = (((!g2621) & (!g2653) & (!g2668) & (g2721)) + ((!g2621) & (g2653) & (!g2668) & (g2721)) + ((!g2621) & (g2653) & (g2668) & (g2721)) + ((g2621) & (!g2653) & (!g2668) & (!g2721)) + ((g2621) & (!g2653) & (g2668) & (!g2721)) + ((g2621) & (!g2653) & (g2668) & (g2721)) + ((g2621) & (g2653) & (!g2668) & (!g2721)) + ((g2621) & (g2653) & (g2668) & (!g2721)));
	assign g2723 = (((!g1879) & (!g2622) & (g2634) & (!g2653) & (!g2668)) + ((!g1879) & (!g2622) & (g2634) & (g2653) & (!g2668)) + ((!g1879) & (!g2622) & (g2634) & (g2653) & (g2668)) + ((!g1879) & (g2622) & (!g2634) & (!g2653) & (!g2668)) + ((!g1879) & (g2622) & (!g2634) & (!g2653) & (g2668)) + ((!g1879) & (g2622) & (!g2634) & (g2653) & (!g2668)) + ((!g1879) & (g2622) & (!g2634) & (g2653) & (g2668)) + ((!g1879) & (g2622) & (g2634) & (!g2653) & (g2668)) + ((g1879) & (!g2622) & (!g2634) & (!g2653) & (!g2668)) + ((g1879) & (!g2622) & (!g2634) & (g2653) & (!g2668)) + ((g1879) & (!g2622) & (!g2634) & (g2653) & (g2668)) + ((g1879) & (g2622) & (!g2634) & (!g2653) & (g2668)) + ((g1879) & (g2622) & (g2634) & (!g2653) & (!g2668)) + ((g1879) & (g2622) & (g2634) & (!g2653) & (g2668)) + ((g1879) & (g2622) & (g2634) & (g2653) & (!g2668)) + ((g1879) & (g2622) & (g2634) & (g2653) & (g2668)));
	assign g2724 = (((!g2075) & (!g2045) & (g2624) & (g2633)) + ((!g2075) & (g2045) & (!g2624) & (g2633)) + ((!g2075) & (g2045) & (g2624) & (!g2633)) + ((!g2075) & (g2045) & (g2624) & (g2633)) + ((g2075) & (!g2045) & (!g2624) & (!g2633)) + ((g2075) & (!g2045) & (!g2624) & (g2633)) + ((g2075) & (!g2045) & (g2624) & (!g2633)) + ((g2075) & (g2045) & (!g2624) & (!g2633)));
	assign g2725 = (((!g2623) & (!g2653) & (!g2668) & (g2724)) + ((!g2623) & (g2653) & (!g2668) & (g2724)) + ((!g2623) & (g2653) & (g2668) & (g2724)) + ((g2623) & (!g2653) & (!g2668) & (!g2724)) + ((g2623) & (!g2653) & (g2668) & (!g2724)) + ((g2623) & (!g2653) & (g2668) & (g2724)) + ((g2623) & (g2653) & (!g2668) & (!g2724)) + ((g2623) & (g2653) & (g2668) & (!g2724)));
	assign g2726 = (((!g2045) & (!g2624) & (g2633) & (!g2653) & (!g2668)) + ((!g2045) & (!g2624) & (g2633) & (g2653) & (!g2668)) + ((!g2045) & (!g2624) & (g2633) & (g2653) & (g2668)) + ((!g2045) & (g2624) & (!g2633) & (!g2653) & (!g2668)) + ((!g2045) & (g2624) & (!g2633) & (!g2653) & (g2668)) + ((!g2045) & (g2624) & (!g2633) & (g2653) & (!g2668)) + ((!g2045) & (g2624) & (!g2633) & (g2653) & (g2668)) + ((!g2045) & (g2624) & (g2633) & (!g2653) & (g2668)) + ((g2045) & (!g2624) & (!g2633) & (!g2653) & (!g2668)) + ((g2045) & (!g2624) & (!g2633) & (g2653) & (!g2668)) + ((g2045) & (!g2624) & (!g2633) & (g2653) & (g2668)) + ((g2045) & (g2624) & (!g2633) & (!g2653) & (g2668)) + ((g2045) & (g2624) & (g2633) & (!g2653) & (!g2668)) + ((g2045) & (g2624) & (g2633) & (!g2653) & (g2668)) + ((g2045) & (g2624) & (g2633) & (g2653) & (!g2668)) + ((g2045) & (g2624) & (g2633) & (g2653) & (g2668)));
	assign g2727 = (((!g2252) & (!g2218) & (g2626) & (g2632)) + ((!g2252) & (g2218) & (!g2626) & (g2632)) + ((!g2252) & (g2218) & (g2626) & (!g2632)) + ((!g2252) & (g2218) & (g2626) & (g2632)) + ((g2252) & (!g2218) & (!g2626) & (!g2632)) + ((g2252) & (!g2218) & (!g2626) & (g2632)) + ((g2252) & (!g2218) & (g2626) & (!g2632)) + ((g2252) & (g2218) & (!g2626) & (!g2632)));
	assign g2728 = (((!g2625) & (!g2653) & (!g2668) & (g2727)) + ((!g2625) & (g2653) & (!g2668) & (g2727)) + ((!g2625) & (g2653) & (g2668) & (g2727)) + ((g2625) & (!g2653) & (!g2668) & (!g2727)) + ((g2625) & (!g2653) & (g2668) & (!g2727)) + ((g2625) & (!g2653) & (g2668) & (g2727)) + ((g2625) & (g2653) & (!g2668) & (!g2727)) + ((g2625) & (g2653) & (g2668) & (!g2727)));
	assign g2729 = (((!g2218) & (!g2626) & (g2632) & (!g2653) & (!g2668)) + ((!g2218) & (!g2626) & (g2632) & (g2653) & (!g2668)) + ((!g2218) & (!g2626) & (g2632) & (g2653) & (g2668)) + ((!g2218) & (g2626) & (!g2632) & (!g2653) & (!g2668)) + ((!g2218) & (g2626) & (!g2632) & (!g2653) & (g2668)) + ((!g2218) & (g2626) & (!g2632) & (g2653) & (!g2668)) + ((!g2218) & (g2626) & (!g2632) & (g2653) & (g2668)) + ((!g2218) & (g2626) & (g2632) & (!g2653) & (g2668)) + ((g2218) & (!g2626) & (!g2632) & (!g2653) & (!g2668)) + ((g2218) & (!g2626) & (!g2632) & (g2653) & (!g2668)) + ((g2218) & (!g2626) & (!g2632) & (g2653) & (g2668)) + ((g2218) & (g2626) & (!g2632) & (!g2653) & (g2668)) + ((g2218) & (g2626) & (g2632) & (!g2653) & (!g2668)) + ((g2218) & (g2626) & (g2632) & (!g2653) & (g2668)) + ((g2218) & (g2626) & (g2632) & (g2653) & (!g2668)) + ((g2218) & (g2626) & (g2632) & (g2653) & (g2668)));
	assign g2730 = (((!g2436) & (!g2398) & (g2629) & (g2631)) + ((!g2436) & (g2398) & (!g2629) & (g2631)) + ((!g2436) & (g2398) & (g2629) & (!g2631)) + ((!g2436) & (g2398) & (g2629) & (g2631)) + ((g2436) & (!g2398) & (!g2629) & (!g2631)) + ((g2436) & (!g2398) & (!g2629) & (g2631)) + ((g2436) & (!g2398) & (g2629) & (!g2631)) + ((g2436) & (g2398) & (!g2629) & (!g2631)));
	assign g2731 = (((!g2628) & (!g2653) & (!g2668) & (g2730)) + ((!g2628) & (g2653) & (!g2668) & (g2730)) + ((!g2628) & (g2653) & (g2668) & (g2730)) + ((g2628) & (!g2653) & (!g2668) & (!g2730)) + ((g2628) & (!g2653) & (g2668) & (!g2730)) + ((g2628) & (!g2653) & (g2668) & (g2730)) + ((g2628) & (g2653) & (!g2668) & (!g2730)) + ((g2628) & (g2653) & (g2668) & (!g2730)));
	assign g2732 = (((!g2398) & (!g2629) & (g2631) & (!g2653) & (!g2668)) + ((!g2398) & (!g2629) & (g2631) & (g2653) & (!g2668)) + ((!g2398) & (!g2629) & (g2631) & (g2653) & (g2668)) + ((!g2398) & (g2629) & (!g2631) & (!g2653) & (!g2668)) + ((!g2398) & (g2629) & (!g2631) & (!g2653) & (g2668)) + ((!g2398) & (g2629) & (!g2631) & (g2653) & (!g2668)) + ((!g2398) & (g2629) & (!g2631) & (g2653) & (g2668)) + ((!g2398) & (g2629) & (g2631) & (!g2653) & (g2668)) + ((g2398) & (!g2629) & (!g2631) & (!g2653) & (!g2668)) + ((g2398) & (!g2629) & (!g2631) & (g2653) & (!g2668)) + ((g2398) & (!g2629) & (!g2631) & (g2653) & (g2668)) + ((g2398) & (g2629) & (!g2631) & (!g2653) & (g2668)) + ((g2398) & (g2629) & (g2631) & (!g2653) & (!g2668)) + ((g2398) & (g2629) & (g2631) & (!g2653) & (g2668)) + ((g2398) & (g2629) & (g2631) & (g2653) & (!g2668)) + ((g2398) & (g2629) & (g2631) & (g2653) & (g2668)));
	assign g2733 = (((!g2627) & (!ax20x) & (!g2585) & (g2630)) + ((!g2627) & (!ax20x) & (g2585) & (g2630)) + ((!g2627) & (ax20x) & (!g2585) & (!g2630)) + ((!g2627) & (ax20x) & (!g2585) & (g2630)) + ((g2627) & (!ax20x) & (!g2585) & (!g2630)) + ((g2627) & (!ax20x) & (g2585) & (!g2630)) + ((g2627) & (ax20x) & (g2585) & (!g2630)) + ((g2627) & (ax20x) & (g2585) & (g2630)));
	assign g2734 = (((!ax20x) & (!ax21x) & (!g2585) & (!g2653) & (!g2668) & (g2733)) + ((!ax20x) & (!ax21x) & (!g2585) & (!g2653) & (g2668) & (!g2733)) + ((!ax20x) & (!ax21x) & (!g2585) & (!g2653) & (g2668) & (g2733)) + ((!ax20x) & (!ax21x) & (!g2585) & (g2653) & (!g2668) & (g2733)) + ((!ax20x) & (!ax21x) & (!g2585) & (g2653) & (g2668) & (g2733)) + ((!ax20x) & (!ax21x) & (g2585) & (!g2653) & (!g2668) & (!g2733)) + ((!ax20x) & (!ax21x) & (g2585) & (g2653) & (!g2668) & (!g2733)) + ((!ax20x) & (!ax21x) & (g2585) & (g2653) & (g2668) & (!g2733)) + ((!ax20x) & (ax21x) & (!g2585) & (!g2653) & (!g2668) & (!g2733)) + ((!ax20x) & (ax21x) & (!g2585) & (g2653) & (!g2668) & (!g2733)) + ((!ax20x) & (ax21x) & (!g2585) & (g2653) & (g2668) & (!g2733)) + ((!ax20x) & (ax21x) & (g2585) & (!g2653) & (!g2668) & (g2733)) + ((!ax20x) & (ax21x) & (g2585) & (!g2653) & (g2668) & (!g2733)) + ((!ax20x) & (ax21x) & (g2585) & (!g2653) & (g2668) & (g2733)) + ((!ax20x) & (ax21x) & (g2585) & (g2653) & (!g2668) & (g2733)) + ((!ax20x) & (ax21x) & (g2585) & (g2653) & (g2668) & (g2733)) + ((ax20x) & (!ax21x) & (!g2585) & (!g2653) & (!g2668) & (!g2733)) + ((ax20x) & (!ax21x) & (!g2585) & (g2653) & (!g2668) & (!g2733)) + ((ax20x) & (!ax21x) & (!g2585) & (g2653) & (g2668) & (!g2733)) + ((ax20x) & (!ax21x) & (g2585) & (!g2653) & (!g2668) & (!g2733)) + ((ax20x) & (!ax21x) & (g2585) & (g2653) & (!g2668) & (!g2733)) + ((ax20x) & (!ax21x) & (g2585) & (g2653) & (g2668) & (!g2733)) + ((ax20x) & (ax21x) & (!g2585) & (!g2653) & (!g2668) & (g2733)) + ((ax20x) & (ax21x) & (!g2585) & (!g2653) & (g2668) & (!g2733)) + ((ax20x) & (ax21x) & (!g2585) & (!g2653) & (g2668) & (g2733)) + ((ax20x) & (ax21x) & (!g2585) & (g2653) & (!g2668) & (g2733)) + ((ax20x) & (ax21x) & (!g2585) & (g2653) & (g2668) & (g2733)) + ((ax20x) & (ax21x) & (g2585) & (!g2653) & (!g2668) & (g2733)) + ((ax20x) & (ax21x) & (g2585) & (!g2653) & (g2668) & (!g2733)) + ((ax20x) & (ax21x) & (g2585) & (!g2653) & (g2668) & (g2733)) + ((ax20x) & (ax21x) & (g2585) & (g2653) & (!g2668) & (g2733)) + ((ax20x) & (ax21x) & (g2585) & (g2653) & (g2668) & (g2733)));
	assign g2735 = (((!ax20x) & (!g2585) & (!g2630) & (!g2653) & (g2668)) + ((!ax20x) & (!g2585) & (g2630) & (!g2653) & (!g2668)) + ((!ax20x) & (!g2585) & (g2630) & (!g2653) & (g2668)) + ((!ax20x) & (!g2585) & (g2630) & (g2653) & (!g2668)) + ((!ax20x) & (!g2585) & (g2630) & (g2653) & (g2668)) + ((!ax20x) & (g2585) & (g2630) & (!g2653) & (!g2668)) + ((!ax20x) & (g2585) & (g2630) & (g2653) & (!g2668)) + ((!ax20x) & (g2585) & (g2630) & (g2653) & (g2668)) + ((ax20x) & (!g2585) & (!g2630) & (!g2653) & (!g2668)) + ((ax20x) & (!g2585) & (!g2630) & (g2653) & (!g2668)) + ((ax20x) & (!g2585) & (!g2630) & (g2653) & (g2668)) + ((ax20x) & (g2585) & (!g2630) & (!g2653) & (!g2668)) + ((ax20x) & (g2585) & (!g2630) & (!g2653) & (g2668)) + ((ax20x) & (g2585) & (!g2630) & (g2653) & (!g2668)) + ((ax20x) & (g2585) & (!g2630) & (g2653) & (g2668)) + ((ax20x) & (g2585) & (g2630) & (!g2653) & (g2668)));
	assign g2736 = (((!ax16x) & (!ax17x)));
	assign g2737 = (((!g2585) & (!ax18x) & (!ax19x) & (!g2653) & (!g2668) & (!g2736)) + ((!g2585) & (!ax18x) & (!ax19x) & (g2653) & (!g2668) & (!g2736)) + ((!g2585) & (!ax18x) & (!ax19x) & (g2653) & (g2668) & (!g2736)) + ((!g2585) & (!ax18x) & (ax19x) & (!g2653) & (g2668) & (!g2736)) + ((!g2585) & (ax18x) & (ax19x) & (!g2653) & (g2668) & (!g2736)) + ((!g2585) & (ax18x) & (ax19x) & (!g2653) & (g2668) & (g2736)) + ((g2585) & (!ax18x) & (!ax19x) & (!g2653) & (!g2668) & (!g2736)) + ((g2585) & (!ax18x) & (!ax19x) & (!g2653) & (!g2668) & (g2736)) + ((g2585) & (!ax18x) & (!ax19x) & (!g2653) & (g2668) & (!g2736)) + ((g2585) & (!ax18x) & (!ax19x) & (g2653) & (!g2668) & (!g2736)) + ((g2585) & (!ax18x) & (!ax19x) & (g2653) & (!g2668) & (g2736)) + ((g2585) & (!ax18x) & (!ax19x) & (g2653) & (g2668) & (!g2736)) + ((g2585) & (!ax18x) & (!ax19x) & (g2653) & (g2668) & (g2736)) + ((g2585) & (!ax18x) & (ax19x) & (!g2653) & (!g2668) & (!g2736)) + ((g2585) & (!ax18x) & (ax19x) & (!g2653) & (g2668) & (!g2736)) + ((g2585) & (!ax18x) & (ax19x) & (!g2653) & (g2668) & (g2736)) + ((g2585) & (!ax18x) & (ax19x) & (g2653) & (!g2668) & (!g2736)) + ((g2585) & (!ax18x) & (ax19x) & (g2653) & (g2668) & (!g2736)) + ((g2585) & (ax18x) & (!ax19x) & (!g2653) & (g2668) & (!g2736)) + ((g2585) & (ax18x) & (!ax19x) & (!g2653) & (g2668) & (g2736)) + ((g2585) & (ax18x) & (ax19x) & (!g2653) & (!g2668) & (!g2736)) + ((g2585) & (ax18x) & (ax19x) & (!g2653) & (!g2668) & (g2736)) + ((g2585) & (ax18x) & (ax19x) & (!g2653) & (g2668) & (!g2736)) + ((g2585) & (ax18x) & (ax19x) & (!g2653) & (g2668) & (g2736)) + ((g2585) & (ax18x) & (ax19x) & (g2653) & (!g2668) & (!g2736)) + ((g2585) & (ax18x) & (ax19x) & (g2653) & (!g2668) & (g2736)) + ((g2585) & (ax18x) & (ax19x) & (g2653) & (g2668) & (!g2736)) + ((g2585) & (ax18x) & (ax19x) & (g2653) & (g2668) & (g2736)));
	assign g2738 = (((!g2398) & (!g2627) & (g2734) & (g2735) & (g2737)) + ((!g2398) & (g2627) & (g2734) & (!g2735) & (g2737)) + ((!g2398) & (g2627) & (g2734) & (g2735) & (!g2737)) + ((!g2398) & (g2627) & (g2734) & (g2735) & (g2737)) + ((g2398) & (!g2627) & (!g2734) & (g2735) & (g2737)) + ((g2398) & (!g2627) & (g2734) & (!g2735) & (!g2737)) + ((g2398) & (!g2627) & (g2734) & (!g2735) & (g2737)) + ((g2398) & (!g2627) & (g2734) & (g2735) & (!g2737)) + ((g2398) & (!g2627) & (g2734) & (g2735) & (g2737)) + ((g2398) & (g2627) & (!g2734) & (!g2735) & (g2737)) + ((g2398) & (g2627) & (!g2734) & (g2735) & (!g2737)) + ((g2398) & (g2627) & (!g2734) & (g2735) & (g2737)) + ((g2398) & (g2627) & (g2734) & (!g2735) & (!g2737)) + ((g2398) & (g2627) & (g2734) & (!g2735) & (g2737)) + ((g2398) & (g2627) & (g2734) & (g2735) & (!g2737)) + ((g2398) & (g2627) & (g2734) & (g2735) & (g2737)));
	assign g2739 = (((!g2218) & (!g2436) & (g2731) & (g2732) & (g2738)) + ((!g2218) & (g2436) & (g2731) & (!g2732) & (g2738)) + ((!g2218) & (g2436) & (g2731) & (g2732) & (!g2738)) + ((!g2218) & (g2436) & (g2731) & (g2732) & (g2738)) + ((g2218) & (!g2436) & (!g2731) & (g2732) & (g2738)) + ((g2218) & (!g2436) & (g2731) & (!g2732) & (!g2738)) + ((g2218) & (!g2436) & (g2731) & (!g2732) & (g2738)) + ((g2218) & (!g2436) & (g2731) & (g2732) & (!g2738)) + ((g2218) & (!g2436) & (g2731) & (g2732) & (g2738)) + ((g2218) & (g2436) & (!g2731) & (!g2732) & (g2738)) + ((g2218) & (g2436) & (!g2731) & (g2732) & (!g2738)) + ((g2218) & (g2436) & (!g2731) & (g2732) & (g2738)) + ((g2218) & (g2436) & (g2731) & (!g2732) & (!g2738)) + ((g2218) & (g2436) & (g2731) & (!g2732) & (g2738)) + ((g2218) & (g2436) & (g2731) & (g2732) & (!g2738)) + ((g2218) & (g2436) & (g2731) & (g2732) & (g2738)));
	assign g2740 = (((!g2045) & (!g2252) & (g2728) & (g2729) & (g2739)) + ((!g2045) & (g2252) & (g2728) & (!g2729) & (g2739)) + ((!g2045) & (g2252) & (g2728) & (g2729) & (!g2739)) + ((!g2045) & (g2252) & (g2728) & (g2729) & (g2739)) + ((g2045) & (!g2252) & (!g2728) & (g2729) & (g2739)) + ((g2045) & (!g2252) & (g2728) & (!g2729) & (!g2739)) + ((g2045) & (!g2252) & (g2728) & (!g2729) & (g2739)) + ((g2045) & (!g2252) & (g2728) & (g2729) & (!g2739)) + ((g2045) & (!g2252) & (g2728) & (g2729) & (g2739)) + ((g2045) & (g2252) & (!g2728) & (!g2729) & (g2739)) + ((g2045) & (g2252) & (!g2728) & (g2729) & (!g2739)) + ((g2045) & (g2252) & (!g2728) & (g2729) & (g2739)) + ((g2045) & (g2252) & (g2728) & (!g2729) & (!g2739)) + ((g2045) & (g2252) & (g2728) & (!g2729) & (g2739)) + ((g2045) & (g2252) & (g2728) & (g2729) & (!g2739)) + ((g2045) & (g2252) & (g2728) & (g2729) & (g2739)));
	assign g2741 = (((!g1879) & (!g2075) & (g2725) & (g2726) & (g2740)) + ((!g1879) & (g2075) & (g2725) & (!g2726) & (g2740)) + ((!g1879) & (g2075) & (g2725) & (g2726) & (!g2740)) + ((!g1879) & (g2075) & (g2725) & (g2726) & (g2740)) + ((g1879) & (!g2075) & (!g2725) & (g2726) & (g2740)) + ((g1879) & (!g2075) & (g2725) & (!g2726) & (!g2740)) + ((g1879) & (!g2075) & (g2725) & (!g2726) & (g2740)) + ((g1879) & (!g2075) & (g2725) & (g2726) & (!g2740)) + ((g1879) & (!g2075) & (g2725) & (g2726) & (g2740)) + ((g1879) & (g2075) & (!g2725) & (!g2726) & (g2740)) + ((g1879) & (g2075) & (!g2725) & (g2726) & (!g2740)) + ((g1879) & (g2075) & (!g2725) & (g2726) & (g2740)) + ((g1879) & (g2075) & (g2725) & (!g2726) & (!g2740)) + ((g1879) & (g2075) & (g2725) & (!g2726) & (g2740)) + ((g1879) & (g2075) & (g2725) & (g2726) & (!g2740)) + ((g1879) & (g2075) & (g2725) & (g2726) & (g2740)));
	assign g2742 = (((!g1720) & (!g1905) & (g2722) & (g2723) & (g2741)) + ((!g1720) & (g1905) & (g2722) & (!g2723) & (g2741)) + ((!g1720) & (g1905) & (g2722) & (g2723) & (!g2741)) + ((!g1720) & (g1905) & (g2722) & (g2723) & (g2741)) + ((g1720) & (!g1905) & (!g2722) & (g2723) & (g2741)) + ((g1720) & (!g1905) & (g2722) & (!g2723) & (!g2741)) + ((g1720) & (!g1905) & (g2722) & (!g2723) & (g2741)) + ((g1720) & (!g1905) & (g2722) & (g2723) & (!g2741)) + ((g1720) & (!g1905) & (g2722) & (g2723) & (g2741)) + ((g1720) & (g1905) & (!g2722) & (!g2723) & (g2741)) + ((g1720) & (g1905) & (!g2722) & (g2723) & (!g2741)) + ((g1720) & (g1905) & (!g2722) & (g2723) & (g2741)) + ((g1720) & (g1905) & (g2722) & (!g2723) & (!g2741)) + ((g1720) & (g1905) & (g2722) & (!g2723) & (g2741)) + ((g1720) & (g1905) & (g2722) & (g2723) & (!g2741)) + ((g1720) & (g1905) & (g2722) & (g2723) & (g2741)));
	assign g2743 = (((!g1568) & (!g1742) & (g2719) & (g2720) & (g2742)) + ((!g1568) & (g1742) & (g2719) & (!g2720) & (g2742)) + ((!g1568) & (g1742) & (g2719) & (g2720) & (!g2742)) + ((!g1568) & (g1742) & (g2719) & (g2720) & (g2742)) + ((g1568) & (!g1742) & (!g2719) & (g2720) & (g2742)) + ((g1568) & (!g1742) & (g2719) & (!g2720) & (!g2742)) + ((g1568) & (!g1742) & (g2719) & (!g2720) & (g2742)) + ((g1568) & (!g1742) & (g2719) & (g2720) & (!g2742)) + ((g1568) & (!g1742) & (g2719) & (g2720) & (g2742)) + ((g1568) & (g1742) & (!g2719) & (!g2720) & (g2742)) + ((g1568) & (g1742) & (!g2719) & (g2720) & (!g2742)) + ((g1568) & (g1742) & (!g2719) & (g2720) & (g2742)) + ((g1568) & (g1742) & (g2719) & (!g2720) & (!g2742)) + ((g1568) & (g1742) & (g2719) & (!g2720) & (g2742)) + ((g1568) & (g1742) & (g2719) & (g2720) & (!g2742)) + ((g1568) & (g1742) & (g2719) & (g2720) & (g2742)));
	assign g2744 = (((!g1423) & (!g1586) & (g2716) & (g2717) & (g2743)) + ((!g1423) & (g1586) & (g2716) & (!g2717) & (g2743)) + ((!g1423) & (g1586) & (g2716) & (g2717) & (!g2743)) + ((!g1423) & (g1586) & (g2716) & (g2717) & (g2743)) + ((g1423) & (!g1586) & (!g2716) & (g2717) & (g2743)) + ((g1423) & (!g1586) & (g2716) & (!g2717) & (!g2743)) + ((g1423) & (!g1586) & (g2716) & (!g2717) & (g2743)) + ((g1423) & (!g1586) & (g2716) & (g2717) & (!g2743)) + ((g1423) & (!g1586) & (g2716) & (g2717) & (g2743)) + ((g1423) & (g1586) & (!g2716) & (!g2717) & (g2743)) + ((g1423) & (g1586) & (!g2716) & (g2717) & (!g2743)) + ((g1423) & (g1586) & (!g2716) & (g2717) & (g2743)) + ((g1423) & (g1586) & (g2716) & (!g2717) & (!g2743)) + ((g1423) & (g1586) & (g2716) & (!g2717) & (g2743)) + ((g1423) & (g1586) & (g2716) & (g2717) & (!g2743)) + ((g1423) & (g1586) & (g2716) & (g2717) & (g2743)));
	assign g2745 = (((!g1285) & (!g1437) & (g2713) & (g2714) & (g2744)) + ((!g1285) & (g1437) & (g2713) & (!g2714) & (g2744)) + ((!g1285) & (g1437) & (g2713) & (g2714) & (!g2744)) + ((!g1285) & (g1437) & (g2713) & (g2714) & (g2744)) + ((g1285) & (!g1437) & (!g2713) & (g2714) & (g2744)) + ((g1285) & (!g1437) & (g2713) & (!g2714) & (!g2744)) + ((g1285) & (!g1437) & (g2713) & (!g2714) & (g2744)) + ((g1285) & (!g1437) & (g2713) & (g2714) & (!g2744)) + ((g1285) & (!g1437) & (g2713) & (g2714) & (g2744)) + ((g1285) & (g1437) & (!g2713) & (!g2714) & (g2744)) + ((g1285) & (g1437) & (!g2713) & (g2714) & (!g2744)) + ((g1285) & (g1437) & (!g2713) & (g2714) & (g2744)) + ((g1285) & (g1437) & (g2713) & (!g2714) & (!g2744)) + ((g1285) & (g1437) & (g2713) & (!g2714) & (g2744)) + ((g1285) & (g1437) & (g2713) & (g2714) & (!g2744)) + ((g1285) & (g1437) & (g2713) & (g2714) & (g2744)));
	assign g2746 = (((!g1154) & (!g1295) & (g2710) & (g2711) & (g2745)) + ((!g1154) & (g1295) & (g2710) & (!g2711) & (g2745)) + ((!g1154) & (g1295) & (g2710) & (g2711) & (!g2745)) + ((!g1154) & (g1295) & (g2710) & (g2711) & (g2745)) + ((g1154) & (!g1295) & (!g2710) & (g2711) & (g2745)) + ((g1154) & (!g1295) & (g2710) & (!g2711) & (!g2745)) + ((g1154) & (!g1295) & (g2710) & (!g2711) & (g2745)) + ((g1154) & (!g1295) & (g2710) & (g2711) & (!g2745)) + ((g1154) & (!g1295) & (g2710) & (g2711) & (g2745)) + ((g1154) & (g1295) & (!g2710) & (!g2711) & (g2745)) + ((g1154) & (g1295) & (!g2710) & (g2711) & (!g2745)) + ((g1154) & (g1295) & (!g2710) & (g2711) & (g2745)) + ((g1154) & (g1295) & (g2710) & (!g2711) & (!g2745)) + ((g1154) & (g1295) & (g2710) & (!g2711) & (g2745)) + ((g1154) & (g1295) & (g2710) & (g2711) & (!g2745)) + ((g1154) & (g1295) & (g2710) & (g2711) & (g2745)));
	assign g2747 = (((!g1030) & (!g1160) & (g2707) & (g2708) & (g2746)) + ((!g1030) & (g1160) & (g2707) & (!g2708) & (g2746)) + ((!g1030) & (g1160) & (g2707) & (g2708) & (!g2746)) + ((!g1030) & (g1160) & (g2707) & (g2708) & (g2746)) + ((g1030) & (!g1160) & (!g2707) & (g2708) & (g2746)) + ((g1030) & (!g1160) & (g2707) & (!g2708) & (!g2746)) + ((g1030) & (!g1160) & (g2707) & (!g2708) & (g2746)) + ((g1030) & (!g1160) & (g2707) & (g2708) & (!g2746)) + ((g1030) & (!g1160) & (g2707) & (g2708) & (g2746)) + ((g1030) & (g1160) & (!g2707) & (!g2708) & (g2746)) + ((g1030) & (g1160) & (!g2707) & (g2708) & (!g2746)) + ((g1030) & (g1160) & (!g2707) & (g2708) & (g2746)) + ((g1030) & (g1160) & (g2707) & (!g2708) & (!g2746)) + ((g1030) & (g1160) & (g2707) & (!g2708) & (g2746)) + ((g1030) & (g1160) & (g2707) & (g2708) & (!g2746)) + ((g1030) & (g1160) & (g2707) & (g2708) & (g2746)));
	assign g2748 = (((!g914) & (!g1032) & (g2704) & (g2705) & (g2747)) + ((!g914) & (g1032) & (g2704) & (!g2705) & (g2747)) + ((!g914) & (g1032) & (g2704) & (g2705) & (!g2747)) + ((!g914) & (g1032) & (g2704) & (g2705) & (g2747)) + ((g914) & (!g1032) & (!g2704) & (g2705) & (g2747)) + ((g914) & (!g1032) & (g2704) & (!g2705) & (!g2747)) + ((g914) & (!g1032) & (g2704) & (!g2705) & (g2747)) + ((g914) & (!g1032) & (g2704) & (g2705) & (!g2747)) + ((g914) & (!g1032) & (g2704) & (g2705) & (g2747)) + ((g914) & (g1032) & (!g2704) & (!g2705) & (g2747)) + ((g914) & (g1032) & (!g2704) & (g2705) & (!g2747)) + ((g914) & (g1032) & (!g2704) & (g2705) & (g2747)) + ((g914) & (g1032) & (g2704) & (!g2705) & (!g2747)) + ((g914) & (g1032) & (g2704) & (!g2705) & (g2747)) + ((g914) & (g1032) & (g2704) & (g2705) & (!g2747)) + ((g914) & (g1032) & (g2704) & (g2705) & (g2747)));
	assign g2749 = (((!g803) & (!g851) & (g2701) & (g2702) & (g2748)) + ((!g803) & (g851) & (g2701) & (!g2702) & (g2748)) + ((!g803) & (g851) & (g2701) & (g2702) & (!g2748)) + ((!g803) & (g851) & (g2701) & (g2702) & (g2748)) + ((g803) & (!g851) & (!g2701) & (g2702) & (g2748)) + ((g803) & (!g851) & (g2701) & (!g2702) & (!g2748)) + ((g803) & (!g851) & (g2701) & (!g2702) & (g2748)) + ((g803) & (!g851) & (g2701) & (g2702) & (!g2748)) + ((g803) & (!g851) & (g2701) & (g2702) & (g2748)) + ((g803) & (g851) & (!g2701) & (!g2702) & (g2748)) + ((g803) & (g851) & (!g2701) & (g2702) & (!g2748)) + ((g803) & (g851) & (!g2701) & (g2702) & (g2748)) + ((g803) & (g851) & (g2701) & (!g2702) & (!g2748)) + ((g803) & (g851) & (g2701) & (!g2702) & (g2748)) + ((g803) & (g851) & (g2701) & (g2702) & (!g2748)) + ((g803) & (g851) & (g2701) & (g2702) & (g2748)));
	assign g2750 = (((!g700) & (!g744) & (g2698) & (g2699) & (g2749)) + ((!g700) & (g744) & (g2698) & (!g2699) & (g2749)) + ((!g700) & (g744) & (g2698) & (g2699) & (!g2749)) + ((!g700) & (g744) & (g2698) & (g2699) & (g2749)) + ((g700) & (!g744) & (!g2698) & (g2699) & (g2749)) + ((g700) & (!g744) & (g2698) & (!g2699) & (!g2749)) + ((g700) & (!g744) & (g2698) & (!g2699) & (g2749)) + ((g700) & (!g744) & (g2698) & (g2699) & (!g2749)) + ((g700) & (!g744) & (g2698) & (g2699) & (g2749)) + ((g700) & (g744) & (!g2698) & (!g2699) & (g2749)) + ((g700) & (g744) & (!g2698) & (g2699) & (!g2749)) + ((g700) & (g744) & (!g2698) & (g2699) & (g2749)) + ((g700) & (g744) & (g2698) & (!g2699) & (!g2749)) + ((g700) & (g744) & (g2698) & (!g2699) & (g2749)) + ((g700) & (g744) & (g2698) & (g2699) & (!g2749)) + ((g700) & (g744) & (g2698) & (g2699) & (g2749)));
	assign g2751 = (((!g604) & (!g645) & (g2695) & (g2696) & (g2750)) + ((!g604) & (g645) & (g2695) & (!g2696) & (g2750)) + ((!g604) & (g645) & (g2695) & (g2696) & (!g2750)) + ((!g604) & (g645) & (g2695) & (g2696) & (g2750)) + ((g604) & (!g645) & (!g2695) & (g2696) & (g2750)) + ((g604) & (!g645) & (g2695) & (!g2696) & (!g2750)) + ((g604) & (!g645) & (g2695) & (!g2696) & (g2750)) + ((g604) & (!g645) & (g2695) & (g2696) & (!g2750)) + ((g604) & (!g645) & (g2695) & (g2696) & (g2750)) + ((g604) & (g645) & (!g2695) & (!g2696) & (g2750)) + ((g604) & (g645) & (!g2695) & (g2696) & (!g2750)) + ((g604) & (g645) & (!g2695) & (g2696) & (g2750)) + ((g604) & (g645) & (g2695) & (!g2696) & (!g2750)) + ((g604) & (g645) & (g2695) & (!g2696) & (g2750)) + ((g604) & (g645) & (g2695) & (g2696) & (!g2750)) + ((g604) & (g645) & (g2695) & (g2696) & (g2750)));
	assign g2752 = (((!g515) & (!g553) & (g2692) & (g2693) & (g2751)) + ((!g515) & (g553) & (g2692) & (!g2693) & (g2751)) + ((!g515) & (g553) & (g2692) & (g2693) & (!g2751)) + ((!g515) & (g553) & (g2692) & (g2693) & (g2751)) + ((g515) & (!g553) & (!g2692) & (g2693) & (g2751)) + ((g515) & (!g553) & (g2692) & (!g2693) & (!g2751)) + ((g515) & (!g553) & (g2692) & (!g2693) & (g2751)) + ((g515) & (!g553) & (g2692) & (g2693) & (!g2751)) + ((g515) & (!g553) & (g2692) & (g2693) & (g2751)) + ((g515) & (g553) & (!g2692) & (!g2693) & (g2751)) + ((g515) & (g553) & (!g2692) & (g2693) & (!g2751)) + ((g515) & (g553) & (!g2692) & (g2693) & (g2751)) + ((g515) & (g553) & (g2692) & (!g2693) & (!g2751)) + ((g515) & (g553) & (g2692) & (!g2693) & (g2751)) + ((g515) & (g553) & (g2692) & (g2693) & (!g2751)) + ((g515) & (g553) & (g2692) & (g2693) & (g2751)));
	assign g2753 = (((!g433) & (!g468) & (g2689) & (g2690) & (g2752)) + ((!g433) & (g468) & (g2689) & (!g2690) & (g2752)) + ((!g433) & (g468) & (g2689) & (g2690) & (!g2752)) + ((!g433) & (g468) & (g2689) & (g2690) & (g2752)) + ((g433) & (!g468) & (!g2689) & (g2690) & (g2752)) + ((g433) & (!g468) & (g2689) & (!g2690) & (!g2752)) + ((g433) & (!g468) & (g2689) & (!g2690) & (g2752)) + ((g433) & (!g468) & (g2689) & (g2690) & (!g2752)) + ((g433) & (!g468) & (g2689) & (g2690) & (g2752)) + ((g433) & (g468) & (!g2689) & (!g2690) & (g2752)) + ((g433) & (g468) & (!g2689) & (g2690) & (!g2752)) + ((g433) & (g468) & (!g2689) & (g2690) & (g2752)) + ((g433) & (g468) & (g2689) & (!g2690) & (!g2752)) + ((g433) & (g468) & (g2689) & (!g2690) & (g2752)) + ((g433) & (g468) & (g2689) & (g2690) & (!g2752)) + ((g433) & (g468) & (g2689) & (g2690) & (g2752)));
	assign g2754 = (((!g358) & (!g390) & (g2686) & (g2687) & (g2753)) + ((!g358) & (g390) & (g2686) & (!g2687) & (g2753)) + ((!g358) & (g390) & (g2686) & (g2687) & (!g2753)) + ((!g358) & (g390) & (g2686) & (g2687) & (g2753)) + ((g358) & (!g390) & (!g2686) & (g2687) & (g2753)) + ((g358) & (!g390) & (g2686) & (!g2687) & (!g2753)) + ((g358) & (!g390) & (g2686) & (!g2687) & (g2753)) + ((g358) & (!g390) & (g2686) & (g2687) & (!g2753)) + ((g358) & (!g390) & (g2686) & (g2687) & (g2753)) + ((g358) & (g390) & (!g2686) & (!g2687) & (g2753)) + ((g358) & (g390) & (!g2686) & (g2687) & (!g2753)) + ((g358) & (g390) & (!g2686) & (g2687) & (g2753)) + ((g358) & (g390) & (g2686) & (!g2687) & (!g2753)) + ((g358) & (g390) & (g2686) & (!g2687) & (g2753)) + ((g358) & (g390) & (g2686) & (g2687) & (!g2753)) + ((g358) & (g390) & (g2686) & (g2687) & (g2753)));
	assign g2755 = (((!g290) & (!g319) & (g2683) & (g2684) & (g2754)) + ((!g290) & (g319) & (g2683) & (!g2684) & (g2754)) + ((!g290) & (g319) & (g2683) & (g2684) & (!g2754)) + ((!g290) & (g319) & (g2683) & (g2684) & (g2754)) + ((g290) & (!g319) & (!g2683) & (g2684) & (g2754)) + ((g290) & (!g319) & (g2683) & (!g2684) & (!g2754)) + ((g290) & (!g319) & (g2683) & (!g2684) & (g2754)) + ((g290) & (!g319) & (g2683) & (g2684) & (!g2754)) + ((g290) & (!g319) & (g2683) & (g2684) & (g2754)) + ((g290) & (g319) & (!g2683) & (!g2684) & (g2754)) + ((g290) & (g319) & (!g2683) & (g2684) & (!g2754)) + ((g290) & (g319) & (!g2683) & (g2684) & (g2754)) + ((g290) & (g319) & (g2683) & (!g2684) & (!g2754)) + ((g290) & (g319) & (g2683) & (!g2684) & (g2754)) + ((g290) & (g319) & (g2683) & (g2684) & (!g2754)) + ((g290) & (g319) & (g2683) & (g2684) & (g2754)));
	assign g2756 = (((!g229) & (!g255) & (g2680) & (g2681) & (g2755)) + ((!g229) & (g255) & (g2680) & (!g2681) & (g2755)) + ((!g229) & (g255) & (g2680) & (g2681) & (!g2755)) + ((!g229) & (g255) & (g2680) & (g2681) & (g2755)) + ((g229) & (!g255) & (!g2680) & (g2681) & (g2755)) + ((g229) & (!g255) & (g2680) & (!g2681) & (!g2755)) + ((g229) & (!g255) & (g2680) & (!g2681) & (g2755)) + ((g229) & (!g255) & (g2680) & (g2681) & (!g2755)) + ((g229) & (!g255) & (g2680) & (g2681) & (g2755)) + ((g229) & (g255) & (!g2680) & (!g2681) & (g2755)) + ((g229) & (g255) & (!g2680) & (g2681) & (!g2755)) + ((g229) & (g255) & (!g2680) & (g2681) & (g2755)) + ((g229) & (g255) & (g2680) & (!g2681) & (!g2755)) + ((g229) & (g255) & (g2680) & (!g2681) & (g2755)) + ((g229) & (g255) & (g2680) & (g2681) & (!g2755)) + ((g229) & (g255) & (g2680) & (g2681) & (g2755)));
	assign g2757 = (((!g174) & (!g198) & (g2677) & (g2678) & (g2756)) + ((!g174) & (g198) & (g2677) & (!g2678) & (g2756)) + ((!g174) & (g198) & (g2677) & (g2678) & (!g2756)) + ((!g174) & (g198) & (g2677) & (g2678) & (g2756)) + ((g174) & (!g198) & (!g2677) & (g2678) & (g2756)) + ((g174) & (!g198) & (g2677) & (!g2678) & (!g2756)) + ((g174) & (!g198) & (g2677) & (!g2678) & (g2756)) + ((g174) & (!g198) & (g2677) & (g2678) & (!g2756)) + ((g174) & (!g198) & (g2677) & (g2678) & (g2756)) + ((g174) & (g198) & (!g2677) & (!g2678) & (g2756)) + ((g174) & (g198) & (!g2677) & (g2678) & (!g2756)) + ((g174) & (g198) & (!g2677) & (g2678) & (g2756)) + ((g174) & (g198) & (g2677) & (!g2678) & (!g2756)) + ((g174) & (g198) & (g2677) & (!g2678) & (g2756)) + ((g174) & (g198) & (g2677) & (g2678) & (!g2756)) + ((g174) & (g198) & (g2677) & (g2678) & (g2756)));
	assign g2758 = (((!g127) & (!g147) & (g2674) & (g2675) & (g2757)) + ((!g127) & (g147) & (g2674) & (!g2675) & (g2757)) + ((!g127) & (g147) & (g2674) & (g2675) & (!g2757)) + ((!g127) & (g147) & (g2674) & (g2675) & (g2757)) + ((g127) & (!g147) & (!g2674) & (g2675) & (g2757)) + ((g127) & (!g147) & (g2674) & (!g2675) & (!g2757)) + ((g127) & (!g147) & (g2674) & (!g2675) & (g2757)) + ((g127) & (!g147) & (g2674) & (g2675) & (!g2757)) + ((g127) & (!g147) & (g2674) & (g2675) & (g2757)) + ((g127) & (g147) & (!g2674) & (!g2675) & (g2757)) + ((g127) & (g147) & (!g2674) & (g2675) & (!g2757)) + ((g127) & (g147) & (!g2674) & (g2675) & (g2757)) + ((g127) & (g147) & (g2674) & (!g2675) & (!g2757)) + ((g127) & (g147) & (g2674) & (!g2675) & (g2757)) + ((g127) & (g147) & (g2674) & (g2675) & (!g2757)) + ((g127) & (g147) & (g2674) & (g2675) & (g2757)));
	assign g2759 = (((!g87) & (!g104) & (g2671) & (g2672) & (g2758)) + ((!g87) & (g104) & (g2671) & (!g2672) & (g2758)) + ((!g87) & (g104) & (g2671) & (g2672) & (!g2758)) + ((!g87) & (g104) & (g2671) & (g2672) & (g2758)) + ((g87) & (!g104) & (!g2671) & (g2672) & (g2758)) + ((g87) & (!g104) & (g2671) & (!g2672) & (!g2758)) + ((g87) & (!g104) & (g2671) & (!g2672) & (g2758)) + ((g87) & (!g104) & (g2671) & (g2672) & (!g2758)) + ((g87) & (!g104) & (g2671) & (g2672) & (g2758)) + ((g87) & (g104) & (!g2671) & (!g2672) & (g2758)) + ((g87) & (g104) & (!g2671) & (g2672) & (!g2758)) + ((g87) & (g104) & (!g2671) & (g2672) & (g2758)) + ((g87) & (g104) & (g2671) & (!g2672) & (!g2758)) + ((g87) & (g104) & (g2671) & (!g2672) & (g2758)) + ((g87) & (g104) & (g2671) & (g2672) & (!g2758)) + ((g87) & (g104) & (g2671) & (g2672) & (g2758)));
	assign g2760 = (((!g4) & (!g2665) & (!g2666) & (!g2653) & (!g2668)) + ((!g4) & (!g2665) & (!g2666) & (g2653) & (!g2668)) + ((!g4) & (!g2665) & (!g2666) & (g2653) & (g2668)) + ((!g4) & (!g2665) & (g2666) & (!g2653) & (g2668)) + ((!g4) & (g2665) & (g2666) & (!g2653) & (!g2668)) + ((!g4) & (g2665) & (g2666) & (!g2653) & (g2668)) + ((!g4) & (g2665) & (g2666) & (g2653) & (!g2668)) + ((!g4) & (g2665) & (g2666) & (g2653) & (g2668)) + ((g4) & (!g2665) & (g2666) & (!g2653) & (!g2668)) + ((g4) & (!g2665) & (g2666) & (!g2653) & (g2668)) + ((g4) & (!g2665) & (g2666) & (g2653) & (!g2668)) + ((g4) & (!g2665) & (g2666) & (g2653) & (g2668)) + ((g4) & (g2665) & (!g2666) & (!g2653) & (!g2668)) + ((g4) & (g2665) & (!g2666) & (g2653) & (!g2668)) + ((g4) & (g2665) & (!g2666) & (g2653) & (g2668)) + ((g4) & (g2665) & (g2666) & (!g2653) & (g2668)));
	assign g2761 = (((!g8) & (!g2656) & (g2664) & (!g2653) & (!g2668)) + ((!g8) & (!g2656) & (g2664) & (g2653) & (!g2668)) + ((!g8) & (!g2656) & (g2664) & (g2653) & (g2668)) + ((!g8) & (g2656) & (!g2664) & (!g2653) & (!g2668)) + ((!g8) & (g2656) & (!g2664) & (!g2653) & (g2668)) + ((!g8) & (g2656) & (!g2664) & (g2653) & (!g2668)) + ((!g8) & (g2656) & (!g2664) & (g2653) & (g2668)) + ((!g8) & (g2656) & (g2664) & (!g2653) & (g2668)) + ((g8) & (!g2656) & (!g2664) & (!g2653) & (!g2668)) + ((g8) & (!g2656) & (!g2664) & (g2653) & (!g2668)) + ((g8) & (!g2656) & (!g2664) & (g2653) & (g2668)) + ((g8) & (g2656) & (!g2664) & (!g2653) & (g2668)) + ((g8) & (g2656) & (g2664) & (!g2653) & (!g2668)) + ((g8) & (g2656) & (g2664) & (!g2653) & (g2668)) + ((g8) & (g2656) & (g2664) & (g2653) & (!g2668)) + ((g8) & (g2656) & (g2664) & (g2653) & (g2668)));
	assign g2762 = (((!g18) & (!g27) & (g2658) & (g2663)) + ((!g18) & (g27) & (!g2658) & (g2663)) + ((!g18) & (g27) & (g2658) & (!g2663)) + ((!g18) & (g27) & (g2658) & (g2663)) + ((g18) & (!g27) & (!g2658) & (!g2663)) + ((g18) & (!g27) & (!g2658) & (g2663)) + ((g18) & (!g27) & (g2658) & (!g2663)) + ((g18) & (g27) & (!g2658) & (!g2663)));
	assign g2763 = (((!g2657) & (!g2653) & (!g2668) & (g2762)) + ((!g2657) & (g2653) & (!g2668) & (g2762)) + ((!g2657) & (g2653) & (g2668) & (g2762)) + ((g2657) & (!g2653) & (!g2668) & (!g2762)) + ((g2657) & (!g2653) & (g2668) & (!g2762)) + ((g2657) & (!g2653) & (g2668) & (g2762)) + ((g2657) & (g2653) & (!g2668) & (!g2762)) + ((g2657) & (g2653) & (g2668) & (!g2762)));
	assign g2764 = (((!g27) & (!g2658) & (g2663) & (!g2653) & (!g2668)) + ((!g27) & (!g2658) & (g2663) & (g2653) & (!g2668)) + ((!g27) & (!g2658) & (g2663) & (g2653) & (g2668)) + ((!g27) & (g2658) & (!g2663) & (!g2653) & (!g2668)) + ((!g27) & (g2658) & (!g2663) & (!g2653) & (g2668)) + ((!g27) & (g2658) & (!g2663) & (g2653) & (!g2668)) + ((!g27) & (g2658) & (!g2663) & (g2653) & (g2668)) + ((!g27) & (g2658) & (g2663) & (!g2653) & (g2668)) + ((g27) & (!g2658) & (!g2663) & (!g2653) & (!g2668)) + ((g27) & (!g2658) & (!g2663) & (g2653) & (!g2668)) + ((g27) & (!g2658) & (!g2663) & (g2653) & (g2668)) + ((g27) & (g2658) & (!g2663) & (!g2653) & (g2668)) + ((g27) & (g2658) & (g2663) & (!g2653) & (!g2668)) + ((g27) & (g2658) & (g2663) & (!g2653) & (g2668)) + ((g27) & (g2658) & (g2663) & (g2653) & (!g2668)) + ((g27) & (g2658) & (g2663) & (g2653) & (g2668)));
	assign g2765 = (((!g39) & (!g54) & (g2660) & (g2662)) + ((!g39) & (g54) & (!g2660) & (g2662)) + ((!g39) & (g54) & (g2660) & (!g2662)) + ((!g39) & (g54) & (g2660) & (g2662)) + ((g39) & (!g54) & (!g2660) & (!g2662)) + ((g39) & (!g54) & (!g2660) & (g2662)) + ((g39) & (!g54) & (g2660) & (!g2662)) + ((g39) & (g54) & (!g2660) & (!g2662)));
	assign g2766 = (((!g2659) & (!g2653) & (!g2668) & (g2765)) + ((!g2659) & (g2653) & (!g2668) & (g2765)) + ((!g2659) & (g2653) & (g2668) & (g2765)) + ((g2659) & (!g2653) & (!g2668) & (!g2765)) + ((g2659) & (!g2653) & (g2668) & (!g2765)) + ((g2659) & (!g2653) & (g2668) & (g2765)) + ((g2659) & (g2653) & (!g2668) & (!g2765)) + ((g2659) & (g2653) & (g2668) & (!g2765)));
	assign g2767 = (((!g54) & (!g2660) & (g2662) & (!g2653) & (!g2668)) + ((!g54) & (!g2660) & (g2662) & (g2653) & (!g2668)) + ((!g54) & (!g2660) & (g2662) & (g2653) & (g2668)) + ((!g54) & (g2660) & (!g2662) & (!g2653) & (!g2668)) + ((!g54) & (g2660) & (!g2662) & (!g2653) & (g2668)) + ((!g54) & (g2660) & (!g2662) & (g2653) & (!g2668)) + ((!g54) & (g2660) & (!g2662) & (g2653) & (g2668)) + ((!g54) & (g2660) & (g2662) & (!g2653) & (g2668)) + ((g54) & (!g2660) & (!g2662) & (!g2653) & (!g2668)) + ((g54) & (!g2660) & (!g2662) & (g2653) & (!g2668)) + ((g54) & (!g2660) & (!g2662) & (g2653) & (g2668)) + ((g54) & (g2660) & (!g2662) & (!g2653) & (g2668)) + ((g54) & (g2660) & (g2662) & (!g2653) & (!g2668)) + ((g54) & (g2660) & (g2662) & (!g2653) & (g2668)) + ((g54) & (g2660) & (g2662) & (g2653) & (!g2668)) + ((g54) & (g2660) & (g2662) & (g2653) & (g2668)));
	assign g2768 = (((!g68) & (!g87) & (g2586) & (g2652)) + ((!g68) & (g87) & (!g2586) & (g2652)) + ((!g68) & (g87) & (g2586) & (!g2652)) + ((!g68) & (g87) & (g2586) & (g2652)) + ((g68) & (!g87) & (!g2586) & (!g2652)) + ((g68) & (!g87) & (!g2586) & (g2652)) + ((g68) & (!g87) & (g2586) & (!g2652)) + ((g68) & (g87) & (!g2586) & (!g2652)));
	assign g2769 = (((!g2661) & (!g2653) & (!g2668) & (g2768)) + ((!g2661) & (g2653) & (!g2668) & (g2768)) + ((!g2661) & (g2653) & (g2668) & (g2768)) + ((g2661) & (!g2653) & (!g2668) & (!g2768)) + ((g2661) & (!g2653) & (g2668) & (!g2768)) + ((g2661) & (!g2653) & (g2668) & (g2768)) + ((g2661) & (g2653) & (!g2668) & (!g2768)) + ((g2661) & (g2653) & (g2668) & (!g2768)));
	assign g2770 = (((!g54) & (!g68) & (g2769) & (g2669) & (g2759)) + ((!g54) & (g68) & (g2769) & (!g2669) & (g2759)) + ((!g54) & (g68) & (g2769) & (g2669) & (!g2759)) + ((!g54) & (g68) & (g2769) & (g2669) & (g2759)) + ((g54) & (!g68) & (!g2769) & (g2669) & (g2759)) + ((g54) & (!g68) & (g2769) & (!g2669) & (!g2759)) + ((g54) & (!g68) & (g2769) & (!g2669) & (g2759)) + ((g54) & (!g68) & (g2769) & (g2669) & (!g2759)) + ((g54) & (!g68) & (g2769) & (g2669) & (g2759)) + ((g54) & (g68) & (!g2769) & (!g2669) & (g2759)) + ((g54) & (g68) & (!g2769) & (g2669) & (!g2759)) + ((g54) & (g68) & (!g2769) & (g2669) & (g2759)) + ((g54) & (g68) & (g2769) & (!g2669) & (!g2759)) + ((g54) & (g68) & (g2769) & (!g2669) & (g2759)) + ((g54) & (g68) & (g2769) & (g2669) & (!g2759)) + ((g54) & (g68) & (g2769) & (g2669) & (g2759)));
	assign g2771 = (((!g27) & (!g39) & (g2766) & (g2767) & (g2770)) + ((!g27) & (g39) & (g2766) & (!g2767) & (g2770)) + ((!g27) & (g39) & (g2766) & (g2767) & (!g2770)) + ((!g27) & (g39) & (g2766) & (g2767) & (g2770)) + ((g27) & (!g39) & (!g2766) & (g2767) & (g2770)) + ((g27) & (!g39) & (g2766) & (!g2767) & (!g2770)) + ((g27) & (!g39) & (g2766) & (!g2767) & (g2770)) + ((g27) & (!g39) & (g2766) & (g2767) & (!g2770)) + ((g27) & (!g39) & (g2766) & (g2767) & (g2770)) + ((g27) & (g39) & (!g2766) & (!g2767) & (g2770)) + ((g27) & (g39) & (!g2766) & (g2767) & (!g2770)) + ((g27) & (g39) & (!g2766) & (g2767) & (g2770)) + ((g27) & (g39) & (g2766) & (!g2767) & (!g2770)) + ((g27) & (g39) & (g2766) & (!g2767) & (g2770)) + ((g27) & (g39) & (g2766) & (g2767) & (!g2770)) + ((g27) & (g39) & (g2766) & (g2767) & (g2770)));
	assign g2772 = (((!g8) & (!g18) & (g2763) & (g2764) & (g2771)) + ((!g8) & (g18) & (g2763) & (!g2764) & (g2771)) + ((!g8) & (g18) & (g2763) & (g2764) & (!g2771)) + ((!g8) & (g18) & (g2763) & (g2764) & (g2771)) + ((g8) & (!g18) & (!g2763) & (g2764) & (g2771)) + ((g8) & (!g18) & (g2763) & (!g2764) & (!g2771)) + ((g8) & (!g18) & (g2763) & (!g2764) & (g2771)) + ((g8) & (!g18) & (g2763) & (g2764) & (!g2771)) + ((g8) & (!g18) & (g2763) & (g2764) & (g2771)) + ((g8) & (g18) & (!g2763) & (!g2764) & (g2771)) + ((g8) & (g18) & (!g2763) & (g2764) & (!g2771)) + ((g8) & (g18) & (!g2763) & (g2764) & (g2771)) + ((g8) & (g18) & (g2763) & (!g2764) & (!g2771)) + ((g8) & (g18) & (g2763) & (!g2764) & (g2771)) + ((g8) & (g18) & (g2763) & (g2764) & (!g2771)) + ((g8) & (g18) & (g2763) & (g2764) & (g2771)));
	assign g2773 = (((!g2) & (!g8) & (g2656) & (g2664)) + ((!g2) & (g8) & (!g2656) & (g2664)) + ((!g2) & (g8) & (g2656) & (!g2664)) + ((!g2) & (g8) & (g2656) & (g2664)) + ((g2) & (!g8) & (!g2656) & (!g2664)) + ((g2) & (!g8) & (!g2656) & (g2664)) + ((g2) & (!g8) & (g2656) & (!g2664)) + ((g2) & (g8) & (!g2656) & (!g2664)));
	assign g2774 = (((!g2655) & (!g2653) & (!g2668) & (g2773)) + ((!g2655) & (g2653) & (!g2668) & (g2773)) + ((!g2655) & (g2653) & (g2668) & (g2773)) + ((g2655) & (!g2653) & (!g2668) & (!g2773)) + ((g2655) & (!g2653) & (g2668) & (!g2773)) + ((g2655) & (!g2653) & (g2668) & (g2773)) + ((g2655) & (g2653) & (!g2668) & (!g2773)) + ((g2655) & (g2653) & (g2668) & (!g2773)));
	assign g2775 = (((!g4) & (!g2) & (!g2761) & (!g2772) & (g2774)) + ((!g4) & (!g2) & (!g2761) & (g2772) & (g2774)) + ((!g4) & (!g2) & (g2761) & (!g2772) & (g2774)) + ((!g4) & (!g2) & (g2761) & (g2772) & (!g2774)) + ((!g4) & (!g2) & (g2761) & (g2772) & (g2774)) + ((!g4) & (g2) & (!g2761) & (!g2772) & (g2774)) + ((!g4) & (g2) & (!g2761) & (g2772) & (!g2774)) + ((!g4) & (g2) & (!g2761) & (g2772) & (g2774)) + ((!g4) & (g2) & (g2761) & (!g2772) & (!g2774)) + ((!g4) & (g2) & (g2761) & (!g2772) & (g2774)) + ((!g4) & (g2) & (g2761) & (g2772) & (!g2774)) + ((!g4) & (g2) & (g2761) & (g2772) & (g2774)) + ((g4) & (!g2) & (g2761) & (g2772) & (g2774)) + ((g4) & (g2) & (!g2761) & (g2772) & (g2774)) + ((g4) & (g2) & (g2761) & (!g2772) & (g2774)) + ((g4) & (g2) & (g2761) & (g2772) & (g2774)));
	assign g2776 = (((!g4) & (!g2665) & (g2666)) + ((!g4) & (g2665) & (!g2666)) + ((!g4) & (g2665) & (g2666)) + ((g4) & (g2665) & (g2666)));
	assign g2777 = (((!g2654) & (!g2776) & (!g2653) & (!g2668)) + ((!g2654) & (!g2776) & (g2653) & (!g2668)) + ((!g2654) & (!g2776) & (g2653) & (g2668)) + ((g2654) & (g2776) & (!g2653) & (!g2668)) + ((g2654) & (g2776) & (!g2653) & (g2668)) + ((g2654) & (g2776) & (g2653) & (!g2668)) + ((g2654) & (g2776) & (g2653) & (g2668)));
	assign g2778 = (((!g1) & (g2654) & (!g2776) & (!g2653) & (g2668)) + ((!g1) & (g2654) & (g2776) & (!g2653) & (g2668)) + ((g1) & (!g2654) & (g2776) & (g2653) & (!g2668)) + ((g1) & (!g2654) & (g2776) & (g2653) & (g2668)) + ((g1) & (g2654) & (!g2776) & (!g2653) & (!g2668)) + ((g1) & (g2654) & (!g2776) & (!g2653) & (g2668)) + ((g1) & (g2654) & (!g2776) & (g2653) & (!g2668)) + ((g1) & (g2654) & (!g2776) & (g2653) & (g2668)) + ((g1) & (g2654) & (g2776) & (!g2653) & (g2668)));
	assign g2779 = (((!g1) & (!g2760) & (!g2775) & (!g2777) & (!g2778)) + ((g1) & (!g2760) & (!g2775) & (!g2777) & (!g2778)) + ((g1) & (!g2760) & (!g2775) & (g2777) & (!g2778)) + ((g1) & (!g2760) & (g2775) & (!g2777) & (!g2778)) + ((g1) & (!g2760) & (g2775) & (g2777) & (!g2778)) + ((g1) & (g2760) & (!g2775) & (!g2777) & (!g2778)) + ((g1) & (g2760) & (!g2775) & (g2777) & (!g2778)));
	assign g2780 = (((!g68) & (!g2669) & (g2759) & (!g2779)) + ((!g68) & (g2669) & (!g2759) & (!g2779)) + ((!g68) & (g2669) & (!g2759) & (g2779)) + ((!g68) & (g2669) & (g2759) & (g2779)) + ((g68) & (!g2669) & (!g2759) & (!g2779)) + ((g68) & (g2669) & (!g2759) & (g2779)) + ((g68) & (g2669) & (g2759) & (!g2779)) + ((g68) & (g2669) & (g2759) & (g2779)));
	assign g2781 = (((!g87) & (!g104) & (!g2671) & (g2672) & (g2758) & (!g2779)) + ((!g87) & (!g104) & (g2671) & (!g2672) & (!g2758) & (!g2779)) + ((!g87) & (!g104) & (g2671) & (!g2672) & (!g2758) & (g2779)) + ((!g87) & (!g104) & (g2671) & (!g2672) & (g2758) & (!g2779)) + ((!g87) & (!g104) & (g2671) & (!g2672) & (g2758) & (g2779)) + ((!g87) & (!g104) & (g2671) & (g2672) & (!g2758) & (!g2779)) + ((!g87) & (!g104) & (g2671) & (g2672) & (!g2758) & (g2779)) + ((!g87) & (!g104) & (g2671) & (g2672) & (g2758) & (g2779)) + ((!g87) & (g104) & (!g2671) & (!g2672) & (g2758) & (!g2779)) + ((!g87) & (g104) & (!g2671) & (g2672) & (!g2758) & (!g2779)) + ((!g87) & (g104) & (!g2671) & (g2672) & (g2758) & (!g2779)) + ((!g87) & (g104) & (g2671) & (!g2672) & (!g2758) & (!g2779)) + ((!g87) & (g104) & (g2671) & (!g2672) & (!g2758) & (g2779)) + ((!g87) & (g104) & (g2671) & (!g2672) & (g2758) & (g2779)) + ((!g87) & (g104) & (g2671) & (g2672) & (!g2758) & (g2779)) + ((!g87) & (g104) & (g2671) & (g2672) & (g2758) & (g2779)) + ((g87) & (!g104) & (!g2671) & (!g2672) & (!g2758) & (!g2779)) + ((g87) & (!g104) & (!g2671) & (!g2672) & (g2758) & (!g2779)) + ((g87) & (!g104) & (!g2671) & (g2672) & (!g2758) & (!g2779)) + ((g87) & (!g104) & (g2671) & (!g2672) & (!g2758) & (g2779)) + ((g87) & (!g104) & (g2671) & (!g2672) & (g2758) & (g2779)) + ((g87) & (!g104) & (g2671) & (g2672) & (!g2758) & (g2779)) + ((g87) & (!g104) & (g2671) & (g2672) & (g2758) & (!g2779)) + ((g87) & (!g104) & (g2671) & (g2672) & (g2758) & (g2779)) + ((g87) & (g104) & (!g2671) & (!g2672) & (!g2758) & (!g2779)) + ((g87) & (g104) & (g2671) & (!g2672) & (!g2758) & (g2779)) + ((g87) & (g104) & (g2671) & (!g2672) & (g2758) & (!g2779)) + ((g87) & (g104) & (g2671) & (!g2672) & (g2758) & (g2779)) + ((g87) & (g104) & (g2671) & (g2672) & (!g2758) & (!g2779)) + ((g87) & (g104) & (g2671) & (g2672) & (!g2758) & (g2779)) + ((g87) & (g104) & (g2671) & (g2672) & (g2758) & (!g2779)) + ((g87) & (g104) & (g2671) & (g2672) & (g2758) & (g2779)));
	assign g2782 = (((!g104) & (!g2672) & (g2758) & (!g2779)) + ((!g104) & (g2672) & (!g2758) & (!g2779)) + ((!g104) & (g2672) & (!g2758) & (g2779)) + ((!g104) & (g2672) & (g2758) & (g2779)) + ((g104) & (!g2672) & (!g2758) & (!g2779)) + ((g104) & (g2672) & (!g2758) & (g2779)) + ((g104) & (g2672) & (g2758) & (!g2779)) + ((g104) & (g2672) & (g2758) & (g2779)));
	assign g2783 = (((!g127) & (!g147) & (!g2674) & (g2675) & (g2757) & (!g2779)) + ((!g127) & (!g147) & (g2674) & (!g2675) & (!g2757) & (!g2779)) + ((!g127) & (!g147) & (g2674) & (!g2675) & (!g2757) & (g2779)) + ((!g127) & (!g147) & (g2674) & (!g2675) & (g2757) & (!g2779)) + ((!g127) & (!g147) & (g2674) & (!g2675) & (g2757) & (g2779)) + ((!g127) & (!g147) & (g2674) & (g2675) & (!g2757) & (!g2779)) + ((!g127) & (!g147) & (g2674) & (g2675) & (!g2757) & (g2779)) + ((!g127) & (!g147) & (g2674) & (g2675) & (g2757) & (g2779)) + ((!g127) & (g147) & (!g2674) & (!g2675) & (g2757) & (!g2779)) + ((!g127) & (g147) & (!g2674) & (g2675) & (!g2757) & (!g2779)) + ((!g127) & (g147) & (!g2674) & (g2675) & (g2757) & (!g2779)) + ((!g127) & (g147) & (g2674) & (!g2675) & (!g2757) & (!g2779)) + ((!g127) & (g147) & (g2674) & (!g2675) & (!g2757) & (g2779)) + ((!g127) & (g147) & (g2674) & (!g2675) & (g2757) & (g2779)) + ((!g127) & (g147) & (g2674) & (g2675) & (!g2757) & (g2779)) + ((!g127) & (g147) & (g2674) & (g2675) & (g2757) & (g2779)) + ((g127) & (!g147) & (!g2674) & (!g2675) & (!g2757) & (!g2779)) + ((g127) & (!g147) & (!g2674) & (!g2675) & (g2757) & (!g2779)) + ((g127) & (!g147) & (!g2674) & (g2675) & (!g2757) & (!g2779)) + ((g127) & (!g147) & (g2674) & (!g2675) & (!g2757) & (g2779)) + ((g127) & (!g147) & (g2674) & (!g2675) & (g2757) & (g2779)) + ((g127) & (!g147) & (g2674) & (g2675) & (!g2757) & (g2779)) + ((g127) & (!g147) & (g2674) & (g2675) & (g2757) & (!g2779)) + ((g127) & (!g147) & (g2674) & (g2675) & (g2757) & (g2779)) + ((g127) & (g147) & (!g2674) & (!g2675) & (!g2757) & (!g2779)) + ((g127) & (g147) & (g2674) & (!g2675) & (!g2757) & (g2779)) + ((g127) & (g147) & (g2674) & (!g2675) & (g2757) & (!g2779)) + ((g127) & (g147) & (g2674) & (!g2675) & (g2757) & (g2779)) + ((g127) & (g147) & (g2674) & (g2675) & (!g2757) & (!g2779)) + ((g127) & (g147) & (g2674) & (g2675) & (!g2757) & (g2779)) + ((g127) & (g147) & (g2674) & (g2675) & (g2757) & (!g2779)) + ((g127) & (g147) & (g2674) & (g2675) & (g2757) & (g2779)));
	assign g2784 = (((!g147) & (!g2675) & (g2757) & (!g2779)) + ((!g147) & (g2675) & (!g2757) & (!g2779)) + ((!g147) & (g2675) & (!g2757) & (g2779)) + ((!g147) & (g2675) & (g2757) & (g2779)) + ((g147) & (!g2675) & (!g2757) & (!g2779)) + ((g147) & (g2675) & (!g2757) & (g2779)) + ((g147) & (g2675) & (g2757) & (!g2779)) + ((g147) & (g2675) & (g2757) & (g2779)));
	assign g2785 = (((!g174) & (!g198) & (!g2677) & (g2678) & (g2756) & (!g2779)) + ((!g174) & (!g198) & (g2677) & (!g2678) & (!g2756) & (!g2779)) + ((!g174) & (!g198) & (g2677) & (!g2678) & (!g2756) & (g2779)) + ((!g174) & (!g198) & (g2677) & (!g2678) & (g2756) & (!g2779)) + ((!g174) & (!g198) & (g2677) & (!g2678) & (g2756) & (g2779)) + ((!g174) & (!g198) & (g2677) & (g2678) & (!g2756) & (!g2779)) + ((!g174) & (!g198) & (g2677) & (g2678) & (!g2756) & (g2779)) + ((!g174) & (!g198) & (g2677) & (g2678) & (g2756) & (g2779)) + ((!g174) & (g198) & (!g2677) & (!g2678) & (g2756) & (!g2779)) + ((!g174) & (g198) & (!g2677) & (g2678) & (!g2756) & (!g2779)) + ((!g174) & (g198) & (!g2677) & (g2678) & (g2756) & (!g2779)) + ((!g174) & (g198) & (g2677) & (!g2678) & (!g2756) & (!g2779)) + ((!g174) & (g198) & (g2677) & (!g2678) & (!g2756) & (g2779)) + ((!g174) & (g198) & (g2677) & (!g2678) & (g2756) & (g2779)) + ((!g174) & (g198) & (g2677) & (g2678) & (!g2756) & (g2779)) + ((!g174) & (g198) & (g2677) & (g2678) & (g2756) & (g2779)) + ((g174) & (!g198) & (!g2677) & (!g2678) & (!g2756) & (!g2779)) + ((g174) & (!g198) & (!g2677) & (!g2678) & (g2756) & (!g2779)) + ((g174) & (!g198) & (!g2677) & (g2678) & (!g2756) & (!g2779)) + ((g174) & (!g198) & (g2677) & (!g2678) & (!g2756) & (g2779)) + ((g174) & (!g198) & (g2677) & (!g2678) & (g2756) & (g2779)) + ((g174) & (!g198) & (g2677) & (g2678) & (!g2756) & (g2779)) + ((g174) & (!g198) & (g2677) & (g2678) & (g2756) & (!g2779)) + ((g174) & (!g198) & (g2677) & (g2678) & (g2756) & (g2779)) + ((g174) & (g198) & (!g2677) & (!g2678) & (!g2756) & (!g2779)) + ((g174) & (g198) & (g2677) & (!g2678) & (!g2756) & (g2779)) + ((g174) & (g198) & (g2677) & (!g2678) & (g2756) & (!g2779)) + ((g174) & (g198) & (g2677) & (!g2678) & (g2756) & (g2779)) + ((g174) & (g198) & (g2677) & (g2678) & (!g2756) & (!g2779)) + ((g174) & (g198) & (g2677) & (g2678) & (!g2756) & (g2779)) + ((g174) & (g198) & (g2677) & (g2678) & (g2756) & (!g2779)) + ((g174) & (g198) & (g2677) & (g2678) & (g2756) & (g2779)));
	assign g2786 = (((!g198) & (!g2678) & (g2756) & (!g2779)) + ((!g198) & (g2678) & (!g2756) & (!g2779)) + ((!g198) & (g2678) & (!g2756) & (g2779)) + ((!g198) & (g2678) & (g2756) & (g2779)) + ((g198) & (!g2678) & (!g2756) & (!g2779)) + ((g198) & (g2678) & (!g2756) & (g2779)) + ((g198) & (g2678) & (g2756) & (!g2779)) + ((g198) & (g2678) & (g2756) & (g2779)));
	assign g2787 = (((!g229) & (!g255) & (!g2680) & (g2681) & (g2755) & (!g2779)) + ((!g229) & (!g255) & (g2680) & (!g2681) & (!g2755) & (!g2779)) + ((!g229) & (!g255) & (g2680) & (!g2681) & (!g2755) & (g2779)) + ((!g229) & (!g255) & (g2680) & (!g2681) & (g2755) & (!g2779)) + ((!g229) & (!g255) & (g2680) & (!g2681) & (g2755) & (g2779)) + ((!g229) & (!g255) & (g2680) & (g2681) & (!g2755) & (!g2779)) + ((!g229) & (!g255) & (g2680) & (g2681) & (!g2755) & (g2779)) + ((!g229) & (!g255) & (g2680) & (g2681) & (g2755) & (g2779)) + ((!g229) & (g255) & (!g2680) & (!g2681) & (g2755) & (!g2779)) + ((!g229) & (g255) & (!g2680) & (g2681) & (!g2755) & (!g2779)) + ((!g229) & (g255) & (!g2680) & (g2681) & (g2755) & (!g2779)) + ((!g229) & (g255) & (g2680) & (!g2681) & (!g2755) & (!g2779)) + ((!g229) & (g255) & (g2680) & (!g2681) & (!g2755) & (g2779)) + ((!g229) & (g255) & (g2680) & (!g2681) & (g2755) & (g2779)) + ((!g229) & (g255) & (g2680) & (g2681) & (!g2755) & (g2779)) + ((!g229) & (g255) & (g2680) & (g2681) & (g2755) & (g2779)) + ((g229) & (!g255) & (!g2680) & (!g2681) & (!g2755) & (!g2779)) + ((g229) & (!g255) & (!g2680) & (!g2681) & (g2755) & (!g2779)) + ((g229) & (!g255) & (!g2680) & (g2681) & (!g2755) & (!g2779)) + ((g229) & (!g255) & (g2680) & (!g2681) & (!g2755) & (g2779)) + ((g229) & (!g255) & (g2680) & (!g2681) & (g2755) & (g2779)) + ((g229) & (!g255) & (g2680) & (g2681) & (!g2755) & (g2779)) + ((g229) & (!g255) & (g2680) & (g2681) & (g2755) & (!g2779)) + ((g229) & (!g255) & (g2680) & (g2681) & (g2755) & (g2779)) + ((g229) & (g255) & (!g2680) & (!g2681) & (!g2755) & (!g2779)) + ((g229) & (g255) & (g2680) & (!g2681) & (!g2755) & (g2779)) + ((g229) & (g255) & (g2680) & (!g2681) & (g2755) & (!g2779)) + ((g229) & (g255) & (g2680) & (!g2681) & (g2755) & (g2779)) + ((g229) & (g255) & (g2680) & (g2681) & (!g2755) & (!g2779)) + ((g229) & (g255) & (g2680) & (g2681) & (!g2755) & (g2779)) + ((g229) & (g255) & (g2680) & (g2681) & (g2755) & (!g2779)) + ((g229) & (g255) & (g2680) & (g2681) & (g2755) & (g2779)));
	assign g2788 = (((!g255) & (!g2681) & (g2755) & (!g2779)) + ((!g255) & (g2681) & (!g2755) & (!g2779)) + ((!g255) & (g2681) & (!g2755) & (g2779)) + ((!g255) & (g2681) & (g2755) & (g2779)) + ((g255) & (!g2681) & (!g2755) & (!g2779)) + ((g255) & (g2681) & (!g2755) & (g2779)) + ((g255) & (g2681) & (g2755) & (!g2779)) + ((g255) & (g2681) & (g2755) & (g2779)));
	assign g2789 = (((!g290) & (!g319) & (!g2683) & (g2684) & (g2754) & (!g2779)) + ((!g290) & (!g319) & (g2683) & (!g2684) & (!g2754) & (!g2779)) + ((!g290) & (!g319) & (g2683) & (!g2684) & (!g2754) & (g2779)) + ((!g290) & (!g319) & (g2683) & (!g2684) & (g2754) & (!g2779)) + ((!g290) & (!g319) & (g2683) & (!g2684) & (g2754) & (g2779)) + ((!g290) & (!g319) & (g2683) & (g2684) & (!g2754) & (!g2779)) + ((!g290) & (!g319) & (g2683) & (g2684) & (!g2754) & (g2779)) + ((!g290) & (!g319) & (g2683) & (g2684) & (g2754) & (g2779)) + ((!g290) & (g319) & (!g2683) & (!g2684) & (g2754) & (!g2779)) + ((!g290) & (g319) & (!g2683) & (g2684) & (!g2754) & (!g2779)) + ((!g290) & (g319) & (!g2683) & (g2684) & (g2754) & (!g2779)) + ((!g290) & (g319) & (g2683) & (!g2684) & (!g2754) & (!g2779)) + ((!g290) & (g319) & (g2683) & (!g2684) & (!g2754) & (g2779)) + ((!g290) & (g319) & (g2683) & (!g2684) & (g2754) & (g2779)) + ((!g290) & (g319) & (g2683) & (g2684) & (!g2754) & (g2779)) + ((!g290) & (g319) & (g2683) & (g2684) & (g2754) & (g2779)) + ((g290) & (!g319) & (!g2683) & (!g2684) & (!g2754) & (!g2779)) + ((g290) & (!g319) & (!g2683) & (!g2684) & (g2754) & (!g2779)) + ((g290) & (!g319) & (!g2683) & (g2684) & (!g2754) & (!g2779)) + ((g290) & (!g319) & (g2683) & (!g2684) & (!g2754) & (g2779)) + ((g290) & (!g319) & (g2683) & (!g2684) & (g2754) & (g2779)) + ((g290) & (!g319) & (g2683) & (g2684) & (!g2754) & (g2779)) + ((g290) & (!g319) & (g2683) & (g2684) & (g2754) & (!g2779)) + ((g290) & (!g319) & (g2683) & (g2684) & (g2754) & (g2779)) + ((g290) & (g319) & (!g2683) & (!g2684) & (!g2754) & (!g2779)) + ((g290) & (g319) & (g2683) & (!g2684) & (!g2754) & (g2779)) + ((g290) & (g319) & (g2683) & (!g2684) & (g2754) & (!g2779)) + ((g290) & (g319) & (g2683) & (!g2684) & (g2754) & (g2779)) + ((g290) & (g319) & (g2683) & (g2684) & (!g2754) & (!g2779)) + ((g290) & (g319) & (g2683) & (g2684) & (!g2754) & (g2779)) + ((g290) & (g319) & (g2683) & (g2684) & (g2754) & (!g2779)) + ((g290) & (g319) & (g2683) & (g2684) & (g2754) & (g2779)));
	assign g2790 = (((!g319) & (!g2684) & (g2754) & (!g2779)) + ((!g319) & (g2684) & (!g2754) & (!g2779)) + ((!g319) & (g2684) & (!g2754) & (g2779)) + ((!g319) & (g2684) & (g2754) & (g2779)) + ((g319) & (!g2684) & (!g2754) & (!g2779)) + ((g319) & (g2684) & (!g2754) & (g2779)) + ((g319) & (g2684) & (g2754) & (!g2779)) + ((g319) & (g2684) & (g2754) & (g2779)));
	assign g2791 = (((!g358) & (!g390) & (!g2686) & (g2687) & (g2753) & (!g2779)) + ((!g358) & (!g390) & (g2686) & (!g2687) & (!g2753) & (!g2779)) + ((!g358) & (!g390) & (g2686) & (!g2687) & (!g2753) & (g2779)) + ((!g358) & (!g390) & (g2686) & (!g2687) & (g2753) & (!g2779)) + ((!g358) & (!g390) & (g2686) & (!g2687) & (g2753) & (g2779)) + ((!g358) & (!g390) & (g2686) & (g2687) & (!g2753) & (!g2779)) + ((!g358) & (!g390) & (g2686) & (g2687) & (!g2753) & (g2779)) + ((!g358) & (!g390) & (g2686) & (g2687) & (g2753) & (g2779)) + ((!g358) & (g390) & (!g2686) & (!g2687) & (g2753) & (!g2779)) + ((!g358) & (g390) & (!g2686) & (g2687) & (!g2753) & (!g2779)) + ((!g358) & (g390) & (!g2686) & (g2687) & (g2753) & (!g2779)) + ((!g358) & (g390) & (g2686) & (!g2687) & (!g2753) & (!g2779)) + ((!g358) & (g390) & (g2686) & (!g2687) & (!g2753) & (g2779)) + ((!g358) & (g390) & (g2686) & (!g2687) & (g2753) & (g2779)) + ((!g358) & (g390) & (g2686) & (g2687) & (!g2753) & (g2779)) + ((!g358) & (g390) & (g2686) & (g2687) & (g2753) & (g2779)) + ((g358) & (!g390) & (!g2686) & (!g2687) & (!g2753) & (!g2779)) + ((g358) & (!g390) & (!g2686) & (!g2687) & (g2753) & (!g2779)) + ((g358) & (!g390) & (!g2686) & (g2687) & (!g2753) & (!g2779)) + ((g358) & (!g390) & (g2686) & (!g2687) & (!g2753) & (g2779)) + ((g358) & (!g390) & (g2686) & (!g2687) & (g2753) & (g2779)) + ((g358) & (!g390) & (g2686) & (g2687) & (!g2753) & (g2779)) + ((g358) & (!g390) & (g2686) & (g2687) & (g2753) & (!g2779)) + ((g358) & (!g390) & (g2686) & (g2687) & (g2753) & (g2779)) + ((g358) & (g390) & (!g2686) & (!g2687) & (!g2753) & (!g2779)) + ((g358) & (g390) & (g2686) & (!g2687) & (!g2753) & (g2779)) + ((g358) & (g390) & (g2686) & (!g2687) & (g2753) & (!g2779)) + ((g358) & (g390) & (g2686) & (!g2687) & (g2753) & (g2779)) + ((g358) & (g390) & (g2686) & (g2687) & (!g2753) & (!g2779)) + ((g358) & (g390) & (g2686) & (g2687) & (!g2753) & (g2779)) + ((g358) & (g390) & (g2686) & (g2687) & (g2753) & (!g2779)) + ((g358) & (g390) & (g2686) & (g2687) & (g2753) & (g2779)));
	assign g2792 = (((!g390) & (!g2687) & (g2753) & (!g2779)) + ((!g390) & (g2687) & (!g2753) & (!g2779)) + ((!g390) & (g2687) & (!g2753) & (g2779)) + ((!g390) & (g2687) & (g2753) & (g2779)) + ((g390) & (!g2687) & (!g2753) & (!g2779)) + ((g390) & (g2687) & (!g2753) & (g2779)) + ((g390) & (g2687) & (g2753) & (!g2779)) + ((g390) & (g2687) & (g2753) & (g2779)));
	assign g2793 = (((!g433) & (!g468) & (!g2689) & (g2690) & (g2752) & (!g2779)) + ((!g433) & (!g468) & (g2689) & (!g2690) & (!g2752) & (!g2779)) + ((!g433) & (!g468) & (g2689) & (!g2690) & (!g2752) & (g2779)) + ((!g433) & (!g468) & (g2689) & (!g2690) & (g2752) & (!g2779)) + ((!g433) & (!g468) & (g2689) & (!g2690) & (g2752) & (g2779)) + ((!g433) & (!g468) & (g2689) & (g2690) & (!g2752) & (!g2779)) + ((!g433) & (!g468) & (g2689) & (g2690) & (!g2752) & (g2779)) + ((!g433) & (!g468) & (g2689) & (g2690) & (g2752) & (g2779)) + ((!g433) & (g468) & (!g2689) & (!g2690) & (g2752) & (!g2779)) + ((!g433) & (g468) & (!g2689) & (g2690) & (!g2752) & (!g2779)) + ((!g433) & (g468) & (!g2689) & (g2690) & (g2752) & (!g2779)) + ((!g433) & (g468) & (g2689) & (!g2690) & (!g2752) & (!g2779)) + ((!g433) & (g468) & (g2689) & (!g2690) & (!g2752) & (g2779)) + ((!g433) & (g468) & (g2689) & (!g2690) & (g2752) & (g2779)) + ((!g433) & (g468) & (g2689) & (g2690) & (!g2752) & (g2779)) + ((!g433) & (g468) & (g2689) & (g2690) & (g2752) & (g2779)) + ((g433) & (!g468) & (!g2689) & (!g2690) & (!g2752) & (!g2779)) + ((g433) & (!g468) & (!g2689) & (!g2690) & (g2752) & (!g2779)) + ((g433) & (!g468) & (!g2689) & (g2690) & (!g2752) & (!g2779)) + ((g433) & (!g468) & (g2689) & (!g2690) & (!g2752) & (g2779)) + ((g433) & (!g468) & (g2689) & (!g2690) & (g2752) & (g2779)) + ((g433) & (!g468) & (g2689) & (g2690) & (!g2752) & (g2779)) + ((g433) & (!g468) & (g2689) & (g2690) & (g2752) & (!g2779)) + ((g433) & (!g468) & (g2689) & (g2690) & (g2752) & (g2779)) + ((g433) & (g468) & (!g2689) & (!g2690) & (!g2752) & (!g2779)) + ((g433) & (g468) & (g2689) & (!g2690) & (!g2752) & (g2779)) + ((g433) & (g468) & (g2689) & (!g2690) & (g2752) & (!g2779)) + ((g433) & (g468) & (g2689) & (!g2690) & (g2752) & (g2779)) + ((g433) & (g468) & (g2689) & (g2690) & (!g2752) & (!g2779)) + ((g433) & (g468) & (g2689) & (g2690) & (!g2752) & (g2779)) + ((g433) & (g468) & (g2689) & (g2690) & (g2752) & (!g2779)) + ((g433) & (g468) & (g2689) & (g2690) & (g2752) & (g2779)));
	assign g2794 = (((!g468) & (!g2690) & (g2752) & (!g2779)) + ((!g468) & (g2690) & (!g2752) & (!g2779)) + ((!g468) & (g2690) & (!g2752) & (g2779)) + ((!g468) & (g2690) & (g2752) & (g2779)) + ((g468) & (!g2690) & (!g2752) & (!g2779)) + ((g468) & (g2690) & (!g2752) & (g2779)) + ((g468) & (g2690) & (g2752) & (!g2779)) + ((g468) & (g2690) & (g2752) & (g2779)));
	assign g2795 = (((!g515) & (!g553) & (!g2692) & (g2693) & (g2751) & (!g2779)) + ((!g515) & (!g553) & (g2692) & (!g2693) & (!g2751) & (!g2779)) + ((!g515) & (!g553) & (g2692) & (!g2693) & (!g2751) & (g2779)) + ((!g515) & (!g553) & (g2692) & (!g2693) & (g2751) & (!g2779)) + ((!g515) & (!g553) & (g2692) & (!g2693) & (g2751) & (g2779)) + ((!g515) & (!g553) & (g2692) & (g2693) & (!g2751) & (!g2779)) + ((!g515) & (!g553) & (g2692) & (g2693) & (!g2751) & (g2779)) + ((!g515) & (!g553) & (g2692) & (g2693) & (g2751) & (g2779)) + ((!g515) & (g553) & (!g2692) & (!g2693) & (g2751) & (!g2779)) + ((!g515) & (g553) & (!g2692) & (g2693) & (!g2751) & (!g2779)) + ((!g515) & (g553) & (!g2692) & (g2693) & (g2751) & (!g2779)) + ((!g515) & (g553) & (g2692) & (!g2693) & (!g2751) & (!g2779)) + ((!g515) & (g553) & (g2692) & (!g2693) & (!g2751) & (g2779)) + ((!g515) & (g553) & (g2692) & (!g2693) & (g2751) & (g2779)) + ((!g515) & (g553) & (g2692) & (g2693) & (!g2751) & (g2779)) + ((!g515) & (g553) & (g2692) & (g2693) & (g2751) & (g2779)) + ((g515) & (!g553) & (!g2692) & (!g2693) & (!g2751) & (!g2779)) + ((g515) & (!g553) & (!g2692) & (!g2693) & (g2751) & (!g2779)) + ((g515) & (!g553) & (!g2692) & (g2693) & (!g2751) & (!g2779)) + ((g515) & (!g553) & (g2692) & (!g2693) & (!g2751) & (g2779)) + ((g515) & (!g553) & (g2692) & (!g2693) & (g2751) & (g2779)) + ((g515) & (!g553) & (g2692) & (g2693) & (!g2751) & (g2779)) + ((g515) & (!g553) & (g2692) & (g2693) & (g2751) & (!g2779)) + ((g515) & (!g553) & (g2692) & (g2693) & (g2751) & (g2779)) + ((g515) & (g553) & (!g2692) & (!g2693) & (!g2751) & (!g2779)) + ((g515) & (g553) & (g2692) & (!g2693) & (!g2751) & (g2779)) + ((g515) & (g553) & (g2692) & (!g2693) & (g2751) & (!g2779)) + ((g515) & (g553) & (g2692) & (!g2693) & (g2751) & (g2779)) + ((g515) & (g553) & (g2692) & (g2693) & (!g2751) & (!g2779)) + ((g515) & (g553) & (g2692) & (g2693) & (!g2751) & (g2779)) + ((g515) & (g553) & (g2692) & (g2693) & (g2751) & (!g2779)) + ((g515) & (g553) & (g2692) & (g2693) & (g2751) & (g2779)));
	assign g2796 = (((!g553) & (!g2693) & (g2751) & (!g2779)) + ((!g553) & (g2693) & (!g2751) & (!g2779)) + ((!g553) & (g2693) & (!g2751) & (g2779)) + ((!g553) & (g2693) & (g2751) & (g2779)) + ((g553) & (!g2693) & (!g2751) & (!g2779)) + ((g553) & (g2693) & (!g2751) & (g2779)) + ((g553) & (g2693) & (g2751) & (!g2779)) + ((g553) & (g2693) & (g2751) & (g2779)));
	assign g2797 = (((!g604) & (!g645) & (!g2695) & (g2696) & (g2750) & (!g2779)) + ((!g604) & (!g645) & (g2695) & (!g2696) & (!g2750) & (!g2779)) + ((!g604) & (!g645) & (g2695) & (!g2696) & (!g2750) & (g2779)) + ((!g604) & (!g645) & (g2695) & (!g2696) & (g2750) & (!g2779)) + ((!g604) & (!g645) & (g2695) & (!g2696) & (g2750) & (g2779)) + ((!g604) & (!g645) & (g2695) & (g2696) & (!g2750) & (!g2779)) + ((!g604) & (!g645) & (g2695) & (g2696) & (!g2750) & (g2779)) + ((!g604) & (!g645) & (g2695) & (g2696) & (g2750) & (g2779)) + ((!g604) & (g645) & (!g2695) & (!g2696) & (g2750) & (!g2779)) + ((!g604) & (g645) & (!g2695) & (g2696) & (!g2750) & (!g2779)) + ((!g604) & (g645) & (!g2695) & (g2696) & (g2750) & (!g2779)) + ((!g604) & (g645) & (g2695) & (!g2696) & (!g2750) & (!g2779)) + ((!g604) & (g645) & (g2695) & (!g2696) & (!g2750) & (g2779)) + ((!g604) & (g645) & (g2695) & (!g2696) & (g2750) & (g2779)) + ((!g604) & (g645) & (g2695) & (g2696) & (!g2750) & (g2779)) + ((!g604) & (g645) & (g2695) & (g2696) & (g2750) & (g2779)) + ((g604) & (!g645) & (!g2695) & (!g2696) & (!g2750) & (!g2779)) + ((g604) & (!g645) & (!g2695) & (!g2696) & (g2750) & (!g2779)) + ((g604) & (!g645) & (!g2695) & (g2696) & (!g2750) & (!g2779)) + ((g604) & (!g645) & (g2695) & (!g2696) & (!g2750) & (g2779)) + ((g604) & (!g645) & (g2695) & (!g2696) & (g2750) & (g2779)) + ((g604) & (!g645) & (g2695) & (g2696) & (!g2750) & (g2779)) + ((g604) & (!g645) & (g2695) & (g2696) & (g2750) & (!g2779)) + ((g604) & (!g645) & (g2695) & (g2696) & (g2750) & (g2779)) + ((g604) & (g645) & (!g2695) & (!g2696) & (!g2750) & (!g2779)) + ((g604) & (g645) & (g2695) & (!g2696) & (!g2750) & (g2779)) + ((g604) & (g645) & (g2695) & (!g2696) & (g2750) & (!g2779)) + ((g604) & (g645) & (g2695) & (!g2696) & (g2750) & (g2779)) + ((g604) & (g645) & (g2695) & (g2696) & (!g2750) & (!g2779)) + ((g604) & (g645) & (g2695) & (g2696) & (!g2750) & (g2779)) + ((g604) & (g645) & (g2695) & (g2696) & (g2750) & (!g2779)) + ((g604) & (g645) & (g2695) & (g2696) & (g2750) & (g2779)));
	assign g2798 = (((!g645) & (!g2696) & (g2750) & (!g2779)) + ((!g645) & (g2696) & (!g2750) & (!g2779)) + ((!g645) & (g2696) & (!g2750) & (g2779)) + ((!g645) & (g2696) & (g2750) & (g2779)) + ((g645) & (!g2696) & (!g2750) & (!g2779)) + ((g645) & (g2696) & (!g2750) & (g2779)) + ((g645) & (g2696) & (g2750) & (!g2779)) + ((g645) & (g2696) & (g2750) & (g2779)));
	assign g2799 = (((!g700) & (!g744) & (!g2698) & (g2699) & (g2749) & (!g2779)) + ((!g700) & (!g744) & (g2698) & (!g2699) & (!g2749) & (!g2779)) + ((!g700) & (!g744) & (g2698) & (!g2699) & (!g2749) & (g2779)) + ((!g700) & (!g744) & (g2698) & (!g2699) & (g2749) & (!g2779)) + ((!g700) & (!g744) & (g2698) & (!g2699) & (g2749) & (g2779)) + ((!g700) & (!g744) & (g2698) & (g2699) & (!g2749) & (!g2779)) + ((!g700) & (!g744) & (g2698) & (g2699) & (!g2749) & (g2779)) + ((!g700) & (!g744) & (g2698) & (g2699) & (g2749) & (g2779)) + ((!g700) & (g744) & (!g2698) & (!g2699) & (g2749) & (!g2779)) + ((!g700) & (g744) & (!g2698) & (g2699) & (!g2749) & (!g2779)) + ((!g700) & (g744) & (!g2698) & (g2699) & (g2749) & (!g2779)) + ((!g700) & (g744) & (g2698) & (!g2699) & (!g2749) & (!g2779)) + ((!g700) & (g744) & (g2698) & (!g2699) & (!g2749) & (g2779)) + ((!g700) & (g744) & (g2698) & (!g2699) & (g2749) & (g2779)) + ((!g700) & (g744) & (g2698) & (g2699) & (!g2749) & (g2779)) + ((!g700) & (g744) & (g2698) & (g2699) & (g2749) & (g2779)) + ((g700) & (!g744) & (!g2698) & (!g2699) & (!g2749) & (!g2779)) + ((g700) & (!g744) & (!g2698) & (!g2699) & (g2749) & (!g2779)) + ((g700) & (!g744) & (!g2698) & (g2699) & (!g2749) & (!g2779)) + ((g700) & (!g744) & (g2698) & (!g2699) & (!g2749) & (g2779)) + ((g700) & (!g744) & (g2698) & (!g2699) & (g2749) & (g2779)) + ((g700) & (!g744) & (g2698) & (g2699) & (!g2749) & (g2779)) + ((g700) & (!g744) & (g2698) & (g2699) & (g2749) & (!g2779)) + ((g700) & (!g744) & (g2698) & (g2699) & (g2749) & (g2779)) + ((g700) & (g744) & (!g2698) & (!g2699) & (!g2749) & (!g2779)) + ((g700) & (g744) & (g2698) & (!g2699) & (!g2749) & (g2779)) + ((g700) & (g744) & (g2698) & (!g2699) & (g2749) & (!g2779)) + ((g700) & (g744) & (g2698) & (!g2699) & (g2749) & (g2779)) + ((g700) & (g744) & (g2698) & (g2699) & (!g2749) & (!g2779)) + ((g700) & (g744) & (g2698) & (g2699) & (!g2749) & (g2779)) + ((g700) & (g744) & (g2698) & (g2699) & (g2749) & (!g2779)) + ((g700) & (g744) & (g2698) & (g2699) & (g2749) & (g2779)));
	assign g2800 = (((!g744) & (!g2699) & (g2749) & (!g2779)) + ((!g744) & (g2699) & (!g2749) & (!g2779)) + ((!g744) & (g2699) & (!g2749) & (g2779)) + ((!g744) & (g2699) & (g2749) & (g2779)) + ((g744) & (!g2699) & (!g2749) & (!g2779)) + ((g744) & (g2699) & (!g2749) & (g2779)) + ((g744) & (g2699) & (g2749) & (!g2779)) + ((g744) & (g2699) & (g2749) & (g2779)));
	assign g2801 = (((!g803) & (!g851) & (!g2701) & (g2702) & (g2748) & (!g2779)) + ((!g803) & (!g851) & (g2701) & (!g2702) & (!g2748) & (!g2779)) + ((!g803) & (!g851) & (g2701) & (!g2702) & (!g2748) & (g2779)) + ((!g803) & (!g851) & (g2701) & (!g2702) & (g2748) & (!g2779)) + ((!g803) & (!g851) & (g2701) & (!g2702) & (g2748) & (g2779)) + ((!g803) & (!g851) & (g2701) & (g2702) & (!g2748) & (!g2779)) + ((!g803) & (!g851) & (g2701) & (g2702) & (!g2748) & (g2779)) + ((!g803) & (!g851) & (g2701) & (g2702) & (g2748) & (g2779)) + ((!g803) & (g851) & (!g2701) & (!g2702) & (g2748) & (!g2779)) + ((!g803) & (g851) & (!g2701) & (g2702) & (!g2748) & (!g2779)) + ((!g803) & (g851) & (!g2701) & (g2702) & (g2748) & (!g2779)) + ((!g803) & (g851) & (g2701) & (!g2702) & (!g2748) & (!g2779)) + ((!g803) & (g851) & (g2701) & (!g2702) & (!g2748) & (g2779)) + ((!g803) & (g851) & (g2701) & (!g2702) & (g2748) & (g2779)) + ((!g803) & (g851) & (g2701) & (g2702) & (!g2748) & (g2779)) + ((!g803) & (g851) & (g2701) & (g2702) & (g2748) & (g2779)) + ((g803) & (!g851) & (!g2701) & (!g2702) & (!g2748) & (!g2779)) + ((g803) & (!g851) & (!g2701) & (!g2702) & (g2748) & (!g2779)) + ((g803) & (!g851) & (!g2701) & (g2702) & (!g2748) & (!g2779)) + ((g803) & (!g851) & (g2701) & (!g2702) & (!g2748) & (g2779)) + ((g803) & (!g851) & (g2701) & (!g2702) & (g2748) & (g2779)) + ((g803) & (!g851) & (g2701) & (g2702) & (!g2748) & (g2779)) + ((g803) & (!g851) & (g2701) & (g2702) & (g2748) & (!g2779)) + ((g803) & (!g851) & (g2701) & (g2702) & (g2748) & (g2779)) + ((g803) & (g851) & (!g2701) & (!g2702) & (!g2748) & (!g2779)) + ((g803) & (g851) & (g2701) & (!g2702) & (!g2748) & (g2779)) + ((g803) & (g851) & (g2701) & (!g2702) & (g2748) & (!g2779)) + ((g803) & (g851) & (g2701) & (!g2702) & (g2748) & (g2779)) + ((g803) & (g851) & (g2701) & (g2702) & (!g2748) & (!g2779)) + ((g803) & (g851) & (g2701) & (g2702) & (!g2748) & (g2779)) + ((g803) & (g851) & (g2701) & (g2702) & (g2748) & (!g2779)) + ((g803) & (g851) & (g2701) & (g2702) & (g2748) & (g2779)));
	assign g2802 = (((!g851) & (!g2702) & (g2748) & (!g2779)) + ((!g851) & (g2702) & (!g2748) & (!g2779)) + ((!g851) & (g2702) & (!g2748) & (g2779)) + ((!g851) & (g2702) & (g2748) & (g2779)) + ((g851) & (!g2702) & (!g2748) & (!g2779)) + ((g851) & (g2702) & (!g2748) & (g2779)) + ((g851) & (g2702) & (g2748) & (!g2779)) + ((g851) & (g2702) & (g2748) & (g2779)));
	assign g2803 = (((!g914) & (!g1032) & (!g2704) & (g2705) & (g2747) & (!g2779)) + ((!g914) & (!g1032) & (g2704) & (!g2705) & (!g2747) & (!g2779)) + ((!g914) & (!g1032) & (g2704) & (!g2705) & (!g2747) & (g2779)) + ((!g914) & (!g1032) & (g2704) & (!g2705) & (g2747) & (!g2779)) + ((!g914) & (!g1032) & (g2704) & (!g2705) & (g2747) & (g2779)) + ((!g914) & (!g1032) & (g2704) & (g2705) & (!g2747) & (!g2779)) + ((!g914) & (!g1032) & (g2704) & (g2705) & (!g2747) & (g2779)) + ((!g914) & (!g1032) & (g2704) & (g2705) & (g2747) & (g2779)) + ((!g914) & (g1032) & (!g2704) & (!g2705) & (g2747) & (!g2779)) + ((!g914) & (g1032) & (!g2704) & (g2705) & (!g2747) & (!g2779)) + ((!g914) & (g1032) & (!g2704) & (g2705) & (g2747) & (!g2779)) + ((!g914) & (g1032) & (g2704) & (!g2705) & (!g2747) & (!g2779)) + ((!g914) & (g1032) & (g2704) & (!g2705) & (!g2747) & (g2779)) + ((!g914) & (g1032) & (g2704) & (!g2705) & (g2747) & (g2779)) + ((!g914) & (g1032) & (g2704) & (g2705) & (!g2747) & (g2779)) + ((!g914) & (g1032) & (g2704) & (g2705) & (g2747) & (g2779)) + ((g914) & (!g1032) & (!g2704) & (!g2705) & (!g2747) & (!g2779)) + ((g914) & (!g1032) & (!g2704) & (!g2705) & (g2747) & (!g2779)) + ((g914) & (!g1032) & (!g2704) & (g2705) & (!g2747) & (!g2779)) + ((g914) & (!g1032) & (g2704) & (!g2705) & (!g2747) & (g2779)) + ((g914) & (!g1032) & (g2704) & (!g2705) & (g2747) & (g2779)) + ((g914) & (!g1032) & (g2704) & (g2705) & (!g2747) & (g2779)) + ((g914) & (!g1032) & (g2704) & (g2705) & (g2747) & (!g2779)) + ((g914) & (!g1032) & (g2704) & (g2705) & (g2747) & (g2779)) + ((g914) & (g1032) & (!g2704) & (!g2705) & (!g2747) & (!g2779)) + ((g914) & (g1032) & (g2704) & (!g2705) & (!g2747) & (g2779)) + ((g914) & (g1032) & (g2704) & (!g2705) & (g2747) & (!g2779)) + ((g914) & (g1032) & (g2704) & (!g2705) & (g2747) & (g2779)) + ((g914) & (g1032) & (g2704) & (g2705) & (!g2747) & (!g2779)) + ((g914) & (g1032) & (g2704) & (g2705) & (!g2747) & (g2779)) + ((g914) & (g1032) & (g2704) & (g2705) & (g2747) & (!g2779)) + ((g914) & (g1032) & (g2704) & (g2705) & (g2747) & (g2779)));
	assign g2804 = (((!g1032) & (!g2705) & (g2747) & (!g2779)) + ((!g1032) & (g2705) & (!g2747) & (!g2779)) + ((!g1032) & (g2705) & (!g2747) & (g2779)) + ((!g1032) & (g2705) & (g2747) & (g2779)) + ((g1032) & (!g2705) & (!g2747) & (!g2779)) + ((g1032) & (g2705) & (!g2747) & (g2779)) + ((g1032) & (g2705) & (g2747) & (!g2779)) + ((g1032) & (g2705) & (g2747) & (g2779)));
	assign g2805 = (((!g1030) & (!g1160) & (!g2707) & (g2708) & (g2746) & (!g2779)) + ((!g1030) & (!g1160) & (g2707) & (!g2708) & (!g2746) & (!g2779)) + ((!g1030) & (!g1160) & (g2707) & (!g2708) & (!g2746) & (g2779)) + ((!g1030) & (!g1160) & (g2707) & (!g2708) & (g2746) & (!g2779)) + ((!g1030) & (!g1160) & (g2707) & (!g2708) & (g2746) & (g2779)) + ((!g1030) & (!g1160) & (g2707) & (g2708) & (!g2746) & (!g2779)) + ((!g1030) & (!g1160) & (g2707) & (g2708) & (!g2746) & (g2779)) + ((!g1030) & (!g1160) & (g2707) & (g2708) & (g2746) & (g2779)) + ((!g1030) & (g1160) & (!g2707) & (!g2708) & (g2746) & (!g2779)) + ((!g1030) & (g1160) & (!g2707) & (g2708) & (!g2746) & (!g2779)) + ((!g1030) & (g1160) & (!g2707) & (g2708) & (g2746) & (!g2779)) + ((!g1030) & (g1160) & (g2707) & (!g2708) & (!g2746) & (!g2779)) + ((!g1030) & (g1160) & (g2707) & (!g2708) & (!g2746) & (g2779)) + ((!g1030) & (g1160) & (g2707) & (!g2708) & (g2746) & (g2779)) + ((!g1030) & (g1160) & (g2707) & (g2708) & (!g2746) & (g2779)) + ((!g1030) & (g1160) & (g2707) & (g2708) & (g2746) & (g2779)) + ((g1030) & (!g1160) & (!g2707) & (!g2708) & (!g2746) & (!g2779)) + ((g1030) & (!g1160) & (!g2707) & (!g2708) & (g2746) & (!g2779)) + ((g1030) & (!g1160) & (!g2707) & (g2708) & (!g2746) & (!g2779)) + ((g1030) & (!g1160) & (g2707) & (!g2708) & (!g2746) & (g2779)) + ((g1030) & (!g1160) & (g2707) & (!g2708) & (g2746) & (g2779)) + ((g1030) & (!g1160) & (g2707) & (g2708) & (!g2746) & (g2779)) + ((g1030) & (!g1160) & (g2707) & (g2708) & (g2746) & (!g2779)) + ((g1030) & (!g1160) & (g2707) & (g2708) & (g2746) & (g2779)) + ((g1030) & (g1160) & (!g2707) & (!g2708) & (!g2746) & (!g2779)) + ((g1030) & (g1160) & (g2707) & (!g2708) & (!g2746) & (g2779)) + ((g1030) & (g1160) & (g2707) & (!g2708) & (g2746) & (!g2779)) + ((g1030) & (g1160) & (g2707) & (!g2708) & (g2746) & (g2779)) + ((g1030) & (g1160) & (g2707) & (g2708) & (!g2746) & (!g2779)) + ((g1030) & (g1160) & (g2707) & (g2708) & (!g2746) & (g2779)) + ((g1030) & (g1160) & (g2707) & (g2708) & (g2746) & (!g2779)) + ((g1030) & (g1160) & (g2707) & (g2708) & (g2746) & (g2779)));
	assign g2806 = (((!g1160) & (!g2708) & (g2746) & (!g2779)) + ((!g1160) & (g2708) & (!g2746) & (!g2779)) + ((!g1160) & (g2708) & (!g2746) & (g2779)) + ((!g1160) & (g2708) & (g2746) & (g2779)) + ((g1160) & (!g2708) & (!g2746) & (!g2779)) + ((g1160) & (g2708) & (!g2746) & (g2779)) + ((g1160) & (g2708) & (g2746) & (!g2779)) + ((g1160) & (g2708) & (g2746) & (g2779)));
	assign g2807 = (((!g1154) & (!g1295) & (!g2710) & (g2711) & (g2745) & (!g2779)) + ((!g1154) & (!g1295) & (g2710) & (!g2711) & (!g2745) & (!g2779)) + ((!g1154) & (!g1295) & (g2710) & (!g2711) & (!g2745) & (g2779)) + ((!g1154) & (!g1295) & (g2710) & (!g2711) & (g2745) & (!g2779)) + ((!g1154) & (!g1295) & (g2710) & (!g2711) & (g2745) & (g2779)) + ((!g1154) & (!g1295) & (g2710) & (g2711) & (!g2745) & (!g2779)) + ((!g1154) & (!g1295) & (g2710) & (g2711) & (!g2745) & (g2779)) + ((!g1154) & (!g1295) & (g2710) & (g2711) & (g2745) & (g2779)) + ((!g1154) & (g1295) & (!g2710) & (!g2711) & (g2745) & (!g2779)) + ((!g1154) & (g1295) & (!g2710) & (g2711) & (!g2745) & (!g2779)) + ((!g1154) & (g1295) & (!g2710) & (g2711) & (g2745) & (!g2779)) + ((!g1154) & (g1295) & (g2710) & (!g2711) & (!g2745) & (!g2779)) + ((!g1154) & (g1295) & (g2710) & (!g2711) & (!g2745) & (g2779)) + ((!g1154) & (g1295) & (g2710) & (!g2711) & (g2745) & (g2779)) + ((!g1154) & (g1295) & (g2710) & (g2711) & (!g2745) & (g2779)) + ((!g1154) & (g1295) & (g2710) & (g2711) & (g2745) & (g2779)) + ((g1154) & (!g1295) & (!g2710) & (!g2711) & (!g2745) & (!g2779)) + ((g1154) & (!g1295) & (!g2710) & (!g2711) & (g2745) & (!g2779)) + ((g1154) & (!g1295) & (!g2710) & (g2711) & (!g2745) & (!g2779)) + ((g1154) & (!g1295) & (g2710) & (!g2711) & (!g2745) & (g2779)) + ((g1154) & (!g1295) & (g2710) & (!g2711) & (g2745) & (g2779)) + ((g1154) & (!g1295) & (g2710) & (g2711) & (!g2745) & (g2779)) + ((g1154) & (!g1295) & (g2710) & (g2711) & (g2745) & (!g2779)) + ((g1154) & (!g1295) & (g2710) & (g2711) & (g2745) & (g2779)) + ((g1154) & (g1295) & (!g2710) & (!g2711) & (!g2745) & (!g2779)) + ((g1154) & (g1295) & (g2710) & (!g2711) & (!g2745) & (g2779)) + ((g1154) & (g1295) & (g2710) & (!g2711) & (g2745) & (!g2779)) + ((g1154) & (g1295) & (g2710) & (!g2711) & (g2745) & (g2779)) + ((g1154) & (g1295) & (g2710) & (g2711) & (!g2745) & (!g2779)) + ((g1154) & (g1295) & (g2710) & (g2711) & (!g2745) & (g2779)) + ((g1154) & (g1295) & (g2710) & (g2711) & (g2745) & (!g2779)) + ((g1154) & (g1295) & (g2710) & (g2711) & (g2745) & (g2779)));
	assign g2808 = (((!g1295) & (!g2711) & (g2745) & (!g2779)) + ((!g1295) & (g2711) & (!g2745) & (!g2779)) + ((!g1295) & (g2711) & (!g2745) & (g2779)) + ((!g1295) & (g2711) & (g2745) & (g2779)) + ((g1295) & (!g2711) & (!g2745) & (!g2779)) + ((g1295) & (g2711) & (!g2745) & (g2779)) + ((g1295) & (g2711) & (g2745) & (!g2779)) + ((g1295) & (g2711) & (g2745) & (g2779)));
	assign g2809 = (((!g1285) & (!g1437) & (!g2713) & (g2714) & (g2744) & (!g2779)) + ((!g1285) & (!g1437) & (g2713) & (!g2714) & (!g2744) & (!g2779)) + ((!g1285) & (!g1437) & (g2713) & (!g2714) & (!g2744) & (g2779)) + ((!g1285) & (!g1437) & (g2713) & (!g2714) & (g2744) & (!g2779)) + ((!g1285) & (!g1437) & (g2713) & (!g2714) & (g2744) & (g2779)) + ((!g1285) & (!g1437) & (g2713) & (g2714) & (!g2744) & (!g2779)) + ((!g1285) & (!g1437) & (g2713) & (g2714) & (!g2744) & (g2779)) + ((!g1285) & (!g1437) & (g2713) & (g2714) & (g2744) & (g2779)) + ((!g1285) & (g1437) & (!g2713) & (!g2714) & (g2744) & (!g2779)) + ((!g1285) & (g1437) & (!g2713) & (g2714) & (!g2744) & (!g2779)) + ((!g1285) & (g1437) & (!g2713) & (g2714) & (g2744) & (!g2779)) + ((!g1285) & (g1437) & (g2713) & (!g2714) & (!g2744) & (!g2779)) + ((!g1285) & (g1437) & (g2713) & (!g2714) & (!g2744) & (g2779)) + ((!g1285) & (g1437) & (g2713) & (!g2714) & (g2744) & (g2779)) + ((!g1285) & (g1437) & (g2713) & (g2714) & (!g2744) & (g2779)) + ((!g1285) & (g1437) & (g2713) & (g2714) & (g2744) & (g2779)) + ((g1285) & (!g1437) & (!g2713) & (!g2714) & (!g2744) & (!g2779)) + ((g1285) & (!g1437) & (!g2713) & (!g2714) & (g2744) & (!g2779)) + ((g1285) & (!g1437) & (!g2713) & (g2714) & (!g2744) & (!g2779)) + ((g1285) & (!g1437) & (g2713) & (!g2714) & (!g2744) & (g2779)) + ((g1285) & (!g1437) & (g2713) & (!g2714) & (g2744) & (g2779)) + ((g1285) & (!g1437) & (g2713) & (g2714) & (!g2744) & (g2779)) + ((g1285) & (!g1437) & (g2713) & (g2714) & (g2744) & (!g2779)) + ((g1285) & (!g1437) & (g2713) & (g2714) & (g2744) & (g2779)) + ((g1285) & (g1437) & (!g2713) & (!g2714) & (!g2744) & (!g2779)) + ((g1285) & (g1437) & (g2713) & (!g2714) & (!g2744) & (g2779)) + ((g1285) & (g1437) & (g2713) & (!g2714) & (g2744) & (!g2779)) + ((g1285) & (g1437) & (g2713) & (!g2714) & (g2744) & (g2779)) + ((g1285) & (g1437) & (g2713) & (g2714) & (!g2744) & (!g2779)) + ((g1285) & (g1437) & (g2713) & (g2714) & (!g2744) & (g2779)) + ((g1285) & (g1437) & (g2713) & (g2714) & (g2744) & (!g2779)) + ((g1285) & (g1437) & (g2713) & (g2714) & (g2744) & (g2779)));
	assign g2810 = (((!g1437) & (!g2714) & (g2744) & (!g2779)) + ((!g1437) & (g2714) & (!g2744) & (!g2779)) + ((!g1437) & (g2714) & (!g2744) & (g2779)) + ((!g1437) & (g2714) & (g2744) & (g2779)) + ((g1437) & (!g2714) & (!g2744) & (!g2779)) + ((g1437) & (g2714) & (!g2744) & (g2779)) + ((g1437) & (g2714) & (g2744) & (!g2779)) + ((g1437) & (g2714) & (g2744) & (g2779)));
	assign g2811 = (((!g1423) & (!g1586) & (!g2716) & (g2717) & (g2743) & (!g2779)) + ((!g1423) & (!g1586) & (g2716) & (!g2717) & (!g2743) & (!g2779)) + ((!g1423) & (!g1586) & (g2716) & (!g2717) & (!g2743) & (g2779)) + ((!g1423) & (!g1586) & (g2716) & (!g2717) & (g2743) & (!g2779)) + ((!g1423) & (!g1586) & (g2716) & (!g2717) & (g2743) & (g2779)) + ((!g1423) & (!g1586) & (g2716) & (g2717) & (!g2743) & (!g2779)) + ((!g1423) & (!g1586) & (g2716) & (g2717) & (!g2743) & (g2779)) + ((!g1423) & (!g1586) & (g2716) & (g2717) & (g2743) & (g2779)) + ((!g1423) & (g1586) & (!g2716) & (!g2717) & (g2743) & (!g2779)) + ((!g1423) & (g1586) & (!g2716) & (g2717) & (!g2743) & (!g2779)) + ((!g1423) & (g1586) & (!g2716) & (g2717) & (g2743) & (!g2779)) + ((!g1423) & (g1586) & (g2716) & (!g2717) & (!g2743) & (!g2779)) + ((!g1423) & (g1586) & (g2716) & (!g2717) & (!g2743) & (g2779)) + ((!g1423) & (g1586) & (g2716) & (!g2717) & (g2743) & (g2779)) + ((!g1423) & (g1586) & (g2716) & (g2717) & (!g2743) & (g2779)) + ((!g1423) & (g1586) & (g2716) & (g2717) & (g2743) & (g2779)) + ((g1423) & (!g1586) & (!g2716) & (!g2717) & (!g2743) & (!g2779)) + ((g1423) & (!g1586) & (!g2716) & (!g2717) & (g2743) & (!g2779)) + ((g1423) & (!g1586) & (!g2716) & (g2717) & (!g2743) & (!g2779)) + ((g1423) & (!g1586) & (g2716) & (!g2717) & (!g2743) & (g2779)) + ((g1423) & (!g1586) & (g2716) & (!g2717) & (g2743) & (g2779)) + ((g1423) & (!g1586) & (g2716) & (g2717) & (!g2743) & (g2779)) + ((g1423) & (!g1586) & (g2716) & (g2717) & (g2743) & (!g2779)) + ((g1423) & (!g1586) & (g2716) & (g2717) & (g2743) & (g2779)) + ((g1423) & (g1586) & (!g2716) & (!g2717) & (!g2743) & (!g2779)) + ((g1423) & (g1586) & (g2716) & (!g2717) & (!g2743) & (g2779)) + ((g1423) & (g1586) & (g2716) & (!g2717) & (g2743) & (!g2779)) + ((g1423) & (g1586) & (g2716) & (!g2717) & (g2743) & (g2779)) + ((g1423) & (g1586) & (g2716) & (g2717) & (!g2743) & (!g2779)) + ((g1423) & (g1586) & (g2716) & (g2717) & (!g2743) & (g2779)) + ((g1423) & (g1586) & (g2716) & (g2717) & (g2743) & (!g2779)) + ((g1423) & (g1586) & (g2716) & (g2717) & (g2743) & (g2779)));
	assign g2812 = (((!g1586) & (!g2717) & (g2743) & (!g2779)) + ((!g1586) & (g2717) & (!g2743) & (!g2779)) + ((!g1586) & (g2717) & (!g2743) & (g2779)) + ((!g1586) & (g2717) & (g2743) & (g2779)) + ((g1586) & (!g2717) & (!g2743) & (!g2779)) + ((g1586) & (g2717) & (!g2743) & (g2779)) + ((g1586) & (g2717) & (g2743) & (!g2779)) + ((g1586) & (g2717) & (g2743) & (g2779)));
	assign g2813 = (((!g1568) & (!g1742) & (!g2719) & (g2720) & (g2742) & (!g2779)) + ((!g1568) & (!g1742) & (g2719) & (!g2720) & (!g2742) & (!g2779)) + ((!g1568) & (!g1742) & (g2719) & (!g2720) & (!g2742) & (g2779)) + ((!g1568) & (!g1742) & (g2719) & (!g2720) & (g2742) & (!g2779)) + ((!g1568) & (!g1742) & (g2719) & (!g2720) & (g2742) & (g2779)) + ((!g1568) & (!g1742) & (g2719) & (g2720) & (!g2742) & (!g2779)) + ((!g1568) & (!g1742) & (g2719) & (g2720) & (!g2742) & (g2779)) + ((!g1568) & (!g1742) & (g2719) & (g2720) & (g2742) & (g2779)) + ((!g1568) & (g1742) & (!g2719) & (!g2720) & (g2742) & (!g2779)) + ((!g1568) & (g1742) & (!g2719) & (g2720) & (!g2742) & (!g2779)) + ((!g1568) & (g1742) & (!g2719) & (g2720) & (g2742) & (!g2779)) + ((!g1568) & (g1742) & (g2719) & (!g2720) & (!g2742) & (!g2779)) + ((!g1568) & (g1742) & (g2719) & (!g2720) & (!g2742) & (g2779)) + ((!g1568) & (g1742) & (g2719) & (!g2720) & (g2742) & (g2779)) + ((!g1568) & (g1742) & (g2719) & (g2720) & (!g2742) & (g2779)) + ((!g1568) & (g1742) & (g2719) & (g2720) & (g2742) & (g2779)) + ((g1568) & (!g1742) & (!g2719) & (!g2720) & (!g2742) & (!g2779)) + ((g1568) & (!g1742) & (!g2719) & (!g2720) & (g2742) & (!g2779)) + ((g1568) & (!g1742) & (!g2719) & (g2720) & (!g2742) & (!g2779)) + ((g1568) & (!g1742) & (g2719) & (!g2720) & (!g2742) & (g2779)) + ((g1568) & (!g1742) & (g2719) & (!g2720) & (g2742) & (g2779)) + ((g1568) & (!g1742) & (g2719) & (g2720) & (!g2742) & (g2779)) + ((g1568) & (!g1742) & (g2719) & (g2720) & (g2742) & (!g2779)) + ((g1568) & (!g1742) & (g2719) & (g2720) & (g2742) & (g2779)) + ((g1568) & (g1742) & (!g2719) & (!g2720) & (!g2742) & (!g2779)) + ((g1568) & (g1742) & (g2719) & (!g2720) & (!g2742) & (g2779)) + ((g1568) & (g1742) & (g2719) & (!g2720) & (g2742) & (!g2779)) + ((g1568) & (g1742) & (g2719) & (!g2720) & (g2742) & (g2779)) + ((g1568) & (g1742) & (g2719) & (g2720) & (!g2742) & (!g2779)) + ((g1568) & (g1742) & (g2719) & (g2720) & (!g2742) & (g2779)) + ((g1568) & (g1742) & (g2719) & (g2720) & (g2742) & (!g2779)) + ((g1568) & (g1742) & (g2719) & (g2720) & (g2742) & (g2779)));
	assign g2814 = (((!g1742) & (!g2720) & (g2742) & (!g2779)) + ((!g1742) & (g2720) & (!g2742) & (!g2779)) + ((!g1742) & (g2720) & (!g2742) & (g2779)) + ((!g1742) & (g2720) & (g2742) & (g2779)) + ((g1742) & (!g2720) & (!g2742) & (!g2779)) + ((g1742) & (g2720) & (!g2742) & (g2779)) + ((g1742) & (g2720) & (g2742) & (!g2779)) + ((g1742) & (g2720) & (g2742) & (g2779)));
	assign g2815 = (((!g1720) & (!g1905) & (!g2722) & (g2723) & (g2741) & (!g2779)) + ((!g1720) & (!g1905) & (g2722) & (!g2723) & (!g2741) & (!g2779)) + ((!g1720) & (!g1905) & (g2722) & (!g2723) & (!g2741) & (g2779)) + ((!g1720) & (!g1905) & (g2722) & (!g2723) & (g2741) & (!g2779)) + ((!g1720) & (!g1905) & (g2722) & (!g2723) & (g2741) & (g2779)) + ((!g1720) & (!g1905) & (g2722) & (g2723) & (!g2741) & (!g2779)) + ((!g1720) & (!g1905) & (g2722) & (g2723) & (!g2741) & (g2779)) + ((!g1720) & (!g1905) & (g2722) & (g2723) & (g2741) & (g2779)) + ((!g1720) & (g1905) & (!g2722) & (!g2723) & (g2741) & (!g2779)) + ((!g1720) & (g1905) & (!g2722) & (g2723) & (!g2741) & (!g2779)) + ((!g1720) & (g1905) & (!g2722) & (g2723) & (g2741) & (!g2779)) + ((!g1720) & (g1905) & (g2722) & (!g2723) & (!g2741) & (!g2779)) + ((!g1720) & (g1905) & (g2722) & (!g2723) & (!g2741) & (g2779)) + ((!g1720) & (g1905) & (g2722) & (!g2723) & (g2741) & (g2779)) + ((!g1720) & (g1905) & (g2722) & (g2723) & (!g2741) & (g2779)) + ((!g1720) & (g1905) & (g2722) & (g2723) & (g2741) & (g2779)) + ((g1720) & (!g1905) & (!g2722) & (!g2723) & (!g2741) & (!g2779)) + ((g1720) & (!g1905) & (!g2722) & (!g2723) & (g2741) & (!g2779)) + ((g1720) & (!g1905) & (!g2722) & (g2723) & (!g2741) & (!g2779)) + ((g1720) & (!g1905) & (g2722) & (!g2723) & (!g2741) & (g2779)) + ((g1720) & (!g1905) & (g2722) & (!g2723) & (g2741) & (g2779)) + ((g1720) & (!g1905) & (g2722) & (g2723) & (!g2741) & (g2779)) + ((g1720) & (!g1905) & (g2722) & (g2723) & (g2741) & (!g2779)) + ((g1720) & (!g1905) & (g2722) & (g2723) & (g2741) & (g2779)) + ((g1720) & (g1905) & (!g2722) & (!g2723) & (!g2741) & (!g2779)) + ((g1720) & (g1905) & (g2722) & (!g2723) & (!g2741) & (g2779)) + ((g1720) & (g1905) & (g2722) & (!g2723) & (g2741) & (!g2779)) + ((g1720) & (g1905) & (g2722) & (!g2723) & (g2741) & (g2779)) + ((g1720) & (g1905) & (g2722) & (g2723) & (!g2741) & (!g2779)) + ((g1720) & (g1905) & (g2722) & (g2723) & (!g2741) & (g2779)) + ((g1720) & (g1905) & (g2722) & (g2723) & (g2741) & (!g2779)) + ((g1720) & (g1905) & (g2722) & (g2723) & (g2741) & (g2779)));
	assign g2816 = (((!g1905) & (!g2723) & (g2741) & (!g2779)) + ((!g1905) & (g2723) & (!g2741) & (!g2779)) + ((!g1905) & (g2723) & (!g2741) & (g2779)) + ((!g1905) & (g2723) & (g2741) & (g2779)) + ((g1905) & (!g2723) & (!g2741) & (!g2779)) + ((g1905) & (g2723) & (!g2741) & (g2779)) + ((g1905) & (g2723) & (g2741) & (!g2779)) + ((g1905) & (g2723) & (g2741) & (g2779)));
	assign g2817 = (((!g1879) & (!g2075) & (!g2725) & (g2726) & (g2740) & (!g2779)) + ((!g1879) & (!g2075) & (g2725) & (!g2726) & (!g2740) & (!g2779)) + ((!g1879) & (!g2075) & (g2725) & (!g2726) & (!g2740) & (g2779)) + ((!g1879) & (!g2075) & (g2725) & (!g2726) & (g2740) & (!g2779)) + ((!g1879) & (!g2075) & (g2725) & (!g2726) & (g2740) & (g2779)) + ((!g1879) & (!g2075) & (g2725) & (g2726) & (!g2740) & (!g2779)) + ((!g1879) & (!g2075) & (g2725) & (g2726) & (!g2740) & (g2779)) + ((!g1879) & (!g2075) & (g2725) & (g2726) & (g2740) & (g2779)) + ((!g1879) & (g2075) & (!g2725) & (!g2726) & (g2740) & (!g2779)) + ((!g1879) & (g2075) & (!g2725) & (g2726) & (!g2740) & (!g2779)) + ((!g1879) & (g2075) & (!g2725) & (g2726) & (g2740) & (!g2779)) + ((!g1879) & (g2075) & (g2725) & (!g2726) & (!g2740) & (!g2779)) + ((!g1879) & (g2075) & (g2725) & (!g2726) & (!g2740) & (g2779)) + ((!g1879) & (g2075) & (g2725) & (!g2726) & (g2740) & (g2779)) + ((!g1879) & (g2075) & (g2725) & (g2726) & (!g2740) & (g2779)) + ((!g1879) & (g2075) & (g2725) & (g2726) & (g2740) & (g2779)) + ((g1879) & (!g2075) & (!g2725) & (!g2726) & (!g2740) & (!g2779)) + ((g1879) & (!g2075) & (!g2725) & (!g2726) & (g2740) & (!g2779)) + ((g1879) & (!g2075) & (!g2725) & (g2726) & (!g2740) & (!g2779)) + ((g1879) & (!g2075) & (g2725) & (!g2726) & (!g2740) & (g2779)) + ((g1879) & (!g2075) & (g2725) & (!g2726) & (g2740) & (g2779)) + ((g1879) & (!g2075) & (g2725) & (g2726) & (!g2740) & (g2779)) + ((g1879) & (!g2075) & (g2725) & (g2726) & (g2740) & (!g2779)) + ((g1879) & (!g2075) & (g2725) & (g2726) & (g2740) & (g2779)) + ((g1879) & (g2075) & (!g2725) & (!g2726) & (!g2740) & (!g2779)) + ((g1879) & (g2075) & (g2725) & (!g2726) & (!g2740) & (g2779)) + ((g1879) & (g2075) & (g2725) & (!g2726) & (g2740) & (!g2779)) + ((g1879) & (g2075) & (g2725) & (!g2726) & (g2740) & (g2779)) + ((g1879) & (g2075) & (g2725) & (g2726) & (!g2740) & (!g2779)) + ((g1879) & (g2075) & (g2725) & (g2726) & (!g2740) & (g2779)) + ((g1879) & (g2075) & (g2725) & (g2726) & (g2740) & (!g2779)) + ((g1879) & (g2075) & (g2725) & (g2726) & (g2740) & (g2779)));
	assign g2818 = (((!g2075) & (!g2726) & (g2740) & (!g2779)) + ((!g2075) & (g2726) & (!g2740) & (!g2779)) + ((!g2075) & (g2726) & (!g2740) & (g2779)) + ((!g2075) & (g2726) & (g2740) & (g2779)) + ((g2075) & (!g2726) & (!g2740) & (!g2779)) + ((g2075) & (g2726) & (!g2740) & (g2779)) + ((g2075) & (g2726) & (g2740) & (!g2779)) + ((g2075) & (g2726) & (g2740) & (g2779)));
	assign g2819 = (((!g2045) & (!g2252) & (!g2728) & (g2729) & (g2739) & (!g2779)) + ((!g2045) & (!g2252) & (g2728) & (!g2729) & (!g2739) & (!g2779)) + ((!g2045) & (!g2252) & (g2728) & (!g2729) & (!g2739) & (g2779)) + ((!g2045) & (!g2252) & (g2728) & (!g2729) & (g2739) & (!g2779)) + ((!g2045) & (!g2252) & (g2728) & (!g2729) & (g2739) & (g2779)) + ((!g2045) & (!g2252) & (g2728) & (g2729) & (!g2739) & (!g2779)) + ((!g2045) & (!g2252) & (g2728) & (g2729) & (!g2739) & (g2779)) + ((!g2045) & (!g2252) & (g2728) & (g2729) & (g2739) & (g2779)) + ((!g2045) & (g2252) & (!g2728) & (!g2729) & (g2739) & (!g2779)) + ((!g2045) & (g2252) & (!g2728) & (g2729) & (!g2739) & (!g2779)) + ((!g2045) & (g2252) & (!g2728) & (g2729) & (g2739) & (!g2779)) + ((!g2045) & (g2252) & (g2728) & (!g2729) & (!g2739) & (!g2779)) + ((!g2045) & (g2252) & (g2728) & (!g2729) & (!g2739) & (g2779)) + ((!g2045) & (g2252) & (g2728) & (!g2729) & (g2739) & (g2779)) + ((!g2045) & (g2252) & (g2728) & (g2729) & (!g2739) & (g2779)) + ((!g2045) & (g2252) & (g2728) & (g2729) & (g2739) & (g2779)) + ((g2045) & (!g2252) & (!g2728) & (!g2729) & (!g2739) & (!g2779)) + ((g2045) & (!g2252) & (!g2728) & (!g2729) & (g2739) & (!g2779)) + ((g2045) & (!g2252) & (!g2728) & (g2729) & (!g2739) & (!g2779)) + ((g2045) & (!g2252) & (g2728) & (!g2729) & (!g2739) & (g2779)) + ((g2045) & (!g2252) & (g2728) & (!g2729) & (g2739) & (g2779)) + ((g2045) & (!g2252) & (g2728) & (g2729) & (!g2739) & (g2779)) + ((g2045) & (!g2252) & (g2728) & (g2729) & (g2739) & (!g2779)) + ((g2045) & (!g2252) & (g2728) & (g2729) & (g2739) & (g2779)) + ((g2045) & (g2252) & (!g2728) & (!g2729) & (!g2739) & (!g2779)) + ((g2045) & (g2252) & (g2728) & (!g2729) & (!g2739) & (g2779)) + ((g2045) & (g2252) & (g2728) & (!g2729) & (g2739) & (!g2779)) + ((g2045) & (g2252) & (g2728) & (!g2729) & (g2739) & (g2779)) + ((g2045) & (g2252) & (g2728) & (g2729) & (!g2739) & (!g2779)) + ((g2045) & (g2252) & (g2728) & (g2729) & (!g2739) & (g2779)) + ((g2045) & (g2252) & (g2728) & (g2729) & (g2739) & (!g2779)) + ((g2045) & (g2252) & (g2728) & (g2729) & (g2739) & (g2779)));
	assign g2820 = (((!g2252) & (!g2729) & (g2739) & (!g2779)) + ((!g2252) & (g2729) & (!g2739) & (!g2779)) + ((!g2252) & (g2729) & (!g2739) & (g2779)) + ((!g2252) & (g2729) & (g2739) & (g2779)) + ((g2252) & (!g2729) & (!g2739) & (!g2779)) + ((g2252) & (g2729) & (!g2739) & (g2779)) + ((g2252) & (g2729) & (g2739) & (!g2779)) + ((g2252) & (g2729) & (g2739) & (g2779)));
	assign g2821 = (((!g2218) & (!g2436) & (!g2731) & (g2732) & (g2738) & (!g2779)) + ((!g2218) & (!g2436) & (g2731) & (!g2732) & (!g2738) & (!g2779)) + ((!g2218) & (!g2436) & (g2731) & (!g2732) & (!g2738) & (g2779)) + ((!g2218) & (!g2436) & (g2731) & (!g2732) & (g2738) & (!g2779)) + ((!g2218) & (!g2436) & (g2731) & (!g2732) & (g2738) & (g2779)) + ((!g2218) & (!g2436) & (g2731) & (g2732) & (!g2738) & (!g2779)) + ((!g2218) & (!g2436) & (g2731) & (g2732) & (!g2738) & (g2779)) + ((!g2218) & (!g2436) & (g2731) & (g2732) & (g2738) & (g2779)) + ((!g2218) & (g2436) & (!g2731) & (!g2732) & (g2738) & (!g2779)) + ((!g2218) & (g2436) & (!g2731) & (g2732) & (!g2738) & (!g2779)) + ((!g2218) & (g2436) & (!g2731) & (g2732) & (g2738) & (!g2779)) + ((!g2218) & (g2436) & (g2731) & (!g2732) & (!g2738) & (!g2779)) + ((!g2218) & (g2436) & (g2731) & (!g2732) & (!g2738) & (g2779)) + ((!g2218) & (g2436) & (g2731) & (!g2732) & (g2738) & (g2779)) + ((!g2218) & (g2436) & (g2731) & (g2732) & (!g2738) & (g2779)) + ((!g2218) & (g2436) & (g2731) & (g2732) & (g2738) & (g2779)) + ((g2218) & (!g2436) & (!g2731) & (!g2732) & (!g2738) & (!g2779)) + ((g2218) & (!g2436) & (!g2731) & (!g2732) & (g2738) & (!g2779)) + ((g2218) & (!g2436) & (!g2731) & (g2732) & (!g2738) & (!g2779)) + ((g2218) & (!g2436) & (g2731) & (!g2732) & (!g2738) & (g2779)) + ((g2218) & (!g2436) & (g2731) & (!g2732) & (g2738) & (g2779)) + ((g2218) & (!g2436) & (g2731) & (g2732) & (!g2738) & (g2779)) + ((g2218) & (!g2436) & (g2731) & (g2732) & (g2738) & (!g2779)) + ((g2218) & (!g2436) & (g2731) & (g2732) & (g2738) & (g2779)) + ((g2218) & (g2436) & (!g2731) & (!g2732) & (!g2738) & (!g2779)) + ((g2218) & (g2436) & (g2731) & (!g2732) & (!g2738) & (g2779)) + ((g2218) & (g2436) & (g2731) & (!g2732) & (g2738) & (!g2779)) + ((g2218) & (g2436) & (g2731) & (!g2732) & (g2738) & (g2779)) + ((g2218) & (g2436) & (g2731) & (g2732) & (!g2738) & (!g2779)) + ((g2218) & (g2436) & (g2731) & (g2732) & (!g2738) & (g2779)) + ((g2218) & (g2436) & (g2731) & (g2732) & (g2738) & (!g2779)) + ((g2218) & (g2436) & (g2731) & (g2732) & (g2738) & (g2779)));
	assign g2822 = (((!g2436) & (!g2732) & (g2738) & (!g2779)) + ((!g2436) & (g2732) & (!g2738) & (!g2779)) + ((!g2436) & (g2732) & (!g2738) & (g2779)) + ((!g2436) & (g2732) & (g2738) & (g2779)) + ((g2436) & (!g2732) & (!g2738) & (!g2779)) + ((g2436) & (g2732) & (!g2738) & (g2779)) + ((g2436) & (g2732) & (g2738) & (!g2779)) + ((g2436) & (g2732) & (g2738) & (g2779)));
	assign g2823 = (((!g2398) & (!g2627) & (!g2734) & (g2735) & (g2737) & (!g2779)) + ((!g2398) & (!g2627) & (g2734) & (!g2735) & (!g2737) & (!g2779)) + ((!g2398) & (!g2627) & (g2734) & (!g2735) & (!g2737) & (g2779)) + ((!g2398) & (!g2627) & (g2734) & (!g2735) & (g2737) & (!g2779)) + ((!g2398) & (!g2627) & (g2734) & (!g2735) & (g2737) & (g2779)) + ((!g2398) & (!g2627) & (g2734) & (g2735) & (!g2737) & (!g2779)) + ((!g2398) & (!g2627) & (g2734) & (g2735) & (!g2737) & (g2779)) + ((!g2398) & (!g2627) & (g2734) & (g2735) & (g2737) & (g2779)) + ((!g2398) & (g2627) & (!g2734) & (!g2735) & (g2737) & (!g2779)) + ((!g2398) & (g2627) & (!g2734) & (g2735) & (!g2737) & (!g2779)) + ((!g2398) & (g2627) & (!g2734) & (g2735) & (g2737) & (!g2779)) + ((!g2398) & (g2627) & (g2734) & (!g2735) & (!g2737) & (!g2779)) + ((!g2398) & (g2627) & (g2734) & (!g2735) & (!g2737) & (g2779)) + ((!g2398) & (g2627) & (g2734) & (!g2735) & (g2737) & (g2779)) + ((!g2398) & (g2627) & (g2734) & (g2735) & (!g2737) & (g2779)) + ((!g2398) & (g2627) & (g2734) & (g2735) & (g2737) & (g2779)) + ((g2398) & (!g2627) & (!g2734) & (!g2735) & (!g2737) & (!g2779)) + ((g2398) & (!g2627) & (!g2734) & (!g2735) & (g2737) & (!g2779)) + ((g2398) & (!g2627) & (!g2734) & (g2735) & (!g2737) & (!g2779)) + ((g2398) & (!g2627) & (g2734) & (!g2735) & (!g2737) & (g2779)) + ((g2398) & (!g2627) & (g2734) & (!g2735) & (g2737) & (g2779)) + ((g2398) & (!g2627) & (g2734) & (g2735) & (!g2737) & (g2779)) + ((g2398) & (!g2627) & (g2734) & (g2735) & (g2737) & (!g2779)) + ((g2398) & (!g2627) & (g2734) & (g2735) & (g2737) & (g2779)) + ((g2398) & (g2627) & (!g2734) & (!g2735) & (!g2737) & (!g2779)) + ((g2398) & (g2627) & (g2734) & (!g2735) & (!g2737) & (g2779)) + ((g2398) & (g2627) & (g2734) & (!g2735) & (g2737) & (!g2779)) + ((g2398) & (g2627) & (g2734) & (!g2735) & (g2737) & (g2779)) + ((g2398) & (g2627) & (g2734) & (g2735) & (!g2737) & (!g2779)) + ((g2398) & (g2627) & (g2734) & (g2735) & (!g2737) & (g2779)) + ((g2398) & (g2627) & (g2734) & (g2735) & (g2737) & (!g2779)) + ((g2398) & (g2627) & (g2734) & (g2735) & (g2737) & (g2779)));
	assign g2824 = (((!g2627) & (!g2735) & (g2737) & (!g2779)) + ((!g2627) & (g2735) & (!g2737) & (!g2779)) + ((!g2627) & (g2735) & (!g2737) & (g2779)) + ((!g2627) & (g2735) & (g2737) & (g2779)) + ((g2627) & (!g2735) & (!g2737) & (!g2779)) + ((g2627) & (g2735) & (!g2737) & (g2779)) + ((g2627) & (g2735) & (g2737) & (!g2779)) + ((g2627) & (g2735) & (g2737) & (g2779)));
	assign g2825 = (((!g2653) & (g2668)));
	assign g2826 = (((!g2585) & (!ax18x) & (!ax19x) & (!g2825) & (!g2736) & (g2779)) + ((!g2585) & (!ax18x) & (!ax19x) & (!g2825) & (g2736) & (!g2779)) + ((!g2585) & (!ax18x) & (!ax19x) & (!g2825) & (g2736) & (g2779)) + ((!g2585) & (!ax18x) & (!ax19x) & (g2825) & (!g2736) & (!g2779)) + ((!g2585) & (!ax18x) & (ax19x) & (!g2825) & (!g2736) & (!g2779)) + ((!g2585) & (!ax18x) & (ax19x) & (g2825) & (!g2736) & (g2779)) + ((!g2585) & (!ax18x) & (ax19x) & (g2825) & (g2736) & (!g2779)) + ((!g2585) & (!ax18x) & (ax19x) & (g2825) & (g2736) & (g2779)) + ((!g2585) & (ax18x) & (!ax19x) & (g2825) & (!g2736) & (!g2779)) + ((!g2585) & (ax18x) & (!ax19x) & (g2825) & (g2736) & (!g2779)) + ((!g2585) & (ax18x) & (ax19x) & (!g2825) & (!g2736) & (!g2779)) + ((!g2585) & (ax18x) & (ax19x) & (!g2825) & (!g2736) & (g2779)) + ((!g2585) & (ax18x) & (ax19x) & (!g2825) & (g2736) & (!g2779)) + ((!g2585) & (ax18x) & (ax19x) & (!g2825) & (g2736) & (g2779)) + ((!g2585) & (ax18x) & (ax19x) & (g2825) & (!g2736) & (g2779)) + ((!g2585) & (ax18x) & (ax19x) & (g2825) & (g2736) & (g2779)) + ((g2585) & (!ax18x) & (!ax19x) & (!g2825) & (!g2736) & (!g2779)) + ((g2585) & (!ax18x) & (!ax19x) & (!g2825) & (!g2736) & (g2779)) + ((g2585) & (!ax18x) & (!ax19x) & (!g2825) & (g2736) & (g2779)) + ((g2585) & (!ax18x) & (!ax19x) & (g2825) & (g2736) & (!g2779)) + ((g2585) & (!ax18x) & (ax19x) & (!g2825) & (g2736) & (!g2779)) + ((g2585) & (!ax18x) & (ax19x) & (g2825) & (!g2736) & (!g2779)) + ((g2585) & (!ax18x) & (ax19x) & (g2825) & (!g2736) & (g2779)) + ((g2585) & (!ax18x) & (ax19x) & (g2825) & (g2736) & (g2779)) + ((g2585) & (ax18x) & (!ax19x) & (!g2825) & (!g2736) & (!g2779)) + ((g2585) & (ax18x) & (!ax19x) & (!g2825) & (g2736) & (!g2779)) + ((g2585) & (ax18x) & (ax19x) & (!g2825) & (!g2736) & (g2779)) + ((g2585) & (ax18x) & (ax19x) & (!g2825) & (g2736) & (g2779)) + ((g2585) & (ax18x) & (ax19x) & (g2825) & (!g2736) & (!g2779)) + ((g2585) & (ax18x) & (ax19x) & (g2825) & (!g2736) & (g2779)) + ((g2585) & (ax18x) & (ax19x) & (g2825) & (g2736) & (!g2779)) + ((g2585) & (ax18x) & (ax19x) & (g2825) & (g2736) & (g2779)));
	assign g2827 = (((!ax18x) & (!g2825) & (!g2736) & (g2779)) + ((!ax18x) & (!g2825) & (g2736) & (!g2779)) + ((!ax18x) & (!g2825) & (g2736) & (g2779)) + ((!ax18x) & (g2825) & (g2736) & (!g2779)) + ((ax18x) & (!g2825) & (!g2736) & (!g2779)) + ((ax18x) & (g2825) & (!g2736) & (!g2779)) + ((ax18x) & (g2825) & (!g2736) & (g2779)) + ((ax18x) & (g2825) & (g2736) & (g2779)));
	assign g2828 = (((!ax14x) & (!ax15x)));
	assign g2829 = (((!g2825) & (!ax16x) & (!ax17x) & (!g2779) & (!g2828)) + ((!g2825) & (!ax16x) & (ax17x) & (g2779) & (!g2828)) + ((!g2825) & (ax16x) & (ax17x) & (g2779) & (!g2828)) + ((!g2825) & (ax16x) & (ax17x) & (g2779) & (g2828)) + ((g2825) & (!ax16x) & (!ax17x) & (!g2779) & (!g2828)) + ((g2825) & (!ax16x) & (!ax17x) & (!g2779) & (g2828)) + ((g2825) & (!ax16x) & (!ax17x) & (g2779) & (!g2828)) + ((g2825) & (!ax16x) & (ax17x) & (!g2779) & (!g2828)) + ((g2825) & (!ax16x) & (ax17x) & (g2779) & (!g2828)) + ((g2825) & (!ax16x) & (ax17x) & (g2779) & (g2828)) + ((g2825) & (ax16x) & (!ax17x) & (g2779) & (!g2828)) + ((g2825) & (ax16x) & (!ax17x) & (g2779) & (g2828)) + ((g2825) & (ax16x) & (ax17x) & (!g2779) & (!g2828)) + ((g2825) & (ax16x) & (ax17x) & (!g2779) & (g2828)) + ((g2825) & (ax16x) & (ax17x) & (g2779) & (!g2828)) + ((g2825) & (ax16x) & (ax17x) & (g2779) & (g2828)));
	assign g2830 = (((!g2627) & (!g2585) & (g2826) & (g2827) & (g2829)) + ((!g2627) & (g2585) & (g2826) & (!g2827) & (g2829)) + ((!g2627) & (g2585) & (g2826) & (g2827) & (!g2829)) + ((!g2627) & (g2585) & (g2826) & (g2827) & (g2829)) + ((g2627) & (!g2585) & (!g2826) & (g2827) & (g2829)) + ((g2627) & (!g2585) & (g2826) & (!g2827) & (!g2829)) + ((g2627) & (!g2585) & (g2826) & (!g2827) & (g2829)) + ((g2627) & (!g2585) & (g2826) & (g2827) & (!g2829)) + ((g2627) & (!g2585) & (g2826) & (g2827) & (g2829)) + ((g2627) & (g2585) & (!g2826) & (!g2827) & (g2829)) + ((g2627) & (g2585) & (!g2826) & (g2827) & (!g2829)) + ((g2627) & (g2585) & (!g2826) & (g2827) & (g2829)) + ((g2627) & (g2585) & (g2826) & (!g2827) & (!g2829)) + ((g2627) & (g2585) & (g2826) & (!g2827) & (g2829)) + ((g2627) & (g2585) & (g2826) & (g2827) & (!g2829)) + ((g2627) & (g2585) & (g2826) & (g2827) & (g2829)));
	assign g2831 = (((!g2436) & (!g2398) & (g2823) & (g2824) & (g2830)) + ((!g2436) & (g2398) & (g2823) & (!g2824) & (g2830)) + ((!g2436) & (g2398) & (g2823) & (g2824) & (!g2830)) + ((!g2436) & (g2398) & (g2823) & (g2824) & (g2830)) + ((g2436) & (!g2398) & (!g2823) & (g2824) & (g2830)) + ((g2436) & (!g2398) & (g2823) & (!g2824) & (!g2830)) + ((g2436) & (!g2398) & (g2823) & (!g2824) & (g2830)) + ((g2436) & (!g2398) & (g2823) & (g2824) & (!g2830)) + ((g2436) & (!g2398) & (g2823) & (g2824) & (g2830)) + ((g2436) & (g2398) & (!g2823) & (!g2824) & (g2830)) + ((g2436) & (g2398) & (!g2823) & (g2824) & (!g2830)) + ((g2436) & (g2398) & (!g2823) & (g2824) & (g2830)) + ((g2436) & (g2398) & (g2823) & (!g2824) & (!g2830)) + ((g2436) & (g2398) & (g2823) & (!g2824) & (g2830)) + ((g2436) & (g2398) & (g2823) & (g2824) & (!g2830)) + ((g2436) & (g2398) & (g2823) & (g2824) & (g2830)));
	assign g2832 = (((!g2252) & (!g2218) & (g2821) & (g2822) & (g2831)) + ((!g2252) & (g2218) & (g2821) & (!g2822) & (g2831)) + ((!g2252) & (g2218) & (g2821) & (g2822) & (!g2831)) + ((!g2252) & (g2218) & (g2821) & (g2822) & (g2831)) + ((g2252) & (!g2218) & (!g2821) & (g2822) & (g2831)) + ((g2252) & (!g2218) & (g2821) & (!g2822) & (!g2831)) + ((g2252) & (!g2218) & (g2821) & (!g2822) & (g2831)) + ((g2252) & (!g2218) & (g2821) & (g2822) & (!g2831)) + ((g2252) & (!g2218) & (g2821) & (g2822) & (g2831)) + ((g2252) & (g2218) & (!g2821) & (!g2822) & (g2831)) + ((g2252) & (g2218) & (!g2821) & (g2822) & (!g2831)) + ((g2252) & (g2218) & (!g2821) & (g2822) & (g2831)) + ((g2252) & (g2218) & (g2821) & (!g2822) & (!g2831)) + ((g2252) & (g2218) & (g2821) & (!g2822) & (g2831)) + ((g2252) & (g2218) & (g2821) & (g2822) & (!g2831)) + ((g2252) & (g2218) & (g2821) & (g2822) & (g2831)));
	assign g2833 = (((!g2075) & (!g2045) & (g2819) & (g2820) & (g2832)) + ((!g2075) & (g2045) & (g2819) & (!g2820) & (g2832)) + ((!g2075) & (g2045) & (g2819) & (g2820) & (!g2832)) + ((!g2075) & (g2045) & (g2819) & (g2820) & (g2832)) + ((g2075) & (!g2045) & (!g2819) & (g2820) & (g2832)) + ((g2075) & (!g2045) & (g2819) & (!g2820) & (!g2832)) + ((g2075) & (!g2045) & (g2819) & (!g2820) & (g2832)) + ((g2075) & (!g2045) & (g2819) & (g2820) & (!g2832)) + ((g2075) & (!g2045) & (g2819) & (g2820) & (g2832)) + ((g2075) & (g2045) & (!g2819) & (!g2820) & (g2832)) + ((g2075) & (g2045) & (!g2819) & (g2820) & (!g2832)) + ((g2075) & (g2045) & (!g2819) & (g2820) & (g2832)) + ((g2075) & (g2045) & (g2819) & (!g2820) & (!g2832)) + ((g2075) & (g2045) & (g2819) & (!g2820) & (g2832)) + ((g2075) & (g2045) & (g2819) & (g2820) & (!g2832)) + ((g2075) & (g2045) & (g2819) & (g2820) & (g2832)));
	assign g2834 = (((!g1905) & (!g1879) & (g2817) & (g2818) & (g2833)) + ((!g1905) & (g1879) & (g2817) & (!g2818) & (g2833)) + ((!g1905) & (g1879) & (g2817) & (g2818) & (!g2833)) + ((!g1905) & (g1879) & (g2817) & (g2818) & (g2833)) + ((g1905) & (!g1879) & (!g2817) & (g2818) & (g2833)) + ((g1905) & (!g1879) & (g2817) & (!g2818) & (!g2833)) + ((g1905) & (!g1879) & (g2817) & (!g2818) & (g2833)) + ((g1905) & (!g1879) & (g2817) & (g2818) & (!g2833)) + ((g1905) & (!g1879) & (g2817) & (g2818) & (g2833)) + ((g1905) & (g1879) & (!g2817) & (!g2818) & (g2833)) + ((g1905) & (g1879) & (!g2817) & (g2818) & (!g2833)) + ((g1905) & (g1879) & (!g2817) & (g2818) & (g2833)) + ((g1905) & (g1879) & (g2817) & (!g2818) & (!g2833)) + ((g1905) & (g1879) & (g2817) & (!g2818) & (g2833)) + ((g1905) & (g1879) & (g2817) & (g2818) & (!g2833)) + ((g1905) & (g1879) & (g2817) & (g2818) & (g2833)));
	assign g2835 = (((!g1742) & (!g1720) & (g2815) & (g2816) & (g2834)) + ((!g1742) & (g1720) & (g2815) & (!g2816) & (g2834)) + ((!g1742) & (g1720) & (g2815) & (g2816) & (!g2834)) + ((!g1742) & (g1720) & (g2815) & (g2816) & (g2834)) + ((g1742) & (!g1720) & (!g2815) & (g2816) & (g2834)) + ((g1742) & (!g1720) & (g2815) & (!g2816) & (!g2834)) + ((g1742) & (!g1720) & (g2815) & (!g2816) & (g2834)) + ((g1742) & (!g1720) & (g2815) & (g2816) & (!g2834)) + ((g1742) & (!g1720) & (g2815) & (g2816) & (g2834)) + ((g1742) & (g1720) & (!g2815) & (!g2816) & (g2834)) + ((g1742) & (g1720) & (!g2815) & (g2816) & (!g2834)) + ((g1742) & (g1720) & (!g2815) & (g2816) & (g2834)) + ((g1742) & (g1720) & (g2815) & (!g2816) & (!g2834)) + ((g1742) & (g1720) & (g2815) & (!g2816) & (g2834)) + ((g1742) & (g1720) & (g2815) & (g2816) & (!g2834)) + ((g1742) & (g1720) & (g2815) & (g2816) & (g2834)));
	assign g2836 = (((!g1586) & (!g1568) & (g2813) & (g2814) & (g2835)) + ((!g1586) & (g1568) & (g2813) & (!g2814) & (g2835)) + ((!g1586) & (g1568) & (g2813) & (g2814) & (!g2835)) + ((!g1586) & (g1568) & (g2813) & (g2814) & (g2835)) + ((g1586) & (!g1568) & (!g2813) & (g2814) & (g2835)) + ((g1586) & (!g1568) & (g2813) & (!g2814) & (!g2835)) + ((g1586) & (!g1568) & (g2813) & (!g2814) & (g2835)) + ((g1586) & (!g1568) & (g2813) & (g2814) & (!g2835)) + ((g1586) & (!g1568) & (g2813) & (g2814) & (g2835)) + ((g1586) & (g1568) & (!g2813) & (!g2814) & (g2835)) + ((g1586) & (g1568) & (!g2813) & (g2814) & (!g2835)) + ((g1586) & (g1568) & (!g2813) & (g2814) & (g2835)) + ((g1586) & (g1568) & (g2813) & (!g2814) & (!g2835)) + ((g1586) & (g1568) & (g2813) & (!g2814) & (g2835)) + ((g1586) & (g1568) & (g2813) & (g2814) & (!g2835)) + ((g1586) & (g1568) & (g2813) & (g2814) & (g2835)));
	assign g2837 = (((!g1437) & (!g1423) & (g2811) & (g2812) & (g2836)) + ((!g1437) & (g1423) & (g2811) & (!g2812) & (g2836)) + ((!g1437) & (g1423) & (g2811) & (g2812) & (!g2836)) + ((!g1437) & (g1423) & (g2811) & (g2812) & (g2836)) + ((g1437) & (!g1423) & (!g2811) & (g2812) & (g2836)) + ((g1437) & (!g1423) & (g2811) & (!g2812) & (!g2836)) + ((g1437) & (!g1423) & (g2811) & (!g2812) & (g2836)) + ((g1437) & (!g1423) & (g2811) & (g2812) & (!g2836)) + ((g1437) & (!g1423) & (g2811) & (g2812) & (g2836)) + ((g1437) & (g1423) & (!g2811) & (!g2812) & (g2836)) + ((g1437) & (g1423) & (!g2811) & (g2812) & (!g2836)) + ((g1437) & (g1423) & (!g2811) & (g2812) & (g2836)) + ((g1437) & (g1423) & (g2811) & (!g2812) & (!g2836)) + ((g1437) & (g1423) & (g2811) & (!g2812) & (g2836)) + ((g1437) & (g1423) & (g2811) & (g2812) & (!g2836)) + ((g1437) & (g1423) & (g2811) & (g2812) & (g2836)));
	assign g2838 = (((!g1295) & (!g1285) & (g2809) & (g2810) & (g2837)) + ((!g1295) & (g1285) & (g2809) & (!g2810) & (g2837)) + ((!g1295) & (g1285) & (g2809) & (g2810) & (!g2837)) + ((!g1295) & (g1285) & (g2809) & (g2810) & (g2837)) + ((g1295) & (!g1285) & (!g2809) & (g2810) & (g2837)) + ((g1295) & (!g1285) & (g2809) & (!g2810) & (!g2837)) + ((g1295) & (!g1285) & (g2809) & (!g2810) & (g2837)) + ((g1295) & (!g1285) & (g2809) & (g2810) & (!g2837)) + ((g1295) & (!g1285) & (g2809) & (g2810) & (g2837)) + ((g1295) & (g1285) & (!g2809) & (!g2810) & (g2837)) + ((g1295) & (g1285) & (!g2809) & (g2810) & (!g2837)) + ((g1295) & (g1285) & (!g2809) & (g2810) & (g2837)) + ((g1295) & (g1285) & (g2809) & (!g2810) & (!g2837)) + ((g1295) & (g1285) & (g2809) & (!g2810) & (g2837)) + ((g1295) & (g1285) & (g2809) & (g2810) & (!g2837)) + ((g1295) & (g1285) & (g2809) & (g2810) & (g2837)));
	assign g2839 = (((!g1160) & (!g1154) & (g2807) & (g2808) & (g2838)) + ((!g1160) & (g1154) & (g2807) & (!g2808) & (g2838)) + ((!g1160) & (g1154) & (g2807) & (g2808) & (!g2838)) + ((!g1160) & (g1154) & (g2807) & (g2808) & (g2838)) + ((g1160) & (!g1154) & (!g2807) & (g2808) & (g2838)) + ((g1160) & (!g1154) & (g2807) & (!g2808) & (!g2838)) + ((g1160) & (!g1154) & (g2807) & (!g2808) & (g2838)) + ((g1160) & (!g1154) & (g2807) & (g2808) & (!g2838)) + ((g1160) & (!g1154) & (g2807) & (g2808) & (g2838)) + ((g1160) & (g1154) & (!g2807) & (!g2808) & (g2838)) + ((g1160) & (g1154) & (!g2807) & (g2808) & (!g2838)) + ((g1160) & (g1154) & (!g2807) & (g2808) & (g2838)) + ((g1160) & (g1154) & (g2807) & (!g2808) & (!g2838)) + ((g1160) & (g1154) & (g2807) & (!g2808) & (g2838)) + ((g1160) & (g1154) & (g2807) & (g2808) & (!g2838)) + ((g1160) & (g1154) & (g2807) & (g2808) & (g2838)));
	assign g2840 = (((!g1032) & (!g1030) & (g2805) & (g2806) & (g2839)) + ((!g1032) & (g1030) & (g2805) & (!g2806) & (g2839)) + ((!g1032) & (g1030) & (g2805) & (g2806) & (!g2839)) + ((!g1032) & (g1030) & (g2805) & (g2806) & (g2839)) + ((g1032) & (!g1030) & (!g2805) & (g2806) & (g2839)) + ((g1032) & (!g1030) & (g2805) & (!g2806) & (!g2839)) + ((g1032) & (!g1030) & (g2805) & (!g2806) & (g2839)) + ((g1032) & (!g1030) & (g2805) & (g2806) & (!g2839)) + ((g1032) & (!g1030) & (g2805) & (g2806) & (g2839)) + ((g1032) & (g1030) & (!g2805) & (!g2806) & (g2839)) + ((g1032) & (g1030) & (!g2805) & (g2806) & (!g2839)) + ((g1032) & (g1030) & (!g2805) & (g2806) & (g2839)) + ((g1032) & (g1030) & (g2805) & (!g2806) & (!g2839)) + ((g1032) & (g1030) & (g2805) & (!g2806) & (g2839)) + ((g1032) & (g1030) & (g2805) & (g2806) & (!g2839)) + ((g1032) & (g1030) & (g2805) & (g2806) & (g2839)));
	assign g2841 = (((!g851) & (!g914) & (g2803) & (g2804) & (g2840)) + ((!g851) & (g914) & (g2803) & (!g2804) & (g2840)) + ((!g851) & (g914) & (g2803) & (g2804) & (!g2840)) + ((!g851) & (g914) & (g2803) & (g2804) & (g2840)) + ((g851) & (!g914) & (!g2803) & (g2804) & (g2840)) + ((g851) & (!g914) & (g2803) & (!g2804) & (!g2840)) + ((g851) & (!g914) & (g2803) & (!g2804) & (g2840)) + ((g851) & (!g914) & (g2803) & (g2804) & (!g2840)) + ((g851) & (!g914) & (g2803) & (g2804) & (g2840)) + ((g851) & (g914) & (!g2803) & (!g2804) & (g2840)) + ((g851) & (g914) & (!g2803) & (g2804) & (!g2840)) + ((g851) & (g914) & (!g2803) & (g2804) & (g2840)) + ((g851) & (g914) & (g2803) & (!g2804) & (!g2840)) + ((g851) & (g914) & (g2803) & (!g2804) & (g2840)) + ((g851) & (g914) & (g2803) & (g2804) & (!g2840)) + ((g851) & (g914) & (g2803) & (g2804) & (g2840)));
	assign g2842 = (((!g744) & (!g803) & (g2801) & (g2802) & (g2841)) + ((!g744) & (g803) & (g2801) & (!g2802) & (g2841)) + ((!g744) & (g803) & (g2801) & (g2802) & (!g2841)) + ((!g744) & (g803) & (g2801) & (g2802) & (g2841)) + ((g744) & (!g803) & (!g2801) & (g2802) & (g2841)) + ((g744) & (!g803) & (g2801) & (!g2802) & (!g2841)) + ((g744) & (!g803) & (g2801) & (!g2802) & (g2841)) + ((g744) & (!g803) & (g2801) & (g2802) & (!g2841)) + ((g744) & (!g803) & (g2801) & (g2802) & (g2841)) + ((g744) & (g803) & (!g2801) & (!g2802) & (g2841)) + ((g744) & (g803) & (!g2801) & (g2802) & (!g2841)) + ((g744) & (g803) & (!g2801) & (g2802) & (g2841)) + ((g744) & (g803) & (g2801) & (!g2802) & (!g2841)) + ((g744) & (g803) & (g2801) & (!g2802) & (g2841)) + ((g744) & (g803) & (g2801) & (g2802) & (!g2841)) + ((g744) & (g803) & (g2801) & (g2802) & (g2841)));
	assign g2843 = (((!g645) & (!g700) & (g2799) & (g2800) & (g2842)) + ((!g645) & (g700) & (g2799) & (!g2800) & (g2842)) + ((!g645) & (g700) & (g2799) & (g2800) & (!g2842)) + ((!g645) & (g700) & (g2799) & (g2800) & (g2842)) + ((g645) & (!g700) & (!g2799) & (g2800) & (g2842)) + ((g645) & (!g700) & (g2799) & (!g2800) & (!g2842)) + ((g645) & (!g700) & (g2799) & (!g2800) & (g2842)) + ((g645) & (!g700) & (g2799) & (g2800) & (!g2842)) + ((g645) & (!g700) & (g2799) & (g2800) & (g2842)) + ((g645) & (g700) & (!g2799) & (!g2800) & (g2842)) + ((g645) & (g700) & (!g2799) & (g2800) & (!g2842)) + ((g645) & (g700) & (!g2799) & (g2800) & (g2842)) + ((g645) & (g700) & (g2799) & (!g2800) & (!g2842)) + ((g645) & (g700) & (g2799) & (!g2800) & (g2842)) + ((g645) & (g700) & (g2799) & (g2800) & (!g2842)) + ((g645) & (g700) & (g2799) & (g2800) & (g2842)));
	assign g2844 = (((!g553) & (!g604) & (g2797) & (g2798) & (g2843)) + ((!g553) & (g604) & (g2797) & (!g2798) & (g2843)) + ((!g553) & (g604) & (g2797) & (g2798) & (!g2843)) + ((!g553) & (g604) & (g2797) & (g2798) & (g2843)) + ((g553) & (!g604) & (!g2797) & (g2798) & (g2843)) + ((g553) & (!g604) & (g2797) & (!g2798) & (!g2843)) + ((g553) & (!g604) & (g2797) & (!g2798) & (g2843)) + ((g553) & (!g604) & (g2797) & (g2798) & (!g2843)) + ((g553) & (!g604) & (g2797) & (g2798) & (g2843)) + ((g553) & (g604) & (!g2797) & (!g2798) & (g2843)) + ((g553) & (g604) & (!g2797) & (g2798) & (!g2843)) + ((g553) & (g604) & (!g2797) & (g2798) & (g2843)) + ((g553) & (g604) & (g2797) & (!g2798) & (!g2843)) + ((g553) & (g604) & (g2797) & (!g2798) & (g2843)) + ((g553) & (g604) & (g2797) & (g2798) & (!g2843)) + ((g553) & (g604) & (g2797) & (g2798) & (g2843)));
	assign g2845 = (((!g468) & (!g515) & (g2795) & (g2796) & (g2844)) + ((!g468) & (g515) & (g2795) & (!g2796) & (g2844)) + ((!g468) & (g515) & (g2795) & (g2796) & (!g2844)) + ((!g468) & (g515) & (g2795) & (g2796) & (g2844)) + ((g468) & (!g515) & (!g2795) & (g2796) & (g2844)) + ((g468) & (!g515) & (g2795) & (!g2796) & (!g2844)) + ((g468) & (!g515) & (g2795) & (!g2796) & (g2844)) + ((g468) & (!g515) & (g2795) & (g2796) & (!g2844)) + ((g468) & (!g515) & (g2795) & (g2796) & (g2844)) + ((g468) & (g515) & (!g2795) & (!g2796) & (g2844)) + ((g468) & (g515) & (!g2795) & (g2796) & (!g2844)) + ((g468) & (g515) & (!g2795) & (g2796) & (g2844)) + ((g468) & (g515) & (g2795) & (!g2796) & (!g2844)) + ((g468) & (g515) & (g2795) & (!g2796) & (g2844)) + ((g468) & (g515) & (g2795) & (g2796) & (!g2844)) + ((g468) & (g515) & (g2795) & (g2796) & (g2844)));
	assign g2846 = (((!g390) & (!g433) & (g2793) & (g2794) & (g2845)) + ((!g390) & (g433) & (g2793) & (!g2794) & (g2845)) + ((!g390) & (g433) & (g2793) & (g2794) & (!g2845)) + ((!g390) & (g433) & (g2793) & (g2794) & (g2845)) + ((g390) & (!g433) & (!g2793) & (g2794) & (g2845)) + ((g390) & (!g433) & (g2793) & (!g2794) & (!g2845)) + ((g390) & (!g433) & (g2793) & (!g2794) & (g2845)) + ((g390) & (!g433) & (g2793) & (g2794) & (!g2845)) + ((g390) & (!g433) & (g2793) & (g2794) & (g2845)) + ((g390) & (g433) & (!g2793) & (!g2794) & (g2845)) + ((g390) & (g433) & (!g2793) & (g2794) & (!g2845)) + ((g390) & (g433) & (!g2793) & (g2794) & (g2845)) + ((g390) & (g433) & (g2793) & (!g2794) & (!g2845)) + ((g390) & (g433) & (g2793) & (!g2794) & (g2845)) + ((g390) & (g433) & (g2793) & (g2794) & (!g2845)) + ((g390) & (g433) & (g2793) & (g2794) & (g2845)));
	assign g2847 = (((!g319) & (!g358) & (g2791) & (g2792) & (g2846)) + ((!g319) & (g358) & (g2791) & (!g2792) & (g2846)) + ((!g319) & (g358) & (g2791) & (g2792) & (!g2846)) + ((!g319) & (g358) & (g2791) & (g2792) & (g2846)) + ((g319) & (!g358) & (!g2791) & (g2792) & (g2846)) + ((g319) & (!g358) & (g2791) & (!g2792) & (!g2846)) + ((g319) & (!g358) & (g2791) & (!g2792) & (g2846)) + ((g319) & (!g358) & (g2791) & (g2792) & (!g2846)) + ((g319) & (!g358) & (g2791) & (g2792) & (g2846)) + ((g319) & (g358) & (!g2791) & (!g2792) & (g2846)) + ((g319) & (g358) & (!g2791) & (g2792) & (!g2846)) + ((g319) & (g358) & (!g2791) & (g2792) & (g2846)) + ((g319) & (g358) & (g2791) & (!g2792) & (!g2846)) + ((g319) & (g358) & (g2791) & (!g2792) & (g2846)) + ((g319) & (g358) & (g2791) & (g2792) & (!g2846)) + ((g319) & (g358) & (g2791) & (g2792) & (g2846)));
	assign g2848 = (((!g255) & (!g290) & (g2789) & (g2790) & (g2847)) + ((!g255) & (g290) & (g2789) & (!g2790) & (g2847)) + ((!g255) & (g290) & (g2789) & (g2790) & (!g2847)) + ((!g255) & (g290) & (g2789) & (g2790) & (g2847)) + ((g255) & (!g290) & (!g2789) & (g2790) & (g2847)) + ((g255) & (!g290) & (g2789) & (!g2790) & (!g2847)) + ((g255) & (!g290) & (g2789) & (!g2790) & (g2847)) + ((g255) & (!g290) & (g2789) & (g2790) & (!g2847)) + ((g255) & (!g290) & (g2789) & (g2790) & (g2847)) + ((g255) & (g290) & (!g2789) & (!g2790) & (g2847)) + ((g255) & (g290) & (!g2789) & (g2790) & (!g2847)) + ((g255) & (g290) & (!g2789) & (g2790) & (g2847)) + ((g255) & (g290) & (g2789) & (!g2790) & (!g2847)) + ((g255) & (g290) & (g2789) & (!g2790) & (g2847)) + ((g255) & (g290) & (g2789) & (g2790) & (!g2847)) + ((g255) & (g290) & (g2789) & (g2790) & (g2847)));
	assign g2849 = (((!g198) & (!g229) & (g2787) & (g2788) & (g2848)) + ((!g198) & (g229) & (g2787) & (!g2788) & (g2848)) + ((!g198) & (g229) & (g2787) & (g2788) & (!g2848)) + ((!g198) & (g229) & (g2787) & (g2788) & (g2848)) + ((g198) & (!g229) & (!g2787) & (g2788) & (g2848)) + ((g198) & (!g229) & (g2787) & (!g2788) & (!g2848)) + ((g198) & (!g229) & (g2787) & (!g2788) & (g2848)) + ((g198) & (!g229) & (g2787) & (g2788) & (!g2848)) + ((g198) & (!g229) & (g2787) & (g2788) & (g2848)) + ((g198) & (g229) & (!g2787) & (!g2788) & (g2848)) + ((g198) & (g229) & (!g2787) & (g2788) & (!g2848)) + ((g198) & (g229) & (!g2787) & (g2788) & (g2848)) + ((g198) & (g229) & (g2787) & (!g2788) & (!g2848)) + ((g198) & (g229) & (g2787) & (!g2788) & (g2848)) + ((g198) & (g229) & (g2787) & (g2788) & (!g2848)) + ((g198) & (g229) & (g2787) & (g2788) & (g2848)));
	assign g2850 = (((!g147) & (!g174) & (g2785) & (g2786) & (g2849)) + ((!g147) & (g174) & (g2785) & (!g2786) & (g2849)) + ((!g147) & (g174) & (g2785) & (g2786) & (!g2849)) + ((!g147) & (g174) & (g2785) & (g2786) & (g2849)) + ((g147) & (!g174) & (!g2785) & (g2786) & (g2849)) + ((g147) & (!g174) & (g2785) & (!g2786) & (!g2849)) + ((g147) & (!g174) & (g2785) & (!g2786) & (g2849)) + ((g147) & (!g174) & (g2785) & (g2786) & (!g2849)) + ((g147) & (!g174) & (g2785) & (g2786) & (g2849)) + ((g147) & (g174) & (!g2785) & (!g2786) & (g2849)) + ((g147) & (g174) & (!g2785) & (g2786) & (!g2849)) + ((g147) & (g174) & (!g2785) & (g2786) & (g2849)) + ((g147) & (g174) & (g2785) & (!g2786) & (!g2849)) + ((g147) & (g174) & (g2785) & (!g2786) & (g2849)) + ((g147) & (g174) & (g2785) & (g2786) & (!g2849)) + ((g147) & (g174) & (g2785) & (g2786) & (g2849)));
	assign g2851 = (((!g104) & (!g127) & (g2783) & (g2784) & (g2850)) + ((!g104) & (g127) & (g2783) & (!g2784) & (g2850)) + ((!g104) & (g127) & (g2783) & (g2784) & (!g2850)) + ((!g104) & (g127) & (g2783) & (g2784) & (g2850)) + ((g104) & (!g127) & (!g2783) & (g2784) & (g2850)) + ((g104) & (!g127) & (g2783) & (!g2784) & (!g2850)) + ((g104) & (!g127) & (g2783) & (!g2784) & (g2850)) + ((g104) & (!g127) & (g2783) & (g2784) & (!g2850)) + ((g104) & (!g127) & (g2783) & (g2784) & (g2850)) + ((g104) & (g127) & (!g2783) & (!g2784) & (g2850)) + ((g104) & (g127) & (!g2783) & (g2784) & (!g2850)) + ((g104) & (g127) & (!g2783) & (g2784) & (g2850)) + ((g104) & (g127) & (g2783) & (!g2784) & (!g2850)) + ((g104) & (g127) & (g2783) & (!g2784) & (g2850)) + ((g104) & (g127) & (g2783) & (g2784) & (!g2850)) + ((g104) & (g127) & (g2783) & (g2784) & (g2850)));
	assign g2852 = (((!g68) & (!g87) & (g2781) & (g2782) & (g2851)) + ((!g68) & (g87) & (g2781) & (!g2782) & (g2851)) + ((!g68) & (g87) & (g2781) & (g2782) & (!g2851)) + ((!g68) & (g87) & (g2781) & (g2782) & (g2851)) + ((g68) & (!g87) & (!g2781) & (g2782) & (g2851)) + ((g68) & (!g87) & (g2781) & (!g2782) & (!g2851)) + ((g68) & (!g87) & (g2781) & (!g2782) & (g2851)) + ((g68) & (!g87) & (g2781) & (g2782) & (!g2851)) + ((g68) & (!g87) & (g2781) & (g2782) & (g2851)) + ((g68) & (g87) & (!g2781) & (!g2782) & (g2851)) + ((g68) & (g87) & (!g2781) & (g2782) & (!g2851)) + ((g68) & (g87) & (!g2781) & (g2782) & (g2851)) + ((g68) & (g87) & (g2781) & (!g2782) & (!g2851)) + ((g68) & (g87) & (g2781) & (!g2782) & (g2851)) + ((g68) & (g87) & (g2781) & (g2782) & (!g2851)) + ((g68) & (g87) & (g2781) & (g2782) & (g2851)));
	assign g2853 = (((g1) & (!g2760) & (g2775) & (g2778)) + ((g1) & (g2760) & (!g2775) & (!g2778)) + ((g1) & (g2760) & (!g2775) & (g2778)));
	assign g2854 = (((!g4) & (!g2) & (!g2761) & (!g2772) & (!g2774) & (!g2779)) + ((!g4) & (!g2) & (!g2761) & (!g2772) & (g2774) & (g2779)) + ((!g4) & (!g2) & (!g2761) & (g2772) & (!g2774) & (!g2779)) + ((!g4) & (!g2) & (!g2761) & (g2772) & (g2774) & (g2779)) + ((!g4) & (!g2) & (g2761) & (!g2772) & (!g2774) & (!g2779)) + ((!g4) & (!g2) & (g2761) & (!g2772) & (g2774) & (g2779)) + ((!g4) & (!g2) & (g2761) & (g2772) & (g2774) & (!g2779)) + ((!g4) & (!g2) & (g2761) & (g2772) & (g2774) & (g2779)) + ((!g4) & (g2) & (!g2761) & (!g2772) & (!g2774) & (!g2779)) + ((!g4) & (g2) & (!g2761) & (!g2772) & (g2774) & (g2779)) + ((!g4) & (g2) & (!g2761) & (g2772) & (g2774) & (!g2779)) + ((!g4) & (g2) & (!g2761) & (g2772) & (g2774) & (g2779)) + ((!g4) & (g2) & (g2761) & (!g2772) & (g2774) & (!g2779)) + ((!g4) & (g2) & (g2761) & (!g2772) & (g2774) & (g2779)) + ((!g4) & (g2) & (g2761) & (g2772) & (g2774) & (!g2779)) + ((!g4) & (g2) & (g2761) & (g2772) & (g2774) & (g2779)) + ((g4) & (!g2) & (!g2761) & (!g2772) & (g2774) & (!g2779)) + ((g4) & (!g2) & (!g2761) & (!g2772) & (g2774) & (g2779)) + ((g4) & (!g2) & (!g2761) & (g2772) & (g2774) & (!g2779)) + ((g4) & (!g2) & (!g2761) & (g2772) & (g2774) & (g2779)) + ((g4) & (!g2) & (g2761) & (!g2772) & (g2774) & (!g2779)) + ((g4) & (!g2) & (g2761) & (!g2772) & (g2774) & (g2779)) + ((g4) & (!g2) & (g2761) & (g2772) & (!g2774) & (!g2779)) + ((g4) & (!g2) & (g2761) & (g2772) & (g2774) & (g2779)) + ((g4) & (g2) & (!g2761) & (!g2772) & (g2774) & (!g2779)) + ((g4) & (g2) & (!g2761) & (!g2772) & (g2774) & (g2779)) + ((g4) & (g2) & (!g2761) & (g2772) & (!g2774) & (!g2779)) + ((g4) & (g2) & (!g2761) & (g2772) & (g2774) & (g2779)) + ((g4) & (g2) & (g2761) & (!g2772) & (!g2774) & (!g2779)) + ((g4) & (g2) & (g2761) & (!g2772) & (g2774) & (g2779)) + ((g4) & (g2) & (g2761) & (g2772) & (!g2774) & (!g2779)) + ((g4) & (g2) & (g2761) & (g2772) & (g2774) & (g2779)));
	assign g2855 = (((!g8) & (!g18) & (!g2763) & (g2764) & (g2771) & (!g2779)) + ((!g8) & (!g18) & (g2763) & (!g2764) & (!g2771) & (!g2779)) + ((!g8) & (!g18) & (g2763) & (!g2764) & (!g2771) & (g2779)) + ((!g8) & (!g18) & (g2763) & (!g2764) & (g2771) & (!g2779)) + ((!g8) & (!g18) & (g2763) & (!g2764) & (g2771) & (g2779)) + ((!g8) & (!g18) & (g2763) & (g2764) & (!g2771) & (!g2779)) + ((!g8) & (!g18) & (g2763) & (g2764) & (!g2771) & (g2779)) + ((!g8) & (!g18) & (g2763) & (g2764) & (g2771) & (g2779)) + ((!g8) & (g18) & (!g2763) & (!g2764) & (g2771) & (!g2779)) + ((!g8) & (g18) & (!g2763) & (g2764) & (!g2771) & (!g2779)) + ((!g8) & (g18) & (!g2763) & (g2764) & (g2771) & (!g2779)) + ((!g8) & (g18) & (g2763) & (!g2764) & (!g2771) & (!g2779)) + ((!g8) & (g18) & (g2763) & (!g2764) & (!g2771) & (g2779)) + ((!g8) & (g18) & (g2763) & (!g2764) & (g2771) & (g2779)) + ((!g8) & (g18) & (g2763) & (g2764) & (!g2771) & (g2779)) + ((!g8) & (g18) & (g2763) & (g2764) & (g2771) & (g2779)) + ((g8) & (!g18) & (!g2763) & (!g2764) & (!g2771) & (!g2779)) + ((g8) & (!g18) & (!g2763) & (!g2764) & (g2771) & (!g2779)) + ((g8) & (!g18) & (!g2763) & (g2764) & (!g2771) & (!g2779)) + ((g8) & (!g18) & (g2763) & (!g2764) & (!g2771) & (g2779)) + ((g8) & (!g18) & (g2763) & (!g2764) & (g2771) & (g2779)) + ((g8) & (!g18) & (g2763) & (g2764) & (!g2771) & (g2779)) + ((g8) & (!g18) & (g2763) & (g2764) & (g2771) & (!g2779)) + ((g8) & (!g18) & (g2763) & (g2764) & (g2771) & (g2779)) + ((g8) & (g18) & (!g2763) & (!g2764) & (!g2771) & (!g2779)) + ((g8) & (g18) & (g2763) & (!g2764) & (!g2771) & (g2779)) + ((g8) & (g18) & (g2763) & (!g2764) & (g2771) & (!g2779)) + ((g8) & (g18) & (g2763) & (!g2764) & (g2771) & (g2779)) + ((g8) & (g18) & (g2763) & (g2764) & (!g2771) & (!g2779)) + ((g8) & (g18) & (g2763) & (g2764) & (!g2771) & (g2779)) + ((g8) & (g18) & (g2763) & (g2764) & (g2771) & (!g2779)) + ((g8) & (g18) & (g2763) & (g2764) & (g2771) & (g2779)));
	assign g2856 = (((!g18) & (!g2764) & (g2771) & (!g2779)) + ((!g18) & (g2764) & (!g2771) & (!g2779)) + ((!g18) & (g2764) & (!g2771) & (g2779)) + ((!g18) & (g2764) & (g2771) & (g2779)) + ((g18) & (!g2764) & (!g2771) & (!g2779)) + ((g18) & (g2764) & (!g2771) & (g2779)) + ((g18) & (g2764) & (g2771) & (!g2779)) + ((g18) & (g2764) & (g2771) & (g2779)));
	assign g2857 = (((!g27) & (!g39) & (!g2766) & (g2767) & (g2770) & (!g2779)) + ((!g27) & (!g39) & (g2766) & (!g2767) & (!g2770) & (!g2779)) + ((!g27) & (!g39) & (g2766) & (!g2767) & (!g2770) & (g2779)) + ((!g27) & (!g39) & (g2766) & (!g2767) & (g2770) & (!g2779)) + ((!g27) & (!g39) & (g2766) & (!g2767) & (g2770) & (g2779)) + ((!g27) & (!g39) & (g2766) & (g2767) & (!g2770) & (!g2779)) + ((!g27) & (!g39) & (g2766) & (g2767) & (!g2770) & (g2779)) + ((!g27) & (!g39) & (g2766) & (g2767) & (g2770) & (g2779)) + ((!g27) & (g39) & (!g2766) & (!g2767) & (g2770) & (!g2779)) + ((!g27) & (g39) & (!g2766) & (g2767) & (!g2770) & (!g2779)) + ((!g27) & (g39) & (!g2766) & (g2767) & (g2770) & (!g2779)) + ((!g27) & (g39) & (g2766) & (!g2767) & (!g2770) & (!g2779)) + ((!g27) & (g39) & (g2766) & (!g2767) & (!g2770) & (g2779)) + ((!g27) & (g39) & (g2766) & (!g2767) & (g2770) & (g2779)) + ((!g27) & (g39) & (g2766) & (g2767) & (!g2770) & (g2779)) + ((!g27) & (g39) & (g2766) & (g2767) & (g2770) & (g2779)) + ((g27) & (!g39) & (!g2766) & (!g2767) & (!g2770) & (!g2779)) + ((g27) & (!g39) & (!g2766) & (!g2767) & (g2770) & (!g2779)) + ((g27) & (!g39) & (!g2766) & (g2767) & (!g2770) & (!g2779)) + ((g27) & (!g39) & (g2766) & (!g2767) & (!g2770) & (g2779)) + ((g27) & (!g39) & (g2766) & (!g2767) & (g2770) & (g2779)) + ((g27) & (!g39) & (g2766) & (g2767) & (!g2770) & (g2779)) + ((g27) & (!g39) & (g2766) & (g2767) & (g2770) & (!g2779)) + ((g27) & (!g39) & (g2766) & (g2767) & (g2770) & (g2779)) + ((g27) & (g39) & (!g2766) & (!g2767) & (!g2770) & (!g2779)) + ((g27) & (g39) & (g2766) & (!g2767) & (!g2770) & (g2779)) + ((g27) & (g39) & (g2766) & (!g2767) & (g2770) & (!g2779)) + ((g27) & (g39) & (g2766) & (!g2767) & (g2770) & (g2779)) + ((g27) & (g39) & (g2766) & (g2767) & (!g2770) & (!g2779)) + ((g27) & (g39) & (g2766) & (g2767) & (!g2770) & (g2779)) + ((g27) & (g39) & (g2766) & (g2767) & (g2770) & (!g2779)) + ((g27) & (g39) & (g2766) & (g2767) & (g2770) & (g2779)));
	assign g2858 = (((!g39) & (!g2767) & (g2770) & (!g2779)) + ((!g39) & (g2767) & (!g2770) & (!g2779)) + ((!g39) & (g2767) & (!g2770) & (g2779)) + ((!g39) & (g2767) & (g2770) & (g2779)) + ((g39) & (!g2767) & (!g2770) & (!g2779)) + ((g39) & (g2767) & (!g2770) & (g2779)) + ((g39) & (g2767) & (g2770) & (!g2779)) + ((g39) & (g2767) & (g2770) & (g2779)));
	assign g2859 = (((!g54) & (!g68) & (!g2769) & (g2669) & (g2759) & (!g2779)) + ((!g54) & (!g68) & (g2769) & (!g2669) & (!g2759) & (!g2779)) + ((!g54) & (!g68) & (g2769) & (!g2669) & (!g2759) & (g2779)) + ((!g54) & (!g68) & (g2769) & (!g2669) & (g2759) & (!g2779)) + ((!g54) & (!g68) & (g2769) & (!g2669) & (g2759) & (g2779)) + ((!g54) & (!g68) & (g2769) & (g2669) & (!g2759) & (!g2779)) + ((!g54) & (!g68) & (g2769) & (g2669) & (!g2759) & (g2779)) + ((!g54) & (!g68) & (g2769) & (g2669) & (g2759) & (g2779)) + ((!g54) & (g68) & (!g2769) & (!g2669) & (g2759) & (!g2779)) + ((!g54) & (g68) & (!g2769) & (g2669) & (!g2759) & (!g2779)) + ((!g54) & (g68) & (!g2769) & (g2669) & (g2759) & (!g2779)) + ((!g54) & (g68) & (g2769) & (!g2669) & (!g2759) & (!g2779)) + ((!g54) & (g68) & (g2769) & (!g2669) & (!g2759) & (g2779)) + ((!g54) & (g68) & (g2769) & (!g2669) & (g2759) & (g2779)) + ((!g54) & (g68) & (g2769) & (g2669) & (!g2759) & (g2779)) + ((!g54) & (g68) & (g2769) & (g2669) & (g2759) & (g2779)) + ((g54) & (!g68) & (!g2769) & (!g2669) & (!g2759) & (!g2779)) + ((g54) & (!g68) & (!g2769) & (!g2669) & (g2759) & (!g2779)) + ((g54) & (!g68) & (!g2769) & (g2669) & (!g2759) & (!g2779)) + ((g54) & (!g68) & (g2769) & (!g2669) & (!g2759) & (g2779)) + ((g54) & (!g68) & (g2769) & (!g2669) & (g2759) & (g2779)) + ((g54) & (!g68) & (g2769) & (g2669) & (!g2759) & (g2779)) + ((g54) & (!g68) & (g2769) & (g2669) & (g2759) & (!g2779)) + ((g54) & (!g68) & (g2769) & (g2669) & (g2759) & (g2779)) + ((g54) & (g68) & (!g2769) & (!g2669) & (!g2759) & (!g2779)) + ((g54) & (g68) & (g2769) & (!g2669) & (!g2759) & (g2779)) + ((g54) & (g68) & (g2769) & (!g2669) & (g2759) & (!g2779)) + ((g54) & (g68) & (g2769) & (!g2669) & (g2759) & (g2779)) + ((g54) & (g68) & (g2769) & (g2669) & (!g2759) & (!g2779)) + ((g54) & (g68) & (g2769) & (g2669) & (!g2759) & (g2779)) + ((g54) & (g68) & (g2769) & (g2669) & (g2759) & (!g2779)) + ((g54) & (g68) & (g2769) & (g2669) & (g2759) & (g2779)));
	assign g2860 = (((!g39) & (!g54) & (g2859) & (g2780) & (g2852)) + ((!g39) & (g54) & (g2859) & (!g2780) & (g2852)) + ((!g39) & (g54) & (g2859) & (g2780) & (!g2852)) + ((!g39) & (g54) & (g2859) & (g2780) & (g2852)) + ((g39) & (!g54) & (!g2859) & (g2780) & (g2852)) + ((g39) & (!g54) & (g2859) & (!g2780) & (!g2852)) + ((g39) & (!g54) & (g2859) & (!g2780) & (g2852)) + ((g39) & (!g54) & (g2859) & (g2780) & (!g2852)) + ((g39) & (!g54) & (g2859) & (g2780) & (g2852)) + ((g39) & (g54) & (!g2859) & (!g2780) & (g2852)) + ((g39) & (g54) & (!g2859) & (g2780) & (!g2852)) + ((g39) & (g54) & (!g2859) & (g2780) & (g2852)) + ((g39) & (g54) & (g2859) & (!g2780) & (!g2852)) + ((g39) & (g54) & (g2859) & (!g2780) & (g2852)) + ((g39) & (g54) & (g2859) & (g2780) & (!g2852)) + ((g39) & (g54) & (g2859) & (g2780) & (g2852)));
	assign g2861 = (((!g18) & (!g27) & (g2857) & (g2858) & (g2860)) + ((!g18) & (g27) & (g2857) & (!g2858) & (g2860)) + ((!g18) & (g27) & (g2857) & (g2858) & (!g2860)) + ((!g18) & (g27) & (g2857) & (g2858) & (g2860)) + ((g18) & (!g27) & (!g2857) & (g2858) & (g2860)) + ((g18) & (!g27) & (g2857) & (!g2858) & (!g2860)) + ((g18) & (!g27) & (g2857) & (!g2858) & (g2860)) + ((g18) & (!g27) & (g2857) & (g2858) & (!g2860)) + ((g18) & (!g27) & (g2857) & (g2858) & (g2860)) + ((g18) & (g27) & (!g2857) & (!g2858) & (g2860)) + ((g18) & (g27) & (!g2857) & (g2858) & (!g2860)) + ((g18) & (g27) & (!g2857) & (g2858) & (g2860)) + ((g18) & (g27) & (g2857) & (!g2858) & (!g2860)) + ((g18) & (g27) & (g2857) & (!g2858) & (g2860)) + ((g18) & (g27) & (g2857) & (g2858) & (!g2860)) + ((g18) & (g27) & (g2857) & (g2858) & (g2860)));
	assign g2862 = (((!g2) & (!g8) & (g2855) & (g2856) & (g2861)) + ((!g2) & (g8) & (g2855) & (!g2856) & (g2861)) + ((!g2) & (g8) & (g2855) & (g2856) & (!g2861)) + ((!g2) & (g8) & (g2855) & (g2856) & (g2861)) + ((g2) & (!g8) & (!g2855) & (g2856) & (g2861)) + ((g2) & (!g8) & (g2855) & (!g2856) & (!g2861)) + ((g2) & (!g8) & (g2855) & (!g2856) & (g2861)) + ((g2) & (!g8) & (g2855) & (g2856) & (!g2861)) + ((g2) & (!g8) & (g2855) & (g2856) & (g2861)) + ((g2) & (g8) & (!g2855) & (!g2856) & (g2861)) + ((g2) & (g8) & (!g2855) & (g2856) & (!g2861)) + ((g2) & (g8) & (!g2855) & (g2856) & (g2861)) + ((g2) & (g8) & (g2855) & (!g2856) & (!g2861)) + ((g2) & (g8) & (g2855) & (!g2856) & (g2861)) + ((g2) & (g8) & (g2855) & (g2856) & (!g2861)) + ((g2) & (g8) & (g2855) & (g2856) & (g2861)));
	assign g2863 = (((!g2) & (!g2761) & (g2772) & (!g2779)) + ((!g2) & (g2761) & (!g2772) & (!g2779)) + ((!g2) & (g2761) & (!g2772) & (g2779)) + ((!g2) & (g2761) & (g2772) & (g2779)) + ((g2) & (!g2761) & (!g2772) & (!g2779)) + ((g2) & (g2761) & (!g2772) & (g2779)) + ((g2) & (g2761) & (g2772) & (!g2779)) + ((g2) & (g2761) & (g2772) & (g2779)));
	assign g2864 = (((!g1) & (!g2760) & (!g2775) & (!g2777) & (g2778)) + ((!g1) & (!g2760) & (!g2775) & (g2777) & (!g2778)) + ((!g1) & (!g2760) & (!g2775) & (g2777) & (g2778)) + ((!g1) & (g2760) & (g2775) & (!g2777) & (!g2778)) + ((!g1) & (g2760) & (g2775) & (!g2777) & (g2778)) + ((!g1) & (g2760) & (g2775) & (g2777) & (!g2778)) + ((!g1) & (g2760) & (g2775) & (g2777) & (g2778)) + ((g1) & (!g2760) & (!g2775) & (!g2777) & (g2778)) + ((g1) & (!g2760) & (!g2775) & (g2777) & (g2778)) + ((g1) & (g2760) & (g2775) & (!g2777) & (!g2778)) + ((g1) & (g2760) & (g2775) & (!g2777) & (g2778)) + ((g1) & (g2760) & (g2775) & (g2777) & (!g2778)) + ((g1) & (g2760) & (g2775) & (g2777) & (g2778)));
	assign g2865 = (((!g4) & (!g1) & (!g2854) & (!g2862) & (!g2863) & (!g2864)) + ((!g4) & (g1) & (!g2854) & (!g2862) & (!g2863) & (!g2864)) + ((!g4) & (g1) & (!g2854) & (!g2862) & (!g2863) & (g2864)) + ((!g4) & (g1) & (!g2854) & (!g2862) & (g2863) & (!g2864)) + ((!g4) & (g1) & (!g2854) & (!g2862) & (g2863) & (g2864)) + ((!g4) & (g1) & (!g2854) & (g2862) & (!g2863) & (!g2864)) + ((!g4) & (g1) & (!g2854) & (g2862) & (!g2863) & (g2864)) + ((!g4) & (g1) & (!g2854) & (g2862) & (g2863) & (!g2864)) + ((!g4) & (g1) & (!g2854) & (g2862) & (g2863) & (g2864)) + ((!g4) & (g1) & (g2854) & (!g2862) & (!g2863) & (!g2864)) + ((!g4) & (g1) & (g2854) & (!g2862) & (!g2863) & (g2864)) + ((g4) & (!g1) & (!g2854) & (!g2862) & (!g2863) & (!g2864)) + ((g4) & (!g1) & (!g2854) & (!g2862) & (g2863) & (!g2864)) + ((g4) & (!g1) & (!g2854) & (g2862) & (!g2863) & (!g2864)) + ((g4) & (g1) & (!g2854) & (!g2862) & (!g2863) & (!g2864)) + ((g4) & (g1) & (!g2854) & (!g2862) & (!g2863) & (g2864)) + ((g4) & (g1) & (!g2854) & (!g2862) & (g2863) & (!g2864)) + ((g4) & (g1) & (!g2854) & (!g2862) & (g2863) & (g2864)) + ((g4) & (g1) & (!g2854) & (g2862) & (!g2863) & (!g2864)) + ((g4) & (g1) & (!g2854) & (g2862) & (!g2863) & (g2864)) + ((g4) & (g1) & (!g2854) & (g2862) & (g2863) & (!g2864)) + ((g4) & (g1) & (!g2854) & (g2862) & (g2863) & (g2864)) + ((g4) & (g1) & (g2854) & (!g2862) & (!g2863) & (!g2864)) + ((g4) & (g1) & (g2854) & (!g2862) & (!g2863) & (g2864)) + ((g4) & (g1) & (g2854) & (!g2862) & (g2863) & (!g2864)) + ((g4) & (g1) & (g2854) & (!g2862) & (g2863) & (g2864)) + ((g4) & (g1) & (g2854) & (g2862) & (!g2863) & (!g2864)) + ((g4) & (g1) & (g2854) & (g2862) & (!g2863) & (g2864)));
	assign g2866 = (((!g54) & (!g2780) & (g2852) & (!g2853) & (!g2865)) + ((!g54) & (!g2780) & (g2852) & (g2853) & (!g2865)) + ((!g54) & (!g2780) & (g2852) & (g2853) & (g2865)) + ((!g54) & (g2780) & (!g2852) & (!g2853) & (!g2865)) + ((!g54) & (g2780) & (!g2852) & (!g2853) & (g2865)) + ((!g54) & (g2780) & (!g2852) & (g2853) & (!g2865)) + ((!g54) & (g2780) & (!g2852) & (g2853) & (g2865)) + ((!g54) & (g2780) & (g2852) & (!g2853) & (g2865)) + ((g54) & (!g2780) & (!g2852) & (!g2853) & (!g2865)) + ((g54) & (!g2780) & (!g2852) & (g2853) & (!g2865)) + ((g54) & (!g2780) & (!g2852) & (g2853) & (g2865)) + ((g54) & (g2780) & (!g2852) & (!g2853) & (g2865)) + ((g54) & (g2780) & (g2852) & (!g2853) & (!g2865)) + ((g54) & (g2780) & (g2852) & (!g2853) & (g2865)) + ((g54) & (g2780) & (g2852) & (g2853) & (!g2865)) + ((g54) & (g2780) & (g2852) & (g2853) & (g2865)));
	assign g2867 = (((!g68) & (!g87) & (g2782) & (g2851)) + ((!g68) & (g87) & (!g2782) & (g2851)) + ((!g68) & (g87) & (g2782) & (!g2851)) + ((!g68) & (g87) & (g2782) & (g2851)) + ((g68) & (!g87) & (!g2782) & (!g2851)) + ((g68) & (!g87) & (!g2782) & (g2851)) + ((g68) & (!g87) & (g2782) & (!g2851)) + ((g68) & (g87) & (!g2782) & (!g2851)));
	assign g2868 = (((!g2781) & (!g2853) & (!g2865) & (g2867)) + ((!g2781) & (g2853) & (!g2865) & (g2867)) + ((!g2781) & (g2853) & (g2865) & (g2867)) + ((g2781) & (!g2853) & (!g2865) & (!g2867)) + ((g2781) & (!g2853) & (g2865) & (!g2867)) + ((g2781) & (!g2853) & (g2865) & (g2867)) + ((g2781) & (g2853) & (!g2865) & (!g2867)) + ((g2781) & (g2853) & (g2865) & (!g2867)));
	assign g2869 = (((!g87) & (!g2782) & (g2851) & (!g2853) & (!g2865)) + ((!g87) & (!g2782) & (g2851) & (g2853) & (!g2865)) + ((!g87) & (!g2782) & (g2851) & (g2853) & (g2865)) + ((!g87) & (g2782) & (!g2851) & (!g2853) & (!g2865)) + ((!g87) & (g2782) & (!g2851) & (!g2853) & (g2865)) + ((!g87) & (g2782) & (!g2851) & (g2853) & (!g2865)) + ((!g87) & (g2782) & (!g2851) & (g2853) & (g2865)) + ((!g87) & (g2782) & (g2851) & (!g2853) & (g2865)) + ((g87) & (!g2782) & (!g2851) & (!g2853) & (!g2865)) + ((g87) & (!g2782) & (!g2851) & (g2853) & (!g2865)) + ((g87) & (!g2782) & (!g2851) & (g2853) & (g2865)) + ((g87) & (g2782) & (!g2851) & (!g2853) & (g2865)) + ((g87) & (g2782) & (g2851) & (!g2853) & (!g2865)) + ((g87) & (g2782) & (g2851) & (!g2853) & (g2865)) + ((g87) & (g2782) & (g2851) & (g2853) & (!g2865)) + ((g87) & (g2782) & (g2851) & (g2853) & (g2865)));
	assign g2870 = (((!g104) & (!g127) & (g2784) & (g2850)) + ((!g104) & (g127) & (!g2784) & (g2850)) + ((!g104) & (g127) & (g2784) & (!g2850)) + ((!g104) & (g127) & (g2784) & (g2850)) + ((g104) & (!g127) & (!g2784) & (!g2850)) + ((g104) & (!g127) & (!g2784) & (g2850)) + ((g104) & (!g127) & (g2784) & (!g2850)) + ((g104) & (g127) & (!g2784) & (!g2850)));
	assign g2871 = (((!g2783) & (!g2853) & (!g2865) & (g2870)) + ((!g2783) & (g2853) & (!g2865) & (g2870)) + ((!g2783) & (g2853) & (g2865) & (g2870)) + ((g2783) & (!g2853) & (!g2865) & (!g2870)) + ((g2783) & (!g2853) & (g2865) & (!g2870)) + ((g2783) & (!g2853) & (g2865) & (g2870)) + ((g2783) & (g2853) & (!g2865) & (!g2870)) + ((g2783) & (g2853) & (g2865) & (!g2870)));
	assign g2872 = (((!g127) & (!g2784) & (g2850) & (!g2853) & (!g2865)) + ((!g127) & (!g2784) & (g2850) & (g2853) & (!g2865)) + ((!g127) & (!g2784) & (g2850) & (g2853) & (g2865)) + ((!g127) & (g2784) & (!g2850) & (!g2853) & (!g2865)) + ((!g127) & (g2784) & (!g2850) & (!g2853) & (g2865)) + ((!g127) & (g2784) & (!g2850) & (g2853) & (!g2865)) + ((!g127) & (g2784) & (!g2850) & (g2853) & (g2865)) + ((!g127) & (g2784) & (g2850) & (!g2853) & (g2865)) + ((g127) & (!g2784) & (!g2850) & (!g2853) & (!g2865)) + ((g127) & (!g2784) & (!g2850) & (g2853) & (!g2865)) + ((g127) & (!g2784) & (!g2850) & (g2853) & (g2865)) + ((g127) & (g2784) & (!g2850) & (!g2853) & (g2865)) + ((g127) & (g2784) & (g2850) & (!g2853) & (!g2865)) + ((g127) & (g2784) & (g2850) & (!g2853) & (g2865)) + ((g127) & (g2784) & (g2850) & (g2853) & (!g2865)) + ((g127) & (g2784) & (g2850) & (g2853) & (g2865)));
	assign g2873 = (((!g147) & (!g174) & (g2786) & (g2849)) + ((!g147) & (g174) & (!g2786) & (g2849)) + ((!g147) & (g174) & (g2786) & (!g2849)) + ((!g147) & (g174) & (g2786) & (g2849)) + ((g147) & (!g174) & (!g2786) & (!g2849)) + ((g147) & (!g174) & (!g2786) & (g2849)) + ((g147) & (!g174) & (g2786) & (!g2849)) + ((g147) & (g174) & (!g2786) & (!g2849)));
	assign g2874 = (((!g2785) & (!g2853) & (!g2865) & (g2873)) + ((!g2785) & (g2853) & (!g2865) & (g2873)) + ((!g2785) & (g2853) & (g2865) & (g2873)) + ((g2785) & (!g2853) & (!g2865) & (!g2873)) + ((g2785) & (!g2853) & (g2865) & (!g2873)) + ((g2785) & (!g2853) & (g2865) & (g2873)) + ((g2785) & (g2853) & (!g2865) & (!g2873)) + ((g2785) & (g2853) & (g2865) & (!g2873)));
	assign g2875 = (((!g174) & (!g2786) & (g2849) & (!g2853) & (!g2865)) + ((!g174) & (!g2786) & (g2849) & (g2853) & (!g2865)) + ((!g174) & (!g2786) & (g2849) & (g2853) & (g2865)) + ((!g174) & (g2786) & (!g2849) & (!g2853) & (!g2865)) + ((!g174) & (g2786) & (!g2849) & (!g2853) & (g2865)) + ((!g174) & (g2786) & (!g2849) & (g2853) & (!g2865)) + ((!g174) & (g2786) & (!g2849) & (g2853) & (g2865)) + ((!g174) & (g2786) & (g2849) & (!g2853) & (g2865)) + ((g174) & (!g2786) & (!g2849) & (!g2853) & (!g2865)) + ((g174) & (!g2786) & (!g2849) & (g2853) & (!g2865)) + ((g174) & (!g2786) & (!g2849) & (g2853) & (g2865)) + ((g174) & (g2786) & (!g2849) & (!g2853) & (g2865)) + ((g174) & (g2786) & (g2849) & (!g2853) & (!g2865)) + ((g174) & (g2786) & (g2849) & (!g2853) & (g2865)) + ((g174) & (g2786) & (g2849) & (g2853) & (!g2865)) + ((g174) & (g2786) & (g2849) & (g2853) & (g2865)));
	assign g2876 = (((!g198) & (!g229) & (g2788) & (g2848)) + ((!g198) & (g229) & (!g2788) & (g2848)) + ((!g198) & (g229) & (g2788) & (!g2848)) + ((!g198) & (g229) & (g2788) & (g2848)) + ((g198) & (!g229) & (!g2788) & (!g2848)) + ((g198) & (!g229) & (!g2788) & (g2848)) + ((g198) & (!g229) & (g2788) & (!g2848)) + ((g198) & (g229) & (!g2788) & (!g2848)));
	assign g2877 = (((!g2787) & (!g2853) & (!g2865) & (g2876)) + ((!g2787) & (g2853) & (!g2865) & (g2876)) + ((!g2787) & (g2853) & (g2865) & (g2876)) + ((g2787) & (!g2853) & (!g2865) & (!g2876)) + ((g2787) & (!g2853) & (g2865) & (!g2876)) + ((g2787) & (!g2853) & (g2865) & (g2876)) + ((g2787) & (g2853) & (!g2865) & (!g2876)) + ((g2787) & (g2853) & (g2865) & (!g2876)));
	assign g2878 = (((!g229) & (!g2788) & (g2848) & (!g2853) & (!g2865)) + ((!g229) & (!g2788) & (g2848) & (g2853) & (!g2865)) + ((!g229) & (!g2788) & (g2848) & (g2853) & (g2865)) + ((!g229) & (g2788) & (!g2848) & (!g2853) & (!g2865)) + ((!g229) & (g2788) & (!g2848) & (!g2853) & (g2865)) + ((!g229) & (g2788) & (!g2848) & (g2853) & (!g2865)) + ((!g229) & (g2788) & (!g2848) & (g2853) & (g2865)) + ((!g229) & (g2788) & (g2848) & (!g2853) & (g2865)) + ((g229) & (!g2788) & (!g2848) & (!g2853) & (!g2865)) + ((g229) & (!g2788) & (!g2848) & (g2853) & (!g2865)) + ((g229) & (!g2788) & (!g2848) & (g2853) & (g2865)) + ((g229) & (g2788) & (!g2848) & (!g2853) & (g2865)) + ((g229) & (g2788) & (g2848) & (!g2853) & (!g2865)) + ((g229) & (g2788) & (g2848) & (!g2853) & (g2865)) + ((g229) & (g2788) & (g2848) & (g2853) & (!g2865)) + ((g229) & (g2788) & (g2848) & (g2853) & (g2865)));
	assign g2879 = (((!g255) & (!g290) & (g2790) & (g2847)) + ((!g255) & (g290) & (!g2790) & (g2847)) + ((!g255) & (g290) & (g2790) & (!g2847)) + ((!g255) & (g290) & (g2790) & (g2847)) + ((g255) & (!g290) & (!g2790) & (!g2847)) + ((g255) & (!g290) & (!g2790) & (g2847)) + ((g255) & (!g290) & (g2790) & (!g2847)) + ((g255) & (g290) & (!g2790) & (!g2847)));
	assign g2880 = (((!g2789) & (!g2853) & (!g2865) & (g2879)) + ((!g2789) & (g2853) & (!g2865) & (g2879)) + ((!g2789) & (g2853) & (g2865) & (g2879)) + ((g2789) & (!g2853) & (!g2865) & (!g2879)) + ((g2789) & (!g2853) & (g2865) & (!g2879)) + ((g2789) & (!g2853) & (g2865) & (g2879)) + ((g2789) & (g2853) & (!g2865) & (!g2879)) + ((g2789) & (g2853) & (g2865) & (!g2879)));
	assign g2881 = (((!g290) & (!g2790) & (g2847) & (!g2853) & (!g2865)) + ((!g290) & (!g2790) & (g2847) & (g2853) & (!g2865)) + ((!g290) & (!g2790) & (g2847) & (g2853) & (g2865)) + ((!g290) & (g2790) & (!g2847) & (!g2853) & (!g2865)) + ((!g290) & (g2790) & (!g2847) & (!g2853) & (g2865)) + ((!g290) & (g2790) & (!g2847) & (g2853) & (!g2865)) + ((!g290) & (g2790) & (!g2847) & (g2853) & (g2865)) + ((!g290) & (g2790) & (g2847) & (!g2853) & (g2865)) + ((g290) & (!g2790) & (!g2847) & (!g2853) & (!g2865)) + ((g290) & (!g2790) & (!g2847) & (g2853) & (!g2865)) + ((g290) & (!g2790) & (!g2847) & (g2853) & (g2865)) + ((g290) & (g2790) & (!g2847) & (!g2853) & (g2865)) + ((g290) & (g2790) & (g2847) & (!g2853) & (!g2865)) + ((g290) & (g2790) & (g2847) & (!g2853) & (g2865)) + ((g290) & (g2790) & (g2847) & (g2853) & (!g2865)) + ((g290) & (g2790) & (g2847) & (g2853) & (g2865)));
	assign g2882 = (((!g319) & (!g358) & (g2792) & (g2846)) + ((!g319) & (g358) & (!g2792) & (g2846)) + ((!g319) & (g358) & (g2792) & (!g2846)) + ((!g319) & (g358) & (g2792) & (g2846)) + ((g319) & (!g358) & (!g2792) & (!g2846)) + ((g319) & (!g358) & (!g2792) & (g2846)) + ((g319) & (!g358) & (g2792) & (!g2846)) + ((g319) & (g358) & (!g2792) & (!g2846)));
	assign g2883 = (((!g2791) & (!g2853) & (!g2865) & (g2882)) + ((!g2791) & (g2853) & (!g2865) & (g2882)) + ((!g2791) & (g2853) & (g2865) & (g2882)) + ((g2791) & (!g2853) & (!g2865) & (!g2882)) + ((g2791) & (!g2853) & (g2865) & (!g2882)) + ((g2791) & (!g2853) & (g2865) & (g2882)) + ((g2791) & (g2853) & (!g2865) & (!g2882)) + ((g2791) & (g2853) & (g2865) & (!g2882)));
	assign g2884 = (((!g358) & (!g2792) & (g2846) & (!g2853) & (!g2865)) + ((!g358) & (!g2792) & (g2846) & (g2853) & (!g2865)) + ((!g358) & (!g2792) & (g2846) & (g2853) & (g2865)) + ((!g358) & (g2792) & (!g2846) & (!g2853) & (!g2865)) + ((!g358) & (g2792) & (!g2846) & (!g2853) & (g2865)) + ((!g358) & (g2792) & (!g2846) & (g2853) & (!g2865)) + ((!g358) & (g2792) & (!g2846) & (g2853) & (g2865)) + ((!g358) & (g2792) & (g2846) & (!g2853) & (g2865)) + ((g358) & (!g2792) & (!g2846) & (!g2853) & (!g2865)) + ((g358) & (!g2792) & (!g2846) & (g2853) & (!g2865)) + ((g358) & (!g2792) & (!g2846) & (g2853) & (g2865)) + ((g358) & (g2792) & (!g2846) & (!g2853) & (g2865)) + ((g358) & (g2792) & (g2846) & (!g2853) & (!g2865)) + ((g358) & (g2792) & (g2846) & (!g2853) & (g2865)) + ((g358) & (g2792) & (g2846) & (g2853) & (!g2865)) + ((g358) & (g2792) & (g2846) & (g2853) & (g2865)));
	assign g2885 = (((!g390) & (!g433) & (g2794) & (g2845)) + ((!g390) & (g433) & (!g2794) & (g2845)) + ((!g390) & (g433) & (g2794) & (!g2845)) + ((!g390) & (g433) & (g2794) & (g2845)) + ((g390) & (!g433) & (!g2794) & (!g2845)) + ((g390) & (!g433) & (!g2794) & (g2845)) + ((g390) & (!g433) & (g2794) & (!g2845)) + ((g390) & (g433) & (!g2794) & (!g2845)));
	assign g2886 = (((!g2793) & (!g2853) & (!g2865) & (g2885)) + ((!g2793) & (g2853) & (!g2865) & (g2885)) + ((!g2793) & (g2853) & (g2865) & (g2885)) + ((g2793) & (!g2853) & (!g2865) & (!g2885)) + ((g2793) & (!g2853) & (g2865) & (!g2885)) + ((g2793) & (!g2853) & (g2865) & (g2885)) + ((g2793) & (g2853) & (!g2865) & (!g2885)) + ((g2793) & (g2853) & (g2865) & (!g2885)));
	assign g2887 = (((!g433) & (!g2794) & (g2845) & (!g2853) & (!g2865)) + ((!g433) & (!g2794) & (g2845) & (g2853) & (!g2865)) + ((!g433) & (!g2794) & (g2845) & (g2853) & (g2865)) + ((!g433) & (g2794) & (!g2845) & (!g2853) & (!g2865)) + ((!g433) & (g2794) & (!g2845) & (!g2853) & (g2865)) + ((!g433) & (g2794) & (!g2845) & (g2853) & (!g2865)) + ((!g433) & (g2794) & (!g2845) & (g2853) & (g2865)) + ((!g433) & (g2794) & (g2845) & (!g2853) & (g2865)) + ((g433) & (!g2794) & (!g2845) & (!g2853) & (!g2865)) + ((g433) & (!g2794) & (!g2845) & (g2853) & (!g2865)) + ((g433) & (!g2794) & (!g2845) & (g2853) & (g2865)) + ((g433) & (g2794) & (!g2845) & (!g2853) & (g2865)) + ((g433) & (g2794) & (g2845) & (!g2853) & (!g2865)) + ((g433) & (g2794) & (g2845) & (!g2853) & (g2865)) + ((g433) & (g2794) & (g2845) & (g2853) & (!g2865)) + ((g433) & (g2794) & (g2845) & (g2853) & (g2865)));
	assign g2888 = (((!g468) & (!g515) & (g2796) & (g2844)) + ((!g468) & (g515) & (!g2796) & (g2844)) + ((!g468) & (g515) & (g2796) & (!g2844)) + ((!g468) & (g515) & (g2796) & (g2844)) + ((g468) & (!g515) & (!g2796) & (!g2844)) + ((g468) & (!g515) & (!g2796) & (g2844)) + ((g468) & (!g515) & (g2796) & (!g2844)) + ((g468) & (g515) & (!g2796) & (!g2844)));
	assign g2889 = (((!g2795) & (!g2853) & (!g2865) & (g2888)) + ((!g2795) & (g2853) & (!g2865) & (g2888)) + ((!g2795) & (g2853) & (g2865) & (g2888)) + ((g2795) & (!g2853) & (!g2865) & (!g2888)) + ((g2795) & (!g2853) & (g2865) & (!g2888)) + ((g2795) & (!g2853) & (g2865) & (g2888)) + ((g2795) & (g2853) & (!g2865) & (!g2888)) + ((g2795) & (g2853) & (g2865) & (!g2888)));
	assign g2890 = (((!g515) & (!g2796) & (g2844) & (!g2853) & (!g2865)) + ((!g515) & (!g2796) & (g2844) & (g2853) & (!g2865)) + ((!g515) & (!g2796) & (g2844) & (g2853) & (g2865)) + ((!g515) & (g2796) & (!g2844) & (!g2853) & (!g2865)) + ((!g515) & (g2796) & (!g2844) & (!g2853) & (g2865)) + ((!g515) & (g2796) & (!g2844) & (g2853) & (!g2865)) + ((!g515) & (g2796) & (!g2844) & (g2853) & (g2865)) + ((!g515) & (g2796) & (g2844) & (!g2853) & (g2865)) + ((g515) & (!g2796) & (!g2844) & (!g2853) & (!g2865)) + ((g515) & (!g2796) & (!g2844) & (g2853) & (!g2865)) + ((g515) & (!g2796) & (!g2844) & (g2853) & (g2865)) + ((g515) & (g2796) & (!g2844) & (!g2853) & (g2865)) + ((g515) & (g2796) & (g2844) & (!g2853) & (!g2865)) + ((g515) & (g2796) & (g2844) & (!g2853) & (g2865)) + ((g515) & (g2796) & (g2844) & (g2853) & (!g2865)) + ((g515) & (g2796) & (g2844) & (g2853) & (g2865)));
	assign g2891 = (((!g553) & (!g604) & (g2798) & (g2843)) + ((!g553) & (g604) & (!g2798) & (g2843)) + ((!g553) & (g604) & (g2798) & (!g2843)) + ((!g553) & (g604) & (g2798) & (g2843)) + ((g553) & (!g604) & (!g2798) & (!g2843)) + ((g553) & (!g604) & (!g2798) & (g2843)) + ((g553) & (!g604) & (g2798) & (!g2843)) + ((g553) & (g604) & (!g2798) & (!g2843)));
	assign g2892 = (((!g2797) & (!g2853) & (!g2865) & (g2891)) + ((!g2797) & (g2853) & (!g2865) & (g2891)) + ((!g2797) & (g2853) & (g2865) & (g2891)) + ((g2797) & (!g2853) & (!g2865) & (!g2891)) + ((g2797) & (!g2853) & (g2865) & (!g2891)) + ((g2797) & (!g2853) & (g2865) & (g2891)) + ((g2797) & (g2853) & (!g2865) & (!g2891)) + ((g2797) & (g2853) & (g2865) & (!g2891)));
	assign g2893 = (((!g604) & (!g2798) & (g2843) & (!g2853) & (!g2865)) + ((!g604) & (!g2798) & (g2843) & (g2853) & (!g2865)) + ((!g604) & (!g2798) & (g2843) & (g2853) & (g2865)) + ((!g604) & (g2798) & (!g2843) & (!g2853) & (!g2865)) + ((!g604) & (g2798) & (!g2843) & (!g2853) & (g2865)) + ((!g604) & (g2798) & (!g2843) & (g2853) & (!g2865)) + ((!g604) & (g2798) & (!g2843) & (g2853) & (g2865)) + ((!g604) & (g2798) & (g2843) & (!g2853) & (g2865)) + ((g604) & (!g2798) & (!g2843) & (!g2853) & (!g2865)) + ((g604) & (!g2798) & (!g2843) & (g2853) & (!g2865)) + ((g604) & (!g2798) & (!g2843) & (g2853) & (g2865)) + ((g604) & (g2798) & (!g2843) & (!g2853) & (g2865)) + ((g604) & (g2798) & (g2843) & (!g2853) & (!g2865)) + ((g604) & (g2798) & (g2843) & (!g2853) & (g2865)) + ((g604) & (g2798) & (g2843) & (g2853) & (!g2865)) + ((g604) & (g2798) & (g2843) & (g2853) & (g2865)));
	assign g2894 = (((!g645) & (!g700) & (g2800) & (g2842)) + ((!g645) & (g700) & (!g2800) & (g2842)) + ((!g645) & (g700) & (g2800) & (!g2842)) + ((!g645) & (g700) & (g2800) & (g2842)) + ((g645) & (!g700) & (!g2800) & (!g2842)) + ((g645) & (!g700) & (!g2800) & (g2842)) + ((g645) & (!g700) & (g2800) & (!g2842)) + ((g645) & (g700) & (!g2800) & (!g2842)));
	assign g2895 = (((!g2799) & (!g2853) & (!g2865) & (g2894)) + ((!g2799) & (g2853) & (!g2865) & (g2894)) + ((!g2799) & (g2853) & (g2865) & (g2894)) + ((g2799) & (!g2853) & (!g2865) & (!g2894)) + ((g2799) & (!g2853) & (g2865) & (!g2894)) + ((g2799) & (!g2853) & (g2865) & (g2894)) + ((g2799) & (g2853) & (!g2865) & (!g2894)) + ((g2799) & (g2853) & (g2865) & (!g2894)));
	assign g2896 = (((!g700) & (!g2800) & (g2842) & (!g2853) & (!g2865)) + ((!g700) & (!g2800) & (g2842) & (g2853) & (!g2865)) + ((!g700) & (!g2800) & (g2842) & (g2853) & (g2865)) + ((!g700) & (g2800) & (!g2842) & (!g2853) & (!g2865)) + ((!g700) & (g2800) & (!g2842) & (!g2853) & (g2865)) + ((!g700) & (g2800) & (!g2842) & (g2853) & (!g2865)) + ((!g700) & (g2800) & (!g2842) & (g2853) & (g2865)) + ((!g700) & (g2800) & (g2842) & (!g2853) & (g2865)) + ((g700) & (!g2800) & (!g2842) & (!g2853) & (!g2865)) + ((g700) & (!g2800) & (!g2842) & (g2853) & (!g2865)) + ((g700) & (!g2800) & (!g2842) & (g2853) & (g2865)) + ((g700) & (g2800) & (!g2842) & (!g2853) & (g2865)) + ((g700) & (g2800) & (g2842) & (!g2853) & (!g2865)) + ((g700) & (g2800) & (g2842) & (!g2853) & (g2865)) + ((g700) & (g2800) & (g2842) & (g2853) & (!g2865)) + ((g700) & (g2800) & (g2842) & (g2853) & (g2865)));
	assign g2897 = (((!g744) & (!g803) & (g2802) & (g2841)) + ((!g744) & (g803) & (!g2802) & (g2841)) + ((!g744) & (g803) & (g2802) & (!g2841)) + ((!g744) & (g803) & (g2802) & (g2841)) + ((g744) & (!g803) & (!g2802) & (!g2841)) + ((g744) & (!g803) & (!g2802) & (g2841)) + ((g744) & (!g803) & (g2802) & (!g2841)) + ((g744) & (g803) & (!g2802) & (!g2841)));
	assign g2898 = (((!g2801) & (!g2853) & (!g2865) & (g2897)) + ((!g2801) & (g2853) & (!g2865) & (g2897)) + ((!g2801) & (g2853) & (g2865) & (g2897)) + ((g2801) & (!g2853) & (!g2865) & (!g2897)) + ((g2801) & (!g2853) & (g2865) & (!g2897)) + ((g2801) & (!g2853) & (g2865) & (g2897)) + ((g2801) & (g2853) & (!g2865) & (!g2897)) + ((g2801) & (g2853) & (g2865) & (!g2897)));
	assign g2899 = (((!g803) & (!g2802) & (g2841) & (!g2853) & (!g2865)) + ((!g803) & (!g2802) & (g2841) & (g2853) & (!g2865)) + ((!g803) & (!g2802) & (g2841) & (g2853) & (g2865)) + ((!g803) & (g2802) & (!g2841) & (!g2853) & (!g2865)) + ((!g803) & (g2802) & (!g2841) & (!g2853) & (g2865)) + ((!g803) & (g2802) & (!g2841) & (g2853) & (!g2865)) + ((!g803) & (g2802) & (!g2841) & (g2853) & (g2865)) + ((!g803) & (g2802) & (g2841) & (!g2853) & (g2865)) + ((g803) & (!g2802) & (!g2841) & (!g2853) & (!g2865)) + ((g803) & (!g2802) & (!g2841) & (g2853) & (!g2865)) + ((g803) & (!g2802) & (!g2841) & (g2853) & (g2865)) + ((g803) & (g2802) & (!g2841) & (!g2853) & (g2865)) + ((g803) & (g2802) & (g2841) & (!g2853) & (!g2865)) + ((g803) & (g2802) & (g2841) & (!g2853) & (g2865)) + ((g803) & (g2802) & (g2841) & (g2853) & (!g2865)) + ((g803) & (g2802) & (g2841) & (g2853) & (g2865)));
	assign g2900 = (((!g851) & (!g914) & (g2804) & (g2840)) + ((!g851) & (g914) & (!g2804) & (g2840)) + ((!g851) & (g914) & (g2804) & (!g2840)) + ((!g851) & (g914) & (g2804) & (g2840)) + ((g851) & (!g914) & (!g2804) & (!g2840)) + ((g851) & (!g914) & (!g2804) & (g2840)) + ((g851) & (!g914) & (g2804) & (!g2840)) + ((g851) & (g914) & (!g2804) & (!g2840)));
	assign g2901 = (((!g2803) & (!g2853) & (!g2865) & (g2900)) + ((!g2803) & (g2853) & (!g2865) & (g2900)) + ((!g2803) & (g2853) & (g2865) & (g2900)) + ((g2803) & (!g2853) & (!g2865) & (!g2900)) + ((g2803) & (!g2853) & (g2865) & (!g2900)) + ((g2803) & (!g2853) & (g2865) & (g2900)) + ((g2803) & (g2853) & (!g2865) & (!g2900)) + ((g2803) & (g2853) & (g2865) & (!g2900)));
	assign g2902 = (((!g914) & (!g2804) & (g2840) & (!g2853) & (!g2865)) + ((!g914) & (!g2804) & (g2840) & (g2853) & (!g2865)) + ((!g914) & (!g2804) & (g2840) & (g2853) & (g2865)) + ((!g914) & (g2804) & (!g2840) & (!g2853) & (!g2865)) + ((!g914) & (g2804) & (!g2840) & (!g2853) & (g2865)) + ((!g914) & (g2804) & (!g2840) & (g2853) & (!g2865)) + ((!g914) & (g2804) & (!g2840) & (g2853) & (g2865)) + ((!g914) & (g2804) & (g2840) & (!g2853) & (g2865)) + ((g914) & (!g2804) & (!g2840) & (!g2853) & (!g2865)) + ((g914) & (!g2804) & (!g2840) & (g2853) & (!g2865)) + ((g914) & (!g2804) & (!g2840) & (g2853) & (g2865)) + ((g914) & (g2804) & (!g2840) & (!g2853) & (g2865)) + ((g914) & (g2804) & (g2840) & (!g2853) & (!g2865)) + ((g914) & (g2804) & (g2840) & (!g2853) & (g2865)) + ((g914) & (g2804) & (g2840) & (g2853) & (!g2865)) + ((g914) & (g2804) & (g2840) & (g2853) & (g2865)));
	assign g2903 = (((!g1032) & (!g1030) & (g2806) & (g2839)) + ((!g1032) & (g1030) & (!g2806) & (g2839)) + ((!g1032) & (g1030) & (g2806) & (!g2839)) + ((!g1032) & (g1030) & (g2806) & (g2839)) + ((g1032) & (!g1030) & (!g2806) & (!g2839)) + ((g1032) & (!g1030) & (!g2806) & (g2839)) + ((g1032) & (!g1030) & (g2806) & (!g2839)) + ((g1032) & (g1030) & (!g2806) & (!g2839)));
	assign g2904 = (((!g2805) & (!g2853) & (!g2865) & (g2903)) + ((!g2805) & (g2853) & (!g2865) & (g2903)) + ((!g2805) & (g2853) & (g2865) & (g2903)) + ((g2805) & (!g2853) & (!g2865) & (!g2903)) + ((g2805) & (!g2853) & (g2865) & (!g2903)) + ((g2805) & (!g2853) & (g2865) & (g2903)) + ((g2805) & (g2853) & (!g2865) & (!g2903)) + ((g2805) & (g2853) & (g2865) & (!g2903)));
	assign g2905 = (((!g1030) & (!g2806) & (g2839) & (!g2853) & (!g2865)) + ((!g1030) & (!g2806) & (g2839) & (g2853) & (!g2865)) + ((!g1030) & (!g2806) & (g2839) & (g2853) & (g2865)) + ((!g1030) & (g2806) & (!g2839) & (!g2853) & (!g2865)) + ((!g1030) & (g2806) & (!g2839) & (!g2853) & (g2865)) + ((!g1030) & (g2806) & (!g2839) & (g2853) & (!g2865)) + ((!g1030) & (g2806) & (!g2839) & (g2853) & (g2865)) + ((!g1030) & (g2806) & (g2839) & (!g2853) & (g2865)) + ((g1030) & (!g2806) & (!g2839) & (!g2853) & (!g2865)) + ((g1030) & (!g2806) & (!g2839) & (g2853) & (!g2865)) + ((g1030) & (!g2806) & (!g2839) & (g2853) & (g2865)) + ((g1030) & (g2806) & (!g2839) & (!g2853) & (g2865)) + ((g1030) & (g2806) & (g2839) & (!g2853) & (!g2865)) + ((g1030) & (g2806) & (g2839) & (!g2853) & (g2865)) + ((g1030) & (g2806) & (g2839) & (g2853) & (!g2865)) + ((g1030) & (g2806) & (g2839) & (g2853) & (g2865)));
	assign g2906 = (((!g1160) & (!g1154) & (g2808) & (g2838)) + ((!g1160) & (g1154) & (!g2808) & (g2838)) + ((!g1160) & (g1154) & (g2808) & (!g2838)) + ((!g1160) & (g1154) & (g2808) & (g2838)) + ((g1160) & (!g1154) & (!g2808) & (!g2838)) + ((g1160) & (!g1154) & (!g2808) & (g2838)) + ((g1160) & (!g1154) & (g2808) & (!g2838)) + ((g1160) & (g1154) & (!g2808) & (!g2838)));
	assign g2907 = (((!g2807) & (!g2853) & (!g2865) & (g2906)) + ((!g2807) & (g2853) & (!g2865) & (g2906)) + ((!g2807) & (g2853) & (g2865) & (g2906)) + ((g2807) & (!g2853) & (!g2865) & (!g2906)) + ((g2807) & (!g2853) & (g2865) & (!g2906)) + ((g2807) & (!g2853) & (g2865) & (g2906)) + ((g2807) & (g2853) & (!g2865) & (!g2906)) + ((g2807) & (g2853) & (g2865) & (!g2906)));
	assign g2908 = (((!g1154) & (!g2808) & (g2838) & (!g2853) & (!g2865)) + ((!g1154) & (!g2808) & (g2838) & (g2853) & (!g2865)) + ((!g1154) & (!g2808) & (g2838) & (g2853) & (g2865)) + ((!g1154) & (g2808) & (!g2838) & (!g2853) & (!g2865)) + ((!g1154) & (g2808) & (!g2838) & (!g2853) & (g2865)) + ((!g1154) & (g2808) & (!g2838) & (g2853) & (!g2865)) + ((!g1154) & (g2808) & (!g2838) & (g2853) & (g2865)) + ((!g1154) & (g2808) & (g2838) & (!g2853) & (g2865)) + ((g1154) & (!g2808) & (!g2838) & (!g2853) & (!g2865)) + ((g1154) & (!g2808) & (!g2838) & (g2853) & (!g2865)) + ((g1154) & (!g2808) & (!g2838) & (g2853) & (g2865)) + ((g1154) & (g2808) & (!g2838) & (!g2853) & (g2865)) + ((g1154) & (g2808) & (g2838) & (!g2853) & (!g2865)) + ((g1154) & (g2808) & (g2838) & (!g2853) & (g2865)) + ((g1154) & (g2808) & (g2838) & (g2853) & (!g2865)) + ((g1154) & (g2808) & (g2838) & (g2853) & (g2865)));
	assign g2909 = (((!g1295) & (!g1285) & (g2810) & (g2837)) + ((!g1295) & (g1285) & (!g2810) & (g2837)) + ((!g1295) & (g1285) & (g2810) & (!g2837)) + ((!g1295) & (g1285) & (g2810) & (g2837)) + ((g1295) & (!g1285) & (!g2810) & (!g2837)) + ((g1295) & (!g1285) & (!g2810) & (g2837)) + ((g1295) & (!g1285) & (g2810) & (!g2837)) + ((g1295) & (g1285) & (!g2810) & (!g2837)));
	assign g2910 = (((!g2809) & (!g2853) & (!g2865) & (g2909)) + ((!g2809) & (g2853) & (!g2865) & (g2909)) + ((!g2809) & (g2853) & (g2865) & (g2909)) + ((g2809) & (!g2853) & (!g2865) & (!g2909)) + ((g2809) & (!g2853) & (g2865) & (!g2909)) + ((g2809) & (!g2853) & (g2865) & (g2909)) + ((g2809) & (g2853) & (!g2865) & (!g2909)) + ((g2809) & (g2853) & (g2865) & (!g2909)));
	assign g2911 = (((!g1285) & (!g2810) & (g2837) & (!g2853) & (!g2865)) + ((!g1285) & (!g2810) & (g2837) & (g2853) & (!g2865)) + ((!g1285) & (!g2810) & (g2837) & (g2853) & (g2865)) + ((!g1285) & (g2810) & (!g2837) & (!g2853) & (!g2865)) + ((!g1285) & (g2810) & (!g2837) & (!g2853) & (g2865)) + ((!g1285) & (g2810) & (!g2837) & (g2853) & (!g2865)) + ((!g1285) & (g2810) & (!g2837) & (g2853) & (g2865)) + ((!g1285) & (g2810) & (g2837) & (!g2853) & (g2865)) + ((g1285) & (!g2810) & (!g2837) & (!g2853) & (!g2865)) + ((g1285) & (!g2810) & (!g2837) & (g2853) & (!g2865)) + ((g1285) & (!g2810) & (!g2837) & (g2853) & (g2865)) + ((g1285) & (g2810) & (!g2837) & (!g2853) & (g2865)) + ((g1285) & (g2810) & (g2837) & (!g2853) & (!g2865)) + ((g1285) & (g2810) & (g2837) & (!g2853) & (g2865)) + ((g1285) & (g2810) & (g2837) & (g2853) & (!g2865)) + ((g1285) & (g2810) & (g2837) & (g2853) & (g2865)));
	assign g2912 = (((!g1437) & (!g1423) & (g2812) & (g2836)) + ((!g1437) & (g1423) & (!g2812) & (g2836)) + ((!g1437) & (g1423) & (g2812) & (!g2836)) + ((!g1437) & (g1423) & (g2812) & (g2836)) + ((g1437) & (!g1423) & (!g2812) & (!g2836)) + ((g1437) & (!g1423) & (!g2812) & (g2836)) + ((g1437) & (!g1423) & (g2812) & (!g2836)) + ((g1437) & (g1423) & (!g2812) & (!g2836)));
	assign g2913 = (((!g2811) & (!g2853) & (!g2865) & (g2912)) + ((!g2811) & (g2853) & (!g2865) & (g2912)) + ((!g2811) & (g2853) & (g2865) & (g2912)) + ((g2811) & (!g2853) & (!g2865) & (!g2912)) + ((g2811) & (!g2853) & (g2865) & (!g2912)) + ((g2811) & (!g2853) & (g2865) & (g2912)) + ((g2811) & (g2853) & (!g2865) & (!g2912)) + ((g2811) & (g2853) & (g2865) & (!g2912)));
	assign g2914 = (((!g1423) & (!g2812) & (g2836) & (!g2853) & (!g2865)) + ((!g1423) & (!g2812) & (g2836) & (g2853) & (!g2865)) + ((!g1423) & (!g2812) & (g2836) & (g2853) & (g2865)) + ((!g1423) & (g2812) & (!g2836) & (!g2853) & (!g2865)) + ((!g1423) & (g2812) & (!g2836) & (!g2853) & (g2865)) + ((!g1423) & (g2812) & (!g2836) & (g2853) & (!g2865)) + ((!g1423) & (g2812) & (!g2836) & (g2853) & (g2865)) + ((!g1423) & (g2812) & (g2836) & (!g2853) & (g2865)) + ((g1423) & (!g2812) & (!g2836) & (!g2853) & (!g2865)) + ((g1423) & (!g2812) & (!g2836) & (g2853) & (!g2865)) + ((g1423) & (!g2812) & (!g2836) & (g2853) & (g2865)) + ((g1423) & (g2812) & (!g2836) & (!g2853) & (g2865)) + ((g1423) & (g2812) & (g2836) & (!g2853) & (!g2865)) + ((g1423) & (g2812) & (g2836) & (!g2853) & (g2865)) + ((g1423) & (g2812) & (g2836) & (g2853) & (!g2865)) + ((g1423) & (g2812) & (g2836) & (g2853) & (g2865)));
	assign g2915 = (((!g1586) & (!g1568) & (g2814) & (g2835)) + ((!g1586) & (g1568) & (!g2814) & (g2835)) + ((!g1586) & (g1568) & (g2814) & (!g2835)) + ((!g1586) & (g1568) & (g2814) & (g2835)) + ((g1586) & (!g1568) & (!g2814) & (!g2835)) + ((g1586) & (!g1568) & (!g2814) & (g2835)) + ((g1586) & (!g1568) & (g2814) & (!g2835)) + ((g1586) & (g1568) & (!g2814) & (!g2835)));
	assign g2916 = (((!g2813) & (!g2853) & (!g2865) & (g2915)) + ((!g2813) & (g2853) & (!g2865) & (g2915)) + ((!g2813) & (g2853) & (g2865) & (g2915)) + ((g2813) & (!g2853) & (!g2865) & (!g2915)) + ((g2813) & (!g2853) & (g2865) & (!g2915)) + ((g2813) & (!g2853) & (g2865) & (g2915)) + ((g2813) & (g2853) & (!g2865) & (!g2915)) + ((g2813) & (g2853) & (g2865) & (!g2915)));
	assign g2917 = (((!g1568) & (!g2814) & (g2835) & (!g2853) & (!g2865)) + ((!g1568) & (!g2814) & (g2835) & (g2853) & (!g2865)) + ((!g1568) & (!g2814) & (g2835) & (g2853) & (g2865)) + ((!g1568) & (g2814) & (!g2835) & (!g2853) & (!g2865)) + ((!g1568) & (g2814) & (!g2835) & (!g2853) & (g2865)) + ((!g1568) & (g2814) & (!g2835) & (g2853) & (!g2865)) + ((!g1568) & (g2814) & (!g2835) & (g2853) & (g2865)) + ((!g1568) & (g2814) & (g2835) & (!g2853) & (g2865)) + ((g1568) & (!g2814) & (!g2835) & (!g2853) & (!g2865)) + ((g1568) & (!g2814) & (!g2835) & (g2853) & (!g2865)) + ((g1568) & (!g2814) & (!g2835) & (g2853) & (g2865)) + ((g1568) & (g2814) & (!g2835) & (!g2853) & (g2865)) + ((g1568) & (g2814) & (g2835) & (!g2853) & (!g2865)) + ((g1568) & (g2814) & (g2835) & (!g2853) & (g2865)) + ((g1568) & (g2814) & (g2835) & (g2853) & (!g2865)) + ((g1568) & (g2814) & (g2835) & (g2853) & (g2865)));
	assign g2918 = (((!g1742) & (!g1720) & (g2816) & (g2834)) + ((!g1742) & (g1720) & (!g2816) & (g2834)) + ((!g1742) & (g1720) & (g2816) & (!g2834)) + ((!g1742) & (g1720) & (g2816) & (g2834)) + ((g1742) & (!g1720) & (!g2816) & (!g2834)) + ((g1742) & (!g1720) & (!g2816) & (g2834)) + ((g1742) & (!g1720) & (g2816) & (!g2834)) + ((g1742) & (g1720) & (!g2816) & (!g2834)));
	assign g2919 = (((!g2815) & (!g2853) & (!g2865) & (g2918)) + ((!g2815) & (g2853) & (!g2865) & (g2918)) + ((!g2815) & (g2853) & (g2865) & (g2918)) + ((g2815) & (!g2853) & (!g2865) & (!g2918)) + ((g2815) & (!g2853) & (g2865) & (!g2918)) + ((g2815) & (!g2853) & (g2865) & (g2918)) + ((g2815) & (g2853) & (!g2865) & (!g2918)) + ((g2815) & (g2853) & (g2865) & (!g2918)));
	assign g2920 = (((!g1720) & (!g2816) & (g2834) & (!g2853) & (!g2865)) + ((!g1720) & (!g2816) & (g2834) & (g2853) & (!g2865)) + ((!g1720) & (!g2816) & (g2834) & (g2853) & (g2865)) + ((!g1720) & (g2816) & (!g2834) & (!g2853) & (!g2865)) + ((!g1720) & (g2816) & (!g2834) & (!g2853) & (g2865)) + ((!g1720) & (g2816) & (!g2834) & (g2853) & (!g2865)) + ((!g1720) & (g2816) & (!g2834) & (g2853) & (g2865)) + ((!g1720) & (g2816) & (g2834) & (!g2853) & (g2865)) + ((g1720) & (!g2816) & (!g2834) & (!g2853) & (!g2865)) + ((g1720) & (!g2816) & (!g2834) & (g2853) & (!g2865)) + ((g1720) & (!g2816) & (!g2834) & (g2853) & (g2865)) + ((g1720) & (g2816) & (!g2834) & (!g2853) & (g2865)) + ((g1720) & (g2816) & (g2834) & (!g2853) & (!g2865)) + ((g1720) & (g2816) & (g2834) & (!g2853) & (g2865)) + ((g1720) & (g2816) & (g2834) & (g2853) & (!g2865)) + ((g1720) & (g2816) & (g2834) & (g2853) & (g2865)));
	assign g2921 = (((!g1905) & (!g1879) & (g2818) & (g2833)) + ((!g1905) & (g1879) & (!g2818) & (g2833)) + ((!g1905) & (g1879) & (g2818) & (!g2833)) + ((!g1905) & (g1879) & (g2818) & (g2833)) + ((g1905) & (!g1879) & (!g2818) & (!g2833)) + ((g1905) & (!g1879) & (!g2818) & (g2833)) + ((g1905) & (!g1879) & (g2818) & (!g2833)) + ((g1905) & (g1879) & (!g2818) & (!g2833)));
	assign g2922 = (((!g2817) & (!g2853) & (!g2865) & (g2921)) + ((!g2817) & (g2853) & (!g2865) & (g2921)) + ((!g2817) & (g2853) & (g2865) & (g2921)) + ((g2817) & (!g2853) & (!g2865) & (!g2921)) + ((g2817) & (!g2853) & (g2865) & (!g2921)) + ((g2817) & (!g2853) & (g2865) & (g2921)) + ((g2817) & (g2853) & (!g2865) & (!g2921)) + ((g2817) & (g2853) & (g2865) & (!g2921)));
	assign g2923 = (((!g1879) & (!g2818) & (g2833) & (!g2853) & (!g2865)) + ((!g1879) & (!g2818) & (g2833) & (g2853) & (!g2865)) + ((!g1879) & (!g2818) & (g2833) & (g2853) & (g2865)) + ((!g1879) & (g2818) & (!g2833) & (!g2853) & (!g2865)) + ((!g1879) & (g2818) & (!g2833) & (!g2853) & (g2865)) + ((!g1879) & (g2818) & (!g2833) & (g2853) & (!g2865)) + ((!g1879) & (g2818) & (!g2833) & (g2853) & (g2865)) + ((!g1879) & (g2818) & (g2833) & (!g2853) & (g2865)) + ((g1879) & (!g2818) & (!g2833) & (!g2853) & (!g2865)) + ((g1879) & (!g2818) & (!g2833) & (g2853) & (!g2865)) + ((g1879) & (!g2818) & (!g2833) & (g2853) & (g2865)) + ((g1879) & (g2818) & (!g2833) & (!g2853) & (g2865)) + ((g1879) & (g2818) & (g2833) & (!g2853) & (!g2865)) + ((g1879) & (g2818) & (g2833) & (!g2853) & (g2865)) + ((g1879) & (g2818) & (g2833) & (g2853) & (!g2865)) + ((g1879) & (g2818) & (g2833) & (g2853) & (g2865)));
	assign g2924 = (((!g2075) & (!g2045) & (g2820) & (g2832)) + ((!g2075) & (g2045) & (!g2820) & (g2832)) + ((!g2075) & (g2045) & (g2820) & (!g2832)) + ((!g2075) & (g2045) & (g2820) & (g2832)) + ((g2075) & (!g2045) & (!g2820) & (!g2832)) + ((g2075) & (!g2045) & (!g2820) & (g2832)) + ((g2075) & (!g2045) & (g2820) & (!g2832)) + ((g2075) & (g2045) & (!g2820) & (!g2832)));
	assign g2925 = (((!g2819) & (!g2853) & (!g2865) & (g2924)) + ((!g2819) & (g2853) & (!g2865) & (g2924)) + ((!g2819) & (g2853) & (g2865) & (g2924)) + ((g2819) & (!g2853) & (!g2865) & (!g2924)) + ((g2819) & (!g2853) & (g2865) & (!g2924)) + ((g2819) & (!g2853) & (g2865) & (g2924)) + ((g2819) & (g2853) & (!g2865) & (!g2924)) + ((g2819) & (g2853) & (g2865) & (!g2924)));
	assign g2926 = (((!g2045) & (!g2820) & (g2832) & (!g2853) & (!g2865)) + ((!g2045) & (!g2820) & (g2832) & (g2853) & (!g2865)) + ((!g2045) & (!g2820) & (g2832) & (g2853) & (g2865)) + ((!g2045) & (g2820) & (!g2832) & (!g2853) & (!g2865)) + ((!g2045) & (g2820) & (!g2832) & (!g2853) & (g2865)) + ((!g2045) & (g2820) & (!g2832) & (g2853) & (!g2865)) + ((!g2045) & (g2820) & (!g2832) & (g2853) & (g2865)) + ((!g2045) & (g2820) & (g2832) & (!g2853) & (g2865)) + ((g2045) & (!g2820) & (!g2832) & (!g2853) & (!g2865)) + ((g2045) & (!g2820) & (!g2832) & (g2853) & (!g2865)) + ((g2045) & (!g2820) & (!g2832) & (g2853) & (g2865)) + ((g2045) & (g2820) & (!g2832) & (!g2853) & (g2865)) + ((g2045) & (g2820) & (g2832) & (!g2853) & (!g2865)) + ((g2045) & (g2820) & (g2832) & (!g2853) & (g2865)) + ((g2045) & (g2820) & (g2832) & (g2853) & (!g2865)) + ((g2045) & (g2820) & (g2832) & (g2853) & (g2865)));
	assign g2927 = (((!g2252) & (!g2218) & (g2822) & (g2831)) + ((!g2252) & (g2218) & (!g2822) & (g2831)) + ((!g2252) & (g2218) & (g2822) & (!g2831)) + ((!g2252) & (g2218) & (g2822) & (g2831)) + ((g2252) & (!g2218) & (!g2822) & (!g2831)) + ((g2252) & (!g2218) & (!g2822) & (g2831)) + ((g2252) & (!g2218) & (g2822) & (!g2831)) + ((g2252) & (g2218) & (!g2822) & (!g2831)));
	assign g2928 = (((!g2821) & (!g2853) & (!g2865) & (g2927)) + ((!g2821) & (g2853) & (!g2865) & (g2927)) + ((!g2821) & (g2853) & (g2865) & (g2927)) + ((g2821) & (!g2853) & (!g2865) & (!g2927)) + ((g2821) & (!g2853) & (g2865) & (!g2927)) + ((g2821) & (!g2853) & (g2865) & (g2927)) + ((g2821) & (g2853) & (!g2865) & (!g2927)) + ((g2821) & (g2853) & (g2865) & (!g2927)));
	assign g2929 = (((!g2218) & (!g2822) & (g2831) & (!g2853) & (!g2865)) + ((!g2218) & (!g2822) & (g2831) & (g2853) & (!g2865)) + ((!g2218) & (!g2822) & (g2831) & (g2853) & (g2865)) + ((!g2218) & (g2822) & (!g2831) & (!g2853) & (!g2865)) + ((!g2218) & (g2822) & (!g2831) & (!g2853) & (g2865)) + ((!g2218) & (g2822) & (!g2831) & (g2853) & (!g2865)) + ((!g2218) & (g2822) & (!g2831) & (g2853) & (g2865)) + ((!g2218) & (g2822) & (g2831) & (!g2853) & (g2865)) + ((g2218) & (!g2822) & (!g2831) & (!g2853) & (!g2865)) + ((g2218) & (!g2822) & (!g2831) & (g2853) & (!g2865)) + ((g2218) & (!g2822) & (!g2831) & (g2853) & (g2865)) + ((g2218) & (g2822) & (!g2831) & (!g2853) & (g2865)) + ((g2218) & (g2822) & (g2831) & (!g2853) & (!g2865)) + ((g2218) & (g2822) & (g2831) & (!g2853) & (g2865)) + ((g2218) & (g2822) & (g2831) & (g2853) & (!g2865)) + ((g2218) & (g2822) & (g2831) & (g2853) & (g2865)));
	assign g2930 = (((!g2436) & (!g2398) & (g2824) & (g2830)) + ((!g2436) & (g2398) & (!g2824) & (g2830)) + ((!g2436) & (g2398) & (g2824) & (!g2830)) + ((!g2436) & (g2398) & (g2824) & (g2830)) + ((g2436) & (!g2398) & (!g2824) & (!g2830)) + ((g2436) & (!g2398) & (!g2824) & (g2830)) + ((g2436) & (!g2398) & (g2824) & (!g2830)) + ((g2436) & (g2398) & (!g2824) & (!g2830)));
	assign g2931 = (((!g2823) & (!g2853) & (!g2865) & (g2930)) + ((!g2823) & (g2853) & (!g2865) & (g2930)) + ((!g2823) & (g2853) & (g2865) & (g2930)) + ((g2823) & (!g2853) & (!g2865) & (!g2930)) + ((g2823) & (!g2853) & (g2865) & (!g2930)) + ((g2823) & (!g2853) & (g2865) & (g2930)) + ((g2823) & (g2853) & (!g2865) & (!g2930)) + ((g2823) & (g2853) & (g2865) & (!g2930)));
	assign g2932 = (((!g2398) & (!g2824) & (g2830) & (!g2853) & (!g2865)) + ((!g2398) & (!g2824) & (g2830) & (g2853) & (!g2865)) + ((!g2398) & (!g2824) & (g2830) & (g2853) & (g2865)) + ((!g2398) & (g2824) & (!g2830) & (!g2853) & (!g2865)) + ((!g2398) & (g2824) & (!g2830) & (!g2853) & (g2865)) + ((!g2398) & (g2824) & (!g2830) & (g2853) & (!g2865)) + ((!g2398) & (g2824) & (!g2830) & (g2853) & (g2865)) + ((!g2398) & (g2824) & (g2830) & (!g2853) & (g2865)) + ((g2398) & (!g2824) & (!g2830) & (!g2853) & (!g2865)) + ((g2398) & (!g2824) & (!g2830) & (g2853) & (!g2865)) + ((g2398) & (!g2824) & (!g2830) & (g2853) & (g2865)) + ((g2398) & (g2824) & (!g2830) & (!g2853) & (g2865)) + ((g2398) & (g2824) & (g2830) & (!g2853) & (!g2865)) + ((g2398) & (g2824) & (g2830) & (!g2853) & (g2865)) + ((g2398) & (g2824) & (g2830) & (g2853) & (!g2865)) + ((g2398) & (g2824) & (g2830) & (g2853) & (g2865)));
	assign g2933 = (((!g2627) & (!g2585) & (g2827) & (g2829)) + ((!g2627) & (g2585) & (!g2827) & (g2829)) + ((!g2627) & (g2585) & (g2827) & (!g2829)) + ((!g2627) & (g2585) & (g2827) & (g2829)) + ((g2627) & (!g2585) & (!g2827) & (!g2829)) + ((g2627) & (!g2585) & (!g2827) & (g2829)) + ((g2627) & (!g2585) & (g2827) & (!g2829)) + ((g2627) & (g2585) & (!g2827) & (!g2829)));
	assign g2934 = (((!g2826) & (!g2853) & (!g2865) & (g2933)) + ((!g2826) & (g2853) & (!g2865) & (g2933)) + ((!g2826) & (g2853) & (g2865) & (g2933)) + ((g2826) & (!g2853) & (!g2865) & (!g2933)) + ((g2826) & (!g2853) & (g2865) & (!g2933)) + ((g2826) & (!g2853) & (g2865) & (g2933)) + ((g2826) & (g2853) & (!g2865) & (!g2933)) + ((g2826) & (g2853) & (g2865) & (!g2933)));
	assign g2935 = (((!g2585) & (!g2827) & (g2829) & (!g2853) & (!g2865)) + ((!g2585) & (!g2827) & (g2829) & (g2853) & (!g2865)) + ((!g2585) & (!g2827) & (g2829) & (g2853) & (g2865)) + ((!g2585) & (g2827) & (!g2829) & (!g2853) & (!g2865)) + ((!g2585) & (g2827) & (!g2829) & (!g2853) & (g2865)) + ((!g2585) & (g2827) & (!g2829) & (g2853) & (!g2865)) + ((!g2585) & (g2827) & (!g2829) & (g2853) & (g2865)) + ((!g2585) & (g2827) & (g2829) & (!g2853) & (g2865)) + ((g2585) & (!g2827) & (!g2829) & (!g2853) & (!g2865)) + ((g2585) & (!g2827) & (!g2829) & (g2853) & (!g2865)) + ((g2585) & (!g2827) & (!g2829) & (g2853) & (g2865)) + ((g2585) & (g2827) & (!g2829) & (!g2853) & (g2865)) + ((g2585) & (g2827) & (g2829) & (!g2853) & (!g2865)) + ((g2585) & (g2827) & (g2829) & (!g2853) & (g2865)) + ((g2585) & (g2827) & (g2829) & (g2853) & (!g2865)) + ((g2585) & (g2827) & (g2829) & (g2853) & (g2865)));
	assign g2936 = (((!g2825) & (!ax16x) & (!g2779) & (g2828)) + ((!g2825) & (!ax16x) & (g2779) & (g2828)) + ((!g2825) & (ax16x) & (!g2779) & (!g2828)) + ((!g2825) & (ax16x) & (!g2779) & (g2828)) + ((g2825) & (!ax16x) & (!g2779) & (!g2828)) + ((g2825) & (!ax16x) & (g2779) & (!g2828)) + ((g2825) & (ax16x) & (g2779) & (!g2828)) + ((g2825) & (ax16x) & (g2779) & (g2828)));
	assign g2937 = (((!ax16x) & (!ax17x) & (!g2779) & (!g2853) & (!g2865) & (g2936)) + ((!ax16x) & (!ax17x) & (!g2779) & (!g2853) & (g2865) & (!g2936)) + ((!ax16x) & (!ax17x) & (!g2779) & (!g2853) & (g2865) & (g2936)) + ((!ax16x) & (!ax17x) & (!g2779) & (g2853) & (!g2865) & (g2936)) + ((!ax16x) & (!ax17x) & (!g2779) & (g2853) & (g2865) & (g2936)) + ((!ax16x) & (!ax17x) & (g2779) & (!g2853) & (!g2865) & (!g2936)) + ((!ax16x) & (!ax17x) & (g2779) & (g2853) & (!g2865) & (!g2936)) + ((!ax16x) & (!ax17x) & (g2779) & (g2853) & (g2865) & (!g2936)) + ((!ax16x) & (ax17x) & (!g2779) & (!g2853) & (!g2865) & (!g2936)) + ((!ax16x) & (ax17x) & (!g2779) & (g2853) & (!g2865) & (!g2936)) + ((!ax16x) & (ax17x) & (!g2779) & (g2853) & (g2865) & (!g2936)) + ((!ax16x) & (ax17x) & (g2779) & (!g2853) & (!g2865) & (g2936)) + ((!ax16x) & (ax17x) & (g2779) & (!g2853) & (g2865) & (!g2936)) + ((!ax16x) & (ax17x) & (g2779) & (!g2853) & (g2865) & (g2936)) + ((!ax16x) & (ax17x) & (g2779) & (g2853) & (!g2865) & (g2936)) + ((!ax16x) & (ax17x) & (g2779) & (g2853) & (g2865) & (g2936)) + ((ax16x) & (!ax17x) & (!g2779) & (!g2853) & (!g2865) & (!g2936)) + ((ax16x) & (!ax17x) & (!g2779) & (g2853) & (!g2865) & (!g2936)) + ((ax16x) & (!ax17x) & (!g2779) & (g2853) & (g2865) & (!g2936)) + ((ax16x) & (!ax17x) & (g2779) & (!g2853) & (!g2865) & (!g2936)) + ((ax16x) & (!ax17x) & (g2779) & (g2853) & (!g2865) & (!g2936)) + ((ax16x) & (!ax17x) & (g2779) & (g2853) & (g2865) & (!g2936)) + ((ax16x) & (ax17x) & (!g2779) & (!g2853) & (!g2865) & (g2936)) + ((ax16x) & (ax17x) & (!g2779) & (!g2853) & (g2865) & (!g2936)) + ((ax16x) & (ax17x) & (!g2779) & (!g2853) & (g2865) & (g2936)) + ((ax16x) & (ax17x) & (!g2779) & (g2853) & (!g2865) & (g2936)) + ((ax16x) & (ax17x) & (!g2779) & (g2853) & (g2865) & (g2936)) + ((ax16x) & (ax17x) & (g2779) & (!g2853) & (!g2865) & (g2936)) + ((ax16x) & (ax17x) & (g2779) & (!g2853) & (g2865) & (!g2936)) + ((ax16x) & (ax17x) & (g2779) & (!g2853) & (g2865) & (g2936)) + ((ax16x) & (ax17x) & (g2779) & (g2853) & (!g2865) & (g2936)) + ((ax16x) & (ax17x) & (g2779) & (g2853) & (g2865) & (g2936)));
	assign g2938 = (((!ax16x) & (!g2779) & (!g2828) & (!g2853) & (g2865)) + ((!ax16x) & (!g2779) & (g2828) & (!g2853) & (!g2865)) + ((!ax16x) & (!g2779) & (g2828) & (!g2853) & (g2865)) + ((!ax16x) & (!g2779) & (g2828) & (g2853) & (!g2865)) + ((!ax16x) & (!g2779) & (g2828) & (g2853) & (g2865)) + ((!ax16x) & (g2779) & (g2828) & (!g2853) & (!g2865)) + ((!ax16x) & (g2779) & (g2828) & (g2853) & (!g2865)) + ((!ax16x) & (g2779) & (g2828) & (g2853) & (g2865)) + ((ax16x) & (!g2779) & (!g2828) & (!g2853) & (!g2865)) + ((ax16x) & (!g2779) & (!g2828) & (g2853) & (!g2865)) + ((ax16x) & (!g2779) & (!g2828) & (g2853) & (g2865)) + ((ax16x) & (g2779) & (!g2828) & (!g2853) & (!g2865)) + ((ax16x) & (g2779) & (!g2828) & (!g2853) & (g2865)) + ((ax16x) & (g2779) & (!g2828) & (g2853) & (!g2865)) + ((ax16x) & (g2779) & (!g2828) & (g2853) & (g2865)) + ((ax16x) & (g2779) & (g2828) & (!g2853) & (g2865)));
	assign g2939 = (((!ax12x) & (!ax13x)));
	assign g2940 = (((!g2779) & (!ax14x) & (!ax15x) & (!g2853) & (!g2865) & (!g2939)) + ((!g2779) & (!ax14x) & (!ax15x) & (g2853) & (!g2865) & (!g2939)) + ((!g2779) & (!ax14x) & (!ax15x) & (g2853) & (g2865) & (!g2939)) + ((!g2779) & (!ax14x) & (ax15x) & (!g2853) & (g2865) & (!g2939)) + ((!g2779) & (ax14x) & (ax15x) & (!g2853) & (g2865) & (!g2939)) + ((!g2779) & (ax14x) & (ax15x) & (!g2853) & (g2865) & (g2939)) + ((g2779) & (!ax14x) & (!ax15x) & (!g2853) & (!g2865) & (!g2939)) + ((g2779) & (!ax14x) & (!ax15x) & (!g2853) & (!g2865) & (g2939)) + ((g2779) & (!ax14x) & (!ax15x) & (!g2853) & (g2865) & (!g2939)) + ((g2779) & (!ax14x) & (!ax15x) & (g2853) & (!g2865) & (!g2939)) + ((g2779) & (!ax14x) & (!ax15x) & (g2853) & (!g2865) & (g2939)) + ((g2779) & (!ax14x) & (!ax15x) & (g2853) & (g2865) & (!g2939)) + ((g2779) & (!ax14x) & (!ax15x) & (g2853) & (g2865) & (g2939)) + ((g2779) & (!ax14x) & (ax15x) & (!g2853) & (!g2865) & (!g2939)) + ((g2779) & (!ax14x) & (ax15x) & (!g2853) & (g2865) & (!g2939)) + ((g2779) & (!ax14x) & (ax15x) & (!g2853) & (g2865) & (g2939)) + ((g2779) & (!ax14x) & (ax15x) & (g2853) & (!g2865) & (!g2939)) + ((g2779) & (!ax14x) & (ax15x) & (g2853) & (g2865) & (!g2939)) + ((g2779) & (ax14x) & (!ax15x) & (!g2853) & (g2865) & (!g2939)) + ((g2779) & (ax14x) & (!ax15x) & (!g2853) & (g2865) & (g2939)) + ((g2779) & (ax14x) & (ax15x) & (!g2853) & (!g2865) & (!g2939)) + ((g2779) & (ax14x) & (ax15x) & (!g2853) & (!g2865) & (g2939)) + ((g2779) & (ax14x) & (ax15x) & (!g2853) & (g2865) & (!g2939)) + ((g2779) & (ax14x) & (ax15x) & (!g2853) & (g2865) & (g2939)) + ((g2779) & (ax14x) & (ax15x) & (g2853) & (!g2865) & (!g2939)) + ((g2779) & (ax14x) & (ax15x) & (g2853) & (!g2865) & (g2939)) + ((g2779) & (ax14x) & (ax15x) & (g2853) & (g2865) & (!g2939)) + ((g2779) & (ax14x) & (ax15x) & (g2853) & (g2865) & (g2939)));
	assign g2941 = (((!g2585) & (!g2825) & (g2937) & (g2938) & (g2940)) + ((!g2585) & (g2825) & (g2937) & (!g2938) & (g2940)) + ((!g2585) & (g2825) & (g2937) & (g2938) & (!g2940)) + ((!g2585) & (g2825) & (g2937) & (g2938) & (g2940)) + ((g2585) & (!g2825) & (!g2937) & (g2938) & (g2940)) + ((g2585) & (!g2825) & (g2937) & (!g2938) & (!g2940)) + ((g2585) & (!g2825) & (g2937) & (!g2938) & (g2940)) + ((g2585) & (!g2825) & (g2937) & (g2938) & (!g2940)) + ((g2585) & (!g2825) & (g2937) & (g2938) & (g2940)) + ((g2585) & (g2825) & (!g2937) & (!g2938) & (g2940)) + ((g2585) & (g2825) & (!g2937) & (g2938) & (!g2940)) + ((g2585) & (g2825) & (!g2937) & (g2938) & (g2940)) + ((g2585) & (g2825) & (g2937) & (!g2938) & (!g2940)) + ((g2585) & (g2825) & (g2937) & (!g2938) & (g2940)) + ((g2585) & (g2825) & (g2937) & (g2938) & (!g2940)) + ((g2585) & (g2825) & (g2937) & (g2938) & (g2940)));
	assign g2942 = (((!g2398) & (!g2627) & (g2934) & (g2935) & (g2941)) + ((!g2398) & (g2627) & (g2934) & (!g2935) & (g2941)) + ((!g2398) & (g2627) & (g2934) & (g2935) & (!g2941)) + ((!g2398) & (g2627) & (g2934) & (g2935) & (g2941)) + ((g2398) & (!g2627) & (!g2934) & (g2935) & (g2941)) + ((g2398) & (!g2627) & (g2934) & (!g2935) & (!g2941)) + ((g2398) & (!g2627) & (g2934) & (!g2935) & (g2941)) + ((g2398) & (!g2627) & (g2934) & (g2935) & (!g2941)) + ((g2398) & (!g2627) & (g2934) & (g2935) & (g2941)) + ((g2398) & (g2627) & (!g2934) & (!g2935) & (g2941)) + ((g2398) & (g2627) & (!g2934) & (g2935) & (!g2941)) + ((g2398) & (g2627) & (!g2934) & (g2935) & (g2941)) + ((g2398) & (g2627) & (g2934) & (!g2935) & (!g2941)) + ((g2398) & (g2627) & (g2934) & (!g2935) & (g2941)) + ((g2398) & (g2627) & (g2934) & (g2935) & (!g2941)) + ((g2398) & (g2627) & (g2934) & (g2935) & (g2941)));
	assign g2943 = (((!g2218) & (!g2436) & (g2931) & (g2932) & (g2942)) + ((!g2218) & (g2436) & (g2931) & (!g2932) & (g2942)) + ((!g2218) & (g2436) & (g2931) & (g2932) & (!g2942)) + ((!g2218) & (g2436) & (g2931) & (g2932) & (g2942)) + ((g2218) & (!g2436) & (!g2931) & (g2932) & (g2942)) + ((g2218) & (!g2436) & (g2931) & (!g2932) & (!g2942)) + ((g2218) & (!g2436) & (g2931) & (!g2932) & (g2942)) + ((g2218) & (!g2436) & (g2931) & (g2932) & (!g2942)) + ((g2218) & (!g2436) & (g2931) & (g2932) & (g2942)) + ((g2218) & (g2436) & (!g2931) & (!g2932) & (g2942)) + ((g2218) & (g2436) & (!g2931) & (g2932) & (!g2942)) + ((g2218) & (g2436) & (!g2931) & (g2932) & (g2942)) + ((g2218) & (g2436) & (g2931) & (!g2932) & (!g2942)) + ((g2218) & (g2436) & (g2931) & (!g2932) & (g2942)) + ((g2218) & (g2436) & (g2931) & (g2932) & (!g2942)) + ((g2218) & (g2436) & (g2931) & (g2932) & (g2942)));
	assign g2944 = (((!g2045) & (!g2252) & (g2928) & (g2929) & (g2943)) + ((!g2045) & (g2252) & (g2928) & (!g2929) & (g2943)) + ((!g2045) & (g2252) & (g2928) & (g2929) & (!g2943)) + ((!g2045) & (g2252) & (g2928) & (g2929) & (g2943)) + ((g2045) & (!g2252) & (!g2928) & (g2929) & (g2943)) + ((g2045) & (!g2252) & (g2928) & (!g2929) & (!g2943)) + ((g2045) & (!g2252) & (g2928) & (!g2929) & (g2943)) + ((g2045) & (!g2252) & (g2928) & (g2929) & (!g2943)) + ((g2045) & (!g2252) & (g2928) & (g2929) & (g2943)) + ((g2045) & (g2252) & (!g2928) & (!g2929) & (g2943)) + ((g2045) & (g2252) & (!g2928) & (g2929) & (!g2943)) + ((g2045) & (g2252) & (!g2928) & (g2929) & (g2943)) + ((g2045) & (g2252) & (g2928) & (!g2929) & (!g2943)) + ((g2045) & (g2252) & (g2928) & (!g2929) & (g2943)) + ((g2045) & (g2252) & (g2928) & (g2929) & (!g2943)) + ((g2045) & (g2252) & (g2928) & (g2929) & (g2943)));
	assign g2945 = (((!g1879) & (!g2075) & (g2925) & (g2926) & (g2944)) + ((!g1879) & (g2075) & (g2925) & (!g2926) & (g2944)) + ((!g1879) & (g2075) & (g2925) & (g2926) & (!g2944)) + ((!g1879) & (g2075) & (g2925) & (g2926) & (g2944)) + ((g1879) & (!g2075) & (!g2925) & (g2926) & (g2944)) + ((g1879) & (!g2075) & (g2925) & (!g2926) & (!g2944)) + ((g1879) & (!g2075) & (g2925) & (!g2926) & (g2944)) + ((g1879) & (!g2075) & (g2925) & (g2926) & (!g2944)) + ((g1879) & (!g2075) & (g2925) & (g2926) & (g2944)) + ((g1879) & (g2075) & (!g2925) & (!g2926) & (g2944)) + ((g1879) & (g2075) & (!g2925) & (g2926) & (!g2944)) + ((g1879) & (g2075) & (!g2925) & (g2926) & (g2944)) + ((g1879) & (g2075) & (g2925) & (!g2926) & (!g2944)) + ((g1879) & (g2075) & (g2925) & (!g2926) & (g2944)) + ((g1879) & (g2075) & (g2925) & (g2926) & (!g2944)) + ((g1879) & (g2075) & (g2925) & (g2926) & (g2944)));
	assign g2946 = (((!g1720) & (!g1905) & (g2922) & (g2923) & (g2945)) + ((!g1720) & (g1905) & (g2922) & (!g2923) & (g2945)) + ((!g1720) & (g1905) & (g2922) & (g2923) & (!g2945)) + ((!g1720) & (g1905) & (g2922) & (g2923) & (g2945)) + ((g1720) & (!g1905) & (!g2922) & (g2923) & (g2945)) + ((g1720) & (!g1905) & (g2922) & (!g2923) & (!g2945)) + ((g1720) & (!g1905) & (g2922) & (!g2923) & (g2945)) + ((g1720) & (!g1905) & (g2922) & (g2923) & (!g2945)) + ((g1720) & (!g1905) & (g2922) & (g2923) & (g2945)) + ((g1720) & (g1905) & (!g2922) & (!g2923) & (g2945)) + ((g1720) & (g1905) & (!g2922) & (g2923) & (!g2945)) + ((g1720) & (g1905) & (!g2922) & (g2923) & (g2945)) + ((g1720) & (g1905) & (g2922) & (!g2923) & (!g2945)) + ((g1720) & (g1905) & (g2922) & (!g2923) & (g2945)) + ((g1720) & (g1905) & (g2922) & (g2923) & (!g2945)) + ((g1720) & (g1905) & (g2922) & (g2923) & (g2945)));
	assign g2947 = (((!g1568) & (!g1742) & (g2919) & (g2920) & (g2946)) + ((!g1568) & (g1742) & (g2919) & (!g2920) & (g2946)) + ((!g1568) & (g1742) & (g2919) & (g2920) & (!g2946)) + ((!g1568) & (g1742) & (g2919) & (g2920) & (g2946)) + ((g1568) & (!g1742) & (!g2919) & (g2920) & (g2946)) + ((g1568) & (!g1742) & (g2919) & (!g2920) & (!g2946)) + ((g1568) & (!g1742) & (g2919) & (!g2920) & (g2946)) + ((g1568) & (!g1742) & (g2919) & (g2920) & (!g2946)) + ((g1568) & (!g1742) & (g2919) & (g2920) & (g2946)) + ((g1568) & (g1742) & (!g2919) & (!g2920) & (g2946)) + ((g1568) & (g1742) & (!g2919) & (g2920) & (!g2946)) + ((g1568) & (g1742) & (!g2919) & (g2920) & (g2946)) + ((g1568) & (g1742) & (g2919) & (!g2920) & (!g2946)) + ((g1568) & (g1742) & (g2919) & (!g2920) & (g2946)) + ((g1568) & (g1742) & (g2919) & (g2920) & (!g2946)) + ((g1568) & (g1742) & (g2919) & (g2920) & (g2946)));
	assign g2948 = (((!g1423) & (!g1586) & (g2916) & (g2917) & (g2947)) + ((!g1423) & (g1586) & (g2916) & (!g2917) & (g2947)) + ((!g1423) & (g1586) & (g2916) & (g2917) & (!g2947)) + ((!g1423) & (g1586) & (g2916) & (g2917) & (g2947)) + ((g1423) & (!g1586) & (!g2916) & (g2917) & (g2947)) + ((g1423) & (!g1586) & (g2916) & (!g2917) & (!g2947)) + ((g1423) & (!g1586) & (g2916) & (!g2917) & (g2947)) + ((g1423) & (!g1586) & (g2916) & (g2917) & (!g2947)) + ((g1423) & (!g1586) & (g2916) & (g2917) & (g2947)) + ((g1423) & (g1586) & (!g2916) & (!g2917) & (g2947)) + ((g1423) & (g1586) & (!g2916) & (g2917) & (!g2947)) + ((g1423) & (g1586) & (!g2916) & (g2917) & (g2947)) + ((g1423) & (g1586) & (g2916) & (!g2917) & (!g2947)) + ((g1423) & (g1586) & (g2916) & (!g2917) & (g2947)) + ((g1423) & (g1586) & (g2916) & (g2917) & (!g2947)) + ((g1423) & (g1586) & (g2916) & (g2917) & (g2947)));
	assign g2949 = (((!g1285) & (!g1437) & (g2913) & (g2914) & (g2948)) + ((!g1285) & (g1437) & (g2913) & (!g2914) & (g2948)) + ((!g1285) & (g1437) & (g2913) & (g2914) & (!g2948)) + ((!g1285) & (g1437) & (g2913) & (g2914) & (g2948)) + ((g1285) & (!g1437) & (!g2913) & (g2914) & (g2948)) + ((g1285) & (!g1437) & (g2913) & (!g2914) & (!g2948)) + ((g1285) & (!g1437) & (g2913) & (!g2914) & (g2948)) + ((g1285) & (!g1437) & (g2913) & (g2914) & (!g2948)) + ((g1285) & (!g1437) & (g2913) & (g2914) & (g2948)) + ((g1285) & (g1437) & (!g2913) & (!g2914) & (g2948)) + ((g1285) & (g1437) & (!g2913) & (g2914) & (!g2948)) + ((g1285) & (g1437) & (!g2913) & (g2914) & (g2948)) + ((g1285) & (g1437) & (g2913) & (!g2914) & (!g2948)) + ((g1285) & (g1437) & (g2913) & (!g2914) & (g2948)) + ((g1285) & (g1437) & (g2913) & (g2914) & (!g2948)) + ((g1285) & (g1437) & (g2913) & (g2914) & (g2948)));
	assign g2950 = (((!g1154) & (!g1295) & (g2910) & (g2911) & (g2949)) + ((!g1154) & (g1295) & (g2910) & (!g2911) & (g2949)) + ((!g1154) & (g1295) & (g2910) & (g2911) & (!g2949)) + ((!g1154) & (g1295) & (g2910) & (g2911) & (g2949)) + ((g1154) & (!g1295) & (!g2910) & (g2911) & (g2949)) + ((g1154) & (!g1295) & (g2910) & (!g2911) & (!g2949)) + ((g1154) & (!g1295) & (g2910) & (!g2911) & (g2949)) + ((g1154) & (!g1295) & (g2910) & (g2911) & (!g2949)) + ((g1154) & (!g1295) & (g2910) & (g2911) & (g2949)) + ((g1154) & (g1295) & (!g2910) & (!g2911) & (g2949)) + ((g1154) & (g1295) & (!g2910) & (g2911) & (!g2949)) + ((g1154) & (g1295) & (!g2910) & (g2911) & (g2949)) + ((g1154) & (g1295) & (g2910) & (!g2911) & (!g2949)) + ((g1154) & (g1295) & (g2910) & (!g2911) & (g2949)) + ((g1154) & (g1295) & (g2910) & (g2911) & (!g2949)) + ((g1154) & (g1295) & (g2910) & (g2911) & (g2949)));
	assign g2951 = (((!g1030) & (!g1160) & (g2907) & (g2908) & (g2950)) + ((!g1030) & (g1160) & (g2907) & (!g2908) & (g2950)) + ((!g1030) & (g1160) & (g2907) & (g2908) & (!g2950)) + ((!g1030) & (g1160) & (g2907) & (g2908) & (g2950)) + ((g1030) & (!g1160) & (!g2907) & (g2908) & (g2950)) + ((g1030) & (!g1160) & (g2907) & (!g2908) & (!g2950)) + ((g1030) & (!g1160) & (g2907) & (!g2908) & (g2950)) + ((g1030) & (!g1160) & (g2907) & (g2908) & (!g2950)) + ((g1030) & (!g1160) & (g2907) & (g2908) & (g2950)) + ((g1030) & (g1160) & (!g2907) & (!g2908) & (g2950)) + ((g1030) & (g1160) & (!g2907) & (g2908) & (!g2950)) + ((g1030) & (g1160) & (!g2907) & (g2908) & (g2950)) + ((g1030) & (g1160) & (g2907) & (!g2908) & (!g2950)) + ((g1030) & (g1160) & (g2907) & (!g2908) & (g2950)) + ((g1030) & (g1160) & (g2907) & (g2908) & (!g2950)) + ((g1030) & (g1160) & (g2907) & (g2908) & (g2950)));
	assign g2952 = (((!g914) & (!g1032) & (g2904) & (g2905) & (g2951)) + ((!g914) & (g1032) & (g2904) & (!g2905) & (g2951)) + ((!g914) & (g1032) & (g2904) & (g2905) & (!g2951)) + ((!g914) & (g1032) & (g2904) & (g2905) & (g2951)) + ((g914) & (!g1032) & (!g2904) & (g2905) & (g2951)) + ((g914) & (!g1032) & (g2904) & (!g2905) & (!g2951)) + ((g914) & (!g1032) & (g2904) & (!g2905) & (g2951)) + ((g914) & (!g1032) & (g2904) & (g2905) & (!g2951)) + ((g914) & (!g1032) & (g2904) & (g2905) & (g2951)) + ((g914) & (g1032) & (!g2904) & (!g2905) & (g2951)) + ((g914) & (g1032) & (!g2904) & (g2905) & (!g2951)) + ((g914) & (g1032) & (!g2904) & (g2905) & (g2951)) + ((g914) & (g1032) & (g2904) & (!g2905) & (!g2951)) + ((g914) & (g1032) & (g2904) & (!g2905) & (g2951)) + ((g914) & (g1032) & (g2904) & (g2905) & (!g2951)) + ((g914) & (g1032) & (g2904) & (g2905) & (g2951)));
	assign g2953 = (((!g803) & (!g851) & (g2901) & (g2902) & (g2952)) + ((!g803) & (g851) & (g2901) & (!g2902) & (g2952)) + ((!g803) & (g851) & (g2901) & (g2902) & (!g2952)) + ((!g803) & (g851) & (g2901) & (g2902) & (g2952)) + ((g803) & (!g851) & (!g2901) & (g2902) & (g2952)) + ((g803) & (!g851) & (g2901) & (!g2902) & (!g2952)) + ((g803) & (!g851) & (g2901) & (!g2902) & (g2952)) + ((g803) & (!g851) & (g2901) & (g2902) & (!g2952)) + ((g803) & (!g851) & (g2901) & (g2902) & (g2952)) + ((g803) & (g851) & (!g2901) & (!g2902) & (g2952)) + ((g803) & (g851) & (!g2901) & (g2902) & (!g2952)) + ((g803) & (g851) & (!g2901) & (g2902) & (g2952)) + ((g803) & (g851) & (g2901) & (!g2902) & (!g2952)) + ((g803) & (g851) & (g2901) & (!g2902) & (g2952)) + ((g803) & (g851) & (g2901) & (g2902) & (!g2952)) + ((g803) & (g851) & (g2901) & (g2902) & (g2952)));
	assign g2954 = (((!g700) & (!g744) & (g2898) & (g2899) & (g2953)) + ((!g700) & (g744) & (g2898) & (!g2899) & (g2953)) + ((!g700) & (g744) & (g2898) & (g2899) & (!g2953)) + ((!g700) & (g744) & (g2898) & (g2899) & (g2953)) + ((g700) & (!g744) & (!g2898) & (g2899) & (g2953)) + ((g700) & (!g744) & (g2898) & (!g2899) & (!g2953)) + ((g700) & (!g744) & (g2898) & (!g2899) & (g2953)) + ((g700) & (!g744) & (g2898) & (g2899) & (!g2953)) + ((g700) & (!g744) & (g2898) & (g2899) & (g2953)) + ((g700) & (g744) & (!g2898) & (!g2899) & (g2953)) + ((g700) & (g744) & (!g2898) & (g2899) & (!g2953)) + ((g700) & (g744) & (!g2898) & (g2899) & (g2953)) + ((g700) & (g744) & (g2898) & (!g2899) & (!g2953)) + ((g700) & (g744) & (g2898) & (!g2899) & (g2953)) + ((g700) & (g744) & (g2898) & (g2899) & (!g2953)) + ((g700) & (g744) & (g2898) & (g2899) & (g2953)));
	assign g2955 = (((!g604) & (!g645) & (g2895) & (g2896) & (g2954)) + ((!g604) & (g645) & (g2895) & (!g2896) & (g2954)) + ((!g604) & (g645) & (g2895) & (g2896) & (!g2954)) + ((!g604) & (g645) & (g2895) & (g2896) & (g2954)) + ((g604) & (!g645) & (!g2895) & (g2896) & (g2954)) + ((g604) & (!g645) & (g2895) & (!g2896) & (!g2954)) + ((g604) & (!g645) & (g2895) & (!g2896) & (g2954)) + ((g604) & (!g645) & (g2895) & (g2896) & (!g2954)) + ((g604) & (!g645) & (g2895) & (g2896) & (g2954)) + ((g604) & (g645) & (!g2895) & (!g2896) & (g2954)) + ((g604) & (g645) & (!g2895) & (g2896) & (!g2954)) + ((g604) & (g645) & (!g2895) & (g2896) & (g2954)) + ((g604) & (g645) & (g2895) & (!g2896) & (!g2954)) + ((g604) & (g645) & (g2895) & (!g2896) & (g2954)) + ((g604) & (g645) & (g2895) & (g2896) & (!g2954)) + ((g604) & (g645) & (g2895) & (g2896) & (g2954)));
	assign g2956 = (((!g515) & (!g553) & (g2892) & (g2893) & (g2955)) + ((!g515) & (g553) & (g2892) & (!g2893) & (g2955)) + ((!g515) & (g553) & (g2892) & (g2893) & (!g2955)) + ((!g515) & (g553) & (g2892) & (g2893) & (g2955)) + ((g515) & (!g553) & (!g2892) & (g2893) & (g2955)) + ((g515) & (!g553) & (g2892) & (!g2893) & (!g2955)) + ((g515) & (!g553) & (g2892) & (!g2893) & (g2955)) + ((g515) & (!g553) & (g2892) & (g2893) & (!g2955)) + ((g515) & (!g553) & (g2892) & (g2893) & (g2955)) + ((g515) & (g553) & (!g2892) & (!g2893) & (g2955)) + ((g515) & (g553) & (!g2892) & (g2893) & (!g2955)) + ((g515) & (g553) & (!g2892) & (g2893) & (g2955)) + ((g515) & (g553) & (g2892) & (!g2893) & (!g2955)) + ((g515) & (g553) & (g2892) & (!g2893) & (g2955)) + ((g515) & (g553) & (g2892) & (g2893) & (!g2955)) + ((g515) & (g553) & (g2892) & (g2893) & (g2955)));
	assign g2957 = (((!g433) & (!g468) & (g2889) & (g2890) & (g2956)) + ((!g433) & (g468) & (g2889) & (!g2890) & (g2956)) + ((!g433) & (g468) & (g2889) & (g2890) & (!g2956)) + ((!g433) & (g468) & (g2889) & (g2890) & (g2956)) + ((g433) & (!g468) & (!g2889) & (g2890) & (g2956)) + ((g433) & (!g468) & (g2889) & (!g2890) & (!g2956)) + ((g433) & (!g468) & (g2889) & (!g2890) & (g2956)) + ((g433) & (!g468) & (g2889) & (g2890) & (!g2956)) + ((g433) & (!g468) & (g2889) & (g2890) & (g2956)) + ((g433) & (g468) & (!g2889) & (!g2890) & (g2956)) + ((g433) & (g468) & (!g2889) & (g2890) & (!g2956)) + ((g433) & (g468) & (!g2889) & (g2890) & (g2956)) + ((g433) & (g468) & (g2889) & (!g2890) & (!g2956)) + ((g433) & (g468) & (g2889) & (!g2890) & (g2956)) + ((g433) & (g468) & (g2889) & (g2890) & (!g2956)) + ((g433) & (g468) & (g2889) & (g2890) & (g2956)));
	assign g2958 = (((!g358) & (!g390) & (g2886) & (g2887) & (g2957)) + ((!g358) & (g390) & (g2886) & (!g2887) & (g2957)) + ((!g358) & (g390) & (g2886) & (g2887) & (!g2957)) + ((!g358) & (g390) & (g2886) & (g2887) & (g2957)) + ((g358) & (!g390) & (!g2886) & (g2887) & (g2957)) + ((g358) & (!g390) & (g2886) & (!g2887) & (!g2957)) + ((g358) & (!g390) & (g2886) & (!g2887) & (g2957)) + ((g358) & (!g390) & (g2886) & (g2887) & (!g2957)) + ((g358) & (!g390) & (g2886) & (g2887) & (g2957)) + ((g358) & (g390) & (!g2886) & (!g2887) & (g2957)) + ((g358) & (g390) & (!g2886) & (g2887) & (!g2957)) + ((g358) & (g390) & (!g2886) & (g2887) & (g2957)) + ((g358) & (g390) & (g2886) & (!g2887) & (!g2957)) + ((g358) & (g390) & (g2886) & (!g2887) & (g2957)) + ((g358) & (g390) & (g2886) & (g2887) & (!g2957)) + ((g358) & (g390) & (g2886) & (g2887) & (g2957)));
	assign g2959 = (((!g290) & (!g319) & (g2883) & (g2884) & (g2958)) + ((!g290) & (g319) & (g2883) & (!g2884) & (g2958)) + ((!g290) & (g319) & (g2883) & (g2884) & (!g2958)) + ((!g290) & (g319) & (g2883) & (g2884) & (g2958)) + ((g290) & (!g319) & (!g2883) & (g2884) & (g2958)) + ((g290) & (!g319) & (g2883) & (!g2884) & (!g2958)) + ((g290) & (!g319) & (g2883) & (!g2884) & (g2958)) + ((g290) & (!g319) & (g2883) & (g2884) & (!g2958)) + ((g290) & (!g319) & (g2883) & (g2884) & (g2958)) + ((g290) & (g319) & (!g2883) & (!g2884) & (g2958)) + ((g290) & (g319) & (!g2883) & (g2884) & (!g2958)) + ((g290) & (g319) & (!g2883) & (g2884) & (g2958)) + ((g290) & (g319) & (g2883) & (!g2884) & (!g2958)) + ((g290) & (g319) & (g2883) & (!g2884) & (g2958)) + ((g290) & (g319) & (g2883) & (g2884) & (!g2958)) + ((g290) & (g319) & (g2883) & (g2884) & (g2958)));
	assign g2960 = (((!g229) & (!g255) & (g2880) & (g2881) & (g2959)) + ((!g229) & (g255) & (g2880) & (!g2881) & (g2959)) + ((!g229) & (g255) & (g2880) & (g2881) & (!g2959)) + ((!g229) & (g255) & (g2880) & (g2881) & (g2959)) + ((g229) & (!g255) & (!g2880) & (g2881) & (g2959)) + ((g229) & (!g255) & (g2880) & (!g2881) & (!g2959)) + ((g229) & (!g255) & (g2880) & (!g2881) & (g2959)) + ((g229) & (!g255) & (g2880) & (g2881) & (!g2959)) + ((g229) & (!g255) & (g2880) & (g2881) & (g2959)) + ((g229) & (g255) & (!g2880) & (!g2881) & (g2959)) + ((g229) & (g255) & (!g2880) & (g2881) & (!g2959)) + ((g229) & (g255) & (!g2880) & (g2881) & (g2959)) + ((g229) & (g255) & (g2880) & (!g2881) & (!g2959)) + ((g229) & (g255) & (g2880) & (!g2881) & (g2959)) + ((g229) & (g255) & (g2880) & (g2881) & (!g2959)) + ((g229) & (g255) & (g2880) & (g2881) & (g2959)));
	assign g2961 = (((!g174) & (!g198) & (g2877) & (g2878) & (g2960)) + ((!g174) & (g198) & (g2877) & (!g2878) & (g2960)) + ((!g174) & (g198) & (g2877) & (g2878) & (!g2960)) + ((!g174) & (g198) & (g2877) & (g2878) & (g2960)) + ((g174) & (!g198) & (!g2877) & (g2878) & (g2960)) + ((g174) & (!g198) & (g2877) & (!g2878) & (!g2960)) + ((g174) & (!g198) & (g2877) & (!g2878) & (g2960)) + ((g174) & (!g198) & (g2877) & (g2878) & (!g2960)) + ((g174) & (!g198) & (g2877) & (g2878) & (g2960)) + ((g174) & (g198) & (!g2877) & (!g2878) & (g2960)) + ((g174) & (g198) & (!g2877) & (g2878) & (!g2960)) + ((g174) & (g198) & (!g2877) & (g2878) & (g2960)) + ((g174) & (g198) & (g2877) & (!g2878) & (!g2960)) + ((g174) & (g198) & (g2877) & (!g2878) & (g2960)) + ((g174) & (g198) & (g2877) & (g2878) & (!g2960)) + ((g174) & (g198) & (g2877) & (g2878) & (g2960)));
	assign g2962 = (((!g127) & (!g147) & (g2874) & (g2875) & (g2961)) + ((!g127) & (g147) & (g2874) & (!g2875) & (g2961)) + ((!g127) & (g147) & (g2874) & (g2875) & (!g2961)) + ((!g127) & (g147) & (g2874) & (g2875) & (g2961)) + ((g127) & (!g147) & (!g2874) & (g2875) & (g2961)) + ((g127) & (!g147) & (g2874) & (!g2875) & (!g2961)) + ((g127) & (!g147) & (g2874) & (!g2875) & (g2961)) + ((g127) & (!g147) & (g2874) & (g2875) & (!g2961)) + ((g127) & (!g147) & (g2874) & (g2875) & (g2961)) + ((g127) & (g147) & (!g2874) & (!g2875) & (g2961)) + ((g127) & (g147) & (!g2874) & (g2875) & (!g2961)) + ((g127) & (g147) & (!g2874) & (g2875) & (g2961)) + ((g127) & (g147) & (g2874) & (!g2875) & (!g2961)) + ((g127) & (g147) & (g2874) & (!g2875) & (g2961)) + ((g127) & (g147) & (g2874) & (g2875) & (!g2961)) + ((g127) & (g147) & (g2874) & (g2875) & (g2961)));
	assign g2963 = (((!g87) & (!g104) & (g2871) & (g2872) & (g2962)) + ((!g87) & (g104) & (g2871) & (!g2872) & (g2962)) + ((!g87) & (g104) & (g2871) & (g2872) & (!g2962)) + ((!g87) & (g104) & (g2871) & (g2872) & (g2962)) + ((g87) & (!g104) & (!g2871) & (g2872) & (g2962)) + ((g87) & (!g104) & (g2871) & (!g2872) & (!g2962)) + ((g87) & (!g104) & (g2871) & (!g2872) & (g2962)) + ((g87) & (!g104) & (g2871) & (g2872) & (!g2962)) + ((g87) & (!g104) & (g2871) & (g2872) & (g2962)) + ((g87) & (g104) & (!g2871) & (!g2872) & (g2962)) + ((g87) & (g104) & (!g2871) & (g2872) & (!g2962)) + ((g87) & (g104) & (!g2871) & (g2872) & (g2962)) + ((g87) & (g104) & (g2871) & (!g2872) & (!g2962)) + ((g87) & (g104) & (g2871) & (!g2872) & (g2962)) + ((g87) & (g104) & (g2871) & (g2872) & (!g2962)) + ((g87) & (g104) & (g2871) & (g2872) & (g2962)));
	assign g2964 = (((!g54) & (!g68) & (g2868) & (g2869) & (g2963)) + ((!g54) & (g68) & (g2868) & (!g2869) & (g2963)) + ((!g54) & (g68) & (g2868) & (g2869) & (!g2963)) + ((!g54) & (g68) & (g2868) & (g2869) & (g2963)) + ((g54) & (!g68) & (!g2868) & (g2869) & (g2963)) + ((g54) & (!g68) & (g2868) & (!g2869) & (!g2963)) + ((g54) & (!g68) & (g2868) & (!g2869) & (g2963)) + ((g54) & (!g68) & (g2868) & (g2869) & (!g2963)) + ((g54) & (!g68) & (g2868) & (g2869) & (g2963)) + ((g54) & (g68) & (!g2868) & (!g2869) & (g2963)) + ((g54) & (g68) & (!g2868) & (g2869) & (!g2963)) + ((g54) & (g68) & (!g2868) & (g2869) & (g2963)) + ((g54) & (g68) & (g2868) & (!g2869) & (!g2963)) + ((g54) & (g68) & (g2868) & (!g2869) & (g2963)) + ((g54) & (g68) & (g2868) & (g2869) & (!g2963)) + ((g54) & (g68) & (g2868) & (g2869) & (g2963)));
	assign g2965 = (((!g4) & (!g2862) & (!g2863) & (!g2853) & (!g2865)) + ((!g4) & (!g2862) & (!g2863) & (g2853) & (!g2865)) + ((!g4) & (!g2862) & (!g2863) & (g2853) & (g2865)) + ((!g4) & (!g2862) & (g2863) & (!g2853) & (g2865)) + ((!g4) & (g2862) & (g2863) & (!g2853) & (!g2865)) + ((!g4) & (g2862) & (g2863) & (!g2853) & (g2865)) + ((!g4) & (g2862) & (g2863) & (g2853) & (!g2865)) + ((!g4) & (g2862) & (g2863) & (g2853) & (g2865)) + ((g4) & (!g2862) & (g2863) & (!g2853) & (!g2865)) + ((g4) & (!g2862) & (g2863) & (!g2853) & (g2865)) + ((g4) & (!g2862) & (g2863) & (g2853) & (!g2865)) + ((g4) & (!g2862) & (g2863) & (g2853) & (g2865)) + ((g4) & (g2862) & (!g2863) & (!g2853) & (!g2865)) + ((g4) & (g2862) & (!g2863) & (g2853) & (!g2865)) + ((g4) & (g2862) & (!g2863) & (g2853) & (g2865)) + ((g4) & (g2862) & (g2863) & (!g2853) & (g2865)));
	assign g2966 = (((!g8) & (!g2856) & (g2861) & (!g2853) & (!g2865)) + ((!g8) & (!g2856) & (g2861) & (g2853) & (!g2865)) + ((!g8) & (!g2856) & (g2861) & (g2853) & (g2865)) + ((!g8) & (g2856) & (!g2861) & (!g2853) & (!g2865)) + ((!g8) & (g2856) & (!g2861) & (!g2853) & (g2865)) + ((!g8) & (g2856) & (!g2861) & (g2853) & (!g2865)) + ((!g8) & (g2856) & (!g2861) & (g2853) & (g2865)) + ((!g8) & (g2856) & (g2861) & (!g2853) & (g2865)) + ((g8) & (!g2856) & (!g2861) & (!g2853) & (!g2865)) + ((g8) & (!g2856) & (!g2861) & (g2853) & (!g2865)) + ((g8) & (!g2856) & (!g2861) & (g2853) & (g2865)) + ((g8) & (g2856) & (!g2861) & (!g2853) & (g2865)) + ((g8) & (g2856) & (g2861) & (!g2853) & (!g2865)) + ((g8) & (g2856) & (g2861) & (!g2853) & (g2865)) + ((g8) & (g2856) & (g2861) & (g2853) & (!g2865)) + ((g8) & (g2856) & (g2861) & (g2853) & (g2865)));
	assign g2967 = (((!g18) & (!g27) & (g2858) & (g2860)) + ((!g18) & (g27) & (!g2858) & (g2860)) + ((!g18) & (g27) & (g2858) & (!g2860)) + ((!g18) & (g27) & (g2858) & (g2860)) + ((g18) & (!g27) & (!g2858) & (!g2860)) + ((g18) & (!g27) & (!g2858) & (g2860)) + ((g18) & (!g27) & (g2858) & (!g2860)) + ((g18) & (g27) & (!g2858) & (!g2860)));
	assign g2968 = (((!g2857) & (!g2853) & (!g2865) & (g2967)) + ((!g2857) & (g2853) & (!g2865) & (g2967)) + ((!g2857) & (g2853) & (g2865) & (g2967)) + ((g2857) & (!g2853) & (!g2865) & (!g2967)) + ((g2857) & (!g2853) & (g2865) & (!g2967)) + ((g2857) & (!g2853) & (g2865) & (g2967)) + ((g2857) & (g2853) & (!g2865) & (!g2967)) + ((g2857) & (g2853) & (g2865) & (!g2967)));
	assign g2969 = (((!g27) & (!g2858) & (g2860) & (!g2853) & (!g2865)) + ((!g27) & (!g2858) & (g2860) & (g2853) & (!g2865)) + ((!g27) & (!g2858) & (g2860) & (g2853) & (g2865)) + ((!g27) & (g2858) & (!g2860) & (!g2853) & (!g2865)) + ((!g27) & (g2858) & (!g2860) & (!g2853) & (g2865)) + ((!g27) & (g2858) & (!g2860) & (g2853) & (!g2865)) + ((!g27) & (g2858) & (!g2860) & (g2853) & (g2865)) + ((!g27) & (g2858) & (g2860) & (!g2853) & (g2865)) + ((g27) & (!g2858) & (!g2860) & (!g2853) & (!g2865)) + ((g27) & (!g2858) & (!g2860) & (g2853) & (!g2865)) + ((g27) & (!g2858) & (!g2860) & (g2853) & (g2865)) + ((g27) & (g2858) & (!g2860) & (!g2853) & (g2865)) + ((g27) & (g2858) & (g2860) & (!g2853) & (!g2865)) + ((g27) & (g2858) & (g2860) & (!g2853) & (g2865)) + ((g27) & (g2858) & (g2860) & (g2853) & (!g2865)) + ((g27) & (g2858) & (g2860) & (g2853) & (g2865)));
	assign g2970 = (((!g39) & (!g54) & (g2780) & (g2852)) + ((!g39) & (g54) & (!g2780) & (g2852)) + ((!g39) & (g54) & (g2780) & (!g2852)) + ((!g39) & (g54) & (g2780) & (g2852)) + ((g39) & (!g54) & (!g2780) & (!g2852)) + ((g39) & (!g54) & (!g2780) & (g2852)) + ((g39) & (!g54) & (g2780) & (!g2852)) + ((g39) & (g54) & (!g2780) & (!g2852)));
	assign g2971 = (((!g2859) & (!g2853) & (!g2865) & (g2970)) + ((!g2859) & (g2853) & (!g2865) & (g2970)) + ((!g2859) & (g2853) & (g2865) & (g2970)) + ((g2859) & (!g2853) & (!g2865) & (!g2970)) + ((g2859) & (!g2853) & (g2865) & (!g2970)) + ((g2859) & (!g2853) & (g2865) & (g2970)) + ((g2859) & (g2853) & (!g2865) & (!g2970)) + ((g2859) & (g2853) & (g2865) & (!g2970)));
	assign g2972 = (((!g27) & (!g39) & (g2971) & (g2866) & (g2964)) + ((!g27) & (g39) & (g2971) & (!g2866) & (g2964)) + ((!g27) & (g39) & (g2971) & (g2866) & (!g2964)) + ((!g27) & (g39) & (g2971) & (g2866) & (g2964)) + ((g27) & (!g39) & (!g2971) & (g2866) & (g2964)) + ((g27) & (!g39) & (g2971) & (!g2866) & (!g2964)) + ((g27) & (!g39) & (g2971) & (!g2866) & (g2964)) + ((g27) & (!g39) & (g2971) & (g2866) & (!g2964)) + ((g27) & (!g39) & (g2971) & (g2866) & (g2964)) + ((g27) & (g39) & (!g2971) & (!g2866) & (g2964)) + ((g27) & (g39) & (!g2971) & (g2866) & (!g2964)) + ((g27) & (g39) & (!g2971) & (g2866) & (g2964)) + ((g27) & (g39) & (g2971) & (!g2866) & (!g2964)) + ((g27) & (g39) & (g2971) & (!g2866) & (g2964)) + ((g27) & (g39) & (g2971) & (g2866) & (!g2964)) + ((g27) & (g39) & (g2971) & (g2866) & (g2964)));
	assign g2973 = (((!g8) & (!g18) & (g2968) & (g2969) & (g2972)) + ((!g8) & (g18) & (g2968) & (!g2969) & (g2972)) + ((!g8) & (g18) & (g2968) & (g2969) & (!g2972)) + ((!g8) & (g18) & (g2968) & (g2969) & (g2972)) + ((g8) & (!g18) & (!g2968) & (g2969) & (g2972)) + ((g8) & (!g18) & (g2968) & (!g2969) & (!g2972)) + ((g8) & (!g18) & (g2968) & (!g2969) & (g2972)) + ((g8) & (!g18) & (g2968) & (g2969) & (!g2972)) + ((g8) & (!g18) & (g2968) & (g2969) & (g2972)) + ((g8) & (g18) & (!g2968) & (!g2969) & (g2972)) + ((g8) & (g18) & (!g2968) & (g2969) & (!g2972)) + ((g8) & (g18) & (!g2968) & (g2969) & (g2972)) + ((g8) & (g18) & (g2968) & (!g2969) & (!g2972)) + ((g8) & (g18) & (g2968) & (!g2969) & (g2972)) + ((g8) & (g18) & (g2968) & (g2969) & (!g2972)) + ((g8) & (g18) & (g2968) & (g2969) & (g2972)));
	assign g2974 = (((!g2) & (!g8) & (g2856) & (g2861)) + ((!g2) & (g8) & (!g2856) & (g2861)) + ((!g2) & (g8) & (g2856) & (!g2861)) + ((!g2) & (g8) & (g2856) & (g2861)) + ((g2) & (!g8) & (!g2856) & (!g2861)) + ((g2) & (!g8) & (!g2856) & (g2861)) + ((g2) & (!g8) & (g2856) & (!g2861)) + ((g2) & (g8) & (!g2856) & (!g2861)));
	assign g2975 = (((!g2855) & (!g2853) & (!g2865) & (g2974)) + ((!g2855) & (g2853) & (!g2865) & (g2974)) + ((!g2855) & (g2853) & (g2865) & (g2974)) + ((g2855) & (!g2853) & (!g2865) & (!g2974)) + ((g2855) & (!g2853) & (g2865) & (!g2974)) + ((g2855) & (!g2853) & (g2865) & (g2974)) + ((g2855) & (g2853) & (!g2865) & (!g2974)) + ((g2855) & (g2853) & (g2865) & (!g2974)));
	assign g2976 = (((!g4) & (!g2) & (!g2966) & (!g2973) & (g2975)) + ((!g4) & (!g2) & (!g2966) & (g2973) & (g2975)) + ((!g4) & (!g2) & (g2966) & (!g2973) & (g2975)) + ((!g4) & (!g2) & (g2966) & (g2973) & (!g2975)) + ((!g4) & (!g2) & (g2966) & (g2973) & (g2975)) + ((!g4) & (g2) & (!g2966) & (!g2973) & (g2975)) + ((!g4) & (g2) & (!g2966) & (g2973) & (!g2975)) + ((!g4) & (g2) & (!g2966) & (g2973) & (g2975)) + ((!g4) & (g2) & (g2966) & (!g2973) & (!g2975)) + ((!g4) & (g2) & (g2966) & (!g2973) & (g2975)) + ((!g4) & (g2) & (g2966) & (g2973) & (!g2975)) + ((!g4) & (g2) & (g2966) & (g2973) & (g2975)) + ((g4) & (!g2) & (g2966) & (g2973) & (g2975)) + ((g4) & (g2) & (!g2966) & (g2973) & (g2975)) + ((g4) & (g2) & (g2966) & (!g2973) & (g2975)) + ((g4) & (g2) & (g2966) & (g2973) & (g2975)));
	assign g2977 = (((!g4) & (!g2862) & (g2863)) + ((!g4) & (g2862) & (!g2863)) + ((!g4) & (g2862) & (g2863)) + ((g4) & (g2862) & (g2863)));
	assign g2978 = (((!g2854) & (!g2977) & (!g2853) & (!g2865)) + ((!g2854) & (!g2977) & (g2853) & (!g2865)) + ((!g2854) & (!g2977) & (g2853) & (g2865)) + ((g2854) & (g2977) & (!g2853) & (!g2865)) + ((g2854) & (g2977) & (!g2853) & (g2865)) + ((g2854) & (g2977) & (g2853) & (!g2865)) + ((g2854) & (g2977) & (g2853) & (g2865)));
	assign g2979 = (((!g1) & (g2854) & (!g2977) & (!g2853) & (g2865)) + ((!g1) & (g2854) & (g2977) & (!g2853) & (g2865)) + ((g1) & (!g2854) & (g2977) & (g2853) & (!g2865)) + ((g1) & (!g2854) & (g2977) & (g2853) & (g2865)) + ((g1) & (g2854) & (!g2977) & (!g2853) & (!g2865)) + ((g1) & (g2854) & (!g2977) & (!g2853) & (g2865)) + ((g1) & (g2854) & (!g2977) & (g2853) & (!g2865)) + ((g1) & (g2854) & (!g2977) & (g2853) & (g2865)) + ((g1) & (g2854) & (g2977) & (!g2853) & (g2865)));
	assign g2980 = (((!g1) & (!g2965) & (!g2976) & (!g2978) & (!g2979)) + ((g1) & (!g2965) & (!g2976) & (!g2978) & (!g2979)) + ((g1) & (!g2965) & (!g2976) & (g2978) & (!g2979)) + ((g1) & (!g2965) & (g2976) & (!g2978) & (!g2979)) + ((g1) & (!g2965) & (g2976) & (g2978) & (!g2979)) + ((g1) & (g2965) & (!g2976) & (!g2978) & (!g2979)) + ((g1) & (g2965) & (!g2976) & (g2978) & (!g2979)));
	assign g2981 = (((!g39) & (!g2866) & (g2964) & (!g2980)) + ((!g39) & (g2866) & (!g2964) & (!g2980)) + ((!g39) & (g2866) & (!g2964) & (g2980)) + ((!g39) & (g2866) & (g2964) & (g2980)) + ((g39) & (!g2866) & (!g2964) & (!g2980)) + ((g39) & (g2866) & (!g2964) & (g2980)) + ((g39) & (g2866) & (g2964) & (!g2980)) + ((g39) & (g2866) & (g2964) & (g2980)));
	assign g2982 = (((!g54) & (!g68) & (!g2868) & (g2869) & (g2963) & (!g2980)) + ((!g54) & (!g68) & (g2868) & (!g2869) & (!g2963) & (!g2980)) + ((!g54) & (!g68) & (g2868) & (!g2869) & (!g2963) & (g2980)) + ((!g54) & (!g68) & (g2868) & (!g2869) & (g2963) & (!g2980)) + ((!g54) & (!g68) & (g2868) & (!g2869) & (g2963) & (g2980)) + ((!g54) & (!g68) & (g2868) & (g2869) & (!g2963) & (!g2980)) + ((!g54) & (!g68) & (g2868) & (g2869) & (!g2963) & (g2980)) + ((!g54) & (!g68) & (g2868) & (g2869) & (g2963) & (g2980)) + ((!g54) & (g68) & (!g2868) & (!g2869) & (g2963) & (!g2980)) + ((!g54) & (g68) & (!g2868) & (g2869) & (!g2963) & (!g2980)) + ((!g54) & (g68) & (!g2868) & (g2869) & (g2963) & (!g2980)) + ((!g54) & (g68) & (g2868) & (!g2869) & (!g2963) & (!g2980)) + ((!g54) & (g68) & (g2868) & (!g2869) & (!g2963) & (g2980)) + ((!g54) & (g68) & (g2868) & (!g2869) & (g2963) & (g2980)) + ((!g54) & (g68) & (g2868) & (g2869) & (!g2963) & (g2980)) + ((!g54) & (g68) & (g2868) & (g2869) & (g2963) & (g2980)) + ((g54) & (!g68) & (!g2868) & (!g2869) & (!g2963) & (!g2980)) + ((g54) & (!g68) & (!g2868) & (!g2869) & (g2963) & (!g2980)) + ((g54) & (!g68) & (!g2868) & (g2869) & (!g2963) & (!g2980)) + ((g54) & (!g68) & (g2868) & (!g2869) & (!g2963) & (g2980)) + ((g54) & (!g68) & (g2868) & (!g2869) & (g2963) & (g2980)) + ((g54) & (!g68) & (g2868) & (g2869) & (!g2963) & (g2980)) + ((g54) & (!g68) & (g2868) & (g2869) & (g2963) & (!g2980)) + ((g54) & (!g68) & (g2868) & (g2869) & (g2963) & (g2980)) + ((g54) & (g68) & (!g2868) & (!g2869) & (!g2963) & (!g2980)) + ((g54) & (g68) & (g2868) & (!g2869) & (!g2963) & (g2980)) + ((g54) & (g68) & (g2868) & (!g2869) & (g2963) & (!g2980)) + ((g54) & (g68) & (g2868) & (!g2869) & (g2963) & (g2980)) + ((g54) & (g68) & (g2868) & (g2869) & (!g2963) & (!g2980)) + ((g54) & (g68) & (g2868) & (g2869) & (!g2963) & (g2980)) + ((g54) & (g68) & (g2868) & (g2869) & (g2963) & (!g2980)) + ((g54) & (g68) & (g2868) & (g2869) & (g2963) & (g2980)));
	assign g2983 = (((!g68) & (!g2869) & (g2963) & (!g2980)) + ((!g68) & (g2869) & (!g2963) & (!g2980)) + ((!g68) & (g2869) & (!g2963) & (g2980)) + ((!g68) & (g2869) & (g2963) & (g2980)) + ((g68) & (!g2869) & (!g2963) & (!g2980)) + ((g68) & (g2869) & (!g2963) & (g2980)) + ((g68) & (g2869) & (g2963) & (!g2980)) + ((g68) & (g2869) & (g2963) & (g2980)));
	assign g2984 = (((!g87) & (!g104) & (!g2871) & (g2872) & (g2962) & (!g2980)) + ((!g87) & (!g104) & (g2871) & (!g2872) & (!g2962) & (!g2980)) + ((!g87) & (!g104) & (g2871) & (!g2872) & (!g2962) & (g2980)) + ((!g87) & (!g104) & (g2871) & (!g2872) & (g2962) & (!g2980)) + ((!g87) & (!g104) & (g2871) & (!g2872) & (g2962) & (g2980)) + ((!g87) & (!g104) & (g2871) & (g2872) & (!g2962) & (!g2980)) + ((!g87) & (!g104) & (g2871) & (g2872) & (!g2962) & (g2980)) + ((!g87) & (!g104) & (g2871) & (g2872) & (g2962) & (g2980)) + ((!g87) & (g104) & (!g2871) & (!g2872) & (g2962) & (!g2980)) + ((!g87) & (g104) & (!g2871) & (g2872) & (!g2962) & (!g2980)) + ((!g87) & (g104) & (!g2871) & (g2872) & (g2962) & (!g2980)) + ((!g87) & (g104) & (g2871) & (!g2872) & (!g2962) & (!g2980)) + ((!g87) & (g104) & (g2871) & (!g2872) & (!g2962) & (g2980)) + ((!g87) & (g104) & (g2871) & (!g2872) & (g2962) & (g2980)) + ((!g87) & (g104) & (g2871) & (g2872) & (!g2962) & (g2980)) + ((!g87) & (g104) & (g2871) & (g2872) & (g2962) & (g2980)) + ((g87) & (!g104) & (!g2871) & (!g2872) & (!g2962) & (!g2980)) + ((g87) & (!g104) & (!g2871) & (!g2872) & (g2962) & (!g2980)) + ((g87) & (!g104) & (!g2871) & (g2872) & (!g2962) & (!g2980)) + ((g87) & (!g104) & (g2871) & (!g2872) & (!g2962) & (g2980)) + ((g87) & (!g104) & (g2871) & (!g2872) & (g2962) & (g2980)) + ((g87) & (!g104) & (g2871) & (g2872) & (!g2962) & (g2980)) + ((g87) & (!g104) & (g2871) & (g2872) & (g2962) & (!g2980)) + ((g87) & (!g104) & (g2871) & (g2872) & (g2962) & (g2980)) + ((g87) & (g104) & (!g2871) & (!g2872) & (!g2962) & (!g2980)) + ((g87) & (g104) & (g2871) & (!g2872) & (!g2962) & (g2980)) + ((g87) & (g104) & (g2871) & (!g2872) & (g2962) & (!g2980)) + ((g87) & (g104) & (g2871) & (!g2872) & (g2962) & (g2980)) + ((g87) & (g104) & (g2871) & (g2872) & (!g2962) & (!g2980)) + ((g87) & (g104) & (g2871) & (g2872) & (!g2962) & (g2980)) + ((g87) & (g104) & (g2871) & (g2872) & (g2962) & (!g2980)) + ((g87) & (g104) & (g2871) & (g2872) & (g2962) & (g2980)));
	assign g2985 = (((!g104) & (!g2872) & (g2962) & (!g2980)) + ((!g104) & (g2872) & (!g2962) & (!g2980)) + ((!g104) & (g2872) & (!g2962) & (g2980)) + ((!g104) & (g2872) & (g2962) & (g2980)) + ((g104) & (!g2872) & (!g2962) & (!g2980)) + ((g104) & (g2872) & (!g2962) & (g2980)) + ((g104) & (g2872) & (g2962) & (!g2980)) + ((g104) & (g2872) & (g2962) & (g2980)));
	assign g2986 = (((!g127) & (!g147) & (!g2874) & (g2875) & (g2961) & (!g2980)) + ((!g127) & (!g147) & (g2874) & (!g2875) & (!g2961) & (!g2980)) + ((!g127) & (!g147) & (g2874) & (!g2875) & (!g2961) & (g2980)) + ((!g127) & (!g147) & (g2874) & (!g2875) & (g2961) & (!g2980)) + ((!g127) & (!g147) & (g2874) & (!g2875) & (g2961) & (g2980)) + ((!g127) & (!g147) & (g2874) & (g2875) & (!g2961) & (!g2980)) + ((!g127) & (!g147) & (g2874) & (g2875) & (!g2961) & (g2980)) + ((!g127) & (!g147) & (g2874) & (g2875) & (g2961) & (g2980)) + ((!g127) & (g147) & (!g2874) & (!g2875) & (g2961) & (!g2980)) + ((!g127) & (g147) & (!g2874) & (g2875) & (!g2961) & (!g2980)) + ((!g127) & (g147) & (!g2874) & (g2875) & (g2961) & (!g2980)) + ((!g127) & (g147) & (g2874) & (!g2875) & (!g2961) & (!g2980)) + ((!g127) & (g147) & (g2874) & (!g2875) & (!g2961) & (g2980)) + ((!g127) & (g147) & (g2874) & (!g2875) & (g2961) & (g2980)) + ((!g127) & (g147) & (g2874) & (g2875) & (!g2961) & (g2980)) + ((!g127) & (g147) & (g2874) & (g2875) & (g2961) & (g2980)) + ((g127) & (!g147) & (!g2874) & (!g2875) & (!g2961) & (!g2980)) + ((g127) & (!g147) & (!g2874) & (!g2875) & (g2961) & (!g2980)) + ((g127) & (!g147) & (!g2874) & (g2875) & (!g2961) & (!g2980)) + ((g127) & (!g147) & (g2874) & (!g2875) & (!g2961) & (g2980)) + ((g127) & (!g147) & (g2874) & (!g2875) & (g2961) & (g2980)) + ((g127) & (!g147) & (g2874) & (g2875) & (!g2961) & (g2980)) + ((g127) & (!g147) & (g2874) & (g2875) & (g2961) & (!g2980)) + ((g127) & (!g147) & (g2874) & (g2875) & (g2961) & (g2980)) + ((g127) & (g147) & (!g2874) & (!g2875) & (!g2961) & (!g2980)) + ((g127) & (g147) & (g2874) & (!g2875) & (!g2961) & (g2980)) + ((g127) & (g147) & (g2874) & (!g2875) & (g2961) & (!g2980)) + ((g127) & (g147) & (g2874) & (!g2875) & (g2961) & (g2980)) + ((g127) & (g147) & (g2874) & (g2875) & (!g2961) & (!g2980)) + ((g127) & (g147) & (g2874) & (g2875) & (!g2961) & (g2980)) + ((g127) & (g147) & (g2874) & (g2875) & (g2961) & (!g2980)) + ((g127) & (g147) & (g2874) & (g2875) & (g2961) & (g2980)));
	assign g2987 = (((!g147) & (!g2875) & (g2961) & (!g2980)) + ((!g147) & (g2875) & (!g2961) & (!g2980)) + ((!g147) & (g2875) & (!g2961) & (g2980)) + ((!g147) & (g2875) & (g2961) & (g2980)) + ((g147) & (!g2875) & (!g2961) & (!g2980)) + ((g147) & (g2875) & (!g2961) & (g2980)) + ((g147) & (g2875) & (g2961) & (!g2980)) + ((g147) & (g2875) & (g2961) & (g2980)));
	assign g2988 = (((!g174) & (!g198) & (!g2877) & (g2878) & (g2960) & (!g2980)) + ((!g174) & (!g198) & (g2877) & (!g2878) & (!g2960) & (!g2980)) + ((!g174) & (!g198) & (g2877) & (!g2878) & (!g2960) & (g2980)) + ((!g174) & (!g198) & (g2877) & (!g2878) & (g2960) & (!g2980)) + ((!g174) & (!g198) & (g2877) & (!g2878) & (g2960) & (g2980)) + ((!g174) & (!g198) & (g2877) & (g2878) & (!g2960) & (!g2980)) + ((!g174) & (!g198) & (g2877) & (g2878) & (!g2960) & (g2980)) + ((!g174) & (!g198) & (g2877) & (g2878) & (g2960) & (g2980)) + ((!g174) & (g198) & (!g2877) & (!g2878) & (g2960) & (!g2980)) + ((!g174) & (g198) & (!g2877) & (g2878) & (!g2960) & (!g2980)) + ((!g174) & (g198) & (!g2877) & (g2878) & (g2960) & (!g2980)) + ((!g174) & (g198) & (g2877) & (!g2878) & (!g2960) & (!g2980)) + ((!g174) & (g198) & (g2877) & (!g2878) & (!g2960) & (g2980)) + ((!g174) & (g198) & (g2877) & (!g2878) & (g2960) & (g2980)) + ((!g174) & (g198) & (g2877) & (g2878) & (!g2960) & (g2980)) + ((!g174) & (g198) & (g2877) & (g2878) & (g2960) & (g2980)) + ((g174) & (!g198) & (!g2877) & (!g2878) & (!g2960) & (!g2980)) + ((g174) & (!g198) & (!g2877) & (!g2878) & (g2960) & (!g2980)) + ((g174) & (!g198) & (!g2877) & (g2878) & (!g2960) & (!g2980)) + ((g174) & (!g198) & (g2877) & (!g2878) & (!g2960) & (g2980)) + ((g174) & (!g198) & (g2877) & (!g2878) & (g2960) & (g2980)) + ((g174) & (!g198) & (g2877) & (g2878) & (!g2960) & (g2980)) + ((g174) & (!g198) & (g2877) & (g2878) & (g2960) & (!g2980)) + ((g174) & (!g198) & (g2877) & (g2878) & (g2960) & (g2980)) + ((g174) & (g198) & (!g2877) & (!g2878) & (!g2960) & (!g2980)) + ((g174) & (g198) & (g2877) & (!g2878) & (!g2960) & (g2980)) + ((g174) & (g198) & (g2877) & (!g2878) & (g2960) & (!g2980)) + ((g174) & (g198) & (g2877) & (!g2878) & (g2960) & (g2980)) + ((g174) & (g198) & (g2877) & (g2878) & (!g2960) & (!g2980)) + ((g174) & (g198) & (g2877) & (g2878) & (!g2960) & (g2980)) + ((g174) & (g198) & (g2877) & (g2878) & (g2960) & (!g2980)) + ((g174) & (g198) & (g2877) & (g2878) & (g2960) & (g2980)));
	assign g2989 = (((!g198) & (!g2878) & (g2960) & (!g2980)) + ((!g198) & (g2878) & (!g2960) & (!g2980)) + ((!g198) & (g2878) & (!g2960) & (g2980)) + ((!g198) & (g2878) & (g2960) & (g2980)) + ((g198) & (!g2878) & (!g2960) & (!g2980)) + ((g198) & (g2878) & (!g2960) & (g2980)) + ((g198) & (g2878) & (g2960) & (!g2980)) + ((g198) & (g2878) & (g2960) & (g2980)));
	assign g2990 = (((!g229) & (!g255) & (!g2880) & (g2881) & (g2959) & (!g2980)) + ((!g229) & (!g255) & (g2880) & (!g2881) & (!g2959) & (!g2980)) + ((!g229) & (!g255) & (g2880) & (!g2881) & (!g2959) & (g2980)) + ((!g229) & (!g255) & (g2880) & (!g2881) & (g2959) & (!g2980)) + ((!g229) & (!g255) & (g2880) & (!g2881) & (g2959) & (g2980)) + ((!g229) & (!g255) & (g2880) & (g2881) & (!g2959) & (!g2980)) + ((!g229) & (!g255) & (g2880) & (g2881) & (!g2959) & (g2980)) + ((!g229) & (!g255) & (g2880) & (g2881) & (g2959) & (g2980)) + ((!g229) & (g255) & (!g2880) & (!g2881) & (g2959) & (!g2980)) + ((!g229) & (g255) & (!g2880) & (g2881) & (!g2959) & (!g2980)) + ((!g229) & (g255) & (!g2880) & (g2881) & (g2959) & (!g2980)) + ((!g229) & (g255) & (g2880) & (!g2881) & (!g2959) & (!g2980)) + ((!g229) & (g255) & (g2880) & (!g2881) & (!g2959) & (g2980)) + ((!g229) & (g255) & (g2880) & (!g2881) & (g2959) & (g2980)) + ((!g229) & (g255) & (g2880) & (g2881) & (!g2959) & (g2980)) + ((!g229) & (g255) & (g2880) & (g2881) & (g2959) & (g2980)) + ((g229) & (!g255) & (!g2880) & (!g2881) & (!g2959) & (!g2980)) + ((g229) & (!g255) & (!g2880) & (!g2881) & (g2959) & (!g2980)) + ((g229) & (!g255) & (!g2880) & (g2881) & (!g2959) & (!g2980)) + ((g229) & (!g255) & (g2880) & (!g2881) & (!g2959) & (g2980)) + ((g229) & (!g255) & (g2880) & (!g2881) & (g2959) & (g2980)) + ((g229) & (!g255) & (g2880) & (g2881) & (!g2959) & (g2980)) + ((g229) & (!g255) & (g2880) & (g2881) & (g2959) & (!g2980)) + ((g229) & (!g255) & (g2880) & (g2881) & (g2959) & (g2980)) + ((g229) & (g255) & (!g2880) & (!g2881) & (!g2959) & (!g2980)) + ((g229) & (g255) & (g2880) & (!g2881) & (!g2959) & (g2980)) + ((g229) & (g255) & (g2880) & (!g2881) & (g2959) & (!g2980)) + ((g229) & (g255) & (g2880) & (!g2881) & (g2959) & (g2980)) + ((g229) & (g255) & (g2880) & (g2881) & (!g2959) & (!g2980)) + ((g229) & (g255) & (g2880) & (g2881) & (!g2959) & (g2980)) + ((g229) & (g255) & (g2880) & (g2881) & (g2959) & (!g2980)) + ((g229) & (g255) & (g2880) & (g2881) & (g2959) & (g2980)));
	assign g2991 = (((!g255) & (!g2881) & (g2959) & (!g2980)) + ((!g255) & (g2881) & (!g2959) & (!g2980)) + ((!g255) & (g2881) & (!g2959) & (g2980)) + ((!g255) & (g2881) & (g2959) & (g2980)) + ((g255) & (!g2881) & (!g2959) & (!g2980)) + ((g255) & (g2881) & (!g2959) & (g2980)) + ((g255) & (g2881) & (g2959) & (!g2980)) + ((g255) & (g2881) & (g2959) & (g2980)));
	assign g2992 = (((!g290) & (!g319) & (!g2883) & (g2884) & (g2958) & (!g2980)) + ((!g290) & (!g319) & (g2883) & (!g2884) & (!g2958) & (!g2980)) + ((!g290) & (!g319) & (g2883) & (!g2884) & (!g2958) & (g2980)) + ((!g290) & (!g319) & (g2883) & (!g2884) & (g2958) & (!g2980)) + ((!g290) & (!g319) & (g2883) & (!g2884) & (g2958) & (g2980)) + ((!g290) & (!g319) & (g2883) & (g2884) & (!g2958) & (!g2980)) + ((!g290) & (!g319) & (g2883) & (g2884) & (!g2958) & (g2980)) + ((!g290) & (!g319) & (g2883) & (g2884) & (g2958) & (g2980)) + ((!g290) & (g319) & (!g2883) & (!g2884) & (g2958) & (!g2980)) + ((!g290) & (g319) & (!g2883) & (g2884) & (!g2958) & (!g2980)) + ((!g290) & (g319) & (!g2883) & (g2884) & (g2958) & (!g2980)) + ((!g290) & (g319) & (g2883) & (!g2884) & (!g2958) & (!g2980)) + ((!g290) & (g319) & (g2883) & (!g2884) & (!g2958) & (g2980)) + ((!g290) & (g319) & (g2883) & (!g2884) & (g2958) & (g2980)) + ((!g290) & (g319) & (g2883) & (g2884) & (!g2958) & (g2980)) + ((!g290) & (g319) & (g2883) & (g2884) & (g2958) & (g2980)) + ((g290) & (!g319) & (!g2883) & (!g2884) & (!g2958) & (!g2980)) + ((g290) & (!g319) & (!g2883) & (!g2884) & (g2958) & (!g2980)) + ((g290) & (!g319) & (!g2883) & (g2884) & (!g2958) & (!g2980)) + ((g290) & (!g319) & (g2883) & (!g2884) & (!g2958) & (g2980)) + ((g290) & (!g319) & (g2883) & (!g2884) & (g2958) & (g2980)) + ((g290) & (!g319) & (g2883) & (g2884) & (!g2958) & (g2980)) + ((g290) & (!g319) & (g2883) & (g2884) & (g2958) & (!g2980)) + ((g290) & (!g319) & (g2883) & (g2884) & (g2958) & (g2980)) + ((g290) & (g319) & (!g2883) & (!g2884) & (!g2958) & (!g2980)) + ((g290) & (g319) & (g2883) & (!g2884) & (!g2958) & (g2980)) + ((g290) & (g319) & (g2883) & (!g2884) & (g2958) & (!g2980)) + ((g290) & (g319) & (g2883) & (!g2884) & (g2958) & (g2980)) + ((g290) & (g319) & (g2883) & (g2884) & (!g2958) & (!g2980)) + ((g290) & (g319) & (g2883) & (g2884) & (!g2958) & (g2980)) + ((g290) & (g319) & (g2883) & (g2884) & (g2958) & (!g2980)) + ((g290) & (g319) & (g2883) & (g2884) & (g2958) & (g2980)));
	assign g2993 = (((!g319) & (!g2884) & (g2958) & (!g2980)) + ((!g319) & (g2884) & (!g2958) & (!g2980)) + ((!g319) & (g2884) & (!g2958) & (g2980)) + ((!g319) & (g2884) & (g2958) & (g2980)) + ((g319) & (!g2884) & (!g2958) & (!g2980)) + ((g319) & (g2884) & (!g2958) & (g2980)) + ((g319) & (g2884) & (g2958) & (!g2980)) + ((g319) & (g2884) & (g2958) & (g2980)));
	assign g2994 = (((!g358) & (!g390) & (!g2886) & (g2887) & (g2957) & (!g2980)) + ((!g358) & (!g390) & (g2886) & (!g2887) & (!g2957) & (!g2980)) + ((!g358) & (!g390) & (g2886) & (!g2887) & (!g2957) & (g2980)) + ((!g358) & (!g390) & (g2886) & (!g2887) & (g2957) & (!g2980)) + ((!g358) & (!g390) & (g2886) & (!g2887) & (g2957) & (g2980)) + ((!g358) & (!g390) & (g2886) & (g2887) & (!g2957) & (!g2980)) + ((!g358) & (!g390) & (g2886) & (g2887) & (!g2957) & (g2980)) + ((!g358) & (!g390) & (g2886) & (g2887) & (g2957) & (g2980)) + ((!g358) & (g390) & (!g2886) & (!g2887) & (g2957) & (!g2980)) + ((!g358) & (g390) & (!g2886) & (g2887) & (!g2957) & (!g2980)) + ((!g358) & (g390) & (!g2886) & (g2887) & (g2957) & (!g2980)) + ((!g358) & (g390) & (g2886) & (!g2887) & (!g2957) & (!g2980)) + ((!g358) & (g390) & (g2886) & (!g2887) & (!g2957) & (g2980)) + ((!g358) & (g390) & (g2886) & (!g2887) & (g2957) & (g2980)) + ((!g358) & (g390) & (g2886) & (g2887) & (!g2957) & (g2980)) + ((!g358) & (g390) & (g2886) & (g2887) & (g2957) & (g2980)) + ((g358) & (!g390) & (!g2886) & (!g2887) & (!g2957) & (!g2980)) + ((g358) & (!g390) & (!g2886) & (!g2887) & (g2957) & (!g2980)) + ((g358) & (!g390) & (!g2886) & (g2887) & (!g2957) & (!g2980)) + ((g358) & (!g390) & (g2886) & (!g2887) & (!g2957) & (g2980)) + ((g358) & (!g390) & (g2886) & (!g2887) & (g2957) & (g2980)) + ((g358) & (!g390) & (g2886) & (g2887) & (!g2957) & (g2980)) + ((g358) & (!g390) & (g2886) & (g2887) & (g2957) & (!g2980)) + ((g358) & (!g390) & (g2886) & (g2887) & (g2957) & (g2980)) + ((g358) & (g390) & (!g2886) & (!g2887) & (!g2957) & (!g2980)) + ((g358) & (g390) & (g2886) & (!g2887) & (!g2957) & (g2980)) + ((g358) & (g390) & (g2886) & (!g2887) & (g2957) & (!g2980)) + ((g358) & (g390) & (g2886) & (!g2887) & (g2957) & (g2980)) + ((g358) & (g390) & (g2886) & (g2887) & (!g2957) & (!g2980)) + ((g358) & (g390) & (g2886) & (g2887) & (!g2957) & (g2980)) + ((g358) & (g390) & (g2886) & (g2887) & (g2957) & (!g2980)) + ((g358) & (g390) & (g2886) & (g2887) & (g2957) & (g2980)));
	assign g2995 = (((!g390) & (!g2887) & (g2957) & (!g2980)) + ((!g390) & (g2887) & (!g2957) & (!g2980)) + ((!g390) & (g2887) & (!g2957) & (g2980)) + ((!g390) & (g2887) & (g2957) & (g2980)) + ((g390) & (!g2887) & (!g2957) & (!g2980)) + ((g390) & (g2887) & (!g2957) & (g2980)) + ((g390) & (g2887) & (g2957) & (!g2980)) + ((g390) & (g2887) & (g2957) & (g2980)));
	assign g2996 = (((!g433) & (!g468) & (!g2889) & (g2890) & (g2956) & (!g2980)) + ((!g433) & (!g468) & (g2889) & (!g2890) & (!g2956) & (!g2980)) + ((!g433) & (!g468) & (g2889) & (!g2890) & (!g2956) & (g2980)) + ((!g433) & (!g468) & (g2889) & (!g2890) & (g2956) & (!g2980)) + ((!g433) & (!g468) & (g2889) & (!g2890) & (g2956) & (g2980)) + ((!g433) & (!g468) & (g2889) & (g2890) & (!g2956) & (!g2980)) + ((!g433) & (!g468) & (g2889) & (g2890) & (!g2956) & (g2980)) + ((!g433) & (!g468) & (g2889) & (g2890) & (g2956) & (g2980)) + ((!g433) & (g468) & (!g2889) & (!g2890) & (g2956) & (!g2980)) + ((!g433) & (g468) & (!g2889) & (g2890) & (!g2956) & (!g2980)) + ((!g433) & (g468) & (!g2889) & (g2890) & (g2956) & (!g2980)) + ((!g433) & (g468) & (g2889) & (!g2890) & (!g2956) & (!g2980)) + ((!g433) & (g468) & (g2889) & (!g2890) & (!g2956) & (g2980)) + ((!g433) & (g468) & (g2889) & (!g2890) & (g2956) & (g2980)) + ((!g433) & (g468) & (g2889) & (g2890) & (!g2956) & (g2980)) + ((!g433) & (g468) & (g2889) & (g2890) & (g2956) & (g2980)) + ((g433) & (!g468) & (!g2889) & (!g2890) & (!g2956) & (!g2980)) + ((g433) & (!g468) & (!g2889) & (!g2890) & (g2956) & (!g2980)) + ((g433) & (!g468) & (!g2889) & (g2890) & (!g2956) & (!g2980)) + ((g433) & (!g468) & (g2889) & (!g2890) & (!g2956) & (g2980)) + ((g433) & (!g468) & (g2889) & (!g2890) & (g2956) & (g2980)) + ((g433) & (!g468) & (g2889) & (g2890) & (!g2956) & (g2980)) + ((g433) & (!g468) & (g2889) & (g2890) & (g2956) & (!g2980)) + ((g433) & (!g468) & (g2889) & (g2890) & (g2956) & (g2980)) + ((g433) & (g468) & (!g2889) & (!g2890) & (!g2956) & (!g2980)) + ((g433) & (g468) & (g2889) & (!g2890) & (!g2956) & (g2980)) + ((g433) & (g468) & (g2889) & (!g2890) & (g2956) & (!g2980)) + ((g433) & (g468) & (g2889) & (!g2890) & (g2956) & (g2980)) + ((g433) & (g468) & (g2889) & (g2890) & (!g2956) & (!g2980)) + ((g433) & (g468) & (g2889) & (g2890) & (!g2956) & (g2980)) + ((g433) & (g468) & (g2889) & (g2890) & (g2956) & (!g2980)) + ((g433) & (g468) & (g2889) & (g2890) & (g2956) & (g2980)));
	assign g2997 = (((!g468) & (!g2890) & (g2956) & (!g2980)) + ((!g468) & (g2890) & (!g2956) & (!g2980)) + ((!g468) & (g2890) & (!g2956) & (g2980)) + ((!g468) & (g2890) & (g2956) & (g2980)) + ((g468) & (!g2890) & (!g2956) & (!g2980)) + ((g468) & (g2890) & (!g2956) & (g2980)) + ((g468) & (g2890) & (g2956) & (!g2980)) + ((g468) & (g2890) & (g2956) & (g2980)));
	assign g2998 = (((!g515) & (!g553) & (!g2892) & (g2893) & (g2955) & (!g2980)) + ((!g515) & (!g553) & (g2892) & (!g2893) & (!g2955) & (!g2980)) + ((!g515) & (!g553) & (g2892) & (!g2893) & (!g2955) & (g2980)) + ((!g515) & (!g553) & (g2892) & (!g2893) & (g2955) & (!g2980)) + ((!g515) & (!g553) & (g2892) & (!g2893) & (g2955) & (g2980)) + ((!g515) & (!g553) & (g2892) & (g2893) & (!g2955) & (!g2980)) + ((!g515) & (!g553) & (g2892) & (g2893) & (!g2955) & (g2980)) + ((!g515) & (!g553) & (g2892) & (g2893) & (g2955) & (g2980)) + ((!g515) & (g553) & (!g2892) & (!g2893) & (g2955) & (!g2980)) + ((!g515) & (g553) & (!g2892) & (g2893) & (!g2955) & (!g2980)) + ((!g515) & (g553) & (!g2892) & (g2893) & (g2955) & (!g2980)) + ((!g515) & (g553) & (g2892) & (!g2893) & (!g2955) & (!g2980)) + ((!g515) & (g553) & (g2892) & (!g2893) & (!g2955) & (g2980)) + ((!g515) & (g553) & (g2892) & (!g2893) & (g2955) & (g2980)) + ((!g515) & (g553) & (g2892) & (g2893) & (!g2955) & (g2980)) + ((!g515) & (g553) & (g2892) & (g2893) & (g2955) & (g2980)) + ((g515) & (!g553) & (!g2892) & (!g2893) & (!g2955) & (!g2980)) + ((g515) & (!g553) & (!g2892) & (!g2893) & (g2955) & (!g2980)) + ((g515) & (!g553) & (!g2892) & (g2893) & (!g2955) & (!g2980)) + ((g515) & (!g553) & (g2892) & (!g2893) & (!g2955) & (g2980)) + ((g515) & (!g553) & (g2892) & (!g2893) & (g2955) & (g2980)) + ((g515) & (!g553) & (g2892) & (g2893) & (!g2955) & (g2980)) + ((g515) & (!g553) & (g2892) & (g2893) & (g2955) & (!g2980)) + ((g515) & (!g553) & (g2892) & (g2893) & (g2955) & (g2980)) + ((g515) & (g553) & (!g2892) & (!g2893) & (!g2955) & (!g2980)) + ((g515) & (g553) & (g2892) & (!g2893) & (!g2955) & (g2980)) + ((g515) & (g553) & (g2892) & (!g2893) & (g2955) & (!g2980)) + ((g515) & (g553) & (g2892) & (!g2893) & (g2955) & (g2980)) + ((g515) & (g553) & (g2892) & (g2893) & (!g2955) & (!g2980)) + ((g515) & (g553) & (g2892) & (g2893) & (!g2955) & (g2980)) + ((g515) & (g553) & (g2892) & (g2893) & (g2955) & (!g2980)) + ((g515) & (g553) & (g2892) & (g2893) & (g2955) & (g2980)));
	assign g2999 = (((!g553) & (!g2893) & (g2955) & (!g2980)) + ((!g553) & (g2893) & (!g2955) & (!g2980)) + ((!g553) & (g2893) & (!g2955) & (g2980)) + ((!g553) & (g2893) & (g2955) & (g2980)) + ((g553) & (!g2893) & (!g2955) & (!g2980)) + ((g553) & (g2893) & (!g2955) & (g2980)) + ((g553) & (g2893) & (g2955) & (!g2980)) + ((g553) & (g2893) & (g2955) & (g2980)));
	assign g3000 = (((!g604) & (!g645) & (!g2895) & (g2896) & (g2954) & (!g2980)) + ((!g604) & (!g645) & (g2895) & (!g2896) & (!g2954) & (!g2980)) + ((!g604) & (!g645) & (g2895) & (!g2896) & (!g2954) & (g2980)) + ((!g604) & (!g645) & (g2895) & (!g2896) & (g2954) & (!g2980)) + ((!g604) & (!g645) & (g2895) & (!g2896) & (g2954) & (g2980)) + ((!g604) & (!g645) & (g2895) & (g2896) & (!g2954) & (!g2980)) + ((!g604) & (!g645) & (g2895) & (g2896) & (!g2954) & (g2980)) + ((!g604) & (!g645) & (g2895) & (g2896) & (g2954) & (g2980)) + ((!g604) & (g645) & (!g2895) & (!g2896) & (g2954) & (!g2980)) + ((!g604) & (g645) & (!g2895) & (g2896) & (!g2954) & (!g2980)) + ((!g604) & (g645) & (!g2895) & (g2896) & (g2954) & (!g2980)) + ((!g604) & (g645) & (g2895) & (!g2896) & (!g2954) & (!g2980)) + ((!g604) & (g645) & (g2895) & (!g2896) & (!g2954) & (g2980)) + ((!g604) & (g645) & (g2895) & (!g2896) & (g2954) & (g2980)) + ((!g604) & (g645) & (g2895) & (g2896) & (!g2954) & (g2980)) + ((!g604) & (g645) & (g2895) & (g2896) & (g2954) & (g2980)) + ((g604) & (!g645) & (!g2895) & (!g2896) & (!g2954) & (!g2980)) + ((g604) & (!g645) & (!g2895) & (!g2896) & (g2954) & (!g2980)) + ((g604) & (!g645) & (!g2895) & (g2896) & (!g2954) & (!g2980)) + ((g604) & (!g645) & (g2895) & (!g2896) & (!g2954) & (g2980)) + ((g604) & (!g645) & (g2895) & (!g2896) & (g2954) & (g2980)) + ((g604) & (!g645) & (g2895) & (g2896) & (!g2954) & (g2980)) + ((g604) & (!g645) & (g2895) & (g2896) & (g2954) & (!g2980)) + ((g604) & (!g645) & (g2895) & (g2896) & (g2954) & (g2980)) + ((g604) & (g645) & (!g2895) & (!g2896) & (!g2954) & (!g2980)) + ((g604) & (g645) & (g2895) & (!g2896) & (!g2954) & (g2980)) + ((g604) & (g645) & (g2895) & (!g2896) & (g2954) & (!g2980)) + ((g604) & (g645) & (g2895) & (!g2896) & (g2954) & (g2980)) + ((g604) & (g645) & (g2895) & (g2896) & (!g2954) & (!g2980)) + ((g604) & (g645) & (g2895) & (g2896) & (!g2954) & (g2980)) + ((g604) & (g645) & (g2895) & (g2896) & (g2954) & (!g2980)) + ((g604) & (g645) & (g2895) & (g2896) & (g2954) & (g2980)));
	assign g3001 = (((!g645) & (!g2896) & (g2954) & (!g2980)) + ((!g645) & (g2896) & (!g2954) & (!g2980)) + ((!g645) & (g2896) & (!g2954) & (g2980)) + ((!g645) & (g2896) & (g2954) & (g2980)) + ((g645) & (!g2896) & (!g2954) & (!g2980)) + ((g645) & (g2896) & (!g2954) & (g2980)) + ((g645) & (g2896) & (g2954) & (!g2980)) + ((g645) & (g2896) & (g2954) & (g2980)));
	assign g3002 = (((!g700) & (!g744) & (!g2898) & (g2899) & (g2953) & (!g2980)) + ((!g700) & (!g744) & (g2898) & (!g2899) & (!g2953) & (!g2980)) + ((!g700) & (!g744) & (g2898) & (!g2899) & (!g2953) & (g2980)) + ((!g700) & (!g744) & (g2898) & (!g2899) & (g2953) & (!g2980)) + ((!g700) & (!g744) & (g2898) & (!g2899) & (g2953) & (g2980)) + ((!g700) & (!g744) & (g2898) & (g2899) & (!g2953) & (!g2980)) + ((!g700) & (!g744) & (g2898) & (g2899) & (!g2953) & (g2980)) + ((!g700) & (!g744) & (g2898) & (g2899) & (g2953) & (g2980)) + ((!g700) & (g744) & (!g2898) & (!g2899) & (g2953) & (!g2980)) + ((!g700) & (g744) & (!g2898) & (g2899) & (!g2953) & (!g2980)) + ((!g700) & (g744) & (!g2898) & (g2899) & (g2953) & (!g2980)) + ((!g700) & (g744) & (g2898) & (!g2899) & (!g2953) & (!g2980)) + ((!g700) & (g744) & (g2898) & (!g2899) & (!g2953) & (g2980)) + ((!g700) & (g744) & (g2898) & (!g2899) & (g2953) & (g2980)) + ((!g700) & (g744) & (g2898) & (g2899) & (!g2953) & (g2980)) + ((!g700) & (g744) & (g2898) & (g2899) & (g2953) & (g2980)) + ((g700) & (!g744) & (!g2898) & (!g2899) & (!g2953) & (!g2980)) + ((g700) & (!g744) & (!g2898) & (!g2899) & (g2953) & (!g2980)) + ((g700) & (!g744) & (!g2898) & (g2899) & (!g2953) & (!g2980)) + ((g700) & (!g744) & (g2898) & (!g2899) & (!g2953) & (g2980)) + ((g700) & (!g744) & (g2898) & (!g2899) & (g2953) & (g2980)) + ((g700) & (!g744) & (g2898) & (g2899) & (!g2953) & (g2980)) + ((g700) & (!g744) & (g2898) & (g2899) & (g2953) & (!g2980)) + ((g700) & (!g744) & (g2898) & (g2899) & (g2953) & (g2980)) + ((g700) & (g744) & (!g2898) & (!g2899) & (!g2953) & (!g2980)) + ((g700) & (g744) & (g2898) & (!g2899) & (!g2953) & (g2980)) + ((g700) & (g744) & (g2898) & (!g2899) & (g2953) & (!g2980)) + ((g700) & (g744) & (g2898) & (!g2899) & (g2953) & (g2980)) + ((g700) & (g744) & (g2898) & (g2899) & (!g2953) & (!g2980)) + ((g700) & (g744) & (g2898) & (g2899) & (!g2953) & (g2980)) + ((g700) & (g744) & (g2898) & (g2899) & (g2953) & (!g2980)) + ((g700) & (g744) & (g2898) & (g2899) & (g2953) & (g2980)));
	assign g3003 = (((!g744) & (!g2899) & (g2953) & (!g2980)) + ((!g744) & (g2899) & (!g2953) & (!g2980)) + ((!g744) & (g2899) & (!g2953) & (g2980)) + ((!g744) & (g2899) & (g2953) & (g2980)) + ((g744) & (!g2899) & (!g2953) & (!g2980)) + ((g744) & (g2899) & (!g2953) & (g2980)) + ((g744) & (g2899) & (g2953) & (!g2980)) + ((g744) & (g2899) & (g2953) & (g2980)));
	assign g3004 = (((!g803) & (!g851) & (!g2901) & (g2902) & (g2952) & (!g2980)) + ((!g803) & (!g851) & (g2901) & (!g2902) & (!g2952) & (!g2980)) + ((!g803) & (!g851) & (g2901) & (!g2902) & (!g2952) & (g2980)) + ((!g803) & (!g851) & (g2901) & (!g2902) & (g2952) & (!g2980)) + ((!g803) & (!g851) & (g2901) & (!g2902) & (g2952) & (g2980)) + ((!g803) & (!g851) & (g2901) & (g2902) & (!g2952) & (!g2980)) + ((!g803) & (!g851) & (g2901) & (g2902) & (!g2952) & (g2980)) + ((!g803) & (!g851) & (g2901) & (g2902) & (g2952) & (g2980)) + ((!g803) & (g851) & (!g2901) & (!g2902) & (g2952) & (!g2980)) + ((!g803) & (g851) & (!g2901) & (g2902) & (!g2952) & (!g2980)) + ((!g803) & (g851) & (!g2901) & (g2902) & (g2952) & (!g2980)) + ((!g803) & (g851) & (g2901) & (!g2902) & (!g2952) & (!g2980)) + ((!g803) & (g851) & (g2901) & (!g2902) & (!g2952) & (g2980)) + ((!g803) & (g851) & (g2901) & (!g2902) & (g2952) & (g2980)) + ((!g803) & (g851) & (g2901) & (g2902) & (!g2952) & (g2980)) + ((!g803) & (g851) & (g2901) & (g2902) & (g2952) & (g2980)) + ((g803) & (!g851) & (!g2901) & (!g2902) & (!g2952) & (!g2980)) + ((g803) & (!g851) & (!g2901) & (!g2902) & (g2952) & (!g2980)) + ((g803) & (!g851) & (!g2901) & (g2902) & (!g2952) & (!g2980)) + ((g803) & (!g851) & (g2901) & (!g2902) & (!g2952) & (g2980)) + ((g803) & (!g851) & (g2901) & (!g2902) & (g2952) & (g2980)) + ((g803) & (!g851) & (g2901) & (g2902) & (!g2952) & (g2980)) + ((g803) & (!g851) & (g2901) & (g2902) & (g2952) & (!g2980)) + ((g803) & (!g851) & (g2901) & (g2902) & (g2952) & (g2980)) + ((g803) & (g851) & (!g2901) & (!g2902) & (!g2952) & (!g2980)) + ((g803) & (g851) & (g2901) & (!g2902) & (!g2952) & (g2980)) + ((g803) & (g851) & (g2901) & (!g2902) & (g2952) & (!g2980)) + ((g803) & (g851) & (g2901) & (!g2902) & (g2952) & (g2980)) + ((g803) & (g851) & (g2901) & (g2902) & (!g2952) & (!g2980)) + ((g803) & (g851) & (g2901) & (g2902) & (!g2952) & (g2980)) + ((g803) & (g851) & (g2901) & (g2902) & (g2952) & (!g2980)) + ((g803) & (g851) & (g2901) & (g2902) & (g2952) & (g2980)));
	assign g3005 = (((!g851) & (!g2902) & (g2952) & (!g2980)) + ((!g851) & (g2902) & (!g2952) & (!g2980)) + ((!g851) & (g2902) & (!g2952) & (g2980)) + ((!g851) & (g2902) & (g2952) & (g2980)) + ((g851) & (!g2902) & (!g2952) & (!g2980)) + ((g851) & (g2902) & (!g2952) & (g2980)) + ((g851) & (g2902) & (g2952) & (!g2980)) + ((g851) & (g2902) & (g2952) & (g2980)));
	assign g3006 = (((!g914) & (!g1032) & (!g2904) & (g2905) & (g2951) & (!g2980)) + ((!g914) & (!g1032) & (g2904) & (!g2905) & (!g2951) & (!g2980)) + ((!g914) & (!g1032) & (g2904) & (!g2905) & (!g2951) & (g2980)) + ((!g914) & (!g1032) & (g2904) & (!g2905) & (g2951) & (!g2980)) + ((!g914) & (!g1032) & (g2904) & (!g2905) & (g2951) & (g2980)) + ((!g914) & (!g1032) & (g2904) & (g2905) & (!g2951) & (!g2980)) + ((!g914) & (!g1032) & (g2904) & (g2905) & (!g2951) & (g2980)) + ((!g914) & (!g1032) & (g2904) & (g2905) & (g2951) & (g2980)) + ((!g914) & (g1032) & (!g2904) & (!g2905) & (g2951) & (!g2980)) + ((!g914) & (g1032) & (!g2904) & (g2905) & (!g2951) & (!g2980)) + ((!g914) & (g1032) & (!g2904) & (g2905) & (g2951) & (!g2980)) + ((!g914) & (g1032) & (g2904) & (!g2905) & (!g2951) & (!g2980)) + ((!g914) & (g1032) & (g2904) & (!g2905) & (!g2951) & (g2980)) + ((!g914) & (g1032) & (g2904) & (!g2905) & (g2951) & (g2980)) + ((!g914) & (g1032) & (g2904) & (g2905) & (!g2951) & (g2980)) + ((!g914) & (g1032) & (g2904) & (g2905) & (g2951) & (g2980)) + ((g914) & (!g1032) & (!g2904) & (!g2905) & (!g2951) & (!g2980)) + ((g914) & (!g1032) & (!g2904) & (!g2905) & (g2951) & (!g2980)) + ((g914) & (!g1032) & (!g2904) & (g2905) & (!g2951) & (!g2980)) + ((g914) & (!g1032) & (g2904) & (!g2905) & (!g2951) & (g2980)) + ((g914) & (!g1032) & (g2904) & (!g2905) & (g2951) & (g2980)) + ((g914) & (!g1032) & (g2904) & (g2905) & (!g2951) & (g2980)) + ((g914) & (!g1032) & (g2904) & (g2905) & (g2951) & (!g2980)) + ((g914) & (!g1032) & (g2904) & (g2905) & (g2951) & (g2980)) + ((g914) & (g1032) & (!g2904) & (!g2905) & (!g2951) & (!g2980)) + ((g914) & (g1032) & (g2904) & (!g2905) & (!g2951) & (g2980)) + ((g914) & (g1032) & (g2904) & (!g2905) & (g2951) & (!g2980)) + ((g914) & (g1032) & (g2904) & (!g2905) & (g2951) & (g2980)) + ((g914) & (g1032) & (g2904) & (g2905) & (!g2951) & (!g2980)) + ((g914) & (g1032) & (g2904) & (g2905) & (!g2951) & (g2980)) + ((g914) & (g1032) & (g2904) & (g2905) & (g2951) & (!g2980)) + ((g914) & (g1032) & (g2904) & (g2905) & (g2951) & (g2980)));
	assign g3007 = (((!g1032) & (!g2905) & (g2951) & (!g2980)) + ((!g1032) & (g2905) & (!g2951) & (!g2980)) + ((!g1032) & (g2905) & (!g2951) & (g2980)) + ((!g1032) & (g2905) & (g2951) & (g2980)) + ((g1032) & (!g2905) & (!g2951) & (!g2980)) + ((g1032) & (g2905) & (!g2951) & (g2980)) + ((g1032) & (g2905) & (g2951) & (!g2980)) + ((g1032) & (g2905) & (g2951) & (g2980)));
	assign g3008 = (((!g1030) & (!g1160) & (!g2907) & (g2908) & (g2950) & (!g2980)) + ((!g1030) & (!g1160) & (g2907) & (!g2908) & (!g2950) & (!g2980)) + ((!g1030) & (!g1160) & (g2907) & (!g2908) & (!g2950) & (g2980)) + ((!g1030) & (!g1160) & (g2907) & (!g2908) & (g2950) & (!g2980)) + ((!g1030) & (!g1160) & (g2907) & (!g2908) & (g2950) & (g2980)) + ((!g1030) & (!g1160) & (g2907) & (g2908) & (!g2950) & (!g2980)) + ((!g1030) & (!g1160) & (g2907) & (g2908) & (!g2950) & (g2980)) + ((!g1030) & (!g1160) & (g2907) & (g2908) & (g2950) & (g2980)) + ((!g1030) & (g1160) & (!g2907) & (!g2908) & (g2950) & (!g2980)) + ((!g1030) & (g1160) & (!g2907) & (g2908) & (!g2950) & (!g2980)) + ((!g1030) & (g1160) & (!g2907) & (g2908) & (g2950) & (!g2980)) + ((!g1030) & (g1160) & (g2907) & (!g2908) & (!g2950) & (!g2980)) + ((!g1030) & (g1160) & (g2907) & (!g2908) & (!g2950) & (g2980)) + ((!g1030) & (g1160) & (g2907) & (!g2908) & (g2950) & (g2980)) + ((!g1030) & (g1160) & (g2907) & (g2908) & (!g2950) & (g2980)) + ((!g1030) & (g1160) & (g2907) & (g2908) & (g2950) & (g2980)) + ((g1030) & (!g1160) & (!g2907) & (!g2908) & (!g2950) & (!g2980)) + ((g1030) & (!g1160) & (!g2907) & (!g2908) & (g2950) & (!g2980)) + ((g1030) & (!g1160) & (!g2907) & (g2908) & (!g2950) & (!g2980)) + ((g1030) & (!g1160) & (g2907) & (!g2908) & (!g2950) & (g2980)) + ((g1030) & (!g1160) & (g2907) & (!g2908) & (g2950) & (g2980)) + ((g1030) & (!g1160) & (g2907) & (g2908) & (!g2950) & (g2980)) + ((g1030) & (!g1160) & (g2907) & (g2908) & (g2950) & (!g2980)) + ((g1030) & (!g1160) & (g2907) & (g2908) & (g2950) & (g2980)) + ((g1030) & (g1160) & (!g2907) & (!g2908) & (!g2950) & (!g2980)) + ((g1030) & (g1160) & (g2907) & (!g2908) & (!g2950) & (g2980)) + ((g1030) & (g1160) & (g2907) & (!g2908) & (g2950) & (!g2980)) + ((g1030) & (g1160) & (g2907) & (!g2908) & (g2950) & (g2980)) + ((g1030) & (g1160) & (g2907) & (g2908) & (!g2950) & (!g2980)) + ((g1030) & (g1160) & (g2907) & (g2908) & (!g2950) & (g2980)) + ((g1030) & (g1160) & (g2907) & (g2908) & (g2950) & (!g2980)) + ((g1030) & (g1160) & (g2907) & (g2908) & (g2950) & (g2980)));
	assign g3009 = (((!g1160) & (!g2908) & (g2950) & (!g2980)) + ((!g1160) & (g2908) & (!g2950) & (!g2980)) + ((!g1160) & (g2908) & (!g2950) & (g2980)) + ((!g1160) & (g2908) & (g2950) & (g2980)) + ((g1160) & (!g2908) & (!g2950) & (!g2980)) + ((g1160) & (g2908) & (!g2950) & (g2980)) + ((g1160) & (g2908) & (g2950) & (!g2980)) + ((g1160) & (g2908) & (g2950) & (g2980)));
	assign g3010 = (((!g1154) & (!g1295) & (!g2910) & (g2911) & (g2949) & (!g2980)) + ((!g1154) & (!g1295) & (g2910) & (!g2911) & (!g2949) & (!g2980)) + ((!g1154) & (!g1295) & (g2910) & (!g2911) & (!g2949) & (g2980)) + ((!g1154) & (!g1295) & (g2910) & (!g2911) & (g2949) & (!g2980)) + ((!g1154) & (!g1295) & (g2910) & (!g2911) & (g2949) & (g2980)) + ((!g1154) & (!g1295) & (g2910) & (g2911) & (!g2949) & (!g2980)) + ((!g1154) & (!g1295) & (g2910) & (g2911) & (!g2949) & (g2980)) + ((!g1154) & (!g1295) & (g2910) & (g2911) & (g2949) & (g2980)) + ((!g1154) & (g1295) & (!g2910) & (!g2911) & (g2949) & (!g2980)) + ((!g1154) & (g1295) & (!g2910) & (g2911) & (!g2949) & (!g2980)) + ((!g1154) & (g1295) & (!g2910) & (g2911) & (g2949) & (!g2980)) + ((!g1154) & (g1295) & (g2910) & (!g2911) & (!g2949) & (!g2980)) + ((!g1154) & (g1295) & (g2910) & (!g2911) & (!g2949) & (g2980)) + ((!g1154) & (g1295) & (g2910) & (!g2911) & (g2949) & (g2980)) + ((!g1154) & (g1295) & (g2910) & (g2911) & (!g2949) & (g2980)) + ((!g1154) & (g1295) & (g2910) & (g2911) & (g2949) & (g2980)) + ((g1154) & (!g1295) & (!g2910) & (!g2911) & (!g2949) & (!g2980)) + ((g1154) & (!g1295) & (!g2910) & (!g2911) & (g2949) & (!g2980)) + ((g1154) & (!g1295) & (!g2910) & (g2911) & (!g2949) & (!g2980)) + ((g1154) & (!g1295) & (g2910) & (!g2911) & (!g2949) & (g2980)) + ((g1154) & (!g1295) & (g2910) & (!g2911) & (g2949) & (g2980)) + ((g1154) & (!g1295) & (g2910) & (g2911) & (!g2949) & (g2980)) + ((g1154) & (!g1295) & (g2910) & (g2911) & (g2949) & (!g2980)) + ((g1154) & (!g1295) & (g2910) & (g2911) & (g2949) & (g2980)) + ((g1154) & (g1295) & (!g2910) & (!g2911) & (!g2949) & (!g2980)) + ((g1154) & (g1295) & (g2910) & (!g2911) & (!g2949) & (g2980)) + ((g1154) & (g1295) & (g2910) & (!g2911) & (g2949) & (!g2980)) + ((g1154) & (g1295) & (g2910) & (!g2911) & (g2949) & (g2980)) + ((g1154) & (g1295) & (g2910) & (g2911) & (!g2949) & (!g2980)) + ((g1154) & (g1295) & (g2910) & (g2911) & (!g2949) & (g2980)) + ((g1154) & (g1295) & (g2910) & (g2911) & (g2949) & (!g2980)) + ((g1154) & (g1295) & (g2910) & (g2911) & (g2949) & (g2980)));
	assign g3011 = (((!g1295) & (!g2911) & (g2949) & (!g2980)) + ((!g1295) & (g2911) & (!g2949) & (!g2980)) + ((!g1295) & (g2911) & (!g2949) & (g2980)) + ((!g1295) & (g2911) & (g2949) & (g2980)) + ((g1295) & (!g2911) & (!g2949) & (!g2980)) + ((g1295) & (g2911) & (!g2949) & (g2980)) + ((g1295) & (g2911) & (g2949) & (!g2980)) + ((g1295) & (g2911) & (g2949) & (g2980)));
	assign g3012 = (((!g1285) & (!g1437) & (!g2913) & (g2914) & (g2948) & (!g2980)) + ((!g1285) & (!g1437) & (g2913) & (!g2914) & (!g2948) & (!g2980)) + ((!g1285) & (!g1437) & (g2913) & (!g2914) & (!g2948) & (g2980)) + ((!g1285) & (!g1437) & (g2913) & (!g2914) & (g2948) & (!g2980)) + ((!g1285) & (!g1437) & (g2913) & (!g2914) & (g2948) & (g2980)) + ((!g1285) & (!g1437) & (g2913) & (g2914) & (!g2948) & (!g2980)) + ((!g1285) & (!g1437) & (g2913) & (g2914) & (!g2948) & (g2980)) + ((!g1285) & (!g1437) & (g2913) & (g2914) & (g2948) & (g2980)) + ((!g1285) & (g1437) & (!g2913) & (!g2914) & (g2948) & (!g2980)) + ((!g1285) & (g1437) & (!g2913) & (g2914) & (!g2948) & (!g2980)) + ((!g1285) & (g1437) & (!g2913) & (g2914) & (g2948) & (!g2980)) + ((!g1285) & (g1437) & (g2913) & (!g2914) & (!g2948) & (!g2980)) + ((!g1285) & (g1437) & (g2913) & (!g2914) & (!g2948) & (g2980)) + ((!g1285) & (g1437) & (g2913) & (!g2914) & (g2948) & (g2980)) + ((!g1285) & (g1437) & (g2913) & (g2914) & (!g2948) & (g2980)) + ((!g1285) & (g1437) & (g2913) & (g2914) & (g2948) & (g2980)) + ((g1285) & (!g1437) & (!g2913) & (!g2914) & (!g2948) & (!g2980)) + ((g1285) & (!g1437) & (!g2913) & (!g2914) & (g2948) & (!g2980)) + ((g1285) & (!g1437) & (!g2913) & (g2914) & (!g2948) & (!g2980)) + ((g1285) & (!g1437) & (g2913) & (!g2914) & (!g2948) & (g2980)) + ((g1285) & (!g1437) & (g2913) & (!g2914) & (g2948) & (g2980)) + ((g1285) & (!g1437) & (g2913) & (g2914) & (!g2948) & (g2980)) + ((g1285) & (!g1437) & (g2913) & (g2914) & (g2948) & (!g2980)) + ((g1285) & (!g1437) & (g2913) & (g2914) & (g2948) & (g2980)) + ((g1285) & (g1437) & (!g2913) & (!g2914) & (!g2948) & (!g2980)) + ((g1285) & (g1437) & (g2913) & (!g2914) & (!g2948) & (g2980)) + ((g1285) & (g1437) & (g2913) & (!g2914) & (g2948) & (!g2980)) + ((g1285) & (g1437) & (g2913) & (!g2914) & (g2948) & (g2980)) + ((g1285) & (g1437) & (g2913) & (g2914) & (!g2948) & (!g2980)) + ((g1285) & (g1437) & (g2913) & (g2914) & (!g2948) & (g2980)) + ((g1285) & (g1437) & (g2913) & (g2914) & (g2948) & (!g2980)) + ((g1285) & (g1437) & (g2913) & (g2914) & (g2948) & (g2980)));
	assign g3013 = (((!g1437) & (!g2914) & (g2948) & (!g2980)) + ((!g1437) & (g2914) & (!g2948) & (!g2980)) + ((!g1437) & (g2914) & (!g2948) & (g2980)) + ((!g1437) & (g2914) & (g2948) & (g2980)) + ((g1437) & (!g2914) & (!g2948) & (!g2980)) + ((g1437) & (g2914) & (!g2948) & (g2980)) + ((g1437) & (g2914) & (g2948) & (!g2980)) + ((g1437) & (g2914) & (g2948) & (g2980)));
	assign g3014 = (((!g1423) & (!g1586) & (!g2916) & (g2917) & (g2947) & (!g2980)) + ((!g1423) & (!g1586) & (g2916) & (!g2917) & (!g2947) & (!g2980)) + ((!g1423) & (!g1586) & (g2916) & (!g2917) & (!g2947) & (g2980)) + ((!g1423) & (!g1586) & (g2916) & (!g2917) & (g2947) & (!g2980)) + ((!g1423) & (!g1586) & (g2916) & (!g2917) & (g2947) & (g2980)) + ((!g1423) & (!g1586) & (g2916) & (g2917) & (!g2947) & (!g2980)) + ((!g1423) & (!g1586) & (g2916) & (g2917) & (!g2947) & (g2980)) + ((!g1423) & (!g1586) & (g2916) & (g2917) & (g2947) & (g2980)) + ((!g1423) & (g1586) & (!g2916) & (!g2917) & (g2947) & (!g2980)) + ((!g1423) & (g1586) & (!g2916) & (g2917) & (!g2947) & (!g2980)) + ((!g1423) & (g1586) & (!g2916) & (g2917) & (g2947) & (!g2980)) + ((!g1423) & (g1586) & (g2916) & (!g2917) & (!g2947) & (!g2980)) + ((!g1423) & (g1586) & (g2916) & (!g2917) & (!g2947) & (g2980)) + ((!g1423) & (g1586) & (g2916) & (!g2917) & (g2947) & (g2980)) + ((!g1423) & (g1586) & (g2916) & (g2917) & (!g2947) & (g2980)) + ((!g1423) & (g1586) & (g2916) & (g2917) & (g2947) & (g2980)) + ((g1423) & (!g1586) & (!g2916) & (!g2917) & (!g2947) & (!g2980)) + ((g1423) & (!g1586) & (!g2916) & (!g2917) & (g2947) & (!g2980)) + ((g1423) & (!g1586) & (!g2916) & (g2917) & (!g2947) & (!g2980)) + ((g1423) & (!g1586) & (g2916) & (!g2917) & (!g2947) & (g2980)) + ((g1423) & (!g1586) & (g2916) & (!g2917) & (g2947) & (g2980)) + ((g1423) & (!g1586) & (g2916) & (g2917) & (!g2947) & (g2980)) + ((g1423) & (!g1586) & (g2916) & (g2917) & (g2947) & (!g2980)) + ((g1423) & (!g1586) & (g2916) & (g2917) & (g2947) & (g2980)) + ((g1423) & (g1586) & (!g2916) & (!g2917) & (!g2947) & (!g2980)) + ((g1423) & (g1586) & (g2916) & (!g2917) & (!g2947) & (g2980)) + ((g1423) & (g1586) & (g2916) & (!g2917) & (g2947) & (!g2980)) + ((g1423) & (g1586) & (g2916) & (!g2917) & (g2947) & (g2980)) + ((g1423) & (g1586) & (g2916) & (g2917) & (!g2947) & (!g2980)) + ((g1423) & (g1586) & (g2916) & (g2917) & (!g2947) & (g2980)) + ((g1423) & (g1586) & (g2916) & (g2917) & (g2947) & (!g2980)) + ((g1423) & (g1586) & (g2916) & (g2917) & (g2947) & (g2980)));
	assign g3015 = (((!g1586) & (!g2917) & (g2947) & (!g2980)) + ((!g1586) & (g2917) & (!g2947) & (!g2980)) + ((!g1586) & (g2917) & (!g2947) & (g2980)) + ((!g1586) & (g2917) & (g2947) & (g2980)) + ((g1586) & (!g2917) & (!g2947) & (!g2980)) + ((g1586) & (g2917) & (!g2947) & (g2980)) + ((g1586) & (g2917) & (g2947) & (!g2980)) + ((g1586) & (g2917) & (g2947) & (g2980)));
	assign g3016 = (((!g1568) & (!g1742) & (!g2919) & (g2920) & (g2946) & (!g2980)) + ((!g1568) & (!g1742) & (g2919) & (!g2920) & (!g2946) & (!g2980)) + ((!g1568) & (!g1742) & (g2919) & (!g2920) & (!g2946) & (g2980)) + ((!g1568) & (!g1742) & (g2919) & (!g2920) & (g2946) & (!g2980)) + ((!g1568) & (!g1742) & (g2919) & (!g2920) & (g2946) & (g2980)) + ((!g1568) & (!g1742) & (g2919) & (g2920) & (!g2946) & (!g2980)) + ((!g1568) & (!g1742) & (g2919) & (g2920) & (!g2946) & (g2980)) + ((!g1568) & (!g1742) & (g2919) & (g2920) & (g2946) & (g2980)) + ((!g1568) & (g1742) & (!g2919) & (!g2920) & (g2946) & (!g2980)) + ((!g1568) & (g1742) & (!g2919) & (g2920) & (!g2946) & (!g2980)) + ((!g1568) & (g1742) & (!g2919) & (g2920) & (g2946) & (!g2980)) + ((!g1568) & (g1742) & (g2919) & (!g2920) & (!g2946) & (!g2980)) + ((!g1568) & (g1742) & (g2919) & (!g2920) & (!g2946) & (g2980)) + ((!g1568) & (g1742) & (g2919) & (!g2920) & (g2946) & (g2980)) + ((!g1568) & (g1742) & (g2919) & (g2920) & (!g2946) & (g2980)) + ((!g1568) & (g1742) & (g2919) & (g2920) & (g2946) & (g2980)) + ((g1568) & (!g1742) & (!g2919) & (!g2920) & (!g2946) & (!g2980)) + ((g1568) & (!g1742) & (!g2919) & (!g2920) & (g2946) & (!g2980)) + ((g1568) & (!g1742) & (!g2919) & (g2920) & (!g2946) & (!g2980)) + ((g1568) & (!g1742) & (g2919) & (!g2920) & (!g2946) & (g2980)) + ((g1568) & (!g1742) & (g2919) & (!g2920) & (g2946) & (g2980)) + ((g1568) & (!g1742) & (g2919) & (g2920) & (!g2946) & (g2980)) + ((g1568) & (!g1742) & (g2919) & (g2920) & (g2946) & (!g2980)) + ((g1568) & (!g1742) & (g2919) & (g2920) & (g2946) & (g2980)) + ((g1568) & (g1742) & (!g2919) & (!g2920) & (!g2946) & (!g2980)) + ((g1568) & (g1742) & (g2919) & (!g2920) & (!g2946) & (g2980)) + ((g1568) & (g1742) & (g2919) & (!g2920) & (g2946) & (!g2980)) + ((g1568) & (g1742) & (g2919) & (!g2920) & (g2946) & (g2980)) + ((g1568) & (g1742) & (g2919) & (g2920) & (!g2946) & (!g2980)) + ((g1568) & (g1742) & (g2919) & (g2920) & (!g2946) & (g2980)) + ((g1568) & (g1742) & (g2919) & (g2920) & (g2946) & (!g2980)) + ((g1568) & (g1742) & (g2919) & (g2920) & (g2946) & (g2980)));
	assign g3017 = (((!g1742) & (!g2920) & (g2946) & (!g2980)) + ((!g1742) & (g2920) & (!g2946) & (!g2980)) + ((!g1742) & (g2920) & (!g2946) & (g2980)) + ((!g1742) & (g2920) & (g2946) & (g2980)) + ((g1742) & (!g2920) & (!g2946) & (!g2980)) + ((g1742) & (g2920) & (!g2946) & (g2980)) + ((g1742) & (g2920) & (g2946) & (!g2980)) + ((g1742) & (g2920) & (g2946) & (g2980)));
	assign g3018 = (((!g1720) & (!g1905) & (!g2922) & (g2923) & (g2945) & (!g2980)) + ((!g1720) & (!g1905) & (g2922) & (!g2923) & (!g2945) & (!g2980)) + ((!g1720) & (!g1905) & (g2922) & (!g2923) & (!g2945) & (g2980)) + ((!g1720) & (!g1905) & (g2922) & (!g2923) & (g2945) & (!g2980)) + ((!g1720) & (!g1905) & (g2922) & (!g2923) & (g2945) & (g2980)) + ((!g1720) & (!g1905) & (g2922) & (g2923) & (!g2945) & (!g2980)) + ((!g1720) & (!g1905) & (g2922) & (g2923) & (!g2945) & (g2980)) + ((!g1720) & (!g1905) & (g2922) & (g2923) & (g2945) & (g2980)) + ((!g1720) & (g1905) & (!g2922) & (!g2923) & (g2945) & (!g2980)) + ((!g1720) & (g1905) & (!g2922) & (g2923) & (!g2945) & (!g2980)) + ((!g1720) & (g1905) & (!g2922) & (g2923) & (g2945) & (!g2980)) + ((!g1720) & (g1905) & (g2922) & (!g2923) & (!g2945) & (!g2980)) + ((!g1720) & (g1905) & (g2922) & (!g2923) & (!g2945) & (g2980)) + ((!g1720) & (g1905) & (g2922) & (!g2923) & (g2945) & (g2980)) + ((!g1720) & (g1905) & (g2922) & (g2923) & (!g2945) & (g2980)) + ((!g1720) & (g1905) & (g2922) & (g2923) & (g2945) & (g2980)) + ((g1720) & (!g1905) & (!g2922) & (!g2923) & (!g2945) & (!g2980)) + ((g1720) & (!g1905) & (!g2922) & (!g2923) & (g2945) & (!g2980)) + ((g1720) & (!g1905) & (!g2922) & (g2923) & (!g2945) & (!g2980)) + ((g1720) & (!g1905) & (g2922) & (!g2923) & (!g2945) & (g2980)) + ((g1720) & (!g1905) & (g2922) & (!g2923) & (g2945) & (g2980)) + ((g1720) & (!g1905) & (g2922) & (g2923) & (!g2945) & (g2980)) + ((g1720) & (!g1905) & (g2922) & (g2923) & (g2945) & (!g2980)) + ((g1720) & (!g1905) & (g2922) & (g2923) & (g2945) & (g2980)) + ((g1720) & (g1905) & (!g2922) & (!g2923) & (!g2945) & (!g2980)) + ((g1720) & (g1905) & (g2922) & (!g2923) & (!g2945) & (g2980)) + ((g1720) & (g1905) & (g2922) & (!g2923) & (g2945) & (!g2980)) + ((g1720) & (g1905) & (g2922) & (!g2923) & (g2945) & (g2980)) + ((g1720) & (g1905) & (g2922) & (g2923) & (!g2945) & (!g2980)) + ((g1720) & (g1905) & (g2922) & (g2923) & (!g2945) & (g2980)) + ((g1720) & (g1905) & (g2922) & (g2923) & (g2945) & (!g2980)) + ((g1720) & (g1905) & (g2922) & (g2923) & (g2945) & (g2980)));
	assign g3019 = (((!g1905) & (!g2923) & (g2945) & (!g2980)) + ((!g1905) & (g2923) & (!g2945) & (!g2980)) + ((!g1905) & (g2923) & (!g2945) & (g2980)) + ((!g1905) & (g2923) & (g2945) & (g2980)) + ((g1905) & (!g2923) & (!g2945) & (!g2980)) + ((g1905) & (g2923) & (!g2945) & (g2980)) + ((g1905) & (g2923) & (g2945) & (!g2980)) + ((g1905) & (g2923) & (g2945) & (g2980)));
	assign g3020 = (((!g1879) & (!g2075) & (!g2925) & (g2926) & (g2944) & (!g2980)) + ((!g1879) & (!g2075) & (g2925) & (!g2926) & (!g2944) & (!g2980)) + ((!g1879) & (!g2075) & (g2925) & (!g2926) & (!g2944) & (g2980)) + ((!g1879) & (!g2075) & (g2925) & (!g2926) & (g2944) & (!g2980)) + ((!g1879) & (!g2075) & (g2925) & (!g2926) & (g2944) & (g2980)) + ((!g1879) & (!g2075) & (g2925) & (g2926) & (!g2944) & (!g2980)) + ((!g1879) & (!g2075) & (g2925) & (g2926) & (!g2944) & (g2980)) + ((!g1879) & (!g2075) & (g2925) & (g2926) & (g2944) & (g2980)) + ((!g1879) & (g2075) & (!g2925) & (!g2926) & (g2944) & (!g2980)) + ((!g1879) & (g2075) & (!g2925) & (g2926) & (!g2944) & (!g2980)) + ((!g1879) & (g2075) & (!g2925) & (g2926) & (g2944) & (!g2980)) + ((!g1879) & (g2075) & (g2925) & (!g2926) & (!g2944) & (!g2980)) + ((!g1879) & (g2075) & (g2925) & (!g2926) & (!g2944) & (g2980)) + ((!g1879) & (g2075) & (g2925) & (!g2926) & (g2944) & (g2980)) + ((!g1879) & (g2075) & (g2925) & (g2926) & (!g2944) & (g2980)) + ((!g1879) & (g2075) & (g2925) & (g2926) & (g2944) & (g2980)) + ((g1879) & (!g2075) & (!g2925) & (!g2926) & (!g2944) & (!g2980)) + ((g1879) & (!g2075) & (!g2925) & (!g2926) & (g2944) & (!g2980)) + ((g1879) & (!g2075) & (!g2925) & (g2926) & (!g2944) & (!g2980)) + ((g1879) & (!g2075) & (g2925) & (!g2926) & (!g2944) & (g2980)) + ((g1879) & (!g2075) & (g2925) & (!g2926) & (g2944) & (g2980)) + ((g1879) & (!g2075) & (g2925) & (g2926) & (!g2944) & (g2980)) + ((g1879) & (!g2075) & (g2925) & (g2926) & (g2944) & (!g2980)) + ((g1879) & (!g2075) & (g2925) & (g2926) & (g2944) & (g2980)) + ((g1879) & (g2075) & (!g2925) & (!g2926) & (!g2944) & (!g2980)) + ((g1879) & (g2075) & (g2925) & (!g2926) & (!g2944) & (g2980)) + ((g1879) & (g2075) & (g2925) & (!g2926) & (g2944) & (!g2980)) + ((g1879) & (g2075) & (g2925) & (!g2926) & (g2944) & (g2980)) + ((g1879) & (g2075) & (g2925) & (g2926) & (!g2944) & (!g2980)) + ((g1879) & (g2075) & (g2925) & (g2926) & (!g2944) & (g2980)) + ((g1879) & (g2075) & (g2925) & (g2926) & (g2944) & (!g2980)) + ((g1879) & (g2075) & (g2925) & (g2926) & (g2944) & (g2980)));
	assign g3021 = (((!g2075) & (!g2926) & (g2944) & (!g2980)) + ((!g2075) & (g2926) & (!g2944) & (!g2980)) + ((!g2075) & (g2926) & (!g2944) & (g2980)) + ((!g2075) & (g2926) & (g2944) & (g2980)) + ((g2075) & (!g2926) & (!g2944) & (!g2980)) + ((g2075) & (g2926) & (!g2944) & (g2980)) + ((g2075) & (g2926) & (g2944) & (!g2980)) + ((g2075) & (g2926) & (g2944) & (g2980)));
	assign g3022 = (((!g2045) & (!g2252) & (!g2928) & (g2929) & (g2943) & (!g2980)) + ((!g2045) & (!g2252) & (g2928) & (!g2929) & (!g2943) & (!g2980)) + ((!g2045) & (!g2252) & (g2928) & (!g2929) & (!g2943) & (g2980)) + ((!g2045) & (!g2252) & (g2928) & (!g2929) & (g2943) & (!g2980)) + ((!g2045) & (!g2252) & (g2928) & (!g2929) & (g2943) & (g2980)) + ((!g2045) & (!g2252) & (g2928) & (g2929) & (!g2943) & (!g2980)) + ((!g2045) & (!g2252) & (g2928) & (g2929) & (!g2943) & (g2980)) + ((!g2045) & (!g2252) & (g2928) & (g2929) & (g2943) & (g2980)) + ((!g2045) & (g2252) & (!g2928) & (!g2929) & (g2943) & (!g2980)) + ((!g2045) & (g2252) & (!g2928) & (g2929) & (!g2943) & (!g2980)) + ((!g2045) & (g2252) & (!g2928) & (g2929) & (g2943) & (!g2980)) + ((!g2045) & (g2252) & (g2928) & (!g2929) & (!g2943) & (!g2980)) + ((!g2045) & (g2252) & (g2928) & (!g2929) & (!g2943) & (g2980)) + ((!g2045) & (g2252) & (g2928) & (!g2929) & (g2943) & (g2980)) + ((!g2045) & (g2252) & (g2928) & (g2929) & (!g2943) & (g2980)) + ((!g2045) & (g2252) & (g2928) & (g2929) & (g2943) & (g2980)) + ((g2045) & (!g2252) & (!g2928) & (!g2929) & (!g2943) & (!g2980)) + ((g2045) & (!g2252) & (!g2928) & (!g2929) & (g2943) & (!g2980)) + ((g2045) & (!g2252) & (!g2928) & (g2929) & (!g2943) & (!g2980)) + ((g2045) & (!g2252) & (g2928) & (!g2929) & (!g2943) & (g2980)) + ((g2045) & (!g2252) & (g2928) & (!g2929) & (g2943) & (g2980)) + ((g2045) & (!g2252) & (g2928) & (g2929) & (!g2943) & (g2980)) + ((g2045) & (!g2252) & (g2928) & (g2929) & (g2943) & (!g2980)) + ((g2045) & (!g2252) & (g2928) & (g2929) & (g2943) & (g2980)) + ((g2045) & (g2252) & (!g2928) & (!g2929) & (!g2943) & (!g2980)) + ((g2045) & (g2252) & (g2928) & (!g2929) & (!g2943) & (g2980)) + ((g2045) & (g2252) & (g2928) & (!g2929) & (g2943) & (!g2980)) + ((g2045) & (g2252) & (g2928) & (!g2929) & (g2943) & (g2980)) + ((g2045) & (g2252) & (g2928) & (g2929) & (!g2943) & (!g2980)) + ((g2045) & (g2252) & (g2928) & (g2929) & (!g2943) & (g2980)) + ((g2045) & (g2252) & (g2928) & (g2929) & (g2943) & (!g2980)) + ((g2045) & (g2252) & (g2928) & (g2929) & (g2943) & (g2980)));
	assign g3023 = (((!g2252) & (!g2929) & (g2943) & (!g2980)) + ((!g2252) & (g2929) & (!g2943) & (!g2980)) + ((!g2252) & (g2929) & (!g2943) & (g2980)) + ((!g2252) & (g2929) & (g2943) & (g2980)) + ((g2252) & (!g2929) & (!g2943) & (!g2980)) + ((g2252) & (g2929) & (!g2943) & (g2980)) + ((g2252) & (g2929) & (g2943) & (!g2980)) + ((g2252) & (g2929) & (g2943) & (g2980)));
	assign g3024 = (((!g2218) & (!g2436) & (!g2931) & (g2932) & (g2942) & (!g2980)) + ((!g2218) & (!g2436) & (g2931) & (!g2932) & (!g2942) & (!g2980)) + ((!g2218) & (!g2436) & (g2931) & (!g2932) & (!g2942) & (g2980)) + ((!g2218) & (!g2436) & (g2931) & (!g2932) & (g2942) & (!g2980)) + ((!g2218) & (!g2436) & (g2931) & (!g2932) & (g2942) & (g2980)) + ((!g2218) & (!g2436) & (g2931) & (g2932) & (!g2942) & (!g2980)) + ((!g2218) & (!g2436) & (g2931) & (g2932) & (!g2942) & (g2980)) + ((!g2218) & (!g2436) & (g2931) & (g2932) & (g2942) & (g2980)) + ((!g2218) & (g2436) & (!g2931) & (!g2932) & (g2942) & (!g2980)) + ((!g2218) & (g2436) & (!g2931) & (g2932) & (!g2942) & (!g2980)) + ((!g2218) & (g2436) & (!g2931) & (g2932) & (g2942) & (!g2980)) + ((!g2218) & (g2436) & (g2931) & (!g2932) & (!g2942) & (!g2980)) + ((!g2218) & (g2436) & (g2931) & (!g2932) & (!g2942) & (g2980)) + ((!g2218) & (g2436) & (g2931) & (!g2932) & (g2942) & (g2980)) + ((!g2218) & (g2436) & (g2931) & (g2932) & (!g2942) & (g2980)) + ((!g2218) & (g2436) & (g2931) & (g2932) & (g2942) & (g2980)) + ((g2218) & (!g2436) & (!g2931) & (!g2932) & (!g2942) & (!g2980)) + ((g2218) & (!g2436) & (!g2931) & (!g2932) & (g2942) & (!g2980)) + ((g2218) & (!g2436) & (!g2931) & (g2932) & (!g2942) & (!g2980)) + ((g2218) & (!g2436) & (g2931) & (!g2932) & (!g2942) & (g2980)) + ((g2218) & (!g2436) & (g2931) & (!g2932) & (g2942) & (g2980)) + ((g2218) & (!g2436) & (g2931) & (g2932) & (!g2942) & (g2980)) + ((g2218) & (!g2436) & (g2931) & (g2932) & (g2942) & (!g2980)) + ((g2218) & (!g2436) & (g2931) & (g2932) & (g2942) & (g2980)) + ((g2218) & (g2436) & (!g2931) & (!g2932) & (!g2942) & (!g2980)) + ((g2218) & (g2436) & (g2931) & (!g2932) & (!g2942) & (g2980)) + ((g2218) & (g2436) & (g2931) & (!g2932) & (g2942) & (!g2980)) + ((g2218) & (g2436) & (g2931) & (!g2932) & (g2942) & (g2980)) + ((g2218) & (g2436) & (g2931) & (g2932) & (!g2942) & (!g2980)) + ((g2218) & (g2436) & (g2931) & (g2932) & (!g2942) & (g2980)) + ((g2218) & (g2436) & (g2931) & (g2932) & (g2942) & (!g2980)) + ((g2218) & (g2436) & (g2931) & (g2932) & (g2942) & (g2980)));
	assign g3025 = (((!g2436) & (!g2932) & (g2942) & (!g2980)) + ((!g2436) & (g2932) & (!g2942) & (!g2980)) + ((!g2436) & (g2932) & (!g2942) & (g2980)) + ((!g2436) & (g2932) & (g2942) & (g2980)) + ((g2436) & (!g2932) & (!g2942) & (!g2980)) + ((g2436) & (g2932) & (!g2942) & (g2980)) + ((g2436) & (g2932) & (g2942) & (!g2980)) + ((g2436) & (g2932) & (g2942) & (g2980)));
	assign g3026 = (((!g2398) & (!g2627) & (!g2934) & (g2935) & (g2941) & (!g2980)) + ((!g2398) & (!g2627) & (g2934) & (!g2935) & (!g2941) & (!g2980)) + ((!g2398) & (!g2627) & (g2934) & (!g2935) & (!g2941) & (g2980)) + ((!g2398) & (!g2627) & (g2934) & (!g2935) & (g2941) & (!g2980)) + ((!g2398) & (!g2627) & (g2934) & (!g2935) & (g2941) & (g2980)) + ((!g2398) & (!g2627) & (g2934) & (g2935) & (!g2941) & (!g2980)) + ((!g2398) & (!g2627) & (g2934) & (g2935) & (!g2941) & (g2980)) + ((!g2398) & (!g2627) & (g2934) & (g2935) & (g2941) & (g2980)) + ((!g2398) & (g2627) & (!g2934) & (!g2935) & (g2941) & (!g2980)) + ((!g2398) & (g2627) & (!g2934) & (g2935) & (!g2941) & (!g2980)) + ((!g2398) & (g2627) & (!g2934) & (g2935) & (g2941) & (!g2980)) + ((!g2398) & (g2627) & (g2934) & (!g2935) & (!g2941) & (!g2980)) + ((!g2398) & (g2627) & (g2934) & (!g2935) & (!g2941) & (g2980)) + ((!g2398) & (g2627) & (g2934) & (!g2935) & (g2941) & (g2980)) + ((!g2398) & (g2627) & (g2934) & (g2935) & (!g2941) & (g2980)) + ((!g2398) & (g2627) & (g2934) & (g2935) & (g2941) & (g2980)) + ((g2398) & (!g2627) & (!g2934) & (!g2935) & (!g2941) & (!g2980)) + ((g2398) & (!g2627) & (!g2934) & (!g2935) & (g2941) & (!g2980)) + ((g2398) & (!g2627) & (!g2934) & (g2935) & (!g2941) & (!g2980)) + ((g2398) & (!g2627) & (g2934) & (!g2935) & (!g2941) & (g2980)) + ((g2398) & (!g2627) & (g2934) & (!g2935) & (g2941) & (g2980)) + ((g2398) & (!g2627) & (g2934) & (g2935) & (!g2941) & (g2980)) + ((g2398) & (!g2627) & (g2934) & (g2935) & (g2941) & (!g2980)) + ((g2398) & (!g2627) & (g2934) & (g2935) & (g2941) & (g2980)) + ((g2398) & (g2627) & (!g2934) & (!g2935) & (!g2941) & (!g2980)) + ((g2398) & (g2627) & (g2934) & (!g2935) & (!g2941) & (g2980)) + ((g2398) & (g2627) & (g2934) & (!g2935) & (g2941) & (!g2980)) + ((g2398) & (g2627) & (g2934) & (!g2935) & (g2941) & (g2980)) + ((g2398) & (g2627) & (g2934) & (g2935) & (!g2941) & (!g2980)) + ((g2398) & (g2627) & (g2934) & (g2935) & (!g2941) & (g2980)) + ((g2398) & (g2627) & (g2934) & (g2935) & (g2941) & (!g2980)) + ((g2398) & (g2627) & (g2934) & (g2935) & (g2941) & (g2980)));
	assign g3027 = (((!g2627) & (!g2935) & (g2941) & (!g2980)) + ((!g2627) & (g2935) & (!g2941) & (!g2980)) + ((!g2627) & (g2935) & (!g2941) & (g2980)) + ((!g2627) & (g2935) & (g2941) & (g2980)) + ((g2627) & (!g2935) & (!g2941) & (!g2980)) + ((g2627) & (g2935) & (!g2941) & (g2980)) + ((g2627) & (g2935) & (g2941) & (!g2980)) + ((g2627) & (g2935) & (g2941) & (g2980)));
	assign g3028 = (((!g2585) & (!g2825) & (!g2937) & (g2938) & (g2940) & (!g2980)) + ((!g2585) & (!g2825) & (g2937) & (!g2938) & (!g2940) & (!g2980)) + ((!g2585) & (!g2825) & (g2937) & (!g2938) & (!g2940) & (g2980)) + ((!g2585) & (!g2825) & (g2937) & (!g2938) & (g2940) & (!g2980)) + ((!g2585) & (!g2825) & (g2937) & (!g2938) & (g2940) & (g2980)) + ((!g2585) & (!g2825) & (g2937) & (g2938) & (!g2940) & (!g2980)) + ((!g2585) & (!g2825) & (g2937) & (g2938) & (!g2940) & (g2980)) + ((!g2585) & (!g2825) & (g2937) & (g2938) & (g2940) & (g2980)) + ((!g2585) & (g2825) & (!g2937) & (!g2938) & (g2940) & (!g2980)) + ((!g2585) & (g2825) & (!g2937) & (g2938) & (!g2940) & (!g2980)) + ((!g2585) & (g2825) & (!g2937) & (g2938) & (g2940) & (!g2980)) + ((!g2585) & (g2825) & (g2937) & (!g2938) & (!g2940) & (!g2980)) + ((!g2585) & (g2825) & (g2937) & (!g2938) & (!g2940) & (g2980)) + ((!g2585) & (g2825) & (g2937) & (!g2938) & (g2940) & (g2980)) + ((!g2585) & (g2825) & (g2937) & (g2938) & (!g2940) & (g2980)) + ((!g2585) & (g2825) & (g2937) & (g2938) & (g2940) & (g2980)) + ((g2585) & (!g2825) & (!g2937) & (!g2938) & (!g2940) & (!g2980)) + ((g2585) & (!g2825) & (!g2937) & (!g2938) & (g2940) & (!g2980)) + ((g2585) & (!g2825) & (!g2937) & (g2938) & (!g2940) & (!g2980)) + ((g2585) & (!g2825) & (g2937) & (!g2938) & (!g2940) & (g2980)) + ((g2585) & (!g2825) & (g2937) & (!g2938) & (g2940) & (g2980)) + ((g2585) & (!g2825) & (g2937) & (g2938) & (!g2940) & (g2980)) + ((g2585) & (!g2825) & (g2937) & (g2938) & (g2940) & (!g2980)) + ((g2585) & (!g2825) & (g2937) & (g2938) & (g2940) & (g2980)) + ((g2585) & (g2825) & (!g2937) & (!g2938) & (!g2940) & (!g2980)) + ((g2585) & (g2825) & (g2937) & (!g2938) & (!g2940) & (g2980)) + ((g2585) & (g2825) & (g2937) & (!g2938) & (g2940) & (!g2980)) + ((g2585) & (g2825) & (g2937) & (!g2938) & (g2940) & (g2980)) + ((g2585) & (g2825) & (g2937) & (g2938) & (!g2940) & (!g2980)) + ((g2585) & (g2825) & (g2937) & (g2938) & (!g2940) & (g2980)) + ((g2585) & (g2825) & (g2937) & (g2938) & (g2940) & (!g2980)) + ((g2585) & (g2825) & (g2937) & (g2938) & (g2940) & (g2980)));
	assign g3029 = (((!g2825) & (!g2938) & (g2940) & (!g2980)) + ((!g2825) & (g2938) & (!g2940) & (!g2980)) + ((!g2825) & (g2938) & (!g2940) & (g2980)) + ((!g2825) & (g2938) & (g2940) & (g2980)) + ((g2825) & (!g2938) & (!g2940) & (!g2980)) + ((g2825) & (g2938) & (!g2940) & (g2980)) + ((g2825) & (g2938) & (g2940) & (!g2980)) + ((g2825) & (g2938) & (g2940) & (g2980)));
	assign g3030 = (((!g2853) & (g2865)));
	assign g3031 = (((!g2779) & (!ax14x) & (!ax15x) & (!g3030) & (!g2939) & (g2980)) + ((!g2779) & (!ax14x) & (!ax15x) & (!g3030) & (g2939) & (!g2980)) + ((!g2779) & (!ax14x) & (!ax15x) & (!g3030) & (g2939) & (g2980)) + ((!g2779) & (!ax14x) & (!ax15x) & (g3030) & (!g2939) & (!g2980)) + ((!g2779) & (!ax14x) & (ax15x) & (!g3030) & (!g2939) & (!g2980)) + ((!g2779) & (!ax14x) & (ax15x) & (g3030) & (!g2939) & (g2980)) + ((!g2779) & (!ax14x) & (ax15x) & (g3030) & (g2939) & (!g2980)) + ((!g2779) & (!ax14x) & (ax15x) & (g3030) & (g2939) & (g2980)) + ((!g2779) & (ax14x) & (!ax15x) & (g3030) & (!g2939) & (!g2980)) + ((!g2779) & (ax14x) & (!ax15x) & (g3030) & (g2939) & (!g2980)) + ((!g2779) & (ax14x) & (ax15x) & (!g3030) & (!g2939) & (!g2980)) + ((!g2779) & (ax14x) & (ax15x) & (!g3030) & (!g2939) & (g2980)) + ((!g2779) & (ax14x) & (ax15x) & (!g3030) & (g2939) & (!g2980)) + ((!g2779) & (ax14x) & (ax15x) & (!g3030) & (g2939) & (g2980)) + ((!g2779) & (ax14x) & (ax15x) & (g3030) & (!g2939) & (g2980)) + ((!g2779) & (ax14x) & (ax15x) & (g3030) & (g2939) & (g2980)) + ((g2779) & (!ax14x) & (!ax15x) & (!g3030) & (!g2939) & (!g2980)) + ((g2779) & (!ax14x) & (!ax15x) & (!g3030) & (!g2939) & (g2980)) + ((g2779) & (!ax14x) & (!ax15x) & (!g3030) & (g2939) & (g2980)) + ((g2779) & (!ax14x) & (!ax15x) & (g3030) & (g2939) & (!g2980)) + ((g2779) & (!ax14x) & (ax15x) & (!g3030) & (g2939) & (!g2980)) + ((g2779) & (!ax14x) & (ax15x) & (g3030) & (!g2939) & (!g2980)) + ((g2779) & (!ax14x) & (ax15x) & (g3030) & (!g2939) & (g2980)) + ((g2779) & (!ax14x) & (ax15x) & (g3030) & (g2939) & (g2980)) + ((g2779) & (ax14x) & (!ax15x) & (!g3030) & (!g2939) & (!g2980)) + ((g2779) & (ax14x) & (!ax15x) & (!g3030) & (g2939) & (!g2980)) + ((g2779) & (ax14x) & (ax15x) & (!g3030) & (!g2939) & (g2980)) + ((g2779) & (ax14x) & (ax15x) & (!g3030) & (g2939) & (g2980)) + ((g2779) & (ax14x) & (ax15x) & (g3030) & (!g2939) & (!g2980)) + ((g2779) & (ax14x) & (ax15x) & (g3030) & (!g2939) & (g2980)) + ((g2779) & (ax14x) & (ax15x) & (g3030) & (g2939) & (!g2980)) + ((g2779) & (ax14x) & (ax15x) & (g3030) & (g2939) & (g2980)));
	assign g3032 = (((!ax14x) & (!g3030) & (!g2939) & (g2980)) + ((!ax14x) & (!g3030) & (g2939) & (!g2980)) + ((!ax14x) & (!g3030) & (g2939) & (g2980)) + ((!ax14x) & (g3030) & (g2939) & (!g2980)) + ((ax14x) & (!g3030) & (!g2939) & (!g2980)) + ((ax14x) & (g3030) & (!g2939) & (!g2980)) + ((ax14x) & (g3030) & (!g2939) & (g2980)) + ((ax14x) & (g3030) & (g2939) & (g2980)));
	assign g3033 = (((!ax10x) & (!ax11x)));
	assign g3034 = (((!g3030) & (!ax12x) & (!ax13x) & (!g2980) & (!g3033)) + ((!g3030) & (!ax12x) & (ax13x) & (g2980) & (!g3033)) + ((!g3030) & (ax12x) & (ax13x) & (g2980) & (!g3033)) + ((!g3030) & (ax12x) & (ax13x) & (g2980) & (g3033)) + ((g3030) & (!ax12x) & (!ax13x) & (!g2980) & (!g3033)) + ((g3030) & (!ax12x) & (!ax13x) & (!g2980) & (g3033)) + ((g3030) & (!ax12x) & (!ax13x) & (g2980) & (!g3033)) + ((g3030) & (!ax12x) & (ax13x) & (!g2980) & (!g3033)) + ((g3030) & (!ax12x) & (ax13x) & (g2980) & (!g3033)) + ((g3030) & (!ax12x) & (ax13x) & (g2980) & (g3033)) + ((g3030) & (ax12x) & (!ax13x) & (g2980) & (!g3033)) + ((g3030) & (ax12x) & (!ax13x) & (g2980) & (g3033)) + ((g3030) & (ax12x) & (ax13x) & (!g2980) & (!g3033)) + ((g3030) & (ax12x) & (ax13x) & (!g2980) & (g3033)) + ((g3030) & (ax12x) & (ax13x) & (g2980) & (!g3033)) + ((g3030) & (ax12x) & (ax13x) & (g2980) & (g3033)));
	assign g3035 = (((!g2825) & (!g2779) & (g3031) & (g3032) & (g3034)) + ((!g2825) & (g2779) & (g3031) & (!g3032) & (g3034)) + ((!g2825) & (g2779) & (g3031) & (g3032) & (!g3034)) + ((!g2825) & (g2779) & (g3031) & (g3032) & (g3034)) + ((g2825) & (!g2779) & (!g3031) & (g3032) & (g3034)) + ((g2825) & (!g2779) & (g3031) & (!g3032) & (!g3034)) + ((g2825) & (!g2779) & (g3031) & (!g3032) & (g3034)) + ((g2825) & (!g2779) & (g3031) & (g3032) & (!g3034)) + ((g2825) & (!g2779) & (g3031) & (g3032) & (g3034)) + ((g2825) & (g2779) & (!g3031) & (!g3032) & (g3034)) + ((g2825) & (g2779) & (!g3031) & (g3032) & (!g3034)) + ((g2825) & (g2779) & (!g3031) & (g3032) & (g3034)) + ((g2825) & (g2779) & (g3031) & (!g3032) & (!g3034)) + ((g2825) & (g2779) & (g3031) & (!g3032) & (g3034)) + ((g2825) & (g2779) & (g3031) & (g3032) & (!g3034)) + ((g2825) & (g2779) & (g3031) & (g3032) & (g3034)));
	assign g3036 = (((!g2627) & (!g2585) & (g3028) & (g3029) & (g3035)) + ((!g2627) & (g2585) & (g3028) & (!g3029) & (g3035)) + ((!g2627) & (g2585) & (g3028) & (g3029) & (!g3035)) + ((!g2627) & (g2585) & (g3028) & (g3029) & (g3035)) + ((g2627) & (!g2585) & (!g3028) & (g3029) & (g3035)) + ((g2627) & (!g2585) & (g3028) & (!g3029) & (!g3035)) + ((g2627) & (!g2585) & (g3028) & (!g3029) & (g3035)) + ((g2627) & (!g2585) & (g3028) & (g3029) & (!g3035)) + ((g2627) & (!g2585) & (g3028) & (g3029) & (g3035)) + ((g2627) & (g2585) & (!g3028) & (!g3029) & (g3035)) + ((g2627) & (g2585) & (!g3028) & (g3029) & (!g3035)) + ((g2627) & (g2585) & (!g3028) & (g3029) & (g3035)) + ((g2627) & (g2585) & (g3028) & (!g3029) & (!g3035)) + ((g2627) & (g2585) & (g3028) & (!g3029) & (g3035)) + ((g2627) & (g2585) & (g3028) & (g3029) & (!g3035)) + ((g2627) & (g2585) & (g3028) & (g3029) & (g3035)));
	assign g3037 = (((!g2436) & (!g2398) & (g3026) & (g3027) & (g3036)) + ((!g2436) & (g2398) & (g3026) & (!g3027) & (g3036)) + ((!g2436) & (g2398) & (g3026) & (g3027) & (!g3036)) + ((!g2436) & (g2398) & (g3026) & (g3027) & (g3036)) + ((g2436) & (!g2398) & (!g3026) & (g3027) & (g3036)) + ((g2436) & (!g2398) & (g3026) & (!g3027) & (!g3036)) + ((g2436) & (!g2398) & (g3026) & (!g3027) & (g3036)) + ((g2436) & (!g2398) & (g3026) & (g3027) & (!g3036)) + ((g2436) & (!g2398) & (g3026) & (g3027) & (g3036)) + ((g2436) & (g2398) & (!g3026) & (!g3027) & (g3036)) + ((g2436) & (g2398) & (!g3026) & (g3027) & (!g3036)) + ((g2436) & (g2398) & (!g3026) & (g3027) & (g3036)) + ((g2436) & (g2398) & (g3026) & (!g3027) & (!g3036)) + ((g2436) & (g2398) & (g3026) & (!g3027) & (g3036)) + ((g2436) & (g2398) & (g3026) & (g3027) & (!g3036)) + ((g2436) & (g2398) & (g3026) & (g3027) & (g3036)));
	assign g3038 = (((!g2252) & (!g2218) & (g3024) & (g3025) & (g3037)) + ((!g2252) & (g2218) & (g3024) & (!g3025) & (g3037)) + ((!g2252) & (g2218) & (g3024) & (g3025) & (!g3037)) + ((!g2252) & (g2218) & (g3024) & (g3025) & (g3037)) + ((g2252) & (!g2218) & (!g3024) & (g3025) & (g3037)) + ((g2252) & (!g2218) & (g3024) & (!g3025) & (!g3037)) + ((g2252) & (!g2218) & (g3024) & (!g3025) & (g3037)) + ((g2252) & (!g2218) & (g3024) & (g3025) & (!g3037)) + ((g2252) & (!g2218) & (g3024) & (g3025) & (g3037)) + ((g2252) & (g2218) & (!g3024) & (!g3025) & (g3037)) + ((g2252) & (g2218) & (!g3024) & (g3025) & (!g3037)) + ((g2252) & (g2218) & (!g3024) & (g3025) & (g3037)) + ((g2252) & (g2218) & (g3024) & (!g3025) & (!g3037)) + ((g2252) & (g2218) & (g3024) & (!g3025) & (g3037)) + ((g2252) & (g2218) & (g3024) & (g3025) & (!g3037)) + ((g2252) & (g2218) & (g3024) & (g3025) & (g3037)));
	assign g3039 = (((!g2075) & (!g2045) & (g3022) & (g3023) & (g3038)) + ((!g2075) & (g2045) & (g3022) & (!g3023) & (g3038)) + ((!g2075) & (g2045) & (g3022) & (g3023) & (!g3038)) + ((!g2075) & (g2045) & (g3022) & (g3023) & (g3038)) + ((g2075) & (!g2045) & (!g3022) & (g3023) & (g3038)) + ((g2075) & (!g2045) & (g3022) & (!g3023) & (!g3038)) + ((g2075) & (!g2045) & (g3022) & (!g3023) & (g3038)) + ((g2075) & (!g2045) & (g3022) & (g3023) & (!g3038)) + ((g2075) & (!g2045) & (g3022) & (g3023) & (g3038)) + ((g2075) & (g2045) & (!g3022) & (!g3023) & (g3038)) + ((g2075) & (g2045) & (!g3022) & (g3023) & (!g3038)) + ((g2075) & (g2045) & (!g3022) & (g3023) & (g3038)) + ((g2075) & (g2045) & (g3022) & (!g3023) & (!g3038)) + ((g2075) & (g2045) & (g3022) & (!g3023) & (g3038)) + ((g2075) & (g2045) & (g3022) & (g3023) & (!g3038)) + ((g2075) & (g2045) & (g3022) & (g3023) & (g3038)));
	assign g3040 = (((!g1905) & (!g1879) & (g3020) & (g3021) & (g3039)) + ((!g1905) & (g1879) & (g3020) & (!g3021) & (g3039)) + ((!g1905) & (g1879) & (g3020) & (g3021) & (!g3039)) + ((!g1905) & (g1879) & (g3020) & (g3021) & (g3039)) + ((g1905) & (!g1879) & (!g3020) & (g3021) & (g3039)) + ((g1905) & (!g1879) & (g3020) & (!g3021) & (!g3039)) + ((g1905) & (!g1879) & (g3020) & (!g3021) & (g3039)) + ((g1905) & (!g1879) & (g3020) & (g3021) & (!g3039)) + ((g1905) & (!g1879) & (g3020) & (g3021) & (g3039)) + ((g1905) & (g1879) & (!g3020) & (!g3021) & (g3039)) + ((g1905) & (g1879) & (!g3020) & (g3021) & (!g3039)) + ((g1905) & (g1879) & (!g3020) & (g3021) & (g3039)) + ((g1905) & (g1879) & (g3020) & (!g3021) & (!g3039)) + ((g1905) & (g1879) & (g3020) & (!g3021) & (g3039)) + ((g1905) & (g1879) & (g3020) & (g3021) & (!g3039)) + ((g1905) & (g1879) & (g3020) & (g3021) & (g3039)));
	assign g3041 = (((!g1742) & (!g1720) & (g3018) & (g3019) & (g3040)) + ((!g1742) & (g1720) & (g3018) & (!g3019) & (g3040)) + ((!g1742) & (g1720) & (g3018) & (g3019) & (!g3040)) + ((!g1742) & (g1720) & (g3018) & (g3019) & (g3040)) + ((g1742) & (!g1720) & (!g3018) & (g3019) & (g3040)) + ((g1742) & (!g1720) & (g3018) & (!g3019) & (!g3040)) + ((g1742) & (!g1720) & (g3018) & (!g3019) & (g3040)) + ((g1742) & (!g1720) & (g3018) & (g3019) & (!g3040)) + ((g1742) & (!g1720) & (g3018) & (g3019) & (g3040)) + ((g1742) & (g1720) & (!g3018) & (!g3019) & (g3040)) + ((g1742) & (g1720) & (!g3018) & (g3019) & (!g3040)) + ((g1742) & (g1720) & (!g3018) & (g3019) & (g3040)) + ((g1742) & (g1720) & (g3018) & (!g3019) & (!g3040)) + ((g1742) & (g1720) & (g3018) & (!g3019) & (g3040)) + ((g1742) & (g1720) & (g3018) & (g3019) & (!g3040)) + ((g1742) & (g1720) & (g3018) & (g3019) & (g3040)));
	assign g3042 = (((!g1586) & (!g1568) & (g3016) & (g3017) & (g3041)) + ((!g1586) & (g1568) & (g3016) & (!g3017) & (g3041)) + ((!g1586) & (g1568) & (g3016) & (g3017) & (!g3041)) + ((!g1586) & (g1568) & (g3016) & (g3017) & (g3041)) + ((g1586) & (!g1568) & (!g3016) & (g3017) & (g3041)) + ((g1586) & (!g1568) & (g3016) & (!g3017) & (!g3041)) + ((g1586) & (!g1568) & (g3016) & (!g3017) & (g3041)) + ((g1586) & (!g1568) & (g3016) & (g3017) & (!g3041)) + ((g1586) & (!g1568) & (g3016) & (g3017) & (g3041)) + ((g1586) & (g1568) & (!g3016) & (!g3017) & (g3041)) + ((g1586) & (g1568) & (!g3016) & (g3017) & (!g3041)) + ((g1586) & (g1568) & (!g3016) & (g3017) & (g3041)) + ((g1586) & (g1568) & (g3016) & (!g3017) & (!g3041)) + ((g1586) & (g1568) & (g3016) & (!g3017) & (g3041)) + ((g1586) & (g1568) & (g3016) & (g3017) & (!g3041)) + ((g1586) & (g1568) & (g3016) & (g3017) & (g3041)));
	assign g3043 = (((!g1437) & (!g1423) & (g3014) & (g3015) & (g3042)) + ((!g1437) & (g1423) & (g3014) & (!g3015) & (g3042)) + ((!g1437) & (g1423) & (g3014) & (g3015) & (!g3042)) + ((!g1437) & (g1423) & (g3014) & (g3015) & (g3042)) + ((g1437) & (!g1423) & (!g3014) & (g3015) & (g3042)) + ((g1437) & (!g1423) & (g3014) & (!g3015) & (!g3042)) + ((g1437) & (!g1423) & (g3014) & (!g3015) & (g3042)) + ((g1437) & (!g1423) & (g3014) & (g3015) & (!g3042)) + ((g1437) & (!g1423) & (g3014) & (g3015) & (g3042)) + ((g1437) & (g1423) & (!g3014) & (!g3015) & (g3042)) + ((g1437) & (g1423) & (!g3014) & (g3015) & (!g3042)) + ((g1437) & (g1423) & (!g3014) & (g3015) & (g3042)) + ((g1437) & (g1423) & (g3014) & (!g3015) & (!g3042)) + ((g1437) & (g1423) & (g3014) & (!g3015) & (g3042)) + ((g1437) & (g1423) & (g3014) & (g3015) & (!g3042)) + ((g1437) & (g1423) & (g3014) & (g3015) & (g3042)));
	assign g3044 = (((!g1295) & (!g1285) & (g3012) & (g3013) & (g3043)) + ((!g1295) & (g1285) & (g3012) & (!g3013) & (g3043)) + ((!g1295) & (g1285) & (g3012) & (g3013) & (!g3043)) + ((!g1295) & (g1285) & (g3012) & (g3013) & (g3043)) + ((g1295) & (!g1285) & (!g3012) & (g3013) & (g3043)) + ((g1295) & (!g1285) & (g3012) & (!g3013) & (!g3043)) + ((g1295) & (!g1285) & (g3012) & (!g3013) & (g3043)) + ((g1295) & (!g1285) & (g3012) & (g3013) & (!g3043)) + ((g1295) & (!g1285) & (g3012) & (g3013) & (g3043)) + ((g1295) & (g1285) & (!g3012) & (!g3013) & (g3043)) + ((g1295) & (g1285) & (!g3012) & (g3013) & (!g3043)) + ((g1295) & (g1285) & (!g3012) & (g3013) & (g3043)) + ((g1295) & (g1285) & (g3012) & (!g3013) & (!g3043)) + ((g1295) & (g1285) & (g3012) & (!g3013) & (g3043)) + ((g1295) & (g1285) & (g3012) & (g3013) & (!g3043)) + ((g1295) & (g1285) & (g3012) & (g3013) & (g3043)));
	assign g3045 = (((!g1160) & (!g1154) & (g3010) & (g3011) & (g3044)) + ((!g1160) & (g1154) & (g3010) & (!g3011) & (g3044)) + ((!g1160) & (g1154) & (g3010) & (g3011) & (!g3044)) + ((!g1160) & (g1154) & (g3010) & (g3011) & (g3044)) + ((g1160) & (!g1154) & (!g3010) & (g3011) & (g3044)) + ((g1160) & (!g1154) & (g3010) & (!g3011) & (!g3044)) + ((g1160) & (!g1154) & (g3010) & (!g3011) & (g3044)) + ((g1160) & (!g1154) & (g3010) & (g3011) & (!g3044)) + ((g1160) & (!g1154) & (g3010) & (g3011) & (g3044)) + ((g1160) & (g1154) & (!g3010) & (!g3011) & (g3044)) + ((g1160) & (g1154) & (!g3010) & (g3011) & (!g3044)) + ((g1160) & (g1154) & (!g3010) & (g3011) & (g3044)) + ((g1160) & (g1154) & (g3010) & (!g3011) & (!g3044)) + ((g1160) & (g1154) & (g3010) & (!g3011) & (g3044)) + ((g1160) & (g1154) & (g3010) & (g3011) & (!g3044)) + ((g1160) & (g1154) & (g3010) & (g3011) & (g3044)));
	assign g3046 = (((!g1032) & (!g1030) & (g3008) & (g3009) & (g3045)) + ((!g1032) & (g1030) & (g3008) & (!g3009) & (g3045)) + ((!g1032) & (g1030) & (g3008) & (g3009) & (!g3045)) + ((!g1032) & (g1030) & (g3008) & (g3009) & (g3045)) + ((g1032) & (!g1030) & (!g3008) & (g3009) & (g3045)) + ((g1032) & (!g1030) & (g3008) & (!g3009) & (!g3045)) + ((g1032) & (!g1030) & (g3008) & (!g3009) & (g3045)) + ((g1032) & (!g1030) & (g3008) & (g3009) & (!g3045)) + ((g1032) & (!g1030) & (g3008) & (g3009) & (g3045)) + ((g1032) & (g1030) & (!g3008) & (!g3009) & (g3045)) + ((g1032) & (g1030) & (!g3008) & (g3009) & (!g3045)) + ((g1032) & (g1030) & (!g3008) & (g3009) & (g3045)) + ((g1032) & (g1030) & (g3008) & (!g3009) & (!g3045)) + ((g1032) & (g1030) & (g3008) & (!g3009) & (g3045)) + ((g1032) & (g1030) & (g3008) & (g3009) & (!g3045)) + ((g1032) & (g1030) & (g3008) & (g3009) & (g3045)));
	assign g3047 = (((!g851) & (!g914) & (g3006) & (g3007) & (g3046)) + ((!g851) & (g914) & (g3006) & (!g3007) & (g3046)) + ((!g851) & (g914) & (g3006) & (g3007) & (!g3046)) + ((!g851) & (g914) & (g3006) & (g3007) & (g3046)) + ((g851) & (!g914) & (!g3006) & (g3007) & (g3046)) + ((g851) & (!g914) & (g3006) & (!g3007) & (!g3046)) + ((g851) & (!g914) & (g3006) & (!g3007) & (g3046)) + ((g851) & (!g914) & (g3006) & (g3007) & (!g3046)) + ((g851) & (!g914) & (g3006) & (g3007) & (g3046)) + ((g851) & (g914) & (!g3006) & (!g3007) & (g3046)) + ((g851) & (g914) & (!g3006) & (g3007) & (!g3046)) + ((g851) & (g914) & (!g3006) & (g3007) & (g3046)) + ((g851) & (g914) & (g3006) & (!g3007) & (!g3046)) + ((g851) & (g914) & (g3006) & (!g3007) & (g3046)) + ((g851) & (g914) & (g3006) & (g3007) & (!g3046)) + ((g851) & (g914) & (g3006) & (g3007) & (g3046)));
	assign g3048 = (((!g744) & (!g803) & (g3004) & (g3005) & (g3047)) + ((!g744) & (g803) & (g3004) & (!g3005) & (g3047)) + ((!g744) & (g803) & (g3004) & (g3005) & (!g3047)) + ((!g744) & (g803) & (g3004) & (g3005) & (g3047)) + ((g744) & (!g803) & (!g3004) & (g3005) & (g3047)) + ((g744) & (!g803) & (g3004) & (!g3005) & (!g3047)) + ((g744) & (!g803) & (g3004) & (!g3005) & (g3047)) + ((g744) & (!g803) & (g3004) & (g3005) & (!g3047)) + ((g744) & (!g803) & (g3004) & (g3005) & (g3047)) + ((g744) & (g803) & (!g3004) & (!g3005) & (g3047)) + ((g744) & (g803) & (!g3004) & (g3005) & (!g3047)) + ((g744) & (g803) & (!g3004) & (g3005) & (g3047)) + ((g744) & (g803) & (g3004) & (!g3005) & (!g3047)) + ((g744) & (g803) & (g3004) & (!g3005) & (g3047)) + ((g744) & (g803) & (g3004) & (g3005) & (!g3047)) + ((g744) & (g803) & (g3004) & (g3005) & (g3047)));
	assign g3049 = (((!g645) & (!g700) & (g3002) & (g3003) & (g3048)) + ((!g645) & (g700) & (g3002) & (!g3003) & (g3048)) + ((!g645) & (g700) & (g3002) & (g3003) & (!g3048)) + ((!g645) & (g700) & (g3002) & (g3003) & (g3048)) + ((g645) & (!g700) & (!g3002) & (g3003) & (g3048)) + ((g645) & (!g700) & (g3002) & (!g3003) & (!g3048)) + ((g645) & (!g700) & (g3002) & (!g3003) & (g3048)) + ((g645) & (!g700) & (g3002) & (g3003) & (!g3048)) + ((g645) & (!g700) & (g3002) & (g3003) & (g3048)) + ((g645) & (g700) & (!g3002) & (!g3003) & (g3048)) + ((g645) & (g700) & (!g3002) & (g3003) & (!g3048)) + ((g645) & (g700) & (!g3002) & (g3003) & (g3048)) + ((g645) & (g700) & (g3002) & (!g3003) & (!g3048)) + ((g645) & (g700) & (g3002) & (!g3003) & (g3048)) + ((g645) & (g700) & (g3002) & (g3003) & (!g3048)) + ((g645) & (g700) & (g3002) & (g3003) & (g3048)));
	assign g3050 = (((!g553) & (!g604) & (g3000) & (g3001) & (g3049)) + ((!g553) & (g604) & (g3000) & (!g3001) & (g3049)) + ((!g553) & (g604) & (g3000) & (g3001) & (!g3049)) + ((!g553) & (g604) & (g3000) & (g3001) & (g3049)) + ((g553) & (!g604) & (!g3000) & (g3001) & (g3049)) + ((g553) & (!g604) & (g3000) & (!g3001) & (!g3049)) + ((g553) & (!g604) & (g3000) & (!g3001) & (g3049)) + ((g553) & (!g604) & (g3000) & (g3001) & (!g3049)) + ((g553) & (!g604) & (g3000) & (g3001) & (g3049)) + ((g553) & (g604) & (!g3000) & (!g3001) & (g3049)) + ((g553) & (g604) & (!g3000) & (g3001) & (!g3049)) + ((g553) & (g604) & (!g3000) & (g3001) & (g3049)) + ((g553) & (g604) & (g3000) & (!g3001) & (!g3049)) + ((g553) & (g604) & (g3000) & (!g3001) & (g3049)) + ((g553) & (g604) & (g3000) & (g3001) & (!g3049)) + ((g553) & (g604) & (g3000) & (g3001) & (g3049)));
	assign g3051 = (((!g468) & (!g515) & (g2998) & (g2999) & (g3050)) + ((!g468) & (g515) & (g2998) & (!g2999) & (g3050)) + ((!g468) & (g515) & (g2998) & (g2999) & (!g3050)) + ((!g468) & (g515) & (g2998) & (g2999) & (g3050)) + ((g468) & (!g515) & (!g2998) & (g2999) & (g3050)) + ((g468) & (!g515) & (g2998) & (!g2999) & (!g3050)) + ((g468) & (!g515) & (g2998) & (!g2999) & (g3050)) + ((g468) & (!g515) & (g2998) & (g2999) & (!g3050)) + ((g468) & (!g515) & (g2998) & (g2999) & (g3050)) + ((g468) & (g515) & (!g2998) & (!g2999) & (g3050)) + ((g468) & (g515) & (!g2998) & (g2999) & (!g3050)) + ((g468) & (g515) & (!g2998) & (g2999) & (g3050)) + ((g468) & (g515) & (g2998) & (!g2999) & (!g3050)) + ((g468) & (g515) & (g2998) & (!g2999) & (g3050)) + ((g468) & (g515) & (g2998) & (g2999) & (!g3050)) + ((g468) & (g515) & (g2998) & (g2999) & (g3050)));
	assign g3052 = (((!g390) & (!g433) & (g2996) & (g2997) & (g3051)) + ((!g390) & (g433) & (g2996) & (!g2997) & (g3051)) + ((!g390) & (g433) & (g2996) & (g2997) & (!g3051)) + ((!g390) & (g433) & (g2996) & (g2997) & (g3051)) + ((g390) & (!g433) & (!g2996) & (g2997) & (g3051)) + ((g390) & (!g433) & (g2996) & (!g2997) & (!g3051)) + ((g390) & (!g433) & (g2996) & (!g2997) & (g3051)) + ((g390) & (!g433) & (g2996) & (g2997) & (!g3051)) + ((g390) & (!g433) & (g2996) & (g2997) & (g3051)) + ((g390) & (g433) & (!g2996) & (!g2997) & (g3051)) + ((g390) & (g433) & (!g2996) & (g2997) & (!g3051)) + ((g390) & (g433) & (!g2996) & (g2997) & (g3051)) + ((g390) & (g433) & (g2996) & (!g2997) & (!g3051)) + ((g390) & (g433) & (g2996) & (!g2997) & (g3051)) + ((g390) & (g433) & (g2996) & (g2997) & (!g3051)) + ((g390) & (g433) & (g2996) & (g2997) & (g3051)));
	assign g3053 = (((!g319) & (!g358) & (g2994) & (g2995) & (g3052)) + ((!g319) & (g358) & (g2994) & (!g2995) & (g3052)) + ((!g319) & (g358) & (g2994) & (g2995) & (!g3052)) + ((!g319) & (g358) & (g2994) & (g2995) & (g3052)) + ((g319) & (!g358) & (!g2994) & (g2995) & (g3052)) + ((g319) & (!g358) & (g2994) & (!g2995) & (!g3052)) + ((g319) & (!g358) & (g2994) & (!g2995) & (g3052)) + ((g319) & (!g358) & (g2994) & (g2995) & (!g3052)) + ((g319) & (!g358) & (g2994) & (g2995) & (g3052)) + ((g319) & (g358) & (!g2994) & (!g2995) & (g3052)) + ((g319) & (g358) & (!g2994) & (g2995) & (!g3052)) + ((g319) & (g358) & (!g2994) & (g2995) & (g3052)) + ((g319) & (g358) & (g2994) & (!g2995) & (!g3052)) + ((g319) & (g358) & (g2994) & (!g2995) & (g3052)) + ((g319) & (g358) & (g2994) & (g2995) & (!g3052)) + ((g319) & (g358) & (g2994) & (g2995) & (g3052)));
	assign g3054 = (((!g255) & (!g290) & (g2992) & (g2993) & (g3053)) + ((!g255) & (g290) & (g2992) & (!g2993) & (g3053)) + ((!g255) & (g290) & (g2992) & (g2993) & (!g3053)) + ((!g255) & (g290) & (g2992) & (g2993) & (g3053)) + ((g255) & (!g290) & (!g2992) & (g2993) & (g3053)) + ((g255) & (!g290) & (g2992) & (!g2993) & (!g3053)) + ((g255) & (!g290) & (g2992) & (!g2993) & (g3053)) + ((g255) & (!g290) & (g2992) & (g2993) & (!g3053)) + ((g255) & (!g290) & (g2992) & (g2993) & (g3053)) + ((g255) & (g290) & (!g2992) & (!g2993) & (g3053)) + ((g255) & (g290) & (!g2992) & (g2993) & (!g3053)) + ((g255) & (g290) & (!g2992) & (g2993) & (g3053)) + ((g255) & (g290) & (g2992) & (!g2993) & (!g3053)) + ((g255) & (g290) & (g2992) & (!g2993) & (g3053)) + ((g255) & (g290) & (g2992) & (g2993) & (!g3053)) + ((g255) & (g290) & (g2992) & (g2993) & (g3053)));
	assign g3055 = (((!g198) & (!g229) & (g2990) & (g2991) & (g3054)) + ((!g198) & (g229) & (g2990) & (!g2991) & (g3054)) + ((!g198) & (g229) & (g2990) & (g2991) & (!g3054)) + ((!g198) & (g229) & (g2990) & (g2991) & (g3054)) + ((g198) & (!g229) & (!g2990) & (g2991) & (g3054)) + ((g198) & (!g229) & (g2990) & (!g2991) & (!g3054)) + ((g198) & (!g229) & (g2990) & (!g2991) & (g3054)) + ((g198) & (!g229) & (g2990) & (g2991) & (!g3054)) + ((g198) & (!g229) & (g2990) & (g2991) & (g3054)) + ((g198) & (g229) & (!g2990) & (!g2991) & (g3054)) + ((g198) & (g229) & (!g2990) & (g2991) & (!g3054)) + ((g198) & (g229) & (!g2990) & (g2991) & (g3054)) + ((g198) & (g229) & (g2990) & (!g2991) & (!g3054)) + ((g198) & (g229) & (g2990) & (!g2991) & (g3054)) + ((g198) & (g229) & (g2990) & (g2991) & (!g3054)) + ((g198) & (g229) & (g2990) & (g2991) & (g3054)));
	assign g3056 = (((!g147) & (!g174) & (g2988) & (g2989) & (g3055)) + ((!g147) & (g174) & (g2988) & (!g2989) & (g3055)) + ((!g147) & (g174) & (g2988) & (g2989) & (!g3055)) + ((!g147) & (g174) & (g2988) & (g2989) & (g3055)) + ((g147) & (!g174) & (!g2988) & (g2989) & (g3055)) + ((g147) & (!g174) & (g2988) & (!g2989) & (!g3055)) + ((g147) & (!g174) & (g2988) & (!g2989) & (g3055)) + ((g147) & (!g174) & (g2988) & (g2989) & (!g3055)) + ((g147) & (!g174) & (g2988) & (g2989) & (g3055)) + ((g147) & (g174) & (!g2988) & (!g2989) & (g3055)) + ((g147) & (g174) & (!g2988) & (g2989) & (!g3055)) + ((g147) & (g174) & (!g2988) & (g2989) & (g3055)) + ((g147) & (g174) & (g2988) & (!g2989) & (!g3055)) + ((g147) & (g174) & (g2988) & (!g2989) & (g3055)) + ((g147) & (g174) & (g2988) & (g2989) & (!g3055)) + ((g147) & (g174) & (g2988) & (g2989) & (g3055)));
	assign g3057 = (((!g104) & (!g127) & (g2986) & (g2987) & (g3056)) + ((!g104) & (g127) & (g2986) & (!g2987) & (g3056)) + ((!g104) & (g127) & (g2986) & (g2987) & (!g3056)) + ((!g104) & (g127) & (g2986) & (g2987) & (g3056)) + ((g104) & (!g127) & (!g2986) & (g2987) & (g3056)) + ((g104) & (!g127) & (g2986) & (!g2987) & (!g3056)) + ((g104) & (!g127) & (g2986) & (!g2987) & (g3056)) + ((g104) & (!g127) & (g2986) & (g2987) & (!g3056)) + ((g104) & (!g127) & (g2986) & (g2987) & (g3056)) + ((g104) & (g127) & (!g2986) & (!g2987) & (g3056)) + ((g104) & (g127) & (!g2986) & (g2987) & (!g3056)) + ((g104) & (g127) & (!g2986) & (g2987) & (g3056)) + ((g104) & (g127) & (g2986) & (!g2987) & (!g3056)) + ((g104) & (g127) & (g2986) & (!g2987) & (g3056)) + ((g104) & (g127) & (g2986) & (g2987) & (!g3056)) + ((g104) & (g127) & (g2986) & (g2987) & (g3056)));
	assign g3058 = (((!g68) & (!g87) & (g2984) & (g2985) & (g3057)) + ((!g68) & (g87) & (g2984) & (!g2985) & (g3057)) + ((!g68) & (g87) & (g2984) & (g2985) & (!g3057)) + ((!g68) & (g87) & (g2984) & (g2985) & (g3057)) + ((g68) & (!g87) & (!g2984) & (g2985) & (g3057)) + ((g68) & (!g87) & (g2984) & (!g2985) & (!g3057)) + ((g68) & (!g87) & (g2984) & (!g2985) & (g3057)) + ((g68) & (!g87) & (g2984) & (g2985) & (!g3057)) + ((g68) & (!g87) & (g2984) & (g2985) & (g3057)) + ((g68) & (g87) & (!g2984) & (!g2985) & (g3057)) + ((g68) & (g87) & (!g2984) & (g2985) & (!g3057)) + ((g68) & (g87) & (!g2984) & (g2985) & (g3057)) + ((g68) & (g87) & (g2984) & (!g2985) & (!g3057)) + ((g68) & (g87) & (g2984) & (!g2985) & (g3057)) + ((g68) & (g87) & (g2984) & (g2985) & (!g3057)) + ((g68) & (g87) & (g2984) & (g2985) & (g3057)));
	assign g3059 = (((!g39) & (!g54) & (g2982) & (g2983) & (g3058)) + ((!g39) & (g54) & (g2982) & (!g2983) & (g3058)) + ((!g39) & (g54) & (g2982) & (g2983) & (!g3058)) + ((!g39) & (g54) & (g2982) & (g2983) & (g3058)) + ((g39) & (!g54) & (!g2982) & (g2983) & (g3058)) + ((g39) & (!g54) & (g2982) & (!g2983) & (!g3058)) + ((g39) & (!g54) & (g2982) & (!g2983) & (g3058)) + ((g39) & (!g54) & (g2982) & (g2983) & (!g3058)) + ((g39) & (!g54) & (g2982) & (g2983) & (g3058)) + ((g39) & (g54) & (!g2982) & (!g2983) & (g3058)) + ((g39) & (g54) & (!g2982) & (g2983) & (!g3058)) + ((g39) & (g54) & (!g2982) & (g2983) & (g3058)) + ((g39) & (g54) & (g2982) & (!g2983) & (!g3058)) + ((g39) & (g54) & (g2982) & (!g2983) & (g3058)) + ((g39) & (g54) & (g2982) & (g2983) & (!g3058)) + ((g39) & (g54) & (g2982) & (g2983) & (g3058)));
	assign g3060 = (((g1) & (!g2965) & (g2976) & (g2979)) + ((g1) & (g2965) & (!g2976) & (!g2979)) + ((g1) & (g2965) & (!g2976) & (g2979)));
	assign g3061 = (((!g4) & (!g2) & (!g2966) & (!g2973) & (!g2975) & (!g2980)) + ((!g4) & (!g2) & (!g2966) & (!g2973) & (g2975) & (g2980)) + ((!g4) & (!g2) & (!g2966) & (g2973) & (!g2975) & (!g2980)) + ((!g4) & (!g2) & (!g2966) & (g2973) & (g2975) & (g2980)) + ((!g4) & (!g2) & (g2966) & (!g2973) & (!g2975) & (!g2980)) + ((!g4) & (!g2) & (g2966) & (!g2973) & (g2975) & (g2980)) + ((!g4) & (!g2) & (g2966) & (g2973) & (g2975) & (!g2980)) + ((!g4) & (!g2) & (g2966) & (g2973) & (g2975) & (g2980)) + ((!g4) & (g2) & (!g2966) & (!g2973) & (!g2975) & (!g2980)) + ((!g4) & (g2) & (!g2966) & (!g2973) & (g2975) & (g2980)) + ((!g4) & (g2) & (!g2966) & (g2973) & (g2975) & (!g2980)) + ((!g4) & (g2) & (!g2966) & (g2973) & (g2975) & (g2980)) + ((!g4) & (g2) & (g2966) & (!g2973) & (g2975) & (!g2980)) + ((!g4) & (g2) & (g2966) & (!g2973) & (g2975) & (g2980)) + ((!g4) & (g2) & (g2966) & (g2973) & (g2975) & (!g2980)) + ((!g4) & (g2) & (g2966) & (g2973) & (g2975) & (g2980)) + ((g4) & (!g2) & (!g2966) & (!g2973) & (g2975) & (!g2980)) + ((g4) & (!g2) & (!g2966) & (!g2973) & (g2975) & (g2980)) + ((g4) & (!g2) & (!g2966) & (g2973) & (g2975) & (!g2980)) + ((g4) & (!g2) & (!g2966) & (g2973) & (g2975) & (g2980)) + ((g4) & (!g2) & (g2966) & (!g2973) & (g2975) & (!g2980)) + ((g4) & (!g2) & (g2966) & (!g2973) & (g2975) & (g2980)) + ((g4) & (!g2) & (g2966) & (g2973) & (!g2975) & (!g2980)) + ((g4) & (!g2) & (g2966) & (g2973) & (g2975) & (g2980)) + ((g4) & (g2) & (!g2966) & (!g2973) & (g2975) & (!g2980)) + ((g4) & (g2) & (!g2966) & (!g2973) & (g2975) & (g2980)) + ((g4) & (g2) & (!g2966) & (g2973) & (!g2975) & (!g2980)) + ((g4) & (g2) & (!g2966) & (g2973) & (g2975) & (g2980)) + ((g4) & (g2) & (g2966) & (!g2973) & (!g2975) & (!g2980)) + ((g4) & (g2) & (g2966) & (!g2973) & (g2975) & (g2980)) + ((g4) & (g2) & (g2966) & (g2973) & (!g2975) & (!g2980)) + ((g4) & (g2) & (g2966) & (g2973) & (g2975) & (g2980)));
	assign g3062 = (((!g8) & (!g18) & (!g2968) & (g2969) & (g2972) & (!g2980)) + ((!g8) & (!g18) & (g2968) & (!g2969) & (!g2972) & (!g2980)) + ((!g8) & (!g18) & (g2968) & (!g2969) & (!g2972) & (g2980)) + ((!g8) & (!g18) & (g2968) & (!g2969) & (g2972) & (!g2980)) + ((!g8) & (!g18) & (g2968) & (!g2969) & (g2972) & (g2980)) + ((!g8) & (!g18) & (g2968) & (g2969) & (!g2972) & (!g2980)) + ((!g8) & (!g18) & (g2968) & (g2969) & (!g2972) & (g2980)) + ((!g8) & (!g18) & (g2968) & (g2969) & (g2972) & (g2980)) + ((!g8) & (g18) & (!g2968) & (!g2969) & (g2972) & (!g2980)) + ((!g8) & (g18) & (!g2968) & (g2969) & (!g2972) & (!g2980)) + ((!g8) & (g18) & (!g2968) & (g2969) & (g2972) & (!g2980)) + ((!g8) & (g18) & (g2968) & (!g2969) & (!g2972) & (!g2980)) + ((!g8) & (g18) & (g2968) & (!g2969) & (!g2972) & (g2980)) + ((!g8) & (g18) & (g2968) & (!g2969) & (g2972) & (g2980)) + ((!g8) & (g18) & (g2968) & (g2969) & (!g2972) & (g2980)) + ((!g8) & (g18) & (g2968) & (g2969) & (g2972) & (g2980)) + ((g8) & (!g18) & (!g2968) & (!g2969) & (!g2972) & (!g2980)) + ((g8) & (!g18) & (!g2968) & (!g2969) & (g2972) & (!g2980)) + ((g8) & (!g18) & (!g2968) & (g2969) & (!g2972) & (!g2980)) + ((g8) & (!g18) & (g2968) & (!g2969) & (!g2972) & (g2980)) + ((g8) & (!g18) & (g2968) & (!g2969) & (g2972) & (g2980)) + ((g8) & (!g18) & (g2968) & (g2969) & (!g2972) & (g2980)) + ((g8) & (!g18) & (g2968) & (g2969) & (g2972) & (!g2980)) + ((g8) & (!g18) & (g2968) & (g2969) & (g2972) & (g2980)) + ((g8) & (g18) & (!g2968) & (!g2969) & (!g2972) & (!g2980)) + ((g8) & (g18) & (g2968) & (!g2969) & (!g2972) & (g2980)) + ((g8) & (g18) & (g2968) & (!g2969) & (g2972) & (!g2980)) + ((g8) & (g18) & (g2968) & (!g2969) & (g2972) & (g2980)) + ((g8) & (g18) & (g2968) & (g2969) & (!g2972) & (!g2980)) + ((g8) & (g18) & (g2968) & (g2969) & (!g2972) & (g2980)) + ((g8) & (g18) & (g2968) & (g2969) & (g2972) & (!g2980)) + ((g8) & (g18) & (g2968) & (g2969) & (g2972) & (g2980)));
	assign g3063 = (((!g18) & (!g2969) & (g2972) & (!g2980)) + ((!g18) & (g2969) & (!g2972) & (!g2980)) + ((!g18) & (g2969) & (!g2972) & (g2980)) + ((!g18) & (g2969) & (g2972) & (g2980)) + ((g18) & (!g2969) & (!g2972) & (!g2980)) + ((g18) & (g2969) & (!g2972) & (g2980)) + ((g18) & (g2969) & (g2972) & (!g2980)) + ((g18) & (g2969) & (g2972) & (g2980)));
	assign g3064 = (((!g27) & (!g39) & (!g2971) & (g2866) & (g2964) & (!g2980)) + ((!g27) & (!g39) & (g2971) & (!g2866) & (!g2964) & (!g2980)) + ((!g27) & (!g39) & (g2971) & (!g2866) & (!g2964) & (g2980)) + ((!g27) & (!g39) & (g2971) & (!g2866) & (g2964) & (!g2980)) + ((!g27) & (!g39) & (g2971) & (!g2866) & (g2964) & (g2980)) + ((!g27) & (!g39) & (g2971) & (g2866) & (!g2964) & (!g2980)) + ((!g27) & (!g39) & (g2971) & (g2866) & (!g2964) & (g2980)) + ((!g27) & (!g39) & (g2971) & (g2866) & (g2964) & (g2980)) + ((!g27) & (g39) & (!g2971) & (!g2866) & (g2964) & (!g2980)) + ((!g27) & (g39) & (!g2971) & (g2866) & (!g2964) & (!g2980)) + ((!g27) & (g39) & (!g2971) & (g2866) & (g2964) & (!g2980)) + ((!g27) & (g39) & (g2971) & (!g2866) & (!g2964) & (!g2980)) + ((!g27) & (g39) & (g2971) & (!g2866) & (!g2964) & (g2980)) + ((!g27) & (g39) & (g2971) & (!g2866) & (g2964) & (g2980)) + ((!g27) & (g39) & (g2971) & (g2866) & (!g2964) & (g2980)) + ((!g27) & (g39) & (g2971) & (g2866) & (g2964) & (g2980)) + ((g27) & (!g39) & (!g2971) & (!g2866) & (!g2964) & (!g2980)) + ((g27) & (!g39) & (!g2971) & (!g2866) & (g2964) & (!g2980)) + ((g27) & (!g39) & (!g2971) & (g2866) & (!g2964) & (!g2980)) + ((g27) & (!g39) & (g2971) & (!g2866) & (!g2964) & (g2980)) + ((g27) & (!g39) & (g2971) & (!g2866) & (g2964) & (g2980)) + ((g27) & (!g39) & (g2971) & (g2866) & (!g2964) & (g2980)) + ((g27) & (!g39) & (g2971) & (g2866) & (g2964) & (!g2980)) + ((g27) & (!g39) & (g2971) & (g2866) & (g2964) & (g2980)) + ((g27) & (g39) & (!g2971) & (!g2866) & (!g2964) & (!g2980)) + ((g27) & (g39) & (g2971) & (!g2866) & (!g2964) & (g2980)) + ((g27) & (g39) & (g2971) & (!g2866) & (g2964) & (!g2980)) + ((g27) & (g39) & (g2971) & (!g2866) & (g2964) & (g2980)) + ((g27) & (g39) & (g2971) & (g2866) & (!g2964) & (!g2980)) + ((g27) & (g39) & (g2971) & (g2866) & (!g2964) & (g2980)) + ((g27) & (g39) & (g2971) & (g2866) & (g2964) & (!g2980)) + ((g27) & (g39) & (g2971) & (g2866) & (g2964) & (g2980)));
	assign g3065 = (((!g18) & (!g27) & (g3064) & (g2981) & (g3059)) + ((!g18) & (g27) & (g3064) & (!g2981) & (g3059)) + ((!g18) & (g27) & (g3064) & (g2981) & (!g3059)) + ((!g18) & (g27) & (g3064) & (g2981) & (g3059)) + ((g18) & (!g27) & (!g3064) & (g2981) & (g3059)) + ((g18) & (!g27) & (g3064) & (!g2981) & (!g3059)) + ((g18) & (!g27) & (g3064) & (!g2981) & (g3059)) + ((g18) & (!g27) & (g3064) & (g2981) & (!g3059)) + ((g18) & (!g27) & (g3064) & (g2981) & (g3059)) + ((g18) & (g27) & (!g3064) & (!g2981) & (g3059)) + ((g18) & (g27) & (!g3064) & (g2981) & (!g3059)) + ((g18) & (g27) & (!g3064) & (g2981) & (g3059)) + ((g18) & (g27) & (g3064) & (!g2981) & (!g3059)) + ((g18) & (g27) & (g3064) & (!g2981) & (g3059)) + ((g18) & (g27) & (g3064) & (g2981) & (!g3059)) + ((g18) & (g27) & (g3064) & (g2981) & (g3059)));
	assign g3066 = (((!g2) & (!g8) & (g3062) & (g3063) & (g3065)) + ((!g2) & (g8) & (g3062) & (!g3063) & (g3065)) + ((!g2) & (g8) & (g3062) & (g3063) & (!g3065)) + ((!g2) & (g8) & (g3062) & (g3063) & (g3065)) + ((g2) & (!g8) & (!g3062) & (g3063) & (g3065)) + ((g2) & (!g8) & (g3062) & (!g3063) & (!g3065)) + ((g2) & (!g8) & (g3062) & (!g3063) & (g3065)) + ((g2) & (!g8) & (g3062) & (g3063) & (!g3065)) + ((g2) & (!g8) & (g3062) & (g3063) & (g3065)) + ((g2) & (g8) & (!g3062) & (!g3063) & (g3065)) + ((g2) & (g8) & (!g3062) & (g3063) & (!g3065)) + ((g2) & (g8) & (!g3062) & (g3063) & (g3065)) + ((g2) & (g8) & (g3062) & (!g3063) & (!g3065)) + ((g2) & (g8) & (g3062) & (!g3063) & (g3065)) + ((g2) & (g8) & (g3062) & (g3063) & (!g3065)) + ((g2) & (g8) & (g3062) & (g3063) & (g3065)));
	assign g3067 = (((!g2) & (!g2966) & (g2973) & (!g2980)) + ((!g2) & (g2966) & (!g2973) & (!g2980)) + ((!g2) & (g2966) & (!g2973) & (g2980)) + ((!g2) & (g2966) & (g2973) & (g2980)) + ((g2) & (!g2966) & (!g2973) & (!g2980)) + ((g2) & (g2966) & (!g2973) & (g2980)) + ((g2) & (g2966) & (g2973) & (!g2980)) + ((g2) & (g2966) & (g2973) & (g2980)));
	assign g3068 = (((!g1) & (!g2965) & (!g2976) & (!g2978) & (g2979)) + ((!g1) & (!g2965) & (!g2976) & (g2978) & (!g2979)) + ((!g1) & (!g2965) & (!g2976) & (g2978) & (g2979)) + ((!g1) & (g2965) & (g2976) & (!g2978) & (!g2979)) + ((!g1) & (g2965) & (g2976) & (!g2978) & (g2979)) + ((!g1) & (g2965) & (g2976) & (g2978) & (!g2979)) + ((!g1) & (g2965) & (g2976) & (g2978) & (g2979)) + ((g1) & (!g2965) & (!g2976) & (!g2978) & (g2979)) + ((g1) & (!g2965) & (!g2976) & (g2978) & (g2979)) + ((g1) & (g2965) & (g2976) & (!g2978) & (!g2979)) + ((g1) & (g2965) & (g2976) & (!g2978) & (g2979)) + ((g1) & (g2965) & (g2976) & (g2978) & (!g2979)) + ((g1) & (g2965) & (g2976) & (g2978) & (g2979)));
	assign g3069 = (((!g4) & (!g1) & (!g3061) & (!g3066) & (!g3067) & (!g3068)) + ((!g4) & (g1) & (!g3061) & (!g3066) & (!g3067) & (!g3068)) + ((!g4) & (g1) & (!g3061) & (!g3066) & (!g3067) & (g3068)) + ((!g4) & (g1) & (!g3061) & (!g3066) & (g3067) & (!g3068)) + ((!g4) & (g1) & (!g3061) & (!g3066) & (g3067) & (g3068)) + ((!g4) & (g1) & (!g3061) & (g3066) & (!g3067) & (!g3068)) + ((!g4) & (g1) & (!g3061) & (g3066) & (!g3067) & (g3068)) + ((!g4) & (g1) & (!g3061) & (g3066) & (g3067) & (!g3068)) + ((!g4) & (g1) & (!g3061) & (g3066) & (g3067) & (g3068)) + ((!g4) & (g1) & (g3061) & (!g3066) & (!g3067) & (!g3068)) + ((!g4) & (g1) & (g3061) & (!g3066) & (!g3067) & (g3068)) + ((g4) & (!g1) & (!g3061) & (!g3066) & (!g3067) & (!g3068)) + ((g4) & (!g1) & (!g3061) & (!g3066) & (g3067) & (!g3068)) + ((g4) & (!g1) & (!g3061) & (g3066) & (!g3067) & (!g3068)) + ((g4) & (g1) & (!g3061) & (!g3066) & (!g3067) & (!g3068)) + ((g4) & (g1) & (!g3061) & (!g3066) & (!g3067) & (g3068)) + ((g4) & (g1) & (!g3061) & (!g3066) & (g3067) & (!g3068)) + ((g4) & (g1) & (!g3061) & (!g3066) & (g3067) & (g3068)) + ((g4) & (g1) & (!g3061) & (g3066) & (!g3067) & (!g3068)) + ((g4) & (g1) & (!g3061) & (g3066) & (!g3067) & (g3068)) + ((g4) & (g1) & (!g3061) & (g3066) & (g3067) & (!g3068)) + ((g4) & (g1) & (!g3061) & (g3066) & (g3067) & (g3068)) + ((g4) & (g1) & (g3061) & (!g3066) & (!g3067) & (!g3068)) + ((g4) & (g1) & (g3061) & (!g3066) & (!g3067) & (g3068)) + ((g4) & (g1) & (g3061) & (!g3066) & (g3067) & (!g3068)) + ((g4) & (g1) & (g3061) & (!g3066) & (g3067) & (g3068)) + ((g4) & (g1) & (g3061) & (g3066) & (!g3067) & (!g3068)) + ((g4) & (g1) & (g3061) & (g3066) & (!g3067) & (g3068)));
	assign g3070 = (((!g27) & (!g2981) & (g3059) & (!g3060) & (!g3069)) + ((!g27) & (!g2981) & (g3059) & (g3060) & (!g3069)) + ((!g27) & (!g2981) & (g3059) & (g3060) & (g3069)) + ((!g27) & (g2981) & (!g3059) & (!g3060) & (!g3069)) + ((!g27) & (g2981) & (!g3059) & (!g3060) & (g3069)) + ((!g27) & (g2981) & (!g3059) & (g3060) & (!g3069)) + ((!g27) & (g2981) & (!g3059) & (g3060) & (g3069)) + ((!g27) & (g2981) & (g3059) & (!g3060) & (g3069)) + ((g27) & (!g2981) & (!g3059) & (!g3060) & (!g3069)) + ((g27) & (!g2981) & (!g3059) & (g3060) & (!g3069)) + ((g27) & (!g2981) & (!g3059) & (g3060) & (g3069)) + ((g27) & (g2981) & (!g3059) & (!g3060) & (g3069)) + ((g27) & (g2981) & (g3059) & (!g3060) & (!g3069)) + ((g27) & (g2981) & (g3059) & (!g3060) & (g3069)) + ((g27) & (g2981) & (g3059) & (g3060) & (!g3069)) + ((g27) & (g2981) & (g3059) & (g3060) & (g3069)));
	assign g3071 = (((!g39) & (!g54) & (g2983) & (g3058)) + ((!g39) & (g54) & (!g2983) & (g3058)) + ((!g39) & (g54) & (g2983) & (!g3058)) + ((!g39) & (g54) & (g2983) & (g3058)) + ((g39) & (!g54) & (!g2983) & (!g3058)) + ((g39) & (!g54) & (!g2983) & (g3058)) + ((g39) & (!g54) & (g2983) & (!g3058)) + ((g39) & (g54) & (!g2983) & (!g3058)));
	assign g3072 = (((!g2982) & (!g3060) & (!g3069) & (g3071)) + ((!g2982) & (g3060) & (!g3069) & (g3071)) + ((!g2982) & (g3060) & (g3069) & (g3071)) + ((g2982) & (!g3060) & (!g3069) & (!g3071)) + ((g2982) & (!g3060) & (g3069) & (!g3071)) + ((g2982) & (!g3060) & (g3069) & (g3071)) + ((g2982) & (g3060) & (!g3069) & (!g3071)) + ((g2982) & (g3060) & (g3069) & (!g3071)));
	assign g3073 = (((!g54) & (!g2983) & (g3058) & (!g3060) & (!g3069)) + ((!g54) & (!g2983) & (g3058) & (g3060) & (!g3069)) + ((!g54) & (!g2983) & (g3058) & (g3060) & (g3069)) + ((!g54) & (g2983) & (!g3058) & (!g3060) & (!g3069)) + ((!g54) & (g2983) & (!g3058) & (!g3060) & (g3069)) + ((!g54) & (g2983) & (!g3058) & (g3060) & (!g3069)) + ((!g54) & (g2983) & (!g3058) & (g3060) & (g3069)) + ((!g54) & (g2983) & (g3058) & (!g3060) & (g3069)) + ((g54) & (!g2983) & (!g3058) & (!g3060) & (!g3069)) + ((g54) & (!g2983) & (!g3058) & (g3060) & (!g3069)) + ((g54) & (!g2983) & (!g3058) & (g3060) & (g3069)) + ((g54) & (g2983) & (!g3058) & (!g3060) & (g3069)) + ((g54) & (g2983) & (g3058) & (!g3060) & (!g3069)) + ((g54) & (g2983) & (g3058) & (!g3060) & (g3069)) + ((g54) & (g2983) & (g3058) & (g3060) & (!g3069)) + ((g54) & (g2983) & (g3058) & (g3060) & (g3069)));
	assign g3074 = (((!g68) & (!g87) & (g2985) & (g3057)) + ((!g68) & (g87) & (!g2985) & (g3057)) + ((!g68) & (g87) & (g2985) & (!g3057)) + ((!g68) & (g87) & (g2985) & (g3057)) + ((g68) & (!g87) & (!g2985) & (!g3057)) + ((g68) & (!g87) & (!g2985) & (g3057)) + ((g68) & (!g87) & (g2985) & (!g3057)) + ((g68) & (g87) & (!g2985) & (!g3057)));
	assign g3075 = (((!g2984) & (!g3060) & (!g3069) & (g3074)) + ((!g2984) & (g3060) & (!g3069) & (g3074)) + ((!g2984) & (g3060) & (g3069) & (g3074)) + ((g2984) & (!g3060) & (!g3069) & (!g3074)) + ((g2984) & (!g3060) & (g3069) & (!g3074)) + ((g2984) & (!g3060) & (g3069) & (g3074)) + ((g2984) & (g3060) & (!g3069) & (!g3074)) + ((g2984) & (g3060) & (g3069) & (!g3074)));
	assign g3076 = (((!g87) & (!g2985) & (g3057) & (!g3060) & (!g3069)) + ((!g87) & (!g2985) & (g3057) & (g3060) & (!g3069)) + ((!g87) & (!g2985) & (g3057) & (g3060) & (g3069)) + ((!g87) & (g2985) & (!g3057) & (!g3060) & (!g3069)) + ((!g87) & (g2985) & (!g3057) & (!g3060) & (g3069)) + ((!g87) & (g2985) & (!g3057) & (g3060) & (!g3069)) + ((!g87) & (g2985) & (!g3057) & (g3060) & (g3069)) + ((!g87) & (g2985) & (g3057) & (!g3060) & (g3069)) + ((g87) & (!g2985) & (!g3057) & (!g3060) & (!g3069)) + ((g87) & (!g2985) & (!g3057) & (g3060) & (!g3069)) + ((g87) & (!g2985) & (!g3057) & (g3060) & (g3069)) + ((g87) & (g2985) & (!g3057) & (!g3060) & (g3069)) + ((g87) & (g2985) & (g3057) & (!g3060) & (!g3069)) + ((g87) & (g2985) & (g3057) & (!g3060) & (g3069)) + ((g87) & (g2985) & (g3057) & (g3060) & (!g3069)) + ((g87) & (g2985) & (g3057) & (g3060) & (g3069)));
	assign g3077 = (((!g104) & (!g127) & (g2987) & (g3056)) + ((!g104) & (g127) & (!g2987) & (g3056)) + ((!g104) & (g127) & (g2987) & (!g3056)) + ((!g104) & (g127) & (g2987) & (g3056)) + ((g104) & (!g127) & (!g2987) & (!g3056)) + ((g104) & (!g127) & (!g2987) & (g3056)) + ((g104) & (!g127) & (g2987) & (!g3056)) + ((g104) & (g127) & (!g2987) & (!g3056)));
	assign g3078 = (((!g2986) & (!g3060) & (!g3069) & (g3077)) + ((!g2986) & (g3060) & (!g3069) & (g3077)) + ((!g2986) & (g3060) & (g3069) & (g3077)) + ((g2986) & (!g3060) & (!g3069) & (!g3077)) + ((g2986) & (!g3060) & (g3069) & (!g3077)) + ((g2986) & (!g3060) & (g3069) & (g3077)) + ((g2986) & (g3060) & (!g3069) & (!g3077)) + ((g2986) & (g3060) & (g3069) & (!g3077)));
	assign g3079 = (((!g127) & (!g2987) & (g3056) & (!g3060) & (!g3069)) + ((!g127) & (!g2987) & (g3056) & (g3060) & (!g3069)) + ((!g127) & (!g2987) & (g3056) & (g3060) & (g3069)) + ((!g127) & (g2987) & (!g3056) & (!g3060) & (!g3069)) + ((!g127) & (g2987) & (!g3056) & (!g3060) & (g3069)) + ((!g127) & (g2987) & (!g3056) & (g3060) & (!g3069)) + ((!g127) & (g2987) & (!g3056) & (g3060) & (g3069)) + ((!g127) & (g2987) & (g3056) & (!g3060) & (g3069)) + ((g127) & (!g2987) & (!g3056) & (!g3060) & (!g3069)) + ((g127) & (!g2987) & (!g3056) & (g3060) & (!g3069)) + ((g127) & (!g2987) & (!g3056) & (g3060) & (g3069)) + ((g127) & (g2987) & (!g3056) & (!g3060) & (g3069)) + ((g127) & (g2987) & (g3056) & (!g3060) & (!g3069)) + ((g127) & (g2987) & (g3056) & (!g3060) & (g3069)) + ((g127) & (g2987) & (g3056) & (g3060) & (!g3069)) + ((g127) & (g2987) & (g3056) & (g3060) & (g3069)));
	assign g3080 = (((!g147) & (!g174) & (g2989) & (g3055)) + ((!g147) & (g174) & (!g2989) & (g3055)) + ((!g147) & (g174) & (g2989) & (!g3055)) + ((!g147) & (g174) & (g2989) & (g3055)) + ((g147) & (!g174) & (!g2989) & (!g3055)) + ((g147) & (!g174) & (!g2989) & (g3055)) + ((g147) & (!g174) & (g2989) & (!g3055)) + ((g147) & (g174) & (!g2989) & (!g3055)));
	assign g3081 = (((!g2988) & (!g3060) & (!g3069) & (g3080)) + ((!g2988) & (g3060) & (!g3069) & (g3080)) + ((!g2988) & (g3060) & (g3069) & (g3080)) + ((g2988) & (!g3060) & (!g3069) & (!g3080)) + ((g2988) & (!g3060) & (g3069) & (!g3080)) + ((g2988) & (!g3060) & (g3069) & (g3080)) + ((g2988) & (g3060) & (!g3069) & (!g3080)) + ((g2988) & (g3060) & (g3069) & (!g3080)));
	assign g3082 = (((!g174) & (!g2989) & (g3055) & (!g3060) & (!g3069)) + ((!g174) & (!g2989) & (g3055) & (g3060) & (!g3069)) + ((!g174) & (!g2989) & (g3055) & (g3060) & (g3069)) + ((!g174) & (g2989) & (!g3055) & (!g3060) & (!g3069)) + ((!g174) & (g2989) & (!g3055) & (!g3060) & (g3069)) + ((!g174) & (g2989) & (!g3055) & (g3060) & (!g3069)) + ((!g174) & (g2989) & (!g3055) & (g3060) & (g3069)) + ((!g174) & (g2989) & (g3055) & (!g3060) & (g3069)) + ((g174) & (!g2989) & (!g3055) & (!g3060) & (!g3069)) + ((g174) & (!g2989) & (!g3055) & (g3060) & (!g3069)) + ((g174) & (!g2989) & (!g3055) & (g3060) & (g3069)) + ((g174) & (g2989) & (!g3055) & (!g3060) & (g3069)) + ((g174) & (g2989) & (g3055) & (!g3060) & (!g3069)) + ((g174) & (g2989) & (g3055) & (!g3060) & (g3069)) + ((g174) & (g2989) & (g3055) & (g3060) & (!g3069)) + ((g174) & (g2989) & (g3055) & (g3060) & (g3069)));
	assign g3083 = (((!g198) & (!g229) & (g2991) & (g3054)) + ((!g198) & (g229) & (!g2991) & (g3054)) + ((!g198) & (g229) & (g2991) & (!g3054)) + ((!g198) & (g229) & (g2991) & (g3054)) + ((g198) & (!g229) & (!g2991) & (!g3054)) + ((g198) & (!g229) & (!g2991) & (g3054)) + ((g198) & (!g229) & (g2991) & (!g3054)) + ((g198) & (g229) & (!g2991) & (!g3054)));
	assign g3084 = (((!g2990) & (!g3060) & (!g3069) & (g3083)) + ((!g2990) & (g3060) & (!g3069) & (g3083)) + ((!g2990) & (g3060) & (g3069) & (g3083)) + ((g2990) & (!g3060) & (!g3069) & (!g3083)) + ((g2990) & (!g3060) & (g3069) & (!g3083)) + ((g2990) & (!g3060) & (g3069) & (g3083)) + ((g2990) & (g3060) & (!g3069) & (!g3083)) + ((g2990) & (g3060) & (g3069) & (!g3083)));
	assign g3085 = (((!g229) & (!g2991) & (g3054) & (!g3060) & (!g3069)) + ((!g229) & (!g2991) & (g3054) & (g3060) & (!g3069)) + ((!g229) & (!g2991) & (g3054) & (g3060) & (g3069)) + ((!g229) & (g2991) & (!g3054) & (!g3060) & (!g3069)) + ((!g229) & (g2991) & (!g3054) & (!g3060) & (g3069)) + ((!g229) & (g2991) & (!g3054) & (g3060) & (!g3069)) + ((!g229) & (g2991) & (!g3054) & (g3060) & (g3069)) + ((!g229) & (g2991) & (g3054) & (!g3060) & (g3069)) + ((g229) & (!g2991) & (!g3054) & (!g3060) & (!g3069)) + ((g229) & (!g2991) & (!g3054) & (g3060) & (!g3069)) + ((g229) & (!g2991) & (!g3054) & (g3060) & (g3069)) + ((g229) & (g2991) & (!g3054) & (!g3060) & (g3069)) + ((g229) & (g2991) & (g3054) & (!g3060) & (!g3069)) + ((g229) & (g2991) & (g3054) & (!g3060) & (g3069)) + ((g229) & (g2991) & (g3054) & (g3060) & (!g3069)) + ((g229) & (g2991) & (g3054) & (g3060) & (g3069)));
	assign g3086 = (((!g255) & (!g290) & (g2993) & (g3053)) + ((!g255) & (g290) & (!g2993) & (g3053)) + ((!g255) & (g290) & (g2993) & (!g3053)) + ((!g255) & (g290) & (g2993) & (g3053)) + ((g255) & (!g290) & (!g2993) & (!g3053)) + ((g255) & (!g290) & (!g2993) & (g3053)) + ((g255) & (!g290) & (g2993) & (!g3053)) + ((g255) & (g290) & (!g2993) & (!g3053)));
	assign g3087 = (((!g2992) & (!g3060) & (!g3069) & (g3086)) + ((!g2992) & (g3060) & (!g3069) & (g3086)) + ((!g2992) & (g3060) & (g3069) & (g3086)) + ((g2992) & (!g3060) & (!g3069) & (!g3086)) + ((g2992) & (!g3060) & (g3069) & (!g3086)) + ((g2992) & (!g3060) & (g3069) & (g3086)) + ((g2992) & (g3060) & (!g3069) & (!g3086)) + ((g2992) & (g3060) & (g3069) & (!g3086)));
	assign g3088 = (((!g290) & (!g2993) & (g3053) & (!g3060) & (!g3069)) + ((!g290) & (!g2993) & (g3053) & (g3060) & (!g3069)) + ((!g290) & (!g2993) & (g3053) & (g3060) & (g3069)) + ((!g290) & (g2993) & (!g3053) & (!g3060) & (!g3069)) + ((!g290) & (g2993) & (!g3053) & (!g3060) & (g3069)) + ((!g290) & (g2993) & (!g3053) & (g3060) & (!g3069)) + ((!g290) & (g2993) & (!g3053) & (g3060) & (g3069)) + ((!g290) & (g2993) & (g3053) & (!g3060) & (g3069)) + ((g290) & (!g2993) & (!g3053) & (!g3060) & (!g3069)) + ((g290) & (!g2993) & (!g3053) & (g3060) & (!g3069)) + ((g290) & (!g2993) & (!g3053) & (g3060) & (g3069)) + ((g290) & (g2993) & (!g3053) & (!g3060) & (g3069)) + ((g290) & (g2993) & (g3053) & (!g3060) & (!g3069)) + ((g290) & (g2993) & (g3053) & (!g3060) & (g3069)) + ((g290) & (g2993) & (g3053) & (g3060) & (!g3069)) + ((g290) & (g2993) & (g3053) & (g3060) & (g3069)));
	assign g3089 = (((!g319) & (!g358) & (g2995) & (g3052)) + ((!g319) & (g358) & (!g2995) & (g3052)) + ((!g319) & (g358) & (g2995) & (!g3052)) + ((!g319) & (g358) & (g2995) & (g3052)) + ((g319) & (!g358) & (!g2995) & (!g3052)) + ((g319) & (!g358) & (!g2995) & (g3052)) + ((g319) & (!g358) & (g2995) & (!g3052)) + ((g319) & (g358) & (!g2995) & (!g3052)));
	assign g3090 = (((!g2994) & (!g3060) & (!g3069) & (g3089)) + ((!g2994) & (g3060) & (!g3069) & (g3089)) + ((!g2994) & (g3060) & (g3069) & (g3089)) + ((g2994) & (!g3060) & (!g3069) & (!g3089)) + ((g2994) & (!g3060) & (g3069) & (!g3089)) + ((g2994) & (!g3060) & (g3069) & (g3089)) + ((g2994) & (g3060) & (!g3069) & (!g3089)) + ((g2994) & (g3060) & (g3069) & (!g3089)));
	assign g3091 = (((!g358) & (!g2995) & (g3052) & (!g3060) & (!g3069)) + ((!g358) & (!g2995) & (g3052) & (g3060) & (!g3069)) + ((!g358) & (!g2995) & (g3052) & (g3060) & (g3069)) + ((!g358) & (g2995) & (!g3052) & (!g3060) & (!g3069)) + ((!g358) & (g2995) & (!g3052) & (!g3060) & (g3069)) + ((!g358) & (g2995) & (!g3052) & (g3060) & (!g3069)) + ((!g358) & (g2995) & (!g3052) & (g3060) & (g3069)) + ((!g358) & (g2995) & (g3052) & (!g3060) & (g3069)) + ((g358) & (!g2995) & (!g3052) & (!g3060) & (!g3069)) + ((g358) & (!g2995) & (!g3052) & (g3060) & (!g3069)) + ((g358) & (!g2995) & (!g3052) & (g3060) & (g3069)) + ((g358) & (g2995) & (!g3052) & (!g3060) & (g3069)) + ((g358) & (g2995) & (g3052) & (!g3060) & (!g3069)) + ((g358) & (g2995) & (g3052) & (!g3060) & (g3069)) + ((g358) & (g2995) & (g3052) & (g3060) & (!g3069)) + ((g358) & (g2995) & (g3052) & (g3060) & (g3069)));
	assign g3092 = (((!g390) & (!g433) & (g2997) & (g3051)) + ((!g390) & (g433) & (!g2997) & (g3051)) + ((!g390) & (g433) & (g2997) & (!g3051)) + ((!g390) & (g433) & (g2997) & (g3051)) + ((g390) & (!g433) & (!g2997) & (!g3051)) + ((g390) & (!g433) & (!g2997) & (g3051)) + ((g390) & (!g433) & (g2997) & (!g3051)) + ((g390) & (g433) & (!g2997) & (!g3051)));
	assign g3093 = (((!g2996) & (!g3060) & (!g3069) & (g3092)) + ((!g2996) & (g3060) & (!g3069) & (g3092)) + ((!g2996) & (g3060) & (g3069) & (g3092)) + ((g2996) & (!g3060) & (!g3069) & (!g3092)) + ((g2996) & (!g3060) & (g3069) & (!g3092)) + ((g2996) & (!g3060) & (g3069) & (g3092)) + ((g2996) & (g3060) & (!g3069) & (!g3092)) + ((g2996) & (g3060) & (g3069) & (!g3092)));
	assign g3094 = (((!g433) & (!g2997) & (g3051) & (!g3060) & (!g3069)) + ((!g433) & (!g2997) & (g3051) & (g3060) & (!g3069)) + ((!g433) & (!g2997) & (g3051) & (g3060) & (g3069)) + ((!g433) & (g2997) & (!g3051) & (!g3060) & (!g3069)) + ((!g433) & (g2997) & (!g3051) & (!g3060) & (g3069)) + ((!g433) & (g2997) & (!g3051) & (g3060) & (!g3069)) + ((!g433) & (g2997) & (!g3051) & (g3060) & (g3069)) + ((!g433) & (g2997) & (g3051) & (!g3060) & (g3069)) + ((g433) & (!g2997) & (!g3051) & (!g3060) & (!g3069)) + ((g433) & (!g2997) & (!g3051) & (g3060) & (!g3069)) + ((g433) & (!g2997) & (!g3051) & (g3060) & (g3069)) + ((g433) & (g2997) & (!g3051) & (!g3060) & (g3069)) + ((g433) & (g2997) & (g3051) & (!g3060) & (!g3069)) + ((g433) & (g2997) & (g3051) & (!g3060) & (g3069)) + ((g433) & (g2997) & (g3051) & (g3060) & (!g3069)) + ((g433) & (g2997) & (g3051) & (g3060) & (g3069)));
	assign g3095 = (((!g468) & (!g515) & (g2999) & (g3050)) + ((!g468) & (g515) & (!g2999) & (g3050)) + ((!g468) & (g515) & (g2999) & (!g3050)) + ((!g468) & (g515) & (g2999) & (g3050)) + ((g468) & (!g515) & (!g2999) & (!g3050)) + ((g468) & (!g515) & (!g2999) & (g3050)) + ((g468) & (!g515) & (g2999) & (!g3050)) + ((g468) & (g515) & (!g2999) & (!g3050)));
	assign g3096 = (((!g2998) & (!g3060) & (!g3069) & (g3095)) + ((!g2998) & (g3060) & (!g3069) & (g3095)) + ((!g2998) & (g3060) & (g3069) & (g3095)) + ((g2998) & (!g3060) & (!g3069) & (!g3095)) + ((g2998) & (!g3060) & (g3069) & (!g3095)) + ((g2998) & (!g3060) & (g3069) & (g3095)) + ((g2998) & (g3060) & (!g3069) & (!g3095)) + ((g2998) & (g3060) & (g3069) & (!g3095)));
	assign g3097 = (((!g515) & (!g2999) & (g3050) & (!g3060) & (!g3069)) + ((!g515) & (!g2999) & (g3050) & (g3060) & (!g3069)) + ((!g515) & (!g2999) & (g3050) & (g3060) & (g3069)) + ((!g515) & (g2999) & (!g3050) & (!g3060) & (!g3069)) + ((!g515) & (g2999) & (!g3050) & (!g3060) & (g3069)) + ((!g515) & (g2999) & (!g3050) & (g3060) & (!g3069)) + ((!g515) & (g2999) & (!g3050) & (g3060) & (g3069)) + ((!g515) & (g2999) & (g3050) & (!g3060) & (g3069)) + ((g515) & (!g2999) & (!g3050) & (!g3060) & (!g3069)) + ((g515) & (!g2999) & (!g3050) & (g3060) & (!g3069)) + ((g515) & (!g2999) & (!g3050) & (g3060) & (g3069)) + ((g515) & (g2999) & (!g3050) & (!g3060) & (g3069)) + ((g515) & (g2999) & (g3050) & (!g3060) & (!g3069)) + ((g515) & (g2999) & (g3050) & (!g3060) & (g3069)) + ((g515) & (g2999) & (g3050) & (g3060) & (!g3069)) + ((g515) & (g2999) & (g3050) & (g3060) & (g3069)));
	assign g3098 = (((!g553) & (!g604) & (g3001) & (g3049)) + ((!g553) & (g604) & (!g3001) & (g3049)) + ((!g553) & (g604) & (g3001) & (!g3049)) + ((!g553) & (g604) & (g3001) & (g3049)) + ((g553) & (!g604) & (!g3001) & (!g3049)) + ((g553) & (!g604) & (!g3001) & (g3049)) + ((g553) & (!g604) & (g3001) & (!g3049)) + ((g553) & (g604) & (!g3001) & (!g3049)));
	assign g3099 = (((!g3000) & (!g3060) & (!g3069) & (g3098)) + ((!g3000) & (g3060) & (!g3069) & (g3098)) + ((!g3000) & (g3060) & (g3069) & (g3098)) + ((g3000) & (!g3060) & (!g3069) & (!g3098)) + ((g3000) & (!g3060) & (g3069) & (!g3098)) + ((g3000) & (!g3060) & (g3069) & (g3098)) + ((g3000) & (g3060) & (!g3069) & (!g3098)) + ((g3000) & (g3060) & (g3069) & (!g3098)));
	assign g3100 = (((!g604) & (!g3001) & (g3049) & (!g3060) & (!g3069)) + ((!g604) & (!g3001) & (g3049) & (g3060) & (!g3069)) + ((!g604) & (!g3001) & (g3049) & (g3060) & (g3069)) + ((!g604) & (g3001) & (!g3049) & (!g3060) & (!g3069)) + ((!g604) & (g3001) & (!g3049) & (!g3060) & (g3069)) + ((!g604) & (g3001) & (!g3049) & (g3060) & (!g3069)) + ((!g604) & (g3001) & (!g3049) & (g3060) & (g3069)) + ((!g604) & (g3001) & (g3049) & (!g3060) & (g3069)) + ((g604) & (!g3001) & (!g3049) & (!g3060) & (!g3069)) + ((g604) & (!g3001) & (!g3049) & (g3060) & (!g3069)) + ((g604) & (!g3001) & (!g3049) & (g3060) & (g3069)) + ((g604) & (g3001) & (!g3049) & (!g3060) & (g3069)) + ((g604) & (g3001) & (g3049) & (!g3060) & (!g3069)) + ((g604) & (g3001) & (g3049) & (!g3060) & (g3069)) + ((g604) & (g3001) & (g3049) & (g3060) & (!g3069)) + ((g604) & (g3001) & (g3049) & (g3060) & (g3069)));
	assign g3101 = (((!g645) & (!g700) & (g3003) & (g3048)) + ((!g645) & (g700) & (!g3003) & (g3048)) + ((!g645) & (g700) & (g3003) & (!g3048)) + ((!g645) & (g700) & (g3003) & (g3048)) + ((g645) & (!g700) & (!g3003) & (!g3048)) + ((g645) & (!g700) & (!g3003) & (g3048)) + ((g645) & (!g700) & (g3003) & (!g3048)) + ((g645) & (g700) & (!g3003) & (!g3048)));
	assign g3102 = (((!g3002) & (!g3060) & (!g3069) & (g3101)) + ((!g3002) & (g3060) & (!g3069) & (g3101)) + ((!g3002) & (g3060) & (g3069) & (g3101)) + ((g3002) & (!g3060) & (!g3069) & (!g3101)) + ((g3002) & (!g3060) & (g3069) & (!g3101)) + ((g3002) & (!g3060) & (g3069) & (g3101)) + ((g3002) & (g3060) & (!g3069) & (!g3101)) + ((g3002) & (g3060) & (g3069) & (!g3101)));
	assign g3103 = (((!g700) & (!g3003) & (g3048) & (!g3060) & (!g3069)) + ((!g700) & (!g3003) & (g3048) & (g3060) & (!g3069)) + ((!g700) & (!g3003) & (g3048) & (g3060) & (g3069)) + ((!g700) & (g3003) & (!g3048) & (!g3060) & (!g3069)) + ((!g700) & (g3003) & (!g3048) & (!g3060) & (g3069)) + ((!g700) & (g3003) & (!g3048) & (g3060) & (!g3069)) + ((!g700) & (g3003) & (!g3048) & (g3060) & (g3069)) + ((!g700) & (g3003) & (g3048) & (!g3060) & (g3069)) + ((g700) & (!g3003) & (!g3048) & (!g3060) & (!g3069)) + ((g700) & (!g3003) & (!g3048) & (g3060) & (!g3069)) + ((g700) & (!g3003) & (!g3048) & (g3060) & (g3069)) + ((g700) & (g3003) & (!g3048) & (!g3060) & (g3069)) + ((g700) & (g3003) & (g3048) & (!g3060) & (!g3069)) + ((g700) & (g3003) & (g3048) & (!g3060) & (g3069)) + ((g700) & (g3003) & (g3048) & (g3060) & (!g3069)) + ((g700) & (g3003) & (g3048) & (g3060) & (g3069)));
	assign g3104 = (((!g744) & (!g803) & (g3005) & (g3047)) + ((!g744) & (g803) & (!g3005) & (g3047)) + ((!g744) & (g803) & (g3005) & (!g3047)) + ((!g744) & (g803) & (g3005) & (g3047)) + ((g744) & (!g803) & (!g3005) & (!g3047)) + ((g744) & (!g803) & (!g3005) & (g3047)) + ((g744) & (!g803) & (g3005) & (!g3047)) + ((g744) & (g803) & (!g3005) & (!g3047)));
	assign g3105 = (((!g3004) & (!g3060) & (!g3069) & (g3104)) + ((!g3004) & (g3060) & (!g3069) & (g3104)) + ((!g3004) & (g3060) & (g3069) & (g3104)) + ((g3004) & (!g3060) & (!g3069) & (!g3104)) + ((g3004) & (!g3060) & (g3069) & (!g3104)) + ((g3004) & (!g3060) & (g3069) & (g3104)) + ((g3004) & (g3060) & (!g3069) & (!g3104)) + ((g3004) & (g3060) & (g3069) & (!g3104)));
	assign g3106 = (((!g803) & (!g3005) & (g3047) & (!g3060) & (!g3069)) + ((!g803) & (!g3005) & (g3047) & (g3060) & (!g3069)) + ((!g803) & (!g3005) & (g3047) & (g3060) & (g3069)) + ((!g803) & (g3005) & (!g3047) & (!g3060) & (!g3069)) + ((!g803) & (g3005) & (!g3047) & (!g3060) & (g3069)) + ((!g803) & (g3005) & (!g3047) & (g3060) & (!g3069)) + ((!g803) & (g3005) & (!g3047) & (g3060) & (g3069)) + ((!g803) & (g3005) & (g3047) & (!g3060) & (g3069)) + ((g803) & (!g3005) & (!g3047) & (!g3060) & (!g3069)) + ((g803) & (!g3005) & (!g3047) & (g3060) & (!g3069)) + ((g803) & (!g3005) & (!g3047) & (g3060) & (g3069)) + ((g803) & (g3005) & (!g3047) & (!g3060) & (g3069)) + ((g803) & (g3005) & (g3047) & (!g3060) & (!g3069)) + ((g803) & (g3005) & (g3047) & (!g3060) & (g3069)) + ((g803) & (g3005) & (g3047) & (g3060) & (!g3069)) + ((g803) & (g3005) & (g3047) & (g3060) & (g3069)));
	assign g3107 = (((!g851) & (!g914) & (g3007) & (g3046)) + ((!g851) & (g914) & (!g3007) & (g3046)) + ((!g851) & (g914) & (g3007) & (!g3046)) + ((!g851) & (g914) & (g3007) & (g3046)) + ((g851) & (!g914) & (!g3007) & (!g3046)) + ((g851) & (!g914) & (!g3007) & (g3046)) + ((g851) & (!g914) & (g3007) & (!g3046)) + ((g851) & (g914) & (!g3007) & (!g3046)));
	assign g3108 = (((!g3006) & (!g3060) & (!g3069) & (g3107)) + ((!g3006) & (g3060) & (!g3069) & (g3107)) + ((!g3006) & (g3060) & (g3069) & (g3107)) + ((g3006) & (!g3060) & (!g3069) & (!g3107)) + ((g3006) & (!g3060) & (g3069) & (!g3107)) + ((g3006) & (!g3060) & (g3069) & (g3107)) + ((g3006) & (g3060) & (!g3069) & (!g3107)) + ((g3006) & (g3060) & (g3069) & (!g3107)));
	assign g3109 = (((!g914) & (!g3007) & (g3046) & (!g3060) & (!g3069)) + ((!g914) & (!g3007) & (g3046) & (g3060) & (!g3069)) + ((!g914) & (!g3007) & (g3046) & (g3060) & (g3069)) + ((!g914) & (g3007) & (!g3046) & (!g3060) & (!g3069)) + ((!g914) & (g3007) & (!g3046) & (!g3060) & (g3069)) + ((!g914) & (g3007) & (!g3046) & (g3060) & (!g3069)) + ((!g914) & (g3007) & (!g3046) & (g3060) & (g3069)) + ((!g914) & (g3007) & (g3046) & (!g3060) & (g3069)) + ((g914) & (!g3007) & (!g3046) & (!g3060) & (!g3069)) + ((g914) & (!g3007) & (!g3046) & (g3060) & (!g3069)) + ((g914) & (!g3007) & (!g3046) & (g3060) & (g3069)) + ((g914) & (g3007) & (!g3046) & (!g3060) & (g3069)) + ((g914) & (g3007) & (g3046) & (!g3060) & (!g3069)) + ((g914) & (g3007) & (g3046) & (!g3060) & (g3069)) + ((g914) & (g3007) & (g3046) & (g3060) & (!g3069)) + ((g914) & (g3007) & (g3046) & (g3060) & (g3069)));
	assign g3110 = (((!g1032) & (!g1030) & (g3009) & (g3045)) + ((!g1032) & (g1030) & (!g3009) & (g3045)) + ((!g1032) & (g1030) & (g3009) & (!g3045)) + ((!g1032) & (g1030) & (g3009) & (g3045)) + ((g1032) & (!g1030) & (!g3009) & (!g3045)) + ((g1032) & (!g1030) & (!g3009) & (g3045)) + ((g1032) & (!g1030) & (g3009) & (!g3045)) + ((g1032) & (g1030) & (!g3009) & (!g3045)));
	assign g3111 = (((!g3008) & (!g3060) & (!g3069) & (g3110)) + ((!g3008) & (g3060) & (!g3069) & (g3110)) + ((!g3008) & (g3060) & (g3069) & (g3110)) + ((g3008) & (!g3060) & (!g3069) & (!g3110)) + ((g3008) & (!g3060) & (g3069) & (!g3110)) + ((g3008) & (!g3060) & (g3069) & (g3110)) + ((g3008) & (g3060) & (!g3069) & (!g3110)) + ((g3008) & (g3060) & (g3069) & (!g3110)));
	assign g3112 = (((!g1030) & (!g3009) & (g3045) & (!g3060) & (!g3069)) + ((!g1030) & (!g3009) & (g3045) & (g3060) & (!g3069)) + ((!g1030) & (!g3009) & (g3045) & (g3060) & (g3069)) + ((!g1030) & (g3009) & (!g3045) & (!g3060) & (!g3069)) + ((!g1030) & (g3009) & (!g3045) & (!g3060) & (g3069)) + ((!g1030) & (g3009) & (!g3045) & (g3060) & (!g3069)) + ((!g1030) & (g3009) & (!g3045) & (g3060) & (g3069)) + ((!g1030) & (g3009) & (g3045) & (!g3060) & (g3069)) + ((g1030) & (!g3009) & (!g3045) & (!g3060) & (!g3069)) + ((g1030) & (!g3009) & (!g3045) & (g3060) & (!g3069)) + ((g1030) & (!g3009) & (!g3045) & (g3060) & (g3069)) + ((g1030) & (g3009) & (!g3045) & (!g3060) & (g3069)) + ((g1030) & (g3009) & (g3045) & (!g3060) & (!g3069)) + ((g1030) & (g3009) & (g3045) & (!g3060) & (g3069)) + ((g1030) & (g3009) & (g3045) & (g3060) & (!g3069)) + ((g1030) & (g3009) & (g3045) & (g3060) & (g3069)));
	assign g3113 = (((!g1160) & (!g1154) & (g3011) & (g3044)) + ((!g1160) & (g1154) & (!g3011) & (g3044)) + ((!g1160) & (g1154) & (g3011) & (!g3044)) + ((!g1160) & (g1154) & (g3011) & (g3044)) + ((g1160) & (!g1154) & (!g3011) & (!g3044)) + ((g1160) & (!g1154) & (!g3011) & (g3044)) + ((g1160) & (!g1154) & (g3011) & (!g3044)) + ((g1160) & (g1154) & (!g3011) & (!g3044)));
	assign g3114 = (((!g3010) & (!g3060) & (!g3069) & (g3113)) + ((!g3010) & (g3060) & (!g3069) & (g3113)) + ((!g3010) & (g3060) & (g3069) & (g3113)) + ((g3010) & (!g3060) & (!g3069) & (!g3113)) + ((g3010) & (!g3060) & (g3069) & (!g3113)) + ((g3010) & (!g3060) & (g3069) & (g3113)) + ((g3010) & (g3060) & (!g3069) & (!g3113)) + ((g3010) & (g3060) & (g3069) & (!g3113)));
	assign g3115 = (((!g1154) & (!g3011) & (g3044) & (!g3060) & (!g3069)) + ((!g1154) & (!g3011) & (g3044) & (g3060) & (!g3069)) + ((!g1154) & (!g3011) & (g3044) & (g3060) & (g3069)) + ((!g1154) & (g3011) & (!g3044) & (!g3060) & (!g3069)) + ((!g1154) & (g3011) & (!g3044) & (!g3060) & (g3069)) + ((!g1154) & (g3011) & (!g3044) & (g3060) & (!g3069)) + ((!g1154) & (g3011) & (!g3044) & (g3060) & (g3069)) + ((!g1154) & (g3011) & (g3044) & (!g3060) & (g3069)) + ((g1154) & (!g3011) & (!g3044) & (!g3060) & (!g3069)) + ((g1154) & (!g3011) & (!g3044) & (g3060) & (!g3069)) + ((g1154) & (!g3011) & (!g3044) & (g3060) & (g3069)) + ((g1154) & (g3011) & (!g3044) & (!g3060) & (g3069)) + ((g1154) & (g3011) & (g3044) & (!g3060) & (!g3069)) + ((g1154) & (g3011) & (g3044) & (!g3060) & (g3069)) + ((g1154) & (g3011) & (g3044) & (g3060) & (!g3069)) + ((g1154) & (g3011) & (g3044) & (g3060) & (g3069)));
	assign g3116 = (((!g1295) & (!g1285) & (g3013) & (g3043)) + ((!g1295) & (g1285) & (!g3013) & (g3043)) + ((!g1295) & (g1285) & (g3013) & (!g3043)) + ((!g1295) & (g1285) & (g3013) & (g3043)) + ((g1295) & (!g1285) & (!g3013) & (!g3043)) + ((g1295) & (!g1285) & (!g3013) & (g3043)) + ((g1295) & (!g1285) & (g3013) & (!g3043)) + ((g1295) & (g1285) & (!g3013) & (!g3043)));
	assign g3117 = (((!g3012) & (!g3060) & (!g3069) & (g3116)) + ((!g3012) & (g3060) & (!g3069) & (g3116)) + ((!g3012) & (g3060) & (g3069) & (g3116)) + ((g3012) & (!g3060) & (!g3069) & (!g3116)) + ((g3012) & (!g3060) & (g3069) & (!g3116)) + ((g3012) & (!g3060) & (g3069) & (g3116)) + ((g3012) & (g3060) & (!g3069) & (!g3116)) + ((g3012) & (g3060) & (g3069) & (!g3116)));
	assign g3118 = (((!g1285) & (!g3013) & (g3043) & (!g3060) & (!g3069)) + ((!g1285) & (!g3013) & (g3043) & (g3060) & (!g3069)) + ((!g1285) & (!g3013) & (g3043) & (g3060) & (g3069)) + ((!g1285) & (g3013) & (!g3043) & (!g3060) & (!g3069)) + ((!g1285) & (g3013) & (!g3043) & (!g3060) & (g3069)) + ((!g1285) & (g3013) & (!g3043) & (g3060) & (!g3069)) + ((!g1285) & (g3013) & (!g3043) & (g3060) & (g3069)) + ((!g1285) & (g3013) & (g3043) & (!g3060) & (g3069)) + ((g1285) & (!g3013) & (!g3043) & (!g3060) & (!g3069)) + ((g1285) & (!g3013) & (!g3043) & (g3060) & (!g3069)) + ((g1285) & (!g3013) & (!g3043) & (g3060) & (g3069)) + ((g1285) & (g3013) & (!g3043) & (!g3060) & (g3069)) + ((g1285) & (g3013) & (g3043) & (!g3060) & (!g3069)) + ((g1285) & (g3013) & (g3043) & (!g3060) & (g3069)) + ((g1285) & (g3013) & (g3043) & (g3060) & (!g3069)) + ((g1285) & (g3013) & (g3043) & (g3060) & (g3069)));
	assign g3119 = (((!g1437) & (!g1423) & (g3015) & (g3042)) + ((!g1437) & (g1423) & (!g3015) & (g3042)) + ((!g1437) & (g1423) & (g3015) & (!g3042)) + ((!g1437) & (g1423) & (g3015) & (g3042)) + ((g1437) & (!g1423) & (!g3015) & (!g3042)) + ((g1437) & (!g1423) & (!g3015) & (g3042)) + ((g1437) & (!g1423) & (g3015) & (!g3042)) + ((g1437) & (g1423) & (!g3015) & (!g3042)));
	assign g3120 = (((!g3014) & (!g3060) & (!g3069) & (g3119)) + ((!g3014) & (g3060) & (!g3069) & (g3119)) + ((!g3014) & (g3060) & (g3069) & (g3119)) + ((g3014) & (!g3060) & (!g3069) & (!g3119)) + ((g3014) & (!g3060) & (g3069) & (!g3119)) + ((g3014) & (!g3060) & (g3069) & (g3119)) + ((g3014) & (g3060) & (!g3069) & (!g3119)) + ((g3014) & (g3060) & (g3069) & (!g3119)));
	assign g3121 = (((!g1423) & (!g3015) & (g3042) & (!g3060) & (!g3069)) + ((!g1423) & (!g3015) & (g3042) & (g3060) & (!g3069)) + ((!g1423) & (!g3015) & (g3042) & (g3060) & (g3069)) + ((!g1423) & (g3015) & (!g3042) & (!g3060) & (!g3069)) + ((!g1423) & (g3015) & (!g3042) & (!g3060) & (g3069)) + ((!g1423) & (g3015) & (!g3042) & (g3060) & (!g3069)) + ((!g1423) & (g3015) & (!g3042) & (g3060) & (g3069)) + ((!g1423) & (g3015) & (g3042) & (!g3060) & (g3069)) + ((g1423) & (!g3015) & (!g3042) & (!g3060) & (!g3069)) + ((g1423) & (!g3015) & (!g3042) & (g3060) & (!g3069)) + ((g1423) & (!g3015) & (!g3042) & (g3060) & (g3069)) + ((g1423) & (g3015) & (!g3042) & (!g3060) & (g3069)) + ((g1423) & (g3015) & (g3042) & (!g3060) & (!g3069)) + ((g1423) & (g3015) & (g3042) & (!g3060) & (g3069)) + ((g1423) & (g3015) & (g3042) & (g3060) & (!g3069)) + ((g1423) & (g3015) & (g3042) & (g3060) & (g3069)));
	assign g3122 = (((!g1586) & (!g1568) & (g3017) & (g3041)) + ((!g1586) & (g1568) & (!g3017) & (g3041)) + ((!g1586) & (g1568) & (g3017) & (!g3041)) + ((!g1586) & (g1568) & (g3017) & (g3041)) + ((g1586) & (!g1568) & (!g3017) & (!g3041)) + ((g1586) & (!g1568) & (!g3017) & (g3041)) + ((g1586) & (!g1568) & (g3017) & (!g3041)) + ((g1586) & (g1568) & (!g3017) & (!g3041)));
	assign g3123 = (((!g3016) & (!g3060) & (!g3069) & (g3122)) + ((!g3016) & (g3060) & (!g3069) & (g3122)) + ((!g3016) & (g3060) & (g3069) & (g3122)) + ((g3016) & (!g3060) & (!g3069) & (!g3122)) + ((g3016) & (!g3060) & (g3069) & (!g3122)) + ((g3016) & (!g3060) & (g3069) & (g3122)) + ((g3016) & (g3060) & (!g3069) & (!g3122)) + ((g3016) & (g3060) & (g3069) & (!g3122)));
	assign g3124 = (((!g1568) & (!g3017) & (g3041) & (!g3060) & (!g3069)) + ((!g1568) & (!g3017) & (g3041) & (g3060) & (!g3069)) + ((!g1568) & (!g3017) & (g3041) & (g3060) & (g3069)) + ((!g1568) & (g3017) & (!g3041) & (!g3060) & (!g3069)) + ((!g1568) & (g3017) & (!g3041) & (!g3060) & (g3069)) + ((!g1568) & (g3017) & (!g3041) & (g3060) & (!g3069)) + ((!g1568) & (g3017) & (!g3041) & (g3060) & (g3069)) + ((!g1568) & (g3017) & (g3041) & (!g3060) & (g3069)) + ((g1568) & (!g3017) & (!g3041) & (!g3060) & (!g3069)) + ((g1568) & (!g3017) & (!g3041) & (g3060) & (!g3069)) + ((g1568) & (!g3017) & (!g3041) & (g3060) & (g3069)) + ((g1568) & (g3017) & (!g3041) & (!g3060) & (g3069)) + ((g1568) & (g3017) & (g3041) & (!g3060) & (!g3069)) + ((g1568) & (g3017) & (g3041) & (!g3060) & (g3069)) + ((g1568) & (g3017) & (g3041) & (g3060) & (!g3069)) + ((g1568) & (g3017) & (g3041) & (g3060) & (g3069)));
	assign g3125 = (((!g1742) & (!g1720) & (g3019) & (g3040)) + ((!g1742) & (g1720) & (!g3019) & (g3040)) + ((!g1742) & (g1720) & (g3019) & (!g3040)) + ((!g1742) & (g1720) & (g3019) & (g3040)) + ((g1742) & (!g1720) & (!g3019) & (!g3040)) + ((g1742) & (!g1720) & (!g3019) & (g3040)) + ((g1742) & (!g1720) & (g3019) & (!g3040)) + ((g1742) & (g1720) & (!g3019) & (!g3040)));
	assign g3126 = (((!g3018) & (!g3060) & (!g3069) & (g3125)) + ((!g3018) & (g3060) & (!g3069) & (g3125)) + ((!g3018) & (g3060) & (g3069) & (g3125)) + ((g3018) & (!g3060) & (!g3069) & (!g3125)) + ((g3018) & (!g3060) & (g3069) & (!g3125)) + ((g3018) & (!g3060) & (g3069) & (g3125)) + ((g3018) & (g3060) & (!g3069) & (!g3125)) + ((g3018) & (g3060) & (g3069) & (!g3125)));
	assign g3127 = (((!g1720) & (!g3019) & (g3040) & (!g3060) & (!g3069)) + ((!g1720) & (!g3019) & (g3040) & (g3060) & (!g3069)) + ((!g1720) & (!g3019) & (g3040) & (g3060) & (g3069)) + ((!g1720) & (g3019) & (!g3040) & (!g3060) & (!g3069)) + ((!g1720) & (g3019) & (!g3040) & (!g3060) & (g3069)) + ((!g1720) & (g3019) & (!g3040) & (g3060) & (!g3069)) + ((!g1720) & (g3019) & (!g3040) & (g3060) & (g3069)) + ((!g1720) & (g3019) & (g3040) & (!g3060) & (g3069)) + ((g1720) & (!g3019) & (!g3040) & (!g3060) & (!g3069)) + ((g1720) & (!g3019) & (!g3040) & (g3060) & (!g3069)) + ((g1720) & (!g3019) & (!g3040) & (g3060) & (g3069)) + ((g1720) & (g3019) & (!g3040) & (!g3060) & (g3069)) + ((g1720) & (g3019) & (g3040) & (!g3060) & (!g3069)) + ((g1720) & (g3019) & (g3040) & (!g3060) & (g3069)) + ((g1720) & (g3019) & (g3040) & (g3060) & (!g3069)) + ((g1720) & (g3019) & (g3040) & (g3060) & (g3069)));
	assign g3128 = (((!g1905) & (!g1879) & (g3021) & (g3039)) + ((!g1905) & (g1879) & (!g3021) & (g3039)) + ((!g1905) & (g1879) & (g3021) & (!g3039)) + ((!g1905) & (g1879) & (g3021) & (g3039)) + ((g1905) & (!g1879) & (!g3021) & (!g3039)) + ((g1905) & (!g1879) & (!g3021) & (g3039)) + ((g1905) & (!g1879) & (g3021) & (!g3039)) + ((g1905) & (g1879) & (!g3021) & (!g3039)));
	assign g3129 = (((!g3020) & (!g3060) & (!g3069) & (g3128)) + ((!g3020) & (g3060) & (!g3069) & (g3128)) + ((!g3020) & (g3060) & (g3069) & (g3128)) + ((g3020) & (!g3060) & (!g3069) & (!g3128)) + ((g3020) & (!g3060) & (g3069) & (!g3128)) + ((g3020) & (!g3060) & (g3069) & (g3128)) + ((g3020) & (g3060) & (!g3069) & (!g3128)) + ((g3020) & (g3060) & (g3069) & (!g3128)));
	assign g3130 = (((!g1879) & (!g3021) & (g3039) & (!g3060) & (!g3069)) + ((!g1879) & (!g3021) & (g3039) & (g3060) & (!g3069)) + ((!g1879) & (!g3021) & (g3039) & (g3060) & (g3069)) + ((!g1879) & (g3021) & (!g3039) & (!g3060) & (!g3069)) + ((!g1879) & (g3021) & (!g3039) & (!g3060) & (g3069)) + ((!g1879) & (g3021) & (!g3039) & (g3060) & (!g3069)) + ((!g1879) & (g3021) & (!g3039) & (g3060) & (g3069)) + ((!g1879) & (g3021) & (g3039) & (!g3060) & (g3069)) + ((g1879) & (!g3021) & (!g3039) & (!g3060) & (!g3069)) + ((g1879) & (!g3021) & (!g3039) & (g3060) & (!g3069)) + ((g1879) & (!g3021) & (!g3039) & (g3060) & (g3069)) + ((g1879) & (g3021) & (!g3039) & (!g3060) & (g3069)) + ((g1879) & (g3021) & (g3039) & (!g3060) & (!g3069)) + ((g1879) & (g3021) & (g3039) & (!g3060) & (g3069)) + ((g1879) & (g3021) & (g3039) & (g3060) & (!g3069)) + ((g1879) & (g3021) & (g3039) & (g3060) & (g3069)));
	assign g3131 = (((!g2075) & (!g2045) & (g3023) & (g3038)) + ((!g2075) & (g2045) & (!g3023) & (g3038)) + ((!g2075) & (g2045) & (g3023) & (!g3038)) + ((!g2075) & (g2045) & (g3023) & (g3038)) + ((g2075) & (!g2045) & (!g3023) & (!g3038)) + ((g2075) & (!g2045) & (!g3023) & (g3038)) + ((g2075) & (!g2045) & (g3023) & (!g3038)) + ((g2075) & (g2045) & (!g3023) & (!g3038)));
	assign g3132 = (((!g3022) & (!g3060) & (!g3069) & (g3131)) + ((!g3022) & (g3060) & (!g3069) & (g3131)) + ((!g3022) & (g3060) & (g3069) & (g3131)) + ((g3022) & (!g3060) & (!g3069) & (!g3131)) + ((g3022) & (!g3060) & (g3069) & (!g3131)) + ((g3022) & (!g3060) & (g3069) & (g3131)) + ((g3022) & (g3060) & (!g3069) & (!g3131)) + ((g3022) & (g3060) & (g3069) & (!g3131)));
	assign g3133 = (((!g2045) & (!g3023) & (g3038) & (!g3060) & (!g3069)) + ((!g2045) & (!g3023) & (g3038) & (g3060) & (!g3069)) + ((!g2045) & (!g3023) & (g3038) & (g3060) & (g3069)) + ((!g2045) & (g3023) & (!g3038) & (!g3060) & (!g3069)) + ((!g2045) & (g3023) & (!g3038) & (!g3060) & (g3069)) + ((!g2045) & (g3023) & (!g3038) & (g3060) & (!g3069)) + ((!g2045) & (g3023) & (!g3038) & (g3060) & (g3069)) + ((!g2045) & (g3023) & (g3038) & (!g3060) & (g3069)) + ((g2045) & (!g3023) & (!g3038) & (!g3060) & (!g3069)) + ((g2045) & (!g3023) & (!g3038) & (g3060) & (!g3069)) + ((g2045) & (!g3023) & (!g3038) & (g3060) & (g3069)) + ((g2045) & (g3023) & (!g3038) & (!g3060) & (g3069)) + ((g2045) & (g3023) & (g3038) & (!g3060) & (!g3069)) + ((g2045) & (g3023) & (g3038) & (!g3060) & (g3069)) + ((g2045) & (g3023) & (g3038) & (g3060) & (!g3069)) + ((g2045) & (g3023) & (g3038) & (g3060) & (g3069)));
	assign g3134 = (((!g2252) & (!g2218) & (g3025) & (g3037)) + ((!g2252) & (g2218) & (!g3025) & (g3037)) + ((!g2252) & (g2218) & (g3025) & (!g3037)) + ((!g2252) & (g2218) & (g3025) & (g3037)) + ((g2252) & (!g2218) & (!g3025) & (!g3037)) + ((g2252) & (!g2218) & (!g3025) & (g3037)) + ((g2252) & (!g2218) & (g3025) & (!g3037)) + ((g2252) & (g2218) & (!g3025) & (!g3037)));
	assign g3135 = (((!g3024) & (!g3060) & (!g3069) & (g3134)) + ((!g3024) & (g3060) & (!g3069) & (g3134)) + ((!g3024) & (g3060) & (g3069) & (g3134)) + ((g3024) & (!g3060) & (!g3069) & (!g3134)) + ((g3024) & (!g3060) & (g3069) & (!g3134)) + ((g3024) & (!g3060) & (g3069) & (g3134)) + ((g3024) & (g3060) & (!g3069) & (!g3134)) + ((g3024) & (g3060) & (g3069) & (!g3134)));
	assign g3136 = (((!g2218) & (!g3025) & (g3037) & (!g3060) & (!g3069)) + ((!g2218) & (!g3025) & (g3037) & (g3060) & (!g3069)) + ((!g2218) & (!g3025) & (g3037) & (g3060) & (g3069)) + ((!g2218) & (g3025) & (!g3037) & (!g3060) & (!g3069)) + ((!g2218) & (g3025) & (!g3037) & (!g3060) & (g3069)) + ((!g2218) & (g3025) & (!g3037) & (g3060) & (!g3069)) + ((!g2218) & (g3025) & (!g3037) & (g3060) & (g3069)) + ((!g2218) & (g3025) & (g3037) & (!g3060) & (g3069)) + ((g2218) & (!g3025) & (!g3037) & (!g3060) & (!g3069)) + ((g2218) & (!g3025) & (!g3037) & (g3060) & (!g3069)) + ((g2218) & (!g3025) & (!g3037) & (g3060) & (g3069)) + ((g2218) & (g3025) & (!g3037) & (!g3060) & (g3069)) + ((g2218) & (g3025) & (g3037) & (!g3060) & (!g3069)) + ((g2218) & (g3025) & (g3037) & (!g3060) & (g3069)) + ((g2218) & (g3025) & (g3037) & (g3060) & (!g3069)) + ((g2218) & (g3025) & (g3037) & (g3060) & (g3069)));
	assign g3137 = (((!g2436) & (!g2398) & (g3027) & (g3036)) + ((!g2436) & (g2398) & (!g3027) & (g3036)) + ((!g2436) & (g2398) & (g3027) & (!g3036)) + ((!g2436) & (g2398) & (g3027) & (g3036)) + ((g2436) & (!g2398) & (!g3027) & (!g3036)) + ((g2436) & (!g2398) & (!g3027) & (g3036)) + ((g2436) & (!g2398) & (g3027) & (!g3036)) + ((g2436) & (g2398) & (!g3027) & (!g3036)));
	assign g3138 = (((!g3026) & (!g3060) & (!g3069) & (g3137)) + ((!g3026) & (g3060) & (!g3069) & (g3137)) + ((!g3026) & (g3060) & (g3069) & (g3137)) + ((g3026) & (!g3060) & (!g3069) & (!g3137)) + ((g3026) & (!g3060) & (g3069) & (!g3137)) + ((g3026) & (!g3060) & (g3069) & (g3137)) + ((g3026) & (g3060) & (!g3069) & (!g3137)) + ((g3026) & (g3060) & (g3069) & (!g3137)));
	assign g3139 = (((!g2398) & (!g3027) & (g3036) & (!g3060) & (!g3069)) + ((!g2398) & (!g3027) & (g3036) & (g3060) & (!g3069)) + ((!g2398) & (!g3027) & (g3036) & (g3060) & (g3069)) + ((!g2398) & (g3027) & (!g3036) & (!g3060) & (!g3069)) + ((!g2398) & (g3027) & (!g3036) & (!g3060) & (g3069)) + ((!g2398) & (g3027) & (!g3036) & (g3060) & (!g3069)) + ((!g2398) & (g3027) & (!g3036) & (g3060) & (g3069)) + ((!g2398) & (g3027) & (g3036) & (!g3060) & (g3069)) + ((g2398) & (!g3027) & (!g3036) & (!g3060) & (!g3069)) + ((g2398) & (!g3027) & (!g3036) & (g3060) & (!g3069)) + ((g2398) & (!g3027) & (!g3036) & (g3060) & (g3069)) + ((g2398) & (g3027) & (!g3036) & (!g3060) & (g3069)) + ((g2398) & (g3027) & (g3036) & (!g3060) & (!g3069)) + ((g2398) & (g3027) & (g3036) & (!g3060) & (g3069)) + ((g2398) & (g3027) & (g3036) & (g3060) & (!g3069)) + ((g2398) & (g3027) & (g3036) & (g3060) & (g3069)));
	assign g3140 = (((!g2627) & (!g2585) & (g3029) & (g3035)) + ((!g2627) & (g2585) & (!g3029) & (g3035)) + ((!g2627) & (g2585) & (g3029) & (!g3035)) + ((!g2627) & (g2585) & (g3029) & (g3035)) + ((g2627) & (!g2585) & (!g3029) & (!g3035)) + ((g2627) & (!g2585) & (!g3029) & (g3035)) + ((g2627) & (!g2585) & (g3029) & (!g3035)) + ((g2627) & (g2585) & (!g3029) & (!g3035)));
	assign g3141 = (((!g3028) & (!g3060) & (!g3069) & (g3140)) + ((!g3028) & (g3060) & (!g3069) & (g3140)) + ((!g3028) & (g3060) & (g3069) & (g3140)) + ((g3028) & (!g3060) & (!g3069) & (!g3140)) + ((g3028) & (!g3060) & (g3069) & (!g3140)) + ((g3028) & (!g3060) & (g3069) & (g3140)) + ((g3028) & (g3060) & (!g3069) & (!g3140)) + ((g3028) & (g3060) & (g3069) & (!g3140)));
	assign g3142 = (((!g2585) & (!g3029) & (g3035) & (!g3060) & (!g3069)) + ((!g2585) & (!g3029) & (g3035) & (g3060) & (!g3069)) + ((!g2585) & (!g3029) & (g3035) & (g3060) & (g3069)) + ((!g2585) & (g3029) & (!g3035) & (!g3060) & (!g3069)) + ((!g2585) & (g3029) & (!g3035) & (!g3060) & (g3069)) + ((!g2585) & (g3029) & (!g3035) & (g3060) & (!g3069)) + ((!g2585) & (g3029) & (!g3035) & (g3060) & (g3069)) + ((!g2585) & (g3029) & (g3035) & (!g3060) & (g3069)) + ((g2585) & (!g3029) & (!g3035) & (!g3060) & (!g3069)) + ((g2585) & (!g3029) & (!g3035) & (g3060) & (!g3069)) + ((g2585) & (!g3029) & (!g3035) & (g3060) & (g3069)) + ((g2585) & (g3029) & (!g3035) & (!g3060) & (g3069)) + ((g2585) & (g3029) & (g3035) & (!g3060) & (!g3069)) + ((g2585) & (g3029) & (g3035) & (!g3060) & (g3069)) + ((g2585) & (g3029) & (g3035) & (g3060) & (!g3069)) + ((g2585) & (g3029) & (g3035) & (g3060) & (g3069)));
	assign g3143 = (((!g2825) & (!g2779) & (g3032) & (g3034)) + ((!g2825) & (g2779) & (!g3032) & (g3034)) + ((!g2825) & (g2779) & (g3032) & (!g3034)) + ((!g2825) & (g2779) & (g3032) & (g3034)) + ((g2825) & (!g2779) & (!g3032) & (!g3034)) + ((g2825) & (!g2779) & (!g3032) & (g3034)) + ((g2825) & (!g2779) & (g3032) & (!g3034)) + ((g2825) & (g2779) & (!g3032) & (!g3034)));
	assign g3144 = (((!g3031) & (!g3060) & (!g3069) & (g3143)) + ((!g3031) & (g3060) & (!g3069) & (g3143)) + ((!g3031) & (g3060) & (g3069) & (g3143)) + ((g3031) & (!g3060) & (!g3069) & (!g3143)) + ((g3031) & (!g3060) & (g3069) & (!g3143)) + ((g3031) & (!g3060) & (g3069) & (g3143)) + ((g3031) & (g3060) & (!g3069) & (!g3143)) + ((g3031) & (g3060) & (g3069) & (!g3143)));
	assign g3145 = (((!g2779) & (!g3032) & (g3034) & (!g3060) & (!g3069)) + ((!g2779) & (!g3032) & (g3034) & (g3060) & (!g3069)) + ((!g2779) & (!g3032) & (g3034) & (g3060) & (g3069)) + ((!g2779) & (g3032) & (!g3034) & (!g3060) & (!g3069)) + ((!g2779) & (g3032) & (!g3034) & (!g3060) & (g3069)) + ((!g2779) & (g3032) & (!g3034) & (g3060) & (!g3069)) + ((!g2779) & (g3032) & (!g3034) & (g3060) & (g3069)) + ((!g2779) & (g3032) & (g3034) & (!g3060) & (g3069)) + ((g2779) & (!g3032) & (!g3034) & (!g3060) & (!g3069)) + ((g2779) & (!g3032) & (!g3034) & (g3060) & (!g3069)) + ((g2779) & (!g3032) & (!g3034) & (g3060) & (g3069)) + ((g2779) & (g3032) & (!g3034) & (!g3060) & (g3069)) + ((g2779) & (g3032) & (g3034) & (!g3060) & (!g3069)) + ((g2779) & (g3032) & (g3034) & (!g3060) & (g3069)) + ((g2779) & (g3032) & (g3034) & (g3060) & (!g3069)) + ((g2779) & (g3032) & (g3034) & (g3060) & (g3069)));
	assign g3146 = (((!g3030) & (!ax12x) & (!g2980) & (g3033)) + ((!g3030) & (!ax12x) & (g2980) & (g3033)) + ((!g3030) & (ax12x) & (!g2980) & (!g3033)) + ((!g3030) & (ax12x) & (!g2980) & (g3033)) + ((g3030) & (!ax12x) & (!g2980) & (!g3033)) + ((g3030) & (!ax12x) & (g2980) & (!g3033)) + ((g3030) & (ax12x) & (g2980) & (!g3033)) + ((g3030) & (ax12x) & (g2980) & (g3033)));
	assign g3147 = (((!ax12x) & (!ax13x) & (!g2980) & (!g3060) & (!g3069) & (g3146)) + ((!ax12x) & (!ax13x) & (!g2980) & (!g3060) & (g3069) & (!g3146)) + ((!ax12x) & (!ax13x) & (!g2980) & (!g3060) & (g3069) & (g3146)) + ((!ax12x) & (!ax13x) & (!g2980) & (g3060) & (!g3069) & (g3146)) + ((!ax12x) & (!ax13x) & (!g2980) & (g3060) & (g3069) & (g3146)) + ((!ax12x) & (!ax13x) & (g2980) & (!g3060) & (!g3069) & (!g3146)) + ((!ax12x) & (!ax13x) & (g2980) & (g3060) & (!g3069) & (!g3146)) + ((!ax12x) & (!ax13x) & (g2980) & (g3060) & (g3069) & (!g3146)) + ((!ax12x) & (ax13x) & (!g2980) & (!g3060) & (!g3069) & (!g3146)) + ((!ax12x) & (ax13x) & (!g2980) & (g3060) & (!g3069) & (!g3146)) + ((!ax12x) & (ax13x) & (!g2980) & (g3060) & (g3069) & (!g3146)) + ((!ax12x) & (ax13x) & (g2980) & (!g3060) & (!g3069) & (g3146)) + ((!ax12x) & (ax13x) & (g2980) & (!g3060) & (g3069) & (!g3146)) + ((!ax12x) & (ax13x) & (g2980) & (!g3060) & (g3069) & (g3146)) + ((!ax12x) & (ax13x) & (g2980) & (g3060) & (!g3069) & (g3146)) + ((!ax12x) & (ax13x) & (g2980) & (g3060) & (g3069) & (g3146)) + ((ax12x) & (!ax13x) & (!g2980) & (!g3060) & (!g3069) & (!g3146)) + ((ax12x) & (!ax13x) & (!g2980) & (g3060) & (!g3069) & (!g3146)) + ((ax12x) & (!ax13x) & (!g2980) & (g3060) & (g3069) & (!g3146)) + ((ax12x) & (!ax13x) & (g2980) & (!g3060) & (!g3069) & (!g3146)) + ((ax12x) & (!ax13x) & (g2980) & (g3060) & (!g3069) & (!g3146)) + ((ax12x) & (!ax13x) & (g2980) & (g3060) & (g3069) & (!g3146)) + ((ax12x) & (ax13x) & (!g2980) & (!g3060) & (!g3069) & (g3146)) + ((ax12x) & (ax13x) & (!g2980) & (!g3060) & (g3069) & (!g3146)) + ((ax12x) & (ax13x) & (!g2980) & (!g3060) & (g3069) & (g3146)) + ((ax12x) & (ax13x) & (!g2980) & (g3060) & (!g3069) & (g3146)) + ((ax12x) & (ax13x) & (!g2980) & (g3060) & (g3069) & (g3146)) + ((ax12x) & (ax13x) & (g2980) & (!g3060) & (!g3069) & (g3146)) + ((ax12x) & (ax13x) & (g2980) & (!g3060) & (g3069) & (!g3146)) + ((ax12x) & (ax13x) & (g2980) & (!g3060) & (g3069) & (g3146)) + ((ax12x) & (ax13x) & (g2980) & (g3060) & (!g3069) & (g3146)) + ((ax12x) & (ax13x) & (g2980) & (g3060) & (g3069) & (g3146)));
	assign g3148 = (((!ax12x) & (!g2980) & (!g3033) & (!g3060) & (g3069)) + ((!ax12x) & (!g2980) & (g3033) & (!g3060) & (!g3069)) + ((!ax12x) & (!g2980) & (g3033) & (!g3060) & (g3069)) + ((!ax12x) & (!g2980) & (g3033) & (g3060) & (!g3069)) + ((!ax12x) & (!g2980) & (g3033) & (g3060) & (g3069)) + ((!ax12x) & (g2980) & (g3033) & (!g3060) & (!g3069)) + ((!ax12x) & (g2980) & (g3033) & (g3060) & (!g3069)) + ((!ax12x) & (g2980) & (g3033) & (g3060) & (g3069)) + ((ax12x) & (!g2980) & (!g3033) & (!g3060) & (!g3069)) + ((ax12x) & (!g2980) & (!g3033) & (g3060) & (!g3069)) + ((ax12x) & (!g2980) & (!g3033) & (g3060) & (g3069)) + ((ax12x) & (g2980) & (!g3033) & (!g3060) & (!g3069)) + ((ax12x) & (g2980) & (!g3033) & (!g3060) & (g3069)) + ((ax12x) & (g2980) & (!g3033) & (g3060) & (!g3069)) + ((ax12x) & (g2980) & (!g3033) & (g3060) & (g3069)) + ((ax12x) & (g2980) & (g3033) & (!g3060) & (g3069)));
	assign g3149 = (((!ax8x) & (!ax9x)));
	assign g3150 = (((!g2980) & (!ax10x) & (!ax11x) & (!g3060) & (!g3069) & (!g3149)) + ((!g2980) & (!ax10x) & (!ax11x) & (g3060) & (!g3069) & (!g3149)) + ((!g2980) & (!ax10x) & (!ax11x) & (g3060) & (g3069) & (!g3149)) + ((!g2980) & (!ax10x) & (ax11x) & (!g3060) & (g3069) & (!g3149)) + ((!g2980) & (ax10x) & (ax11x) & (!g3060) & (g3069) & (!g3149)) + ((!g2980) & (ax10x) & (ax11x) & (!g3060) & (g3069) & (g3149)) + ((g2980) & (!ax10x) & (!ax11x) & (!g3060) & (!g3069) & (!g3149)) + ((g2980) & (!ax10x) & (!ax11x) & (!g3060) & (!g3069) & (g3149)) + ((g2980) & (!ax10x) & (!ax11x) & (!g3060) & (g3069) & (!g3149)) + ((g2980) & (!ax10x) & (!ax11x) & (g3060) & (!g3069) & (!g3149)) + ((g2980) & (!ax10x) & (!ax11x) & (g3060) & (!g3069) & (g3149)) + ((g2980) & (!ax10x) & (!ax11x) & (g3060) & (g3069) & (!g3149)) + ((g2980) & (!ax10x) & (!ax11x) & (g3060) & (g3069) & (g3149)) + ((g2980) & (!ax10x) & (ax11x) & (!g3060) & (!g3069) & (!g3149)) + ((g2980) & (!ax10x) & (ax11x) & (!g3060) & (g3069) & (!g3149)) + ((g2980) & (!ax10x) & (ax11x) & (!g3060) & (g3069) & (g3149)) + ((g2980) & (!ax10x) & (ax11x) & (g3060) & (!g3069) & (!g3149)) + ((g2980) & (!ax10x) & (ax11x) & (g3060) & (g3069) & (!g3149)) + ((g2980) & (ax10x) & (!ax11x) & (!g3060) & (g3069) & (!g3149)) + ((g2980) & (ax10x) & (!ax11x) & (!g3060) & (g3069) & (g3149)) + ((g2980) & (ax10x) & (ax11x) & (!g3060) & (!g3069) & (!g3149)) + ((g2980) & (ax10x) & (ax11x) & (!g3060) & (!g3069) & (g3149)) + ((g2980) & (ax10x) & (ax11x) & (!g3060) & (g3069) & (!g3149)) + ((g2980) & (ax10x) & (ax11x) & (!g3060) & (g3069) & (g3149)) + ((g2980) & (ax10x) & (ax11x) & (g3060) & (!g3069) & (!g3149)) + ((g2980) & (ax10x) & (ax11x) & (g3060) & (!g3069) & (g3149)) + ((g2980) & (ax10x) & (ax11x) & (g3060) & (g3069) & (!g3149)) + ((g2980) & (ax10x) & (ax11x) & (g3060) & (g3069) & (g3149)));
	assign g3151 = (((!g2779) & (!g3030) & (g3147) & (g3148) & (g3150)) + ((!g2779) & (g3030) & (g3147) & (!g3148) & (g3150)) + ((!g2779) & (g3030) & (g3147) & (g3148) & (!g3150)) + ((!g2779) & (g3030) & (g3147) & (g3148) & (g3150)) + ((g2779) & (!g3030) & (!g3147) & (g3148) & (g3150)) + ((g2779) & (!g3030) & (g3147) & (!g3148) & (!g3150)) + ((g2779) & (!g3030) & (g3147) & (!g3148) & (g3150)) + ((g2779) & (!g3030) & (g3147) & (g3148) & (!g3150)) + ((g2779) & (!g3030) & (g3147) & (g3148) & (g3150)) + ((g2779) & (g3030) & (!g3147) & (!g3148) & (g3150)) + ((g2779) & (g3030) & (!g3147) & (g3148) & (!g3150)) + ((g2779) & (g3030) & (!g3147) & (g3148) & (g3150)) + ((g2779) & (g3030) & (g3147) & (!g3148) & (!g3150)) + ((g2779) & (g3030) & (g3147) & (!g3148) & (g3150)) + ((g2779) & (g3030) & (g3147) & (g3148) & (!g3150)) + ((g2779) & (g3030) & (g3147) & (g3148) & (g3150)));
	assign g3152 = (((!g2585) & (!g2825) & (g3144) & (g3145) & (g3151)) + ((!g2585) & (g2825) & (g3144) & (!g3145) & (g3151)) + ((!g2585) & (g2825) & (g3144) & (g3145) & (!g3151)) + ((!g2585) & (g2825) & (g3144) & (g3145) & (g3151)) + ((g2585) & (!g2825) & (!g3144) & (g3145) & (g3151)) + ((g2585) & (!g2825) & (g3144) & (!g3145) & (!g3151)) + ((g2585) & (!g2825) & (g3144) & (!g3145) & (g3151)) + ((g2585) & (!g2825) & (g3144) & (g3145) & (!g3151)) + ((g2585) & (!g2825) & (g3144) & (g3145) & (g3151)) + ((g2585) & (g2825) & (!g3144) & (!g3145) & (g3151)) + ((g2585) & (g2825) & (!g3144) & (g3145) & (!g3151)) + ((g2585) & (g2825) & (!g3144) & (g3145) & (g3151)) + ((g2585) & (g2825) & (g3144) & (!g3145) & (!g3151)) + ((g2585) & (g2825) & (g3144) & (!g3145) & (g3151)) + ((g2585) & (g2825) & (g3144) & (g3145) & (!g3151)) + ((g2585) & (g2825) & (g3144) & (g3145) & (g3151)));
	assign g3153 = (((!g2398) & (!g2627) & (g3141) & (g3142) & (g3152)) + ((!g2398) & (g2627) & (g3141) & (!g3142) & (g3152)) + ((!g2398) & (g2627) & (g3141) & (g3142) & (!g3152)) + ((!g2398) & (g2627) & (g3141) & (g3142) & (g3152)) + ((g2398) & (!g2627) & (!g3141) & (g3142) & (g3152)) + ((g2398) & (!g2627) & (g3141) & (!g3142) & (!g3152)) + ((g2398) & (!g2627) & (g3141) & (!g3142) & (g3152)) + ((g2398) & (!g2627) & (g3141) & (g3142) & (!g3152)) + ((g2398) & (!g2627) & (g3141) & (g3142) & (g3152)) + ((g2398) & (g2627) & (!g3141) & (!g3142) & (g3152)) + ((g2398) & (g2627) & (!g3141) & (g3142) & (!g3152)) + ((g2398) & (g2627) & (!g3141) & (g3142) & (g3152)) + ((g2398) & (g2627) & (g3141) & (!g3142) & (!g3152)) + ((g2398) & (g2627) & (g3141) & (!g3142) & (g3152)) + ((g2398) & (g2627) & (g3141) & (g3142) & (!g3152)) + ((g2398) & (g2627) & (g3141) & (g3142) & (g3152)));
	assign g3154 = (((!g2218) & (!g2436) & (g3138) & (g3139) & (g3153)) + ((!g2218) & (g2436) & (g3138) & (!g3139) & (g3153)) + ((!g2218) & (g2436) & (g3138) & (g3139) & (!g3153)) + ((!g2218) & (g2436) & (g3138) & (g3139) & (g3153)) + ((g2218) & (!g2436) & (!g3138) & (g3139) & (g3153)) + ((g2218) & (!g2436) & (g3138) & (!g3139) & (!g3153)) + ((g2218) & (!g2436) & (g3138) & (!g3139) & (g3153)) + ((g2218) & (!g2436) & (g3138) & (g3139) & (!g3153)) + ((g2218) & (!g2436) & (g3138) & (g3139) & (g3153)) + ((g2218) & (g2436) & (!g3138) & (!g3139) & (g3153)) + ((g2218) & (g2436) & (!g3138) & (g3139) & (!g3153)) + ((g2218) & (g2436) & (!g3138) & (g3139) & (g3153)) + ((g2218) & (g2436) & (g3138) & (!g3139) & (!g3153)) + ((g2218) & (g2436) & (g3138) & (!g3139) & (g3153)) + ((g2218) & (g2436) & (g3138) & (g3139) & (!g3153)) + ((g2218) & (g2436) & (g3138) & (g3139) & (g3153)));
	assign g3155 = (((!g2045) & (!g2252) & (g3135) & (g3136) & (g3154)) + ((!g2045) & (g2252) & (g3135) & (!g3136) & (g3154)) + ((!g2045) & (g2252) & (g3135) & (g3136) & (!g3154)) + ((!g2045) & (g2252) & (g3135) & (g3136) & (g3154)) + ((g2045) & (!g2252) & (!g3135) & (g3136) & (g3154)) + ((g2045) & (!g2252) & (g3135) & (!g3136) & (!g3154)) + ((g2045) & (!g2252) & (g3135) & (!g3136) & (g3154)) + ((g2045) & (!g2252) & (g3135) & (g3136) & (!g3154)) + ((g2045) & (!g2252) & (g3135) & (g3136) & (g3154)) + ((g2045) & (g2252) & (!g3135) & (!g3136) & (g3154)) + ((g2045) & (g2252) & (!g3135) & (g3136) & (!g3154)) + ((g2045) & (g2252) & (!g3135) & (g3136) & (g3154)) + ((g2045) & (g2252) & (g3135) & (!g3136) & (!g3154)) + ((g2045) & (g2252) & (g3135) & (!g3136) & (g3154)) + ((g2045) & (g2252) & (g3135) & (g3136) & (!g3154)) + ((g2045) & (g2252) & (g3135) & (g3136) & (g3154)));
	assign g3156 = (((!g1879) & (!g2075) & (g3132) & (g3133) & (g3155)) + ((!g1879) & (g2075) & (g3132) & (!g3133) & (g3155)) + ((!g1879) & (g2075) & (g3132) & (g3133) & (!g3155)) + ((!g1879) & (g2075) & (g3132) & (g3133) & (g3155)) + ((g1879) & (!g2075) & (!g3132) & (g3133) & (g3155)) + ((g1879) & (!g2075) & (g3132) & (!g3133) & (!g3155)) + ((g1879) & (!g2075) & (g3132) & (!g3133) & (g3155)) + ((g1879) & (!g2075) & (g3132) & (g3133) & (!g3155)) + ((g1879) & (!g2075) & (g3132) & (g3133) & (g3155)) + ((g1879) & (g2075) & (!g3132) & (!g3133) & (g3155)) + ((g1879) & (g2075) & (!g3132) & (g3133) & (!g3155)) + ((g1879) & (g2075) & (!g3132) & (g3133) & (g3155)) + ((g1879) & (g2075) & (g3132) & (!g3133) & (!g3155)) + ((g1879) & (g2075) & (g3132) & (!g3133) & (g3155)) + ((g1879) & (g2075) & (g3132) & (g3133) & (!g3155)) + ((g1879) & (g2075) & (g3132) & (g3133) & (g3155)));
	assign g3157 = (((!g1720) & (!g1905) & (g3129) & (g3130) & (g3156)) + ((!g1720) & (g1905) & (g3129) & (!g3130) & (g3156)) + ((!g1720) & (g1905) & (g3129) & (g3130) & (!g3156)) + ((!g1720) & (g1905) & (g3129) & (g3130) & (g3156)) + ((g1720) & (!g1905) & (!g3129) & (g3130) & (g3156)) + ((g1720) & (!g1905) & (g3129) & (!g3130) & (!g3156)) + ((g1720) & (!g1905) & (g3129) & (!g3130) & (g3156)) + ((g1720) & (!g1905) & (g3129) & (g3130) & (!g3156)) + ((g1720) & (!g1905) & (g3129) & (g3130) & (g3156)) + ((g1720) & (g1905) & (!g3129) & (!g3130) & (g3156)) + ((g1720) & (g1905) & (!g3129) & (g3130) & (!g3156)) + ((g1720) & (g1905) & (!g3129) & (g3130) & (g3156)) + ((g1720) & (g1905) & (g3129) & (!g3130) & (!g3156)) + ((g1720) & (g1905) & (g3129) & (!g3130) & (g3156)) + ((g1720) & (g1905) & (g3129) & (g3130) & (!g3156)) + ((g1720) & (g1905) & (g3129) & (g3130) & (g3156)));
	assign g3158 = (((!g1568) & (!g1742) & (g3126) & (g3127) & (g3157)) + ((!g1568) & (g1742) & (g3126) & (!g3127) & (g3157)) + ((!g1568) & (g1742) & (g3126) & (g3127) & (!g3157)) + ((!g1568) & (g1742) & (g3126) & (g3127) & (g3157)) + ((g1568) & (!g1742) & (!g3126) & (g3127) & (g3157)) + ((g1568) & (!g1742) & (g3126) & (!g3127) & (!g3157)) + ((g1568) & (!g1742) & (g3126) & (!g3127) & (g3157)) + ((g1568) & (!g1742) & (g3126) & (g3127) & (!g3157)) + ((g1568) & (!g1742) & (g3126) & (g3127) & (g3157)) + ((g1568) & (g1742) & (!g3126) & (!g3127) & (g3157)) + ((g1568) & (g1742) & (!g3126) & (g3127) & (!g3157)) + ((g1568) & (g1742) & (!g3126) & (g3127) & (g3157)) + ((g1568) & (g1742) & (g3126) & (!g3127) & (!g3157)) + ((g1568) & (g1742) & (g3126) & (!g3127) & (g3157)) + ((g1568) & (g1742) & (g3126) & (g3127) & (!g3157)) + ((g1568) & (g1742) & (g3126) & (g3127) & (g3157)));
	assign g3159 = (((!g1423) & (!g1586) & (g3123) & (g3124) & (g3158)) + ((!g1423) & (g1586) & (g3123) & (!g3124) & (g3158)) + ((!g1423) & (g1586) & (g3123) & (g3124) & (!g3158)) + ((!g1423) & (g1586) & (g3123) & (g3124) & (g3158)) + ((g1423) & (!g1586) & (!g3123) & (g3124) & (g3158)) + ((g1423) & (!g1586) & (g3123) & (!g3124) & (!g3158)) + ((g1423) & (!g1586) & (g3123) & (!g3124) & (g3158)) + ((g1423) & (!g1586) & (g3123) & (g3124) & (!g3158)) + ((g1423) & (!g1586) & (g3123) & (g3124) & (g3158)) + ((g1423) & (g1586) & (!g3123) & (!g3124) & (g3158)) + ((g1423) & (g1586) & (!g3123) & (g3124) & (!g3158)) + ((g1423) & (g1586) & (!g3123) & (g3124) & (g3158)) + ((g1423) & (g1586) & (g3123) & (!g3124) & (!g3158)) + ((g1423) & (g1586) & (g3123) & (!g3124) & (g3158)) + ((g1423) & (g1586) & (g3123) & (g3124) & (!g3158)) + ((g1423) & (g1586) & (g3123) & (g3124) & (g3158)));
	assign g3160 = (((!g1285) & (!g1437) & (g3120) & (g3121) & (g3159)) + ((!g1285) & (g1437) & (g3120) & (!g3121) & (g3159)) + ((!g1285) & (g1437) & (g3120) & (g3121) & (!g3159)) + ((!g1285) & (g1437) & (g3120) & (g3121) & (g3159)) + ((g1285) & (!g1437) & (!g3120) & (g3121) & (g3159)) + ((g1285) & (!g1437) & (g3120) & (!g3121) & (!g3159)) + ((g1285) & (!g1437) & (g3120) & (!g3121) & (g3159)) + ((g1285) & (!g1437) & (g3120) & (g3121) & (!g3159)) + ((g1285) & (!g1437) & (g3120) & (g3121) & (g3159)) + ((g1285) & (g1437) & (!g3120) & (!g3121) & (g3159)) + ((g1285) & (g1437) & (!g3120) & (g3121) & (!g3159)) + ((g1285) & (g1437) & (!g3120) & (g3121) & (g3159)) + ((g1285) & (g1437) & (g3120) & (!g3121) & (!g3159)) + ((g1285) & (g1437) & (g3120) & (!g3121) & (g3159)) + ((g1285) & (g1437) & (g3120) & (g3121) & (!g3159)) + ((g1285) & (g1437) & (g3120) & (g3121) & (g3159)));
	assign g3161 = (((!g1154) & (!g1295) & (g3117) & (g3118) & (g3160)) + ((!g1154) & (g1295) & (g3117) & (!g3118) & (g3160)) + ((!g1154) & (g1295) & (g3117) & (g3118) & (!g3160)) + ((!g1154) & (g1295) & (g3117) & (g3118) & (g3160)) + ((g1154) & (!g1295) & (!g3117) & (g3118) & (g3160)) + ((g1154) & (!g1295) & (g3117) & (!g3118) & (!g3160)) + ((g1154) & (!g1295) & (g3117) & (!g3118) & (g3160)) + ((g1154) & (!g1295) & (g3117) & (g3118) & (!g3160)) + ((g1154) & (!g1295) & (g3117) & (g3118) & (g3160)) + ((g1154) & (g1295) & (!g3117) & (!g3118) & (g3160)) + ((g1154) & (g1295) & (!g3117) & (g3118) & (!g3160)) + ((g1154) & (g1295) & (!g3117) & (g3118) & (g3160)) + ((g1154) & (g1295) & (g3117) & (!g3118) & (!g3160)) + ((g1154) & (g1295) & (g3117) & (!g3118) & (g3160)) + ((g1154) & (g1295) & (g3117) & (g3118) & (!g3160)) + ((g1154) & (g1295) & (g3117) & (g3118) & (g3160)));
	assign g3162 = (((!g1030) & (!g1160) & (g3114) & (g3115) & (g3161)) + ((!g1030) & (g1160) & (g3114) & (!g3115) & (g3161)) + ((!g1030) & (g1160) & (g3114) & (g3115) & (!g3161)) + ((!g1030) & (g1160) & (g3114) & (g3115) & (g3161)) + ((g1030) & (!g1160) & (!g3114) & (g3115) & (g3161)) + ((g1030) & (!g1160) & (g3114) & (!g3115) & (!g3161)) + ((g1030) & (!g1160) & (g3114) & (!g3115) & (g3161)) + ((g1030) & (!g1160) & (g3114) & (g3115) & (!g3161)) + ((g1030) & (!g1160) & (g3114) & (g3115) & (g3161)) + ((g1030) & (g1160) & (!g3114) & (!g3115) & (g3161)) + ((g1030) & (g1160) & (!g3114) & (g3115) & (!g3161)) + ((g1030) & (g1160) & (!g3114) & (g3115) & (g3161)) + ((g1030) & (g1160) & (g3114) & (!g3115) & (!g3161)) + ((g1030) & (g1160) & (g3114) & (!g3115) & (g3161)) + ((g1030) & (g1160) & (g3114) & (g3115) & (!g3161)) + ((g1030) & (g1160) & (g3114) & (g3115) & (g3161)));
	assign g3163 = (((!g914) & (!g1032) & (g3111) & (g3112) & (g3162)) + ((!g914) & (g1032) & (g3111) & (!g3112) & (g3162)) + ((!g914) & (g1032) & (g3111) & (g3112) & (!g3162)) + ((!g914) & (g1032) & (g3111) & (g3112) & (g3162)) + ((g914) & (!g1032) & (!g3111) & (g3112) & (g3162)) + ((g914) & (!g1032) & (g3111) & (!g3112) & (!g3162)) + ((g914) & (!g1032) & (g3111) & (!g3112) & (g3162)) + ((g914) & (!g1032) & (g3111) & (g3112) & (!g3162)) + ((g914) & (!g1032) & (g3111) & (g3112) & (g3162)) + ((g914) & (g1032) & (!g3111) & (!g3112) & (g3162)) + ((g914) & (g1032) & (!g3111) & (g3112) & (!g3162)) + ((g914) & (g1032) & (!g3111) & (g3112) & (g3162)) + ((g914) & (g1032) & (g3111) & (!g3112) & (!g3162)) + ((g914) & (g1032) & (g3111) & (!g3112) & (g3162)) + ((g914) & (g1032) & (g3111) & (g3112) & (!g3162)) + ((g914) & (g1032) & (g3111) & (g3112) & (g3162)));
	assign g3164 = (((!g803) & (!g851) & (g3108) & (g3109) & (g3163)) + ((!g803) & (g851) & (g3108) & (!g3109) & (g3163)) + ((!g803) & (g851) & (g3108) & (g3109) & (!g3163)) + ((!g803) & (g851) & (g3108) & (g3109) & (g3163)) + ((g803) & (!g851) & (!g3108) & (g3109) & (g3163)) + ((g803) & (!g851) & (g3108) & (!g3109) & (!g3163)) + ((g803) & (!g851) & (g3108) & (!g3109) & (g3163)) + ((g803) & (!g851) & (g3108) & (g3109) & (!g3163)) + ((g803) & (!g851) & (g3108) & (g3109) & (g3163)) + ((g803) & (g851) & (!g3108) & (!g3109) & (g3163)) + ((g803) & (g851) & (!g3108) & (g3109) & (!g3163)) + ((g803) & (g851) & (!g3108) & (g3109) & (g3163)) + ((g803) & (g851) & (g3108) & (!g3109) & (!g3163)) + ((g803) & (g851) & (g3108) & (!g3109) & (g3163)) + ((g803) & (g851) & (g3108) & (g3109) & (!g3163)) + ((g803) & (g851) & (g3108) & (g3109) & (g3163)));
	assign g3165 = (((!g700) & (!g744) & (g3105) & (g3106) & (g3164)) + ((!g700) & (g744) & (g3105) & (!g3106) & (g3164)) + ((!g700) & (g744) & (g3105) & (g3106) & (!g3164)) + ((!g700) & (g744) & (g3105) & (g3106) & (g3164)) + ((g700) & (!g744) & (!g3105) & (g3106) & (g3164)) + ((g700) & (!g744) & (g3105) & (!g3106) & (!g3164)) + ((g700) & (!g744) & (g3105) & (!g3106) & (g3164)) + ((g700) & (!g744) & (g3105) & (g3106) & (!g3164)) + ((g700) & (!g744) & (g3105) & (g3106) & (g3164)) + ((g700) & (g744) & (!g3105) & (!g3106) & (g3164)) + ((g700) & (g744) & (!g3105) & (g3106) & (!g3164)) + ((g700) & (g744) & (!g3105) & (g3106) & (g3164)) + ((g700) & (g744) & (g3105) & (!g3106) & (!g3164)) + ((g700) & (g744) & (g3105) & (!g3106) & (g3164)) + ((g700) & (g744) & (g3105) & (g3106) & (!g3164)) + ((g700) & (g744) & (g3105) & (g3106) & (g3164)));
	assign g3166 = (((!g604) & (!g645) & (g3102) & (g3103) & (g3165)) + ((!g604) & (g645) & (g3102) & (!g3103) & (g3165)) + ((!g604) & (g645) & (g3102) & (g3103) & (!g3165)) + ((!g604) & (g645) & (g3102) & (g3103) & (g3165)) + ((g604) & (!g645) & (!g3102) & (g3103) & (g3165)) + ((g604) & (!g645) & (g3102) & (!g3103) & (!g3165)) + ((g604) & (!g645) & (g3102) & (!g3103) & (g3165)) + ((g604) & (!g645) & (g3102) & (g3103) & (!g3165)) + ((g604) & (!g645) & (g3102) & (g3103) & (g3165)) + ((g604) & (g645) & (!g3102) & (!g3103) & (g3165)) + ((g604) & (g645) & (!g3102) & (g3103) & (!g3165)) + ((g604) & (g645) & (!g3102) & (g3103) & (g3165)) + ((g604) & (g645) & (g3102) & (!g3103) & (!g3165)) + ((g604) & (g645) & (g3102) & (!g3103) & (g3165)) + ((g604) & (g645) & (g3102) & (g3103) & (!g3165)) + ((g604) & (g645) & (g3102) & (g3103) & (g3165)));
	assign g3167 = (((!g515) & (!g553) & (g3099) & (g3100) & (g3166)) + ((!g515) & (g553) & (g3099) & (!g3100) & (g3166)) + ((!g515) & (g553) & (g3099) & (g3100) & (!g3166)) + ((!g515) & (g553) & (g3099) & (g3100) & (g3166)) + ((g515) & (!g553) & (!g3099) & (g3100) & (g3166)) + ((g515) & (!g553) & (g3099) & (!g3100) & (!g3166)) + ((g515) & (!g553) & (g3099) & (!g3100) & (g3166)) + ((g515) & (!g553) & (g3099) & (g3100) & (!g3166)) + ((g515) & (!g553) & (g3099) & (g3100) & (g3166)) + ((g515) & (g553) & (!g3099) & (!g3100) & (g3166)) + ((g515) & (g553) & (!g3099) & (g3100) & (!g3166)) + ((g515) & (g553) & (!g3099) & (g3100) & (g3166)) + ((g515) & (g553) & (g3099) & (!g3100) & (!g3166)) + ((g515) & (g553) & (g3099) & (!g3100) & (g3166)) + ((g515) & (g553) & (g3099) & (g3100) & (!g3166)) + ((g515) & (g553) & (g3099) & (g3100) & (g3166)));
	assign g3168 = (((!g433) & (!g468) & (g3096) & (g3097) & (g3167)) + ((!g433) & (g468) & (g3096) & (!g3097) & (g3167)) + ((!g433) & (g468) & (g3096) & (g3097) & (!g3167)) + ((!g433) & (g468) & (g3096) & (g3097) & (g3167)) + ((g433) & (!g468) & (!g3096) & (g3097) & (g3167)) + ((g433) & (!g468) & (g3096) & (!g3097) & (!g3167)) + ((g433) & (!g468) & (g3096) & (!g3097) & (g3167)) + ((g433) & (!g468) & (g3096) & (g3097) & (!g3167)) + ((g433) & (!g468) & (g3096) & (g3097) & (g3167)) + ((g433) & (g468) & (!g3096) & (!g3097) & (g3167)) + ((g433) & (g468) & (!g3096) & (g3097) & (!g3167)) + ((g433) & (g468) & (!g3096) & (g3097) & (g3167)) + ((g433) & (g468) & (g3096) & (!g3097) & (!g3167)) + ((g433) & (g468) & (g3096) & (!g3097) & (g3167)) + ((g433) & (g468) & (g3096) & (g3097) & (!g3167)) + ((g433) & (g468) & (g3096) & (g3097) & (g3167)));
	assign g3169 = (((!g358) & (!g390) & (g3093) & (g3094) & (g3168)) + ((!g358) & (g390) & (g3093) & (!g3094) & (g3168)) + ((!g358) & (g390) & (g3093) & (g3094) & (!g3168)) + ((!g358) & (g390) & (g3093) & (g3094) & (g3168)) + ((g358) & (!g390) & (!g3093) & (g3094) & (g3168)) + ((g358) & (!g390) & (g3093) & (!g3094) & (!g3168)) + ((g358) & (!g390) & (g3093) & (!g3094) & (g3168)) + ((g358) & (!g390) & (g3093) & (g3094) & (!g3168)) + ((g358) & (!g390) & (g3093) & (g3094) & (g3168)) + ((g358) & (g390) & (!g3093) & (!g3094) & (g3168)) + ((g358) & (g390) & (!g3093) & (g3094) & (!g3168)) + ((g358) & (g390) & (!g3093) & (g3094) & (g3168)) + ((g358) & (g390) & (g3093) & (!g3094) & (!g3168)) + ((g358) & (g390) & (g3093) & (!g3094) & (g3168)) + ((g358) & (g390) & (g3093) & (g3094) & (!g3168)) + ((g358) & (g390) & (g3093) & (g3094) & (g3168)));
	assign g3170 = (((!g290) & (!g319) & (g3090) & (g3091) & (g3169)) + ((!g290) & (g319) & (g3090) & (!g3091) & (g3169)) + ((!g290) & (g319) & (g3090) & (g3091) & (!g3169)) + ((!g290) & (g319) & (g3090) & (g3091) & (g3169)) + ((g290) & (!g319) & (!g3090) & (g3091) & (g3169)) + ((g290) & (!g319) & (g3090) & (!g3091) & (!g3169)) + ((g290) & (!g319) & (g3090) & (!g3091) & (g3169)) + ((g290) & (!g319) & (g3090) & (g3091) & (!g3169)) + ((g290) & (!g319) & (g3090) & (g3091) & (g3169)) + ((g290) & (g319) & (!g3090) & (!g3091) & (g3169)) + ((g290) & (g319) & (!g3090) & (g3091) & (!g3169)) + ((g290) & (g319) & (!g3090) & (g3091) & (g3169)) + ((g290) & (g319) & (g3090) & (!g3091) & (!g3169)) + ((g290) & (g319) & (g3090) & (!g3091) & (g3169)) + ((g290) & (g319) & (g3090) & (g3091) & (!g3169)) + ((g290) & (g319) & (g3090) & (g3091) & (g3169)));
	assign g3171 = (((!g229) & (!g255) & (g3087) & (g3088) & (g3170)) + ((!g229) & (g255) & (g3087) & (!g3088) & (g3170)) + ((!g229) & (g255) & (g3087) & (g3088) & (!g3170)) + ((!g229) & (g255) & (g3087) & (g3088) & (g3170)) + ((g229) & (!g255) & (!g3087) & (g3088) & (g3170)) + ((g229) & (!g255) & (g3087) & (!g3088) & (!g3170)) + ((g229) & (!g255) & (g3087) & (!g3088) & (g3170)) + ((g229) & (!g255) & (g3087) & (g3088) & (!g3170)) + ((g229) & (!g255) & (g3087) & (g3088) & (g3170)) + ((g229) & (g255) & (!g3087) & (!g3088) & (g3170)) + ((g229) & (g255) & (!g3087) & (g3088) & (!g3170)) + ((g229) & (g255) & (!g3087) & (g3088) & (g3170)) + ((g229) & (g255) & (g3087) & (!g3088) & (!g3170)) + ((g229) & (g255) & (g3087) & (!g3088) & (g3170)) + ((g229) & (g255) & (g3087) & (g3088) & (!g3170)) + ((g229) & (g255) & (g3087) & (g3088) & (g3170)));
	assign g3172 = (((!g174) & (!g198) & (g3084) & (g3085) & (g3171)) + ((!g174) & (g198) & (g3084) & (!g3085) & (g3171)) + ((!g174) & (g198) & (g3084) & (g3085) & (!g3171)) + ((!g174) & (g198) & (g3084) & (g3085) & (g3171)) + ((g174) & (!g198) & (!g3084) & (g3085) & (g3171)) + ((g174) & (!g198) & (g3084) & (!g3085) & (!g3171)) + ((g174) & (!g198) & (g3084) & (!g3085) & (g3171)) + ((g174) & (!g198) & (g3084) & (g3085) & (!g3171)) + ((g174) & (!g198) & (g3084) & (g3085) & (g3171)) + ((g174) & (g198) & (!g3084) & (!g3085) & (g3171)) + ((g174) & (g198) & (!g3084) & (g3085) & (!g3171)) + ((g174) & (g198) & (!g3084) & (g3085) & (g3171)) + ((g174) & (g198) & (g3084) & (!g3085) & (!g3171)) + ((g174) & (g198) & (g3084) & (!g3085) & (g3171)) + ((g174) & (g198) & (g3084) & (g3085) & (!g3171)) + ((g174) & (g198) & (g3084) & (g3085) & (g3171)));
	assign g3173 = (((!g127) & (!g147) & (g3081) & (g3082) & (g3172)) + ((!g127) & (g147) & (g3081) & (!g3082) & (g3172)) + ((!g127) & (g147) & (g3081) & (g3082) & (!g3172)) + ((!g127) & (g147) & (g3081) & (g3082) & (g3172)) + ((g127) & (!g147) & (!g3081) & (g3082) & (g3172)) + ((g127) & (!g147) & (g3081) & (!g3082) & (!g3172)) + ((g127) & (!g147) & (g3081) & (!g3082) & (g3172)) + ((g127) & (!g147) & (g3081) & (g3082) & (!g3172)) + ((g127) & (!g147) & (g3081) & (g3082) & (g3172)) + ((g127) & (g147) & (!g3081) & (!g3082) & (g3172)) + ((g127) & (g147) & (!g3081) & (g3082) & (!g3172)) + ((g127) & (g147) & (!g3081) & (g3082) & (g3172)) + ((g127) & (g147) & (g3081) & (!g3082) & (!g3172)) + ((g127) & (g147) & (g3081) & (!g3082) & (g3172)) + ((g127) & (g147) & (g3081) & (g3082) & (!g3172)) + ((g127) & (g147) & (g3081) & (g3082) & (g3172)));
	assign g3174 = (((!g87) & (!g104) & (g3078) & (g3079) & (g3173)) + ((!g87) & (g104) & (g3078) & (!g3079) & (g3173)) + ((!g87) & (g104) & (g3078) & (g3079) & (!g3173)) + ((!g87) & (g104) & (g3078) & (g3079) & (g3173)) + ((g87) & (!g104) & (!g3078) & (g3079) & (g3173)) + ((g87) & (!g104) & (g3078) & (!g3079) & (!g3173)) + ((g87) & (!g104) & (g3078) & (!g3079) & (g3173)) + ((g87) & (!g104) & (g3078) & (g3079) & (!g3173)) + ((g87) & (!g104) & (g3078) & (g3079) & (g3173)) + ((g87) & (g104) & (!g3078) & (!g3079) & (g3173)) + ((g87) & (g104) & (!g3078) & (g3079) & (!g3173)) + ((g87) & (g104) & (!g3078) & (g3079) & (g3173)) + ((g87) & (g104) & (g3078) & (!g3079) & (!g3173)) + ((g87) & (g104) & (g3078) & (!g3079) & (g3173)) + ((g87) & (g104) & (g3078) & (g3079) & (!g3173)) + ((g87) & (g104) & (g3078) & (g3079) & (g3173)));
	assign g3175 = (((!g54) & (!g68) & (g3075) & (g3076) & (g3174)) + ((!g54) & (g68) & (g3075) & (!g3076) & (g3174)) + ((!g54) & (g68) & (g3075) & (g3076) & (!g3174)) + ((!g54) & (g68) & (g3075) & (g3076) & (g3174)) + ((g54) & (!g68) & (!g3075) & (g3076) & (g3174)) + ((g54) & (!g68) & (g3075) & (!g3076) & (!g3174)) + ((g54) & (!g68) & (g3075) & (!g3076) & (g3174)) + ((g54) & (!g68) & (g3075) & (g3076) & (!g3174)) + ((g54) & (!g68) & (g3075) & (g3076) & (g3174)) + ((g54) & (g68) & (!g3075) & (!g3076) & (g3174)) + ((g54) & (g68) & (!g3075) & (g3076) & (!g3174)) + ((g54) & (g68) & (!g3075) & (g3076) & (g3174)) + ((g54) & (g68) & (g3075) & (!g3076) & (!g3174)) + ((g54) & (g68) & (g3075) & (!g3076) & (g3174)) + ((g54) & (g68) & (g3075) & (g3076) & (!g3174)) + ((g54) & (g68) & (g3075) & (g3076) & (g3174)));
	assign g3176 = (((!g27) & (!g39) & (g3072) & (g3073) & (g3175)) + ((!g27) & (g39) & (g3072) & (!g3073) & (g3175)) + ((!g27) & (g39) & (g3072) & (g3073) & (!g3175)) + ((!g27) & (g39) & (g3072) & (g3073) & (g3175)) + ((g27) & (!g39) & (!g3072) & (g3073) & (g3175)) + ((g27) & (!g39) & (g3072) & (!g3073) & (!g3175)) + ((g27) & (!g39) & (g3072) & (!g3073) & (g3175)) + ((g27) & (!g39) & (g3072) & (g3073) & (!g3175)) + ((g27) & (!g39) & (g3072) & (g3073) & (g3175)) + ((g27) & (g39) & (!g3072) & (!g3073) & (g3175)) + ((g27) & (g39) & (!g3072) & (g3073) & (!g3175)) + ((g27) & (g39) & (!g3072) & (g3073) & (g3175)) + ((g27) & (g39) & (g3072) & (!g3073) & (!g3175)) + ((g27) & (g39) & (g3072) & (!g3073) & (g3175)) + ((g27) & (g39) & (g3072) & (g3073) & (!g3175)) + ((g27) & (g39) & (g3072) & (g3073) & (g3175)));
	assign g3177 = (((!g4) & (!g3066) & (g3067)) + ((!g4) & (g3066) & (!g3067)) + ((!g4) & (g3066) & (g3067)) + ((g4) & (g3066) & (g3067)));
	assign g3178 = (((!g3060) & (g3069)));
	assign g3179 = (((!g4) & (!g3066) & (!g3067) & (!g3060) & (!g3069)) + ((!g4) & (!g3066) & (!g3067) & (g3060) & (!g3069)) + ((!g4) & (!g3066) & (!g3067) & (g3060) & (g3069)) + ((!g4) & (!g3066) & (g3067) & (!g3060) & (g3069)) + ((!g4) & (g3066) & (g3067) & (!g3060) & (!g3069)) + ((!g4) & (g3066) & (g3067) & (!g3060) & (g3069)) + ((!g4) & (g3066) & (g3067) & (g3060) & (!g3069)) + ((!g4) & (g3066) & (g3067) & (g3060) & (g3069)) + ((g4) & (!g3066) & (g3067) & (!g3060) & (!g3069)) + ((g4) & (!g3066) & (g3067) & (!g3060) & (g3069)) + ((g4) & (!g3066) & (g3067) & (g3060) & (!g3069)) + ((g4) & (!g3066) & (g3067) & (g3060) & (g3069)) + ((g4) & (g3066) & (!g3067) & (!g3060) & (!g3069)) + ((g4) & (g3066) & (!g3067) & (g3060) & (!g3069)) + ((g4) & (g3066) & (!g3067) & (g3060) & (g3069)) + ((g4) & (g3066) & (g3067) & (!g3060) & (g3069)));
	assign g3180 = (((!g8) & (!g3063) & (g3065) & (!g3060) & (!g3069)) + ((!g8) & (!g3063) & (g3065) & (g3060) & (!g3069)) + ((!g8) & (!g3063) & (g3065) & (g3060) & (g3069)) + ((!g8) & (g3063) & (!g3065) & (!g3060) & (!g3069)) + ((!g8) & (g3063) & (!g3065) & (!g3060) & (g3069)) + ((!g8) & (g3063) & (!g3065) & (g3060) & (!g3069)) + ((!g8) & (g3063) & (!g3065) & (g3060) & (g3069)) + ((!g8) & (g3063) & (g3065) & (!g3060) & (g3069)) + ((g8) & (!g3063) & (!g3065) & (!g3060) & (!g3069)) + ((g8) & (!g3063) & (!g3065) & (g3060) & (!g3069)) + ((g8) & (!g3063) & (!g3065) & (g3060) & (g3069)) + ((g8) & (g3063) & (!g3065) & (!g3060) & (g3069)) + ((g8) & (g3063) & (g3065) & (!g3060) & (!g3069)) + ((g8) & (g3063) & (g3065) & (!g3060) & (g3069)) + ((g8) & (g3063) & (g3065) & (g3060) & (!g3069)) + ((g8) & (g3063) & (g3065) & (g3060) & (g3069)));
	assign g3181 = (((!g18) & (!g27) & (g2981) & (g3059)) + ((!g18) & (g27) & (!g2981) & (g3059)) + ((!g18) & (g27) & (g2981) & (!g3059)) + ((!g18) & (g27) & (g2981) & (g3059)) + ((g18) & (!g27) & (!g2981) & (!g3059)) + ((g18) & (!g27) & (!g2981) & (g3059)) + ((g18) & (!g27) & (g2981) & (!g3059)) + ((g18) & (g27) & (!g2981) & (!g3059)));
	assign g3182 = (((!g3064) & (!g3060) & (!g3069) & (g3181)) + ((!g3064) & (g3060) & (!g3069) & (g3181)) + ((!g3064) & (g3060) & (g3069) & (g3181)) + ((g3064) & (!g3060) & (!g3069) & (!g3181)) + ((g3064) & (!g3060) & (g3069) & (!g3181)) + ((g3064) & (!g3060) & (g3069) & (g3181)) + ((g3064) & (g3060) & (!g3069) & (!g3181)) + ((g3064) & (g3060) & (g3069) & (!g3181)));
	assign g3183 = (((!g8) & (!g18) & (g3182) & (g3070) & (g3176)) + ((!g8) & (g18) & (g3182) & (!g3070) & (g3176)) + ((!g8) & (g18) & (g3182) & (g3070) & (!g3176)) + ((!g8) & (g18) & (g3182) & (g3070) & (g3176)) + ((g8) & (!g18) & (!g3182) & (g3070) & (g3176)) + ((g8) & (!g18) & (g3182) & (!g3070) & (!g3176)) + ((g8) & (!g18) & (g3182) & (!g3070) & (g3176)) + ((g8) & (!g18) & (g3182) & (g3070) & (!g3176)) + ((g8) & (!g18) & (g3182) & (g3070) & (g3176)) + ((g8) & (g18) & (!g3182) & (!g3070) & (g3176)) + ((g8) & (g18) & (!g3182) & (g3070) & (!g3176)) + ((g8) & (g18) & (!g3182) & (g3070) & (g3176)) + ((g8) & (g18) & (g3182) & (!g3070) & (!g3176)) + ((g8) & (g18) & (g3182) & (!g3070) & (g3176)) + ((g8) & (g18) & (g3182) & (g3070) & (!g3176)) + ((g8) & (g18) & (g3182) & (g3070) & (g3176)));
	assign g3184 = (((!g2) & (!g8) & (g3063) & (g3065)) + ((!g2) & (g8) & (!g3063) & (g3065)) + ((!g2) & (g8) & (g3063) & (!g3065)) + ((!g2) & (g8) & (g3063) & (g3065)) + ((g2) & (!g8) & (!g3063) & (!g3065)) + ((g2) & (!g8) & (!g3063) & (g3065)) + ((g2) & (!g8) & (g3063) & (!g3065)) + ((g2) & (g8) & (!g3063) & (!g3065)));
	assign g3185 = (((!g3062) & (!g3060) & (!g3069) & (g3184)) + ((!g3062) & (g3060) & (!g3069) & (g3184)) + ((!g3062) & (g3060) & (g3069) & (g3184)) + ((g3062) & (!g3060) & (!g3069) & (!g3184)) + ((g3062) & (!g3060) & (g3069) & (!g3184)) + ((g3062) & (!g3060) & (g3069) & (g3184)) + ((g3062) & (g3060) & (!g3069) & (!g3184)) + ((g3062) & (g3060) & (g3069) & (!g3184)));
	assign g3186 = (((!g4) & (!g2) & (!g3180) & (!g3183) & (g3185)) + ((!g4) & (!g2) & (!g3180) & (g3183) & (g3185)) + ((!g4) & (!g2) & (g3180) & (!g3183) & (g3185)) + ((!g4) & (!g2) & (g3180) & (g3183) & (!g3185)) + ((!g4) & (!g2) & (g3180) & (g3183) & (g3185)) + ((!g4) & (g2) & (!g3180) & (!g3183) & (g3185)) + ((!g4) & (g2) & (!g3180) & (g3183) & (!g3185)) + ((!g4) & (g2) & (!g3180) & (g3183) & (g3185)) + ((!g4) & (g2) & (g3180) & (!g3183) & (!g3185)) + ((!g4) & (g2) & (g3180) & (!g3183) & (g3185)) + ((!g4) & (g2) & (g3180) & (g3183) & (!g3185)) + ((!g4) & (g2) & (g3180) & (g3183) & (g3185)) + ((g4) & (!g2) & (g3180) & (g3183) & (g3185)) + ((g4) & (g2) & (!g3180) & (g3183) & (g3185)) + ((g4) & (g2) & (g3180) & (!g3183) & (g3185)) + ((g4) & (g2) & (g3180) & (g3183) & (g3185)));
	assign g3187 = (((!g1) & (!g3061) & (!g3177) & (g3178) & (!g3179) & (!g3186)) + ((!g1) & (!g3061) & (g3177) & (!g3178) & (!g3179) & (!g3186)) + ((!g1) & (!g3061) & (g3177) & (g3178) & (!g3179) & (!g3186)) + ((!g1) & (g3061) & (!g3177) & (!g3178) & (!g3179) & (!g3186)) + ((!g1) & (g3061) & (!g3177) & (g3178) & (!g3179) & (!g3186)) + ((g1) & (!g3061) & (!g3177) & (!g3178) & (!g3179) & (!g3186)) + ((g1) & (!g3061) & (!g3177) & (!g3178) & (!g3179) & (g3186)) + ((g1) & (!g3061) & (!g3177) & (!g3178) & (g3179) & (!g3186)) + ((g1) & (!g3061) & (!g3177) & (g3178) & (!g3179) & (!g3186)) + ((g1) & (!g3061) & (!g3177) & (g3178) & (!g3179) & (g3186)) + ((g1) & (!g3061) & (!g3177) & (g3178) & (g3179) & (!g3186)) + ((g1) & (!g3061) & (g3177) & (g3178) & (!g3179) & (!g3186)) + ((g1) & (!g3061) & (g3177) & (g3178) & (!g3179) & (g3186)) + ((g1) & (!g3061) & (g3177) & (g3178) & (g3179) & (!g3186)) + ((g1) & (g3061) & (g3177) & (!g3178) & (!g3179) & (!g3186)) + ((g1) & (g3061) & (g3177) & (!g3178) & (!g3179) & (g3186)) + ((g1) & (g3061) & (g3177) & (!g3178) & (g3179) & (!g3186)) + ((g1) & (g3061) & (g3177) & (g3178) & (!g3179) & (!g3186)) + ((g1) & (g3061) & (g3177) & (g3178) & (!g3179) & (g3186)) + ((g1) & (g3061) & (g3177) & (g3178) & (g3179) & (!g3186)));
	assign g3188 = (((!g18) & (!g3070) & (g3176) & (!g3187)) + ((!g18) & (g3070) & (!g3176) & (!g3187)) + ((!g18) & (g3070) & (!g3176) & (g3187)) + ((!g18) & (g3070) & (g3176) & (g3187)) + ((g18) & (!g3070) & (!g3176) & (!g3187)) + ((g18) & (g3070) & (!g3176) & (g3187)) + ((g18) & (g3070) & (g3176) & (!g3187)) + ((g18) & (g3070) & (g3176) & (g3187)));
	assign g3189 = (((!g27) & (!g39) & (!g3072) & (g3073) & (g3175) & (!g3187)) + ((!g27) & (!g39) & (g3072) & (!g3073) & (!g3175) & (!g3187)) + ((!g27) & (!g39) & (g3072) & (!g3073) & (!g3175) & (g3187)) + ((!g27) & (!g39) & (g3072) & (!g3073) & (g3175) & (!g3187)) + ((!g27) & (!g39) & (g3072) & (!g3073) & (g3175) & (g3187)) + ((!g27) & (!g39) & (g3072) & (g3073) & (!g3175) & (!g3187)) + ((!g27) & (!g39) & (g3072) & (g3073) & (!g3175) & (g3187)) + ((!g27) & (!g39) & (g3072) & (g3073) & (g3175) & (g3187)) + ((!g27) & (g39) & (!g3072) & (!g3073) & (g3175) & (!g3187)) + ((!g27) & (g39) & (!g3072) & (g3073) & (!g3175) & (!g3187)) + ((!g27) & (g39) & (!g3072) & (g3073) & (g3175) & (!g3187)) + ((!g27) & (g39) & (g3072) & (!g3073) & (!g3175) & (!g3187)) + ((!g27) & (g39) & (g3072) & (!g3073) & (!g3175) & (g3187)) + ((!g27) & (g39) & (g3072) & (!g3073) & (g3175) & (g3187)) + ((!g27) & (g39) & (g3072) & (g3073) & (!g3175) & (g3187)) + ((!g27) & (g39) & (g3072) & (g3073) & (g3175) & (g3187)) + ((g27) & (!g39) & (!g3072) & (!g3073) & (!g3175) & (!g3187)) + ((g27) & (!g39) & (!g3072) & (!g3073) & (g3175) & (!g3187)) + ((g27) & (!g39) & (!g3072) & (g3073) & (!g3175) & (!g3187)) + ((g27) & (!g39) & (g3072) & (!g3073) & (!g3175) & (g3187)) + ((g27) & (!g39) & (g3072) & (!g3073) & (g3175) & (g3187)) + ((g27) & (!g39) & (g3072) & (g3073) & (!g3175) & (g3187)) + ((g27) & (!g39) & (g3072) & (g3073) & (g3175) & (!g3187)) + ((g27) & (!g39) & (g3072) & (g3073) & (g3175) & (g3187)) + ((g27) & (g39) & (!g3072) & (!g3073) & (!g3175) & (!g3187)) + ((g27) & (g39) & (g3072) & (!g3073) & (!g3175) & (g3187)) + ((g27) & (g39) & (g3072) & (!g3073) & (g3175) & (!g3187)) + ((g27) & (g39) & (g3072) & (!g3073) & (g3175) & (g3187)) + ((g27) & (g39) & (g3072) & (g3073) & (!g3175) & (!g3187)) + ((g27) & (g39) & (g3072) & (g3073) & (!g3175) & (g3187)) + ((g27) & (g39) & (g3072) & (g3073) & (g3175) & (!g3187)) + ((g27) & (g39) & (g3072) & (g3073) & (g3175) & (g3187)));
	assign g3190 = (((!g39) & (!g3073) & (g3175) & (!g3187)) + ((!g39) & (g3073) & (!g3175) & (!g3187)) + ((!g39) & (g3073) & (!g3175) & (g3187)) + ((!g39) & (g3073) & (g3175) & (g3187)) + ((g39) & (!g3073) & (!g3175) & (!g3187)) + ((g39) & (g3073) & (!g3175) & (g3187)) + ((g39) & (g3073) & (g3175) & (!g3187)) + ((g39) & (g3073) & (g3175) & (g3187)));
	assign g3191 = (((!g54) & (!g68) & (!g3075) & (g3076) & (g3174) & (!g3187)) + ((!g54) & (!g68) & (g3075) & (!g3076) & (!g3174) & (!g3187)) + ((!g54) & (!g68) & (g3075) & (!g3076) & (!g3174) & (g3187)) + ((!g54) & (!g68) & (g3075) & (!g3076) & (g3174) & (!g3187)) + ((!g54) & (!g68) & (g3075) & (!g3076) & (g3174) & (g3187)) + ((!g54) & (!g68) & (g3075) & (g3076) & (!g3174) & (!g3187)) + ((!g54) & (!g68) & (g3075) & (g3076) & (!g3174) & (g3187)) + ((!g54) & (!g68) & (g3075) & (g3076) & (g3174) & (g3187)) + ((!g54) & (g68) & (!g3075) & (!g3076) & (g3174) & (!g3187)) + ((!g54) & (g68) & (!g3075) & (g3076) & (!g3174) & (!g3187)) + ((!g54) & (g68) & (!g3075) & (g3076) & (g3174) & (!g3187)) + ((!g54) & (g68) & (g3075) & (!g3076) & (!g3174) & (!g3187)) + ((!g54) & (g68) & (g3075) & (!g3076) & (!g3174) & (g3187)) + ((!g54) & (g68) & (g3075) & (!g3076) & (g3174) & (g3187)) + ((!g54) & (g68) & (g3075) & (g3076) & (!g3174) & (g3187)) + ((!g54) & (g68) & (g3075) & (g3076) & (g3174) & (g3187)) + ((g54) & (!g68) & (!g3075) & (!g3076) & (!g3174) & (!g3187)) + ((g54) & (!g68) & (!g3075) & (!g3076) & (g3174) & (!g3187)) + ((g54) & (!g68) & (!g3075) & (g3076) & (!g3174) & (!g3187)) + ((g54) & (!g68) & (g3075) & (!g3076) & (!g3174) & (g3187)) + ((g54) & (!g68) & (g3075) & (!g3076) & (g3174) & (g3187)) + ((g54) & (!g68) & (g3075) & (g3076) & (!g3174) & (g3187)) + ((g54) & (!g68) & (g3075) & (g3076) & (g3174) & (!g3187)) + ((g54) & (!g68) & (g3075) & (g3076) & (g3174) & (g3187)) + ((g54) & (g68) & (!g3075) & (!g3076) & (!g3174) & (!g3187)) + ((g54) & (g68) & (g3075) & (!g3076) & (!g3174) & (g3187)) + ((g54) & (g68) & (g3075) & (!g3076) & (g3174) & (!g3187)) + ((g54) & (g68) & (g3075) & (!g3076) & (g3174) & (g3187)) + ((g54) & (g68) & (g3075) & (g3076) & (!g3174) & (!g3187)) + ((g54) & (g68) & (g3075) & (g3076) & (!g3174) & (g3187)) + ((g54) & (g68) & (g3075) & (g3076) & (g3174) & (!g3187)) + ((g54) & (g68) & (g3075) & (g3076) & (g3174) & (g3187)));
	assign g3192 = (((!g68) & (!g3076) & (g3174) & (!g3187)) + ((!g68) & (g3076) & (!g3174) & (!g3187)) + ((!g68) & (g3076) & (!g3174) & (g3187)) + ((!g68) & (g3076) & (g3174) & (g3187)) + ((g68) & (!g3076) & (!g3174) & (!g3187)) + ((g68) & (g3076) & (!g3174) & (g3187)) + ((g68) & (g3076) & (g3174) & (!g3187)) + ((g68) & (g3076) & (g3174) & (g3187)));
	assign g3193 = (((!g87) & (!g104) & (!g3078) & (g3079) & (g3173) & (!g3187)) + ((!g87) & (!g104) & (g3078) & (!g3079) & (!g3173) & (!g3187)) + ((!g87) & (!g104) & (g3078) & (!g3079) & (!g3173) & (g3187)) + ((!g87) & (!g104) & (g3078) & (!g3079) & (g3173) & (!g3187)) + ((!g87) & (!g104) & (g3078) & (!g3079) & (g3173) & (g3187)) + ((!g87) & (!g104) & (g3078) & (g3079) & (!g3173) & (!g3187)) + ((!g87) & (!g104) & (g3078) & (g3079) & (!g3173) & (g3187)) + ((!g87) & (!g104) & (g3078) & (g3079) & (g3173) & (g3187)) + ((!g87) & (g104) & (!g3078) & (!g3079) & (g3173) & (!g3187)) + ((!g87) & (g104) & (!g3078) & (g3079) & (!g3173) & (!g3187)) + ((!g87) & (g104) & (!g3078) & (g3079) & (g3173) & (!g3187)) + ((!g87) & (g104) & (g3078) & (!g3079) & (!g3173) & (!g3187)) + ((!g87) & (g104) & (g3078) & (!g3079) & (!g3173) & (g3187)) + ((!g87) & (g104) & (g3078) & (!g3079) & (g3173) & (g3187)) + ((!g87) & (g104) & (g3078) & (g3079) & (!g3173) & (g3187)) + ((!g87) & (g104) & (g3078) & (g3079) & (g3173) & (g3187)) + ((g87) & (!g104) & (!g3078) & (!g3079) & (!g3173) & (!g3187)) + ((g87) & (!g104) & (!g3078) & (!g3079) & (g3173) & (!g3187)) + ((g87) & (!g104) & (!g3078) & (g3079) & (!g3173) & (!g3187)) + ((g87) & (!g104) & (g3078) & (!g3079) & (!g3173) & (g3187)) + ((g87) & (!g104) & (g3078) & (!g3079) & (g3173) & (g3187)) + ((g87) & (!g104) & (g3078) & (g3079) & (!g3173) & (g3187)) + ((g87) & (!g104) & (g3078) & (g3079) & (g3173) & (!g3187)) + ((g87) & (!g104) & (g3078) & (g3079) & (g3173) & (g3187)) + ((g87) & (g104) & (!g3078) & (!g3079) & (!g3173) & (!g3187)) + ((g87) & (g104) & (g3078) & (!g3079) & (!g3173) & (g3187)) + ((g87) & (g104) & (g3078) & (!g3079) & (g3173) & (!g3187)) + ((g87) & (g104) & (g3078) & (!g3079) & (g3173) & (g3187)) + ((g87) & (g104) & (g3078) & (g3079) & (!g3173) & (!g3187)) + ((g87) & (g104) & (g3078) & (g3079) & (!g3173) & (g3187)) + ((g87) & (g104) & (g3078) & (g3079) & (g3173) & (!g3187)) + ((g87) & (g104) & (g3078) & (g3079) & (g3173) & (g3187)));
	assign g3194 = (((!g104) & (!g3079) & (g3173) & (!g3187)) + ((!g104) & (g3079) & (!g3173) & (!g3187)) + ((!g104) & (g3079) & (!g3173) & (g3187)) + ((!g104) & (g3079) & (g3173) & (g3187)) + ((g104) & (!g3079) & (!g3173) & (!g3187)) + ((g104) & (g3079) & (!g3173) & (g3187)) + ((g104) & (g3079) & (g3173) & (!g3187)) + ((g104) & (g3079) & (g3173) & (g3187)));
	assign g3195 = (((!g127) & (!g147) & (!g3081) & (g3082) & (g3172) & (!g3187)) + ((!g127) & (!g147) & (g3081) & (!g3082) & (!g3172) & (!g3187)) + ((!g127) & (!g147) & (g3081) & (!g3082) & (!g3172) & (g3187)) + ((!g127) & (!g147) & (g3081) & (!g3082) & (g3172) & (!g3187)) + ((!g127) & (!g147) & (g3081) & (!g3082) & (g3172) & (g3187)) + ((!g127) & (!g147) & (g3081) & (g3082) & (!g3172) & (!g3187)) + ((!g127) & (!g147) & (g3081) & (g3082) & (!g3172) & (g3187)) + ((!g127) & (!g147) & (g3081) & (g3082) & (g3172) & (g3187)) + ((!g127) & (g147) & (!g3081) & (!g3082) & (g3172) & (!g3187)) + ((!g127) & (g147) & (!g3081) & (g3082) & (!g3172) & (!g3187)) + ((!g127) & (g147) & (!g3081) & (g3082) & (g3172) & (!g3187)) + ((!g127) & (g147) & (g3081) & (!g3082) & (!g3172) & (!g3187)) + ((!g127) & (g147) & (g3081) & (!g3082) & (!g3172) & (g3187)) + ((!g127) & (g147) & (g3081) & (!g3082) & (g3172) & (g3187)) + ((!g127) & (g147) & (g3081) & (g3082) & (!g3172) & (g3187)) + ((!g127) & (g147) & (g3081) & (g3082) & (g3172) & (g3187)) + ((g127) & (!g147) & (!g3081) & (!g3082) & (!g3172) & (!g3187)) + ((g127) & (!g147) & (!g3081) & (!g3082) & (g3172) & (!g3187)) + ((g127) & (!g147) & (!g3081) & (g3082) & (!g3172) & (!g3187)) + ((g127) & (!g147) & (g3081) & (!g3082) & (!g3172) & (g3187)) + ((g127) & (!g147) & (g3081) & (!g3082) & (g3172) & (g3187)) + ((g127) & (!g147) & (g3081) & (g3082) & (!g3172) & (g3187)) + ((g127) & (!g147) & (g3081) & (g3082) & (g3172) & (!g3187)) + ((g127) & (!g147) & (g3081) & (g3082) & (g3172) & (g3187)) + ((g127) & (g147) & (!g3081) & (!g3082) & (!g3172) & (!g3187)) + ((g127) & (g147) & (g3081) & (!g3082) & (!g3172) & (g3187)) + ((g127) & (g147) & (g3081) & (!g3082) & (g3172) & (!g3187)) + ((g127) & (g147) & (g3081) & (!g3082) & (g3172) & (g3187)) + ((g127) & (g147) & (g3081) & (g3082) & (!g3172) & (!g3187)) + ((g127) & (g147) & (g3081) & (g3082) & (!g3172) & (g3187)) + ((g127) & (g147) & (g3081) & (g3082) & (g3172) & (!g3187)) + ((g127) & (g147) & (g3081) & (g3082) & (g3172) & (g3187)));
	assign g3196 = (((!g147) & (!g3082) & (g3172) & (!g3187)) + ((!g147) & (g3082) & (!g3172) & (!g3187)) + ((!g147) & (g3082) & (!g3172) & (g3187)) + ((!g147) & (g3082) & (g3172) & (g3187)) + ((g147) & (!g3082) & (!g3172) & (!g3187)) + ((g147) & (g3082) & (!g3172) & (g3187)) + ((g147) & (g3082) & (g3172) & (!g3187)) + ((g147) & (g3082) & (g3172) & (g3187)));
	assign g3197 = (((!g174) & (!g198) & (!g3084) & (g3085) & (g3171) & (!g3187)) + ((!g174) & (!g198) & (g3084) & (!g3085) & (!g3171) & (!g3187)) + ((!g174) & (!g198) & (g3084) & (!g3085) & (!g3171) & (g3187)) + ((!g174) & (!g198) & (g3084) & (!g3085) & (g3171) & (!g3187)) + ((!g174) & (!g198) & (g3084) & (!g3085) & (g3171) & (g3187)) + ((!g174) & (!g198) & (g3084) & (g3085) & (!g3171) & (!g3187)) + ((!g174) & (!g198) & (g3084) & (g3085) & (!g3171) & (g3187)) + ((!g174) & (!g198) & (g3084) & (g3085) & (g3171) & (g3187)) + ((!g174) & (g198) & (!g3084) & (!g3085) & (g3171) & (!g3187)) + ((!g174) & (g198) & (!g3084) & (g3085) & (!g3171) & (!g3187)) + ((!g174) & (g198) & (!g3084) & (g3085) & (g3171) & (!g3187)) + ((!g174) & (g198) & (g3084) & (!g3085) & (!g3171) & (!g3187)) + ((!g174) & (g198) & (g3084) & (!g3085) & (!g3171) & (g3187)) + ((!g174) & (g198) & (g3084) & (!g3085) & (g3171) & (g3187)) + ((!g174) & (g198) & (g3084) & (g3085) & (!g3171) & (g3187)) + ((!g174) & (g198) & (g3084) & (g3085) & (g3171) & (g3187)) + ((g174) & (!g198) & (!g3084) & (!g3085) & (!g3171) & (!g3187)) + ((g174) & (!g198) & (!g3084) & (!g3085) & (g3171) & (!g3187)) + ((g174) & (!g198) & (!g3084) & (g3085) & (!g3171) & (!g3187)) + ((g174) & (!g198) & (g3084) & (!g3085) & (!g3171) & (g3187)) + ((g174) & (!g198) & (g3084) & (!g3085) & (g3171) & (g3187)) + ((g174) & (!g198) & (g3084) & (g3085) & (!g3171) & (g3187)) + ((g174) & (!g198) & (g3084) & (g3085) & (g3171) & (!g3187)) + ((g174) & (!g198) & (g3084) & (g3085) & (g3171) & (g3187)) + ((g174) & (g198) & (!g3084) & (!g3085) & (!g3171) & (!g3187)) + ((g174) & (g198) & (g3084) & (!g3085) & (!g3171) & (g3187)) + ((g174) & (g198) & (g3084) & (!g3085) & (g3171) & (!g3187)) + ((g174) & (g198) & (g3084) & (!g3085) & (g3171) & (g3187)) + ((g174) & (g198) & (g3084) & (g3085) & (!g3171) & (!g3187)) + ((g174) & (g198) & (g3084) & (g3085) & (!g3171) & (g3187)) + ((g174) & (g198) & (g3084) & (g3085) & (g3171) & (!g3187)) + ((g174) & (g198) & (g3084) & (g3085) & (g3171) & (g3187)));
	assign g3198 = (((!g198) & (!g3085) & (g3171) & (!g3187)) + ((!g198) & (g3085) & (!g3171) & (!g3187)) + ((!g198) & (g3085) & (!g3171) & (g3187)) + ((!g198) & (g3085) & (g3171) & (g3187)) + ((g198) & (!g3085) & (!g3171) & (!g3187)) + ((g198) & (g3085) & (!g3171) & (g3187)) + ((g198) & (g3085) & (g3171) & (!g3187)) + ((g198) & (g3085) & (g3171) & (g3187)));
	assign g3199 = (((!g229) & (!g255) & (!g3087) & (g3088) & (g3170) & (!g3187)) + ((!g229) & (!g255) & (g3087) & (!g3088) & (!g3170) & (!g3187)) + ((!g229) & (!g255) & (g3087) & (!g3088) & (!g3170) & (g3187)) + ((!g229) & (!g255) & (g3087) & (!g3088) & (g3170) & (!g3187)) + ((!g229) & (!g255) & (g3087) & (!g3088) & (g3170) & (g3187)) + ((!g229) & (!g255) & (g3087) & (g3088) & (!g3170) & (!g3187)) + ((!g229) & (!g255) & (g3087) & (g3088) & (!g3170) & (g3187)) + ((!g229) & (!g255) & (g3087) & (g3088) & (g3170) & (g3187)) + ((!g229) & (g255) & (!g3087) & (!g3088) & (g3170) & (!g3187)) + ((!g229) & (g255) & (!g3087) & (g3088) & (!g3170) & (!g3187)) + ((!g229) & (g255) & (!g3087) & (g3088) & (g3170) & (!g3187)) + ((!g229) & (g255) & (g3087) & (!g3088) & (!g3170) & (!g3187)) + ((!g229) & (g255) & (g3087) & (!g3088) & (!g3170) & (g3187)) + ((!g229) & (g255) & (g3087) & (!g3088) & (g3170) & (g3187)) + ((!g229) & (g255) & (g3087) & (g3088) & (!g3170) & (g3187)) + ((!g229) & (g255) & (g3087) & (g3088) & (g3170) & (g3187)) + ((g229) & (!g255) & (!g3087) & (!g3088) & (!g3170) & (!g3187)) + ((g229) & (!g255) & (!g3087) & (!g3088) & (g3170) & (!g3187)) + ((g229) & (!g255) & (!g3087) & (g3088) & (!g3170) & (!g3187)) + ((g229) & (!g255) & (g3087) & (!g3088) & (!g3170) & (g3187)) + ((g229) & (!g255) & (g3087) & (!g3088) & (g3170) & (g3187)) + ((g229) & (!g255) & (g3087) & (g3088) & (!g3170) & (g3187)) + ((g229) & (!g255) & (g3087) & (g3088) & (g3170) & (!g3187)) + ((g229) & (!g255) & (g3087) & (g3088) & (g3170) & (g3187)) + ((g229) & (g255) & (!g3087) & (!g3088) & (!g3170) & (!g3187)) + ((g229) & (g255) & (g3087) & (!g3088) & (!g3170) & (g3187)) + ((g229) & (g255) & (g3087) & (!g3088) & (g3170) & (!g3187)) + ((g229) & (g255) & (g3087) & (!g3088) & (g3170) & (g3187)) + ((g229) & (g255) & (g3087) & (g3088) & (!g3170) & (!g3187)) + ((g229) & (g255) & (g3087) & (g3088) & (!g3170) & (g3187)) + ((g229) & (g255) & (g3087) & (g3088) & (g3170) & (!g3187)) + ((g229) & (g255) & (g3087) & (g3088) & (g3170) & (g3187)));
	assign g3200 = (((!g255) & (!g3088) & (g3170) & (!g3187)) + ((!g255) & (g3088) & (!g3170) & (!g3187)) + ((!g255) & (g3088) & (!g3170) & (g3187)) + ((!g255) & (g3088) & (g3170) & (g3187)) + ((g255) & (!g3088) & (!g3170) & (!g3187)) + ((g255) & (g3088) & (!g3170) & (g3187)) + ((g255) & (g3088) & (g3170) & (!g3187)) + ((g255) & (g3088) & (g3170) & (g3187)));
	assign g3201 = (((!g290) & (!g319) & (!g3090) & (g3091) & (g3169) & (!g3187)) + ((!g290) & (!g319) & (g3090) & (!g3091) & (!g3169) & (!g3187)) + ((!g290) & (!g319) & (g3090) & (!g3091) & (!g3169) & (g3187)) + ((!g290) & (!g319) & (g3090) & (!g3091) & (g3169) & (!g3187)) + ((!g290) & (!g319) & (g3090) & (!g3091) & (g3169) & (g3187)) + ((!g290) & (!g319) & (g3090) & (g3091) & (!g3169) & (!g3187)) + ((!g290) & (!g319) & (g3090) & (g3091) & (!g3169) & (g3187)) + ((!g290) & (!g319) & (g3090) & (g3091) & (g3169) & (g3187)) + ((!g290) & (g319) & (!g3090) & (!g3091) & (g3169) & (!g3187)) + ((!g290) & (g319) & (!g3090) & (g3091) & (!g3169) & (!g3187)) + ((!g290) & (g319) & (!g3090) & (g3091) & (g3169) & (!g3187)) + ((!g290) & (g319) & (g3090) & (!g3091) & (!g3169) & (!g3187)) + ((!g290) & (g319) & (g3090) & (!g3091) & (!g3169) & (g3187)) + ((!g290) & (g319) & (g3090) & (!g3091) & (g3169) & (g3187)) + ((!g290) & (g319) & (g3090) & (g3091) & (!g3169) & (g3187)) + ((!g290) & (g319) & (g3090) & (g3091) & (g3169) & (g3187)) + ((g290) & (!g319) & (!g3090) & (!g3091) & (!g3169) & (!g3187)) + ((g290) & (!g319) & (!g3090) & (!g3091) & (g3169) & (!g3187)) + ((g290) & (!g319) & (!g3090) & (g3091) & (!g3169) & (!g3187)) + ((g290) & (!g319) & (g3090) & (!g3091) & (!g3169) & (g3187)) + ((g290) & (!g319) & (g3090) & (!g3091) & (g3169) & (g3187)) + ((g290) & (!g319) & (g3090) & (g3091) & (!g3169) & (g3187)) + ((g290) & (!g319) & (g3090) & (g3091) & (g3169) & (!g3187)) + ((g290) & (!g319) & (g3090) & (g3091) & (g3169) & (g3187)) + ((g290) & (g319) & (!g3090) & (!g3091) & (!g3169) & (!g3187)) + ((g290) & (g319) & (g3090) & (!g3091) & (!g3169) & (g3187)) + ((g290) & (g319) & (g3090) & (!g3091) & (g3169) & (!g3187)) + ((g290) & (g319) & (g3090) & (!g3091) & (g3169) & (g3187)) + ((g290) & (g319) & (g3090) & (g3091) & (!g3169) & (!g3187)) + ((g290) & (g319) & (g3090) & (g3091) & (!g3169) & (g3187)) + ((g290) & (g319) & (g3090) & (g3091) & (g3169) & (!g3187)) + ((g290) & (g319) & (g3090) & (g3091) & (g3169) & (g3187)));
	assign g3202 = (((!g319) & (!g3091) & (g3169) & (!g3187)) + ((!g319) & (g3091) & (!g3169) & (!g3187)) + ((!g319) & (g3091) & (!g3169) & (g3187)) + ((!g319) & (g3091) & (g3169) & (g3187)) + ((g319) & (!g3091) & (!g3169) & (!g3187)) + ((g319) & (g3091) & (!g3169) & (g3187)) + ((g319) & (g3091) & (g3169) & (!g3187)) + ((g319) & (g3091) & (g3169) & (g3187)));
	assign g3203 = (((!g358) & (!g390) & (!g3093) & (g3094) & (g3168) & (!g3187)) + ((!g358) & (!g390) & (g3093) & (!g3094) & (!g3168) & (!g3187)) + ((!g358) & (!g390) & (g3093) & (!g3094) & (!g3168) & (g3187)) + ((!g358) & (!g390) & (g3093) & (!g3094) & (g3168) & (!g3187)) + ((!g358) & (!g390) & (g3093) & (!g3094) & (g3168) & (g3187)) + ((!g358) & (!g390) & (g3093) & (g3094) & (!g3168) & (!g3187)) + ((!g358) & (!g390) & (g3093) & (g3094) & (!g3168) & (g3187)) + ((!g358) & (!g390) & (g3093) & (g3094) & (g3168) & (g3187)) + ((!g358) & (g390) & (!g3093) & (!g3094) & (g3168) & (!g3187)) + ((!g358) & (g390) & (!g3093) & (g3094) & (!g3168) & (!g3187)) + ((!g358) & (g390) & (!g3093) & (g3094) & (g3168) & (!g3187)) + ((!g358) & (g390) & (g3093) & (!g3094) & (!g3168) & (!g3187)) + ((!g358) & (g390) & (g3093) & (!g3094) & (!g3168) & (g3187)) + ((!g358) & (g390) & (g3093) & (!g3094) & (g3168) & (g3187)) + ((!g358) & (g390) & (g3093) & (g3094) & (!g3168) & (g3187)) + ((!g358) & (g390) & (g3093) & (g3094) & (g3168) & (g3187)) + ((g358) & (!g390) & (!g3093) & (!g3094) & (!g3168) & (!g3187)) + ((g358) & (!g390) & (!g3093) & (!g3094) & (g3168) & (!g3187)) + ((g358) & (!g390) & (!g3093) & (g3094) & (!g3168) & (!g3187)) + ((g358) & (!g390) & (g3093) & (!g3094) & (!g3168) & (g3187)) + ((g358) & (!g390) & (g3093) & (!g3094) & (g3168) & (g3187)) + ((g358) & (!g390) & (g3093) & (g3094) & (!g3168) & (g3187)) + ((g358) & (!g390) & (g3093) & (g3094) & (g3168) & (!g3187)) + ((g358) & (!g390) & (g3093) & (g3094) & (g3168) & (g3187)) + ((g358) & (g390) & (!g3093) & (!g3094) & (!g3168) & (!g3187)) + ((g358) & (g390) & (g3093) & (!g3094) & (!g3168) & (g3187)) + ((g358) & (g390) & (g3093) & (!g3094) & (g3168) & (!g3187)) + ((g358) & (g390) & (g3093) & (!g3094) & (g3168) & (g3187)) + ((g358) & (g390) & (g3093) & (g3094) & (!g3168) & (!g3187)) + ((g358) & (g390) & (g3093) & (g3094) & (!g3168) & (g3187)) + ((g358) & (g390) & (g3093) & (g3094) & (g3168) & (!g3187)) + ((g358) & (g390) & (g3093) & (g3094) & (g3168) & (g3187)));
	assign g3204 = (((!g390) & (!g3094) & (g3168) & (!g3187)) + ((!g390) & (g3094) & (!g3168) & (!g3187)) + ((!g390) & (g3094) & (!g3168) & (g3187)) + ((!g390) & (g3094) & (g3168) & (g3187)) + ((g390) & (!g3094) & (!g3168) & (!g3187)) + ((g390) & (g3094) & (!g3168) & (g3187)) + ((g390) & (g3094) & (g3168) & (!g3187)) + ((g390) & (g3094) & (g3168) & (g3187)));
	assign g3205 = (((!g433) & (!g468) & (!g3096) & (g3097) & (g3167) & (!g3187)) + ((!g433) & (!g468) & (g3096) & (!g3097) & (!g3167) & (!g3187)) + ((!g433) & (!g468) & (g3096) & (!g3097) & (!g3167) & (g3187)) + ((!g433) & (!g468) & (g3096) & (!g3097) & (g3167) & (!g3187)) + ((!g433) & (!g468) & (g3096) & (!g3097) & (g3167) & (g3187)) + ((!g433) & (!g468) & (g3096) & (g3097) & (!g3167) & (!g3187)) + ((!g433) & (!g468) & (g3096) & (g3097) & (!g3167) & (g3187)) + ((!g433) & (!g468) & (g3096) & (g3097) & (g3167) & (g3187)) + ((!g433) & (g468) & (!g3096) & (!g3097) & (g3167) & (!g3187)) + ((!g433) & (g468) & (!g3096) & (g3097) & (!g3167) & (!g3187)) + ((!g433) & (g468) & (!g3096) & (g3097) & (g3167) & (!g3187)) + ((!g433) & (g468) & (g3096) & (!g3097) & (!g3167) & (!g3187)) + ((!g433) & (g468) & (g3096) & (!g3097) & (!g3167) & (g3187)) + ((!g433) & (g468) & (g3096) & (!g3097) & (g3167) & (g3187)) + ((!g433) & (g468) & (g3096) & (g3097) & (!g3167) & (g3187)) + ((!g433) & (g468) & (g3096) & (g3097) & (g3167) & (g3187)) + ((g433) & (!g468) & (!g3096) & (!g3097) & (!g3167) & (!g3187)) + ((g433) & (!g468) & (!g3096) & (!g3097) & (g3167) & (!g3187)) + ((g433) & (!g468) & (!g3096) & (g3097) & (!g3167) & (!g3187)) + ((g433) & (!g468) & (g3096) & (!g3097) & (!g3167) & (g3187)) + ((g433) & (!g468) & (g3096) & (!g3097) & (g3167) & (g3187)) + ((g433) & (!g468) & (g3096) & (g3097) & (!g3167) & (g3187)) + ((g433) & (!g468) & (g3096) & (g3097) & (g3167) & (!g3187)) + ((g433) & (!g468) & (g3096) & (g3097) & (g3167) & (g3187)) + ((g433) & (g468) & (!g3096) & (!g3097) & (!g3167) & (!g3187)) + ((g433) & (g468) & (g3096) & (!g3097) & (!g3167) & (g3187)) + ((g433) & (g468) & (g3096) & (!g3097) & (g3167) & (!g3187)) + ((g433) & (g468) & (g3096) & (!g3097) & (g3167) & (g3187)) + ((g433) & (g468) & (g3096) & (g3097) & (!g3167) & (!g3187)) + ((g433) & (g468) & (g3096) & (g3097) & (!g3167) & (g3187)) + ((g433) & (g468) & (g3096) & (g3097) & (g3167) & (!g3187)) + ((g433) & (g468) & (g3096) & (g3097) & (g3167) & (g3187)));
	assign g3206 = (((!g468) & (!g3097) & (g3167) & (!g3187)) + ((!g468) & (g3097) & (!g3167) & (!g3187)) + ((!g468) & (g3097) & (!g3167) & (g3187)) + ((!g468) & (g3097) & (g3167) & (g3187)) + ((g468) & (!g3097) & (!g3167) & (!g3187)) + ((g468) & (g3097) & (!g3167) & (g3187)) + ((g468) & (g3097) & (g3167) & (!g3187)) + ((g468) & (g3097) & (g3167) & (g3187)));
	assign g3207 = (((!g515) & (!g553) & (!g3099) & (g3100) & (g3166) & (!g3187)) + ((!g515) & (!g553) & (g3099) & (!g3100) & (!g3166) & (!g3187)) + ((!g515) & (!g553) & (g3099) & (!g3100) & (!g3166) & (g3187)) + ((!g515) & (!g553) & (g3099) & (!g3100) & (g3166) & (!g3187)) + ((!g515) & (!g553) & (g3099) & (!g3100) & (g3166) & (g3187)) + ((!g515) & (!g553) & (g3099) & (g3100) & (!g3166) & (!g3187)) + ((!g515) & (!g553) & (g3099) & (g3100) & (!g3166) & (g3187)) + ((!g515) & (!g553) & (g3099) & (g3100) & (g3166) & (g3187)) + ((!g515) & (g553) & (!g3099) & (!g3100) & (g3166) & (!g3187)) + ((!g515) & (g553) & (!g3099) & (g3100) & (!g3166) & (!g3187)) + ((!g515) & (g553) & (!g3099) & (g3100) & (g3166) & (!g3187)) + ((!g515) & (g553) & (g3099) & (!g3100) & (!g3166) & (!g3187)) + ((!g515) & (g553) & (g3099) & (!g3100) & (!g3166) & (g3187)) + ((!g515) & (g553) & (g3099) & (!g3100) & (g3166) & (g3187)) + ((!g515) & (g553) & (g3099) & (g3100) & (!g3166) & (g3187)) + ((!g515) & (g553) & (g3099) & (g3100) & (g3166) & (g3187)) + ((g515) & (!g553) & (!g3099) & (!g3100) & (!g3166) & (!g3187)) + ((g515) & (!g553) & (!g3099) & (!g3100) & (g3166) & (!g3187)) + ((g515) & (!g553) & (!g3099) & (g3100) & (!g3166) & (!g3187)) + ((g515) & (!g553) & (g3099) & (!g3100) & (!g3166) & (g3187)) + ((g515) & (!g553) & (g3099) & (!g3100) & (g3166) & (g3187)) + ((g515) & (!g553) & (g3099) & (g3100) & (!g3166) & (g3187)) + ((g515) & (!g553) & (g3099) & (g3100) & (g3166) & (!g3187)) + ((g515) & (!g553) & (g3099) & (g3100) & (g3166) & (g3187)) + ((g515) & (g553) & (!g3099) & (!g3100) & (!g3166) & (!g3187)) + ((g515) & (g553) & (g3099) & (!g3100) & (!g3166) & (g3187)) + ((g515) & (g553) & (g3099) & (!g3100) & (g3166) & (!g3187)) + ((g515) & (g553) & (g3099) & (!g3100) & (g3166) & (g3187)) + ((g515) & (g553) & (g3099) & (g3100) & (!g3166) & (!g3187)) + ((g515) & (g553) & (g3099) & (g3100) & (!g3166) & (g3187)) + ((g515) & (g553) & (g3099) & (g3100) & (g3166) & (!g3187)) + ((g515) & (g553) & (g3099) & (g3100) & (g3166) & (g3187)));
	assign g3208 = (((!g553) & (!g3100) & (g3166) & (!g3187)) + ((!g553) & (g3100) & (!g3166) & (!g3187)) + ((!g553) & (g3100) & (!g3166) & (g3187)) + ((!g553) & (g3100) & (g3166) & (g3187)) + ((g553) & (!g3100) & (!g3166) & (!g3187)) + ((g553) & (g3100) & (!g3166) & (g3187)) + ((g553) & (g3100) & (g3166) & (!g3187)) + ((g553) & (g3100) & (g3166) & (g3187)));
	assign g3209 = (((!g604) & (!g645) & (!g3102) & (g3103) & (g3165) & (!g3187)) + ((!g604) & (!g645) & (g3102) & (!g3103) & (!g3165) & (!g3187)) + ((!g604) & (!g645) & (g3102) & (!g3103) & (!g3165) & (g3187)) + ((!g604) & (!g645) & (g3102) & (!g3103) & (g3165) & (!g3187)) + ((!g604) & (!g645) & (g3102) & (!g3103) & (g3165) & (g3187)) + ((!g604) & (!g645) & (g3102) & (g3103) & (!g3165) & (!g3187)) + ((!g604) & (!g645) & (g3102) & (g3103) & (!g3165) & (g3187)) + ((!g604) & (!g645) & (g3102) & (g3103) & (g3165) & (g3187)) + ((!g604) & (g645) & (!g3102) & (!g3103) & (g3165) & (!g3187)) + ((!g604) & (g645) & (!g3102) & (g3103) & (!g3165) & (!g3187)) + ((!g604) & (g645) & (!g3102) & (g3103) & (g3165) & (!g3187)) + ((!g604) & (g645) & (g3102) & (!g3103) & (!g3165) & (!g3187)) + ((!g604) & (g645) & (g3102) & (!g3103) & (!g3165) & (g3187)) + ((!g604) & (g645) & (g3102) & (!g3103) & (g3165) & (g3187)) + ((!g604) & (g645) & (g3102) & (g3103) & (!g3165) & (g3187)) + ((!g604) & (g645) & (g3102) & (g3103) & (g3165) & (g3187)) + ((g604) & (!g645) & (!g3102) & (!g3103) & (!g3165) & (!g3187)) + ((g604) & (!g645) & (!g3102) & (!g3103) & (g3165) & (!g3187)) + ((g604) & (!g645) & (!g3102) & (g3103) & (!g3165) & (!g3187)) + ((g604) & (!g645) & (g3102) & (!g3103) & (!g3165) & (g3187)) + ((g604) & (!g645) & (g3102) & (!g3103) & (g3165) & (g3187)) + ((g604) & (!g645) & (g3102) & (g3103) & (!g3165) & (g3187)) + ((g604) & (!g645) & (g3102) & (g3103) & (g3165) & (!g3187)) + ((g604) & (!g645) & (g3102) & (g3103) & (g3165) & (g3187)) + ((g604) & (g645) & (!g3102) & (!g3103) & (!g3165) & (!g3187)) + ((g604) & (g645) & (g3102) & (!g3103) & (!g3165) & (g3187)) + ((g604) & (g645) & (g3102) & (!g3103) & (g3165) & (!g3187)) + ((g604) & (g645) & (g3102) & (!g3103) & (g3165) & (g3187)) + ((g604) & (g645) & (g3102) & (g3103) & (!g3165) & (!g3187)) + ((g604) & (g645) & (g3102) & (g3103) & (!g3165) & (g3187)) + ((g604) & (g645) & (g3102) & (g3103) & (g3165) & (!g3187)) + ((g604) & (g645) & (g3102) & (g3103) & (g3165) & (g3187)));
	assign g3210 = (((!g645) & (!g3103) & (g3165) & (!g3187)) + ((!g645) & (g3103) & (!g3165) & (!g3187)) + ((!g645) & (g3103) & (!g3165) & (g3187)) + ((!g645) & (g3103) & (g3165) & (g3187)) + ((g645) & (!g3103) & (!g3165) & (!g3187)) + ((g645) & (g3103) & (!g3165) & (g3187)) + ((g645) & (g3103) & (g3165) & (!g3187)) + ((g645) & (g3103) & (g3165) & (g3187)));
	assign g3211 = (((!g700) & (!g744) & (!g3105) & (g3106) & (g3164) & (!g3187)) + ((!g700) & (!g744) & (g3105) & (!g3106) & (!g3164) & (!g3187)) + ((!g700) & (!g744) & (g3105) & (!g3106) & (!g3164) & (g3187)) + ((!g700) & (!g744) & (g3105) & (!g3106) & (g3164) & (!g3187)) + ((!g700) & (!g744) & (g3105) & (!g3106) & (g3164) & (g3187)) + ((!g700) & (!g744) & (g3105) & (g3106) & (!g3164) & (!g3187)) + ((!g700) & (!g744) & (g3105) & (g3106) & (!g3164) & (g3187)) + ((!g700) & (!g744) & (g3105) & (g3106) & (g3164) & (g3187)) + ((!g700) & (g744) & (!g3105) & (!g3106) & (g3164) & (!g3187)) + ((!g700) & (g744) & (!g3105) & (g3106) & (!g3164) & (!g3187)) + ((!g700) & (g744) & (!g3105) & (g3106) & (g3164) & (!g3187)) + ((!g700) & (g744) & (g3105) & (!g3106) & (!g3164) & (!g3187)) + ((!g700) & (g744) & (g3105) & (!g3106) & (!g3164) & (g3187)) + ((!g700) & (g744) & (g3105) & (!g3106) & (g3164) & (g3187)) + ((!g700) & (g744) & (g3105) & (g3106) & (!g3164) & (g3187)) + ((!g700) & (g744) & (g3105) & (g3106) & (g3164) & (g3187)) + ((g700) & (!g744) & (!g3105) & (!g3106) & (!g3164) & (!g3187)) + ((g700) & (!g744) & (!g3105) & (!g3106) & (g3164) & (!g3187)) + ((g700) & (!g744) & (!g3105) & (g3106) & (!g3164) & (!g3187)) + ((g700) & (!g744) & (g3105) & (!g3106) & (!g3164) & (g3187)) + ((g700) & (!g744) & (g3105) & (!g3106) & (g3164) & (g3187)) + ((g700) & (!g744) & (g3105) & (g3106) & (!g3164) & (g3187)) + ((g700) & (!g744) & (g3105) & (g3106) & (g3164) & (!g3187)) + ((g700) & (!g744) & (g3105) & (g3106) & (g3164) & (g3187)) + ((g700) & (g744) & (!g3105) & (!g3106) & (!g3164) & (!g3187)) + ((g700) & (g744) & (g3105) & (!g3106) & (!g3164) & (g3187)) + ((g700) & (g744) & (g3105) & (!g3106) & (g3164) & (!g3187)) + ((g700) & (g744) & (g3105) & (!g3106) & (g3164) & (g3187)) + ((g700) & (g744) & (g3105) & (g3106) & (!g3164) & (!g3187)) + ((g700) & (g744) & (g3105) & (g3106) & (!g3164) & (g3187)) + ((g700) & (g744) & (g3105) & (g3106) & (g3164) & (!g3187)) + ((g700) & (g744) & (g3105) & (g3106) & (g3164) & (g3187)));
	assign g3212 = (((!g744) & (!g3106) & (g3164) & (!g3187)) + ((!g744) & (g3106) & (!g3164) & (!g3187)) + ((!g744) & (g3106) & (!g3164) & (g3187)) + ((!g744) & (g3106) & (g3164) & (g3187)) + ((g744) & (!g3106) & (!g3164) & (!g3187)) + ((g744) & (g3106) & (!g3164) & (g3187)) + ((g744) & (g3106) & (g3164) & (!g3187)) + ((g744) & (g3106) & (g3164) & (g3187)));
	assign g3213 = (((!g803) & (!g851) & (!g3108) & (g3109) & (g3163) & (!g3187)) + ((!g803) & (!g851) & (g3108) & (!g3109) & (!g3163) & (!g3187)) + ((!g803) & (!g851) & (g3108) & (!g3109) & (!g3163) & (g3187)) + ((!g803) & (!g851) & (g3108) & (!g3109) & (g3163) & (!g3187)) + ((!g803) & (!g851) & (g3108) & (!g3109) & (g3163) & (g3187)) + ((!g803) & (!g851) & (g3108) & (g3109) & (!g3163) & (!g3187)) + ((!g803) & (!g851) & (g3108) & (g3109) & (!g3163) & (g3187)) + ((!g803) & (!g851) & (g3108) & (g3109) & (g3163) & (g3187)) + ((!g803) & (g851) & (!g3108) & (!g3109) & (g3163) & (!g3187)) + ((!g803) & (g851) & (!g3108) & (g3109) & (!g3163) & (!g3187)) + ((!g803) & (g851) & (!g3108) & (g3109) & (g3163) & (!g3187)) + ((!g803) & (g851) & (g3108) & (!g3109) & (!g3163) & (!g3187)) + ((!g803) & (g851) & (g3108) & (!g3109) & (!g3163) & (g3187)) + ((!g803) & (g851) & (g3108) & (!g3109) & (g3163) & (g3187)) + ((!g803) & (g851) & (g3108) & (g3109) & (!g3163) & (g3187)) + ((!g803) & (g851) & (g3108) & (g3109) & (g3163) & (g3187)) + ((g803) & (!g851) & (!g3108) & (!g3109) & (!g3163) & (!g3187)) + ((g803) & (!g851) & (!g3108) & (!g3109) & (g3163) & (!g3187)) + ((g803) & (!g851) & (!g3108) & (g3109) & (!g3163) & (!g3187)) + ((g803) & (!g851) & (g3108) & (!g3109) & (!g3163) & (g3187)) + ((g803) & (!g851) & (g3108) & (!g3109) & (g3163) & (g3187)) + ((g803) & (!g851) & (g3108) & (g3109) & (!g3163) & (g3187)) + ((g803) & (!g851) & (g3108) & (g3109) & (g3163) & (!g3187)) + ((g803) & (!g851) & (g3108) & (g3109) & (g3163) & (g3187)) + ((g803) & (g851) & (!g3108) & (!g3109) & (!g3163) & (!g3187)) + ((g803) & (g851) & (g3108) & (!g3109) & (!g3163) & (g3187)) + ((g803) & (g851) & (g3108) & (!g3109) & (g3163) & (!g3187)) + ((g803) & (g851) & (g3108) & (!g3109) & (g3163) & (g3187)) + ((g803) & (g851) & (g3108) & (g3109) & (!g3163) & (!g3187)) + ((g803) & (g851) & (g3108) & (g3109) & (!g3163) & (g3187)) + ((g803) & (g851) & (g3108) & (g3109) & (g3163) & (!g3187)) + ((g803) & (g851) & (g3108) & (g3109) & (g3163) & (g3187)));
	assign g3214 = (((!g851) & (!g3109) & (g3163) & (!g3187)) + ((!g851) & (g3109) & (!g3163) & (!g3187)) + ((!g851) & (g3109) & (!g3163) & (g3187)) + ((!g851) & (g3109) & (g3163) & (g3187)) + ((g851) & (!g3109) & (!g3163) & (!g3187)) + ((g851) & (g3109) & (!g3163) & (g3187)) + ((g851) & (g3109) & (g3163) & (!g3187)) + ((g851) & (g3109) & (g3163) & (g3187)));
	assign g3215 = (((!g914) & (!g1032) & (!g3111) & (g3112) & (g3162) & (!g3187)) + ((!g914) & (!g1032) & (g3111) & (!g3112) & (!g3162) & (!g3187)) + ((!g914) & (!g1032) & (g3111) & (!g3112) & (!g3162) & (g3187)) + ((!g914) & (!g1032) & (g3111) & (!g3112) & (g3162) & (!g3187)) + ((!g914) & (!g1032) & (g3111) & (!g3112) & (g3162) & (g3187)) + ((!g914) & (!g1032) & (g3111) & (g3112) & (!g3162) & (!g3187)) + ((!g914) & (!g1032) & (g3111) & (g3112) & (!g3162) & (g3187)) + ((!g914) & (!g1032) & (g3111) & (g3112) & (g3162) & (g3187)) + ((!g914) & (g1032) & (!g3111) & (!g3112) & (g3162) & (!g3187)) + ((!g914) & (g1032) & (!g3111) & (g3112) & (!g3162) & (!g3187)) + ((!g914) & (g1032) & (!g3111) & (g3112) & (g3162) & (!g3187)) + ((!g914) & (g1032) & (g3111) & (!g3112) & (!g3162) & (!g3187)) + ((!g914) & (g1032) & (g3111) & (!g3112) & (!g3162) & (g3187)) + ((!g914) & (g1032) & (g3111) & (!g3112) & (g3162) & (g3187)) + ((!g914) & (g1032) & (g3111) & (g3112) & (!g3162) & (g3187)) + ((!g914) & (g1032) & (g3111) & (g3112) & (g3162) & (g3187)) + ((g914) & (!g1032) & (!g3111) & (!g3112) & (!g3162) & (!g3187)) + ((g914) & (!g1032) & (!g3111) & (!g3112) & (g3162) & (!g3187)) + ((g914) & (!g1032) & (!g3111) & (g3112) & (!g3162) & (!g3187)) + ((g914) & (!g1032) & (g3111) & (!g3112) & (!g3162) & (g3187)) + ((g914) & (!g1032) & (g3111) & (!g3112) & (g3162) & (g3187)) + ((g914) & (!g1032) & (g3111) & (g3112) & (!g3162) & (g3187)) + ((g914) & (!g1032) & (g3111) & (g3112) & (g3162) & (!g3187)) + ((g914) & (!g1032) & (g3111) & (g3112) & (g3162) & (g3187)) + ((g914) & (g1032) & (!g3111) & (!g3112) & (!g3162) & (!g3187)) + ((g914) & (g1032) & (g3111) & (!g3112) & (!g3162) & (g3187)) + ((g914) & (g1032) & (g3111) & (!g3112) & (g3162) & (!g3187)) + ((g914) & (g1032) & (g3111) & (!g3112) & (g3162) & (g3187)) + ((g914) & (g1032) & (g3111) & (g3112) & (!g3162) & (!g3187)) + ((g914) & (g1032) & (g3111) & (g3112) & (!g3162) & (g3187)) + ((g914) & (g1032) & (g3111) & (g3112) & (g3162) & (!g3187)) + ((g914) & (g1032) & (g3111) & (g3112) & (g3162) & (g3187)));
	assign g3216 = (((!g1032) & (!g3112) & (g3162) & (!g3187)) + ((!g1032) & (g3112) & (!g3162) & (!g3187)) + ((!g1032) & (g3112) & (!g3162) & (g3187)) + ((!g1032) & (g3112) & (g3162) & (g3187)) + ((g1032) & (!g3112) & (!g3162) & (!g3187)) + ((g1032) & (g3112) & (!g3162) & (g3187)) + ((g1032) & (g3112) & (g3162) & (!g3187)) + ((g1032) & (g3112) & (g3162) & (g3187)));
	assign g3217 = (((!g1030) & (!g1160) & (!g3114) & (g3115) & (g3161) & (!g3187)) + ((!g1030) & (!g1160) & (g3114) & (!g3115) & (!g3161) & (!g3187)) + ((!g1030) & (!g1160) & (g3114) & (!g3115) & (!g3161) & (g3187)) + ((!g1030) & (!g1160) & (g3114) & (!g3115) & (g3161) & (!g3187)) + ((!g1030) & (!g1160) & (g3114) & (!g3115) & (g3161) & (g3187)) + ((!g1030) & (!g1160) & (g3114) & (g3115) & (!g3161) & (!g3187)) + ((!g1030) & (!g1160) & (g3114) & (g3115) & (!g3161) & (g3187)) + ((!g1030) & (!g1160) & (g3114) & (g3115) & (g3161) & (g3187)) + ((!g1030) & (g1160) & (!g3114) & (!g3115) & (g3161) & (!g3187)) + ((!g1030) & (g1160) & (!g3114) & (g3115) & (!g3161) & (!g3187)) + ((!g1030) & (g1160) & (!g3114) & (g3115) & (g3161) & (!g3187)) + ((!g1030) & (g1160) & (g3114) & (!g3115) & (!g3161) & (!g3187)) + ((!g1030) & (g1160) & (g3114) & (!g3115) & (!g3161) & (g3187)) + ((!g1030) & (g1160) & (g3114) & (!g3115) & (g3161) & (g3187)) + ((!g1030) & (g1160) & (g3114) & (g3115) & (!g3161) & (g3187)) + ((!g1030) & (g1160) & (g3114) & (g3115) & (g3161) & (g3187)) + ((g1030) & (!g1160) & (!g3114) & (!g3115) & (!g3161) & (!g3187)) + ((g1030) & (!g1160) & (!g3114) & (!g3115) & (g3161) & (!g3187)) + ((g1030) & (!g1160) & (!g3114) & (g3115) & (!g3161) & (!g3187)) + ((g1030) & (!g1160) & (g3114) & (!g3115) & (!g3161) & (g3187)) + ((g1030) & (!g1160) & (g3114) & (!g3115) & (g3161) & (g3187)) + ((g1030) & (!g1160) & (g3114) & (g3115) & (!g3161) & (g3187)) + ((g1030) & (!g1160) & (g3114) & (g3115) & (g3161) & (!g3187)) + ((g1030) & (!g1160) & (g3114) & (g3115) & (g3161) & (g3187)) + ((g1030) & (g1160) & (!g3114) & (!g3115) & (!g3161) & (!g3187)) + ((g1030) & (g1160) & (g3114) & (!g3115) & (!g3161) & (g3187)) + ((g1030) & (g1160) & (g3114) & (!g3115) & (g3161) & (!g3187)) + ((g1030) & (g1160) & (g3114) & (!g3115) & (g3161) & (g3187)) + ((g1030) & (g1160) & (g3114) & (g3115) & (!g3161) & (!g3187)) + ((g1030) & (g1160) & (g3114) & (g3115) & (!g3161) & (g3187)) + ((g1030) & (g1160) & (g3114) & (g3115) & (g3161) & (!g3187)) + ((g1030) & (g1160) & (g3114) & (g3115) & (g3161) & (g3187)));
	assign g3218 = (((!g1160) & (!g3115) & (g3161) & (!g3187)) + ((!g1160) & (g3115) & (!g3161) & (!g3187)) + ((!g1160) & (g3115) & (!g3161) & (g3187)) + ((!g1160) & (g3115) & (g3161) & (g3187)) + ((g1160) & (!g3115) & (!g3161) & (!g3187)) + ((g1160) & (g3115) & (!g3161) & (g3187)) + ((g1160) & (g3115) & (g3161) & (!g3187)) + ((g1160) & (g3115) & (g3161) & (g3187)));
	assign g3219 = (((!g1154) & (!g1295) & (!g3117) & (g3118) & (g3160) & (!g3187)) + ((!g1154) & (!g1295) & (g3117) & (!g3118) & (!g3160) & (!g3187)) + ((!g1154) & (!g1295) & (g3117) & (!g3118) & (!g3160) & (g3187)) + ((!g1154) & (!g1295) & (g3117) & (!g3118) & (g3160) & (!g3187)) + ((!g1154) & (!g1295) & (g3117) & (!g3118) & (g3160) & (g3187)) + ((!g1154) & (!g1295) & (g3117) & (g3118) & (!g3160) & (!g3187)) + ((!g1154) & (!g1295) & (g3117) & (g3118) & (!g3160) & (g3187)) + ((!g1154) & (!g1295) & (g3117) & (g3118) & (g3160) & (g3187)) + ((!g1154) & (g1295) & (!g3117) & (!g3118) & (g3160) & (!g3187)) + ((!g1154) & (g1295) & (!g3117) & (g3118) & (!g3160) & (!g3187)) + ((!g1154) & (g1295) & (!g3117) & (g3118) & (g3160) & (!g3187)) + ((!g1154) & (g1295) & (g3117) & (!g3118) & (!g3160) & (!g3187)) + ((!g1154) & (g1295) & (g3117) & (!g3118) & (!g3160) & (g3187)) + ((!g1154) & (g1295) & (g3117) & (!g3118) & (g3160) & (g3187)) + ((!g1154) & (g1295) & (g3117) & (g3118) & (!g3160) & (g3187)) + ((!g1154) & (g1295) & (g3117) & (g3118) & (g3160) & (g3187)) + ((g1154) & (!g1295) & (!g3117) & (!g3118) & (!g3160) & (!g3187)) + ((g1154) & (!g1295) & (!g3117) & (!g3118) & (g3160) & (!g3187)) + ((g1154) & (!g1295) & (!g3117) & (g3118) & (!g3160) & (!g3187)) + ((g1154) & (!g1295) & (g3117) & (!g3118) & (!g3160) & (g3187)) + ((g1154) & (!g1295) & (g3117) & (!g3118) & (g3160) & (g3187)) + ((g1154) & (!g1295) & (g3117) & (g3118) & (!g3160) & (g3187)) + ((g1154) & (!g1295) & (g3117) & (g3118) & (g3160) & (!g3187)) + ((g1154) & (!g1295) & (g3117) & (g3118) & (g3160) & (g3187)) + ((g1154) & (g1295) & (!g3117) & (!g3118) & (!g3160) & (!g3187)) + ((g1154) & (g1295) & (g3117) & (!g3118) & (!g3160) & (g3187)) + ((g1154) & (g1295) & (g3117) & (!g3118) & (g3160) & (!g3187)) + ((g1154) & (g1295) & (g3117) & (!g3118) & (g3160) & (g3187)) + ((g1154) & (g1295) & (g3117) & (g3118) & (!g3160) & (!g3187)) + ((g1154) & (g1295) & (g3117) & (g3118) & (!g3160) & (g3187)) + ((g1154) & (g1295) & (g3117) & (g3118) & (g3160) & (!g3187)) + ((g1154) & (g1295) & (g3117) & (g3118) & (g3160) & (g3187)));
	assign g3220 = (((!g1295) & (!g3118) & (g3160) & (!g3187)) + ((!g1295) & (g3118) & (!g3160) & (!g3187)) + ((!g1295) & (g3118) & (!g3160) & (g3187)) + ((!g1295) & (g3118) & (g3160) & (g3187)) + ((g1295) & (!g3118) & (!g3160) & (!g3187)) + ((g1295) & (g3118) & (!g3160) & (g3187)) + ((g1295) & (g3118) & (g3160) & (!g3187)) + ((g1295) & (g3118) & (g3160) & (g3187)));
	assign g3221 = (((!g1285) & (!g1437) & (!g3120) & (g3121) & (g3159) & (!g3187)) + ((!g1285) & (!g1437) & (g3120) & (!g3121) & (!g3159) & (!g3187)) + ((!g1285) & (!g1437) & (g3120) & (!g3121) & (!g3159) & (g3187)) + ((!g1285) & (!g1437) & (g3120) & (!g3121) & (g3159) & (!g3187)) + ((!g1285) & (!g1437) & (g3120) & (!g3121) & (g3159) & (g3187)) + ((!g1285) & (!g1437) & (g3120) & (g3121) & (!g3159) & (!g3187)) + ((!g1285) & (!g1437) & (g3120) & (g3121) & (!g3159) & (g3187)) + ((!g1285) & (!g1437) & (g3120) & (g3121) & (g3159) & (g3187)) + ((!g1285) & (g1437) & (!g3120) & (!g3121) & (g3159) & (!g3187)) + ((!g1285) & (g1437) & (!g3120) & (g3121) & (!g3159) & (!g3187)) + ((!g1285) & (g1437) & (!g3120) & (g3121) & (g3159) & (!g3187)) + ((!g1285) & (g1437) & (g3120) & (!g3121) & (!g3159) & (!g3187)) + ((!g1285) & (g1437) & (g3120) & (!g3121) & (!g3159) & (g3187)) + ((!g1285) & (g1437) & (g3120) & (!g3121) & (g3159) & (g3187)) + ((!g1285) & (g1437) & (g3120) & (g3121) & (!g3159) & (g3187)) + ((!g1285) & (g1437) & (g3120) & (g3121) & (g3159) & (g3187)) + ((g1285) & (!g1437) & (!g3120) & (!g3121) & (!g3159) & (!g3187)) + ((g1285) & (!g1437) & (!g3120) & (!g3121) & (g3159) & (!g3187)) + ((g1285) & (!g1437) & (!g3120) & (g3121) & (!g3159) & (!g3187)) + ((g1285) & (!g1437) & (g3120) & (!g3121) & (!g3159) & (g3187)) + ((g1285) & (!g1437) & (g3120) & (!g3121) & (g3159) & (g3187)) + ((g1285) & (!g1437) & (g3120) & (g3121) & (!g3159) & (g3187)) + ((g1285) & (!g1437) & (g3120) & (g3121) & (g3159) & (!g3187)) + ((g1285) & (!g1437) & (g3120) & (g3121) & (g3159) & (g3187)) + ((g1285) & (g1437) & (!g3120) & (!g3121) & (!g3159) & (!g3187)) + ((g1285) & (g1437) & (g3120) & (!g3121) & (!g3159) & (g3187)) + ((g1285) & (g1437) & (g3120) & (!g3121) & (g3159) & (!g3187)) + ((g1285) & (g1437) & (g3120) & (!g3121) & (g3159) & (g3187)) + ((g1285) & (g1437) & (g3120) & (g3121) & (!g3159) & (!g3187)) + ((g1285) & (g1437) & (g3120) & (g3121) & (!g3159) & (g3187)) + ((g1285) & (g1437) & (g3120) & (g3121) & (g3159) & (!g3187)) + ((g1285) & (g1437) & (g3120) & (g3121) & (g3159) & (g3187)));
	assign g3222 = (((!g1437) & (!g3121) & (g3159) & (!g3187)) + ((!g1437) & (g3121) & (!g3159) & (!g3187)) + ((!g1437) & (g3121) & (!g3159) & (g3187)) + ((!g1437) & (g3121) & (g3159) & (g3187)) + ((g1437) & (!g3121) & (!g3159) & (!g3187)) + ((g1437) & (g3121) & (!g3159) & (g3187)) + ((g1437) & (g3121) & (g3159) & (!g3187)) + ((g1437) & (g3121) & (g3159) & (g3187)));
	assign g3223 = (((!g1423) & (!g1586) & (!g3123) & (g3124) & (g3158) & (!g3187)) + ((!g1423) & (!g1586) & (g3123) & (!g3124) & (!g3158) & (!g3187)) + ((!g1423) & (!g1586) & (g3123) & (!g3124) & (!g3158) & (g3187)) + ((!g1423) & (!g1586) & (g3123) & (!g3124) & (g3158) & (!g3187)) + ((!g1423) & (!g1586) & (g3123) & (!g3124) & (g3158) & (g3187)) + ((!g1423) & (!g1586) & (g3123) & (g3124) & (!g3158) & (!g3187)) + ((!g1423) & (!g1586) & (g3123) & (g3124) & (!g3158) & (g3187)) + ((!g1423) & (!g1586) & (g3123) & (g3124) & (g3158) & (g3187)) + ((!g1423) & (g1586) & (!g3123) & (!g3124) & (g3158) & (!g3187)) + ((!g1423) & (g1586) & (!g3123) & (g3124) & (!g3158) & (!g3187)) + ((!g1423) & (g1586) & (!g3123) & (g3124) & (g3158) & (!g3187)) + ((!g1423) & (g1586) & (g3123) & (!g3124) & (!g3158) & (!g3187)) + ((!g1423) & (g1586) & (g3123) & (!g3124) & (!g3158) & (g3187)) + ((!g1423) & (g1586) & (g3123) & (!g3124) & (g3158) & (g3187)) + ((!g1423) & (g1586) & (g3123) & (g3124) & (!g3158) & (g3187)) + ((!g1423) & (g1586) & (g3123) & (g3124) & (g3158) & (g3187)) + ((g1423) & (!g1586) & (!g3123) & (!g3124) & (!g3158) & (!g3187)) + ((g1423) & (!g1586) & (!g3123) & (!g3124) & (g3158) & (!g3187)) + ((g1423) & (!g1586) & (!g3123) & (g3124) & (!g3158) & (!g3187)) + ((g1423) & (!g1586) & (g3123) & (!g3124) & (!g3158) & (g3187)) + ((g1423) & (!g1586) & (g3123) & (!g3124) & (g3158) & (g3187)) + ((g1423) & (!g1586) & (g3123) & (g3124) & (!g3158) & (g3187)) + ((g1423) & (!g1586) & (g3123) & (g3124) & (g3158) & (!g3187)) + ((g1423) & (!g1586) & (g3123) & (g3124) & (g3158) & (g3187)) + ((g1423) & (g1586) & (!g3123) & (!g3124) & (!g3158) & (!g3187)) + ((g1423) & (g1586) & (g3123) & (!g3124) & (!g3158) & (g3187)) + ((g1423) & (g1586) & (g3123) & (!g3124) & (g3158) & (!g3187)) + ((g1423) & (g1586) & (g3123) & (!g3124) & (g3158) & (g3187)) + ((g1423) & (g1586) & (g3123) & (g3124) & (!g3158) & (!g3187)) + ((g1423) & (g1586) & (g3123) & (g3124) & (!g3158) & (g3187)) + ((g1423) & (g1586) & (g3123) & (g3124) & (g3158) & (!g3187)) + ((g1423) & (g1586) & (g3123) & (g3124) & (g3158) & (g3187)));
	assign g3224 = (((!g1586) & (!g3124) & (g3158) & (!g3187)) + ((!g1586) & (g3124) & (!g3158) & (!g3187)) + ((!g1586) & (g3124) & (!g3158) & (g3187)) + ((!g1586) & (g3124) & (g3158) & (g3187)) + ((g1586) & (!g3124) & (!g3158) & (!g3187)) + ((g1586) & (g3124) & (!g3158) & (g3187)) + ((g1586) & (g3124) & (g3158) & (!g3187)) + ((g1586) & (g3124) & (g3158) & (g3187)));
	assign g3225 = (((!g1568) & (!g1742) & (!g3126) & (g3127) & (g3157) & (!g3187)) + ((!g1568) & (!g1742) & (g3126) & (!g3127) & (!g3157) & (!g3187)) + ((!g1568) & (!g1742) & (g3126) & (!g3127) & (!g3157) & (g3187)) + ((!g1568) & (!g1742) & (g3126) & (!g3127) & (g3157) & (!g3187)) + ((!g1568) & (!g1742) & (g3126) & (!g3127) & (g3157) & (g3187)) + ((!g1568) & (!g1742) & (g3126) & (g3127) & (!g3157) & (!g3187)) + ((!g1568) & (!g1742) & (g3126) & (g3127) & (!g3157) & (g3187)) + ((!g1568) & (!g1742) & (g3126) & (g3127) & (g3157) & (g3187)) + ((!g1568) & (g1742) & (!g3126) & (!g3127) & (g3157) & (!g3187)) + ((!g1568) & (g1742) & (!g3126) & (g3127) & (!g3157) & (!g3187)) + ((!g1568) & (g1742) & (!g3126) & (g3127) & (g3157) & (!g3187)) + ((!g1568) & (g1742) & (g3126) & (!g3127) & (!g3157) & (!g3187)) + ((!g1568) & (g1742) & (g3126) & (!g3127) & (!g3157) & (g3187)) + ((!g1568) & (g1742) & (g3126) & (!g3127) & (g3157) & (g3187)) + ((!g1568) & (g1742) & (g3126) & (g3127) & (!g3157) & (g3187)) + ((!g1568) & (g1742) & (g3126) & (g3127) & (g3157) & (g3187)) + ((g1568) & (!g1742) & (!g3126) & (!g3127) & (!g3157) & (!g3187)) + ((g1568) & (!g1742) & (!g3126) & (!g3127) & (g3157) & (!g3187)) + ((g1568) & (!g1742) & (!g3126) & (g3127) & (!g3157) & (!g3187)) + ((g1568) & (!g1742) & (g3126) & (!g3127) & (!g3157) & (g3187)) + ((g1568) & (!g1742) & (g3126) & (!g3127) & (g3157) & (g3187)) + ((g1568) & (!g1742) & (g3126) & (g3127) & (!g3157) & (g3187)) + ((g1568) & (!g1742) & (g3126) & (g3127) & (g3157) & (!g3187)) + ((g1568) & (!g1742) & (g3126) & (g3127) & (g3157) & (g3187)) + ((g1568) & (g1742) & (!g3126) & (!g3127) & (!g3157) & (!g3187)) + ((g1568) & (g1742) & (g3126) & (!g3127) & (!g3157) & (g3187)) + ((g1568) & (g1742) & (g3126) & (!g3127) & (g3157) & (!g3187)) + ((g1568) & (g1742) & (g3126) & (!g3127) & (g3157) & (g3187)) + ((g1568) & (g1742) & (g3126) & (g3127) & (!g3157) & (!g3187)) + ((g1568) & (g1742) & (g3126) & (g3127) & (!g3157) & (g3187)) + ((g1568) & (g1742) & (g3126) & (g3127) & (g3157) & (!g3187)) + ((g1568) & (g1742) & (g3126) & (g3127) & (g3157) & (g3187)));
	assign g3226 = (((!g1742) & (!g3127) & (g3157) & (!g3187)) + ((!g1742) & (g3127) & (!g3157) & (!g3187)) + ((!g1742) & (g3127) & (!g3157) & (g3187)) + ((!g1742) & (g3127) & (g3157) & (g3187)) + ((g1742) & (!g3127) & (!g3157) & (!g3187)) + ((g1742) & (g3127) & (!g3157) & (g3187)) + ((g1742) & (g3127) & (g3157) & (!g3187)) + ((g1742) & (g3127) & (g3157) & (g3187)));
	assign g3227 = (((!g1720) & (!g1905) & (!g3129) & (g3130) & (g3156) & (!g3187)) + ((!g1720) & (!g1905) & (g3129) & (!g3130) & (!g3156) & (!g3187)) + ((!g1720) & (!g1905) & (g3129) & (!g3130) & (!g3156) & (g3187)) + ((!g1720) & (!g1905) & (g3129) & (!g3130) & (g3156) & (!g3187)) + ((!g1720) & (!g1905) & (g3129) & (!g3130) & (g3156) & (g3187)) + ((!g1720) & (!g1905) & (g3129) & (g3130) & (!g3156) & (!g3187)) + ((!g1720) & (!g1905) & (g3129) & (g3130) & (!g3156) & (g3187)) + ((!g1720) & (!g1905) & (g3129) & (g3130) & (g3156) & (g3187)) + ((!g1720) & (g1905) & (!g3129) & (!g3130) & (g3156) & (!g3187)) + ((!g1720) & (g1905) & (!g3129) & (g3130) & (!g3156) & (!g3187)) + ((!g1720) & (g1905) & (!g3129) & (g3130) & (g3156) & (!g3187)) + ((!g1720) & (g1905) & (g3129) & (!g3130) & (!g3156) & (!g3187)) + ((!g1720) & (g1905) & (g3129) & (!g3130) & (!g3156) & (g3187)) + ((!g1720) & (g1905) & (g3129) & (!g3130) & (g3156) & (g3187)) + ((!g1720) & (g1905) & (g3129) & (g3130) & (!g3156) & (g3187)) + ((!g1720) & (g1905) & (g3129) & (g3130) & (g3156) & (g3187)) + ((g1720) & (!g1905) & (!g3129) & (!g3130) & (!g3156) & (!g3187)) + ((g1720) & (!g1905) & (!g3129) & (!g3130) & (g3156) & (!g3187)) + ((g1720) & (!g1905) & (!g3129) & (g3130) & (!g3156) & (!g3187)) + ((g1720) & (!g1905) & (g3129) & (!g3130) & (!g3156) & (g3187)) + ((g1720) & (!g1905) & (g3129) & (!g3130) & (g3156) & (g3187)) + ((g1720) & (!g1905) & (g3129) & (g3130) & (!g3156) & (g3187)) + ((g1720) & (!g1905) & (g3129) & (g3130) & (g3156) & (!g3187)) + ((g1720) & (!g1905) & (g3129) & (g3130) & (g3156) & (g3187)) + ((g1720) & (g1905) & (!g3129) & (!g3130) & (!g3156) & (!g3187)) + ((g1720) & (g1905) & (g3129) & (!g3130) & (!g3156) & (g3187)) + ((g1720) & (g1905) & (g3129) & (!g3130) & (g3156) & (!g3187)) + ((g1720) & (g1905) & (g3129) & (!g3130) & (g3156) & (g3187)) + ((g1720) & (g1905) & (g3129) & (g3130) & (!g3156) & (!g3187)) + ((g1720) & (g1905) & (g3129) & (g3130) & (!g3156) & (g3187)) + ((g1720) & (g1905) & (g3129) & (g3130) & (g3156) & (!g3187)) + ((g1720) & (g1905) & (g3129) & (g3130) & (g3156) & (g3187)));
	assign g3228 = (((!g1905) & (!g3130) & (g3156) & (!g3187)) + ((!g1905) & (g3130) & (!g3156) & (!g3187)) + ((!g1905) & (g3130) & (!g3156) & (g3187)) + ((!g1905) & (g3130) & (g3156) & (g3187)) + ((g1905) & (!g3130) & (!g3156) & (!g3187)) + ((g1905) & (g3130) & (!g3156) & (g3187)) + ((g1905) & (g3130) & (g3156) & (!g3187)) + ((g1905) & (g3130) & (g3156) & (g3187)));
	assign g3229 = (((!g1879) & (!g2075) & (!g3132) & (g3133) & (g3155) & (!g3187)) + ((!g1879) & (!g2075) & (g3132) & (!g3133) & (!g3155) & (!g3187)) + ((!g1879) & (!g2075) & (g3132) & (!g3133) & (!g3155) & (g3187)) + ((!g1879) & (!g2075) & (g3132) & (!g3133) & (g3155) & (!g3187)) + ((!g1879) & (!g2075) & (g3132) & (!g3133) & (g3155) & (g3187)) + ((!g1879) & (!g2075) & (g3132) & (g3133) & (!g3155) & (!g3187)) + ((!g1879) & (!g2075) & (g3132) & (g3133) & (!g3155) & (g3187)) + ((!g1879) & (!g2075) & (g3132) & (g3133) & (g3155) & (g3187)) + ((!g1879) & (g2075) & (!g3132) & (!g3133) & (g3155) & (!g3187)) + ((!g1879) & (g2075) & (!g3132) & (g3133) & (!g3155) & (!g3187)) + ((!g1879) & (g2075) & (!g3132) & (g3133) & (g3155) & (!g3187)) + ((!g1879) & (g2075) & (g3132) & (!g3133) & (!g3155) & (!g3187)) + ((!g1879) & (g2075) & (g3132) & (!g3133) & (!g3155) & (g3187)) + ((!g1879) & (g2075) & (g3132) & (!g3133) & (g3155) & (g3187)) + ((!g1879) & (g2075) & (g3132) & (g3133) & (!g3155) & (g3187)) + ((!g1879) & (g2075) & (g3132) & (g3133) & (g3155) & (g3187)) + ((g1879) & (!g2075) & (!g3132) & (!g3133) & (!g3155) & (!g3187)) + ((g1879) & (!g2075) & (!g3132) & (!g3133) & (g3155) & (!g3187)) + ((g1879) & (!g2075) & (!g3132) & (g3133) & (!g3155) & (!g3187)) + ((g1879) & (!g2075) & (g3132) & (!g3133) & (!g3155) & (g3187)) + ((g1879) & (!g2075) & (g3132) & (!g3133) & (g3155) & (g3187)) + ((g1879) & (!g2075) & (g3132) & (g3133) & (!g3155) & (g3187)) + ((g1879) & (!g2075) & (g3132) & (g3133) & (g3155) & (!g3187)) + ((g1879) & (!g2075) & (g3132) & (g3133) & (g3155) & (g3187)) + ((g1879) & (g2075) & (!g3132) & (!g3133) & (!g3155) & (!g3187)) + ((g1879) & (g2075) & (g3132) & (!g3133) & (!g3155) & (g3187)) + ((g1879) & (g2075) & (g3132) & (!g3133) & (g3155) & (!g3187)) + ((g1879) & (g2075) & (g3132) & (!g3133) & (g3155) & (g3187)) + ((g1879) & (g2075) & (g3132) & (g3133) & (!g3155) & (!g3187)) + ((g1879) & (g2075) & (g3132) & (g3133) & (!g3155) & (g3187)) + ((g1879) & (g2075) & (g3132) & (g3133) & (g3155) & (!g3187)) + ((g1879) & (g2075) & (g3132) & (g3133) & (g3155) & (g3187)));
	assign g3230 = (((!g2075) & (!g3133) & (g3155) & (!g3187)) + ((!g2075) & (g3133) & (!g3155) & (!g3187)) + ((!g2075) & (g3133) & (!g3155) & (g3187)) + ((!g2075) & (g3133) & (g3155) & (g3187)) + ((g2075) & (!g3133) & (!g3155) & (!g3187)) + ((g2075) & (g3133) & (!g3155) & (g3187)) + ((g2075) & (g3133) & (g3155) & (!g3187)) + ((g2075) & (g3133) & (g3155) & (g3187)));
	assign g3231 = (((!g2045) & (!g2252) & (!g3135) & (g3136) & (g3154) & (!g3187)) + ((!g2045) & (!g2252) & (g3135) & (!g3136) & (!g3154) & (!g3187)) + ((!g2045) & (!g2252) & (g3135) & (!g3136) & (!g3154) & (g3187)) + ((!g2045) & (!g2252) & (g3135) & (!g3136) & (g3154) & (!g3187)) + ((!g2045) & (!g2252) & (g3135) & (!g3136) & (g3154) & (g3187)) + ((!g2045) & (!g2252) & (g3135) & (g3136) & (!g3154) & (!g3187)) + ((!g2045) & (!g2252) & (g3135) & (g3136) & (!g3154) & (g3187)) + ((!g2045) & (!g2252) & (g3135) & (g3136) & (g3154) & (g3187)) + ((!g2045) & (g2252) & (!g3135) & (!g3136) & (g3154) & (!g3187)) + ((!g2045) & (g2252) & (!g3135) & (g3136) & (!g3154) & (!g3187)) + ((!g2045) & (g2252) & (!g3135) & (g3136) & (g3154) & (!g3187)) + ((!g2045) & (g2252) & (g3135) & (!g3136) & (!g3154) & (!g3187)) + ((!g2045) & (g2252) & (g3135) & (!g3136) & (!g3154) & (g3187)) + ((!g2045) & (g2252) & (g3135) & (!g3136) & (g3154) & (g3187)) + ((!g2045) & (g2252) & (g3135) & (g3136) & (!g3154) & (g3187)) + ((!g2045) & (g2252) & (g3135) & (g3136) & (g3154) & (g3187)) + ((g2045) & (!g2252) & (!g3135) & (!g3136) & (!g3154) & (!g3187)) + ((g2045) & (!g2252) & (!g3135) & (!g3136) & (g3154) & (!g3187)) + ((g2045) & (!g2252) & (!g3135) & (g3136) & (!g3154) & (!g3187)) + ((g2045) & (!g2252) & (g3135) & (!g3136) & (!g3154) & (g3187)) + ((g2045) & (!g2252) & (g3135) & (!g3136) & (g3154) & (g3187)) + ((g2045) & (!g2252) & (g3135) & (g3136) & (!g3154) & (g3187)) + ((g2045) & (!g2252) & (g3135) & (g3136) & (g3154) & (!g3187)) + ((g2045) & (!g2252) & (g3135) & (g3136) & (g3154) & (g3187)) + ((g2045) & (g2252) & (!g3135) & (!g3136) & (!g3154) & (!g3187)) + ((g2045) & (g2252) & (g3135) & (!g3136) & (!g3154) & (g3187)) + ((g2045) & (g2252) & (g3135) & (!g3136) & (g3154) & (!g3187)) + ((g2045) & (g2252) & (g3135) & (!g3136) & (g3154) & (g3187)) + ((g2045) & (g2252) & (g3135) & (g3136) & (!g3154) & (!g3187)) + ((g2045) & (g2252) & (g3135) & (g3136) & (!g3154) & (g3187)) + ((g2045) & (g2252) & (g3135) & (g3136) & (g3154) & (!g3187)) + ((g2045) & (g2252) & (g3135) & (g3136) & (g3154) & (g3187)));
	assign g3232 = (((!g2252) & (!g3136) & (g3154) & (!g3187)) + ((!g2252) & (g3136) & (!g3154) & (!g3187)) + ((!g2252) & (g3136) & (!g3154) & (g3187)) + ((!g2252) & (g3136) & (g3154) & (g3187)) + ((g2252) & (!g3136) & (!g3154) & (!g3187)) + ((g2252) & (g3136) & (!g3154) & (g3187)) + ((g2252) & (g3136) & (g3154) & (!g3187)) + ((g2252) & (g3136) & (g3154) & (g3187)));
	assign g3233 = (((!g2218) & (!g2436) & (!g3138) & (g3139) & (g3153) & (!g3187)) + ((!g2218) & (!g2436) & (g3138) & (!g3139) & (!g3153) & (!g3187)) + ((!g2218) & (!g2436) & (g3138) & (!g3139) & (!g3153) & (g3187)) + ((!g2218) & (!g2436) & (g3138) & (!g3139) & (g3153) & (!g3187)) + ((!g2218) & (!g2436) & (g3138) & (!g3139) & (g3153) & (g3187)) + ((!g2218) & (!g2436) & (g3138) & (g3139) & (!g3153) & (!g3187)) + ((!g2218) & (!g2436) & (g3138) & (g3139) & (!g3153) & (g3187)) + ((!g2218) & (!g2436) & (g3138) & (g3139) & (g3153) & (g3187)) + ((!g2218) & (g2436) & (!g3138) & (!g3139) & (g3153) & (!g3187)) + ((!g2218) & (g2436) & (!g3138) & (g3139) & (!g3153) & (!g3187)) + ((!g2218) & (g2436) & (!g3138) & (g3139) & (g3153) & (!g3187)) + ((!g2218) & (g2436) & (g3138) & (!g3139) & (!g3153) & (!g3187)) + ((!g2218) & (g2436) & (g3138) & (!g3139) & (!g3153) & (g3187)) + ((!g2218) & (g2436) & (g3138) & (!g3139) & (g3153) & (g3187)) + ((!g2218) & (g2436) & (g3138) & (g3139) & (!g3153) & (g3187)) + ((!g2218) & (g2436) & (g3138) & (g3139) & (g3153) & (g3187)) + ((g2218) & (!g2436) & (!g3138) & (!g3139) & (!g3153) & (!g3187)) + ((g2218) & (!g2436) & (!g3138) & (!g3139) & (g3153) & (!g3187)) + ((g2218) & (!g2436) & (!g3138) & (g3139) & (!g3153) & (!g3187)) + ((g2218) & (!g2436) & (g3138) & (!g3139) & (!g3153) & (g3187)) + ((g2218) & (!g2436) & (g3138) & (!g3139) & (g3153) & (g3187)) + ((g2218) & (!g2436) & (g3138) & (g3139) & (!g3153) & (g3187)) + ((g2218) & (!g2436) & (g3138) & (g3139) & (g3153) & (!g3187)) + ((g2218) & (!g2436) & (g3138) & (g3139) & (g3153) & (g3187)) + ((g2218) & (g2436) & (!g3138) & (!g3139) & (!g3153) & (!g3187)) + ((g2218) & (g2436) & (g3138) & (!g3139) & (!g3153) & (g3187)) + ((g2218) & (g2436) & (g3138) & (!g3139) & (g3153) & (!g3187)) + ((g2218) & (g2436) & (g3138) & (!g3139) & (g3153) & (g3187)) + ((g2218) & (g2436) & (g3138) & (g3139) & (!g3153) & (!g3187)) + ((g2218) & (g2436) & (g3138) & (g3139) & (!g3153) & (g3187)) + ((g2218) & (g2436) & (g3138) & (g3139) & (g3153) & (!g3187)) + ((g2218) & (g2436) & (g3138) & (g3139) & (g3153) & (g3187)));
	assign g3234 = (((!g2436) & (!g3139) & (g3153) & (!g3187)) + ((!g2436) & (g3139) & (!g3153) & (!g3187)) + ((!g2436) & (g3139) & (!g3153) & (g3187)) + ((!g2436) & (g3139) & (g3153) & (g3187)) + ((g2436) & (!g3139) & (!g3153) & (!g3187)) + ((g2436) & (g3139) & (!g3153) & (g3187)) + ((g2436) & (g3139) & (g3153) & (!g3187)) + ((g2436) & (g3139) & (g3153) & (g3187)));
	assign g3235 = (((!g2398) & (!g2627) & (!g3141) & (g3142) & (g3152) & (!g3187)) + ((!g2398) & (!g2627) & (g3141) & (!g3142) & (!g3152) & (!g3187)) + ((!g2398) & (!g2627) & (g3141) & (!g3142) & (!g3152) & (g3187)) + ((!g2398) & (!g2627) & (g3141) & (!g3142) & (g3152) & (!g3187)) + ((!g2398) & (!g2627) & (g3141) & (!g3142) & (g3152) & (g3187)) + ((!g2398) & (!g2627) & (g3141) & (g3142) & (!g3152) & (!g3187)) + ((!g2398) & (!g2627) & (g3141) & (g3142) & (!g3152) & (g3187)) + ((!g2398) & (!g2627) & (g3141) & (g3142) & (g3152) & (g3187)) + ((!g2398) & (g2627) & (!g3141) & (!g3142) & (g3152) & (!g3187)) + ((!g2398) & (g2627) & (!g3141) & (g3142) & (!g3152) & (!g3187)) + ((!g2398) & (g2627) & (!g3141) & (g3142) & (g3152) & (!g3187)) + ((!g2398) & (g2627) & (g3141) & (!g3142) & (!g3152) & (!g3187)) + ((!g2398) & (g2627) & (g3141) & (!g3142) & (!g3152) & (g3187)) + ((!g2398) & (g2627) & (g3141) & (!g3142) & (g3152) & (g3187)) + ((!g2398) & (g2627) & (g3141) & (g3142) & (!g3152) & (g3187)) + ((!g2398) & (g2627) & (g3141) & (g3142) & (g3152) & (g3187)) + ((g2398) & (!g2627) & (!g3141) & (!g3142) & (!g3152) & (!g3187)) + ((g2398) & (!g2627) & (!g3141) & (!g3142) & (g3152) & (!g3187)) + ((g2398) & (!g2627) & (!g3141) & (g3142) & (!g3152) & (!g3187)) + ((g2398) & (!g2627) & (g3141) & (!g3142) & (!g3152) & (g3187)) + ((g2398) & (!g2627) & (g3141) & (!g3142) & (g3152) & (g3187)) + ((g2398) & (!g2627) & (g3141) & (g3142) & (!g3152) & (g3187)) + ((g2398) & (!g2627) & (g3141) & (g3142) & (g3152) & (!g3187)) + ((g2398) & (!g2627) & (g3141) & (g3142) & (g3152) & (g3187)) + ((g2398) & (g2627) & (!g3141) & (!g3142) & (!g3152) & (!g3187)) + ((g2398) & (g2627) & (g3141) & (!g3142) & (!g3152) & (g3187)) + ((g2398) & (g2627) & (g3141) & (!g3142) & (g3152) & (!g3187)) + ((g2398) & (g2627) & (g3141) & (!g3142) & (g3152) & (g3187)) + ((g2398) & (g2627) & (g3141) & (g3142) & (!g3152) & (!g3187)) + ((g2398) & (g2627) & (g3141) & (g3142) & (!g3152) & (g3187)) + ((g2398) & (g2627) & (g3141) & (g3142) & (g3152) & (!g3187)) + ((g2398) & (g2627) & (g3141) & (g3142) & (g3152) & (g3187)));
	assign g3236 = (((!g2627) & (!g3142) & (g3152) & (!g3187)) + ((!g2627) & (g3142) & (!g3152) & (!g3187)) + ((!g2627) & (g3142) & (!g3152) & (g3187)) + ((!g2627) & (g3142) & (g3152) & (g3187)) + ((g2627) & (!g3142) & (!g3152) & (!g3187)) + ((g2627) & (g3142) & (!g3152) & (g3187)) + ((g2627) & (g3142) & (g3152) & (!g3187)) + ((g2627) & (g3142) & (g3152) & (g3187)));
	assign g3237 = (((!g2585) & (!g2825) & (!g3144) & (g3145) & (g3151) & (!g3187)) + ((!g2585) & (!g2825) & (g3144) & (!g3145) & (!g3151) & (!g3187)) + ((!g2585) & (!g2825) & (g3144) & (!g3145) & (!g3151) & (g3187)) + ((!g2585) & (!g2825) & (g3144) & (!g3145) & (g3151) & (!g3187)) + ((!g2585) & (!g2825) & (g3144) & (!g3145) & (g3151) & (g3187)) + ((!g2585) & (!g2825) & (g3144) & (g3145) & (!g3151) & (!g3187)) + ((!g2585) & (!g2825) & (g3144) & (g3145) & (!g3151) & (g3187)) + ((!g2585) & (!g2825) & (g3144) & (g3145) & (g3151) & (g3187)) + ((!g2585) & (g2825) & (!g3144) & (!g3145) & (g3151) & (!g3187)) + ((!g2585) & (g2825) & (!g3144) & (g3145) & (!g3151) & (!g3187)) + ((!g2585) & (g2825) & (!g3144) & (g3145) & (g3151) & (!g3187)) + ((!g2585) & (g2825) & (g3144) & (!g3145) & (!g3151) & (!g3187)) + ((!g2585) & (g2825) & (g3144) & (!g3145) & (!g3151) & (g3187)) + ((!g2585) & (g2825) & (g3144) & (!g3145) & (g3151) & (g3187)) + ((!g2585) & (g2825) & (g3144) & (g3145) & (!g3151) & (g3187)) + ((!g2585) & (g2825) & (g3144) & (g3145) & (g3151) & (g3187)) + ((g2585) & (!g2825) & (!g3144) & (!g3145) & (!g3151) & (!g3187)) + ((g2585) & (!g2825) & (!g3144) & (!g3145) & (g3151) & (!g3187)) + ((g2585) & (!g2825) & (!g3144) & (g3145) & (!g3151) & (!g3187)) + ((g2585) & (!g2825) & (g3144) & (!g3145) & (!g3151) & (g3187)) + ((g2585) & (!g2825) & (g3144) & (!g3145) & (g3151) & (g3187)) + ((g2585) & (!g2825) & (g3144) & (g3145) & (!g3151) & (g3187)) + ((g2585) & (!g2825) & (g3144) & (g3145) & (g3151) & (!g3187)) + ((g2585) & (!g2825) & (g3144) & (g3145) & (g3151) & (g3187)) + ((g2585) & (g2825) & (!g3144) & (!g3145) & (!g3151) & (!g3187)) + ((g2585) & (g2825) & (g3144) & (!g3145) & (!g3151) & (g3187)) + ((g2585) & (g2825) & (g3144) & (!g3145) & (g3151) & (!g3187)) + ((g2585) & (g2825) & (g3144) & (!g3145) & (g3151) & (g3187)) + ((g2585) & (g2825) & (g3144) & (g3145) & (!g3151) & (!g3187)) + ((g2585) & (g2825) & (g3144) & (g3145) & (!g3151) & (g3187)) + ((g2585) & (g2825) & (g3144) & (g3145) & (g3151) & (!g3187)) + ((g2585) & (g2825) & (g3144) & (g3145) & (g3151) & (g3187)));
	assign g3238 = (((!g2825) & (!g3145) & (g3151) & (!g3187)) + ((!g2825) & (g3145) & (!g3151) & (!g3187)) + ((!g2825) & (g3145) & (!g3151) & (g3187)) + ((!g2825) & (g3145) & (g3151) & (g3187)) + ((g2825) & (!g3145) & (!g3151) & (!g3187)) + ((g2825) & (g3145) & (!g3151) & (g3187)) + ((g2825) & (g3145) & (g3151) & (!g3187)) + ((g2825) & (g3145) & (g3151) & (g3187)));
	assign g3239 = (((!g2779) & (!g3030) & (!g3147) & (g3148) & (g3150) & (!g3187)) + ((!g2779) & (!g3030) & (g3147) & (!g3148) & (!g3150) & (!g3187)) + ((!g2779) & (!g3030) & (g3147) & (!g3148) & (!g3150) & (g3187)) + ((!g2779) & (!g3030) & (g3147) & (!g3148) & (g3150) & (!g3187)) + ((!g2779) & (!g3030) & (g3147) & (!g3148) & (g3150) & (g3187)) + ((!g2779) & (!g3030) & (g3147) & (g3148) & (!g3150) & (!g3187)) + ((!g2779) & (!g3030) & (g3147) & (g3148) & (!g3150) & (g3187)) + ((!g2779) & (!g3030) & (g3147) & (g3148) & (g3150) & (g3187)) + ((!g2779) & (g3030) & (!g3147) & (!g3148) & (g3150) & (!g3187)) + ((!g2779) & (g3030) & (!g3147) & (g3148) & (!g3150) & (!g3187)) + ((!g2779) & (g3030) & (!g3147) & (g3148) & (g3150) & (!g3187)) + ((!g2779) & (g3030) & (g3147) & (!g3148) & (!g3150) & (!g3187)) + ((!g2779) & (g3030) & (g3147) & (!g3148) & (!g3150) & (g3187)) + ((!g2779) & (g3030) & (g3147) & (!g3148) & (g3150) & (g3187)) + ((!g2779) & (g3030) & (g3147) & (g3148) & (!g3150) & (g3187)) + ((!g2779) & (g3030) & (g3147) & (g3148) & (g3150) & (g3187)) + ((g2779) & (!g3030) & (!g3147) & (!g3148) & (!g3150) & (!g3187)) + ((g2779) & (!g3030) & (!g3147) & (!g3148) & (g3150) & (!g3187)) + ((g2779) & (!g3030) & (!g3147) & (g3148) & (!g3150) & (!g3187)) + ((g2779) & (!g3030) & (g3147) & (!g3148) & (!g3150) & (g3187)) + ((g2779) & (!g3030) & (g3147) & (!g3148) & (g3150) & (g3187)) + ((g2779) & (!g3030) & (g3147) & (g3148) & (!g3150) & (g3187)) + ((g2779) & (!g3030) & (g3147) & (g3148) & (g3150) & (!g3187)) + ((g2779) & (!g3030) & (g3147) & (g3148) & (g3150) & (g3187)) + ((g2779) & (g3030) & (!g3147) & (!g3148) & (!g3150) & (!g3187)) + ((g2779) & (g3030) & (g3147) & (!g3148) & (!g3150) & (g3187)) + ((g2779) & (g3030) & (g3147) & (!g3148) & (g3150) & (!g3187)) + ((g2779) & (g3030) & (g3147) & (!g3148) & (g3150) & (g3187)) + ((g2779) & (g3030) & (g3147) & (g3148) & (!g3150) & (!g3187)) + ((g2779) & (g3030) & (g3147) & (g3148) & (!g3150) & (g3187)) + ((g2779) & (g3030) & (g3147) & (g3148) & (g3150) & (!g3187)) + ((g2779) & (g3030) & (g3147) & (g3148) & (g3150) & (g3187)));
	assign g3240 = (((!g3030) & (!g3148) & (g3150) & (!g3187)) + ((!g3030) & (g3148) & (!g3150) & (!g3187)) + ((!g3030) & (g3148) & (!g3150) & (g3187)) + ((!g3030) & (g3148) & (g3150) & (g3187)) + ((g3030) & (!g3148) & (!g3150) & (!g3187)) + ((g3030) & (g3148) & (!g3150) & (g3187)) + ((g3030) & (g3148) & (g3150) & (!g3187)) + ((g3030) & (g3148) & (g3150) & (g3187)));
	assign g3241 = (((!g2980) & (!ax10x) & (!ax11x) & (!g3178) & (!g3149) & (g3187)) + ((!g2980) & (!ax10x) & (!ax11x) & (!g3178) & (g3149) & (!g3187)) + ((!g2980) & (!ax10x) & (!ax11x) & (!g3178) & (g3149) & (g3187)) + ((!g2980) & (!ax10x) & (!ax11x) & (g3178) & (!g3149) & (!g3187)) + ((!g2980) & (!ax10x) & (ax11x) & (!g3178) & (!g3149) & (!g3187)) + ((!g2980) & (!ax10x) & (ax11x) & (g3178) & (!g3149) & (g3187)) + ((!g2980) & (!ax10x) & (ax11x) & (g3178) & (g3149) & (!g3187)) + ((!g2980) & (!ax10x) & (ax11x) & (g3178) & (g3149) & (g3187)) + ((!g2980) & (ax10x) & (!ax11x) & (g3178) & (!g3149) & (!g3187)) + ((!g2980) & (ax10x) & (!ax11x) & (g3178) & (g3149) & (!g3187)) + ((!g2980) & (ax10x) & (ax11x) & (!g3178) & (!g3149) & (!g3187)) + ((!g2980) & (ax10x) & (ax11x) & (!g3178) & (!g3149) & (g3187)) + ((!g2980) & (ax10x) & (ax11x) & (!g3178) & (g3149) & (!g3187)) + ((!g2980) & (ax10x) & (ax11x) & (!g3178) & (g3149) & (g3187)) + ((!g2980) & (ax10x) & (ax11x) & (g3178) & (!g3149) & (g3187)) + ((!g2980) & (ax10x) & (ax11x) & (g3178) & (g3149) & (g3187)) + ((g2980) & (!ax10x) & (!ax11x) & (!g3178) & (!g3149) & (!g3187)) + ((g2980) & (!ax10x) & (!ax11x) & (!g3178) & (!g3149) & (g3187)) + ((g2980) & (!ax10x) & (!ax11x) & (!g3178) & (g3149) & (g3187)) + ((g2980) & (!ax10x) & (!ax11x) & (g3178) & (g3149) & (!g3187)) + ((g2980) & (!ax10x) & (ax11x) & (!g3178) & (g3149) & (!g3187)) + ((g2980) & (!ax10x) & (ax11x) & (g3178) & (!g3149) & (!g3187)) + ((g2980) & (!ax10x) & (ax11x) & (g3178) & (!g3149) & (g3187)) + ((g2980) & (!ax10x) & (ax11x) & (g3178) & (g3149) & (g3187)) + ((g2980) & (ax10x) & (!ax11x) & (!g3178) & (!g3149) & (!g3187)) + ((g2980) & (ax10x) & (!ax11x) & (!g3178) & (g3149) & (!g3187)) + ((g2980) & (ax10x) & (ax11x) & (!g3178) & (!g3149) & (g3187)) + ((g2980) & (ax10x) & (ax11x) & (!g3178) & (g3149) & (g3187)) + ((g2980) & (ax10x) & (ax11x) & (g3178) & (!g3149) & (!g3187)) + ((g2980) & (ax10x) & (ax11x) & (g3178) & (!g3149) & (g3187)) + ((g2980) & (ax10x) & (ax11x) & (g3178) & (g3149) & (!g3187)) + ((g2980) & (ax10x) & (ax11x) & (g3178) & (g3149) & (g3187)));
	assign g3242 = (((!ax10x) & (!g3178) & (!g3149) & (g3187)) + ((!ax10x) & (!g3178) & (g3149) & (!g3187)) + ((!ax10x) & (!g3178) & (g3149) & (g3187)) + ((!ax10x) & (g3178) & (g3149) & (!g3187)) + ((ax10x) & (!g3178) & (!g3149) & (!g3187)) + ((ax10x) & (g3178) & (!g3149) & (!g3187)) + ((ax10x) & (g3178) & (!g3149) & (g3187)) + ((ax10x) & (g3178) & (g3149) & (g3187)));
	assign g3243 = (((!ax6x) & (!ax7x)));
	assign g3244 = (((!g3178) & (!ax8x) & (!ax9x) & (!g3187) & (!g3243)) + ((!g3178) & (!ax8x) & (ax9x) & (g3187) & (!g3243)) + ((!g3178) & (ax8x) & (ax9x) & (g3187) & (!g3243)) + ((!g3178) & (ax8x) & (ax9x) & (g3187) & (g3243)) + ((g3178) & (!ax8x) & (!ax9x) & (!g3187) & (!g3243)) + ((g3178) & (!ax8x) & (!ax9x) & (!g3187) & (g3243)) + ((g3178) & (!ax8x) & (!ax9x) & (g3187) & (!g3243)) + ((g3178) & (!ax8x) & (ax9x) & (!g3187) & (!g3243)) + ((g3178) & (!ax8x) & (ax9x) & (g3187) & (!g3243)) + ((g3178) & (!ax8x) & (ax9x) & (g3187) & (g3243)) + ((g3178) & (ax8x) & (!ax9x) & (g3187) & (!g3243)) + ((g3178) & (ax8x) & (!ax9x) & (g3187) & (g3243)) + ((g3178) & (ax8x) & (ax9x) & (!g3187) & (!g3243)) + ((g3178) & (ax8x) & (ax9x) & (!g3187) & (g3243)) + ((g3178) & (ax8x) & (ax9x) & (g3187) & (!g3243)) + ((g3178) & (ax8x) & (ax9x) & (g3187) & (g3243)));
	assign g3245 = (((!g3030) & (!g2980) & (g3241) & (g3242) & (g3244)) + ((!g3030) & (g2980) & (g3241) & (!g3242) & (g3244)) + ((!g3030) & (g2980) & (g3241) & (g3242) & (!g3244)) + ((!g3030) & (g2980) & (g3241) & (g3242) & (g3244)) + ((g3030) & (!g2980) & (!g3241) & (g3242) & (g3244)) + ((g3030) & (!g2980) & (g3241) & (!g3242) & (!g3244)) + ((g3030) & (!g2980) & (g3241) & (!g3242) & (g3244)) + ((g3030) & (!g2980) & (g3241) & (g3242) & (!g3244)) + ((g3030) & (!g2980) & (g3241) & (g3242) & (g3244)) + ((g3030) & (g2980) & (!g3241) & (!g3242) & (g3244)) + ((g3030) & (g2980) & (!g3241) & (g3242) & (!g3244)) + ((g3030) & (g2980) & (!g3241) & (g3242) & (g3244)) + ((g3030) & (g2980) & (g3241) & (!g3242) & (!g3244)) + ((g3030) & (g2980) & (g3241) & (!g3242) & (g3244)) + ((g3030) & (g2980) & (g3241) & (g3242) & (!g3244)) + ((g3030) & (g2980) & (g3241) & (g3242) & (g3244)));
	assign g3246 = (((!g2825) & (!g2779) & (g3239) & (g3240) & (g3245)) + ((!g2825) & (g2779) & (g3239) & (!g3240) & (g3245)) + ((!g2825) & (g2779) & (g3239) & (g3240) & (!g3245)) + ((!g2825) & (g2779) & (g3239) & (g3240) & (g3245)) + ((g2825) & (!g2779) & (!g3239) & (g3240) & (g3245)) + ((g2825) & (!g2779) & (g3239) & (!g3240) & (!g3245)) + ((g2825) & (!g2779) & (g3239) & (!g3240) & (g3245)) + ((g2825) & (!g2779) & (g3239) & (g3240) & (!g3245)) + ((g2825) & (!g2779) & (g3239) & (g3240) & (g3245)) + ((g2825) & (g2779) & (!g3239) & (!g3240) & (g3245)) + ((g2825) & (g2779) & (!g3239) & (g3240) & (!g3245)) + ((g2825) & (g2779) & (!g3239) & (g3240) & (g3245)) + ((g2825) & (g2779) & (g3239) & (!g3240) & (!g3245)) + ((g2825) & (g2779) & (g3239) & (!g3240) & (g3245)) + ((g2825) & (g2779) & (g3239) & (g3240) & (!g3245)) + ((g2825) & (g2779) & (g3239) & (g3240) & (g3245)));
	assign g3247 = (((!g2627) & (!g2585) & (g3237) & (g3238) & (g3246)) + ((!g2627) & (g2585) & (g3237) & (!g3238) & (g3246)) + ((!g2627) & (g2585) & (g3237) & (g3238) & (!g3246)) + ((!g2627) & (g2585) & (g3237) & (g3238) & (g3246)) + ((g2627) & (!g2585) & (!g3237) & (g3238) & (g3246)) + ((g2627) & (!g2585) & (g3237) & (!g3238) & (!g3246)) + ((g2627) & (!g2585) & (g3237) & (!g3238) & (g3246)) + ((g2627) & (!g2585) & (g3237) & (g3238) & (!g3246)) + ((g2627) & (!g2585) & (g3237) & (g3238) & (g3246)) + ((g2627) & (g2585) & (!g3237) & (!g3238) & (g3246)) + ((g2627) & (g2585) & (!g3237) & (g3238) & (!g3246)) + ((g2627) & (g2585) & (!g3237) & (g3238) & (g3246)) + ((g2627) & (g2585) & (g3237) & (!g3238) & (!g3246)) + ((g2627) & (g2585) & (g3237) & (!g3238) & (g3246)) + ((g2627) & (g2585) & (g3237) & (g3238) & (!g3246)) + ((g2627) & (g2585) & (g3237) & (g3238) & (g3246)));
	assign g3248 = (((!g2436) & (!g2398) & (g3235) & (g3236) & (g3247)) + ((!g2436) & (g2398) & (g3235) & (!g3236) & (g3247)) + ((!g2436) & (g2398) & (g3235) & (g3236) & (!g3247)) + ((!g2436) & (g2398) & (g3235) & (g3236) & (g3247)) + ((g2436) & (!g2398) & (!g3235) & (g3236) & (g3247)) + ((g2436) & (!g2398) & (g3235) & (!g3236) & (!g3247)) + ((g2436) & (!g2398) & (g3235) & (!g3236) & (g3247)) + ((g2436) & (!g2398) & (g3235) & (g3236) & (!g3247)) + ((g2436) & (!g2398) & (g3235) & (g3236) & (g3247)) + ((g2436) & (g2398) & (!g3235) & (!g3236) & (g3247)) + ((g2436) & (g2398) & (!g3235) & (g3236) & (!g3247)) + ((g2436) & (g2398) & (!g3235) & (g3236) & (g3247)) + ((g2436) & (g2398) & (g3235) & (!g3236) & (!g3247)) + ((g2436) & (g2398) & (g3235) & (!g3236) & (g3247)) + ((g2436) & (g2398) & (g3235) & (g3236) & (!g3247)) + ((g2436) & (g2398) & (g3235) & (g3236) & (g3247)));
	assign g3249 = (((!g2252) & (!g2218) & (g3233) & (g3234) & (g3248)) + ((!g2252) & (g2218) & (g3233) & (!g3234) & (g3248)) + ((!g2252) & (g2218) & (g3233) & (g3234) & (!g3248)) + ((!g2252) & (g2218) & (g3233) & (g3234) & (g3248)) + ((g2252) & (!g2218) & (!g3233) & (g3234) & (g3248)) + ((g2252) & (!g2218) & (g3233) & (!g3234) & (!g3248)) + ((g2252) & (!g2218) & (g3233) & (!g3234) & (g3248)) + ((g2252) & (!g2218) & (g3233) & (g3234) & (!g3248)) + ((g2252) & (!g2218) & (g3233) & (g3234) & (g3248)) + ((g2252) & (g2218) & (!g3233) & (!g3234) & (g3248)) + ((g2252) & (g2218) & (!g3233) & (g3234) & (!g3248)) + ((g2252) & (g2218) & (!g3233) & (g3234) & (g3248)) + ((g2252) & (g2218) & (g3233) & (!g3234) & (!g3248)) + ((g2252) & (g2218) & (g3233) & (!g3234) & (g3248)) + ((g2252) & (g2218) & (g3233) & (g3234) & (!g3248)) + ((g2252) & (g2218) & (g3233) & (g3234) & (g3248)));
	assign g3250 = (((!g2075) & (!g2045) & (g3231) & (g3232) & (g3249)) + ((!g2075) & (g2045) & (g3231) & (!g3232) & (g3249)) + ((!g2075) & (g2045) & (g3231) & (g3232) & (!g3249)) + ((!g2075) & (g2045) & (g3231) & (g3232) & (g3249)) + ((g2075) & (!g2045) & (!g3231) & (g3232) & (g3249)) + ((g2075) & (!g2045) & (g3231) & (!g3232) & (!g3249)) + ((g2075) & (!g2045) & (g3231) & (!g3232) & (g3249)) + ((g2075) & (!g2045) & (g3231) & (g3232) & (!g3249)) + ((g2075) & (!g2045) & (g3231) & (g3232) & (g3249)) + ((g2075) & (g2045) & (!g3231) & (!g3232) & (g3249)) + ((g2075) & (g2045) & (!g3231) & (g3232) & (!g3249)) + ((g2075) & (g2045) & (!g3231) & (g3232) & (g3249)) + ((g2075) & (g2045) & (g3231) & (!g3232) & (!g3249)) + ((g2075) & (g2045) & (g3231) & (!g3232) & (g3249)) + ((g2075) & (g2045) & (g3231) & (g3232) & (!g3249)) + ((g2075) & (g2045) & (g3231) & (g3232) & (g3249)));
	assign g3251 = (((!g1905) & (!g1879) & (g3229) & (g3230) & (g3250)) + ((!g1905) & (g1879) & (g3229) & (!g3230) & (g3250)) + ((!g1905) & (g1879) & (g3229) & (g3230) & (!g3250)) + ((!g1905) & (g1879) & (g3229) & (g3230) & (g3250)) + ((g1905) & (!g1879) & (!g3229) & (g3230) & (g3250)) + ((g1905) & (!g1879) & (g3229) & (!g3230) & (!g3250)) + ((g1905) & (!g1879) & (g3229) & (!g3230) & (g3250)) + ((g1905) & (!g1879) & (g3229) & (g3230) & (!g3250)) + ((g1905) & (!g1879) & (g3229) & (g3230) & (g3250)) + ((g1905) & (g1879) & (!g3229) & (!g3230) & (g3250)) + ((g1905) & (g1879) & (!g3229) & (g3230) & (!g3250)) + ((g1905) & (g1879) & (!g3229) & (g3230) & (g3250)) + ((g1905) & (g1879) & (g3229) & (!g3230) & (!g3250)) + ((g1905) & (g1879) & (g3229) & (!g3230) & (g3250)) + ((g1905) & (g1879) & (g3229) & (g3230) & (!g3250)) + ((g1905) & (g1879) & (g3229) & (g3230) & (g3250)));
	assign g3252 = (((!g1742) & (!g1720) & (g3227) & (g3228) & (g3251)) + ((!g1742) & (g1720) & (g3227) & (!g3228) & (g3251)) + ((!g1742) & (g1720) & (g3227) & (g3228) & (!g3251)) + ((!g1742) & (g1720) & (g3227) & (g3228) & (g3251)) + ((g1742) & (!g1720) & (!g3227) & (g3228) & (g3251)) + ((g1742) & (!g1720) & (g3227) & (!g3228) & (!g3251)) + ((g1742) & (!g1720) & (g3227) & (!g3228) & (g3251)) + ((g1742) & (!g1720) & (g3227) & (g3228) & (!g3251)) + ((g1742) & (!g1720) & (g3227) & (g3228) & (g3251)) + ((g1742) & (g1720) & (!g3227) & (!g3228) & (g3251)) + ((g1742) & (g1720) & (!g3227) & (g3228) & (!g3251)) + ((g1742) & (g1720) & (!g3227) & (g3228) & (g3251)) + ((g1742) & (g1720) & (g3227) & (!g3228) & (!g3251)) + ((g1742) & (g1720) & (g3227) & (!g3228) & (g3251)) + ((g1742) & (g1720) & (g3227) & (g3228) & (!g3251)) + ((g1742) & (g1720) & (g3227) & (g3228) & (g3251)));
	assign g3253 = (((!g1586) & (!g1568) & (g3225) & (g3226) & (g3252)) + ((!g1586) & (g1568) & (g3225) & (!g3226) & (g3252)) + ((!g1586) & (g1568) & (g3225) & (g3226) & (!g3252)) + ((!g1586) & (g1568) & (g3225) & (g3226) & (g3252)) + ((g1586) & (!g1568) & (!g3225) & (g3226) & (g3252)) + ((g1586) & (!g1568) & (g3225) & (!g3226) & (!g3252)) + ((g1586) & (!g1568) & (g3225) & (!g3226) & (g3252)) + ((g1586) & (!g1568) & (g3225) & (g3226) & (!g3252)) + ((g1586) & (!g1568) & (g3225) & (g3226) & (g3252)) + ((g1586) & (g1568) & (!g3225) & (!g3226) & (g3252)) + ((g1586) & (g1568) & (!g3225) & (g3226) & (!g3252)) + ((g1586) & (g1568) & (!g3225) & (g3226) & (g3252)) + ((g1586) & (g1568) & (g3225) & (!g3226) & (!g3252)) + ((g1586) & (g1568) & (g3225) & (!g3226) & (g3252)) + ((g1586) & (g1568) & (g3225) & (g3226) & (!g3252)) + ((g1586) & (g1568) & (g3225) & (g3226) & (g3252)));
	assign g3254 = (((!g1437) & (!g1423) & (g3223) & (g3224) & (g3253)) + ((!g1437) & (g1423) & (g3223) & (!g3224) & (g3253)) + ((!g1437) & (g1423) & (g3223) & (g3224) & (!g3253)) + ((!g1437) & (g1423) & (g3223) & (g3224) & (g3253)) + ((g1437) & (!g1423) & (!g3223) & (g3224) & (g3253)) + ((g1437) & (!g1423) & (g3223) & (!g3224) & (!g3253)) + ((g1437) & (!g1423) & (g3223) & (!g3224) & (g3253)) + ((g1437) & (!g1423) & (g3223) & (g3224) & (!g3253)) + ((g1437) & (!g1423) & (g3223) & (g3224) & (g3253)) + ((g1437) & (g1423) & (!g3223) & (!g3224) & (g3253)) + ((g1437) & (g1423) & (!g3223) & (g3224) & (!g3253)) + ((g1437) & (g1423) & (!g3223) & (g3224) & (g3253)) + ((g1437) & (g1423) & (g3223) & (!g3224) & (!g3253)) + ((g1437) & (g1423) & (g3223) & (!g3224) & (g3253)) + ((g1437) & (g1423) & (g3223) & (g3224) & (!g3253)) + ((g1437) & (g1423) & (g3223) & (g3224) & (g3253)));
	assign g3255 = (((!g1295) & (!g1285) & (g3221) & (g3222) & (g3254)) + ((!g1295) & (g1285) & (g3221) & (!g3222) & (g3254)) + ((!g1295) & (g1285) & (g3221) & (g3222) & (!g3254)) + ((!g1295) & (g1285) & (g3221) & (g3222) & (g3254)) + ((g1295) & (!g1285) & (!g3221) & (g3222) & (g3254)) + ((g1295) & (!g1285) & (g3221) & (!g3222) & (!g3254)) + ((g1295) & (!g1285) & (g3221) & (!g3222) & (g3254)) + ((g1295) & (!g1285) & (g3221) & (g3222) & (!g3254)) + ((g1295) & (!g1285) & (g3221) & (g3222) & (g3254)) + ((g1295) & (g1285) & (!g3221) & (!g3222) & (g3254)) + ((g1295) & (g1285) & (!g3221) & (g3222) & (!g3254)) + ((g1295) & (g1285) & (!g3221) & (g3222) & (g3254)) + ((g1295) & (g1285) & (g3221) & (!g3222) & (!g3254)) + ((g1295) & (g1285) & (g3221) & (!g3222) & (g3254)) + ((g1295) & (g1285) & (g3221) & (g3222) & (!g3254)) + ((g1295) & (g1285) & (g3221) & (g3222) & (g3254)));
	assign g3256 = (((!g1160) & (!g1154) & (g3219) & (g3220) & (g3255)) + ((!g1160) & (g1154) & (g3219) & (!g3220) & (g3255)) + ((!g1160) & (g1154) & (g3219) & (g3220) & (!g3255)) + ((!g1160) & (g1154) & (g3219) & (g3220) & (g3255)) + ((g1160) & (!g1154) & (!g3219) & (g3220) & (g3255)) + ((g1160) & (!g1154) & (g3219) & (!g3220) & (!g3255)) + ((g1160) & (!g1154) & (g3219) & (!g3220) & (g3255)) + ((g1160) & (!g1154) & (g3219) & (g3220) & (!g3255)) + ((g1160) & (!g1154) & (g3219) & (g3220) & (g3255)) + ((g1160) & (g1154) & (!g3219) & (!g3220) & (g3255)) + ((g1160) & (g1154) & (!g3219) & (g3220) & (!g3255)) + ((g1160) & (g1154) & (!g3219) & (g3220) & (g3255)) + ((g1160) & (g1154) & (g3219) & (!g3220) & (!g3255)) + ((g1160) & (g1154) & (g3219) & (!g3220) & (g3255)) + ((g1160) & (g1154) & (g3219) & (g3220) & (!g3255)) + ((g1160) & (g1154) & (g3219) & (g3220) & (g3255)));
	assign g3257 = (((!g1032) & (!g1030) & (g3217) & (g3218) & (g3256)) + ((!g1032) & (g1030) & (g3217) & (!g3218) & (g3256)) + ((!g1032) & (g1030) & (g3217) & (g3218) & (!g3256)) + ((!g1032) & (g1030) & (g3217) & (g3218) & (g3256)) + ((g1032) & (!g1030) & (!g3217) & (g3218) & (g3256)) + ((g1032) & (!g1030) & (g3217) & (!g3218) & (!g3256)) + ((g1032) & (!g1030) & (g3217) & (!g3218) & (g3256)) + ((g1032) & (!g1030) & (g3217) & (g3218) & (!g3256)) + ((g1032) & (!g1030) & (g3217) & (g3218) & (g3256)) + ((g1032) & (g1030) & (!g3217) & (!g3218) & (g3256)) + ((g1032) & (g1030) & (!g3217) & (g3218) & (!g3256)) + ((g1032) & (g1030) & (!g3217) & (g3218) & (g3256)) + ((g1032) & (g1030) & (g3217) & (!g3218) & (!g3256)) + ((g1032) & (g1030) & (g3217) & (!g3218) & (g3256)) + ((g1032) & (g1030) & (g3217) & (g3218) & (!g3256)) + ((g1032) & (g1030) & (g3217) & (g3218) & (g3256)));
	assign g3258 = (((!g851) & (!g914) & (g3215) & (g3216) & (g3257)) + ((!g851) & (g914) & (g3215) & (!g3216) & (g3257)) + ((!g851) & (g914) & (g3215) & (g3216) & (!g3257)) + ((!g851) & (g914) & (g3215) & (g3216) & (g3257)) + ((g851) & (!g914) & (!g3215) & (g3216) & (g3257)) + ((g851) & (!g914) & (g3215) & (!g3216) & (!g3257)) + ((g851) & (!g914) & (g3215) & (!g3216) & (g3257)) + ((g851) & (!g914) & (g3215) & (g3216) & (!g3257)) + ((g851) & (!g914) & (g3215) & (g3216) & (g3257)) + ((g851) & (g914) & (!g3215) & (!g3216) & (g3257)) + ((g851) & (g914) & (!g3215) & (g3216) & (!g3257)) + ((g851) & (g914) & (!g3215) & (g3216) & (g3257)) + ((g851) & (g914) & (g3215) & (!g3216) & (!g3257)) + ((g851) & (g914) & (g3215) & (!g3216) & (g3257)) + ((g851) & (g914) & (g3215) & (g3216) & (!g3257)) + ((g851) & (g914) & (g3215) & (g3216) & (g3257)));
	assign g3259 = (((!g744) & (!g803) & (g3213) & (g3214) & (g3258)) + ((!g744) & (g803) & (g3213) & (!g3214) & (g3258)) + ((!g744) & (g803) & (g3213) & (g3214) & (!g3258)) + ((!g744) & (g803) & (g3213) & (g3214) & (g3258)) + ((g744) & (!g803) & (!g3213) & (g3214) & (g3258)) + ((g744) & (!g803) & (g3213) & (!g3214) & (!g3258)) + ((g744) & (!g803) & (g3213) & (!g3214) & (g3258)) + ((g744) & (!g803) & (g3213) & (g3214) & (!g3258)) + ((g744) & (!g803) & (g3213) & (g3214) & (g3258)) + ((g744) & (g803) & (!g3213) & (!g3214) & (g3258)) + ((g744) & (g803) & (!g3213) & (g3214) & (!g3258)) + ((g744) & (g803) & (!g3213) & (g3214) & (g3258)) + ((g744) & (g803) & (g3213) & (!g3214) & (!g3258)) + ((g744) & (g803) & (g3213) & (!g3214) & (g3258)) + ((g744) & (g803) & (g3213) & (g3214) & (!g3258)) + ((g744) & (g803) & (g3213) & (g3214) & (g3258)));
	assign g3260 = (((!g645) & (!g700) & (g3211) & (g3212) & (g3259)) + ((!g645) & (g700) & (g3211) & (!g3212) & (g3259)) + ((!g645) & (g700) & (g3211) & (g3212) & (!g3259)) + ((!g645) & (g700) & (g3211) & (g3212) & (g3259)) + ((g645) & (!g700) & (!g3211) & (g3212) & (g3259)) + ((g645) & (!g700) & (g3211) & (!g3212) & (!g3259)) + ((g645) & (!g700) & (g3211) & (!g3212) & (g3259)) + ((g645) & (!g700) & (g3211) & (g3212) & (!g3259)) + ((g645) & (!g700) & (g3211) & (g3212) & (g3259)) + ((g645) & (g700) & (!g3211) & (!g3212) & (g3259)) + ((g645) & (g700) & (!g3211) & (g3212) & (!g3259)) + ((g645) & (g700) & (!g3211) & (g3212) & (g3259)) + ((g645) & (g700) & (g3211) & (!g3212) & (!g3259)) + ((g645) & (g700) & (g3211) & (!g3212) & (g3259)) + ((g645) & (g700) & (g3211) & (g3212) & (!g3259)) + ((g645) & (g700) & (g3211) & (g3212) & (g3259)));
	assign g3261 = (((!g553) & (!g604) & (g3209) & (g3210) & (g3260)) + ((!g553) & (g604) & (g3209) & (!g3210) & (g3260)) + ((!g553) & (g604) & (g3209) & (g3210) & (!g3260)) + ((!g553) & (g604) & (g3209) & (g3210) & (g3260)) + ((g553) & (!g604) & (!g3209) & (g3210) & (g3260)) + ((g553) & (!g604) & (g3209) & (!g3210) & (!g3260)) + ((g553) & (!g604) & (g3209) & (!g3210) & (g3260)) + ((g553) & (!g604) & (g3209) & (g3210) & (!g3260)) + ((g553) & (!g604) & (g3209) & (g3210) & (g3260)) + ((g553) & (g604) & (!g3209) & (!g3210) & (g3260)) + ((g553) & (g604) & (!g3209) & (g3210) & (!g3260)) + ((g553) & (g604) & (!g3209) & (g3210) & (g3260)) + ((g553) & (g604) & (g3209) & (!g3210) & (!g3260)) + ((g553) & (g604) & (g3209) & (!g3210) & (g3260)) + ((g553) & (g604) & (g3209) & (g3210) & (!g3260)) + ((g553) & (g604) & (g3209) & (g3210) & (g3260)));
	assign g3262 = (((!g468) & (!g515) & (g3207) & (g3208) & (g3261)) + ((!g468) & (g515) & (g3207) & (!g3208) & (g3261)) + ((!g468) & (g515) & (g3207) & (g3208) & (!g3261)) + ((!g468) & (g515) & (g3207) & (g3208) & (g3261)) + ((g468) & (!g515) & (!g3207) & (g3208) & (g3261)) + ((g468) & (!g515) & (g3207) & (!g3208) & (!g3261)) + ((g468) & (!g515) & (g3207) & (!g3208) & (g3261)) + ((g468) & (!g515) & (g3207) & (g3208) & (!g3261)) + ((g468) & (!g515) & (g3207) & (g3208) & (g3261)) + ((g468) & (g515) & (!g3207) & (!g3208) & (g3261)) + ((g468) & (g515) & (!g3207) & (g3208) & (!g3261)) + ((g468) & (g515) & (!g3207) & (g3208) & (g3261)) + ((g468) & (g515) & (g3207) & (!g3208) & (!g3261)) + ((g468) & (g515) & (g3207) & (!g3208) & (g3261)) + ((g468) & (g515) & (g3207) & (g3208) & (!g3261)) + ((g468) & (g515) & (g3207) & (g3208) & (g3261)));
	assign g3263 = (((!g390) & (!g433) & (g3205) & (g3206) & (g3262)) + ((!g390) & (g433) & (g3205) & (!g3206) & (g3262)) + ((!g390) & (g433) & (g3205) & (g3206) & (!g3262)) + ((!g390) & (g433) & (g3205) & (g3206) & (g3262)) + ((g390) & (!g433) & (!g3205) & (g3206) & (g3262)) + ((g390) & (!g433) & (g3205) & (!g3206) & (!g3262)) + ((g390) & (!g433) & (g3205) & (!g3206) & (g3262)) + ((g390) & (!g433) & (g3205) & (g3206) & (!g3262)) + ((g390) & (!g433) & (g3205) & (g3206) & (g3262)) + ((g390) & (g433) & (!g3205) & (!g3206) & (g3262)) + ((g390) & (g433) & (!g3205) & (g3206) & (!g3262)) + ((g390) & (g433) & (!g3205) & (g3206) & (g3262)) + ((g390) & (g433) & (g3205) & (!g3206) & (!g3262)) + ((g390) & (g433) & (g3205) & (!g3206) & (g3262)) + ((g390) & (g433) & (g3205) & (g3206) & (!g3262)) + ((g390) & (g433) & (g3205) & (g3206) & (g3262)));
	assign g3264 = (((!g319) & (!g358) & (g3203) & (g3204) & (g3263)) + ((!g319) & (g358) & (g3203) & (!g3204) & (g3263)) + ((!g319) & (g358) & (g3203) & (g3204) & (!g3263)) + ((!g319) & (g358) & (g3203) & (g3204) & (g3263)) + ((g319) & (!g358) & (!g3203) & (g3204) & (g3263)) + ((g319) & (!g358) & (g3203) & (!g3204) & (!g3263)) + ((g319) & (!g358) & (g3203) & (!g3204) & (g3263)) + ((g319) & (!g358) & (g3203) & (g3204) & (!g3263)) + ((g319) & (!g358) & (g3203) & (g3204) & (g3263)) + ((g319) & (g358) & (!g3203) & (!g3204) & (g3263)) + ((g319) & (g358) & (!g3203) & (g3204) & (!g3263)) + ((g319) & (g358) & (!g3203) & (g3204) & (g3263)) + ((g319) & (g358) & (g3203) & (!g3204) & (!g3263)) + ((g319) & (g358) & (g3203) & (!g3204) & (g3263)) + ((g319) & (g358) & (g3203) & (g3204) & (!g3263)) + ((g319) & (g358) & (g3203) & (g3204) & (g3263)));
	assign g3265 = (((!g255) & (!g290) & (g3201) & (g3202) & (g3264)) + ((!g255) & (g290) & (g3201) & (!g3202) & (g3264)) + ((!g255) & (g290) & (g3201) & (g3202) & (!g3264)) + ((!g255) & (g290) & (g3201) & (g3202) & (g3264)) + ((g255) & (!g290) & (!g3201) & (g3202) & (g3264)) + ((g255) & (!g290) & (g3201) & (!g3202) & (!g3264)) + ((g255) & (!g290) & (g3201) & (!g3202) & (g3264)) + ((g255) & (!g290) & (g3201) & (g3202) & (!g3264)) + ((g255) & (!g290) & (g3201) & (g3202) & (g3264)) + ((g255) & (g290) & (!g3201) & (!g3202) & (g3264)) + ((g255) & (g290) & (!g3201) & (g3202) & (!g3264)) + ((g255) & (g290) & (!g3201) & (g3202) & (g3264)) + ((g255) & (g290) & (g3201) & (!g3202) & (!g3264)) + ((g255) & (g290) & (g3201) & (!g3202) & (g3264)) + ((g255) & (g290) & (g3201) & (g3202) & (!g3264)) + ((g255) & (g290) & (g3201) & (g3202) & (g3264)));
	assign g3266 = (((!g198) & (!g229) & (g3199) & (g3200) & (g3265)) + ((!g198) & (g229) & (g3199) & (!g3200) & (g3265)) + ((!g198) & (g229) & (g3199) & (g3200) & (!g3265)) + ((!g198) & (g229) & (g3199) & (g3200) & (g3265)) + ((g198) & (!g229) & (!g3199) & (g3200) & (g3265)) + ((g198) & (!g229) & (g3199) & (!g3200) & (!g3265)) + ((g198) & (!g229) & (g3199) & (!g3200) & (g3265)) + ((g198) & (!g229) & (g3199) & (g3200) & (!g3265)) + ((g198) & (!g229) & (g3199) & (g3200) & (g3265)) + ((g198) & (g229) & (!g3199) & (!g3200) & (g3265)) + ((g198) & (g229) & (!g3199) & (g3200) & (!g3265)) + ((g198) & (g229) & (!g3199) & (g3200) & (g3265)) + ((g198) & (g229) & (g3199) & (!g3200) & (!g3265)) + ((g198) & (g229) & (g3199) & (!g3200) & (g3265)) + ((g198) & (g229) & (g3199) & (g3200) & (!g3265)) + ((g198) & (g229) & (g3199) & (g3200) & (g3265)));
	assign g3267 = (((!g147) & (!g174) & (g3197) & (g3198) & (g3266)) + ((!g147) & (g174) & (g3197) & (!g3198) & (g3266)) + ((!g147) & (g174) & (g3197) & (g3198) & (!g3266)) + ((!g147) & (g174) & (g3197) & (g3198) & (g3266)) + ((g147) & (!g174) & (!g3197) & (g3198) & (g3266)) + ((g147) & (!g174) & (g3197) & (!g3198) & (!g3266)) + ((g147) & (!g174) & (g3197) & (!g3198) & (g3266)) + ((g147) & (!g174) & (g3197) & (g3198) & (!g3266)) + ((g147) & (!g174) & (g3197) & (g3198) & (g3266)) + ((g147) & (g174) & (!g3197) & (!g3198) & (g3266)) + ((g147) & (g174) & (!g3197) & (g3198) & (!g3266)) + ((g147) & (g174) & (!g3197) & (g3198) & (g3266)) + ((g147) & (g174) & (g3197) & (!g3198) & (!g3266)) + ((g147) & (g174) & (g3197) & (!g3198) & (g3266)) + ((g147) & (g174) & (g3197) & (g3198) & (!g3266)) + ((g147) & (g174) & (g3197) & (g3198) & (g3266)));
	assign g3268 = (((!g104) & (!g127) & (g3195) & (g3196) & (g3267)) + ((!g104) & (g127) & (g3195) & (!g3196) & (g3267)) + ((!g104) & (g127) & (g3195) & (g3196) & (!g3267)) + ((!g104) & (g127) & (g3195) & (g3196) & (g3267)) + ((g104) & (!g127) & (!g3195) & (g3196) & (g3267)) + ((g104) & (!g127) & (g3195) & (!g3196) & (!g3267)) + ((g104) & (!g127) & (g3195) & (!g3196) & (g3267)) + ((g104) & (!g127) & (g3195) & (g3196) & (!g3267)) + ((g104) & (!g127) & (g3195) & (g3196) & (g3267)) + ((g104) & (g127) & (!g3195) & (!g3196) & (g3267)) + ((g104) & (g127) & (!g3195) & (g3196) & (!g3267)) + ((g104) & (g127) & (!g3195) & (g3196) & (g3267)) + ((g104) & (g127) & (g3195) & (!g3196) & (!g3267)) + ((g104) & (g127) & (g3195) & (!g3196) & (g3267)) + ((g104) & (g127) & (g3195) & (g3196) & (!g3267)) + ((g104) & (g127) & (g3195) & (g3196) & (g3267)));
	assign g3269 = (((!g68) & (!g87) & (g3193) & (g3194) & (g3268)) + ((!g68) & (g87) & (g3193) & (!g3194) & (g3268)) + ((!g68) & (g87) & (g3193) & (g3194) & (!g3268)) + ((!g68) & (g87) & (g3193) & (g3194) & (g3268)) + ((g68) & (!g87) & (!g3193) & (g3194) & (g3268)) + ((g68) & (!g87) & (g3193) & (!g3194) & (!g3268)) + ((g68) & (!g87) & (g3193) & (!g3194) & (g3268)) + ((g68) & (!g87) & (g3193) & (g3194) & (!g3268)) + ((g68) & (!g87) & (g3193) & (g3194) & (g3268)) + ((g68) & (g87) & (!g3193) & (!g3194) & (g3268)) + ((g68) & (g87) & (!g3193) & (g3194) & (!g3268)) + ((g68) & (g87) & (!g3193) & (g3194) & (g3268)) + ((g68) & (g87) & (g3193) & (!g3194) & (!g3268)) + ((g68) & (g87) & (g3193) & (!g3194) & (g3268)) + ((g68) & (g87) & (g3193) & (g3194) & (!g3268)) + ((g68) & (g87) & (g3193) & (g3194) & (g3268)));
	assign g3270 = (((!g39) & (!g54) & (g3191) & (g3192) & (g3269)) + ((!g39) & (g54) & (g3191) & (!g3192) & (g3269)) + ((!g39) & (g54) & (g3191) & (g3192) & (!g3269)) + ((!g39) & (g54) & (g3191) & (g3192) & (g3269)) + ((g39) & (!g54) & (!g3191) & (g3192) & (g3269)) + ((g39) & (!g54) & (g3191) & (!g3192) & (!g3269)) + ((g39) & (!g54) & (g3191) & (!g3192) & (g3269)) + ((g39) & (!g54) & (g3191) & (g3192) & (!g3269)) + ((g39) & (!g54) & (g3191) & (g3192) & (g3269)) + ((g39) & (g54) & (!g3191) & (!g3192) & (g3269)) + ((g39) & (g54) & (!g3191) & (g3192) & (!g3269)) + ((g39) & (g54) & (!g3191) & (g3192) & (g3269)) + ((g39) & (g54) & (g3191) & (!g3192) & (!g3269)) + ((g39) & (g54) & (g3191) & (!g3192) & (g3269)) + ((g39) & (g54) & (g3191) & (g3192) & (!g3269)) + ((g39) & (g54) & (g3191) & (g3192) & (g3269)));
	assign g3271 = (((!g18) & (!g27) & (g3189) & (g3190) & (g3270)) + ((!g18) & (g27) & (g3189) & (!g3190) & (g3270)) + ((!g18) & (g27) & (g3189) & (g3190) & (!g3270)) + ((!g18) & (g27) & (g3189) & (g3190) & (g3270)) + ((g18) & (!g27) & (!g3189) & (g3190) & (g3270)) + ((g18) & (!g27) & (g3189) & (!g3190) & (!g3270)) + ((g18) & (!g27) & (g3189) & (!g3190) & (g3270)) + ((g18) & (!g27) & (g3189) & (g3190) & (!g3270)) + ((g18) & (!g27) & (g3189) & (g3190) & (g3270)) + ((g18) & (g27) & (!g3189) & (!g3190) & (g3270)) + ((g18) & (g27) & (!g3189) & (g3190) & (!g3270)) + ((g18) & (g27) & (!g3189) & (g3190) & (g3270)) + ((g18) & (g27) & (g3189) & (!g3190) & (!g3270)) + ((g18) & (g27) & (g3189) & (!g3190) & (g3270)) + ((g18) & (g27) & (g3189) & (g3190) & (!g3270)) + ((g18) & (g27) & (g3189) & (g3190) & (g3270)));
	assign g3272 = (((g1) & (!g3061) & (!g3177) & (!g3178) & (g3179) & (!g3186)) + ((g1) & (!g3061) & (!g3177) & (g3178) & (g3179) & (!g3186)) + ((g1) & (!g3061) & (g3177) & (!g3178) & (!g3179) & (g3186)) + ((g1) & (!g3061) & (g3177) & (!g3178) & (g3179) & (!g3186)) + ((g1) & (!g3061) & (g3177) & (g3178) & (g3179) & (!g3186)) + ((g1) & (g3061) & (!g3177) & (!g3178) & (!g3179) & (g3186)) + ((g1) & (g3061) & (!g3177) & (!g3178) & (g3179) & (!g3186)) + ((g1) & (g3061) & (!g3177) & (g3178) & (!g3179) & (g3186)) + ((g1) & (g3061) & (!g3177) & (g3178) & (g3179) & (!g3186)) + ((g1) & (g3061) & (g3177) & (!g3178) & (g3179) & (!g3186)) + ((g1) & (g3061) & (g3177) & (g3178) & (g3179) & (!g3186)));
	assign g3273 = (((!g4) & (!g2) & (!g3180) & (!g3183) & (!g3185) & (!g3187)) + ((!g4) & (!g2) & (!g3180) & (!g3183) & (g3185) & (g3187)) + ((!g4) & (!g2) & (!g3180) & (g3183) & (!g3185) & (!g3187)) + ((!g4) & (!g2) & (!g3180) & (g3183) & (g3185) & (g3187)) + ((!g4) & (!g2) & (g3180) & (!g3183) & (!g3185) & (!g3187)) + ((!g4) & (!g2) & (g3180) & (!g3183) & (g3185) & (g3187)) + ((!g4) & (!g2) & (g3180) & (g3183) & (g3185) & (!g3187)) + ((!g4) & (!g2) & (g3180) & (g3183) & (g3185) & (g3187)) + ((!g4) & (g2) & (!g3180) & (!g3183) & (!g3185) & (!g3187)) + ((!g4) & (g2) & (!g3180) & (!g3183) & (g3185) & (g3187)) + ((!g4) & (g2) & (!g3180) & (g3183) & (g3185) & (!g3187)) + ((!g4) & (g2) & (!g3180) & (g3183) & (g3185) & (g3187)) + ((!g4) & (g2) & (g3180) & (!g3183) & (g3185) & (!g3187)) + ((!g4) & (g2) & (g3180) & (!g3183) & (g3185) & (g3187)) + ((!g4) & (g2) & (g3180) & (g3183) & (g3185) & (!g3187)) + ((!g4) & (g2) & (g3180) & (g3183) & (g3185) & (g3187)) + ((g4) & (!g2) & (!g3180) & (!g3183) & (g3185) & (!g3187)) + ((g4) & (!g2) & (!g3180) & (!g3183) & (g3185) & (g3187)) + ((g4) & (!g2) & (!g3180) & (g3183) & (g3185) & (!g3187)) + ((g4) & (!g2) & (!g3180) & (g3183) & (g3185) & (g3187)) + ((g4) & (!g2) & (g3180) & (!g3183) & (g3185) & (!g3187)) + ((g4) & (!g2) & (g3180) & (!g3183) & (g3185) & (g3187)) + ((g4) & (!g2) & (g3180) & (g3183) & (!g3185) & (!g3187)) + ((g4) & (!g2) & (g3180) & (g3183) & (g3185) & (g3187)) + ((g4) & (g2) & (!g3180) & (!g3183) & (g3185) & (!g3187)) + ((g4) & (g2) & (!g3180) & (!g3183) & (g3185) & (g3187)) + ((g4) & (g2) & (!g3180) & (g3183) & (!g3185) & (!g3187)) + ((g4) & (g2) & (!g3180) & (g3183) & (g3185) & (g3187)) + ((g4) & (g2) & (g3180) & (!g3183) & (!g3185) & (!g3187)) + ((g4) & (g2) & (g3180) & (!g3183) & (g3185) & (g3187)) + ((g4) & (g2) & (g3180) & (g3183) & (!g3185) & (!g3187)) + ((g4) & (g2) & (g3180) & (g3183) & (g3185) & (g3187)));
	assign g3274 = (((!g8) & (!g18) & (!g3182) & (g3070) & (g3176) & (!g3187)) + ((!g8) & (!g18) & (g3182) & (!g3070) & (!g3176) & (!g3187)) + ((!g8) & (!g18) & (g3182) & (!g3070) & (!g3176) & (g3187)) + ((!g8) & (!g18) & (g3182) & (!g3070) & (g3176) & (!g3187)) + ((!g8) & (!g18) & (g3182) & (!g3070) & (g3176) & (g3187)) + ((!g8) & (!g18) & (g3182) & (g3070) & (!g3176) & (!g3187)) + ((!g8) & (!g18) & (g3182) & (g3070) & (!g3176) & (g3187)) + ((!g8) & (!g18) & (g3182) & (g3070) & (g3176) & (g3187)) + ((!g8) & (g18) & (!g3182) & (!g3070) & (g3176) & (!g3187)) + ((!g8) & (g18) & (!g3182) & (g3070) & (!g3176) & (!g3187)) + ((!g8) & (g18) & (!g3182) & (g3070) & (g3176) & (!g3187)) + ((!g8) & (g18) & (g3182) & (!g3070) & (!g3176) & (!g3187)) + ((!g8) & (g18) & (g3182) & (!g3070) & (!g3176) & (g3187)) + ((!g8) & (g18) & (g3182) & (!g3070) & (g3176) & (g3187)) + ((!g8) & (g18) & (g3182) & (g3070) & (!g3176) & (g3187)) + ((!g8) & (g18) & (g3182) & (g3070) & (g3176) & (g3187)) + ((g8) & (!g18) & (!g3182) & (!g3070) & (!g3176) & (!g3187)) + ((g8) & (!g18) & (!g3182) & (!g3070) & (g3176) & (!g3187)) + ((g8) & (!g18) & (!g3182) & (g3070) & (!g3176) & (!g3187)) + ((g8) & (!g18) & (g3182) & (!g3070) & (!g3176) & (g3187)) + ((g8) & (!g18) & (g3182) & (!g3070) & (g3176) & (g3187)) + ((g8) & (!g18) & (g3182) & (g3070) & (!g3176) & (g3187)) + ((g8) & (!g18) & (g3182) & (g3070) & (g3176) & (!g3187)) + ((g8) & (!g18) & (g3182) & (g3070) & (g3176) & (g3187)) + ((g8) & (g18) & (!g3182) & (!g3070) & (!g3176) & (!g3187)) + ((g8) & (g18) & (g3182) & (!g3070) & (!g3176) & (g3187)) + ((g8) & (g18) & (g3182) & (!g3070) & (g3176) & (!g3187)) + ((g8) & (g18) & (g3182) & (!g3070) & (g3176) & (g3187)) + ((g8) & (g18) & (g3182) & (g3070) & (!g3176) & (!g3187)) + ((g8) & (g18) & (g3182) & (g3070) & (!g3176) & (g3187)) + ((g8) & (g18) & (g3182) & (g3070) & (g3176) & (!g3187)) + ((g8) & (g18) & (g3182) & (g3070) & (g3176) & (g3187)));
	assign g3275 = (((!g2) & (!g8) & (g3274) & (g3188) & (g3271)) + ((!g2) & (g8) & (g3274) & (!g3188) & (g3271)) + ((!g2) & (g8) & (g3274) & (g3188) & (!g3271)) + ((!g2) & (g8) & (g3274) & (g3188) & (g3271)) + ((g2) & (!g8) & (!g3274) & (g3188) & (g3271)) + ((g2) & (!g8) & (g3274) & (!g3188) & (!g3271)) + ((g2) & (!g8) & (g3274) & (!g3188) & (g3271)) + ((g2) & (!g8) & (g3274) & (g3188) & (!g3271)) + ((g2) & (!g8) & (g3274) & (g3188) & (g3271)) + ((g2) & (g8) & (!g3274) & (!g3188) & (g3271)) + ((g2) & (g8) & (!g3274) & (g3188) & (!g3271)) + ((g2) & (g8) & (!g3274) & (g3188) & (g3271)) + ((g2) & (g8) & (g3274) & (!g3188) & (!g3271)) + ((g2) & (g8) & (g3274) & (!g3188) & (g3271)) + ((g2) & (g8) & (g3274) & (g3188) & (!g3271)) + ((g2) & (g8) & (g3274) & (g3188) & (g3271)));
	assign g3276 = (((!g2) & (!g3180) & (g3183) & (!g3187)) + ((!g2) & (g3180) & (!g3183) & (!g3187)) + ((!g2) & (g3180) & (!g3183) & (g3187)) + ((!g2) & (g3180) & (g3183) & (g3187)) + ((g2) & (!g3180) & (!g3183) & (!g3187)) + ((g2) & (g3180) & (!g3183) & (g3187)) + ((g2) & (g3180) & (g3183) & (!g3187)) + ((g2) & (g3180) & (g3183) & (g3187)));
	assign g3277 = (((!g1) & (!g3061) & (!g3177) & (!g3178) & (!g3179) & (!g3186)) + ((!g1) & (!g3061) & (!g3177) & (!g3178) & (g3179) & (g3186)) + ((!g1) & (!g3061) & (!g3177) & (g3178) & (g3179) & (g3186)) + ((!g1) & (!g3061) & (g3177) & (!g3178) & (g3179) & (g3186)) + ((!g1) & (!g3061) & (g3177) & (g3178) & (g3179) & (g3186)) + ((!g1) & (g3061) & (!g3177) & (!g3178) & (g3179) & (g3186)) + ((!g1) & (g3061) & (!g3177) & (g3178) & (g3179) & (g3186)) + ((!g1) & (g3061) & (g3177) & (!g3178) & (!g3179) & (!g3186)) + ((!g1) & (g3061) & (g3177) & (!g3178) & (g3179) & (g3186)) + ((!g1) & (g3061) & (g3177) & (g3178) & (!g3179) & (!g3186)) + ((!g1) & (g3061) & (g3177) & (g3178) & (g3179) & (g3186)) + ((g1) & (!g3061) & (!g3177) & (!g3178) & (g3179) & (g3186)) + ((g1) & (!g3061) & (!g3177) & (g3178) & (g3179) & (g3186)) + ((g1) & (!g3061) & (g3177) & (!g3178) & (!g3179) & (!g3186)) + ((g1) & (!g3061) & (g3177) & (!g3178) & (g3179) & (g3186)) + ((g1) & (!g3061) & (g3177) & (g3178) & (g3179) & (g3186)) + ((g1) & (g3061) & (!g3177) & (!g3178) & (!g3179) & (!g3186)) + ((g1) & (g3061) & (!g3177) & (!g3178) & (g3179) & (g3186)) + ((g1) & (g3061) & (!g3177) & (g3178) & (!g3179) & (!g3186)) + ((g1) & (g3061) & (!g3177) & (g3178) & (g3179) & (g3186)) + ((g1) & (g3061) & (g3177) & (!g3178) & (g3179) & (g3186)) + ((g1) & (g3061) & (g3177) & (g3178) & (g3179) & (g3186)));
	assign g3278 = (((!g4) & (!g1) & (!g3273) & (!g3275) & (!g3276) & (!g3277)) + ((!g4) & (g1) & (!g3273) & (!g3275) & (!g3276) & (!g3277)) + ((!g4) & (g1) & (!g3273) & (!g3275) & (!g3276) & (g3277)) + ((!g4) & (g1) & (!g3273) & (!g3275) & (g3276) & (!g3277)) + ((!g4) & (g1) & (!g3273) & (!g3275) & (g3276) & (g3277)) + ((!g4) & (g1) & (!g3273) & (g3275) & (!g3276) & (!g3277)) + ((!g4) & (g1) & (!g3273) & (g3275) & (!g3276) & (g3277)) + ((!g4) & (g1) & (!g3273) & (g3275) & (g3276) & (!g3277)) + ((!g4) & (g1) & (!g3273) & (g3275) & (g3276) & (g3277)) + ((!g4) & (g1) & (g3273) & (!g3275) & (!g3276) & (!g3277)) + ((!g4) & (g1) & (g3273) & (!g3275) & (!g3276) & (g3277)) + ((g4) & (!g1) & (!g3273) & (!g3275) & (!g3276) & (!g3277)) + ((g4) & (!g1) & (!g3273) & (!g3275) & (g3276) & (!g3277)) + ((g4) & (!g1) & (!g3273) & (g3275) & (!g3276) & (!g3277)) + ((g4) & (g1) & (!g3273) & (!g3275) & (!g3276) & (!g3277)) + ((g4) & (g1) & (!g3273) & (!g3275) & (!g3276) & (g3277)) + ((g4) & (g1) & (!g3273) & (!g3275) & (g3276) & (!g3277)) + ((g4) & (g1) & (!g3273) & (!g3275) & (g3276) & (g3277)) + ((g4) & (g1) & (!g3273) & (g3275) & (!g3276) & (!g3277)) + ((g4) & (g1) & (!g3273) & (g3275) & (!g3276) & (g3277)) + ((g4) & (g1) & (!g3273) & (g3275) & (g3276) & (!g3277)) + ((g4) & (g1) & (!g3273) & (g3275) & (g3276) & (g3277)) + ((g4) & (g1) & (g3273) & (!g3275) & (!g3276) & (!g3277)) + ((g4) & (g1) & (g3273) & (!g3275) & (!g3276) & (g3277)) + ((g4) & (g1) & (g3273) & (!g3275) & (g3276) & (!g3277)) + ((g4) & (g1) & (g3273) & (!g3275) & (g3276) & (g3277)) + ((g4) & (g1) & (g3273) & (g3275) & (!g3276) & (!g3277)) + ((g4) & (g1) & (g3273) & (g3275) & (!g3276) & (g3277)));
	assign g3279 = (((!g8) & (!g3188) & (g3271) & (!g3272) & (!g3278)) + ((!g8) & (!g3188) & (g3271) & (g3272) & (!g3278)) + ((!g8) & (!g3188) & (g3271) & (g3272) & (g3278)) + ((!g8) & (g3188) & (!g3271) & (!g3272) & (!g3278)) + ((!g8) & (g3188) & (!g3271) & (!g3272) & (g3278)) + ((!g8) & (g3188) & (!g3271) & (g3272) & (!g3278)) + ((!g8) & (g3188) & (!g3271) & (g3272) & (g3278)) + ((!g8) & (g3188) & (g3271) & (!g3272) & (g3278)) + ((g8) & (!g3188) & (!g3271) & (!g3272) & (!g3278)) + ((g8) & (!g3188) & (!g3271) & (g3272) & (!g3278)) + ((g8) & (!g3188) & (!g3271) & (g3272) & (g3278)) + ((g8) & (g3188) & (!g3271) & (!g3272) & (g3278)) + ((g8) & (g3188) & (g3271) & (!g3272) & (!g3278)) + ((g8) & (g3188) & (g3271) & (!g3272) & (g3278)) + ((g8) & (g3188) & (g3271) & (g3272) & (!g3278)) + ((g8) & (g3188) & (g3271) & (g3272) & (g3278)));
	assign g3280 = (((!g18) & (!g27) & (g3190) & (g3270)) + ((!g18) & (g27) & (!g3190) & (g3270)) + ((!g18) & (g27) & (g3190) & (!g3270)) + ((!g18) & (g27) & (g3190) & (g3270)) + ((g18) & (!g27) & (!g3190) & (!g3270)) + ((g18) & (!g27) & (!g3190) & (g3270)) + ((g18) & (!g27) & (g3190) & (!g3270)) + ((g18) & (g27) & (!g3190) & (!g3270)));
	assign g3281 = (((!g3189) & (!g3272) & (!g3278) & (g3280)) + ((!g3189) & (g3272) & (!g3278) & (g3280)) + ((!g3189) & (g3272) & (g3278) & (g3280)) + ((g3189) & (!g3272) & (!g3278) & (!g3280)) + ((g3189) & (!g3272) & (g3278) & (!g3280)) + ((g3189) & (!g3272) & (g3278) & (g3280)) + ((g3189) & (g3272) & (!g3278) & (!g3280)) + ((g3189) & (g3272) & (g3278) & (!g3280)));
	assign g3282 = (((!g27) & (!g3190) & (g3270) & (!g3272) & (!g3278)) + ((!g27) & (!g3190) & (g3270) & (g3272) & (!g3278)) + ((!g27) & (!g3190) & (g3270) & (g3272) & (g3278)) + ((!g27) & (g3190) & (!g3270) & (!g3272) & (!g3278)) + ((!g27) & (g3190) & (!g3270) & (!g3272) & (g3278)) + ((!g27) & (g3190) & (!g3270) & (g3272) & (!g3278)) + ((!g27) & (g3190) & (!g3270) & (g3272) & (g3278)) + ((!g27) & (g3190) & (g3270) & (!g3272) & (g3278)) + ((g27) & (!g3190) & (!g3270) & (!g3272) & (!g3278)) + ((g27) & (!g3190) & (!g3270) & (g3272) & (!g3278)) + ((g27) & (!g3190) & (!g3270) & (g3272) & (g3278)) + ((g27) & (g3190) & (!g3270) & (!g3272) & (g3278)) + ((g27) & (g3190) & (g3270) & (!g3272) & (!g3278)) + ((g27) & (g3190) & (g3270) & (!g3272) & (g3278)) + ((g27) & (g3190) & (g3270) & (g3272) & (!g3278)) + ((g27) & (g3190) & (g3270) & (g3272) & (g3278)));
	assign g3283 = (((!g39) & (!g54) & (g3192) & (g3269)) + ((!g39) & (g54) & (!g3192) & (g3269)) + ((!g39) & (g54) & (g3192) & (!g3269)) + ((!g39) & (g54) & (g3192) & (g3269)) + ((g39) & (!g54) & (!g3192) & (!g3269)) + ((g39) & (!g54) & (!g3192) & (g3269)) + ((g39) & (!g54) & (g3192) & (!g3269)) + ((g39) & (g54) & (!g3192) & (!g3269)));
	assign g3284 = (((!g3191) & (!g3272) & (!g3278) & (g3283)) + ((!g3191) & (g3272) & (!g3278) & (g3283)) + ((!g3191) & (g3272) & (g3278) & (g3283)) + ((g3191) & (!g3272) & (!g3278) & (!g3283)) + ((g3191) & (!g3272) & (g3278) & (!g3283)) + ((g3191) & (!g3272) & (g3278) & (g3283)) + ((g3191) & (g3272) & (!g3278) & (!g3283)) + ((g3191) & (g3272) & (g3278) & (!g3283)));
	assign g3285 = (((!g54) & (!g3192) & (g3269) & (!g3272) & (!g3278)) + ((!g54) & (!g3192) & (g3269) & (g3272) & (!g3278)) + ((!g54) & (!g3192) & (g3269) & (g3272) & (g3278)) + ((!g54) & (g3192) & (!g3269) & (!g3272) & (!g3278)) + ((!g54) & (g3192) & (!g3269) & (!g3272) & (g3278)) + ((!g54) & (g3192) & (!g3269) & (g3272) & (!g3278)) + ((!g54) & (g3192) & (!g3269) & (g3272) & (g3278)) + ((!g54) & (g3192) & (g3269) & (!g3272) & (g3278)) + ((g54) & (!g3192) & (!g3269) & (!g3272) & (!g3278)) + ((g54) & (!g3192) & (!g3269) & (g3272) & (!g3278)) + ((g54) & (!g3192) & (!g3269) & (g3272) & (g3278)) + ((g54) & (g3192) & (!g3269) & (!g3272) & (g3278)) + ((g54) & (g3192) & (g3269) & (!g3272) & (!g3278)) + ((g54) & (g3192) & (g3269) & (!g3272) & (g3278)) + ((g54) & (g3192) & (g3269) & (g3272) & (!g3278)) + ((g54) & (g3192) & (g3269) & (g3272) & (g3278)));
	assign g3286 = (((!g68) & (!g87) & (g3194) & (g3268)) + ((!g68) & (g87) & (!g3194) & (g3268)) + ((!g68) & (g87) & (g3194) & (!g3268)) + ((!g68) & (g87) & (g3194) & (g3268)) + ((g68) & (!g87) & (!g3194) & (!g3268)) + ((g68) & (!g87) & (!g3194) & (g3268)) + ((g68) & (!g87) & (g3194) & (!g3268)) + ((g68) & (g87) & (!g3194) & (!g3268)));
	assign g3287 = (((!g3193) & (!g3272) & (!g3278) & (g3286)) + ((!g3193) & (g3272) & (!g3278) & (g3286)) + ((!g3193) & (g3272) & (g3278) & (g3286)) + ((g3193) & (!g3272) & (!g3278) & (!g3286)) + ((g3193) & (!g3272) & (g3278) & (!g3286)) + ((g3193) & (!g3272) & (g3278) & (g3286)) + ((g3193) & (g3272) & (!g3278) & (!g3286)) + ((g3193) & (g3272) & (g3278) & (!g3286)));
	assign g3288 = (((!g87) & (!g3194) & (g3268) & (!g3272) & (!g3278)) + ((!g87) & (!g3194) & (g3268) & (g3272) & (!g3278)) + ((!g87) & (!g3194) & (g3268) & (g3272) & (g3278)) + ((!g87) & (g3194) & (!g3268) & (!g3272) & (!g3278)) + ((!g87) & (g3194) & (!g3268) & (!g3272) & (g3278)) + ((!g87) & (g3194) & (!g3268) & (g3272) & (!g3278)) + ((!g87) & (g3194) & (!g3268) & (g3272) & (g3278)) + ((!g87) & (g3194) & (g3268) & (!g3272) & (g3278)) + ((g87) & (!g3194) & (!g3268) & (!g3272) & (!g3278)) + ((g87) & (!g3194) & (!g3268) & (g3272) & (!g3278)) + ((g87) & (!g3194) & (!g3268) & (g3272) & (g3278)) + ((g87) & (g3194) & (!g3268) & (!g3272) & (g3278)) + ((g87) & (g3194) & (g3268) & (!g3272) & (!g3278)) + ((g87) & (g3194) & (g3268) & (!g3272) & (g3278)) + ((g87) & (g3194) & (g3268) & (g3272) & (!g3278)) + ((g87) & (g3194) & (g3268) & (g3272) & (g3278)));
	assign g3289 = (((!g104) & (!g127) & (g3196) & (g3267)) + ((!g104) & (g127) & (!g3196) & (g3267)) + ((!g104) & (g127) & (g3196) & (!g3267)) + ((!g104) & (g127) & (g3196) & (g3267)) + ((g104) & (!g127) & (!g3196) & (!g3267)) + ((g104) & (!g127) & (!g3196) & (g3267)) + ((g104) & (!g127) & (g3196) & (!g3267)) + ((g104) & (g127) & (!g3196) & (!g3267)));
	assign g3290 = (((!g3195) & (!g3272) & (!g3278) & (g3289)) + ((!g3195) & (g3272) & (!g3278) & (g3289)) + ((!g3195) & (g3272) & (g3278) & (g3289)) + ((g3195) & (!g3272) & (!g3278) & (!g3289)) + ((g3195) & (!g3272) & (g3278) & (!g3289)) + ((g3195) & (!g3272) & (g3278) & (g3289)) + ((g3195) & (g3272) & (!g3278) & (!g3289)) + ((g3195) & (g3272) & (g3278) & (!g3289)));
	assign g3291 = (((!g127) & (!g3196) & (g3267) & (!g3272) & (!g3278)) + ((!g127) & (!g3196) & (g3267) & (g3272) & (!g3278)) + ((!g127) & (!g3196) & (g3267) & (g3272) & (g3278)) + ((!g127) & (g3196) & (!g3267) & (!g3272) & (!g3278)) + ((!g127) & (g3196) & (!g3267) & (!g3272) & (g3278)) + ((!g127) & (g3196) & (!g3267) & (g3272) & (!g3278)) + ((!g127) & (g3196) & (!g3267) & (g3272) & (g3278)) + ((!g127) & (g3196) & (g3267) & (!g3272) & (g3278)) + ((g127) & (!g3196) & (!g3267) & (!g3272) & (!g3278)) + ((g127) & (!g3196) & (!g3267) & (g3272) & (!g3278)) + ((g127) & (!g3196) & (!g3267) & (g3272) & (g3278)) + ((g127) & (g3196) & (!g3267) & (!g3272) & (g3278)) + ((g127) & (g3196) & (g3267) & (!g3272) & (!g3278)) + ((g127) & (g3196) & (g3267) & (!g3272) & (g3278)) + ((g127) & (g3196) & (g3267) & (g3272) & (!g3278)) + ((g127) & (g3196) & (g3267) & (g3272) & (g3278)));
	assign g3292 = (((!g147) & (!g174) & (g3198) & (g3266)) + ((!g147) & (g174) & (!g3198) & (g3266)) + ((!g147) & (g174) & (g3198) & (!g3266)) + ((!g147) & (g174) & (g3198) & (g3266)) + ((g147) & (!g174) & (!g3198) & (!g3266)) + ((g147) & (!g174) & (!g3198) & (g3266)) + ((g147) & (!g174) & (g3198) & (!g3266)) + ((g147) & (g174) & (!g3198) & (!g3266)));
	assign g3293 = (((!g3197) & (!g3272) & (!g3278) & (g3292)) + ((!g3197) & (g3272) & (!g3278) & (g3292)) + ((!g3197) & (g3272) & (g3278) & (g3292)) + ((g3197) & (!g3272) & (!g3278) & (!g3292)) + ((g3197) & (!g3272) & (g3278) & (!g3292)) + ((g3197) & (!g3272) & (g3278) & (g3292)) + ((g3197) & (g3272) & (!g3278) & (!g3292)) + ((g3197) & (g3272) & (g3278) & (!g3292)));
	assign g3294 = (((!g174) & (!g3198) & (g3266) & (!g3272) & (!g3278)) + ((!g174) & (!g3198) & (g3266) & (g3272) & (!g3278)) + ((!g174) & (!g3198) & (g3266) & (g3272) & (g3278)) + ((!g174) & (g3198) & (!g3266) & (!g3272) & (!g3278)) + ((!g174) & (g3198) & (!g3266) & (!g3272) & (g3278)) + ((!g174) & (g3198) & (!g3266) & (g3272) & (!g3278)) + ((!g174) & (g3198) & (!g3266) & (g3272) & (g3278)) + ((!g174) & (g3198) & (g3266) & (!g3272) & (g3278)) + ((g174) & (!g3198) & (!g3266) & (!g3272) & (!g3278)) + ((g174) & (!g3198) & (!g3266) & (g3272) & (!g3278)) + ((g174) & (!g3198) & (!g3266) & (g3272) & (g3278)) + ((g174) & (g3198) & (!g3266) & (!g3272) & (g3278)) + ((g174) & (g3198) & (g3266) & (!g3272) & (!g3278)) + ((g174) & (g3198) & (g3266) & (!g3272) & (g3278)) + ((g174) & (g3198) & (g3266) & (g3272) & (!g3278)) + ((g174) & (g3198) & (g3266) & (g3272) & (g3278)));
	assign g3295 = (((!g198) & (!g229) & (g3200) & (g3265)) + ((!g198) & (g229) & (!g3200) & (g3265)) + ((!g198) & (g229) & (g3200) & (!g3265)) + ((!g198) & (g229) & (g3200) & (g3265)) + ((g198) & (!g229) & (!g3200) & (!g3265)) + ((g198) & (!g229) & (!g3200) & (g3265)) + ((g198) & (!g229) & (g3200) & (!g3265)) + ((g198) & (g229) & (!g3200) & (!g3265)));
	assign g3296 = (((!g3199) & (!g3272) & (!g3278) & (g3295)) + ((!g3199) & (g3272) & (!g3278) & (g3295)) + ((!g3199) & (g3272) & (g3278) & (g3295)) + ((g3199) & (!g3272) & (!g3278) & (!g3295)) + ((g3199) & (!g3272) & (g3278) & (!g3295)) + ((g3199) & (!g3272) & (g3278) & (g3295)) + ((g3199) & (g3272) & (!g3278) & (!g3295)) + ((g3199) & (g3272) & (g3278) & (!g3295)));
	assign g3297 = (((!g229) & (!g3200) & (g3265) & (!g3272) & (!g3278)) + ((!g229) & (!g3200) & (g3265) & (g3272) & (!g3278)) + ((!g229) & (!g3200) & (g3265) & (g3272) & (g3278)) + ((!g229) & (g3200) & (!g3265) & (!g3272) & (!g3278)) + ((!g229) & (g3200) & (!g3265) & (!g3272) & (g3278)) + ((!g229) & (g3200) & (!g3265) & (g3272) & (!g3278)) + ((!g229) & (g3200) & (!g3265) & (g3272) & (g3278)) + ((!g229) & (g3200) & (g3265) & (!g3272) & (g3278)) + ((g229) & (!g3200) & (!g3265) & (!g3272) & (!g3278)) + ((g229) & (!g3200) & (!g3265) & (g3272) & (!g3278)) + ((g229) & (!g3200) & (!g3265) & (g3272) & (g3278)) + ((g229) & (g3200) & (!g3265) & (!g3272) & (g3278)) + ((g229) & (g3200) & (g3265) & (!g3272) & (!g3278)) + ((g229) & (g3200) & (g3265) & (!g3272) & (g3278)) + ((g229) & (g3200) & (g3265) & (g3272) & (!g3278)) + ((g229) & (g3200) & (g3265) & (g3272) & (g3278)));
	assign g3298 = (((!g255) & (!g290) & (g3202) & (g3264)) + ((!g255) & (g290) & (!g3202) & (g3264)) + ((!g255) & (g290) & (g3202) & (!g3264)) + ((!g255) & (g290) & (g3202) & (g3264)) + ((g255) & (!g290) & (!g3202) & (!g3264)) + ((g255) & (!g290) & (!g3202) & (g3264)) + ((g255) & (!g290) & (g3202) & (!g3264)) + ((g255) & (g290) & (!g3202) & (!g3264)));
	assign g3299 = (((!g3201) & (!g3272) & (!g3278) & (g3298)) + ((!g3201) & (g3272) & (!g3278) & (g3298)) + ((!g3201) & (g3272) & (g3278) & (g3298)) + ((g3201) & (!g3272) & (!g3278) & (!g3298)) + ((g3201) & (!g3272) & (g3278) & (!g3298)) + ((g3201) & (!g3272) & (g3278) & (g3298)) + ((g3201) & (g3272) & (!g3278) & (!g3298)) + ((g3201) & (g3272) & (g3278) & (!g3298)));
	assign g3300 = (((!g290) & (!g3202) & (g3264) & (!g3272) & (!g3278)) + ((!g290) & (!g3202) & (g3264) & (g3272) & (!g3278)) + ((!g290) & (!g3202) & (g3264) & (g3272) & (g3278)) + ((!g290) & (g3202) & (!g3264) & (!g3272) & (!g3278)) + ((!g290) & (g3202) & (!g3264) & (!g3272) & (g3278)) + ((!g290) & (g3202) & (!g3264) & (g3272) & (!g3278)) + ((!g290) & (g3202) & (!g3264) & (g3272) & (g3278)) + ((!g290) & (g3202) & (g3264) & (!g3272) & (g3278)) + ((g290) & (!g3202) & (!g3264) & (!g3272) & (!g3278)) + ((g290) & (!g3202) & (!g3264) & (g3272) & (!g3278)) + ((g290) & (!g3202) & (!g3264) & (g3272) & (g3278)) + ((g290) & (g3202) & (!g3264) & (!g3272) & (g3278)) + ((g290) & (g3202) & (g3264) & (!g3272) & (!g3278)) + ((g290) & (g3202) & (g3264) & (!g3272) & (g3278)) + ((g290) & (g3202) & (g3264) & (g3272) & (!g3278)) + ((g290) & (g3202) & (g3264) & (g3272) & (g3278)));
	assign g3301 = (((!g319) & (!g358) & (g3204) & (g3263)) + ((!g319) & (g358) & (!g3204) & (g3263)) + ((!g319) & (g358) & (g3204) & (!g3263)) + ((!g319) & (g358) & (g3204) & (g3263)) + ((g319) & (!g358) & (!g3204) & (!g3263)) + ((g319) & (!g358) & (!g3204) & (g3263)) + ((g319) & (!g358) & (g3204) & (!g3263)) + ((g319) & (g358) & (!g3204) & (!g3263)));
	assign g3302 = (((!g3203) & (!g3272) & (!g3278) & (g3301)) + ((!g3203) & (g3272) & (!g3278) & (g3301)) + ((!g3203) & (g3272) & (g3278) & (g3301)) + ((g3203) & (!g3272) & (!g3278) & (!g3301)) + ((g3203) & (!g3272) & (g3278) & (!g3301)) + ((g3203) & (!g3272) & (g3278) & (g3301)) + ((g3203) & (g3272) & (!g3278) & (!g3301)) + ((g3203) & (g3272) & (g3278) & (!g3301)));
	assign g3303 = (((!g358) & (!g3204) & (g3263) & (!g3272) & (!g3278)) + ((!g358) & (!g3204) & (g3263) & (g3272) & (!g3278)) + ((!g358) & (!g3204) & (g3263) & (g3272) & (g3278)) + ((!g358) & (g3204) & (!g3263) & (!g3272) & (!g3278)) + ((!g358) & (g3204) & (!g3263) & (!g3272) & (g3278)) + ((!g358) & (g3204) & (!g3263) & (g3272) & (!g3278)) + ((!g358) & (g3204) & (!g3263) & (g3272) & (g3278)) + ((!g358) & (g3204) & (g3263) & (!g3272) & (g3278)) + ((g358) & (!g3204) & (!g3263) & (!g3272) & (!g3278)) + ((g358) & (!g3204) & (!g3263) & (g3272) & (!g3278)) + ((g358) & (!g3204) & (!g3263) & (g3272) & (g3278)) + ((g358) & (g3204) & (!g3263) & (!g3272) & (g3278)) + ((g358) & (g3204) & (g3263) & (!g3272) & (!g3278)) + ((g358) & (g3204) & (g3263) & (!g3272) & (g3278)) + ((g358) & (g3204) & (g3263) & (g3272) & (!g3278)) + ((g358) & (g3204) & (g3263) & (g3272) & (g3278)));
	assign g3304 = (((!g390) & (!g433) & (g3206) & (g3262)) + ((!g390) & (g433) & (!g3206) & (g3262)) + ((!g390) & (g433) & (g3206) & (!g3262)) + ((!g390) & (g433) & (g3206) & (g3262)) + ((g390) & (!g433) & (!g3206) & (!g3262)) + ((g390) & (!g433) & (!g3206) & (g3262)) + ((g390) & (!g433) & (g3206) & (!g3262)) + ((g390) & (g433) & (!g3206) & (!g3262)));
	assign g3305 = (((!g3205) & (!g3272) & (!g3278) & (g3304)) + ((!g3205) & (g3272) & (!g3278) & (g3304)) + ((!g3205) & (g3272) & (g3278) & (g3304)) + ((g3205) & (!g3272) & (!g3278) & (!g3304)) + ((g3205) & (!g3272) & (g3278) & (!g3304)) + ((g3205) & (!g3272) & (g3278) & (g3304)) + ((g3205) & (g3272) & (!g3278) & (!g3304)) + ((g3205) & (g3272) & (g3278) & (!g3304)));
	assign g3306 = (((!g433) & (!g3206) & (g3262) & (!g3272) & (!g3278)) + ((!g433) & (!g3206) & (g3262) & (g3272) & (!g3278)) + ((!g433) & (!g3206) & (g3262) & (g3272) & (g3278)) + ((!g433) & (g3206) & (!g3262) & (!g3272) & (!g3278)) + ((!g433) & (g3206) & (!g3262) & (!g3272) & (g3278)) + ((!g433) & (g3206) & (!g3262) & (g3272) & (!g3278)) + ((!g433) & (g3206) & (!g3262) & (g3272) & (g3278)) + ((!g433) & (g3206) & (g3262) & (!g3272) & (g3278)) + ((g433) & (!g3206) & (!g3262) & (!g3272) & (!g3278)) + ((g433) & (!g3206) & (!g3262) & (g3272) & (!g3278)) + ((g433) & (!g3206) & (!g3262) & (g3272) & (g3278)) + ((g433) & (g3206) & (!g3262) & (!g3272) & (g3278)) + ((g433) & (g3206) & (g3262) & (!g3272) & (!g3278)) + ((g433) & (g3206) & (g3262) & (!g3272) & (g3278)) + ((g433) & (g3206) & (g3262) & (g3272) & (!g3278)) + ((g433) & (g3206) & (g3262) & (g3272) & (g3278)));
	assign g3307 = (((!g468) & (!g515) & (g3208) & (g3261)) + ((!g468) & (g515) & (!g3208) & (g3261)) + ((!g468) & (g515) & (g3208) & (!g3261)) + ((!g468) & (g515) & (g3208) & (g3261)) + ((g468) & (!g515) & (!g3208) & (!g3261)) + ((g468) & (!g515) & (!g3208) & (g3261)) + ((g468) & (!g515) & (g3208) & (!g3261)) + ((g468) & (g515) & (!g3208) & (!g3261)));
	assign g3308 = (((!g3207) & (!g3272) & (!g3278) & (g3307)) + ((!g3207) & (g3272) & (!g3278) & (g3307)) + ((!g3207) & (g3272) & (g3278) & (g3307)) + ((g3207) & (!g3272) & (!g3278) & (!g3307)) + ((g3207) & (!g3272) & (g3278) & (!g3307)) + ((g3207) & (!g3272) & (g3278) & (g3307)) + ((g3207) & (g3272) & (!g3278) & (!g3307)) + ((g3207) & (g3272) & (g3278) & (!g3307)));
	assign g3309 = (((!g515) & (!g3208) & (g3261) & (!g3272) & (!g3278)) + ((!g515) & (!g3208) & (g3261) & (g3272) & (!g3278)) + ((!g515) & (!g3208) & (g3261) & (g3272) & (g3278)) + ((!g515) & (g3208) & (!g3261) & (!g3272) & (!g3278)) + ((!g515) & (g3208) & (!g3261) & (!g3272) & (g3278)) + ((!g515) & (g3208) & (!g3261) & (g3272) & (!g3278)) + ((!g515) & (g3208) & (!g3261) & (g3272) & (g3278)) + ((!g515) & (g3208) & (g3261) & (!g3272) & (g3278)) + ((g515) & (!g3208) & (!g3261) & (!g3272) & (!g3278)) + ((g515) & (!g3208) & (!g3261) & (g3272) & (!g3278)) + ((g515) & (!g3208) & (!g3261) & (g3272) & (g3278)) + ((g515) & (g3208) & (!g3261) & (!g3272) & (g3278)) + ((g515) & (g3208) & (g3261) & (!g3272) & (!g3278)) + ((g515) & (g3208) & (g3261) & (!g3272) & (g3278)) + ((g515) & (g3208) & (g3261) & (g3272) & (!g3278)) + ((g515) & (g3208) & (g3261) & (g3272) & (g3278)));
	assign g3310 = (((!g553) & (!g604) & (g3210) & (g3260)) + ((!g553) & (g604) & (!g3210) & (g3260)) + ((!g553) & (g604) & (g3210) & (!g3260)) + ((!g553) & (g604) & (g3210) & (g3260)) + ((g553) & (!g604) & (!g3210) & (!g3260)) + ((g553) & (!g604) & (!g3210) & (g3260)) + ((g553) & (!g604) & (g3210) & (!g3260)) + ((g553) & (g604) & (!g3210) & (!g3260)));
	assign g3311 = (((!g3209) & (!g3272) & (!g3278) & (g3310)) + ((!g3209) & (g3272) & (!g3278) & (g3310)) + ((!g3209) & (g3272) & (g3278) & (g3310)) + ((g3209) & (!g3272) & (!g3278) & (!g3310)) + ((g3209) & (!g3272) & (g3278) & (!g3310)) + ((g3209) & (!g3272) & (g3278) & (g3310)) + ((g3209) & (g3272) & (!g3278) & (!g3310)) + ((g3209) & (g3272) & (g3278) & (!g3310)));
	assign g3312 = (((!g604) & (!g3210) & (g3260) & (!g3272) & (!g3278)) + ((!g604) & (!g3210) & (g3260) & (g3272) & (!g3278)) + ((!g604) & (!g3210) & (g3260) & (g3272) & (g3278)) + ((!g604) & (g3210) & (!g3260) & (!g3272) & (!g3278)) + ((!g604) & (g3210) & (!g3260) & (!g3272) & (g3278)) + ((!g604) & (g3210) & (!g3260) & (g3272) & (!g3278)) + ((!g604) & (g3210) & (!g3260) & (g3272) & (g3278)) + ((!g604) & (g3210) & (g3260) & (!g3272) & (g3278)) + ((g604) & (!g3210) & (!g3260) & (!g3272) & (!g3278)) + ((g604) & (!g3210) & (!g3260) & (g3272) & (!g3278)) + ((g604) & (!g3210) & (!g3260) & (g3272) & (g3278)) + ((g604) & (g3210) & (!g3260) & (!g3272) & (g3278)) + ((g604) & (g3210) & (g3260) & (!g3272) & (!g3278)) + ((g604) & (g3210) & (g3260) & (!g3272) & (g3278)) + ((g604) & (g3210) & (g3260) & (g3272) & (!g3278)) + ((g604) & (g3210) & (g3260) & (g3272) & (g3278)));
	assign g3313 = (((!g645) & (!g700) & (g3212) & (g3259)) + ((!g645) & (g700) & (!g3212) & (g3259)) + ((!g645) & (g700) & (g3212) & (!g3259)) + ((!g645) & (g700) & (g3212) & (g3259)) + ((g645) & (!g700) & (!g3212) & (!g3259)) + ((g645) & (!g700) & (!g3212) & (g3259)) + ((g645) & (!g700) & (g3212) & (!g3259)) + ((g645) & (g700) & (!g3212) & (!g3259)));
	assign g3314 = (((!g3211) & (!g3272) & (!g3278) & (g3313)) + ((!g3211) & (g3272) & (!g3278) & (g3313)) + ((!g3211) & (g3272) & (g3278) & (g3313)) + ((g3211) & (!g3272) & (!g3278) & (!g3313)) + ((g3211) & (!g3272) & (g3278) & (!g3313)) + ((g3211) & (!g3272) & (g3278) & (g3313)) + ((g3211) & (g3272) & (!g3278) & (!g3313)) + ((g3211) & (g3272) & (g3278) & (!g3313)));
	assign g3315 = (((!g700) & (!g3212) & (g3259) & (!g3272) & (!g3278)) + ((!g700) & (!g3212) & (g3259) & (g3272) & (!g3278)) + ((!g700) & (!g3212) & (g3259) & (g3272) & (g3278)) + ((!g700) & (g3212) & (!g3259) & (!g3272) & (!g3278)) + ((!g700) & (g3212) & (!g3259) & (!g3272) & (g3278)) + ((!g700) & (g3212) & (!g3259) & (g3272) & (!g3278)) + ((!g700) & (g3212) & (!g3259) & (g3272) & (g3278)) + ((!g700) & (g3212) & (g3259) & (!g3272) & (g3278)) + ((g700) & (!g3212) & (!g3259) & (!g3272) & (!g3278)) + ((g700) & (!g3212) & (!g3259) & (g3272) & (!g3278)) + ((g700) & (!g3212) & (!g3259) & (g3272) & (g3278)) + ((g700) & (g3212) & (!g3259) & (!g3272) & (g3278)) + ((g700) & (g3212) & (g3259) & (!g3272) & (!g3278)) + ((g700) & (g3212) & (g3259) & (!g3272) & (g3278)) + ((g700) & (g3212) & (g3259) & (g3272) & (!g3278)) + ((g700) & (g3212) & (g3259) & (g3272) & (g3278)));
	assign g3316 = (((!g744) & (!g803) & (g3214) & (g3258)) + ((!g744) & (g803) & (!g3214) & (g3258)) + ((!g744) & (g803) & (g3214) & (!g3258)) + ((!g744) & (g803) & (g3214) & (g3258)) + ((g744) & (!g803) & (!g3214) & (!g3258)) + ((g744) & (!g803) & (!g3214) & (g3258)) + ((g744) & (!g803) & (g3214) & (!g3258)) + ((g744) & (g803) & (!g3214) & (!g3258)));
	assign g3317 = (((!g3213) & (!g3272) & (!g3278) & (g3316)) + ((!g3213) & (g3272) & (!g3278) & (g3316)) + ((!g3213) & (g3272) & (g3278) & (g3316)) + ((g3213) & (!g3272) & (!g3278) & (!g3316)) + ((g3213) & (!g3272) & (g3278) & (!g3316)) + ((g3213) & (!g3272) & (g3278) & (g3316)) + ((g3213) & (g3272) & (!g3278) & (!g3316)) + ((g3213) & (g3272) & (g3278) & (!g3316)));
	assign g3318 = (((!g803) & (!g3214) & (g3258) & (!g3272) & (!g3278)) + ((!g803) & (!g3214) & (g3258) & (g3272) & (!g3278)) + ((!g803) & (!g3214) & (g3258) & (g3272) & (g3278)) + ((!g803) & (g3214) & (!g3258) & (!g3272) & (!g3278)) + ((!g803) & (g3214) & (!g3258) & (!g3272) & (g3278)) + ((!g803) & (g3214) & (!g3258) & (g3272) & (!g3278)) + ((!g803) & (g3214) & (!g3258) & (g3272) & (g3278)) + ((!g803) & (g3214) & (g3258) & (!g3272) & (g3278)) + ((g803) & (!g3214) & (!g3258) & (!g3272) & (!g3278)) + ((g803) & (!g3214) & (!g3258) & (g3272) & (!g3278)) + ((g803) & (!g3214) & (!g3258) & (g3272) & (g3278)) + ((g803) & (g3214) & (!g3258) & (!g3272) & (g3278)) + ((g803) & (g3214) & (g3258) & (!g3272) & (!g3278)) + ((g803) & (g3214) & (g3258) & (!g3272) & (g3278)) + ((g803) & (g3214) & (g3258) & (g3272) & (!g3278)) + ((g803) & (g3214) & (g3258) & (g3272) & (g3278)));
	assign g3319 = (((!g851) & (!g914) & (g3216) & (g3257)) + ((!g851) & (g914) & (!g3216) & (g3257)) + ((!g851) & (g914) & (g3216) & (!g3257)) + ((!g851) & (g914) & (g3216) & (g3257)) + ((g851) & (!g914) & (!g3216) & (!g3257)) + ((g851) & (!g914) & (!g3216) & (g3257)) + ((g851) & (!g914) & (g3216) & (!g3257)) + ((g851) & (g914) & (!g3216) & (!g3257)));
	assign g3320 = (((!g3215) & (!g3272) & (!g3278) & (g3319)) + ((!g3215) & (g3272) & (!g3278) & (g3319)) + ((!g3215) & (g3272) & (g3278) & (g3319)) + ((g3215) & (!g3272) & (!g3278) & (!g3319)) + ((g3215) & (!g3272) & (g3278) & (!g3319)) + ((g3215) & (!g3272) & (g3278) & (g3319)) + ((g3215) & (g3272) & (!g3278) & (!g3319)) + ((g3215) & (g3272) & (g3278) & (!g3319)));
	assign g3321 = (((!g914) & (!g3216) & (g3257) & (!g3272) & (!g3278)) + ((!g914) & (!g3216) & (g3257) & (g3272) & (!g3278)) + ((!g914) & (!g3216) & (g3257) & (g3272) & (g3278)) + ((!g914) & (g3216) & (!g3257) & (!g3272) & (!g3278)) + ((!g914) & (g3216) & (!g3257) & (!g3272) & (g3278)) + ((!g914) & (g3216) & (!g3257) & (g3272) & (!g3278)) + ((!g914) & (g3216) & (!g3257) & (g3272) & (g3278)) + ((!g914) & (g3216) & (g3257) & (!g3272) & (g3278)) + ((g914) & (!g3216) & (!g3257) & (!g3272) & (!g3278)) + ((g914) & (!g3216) & (!g3257) & (g3272) & (!g3278)) + ((g914) & (!g3216) & (!g3257) & (g3272) & (g3278)) + ((g914) & (g3216) & (!g3257) & (!g3272) & (g3278)) + ((g914) & (g3216) & (g3257) & (!g3272) & (!g3278)) + ((g914) & (g3216) & (g3257) & (!g3272) & (g3278)) + ((g914) & (g3216) & (g3257) & (g3272) & (!g3278)) + ((g914) & (g3216) & (g3257) & (g3272) & (g3278)));
	assign g3322 = (((!g1032) & (!g1030) & (g3218) & (g3256)) + ((!g1032) & (g1030) & (!g3218) & (g3256)) + ((!g1032) & (g1030) & (g3218) & (!g3256)) + ((!g1032) & (g1030) & (g3218) & (g3256)) + ((g1032) & (!g1030) & (!g3218) & (!g3256)) + ((g1032) & (!g1030) & (!g3218) & (g3256)) + ((g1032) & (!g1030) & (g3218) & (!g3256)) + ((g1032) & (g1030) & (!g3218) & (!g3256)));
	assign g3323 = (((!g3217) & (!g3272) & (!g3278) & (g3322)) + ((!g3217) & (g3272) & (!g3278) & (g3322)) + ((!g3217) & (g3272) & (g3278) & (g3322)) + ((g3217) & (!g3272) & (!g3278) & (!g3322)) + ((g3217) & (!g3272) & (g3278) & (!g3322)) + ((g3217) & (!g3272) & (g3278) & (g3322)) + ((g3217) & (g3272) & (!g3278) & (!g3322)) + ((g3217) & (g3272) & (g3278) & (!g3322)));
	assign g3324 = (((!g1030) & (!g3218) & (g3256) & (!g3272) & (!g3278)) + ((!g1030) & (!g3218) & (g3256) & (g3272) & (!g3278)) + ((!g1030) & (!g3218) & (g3256) & (g3272) & (g3278)) + ((!g1030) & (g3218) & (!g3256) & (!g3272) & (!g3278)) + ((!g1030) & (g3218) & (!g3256) & (!g3272) & (g3278)) + ((!g1030) & (g3218) & (!g3256) & (g3272) & (!g3278)) + ((!g1030) & (g3218) & (!g3256) & (g3272) & (g3278)) + ((!g1030) & (g3218) & (g3256) & (!g3272) & (g3278)) + ((g1030) & (!g3218) & (!g3256) & (!g3272) & (!g3278)) + ((g1030) & (!g3218) & (!g3256) & (g3272) & (!g3278)) + ((g1030) & (!g3218) & (!g3256) & (g3272) & (g3278)) + ((g1030) & (g3218) & (!g3256) & (!g3272) & (g3278)) + ((g1030) & (g3218) & (g3256) & (!g3272) & (!g3278)) + ((g1030) & (g3218) & (g3256) & (!g3272) & (g3278)) + ((g1030) & (g3218) & (g3256) & (g3272) & (!g3278)) + ((g1030) & (g3218) & (g3256) & (g3272) & (g3278)));
	assign g3325 = (((!g1160) & (!g1154) & (g3220) & (g3255)) + ((!g1160) & (g1154) & (!g3220) & (g3255)) + ((!g1160) & (g1154) & (g3220) & (!g3255)) + ((!g1160) & (g1154) & (g3220) & (g3255)) + ((g1160) & (!g1154) & (!g3220) & (!g3255)) + ((g1160) & (!g1154) & (!g3220) & (g3255)) + ((g1160) & (!g1154) & (g3220) & (!g3255)) + ((g1160) & (g1154) & (!g3220) & (!g3255)));
	assign g3326 = (((!g3219) & (!g3272) & (!g3278) & (g3325)) + ((!g3219) & (g3272) & (!g3278) & (g3325)) + ((!g3219) & (g3272) & (g3278) & (g3325)) + ((g3219) & (!g3272) & (!g3278) & (!g3325)) + ((g3219) & (!g3272) & (g3278) & (!g3325)) + ((g3219) & (!g3272) & (g3278) & (g3325)) + ((g3219) & (g3272) & (!g3278) & (!g3325)) + ((g3219) & (g3272) & (g3278) & (!g3325)));
	assign g3327 = (((!g1154) & (!g3220) & (g3255) & (!g3272) & (!g3278)) + ((!g1154) & (!g3220) & (g3255) & (g3272) & (!g3278)) + ((!g1154) & (!g3220) & (g3255) & (g3272) & (g3278)) + ((!g1154) & (g3220) & (!g3255) & (!g3272) & (!g3278)) + ((!g1154) & (g3220) & (!g3255) & (!g3272) & (g3278)) + ((!g1154) & (g3220) & (!g3255) & (g3272) & (!g3278)) + ((!g1154) & (g3220) & (!g3255) & (g3272) & (g3278)) + ((!g1154) & (g3220) & (g3255) & (!g3272) & (g3278)) + ((g1154) & (!g3220) & (!g3255) & (!g3272) & (!g3278)) + ((g1154) & (!g3220) & (!g3255) & (g3272) & (!g3278)) + ((g1154) & (!g3220) & (!g3255) & (g3272) & (g3278)) + ((g1154) & (g3220) & (!g3255) & (!g3272) & (g3278)) + ((g1154) & (g3220) & (g3255) & (!g3272) & (!g3278)) + ((g1154) & (g3220) & (g3255) & (!g3272) & (g3278)) + ((g1154) & (g3220) & (g3255) & (g3272) & (!g3278)) + ((g1154) & (g3220) & (g3255) & (g3272) & (g3278)));
	assign g3328 = (((!g1295) & (!g1285) & (g3222) & (g3254)) + ((!g1295) & (g1285) & (!g3222) & (g3254)) + ((!g1295) & (g1285) & (g3222) & (!g3254)) + ((!g1295) & (g1285) & (g3222) & (g3254)) + ((g1295) & (!g1285) & (!g3222) & (!g3254)) + ((g1295) & (!g1285) & (!g3222) & (g3254)) + ((g1295) & (!g1285) & (g3222) & (!g3254)) + ((g1295) & (g1285) & (!g3222) & (!g3254)));
	assign g3329 = (((!g3221) & (!g3272) & (!g3278) & (g3328)) + ((!g3221) & (g3272) & (!g3278) & (g3328)) + ((!g3221) & (g3272) & (g3278) & (g3328)) + ((g3221) & (!g3272) & (!g3278) & (!g3328)) + ((g3221) & (!g3272) & (g3278) & (!g3328)) + ((g3221) & (!g3272) & (g3278) & (g3328)) + ((g3221) & (g3272) & (!g3278) & (!g3328)) + ((g3221) & (g3272) & (g3278) & (!g3328)));
	assign g3330 = (((!g1285) & (!g3222) & (g3254) & (!g3272) & (!g3278)) + ((!g1285) & (!g3222) & (g3254) & (g3272) & (!g3278)) + ((!g1285) & (!g3222) & (g3254) & (g3272) & (g3278)) + ((!g1285) & (g3222) & (!g3254) & (!g3272) & (!g3278)) + ((!g1285) & (g3222) & (!g3254) & (!g3272) & (g3278)) + ((!g1285) & (g3222) & (!g3254) & (g3272) & (!g3278)) + ((!g1285) & (g3222) & (!g3254) & (g3272) & (g3278)) + ((!g1285) & (g3222) & (g3254) & (!g3272) & (g3278)) + ((g1285) & (!g3222) & (!g3254) & (!g3272) & (!g3278)) + ((g1285) & (!g3222) & (!g3254) & (g3272) & (!g3278)) + ((g1285) & (!g3222) & (!g3254) & (g3272) & (g3278)) + ((g1285) & (g3222) & (!g3254) & (!g3272) & (g3278)) + ((g1285) & (g3222) & (g3254) & (!g3272) & (!g3278)) + ((g1285) & (g3222) & (g3254) & (!g3272) & (g3278)) + ((g1285) & (g3222) & (g3254) & (g3272) & (!g3278)) + ((g1285) & (g3222) & (g3254) & (g3272) & (g3278)));
	assign g3331 = (((!g1437) & (!g1423) & (g3224) & (g3253)) + ((!g1437) & (g1423) & (!g3224) & (g3253)) + ((!g1437) & (g1423) & (g3224) & (!g3253)) + ((!g1437) & (g1423) & (g3224) & (g3253)) + ((g1437) & (!g1423) & (!g3224) & (!g3253)) + ((g1437) & (!g1423) & (!g3224) & (g3253)) + ((g1437) & (!g1423) & (g3224) & (!g3253)) + ((g1437) & (g1423) & (!g3224) & (!g3253)));
	assign g3332 = (((!g3223) & (!g3272) & (!g3278) & (g3331)) + ((!g3223) & (g3272) & (!g3278) & (g3331)) + ((!g3223) & (g3272) & (g3278) & (g3331)) + ((g3223) & (!g3272) & (!g3278) & (!g3331)) + ((g3223) & (!g3272) & (g3278) & (!g3331)) + ((g3223) & (!g3272) & (g3278) & (g3331)) + ((g3223) & (g3272) & (!g3278) & (!g3331)) + ((g3223) & (g3272) & (g3278) & (!g3331)));
	assign g3333 = (((!g1423) & (!g3224) & (g3253) & (!g3272) & (!g3278)) + ((!g1423) & (!g3224) & (g3253) & (g3272) & (!g3278)) + ((!g1423) & (!g3224) & (g3253) & (g3272) & (g3278)) + ((!g1423) & (g3224) & (!g3253) & (!g3272) & (!g3278)) + ((!g1423) & (g3224) & (!g3253) & (!g3272) & (g3278)) + ((!g1423) & (g3224) & (!g3253) & (g3272) & (!g3278)) + ((!g1423) & (g3224) & (!g3253) & (g3272) & (g3278)) + ((!g1423) & (g3224) & (g3253) & (!g3272) & (g3278)) + ((g1423) & (!g3224) & (!g3253) & (!g3272) & (!g3278)) + ((g1423) & (!g3224) & (!g3253) & (g3272) & (!g3278)) + ((g1423) & (!g3224) & (!g3253) & (g3272) & (g3278)) + ((g1423) & (g3224) & (!g3253) & (!g3272) & (g3278)) + ((g1423) & (g3224) & (g3253) & (!g3272) & (!g3278)) + ((g1423) & (g3224) & (g3253) & (!g3272) & (g3278)) + ((g1423) & (g3224) & (g3253) & (g3272) & (!g3278)) + ((g1423) & (g3224) & (g3253) & (g3272) & (g3278)));
	assign g3334 = (((!g1586) & (!g1568) & (g3226) & (g3252)) + ((!g1586) & (g1568) & (!g3226) & (g3252)) + ((!g1586) & (g1568) & (g3226) & (!g3252)) + ((!g1586) & (g1568) & (g3226) & (g3252)) + ((g1586) & (!g1568) & (!g3226) & (!g3252)) + ((g1586) & (!g1568) & (!g3226) & (g3252)) + ((g1586) & (!g1568) & (g3226) & (!g3252)) + ((g1586) & (g1568) & (!g3226) & (!g3252)));
	assign g3335 = (((!g3225) & (!g3272) & (!g3278) & (g3334)) + ((!g3225) & (g3272) & (!g3278) & (g3334)) + ((!g3225) & (g3272) & (g3278) & (g3334)) + ((g3225) & (!g3272) & (!g3278) & (!g3334)) + ((g3225) & (!g3272) & (g3278) & (!g3334)) + ((g3225) & (!g3272) & (g3278) & (g3334)) + ((g3225) & (g3272) & (!g3278) & (!g3334)) + ((g3225) & (g3272) & (g3278) & (!g3334)));
	assign g3336 = (((!g1568) & (!g3226) & (g3252) & (!g3272) & (!g3278)) + ((!g1568) & (!g3226) & (g3252) & (g3272) & (!g3278)) + ((!g1568) & (!g3226) & (g3252) & (g3272) & (g3278)) + ((!g1568) & (g3226) & (!g3252) & (!g3272) & (!g3278)) + ((!g1568) & (g3226) & (!g3252) & (!g3272) & (g3278)) + ((!g1568) & (g3226) & (!g3252) & (g3272) & (!g3278)) + ((!g1568) & (g3226) & (!g3252) & (g3272) & (g3278)) + ((!g1568) & (g3226) & (g3252) & (!g3272) & (g3278)) + ((g1568) & (!g3226) & (!g3252) & (!g3272) & (!g3278)) + ((g1568) & (!g3226) & (!g3252) & (g3272) & (!g3278)) + ((g1568) & (!g3226) & (!g3252) & (g3272) & (g3278)) + ((g1568) & (g3226) & (!g3252) & (!g3272) & (g3278)) + ((g1568) & (g3226) & (g3252) & (!g3272) & (!g3278)) + ((g1568) & (g3226) & (g3252) & (!g3272) & (g3278)) + ((g1568) & (g3226) & (g3252) & (g3272) & (!g3278)) + ((g1568) & (g3226) & (g3252) & (g3272) & (g3278)));
	assign g3337 = (((!g1742) & (!g1720) & (g3228) & (g3251)) + ((!g1742) & (g1720) & (!g3228) & (g3251)) + ((!g1742) & (g1720) & (g3228) & (!g3251)) + ((!g1742) & (g1720) & (g3228) & (g3251)) + ((g1742) & (!g1720) & (!g3228) & (!g3251)) + ((g1742) & (!g1720) & (!g3228) & (g3251)) + ((g1742) & (!g1720) & (g3228) & (!g3251)) + ((g1742) & (g1720) & (!g3228) & (!g3251)));
	assign g3338 = (((!g3227) & (!g3272) & (!g3278) & (g3337)) + ((!g3227) & (g3272) & (!g3278) & (g3337)) + ((!g3227) & (g3272) & (g3278) & (g3337)) + ((g3227) & (!g3272) & (!g3278) & (!g3337)) + ((g3227) & (!g3272) & (g3278) & (!g3337)) + ((g3227) & (!g3272) & (g3278) & (g3337)) + ((g3227) & (g3272) & (!g3278) & (!g3337)) + ((g3227) & (g3272) & (g3278) & (!g3337)));
	assign g3339 = (((!g1720) & (!g3228) & (g3251) & (!g3272) & (!g3278)) + ((!g1720) & (!g3228) & (g3251) & (g3272) & (!g3278)) + ((!g1720) & (!g3228) & (g3251) & (g3272) & (g3278)) + ((!g1720) & (g3228) & (!g3251) & (!g3272) & (!g3278)) + ((!g1720) & (g3228) & (!g3251) & (!g3272) & (g3278)) + ((!g1720) & (g3228) & (!g3251) & (g3272) & (!g3278)) + ((!g1720) & (g3228) & (!g3251) & (g3272) & (g3278)) + ((!g1720) & (g3228) & (g3251) & (!g3272) & (g3278)) + ((g1720) & (!g3228) & (!g3251) & (!g3272) & (!g3278)) + ((g1720) & (!g3228) & (!g3251) & (g3272) & (!g3278)) + ((g1720) & (!g3228) & (!g3251) & (g3272) & (g3278)) + ((g1720) & (g3228) & (!g3251) & (!g3272) & (g3278)) + ((g1720) & (g3228) & (g3251) & (!g3272) & (!g3278)) + ((g1720) & (g3228) & (g3251) & (!g3272) & (g3278)) + ((g1720) & (g3228) & (g3251) & (g3272) & (!g3278)) + ((g1720) & (g3228) & (g3251) & (g3272) & (g3278)));
	assign g3340 = (((!g1905) & (!g1879) & (g3230) & (g3250)) + ((!g1905) & (g1879) & (!g3230) & (g3250)) + ((!g1905) & (g1879) & (g3230) & (!g3250)) + ((!g1905) & (g1879) & (g3230) & (g3250)) + ((g1905) & (!g1879) & (!g3230) & (!g3250)) + ((g1905) & (!g1879) & (!g3230) & (g3250)) + ((g1905) & (!g1879) & (g3230) & (!g3250)) + ((g1905) & (g1879) & (!g3230) & (!g3250)));
	assign g3341 = (((!g3229) & (!g3272) & (!g3278) & (g3340)) + ((!g3229) & (g3272) & (!g3278) & (g3340)) + ((!g3229) & (g3272) & (g3278) & (g3340)) + ((g3229) & (!g3272) & (!g3278) & (!g3340)) + ((g3229) & (!g3272) & (g3278) & (!g3340)) + ((g3229) & (!g3272) & (g3278) & (g3340)) + ((g3229) & (g3272) & (!g3278) & (!g3340)) + ((g3229) & (g3272) & (g3278) & (!g3340)));
	assign g3342 = (((!g1879) & (!g3230) & (g3250) & (!g3272) & (!g3278)) + ((!g1879) & (!g3230) & (g3250) & (g3272) & (!g3278)) + ((!g1879) & (!g3230) & (g3250) & (g3272) & (g3278)) + ((!g1879) & (g3230) & (!g3250) & (!g3272) & (!g3278)) + ((!g1879) & (g3230) & (!g3250) & (!g3272) & (g3278)) + ((!g1879) & (g3230) & (!g3250) & (g3272) & (!g3278)) + ((!g1879) & (g3230) & (!g3250) & (g3272) & (g3278)) + ((!g1879) & (g3230) & (g3250) & (!g3272) & (g3278)) + ((g1879) & (!g3230) & (!g3250) & (!g3272) & (!g3278)) + ((g1879) & (!g3230) & (!g3250) & (g3272) & (!g3278)) + ((g1879) & (!g3230) & (!g3250) & (g3272) & (g3278)) + ((g1879) & (g3230) & (!g3250) & (!g3272) & (g3278)) + ((g1879) & (g3230) & (g3250) & (!g3272) & (!g3278)) + ((g1879) & (g3230) & (g3250) & (!g3272) & (g3278)) + ((g1879) & (g3230) & (g3250) & (g3272) & (!g3278)) + ((g1879) & (g3230) & (g3250) & (g3272) & (g3278)));
	assign g3343 = (((!g2075) & (!g2045) & (g3232) & (g3249)) + ((!g2075) & (g2045) & (!g3232) & (g3249)) + ((!g2075) & (g2045) & (g3232) & (!g3249)) + ((!g2075) & (g2045) & (g3232) & (g3249)) + ((g2075) & (!g2045) & (!g3232) & (!g3249)) + ((g2075) & (!g2045) & (!g3232) & (g3249)) + ((g2075) & (!g2045) & (g3232) & (!g3249)) + ((g2075) & (g2045) & (!g3232) & (!g3249)));
	assign g3344 = (((!g3231) & (!g3272) & (!g3278) & (g3343)) + ((!g3231) & (g3272) & (!g3278) & (g3343)) + ((!g3231) & (g3272) & (g3278) & (g3343)) + ((g3231) & (!g3272) & (!g3278) & (!g3343)) + ((g3231) & (!g3272) & (g3278) & (!g3343)) + ((g3231) & (!g3272) & (g3278) & (g3343)) + ((g3231) & (g3272) & (!g3278) & (!g3343)) + ((g3231) & (g3272) & (g3278) & (!g3343)));
	assign g3345 = (((!g2045) & (!g3232) & (g3249) & (!g3272) & (!g3278)) + ((!g2045) & (!g3232) & (g3249) & (g3272) & (!g3278)) + ((!g2045) & (!g3232) & (g3249) & (g3272) & (g3278)) + ((!g2045) & (g3232) & (!g3249) & (!g3272) & (!g3278)) + ((!g2045) & (g3232) & (!g3249) & (!g3272) & (g3278)) + ((!g2045) & (g3232) & (!g3249) & (g3272) & (!g3278)) + ((!g2045) & (g3232) & (!g3249) & (g3272) & (g3278)) + ((!g2045) & (g3232) & (g3249) & (!g3272) & (g3278)) + ((g2045) & (!g3232) & (!g3249) & (!g3272) & (!g3278)) + ((g2045) & (!g3232) & (!g3249) & (g3272) & (!g3278)) + ((g2045) & (!g3232) & (!g3249) & (g3272) & (g3278)) + ((g2045) & (g3232) & (!g3249) & (!g3272) & (g3278)) + ((g2045) & (g3232) & (g3249) & (!g3272) & (!g3278)) + ((g2045) & (g3232) & (g3249) & (!g3272) & (g3278)) + ((g2045) & (g3232) & (g3249) & (g3272) & (!g3278)) + ((g2045) & (g3232) & (g3249) & (g3272) & (g3278)));
	assign g3346 = (((!g2252) & (!g2218) & (g3234) & (g3248)) + ((!g2252) & (g2218) & (!g3234) & (g3248)) + ((!g2252) & (g2218) & (g3234) & (!g3248)) + ((!g2252) & (g2218) & (g3234) & (g3248)) + ((g2252) & (!g2218) & (!g3234) & (!g3248)) + ((g2252) & (!g2218) & (!g3234) & (g3248)) + ((g2252) & (!g2218) & (g3234) & (!g3248)) + ((g2252) & (g2218) & (!g3234) & (!g3248)));
	assign g3347 = (((!g3233) & (!g3272) & (!g3278) & (g3346)) + ((!g3233) & (g3272) & (!g3278) & (g3346)) + ((!g3233) & (g3272) & (g3278) & (g3346)) + ((g3233) & (!g3272) & (!g3278) & (!g3346)) + ((g3233) & (!g3272) & (g3278) & (!g3346)) + ((g3233) & (!g3272) & (g3278) & (g3346)) + ((g3233) & (g3272) & (!g3278) & (!g3346)) + ((g3233) & (g3272) & (g3278) & (!g3346)));
	assign g3348 = (((!g2218) & (!g3234) & (g3248) & (!g3272) & (!g3278)) + ((!g2218) & (!g3234) & (g3248) & (g3272) & (!g3278)) + ((!g2218) & (!g3234) & (g3248) & (g3272) & (g3278)) + ((!g2218) & (g3234) & (!g3248) & (!g3272) & (!g3278)) + ((!g2218) & (g3234) & (!g3248) & (!g3272) & (g3278)) + ((!g2218) & (g3234) & (!g3248) & (g3272) & (!g3278)) + ((!g2218) & (g3234) & (!g3248) & (g3272) & (g3278)) + ((!g2218) & (g3234) & (g3248) & (!g3272) & (g3278)) + ((g2218) & (!g3234) & (!g3248) & (!g3272) & (!g3278)) + ((g2218) & (!g3234) & (!g3248) & (g3272) & (!g3278)) + ((g2218) & (!g3234) & (!g3248) & (g3272) & (g3278)) + ((g2218) & (g3234) & (!g3248) & (!g3272) & (g3278)) + ((g2218) & (g3234) & (g3248) & (!g3272) & (!g3278)) + ((g2218) & (g3234) & (g3248) & (!g3272) & (g3278)) + ((g2218) & (g3234) & (g3248) & (g3272) & (!g3278)) + ((g2218) & (g3234) & (g3248) & (g3272) & (g3278)));
	assign g3349 = (((!g2436) & (!g2398) & (g3236) & (g3247)) + ((!g2436) & (g2398) & (!g3236) & (g3247)) + ((!g2436) & (g2398) & (g3236) & (!g3247)) + ((!g2436) & (g2398) & (g3236) & (g3247)) + ((g2436) & (!g2398) & (!g3236) & (!g3247)) + ((g2436) & (!g2398) & (!g3236) & (g3247)) + ((g2436) & (!g2398) & (g3236) & (!g3247)) + ((g2436) & (g2398) & (!g3236) & (!g3247)));
	assign g3350 = (((!g3235) & (!g3272) & (!g3278) & (g3349)) + ((!g3235) & (g3272) & (!g3278) & (g3349)) + ((!g3235) & (g3272) & (g3278) & (g3349)) + ((g3235) & (!g3272) & (!g3278) & (!g3349)) + ((g3235) & (!g3272) & (g3278) & (!g3349)) + ((g3235) & (!g3272) & (g3278) & (g3349)) + ((g3235) & (g3272) & (!g3278) & (!g3349)) + ((g3235) & (g3272) & (g3278) & (!g3349)));
	assign g3351 = (((!g2398) & (!g3236) & (g3247) & (!g3272) & (!g3278)) + ((!g2398) & (!g3236) & (g3247) & (g3272) & (!g3278)) + ((!g2398) & (!g3236) & (g3247) & (g3272) & (g3278)) + ((!g2398) & (g3236) & (!g3247) & (!g3272) & (!g3278)) + ((!g2398) & (g3236) & (!g3247) & (!g3272) & (g3278)) + ((!g2398) & (g3236) & (!g3247) & (g3272) & (!g3278)) + ((!g2398) & (g3236) & (!g3247) & (g3272) & (g3278)) + ((!g2398) & (g3236) & (g3247) & (!g3272) & (g3278)) + ((g2398) & (!g3236) & (!g3247) & (!g3272) & (!g3278)) + ((g2398) & (!g3236) & (!g3247) & (g3272) & (!g3278)) + ((g2398) & (!g3236) & (!g3247) & (g3272) & (g3278)) + ((g2398) & (g3236) & (!g3247) & (!g3272) & (g3278)) + ((g2398) & (g3236) & (g3247) & (!g3272) & (!g3278)) + ((g2398) & (g3236) & (g3247) & (!g3272) & (g3278)) + ((g2398) & (g3236) & (g3247) & (g3272) & (!g3278)) + ((g2398) & (g3236) & (g3247) & (g3272) & (g3278)));
	assign g3352 = (((!g2627) & (!g2585) & (g3238) & (g3246)) + ((!g2627) & (g2585) & (!g3238) & (g3246)) + ((!g2627) & (g2585) & (g3238) & (!g3246)) + ((!g2627) & (g2585) & (g3238) & (g3246)) + ((g2627) & (!g2585) & (!g3238) & (!g3246)) + ((g2627) & (!g2585) & (!g3238) & (g3246)) + ((g2627) & (!g2585) & (g3238) & (!g3246)) + ((g2627) & (g2585) & (!g3238) & (!g3246)));
	assign g3353 = (((!g3237) & (!g3272) & (!g3278) & (g3352)) + ((!g3237) & (g3272) & (!g3278) & (g3352)) + ((!g3237) & (g3272) & (g3278) & (g3352)) + ((g3237) & (!g3272) & (!g3278) & (!g3352)) + ((g3237) & (!g3272) & (g3278) & (!g3352)) + ((g3237) & (!g3272) & (g3278) & (g3352)) + ((g3237) & (g3272) & (!g3278) & (!g3352)) + ((g3237) & (g3272) & (g3278) & (!g3352)));
	assign g3354 = (((!g2585) & (!g3238) & (g3246) & (!g3272) & (!g3278)) + ((!g2585) & (!g3238) & (g3246) & (g3272) & (!g3278)) + ((!g2585) & (!g3238) & (g3246) & (g3272) & (g3278)) + ((!g2585) & (g3238) & (!g3246) & (!g3272) & (!g3278)) + ((!g2585) & (g3238) & (!g3246) & (!g3272) & (g3278)) + ((!g2585) & (g3238) & (!g3246) & (g3272) & (!g3278)) + ((!g2585) & (g3238) & (!g3246) & (g3272) & (g3278)) + ((!g2585) & (g3238) & (g3246) & (!g3272) & (g3278)) + ((g2585) & (!g3238) & (!g3246) & (!g3272) & (!g3278)) + ((g2585) & (!g3238) & (!g3246) & (g3272) & (!g3278)) + ((g2585) & (!g3238) & (!g3246) & (g3272) & (g3278)) + ((g2585) & (g3238) & (!g3246) & (!g3272) & (g3278)) + ((g2585) & (g3238) & (g3246) & (!g3272) & (!g3278)) + ((g2585) & (g3238) & (g3246) & (!g3272) & (g3278)) + ((g2585) & (g3238) & (g3246) & (g3272) & (!g3278)) + ((g2585) & (g3238) & (g3246) & (g3272) & (g3278)));
	assign g3355 = (((!g2825) & (!g2779) & (g3240) & (g3245)) + ((!g2825) & (g2779) & (!g3240) & (g3245)) + ((!g2825) & (g2779) & (g3240) & (!g3245)) + ((!g2825) & (g2779) & (g3240) & (g3245)) + ((g2825) & (!g2779) & (!g3240) & (!g3245)) + ((g2825) & (!g2779) & (!g3240) & (g3245)) + ((g2825) & (!g2779) & (g3240) & (!g3245)) + ((g2825) & (g2779) & (!g3240) & (!g3245)));
	assign g3356 = (((!g3239) & (!g3272) & (!g3278) & (g3355)) + ((!g3239) & (g3272) & (!g3278) & (g3355)) + ((!g3239) & (g3272) & (g3278) & (g3355)) + ((g3239) & (!g3272) & (!g3278) & (!g3355)) + ((g3239) & (!g3272) & (g3278) & (!g3355)) + ((g3239) & (!g3272) & (g3278) & (g3355)) + ((g3239) & (g3272) & (!g3278) & (!g3355)) + ((g3239) & (g3272) & (g3278) & (!g3355)));
	assign g3357 = (((!g2779) & (!g3240) & (g3245) & (!g3272) & (!g3278)) + ((!g2779) & (!g3240) & (g3245) & (g3272) & (!g3278)) + ((!g2779) & (!g3240) & (g3245) & (g3272) & (g3278)) + ((!g2779) & (g3240) & (!g3245) & (!g3272) & (!g3278)) + ((!g2779) & (g3240) & (!g3245) & (!g3272) & (g3278)) + ((!g2779) & (g3240) & (!g3245) & (g3272) & (!g3278)) + ((!g2779) & (g3240) & (!g3245) & (g3272) & (g3278)) + ((!g2779) & (g3240) & (g3245) & (!g3272) & (g3278)) + ((g2779) & (!g3240) & (!g3245) & (!g3272) & (!g3278)) + ((g2779) & (!g3240) & (!g3245) & (g3272) & (!g3278)) + ((g2779) & (!g3240) & (!g3245) & (g3272) & (g3278)) + ((g2779) & (g3240) & (!g3245) & (!g3272) & (g3278)) + ((g2779) & (g3240) & (g3245) & (!g3272) & (!g3278)) + ((g2779) & (g3240) & (g3245) & (!g3272) & (g3278)) + ((g2779) & (g3240) & (g3245) & (g3272) & (!g3278)) + ((g2779) & (g3240) & (g3245) & (g3272) & (g3278)));
	assign g3358 = (((!g3030) & (!g2980) & (g3242) & (g3244)) + ((!g3030) & (g2980) & (!g3242) & (g3244)) + ((!g3030) & (g2980) & (g3242) & (!g3244)) + ((!g3030) & (g2980) & (g3242) & (g3244)) + ((g3030) & (!g2980) & (!g3242) & (!g3244)) + ((g3030) & (!g2980) & (!g3242) & (g3244)) + ((g3030) & (!g2980) & (g3242) & (!g3244)) + ((g3030) & (g2980) & (!g3242) & (!g3244)));
	assign g3359 = (((!g3241) & (!g3272) & (!g3278) & (g3358)) + ((!g3241) & (g3272) & (!g3278) & (g3358)) + ((!g3241) & (g3272) & (g3278) & (g3358)) + ((g3241) & (!g3272) & (!g3278) & (!g3358)) + ((g3241) & (!g3272) & (g3278) & (!g3358)) + ((g3241) & (!g3272) & (g3278) & (g3358)) + ((g3241) & (g3272) & (!g3278) & (!g3358)) + ((g3241) & (g3272) & (g3278) & (!g3358)));
	assign g3360 = (((!g2980) & (!g3242) & (g3244) & (!g3272) & (!g3278)) + ((!g2980) & (!g3242) & (g3244) & (g3272) & (!g3278)) + ((!g2980) & (!g3242) & (g3244) & (g3272) & (g3278)) + ((!g2980) & (g3242) & (!g3244) & (!g3272) & (!g3278)) + ((!g2980) & (g3242) & (!g3244) & (!g3272) & (g3278)) + ((!g2980) & (g3242) & (!g3244) & (g3272) & (!g3278)) + ((!g2980) & (g3242) & (!g3244) & (g3272) & (g3278)) + ((!g2980) & (g3242) & (g3244) & (!g3272) & (g3278)) + ((g2980) & (!g3242) & (!g3244) & (!g3272) & (!g3278)) + ((g2980) & (!g3242) & (!g3244) & (g3272) & (!g3278)) + ((g2980) & (!g3242) & (!g3244) & (g3272) & (g3278)) + ((g2980) & (g3242) & (!g3244) & (!g3272) & (g3278)) + ((g2980) & (g3242) & (g3244) & (!g3272) & (!g3278)) + ((g2980) & (g3242) & (g3244) & (!g3272) & (g3278)) + ((g2980) & (g3242) & (g3244) & (g3272) & (!g3278)) + ((g2980) & (g3242) & (g3244) & (g3272) & (g3278)));
	assign g3361 = (((!g3178) & (!ax8x) & (!g3187) & (g3243)) + ((!g3178) & (!ax8x) & (g3187) & (g3243)) + ((!g3178) & (ax8x) & (!g3187) & (!g3243)) + ((!g3178) & (ax8x) & (!g3187) & (g3243)) + ((g3178) & (!ax8x) & (!g3187) & (!g3243)) + ((g3178) & (!ax8x) & (g3187) & (!g3243)) + ((g3178) & (ax8x) & (g3187) & (!g3243)) + ((g3178) & (ax8x) & (g3187) & (g3243)));
	assign g3362 = (((!ax8x) & (!ax9x) & (!g3187) & (!g3272) & (!g3278) & (g3361)) + ((!ax8x) & (!ax9x) & (!g3187) & (!g3272) & (g3278) & (!g3361)) + ((!ax8x) & (!ax9x) & (!g3187) & (!g3272) & (g3278) & (g3361)) + ((!ax8x) & (!ax9x) & (!g3187) & (g3272) & (!g3278) & (g3361)) + ((!ax8x) & (!ax9x) & (!g3187) & (g3272) & (g3278) & (g3361)) + ((!ax8x) & (!ax9x) & (g3187) & (!g3272) & (!g3278) & (!g3361)) + ((!ax8x) & (!ax9x) & (g3187) & (g3272) & (!g3278) & (!g3361)) + ((!ax8x) & (!ax9x) & (g3187) & (g3272) & (g3278) & (!g3361)) + ((!ax8x) & (ax9x) & (!g3187) & (!g3272) & (!g3278) & (!g3361)) + ((!ax8x) & (ax9x) & (!g3187) & (g3272) & (!g3278) & (!g3361)) + ((!ax8x) & (ax9x) & (!g3187) & (g3272) & (g3278) & (!g3361)) + ((!ax8x) & (ax9x) & (g3187) & (!g3272) & (!g3278) & (g3361)) + ((!ax8x) & (ax9x) & (g3187) & (!g3272) & (g3278) & (!g3361)) + ((!ax8x) & (ax9x) & (g3187) & (!g3272) & (g3278) & (g3361)) + ((!ax8x) & (ax9x) & (g3187) & (g3272) & (!g3278) & (g3361)) + ((!ax8x) & (ax9x) & (g3187) & (g3272) & (g3278) & (g3361)) + ((ax8x) & (!ax9x) & (!g3187) & (!g3272) & (!g3278) & (!g3361)) + ((ax8x) & (!ax9x) & (!g3187) & (g3272) & (!g3278) & (!g3361)) + ((ax8x) & (!ax9x) & (!g3187) & (g3272) & (g3278) & (!g3361)) + ((ax8x) & (!ax9x) & (g3187) & (!g3272) & (!g3278) & (!g3361)) + ((ax8x) & (!ax9x) & (g3187) & (g3272) & (!g3278) & (!g3361)) + ((ax8x) & (!ax9x) & (g3187) & (g3272) & (g3278) & (!g3361)) + ((ax8x) & (ax9x) & (!g3187) & (!g3272) & (!g3278) & (g3361)) + ((ax8x) & (ax9x) & (!g3187) & (!g3272) & (g3278) & (!g3361)) + ((ax8x) & (ax9x) & (!g3187) & (!g3272) & (g3278) & (g3361)) + ((ax8x) & (ax9x) & (!g3187) & (g3272) & (!g3278) & (g3361)) + ((ax8x) & (ax9x) & (!g3187) & (g3272) & (g3278) & (g3361)) + ((ax8x) & (ax9x) & (g3187) & (!g3272) & (!g3278) & (g3361)) + ((ax8x) & (ax9x) & (g3187) & (!g3272) & (g3278) & (!g3361)) + ((ax8x) & (ax9x) & (g3187) & (!g3272) & (g3278) & (g3361)) + ((ax8x) & (ax9x) & (g3187) & (g3272) & (!g3278) & (g3361)) + ((ax8x) & (ax9x) & (g3187) & (g3272) & (g3278) & (g3361)));
	assign g3363 = (((!ax8x) & (!g3187) & (!g3243) & (!g3272) & (g3278)) + ((!ax8x) & (!g3187) & (g3243) & (!g3272) & (!g3278)) + ((!ax8x) & (!g3187) & (g3243) & (!g3272) & (g3278)) + ((!ax8x) & (!g3187) & (g3243) & (g3272) & (!g3278)) + ((!ax8x) & (!g3187) & (g3243) & (g3272) & (g3278)) + ((!ax8x) & (g3187) & (g3243) & (!g3272) & (!g3278)) + ((!ax8x) & (g3187) & (g3243) & (g3272) & (!g3278)) + ((!ax8x) & (g3187) & (g3243) & (g3272) & (g3278)) + ((ax8x) & (!g3187) & (!g3243) & (!g3272) & (!g3278)) + ((ax8x) & (!g3187) & (!g3243) & (g3272) & (!g3278)) + ((ax8x) & (!g3187) & (!g3243) & (g3272) & (g3278)) + ((ax8x) & (g3187) & (!g3243) & (!g3272) & (!g3278)) + ((ax8x) & (g3187) & (!g3243) & (!g3272) & (g3278)) + ((ax8x) & (g3187) & (!g3243) & (g3272) & (!g3278)) + ((ax8x) & (g3187) & (!g3243) & (g3272) & (g3278)) + ((ax8x) & (g3187) & (g3243) & (!g3272) & (g3278)));
	assign g3364 = (((!ax4x) & (!ax5x)));
	assign g3365 = (((!g3187) & (!ax6x) & (!ax7x) & (!g3272) & (!g3278) & (!g3364)) + ((!g3187) & (!ax6x) & (!ax7x) & (g3272) & (!g3278) & (!g3364)) + ((!g3187) & (!ax6x) & (!ax7x) & (g3272) & (g3278) & (!g3364)) + ((!g3187) & (!ax6x) & (ax7x) & (!g3272) & (g3278) & (!g3364)) + ((!g3187) & (ax6x) & (ax7x) & (!g3272) & (g3278) & (!g3364)) + ((!g3187) & (ax6x) & (ax7x) & (!g3272) & (g3278) & (g3364)) + ((g3187) & (!ax6x) & (!ax7x) & (!g3272) & (!g3278) & (!g3364)) + ((g3187) & (!ax6x) & (!ax7x) & (!g3272) & (!g3278) & (g3364)) + ((g3187) & (!ax6x) & (!ax7x) & (!g3272) & (g3278) & (!g3364)) + ((g3187) & (!ax6x) & (!ax7x) & (g3272) & (!g3278) & (!g3364)) + ((g3187) & (!ax6x) & (!ax7x) & (g3272) & (!g3278) & (g3364)) + ((g3187) & (!ax6x) & (!ax7x) & (g3272) & (g3278) & (!g3364)) + ((g3187) & (!ax6x) & (!ax7x) & (g3272) & (g3278) & (g3364)) + ((g3187) & (!ax6x) & (ax7x) & (!g3272) & (!g3278) & (!g3364)) + ((g3187) & (!ax6x) & (ax7x) & (!g3272) & (g3278) & (!g3364)) + ((g3187) & (!ax6x) & (ax7x) & (!g3272) & (g3278) & (g3364)) + ((g3187) & (!ax6x) & (ax7x) & (g3272) & (!g3278) & (!g3364)) + ((g3187) & (!ax6x) & (ax7x) & (g3272) & (g3278) & (!g3364)) + ((g3187) & (ax6x) & (!ax7x) & (!g3272) & (g3278) & (!g3364)) + ((g3187) & (ax6x) & (!ax7x) & (!g3272) & (g3278) & (g3364)) + ((g3187) & (ax6x) & (ax7x) & (!g3272) & (!g3278) & (!g3364)) + ((g3187) & (ax6x) & (ax7x) & (!g3272) & (!g3278) & (g3364)) + ((g3187) & (ax6x) & (ax7x) & (!g3272) & (g3278) & (!g3364)) + ((g3187) & (ax6x) & (ax7x) & (!g3272) & (g3278) & (g3364)) + ((g3187) & (ax6x) & (ax7x) & (g3272) & (!g3278) & (!g3364)) + ((g3187) & (ax6x) & (ax7x) & (g3272) & (!g3278) & (g3364)) + ((g3187) & (ax6x) & (ax7x) & (g3272) & (g3278) & (!g3364)) + ((g3187) & (ax6x) & (ax7x) & (g3272) & (g3278) & (g3364)));
	assign g3366 = (((!g2980) & (!g3178) & (g3362) & (g3363) & (g3365)) + ((!g2980) & (g3178) & (g3362) & (!g3363) & (g3365)) + ((!g2980) & (g3178) & (g3362) & (g3363) & (!g3365)) + ((!g2980) & (g3178) & (g3362) & (g3363) & (g3365)) + ((g2980) & (!g3178) & (!g3362) & (g3363) & (g3365)) + ((g2980) & (!g3178) & (g3362) & (!g3363) & (!g3365)) + ((g2980) & (!g3178) & (g3362) & (!g3363) & (g3365)) + ((g2980) & (!g3178) & (g3362) & (g3363) & (!g3365)) + ((g2980) & (!g3178) & (g3362) & (g3363) & (g3365)) + ((g2980) & (g3178) & (!g3362) & (!g3363) & (g3365)) + ((g2980) & (g3178) & (!g3362) & (g3363) & (!g3365)) + ((g2980) & (g3178) & (!g3362) & (g3363) & (g3365)) + ((g2980) & (g3178) & (g3362) & (!g3363) & (!g3365)) + ((g2980) & (g3178) & (g3362) & (!g3363) & (g3365)) + ((g2980) & (g3178) & (g3362) & (g3363) & (!g3365)) + ((g2980) & (g3178) & (g3362) & (g3363) & (g3365)));
	assign g3367 = (((!g2779) & (!g3030) & (g3359) & (g3360) & (g3366)) + ((!g2779) & (g3030) & (g3359) & (!g3360) & (g3366)) + ((!g2779) & (g3030) & (g3359) & (g3360) & (!g3366)) + ((!g2779) & (g3030) & (g3359) & (g3360) & (g3366)) + ((g2779) & (!g3030) & (!g3359) & (g3360) & (g3366)) + ((g2779) & (!g3030) & (g3359) & (!g3360) & (!g3366)) + ((g2779) & (!g3030) & (g3359) & (!g3360) & (g3366)) + ((g2779) & (!g3030) & (g3359) & (g3360) & (!g3366)) + ((g2779) & (!g3030) & (g3359) & (g3360) & (g3366)) + ((g2779) & (g3030) & (!g3359) & (!g3360) & (g3366)) + ((g2779) & (g3030) & (!g3359) & (g3360) & (!g3366)) + ((g2779) & (g3030) & (!g3359) & (g3360) & (g3366)) + ((g2779) & (g3030) & (g3359) & (!g3360) & (!g3366)) + ((g2779) & (g3030) & (g3359) & (!g3360) & (g3366)) + ((g2779) & (g3030) & (g3359) & (g3360) & (!g3366)) + ((g2779) & (g3030) & (g3359) & (g3360) & (g3366)));
	assign g3368 = (((!g2585) & (!g2825) & (g3356) & (g3357) & (g3367)) + ((!g2585) & (g2825) & (g3356) & (!g3357) & (g3367)) + ((!g2585) & (g2825) & (g3356) & (g3357) & (!g3367)) + ((!g2585) & (g2825) & (g3356) & (g3357) & (g3367)) + ((g2585) & (!g2825) & (!g3356) & (g3357) & (g3367)) + ((g2585) & (!g2825) & (g3356) & (!g3357) & (!g3367)) + ((g2585) & (!g2825) & (g3356) & (!g3357) & (g3367)) + ((g2585) & (!g2825) & (g3356) & (g3357) & (!g3367)) + ((g2585) & (!g2825) & (g3356) & (g3357) & (g3367)) + ((g2585) & (g2825) & (!g3356) & (!g3357) & (g3367)) + ((g2585) & (g2825) & (!g3356) & (g3357) & (!g3367)) + ((g2585) & (g2825) & (!g3356) & (g3357) & (g3367)) + ((g2585) & (g2825) & (g3356) & (!g3357) & (!g3367)) + ((g2585) & (g2825) & (g3356) & (!g3357) & (g3367)) + ((g2585) & (g2825) & (g3356) & (g3357) & (!g3367)) + ((g2585) & (g2825) & (g3356) & (g3357) & (g3367)));
	assign g3369 = (((!g2398) & (!g2627) & (g3353) & (g3354) & (g3368)) + ((!g2398) & (g2627) & (g3353) & (!g3354) & (g3368)) + ((!g2398) & (g2627) & (g3353) & (g3354) & (!g3368)) + ((!g2398) & (g2627) & (g3353) & (g3354) & (g3368)) + ((g2398) & (!g2627) & (!g3353) & (g3354) & (g3368)) + ((g2398) & (!g2627) & (g3353) & (!g3354) & (!g3368)) + ((g2398) & (!g2627) & (g3353) & (!g3354) & (g3368)) + ((g2398) & (!g2627) & (g3353) & (g3354) & (!g3368)) + ((g2398) & (!g2627) & (g3353) & (g3354) & (g3368)) + ((g2398) & (g2627) & (!g3353) & (!g3354) & (g3368)) + ((g2398) & (g2627) & (!g3353) & (g3354) & (!g3368)) + ((g2398) & (g2627) & (!g3353) & (g3354) & (g3368)) + ((g2398) & (g2627) & (g3353) & (!g3354) & (!g3368)) + ((g2398) & (g2627) & (g3353) & (!g3354) & (g3368)) + ((g2398) & (g2627) & (g3353) & (g3354) & (!g3368)) + ((g2398) & (g2627) & (g3353) & (g3354) & (g3368)));
	assign g3370 = (((!g2218) & (!g2436) & (g3350) & (g3351) & (g3369)) + ((!g2218) & (g2436) & (g3350) & (!g3351) & (g3369)) + ((!g2218) & (g2436) & (g3350) & (g3351) & (!g3369)) + ((!g2218) & (g2436) & (g3350) & (g3351) & (g3369)) + ((g2218) & (!g2436) & (!g3350) & (g3351) & (g3369)) + ((g2218) & (!g2436) & (g3350) & (!g3351) & (!g3369)) + ((g2218) & (!g2436) & (g3350) & (!g3351) & (g3369)) + ((g2218) & (!g2436) & (g3350) & (g3351) & (!g3369)) + ((g2218) & (!g2436) & (g3350) & (g3351) & (g3369)) + ((g2218) & (g2436) & (!g3350) & (!g3351) & (g3369)) + ((g2218) & (g2436) & (!g3350) & (g3351) & (!g3369)) + ((g2218) & (g2436) & (!g3350) & (g3351) & (g3369)) + ((g2218) & (g2436) & (g3350) & (!g3351) & (!g3369)) + ((g2218) & (g2436) & (g3350) & (!g3351) & (g3369)) + ((g2218) & (g2436) & (g3350) & (g3351) & (!g3369)) + ((g2218) & (g2436) & (g3350) & (g3351) & (g3369)));
	assign g3371 = (((!g2045) & (!g2252) & (g3347) & (g3348) & (g3370)) + ((!g2045) & (g2252) & (g3347) & (!g3348) & (g3370)) + ((!g2045) & (g2252) & (g3347) & (g3348) & (!g3370)) + ((!g2045) & (g2252) & (g3347) & (g3348) & (g3370)) + ((g2045) & (!g2252) & (!g3347) & (g3348) & (g3370)) + ((g2045) & (!g2252) & (g3347) & (!g3348) & (!g3370)) + ((g2045) & (!g2252) & (g3347) & (!g3348) & (g3370)) + ((g2045) & (!g2252) & (g3347) & (g3348) & (!g3370)) + ((g2045) & (!g2252) & (g3347) & (g3348) & (g3370)) + ((g2045) & (g2252) & (!g3347) & (!g3348) & (g3370)) + ((g2045) & (g2252) & (!g3347) & (g3348) & (!g3370)) + ((g2045) & (g2252) & (!g3347) & (g3348) & (g3370)) + ((g2045) & (g2252) & (g3347) & (!g3348) & (!g3370)) + ((g2045) & (g2252) & (g3347) & (!g3348) & (g3370)) + ((g2045) & (g2252) & (g3347) & (g3348) & (!g3370)) + ((g2045) & (g2252) & (g3347) & (g3348) & (g3370)));
	assign g3372 = (((!g1879) & (!g2075) & (g3344) & (g3345) & (g3371)) + ((!g1879) & (g2075) & (g3344) & (!g3345) & (g3371)) + ((!g1879) & (g2075) & (g3344) & (g3345) & (!g3371)) + ((!g1879) & (g2075) & (g3344) & (g3345) & (g3371)) + ((g1879) & (!g2075) & (!g3344) & (g3345) & (g3371)) + ((g1879) & (!g2075) & (g3344) & (!g3345) & (!g3371)) + ((g1879) & (!g2075) & (g3344) & (!g3345) & (g3371)) + ((g1879) & (!g2075) & (g3344) & (g3345) & (!g3371)) + ((g1879) & (!g2075) & (g3344) & (g3345) & (g3371)) + ((g1879) & (g2075) & (!g3344) & (!g3345) & (g3371)) + ((g1879) & (g2075) & (!g3344) & (g3345) & (!g3371)) + ((g1879) & (g2075) & (!g3344) & (g3345) & (g3371)) + ((g1879) & (g2075) & (g3344) & (!g3345) & (!g3371)) + ((g1879) & (g2075) & (g3344) & (!g3345) & (g3371)) + ((g1879) & (g2075) & (g3344) & (g3345) & (!g3371)) + ((g1879) & (g2075) & (g3344) & (g3345) & (g3371)));
	assign g3373 = (((!g1720) & (!g1905) & (g3341) & (g3342) & (g3372)) + ((!g1720) & (g1905) & (g3341) & (!g3342) & (g3372)) + ((!g1720) & (g1905) & (g3341) & (g3342) & (!g3372)) + ((!g1720) & (g1905) & (g3341) & (g3342) & (g3372)) + ((g1720) & (!g1905) & (!g3341) & (g3342) & (g3372)) + ((g1720) & (!g1905) & (g3341) & (!g3342) & (!g3372)) + ((g1720) & (!g1905) & (g3341) & (!g3342) & (g3372)) + ((g1720) & (!g1905) & (g3341) & (g3342) & (!g3372)) + ((g1720) & (!g1905) & (g3341) & (g3342) & (g3372)) + ((g1720) & (g1905) & (!g3341) & (!g3342) & (g3372)) + ((g1720) & (g1905) & (!g3341) & (g3342) & (!g3372)) + ((g1720) & (g1905) & (!g3341) & (g3342) & (g3372)) + ((g1720) & (g1905) & (g3341) & (!g3342) & (!g3372)) + ((g1720) & (g1905) & (g3341) & (!g3342) & (g3372)) + ((g1720) & (g1905) & (g3341) & (g3342) & (!g3372)) + ((g1720) & (g1905) & (g3341) & (g3342) & (g3372)));
	assign g3374 = (((!g1568) & (!g1742) & (g3338) & (g3339) & (g3373)) + ((!g1568) & (g1742) & (g3338) & (!g3339) & (g3373)) + ((!g1568) & (g1742) & (g3338) & (g3339) & (!g3373)) + ((!g1568) & (g1742) & (g3338) & (g3339) & (g3373)) + ((g1568) & (!g1742) & (!g3338) & (g3339) & (g3373)) + ((g1568) & (!g1742) & (g3338) & (!g3339) & (!g3373)) + ((g1568) & (!g1742) & (g3338) & (!g3339) & (g3373)) + ((g1568) & (!g1742) & (g3338) & (g3339) & (!g3373)) + ((g1568) & (!g1742) & (g3338) & (g3339) & (g3373)) + ((g1568) & (g1742) & (!g3338) & (!g3339) & (g3373)) + ((g1568) & (g1742) & (!g3338) & (g3339) & (!g3373)) + ((g1568) & (g1742) & (!g3338) & (g3339) & (g3373)) + ((g1568) & (g1742) & (g3338) & (!g3339) & (!g3373)) + ((g1568) & (g1742) & (g3338) & (!g3339) & (g3373)) + ((g1568) & (g1742) & (g3338) & (g3339) & (!g3373)) + ((g1568) & (g1742) & (g3338) & (g3339) & (g3373)));
	assign g3375 = (((!g1423) & (!g1586) & (g3335) & (g3336) & (g3374)) + ((!g1423) & (g1586) & (g3335) & (!g3336) & (g3374)) + ((!g1423) & (g1586) & (g3335) & (g3336) & (!g3374)) + ((!g1423) & (g1586) & (g3335) & (g3336) & (g3374)) + ((g1423) & (!g1586) & (!g3335) & (g3336) & (g3374)) + ((g1423) & (!g1586) & (g3335) & (!g3336) & (!g3374)) + ((g1423) & (!g1586) & (g3335) & (!g3336) & (g3374)) + ((g1423) & (!g1586) & (g3335) & (g3336) & (!g3374)) + ((g1423) & (!g1586) & (g3335) & (g3336) & (g3374)) + ((g1423) & (g1586) & (!g3335) & (!g3336) & (g3374)) + ((g1423) & (g1586) & (!g3335) & (g3336) & (!g3374)) + ((g1423) & (g1586) & (!g3335) & (g3336) & (g3374)) + ((g1423) & (g1586) & (g3335) & (!g3336) & (!g3374)) + ((g1423) & (g1586) & (g3335) & (!g3336) & (g3374)) + ((g1423) & (g1586) & (g3335) & (g3336) & (!g3374)) + ((g1423) & (g1586) & (g3335) & (g3336) & (g3374)));
	assign g3376 = (((!g1285) & (!g1437) & (g3332) & (g3333) & (g3375)) + ((!g1285) & (g1437) & (g3332) & (!g3333) & (g3375)) + ((!g1285) & (g1437) & (g3332) & (g3333) & (!g3375)) + ((!g1285) & (g1437) & (g3332) & (g3333) & (g3375)) + ((g1285) & (!g1437) & (!g3332) & (g3333) & (g3375)) + ((g1285) & (!g1437) & (g3332) & (!g3333) & (!g3375)) + ((g1285) & (!g1437) & (g3332) & (!g3333) & (g3375)) + ((g1285) & (!g1437) & (g3332) & (g3333) & (!g3375)) + ((g1285) & (!g1437) & (g3332) & (g3333) & (g3375)) + ((g1285) & (g1437) & (!g3332) & (!g3333) & (g3375)) + ((g1285) & (g1437) & (!g3332) & (g3333) & (!g3375)) + ((g1285) & (g1437) & (!g3332) & (g3333) & (g3375)) + ((g1285) & (g1437) & (g3332) & (!g3333) & (!g3375)) + ((g1285) & (g1437) & (g3332) & (!g3333) & (g3375)) + ((g1285) & (g1437) & (g3332) & (g3333) & (!g3375)) + ((g1285) & (g1437) & (g3332) & (g3333) & (g3375)));
	assign g3377 = (((!g1154) & (!g1295) & (g3329) & (g3330) & (g3376)) + ((!g1154) & (g1295) & (g3329) & (!g3330) & (g3376)) + ((!g1154) & (g1295) & (g3329) & (g3330) & (!g3376)) + ((!g1154) & (g1295) & (g3329) & (g3330) & (g3376)) + ((g1154) & (!g1295) & (!g3329) & (g3330) & (g3376)) + ((g1154) & (!g1295) & (g3329) & (!g3330) & (!g3376)) + ((g1154) & (!g1295) & (g3329) & (!g3330) & (g3376)) + ((g1154) & (!g1295) & (g3329) & (g3330) & (!g3376)) + ((g1154) & (!g1295) & (g3329) & (g3330) & (g3376)) + ((g1154) & (g1295) & (!g3329) & (!g3330) & (g3376)) + ((g1154) & (g1295) & (!g3329) & (g3330) & (!g3376)) + ((g1154) & (g1295) & (!g3329) & (g3330) & (g3376)) + ((g1154) & (g1295) & (g3329) & (!g3330) & (!g3376)) + ((g1154) & (g1295) & (g3329) & (!g3330) & (g3376)) + ((g1154) & (g1295) & (g3329) & (g3330) & (!g3376)) + ((g1154) & (g1295) & (g3329) & (g3330) & (g3376)));
	assign g3378 = (((!g1030) & (!g1160) & (g3326) & (g3327) & (g3377)) + ((!g1030) & (g1160) & (g3326) & (!g3327) & (g3377)) + ((!g1030) & (g1160) & (g3326) & (g3327) & (!g3377)) + ((!g1030) & (g1160) & (g3326) & (g3327) & (g3377)) + ((g1030) & (!g1160) & (!g3326) & (g3327) & (g3377)) + ((g1030) & (!g1160) & (g3326) & (!g3327) & (!g3377)) + ((g1030) & (!g1160) & (g3326) & (!g3327) & (g3377)) + ((g1030) & (!g1160) & (g3326) & (g3327) & (!g3377)) + ((g1030) & (!g1160) & (g3326) & (g3327) & (g3377)) + ((g1030) & (g1160) & (!g3326) & (!g3327) & (g3377)) + ((g1030) & (g1160) & (!g3326) & (g3327) & (!g3377)) + ((g1030) & (g1160) & (!g3326) & (g3327) & (g3377)) + ((g1030) & (g1160) & (g3326) & (!g3327) & (!g3377)) + ((g1030) & (g1160) & (g3326) & (!g3327) & (g3377)) + ((g1030) & (g1160) & (g3326) & (g3327) & (!g3377)) + ((g1030) & (g1160) & (g3326) & (g3327) & (g3377)));
	assign g3379 = (((!g914) & (!g1032) & (g3323) & (g3324) & (g3378)) + ((!g914) & (g1032) & (g3323) & (!g3324) & (g3378)) + ((!g914) & (g1032) & (g3323) & (g3324) & (!g3378)) + ((!g914) & (g1032) & (g3323) & (g3324) & (g3378)) + ((g914) & (!g1032) & (!g3323) & (g3324) & (g3378)) + ((g914) & (!g1032) & (g3323) & (!g3324) & (!g3378)) + ((g914) & (!g1032) & (g3323) & (!g3324) & (g3378)) + ((g914) & (!g1032) & (g3323) & (g3324) & (!g3378)) + ((g914) & (!g1032) & (g3323) & (g3324) & (g3378)) + ((g914) & (g1032) & (!g3323) & (!g3324) & (g3378)) + ((g914) & (g1032) & (!g3323) & (g3324) & (!g3378)) + ((g914) & (g1032) & (!g3323) & (g3324) & (g3378)) + ((g914) & (g1032) & (g3323) & (!g3324) & (!g3378)) + ((g914) & (g1032) & (g3323) & (!g3324) & (g3378)) + ((g914) & (g1032) & (g3323) & (g3324) & (!g3378)) + ((g914) & (g1032) & (g3323) & (g3324) & (g3378)));
	assign g3380 = (((!g803) & (!g851) & (g3320) & (g3321) & (g3379)) + ((!g803) & (g851) & (g3320) & (!g3321) & (g3379)) + ((!g803) & (g851) & (g3320) & (g3321) & (!g3379)) + ((!g803) & (g851) & (g3320) & (g3321) & (g3379)) + ((g803) & (!g851) & (!g3320) & (g3321) & (g3379)) + ((g803) & (!g851) & (g3320) & (!g3321) & (!g3379)) + ((g803) & (!g851) & (g3320) & (!g3321) & (g3379)) + ((g803) & (!g851) & (g3320) & (g3321) & (!g3379)) + ((g803) & (!g851) & (g3320) & (g3321) & (g3379)) + ((g803) & (g851) & (!g3320) & (!g3321) & (g3379)) + ((g803) & (g851) & (!g3320) & (g3321) & (!g3379)) + ((g803) & (g851) & (!g3320) & (g3321) & (g3379)) + ((g803) & (g851) & (g3320) & (!g3321) & (!g3379)) + ((g803) & (g851) & (g3320) & (!g3321) & (g3379)) + ((g803) & (g851) & (g3320) & (g3321) & (!g3379)) + ((g803) & (g851) & (g3320) & (g3321) & (g3379)));
	assign g3381 = (((!g700) & (!g744) & (g3317) & (g3318) & (g3380)) + ((!g700) & (g744) & (g3317) & (!g3318) & (g3380)) + ((!g700) & (g744) & (g3317) & (g3318) & (!g3380)) + ((!g700) & (g744) & (g3317) & (g3318) & (g3380)) + ((g700) & (!g744) & (!g3317) & (g3318) & (g3380)) + ((g700) & (!g744) & (g3317) & (!g3318) & (!g3380)) + ((g700) & (!g744) & (g3317) & (!g3318) & (g3380)) + ((g700) & (!g744) & (g3317) & (g3318) & (!g3380)) + ((g700) & (!g744) & (g3317) & (g3318) & (g3380)) + ((g700) & (g744) & (!g3317) & (!g3318) & (g3380)) + ((g700) & (g744) & (!g3317) & (g3318) & (!g3380)) + ((g700) & (g744) & (!g3317) & (g3318) & (g3380)) + ((g700) & (g744) & (g3317) & (!g3318) & (!g3380)) + ((g700) & (g744) & (g3317) & (!g3318) & (g3380)) + ((g700) & (g744) & (g3317) & (g3318) & (!g3380)) + ((g700) & (g744) & (g3317) & (g3318) & (g3380)));
	assign g3382 = (((!g604) & (!g645) & (g3314) & (g3315) & (g3381)) + ((!g604) & (g645) & (g3314) & (!g3315) & (g3381)) + ((!g604) & (g645) & (g3314) & (g3315) & (!g3381)) + ((!g604) & (g645) & (g3314) & (g3315) & (g3381)) + ((g604) & (!g645) & (!g3314) & (g3315) & (g3381)) + ((g604) & (!g645) & (g3314) & (!g3315) & (!g3381)) + ((g604) & (!g645) & (g3314) & (!g3315) & (g3381)) + ((g604) & (!g645) & (g3314) & (g3315) & (!g3381)) + ((g604) & (!g645) & (g3314) & (g3315) & (g3381)) + ((g604) & (g645) & (!g3314) & (!g3315) & (g3381)) + ((g604) & (g645) & (!g3314) & (g3315) & (!g3381)) + ((g604) & (g645) & (!g3314) & (g3315) & (g3381)) + ((g604) & (g645) & (g3314) & (!g3315) & (!g3381)) + ((g604) & (g645) & (g3314) & (!g3315) & (g3381)) + ((g604) & (g645) & (g3314) & (g3315) & (!g3381)) + ((g604) & (g645) & (g3314) & (g3315) & (g3381)));
	assign g3383 = (((!g515) & (!g553) & (g3311) & (g3312) & (g3382)) + ((!g515) & (g553) & (g3311) & (!g3312) & (g3382)) + ((!g515) & (g553) & (g3311) & (g3312) & (!g3382)) + ((!g515) & (g553) & (g3311) & (g3312) & (g3382)) + ((g515) & (!g553) & (!g3311) & (g3312) & (g3382)) + ((g515) & (!g553) & (g3311) & (!g3312) & (!g3382)) + ((g515) & (!g553) & (g3311) & (!g3312) & (g3382)) + ((g515) & (!g553) & (g3311) & (g3312) & (!g3382)) + ((g515) & (!g553) & (g3311) & (g3312) & (g3382)) + ((g515) & (g553) & (!g3311) & (!g3312) & (g3382)) + ((g515) & (g553) & (!g3311) & (g3312) & (!g3382)) + ((g515) & (g553) & (!g3311) & (g3312) & (g3382)) + ((g515) & (g553) & (g3311) & (!g3312) & (!g3382)) + ((g515) & (g553) & (g3311) & (!g3312) & (g3382)) + ((g515) & (g553) & (g3311) & (g3312) & (!g3382)) + ((g515) & (g553) & (g3311) & (g3312) & (g3382)));
	assign g3384 = (((!g433) & (!g468) & (g3308) & (g3309) & (g3383)) + ((!g433) & (g468) & (g3308) & (!g3309) & (g3383)) + ((!g433) & (g468) & (g3308) & (g3309) & (!g3383)) + ((!g433) & (g468) & (g3308) & (g3309) & (g3383)) + ((g433) & (!g468) & (!g3308) & (g3309) & (g3383)) + ((g433) & (!g468) & (g3308) & (!g3309) & (!g3383)) + ((g433) & (!g468) & (g3308) & (!g3309) & (g3383)) + ((g433) & (!g468) & (g3308) & (g3309) & (!g3383)) + ((g433) & (!g468) & (g3308) & (g3309) & (g3383)) + ((g433) & (g468) & (!g3308) & (!g3309) & (g3383)) + ((g433) & (g468) & (!g3308) & (g3309) & (!g3383)) + ((g433) & (g468) & (!g3308) & (g3309) & (g3383)) + ((g433) & (g468) & (g3308) & (!g3309) & (!g3383)) + ((g433) & (g468) & (g3308) & (!g3309) & (g3383)) + ((g433) & (g468) & (g3308) & (g3309) & (!g3383)) + ((g433) & (g468) & (g3308) & (g3309) & (g3383)));
	assign g3385 = (((!g358) & (!g390) & (g3305) & (g3306) & (g3384)) + ((!g358) & (g390) & (g3305) & (!g3306) & (g3384)) + ((!g358) & (g390) & (g3305) & (g3306) & (!g3384)) + ((!g358) & (g390) & (g3305) & (g3306) & (g3384)) + ((g358) & (!g390) & (!g3305) & (g3306) & (g3384)) + ((g358) & (!g390) & (g3305) & (!g3306) & (!g3384)) + ((g358) & (!g390) & (g3305) & (!g3306) & (g3384)) + ((g358) & (!g390) & (g3305) & (g3306) & (!g3384)) + ((g358) & (!g390) & (g3305) & (g3306) & (g3384)) + ((g358) & (g390) & (!g3305) & (!g3306) & (g3384)) + ((g358) & (g390) & (!g3305) & (g3306) & (!g3384)) + ((g358) & (g390) & (!g3305) & (g3306) & (g3384)) + ((g358) & (g390) & (g3305) & (!g3306) & (!g3384)) + ((g358) & (g390) & (g3305) & (!g3306) & (g3384)) + ((g358) & (g390) & (g3305) & (g3306) & (!g3384)) + ((g358) & (g390) & (g3305) & (g3306) & (g3384)));
	assign g3386 = (((!g290) & (!g319) & (g3302) & (g3303) & (g3385)) + ((!g290) & (g319) & (g3302) & (!g3303) & (g3385)) + ((!g290) & (g319) & (g3302) & (g3303) & (!g3385)) + ((!g290) & (g319) & (g3302) & (g3303) & (g3385)) + ((g290) & (!g319) & (!g3302) & (g3303) & (g3385)) + ((g290) & (!g319) & (g3302) & (!g3303) & (!g3385)) + ((g290) & (!g319) & (g3302) & (!g3303) & (g3385)) + ((g290) & (!g319) & (g3302) & (g3303) & (!g3385)) + ((g290) & (!g319) & (g3302) & (g3303) & (g3385)) + ((g290) & (g319) & (!g3302) & (!g3303) & (g3385)) + ((g290) & (g319) & (!g3302) & (g3303) & (!g3385)) + ((g290) & (g319) & (!g3302) & (g3303) & (g3385)) + ((g290) & (g319) & (g3302) & (!g3303) & (!g3385)) + ((g290) & (g319) & (g3302) & (!g3303) & (g3385)) + ((g290) & (g319) & (g3302) & (g3303) & (!g3385)) + ((g290) & (g319) & (g3302) & (g3303) & (g3385)));
	assign g3387 = (((!g229) & (!g255) & (g3299) & (g3300) & (g3386)) + ((!g229) & (g255) & (g3299) & (!g3300) & (g3386)) + ((!g229) & (g255) & (g3299) & (g3300) & (!g3386)) + ((!g229) & (g255) & (g3299) & (g3300) & (g3386)) + ((g229) & (!g255) & (!g3299) & (g3300) & (g3386)) + ((g229) & (!g255) & (g3299) & (!g3300) & (!g3386)) + ((g229) & (!g255) & (g3299) & (!g3300) & (g3386)) + ((g229) & (!g255) & (g3299) & (g3300) & (!g3386)) + ((g229) & (!g255) & (g3299) & (g3300) & (g3386)) + ((g229) & (g255) & (!g3299) & (!g3300) & (g3386)) + ((g229) & (g255) & (!g3299) & (g3300) & (!g3386)) + ((g229) & (g255) & (!g3299) & (g3300) & (g3386)) + ((g229) & (g255) & (g3299) & (!g3300) & (!g3386)) + ((g229) & (g255) & (g3299) & (!g3300) & (g3386)) + ((g229) & (g255) & (g3299) & (g3300) & (!g3386)) + ((g229) & (g255) & (g3299) & (g3300) & (g3386)));
	assign g3388 = (((!g174) & (!g198) & (g3296) & (g3297) & (g3387)) + ((!g174) & (g198) & (g3296) & (!g3297) & (g3387)) + ((!g174) & (g198) & (g3296) & (g3297) & (!g3387)) + ((!g174) & (g198) & (g3296) & (g3297) & (g3387)) + ((g174) & (!g198) & (!g3296) & (g3297) & (g3387)) + ((g174) & (!g198) & (g3296) & (!g3297) & (!g3387)) + ((g174) & (!g198) & (g3296) & (!g3297) & (g3387)) + ((g174) & (!g198) & (g3296) & (g3297) & (!g3387)) + ((g174) & (!g198) & (g3296) & (g3297) & (g3387)) + ((g174) & (g198) & (!g3296) & (!g3297) & (g3387)) + ((g174) & (g198) & (!g3296) & (g3297) & (!g3387)) + ((g174) & (g198) & (!g3296) & (g3297) & (g3387)) + ((g174) & (g198) & (g3296) & (!g3297) & (!g3387)) + ((g174) & (g198) & (g3296) & (!g3297) & (g3387)) + ((g174) & (g198) & (g3296) & (g3297) & (!g3387)) + ((g174) & (g198) & (g3296) & (g3297) & (g3387)));
	assign g3389 = (((!g127) & (!g147) & (g3293) & (g3294) & (g3388)) + ((!g127) & (g147) & (g3293) & (!g3294) & (g3388)) + ((!g127) & (g147) & (g3293) & (g3294) & (!g3388)) + ((!g127) & (g147) & (g3293) & (g3294) & (g3388)) + ((g127) & (!g147) & (!g3293) & (g3294) & (g3388)) + ((g127) & (!g147) & (g3293) & (!g3294) & (!g3388)) + ((g127) & (!g147) & (g3293) & (!g3294) & (g3388)) + ((g127) & (!g147) & (g3293) & (g3294) & (!g3388)) + ((g127) & (!g147) & (g3293) & (g3294) & (g3388)) + ((g127) & (g147) & (!g3293) & (!g3294) & (g3388)) + ((g127) & (g147) & (!g3293) & (g3294) & (!g3388)) + ((g127) & (g147) & (!g3293) & (g3294) & (g3388)) + ((g127) & (g147) & (g3293) & (!g3294) & (!g3388)) + ((g127) & (g147) & (g3293) & (!g3294) & (g3388)) + ((g127) & (g147) & (g3293) & (g3294) & (!g3388)) + ((g127) & (g147) & (g3293) & (g3294) & (g3388)));
	assign g3390 = (((!g87) & (!g104) & (g3290) & (g3291) & (g3389)) + ((!g87) & (g104) & (g3290) & (!g3291) & (g3389)) + ((!g87) & (g104) & (g3290) & (g3291) & (!g3389)) + ((!g87) & (g104) & (g3290) & (g3291) & (g3389)) + ((g87) & (!g104) & (!g3290) & (g3291) & (g3389)) + ((g87) & (!g104) & (g3290) & (!g3291) & (!g3389)) + ((g87) & (!g104) & (g3290) & (!g3291) & (g3389)) + ((g87) & (!g104) & (g3290) & (g3291) & (!g3389)) + ((g87) & (!g104) & (g3290) & (g3291) & (g3389)) + ((g87) & (g104) & (!g3290) & (!g3291) & (g3389)) + ((g87) & (g104) & (!g3290) & (g3291) & (!g3389)) + ((g87) & (g104) & (!g3290) & (g3291) & (g3389)) + ((g87) & (g104) & (g3290) & (!g3291) & (!g3389)) + ((g87) & (g104) & (g3290) & (!g3291) & (g3389)) + ((g87) & (g104) & (g3290) & (g3291) & (!g3389)) + ((g87) & (g104) & (g3290) & (g3291) & (g3389)));
	assign g3391 = (((!g54) & (!g68) & (g3287) & (g3288) & (g3390)) + ((!g54) & (g68) & (g3287) & (!g3288) & (g3390)) + ((!g54) & (g68) & (g3287) & (g3288) & (!g3390)) + ((!g54) & (g68) & (g3287) & (g3288) & (g3390)) + ((g54) & (!g68) & (!g3287) & (g3288) & (g3390)) + ((g54) & (!g68) & (g3287) & (!g3288) & (!g3390)) + ((g54) & (!g68) & (g3287) & (!g3288) & (g3390)) + ((g54) & (!g68) & (g3287) & (g3288) & (!g3390)) + ((g54) & (!g68) & (g3287) & (g3288) & (g3390)) + ((g54) & (g68) & (!g3287) & (!g3288) & (g3390)) + ((g54) & (g68) & (!g3287) & (g3288) & (!g3390)) + ((g54) & (g68) & (!g3287) & (g3288) & (g3390)) + ((g54) & (g68) & (g3287) & (!g3288) & (!g3390)) + ((g54) & (g68) & (g3287) & (!g3288) & (g3390)) + ((g54) & (g68) & (g3287) & (g3288) & (!g3390)) + ((g54) & (g68) & (g3287) & (g3288) & (g3390)));
	assign g3392 = (((!g27) & (!g39) & (g3284) & (g3285) & (g3391)) + ((!g27) & (g39) & (g3284) & (!g3285) & (g3391)) + ((!g27) & (g39) & (g3284) & (g3285) & (!g3391)) + ((!g27) & (g39) & (g3284) & (g3285) & (g3391)) + ((g27) & (!g39) & (!g3284) & (g3285) & (g3391)) + ((g27) & (!g39) & (g3284) & (!g3285) & (!g3391)) + ((g27) & (!g39) & (g3284) & (!g3285) & (g3391)) + ((g27) & (!g39) & (g3284) & (g3285) & (!g3391)) + ((g27) & (!g39) & (g3284) & (g3285) & (g3391)) + ((g27) & (g39) & (!g3284) & (!g3285) & (g3391)) + ((g27) & (g39) & (!g3284) & (g3285) & (!g3391)) + ((g27) & (g39) & (!g3284) & (g3285) & (g3391)) + ((g27) & (g39) & (g3284) & (!g3285) & (!g3391)) + ((g27) & (g39) & (g3284) & (!g3285) & (g3391)) + ((g27) & (g39) & (g3284) & (g3285) & (!g3391)) + ((g27) & (g39) & (g3284) & (g3285) & (g3391)));
	assign g3393 = (((!g8) & (!g18) & (g3281) & (g3282) & (g3392)) + ((!g8) & (g18) & (g3281) & (!g3282) & (g3392)) + ((!g8) & (g18) & (g3281) & (g3282) & (!g3392)) + ((!g8) & (g18) & (g3281) & (g3282) & (g3392)) + ((g8) & (!g18) & (!g3281) & (g3282) & (g3392)) + ((g8) & (!g18) & (g3281) & (!g3282) & (!g3392)) + ((g8) & (!g18) & (g3281) & (!g3282) & (g3392)) + ((g8) & (!g18) & (g3281) & (g3282) & (!g3392)) + ((g8) & (!g18) & (g3281) & (g3282) & (g3392)) + ((g8) & (g18) & (!g3281) & (!g3282) & (g3392)) + ((g8) & (g18) & (!g3281) & (g3282) & (!g3392)) + ((g8) & (g18) & (!g3281) & (g3282) & (g3392)) + ((g8) & (g18) & (g3281) & (!g3282) & (!g3392)) + ((g8) & (g18) & (g3281) & (!g3282) & (g3392)) + ((g8) & (g18) & (g3281) & (g3282) & (!g3392)) + ((g8) & (g18) & (g3281) & (g3282) & (g3392)));
	assign g3394 = (((!g4) & (!g3275) & (g3276)) + ((!g4) & (g3275) & (!g3276)) + ((!g4) & (g3275) & (g3276)) + ((g4) & (g3275) & (g3276)));
	assign g3395 = (((!g3272) & (g3278)));
	assign g3396 = (((!g4) & (!g3275) & (!g3276) & (!g3272) & (!g3278)) + ((!g4) & (!g3275) & (!g3276) & (g3272) & (!g3278)) + ((!g4) & (!g3275) & (!g3276) & (g3272) & (g3278)) + ((!g4) & (!g3275) & (g3276) & (!g3272) & (g3278)) + ((!g4) & (g3275) & (g3276) & (!g3272) & (!g3278)) + ((!g4) & (g3275) & (g3276) & (!g3272) & (g3278)) + ((!g4) & (g3275) & (g3276) & (g3272) & (!g3278)) + ((!g4) & (g3275) & (g3276) & (g3272) & (g3278)) + ((g4) & (!g3275) & (g3276) & (!g3272) & (!g3278)) + ((g4) & (!g3275) & (g3276) & (!g3272) & (g3278)) + ((g4) & (!g3275) & (g3276) & (g3272) & (!g3278)) + ((g4) & (!g3275) & (g3276) & (g3272) & (g3278)) + ((g4) & (g3275) & (!g3276) & (!g3272) & (!g3278)) + ((g4) & (g3275) & (!g3276) & (g3272) & (!g3278)) + ((g4) & (g3275) & (!g3276) & (g3272) & (g3278)) + ((g4) & (g3275) & (g3276) & (!g3272) & (g3278)));
	assign g3397 = (((!g2) & (!g8) & (g3188) & (g3271)) + ((!g2) & (g8) & (!g3188) & (g3271)) + ((!g2) & (g8) & (g3188) & (!g3271)) + ((!g2) & (g8) & (g3188) & (g3271)) + ((g2) & (!g8) & (!g3188) & (!g3271)) + ((g2) & (!g8) & (!g3188) & (g3271)) + ((g2) & (!g8) & (g3188) & (!g3271)) + ((g2) & (g8) & (!g3188) & (!g3271)));
	assign g3398 = (((!g3274) & (!g3272) & (!g3278) & (g3397)) + ((!g3274) & (g3272) & (!g3278) & (g3397)) + ((!g3274) & (g3272) & (g3278) & (g3397)) + ((g3274) & (!g3272) & (!g3278) & (!g3397)) + ((g3274) & (!g3272) & (g3278) & (!g3397)) + ((g3274) & (!g3272) & (g3278) & (g3397)) + ((g3274) & (g3272) & (!g3278) & (!g3397)) + ((g3274) & (g3272) & (g3278) & (!g3397)));
	assign g3399 = (((!g4) & (!g2) & (!g3398) & (g3279) & (g3393)) + ((!g4) & (!g2) & (g3398) & (!g3279) & (!g3393)) + ((!g4) & (!g2) & (g3398) & (!g3279) & (g3393)) + ((!g4) & (!g2) & (g3398) & (g3279) & (!g3393)) + ((!g4) & (!g2) & (g3398) & (g3279) & (g3393)) + ((!g4) & (g2) & (!g3398) & (!g3279) & (g3393)) + ((!g4) & (g2) & (!g3398) & (g3279) & (!g3393)) + ((!g4) & (g2) & (!g3398) & (g3279) & (g3393)) + ((!g4) & (g2) & (g3398) & (!g3279) & (!g3393)) + ((!g4) & (g2) & (g3398) & (!g3279) & (g3393)) + ((!g4) & (g2) & (g3398) & (g3279) & (!g3393)) + ((!g4) & (g2) & (g3398) & (g3279) & (g3393)) + ((g4) & (!g2) & (g3398) & (g3279) & (g3393)) + ((g4) & (g2) & (g3398) & (!g3279) & (g3393)) + ((g4) & (g2) & (g3398) & (g3279) & (!g3393)) + ((g4) & (g2) & (g3398) & (g3279) & (g3393)));
	assign g3400 = (((!g1) & (!g3273) & (!g3394) & (g3395) & (!g3396) & (!g3399)) + ((!g1) & (!g3273) & (g3394) & (!g3395) & (!g3396) & (!g3399)) + ((!g1) & (!g3273) & (g3394) & (g3395) & (!g3396) & (!g3399)) + ((!g1) & (g3273) & (!g3394) & (!g3395) & (!g3396) & (!g3399)) + ((!g1) & (g3273) & (!g3394) & (g3395) & (!g3396) & (!g3399)) + ((g1) & (!g3273) & (!g3394) & (!g3395) & (!g3396) & (!g3399)) + ((g1) & (!g3273) & (!g3394) & (!g3395) & (!g3396) & (g3399)) + ((g1) & (!g3273) & (!g3394) & (!g3395) & (g3396) & (!g3399)) + ((g1) & (!g3273) & (!g3394) & (g3395) & (!g3396) & (!g3399)) + ((g1) & (!g3273) & (!g3394) & (g3395) & (!g3396) & (g3399)) + ((g1) & (!g3273) & (!g3394) & (g3395) & (g3396) & (!g3399)) + ((g1) & (!g3273) & (g3394) & (g3395) & (!g3396) & (!g3399)) + ((g1) & (!g3273) & (g3394) & (g3395) & (!g3396) & (g3399)) + ((g1) & (!g3273) & (g3394) & (g3395) & (g3396) & (!g3399)) + ((g1) & (g3273) & (g3394) & (!g3395) & (!g3396) & (!g3399)) + ((g1) & (g3273) & (g3394) & (!g3395) & (!g3396) & (g3399)) + ((g1) & (g3273) & (g3394) & (!g3395) & (g3396) & (!g3399)) + ((g1) & (g3273) & (g3394) & (g3395) & (!g3396) & (!g3399)) + ((g1) & (g3273) & (g3394) & (g3395) & (!g3396) & (g3399)) + ((g1) & (g3273) & (g3394) & (g3395) & (g3396) & (!g3399)));
	assign g3401 = (((!g2) & (!g3279) & (g3393) & (!g3400)) + ((!g2) & (g3279) & (!g3393) & (!g3400)) + ((!g2) & (g3279) & (!g3393) & (g3400)) + ((!g2) & (g3279) & (g3393) & (g3400)) + ((g2) & (!g3279) & (!g3393) & (!g3400)) + ((g2) & (g3279) & (!g3393) & (g3400)) + ((g2) & (g3279) & (g3393) & (!g3400)) + ((g2) & (g3279) & (g3393) & (g3400)));
	assign g3402 = (((!g4) & (!g2) & (!g3398) & (!g3279) & (!g3393) & (!g3400)) + ((!g4) & (!g2) & (!g3398) & (!g3279) & (g3393) & (!g3400)) + ((!g4) & (!g2) & (!g3398) & (g3279) & (!g3393) & (!g3400)) + ((!g4) & (!g2) & (g3398) & (!g3279) & (!g3393) & (g3400)) + ((!g4) & (!g2) & (g3398) & (!g3279) & (g3393) & (g3400)) + ((!g4) & (!g2) & (g3398) & (g3279) & (!g3393) & (g3400)) + ((!g4) & (!g2) & (g3398) & (g3279) & (g3393) & (!g3400)) + ((!g4) & (!g2) & (g3398) & (g3279) & (g3393) & (g3400)) + ((!g4) & (g2) & (!g3398) & (!g3279) & (!g3393) & (!g3400)) + ((!g4) & (g2) & (g3398) & (!g3279) & (!g3393) & (g3400)) + ((!g4) & (g2) & (g3398) & (!g3279) & (g3393) & (!g3400)) + ((!g4) & (g2) & (g3398) & (!g3279) & (g3393) & (g3400)) + ((!g4) & (g2) & (g3398) & (g3279) & (!g3393) & (!g3400)) + ((!g4) & (g2) & (g3398) & (g3279) & (!g3393) & (g3400)) + ((!g4) & (g2) & (g3398) & (g3279) & (g3393) & (!g3400)) + ((!g4) & (g2) & (g3398) & (g3279) & (g3393) & (g3400)) + ((g4) & (!g2) & (!g3398) & (g3279) & (g3393) & (!g3400)) + ((g4) & (!g2) & (g3398) & (!g3279) & (!g3393) & (!g3400)) + ((g4) & (!g2) & (g3398) & (!g3279) & (!g3393) & (g3400)) + ((g4) & (!g2) & (g3398) & (!g3279) & (g3393) & (!g3400)) + ((g4) & (!g2) & (g3398) & (!g3279) & (g3393) & (g3400)) + ((g4) & (!g2) & (g3398) & (g3279) & (!g3393) & (!g3400)) + ((g4) & (!g2) & (g3398) & (g3279) & (!g3393) & (g3400)) + ((g4) & (!g2) & (g3398) & (g3279) & (g3393) & (g3400)) + ((g4) & (g2) & (!g3398) & (!g3279) & (g3393) & (!g3400)) + ((g4) & (g2) & (!g3398) & (g3279) & (!g3393) & (!g3400)) + ((g4) & (g2) & (!g3398) & (g3279) & (g3393) & (!g3400)) + ((g4) & (g2) & (g3398) & (!g3279) & (!g3393) & (!g3400)) + ((g4) & (g2) & (g3398) & (!g3279) & (!g3393) & (g3400)) + ((g4) & (g2) & (g3398) & (!g3279) & (g3393) & (g3400)) + ((g4) & (g2) & (g3398) & (g3279) & (!g3393) & (g3400)) + ((g4) & (g2) & (g3398) & (g3279) & (g3393) & (g3400)));
	assign g3403 = (((!g8) & (!g18) & (!g3281) & (g3282) & (g3392) & (!g3400)) + ((!g8) & (!g18) & (g3281) & (!g3282) & (!g3392) & (!g3400)) + ((!g8) & (!g18) & (g3281) & (!g3282) & (!g3392) & (g3400)) + ((!g8) & (!g18) & (g3281) & (!g3282) & (g3392) & (!g3400)) + ((!g8) & (!g18) & (g3281) & (!g3282) & (g3392) & (g3400)) + ((!g8) & (!g18) & (g3281) & (g3282) & (!g3392) & (!g3400)) + ((!g8) & (!g18) & (g3281) & (g3282) & (!g3392) & (g3400)) + ((!g8) & (!g18) & (g3281) & (g3282) & (g3392) & (g3400)) + ((!g8) & (g18) & (!g3281) & (!g3282) & (g3392) & (!g3400)) + ((!g8) & (g18) & (!g3281) & (g3282) & (!g3392) & (!g3400)) + ((!g8) & (g18) & (!g3281) & (g3282) & (g3392) & (!g3400)) + ((!g8) & (g18) & (g3281) & (!g3282) & (!g3392) & (!g3400)) + ((!g8) & (g18) & (g3281) & (!g3282) & (!g3392) & (g3400)) + ((!g8) & (g18) & (g3281) & (!g3282) & (g3392) & (g3400)) + ((!g8) & (g18) & (g3281) & (g3282) & (!g3392) & (g3400)) + ((!g8) & (g18) & (g3281) & (g3282) & (g3392) & (g3400)) + ((g8) & (!g18) & (!g3281) & (!g3282) & (!g3392) & (!g3400)) + ((g8) & (!g18) & (!g3281) & (!g3282) & (g3392) & (!g3400)) + ((g8) & (!g18) & (!g3281) & (g3282) & (!g3392) & (!g3400)) + ((g8) & (!g18) & (g3281) & (!g3282) & (!g3392) & (g3400)) + ((g8) & (!g18) & (g3281) & (!g3282) & (g3392) & (g3400)) + ((g8) & (!g18) & (g3281) & (g3282) & (!g3392) & (g3400)) + ((g8) & (!g18) & (g3281) & (g3282) & (g3392) & (!g3400)) + ((g8) & (!g18) & (g3281) & (g3282) & (g3392) & (g3400)) + ((g8) & (g18) & (!g3281) & (!g3282) & (!g3392) & (!g3400)) + ((g8) & (g18) & (g3281) & (!g3282) & (!g3392) & (g3400)) + ((g8) & (g18) & (g3281) & (!g3282) & (g3392) & (!g3400)) + ((g8) & (g18) & (g3281) & (!g3282) & (g3392) & (g3400)) + ((g8) & (g18) & (g3281) & (g3282) & (!g3392) & (!g3400)) + ((g8) & (g18) & (g3281) & (g3282) & (!g3392) & (g3400)) + ((g8) & (g18) & (g3281) & (g3282) & (g3392) & (!g3400)) + ((g8) & (g18) & (g3281) & (g3282) & (g3392) & (g3400)));
	assign g3404 = (((!g18) & (!g3282) & (g3392) & (!g3400)) + ((!g18) & (g3282) & (!g3392) & (!g3400)) + ((!g18) & (g3282) & (!g3392) & (g3400)) + ((!g18) & (g3282) & (g3392) & (g3400)) + ((g18) & (!g3282) & (!g3392) & (!g3400)) + ((g18) & (g3282) & (!g3392) & (g3400)) + ((g18) & (g3282) & (g3392) & (!g3400)) + ((g18) & (g3282) & (g3392) & (g3400)));
	assign g3405 = (((!g27) & (!g39) & (!g3284) & (g3285) & (g3391) & (!g3400)) + ((!g27) & (!g39) & (g3284) & (!g3285) & (!g3391) & (!g3400)) + ((!g27) & (!g39) & (g3284) & (!g3285) & (!g3391) & (g3400)) + ((!g27) & (!g39) & (g3284) & (!g3285) & (g3391) & (!g3400)) + ((!g27) & (!g39) & (g3284) & (!g3285) & (g3391) & (g3400)) + ((!g27) & (!g39) & (g3284) & (g3285) & (!g3391) & (!g3400)) + ((!g27) & (!g39) & (g3284) & (g3285) & (!g3391) & (g3400)) + ((!g27) & (!g39) & (g3284) & (g3285) & (g3391) & (g3400)) + ((!g27) & (g39) & (!g3284) & (!g3285) & (g3391) & (!g3400)) + ((!g27) & (g39) & (!g3284) & (g3285) & (!g3391) & (!g3400)) + ((!g27) & (g39) & (!g3284) & (g3285) & (g3391) & (!g3400)) + ((!g27) & (g39) & (g3284) & (!g3285) & (!g3391) & (!g3400)) + ((!g27) & (g39) & (g3284) & (!g3285) & (!g3391) & (g3400)) + ((!g27) & (g39) & (g3284) & (!g3285) & (g3391) & (g3400)) + ((!g27) & (g39) & (g3284) & (g3285) & (!g3391) & (g3400)) + ((!g27) & (g39) & (g3284) & (g3285) & (g3391) & (g3400)) + ((g27) & (!g39) & (!g3284) & (!g3285) & (!g3391) & (!g3400)) + ((g27) & (!g39) & (!g3284) & (!g3285) & (g3391) & (!g3400)) + ((g27) & (!g39) & (!g3284) & (g3285) & (!g3391) & (!g3400)) + ((g27) & (!g39) & (g3284) & (!g3285) & (!g3391) & (g3400)) + ((g27) & (!g39) & (g3284) & (!g3285) & (g3391) & (g3400)) + ((g27) & (!g39) & (g3284) & (g3285) & (!g3391) & (g3400)) + ((g27) & (!g39) & (g3284) & (g3285) & (g3391) & (!g3400)) + ((g27) & (!g39) & (g3284) & (g3285) & (g3391) & (g3400)) + ((g27) & (g39) & (!g3284) & (!g3285) & (!g3391) & (!g3400)) + ((g27) & (g39) & (g3284) & (!g3285) & (!g3391) & (g3400)) + ((g27) & (g39) & (g3284) & (!g3285) & (g3391) & (!g3400)) + ((g27) & (g39) & (g3284) & (!g3285) & (g3391) & (g3400)) + ((g27) & (g39) & (g3284) & (g3285) & (!g3391) & (!g3400)) + ((g27) & (g39) & (g3284) & (g3285) & (!g3391) & (g3400)) + ((g27) & (g39) & (g3284) & (g3285) & (g3391) & (!g3400)) + ((g27) & (g39) & (g3284) & (g3285) & (g3391) & (g3400)));
	assign g3406 = (((!g39) & (!g3285) & (g3391) & (!g3400)) + ((!g39) & (g3285) & (!g3391) & (!g3400)) + ((!g39) & (g3285) & (!g3391) & (g3400)) + ((!g39) & (g3285) & (g3391) & (g3400)) + ((g39) & (!g3285) & (!g3391) & (!g3400)) + ((g39) & (g3285) & (!g3391) & (g3400)) + ((g39) & (g3285) & (g3391) & (!g3400)) + ((g39) & (g3285) & (g3391) & (g3400)));
	assign g3407 = (((!g54) & (!g68) & (!g3287) & (g3288) & (g3390) & (!g3400)) + ((!g54) & (!g68) & (g3287) & (!g3288) & (!g3390) & (!g3400)) + ((!g54) & (!g68) & (g3287) & (!g3288) & (!g3390) & (g3400)) + ((!g54) & (!g68) & (g3287) & (!g3288) & (g3390) & (!g3400)) + ((!g54) & (!g68) & (g3287) & (!g3288) & (g3390) & (g3400)) + ((!g54) & (!g68) & (g3287) & (g3288) & (!g3390) & (!g3400)) + ((!g54) & (!g68) & (g3287) & (g3288) & (!g3390) & (g3400)) + ((!g54) & (!g68) & (g3287) & (g3288) & (g3390) & (g3400)) + ((!g54) & (g68) & (!g3287) & (!g3288) & (g3390) & (!g3400)) + ((!g54) & (g68) & (!g3287) & (g3288) & (!g3390) & (!g3400)) + ((!g54) & (g68) & (!g3287) & (g3288) & (g3390) & (!g3400)) + ((!g54) & (g68) & (g3287) & (!g3288) & (!g3390) & (!g3400)) + ((!g54) & (g68) & (g3287) & (!g3288) & (!g3390) & (g3400)) + ((!g54) & (g68) & (g3287) & (!g3288) & (g3390) & (g3400)) + ((!g54) & (g68) & (g3287) & (g3288) & (!g3390) & (g3400)) + ((!g54) & (g68) & (g3287) & (g3288) & (g3390) & (g3400)) + ((g54) & (!g68) & (!g3287) & (!g3288) & (!g3390) & (!g3400)) + ((g54) & (!g68) & (!g3287) & (!g3288) & (g3390) & (!g3400)) + ((g54) & (!g68) & (!g3287) & (g3288) & (!g3390) & (!g3400)) + ((g54) & (!g68) & (g3287) & (!g3288) & (!g3390) & (g3400)) + ((g54) & (!g68) & (g3287) & (!g3288) & (g3390) & (g3400)) + ((g54) & (!g68) & (g3287) & (g3288) & (!g3390) & (g3400)) + ((g54) & (!g68) & (g3287) & (g3288) & (g3390) & (!g3400)) + ((g54) & (!g68) & (g3287) & (g3288) & (g3390) & (g3400)) + ((g54) & (g68) & (!g3287) & (!g3288) & (!g3390) & (!g3400)) + ((g54) & (g68) & (g3287) & (!g3288) & (!g3390) & (g3400)) + ((g54) & (g68) & (g3287) & (!g3288) & (g3390) & (!g3400)) + ((g54) & (g68) & (g3287) & (!g3288) & (g3390) & (g3400)) + ((g54) & (g68) & (g3287) & (g3288) & (!g3390) & (!g3400)) + ((g54) & (g68) & (g3287) & (g3288) & (!g3390) & (g3400)) + ((g54) & (g68) & (g3287) & (g3288) & (g3390) & (!g3400)) + ((g54) & (g68) & (g3287) & (g3288) & (g3390) & (g3400)));
	assign g3408 = (((!g68) & (!g3288) & (g3390) & (!g3400)) + ((!g68) & (g3288) & (!g3390) & (!g3400)) + ((!g68) & (g3288) & (!g3390) & (g3400)) + ((!g68) & (g3288) & (g3390) & (g3400)) + ((g68) & (!g3288) & (!g3390) & (!g3400)) + ((g68) & (g3288) & (!g3390) & (g3400)) + ((g68) & (g3288) & (g3390) & (!g3400)) + ((g68) & (g3288) & (g3390) & (g3400)));
	assign g3409 = (((!g87) & (!g104) & (!g3290) & (g3291) & (g3389) & (!g3400)) + ((!g87) & (!g104) & (g3290) & (!g3291) & (!g3389) & (!g3400)) + ((!g87) & (!g104) & (g3290) & (!g3291) & (!g3389) & (g3400)) + ((!g87) & (!g104) & (g3290) & (!g3291) & (g3389) & (!g3400)) + ((!g87) & (!g104) & (g3290) & (!g3291) & (g3389) & (g3400)) + ((!g87) & (!g104) & (g3290) & (g3291) & (!g3389) & (!g3400)) + ((!g87) & (!g104) & (g3290) & (g3291) & (!g3389) & (g3400)) + ((!g87) & (!g104) & (g3290) & (g3291) & (g3389) & (g3400)) + ((!g87) & (g104) & (!g3290) & (!g3291) & (g3389) & (!g3400)) + ((!g87) & (g104) & (!g3290) & (g3291) & (!g3389) & (!g3400)) + ((!g87) & (g104) & (!g3290) & (g3291) & (g3389) & (!g3400)) + ((!g87) & (g104) & (g3290) & (!g3291) & (!g3389) & (!g3400)) + ((!g87) & (g104) & (g3290) & (!g3291) & (!g3389) & (g3400)) + ((!g87) & (g104) & (g3290) & (!g3291) & (g3389) & (g3400)) + ((!g87) & (g104) & (g3290) & (g3291) & (!g3389) & (g3400)) + ((!g87) & (g104) & (g3290) & (g3291) & (g3389) & (g3400)) + ((g87) & (!g104) & (!g3290) & (!g3291) & (!g3389) & (!g3400)) + ((g87) & (!g104) & (!g3290) & (!g3291) & (g3389) & (!g3400)) + ((g87) & (!g104) & (!g3290) & (g3291) & (!g3389) & (!g3400)) + ((g87) & (!g104) & (g3290) & (!g3291) & (!g3389) & (g3400)) + ((g87) & (!g104) & (g3290) & (!g3291) & (g3389) & (g3400)) + ((g87) & (!g104) & (g3290) & (g3291) & (!g3389) & (g3400)) + ((g87) & (!g104) & (g3290) & (g3291) & (g3389) & (!g3400)) + ((g87) & (!g104) & (g3290) & (g3291) & (g3389) & (g3400)) + ((g87) & (g104) & (!g3290) & (!g3291) & (!g3389) & (!g3400)) + ((g87) & (g104) & (g3290) & (!g3291) & (!g3389) & (g3400)) + ((g87) & (g104) & (g3290) & (!g3291) & (g3389) & (!g3400)) + ((g87) & (g104) & (g3290) & (!g3291) & (g3389) & (g3400)) + ((g87) & (g104) & (g3290) & (g3291) & (!g3389) & (!g3400)) + ((g87) & (g104) & (g3290) & (g3291) & (!g3389) & (g3400)) + ((g87) & (g104) & (g3290) & (g3291) & (g3389) & (!g3400)) + ((g87) & (g104) & (g3290) & (g3291) & (g3389) & (g3400)));
	assign g3410 = (((!g104) & (!g3291) & (g3389) & (!g3400)) + ((!g104) & (g3291) & (!g3389) & (!g3400)) + ((!g104) & (g3291) & (!g3389) & (g3400)) + ((!g104) & (g3291) & (g3389) & (g3400)) + ((g104) & (!g3291) & (!g3389) & (!g3400)) + ((g104) & (g3291) & (!g3389) & (g3400)) + ((g104) & (g3291) & (g3389) & (!g3400)) + ((g104) & (g3291) & (g3389) & (g3400)));
	assign g3411 = (((!g127) & (!g147) & (!g3293) & (g3294) & (g3388) & (!g3400)) + ((!g127) & (!g147) & (g3293) & (!g3294) & (!g3388) & (!g3400)) + ((!g127) & (!g147) & (g3293) & (!g3294) & (!g3388) & (g3400)) + ((!g127) & (!g147) & (g3293) & (!g3294) & (g3388) & (!g3400)) + ((!g127) & (!g147) & (g3293) & (!g3294) & (g3388) & (g3400)) + ((!g127) & (!g147) & (g3293) & (g3294) & (!g3388) & (!g3400)) + ((!g127) & (!g147) & (g3293) & (g3294) & (!g3388) & (g3400)) + ((!g127) & (!g147) & (g3293) & (g3294) & (g3388) & (g3400)) + ((!g127) & (g147) & (!g3293) & (!g3294) & (g3388) & (!g3400)) + ((!g127) & (g147) & (!g3293) & (g3294) & (!g3388) & (!g3400)) + ((!g127) & (g147) & (!g3293) & (g3294) & (g3388) & (!g3400)) + ((!g127) & (g147) & (g3293) & (!g3294) & (!g3388) & (!g3400)) + ((!g127) & (g147) & (g3293) & (!g3294) & (!g3388) & (g3400)) + ((!g127) & (g147) & (g3293) & (!g3294) & (g3388) & (g3400)) + ((!g127) & (g147) & (g3293) & (g3294) & (!g3388) & (g3400)) + ((!g127) & (g147) & (g3293) & (g3294) & (g3388) & (g3400)) + ((g127) & (!g147) & (!g3293) & (!g3294) & (!g3388) & (!g3400)) + ((g127) & (!g147) & (!g3293) & (!g3294) & (g3388) & (!g3400)) + ((g127) & (!g147) & (!g3293) & (g3294) & (!g3388) & (!g3400)) + ((g127) & (!g147) & (g3293) & (!g3294) & (!g3388) & (g3400)) + ((g127) & (!g147) & (g3293) & (!g3294) & (g3388) & (g3400)) + ((g127) & (!g147) & (g3293) & (g3294) & (!g3388) & (g3400)) + ((g127) & (!g147) & (g3293) & (g3294) & (g3388) & (!g3400)) + ((g127) & (!g147) & (g3293) & (g3294) & (g3388) & (g3400)) + ((g127) & (g147) & (!g3293) & (!g3294) & (!g3388) & (!g3400)) + ((g127) & (g147) & (g3293) & (!g3294) & (!g3388) & (g3400)) + ((g127) & (g147) & (g3293) & (!g3294) & (g3388) & (!g3400)) + ((g127) & (g147) & (g3293) & (!g3294) & (g3388) & (g3400)) + ((g127) & (g147) & (g3293) & (g3294) & (!g3388) & (!g3400)) + ((g127) & (g147) & (g3293) & (g3294) & (!g3388) & (g3400)) + ((g127) & (g147) & (g3293) & (g3294) & (g3388) & (!g3400)) + ((g127) & (g147) & (g3293) & (g3294) & (g3388) & (g3400)));
	assign g3412 = (((!g147) & (!g3294) & (g3388) & (!g3400)) + ((!g147) & (g3294) & (!g3388) & (!g3400)) + ((!g147) & (g3294) & (!g3388) & (g3400)) + ((!g147) & (g3294) & (g3388) & (g3400)) + ((g147) & (!g3294) & (!g3388) & (!g3400)) + ((g147) & (g3294) & (!g3388) & (g3400)) + ((g147) & (g3294) & (g3388) & (!g3400)) + ((g147) & (g3294) & (g3388) & (g3400)));
	assign g3413 = (((!g174) & (!g198) & (!g3296) & (g3297) & (g3387) & (!g3400)) + ((!g174) & (!g198) & (g3296) & (!g3297) & (!g3387) & (!g3400)) + ((!g174) & (!g198) & (g3296) & (!g3297) & (!g3387) & (g3400)) + ((!g174) & (!g198) & (g3296) & (!g3297) & (g3387) & (!g3400)) + ((!g174) & (!g198) & (g3296) & (!g3297) & (g3387) & (g3400)) + ((!g174) & (!g198) & (g3296) & (g3297) & (!g3387) & (!g3400)) + ((!g174) & (!g198) & (g3296) & (g3297) & (!g3387) & (g3400)) + ((!g174) & (!g198) & (g3296) & (g3297) & (g3387) & (g3400)) + ((!g174) & (g198) & (!g3296) & (!g3297) & (g3387) & (!g3400)) + ((!g174) & (g198) & (!g3296) & (g3297) & (!g3387) & (!g3400)) + ((!g174) & (g198) & (!g3296) & (g3297) & (g3387) & (!g3400)) + ((!g174) & (g198) & (g3296) & (!g3297) & (!g3387) & (!g3400)) + ((!g174) & (g198) & (g3296) & (!g3297) & (!g3387) & (g3400)) + ((!g174) & (g198) & (g3296) & (!g3297) & (g3387) & (g3400)) + ((!g174) & (g198) & (g3296) & (g3297) & (!g3387) & (g3400)) + ((!g174) & (g198) & (g3296) & (g3297) & (g3387) & (g3400)) + ((g174) & (!g198) & (!g3296) & (!g3297) & (!g3387) & (!g3400)) + ((g174) & (!g198) & (!g3296) & (!g3297) & (g3387) & (!g3400)) + ((g174) & (!g198) & (!g3296) & (g3297) & (!g3387) & (!g3400)) + ((g174) & (!g198) & (g3296) & (!g3297) & (!g3387) & (g3400)) + ((g174) & (!g198) & (g3296) & (!g3297) & (g3387) & (g3400)) + ((g174) & (!g198) & (g3296) & (g3297) & (!g3387) & (g3400)) + ((g174) & (!g198) & (g3296) & (g3297) & (g3387) & (!g3400)) + ((g174) & (!g198) & (g3296) & (g3297) & (g3387) & (g3400)) + ((g174) & (g198) & (!g3296) & (!g3297) & (!g3387) & (!g3400)) + ((g174) & (g198) & (g3296) & (!g3297) & (!g3387) & (g3400)) + ((g174) & (g198) & (g3296) & (!g3297) & (g3387) & (!g3400)) + ((g174) & (g198) & (g3296) & (!g3297) & (g3387) & (g3400)) + ((g174) & (g198) & (g3296) & (g3297) & (!g3387) & (!g3400)) + ((g174) & (g198) & (g3296) & (g3297) & (!g3387) & (g3400)) + ((g174) & (g198) & (g3296) & (g3297) & (g3387) & (!g3400)) + ((g174) & (g198) & (g3296) & (g3297) & (g3387) & (g3400)));
	assign g3414 = (((!g198) & (!g3297) & (g3387) & (!g3400)) + ((!g198) & (g3297) & (!g3387) & (!g3400)) + ((!g198) & (g3297) & (!g3387) & (g3400)) + ((!g198) & (g3297) & (g3387) & (g3400)) + ((g198) & (!g3297) & (!g3387) & (!g3400)) + ((g198) & (g3297) & (!g3387) & (g3400)) + ((g198) & (g3297) & (g3387) & (!g3400)) + ((g198) & (g3297) & (g3387) & (g3400)));
	assign g3415 = (((!g229) & (!g255) & (!g3299) & (g3300) & (g3386) & (!g3400)) + ((!g229) & (!g255) & (g3299) & (!g3300) & (!g3386) & (!g3400)) + ((!g229) & (!g255) & (g3299) & (!g3300) & (!g3386) & (g3400)) + ((!g229) & (!g255) & (g3299) & (!g3300) & (g3386) & (!g3400)) + ((!g229) & (!g255) & (g3299) & (!g3300) & (g3386) & (g3400)) + ((!g229) & (!g255) & (g3299) & (g3300) & (!g3386) & (!g3400)) + ((!g229) & (!g255) & (g3299) & (g3300) & (!g3386) & (g3400)) + ((!g229) & (!g255) & (g3299) & (g3300) & (g3386) & (g3400)) + ((!g229) & (g255) & (!g3299) & (!g3300) & (g3386) & (!g3400)) + ((!g229) & (g255) & (!g3299) & (g3300) & (!g3386) & (!g3400)) + ((!g229) & (g255) & (!g3299) & (g3300) & (g3386) & (!g3400)) + ((!g229) & (g255) & (g3299) & (!g3300) & (!g3386) & (!g3400)) + ((!g229) & (g255) & (g3299) & (!g3300) & (!g3386) & (g3400)) + ((!g229) & (g255) & (g3299) & (!g3300) & (g3386) & (g3400)) + ((!g229) & (g255) & (g3299) & (g3300) & (!g3386) & (g3400)) + ((!g229) & (g255) & (g3299) & (g3300) & (g3386) & (g3400)) + ((g229) & (!g255) & (!g3299) & (!g3300) & (!g3386) & (!g3400)) + ((g229) & (!g255) & (!g3299) & (!g3300) & (g3386) & (!g3400)) + ((g229) & (!g255) & (!g3299) & (g3300) & (!g3386) & (!g3400)) + ((g229) & (!g255) & (g3299) & (!g3300) & (!g3386) & (g3400)) + ((g229) & (!g255) & (g3299) & (!g3300) & (g3386) & (g3400)) + ((g229) & (!g255) & (g3299) & (g3300) & (!g3386) & (g3400)) + ((g229) & (!g255) & (g3299) & (g3300) & (g3386) & (!g3400)) + ((g229) & (!g255) & (g3299) & (g3300) & (g3386) & (g3400)) + ((g229) & (g255) & (!g3299) & (!g3300) & (!g3386) & (!g3400)) + ((g229) & (g255) & (g3299) & (!g3300) & (!g3386) & (g3400)) + ((g229) & (g255) & (g3299) & (!g3300) & (g3386) & (!g3400)) + ((g229) & (g255) & (g3299) & (!g3300) & (g3386) & (g3400)) + ((g229) & (g255) & (g3299) & (g3300) & (!g3386) & (!g3400)) + ((g229) & (g255) & (g3299) & (g3300) & (!g3386) & (g3400)) + ((g229) & (g255) & (g3299) & (g3300) & (g3386) & (!g3400)) + ((g229) & (g255) & (g3299) & (g3300) & (g3386) & (g3400)));
	assign g3416 = (((!g255) & (!g3300) & (g3386) & (!g3400)) + ((!g255) & (g3300) & (!g3386) & (!g3400)) + ((!g255) & (g3300) & (!g3386) & (g3400)) + ((!g255) & (g3300) & (g3386) & (g3400)) + ((g255) & (!g3300) & (!g3386) & (!g3400)) + ((g255) & (g3300) & (!g3386) & (g3400)) + ((g255) & (g3300) & (g3386) & (!g3400)) + ((g255) & (g3300) & (g3386) & (g3400)));
	assign g3417 = (((!g290) & (!g319) & (!g3302) & (g3303) & (g3385) & (!g3400)) + ((!g290) & (!g319) & (g3302) & (!g3303) & (!g3385) & (!g3400)) + ((!g290) & (!g319) & (g3302) & (!g3303) & (!g3385) & (g3400)) + ((!g290) & (!g319) & (g3302) & (!g3303) & (g3385) & (!g3400)) + ((!g290) & (!g319) & (g3302) & (!g3303) & (g3385) & (g3400)) + ((!g290) & (!g319) & (g3302) & (g3303) & (!g3385) & (!g3400)) + ((!g290) & (!g319) & (g3302) & (g3303) & (!g3385) & (g3400)) + ((!g290) & (!g319) & (g3302) & (g3303) & (g3385) & (g3400)) + ((!g290) & (g319) & (!g3302) & (!g3303) & (g3385) & (!g3400)) + ((!g290) & (g319) & (!g3302) & (g3303) & (!g3385) & (!g3400)) + ((!g290) & (g319) & (!g3302) & (g3303) & (g3385) & (!g3400)) + ((!g290) & (g319) & (g3302) & (!g3303) & (!g3385) & (!g3400)) + ((!g290) & (g319) & (g3302) & (!g3303) & (!g3385) & (g3400)) + ((!g290) & (g319) & (g3302) & (!g3303) & (g3385) & (g3400)) + ((!g290) & (g319) & (g3302) & (g3303) & (!g3385) & (g3400)) + ((!g290) & (g319) & (g3302) & (g3303) & (g3385) & (g3400)) + ((g290) & (!g319) & (!g3302) & (!g3303) & (!g3385) & (!g3400)) + ((g290) & (!g319) & (!g3302) & (!g3303) & (g3385) & (!g3400)) + ((g290) & (!g319) & (!g3302) & (g3303) & (!g3385) & (!g3400)) + ((g290) & (!g319) & (g3302) & (!g3303) & (!g3385) & (g3400)) + ((g290) & (!g319) & (g3302) & (!g3303) & (g3385) & (g3400)) + ((g290) & (!g319) & (g3302) & (g3303) & (!g3385) & (g3400)) + ((g290) & (!g319) & (g3302) & (g3303) & (g3385) & (!g3400)) + ((g290) & (!g319) & (g3302) & (g3303) & (g3385) & (g3400)) + ((g290) & (g319) & (!g3302) & (!g3303) & (!g3385) & (!g3400)) + ((g290) & (g319) & (g3302) & (!g3303) & (!g3385) & (g3400)) + ((g290) & (g319) & (g3302) & (!g3303) & (g3385) & (!g3400)) + ((g290) & (g319) & (g3302) & (!g3303) & (g3385) & (g3400)) + ((g290) & (g319) & (g3302) & (g3303) & (!g3385) & (!g3400)) + ((g290) & (g319) & (g3302) & (g3303) & (!g3385) & (g3400)) + ((g290) & (g319) & (g3302) & (g3303) & (g3385) & (!g3400)) + ((g290) & (g319) & (g3302) & (g3303) & (g3385) & (g3400)));
	assign g3418 = (((!g319) & (!g3303) & (g3385) & (!g3400)) + ((!g319) & (g3303) & (!g3385) & (!g3400)) + ((!g319) & (g3303) & (!g3385) & (g3400)) + ((!g319) & (g3303) & (g3385) & (g3400)) + ((g319) & (!g3303) & (!g3385) & (!g3400)) + ((g319) & (g3303) & (!g3385) & (g3400)) + ((g319) & (g3303) & (g3385) & (!g3400)) + ((g319) & (g3303) & (g3385) & (g3400)));
	assign g3419 = (((!g358) & (!g390) & (!g3305) & (g3306) & (g3384) & (!g3400)) + ((!g358) & (!g390) & (g3305) & (!g3306) & (!g3384) & (!g3400)) + ((!g358) & (!g390) & (g3305) & (!g3306) & (!g3384) & (g3400)) + ((!g358) & (!g390) & (g3305) & (!g3306) & (g3384) & (!g3400)) + ((!g358) & (!g390) & (g3305) & (!g3306) & (g3384) & (g3400)) + ((!g358) & (!g390) & (g3305) & (g3306) & (!g3384) & (!g3400)) + ((!g358) & (!g390) & (g3305) & (g3306) & (!g3384) & (g3400)) + ((!g358) & (!g390) & (g3305) & (g3306) & (g3384) & (g3400)) + ((!g358) & (g390) & (!g3305) & (!g3306) & (g3384) & (!g3400)) + ((!g358) & (g390) & (!g3305) & (g3306) & (!g3384) & (!g3400)) + ((!g358) & (g390) & (!g3305) & (g3306) & (g3384) & (!g3400)) + ((!g358) & (g390) & (g3305) & (!g3306) & (!g3384) & (!g3400)) + ((!g358) & (g390) & (g3305) & (!g3306) & (!g3384) & (g3400)) + ((!g358) & (g390) & (g3305) & (!g3306) & (g3384) & (g3400)) + ((!g358) & (g390) & (g3305) & (g3306) & (!g3384) & (g3400)) + ((!g358) & (g390) & (g3305) & (g3306) & (g3384) & (g3400)) + ((g358) & (!g390) & (!g3305) & (!g3306) & (!g3384) & (!g3400)) + ((g358) & (!g390) & (!g3305) & (!g3306) & (g3384) & (!g3400)) + ((g358) & (!g390) & (!g3305) & (g3306) & (!g3384) & (!g3400)) + ((g358) & (!g390) & (g3305) & (!g3306) & (!g3384) & (g3400)) + ((g358) & (!g390) & (g3305) & (!g3306) & (g3384) & (g3400)) + ((g358) & (!g390) & (g3305) & (g3306) & (!g3384) & (g3400)) + ((g358) & (!g390) & (g3305) & (g3306) & (g3384) & (!g3400)) + ((g358) & (!g390) & (g3305) & (g3306) & (g3384) & (g3400)) + ((g358) & (g390) & (!g3305) & (!g3306) & (!g3384) & (!g3400)) + ((g358) & (g390) & (g3305) & (!g3306) & (!g3384) & (g3400)) + ((g358) & (g390) & (g3305) & (!g3306) & (g3384) & (!g3400)) + ((g358) & (g390) & (g3305) & (!g3306) & (g3384) & (g3400)) + ((g358) & (g390) & (g3305) & (g3306) & (!g3384) & (!g3400)) + ((g358) & (g390) & (g3305) & (g3306) & (!g3384) & (g3400)) + ((g358) & (g390) & (g3305) & (g3306) & (g3384) & (!g3400)) + ((g358) & (g390) & (g3305) & (g3306) & (g3384) & (g3400)));
	assign g3420 = (((!g390) & (!g3306) & (g3384) & (!g3400)) + ((!g390) & (g3306) & (!g3384) & (!g3400)) + ((!g390) & (g3306) & (!g3384) & (g3400)) + ((!g390) & (g3306) & (g3384) & (g3400)) + ((g390) & (!g3306) & (!g3384) & (!g3400)) + ((g390) & (g3306) & (!g3384) & (g3400)) + ((g390) & (g3306) & (g3384) & (!g3400)) + ((g390) & (g3306) & (g3384) & (g3400)));
	assign g3421 = (((!g433) & (!g468) & (!g3308) & (g3309) & (g3383) & (!g3400)) + ((!g433) & (!g468) & (g3308) & (!g3309) & (!g3383) & (!g3400)) + ((!g433) & (!g468) & (g3308) & (!g3309) & (!g3383) & (g3400)) + ((!g433) & (!g468) & (g3308) & (!g3309) & (g3383) & (!g3400)) + ((!g433) & (!g468) & (g3308) & (!g3309) & (g3383) & (g3400)) + ((!g433) & (!g468) & (g3308) & (g3309) & (!g3383) & (!g3400)) + ((!g433) & (!g468) & (g3308) & (g3309) & (!g3383) & (g3400)) + ((!g433) & (!g468) & (g3308) & (g3309) & (g3383) & (g3400)) + ((!g433) & (g468) & (!g3308) & (!g3309) & (g3383) & (!g3400)) + ((!g433) & (g468) & (!g3308) & (g3309) & (!g3383) & (!g3400)) + ((!g433) & (g468) & (!g3308) & (g3309) & (g3383) & (!g3400)) + ((!g433) & (g468) & (g3308) & (!g3309) & (!g3383) & (!g3400)) + ((!g433) & (g468) & (g3308) & (!g3309) & (!g3383) & (g3400)) + ((!g433) & (g468) & (g3308) & (!g3309) & (g3383) & (g3400)) + ((!g433) & (g468) & (g3308) & (g3309) & (!g3383) & (g3400)) + ((!g433) & (g468) & (g3308) & (g3309) & (g3383) & (g3400)) + ((g433) & (!g468) & (!g3308) & (!g3309) & (!g3383) & (!g3400)) + ((g433) & (!g468) & (!g3308) & (!g3309) & (g3383) & (!g3400)) + ((g433) & (!g468) & (!g3308) & (g3309) & (!g3383) & (!g3400)) + ((g433) & (!g468) & (g3308) & (!g3309) & (!g3383) & (g3400)) + ((g433) & (!g468) & (g3308) & (!g3309) & (g3383) & (g3400)) + ((g433) & (!g468) & (g3308) & (g3309) & (!g3383) & (g3400)) + ((g433) & (!g468) & (g3308) & (g3309) & (g3383) & (!g3400)) + ((g433) & (!g468) & (g3308) & (g3309) & (g3383) & (g3400)) + ((g433) & (g468) & (!g3308) & (!g3309) & (!g3383) & (!g3400)) + ((g433) & (g468) & (g3308) & (!g3309) & (!g3383) & (g3400)) + ((g433) & (g468) & (g3308) & (!g3309) & (g3383) & (!g3400)) + ((g433) & (g468) & (g3308) & (!g3309) & (g3383) & (g3400)) + ((g433) & (g468) & (g3308) & (g3309) & (!g3383) & (!g3400)) + ((g433) & (g468) & (g3308) & (g3309) & (!g3383) & (g3400)) + ((g433) & (g468) & (g3308) & (g3309) & (g3383) & (!g3400)) + ((g433) & (g468) & (g3308) & (g3309) & (g3383) & (g3400)));
	assign g3422 = (((!g468) & (!g3309) & (g3383) & (!g3400)) + ((!g468) & (g3309) & (!g3383) & (!g3400)) + ((!g468) & (g3309) & (!g3383) & (g3400)) + ((!g468) & (g3309) & (g3383) & (g3400)) + ((g468) & (!g3309) & (!g3383) & (!g3400)) + ((g468) & (g3309) & (!g3383) & (g3400)) + ((g468) & (g3309) & (g3383) & (!g3400)) + ((g468) & (g3309) & (g3383) & (g3400)));
	assign g3423 = (((!g515) & (!g553) & (!g3311) & (g3312) & (g3382) & (!g3400)) + ((!g515) & (!g553) & (g3311) & (!g3312) & (!g3382) & (!g3400)) + ((!g515) & (!g553) & (g3311) & (!g3312) & (!g3382) & (g3400)) + ((!g515) & (!g553) & (g3311) & (!g3312) & (g3382) & (!g3400)) + ((!g515) & (!g553) & (g3311) & (!g3312) & (g3382) & (g3400)) + ((!g515) & (!g553) & (g3311) & (g3312) & (!g3382) & (!g3400)) + ((!g515) & (!g553) & (g3311) & (g3312) & (!g3382) & (g3400)) + ((!g515) & (!g553) & (g3311) & (g3312) & (g3382) & (g3400)) + ((!g515) & (g553) & (!g3311) & (!g3312) & (g3382) & (!g3400)) + ((!g515) & (g553) & (!g3311) & (g3312) & (!g3382) & (!g3400)) + ((!g515) & (g553) & (!g3311) & (g3312) & (g3382) & (!g3400)) + ((!g515) & (g553) & (g3311) & (!g3312) & (!g3382) & (!g3400)) + ((!g515) & (g553) & (g3311) & (!g3312) & (!g3382) & (g3400)) + ((!g515) & (g553) & (g3311) & (!g3312) & (g3382) & (g3400)) + ((!g515) & (g553) & (g3311) & (g3312) & (!g3382) & (g3400)) + ((!g515) & (g553) & (g3311) & (g3312) & (g3382) & (g3400)) + ((g515) & (!g553) & (!g3311) & (!g3312) & (!g3382) & (!g3400)) + ((g515) & (!g553) & (!g3311) & (!g3312) & (g3382) & (!g3400)) + ((g515) & (!g553) & (!g3311) & (g3312) & (!g3382) & (!g3400)) + ((g515) & (!g553) & (g3311) & (!g3312) & (!g3382) & (g3400)) + ((g515) & (!g553) & (g3311) & (!g3312) & (g3382) & (g3400)) + ((g515) & (!g553) & (g3311) & (g3312) & (!g3382) & (g3400)) + ((g515) & (!g553) & (g3311) & (g3312) & (g3382) & (!g3400)) + ((g515) & (!g553) & (g3311) & (g3312) & (g3382) & (g3400)) + ((g515) & (g553) & (!g3311) & (!g3312) & (!g3382) & (!g3400)) + ((g515) & (g553) & (g3311) & (!g3312) & (!g3382) & (g3400)) + ((g515) & (g553) & (g3311) & (!g3312) & (g3382) & (!g3400)) + ((g515) & (g553) & (g3311) & (!g3312) & (g3382) & (g3400)) + ((g515) & (g553) & (g3311) & (g3312) & (!g3382) & (!g3400)) + ((g515) & (g553) & (g3311) & (g3312) & (!g3382) & (g3400)) + ((g515) & (g553) & (g3311) & (g3312) & (g3382) & (!g3400)) + ((g515) & (g553) & (g3311) & (g3312) & (g3382) & (g3400)));
	assign g3424 = (((!g553) & (!g3312) & (g3382) & (!g3400)) + ((!g553) & (g3312) & (!g3382) & (!g3400)) + ((!g553) & (g3312) & (!g3382) & (g3400)) + ((!g553) & (g3312) & (g3382) & (g3400)) + ((g553) & (!g3312) & (!g3382) & (!g3400)) + ((g553) & (g3312) & (!g3382) & (g3400)) + ((g553) & (g3312) & (g3382) & (!g3400)) + ((g553) & (g3312) & (g3382) & (g3400)));
	assign g3425 = (((!g604) & (!g645) & (!g3314) & (g3315) & (g3381) & (!g3400)) + ((!g604) & (!g645) & (g3314) & (!g3315) & (!g3381) & (!g3400)) + ((!g604) & (!g645) & (g3314) & (!g3315) & (!g3381) & (g3400)) + ((!g604) & (!g645) & (g3314) & (!g3315) & (g3381) & (!g3400)) + ((!g604) & (!g645) & (g3314) & (!g3315) & (g3381) & (g3400)) + ((!g604) & (!g645) & (g3314) & (g3315) & (!g3381) & (!g3400)) + ((!g604) & (!g645) & (g3314) & (g3315) & (!g3381) & (g3400)) + ((!g604) & (!g645) & (g3314) & (g3315) & (g3381) & (g3400)) + ((!g604) & (g645) & (!g3314) & (!g3315) & (g3381) & (!g3400)) + ((!g604) & (g645) & (!g3314) & (g3315) & (!g3381) & (!g3400)) + ((!g604) & (g645) & (!g3314) & (g3315) & (g3381) & (!g3400)) + ((!g604) & (g645) & (g3314) & (!g3315) & (!g3381) & (!g3400)) + ((!g604) & (g645) & (g3314) & (!g3315) & (!g3381) & (g3400)) + ((!g604) & (g645) & (g3314) & (!g3315) & (g3381) & (g3400)) + ((!g604) & (g645) & (g3314) & (g3315) & (!g3381) & (g3400)) + ((!g604) & (g645) & (g3314) & (g3315) & (g3381) & (g3400)) + ((g604) & (!g645) & (!g3314) & (!g3315) & (!g3381) & (!g3400)) + ((g604) & (!g645) & (!g3314) & (!g3315) & (g3381) & (!g3400)) + ((g604) & (!g645) & (!g3314) & (g3315) & (!g3381) & (!g3400)) + ((g604) & (!g645) & (g3314) & (!g3315) & (!g3381) & (g3400)) + ((g604) & (!g645) & (g3314) & (!g3315) & (g3381) & (g3400)) + ((g604) & (!g645) & (g3314) & (g3315) & (!g3381) & (g3400)) + ((g604) & (!g645) & (g3314) & (g3315) & (g3381) & (!g3400)) + ((g604) & (!g645) & (g3314) & (g3315) & (g3381) & (g3400)) + ((g604) & (g645) & (!g3314) & (!g3315) & (!g3381) & (!g3400)) + ((g604) & (g645) & (g3314) & (!g3315) & (!g3381) & (g3400)) + ((g604) & (g645) & (g3314) & (!g3315) & (g3381) & (!g3400)) + ((g604) & (g645) & (g3314) & (!g3315) & (g3381) & (g3400)) + ((g604) & (g645) & (g3314) & (g3315) & (!g3381) & (!g3400)) + ((g604) & (g645) & (g3314) & (g3315) & (!g3381) & (g3400)) + ((g604) & (g645) & (g3314) & (g3315) & (g3381) & (!g3400)) + ((g604) & (g645) & (g3314) & (g3315) & (g3381) & (g3400)));
	assign g3426 = (((!g645) & (!g3315) & (g3381) & (!g3400)) + ((!g645) & (g3315) & (!g3381) & (!g3400)) + ((!g645) & (g3315) & (!g3381) & (g3400)) + ((!g645) & (g3315) & (g3381) & (g3400)) + ((g645) & (!g3315) & (!g3381) & (!g3400)) + ((g645) & (g3315) & (!g3381) & (g3400)) + ((g645) & (g3315) & (g3381) & (!g3400)) + ((g645) & (g3315) & (g3381) & (g3400)));
	assign g3427 = (((!g700) & (!g744) & (!g3317) & (g3318) & (g3380) & (!g3400)) + ((!g700) & (!g744) & (g3317) & (!g3318) & (!g3380) & (!g3400)) + ((!g700) & (!g744) & (g3317) & (!g3318) & (!g3380) & (g3400)) + ((!g700) & (!g744) & (g3317) & (!g3318) & (g3380) & (!g3400)) + ((!g700) & (!g744) & (g3317) & (!g3318) & (g3380) & (g3400)) + ((!g700) & (!g744) & (g3317) & (g3318) & (!g3380) & (!g3400)) + ((!g700) & (!g744) & (g3317) & (g3318) & (!g3380) & (g3400)) + ((!g700) & (!g744) & (g3317) & (g3318) & (g3380) & (g3400)) + ((!g700) & (g744) & (!g3317) & (!g3318) & (g3380) & (!g3400)) + ((!g700) & (g744) & (!g3317) & (g3318) & (!g3380) & (!g3400)) + ((!g700) & (g744) & (!g3317) & (g3318) & (g3380) & (!g3400)) + ((!g700) & (g744) & (g3317) & (!g3318) & (!g3380) & (!g3400)) + ((!g700) & (g744) & (g3317) & (!g3318) & (!g3380) & (g3400)) + ((!g700) & (g744) & (g3317) & (!g3318) & (g3380) & (g3400)) + ((!g700) & (g744) & (g3317) & (g3318) & (!g3380) & (g3400)) + ((!g700) & (g744) & (g3317) & (g3318) & (g3380) & (g3400)) + ((g700) & (!g744) & (!g3317) & (!g3318) & (!g3380) & (!g3400)) + ((g700) & (!g744) & (!g3317) & (!g3318) & (g3380) & (!g3400)) + ((g700) & (!g744) & (!g3317) & (g3318) & (!g3380) & (!g3400)) + ((g700) & (!g744) & (g3317) & (!g3318) & (!g3380) & (g3400)) + ((g700) & (!g744) & (g3317) & (!g3318) & (g3380) & (g3400)) + ((g700) & (!g744) & (g3317) & (g3318) & (!g3380) & (g3400)) + ((g700) & (!g744) & (g3317) & (g3318) & (g3380) & (!g3400)) + ((g700) & (!g744) & (g3317) & (g3318) & (g3380) & (g3400)) + ((g700) & (g744) & (!g3317) & (!g3318) & (!g3380) & (!g3400)) + ((g700) & (g744) & (g3317) & (!g3318) & (!g3380) & (g3400)) + ((g700) & (g744) & (g3317) & (!g3318) & (g3380) & (!g3400)) + ((g700) & (g744) & (g3317) & (!g3318) & (g3380) & (g3400)) + ((g700) & (g744) & (g3317) & (g3318) & (!g3380) & (!g3400)) + ((g700) & (g744) & (g3317) & (g3318) & (!g3380) & (g3400)) + ((g700) & (g744) & (g3317) & (g3318) & (g3380) & (!g3400)) + ((g700) & (g744) & (g3317) & (g3318) & (g3380) & (g3400)));
	assign g3428 = (((!g744) & (!g3318) & (g3380) & (!g3400)) + ((!g744) & (g3318) & (!g3380) & (!g3400)) + ((!g744) & (g3318) & (!g3380) & (g3400)) + ((!g744) & (g3318) & (g3380) & (g3400)) + ((g744) & (!g3318) & (!g3380) & (!g3400)) + ((g744) & (g3318) & (!g3380) & (g3400)) + ((g744) & (g3318) & (g3380) & (!g3400)) + ((g744) & (g3318) & (g3380) & (g3400)));
	assign g3429 = (((!g803) & (!g851) & (!g3320) & (g3321) & (g3379) & (!g3400)) + ((!g803) & (!g851) & (g3320) & (!g3321) & (!g3379) & (!g3400)) + ((!g803) & (!g851) & (g3320) & (!g3321) & (!g3379) & (g3400)) + ((!g803) & (!g851) & (g3320) & (!g3321) & (g3379) & (!g3400)) + ((!g803) & (!g851) & (g3320) & (!g3321) & (g3379) & (g3400)) + ((!g803) & (!g851) & (g3320) & (g3321) & (!g3379) & (!g3400)) + ((!g803) & (!g851) & (g3320) & (g3321) & (!g3379) & (g3400)) + ((!g803) & (!g851) & (g3320) & (g3321) & (g3379) & (g3400)) + ((!g803) & (g851) & (!g3320) & (!g3321) & (g3379) & (!g3400)) + ((!g803) & (g851) & (!g3320) & (g3321) & (!g3379) & (!g3400)) + ((!g803) & (g851) & (!g3320) & (g3321) & (g3379) & (!g3400)) + ((!g803) & (g851) & (g3320) & (!g3321) & (!g3379) & (!g3400)) + ((!g803) & (g851) & (g3320) & (!g3321) & (!g3379) & (g3400)) + ((!g803) & (g851) & (g3320) & (!g3321) & (g3379) & (g3400)) + ((!g803) & (g851) & (g3320) & (g3321) & (!g3379) & (g3400)) + ((!g803) & (g851) & (g3320) & (g3321) & (g3379) & (g3400)) + ((g803) & (!g851) & (!g3320) & (!g3321) & (!g3379) & (!g3400)) + ((g803) & (!g851) & (!g3320) & (!g3321) & (g3379) & (!g3400)) + ((g803) & (!g851) & (!g3320) & (g3321) & (!g3379) & (!g3400)) + ((g803) & (!g851) & (g3320) & (!g3321) & (!g3379) & (g3400)) + ((g803) & (!g851) & (g3320) & (!g3321) & (g3379) & (g3400)) + ((g803) & (!g851) & (g3320) & (g3321) & (!g3379) & (g3400)) + ((g803) & (!g851) & (g3320) & (g3321) & (g3379) & (!g3400)) + ((g803) & (!g851) & (g3320) & (g3321) & (g3379) & (g3400)) + ((g803) & (g851) & (!g3320) & (!g3321) & (!g3379) & (!g3400)) + ((g803) & (g851) & (g3320) & (!g3321) & (!g3379) & (g3400)) + ((g803) & (g851) & (g3320) & (!g3321) & (g3379) & (!g3400)) + ((g803) & (g851) & (g3320) & (!g3321) & (g3379) & (g3400)) + ((g803) & (g851) & (g3320) & (g3321) & (!g3379) & (!g3400)) + ((g803) & (g851) & (g3320) & (g3321) & (!g3379) & (g3400)) + ((g803) & (g851) & (g3320) & (g3321) & (g3379) & (!g3400)) + ((g803) & (g851) & (g3320) & (g3321) & (g3379) & (g3400)));
	assign g3430 = (((!g851) & (!g3321) & (g3379) & (!g3400)) + ((!g851) & (g3321) & (!g3379) & (!g3400)) + ((!g851) & (g3321) & (!g3379) & (g3400)) + ((!g851) & (g3321) & (g3379) & (g3400)) + ((g851) & (!g3321) & (!g3379) & (!g3400)) + ((g851) & (g3321) & (!g3379) & (g3400)) + ((g851) & (g3321) & (g3379) & (!g3400)) + ((g851) & (g3321) & (g3379) & (g3400)));
	assign g3431 = (((!g914) & (!g1032) & (!g3323) & (g3324) & (g3378) & (!g3400)) + ((!g914) & (!g1032) & (g3323) & (!g3324) & (!g3378) & (!g3400)) + ((!g914) & (!g1032) & (g3323) & (!g3324) & (!g3378) & (g3400)) + ((!g914) & (!g1032) & (g3323) & (!g3324) & (g3378) & (!g3400)) + ((!g914) & (!g1032) & (g3323) & (!g3324) & (g3378) & (g3400)) + ((!g914) & (!g1032) & (g3323) & (g3324) & (!g3378) & (!g3400)) + ((!g914) & (!g1032) & (g3323) & (g3324) & (!g3378) & (g3400)) + ((!g914) & (!g1032) & (g3323) & (g3324) & (g3378) & (g3400)) + ((!g914) & (g1032) & (!g3323) & (!g3324) & (g3378) & (!g3400)) + ((!g914) & (g1032) & (!g3323) & (g3324) & (!g3378) & (!g3400)) + ((!g914) & (g1032) & (!g3323) & (g3324) & (g3378) & (!g3400)) + ((!g914) & (g1032) & (g3323) & (!g3324) & (!g3378) & (!g3400)) + ((!g914) & (g1032) & (g3323) & (!g3324) & (!g3378) & (g3400)) + ((!g914) & (g1032) & (g3323) & (!g3324) & (g3378) & (g3400)) + ((!g914) & (g1032) & (g3323) & (g3324) & (!g3378) & (g3400)) + ((!g914) & (g1032) & (g3323) & (g3324) & (g3378) & (g3400)) + ((g914) & (!g1032) & (!g3323) & (!g3324) & (!g3378) & (!g3400)) + ((g914) & (!g1032) & (!g3323) & (!g3324) & (g3378) & (!g3400)) + ((g914) & (!g1032) & (!g3323) & (g3324) & (!g3378) & (!g3400)) + ((g914) & (!g1032) & (g3323) & (!g3324) & (!g3378) & (g3400)) + ((g914) & (!g1032) & (g3323) & (!g3324) & (g3378) & (g3400)) + ((g914) & (!g1032) & (g3323) & (g3324) & (!g3378) & (g3400)) + ((g914) & (!g1032) & (g3323) & (g3324) & (g3378) & (!g3400)) + ((g914) & (!g1032) & (g3323) & (g3324) & (g3378) & (g3400)) + ((g914) & (g1032) & (!g3323) & (!g3324) & (!g3378) & (!g3400)) + ((g914) & (g1032) & (g3323) & (!g3324) & (!g3378) & (g3400)) + ((g914) & (g1032) & (g3323) & (!g3324) & (g3378) & (!g3400)) + ((g914) & (g1032) & (g3323) & (!g3324) & (g3378) & (g3400)) + ((g914) & (g1032) & (g3323) & (g3324) & (!g3378) & (!g3400)) + ((g914) & (g1032) & (g3323) & (g3324) & (!g3378) & (g3400)) + ((g914) & (g1032) & (g3323) & (g3324) & (g3378) & (!g3400)) + ((g914) & (g1032) & (g3323) & (g3324) & (g3378) & (g3400)));
	assign g3432 = (((!g1032) & (!g3324) & (g3378) & (!g3400)) + ((!g1032) & (g3324) & (!g3378) & (!g3400)) + ((!g1032) & (g3324) & (!g3378) & (g3400)) + ((!g1032) & (g3324) & (g3378) & (g3400)) + ((g1032) & (!g3324) & (!g3378) & (!g3400)) + ((g1032) & (g3324) & (!g3378) & (g3400)) + ((g1032) & (g3324) & (g3378) & (!g3400)) + ((g1032) & (g3324) & (g3378) & (g3400)));
	assign g3433 = (((!g1030) & (!g1160) & (!g3326) & (g3327) & (g3377) & (!g3400)) + ((!g1030) & (!g1160) & (g3326) & (!g3327) & (!g3377) & (!g3400)) + ((!g1030) & (!g1160) & (g3326) & (!g3327) & (!g3377) & (g3400)) + ((!g1030) & (!g1160) & (g3326) & (!g3327) & (g3377) & (!g3400)) + ((!g1030) & (!g1160) & (g3326) & (!g3327) & (g3377) & (g3400)) + ((!g1030) & (!g1160) & (g3326) & (g3327) & (!g3377) & (!g3400)) + ((!g1030) & (!g1160) & (g3326) & (g3327) & (!g3377) & (g3400)) + ((!g1030) & (!g1160) & (g3326) & (g3327) & (g3377) & (g3400)) + ((!g1030) & (g1160) & (!g3326) & (!g3327) & (g3377) & (!g3400)) + ((!g1030) & (g1160) & (!g3326) & (g3327) & (!g3377) & (!g3400)) + ((!g1030) & (g1160) & (!g3326) & (g3327) & (g3377) & (!g3400)) + ((!g1030) & (g1160) & (g3326) & (!g3327) & (!g3377) & (!g3400)) + ((!g1030) & (g1160) & (g3326) & (!g3327) & (!g3377) & (g3400)) + ((!g1030) & (g1160) & (g3326) & (!g3327) & (g3377) & (g3400)) + ((!g1030) & (g1160) & (g3326) & (g3327) & (!g3377) & (g3400)) + ((!g1030) & (g1160) & (g3326) & (g3327) & (g3377) & (g3400)) + ((g1030) & (!g1160) & (!g3326) & (!g3327) & (!g3377) & (!g3400)) + ((g1030) & (!g1160) & (!g3326) & (!g3327) & (g3377) & (!g3400)) + ((g1030) & (!g1160) & (!g3326) & (g3327) & (!g3377) & (!g3400)) + ((g1030) & (!g1160) & (g3326) & (!g3327) & (!g3377) & (g3400)) + ((g1030) & (!g1160) & (g3326) & (!g3327) & (g3377) & (g3400)) + ((g1030) & (!g1160) & (g3326) & (g3327) & (!g3377) & (g3400)) + ((g1030) & (!g1160) & (g3326) & (g3327) & (g3377) & (!g3400)) + ((g1030) & (!g1160) & (g3326) & (g3327) & (g3377) & (g3400)) + ((g1030) & (g1160) & (!g3326) & (!g3327) & (!g3377) & (!g3400)) + ((g1030) & (g1160) & (g3326) & (!g3327) & (!g3377) & (g3400)) + ((g1030) & (g1160) & (g3326) & (!g3327) & (g3377) & (!g3400)) + ((g1030) & (g1160) & (g3326) & (!g3327) & (g3377) & (g3400)) + ((g1030) & (g1160) & (g3326) & (g3327) & (!g3377) & (!g3400)) + ((g1030) & (g1160) & (g3326) & (g3327) & (!g3377) & (g3400)) + ((g1030) & (g1160) & (g3326) & (g3327) & (g3377) & (!g3400)) + ((g1030) & (g1160) & (g3326) & (g3327) & (g3377) & (g3400)));
	assign g3434 = (((!g1160) & (!g3327) & (g3377) & (!g3400)) + ((!g1160) & (g3327) & (!g3377) & (!g3400)) + ((!g1160) & (g3327) & (!g3377) & (g3400)) + ((!g1160) & (g3327) & (g3377) & (g3400)) + ((g1160) & (!g3327) & (!g3377) & (!g3400)) + ((g1160) & (g3327) & (!g3377) & (g3400)) + ((g1160) & (g3327) & (g3377) & (!g3400)) + ((g1160) & (g3327) & (g3377) & (g3400)));
	assign g3435 = (((!g1154) & (!g1295) & (!g3329) & (g3330) & (g3376) & (!g3400)) + ((!g1154) & (!g1295) & (g3329) & (!g3330) & (!g3376) & (!g3400)) + ((!g1154) & (!g1295) & (g3329) & (!g3330) & (!g3376) & (g3400)) + ((!g1154) & (!g1295) & (g3329) & (!g3330) & (g3376) & (!g3400)) + ((!g1154) & (!g1295) & (g3329) & (!g3330) & (g3376) & (g3400)) + ((!g1154) & (!g1295) & (g3329) & (g3330) & (!g3376) & (!g3400)) + ((!g1154) & (!g1295) & (g3329) & (g3330) & (!g3376) & (g3400)) + ((!g1154) & (!g1295) & (g3329) & (g3330) & (g3376) & (g3400)) + ((!g1154) & (g1295) & (!g3329) & (!g3330) & (g3376) & (!g3400)) + ((!g1154) & (g1295) & (!g3329) & (g3330) & (!g3376) & (!g3400)) + ((!g1154) & (g1295) & (!g3329) & (g3330) & (g3376) & (!g3400)) + ((!g1154) & (g1295) & (g3329) & (!g3330) & (!g3376) & (!g3400)) + ((!g1154) & (g1295) & (g3329) & (!g3330) & (!g3376) & (g3400)) + ((!g1154) & (g1295) & (g3329) & (!g3330) & (g3376) & (g3400)) + ((!g1154) & (g1295) & (g3329) & (g3330) & (!g3376) & (g3400)) + ((!g1154) & (g1295) & (g3329) & (g3330) & (g3376) & (g3400)) + ((g1154) & (!g1295) & (!g3329) & (!g3330) & (!g3376) & (!g3400)) + ((g1154) & (!g1295) & (!g3329) & (!g3330) & (g3376) & (!g3400)) + ((g1154) & (!g1295) & (!g3329) & (g3330) & (!g3376) & (!g3400)) + ((g1154) & (!g1295) & (g3329) & (!g3330) & (!g3376) & (g3400)) + ((g1154) & (!g1295) & (g3329) & (!g3330) & (g3376) & (g3400)) + ((g1154) & (!g1295) & (g3329) & (g3330) & (!g3376) & (g3400)) + ((g1154) & (!g1295) & (g3329) & (g3330) & (g3376) & (!g3400)) + ((g1154) & (!g1295) & (g3329) & (g3330) & (g3376) & (g3400)) + ((g1154) & (g1295) & (!g3329) & (!g3330) & (!g3376) & (!g3400)) + ((g1154) & (g1295) & (g3329) & (!g3330) & (!g3376) & (g3400)) + ((g1154) & (g1295) & (g3329) & (!g3330) & (g3376) & (!g3400)) + ((g1154) & (g1295) & (g3329) & (!g3330) & (g3376) & (g3400)) + ((g1154) & (g1295) & (g3329) & (g3330) & (!g3376) & (!g3400)) + ((g1154) & (g1295) & (g3329) & (g3330) & (!g3376) & (g3400)) + ((g1154) & (g1295) & (g3329) & (g3330) & (g3376) & (!g3400)) + ((g1154) & (g1295) & (g3329) & (g3330) & (g3376) & (g3400)));
	assign g3436 = (((!g1295) & (!g3330) & (g3376) & (!g3400)) + ((!g1295) & (g3330) & (!g3376) & (!g3400)) + ((!g1295) & (g3330) & (!g3376) & (g3400)) + ((!g1295) & (g3330) & (g3376) & (g3400)) + ((g1295) & (!g3330) & (!g3376) & (!g3400)) + ((g1295) & (g3330) & (!g3376) & (g3400)) + ((g1295) & (g3330) & (g3376) & (!g3400)) + ((g1295) & (g3330) & (g3376) & (g3400)));
	assign g3437 = (((!g1285) & (!g1437) & (!g3332) & (g3333) & (g3375) & (!g3400)) + ((!g1285) & (!g1437) & (g3332) & (!g3333) & (!g3375) & (!g3400)) + ((!g1285) & (!g1437) & (g3332) & (!g3333) & (!g3375) & (g3400)) + ((!g1285) & (!g1437) & (g3332) & (!g3333) & (g3375) & (!g3400)) + ((!g1285) & (!g1437) & (g3332) & (!g3333) & (g3375) & (g3400)) + ((!g1285) & (!g1437) & (g3332) & (g3333) & (!g3375) & (!g3400)) + ((!g1285) & (!g1437) & (g3332) & (g3333) & (!g3375) & (g3400)) + ((!g1285) & (!g1437) & (g3332) & (g3333) & (g3375) & (g3400)) + ((!g1285) & (g1437) & (!g3332) & (!g3333) & (g3375) & (!g3400)) + ((!g1285) & (g1437) & (!g3332) & (g3333) & (!g3375) & (!g3400)) + ((!g1285) & (g1437) & (!g3332) & (g3333) & (g3375) & (!g3400)) + ((!g1285) & (g1437) & (g3332) & (!g3333) & (!g3375) & (!g3400)) + ((!g1285) & (g1437) & (g3332) & (!g3333) & (!g3375) & (g3400)) + ((!g1285) & (g1437) & (g3332) & (!g3333) & (g3375) & (g3400)) + ((!g1285) & (g1437) & (g3332) & (g3333) & (!g3375) & (g3400)) + ((!g1285) & (g1437) & (g3332) & (g3333) & (g3375) & (g3400)) + ((g1285) & (!g1437) & (!g3332) & (!g3333) & (!g3375) & (!g3400)) + ((g1285) & (!g1437) & (!g3332) & (!g3333) & (g3375) & (!g3400)) + ((g1285) & (!g1437) & (!g3332) & (g3333) & (!g3375) & (!g3400)) + ((g1285) & (!g1437) & (g3332) & (!g3333) & (!g3375) & (g3400)) + ((g1285) & (!g1437) & (g3332) & (!g3333) & (g3375) & (g3400)) + ((g1285) & (!g1437) & (g3332) & (g3333) & (!g3375) & (g3400)) + ((g1285) & (!g1437) & (g3332) & (g3333) & (g3375) & (!g3400)) + ((g1285) & (!g1437) & (g3332) & (g3333) & (g3375) & (g3400)) + ((g1285) & (g1437) & (!g3332) & (!g3333) & (!g3375) & (!g3400)) + ((g1285) & (g1437) & (g3332) & (!g3333) & (!g3375) & (g3400)) + ((g1285) & (g1437) & (g3332) & (!g3333) & (g3375) & (!g3400)) + ((g1285) & (g1437) & (g3332) & (!g3333) & (g3375) & (g3400)) + ((g1285) & (g1437) & (g3332) & (g3333) & (!g3375) & (!g3400)) + ((g1285) & (g1437) & (g3332) & (g3333) & (!g3375) & (g3400)) + ((g1285) & (g1437) & (g3332) & (g3333) & (g3375) & (!g3400)) + ((g1285) & (g1437) & (g3332) & (g3333) & (g3375) & (g3400)));
	assign g3438 = (((!g1437) & (!g3333) & (g3375) & (!g3400)) + ((!g1437) & (g3333) & (!g3375) & (!g3400)) + ((!g1437) & (g3333) & (!g3375) & (g3400)) + ((!g1437) & (g3333) & (g3375) & (g3400)) + ((g1437) & (!g3333) & (!g3375) & (!g3400)) + ((g1437) & (g3333) & (!g3375) & (g3400)) + ((g1437) & (g3333) & (g3375) & (!g3400)) + ((g1437) & (g3333) & (g3375) & (g3400)));
	assign g3439 = (((!g1423) & (!g1586) & (!g3335) & (g3336) & (g3374) & (!g3400)) + ((!g1423) & (!g1586) & (g3335) & (!g3336) & (!g3374) & (!g3400)) + ((!g1423) & (!g1586) & (g3335) & (!g3336) & (!g3374) & (g3400)) + ((!g1423) & (!g1586) & (g3335) & (!g3336) & (g3374) & (!g3400)) + ((!g1423) & (!g1586) & (g3335) & (!g3336) & (g3374) & (g3400)) + ((!g1423) & (!g1586) & (g3335) & (g3336) & (!g3374) & (!g3400)) + ((!g1423) & (!g1586) & (g3335) & (g3336) & (!g3374) & (g3400)) + ((!g1423) & (!g1586) & (g3335) & (g3336) & (g3374) & (g3400)) + ((!g1423) & (g1586) & (!g3335) & (!g3336) & (g3374) & (!g3400)) + ((!g1423) & (g1586) & (!g3335) & (g3336) & (!g3374) & (!g3400)) + ((!g1423) & (g1586) & (!g3335) & (g3336) & (g3374) & (!g3400)) + ((!g1423) & (g1586) & (g3335) & (!g3336) & (!g3374) & (!g3400)) + ((!g1423) & (g1586) & (g3335) & (!g3336) & (!g3374) & (g3400)) + ((!g1423) & (g1586) & (g3335) & (!g3336) & (g3374) & (g3400)) + ((!g1423) & (g1586) & (g3335) & (g3336) & (!g3374) & (g3400)) + ((!g1423) & (g1586) & (g3335) & (g3336) & (g3374) & (g3400)) + ((g1423) & (!g1586) & (!g3335) & (!g3336) & (!g3374) & (!g3400)) + ((g1423) & (!g1586) & (!g3335) & (!g3336) & (g3374) & (!g3400)) + ((g1423) & (!g1586) & (!g3335) & (g3336) & (!g3374) & (!g3400)) + ((g1423) & (!g1586) & (g3335) & (!g3336) & (!g3374) & (g3400)) + ((g1423) & (!g1586) & (g3335) & (!g3336) & (g3374) & (g3400)) + ((g1423) & (!g1586) & (g3335) & (g3336) & (!g3374) & (g3400)) + ((g1423) & (!g1586) & (g3335) & (g3336) & (g3374) & (!g3400)) + ((g1423) & (!g1586) & (g3335) & (g3336) & (g3374) & (g3400)) + ((g1423) & (g1586) & (!g3335) & (!g3336) & (!g3374) & (!g3400)) + ((g1423) & (g1586) & (g3335) & (!g3336) & (!g3374) & (g3400)) + ((g1423) & (g1586) & (g3335) & (!g3336) & (g3374) & (!g3400)) + ((g1423) & (g1586) & (g3335) & (!g3336) & (g3374) & (g3400)) + ((g1423) & (g1586) & (g3335) & (g3336) & (!g3374) & (!g3400)) + ((g1423) & (g1586) & (g3335) & (g3336) & (!g3374) & (g3400)) + ((g1423) & (g1586) & (g3335) & (g3336) & (g3374) & (!g3400)) + ((g1423) & (g1586) & (g3335) & (g3336) & (g3374) & (g3400)));
	assign g3440 = (((!g1586) & (!g3336) & (g3374) & (!g3400)) + ((!g1586) & (g3336) & (!g3374) & (!g3400)) + ((!g1586) & (g3336) & (!g3374) & (g3400)) + ((!g1586) & (g3336) & (g3374) & (g3400)) + ((g1586) & (!g3336) & (!g3374) & (!g3400)) + ((g1586) & (g3336) & (!g3374) & (g3400)) + ((g1586) & (g3336) & (g3374) & (!g3400)) + ((g1586) & (g3336) & (g3374) & (g3400)));
	assign g3441 = (((!g1568) & (!g1742) & (!g3338) & (g3339) & (g3373) & (!g3400)) + ((!g1568) & (!g1742) & (g3338) & (!g3339) & (!g3373) & (!g3400)) + ((!g1568) & (!g1742) & (g3338) & (!g3339) & (!g3373) & (g3400)) + ((!g1568) & (!g1742) & (g3338) & (!g3339) & (g3373) & (!g3400)) + ((!g1568) & (!g1742) & (g3338) & (!g3339) & (g3373) & (g3400)) + ((!g1568) & (!g1742) & (g3338) & (g3339) & (!g3373) & (!g3400)) + ((!g1568) & (!g1742) & (g3338) & (g3339) & (!g3373) & (g3400)) + ((!g1568) & (!g1742) & (g3338) & (g3339) & (g3373) & (g3400)) + ((!g1568) & (g1742) & (!g3338) & (!g3339) & (g3373) & (!g3400)) + ((!g1568) & (g1742) & (!g3338) & (g3339) & (!g3373) & (!g3400)) + ((!g1568) & (g1742) & (!g3338) & (g3339) & (g3373) & (!g3400)) + ((!g1568) & (g1742) & (g3338) & (!g3339) & (!g3373) & (!g3400)) + ((!g1568) & (g1742) & (g3338) & (!g3339) & (!g3373) & (g3400)) + ((!g1568) & (g1742) & (g3338) & (!g3339) & (g3373) & (g3400)) + ((!g1568) & (g1742) & (g3338) & (g3339) & (!g3373) & (g3400)) + ((!g1568) & (g1742) & (g3338) & (g3339) & (g3373) & (g3400)) + ((g1568) & (!g1742) & (!g3338) & (!g3339) & (!g3373) & (!g3400)) + ((g1568) & (!g1742) & (!g3338) & (!g3339) & (g3373) & (!g3400)) + ((g1568) & (!g1742) & (!g3338) & (g3339) & (!g3373) & (!g3400)) + ((g1568) & (!g1742) & (g3338) & (!g3339) & (!g3373) & (g3400)) + ((g1568) & (!g1742) & (g3338) & (!g3339) & (g3373) & (g3400)) + ((g1568) & (!g1742) & (g3338) & (g3339) & (!g3373) & (g3400)) + ((g1568) & (!g1742) & (g3338) & (g3339) & (g3373) & (!g3400)) + ((g1568) & (!g1742) & (g3338) & (g3339) & (g3373) & (g3400)) + ((g1568) & (g1742) & (!g3338) & (!g3339) & (!g3373) & (!g3400)) + ((g1568) & (g1742) & (g3338) & (!g3339) & (!g3373) & (g3400)) + ((g1568) & (g1742) & (g3338) & (!g3339) & (g3373) & (!g3400)) + ((g1568) & (g1742) & (g3338) & (!g3339) & (g3373) & (g3400)) + ((g1568) & (g1742) & (g3338) & (g3339) & (!g3373) & (!g3400)) + ((g1568) & (g1742) & (g3338) & (g3339) & (!g3373) & (g3400)) + ((g1568) & (g1742) & (g3338) & (g3339) & (g3373) & (!g3400)) + ((g1568) & (g1742) & (g3338) & (g3339) & (g3373) & (g3400)));
	assign g3442 = (((!g1742) & (!g3339) & (g3373) & (!g3400)) + ((!g1742) & (g3339) & (!g3373) & (!g3400)) + ((!g1742) & (g3339) & (!g3373) & (g3400)) + ((!g1742) & (g3339) & (g3373) & (g3400)) + ((g1742) & (!g3339) & (!g3373) & (!g3400)) + ((g1742) & (g3339) & (!g3373) & (g3400)) + ((g1742) & (g3339) & (g3373) & (!g3400)) + ((g1742) & (g3339) & (g3373) & (g3400)));
	assign g3443 = (((!g1720) & (!g1905) & (!g3341) & (g3342) & (g3372) & (!g3400)) + ((!g1720) & (!g1905) & (g3341) & (!g3342) & (!g3372) & (!g3400)) + ((!g1720) & (!g1905) & (g3341) & (!g3342) & (!g3372) & (g3400)) + ((!g1720) & (!g1905) & (g3341) & (!g3342) & (g3372) & (!g3400)) + ((!g1720) & (!g1905) & (g3341) & (!g3342) & (g3372) & (g3400)) + ((!g1720) & (!g1905) & (g3341) & (g3342) & (!g3372) & (!g3400)) + ((!g1720) & (!g1905) & (g3341) & (g3342) & (!g3372) & (g3400)) + ((!g1720) & (!g1905) & (g3341) & (g3342) & (g3372) & (g3400)) + ((!g1720) & (g1905) & (!g3341) & (!g3342) & (g3372) & (!g3400)) + ((!g1720) & (g1905) & (!g3341) & (g3342) & (!g3372) & (!g3400)) + ((!g1720) & (g1905) & (!g3341) & (g3342) & (g3372) & (!g3400)) + ((!g1720) & (g1905) & (g3341) & (!g3342) & (!g3372) & (!g3400)) + ((!g1720) & (g1905) & (g3341) & (!g3342) & (!g3372) & (g3400)) + ((!g1720) & (g1905) & (g3341) & (!g3342) & (g3372) & (g3400)) + ((!g1720) & (g1905) & (g3341) & (g3342) & (!g3372) & (g3400)) + ((!g1720) & (g1905) & (g3341) & (g3342) & (g3372) & (g3400)) + ((g1720) & (!g1905) & (!g3341) & (!g3342) & (!g3372) & (!g3400)) + ((g1720) & (!g1905) & (!g3341) & (!g3342) & (g3372) & (!g3400)) + ((g1720) & (!g1905) & (!g3341) & (g3342) & (!g3372) & (!g3400)) + ((g1720) & (!g1905) & (g3341) & (!g3342) & (!g3372) & (g3400)) + ((g1720) & (!g1905) & (g3341) & (!g3342) & (g3372) & (g3400)) + ((g1720) & (!g1905) & (g3341) & (g3342) & (!g3372) & (g3400)) + ((g1720) & (!g1905) & (g3341) & (g3342) & (g3372) & (!g3400)) + ((g1720) & (!g1905) & (g3341) & (g3342) & (g3372) & (g3400)) + ((g1720) & (g1905) & (!g3341) & (!g3342) & (!g3372) & (!g3400)) + ((g1720) & (g1905) & (g3341) & (!g3342) & (!g3372) & (g3400)) + ((g1720) & (g1905) & (g3341) & (!g3342) & (g3372) & (!g3400)) + ((g1720) & (g1905) & (g3341) & (!g3342) & (g3372) & (g3400)) + ((g1720) & (g1905) & (g3341) & (g3342) & (!g3372) & (!g3400)) + ((g1720) & (g1905) & (g3341) & (g3342) & (!g3372) & (g3400)) + ((g1720) & (g1905) & (g3341) & (g3342) & (g3372) & (!g3400)) + ((g1720) & (g1905) & (g3341) & (g3342) & (g3372) & (g3400)));
	assign g3444 = (((!g1905) & (!g3342) & (g3372) & (!g3400)) + ((!g1905) & (g3342) & (!g3372) & (!g3400)) + ((!g1905) & (g3342) & (!g3372) & (g3400)) + ((!g1905) & (g3342) & (g3372) & (g3400)) + ((g1905) & (!g3342) & (!g3372) & (!g3400)) + ((g1905) & (g3342) & (!g3372) & (g3400)) + ((g1905) & (g3342) & (g3372) & (!g3400)) + ((g1905) & (g3342) & (g3372) & (g3400)));
	assign g3445 = (((!g1879) & (!g2075) & (!g3344) & (g3345) & (g3371) & (!g3400)) + ((!g1879) & (!g2075) & (g3344) & (!g3345) & (!g3371) & (!g3400)) + ((!g1879) & (!g2075) & (g3344) & (!g3345) & (!g3371) & (g3400)) + ((!g1879) & (!g2075) & (g3344) & (!g3345) & (g3371) & (!g3400)) + ((!g1879) & (!g2075) & (g3344) & (!g3345) & (g3371) & (g3400)) + ((!g1879) & (!g2075) & (g3344) & (g3345) & (!g3371) & (!g3400)) + ((!g1879) & (!g2075) & (g3344) & (g3345) & (!g3371) & (g3400)) + ((!g1879) & (!g2075) & (g3344) & (g3345) & (g3371) & (g3400)) + ((!g1879) & (g2075) & (!g3344) & (!g3345) & (g3371) & (!g3400)) + ((!g1879) & (g2075) & (!g3344) & (g3345) & (!g3371) & (!g3400)) + ((!g1879) & (g2075) & (!g3344) & (g3345) & (g3371) & (!g3400)) + ((!g1879) & (g2075) & (g3344) & (!g3345) & (!g3371) & (!g3400)) + ((!g1879) & (g2075) & (g3344) & (!g3345) & (!g3371) & (g3400)) + ((!g1879) & (g2075) & (g3344) & (!g3345) & (g3371) & (g3400)) + ((!g1879) & (g2075) & (g3344) & (g3345) & (!g3371) & (g3400)) + ((!g1879) & (g2075) & (g3344) & (g3345) & (g3371) & (g3400)) + ((g1879) & (!g2075) & (!g3344) & (!g3345) & (!g3371) & (!g3400)) + ((g1879) & (!g2075) & (!g3344) & (!g3345) & (g3371) & (!g3400)) + ((g1879) & (!g2075) & (!g3344) & (g3345) & (!g3371) & (!g3400)) + ((g1879) & (!g2075) & (g3344) & (!g3345) & (!g3371) & (g3400)) + ((g1879) & (!g2075) & (g3344) & (!g3345) & (g3371) & (g3400)) + ((g1879) & (!g2075) & (g3344) & (g3345) & (!g3371) & (g3400)) + ((g1879) & (!g2075) & (g3344) & (g3345) & (g3371) & (!g3400)) + ((g1879) & (!g2075) & (g3344) & (g3345) & (g3371) & (g3400)) + ((g1879) & (g2075) & (!g3344) & (!g3345) & (!g3371) & (!g3400)) + ((g1879) & (g2075) & (g3344) & (!g3345) & (!g3371) & (g3400)) + ((g1879) & (g2075) & (g3344) & (!g3345) & (g3371) & (!g3400)) + ((g1879) & (g2075) & (g3344) & (!g3345) & (g3371) & (g3400)) + ((g1879) & (g2075) & (g3344) & (g3345) & (!g3371) & (!g3400)) + ((g1879) & (g2075) & (g3344) & (g3345) & (!g3371) & (g3400)) + ((g1879) & (g2075) & (g3344) & (g3345) & (g3371) & (!g3400)) + ((g1879) & (g2075) & (g3344) & (g3345) & (g3371) & (g3400)));
	assign g3446 = (((!g2075) & (!g3345) & (g3371) & (!g3400)) + ((!g2075) & (g3345) & (!g3371) & (!g3400)) + ((!g2075) & (g3345) & (!g3371) & (g3400)) + ((!g2075) & (g3345) & (g3371) & (g3400)) + ((g2075) & (!g3345) & (!g3371) & (!g3400)) + ((g2075) & (g3345) & (!g3371) & (g3400)) + ((g2075) & (g3345) & (g3371) & (!g3400)) + ((g2075) & (g3345) & (g3371) & (g3400)));
	assign g3447 = (((!g2045) & (!g2252) & (!g3347) & (g3348) & (g3370) & (!g3400)) + ((!g2045) & (!g2252) & (g3347) & (!g3348) & (!g3370) & (!g3400)) + ((!g2045) & (!g2252) & (g3347) & (!g3348) & (!g3370) & (g3400)) + ((!g2045) & (!g2252) & (g3347) & (!g3348) & (g3370) & (!g3400)) + ((!g2045) & (!g2252) & (g3347) & (!g3348) & (g3370) & (g3400)) + ((!g2045) & (!g2252) & (g3347) & (g3348) & (!g3370) & (!g3400)) + ((!g2045) & (!g2252) & (g3347) & (g3348) & (!g3370) & (g3400)) + ((!g2045) & (!g2252) & (g3347) & (g3348) & (g3370) & (g3400)) + ((!g2045) & (g2252) & (!g3347) & (!g3348) & (g3370) & (!g3400)) + ((!g2045) & (g2252) & (!g3347) & (g3348) & (!g3370) & (!g3400)) + ((!g2045) & (g2252) & (!g3347) & (g3348) & (g3370) & (!g3400)) + ((!g2045) & (g2252) & (g3347) & (!g3348) & (!g3370) & (!g3400)) + ((!g2045) & (g2252) & (g3347) & (!g3348) & (!g3370) & (g3400)) + ((!g2045) & (g2252) & (g3347) & (!g3348) & (g3370) & (g3400)) + ((!g2045) & (g2252) & (g3347) & (g3348) & (!g3370) & (g3400)) + ((!g2045) & (g2252) & (g3347) & (g3348) & (g3370) & (g3400)) + ((g2045) & (!g2252) & (!g3347) & (!g3348) & (!g3370) & (!g3400)) + ((g2045) & (!g2252) & (!g3347) & (!g3348) & (g3370) & (!g3400)) + ((g2045) & (!g2252) & (!g3347) & (g3348) & (!g3370) & (!g3400)) + ((g2045) & (!g2252) & (g3347) & (!g3348) & (!g3370) & (g3400)) + ((g2045) & (!g2252) & (g3347) & (!g3348) & (g3370) & (g3400)) + ((g2045) & (!g2252) & (g3347) & (g3348) & (!g3370) & (g3400)) + ((g2045) & (!g2252) & (g3347) & (g3348) & (g3370) & (!g3400)) + ((g2045) & (!g2252) & (g3347) & (g3348) & (g3370) & (g3400)) + ((g2045) & (g2252) & (!g3347) & (!g3348) & (!g3370) & (!g3400)) + ((g2045) & (g2252) & (g3347) & (!g3348) & (!g3370) & (g3400)) + ((g2045) & (g2252) & (g3347) & (!g3348) & (g3370) & (!g3400)) + ((g2045) & (g2252) & (g3347) & (!g3348) & (g3370) & (g3400)) + ((g2045) & (g2252) & (g3347) & (g3348) & (!g3370) & (!g3400)) + ((g2045) & (g2252) & (g3347) & (g3348) & (!g3370) & (g3400)) + ((g2045) & (g2252) & (g3347) & (g3348) & (g3370) & (!g3400)) + ((g2045) & (g2252) & (g3347) & (g3348) & (g3370) & (g3400)));
	assign g3448 = (((!g2252) & (!g3348) & (g3370) & (!g3400)) + ((!g2252) & (g3348) & (!g3370) & (!g3400)) + ((!g2252) & (g3348) & (!g3370) & (g3400)) + ((!g2252) & (g3348) & (g3370) & (g3400)) + ((g2252) & (!g3348) & (!g3370) & (!g3400)) + ((g2252) & (g3348) & (!g3370) & (g3400)) + ((g2252) & (g3348) & (g3370) & (!g3400)) + ((g2252) & (g3348) & (g3370) & (g3400)));
	assign g3449 = (((!g2218) & (!g2436) & (!g3350) & (g3351) & (g3369) & (!g3400)) + ((!g2218) & (!g2436) & (g3350) & (!g3351) & (!g3369) & (!g3400)) + ((!g2218) & (!g2436) & (g3350) & (!g3351) & (!g3369) & (g3400)) + ((!g2218) & (!g2436) & (g3350) & (!g3351) & (g3369) & (!g3400)) + ((!g2218) & (!g2436) & (g3350) & (!g3351) & (g3369) & (g3400)) + ((!g2218) & (!g2436) & (g3350) & (g3351) & (!g3369) & (!g3400)) + ((!g2218) & (!g2436) & (g3350) & (g3351) & (!g3369) & (g3400)) + ((!g2218) & (!g2436) & (g3350) & (g3351) & (g3369) & (g3400)) + ((!g2218) & (g2436) & (!g3350) & (!g3351) & (g3369) & (!g3400)) + ((!g2218) & (g2436) & (!g3350) & (g3351) & (!g3369) & (!g3400)) + ((!g2218) & (g2436) & (!g3350) & (g3351) & (g3369) & (!g3400)) + ((!g2218) & (g2436) & (g3350) & (!g3351) & (!g3369) & (!g3400)) + ((!g2218) & (g2436) & (g3350) & (!g3351) & (!g3369) & (g3400)) + ((!g2218) & (g2436) & (g3350) & (!g3351) & (g3369) & (g3400)) + ((!g2218) & (g2436) & (g3350) & (g3351) & (!g3369) & (g3400)) + ((!g2218) & (g2436) & (g3350) & (g3351) & (g3369) & (g3400)) + ((g2218) & (!g2436) & (!g3350) & (!g3351) & (!g3369) & (!g3400)) + ((g2218) & (!g2436) & (!g3350) & (!g3351) & (g3369) & (!g3400)) + ((g2218) & (!g2436) & (!g3350) & (g3351) & (!g3369) & (!g3400)) + ((g2218) & (!g2436) & (g3350) & (!g3351) & (!g3369) & (g3400)) + ((g2218) & (!g2436) & (g3350) & (!g3351) & (g3369) & (g3400)) + ((g2218) & (!g2436) & (g3350) & (g3351) & (!g3369) & (g3400)) + ((g2218) & (!g2436) & (g3350) & (g3351) & (g3369) & (!g3400)) + ((g2218) & (!g2436) & (g3350) & (g3351) & (g3369) & (g3400)) + ((g2218) & (g2436) & (!g3350) & (!g3351) & (!g3369) & (!g3400)) + ((g2218) & (g2436) & (g3350) & (!g3351) & (!g3369) & (g3400)) + ((g2218) & (g2436) & (g3350) & (!g3351) & (g3369) & (!g3400)) + ((g2218) & (g2436) & (g3350) & (!g3351) & (g3369) & (g3400)) + ((g2218) & (g2436) & (g3350) & (g3351) & (!g3369) & (!g3400)) + ((g2218) & (g2436) & (g3350) & (g3351) & (!g3369) & (g3400)) + ((g2218) & (g2436) & (g3350) & (g3351) & (g3369) & (!g3400)) + ((g2218) & (g2436) & (g3350) & (g3351) & (g3369) & (g3400)));
	assign g3450 = (((!g2436) & (!g3351) & (g3369) & (!g3400)) + ((!g2436) & (g3351) & (!g3369) & (!g3400)) + ((!g2436) & (g3351) & (!g3369) & (g3400)) + ((!g2436) & (g3351) & (g3369) & (g3400)) + ((g2436) & (!g3351) & (!g3369) & (!g3400)) + ((g2436) & (g3351) & (!g3369) & (g3400)) + ((g2436) & (g3351) & (g3369) & (!g3400)) + ((g2436) & (g3351) & (g3369) & (g3400)));
	assign g3451 = (((!g2398) & (!g2627) & (!g3353) & (g3354) & (g3368) & (!g3400)) + ((!g2398) & (!g2627) & (g3353) & (!g3354) & (!g3368) & (!g3400)) + ((!g2398) & (!g2627) & (g3353) & (!g3354) & (!g3368) & (g3400)) + ((!g2398) & (!g2627) & (g3353) & (!g3354) & (g3368) & (!g3400)) + ((!g2398) & (!g2627) & (g3353) & (!g3354) & (g3368) & (g3400)) + ((!g2398) & (!g2627) & (g3353) & (g3354) & (!g3368) & (!g3400)) + ((!g2398) & (!g2627) & (g3353) & (g3354) & (!g3368) & (g3400)) + ((!g2398) & (!g2627) & (g3353) & (g3354) & (g3368) & (g3400)) + ((!g2398) & (g2627) & (!g3353) & (!g3354) & (g3368) & (!g3400)) + ((!g2398) & (g2627) & (!g3353) & (g3354) & (!g3368) & (!g3400)) + ((!g2398) & (g2627) & (!g3353) & (g3354) & (g3368) & (!g3400)) + ((!g2398) & (g2627) & (g3353) & (!g3354) & (!g3368) & (!g3400)) + ((!g2398) & (g2627) & (g3353) & (!g3354) & (!g3368) & (g3400)) + ((!g2398) & (g2627) & (g3353) & (!g3354) & (g3368) & (g3400)) + ((!g2398) & (g2627) & (g3353) & (g3354) & (!g3368) & (g3400)) + ((!g2398) & (g2627) & (g3353) & (g3354) & (g3368) & (g3400)) + ((g2398) & (!g2627) & (!g3353) & (!g3354) & (!g3368) & (!g3400)) + ((g2398) & (!g2627) & (!g3353) & (!g3354) & (g3368) & (!g3400)) + ((g2398) & (!g2627) & (!g3353) & (g3354) & (!g3368) & (!g3400)) + ((g2398) & (!g2627) & (g3353) & (!g3354) & (!g3368) & (g3400)) + ((g2398) & (!g2627) & (g3353) & (!g3354) & (g3368) & (g3400)) + ((g2398) & (!g2627) & (g3353) & (g3354) & (!g3368) & (g3400)) + ((g2398) & (!g2627) & (g3353) & (g3354) & (g3368) & (!g3400)) + ((g2398) & (!g2627) & (g3353) & (g3354) & (g3368) & (g3400)) + ((g2398) & (g2627) & (!g3353) & (!g3354) & (!g3368) & (!g3400)) + ((g2398) & (g2627) & (g3353) & (!g3354) & (!g3368) & (g3400)) + ((g2398) & (g2627) & (g3353) & (!g3354) & (g3368) & (!g3400)) + ((g2398) & (g2627) & (g3353) & (!g3354) & (g3368) & (g3400)) + ((g2398) & (g2627) & (g3353) & (g3354) & (!g3368) & (!g3400)) + ((g2398) & (g2627) & (g3353) & (g3354) & (!g3368) & (g3400)) + ((g2398) & (g2627) & (g3353) & (g3354) & (g3368) & (!g3400)) + ((g2398) & (g2627) & (g3353) & (g3354) & (g3368) & (g3400)));
	assign g3452 = (((!g2627) & (!g3354) & (g3368) & (!g3400)) + ((!g2627) & (g3354) & (!g3368) & (!g3400)) + ((!g2627) & (g3354) & (!g3368) & (g3400)) + ((!g2627) & (g3354) & (g3368) & (g3400)) + ((g2627) & (!g3354) & (!g3368) & (!g3400)) + ((g2627) & (g3354) & (!g3368) & (g3400)) + ((g2627) & (g3354) & (g3368) & (!g3400)) + ((g2627) & (g3354) & (g3368) & (g3400)));
	assign g3453 = (((!g2585) & (!g2825) & (!g3356) & (g3357) & (g3367) & (!g3400)) + ((!g2585) & (!g2825) & (g3356) & (!g3357) & (!g3367) & (!g3400)) + ((!g2585) & (!g2825) & (g3356) & (!g3357) & (!g3367) & (g3400)) + ((!g2585) & (!g2825) & (g3356) & (!g3357) & (g3367) & (!g3400)) + ((!g2585) & (!g2825) & (g3356) & (!g3357) & (g3367) & (g3400)) + ((!g2585) & (!g2825) & (g3356) & (g3357) & (!g3367) & (!g3400)) + ((!g2585) & (!g2825) & (g3356) & (g3357) & (!g3367) & (g3400)) + ((!g2585) & (!g2825) & (g3356) & (g3357) & (g3367) & (g3400)) + ((!g2585) & (g2825) & (!g3356) & (!g3357) & (g3367) & (!g3400)) + ((!g2585) & (g2825) & (!g3356) & (g3357) & (!g3367) & (!g3400)) + ((!g2585) & (g2825) & (!g3356) & (g3357) & (g3367) & (!g3400)) + ((!g2585) & (g2825) & (g3356) & (!g3357) & (!g3367) & (!g3400)) + ((!g2585) & (g2825) & (g3356) & (!g3357) & (!g3367) & (g3400)) + ((!g2585) & (g2825) & (g3356) & (!g3357) & (g3367) & (g3400)) + ((!g2585) & (g2825) & (g3356) & (g3357) & (!g3367) & (g3400)) + ((!g2585) & (g2825) & (g3356) & (g3357) & (g3367) & (g3400)) + ((g2585) & (!g2825) & (!g3356) & (!g3357) & (!g3367) & (!g3400)) + ((g2585) & (!g2825) & (!g3356) & (!g3357) & (g3367) & (!g3400)) + ((g2585) & (!g2825) & (!g3356) & (g3357) & (!g3367) & (!g3400)) + ((g2585) & (!g2825) & (g3356) & (!g3357) & (!g3367) & (g3400)) + ((g2585) & (!g2825) & (g3356) & (!g3357) & (g3367) & (g3400)) + ((g2585) & (!g2825) & (g3356) & (g3357) & (!g3367) & (g3400)) + ((g2585) & (!g2825) & (g3356) & (g3357) & (g3367) & (!g3400)) + ((g2585) & (!g2825) & (g3356) & (g3357) & (g3367) & (g3400)) + ((g2585) & (g2825) & (!g3356) & (!g3357) & (!g3367) & (!g3400)) + ((g2585) & (g2825) & (g3356) & (!g3357) & (!g3367) & (g3400)) + ((g2585) & (g2825) & (g3356) & (!g3357) & (g3367) & (!g3400)) + ((g2585) & (g2825) & (g3356) & (!g3357) & (g3367) & (g3400)) + ((g2585) & (g2825) & (g3356) & (g3357) & (!g3367) & (!g3400)) + ((g2585) & (g2825) & (g3356) & (g3357) & (!g3367) & (g3400)) + ((g2585) & (g2825) & (g3356) & (g3357) & (g3367) & (!g3400)) + ((g2585) & (g2825) & (g3356) & (g3357) & (g3367) & (g3400)));
	assign g3454 = (((!g2825) & (!g3357) & (g3367) & (!g3400)) + ((!g2825) & (g3357) & (!g3367) & (!g3400)) + ((!g2825) & (g3357) & (!g3367) & (g3400)) + ((!g2825) & (g3357) & (g3367) & (g3400)) + ((g2825) & (!g3357) & (!g3367) & (!g3400)) + ((g2825) & (g3357) & (!g3367) & (g3400)) + ((g2825) & (g3357) & (g3367) & (!g3400)) + ((g2825) & (g3357) & (g3367) & (g3400)));
	assign g3455 = (((!g2779) & (!g3030) & (!g3359) & (g3360) & (g3366) & (!g3400)) + ((!g2779) & (!g3030) & (g3359) & (!g3360) & (!g3366) & (!g3400)) + ((!g2779) & (!g3030) & (g3359) & (!g3360) & (!g3366) & (g3400)) + ((!g2779) & (!g3030) & (g3359) & (!g3360) & (g3366) & (!g3400)) + ((!g2779) & (!g3030) & (g3359) & (!g3360) & (g3366) & (g3400)) + ((!g2779) & (!g3030) & (g3359) & (g3360) & (!g3366) & (!g3400)) + ((!g2779) & (!g3030) & (g3359) & (g3360) & (!g3366) & (g3400)) + ((!g2779) & (!g3030) & (g3359) & (g3360) & (g3366) & (g3400)) + ((!g2779) & (g3030) & (!g3359) & (!g3360) & (g3366) & (!g3400)) + ((!g2779) & (g3030) & (!g3359) & (g3360) & (!g3366) & (!g3400)) + ((!g2779) & (g3030) & (!g3359) & (g3360) & (g3366) & (!g3400)) + ((!g2779) & (g3030) & (g3359) & (!g3360) & (!g3366) & (!g3400)) + ((!g2779) & (g3030) & (g3359) & (!g3360) & (!g3366) & (g3400)) + ((!g2779) & (g3030) & (g3359) & (!g3360) & (g3366) & (g3400)) + ((!g2779) & (g3030) & (g3359) & (g3360) & (!g3366) & (g3400)) + ((!g2779) & (g3030) & (g3359) & (g3360) & (g3366) & (g3400)) + ((g2779) & (!g3030) & (!g3359) & (!g3360) & (!g3366) & (!g3400)) + ((g2779) & (!g3030) & (!g3359) & (!g3360) & (g3366) & (!g3400)) + ((g2779) & (!g3030) & (!g3359) & (g3360) & (!g3366) & (!g3400)) + ((g2779) & (!g3030) & (g3359) & (!g3360) & (!g3366) & (g3400)) + ((g2779) & (!g3030) & (g3359) & (!g3360) & (g3366) & (g3400)) + ((g2779) & (!g3030) & (g3359) & (g3360) & (!g3366) & (g3400)) + ((g2779) & (!g3030) & (g3359) & (g3360) & (g3366) & (!g3400)) + ((g2779) & (!g3030) & (g3359) & (g3360) & (g3366) & (g3400)) + ((g2779) & (g3030) & (!g3359) & (!g3360) & (!g3366) & (!g3400)) + ((g2779) & (g3030) & (g3359) & (!g3360) & (!g3366) & (g3400)) + ((g2779) & (g3030) & (g3359) & (!g3360) & (g3366) & (!g3400)) + ((g2779) & (g3030) & (g3359) & (!g3360) & (g3366) & (g3400)) + ((g2779) & (g3030) & (g3359) & (g3360) & (!g3366) & (!g3400)) + ((g2779) & (g3030) & (g3359) & (g3360) & (!g3366) & (g3400)) + ((g2779) & (g3030) & (g3359) & (g3360) & (g3366) & (!g3400)) + ((g2779) & (g3030) & (g3359) & (g3360) & (g3366) & (g3400)));
	assign g3456 = (((!g3030) & (!g3360) & (g3366) & (!g3400)) + ((!g3030) & (g3360) & (!g3366) & (!g3400)) + ((!g3030) & (g3360) & (!g3366) & (g3400)) + ((!g3030) & (g3360) & (g3366) & (g3400)) + ((g3030) & (!g3360) & (!g3366) & (!g3400)) + ((g3030) & (g3360) & (!g3366) & (g3400)) + ((g3030) & (g3360) & (g3366) & (!g3400)) + ((g3030) & (g3360) & (g3366) & (g3400)));
	assign g3457 = (((!g2980) & (!g3178) & (!g3362) & (g3363) & (g3365) & (!g3400)) + ((!g2980) & (!g3178) & (g3362) & (!g3363) & (!g3365) & (!g3400)) + ((!g2980) & (!g3178) & (g3362) & (!g3363) & (!g3365) & (g3400)) + ((!g2980) & (!g3178) & (g3362) & (!g3363) & (g3365) & (!g3400)) + ((!g2980) & (!g3178) & (g3362) & (!g3363) & (g3365) & (g3400)) + ((!g2980) & (!g3178) & (g3362) & (g3363) & (!g3365) & (!g3400)) + ((!g2980) & (!g3178) & (g3362) & (g3363) & (!g3365) & (g3400)) + ((!g2980) & (!g3178) & (g3362) & (g3363) & (g3365) & (g3400)) + ((!g2980) & (g3178) & (!g3362) & (!g3363) & (g3365) & (!g3400)) + ((!g2980) & (g3178) & (!g3362) & (g3363) & (!g3365) & (!g3400)) + ((!g2980) & (g3178) & (!g3362) & (g3363) & (g3365) & (!g3400)) + ((!g2980) & (g3178) & (g3362) & (!g3363) & (!g3365) & (!g3400)) + ((!g2980) & (g3178) & (g3362) & (!g3363) & (!g3365) & (g3400)) + ((!g2980) & (g3178) & (g3362) & (!g3363) & (g3365) & (g3400)) + ((!g2980) & (g3178) & (g3362) & (g3363) & (!g3365) & (g3400)) + ((!g2980) & (g3178) & (g3362) & (g3363) & (g3365) & (g3400)) + ((g2980) & (!g3178) & (!g3362) & (!g3363) & (!g3365) & (!g3400)) + ((g2980) & (!g3178) & (!g3362) & (!g3363) & (g3365) & (!g3400)) + ((g2980) & (!g3178) & (!g3362) & (g3363) & (!g3365) & (!g3400)) + ((g2980) & (!g3178) & (g3362) & (!g3363) & (!g3365) & (g3400)) + ((g2980) & (!g3178) & (g3362) & (!g3363) & (g3365) & (g3400)) + ((g2980) & (!g3178) & (g3362) & (g3363) & (!g3365) & (g3400)) + ((g2980) & (!g3178) & (g3362) & (g3363) & (g3365) & (!g3400)) + ((g2980) & (!g3178) & (g3362) & (g3363) & (g3365) & (g3400)) + ((g2980) & (g3178) & (!g3362) & (!g3363) & (!g3365) & (!g3400)) + ((g2980) & (g3178) & (g3362) & (!g3363) & (!g3365) & (g3400)) + ((g2980) & (g3178) & (g3362) & (!g3363) & (g3365) & (!g3400)) + ((g2980) & (g3178) & (g3362) & (!g3363) & (g3365) & (g3400)) + ((g2980) & (g3178) & (g3362) & (g3363) & (!g3365) & (!g3400)) + ((g2980) & (g3178) & (g3362) & (g3363) & (!g3365) & (g3400)) + ((g2980) & (g3178) & (g3362) & (g3363) & (g3365) & (!g3400)) + ((g2980) & (g3178) & (g3362) & (g3363) & (g3365) & (g3400)));
	assign g3458 = (((!g3178) & (!g3363) & (g3365) & (!g3400)) + ((!g3178) & (g3363) & (!g3365) & (!g3400)) + ((!g3178) & (g3363) & (!g3365) & (g3400)) + ((!g3178) & (g3363) & (g3365) & (g3400)) + ((g3178) & (!g3363) & (!g3365) & (!g3400)) + ((g3178) & (g3363) & (!g3365) & (g3400)) + ((g3178) & (g3363) & (g3365) & (!g3400)) + ((g3178) & (g3363) & (g3365) & (g3400)));
	assign g3459 = (((!g3187) & (!ax6x) & (!ax7x) & (!g3395) & (!g3364) & (g3400)) + ((!g3187) & (!ax6x) & (!ax7x) & (!g3395) & (g3364) & (!g3400)) + ((!g3187) & (!ax6x) & (!ax7x) & (!g3395) & (g3364) & (g3400)) + ((!g3187) & (!ax6x) & (!ax7x) & (g3395) & (!g3364) & (!g3400)) + ((!g3187) & (!ax6x) & (ax7x) & (!g3395) & (!g3364) & (!g3400)) + ((!g3187) & (!ax6x) & (ax7x) & (g3395) & (!g3364) & (g3400)) + ((!g3187) & (!ax6x) & (ax7x) & (g3395) & (g3364) & (!g3400)) + ((!g3187) & (!ax6x) & (ax7x) & (g3395) & (g3364) & (g3400)) + ((!g3187) & (ax6x) & (!ax7x) & (g3395) & (!g3364) & (!g3400)) + ((!g3187) & (ax6x) & (!ax7x) & (g3395) & (g3364) & (!g3400)) + ((!g3187) & (ax6x) & (ax7x) & (!g3395) & (!g3364) & (!g3400)) + ((!g3187) & (ax6x) & (ax7x) & (!g3395) & (!g3364) & (g3400)) + ((!g3187) & (ax6x) & (ax7x) & (!g3395) & (g3364) & (!g3400)) + ((!g3187) & (ax6x) & (ax7x) & (!g3395) & (g3364) & (g3400)) + ((!g3187) & (ax6x) & (ax7x) & (g3395) & (!g3364) & (g3400)) + ((!g3187) & (ax6x) & (ax7x) & (g3395) & (g3364) & (g3400)) + ((g3187) & (!ax6x) & (!ax7x) & (!g3395) & (!g3364) & (!g3400)) + ((g3187) & (!ax6x) & (!ax7x) & (!g3395) & (!g3364) & (g3400)) + ((g3187) & (!ax6x) & (!ax7x) & (!g3395) & (g3364) & (g3400)) + ((g3187) & (!ax6x) & (!ax7x) & (g3395) & (g3364) & (!g3400)) + ((g3187) & (!ax6x) & (ax7x) & (!g3395) & (g3364) & (!g3400)) + ((g3187) & (!ax6x) & (ax7x) & (g3395) & (!g3364) & (!g3400)) + ((g3187) & (!ax6x) & (ax7x) & (g3395) & (!g3364) & (g3400)) + ((g3187) & (!ax6x) & (ax7x) & (g3395) & (g3364) & (g3400)) + ((g3187) & (ax6x) & (!ax7x) & (!g3395) & (!g3364) & (!g3400)) + ((g3187) & (ax6x) & (!ax7x) & (!g3395) & (g3364) & (!g3400)) + ((g3187) & (ax6x) & (ax7x) & (!g3395) & (!g3364) & (g3400)) + ((g3187) & (ax6x) & (ax7x) & (!g3395) & (g3364) & (g3400)) + ((g3187) & (ax6x) & (ax7x) & (g3395) & (!g3364) & (!g3400)) + ((g3187) & (ax6x) & (ax7x) & (g3395) & (!g3364) & (g3400)) + ((g3187) & (ax6x) & (ax7x) & (g3395) & (g3364) & (!g3400)) + ((g3187) & (ax6x) & (ax7x) & (g3395) & (g3364) & (g3400)));
	assign g3460 = (((!ax6x) & (!g3395) & (!g3364) & (g3400)) + ((!ax6x) & (!g3395) & (g3364) & (!g3400)) + ((!ax6x) & (!g3395) & (g3364) & (g3400)) + ((!ax6x) & (g3395) & (g3364) & (!g3400)) + ((ax6x) & (!g3395) & (!g3364) & (!g3400)) + ((ax6x) & (g3395) & (!g3364) & (!g3400)) + ((ax6x) & (g3395) & (!g3364) & (g3400)) + ((ax6x) & (g3395) & (g3364) & (g3400)));
	assign g3461 = (((!ax2x) & (!ax3x)));
	assign g3462 = (((!g3395) & (!ax4x) & (!ax5x) & (!g3400) & (!g3461)) + ((!g3395) & (!ax4x) & (ax5x) & (g3400) & (!g3461)) + ((!g3395) & (ax4x) & (ax5x) & (g3400) & (!g3461)) + ((!g3395) & (ax4x) & (ax5x) & (g3400) & (g3461)) + ((g3395) & (!ax4x) & (!ax5x) & (!g3400) & (!g3461)) + ((g3395) & (!ax4x) & (!ax5x) & (!g3400) & (g3461)) + ((g3395) & (!ax4x) & (!ax5x) & (g3400) & (!g3461)) + ((g3395) & (!ax4x) & (ax5x) & (!g3400) & (!g3461)) + ((g3395) & (!ax4x) & (ax5x) & (g3400) & (!g3461)) + ((g3395) & (!ax4x) & (ax5x) & (g3400) & (g3461)) + ((g3395) & (ax4x) & (!ax5x) & (g3400) & (!g3461)) + ((g3395) & (ax4x) & (!ax5x) & (g3400) & (g3461)) + ((g3395) & (ax4x) & (ax5x) & (!g3400) & (!g3461)) + ((g3395) & (ax4x) & (ax5x) & (!g3400) & (g3461)) + ((g3395) & (ax4x) & (ax5x) & (g3400) & (!g3461)) + ((g3395) & (ax4x) & (ax5x) & (g3400) & (g3461)));
	assign g3463 = (((!g3178) & (!g3187) & (g3459) & (g3460) & (g3462)) + ((!g3178) & (g3187) & (g3459) & (!g3460) & (g3462)) + ((!g3178) & (g3187) & (g3459) & (g3460) & (!g3462)) + ((!g3178) & (g3187) & (g3459) & (g3460) & (g3462)) + ((g3178) & (!g3187) & (!g3459) & (g3460) & (g3462)) + ((g3178) & (!g3187) & (g3459) & (!g3460) & (!g3462)) + ((g3178) & (!g3187) & (g3459) & (!g3460) & (g3462)) + ((g3178) & (!g3187) & (g3459) & (g3460) & (!g3462)) + ((g3178) & (!g3187) & (g3459) & (g3460) & (g3462)) + ((g3178) & (g3187) & (!g3459) & (!g3460) & (g3462)) + ((g3178) & (g3187) & (!g3459) & (g3460) & (!g3462)) + ((g3178) & (g3187) & (!g3459) & (g3460) & (g3462)) + ((g3178) & (g3187) & (g3459) & (!g3460) & (!g3462)) + ((g3178) & (g3187) & (g3459) & (!g3460) & (g3462)) + ((g3178) & (g3187) & (g3459) & (g3460) & (!g3462)) + ((g3178) & (g3187) & (g3459) & (g3460) & (g3462)));
	assign g3464 = (((!g3030) & (!g2980) & (g3457) & (g3458) & (g3463)) + ((!g3030) & (g2980) & (g3457) & (!g3458) & (g3463)) + ((!g3030) & (g2980) & (g3457) & (g3458) & (!g3463)) + ((!g3030) & (g2980) & (g3457) & (g3458) & (g3463)) + ((g3030) & (!g2980) & (!g3457) & (g3458) & (g3463)) + ((g3030) & (!g2980) & (g3457) & (!g3458) & (!g3463)) + ((g3030) & (!g2980) & (g3457) & (!g3458) & (g3463)) + ((g3030) & (!g2980) & (g3457) & (g3458) & (!g3463)) + ((g3030) & (!g2980) & (g3457) & (g3458) & (g3463)) + ((g3030) & (g2980) & (!g3457) & (!g3458) & (g3463)) + ((g3030) & (g2980) & (!g3457) & (g3458) & (!g3463)) + ((g3030) & (g2980) & (!g3457) & (g3458) & (g3463)) + ((g3030) & (g2980) & (g3457) & (!g3458) & (!g3463)) + ((g3030) & (g2980) & (g3457) & (!g3458) & (g3463)) + ((g3030) & (g2980) & (g3457) & (g3458) & (!g3463)) + ((g3030) & (g2980) & (g3457) & (g3458) & (g3463)));
	assign g3465 = (((!g2825) & (!g2779) & (g3455) & (g3456) & (g3464)) + ((!g2825) & (g2779) & (g3455) & (!g3456) & (g3464)) + ((!g2825) & (g2779) & (g3455) & (g3456) & (!g3464)) + ((!g2825) & (g2779) & (g3455) & (g3456) & (g3464)) + ((g2825) & (!g2779) & (!g3455) & (g3456) & (g3464)) + ((g2825) & (!g2779) & (g3455) & (!g3456) & (!g3464)) + ((g2825) & (!g2779) & (g3455) & (!g3456) & (g3464)) + ((g2825) & (!g2779) & (g3455) & (g3456) & (!g3464)) + ((g2825) & (!g2779) & (g3455) & (g3456) & (g3464)) + ((g2825) & (g2779) & (!g3455) & (!g3456) & (g3464)) + ((g2825) & (g2779) & (!g3455) & (g3456) & (!g3464)) + ((g2825) & (g2779) & (!g3455) & (g3456) & (g3464)) + ((g2825) & (g2779) & (g3455) & (!g3456) & (!g3464)) + ((g2825) & (g2779) & (g3455) & (!g3456) & (g3464)) + ((g2825) & (g2779) & (g3455) & (g3456) & (!g3464)) + ((g2825) & (g2779) & (g3455) & (g3456) & (g3464)));
	assign g3466 = (((!g2627) & (!g2585) & (g3453) & (g3454) & (g3465)) + ((!g2627) & (g2585) & (g3453) & (!g3454) & (g3465)) + ((!g2627) & (g2585) & (g3453) & (g3454) & (!g3465)) + ((!g2627) & (g2585) & (g3453) & (g3454) & (g3465)) + ((g2627) & (!g2585) & (!g3453) & (g3454) & (g3465)) + ((g2627) & (!g2585) & (g3453) & (!g3454) & (!g3465)) + ((g2627) & (!g2585) & (g3453) & (!g3454) & (g3465)) + ((g2627) & (!g2585) & (g3453) & (g3454) & (!g3465)) + ((g2627) & (!g2585) & (g3453) & (g3454) & (g3465)) + ((g2627) & (g2585) & (!g3453) & (!g3454) & (g3465)) + ((g2627) & (g2585) & (!g3453) & (g3454) & (!g3465)) + ((g2627) & (g2585) & (!g3453) & (g3454) & (g3465)) + ((g2627) & (g2585) & (g3453) & (!g3454) & (!g3465)) + ((g2627) & (g2585) & (g3453) & (!g3454) & (g3465)) + ((g2627) & (g2585) & (g3453) & (g3454) & (!g3465)) + ((g2627) & (g2585) & (g3453) & (g3454) & (g3465)));
	assign g3467 = (((!g2436) & (!g2398) & (g3451) & (g3452) & (g3466)) + ((!g2436) & (g2398) & (g3451) & (!g3452) & (g3466)) + ((!g2436) & (g2398) & (g3451) & (g3452) & (!g3466)) + ((!g2436) & (g2398) & (g3451) & (g3452) & (g3466)) + ((g2436) & (!g2398) & (!g3451) & (g3452) & (g3466)) + ((g2436) & (!g2398) & (g3451) & (!g3452) & (!g3466)) + ((g2436) & (!g2398) & (g3451) & (!g3452) & (g3466)) + ((g2436) & (!g2398) & (g3451) & (g3452) & (!g3466)) + ((g2436) & (!g2398) & (g3451) & (g3452) & (g3466)) + ((g2436) & (g2398) & (!g3451) & (!g3452) & (g3466)) + ((g2436) & (g2398) & (!g3451) & (g3452) & (!g3466)) + ((g2436) & (g2398) & (!g3451) & (g3452) & (g3466)) + ((g2436) & (g2398) & (g3451) & (!g3452) & (!g3466)) + ((g2436) & (g2398) & (g3451) & (!g3452) & (g3466)) + ((g2436) & (g2398) & (g3451) & (g3452) & (!g3466)) + ((g2436) & (g2398) & (g3451) & (g3452) & (g3466)));
	assign g3468 = (((!g2252) & (!g2218) & (g3449) & (g3450) & (g3467)) + ((!g2252) & (g2218) & (g3449) & (!g3450) & (g3467)) + ((!g2252) & (g2218) & (g3449) & (g3450) & (!g3467)) + ((!g2252) & (g2218) & (g3449) & (g3450) & (g3467)) + ((g2252) & (!g2218) & (!g3449) & (g3450) & (g3467)) + ((g2252) & (!g2218) & (g3449) & (!g3450) & (!g3467)) + ((g2252) & (!g2218) & (g3449) & (!g3450) & (g3467)) + ((g2252) & (!g2218) & (g3449) & (g3450) & (!g3467)) + ((g2252) & (!g2218) & (g3449) & (g3450) & (g3467)) + ((g2252) & (g2218) & (!g3449) & (!g3450) & (g3467)) + ((g2252) & (g2218) & (!g3449) & (g3450) & (!g3467)) + ((g2252) & (g2218) & (!g3449) & (g3450) & (g3467)) + ((g2252) & (g2218) & (g3449) & (!g3450) & (!g3467)) + ((g2252) & (g2218) & (g3449) & (!g3450) & (g3467)) + ((g2252) & (g2218) & (g3449) & (g3450) & (!g3467)) + ((g2252) & (g2218) & (g3449) & (g3450) & (g3467)));
	assign g3469 = (((!g2075) & (!g2045) & (g3447) & (g3448) & (g3468)) + ((!g2075) & (g2045) & (g3447) & (!g3448) & (g3468)) + ((!g2075) & (g2045) & (g3447) & (g3448) & (!g3468)) + ((!g2075) & (g2045) & (g3447) & (g3448) & (g3468)) + ((g2075) & (!g2045) & (!g3447) & (g3448) & (g3468)) + ((g2075) & (!g2045) & (g3447) & (!g3448) & (!g3468)) + ((g2075) & (!g2045) & (g3447) & (!g3448) & (g3468)) + ((g2075) & (!g2045) & (g3447) & (g3448) & (!g3468)) + ((g2075) & (!g2045) & (g3447) & (g3448) & (g3468)) + ((g2075) & (g2045) & (!g3447) & (!g3448) & (g3468)) + ((g2075) & (g2045) & (!g3447) & (g3448) & (!g3468)) + ((g2075) & (g2045) & (!g3447) & (g3448) & (g3468)) + ((g2075) & (g2045) & (g3447) & (!g3448) & (!g3468)) + ((g2075) & (g2045) & (g3447) & (!g3448) & (g3468)) + ((g2075) & (g2045) & (g3447) & (g3448) & (!g3468)) + ((g2075) & (g2045) & (g3447) & (g3448) & (g3468)));
	assign g3470 = (((!g1905) & (!g1879) & (g3445) & (g3446) & (g3469)) + ((!g1905) & (g1879) & (g3445) & (!g3446) & (g3469)) + ((!g1905) & (g1879) & (g3445) & (g3446) & (!g3469)) + ((!g1905) & (g1879) & (g3445) & (g3446) & (g3469)) + ((g1905) & (!g1879) & (!g3445) & (g3446) & (g3469)) + ((g1905) & (!g1879) & (g3445) & (!g3446) & (!g3469)) + ((g1905) & (!g1879) & (g3445) & (!g3446) & (g3469)) + ((g1905) & (!g1879) & (g3445) & (g3446) & (!g3469)) + ((g1905) & (!g1879) & (g3445) & (g3446) & (g3469)) + ((g1905) & (g1879) & (!g3445) & (!g3446) & (g3469)) + ((g1905) & (g1879) & (!g3445) & (g3446) & (!g3469)) + ((g1905) & (g1879) & (!g3445) & (g3446) & (g3469)) + ((g1905) & (g1879) & (g3445) & (!g3446) & (!g3469)) + ((g1905) & (g1879) & (g3445) & (!g3446) & (g3469)) + ((g1905) & (g1879) & (g3445) & (g3446) & (!g3469)) + ((g1905) & (g1879) & (g3445) & (g3446) & (g3469)));
	assign g3471 = (((!g1742) & (!g1720) & (g3443) & (g3444) & (g3470)) + ((!g1742) & (g1720) & (g3443) & (!g3444) & (g3470)) + ((!g1742) & (g1720) & (g3443) & (g3444) & (!g3470)) + ((!g1742) & (g1720) & (g3443) & (g3444) & (g3470)) + ((g1742) & (!g1720) & (!g3443) & (g3444) & (g3470)) + ((g1742) & (!g1720) & (g3443) & (!g3444) & (!g3470)) + ((g1742) & (!g1720) & (g3443) & (!g3444) & (g3470)) + ((g1742) & (!g1720) & (g3443) & (g3444) & (!g3470)) + ((g1742) & (!g1720) & (g3443) & (g3444) & (g3470)) + ((g1742) & (g1720) & (!g3443) & (!g3444) & (g3470)) + ((g1742) & (g1720) & (!g3443) & (g3444) & (!g3470)) + ((g1742) & (g1720) & (!g3443) & (g3444) & (g3470)) + ((g1742) & (g1720) & (g3443) & (!g3444) & (!g3470)) + ((g1742) & (g1720) & (g3443) & (!g3444) & (g3470)) + ((g1742) & (g1720) & (g3443) & (g3444) & (!g3470)) + ((g1742) & (g1720) & (g3443) & (g3444) & (g3470)));
	assign g3472 = (((!g1586) & (!g1568) & (g3441) & (g3442) & (g3471)) + ((!g1586) & (g1568) & (g3441) & (!g3442) & (g3471)) + ((!g1586) & (g1568) & (g3441) & (g3442) & (!g3471)) + ((!g1586) & (g1568) & (g3441) & (g3442) & (g3471)) + ((g1586) & (!g1568) & (!g3441) & (g3442) & (g3471)) + ((g1586) & (!g1568) & (g3441) & (!g3442) & (!g3471)) + ((g1586) & (!g1568) & (g3441) & (!g3442) & (g3471)) + ((g1586) & (!g1568) & (g3441) & (g3442) & (!g3471)) + ((g1586) & (!g1568) & (g3441) & (g3442) & (g3471)) + ((g1586) & (g1568) & (!g3441) & (!g3442) & (g3471)) + ((g1586) & (g1568) & (!g3441) & (g3442) & (!g3471)) + ((g1586) & (g1568) & (!g3441) & (g3442) & (g3471)) + ((g1586) & (g1568) & (g3441) & (!g3442) & (!g3471)) + ((g1586) & (g1568) & (g3441) & (!g3442) & (g3471)) + ((g1586) & (g1568) & (g3441) & (g3442) & (!g3471)) + ((g1586) & (g1568) & (g3441) & (g3442) & (g3471)));
	assign g3473 = (((!g1437) & (!g1423) & (g3439) & (g3440) & (g3472)) + ((!g1437) & (g1423) & (g3439) & (!g3440) & (g3472)) + ((!g1437) & (g1423) & (g3439) & (g3440) & (!g3472)) + ((!g1437) & (g1423) & (g3439) & (g3440) & (g3472)) + ((g1437) & (!g1423) & (!g3439) & (g3440) & (g3472)) + ((g1437) & (!g1423) & (g3439) & (!g3440) & (!g3472)) + ((g1437) & (!g1423) & (g3439) & (!g3440) & (g3472)) + ((g1437) & (!g1423) & (g3439) & (g3440) & (!g3472)) + ((g1437) & (!g1423) & (g3439) & (g3440) & (g3472)) + ((g1437) & (g1423) & (!g3439) & (!g3440) & (g3472)) + ((g1437) & (g1423) & (!g3439) & (g3440) & (!g3472)) + ((g1437) & (g1423) & (!g3439) & (g3440) & (g3472)) + ((g1437) & (g1423) & (g3439) & (!g3440) & (!g3472)) + ((g1437) & (g1423) & (g3439) & (!g3440) & (g3472)) + ((g1437) & (g1423) & (g3439) & (g3440) & (!g3472)) + ((g1437) & (g1423) & (g3439) & (g3440) & (g3472)));
	assign g3474 = (((!g1295) & (!g1285) & (g3437) & (g3438) & (g3473)) + ((!g1295) & (g1285) & (g3437) & (!g3438) & (g3473)) + ((!g1295) & (g1285) & (g3437) & (g3438) & (!g3473)) + ((!g1295) & (g1285) & (g3437) & (g3438) & (g3473)) + ((g1295) & (!g1285) & (!g3437) & (g3438) & (g3473)) + ((g1295) & (!g1285) & (g3437) & (!g3438) & (!g3473)) + ((g1295) & (!g1285) & (g3437) & (!g3438) & (g3473)) + ((g1295) & (!g1285) & (g3437) & (g3438) & (!g3473)) + ((g1295) & (!g1285) & (g3437) & (g3438) & (g3473)) + ((g1295) & (g1285) & (!g3437) & (!g3438) & (g3473)) + ((g1295) & (g1285) & (!g3437) & (g3438) & (!g3473)) + ((g1295) & (g1285) & (!g3437) & (g3438) & (g3473)) + ((g1295) & (g1285) & (g3437) & (!g3438) & (!g3473)) + ((g1295) & (g1285) & (g3437) & (!g3438) & (g3473)) + ((g1295) & (g1285) & (g3437) & (g3438) & (!g3473)) + ((g1295) & (g1285) & (g3437) & (g3438) & (g3473)));
	assign g3475 = (((!g1160) & (!g1154) & (g3435) & (g3436) & (g3474)) + ((!g1160) & (g1154) & (g3435) & (!g3436) & (g3474)) + ((!g1160) & (g1154) & (g3435) & (g3436) & (!g3474)) + ((!g1160) & (g1154) & (g3435) & (g3436) & (g3474)) + ((g1160) & (!g1154) & (!g3435) & (g3436) & (g3474)) + ((g1160) & (!g1154) & (g3435) & (!g3436) & (!g3474)) + ((g1160) & (!g1154) & (g3435) & (!g3436) & (g3474)) + ((g1160) & (!g1154) & (g3435) & (g3436) & (!g3474)) + ((g1160) & (!g1154) & (g3435) & (g3436) & (g3474)) + ((g1160) & (g1154) & (!g3435) & (!g3436) & (g3474)) + ((g1160) & (g1154) & (!g3435) & (g3436) & (!g3474)) + ((g1160) & (g1154) & (!g3435) & (g3436) & (g3474)) + ((g1160) & (g1154) & (g3435) & (!g3436) & (!g3474)) + ((g1160) & (g1154) & (g3435) & (!g3436) & (g3474)) + ((g1160) & (g1154) & (g3435) & (g3436) & (!g3474)) + ((g1160) & (g1154) & (g3435) & (g3436) & (g3474)));
	assign g3476 = (((!g1032) & (!g1030) & (g3433) & (g3434) & (g3475)) + ((!g1032) & (g1030) & (g3433) & (!g3434) & (g3475)) + ((!g1032) & (g1030) & (g3433) & (g3434) & (!g3475)) + ((!g1032) & (g1030) & (g3433) & (g3434) & (g3475)) + ((g1032) & (!g1030) & (!g3433) & (g3434) & (g3475)) + ((g1032) & (!g1030) & (g3433) & (!g3434) & (!g3475)) + ((g1032) & (!g1030) & (g3433) & (!g3434) & (g3475)) + ((g1032) & (!g1030) & (g3433) & (g3434) & (!g3475)) + ((g1032) & (!g1030) & (g3433) & (g3434) & (g3475)) + ((g1032) & (g1030) & (!g3433) & (!g3434) & (g3475)) + ((g1032) & (g1030) & (!g3433) & (g3434) & (!g3475)) + ((g1032) & (g1030) & (!g3433) & (g3434) & (g3475)) + ((g1032) & (g1030) & (g3433) & (!g3434) & (!g3475)) + ((g1032) & (g1030) & (g3433) & (!g3434) & (g3475)) + ((g1032) & (g1030) & (g3433) & (g3434) & (!g3475)) + ((g1032) & (g1030) & (g3433) & (g3434) & (g3475)));
	assign g3477 = (((!g851) & (!g914) & (g3431) & (g3432) & (g3476)) + ((!g851) & (g914) & (g3431) & (!g3432) & (g3476)) + ((!g851) & (g914) & (g3431) & (g3432) & (!g3476)) + ((!g851) & (g914) & (g3431) & (g3432) & (g3476)) + ((g851) & (!g914) & (!g3431) & (g3432) & (g3476)) + ((g851) & (!g914) & (g3431) & (!g3432) & (!g3476)) + ((g851) & (!g914) & (g3431) & (!g3432) & (g3476)) + ((g851) & (!g914) & (g3431) & (g3432) & (!g3476)) + ((g851) & (!g914) & (g3431) & (g3432) & (g3476)) + ((g851) & (g914) & (!g3431) & (!g3432) & (g3476)) + ((g851) & (g914) & (!g3431) & (g3432) & (!g3476)) + ((g851) & (g914) & (!g3431) & (g3432) & (g3476)) + ((g851) & (g914) & (g3431) & (!g3432) & (!g3476)) + ((g851) & (g914) & (g3431) & (!g3432) & (g3476)) + ((g851) & (g914) & (g3431) & (g3432) & (!g3476)) + ((g851) & (g914) & (g3431) & (g3432) & (g3476)));
	assign g3478 = (((!g744) & (!g803) & (g3429) & (g3430) & (g3477)) + ((!g744) & (g803) & (g3429) & (!g3430) & (g3477)) + ((!g744) & (g803) & (g3429) & (g3430) & (!g3477)) + ((!g744) & (g803) & (g3429) & (g3430) & (g3477)) + ((g744) & (!g803) & (!g3429) & (g3430) & (g3477)) + ((g744) & (!g803) & (g3429) & (!g3430) & (!g3477)) + ((g744) & (!g803) & (g3429) & (!g3430) & (g3477)) + ((g744) & (!g803) & (g3429) & (g3430) & (!g3477)) + ((g744) & (!g803) & (g3429) & (g3430) & (g3477)) + ((g744) & (g803) & (!g3429) & (!g3430) & (g3477)) + ((g744) & (g803) & (!g3429) & (g3430) & (!g3477)) + ((g744) & (g803) & (!g3429) & (g3430) & (g3477)) + ((g744) & (g803) & (g3429) & (!g3430) & (!g3477)) + ((g744) & (g803) & (g3429) & (!g3430) & (g3477)) + ((g744) & (g803) & (g3429) & (g3430) & (!g3477)) + ((g744) & (g803) & (g3429) & (g3430) & (g3477)));
	assign g3479 = (((!g645) & (!g700) & (g3427) & (g3428) & (g3478)) + ((!g645) & (g700) & (g3427) & (!g3428) & (g3478)) + ((!g645) & (g700) & (g3427) & (g3428) & (!g3478)) + ((!g645) & (g700) & (g3427) & (g3428) & (g3478)) + ((g645) & (!g700) & (!g3427) & (g3428) & (g3478)) + ((g645) & (!g700) & (g3427) & (!g3428) & (!g3478)) + ((g645) & (!g700) & (g3427) & (!g3428) & (g3478)) + ((g645) & (!g700) & (g3427) & (g3428) & (!g3478)) + ((g645) & (!g700) & (g3427) & (g3428) & (g3478)) + ((g645) & (g700) & (!g3427) & (!g3428) & (g3478)) + ((g645) & (g700) & (!g3427) & (g3428) & (!g3478)) + ((g645) & (g700) & (!g3427) & (g3428) & (g3478)) + ((g645) & (g700) & (g3427) & (!g3428) & (!g3478)) + ((g645) & (g700) & (g3427) & (!g3428) & (g3478)) + ((g645) & (g700) & (g3427) & (g3428) & (!g3478)) + ((g645) & (g700) & (g3427) & (g3428) & (g3478)));
	assign g3480 = (((!g553) & (!g604) & (g3425) & (g3426) & (g3479)) + ((!g553) & (g604) & (g3425) & (!g3426) & (g3479)) + ((!g553) & (g604) & (g3425) & (g3426) & (!g3479)) + ((!g553) & (g604) & (g3425) & (g3426) & (g3479)) + ((g553) & (!g604) & (!g3425) & (g3426) & (g3479)) + ((g553) & (!g604) & (g3425) & (!g3426) & (!g3479)) + ((g553) & (!g604) & (g3425) & (!g3426) & (g3479)) + ((g553) & (!g604) & (g3425) & (g3426) & (!g3479)) + ((g553) & (!g604) & (g3425) & (g3426) & (g3479)) + ((g553) & (g604) & (!g3425) & (!g3426) & (g3479)) + ((g553) & (g604) & (!g3425) & (g3426) & (!g3479)) + ((g553) & (g604) & (!g3425) & (g3426) & (g3479)) + ((g553) & (g604) & (g3425) & (!g3426) & (!g3479)) + ((g553) & (g604) & (g3425) & (!g3426) & (g3479)) + ((g553) & (g604) & (g3425) & (g3426) & (!g3479)) + ((g553) & (g604) & (g3425) & (g3426) & (g3479)));
	assign g3481 = (((!g468) & (!g515) & (g3423) & (g3424) & (g3480)) + ((!g468) & (g515) & (g3423) & (!g3424) & (g3480)) + ((!g468) & (g515) & (g3423) & (g3424) & (!g3480)) + ((!g468) & (g515) & (g3423) & (g3424) & (g3480)) + ((g468) & (!g515) & (!g3423) & (g3424) & (g3480)) + ((g468) & (!g515) & (g3423) & (!g3424) & (!g3480)) + ((g468) & (!g515) & (g3423) & (!g3424) & (g3480)) + ((g468) & (!g515) & (g3423) & (g3424) & (!g3480)) + ((g468) & (!g515) & (g3423) & (g3424) & (g3480)) + ((g468) & (g515) & (!g3423) & (!g3424) & (g3480)) + ((g468) & (g515) & (!g3423) & (g3424) & (!g3480)) + ((g468) & (g515) & (!g3423) & (g3424) & (g3480)) + ((g468) & (g515) & (g3423) & (!g3424) & (!g3480)) + ((g468) & (g515) & (g3423) & (!g3424) & (g3480)) + ((g468) & (g515) & (g3423) & (g3424) & (!g3480)) + ((g468) & (g515) & (g3423) & (g3424) & (g3480)));
	assign g3482 = (((!g390) & (!g433) & (g3421) & (g3422) & (g3481)) + ((!g390) & (g433) & (g3421) & (!g3422) & (g3481)) + ((!g390) & (g433) & (g3421) & (g3422) & (!g3481)) + ((!g390) & (g433) & (g3421) & (g3422) & (g3481)) + ((g390) & (!g433) & (!g3421) & (g3422) & (g3481)) + ((g390) & (!g433) & (g3421) & (!g3422) & (!g3481)) + ((g390) & (!g433) & (g3421) & (!g3422) & (g3481)) + ((g390) & (!g433) & (g3421) & (g3422) & (!g3481)) + ((g390) & (!g433) & (g3421) & (g3422) & (g3481)) + ((g390) & (g433) & (!g3421) & (!g3422) & (g3481)) + ((g390) & (g433) & (!g3421) & (g3422) & (!g3481)) + ((g390) & (g433) & (!g3421) & (g3422) & (g3481)) + ((g390) & (g433) & (g3421) & (!g3422) & (!g3481)) + ((g390) & (g433) & (g3421) & (!g3422) & (g3481)) + ((g390) & (g433) & (g3421) & (g3422) & (!g3481)) + ((g390) & (g433) & (g3421) & (g3422) & (g3481)));
	assign g3483 = (((!g319) & (!g358) & (g3419) & (g3420) & (g3482)) + ((!g319) & (g358) & (g3419) & (!g3420) & (g3482)) + ((!g319) & (g358) & (g3419) & (g3420) & (!g3482)) + ((!g319) & (g358) & (g3419) & (g3420) & (g3482)) + ((g319) & (!g358) & (!g3419) & (g3420) & (g3482)) + ((g319) & (!g358) & (g3419) & (!g3420) & (!g3482)) + ((g319) & (!g358) & (g3419) & (!g3420) & (g3482)) + ((g319) & (!g358) & (g3419) & (g3420) & (!g3482)) + ((g319) & (!g358) & (g3419) & (g3420) & (g3482)) + ((g319) & (g358) & (!g3419) & (!g3420) & (g3482)) + ((g319) & (g358) & (!g3419) & (g3420) & (!g3482)) + ((g319) & (g358) & (!g3419) & (g3420) & (g3482)) + ((g319) & (g358) & (g3419) & (!g3420) & (!g3482)) + ((g319) & (g358) & (g3419) & (!g3420) & (g3482)) + ((g319) & (g358) & (g3419) & (g3420) & (!g3482)) + ((g319) & (g358) & (g3419) & (g3420) & (g3482)));
	assign g3484 = (((!g255) & (!g290) & (g3417) & (g3418) & (g3483)) + ((!g255) & (g290) & (g3417) & (!g3418) & (g3483)) + ((!g255) & (g290) & (g3417) & (g3418) & (!g3483)) + ((!g255) & (g290) & (g3417) & (g3418) & (g3483)) + ((g255) & (!g290) & (!g3417) & (g3418) & (g3483)) + ((g255) & (!g290) & (g3417) & (!g3418) & (!g3483)) + ((g255) & (!g290) & (g3417) & (!g3418) & (g3483)) + ((g255) & (!g290) & (g3417) & (g3418) & (!g3483)) + ((g255) & (!g290) & (g3417) & (g3418) & (g3483)) + ((g255) & (g290) & (!g3417) & (!g3418) & (g3483)) + ((g255) & (g290) & (!g3417) & (g3418) & (!g3483)) + ((g255) & (g290) & (!g3417) & (g3418) & (g3483)) + ((g255) & (g290) & (g3417) & (!g3418) & (!g3483)) + ((g255) & (g290) & (g3417) & (!g3418) & (g3483)) + ((g255) & (g290) & (g3417) & (g3418) & (!g3483)) + ((g255) & (g290) & (g3417) & (g3418) & (g3483)));
	assign g3485 = (((!g198) & (!g229) & (g3415) & (g3416) & (g3484)) + ((!g198) & (g229) & (g3415) & (!g3416) & (g3484)) + ((!g198) & (g229) & (g3415) & (g3416) & (!g3484)) + ((!g198) & (g229) & (g3415) & (g3416) & (g3484)) + ((g198) & (!g229) & (!g3415) & (g3416) & (g3484)) + ((g198) & (!g229) & (g3415) & (!g3416) & (!g3484)) + ((g198) & (!g229) & (g3415) & (!g3416) & (g3484)) + ((g198) & (!g229) & (g3415) & (g3416) & (!g3484)) + ((g198) & (!g229) & (g3415) & (g3416) & (g3484)) + ((g198) & (g229) & (!g3415) & (!g3416) & (g3484)) + ((g198) & (g229) & (!g3415) & (g3416) & (!g3484)) + ((g198) & (g229) & (!g3415) & (g3416) & (g3484)) + ((g198) & (g229) & (g3415) & (!g3416) & (!g3484)) + ((g198) & (g229) & (g3415) & (!g3416) & (g3484)) + ((g198) & (g229) & (g3415) & (g3416) & (!g3484)) + ((g198) & (g229) & (g3415) & (g3416) & (g3484)));
	assign g3486 = (((!g147) & (!g174) & (g3413) & (g3414) & (g3485)) + ((!g147) & (g174) & (g3413) & (!g3414) & (g3485)) + ((!g147) & (g174) & (g3413) & (g3414) & (!g3485)) + ((!g147) & (g174) & (g3413) & (g3414) & (g3485)) + ((g147) & (!g174) & (!g3413) & (g3414) & (g3485)) + ((g147) & (!g174) & (g3413) & (!g3414) & (!g3485)) + ((g147) & (!g174) & (g3413) & (!g3414) & (g3485)) + ((g147) & (!g174) & (g3413) & (g3414) & (!g3485)) + ((g147) & (!g174) & (g3413) & (g3414) & (g3485)) + ((g147) & (g174) & (!g3413) & (!g3414) & (g3485)) + ((g147) & (g174) & (!g3413) & (g3414) & (!g3485)) + ((g147) & (g174) & (!g3413) & (g3414) & (g3485)) + ((g147) & (g174) & (g3413) & (!g3414) & (!g3485)) + ((g147) & (g174) & (g3413) & (!g3414) & (g3485)) + ((g147) & (g174) & (g3413) & (g3414) & (!g3485)) + ((g147) & (g174) & (g3413) & (g3414) & (g3485)));
	assign g3487 = (((!g104) & (!g127) & (g3411) & (g3412) & (g3486)) + ((!g104) & (g127) & (g3411) & (!g3412) & (g3486)) + ((!g104) & (g127) & (g3411) & (g3412) & (!g3486)) + ((!g104) & (g127) & (g3411) & (g3412) & (g3486)) + ((g104) & (!g127) & (!g3411) & (g3412) & (g3486)) + ((g104) & (!g127) & (g3411) & (!g3412) & (!g3486)) + ((g104) & (!g127) & (g3411) & (!g3412) & (g3486)) + ((g104) & (!g127) & (g3411) & (g3412) & (!g3486)) + ((g104) & (!g127) & (g3411) & (g3412) & (g3486)) + ((g104) & (g127) & (!g3411) & (!g3412) & (g3486)) + ((g104) & (g127) & (!g3411) & (g3412) & (!g3486)) + ((g104) & (g127) & (!g3411) & (g3412) & (g3486)) + ((g104) & (g127) & (g3411) & (!g3412) & (!g3486)) + ((g104) & (g127) & (g3411) & (!g3412) & (g3486)) + ((g104) & (g127) & (g3411) & (g3412) & (!g3486)) + ((g104) & (g127) & (g3411) & (g3412) & (g3486)));
	assign g3488 = (((!g68) & (!g87) & (g3409) & (g3410) & (g3487)) + ((!g68) & (g87) & (g3409) & (!g3410) & (g3487)) + ((!g68) & (g87) & (g3409) & (g3410) & (!g3487)) + ((!g68) & (g87) & (g3409) & (g3410) & (g3487)) + ((g68) & (!g87) & (!g3409) & (g3410) & (g3487)) + ((g68) & (!g87) & (g3409) & (!g3410) & (!g3487)) + ((g68) & (!g87) & (g3409) & (!g3410) & (g3487)) + ((g68) & (!g87) & (g3409) & (g3410) & (!g3487)) + ((g68) & (!g87) & (g3409) & (g3410) & (g3487)) + ((g68) & (g87) & (!g3409) & (!g3410) & (g3487)) + ((g68) & (g87) & (!g3409) & (g3410) & (!g3487)) + ((g68) & (g87) & (!g3409) & (g3410) & (g3487)) + ((g68) & (g87) & (g3409) & (!g3410) & (!g3487)) + ((g68) & (g87) & (g3409) & (!g3410) & (g3487)) + ((g68) & (g87) & (g3409) & (g3410) & (!g3487)) + ((g68) & (g87) & (g3409) & (g3410) & (g3487)));
	assign g3489 = (((!g39) & (!g54) & (g3407) & (g3408) & (g3488)) + ((!g39) & (g54) & (g3407) & (!g3408) & (g3488)) + ((!g39) & (g54) & (g3407) & (g3408) & (!g3488)) + ((!g39) & (g54) & (g3407) & (g3408) & (g3488)) + ((g39) & (!g54) & (!g3407) & (g3408) & (g3488)) + ((g39) & (!g54) & (g3407) & (!g3408) & (!g3488)) + ((g39) & (!g54) & (g3407) & (!g3408) & (g3488)) + ((g39) & (!g54) & (g3407) & (g3408) & (!g3488)) + ((g39) & (!g54) & (g3407) & (g3408) & (g3488)) + ((g39) & (g54) & (!g3407) & (!g3408) & (g3488)) + ((g39) & (g54) & (!g3407) & (g3408) & (!g3488)) + ((g39) & (g54) & (!g3407) & (g3408) & (g3488)) + ((g39) & (g54) & (g3407) & (!g3408) & (!g3488)) + ((g39) & (g54) & (g3407) & (!g3408) & (g3488)) + ((g39) & (g54) & (g3407) & (g3408) & (!g3488)) + ((g39) & (g54) & (g3407) & (g3408) & (g3488)));
	assign g3490 = (((!g18) & (!g27) & (g3405) & (g3406) & (g3489)) + ((!g18) & (g27) & (g3405) & (!g3406) & (g3489)) + ((!g18) & (g27) & (g3405) & (g3406) & (!g3489)) + ((!g18) & (g27) & (g3405) & (g3406) & (g3489)) + ((g18) & (!g27) & (!g3405) & (g3406) & (g3489)) + ((g18) & (!g27) & (g3405) & (!g3406) & (!g3489)) + ((g18) & (!g27) & (g3405) & (!g3406) & (g3489)) + ((g18) & (!g27) & (g3405) & (g3406) & (!g3489)) + ((g18) & (!g27) & (g3405) & (g3406) & (g3489)) + ((g18) & (g27) & (!g3405) & (!g3406) & (g3489)) + ((g18) & (g27) & (!g3405) & (g3406) & (!g3489)) + ((g18) & (g27) & (!g3405) & (g3406) & (g3489)) + ((g18) & (g27) & (g3405) & (!g3406) & (!g3489)) + ((g18) & (g27) & (g3405) & (!g3406) & (g3489)) + ((g18) & (g27) & (g3405) & (g3406) & (!g3489)) + ((g18) & (g27) & (g3405) & (g3406) & (g3489)));
	assign g3491 = (((!g2) & (!g8) & (g3403) & (g3404) & (g3490)) + ((!g2) & (g8) & (g3403) & (!g3404) & (g3490)) + ((!g2) & (g8) & (g3403) & (g3404) & (!g3490)) + ((!g2) & (g8) & (g3403) & (g3404) & (g3490)) + ((g2) & (!g8) & (!g3403) & (g3404) & (g3490)) + ((g2) & (!g8) & (g3403) & (!g3404) & (!g3490)) + ((g2) & (!g8) & (g3403) & (!g3404) & (g3490)) + ((g2) & (!g8) & (g3403) & (g3404) & (!g3490)) + ((g2) & (!g8) & (g3403) & (g3404) & (g3490)) + ((g2) & (g8) & (!g3403) & (!g3404) & (g3490)) + ((g2) & (g8) & (!g3403) & (g3404) & (!g3490)) + ((g2) & (g8) & (!g3403) & (g3404) & (g3490)) + ((g2) & (g8) & (g3403) & (!g3404) & (!g3490)) + ((g2) & (g8) & (g3403) & (!g3404) & (g3490)) + ((g2) & (g8) & (g3403) & (g3404) & (!g3490)) + ((g2) & (g8) & (g3403) & (g3404) & (g3490)));
	assign g3492 = (((!g1) & (!g3273) & (!g3394) & (!g3395) & (!g3396) & (!g3399)) + ((!g1) & (!g3273) & (!g3394) & (!g3395) & (g3396) & (g3399)) + ((!g1) & (!g3273) & (!g3394) & (g3395) & (g3396) & (g3399)) + ((!g1) & (!g3273) & (g3394) & (!g3395) & (g3396) & (g3399)) + ((!g1) & (!g3273) & (g3394) & (g3395) & (g3396) & (g3399)) + ((!g1) & (g3273) & (!g3394) & (!g3395) & (g3396) & (g3399)) + ((!g1) & (g3273) & (!g3394) & (g3395) & (g3396) & (g3399)) + ((!g1) & (g3273) & (g3394) & (!g3395) & (!g3396) & (!g3399)) + ((!g1) & (g3273) & (g3394) & (!g3395) & (g3396) & (g3399)) + ((!g1) & (g3273) & (g3394) & (g3395) & (!g3396) & (!g3399)) + ((!g1) & (g3273) & (g3394) & (g3395) & (g3396) & (g3399)) + ((g1) & (!g3273) & (!g3394) & (!g3395) & (g3396) & (g3399)) + ((g1) & (!g3273) & (!g3394) & (g3395) & (g3396) & (g3399)) + ((g1) & (!g3273) & (g3394) & (!g3395) & (!g3396) & (!g3399)) + ((g1) & (!g3273) & (g3394) & (!g3395) & (g3396) & (g3399)) + ((g1) & (!g3273) & (g3394) & (g3395) & (g3396) & (g3399)) + ((g1) & (g3273) & (!g3394) & (!g3395) & (!g3396) & (!g3399)) + ((g1) & (g3273) & (!g3394) & (!g3395) & (g3396) & (g3399)) + ((g1) & (g3273) & (!g3394) & (g3395) & (!g3396) & (!g3399)) + ((g1) & (g3273) & (!g3394) & (g3395) & (g3396) & (g3399)) + ((g1) & (g3273) & (g3394) & (!g3395) & (g3396) & (g3399)) + ((g1) & (g3273) & (g3394) & (g3395) & (g3396) & (g3399)));
	assign g3493 = (((!g4) & (!g1) & (!g3402) & (!g3491) & (!g3401) & (g3492)) + ((!g4) & (!g1) & (!g3402) & (!g3491) & (g3401) & (!g3492)) + ((!g4) & (!g1) & (!g3402) & (!g3491) & (g3401) & (g3492)) + ((!g4) & (!g1) & (!g3402) & (g3491) & (!g3401) & (!g3492)) + ((!g4) & (!g1) & (!g3402) & (g3491) & (!g3401) & (g3492)) + ((!g4) & (!g1) & (!g3402) & (g3491) & (g3401) & (!g3492)) + ((!g4) & (!g1) & (!g3402) & (g3491) & (g3401) & (g3492)) + ((!g4) & (!g1) & (g3402) & (!g3491) & (!g3401) & (!g3492)) + ((!g4) & (!g1) & (g3402) & (!g3491) & (!g3401) & (g3492)) + ((!g4) & (!g1) & (g3402) & (!g3491) & (g3401) & (!g3492)) + ((!g4) & (!g1) & (g3402) & (!g3491) & (g3401) & (g3492)) + ((!g4) & (!g1) & (g3402) & (g3491) & (!g3401) & (!g3492)) + ((!g4) & (!g1) & (g3402) & (g3491) & (!g3401) & (g3492)) + ((!g4) & (!g1) & (g3402) & (g3491) & (g3401) & (!g3492)) + ((!g4) & (!g1) & (g3402) & (g3491) & (g3401) & (g3492)) + ((g4) & (!g1) & (!g3402) & (!g3491) & (!g3401) & (g3492)) + ((g4) & (!g1) & (!g3402) & (!g3491) & (g3401) & (g3492)) + ((g4) & (!g1) & (!g3402) & (g3491) & (!g3401) & (g3492)) + ((g4) & (!g1) & (!g3402) & (g3491) & (g3401) & (!g3492)) + ((g4) & (!g1) & (!g3402) & (g3491) & (g3401) & (g3492)) + ((g4) & (!g1) & (g3402) & (!g3491) & (!g3401) & (!g3492)) + ((g4) & (!g1) & (g3402) & (!g3491) & (!g3401) & (g3492)) + ((g4) & (!g1) & (g3402) & (!g3491) & (g3401) & (!g3492)) + ((g4) & (!g1) & (g3402) & (!g3491) & (g3401) & (g3492)) + ((g4) & (!g1) & (g3402) & (g3491) & (!g3401) & (!g3492)) + ((g4) & (!g1) & (g3402) & (g3491) & (!g3401) & (g3492)) + ((g4) & (!g1) & (g3402) & (g3491) & (g3401) & (!g3492)) + ((g4) & (!g1) & (g3402) & (g3491) & (g3401) & (g3492)));
	assign g3494 = (((g1) & (!g3273) & (!g3394) & (!g3395) & (g3396) & (!g3399)) + ((g1) & (!g3273) & (!g3394) & (g3395) & (g3396) & (!g3399)) + ((g1) & (!g3273) & (g3394) & (!g3395) & (!g3396) & (g3399)) + ((g1) & (!g3273) & (g3394) & (!g3395) & (g3396) & (!g3399)) + ((g1) & (!g3273) & (g3394) & (g3395) & (g3396) & (!g3399)) + ((g1) & (g3273) & (!g3394) & (!g3395) & (!g3396) & (g3399)) + ((g1) & (g3273) & (!g3394) & (!g3395) & (g3396) & (!g3399)) + ((g1) & (g3273) & (!g3394) & (g3395) & (!g3396) & (g3399)) + ((g1) & (g3273) & (!g3394) & (g3395) & (g3396) & (!g3399)) + ((g1) & (g3273) & (g3394) & (!g3395) & (g3396) & (!g3399)) + ((g1) & (g3273) & (g3394) & (g3395) & (g3396) & (!g3399)));
	assign g3495 = (((!g4) & (!g3402) & (!g3491) & (!g3401) & (!g3494)) + ((!g4) & (!g3402) & (!g3491) & (g3401) & (!g3494)) + ((!g4) & (!g3402) & (g3491) & (!g3401) & (!g3494)) + ((!g4) & (!g3402) & (g3491) & (g3401) & (!g3494)) + ((!g4) & (g3402) & (!g3491) & (!g3401) & (!g3494)) + ((g4) & (!g3402) & (!g3491) & (!g3401) & (!g3494)) + ((g4) & (!g3402) & (!g3491) & (g3401) & (!g3494)) + ((g4) & (!g3402) & (g3491) & (!g3401) & (!g3494)) + ((g4) & (!g3402) & (g3491) & (g3401) & (!g3494)) + ((g4) & (g3402) & (!g3491) & (!g3401) & (!g3494)) + ((g4) & (g3402) & (!g3491) & (g3401) & (!g3494)) + ((g4) & (g3402) & (g3491) & (!g3401) & (!g3494)));
	assign g3496 = (((!g3493) & (g3495)));
	assign g3497 = (((!g2) & (!g8) & (g3404) & (g3490)) + ((!g2) & (g8) & (!g3404) & (g3490)) + ((!g2) & (g8) & (g3404) & (!g3490)) + ((!g2) & (g8) & (g3404) & (g3490)) + ((g2) & (!g8) & (!g3404) & (!g3490)) + ((g2) & (!g8) & (!g3404) & (g3490)) + ((g2) & (!g8) & (g3404) & (!g3490)) + ((g2) & (g8) & (!g3404) & (!g3490)));
	assign g3498 = (((!g3403) & (!g3493) & (!g3495) & (g3497)) + ((!g3403) & (g3493) & (!g3495) & (g3497)) + ((!g3403) & (g3493) & (g3495) & (g3497)) + ((g3403) & (!g3493) & (!g3495) & (!g3497)) + ((g3403) & (!g3493) & (g3495) & (!g3497)) + ((g3403) & (!g3493) & (g3495) & (g3497)) + ((g3403) & (g3493) & (!g3495) & (!g3497)) + ((g3403) & (g3493) & (g3495) & (!g3497)));
	assign g3499 = (((!g8) & (!g3404) & (g3490) & (!g3493) & (!g3495)) + ((!g8) & (!g3404) & (g3490) & (g3493) & (!g3495)) + ((!g8) & (!g3404) & (g3490) & (g3493) & (g3495)) + ((!g8) & (g3404) & (!g3490) & (!g3493) & (!g3495)) + ((!g8) & (g3404) & (!g3490) & (!g3493) & (g3495)) + ((!g8) & (g3404) & (!g3490) & (g3493) & (!g3495)) + ((!g8) & (g3404) & (!g3490) & (g3493) & (g3495)) + ((!g8) & (g3404) & (g3490) & (!g3493) & (g3495)) + ((g8) & (!g3404) & (!g3490) & (!g3493) & (!g3495)) + ((g8) & (!g3404) & (!g3490) & (g3493) & (!g3495)) + ((g8) & (!g3404) & (!g3490) & (g3493) & (g3495)) + ((g8) & (g3404) & (!g3490) & (!g3493) & (g3495)) + ((g8) & (g3404) & (g3490) & (!g3493) & (!g3495)) + ((g8) & (g3404) & (g3490) & (!g3493) & (g3495)) + ((g8) & (g3404) & (g3490) & (g3493) & (!g3495)) + ((g8) & (g3404) & (g3490) & (g3493) & (g3495)));
	assign g3500 = (((!g18) & (!g27) & (g3406) & (g3489)) + ((!g18) & (g27) & (!g3406) & (g3489)) + ((!g18) & (g27) & (g3406) & (!g3489)) + ((!g18) & (g27) & (g3406) & (g3489)) + ((g18) & (!g27) & (!g3406) & (!g3489)) + ((g18) & (!g27) & (!g3406) & (g3489)) + ((g18) & (!g27) & (g3406) & (!g3489)) + ((g18) & (g27) & (!g3406) & (!g3489)));
	assign g3501 = (((!g3405) & (!g3493) & (!g3495) & (g3500)) + ((!g3405) & (g3493) & (!g3495) & (g3500)) + ((!g3405) & (g3493) & (g3495) & (g3500)) + ((g3405) & (!g3493) & (!g3495) & (!g3500)) + ((g3405) & (!g3493) & (g3495) & (!g3500)) + ((g3405) & (!g3493) & (g3495) & (g3500)) + ((g3405) & (g3493) & (!g3495) & (!g3500)) + ((g3405) & (g3493) & (g3495) & (!g3500)));
	assign g3502 = (((!g27) & (!g3406) & (g3489) & (!g3493) & (!g3495)) + ((!g27) & (!g3406) & (g3489) & (g3493) & (!g3495)) + ((!g27) & (!g3406) & (g3489) & (g3493) & (g3495)) + ((!g27) & (g3406) & (!g3489) & (!g3493) & (!g3495)) + ((!g27) & (g3406) & (!g3489) & (!g3493) & (g3495)) + ((!g27) & (g3406) & (!g3489) & (g3493) & (!g3495)) + ((!g27) & (g3406) & (!g3489) & (g3493) & (g3495)) + ((!g27) & (g3406) & (g3489) & (!g3493) & (g3495)) + ((g27) & (!g3406) & (!g3489) & (!g3493) & (!g3495)) + ((g27) & (!g3406) & (!g3489) & (g3493) & (!g3495)) + ((g27) & (!g3406) & (!g3489) & (g3493) & (g3495)) + ((g27) & (g3406) & (!g3489) & (!g3493) & (g3495)) + ((g27) & (g3406) & (g3489) & (!g3493) & (!g3495)) + ((g27) & (g3406) & (g3489) & (!g3493) & (g3495)) + ((g27) & (g3406) & (g3489) & (g3493) & (!g3495)) + ((g27) & (g3406) & (g3489) & (g3493) & (g3495)));
	assign g3503 = (((!g39) & (!g54) & (g3408) & (g3488)) + ((!g39) & (g54) & (!g3408) & (g3488)) + ((!g39) & (g54) & (g3408) & (!g3488)) + ((!g39) & (g54) & (g3408) & (g3488)) + ((g39) & (!g54) & (!g3408) & (!g3488)) + ((g39) & (!g54) & (!g3408) & (g3488)) + ((g39) & (!g54) & (g3408) & (!g3488)) + ((g39) & (g54) & (!g3408) & (!g3488)));
	assign g3504 = (((!g3407) & (!g3493) & (!g3495) & (g3503)) + ((!g3407) & (g3493) & (!g3495) & (g3503)) + ((!g3407) & (g3493) & (g3495) & (g3503)) + ((g3407) & (!g3493) & (!g3495) & (!g3503)) + ((g3407) & (!g3493) & (g3495) & (!g3503)) + ((g3407) & (!g3493) & (g3495) & (g3503)) + ((g3407) & (g3493) & (!g3495) & (!g3503)) + ((g3407) & (g3493) & (g3495) & (!g3503)));
	assign g3505 = (((!g54) & (!g3408) & (g3488) & (!g3493) & (!g3495)) + ((!g54) & (!g3408) & (g3488) & (g3493) & (!g3495)) + ((!g54) & (!g3408) & (g3488) & (g3493) & (g3495)) + ((!g54) & (g3408) & (!g3488) & (!g3493) & (!g3495)) + ((!g54) & (g3408) & (!g3488) & (!g3493) & (g3495)) + ((!g54) & (g3408) & (!g3488) & (g3493) & (!g3495)) + ((!g54) & (g3408) & (!g3488) & (g3493) & (g3495)) + ((!g54) & (g3408) & (g3488) & (!g3493) & (g3495)) + ((g54) & (!g3408) & (!g3488) & (!g3493) & (!g3495)) + ((g54) & (!g3408) & (!g3488) & (g3493) & (!g3495)) + ((g54) & (!g3408) & (!g3488) & (g3493) & (g3495)) + ((g54) & (g3408) & (!g3488) & (!g3493) & (g3495)) + ((g54) & (g3408) & (g3488) & (!g3493) & (!g3495)) + ((g54) & (g3408) & (g3488) & (!g3493) & (g3495)) + ((g54) & (g3408) & (g3488) & (g3493) & (!g3495)) + ((g54) & (g3408) & (g3488) & (g3493) & (g3495)));
	assign g3506 = (((!g68) & (!g87) & (g3410) & (g3487)) + ((!g68) & (g87) & (!g3410) & (g3487)) + ((!g68) & (g87) & (g3410) & (!g3487)) + ((!g68) & (g87) & (g3410) & (g3487)) + ((g68) & (!g87) & (!g3410) & (!g3487)) + ((g68) & (!g87) & (!g3410) & (g3487)) + ((g68) & (!g87) & (g3410) & (!g3487)) + ((g68) & (g87) & (!g3410) & (!g3487)));
	assign g3507 = (((!g3409) & (!g3493) & (!g3495) & (g3506)) + ((!g3409) & (g3493) & (!g3495) & (g3506)) + ((!g3409) & (g3493) & (g3495) & (g3506)) + ((g3409) & (!g3493) & (!g3495) & (!g3506)) + ((g3409) & (!g3493) & (g3495) & (!g3506)) + ((g3409) & (!g3493) & (g3495) & (g3506)) + ((g3409) & (g3493) & (!g3495) & (!g3506)) + ((g3409) & (g3493) & (g3495) & (!g3506)));
	assign g3508 = (((!g87) & (!g3410) & (g3487) & (!g3493) & (!g3495)) + ((!g87) & (!g3410) & (g3487) & (g3493) & (!g3495)) + ((!g87) & (!g3410) & (g3487) & (g3493) & (g3495)) + ((!g87) & (g3410) & (!g3487) & (!g3493) & (!g3495)) + ((!g87) & (g3410) & (!g3487) & (!g3493) & (g3495)) + ((!g87) & (g3410) & (!g3487) & (g3493) & (!g3495)) + ((!g87) & (g3410) & (!g3487) & (g3493) & (g3495)) + ((!g87) & (g3410) & (g3487) & (!g3493) & (g3495)) + ((g87) & (!g3410) & (!g3487) & (!g3493) & (!g3495)) + ((g87) & (!g3410) & (!g3487) & (g3493) & (!g3495)) + ((g87) & (!g3410) & (!g3487) & (g3493) & (g3495)) + ((g87) & (g3410) & (!g3487) & (!g3493) & (g3495)) + ((g87) & (g3410) & (g3487) & (!g3493) & (!g3495)) + ((g87) & (g3410) & (g3487) & (!g3493) & (g3495)) + ((g87) & (g3410) & (g3487) & (g3493) & (!g3495)) + ((g87) & (g3410) & (g3487) & (g3493) & (g3495)));
	assign g3509 = (((!g104) & (!g127) & (g3412) & (g3486)) + ((!g104) & (g127) & (!g3412) & (g3486)) + ((!g104) & (g127) & (g3412) & (!g3486)) + ((!g104) & (g127) & (g3412) & (g3486)) + ((g104) & (!g127) & (!g3412) & (!g3486)) + ((g104) & (!g127) & (!g3412) & (g3486)) + ((g104) & (!g127) & (g3412) & (!g3486)) + ((g104) & (g127) & (!g3412) & (!g3486)));
	assign g3510 = (((!g3411) & (!g3493) & (!g3495) & (g3509)) + ((!g3411) & (g3493) & (!g3495) & (g3509)) + ((!g3411) & (g3493) & (g3495) & (g3509)) + ((g3411) & (!g3493) & (!g3495) & (!g3509)) + ((g3411) & (!g3493) & (g3495) & (!g3509)) + ((g3411) & (!g3493) & (g3495) & (g3509)) + ((g3411) & (g3493) & (!g3495) & (!g3509)) + ((g3411) & (g3493) & (g3495) & (!g3509)));
	assign g3511 = (((!g127) & (!g3412) & (g3486) & (!g3493) & (!g3495)) + ((!g127) & (!g3412) & (g3486) & (g3493) & (!g3495)) + ((!g127) & (!g3412) & (g3486) & (g3493) & (g3495)) + ((!g127) & (g3412) & (!g3486) & (!g3493) & (!g3495)) + ((!g127) & (g3412) & (!g3486) & (!g3493) & (g3495)) + ((!g127) & (g3412) & (!g3486) & (g3493) & (!g3495)) + ((!g127) & (g3412) & (!g3486) & (g3493) & (g3495)) + ((!g127) & (g3412) & (g3486) & (!g3493) & (g3495)) + ((g127) & (!g3412) & (!g3486) & (!g3493) & (!g3495)) + ((g127) & (!g3412) & (!g3486) & (g3493) & (!g3495)) + ((g127) & (!g3412) & (!g3486) & (g3493) & (g3495)) + ((g127) & (g3412) & (!g3486) & (!g3493) & (g3495)) + ((g127) & (g3412) & (g3486) & (!g3493) & (!g3495)) + ((g127) & (g3412) & (g3486) & (!g3493) & (g3495)) + ((g127) & (g3412) & (g3486) & (g3493) & (!g3495)) + ((g127) & (g3412) & (g3486) & (g3493) & (g3495)));
	assign g3512 = (((!g147) & (!g174) & (g3414) & (g3485)) + ((!g147) & (g174) & (!g3414) & (g3485)) + ((!g147) & (g174) & (g3414) & (!g3485)) + ((!g147) & (g174) & (g3414) & (g3485)) + ((g147) & (!g174) & (!g3414) & (!g3485)) + ((g147) & (!g174) & (!g3414) & (g3485)) + ((g147) & (!g174) & (g3414) & (!g3485)) + ((g147) & (g174) & (!g3414) & (!g3485)));
	assign g3513 = (((!g3413) & (!g3493) & (!g3495) & (g3512)) + ((!g3413) & (g3493) & (!g3495) & (g3512)) + ((!g3413) & (g3493) & (g3495) & (g3512)) + ((g3413) & (!g3493) & (!g3495) & (!g3512)) + ((g3413) & (!g3493) & (g3495) & (!g3512)) + ((g3413) & (!g3493) & (g3495) & (g3512)) + ((g3413) & (g3493) & (!g3495) & (!g3512)) + ((g3413) & (g3493) & (g3495) & (!g3512)));
	assign g3514 = (((!g174) & (!g3414) & (g3485) & (!g3493) & (!g3495)) + ((!g174) & (!g3414) & (g3485) & (g3493) & (!g3495)) + ((!g174) & (!g3414) & (g3485) & (g3493) & (g3495)) + ((!g174) & (g3414) & (!g3485) & (!g3493) & (!g3495)) + ((!g174) & (g3414) & (!g3485) & (!g3493) & (g3495)) + ((!g174) & (g3414) & (!g3485) & (g3493) & (!g3495)) + ((!g174) & (g3414) & (!g3485) & (g3493) & (g3495)) + ((!g174) & (g3414) & (g3485) & (!g3493) & (g3495)) + ((g174) & (!g3414) & (!g3485) & (!g3493) & (!g3495)) + ((g174) & (!g3414) & (!g3485) & (g3493) & (!g3495)) + ((g174) & (!g3414) & (!g3485) & (g3493) & (g3495)) + ((g174) & (g3414) & (!g3485) & (!g3493) & (g3495)) + ((g174) & (g3414) & (g3485) & (!g3493) & (!g3495)) + ((g174) & (g3414) & (g3485) & (!g3493) & (g3495)) + ((g174) & (g3414) & (g3485) & (g3493) & (!g3495)) + ((g174) & (g3414) & (g3485) & (g3493) & (g3495)));
	assign g3515 = (((!g198) & (!g229) & (g3416) & (g3484)) + ((!g198) & (g229) & (!g3416) & (g3484)) + ((!g198) & (g229) & (g3416) & (!g3484)) + ((!g198) & (g229) & (g3416) & (g3484)) + ((g198) & (!g229) & (!g3416) & (!g3484)) + ((g198) & (!g229) & (!g3416) & (g3484)) + ((g198) & (!g229) & (g3416) & (!g3484)) + ((g198) & (g229) & (!g3416) & (!g3484)));
	assign g3516 = (((!g3415) & (!g3493) & (!g3495) & (g3515)) + ((!g3415) & (g3493) & (!g3495) & (g3515)) + ((!g3415) & (g3493) & (g3495) & (g3515)) + ((g3415) & (!g3493) & (!g3495) & (!g3515)) + ((g3415) & (!g3493) & (g3495) & (!g3515)) + ((g3415) & (!g3493) & (g3495) & (g3515)) + ((g3415) & (g3493) & (!g3495) & (!g3515)) + ((g3415) & (g3493) & (g3495) & (!g3515)));
	assign g3517 = (((!g229) & (!g3416) & (g3484) & (!g3493) & (!g3495)) + ((!g229) & (!g3416) & (g3484) & (g3493) & (!g3495)) + ((!g229) & (!g3416) & (g3484) & (g3493) & (g3495)) + ((!g229) & (g3416) & (!g3484) & (!g3493) & (!g3495)) + ((!g229) & (g3416) & (!g3484) & (!g3493) & (g3495)) + ((!g229) & (g3416) & (!g3484) & (g3493) & (!g3495)) + ((!g229) & (g3416) & (!g3484) & (g3493) & (g3495)) + ((!g229) & (g3416) & (g3484) & (!g3493) & (g3495)) + ((g229) & (!g3416) & (!g3484) & (!g3493) & (!g3495)) + ((g229) & (!g3416) & (!g3484) & (g3493) & (!g3495)) + ((g229) & (!g3416) & (!g3484) & (g3493) & (g3495)) + ((g229) & (g3416) & (!g3484) & (!g3493) & (g3495)) + ((g229) & (g3416) & (g3484) & (!g3493) & (!g3495)) + ((g229) & (g3416) & (g3484) & (!g3493) & (g3495)) + ((g229) & (g3416) & (g3484) & (g3493) & (!g3495)) + ((g229) & (g3416) & (g3484) & (g3493) & (g3495)));
	assign g3518 = (((!g255) & (!g290) & (g3418) & (g3483)) + ((!g255) & (g290) & (!g3418) & (g3483)) + ((!g255) & (g290) & (g3418) & (!g3483)) + ((!g255) & (g290) & (g3418) & (g3483)) + ((g255) & (!g290) & (!g3418) & (!g3483)) + ((g255) & (!g290) & (!g3418) & (g3483)) + ((g255) & (!g290) & (g3418) & (!g3483)) + ((g255) & (g290) & (!g3418) & (!g3483)));
	assign g3519 = (((!g3417) & (!g3493) & (!g3495) & (g3518)) + ((!g3417) & (g3493) & (!g3495) & (g3518)) + ((!g3417) & (g3493) & (g3495) & (g3518)) + ((g3417) & (!g3493) & (!g3495) & (!g3518)) + ((g3417) & (!g3493) & (g3495) & (!g3518)) + ((g3417) & (!g3493) & (g3495) & (g3518)) + ((g3417) & (g3493) & (!g3495) & (!g3518)) + ((g3417) & (g3493) & (g3495) & (!g3518)));
	assign g3520 = (((!g290) & (!g3418) & (g3483) & (!g3493) & (!g3495)) + ((!g290) & (!g3418) & (g3483) & (g3493) & (!g3495)) + ((!g290) & (!g3418) & (g3483) & (g3493) & (g3495)) + ((!g290) & (g3418) & (!g3483) & (!g3493) & (!g3495)) + ((!g290) & (g3418) & (!g3483) & (!g3493) & (g3495)) + ((!g290) & (g3418) & (!g3483) & (g3493) & (!g3495)) + ((!g290) & (g3418) & (!g3483) & (g3493) & (g3495)) + ((!g290) & (g3418) & (g3483) & (!g3493) & (g3495)) + ((g290) & (!g3418) & (!g3483) & (!g3493) & (!g3495)) + ((g290) & (!g3418) & (!g3483) & (g3493) & (!g3495)) + ((g290) & (!g3418) & (!g3483) & (g3493) & (g3495)) + ((g290) & (g3418) & (!g3483) & (!g3493) & (g3495)) + ((g290) & (g3418) & (g3483) & (!g3493) & (!g3495)) + ((g290) & (g3418) & (g3483) & (!g3493) & (g3495)) + ((g290) & (g3418) & (g3483) & (g3493) & (!g3495)) + ((g290) & (g3418) & (g3483) & (g3493) & (g3495)));
	assign g3521 = (((!g319) & (!g358) & (g3420) & (g3482)) + ((!g319) & (g358) & (!g3420) & (g3482)) + ((!g319) & (g358) & (g3420) & (!g3482)) + ((!g319) & (g358) & (g3420) & (g3482)) + ((g319) & (!g358) & (!g3420) & (!g3482)) + ((g319) & (!g358) & (!g3420) & (g3482)) + ((g319) & (!g358) & (g3420) & (!g3482)) + ((g319) & (g358) & (!g3420) & (!g3482)));
	assign g3522 = (((!g3419) & (!g3493) & (!g3495) & (g3521)) + ((!g3419) & (g3493) & (!g3495) & (g3521)) + ((!g3419) & (g3493) & (g3495) & (g3521)) + ((g3419) & (!g3493) & (!g3495) & (!g3521)) + ((g3419) & (!g3493) & (g3495) & (!g3521)) + ((g3419) & (!g3493) & (g3495) & (g3521)) + ((g3419) & (g3493) & (!g3495) & (!g3521)) + ((g3419) & (g3493) & (g3495) & (!g3521)));
	assign g3523 = (((!g358) & (!g3420) & (g3482) & (!g3493) & (!g3495)) + ((!g358) & (!g3420) & (g3482) & (g3493) & (!g3495)) + ((!g358) & (!g3420) & (g3482) & (g3493) & (g3495)) + ((!g358) & (g3420) & (!g3482) & (!g3493) & (!g3495)) + ((!g358) & (g3420) & (!g3482) & (!g3493) & (g3495)) + ((!g358) & (g3420) & (!g3482) & (g3493) & (!g3495)) + ((!g358) & (g3420) & (!g3482) & (g3493) & (g3495)) + ((!g358) & (g3420) & (g3482) & (!g3493) & (g3495)) + ((g358) & (!g3420) & (!g3482) & (!g3493) & (!g3495)) + ((g358) & (!g3420) & (!g3482) & (g3493) & (!g3495)) + ((g358) & (!g3420) & (!g3482) & (g3493) & (g3495)) + ((g358) & (g3420) & (!g3482) & (!g3493) & (g3495)) + ((g358) & (g3420) & (g3482) & (!g3493) & (!g3495)) + ((g358) & (g3420) & (g3482) & (!g3493) & (g3495)) + ((g358) & (g3420) & (g3482) & (g3493) & (!g3495)) + ((g358) & (g3420) & (g3482) & (g3493) & (g3495)));
	assign g3524 = (((!g390) & (!g433) & (g3422) & (g3481)) + ((!g390) & (g433) & (!g3422) & (g3481)) + ((!g390) & (g433) & (g3422) & (!g3481)) + ((!g390) & (g433) & (g3422) & (g3481)) + ((g390) & (!g433) & (!g3422) & (!g3481)) + ((g390) & (!g433) & (!g3422) & (g3481)) + ((g390) & (!g433) & (g3422) & (!g3481)) + ((g390) & (g433) & (!g3422) & (!g3481)));
	assign g3525 = (((!g3421) & (!g3493) & (!g3495) & (g3524)) + ((!g3421) & (g3493) & (!g3495) & (g3524)) + ((!g3421) & (g3493) & (g3495) & (g3524)) + ((g3421) & (!g3493) & (!g3495) & (!g3524)) + ((g3421) & (!g3493) & (g3495) & (!g3524)) + ((g3421) & (!g3493) & (g3495) & (g3524)) + ((g3421) & (g3493) & (!g3495) & (!g3524)) + ((g3421) & (g3493) & (g3495) & (!g3524)));
	assign g3526 = (((!g433) & (!g3422) & (g3481) & (!g3493) & (!g3495)) + ((!g433) & (!g3422) & (g3481) & (g3493) & (!g3495)) + ((!g433) & (!g3422) & (g3481) & (g3493) & (g3495)) + ((!g433) & (g3422) & (!g3481) & (!g3493) & (!g3495)) + ((!g433) & (g3422) & (!g3481) & (!g3493) & (g3495)) + ((!g433) & (g3422) & (!g3481) & (g3493) & (!g3495)) + ((!g433) & (g3422) & (!g3481) & (g3493) & (g3495)) + ((!g433) & (g3422) & (g3481) & (!g3493) & (g3495)) + ((g433) & (!g3422) & (!g3481) & (!g3493) & (!g3495)) + ((g433) & (!g3422) & (!g3481) & (g3493) & (!g3495)) + ((g433) & (!g3422) & (!g3481) & (g3493) & (g3495)) + ((g433) & (g3422) & (!g3481) & (!g3493) & (g3495)) + ((g433) & (g3422) & (g3481) & (!g3493) & (!g3495)) + ((g433) & (g3422) & (g3481) & (!g3493) & (g3495)) + ((g433) & (g3422) & (g3481) & (g3493) & (!g3495)) + ((g433) & (g3422) & (g3481) & (g3493) & (g3495)));
	assign g3527 = (((!g468) & (!g515) & (g3424) & (g3480)) + ((!g468) & (g515) & (!g3424) & (g3480)) + ((!g468) & (g515) & (g3424) & (!g3480)) + ((!g468) & (g515) & (g3424) & (g3480)) + ((g468) & (!g515) & (!g3424) & (!g3480)) + ((g468) & (!g515) & (!g3424) & (g3480)) + ((g468) & (!g515) & (g3424) & (!g3480)) + ((g468) & (g515) & (!g3424) & (!g3480)));
	assign g3528 = (((!g3423) & (!g3493) & (!g3495) & (g3527)) + ((!g3423) & (g3493) & (!g3495) & (g3527)) + ((!g3423) & (g3493) & (g3495) & (g3527)) + ((g3423) & (!g3493) & (!g3495) & (!g3527)) + ((g3423) & (!g3493) & (g3495) & (!g3527)) + ((g3423) & (!g3493) & (g3495) & (g3527)) + ((g3423) & (g3493) & (!g3495) & (!g3527)) + ((g3423) & (g3493) & (g3495) & (!g3527)));
	assign g3529 = (((!g515) & (!g3424) & (g3480) & (!g3493) & (!g3495)) + ((!g515) & (!g3424) & (g3480) & (g3493) & (!g3495)) + ((!g515) & (!g3424) & (g3480) & (g3493) & (g3495)) + ((!g515) & (g3424) & (!g3480) & (!g3493) & (!g3495)) + ((!g515) & (g3424) & (!g3480) & (!g3493) & (g3495)) + ((!g515) & (g3424) & (!g3480) & (g3493) & (!g3495)) + ((!g515) & (g3424) & (!g3480) & (g3493) & (g3495)) + ((!g515) & (g3424) & (g3480) & (!g3493) & (g3495)) + ((g515) & (!g3424) & (!g3480) & (!g3493) & (!g3495)) + ((g515) & (!g3424) & (!g3480) & (g3493) & (!g3495)) + ((g515) & (!g3424) & (!g3480) & (g3493) & (g3495)) + ((g515) & (g3424) & (!g3480) & (!g3493) & (g3495)) + ((g515) & (g3424) & (g3480) & (!g3493) & (!g3495)) + ((g515) & (g3424) & (g3480) & (!g3493) & (g3495)) + ((g515) & (g3424) & (g3480) & (g3493) & (!g3495)) + ((g515) & (g3424) & (g3480) & (g3493) & (g3495)));
	assign g3530 = (((!g553) & (!g604) & (g3426) & (g3479)) + ((!g553) & (g604) & (!g3426) & (g3479)) + ((!g553) & (g604) & (g3426) & (!g3479)) + ((!g553) & (g604) & (g3426) & (g3479)) + ((g553) & (!g604) & (!g3426) & (!g3479)) + ((g553) & (!g604) & (!g3426) & (g3479)) + ((g553) & (!g604) & (g3426) & (!g3479)) + ((g553) & (g604) & (!g3426) & (!g3479)));
	assign g3531 = (((!g3425) & (!g3493) & (!g3495) & (g3530)) + ((!g3425) & (g3493) & (!g3495) & (g3530)) + ((!g3425) & (g3493) & (g3495) & (g3530)) + ((g3425) & (!g3493) & (!g3495) & (!g3530)) + ((g3425) & (!g3493) & (g3495) & (!g3530)) + ((g3425) & (!g3493) & (g3495) & (g3530)) + ((g3425) & (g3493) & (!g3495) & (!g3530)) + ((g3425) & (g3493) & (g3495) & (!g3530)));
	assign g3532 = (((!g604) & (!g3426) & (g3479) & (!g3493) & (!g3495)) + ((!g604) & (!g3426) & (g3479) & (g3493) & (!g3495)) + ((!g604) & (!g3426) & (g3479) & (g3493) & (g3495)) + ((!g604) & (g3426) & (!g3479) & (!g3493) & (!g3495)) + ((!g604) & (g3426) & (!g3479) & (!g3493) & (g3495)) + ((!g604) & (g3426) & (!g3479) & (g3493) & (!g3495)) + ((!g604) & (g3426) & (!g3479) & (g3493) & (g3495)) + ((!g604) & (g3426) & (g3479) & (!g3493) & (g3495)) + ((g604) & (!g3426) & (!g3479) & (!g3493) & (!g3495)) + ((g604) & (!g3426) & (!g3479) & (g3493) & (!g3495)) + ((g604) & (!g3426) & (!g3479) & (g3493) & (g3495)) + ((g604) & (g3426) & (!g3479) & (!g3493) & (g3495)) + ((g604) & (g3426) & (g3479) & (!g3493) & (!g3495)) + ((g604) & (g3426) & (g3479) & (!g3493) & (g3495)) + ((g604) & (g3426) & (g3479) & (g3493) & (!g3495)) + ((g604) & (g3426) & (g3479) & (g3493) & (g3495)));
	assign g3533 = (((!g645) & (!g700) & (g3428) & (g3478)) + ((!g645) & (g700) & (!g3428) & (g3478)) + ((!g645) & (g700) & (g3428) & (!g3478)) + ((!g645) & (g700) & (g3428) & (g3478)) + ((g645) & (!g700) & (!g3428) & (!g3478)) + ((g645) & (!g700) & (!g3428) & (g3478)) + ((g645) & (!g700) & (g3428) & (!g3478)) + ((g645) & (g700) & (!g3428) & (!g3478)));
	assign g3534 = (((!g3427) & (!g3493) & (!g3495) & (g3533)) + ((!g3427) & (g3493) & (!g3495) & (g3533)) + ((!g3427) & (g3493) & (g3495) & (g3533)) + ((g3427) & (!g3493) & (!g3495) & (!g3533)) + ((g3427) & (!g3493) & (g3495) & (!g3533)) + ((g3427) & (!g3493) & (g3495) & (g3533)) + ((g3427) & (g3493) & (!g3495) & (!g3533)) + ((g3427) & (g3493) & (g3495) & (!g3533)));
	assign g3535 = (((!g700) & (!g3428) & (g3478) & (!g3493) & (!g3495)) + ((!g700) & (!g3428) & (g3478) & (g3493) & (!g3495)) + ((!g700) & (!g3428) & (g3478) & (g3493) & (g3495)) + ((!g700) & (g3428) & (!g3478) & (!g3493) & (!g3495)) + ((!g700) & (g3428) & (!g3478) & (!g3493) & (g3495)) + ((!g700) & (g3428) & (!g3478) & (g3493) & (!g3495)) + ((!g700) & (g3428) & (!g3478) & (g3493) & (g3495)) + ((!g700) & (g3428) & (g3478) & (!g3493) & (g3495)) + ((g700) & (!g3428) & (!g3478) & (!g3493) & (!g3495)) + ((g700) & (!g3428) & (!g3478) & (g3493) & (!g3495)) + ((g700) & (!g3428) & (!g3478) & (g3493) & (g3495)) + ((g700) & (g3428) & (!g3478) & (!g3493) & (g3495)) + ((g700) & (g3428) & (g3478) & (!g3493) & (!g3495)) + ((g700) & (g3428) & (g3478) & (!g3493) & (g3495)) + ((g700) & (g3428) & (g3478) & (g3493) & (!g3495)) + ((g700) & (g3428) & (g3478) & (g3493) & (g3495)));
	assign g3536 = (((!g744) & (!g803) & (g3430) & (g3477)) + ((!g744) & (g803) & (!g3430) & (g3477)) + ((!g744) & (g803) & (g3430) & (!g3477)) + ((!g744) & (g803) & (g3430) & (g3477)) + ((g744) & (!g803) & (!g3430) & (!g3477)) + ((g744) & (!g803) & (!g3430) & (g3477)) + ((g744) & (!g803) & (g3430) & (!g3477)) + ((g744) & (g803) & (!g3430) & (!g3477)));
	assign g3537 = (((!g3429) & (!g3493) & (!g3495) & (g3536)) + ((!g3429) & (g3493) & (!g3495) & (g3536)) + ((!g3429) & (g3493) & (g3495) & (g3536)) + ((g3429) & (!g3493) & (!g3495) & (!g3536)) + ((g3429) & (!g3493) & (g3495) & (!g3536)) + ((g3429) & (!g3493) & (g3495) & (g3536)) + ((g3429) & (g3493) & (!g3495) & (!g3536)) + ((g3429) & (g3493) & (g3495) & (!g3536)));
	assign g3538 = (((!g803) & (!g3430) & (g3477) & (!g3493) & (!g3495)) + ((!g803) & (!g3430) & (g3477) & (g3493) & (!g3495)) + ((!g803) & (!g3430) & (g3477) & (g3493) & (g3495)) + ((!g803) & (g3430) & (!g3477) & (!g3493) & (!g3495)) + ((!g803) & (g3430) & (!g3477) & (!g3493) & (g3495)) + ((!g803) & (g3430) & (!g3477) & (g3493) & (!g3495)) + ((!g803) & (g3430) & (!g3477) & (g3493) & (g3495)) + ((!g803) & (g3430) & (g3477) & (!g3493) & (g3495)) + ((g803) & (!g3430) & (!g3477) & (!g3493) & (!g3495)) + ((g803) & (!g3430) & (!g3477) & (g3493) & (!g3495)) + ((g803) & (!g3430) & (!g3477) & (g3493) & (g3495)) + ((g803) & (g3430) & (!g3477) & (!g3493) & (g3495)) + ((g803) & (g3430) & (g3477) & (!g3493) & (!g3495)) + ((g803) & (g3430) & (g3477) & (!g3493) & (g3495)) + ((g803) & (g3430) & (g3477) & (g3493) & (!g3495)) + ((g803) & (g3430) & (g3477) & (g3493) & (g3495)));
	assign g3539 = (((!g851) & (!g914) & (g3432) & (g3476)) + ((!g851) & (g914) & (!g3432) & (g3476)) + ((!g851) & (g914) & (g3432) & (!g3476)) + ((!g851) & (g914) & (g3432) & (g3476)) + ((g851) & (!g914) & (!g3432) & (!g3476)) + ((g851) & (!g914) & (!g3432) & (g3476)) + ((g851) & (!g914) & (g3432) & (!g3476)) + ((g851) & (g914) & (!g3432) & (!g3476)));
	assign g3540 = (((!g3431) & (!g3493) & (!g3495) & (g3539)) + ((!g3431) & (g3493) & (!g3495) & (g3539)) + ((!g3431) & (g3493) & (g3495) & (g3539)) + ((g3431) & (!g3493) & (!g3495) & (!g3539)) + ((g3431) & (!g3493) & (g3495) & (!g3539)) + ((g3431) & (!g3493) & (g3495) & (g3539)) + ((g3431) & (g3493) & (!g3495) & (!g3539)) + ((g3431) & (g3493) & (g3495) & (!g3539)));
	assign g3541 = (((!g914) & (!g3432) & (g3476) & (!g3493) & (!g3495)) + ((!g914) & (!g3432) & (g3476) & (g3493) & (!g3495)) + ((!g914) & (!g3432) & (g3476) & (g3493) & (g3495)) + ((!g914) & (g3432) & (!g3476) & (!g3493) & (!g3495)) + ((!g914) & (g3432) & (!g3476) & (!g3493) & (g3495)) + ((!g914) & (g3432) & (!g3476) & (g3493) & (!g3495)) + ((!g914) & (g3432) & (!g3476) & (g3493) & (g3495)) + ((!g914) & (g3432) & (g3476) & (!g3493) & (g3495)) + ((g914) & (!g3432) & (!g3476) & (!g3493) & (!g3495)) + ((g914) & (!g3432) & (!g3476) & (g3493) & (!g3495)) + ((g914) & (!g3432) & (!g3476) & (g3493) & (g3495)) + ((g914) & (g3432) & (!g3476) & (!g3493) & (g3495)) + ((g914) & (g3432) & (g3476) & (!g3493) & (!g3495)) + ((g914) & (g3432) & (g3476) & (!g3493) & (g3495)) + ((g914) & (g3432) & (g3476) & (g3493) & (!g3495)) + ((g914) & (g3432) & (g3476) & (g3493) & (g3495)));
	assign g3542 = (((!g1032) & (!g1030) & (g3434) & (g3475)) + ((!g1032) & (g1030) & (!g3434) & (g3475)) + ((!g1032) & (g1030) & (g3434) & (!g3475)) + ((!g1032) & (g1030) & (g3434) & (g3475)) + ((g1032) & (!g1030) & (!g3434) & (!g3475)) + ((g1032) & (!g1030) & (!g3434) & (g3475)) + ((g1032) & (!g1030) & (g3434) & (!g3475)) + ((g1032) & (g1030) & (!g3434) & (!g3475)));
	assign g3543 = (((!g3433) & (!g3493) & (!g3495) & (g3542)) + ((!g3433) & (g3493) & (!g3495) & (g3542)) + ((!g3433) & (g3493) & (g3495) & (g3542)) + ((g3433) & (!g3493) & (!g3495) & (!g3542)) + ((g3433) & (!g3493) & (g3495) & (!g3542)) + ((g3433) & (!g3493) & (g3495) & (g3542)) + ((g3433) & (g3493) & (!g3495) & (!g3542)) + ((g3433) & (g3493) & (g3495) & (!g3542)));
	assign g3544 = (((!g1030) & (!g3434) & (g3475) & (!g3493) & (!g3495)) + ((!g1030) & (!g3434) & (g3475) & (g3493) & (!g3495)) + ((!g1030) & (!g3434) & (g3475) & (g3493) & (g3495)) + ((!g1030) & (g3434) & (!g3475) & (!g3493) & (!g3495)) + ((!g1030) & (g3434) & (!g3475) & (!g3493) & (g3495)) + ((!g1030) & (g3434) & (!g3475) & (g3493) & (!g3495)) + ((!g1030) & (g3434) & (!g3475) & (g3493) & (g3495)) + ((!g1030) & (g3434) & (g3475) & (!g3493) & (g3495)) + ((g1030) & (!g3434) & (!g3475) & (!g3493) & (!g3495)) + ((g1030) & (!g3434) & (!g3475) & (g3493) & (!g3495)) + ((g1030) & (!g3434) & (!g3475) & (g3493) & (g3495)) + ((g1030) & (g3434) & (!g3475) & (!g3493) & (g3495)) + ((g1030) & (g3434) & (g3475) & (!g3493) & (!g3495)) + ((g1030) & (g3434) & (g3475) & (!g3493) & (g3495)) + ((g1030) & (g3434) & (g3475) & (g3493) & (!g3495)) + ((g1030) & (g3434) & (g3475) & (g3493) & (g3495)));
	assign g3545 = (((!g1160) & (!g1154) & (g3436) & (g3474)) + ((!g1160) & (g1154) & (!g3436) & (g3474)) + ((!g1160) & (g1154) & (g3436) & (!g3474)) + ((!g1160) & (g1154) & (g3436) & (g3474)) + ((g1160) & (!g1154) & (!g3436) & (!g3474)) + ((g1160) & (!g1154) & (!g3436) & (g3474)) + ((g1160) & (!g1154) & (g3436) & (!g3474)) + ((g1160) & (g1154) & (!g3436) & (!g3474)));
	assign g3546 = (((!g3435) & (!g3493) & (!g3495) & (g3545)) + ((!g3435) & (g3493) & (!g3495) & (g3545)) + ((!g3435) & (g3493) & (g3495) & (g3545)) + ((g3435) & (!g3493) & (!g3495) & (!g3545)) + ((g3435) & (!g3493) & (g3495) & (!g3545)) + ((g3435) & (!g3493) & (g3495) & (g3545)) + ((g3435) & (g3493) & (!g3495) & (!g3545)) + ((g3435) & (g3493) & (g3495) & (!g3545)));
	assign g3547 = (((!g1154) & (!g3436) & (g3474) & (!g3493) & (!g3495)) + ((!g1154) & (!g3436) & (g3474) & (g3493) & (!g3495)) + ((!g1154) & (!g3436) & (g3474) & (g3493) & (g3495)) + ((!g1154) & (g3436) & (!g3474) & (!g3493) & (!g3495)) + ((!g1154) & (g3436) & (!g3474) & (!g3493) & (g3495)) + ((!g1154) & (g3436) & (!g3474) & (g3493) & (!g3495)) + ((!g1154) & (g3436) & (!g3474) & (g3493) & (g3495)) + ((!g1154) & (g3436) & (g3474) & (!g3493) & (g3495)) + ((g1154) & (!g3436) & (!g3474) & (!g3493) & (!g3495)) + ((g1154) & (!g3436) & (!g3474) & (g3493) & (!g3495)) + ((g1154) & (!g3436) & (!g3474) & (g3493) & (g3495)) + ((g1154) & (g3436) & (!g3474) & (!g3493) & (g3495)) + ((g1154) & (g3436) & (g3474) & (!g3493) & (!g3495)) + ((g1154) & (g3436) & (g3474) & (!g3493) & (g3495)) + ((g1154) & (g3436) & (g3474) & (g3493) & (!g3495)) + ((g1154) & (g3436) & (g3474) & (g3493) & (g3495)));
	assign g3548 = (((!g1295) & (!g1285) & (g3438) & (g3473)) + ((!g1295) & (g1285) & (!g3438) & (g3473)) + ((!g1295) & (g1285) & (g3438) & (!g3473)) + ((!g1295) & (g1285) & (g3438) & (g3473)) + ((g1295) & (!g1285) & (!g3438) & (!g3473)) + ((g1295) & (!g1285) & (!g3438) & (g3473)) + ((g1295) & (!g1285) & (g3438) & (!g3473)) + ((g1295) & (g1285) & (!g3438) & (!g3473)));
	assign g3549 = (((!g3437) & (!g3493) & (!g3495) & (g3548)) + ((!g3437) & (g3493) & (!g3495) & (g3548)) + ((!g3437) & (g3493) & (g3495) & (g3548)) + ((g3437) & (!g3493) & (!g3495) & (!g3548)) + ((g3437) & (!g3493) & (g3495) & (!g3548)) + ((g3437) & (!g3493) & (g3495) & (g3548)) + ((g3437) & (g3493) & (!g3495) & (!g3548)) + ((g3437) & (g3493) & (g3495) & (!g3548)));
	assign g3550 = (((!g1285) & (!g3438) & (g3473) & (!g3493) & (!g3495)) + ((!g1285) & (!g3438) & (g3473) & (g3493) & (!g3495)) + ((!g1285) & (!g3438) & (g3473) & (g3493) & (g3495)) + ((!g1285) & (g3438) & (!g3473) & (!g3493) & (!g3495)) + ((!g1285) & (g3438) & (!g3473) & (!g3493) & (g3495)) + ((!g1285) & (g3438) & (!g3473) & (g3493) & (!g3495)) + ((!g1285) & (g3438) & (!g3473) & (g3493) & (g3495)) + ((!g1285) & (g3438) & (g3473) & (!g3493) & (g3495)) + ((g1285) & (!g3438) & (!g3473) & (!g3493) & (!g3495)) + ((g1285) & (!g3438) & (!g3473) & (g3493) & (!g3495)) + ((g1285) & (!g3438) & (!g3473) & (g3493) & (g3495)) + ((g1285) & (g3438) & (!g3473) & (!g3493) & (g3495)) + ((g1285) & (g3438) & (g3473) & (!g3493) & (!g3495)) + ((g1285) & (g3438) & (g3473) & (!g3493) & (g3495)) + ((g1285) & (g3438) & (g3473) & (g3493) & (!g3495)) + ((g1285) & (g3438) & (g3473) & (g3493) & (g3495)));
	assign g3551 = (((!g1437) & (!g1423) & (g3440) & (g3472)) + ((!g1437) & (g1423) & (!g3440) & (g3472)) + ((!g1437) & (g1423) & (g3440) & (!g3472)) + ((!g1437) & (g1423) & (g3440) & (g3472)) + ((g1437) & (!g1423) & (!g3440) & (!g3472)) + ((g1437) & (!g1423) & (!g3440) & (g3472)) + ((g1437) & (!g1423) & (g3440) & (!g3472)) + ((g1437) & (g1423) & (!g3440) & (!g3472)));
	assign g3552 = (((!g3439) & (!g3493) & (!g3495) & (g3551)) + ((!g3439) & (g3493) & (!g3495) & (g3551)) + ((!g3439) & (g3493) & (g3495) & (g3551)) + ((g3439) & (!g3493) & (!g3495) & (!g3551)) + ((g3439) & (!g3493) & (g3495) & (!g3551)) + ((g3439) & (!g3493) & (g3495) & (g3551)) + ((g3439) & (g3493) & (!g3495) & (!g3551)) + ((g3439) & (g3493) & (g3495) & (!g3551)));
	assign g3553 = (((!g1423) & (!g3440) & (g3472) & (!g3493) & (!g3495)) + ((!g1423) & (!g3440) & (g3472) & (g3493) & (!g3495)) + ((!g1423) & (!g3440) & (g3472) & (g3493) & (g3495)) + ((!g1423) & (g3440) & (!g3472) & (!g3493) & (!g3495)) + ((!g1423) & (g3440) & (!g3472) & (!g3493) & (g3495)) + ((!g1423) & (g3440) & (!g3472) & (g3493) & (!g3495)) + ((!g1423) & (g3440) & (!g3472) & (g3493) & (g3495)) + ((!g1423) & (g3440) & (g3472) & (!g3493) & (g3495)) + ((g1423) & (!g3440) & (!g3472) & (!g3493) & (!g3495)) + ((g1423) & (!g3440) & (!g3472) & (g3493) & (!g3495)) + ((g1423) & (!g3440) & (!g3472) & (g3493) & (g3495)) + ((g1423) & (g3440) & (!g3472) & (!g3493) & (g3495)) + ((g1423) & (g3440) & (g3472) & (!g3493) & (!g3495)) + ((g1423) & (g3440) & (g3472) & (!g3493) & (g3495)) + ((g1423) & (g3440) & (g3472) & (g3493) & (!g3495)) + ((g1423) & (g3440) & (g3472) & (g3493) & (g3495)));
	assign g3554 = (((!g1586) & (!g1568) & (g3442) & (g3471)) + ((!g1586) & (g1568) & (!g3442) & (g3471)) + ((!g1586) & (g1568) & (g3442) & (!g3471)) + ((!g1586) & (g1568) & (g3442) & (g3471)) + ((g1586) & (!g1568) & (!g3442) & (!g3471)) + ((g1586) & (!g1568) & (!g3442) & (g3471)) + ((g1586) & (!g1568) & (g3442) & (!g3471)) + ((g1586) & (g1568) & (!g3442) & (!g3471)));
	assign g3555 = (((!g3441) & (!g3493) & (!g3495) & (g3554)) + ((!g3441) & (g3493) & (!g3495) & (g3554)) + ((!g3441) & (g3493) & (g3495) & (g3554)) + ((g3441) & (!g3493) & (!g3495) & (!g3554)) + ((g3441) & (!g3493) & (g3495) & (!g3554)) + ((g3441) & (!g3493) & (g3495) & (g3554)) + ((g3441) & (g3493) & (!g3495) & (!g3554)) + ((g3441) & (g3493) & (g3495) & (!g3554)));
	assign g3556 = (((!g1568) & (!g3442) & (g3471) & (!g3493) & (!g3495)) + ((!g1568) & (!g3442) & (g3471) & (g3493) & (!g3495)) + ((!g1568) & (!g3442) & (g3471) & (g3493) & (g3495)) + ((!g1568) & (g3442) & (!g3471) & (!g3493) & (!g3495)) + ((!g1568) & (g3442) & (!g3471) & (!g3493) & (g3495)) + ((!g1568) & (g3442) & (!g3471) & (g3493) & (!g3495)) + ((!g1568) & (g3442) & (!g3471) & (g3493) & (g3495)) + ((!g1568) & (g3442) & (g3471) & (!g3493) & (g3495)) + ((g1568) & (!g3442) & (!g3471) & (!g3493) & (!g3495)) + ((g1568) & (!g3442) & (!g3471) & (g3493) & (!g3495)) + ((g1568) & (!g3442) & (!g3471) & (g3493) & (g3495)) + ((g1568) & (g3442) & (!g3471) & (!g3493) & (g3495)) + ((g1568) & (g3442) & (g3471) & (!g3493) & (!g3495)) + ((g1568) & (g3442) & (g3471) & (!g3493) & (g3495)) + ((g1568) & (g3442) & (g3471) & (g3493) & (!g3495)) + ((g1568) & (g3442) & (g3471) & (g3493) & (g3495)));
	assign g3557 = (((!g1742) & (!g1720) & (g3444) & (g3470)) + ((!g1742) & (g1720) & (!g3444) & (g3470)) + ((!g1742) & (g1720) & (g3444) & (!g3470)) + ((!g1742) & (g1720) & (g3444) & (g3470)) + ((g1742) & (!g1720) & (!g3444) & (!g3470)) + ((g1742) & (!g1720) & (!g3444) & (g3470)) + ((g1742) & (!g1720) & (g3444) & (!g3470)) + ((g1742) & (g1720) & (!g3444) & (!g3470)));
	assign g3558 = (((!g3443) & (!g3493) & (!g3495) & (g3557)) + ((!g3443) & (g3493) & (!g3495) & (g3557)) + ((!g3443) & (g3493) & (g3495) & (g3557)) + ((g3443) & (!g3493) & (!g3495) & (!g3557)) + ((g3443) & (!g3493) & (g3495) & (!g3557)) + ((g3443) & (!g3493) & (g3495) & (g3557)) + ((g3443) & (g3493) & (!g3495) & (!g3557)) + ((g3443) & (g3493) & (g3495) & (!g3557)));
	assign g3559 = (((!g1720) & (!g3444) & (g3470) & (!g3493) & (!g3495)) + ((!g1720) & (!g3444) & (g3470) & (g3493) & (!g3495)) + ((!g1720) & (!g3444) & (g3470) & (g3493) & (g3495)) + ((!g1720) & (g3444) & (!g3470) & (!g3493) & (!g3495)) + ((!g1720) & (g3444) & (!g3470) & (!g3493) & (g3495)) + ((!g1720) & (g3444) & (!g3470) & (g3493) & (!g3495)) + ((!g1720) & (g3444) & (!g3470) & (g3493) & (g3495)) + ((!g1720) & (g3444) & (g3470) & (!g3493) & (g3495)) + ((g1720) & (!g3444) & (!g3470) & (!g3493) & (!g3495)) + ((g1720) & (!g3444) & (!g3470) & (g3493) & (!g3495)) + ((g1720) & (!g3444) & (!g3470) & (g3493) & (g3495)) + ((g1720) & (g3444) & (!g3470) & (!g3493) & (g3495)) + ((g1720) & (g3444) & (g3470) & (!g3493) & (!g3495)) + ((g1720) & (g3444) & (g3470) & (!g3493) & (g3495)) + ((g1720) & (g3444) & (g3470) & (g3493) & (!g3495)) + ((g1720) & (g3444) & (g3470) & (g3493) & (g3495)));
	assign g3560 = (((!g1905) & (!g1879) & (g3446) & (g3469)) + ((!g1905) & (g1879) & (!g3446) & (g3469)) + ((!g1905) & (g1879) & (g3446) & (!g3469)) + ((!g1905) & (g1879) & (g3446) & (g3469)) + ((g1905) & (!g1879) & (!g3446) & (!g3469)) + ((g1905) & (!g1879) & (!g3446) & (g3469)) + ((g1905) & (!g1879) & (g3446) & (!g3469)) + ((g1905) & (g1879) & (!g3446) & (!g3469)));
	assign g3561 = (((!g3445) & (!g3493) & (!g3495) & (g3560)) + ((!g3445) & (g3493) & (!g3495) & (g3560)) + ((!g3445) & (g3493) & (g3495) & (g3560)) + ((g3445) & (!g3493) & (!g3495) & (!g3560)) + ((g3445) & (!g3493) & (g3495) & (!g3560)) + ((g3445) & (!g3493) & (g3495) & (g3560)) + ((g3445) & (g3493) & (!g3495) & (!g3560)) + ((g3445) & (g3493) & (g3495) & (!g3560)));
	assign g3562 = (((!g1879) & (!g3446) & (g3469) & (!g3493) & (!g3495)) + ((!g1879) & (!g3446) & (g3469) & (g3493) & (!g3495)) + ((!g1879) & (!g3446) & (g3469) & (g3493) & (g3495)) + ((!g1879) & (g3446) & (!g3469) & (!g3493) & (!g3495)) + ((!g1879) & (g3446) & (!g3469) & (!g3493) & (g3495)) + ((!g1879) & (g3446) & (!g3469) & (g3493) & (!g3495)) + ((!g1879) & (g3446) & (!g3469) & (g3493) & (g3495)) + ((!g1879) & (g3446) & (g3469) & (!g3493) & (g3495)) + ((g1879) & (!g3446) & (!g3469) & (!g3493) & (!g3495)) + ((g1879) & (!g3446) & (!g3469) & (g3493) & (!g3495)) + ((g1879) & (!g3446) & (!g3469) & (g3493) & (g3495)) + ((g1879) & (g3446) & (!g3469) & (!g3493) & (g3495)) + ((g1879) & (g3446) & (g3469) & (!g3493) & (!g3495)) + ((g1879) & (g3446) & (g3469) & (!g3493) & (g3495)) + ((g1879) & (g3446) & (g3469) & (g3493) & (!g3495)) + ((g1879) & (g3446) & (g3469) & (g3493) & (g3495)));
	assign g3563 = (((!g2075) & (!g2045) & (g3448) & (g3468)) + ((!g2075) & (g2045) & (!g3448) & (g3468)) + ((!g2075) & (g2045) & (g3448) & (!g3468)) + ((!g2075) & (g2045) & (g3448) & (g3468)) + ((g2075) & (!g2045) & (!g3448) & (!g3468)) + ((g2075) & (!g2045) & (!g3448) & (g3468)) + ((g2075) & (!g2045) & (g3448) & (!g3468)) + ((g2075) & (g2045) & (!g3448) & (!g3468)));
	assign g3564 = (((!g3447) & (!g3493) & (!g3495) & (g3563)) + ((!g3447) & (g3493) & (!g3495) & (g3563)) + ((!g3447) & (g3493) & (g3495) & (g3563)) + ((g3447) & (!g3493) & (!g3495) & (!g3563)) + ((g3447) & (!g3493) & (g3495) & (!g3563)) + ((g3447) & (!g3493) & (g3495) & (g3563)) + ((g3447) & (g3493) & (!g3495) & (!g3563)) + ((g3447) & (g3493) & (g3495) & (!g3563)));
	assign g3565 = (((!g2045) & (!g3448) & (g3468) & (!g3493) & (!g3495)) + ((!g2045) & (!g3448) & (g3468) & (g3493) & (!g3495)) + ((!g2045) & (!g3448) & (g3468) & (g3493) & (g3495)) + ((!g2045) & (g3448) & (!g3468) & (!g3493) & (!g3495)) + ((!g2045) & (g3448) & (!g3468) & (!g3493) & (g3495)) + ((!g2045) & (g3448) & (!g3468) & (g3493) & (!g3495)) + ((!g2045) & (g3448) & (!g3468) & (g3493) & (g3495)) + ((!g2045) & (g3448) & (g3468) & (!g3493) & (g3495)) + ((g2045) & (!g3448) & (!g3468) & (!g3493) & (!g3495)) + ((g2045) & (!g3448) & (!g3468) & (g3493) & (!g3495)) + ((g2045) & (!g3448) & (!g3468) & (g3493) & (g3495)) + ((g2045) & (g3448) & (!g3468) & (!g3493) & (g3495)) + ((g2045) & (g3448) & (g3468) & (!g3493) & (!g3495)) + ((g2045) & (g3448) & (g3468) & (!g3493) & (g3495)) + ((g2045) & (g3448) & (g3468) & (g3493) & (!g3495)) + ((g2045) & (g3448) & (g3468) & (g3493) & (g3495)));
	assign g3566 = (((!g2252) & (!g2218) & (g3450) & (g3467)) + ((!g2252) & (g2218) & (!g3450) & (g3467)) + ((!g2252) & (g2218) & (g3450) & (!g3467)) + ((!g2252) & (g2218) & (g3450) & (g3467)) + ((g2252) & (!g2218) & (!g3450) & (!g3467)) + ((g2252) & (!g2218) & (!g3450) & (g3467)) + ((g2252) & (!g2218) & (g3450) & (!g3467)) + ((g2252) & (g2218) & (!g3450) & (!g3467)));
	assign g3567 = (((!g3449) & (!g3493) & (!g3495) & (g3566)) + ((!g3449) & (g3493) & (!g3495) & (g3566)) + ((!g3449) & (g3493) & (g3495) & (g3566)) + ((g3449) & (!g3493) & (!g3495) & (!g3566)) + ((g3449) & (!g3493) & (g3495) & (!g3566)) + ((g3449) & (!g3493) & (g3495) & (g3566)) + ((g3449) & (g3493) & (!g3495) & (!g3566)) + ((g3449) & (g3493) & (g3495) & (!g3566)));
	assign g3568 = (((!g2218) & (!g3450) & (g3467) & (!g3493) & (!g3495)) + ((!g2218) & (!g3450) & (g3467) & (g3493) & (!g3495)) + ((!g2218) & (!g3450) & (g3467) & (g3493) & (g3495)) + ((!g2218) & (g3450) & (!g3467) & (!g3493) & (!g3495)) + ((!g2218) & (g3450) & (!g3467) & (!g3493) & (g3495)) + ((!g2218) & (g3450) & (!g3467) & (g3493) & (!g3495)) + ((!g2218) & (g3450) & (!g3467) & (g3493) & (g3495)) + ((!g2218) & (g3450) & (g3467) & (!g3493) & (g3495)) + ((g2218) & (!g3450) & (!g3467) & (!g3493) & (!g3495)) + ((g2218) & (!g3450) & (!g3467) & (g3493) & (!g3495)) + ((g2218) & (!g3450) & (!g3467) & (g3493) & (g3495)) + ((g2218) & (g3450) & (!g3467) & (!g3493) & (g3495)) + ((g2218) & (g3450) & (g3467) & (!g3493) & (!g3495)) + ((g2218) & (g3450) & (g3467) & (!g3493) & (g3495)) + ((g2218) & (g3450) & (g3467) & (g3493) & (!g3495)) + ((g2218) & (g3450) & (g3467) & (g3493) & (g3495)));
	assign g3569 = (((!g2436) & (!g2398) & (g3452) & (g3466)) + ((!g2436) & (g2398) & (!g3452) & (g3466)) + ((!g2436) & (g2398) & (g3452) & (!g3466)) + ((!g2436) & (g2398) & (g3452) & (g3466)) + ((g2436) & (!g2398) & (!g3452) & (!g3466)) + ((g2436) & (!g2398) & (!g3452) & (g3466)) + ((g2436) & (!g2398) & (g3452) & (!g3466)) + ((g2436) & (g2398) & (!g3452) & (!g3466)));
	assign g3570 = (((!g3451) & (!g3493) & (!g3495) & (g3569)) + ((!g3451) & (g3493) & (!g3495) & (g3569)) + ((!g3451) & (g3493) & (g3495) & (g3569)) + ((g3451) & (!g3493) & (!g3495) & (!g3569)) + ((g3451) & (!g3493) & (g3495) & (!g3569)) + ((g3451) & (!g3493) & (g3495) & (g3569)) + ((g3451) & (g3493) & (!g3495) & (!g3569)) + ((g3451) & (g3493) & (g3495) & (!g3569)));
	assign g3571 = (((!g2398) & (!g3452) & (g3466) & (!g3493) & (!g3495)) + ((!g2398) & (!g3452) & (g3466) & (g3493) & (!g3495)) + ((!g2398) & (!g3452) & (g3466) & (g3493) & (g3495)) + ((!g2398) & (g3452) & (!g3466) & (!g3493) & (!g3495)) + ((!g2398) & (g3452) & (!g3466) & (!g3493) & (g3495)) + ((!g2398) & (g3452) & (!g3466) & (g3493) & (!g3495)) + ((!g2398) & (g3452) & (!g3466) & (g3493) & (g3495)) + ((!g2398) & (g3452) & (g3466) & (!g3493) & (g3495)) + ((g2398) & (!g3452) & (!g3466) & (!g3493) & (!g3495)) + ((g2398) & (!g3452) & (!g3466) & (g3493) & (!g3495)) + ((g2398) & (!g3452) & (!g3466) & (g3493) & (g3495)) + ((g2398) & (g3452) & (!g3466) & (!g3493) & (g3495)) + ((g2398) & (g3452) & (g3466) & (!g3493) & (!g3495)) + ((g2398) & (g3452) & (g3466) & (!g3493) & (g3495)) + ((g2398) & (g3452) & (g3466) & (g3493) & (!g3495)) + ((g2398) & (g3452) & (g3466) & (g3493) & (g3495)));
	assign g3572 = (((!g2627) & (!g2585) & (g3454) & (g3465)) + ((!g2627) & (g2585) & (!g3454) & (g3465)) + ((!g2627) & (g2585) & (g3454) & (!g3465)) + ((!g2627) & (g2585) & (g3454) & (g3465)) + ((g2627) & (!g2585) & (!g3454) & (!g3465)) + ((g2627) & (!g2585) & (!g3454) & (g3465)) + ((g2627) & (!g2585) & (g3454) & (!g3465)) + ((g2627) & (g2585) & (!g3454) & (!g3465)));
	assign g3573 = (((!g3453) & (!g3493) & (!g3495) & (g3572)) + ((!g3453) & (g3493) & (!g3495) & (g3572)) + ((!g3453) & (g3493) & (g3495) & (g3572)) + ((g3453) & (!g3493) & (!g3495) & (!g3572)) + ((g3453) & (!g3493) & (g3495) & (!g3572)) + ((g3453) & (!g3493) & (g3495) & (g3572)) + ((g3453) & (g3493) & (!g3495) & (!g3572)) + ((g3453) & (g3493) & (g3495) & (!g3572)));
	assign g3574 = (((!g2585) & (!g3454) & (g3465) & (!g3493) & (!g3495)) + ((!g2585) & (!g3454) & (g3465) & (g3493) & (!g3495)) + ((!g2585) & (!g3454) & (g3465) & (g3493) & (g3495)) + ((!g2585) & (g3454) & (!g3465) & (!g3493) & (!g3495)) + ((!g2585) & (g3454) & (!g3465) & (!g3493) & (g3495)) + ((!g2585) & (g3454) & (!g3465) & (g3493) & (!g3495)) + ((!g2585) & (g3454) & (!g3465) & (g3493) & (g3495)) + ((!g2585) & (g3454) & (g3465) & (!g3493) & (g3495)) + ((g2585) & (!g3454) & (!g3465) & (!g3493) & (!g3495)) + ((g2585) & (!g3454) & (!g3465) & (g3493) & (!g3495)) + ((g2585) & (!g3454) & (!g3465) & (g3493) & (g3495)) + ((g2585) & (g3454) & (!g3465) & (!g3493) & (g3495)) + ((g2585) & (g3454) & (g3465) & (!g3493) & (!g3495)) + ((g2585) & (g3454) & (g3465) & (!g3493) & (g3495)) + ((g2585) & (g3454) & (g3465) & (g3493) & (!g3495)) + ((g2585) & (g3454) & (g3465) & (g3493) & (g3495)));
	assign g3575 = (((!g2825) & (!g2779) & (g3456) & (g3464)) + ((!g2825) & (g2779) & (!g3456) & (g3464)) + ((!g2825) & (g2779) & (g3456) & (!g3464)) + ((!g2825) & (g2779) & (g3456) & (g3464)) + ((g2825) & (!g2779) & (!g3456) & (!g3464)) + ((g2825) & (!g2779) & (!g3456) & (g3464)) + ((g2825) & (!g2779) & (g3456) & (!g3464)) + ((g2825) & (g2779) & (!g3456) & (!g3464)));
	assign g3576 = (((!g3455) & (!g3493) & (!g3495) & (g3575)) + ((!g3455) & (g3493) & (!g3495) & (g3575)) + ((!g3455) & (g3493) & (g3495) & (g3575)) + ((g3455) & (!g3493) & (!g3495) & (!g3575)) + ((g3455) & (!g3493) & (g3495) & (!g3575)) + ((g3455) & (!g3493) & (g3495) & (g3575)) + ((g3455) & (g3493) & (!g3495) & (!g3575)) + ((g3455) & (g3493) & (g3495) & (!g3575)));
	assign g3577 = (((!g2779) & (!g3456) & (g3464) & (!g3493) & (!g3495)) + ((!g2779) & (!g3456) & (g3464) & (g3493) & (!g3495)) + ((!g2779) & (!g3456) & (g3464) & (g3493) & (g3495)) + ((!g2779) & (g3456) & (!g3464) & (!g3493) & (!g3495)) + ((!g2779) & (g3456) & (!g3464) & (!g3493) & (g3495)) + ((!g2779) & (g3456) & (!g3464) & (g3493) & (!g3495)) + ((!g2779) & (g3456) & (!g3464) & (g3493) & (g3495)) + ((!g2779) & (g3456) & (g3464) & (!g3493) & (g3495)) + ((g2779) & (!g3456) & (!g3464) & (!g3493) & (!g3495)) + ((g2779) & (!g3456) & (!g3464) & (g3493) & (!g3495)) + ((g2779) & (!g3456) & (!g3464) & (g3493) & (g3495)) + ((g2779) & (g3456) & (!g3464) & (!g3493) & (g3495)) + ((g2779) & (g3456) & (g3464) & (!g3493) & (!g3495)) + ((g2779) & (g3456) & (g3464) & (!g3493) & (g3495)) + ((g2779) & (g3456) & (g3464) & (g3493) & (!g3495)) + ((g2779) & (g3456) & (g3464) & (g3493) & (g3495)));
	assign g3578 = (((!g3030) & (!g2980) & (g3458) & (g3463)) + ((!g3030) & (g2980) & (!g3458) & (g3463)) + ((!g3030) & (g2980) & (g3458) & (!g3463)) + ((!g3030) & (g2980) & (g3458) & (g3463)) + ((g3030) & (!g2980) & (!g3458) & (!g3463)) + ((g3030) & (!g2980) & (!g3458) & (g3463)) + ((g3030) & (!g2980) & (g3458) & (!g3463)) + ((g3030) & (g2980) & (!g3458) & (!g3463)));
	assign g3579 = (((!g3457) & (!g3493) & (!g3495) & (g3578)) + ((!g3457) & (g3493) & (!g3495) & (g3578)) + ((!g3457) & (g3493) & (g3495) & (g3578)) + ((g3457) & (!g3493) & (!g3495) & (!g3578)) + ((g3457) & (!g3493) & (g3495) & (!g3578)) + ((g3457) & (!g3493) & (g3495) & (g3578)) + ((g3457) & (g3493) & (!g3495) & (!g3578)) + ((g3457) & (g3493) & (g3495) & (!g3578)));
	assign g3580 = (((!g2980) & (!g3458) & (g3463) & (!g3493) & (!g3495)) + ((!g2980) & (!g3458) & (g3463) & (g3493) & (!g3495)) + ((!g2980) & (!g3458) & (g3463) & (g3493) & (g3495)) + ((!g2980) & (g3458) & (!g3463) & (!g3493) & (!g3495)) + ((!g2980) & (g3458) & (!g3463) & (!g3493) & (g3495)) + ((!g2980) & (g3458) & (!g3463) & (g3493) & (!g3495)) + ((!g2980) & (g3458) & (!g3463) & (g3493) & (g3495)) + ((!g2980) & (g3458) & (g3463) & (!g3493) & (g3495)) + ((g2980) & (!g3458) & (!g3463) & (!g3493) & (!g3495)) + ((g2980) & (!g3458) & (!g3463) & (g3493) & (!g3495)) + ((g2980) & (!g3458) & (!g3463) & (g3493) & (g3495)) + ((g2980) & (g3458) & (!g3463) & (!g3493) & (g3495)) + ((g2980) & (g3458) & (g3463) & (!g3493) & (!g3495)) + ((g2980) & (g3458) & (g3463) & (!g3493) & (g3495)) + ((g2980) & (g3458) & (g3463) & (g3493) & (!g3495)) + ((g2980) & (g3458) & (g3463) & (g3493) & (g3495)));
	assign g3581 = (((!g3178) & (!g3187) & (g3460) & (g3462)) + ((!g3178) & (g3187) & (!g3460) & (g3462)) + ((!g3178) & (g3187) & (g3460) & (!g3462)) + ((!g3178) & (g3187) & (g3460) & (g3462)) + ((g3178) & (!g3187) & (!g3460) & (!g3462)) + ((g3178) & (!g3187) & (!g3460) & (g3462)) + ((g3178) & (!g3187) & (g3460) & (!g3462)) + ((g3178) & (g3187) & (!g3460) & (!g3462)));
	assign g3582 = (((!g3459) & (!g3493) & (!g3495) & (g3581)) + ((!g3459) & (g3493) & (!g3495) & (g3581)) + ((!g3459) & (g3493) & (g3495) & (g3581)) + ((g3459) & (!g3493) & (!g3495) & (!g3581)) + ((g3459) & (!g3493) & (g3495) & (!g3581)) + ((g3459) & (!g3493) & (g3495) & (g3581)) + ((g3459) & (g3493) & (!g3495) & (!g3581)) + ((g3459) & (g3493) & (g3495) & (!g3581)));
	assign g3583 = (((!g3187) & (!g3460) & (g3462) & (!g3493) & (!g3495)) + ((!g3187) & (!g3460) & (g3462) & (g3493) & (!g3495)) + ((!g3187) & (!g3460) & (g3462) & (g3493) & (g3495)) + ((!g3187) & (g3460) & (!g3462) & (!g3493) & (!g3495)) + ((!g3187) & (g3460) & (!g3462) & (!g3493) & (g3495)) + ((!g3187) & (g3460) & (!g3462) & (g3493) & (!g3495)) + ((!g3187) & (g3460) & (!g3462) & (g3493) & (g3495)) + ((!g3187) & (g3460) & (g3462) & (!g3493) & (g3495)) + ((g3187) & (!g3460) & (!g3462) & (!g3493) & (!g3495)) + ((g3187) & (!g3460) & (!g3462) & (g3493) & (!g3495)) + ((g3187) & (!g3460) & (!g3462) & (g3493) & (g3495)) + ((g3187) & (g3460) & (!g3462) & (!g3493) & (g3495)) + ((g3187) & (g3460) & (g3462) & (!g3493) & (!g3495)) + ((g3187) & (g3460) & (g3462) & (!g3493) & (g3495)) + ((g3187) & (g3460) & (g3462) & (g3493) & (!g3495)) + ((g3187) & (g3460) & (g3462) & (g3493) & (g3495)));
	assign g3584 = (((!g3395) & (!ax4x) & (!g3400) & (g3461)) + ((!g3395) & (!ax4x) & (g3400) & (g3461)) + ((!g3395) & (ax4x) & (!g3400) & (!g3461)) + ((!g3395) & (ax4x) & (!g3400) & (g3461)) + ((g3395) & (!ax4x) & (!g3400) & (!g3461)) + ((g3395) & (!ax4x) & (g3400) & (!g3461)) + ((g3395) & (ax4x) & (g3400) & (!g3461)) + ((g3395) & (ax4x) & (g3400) & (g3461)));
	assign g3585 = (((!ax4x) & (!ax5x) & (!g3400) & (!g3493) & (!g3495) & (g3584)) + ((!ax4x) & (!ax5x) & (!g3400) & (!g3493) & (g3495) & (!g3584)) + ((!ax4x) & (!ax5x) & (!g3400) & (!g3493) & (g3495) & (g3584)) + ((!ax4x) & (!ax5x) & (!g3400) & (g3493) & (!g3495) & (g3584)) + ((!ax4x) & (!ax5x) & (!g3400) & (g3493) & (g3495) & (g3584)) + ((!ax4x) & (!ax5x) & (g3400) & (!g3493) & (!g3495) & (!g3584)) + ((!ax4x) & (!ax5x) & (g3400) & (g3493) & (!g3495) & (!g3584)) + ((!ax4x) & (!ax5x) & (g3400) & (g3493) & (g3495) & (!g3584)) + ((!ax4x) & (ax5x) & (!g3400) & (!g3493) & (!g3495) & (!g3584)) + ((!ax4x) & (ax5x) & (!g3400) & (g3493) & (!g3495) & (!g3584)) + ((!ax4x) & (ax5x) & (!g3400) & (g3493) & (g3495) & (!g3584)) + ((!ax4x) & (ax5x) & (g3400) & (!g3493) & (!g3495) & (g3584)) + ((!ax4x) & (ax5x) & (g3400) & (!g3493) & (g3495) & (!g3584)) + ((!ax4x) & (ax5x) & (g3400) & (!g3493) & (g3495) & (g3584)) + ((!ax4x) & (ax5x) & (g3400) & (g3493) & (!g3495) & (g3584)) + ((!ax4x) & (ax5x) & (g3400) & (g3493) & (g3495) & (g3584)) + ((ax4x) & (!ax5x) & (!g3400) & (!g3493) & (!g3495) & (!g3584)) + ((ax4x) & (!ax5x) & (!g3400) & (g3493) & (!g3495) & (!g3584)) + ((ax4x) & (!ax5x) & (!g3400) & (g3493) & (g3495) & (!g3584)) + ((ax4x) & (!ax5x) & (g3400) & (!g3493) & (!g3495) & (!g3584)) + ((ax4x) & (!ax5x) & (g3400) & (g3493) & (!g3495) & (!g3584)) + ((ax4x) & (!ax5x) & (g3400) & (g3493) & (g3495) & (!g3584)) + ((ax4x) & (ax5x) & (!g3400) & (!g3493) & (!g3495) & (g3584)) + ((ax4x) & (ax5x) & (!g3400) & (!g3493) & (g3495) & (!g3584)) + ((ax4x) & (ax5x) & (!g3400) & (!g3493) & (g3495) & (g3584)) + ((ax4x) & (ax5x) & (!g3400) & (g3493) & (!g3495) & (g3584)) + ((ax4x) & (ax5x) & (!g3400) & (g3493) & (g3495) & (g3584)) + ((ax4x) & (ax5x) & (g3400) & (!g3493) & (!g3495) & (g3584)) + ((ax4x) & (ax5x) & (g3400) & (!g3493) & (g3495) & (!g3584)) + ((ax4x) & (ax5x) & (g3400) & (!g3493) & (g3495) & (g3584)) + ((ax4x) & (ax5x) & (g3400) & (g3493) & (!g3495) & (g3584)) + ((ax4x) & (ax5x) & (g3400) & (g3493) & (g3495) & (g3584)));
	assign g3586 = (((!ax0x) & (!ax1x)));
	assign g3587 = (((!g3400) & (!ax2x) & (!ax3x) & (!g3493) & (!g3495) & (!g3586)) + ((!g3400) & (!ax2x) & (!ax3x) & (g3493) & (!g3495) & (!g3586)) + ((!g3400) & (!ax2x) & (!ax3x) & (g3493) & (g3495) & (!g3586)) + ((!g3400) & (!ax2x) & (ax3x) & (!g3493) & (g3495) & (!g3586)) + ((!g3400) & (ax2x) & (ax3x) & (!g3493) & (g3495) & (!g3586)) + ((!g3400) & (ax2x) & (ax3x) & (!g3493) & (g3495) & (g3586)) + ((g3400) & (!ax2x) & (!ax3x) & (!g3493) & (!g3495) & (!g3586)) + ((g3400) & (!ax2x) & (!ax3x) & (!g3493) & (!g3495) & (g3586)) + ((g3400) & (!ax2x) & (!ax3x) & (!g3493) & (g3495) & (!g3586)) + ((g3400) & (!ax2x) & (!ax3x) & (g3493) & (!g3495) & (!g3586)) + ((g3400) & (!ax2x) & (!ax3x) & (g3493) & (!g3495) & (g3586)) + ((g3400) & (!ax2x) & (!ax3x) & (g3493) & (g3495) & (!g3586)) + ((g3400) & (!ax2x) & (!ax3x) & (g3493) & (g3495) & (g3586)) + ((g3400) & (!ax2x) & (ax3x) & (!g3493) & (!g3495) & (!g3586)) + ((g3400) & (!ax2x) & (ax3x) & (!g3493) & (g3495) & (!g3586)) + ((g3400) & (!ax2x) & (ax3x) & (!g3493) & (g3495) & (g3586)) + ((g3400) & (!ax2x) & (ax3x) & (g3493) & (!g3495) & (!g3586)) + ((g3400) & (!ax2x) & (ax3x) & (g3493) & (g3495) & (!g3586)) + ((g3400) & (ax2x) & (!ax3x) & (!g3493) & (g3495) & (!g3586)) + ((g3400) & (ax2x) & (!ax3x) & (!g3493) & (g3495) & (g3586)) + ((g3400) & (ax2x) & (ax3x) & (!g3493) & (!g3495) & (!g3586)) + ((g3400) & (ax2x) & (ax3x) & (!g3493) & (!g3495) & (g3586)) + ((g3400) & (ax2x) & (ax3x) & (!g3493) & (g3495) & (!g3586)) + ((g3400) & (ax2x) & (ax3x) & (!g3493) & (g3495) & (g3586)) + ((g3400) & (ax2x) & (ax3x) & (g3493) & (!g3495) & (!g3586)) + ((g3400) & (ax2x) & (ax3x) & (g3493) & (!g3495) & (g3586)) + ((g3400) & (ax2x) & (ax3x) & (g3493) & (g3495) & (!g3586)) + ((g3400) & (ax2x) & (ax3x) & (g3493) & (g3495) & (g3586)));
	assign g3588 = (((!ax4x) & (!g3400) & (!g3461) & (!g3493) & (!g3495)) + ((!ax4x) & (!g3400) & (!g3461) & (g3493) & (!g3495)) + ((!ax4x) & (!g3400) & (!g3461) & (g3493) & (g3495)) + ((!ax4x) & (g3400) & (!g3461) & (!g3493) & (!g3495)) + ((!ax4x) & (g3400) & (!g3461) & (!g3493) & (g3495)) + ((!ax4x) & (g3400) & (!g3461) & (g3493) & (!g3495)) + ((!ax4x) & (g3400) & (!g3461) & (g3493) & (g3495)) + ((!ax4x) & (g3400) & (g3461) & (!g3493) & (g3495)) + ((ax4x) & (!g3400) & (!g3461) & (!g3493) & (g3495)) + ((ax4x) & (!g3400) & (g3461) & (!g3493) & (!g3495)) + ((ax4x) & (!g3400) & (g3461) & (!g3493) & (g3495)) + ((ax4x) & (!g3400) & (g3461) & (g3493) & (!g3495)) + ((ax4x) & (!g3400) & (g3461) & (g3493) & (g3495)) + ((ax4x) & (g3400) & (g3461) & (!g3493) & (!g3495)) + ((ax4x) & (g3400) & (g3461) & (g3493) & (!g3495)) + ((ax4x) & (g3400) & (g3461) & (g3493) & (g3495)));
	assign g3589 = (((!g3187) & (!g3395) & (!g3585) & (!g3587) & (!g3588)) + ((!g3187) & (!g3395) & (!g3585) & (!g3587) & (g3588)) + ((!g3187) & (!g3395) & (!g3585) & (g3587) & (!g3588)) + ((!g3187) & (!g3395) & (!g3585) & (g3587) & (g3588)) + ((!g3187) & (!g3395) & (g3585) & (!g3587) & (!g3588)) + ((!g3187) & (!g3395) & (g3585) & (!g3587) & (g3588)) + ((!g3187) & (!g3395) & (g3585) & (g3587) & (g3588)) + ((!g3187) & (g3395) & (!g3585) & (!g3587) & (!g3588)) + ((!g3187) & (g3395) & (!g3585) & (!g3587) & (g3588)) + ((!g3187) & (g3395) & (!g3585) & (g3587) & (!g3588)) + ((!g3187) & (g3395) & (!g3585) & (g3587) & (g3588)) + ((!g3187) & (g3395) & (g3585) & (!g3587) & (g3588)) + ((g3187) & (!g3395) & (!g3585) & (!g3587) & (!g3588)) + ((g3187) & (!g3395) & (!g3585) & (!g3587) & (g3588)) + ((g3187) & (!g3395) & (!g3585) & (g3587) & (g3588)) + ((g3187) & (g3395) & (!g3585) & (!g3587) & (g3588)));
	assign g3590 = (((!g2980) & (!g3178) & (!g3582) & (!g3583) & (!g3589)) + ((!g2980) & (!g3178) & (!g3582) & (!g3583) & (g3589)) + ((!g2980) & (!g3178) & (!g3582) & (g3583) & (!g3589)) + ((!g2980) & (!g3178) & (!g3582) & (g3583) & (g3589)) + ((!g2980) & (!g3178) & (g3582) & (!g3583) & (!g3589)) + ((!g2980) & (!g3178) & (g3582) & (!g3583) & (g3589)) + ((!g2980) & (!g3178) & (g3582) & (g3583) & (g3589)) + ((!g2980) & (g3178) & (!g3582) & (!g3583) & (!g3589)) + ((!g2980) & (g3178) & (!g3582) & (!g3583) & (g3589)) + ((!g2980) & (g3178) & (!g3582) & (g3583) & (!g3589)) + ((!g2980) & (g3178) & (!g3582) & (g3583) & (g3589)) + ((!g2980) & (g3178) & (g3582) & (!g3583) & (g3589)) + ((g2980) & (!g3178) & (!g3582) & (!g3583) & (!g3589)) + ((g2980) & (!g3178) & (!g3582) & (!g3583) & (g3589)) + ((g2980) & (!g3178) & (!g3582) & (g3583) & (g3589)) + ((g2980) & (g3178) & (!g3582) & (!g3583) & (g3589)));
	assign g3591 = (((!g2779) & (!g3030) & (!g3579) & (!g3580) & (!g3590)) + ((!g2779) & (!g3030) & (!g3579) & (!g3580) & (g3590)) + ((!g2779) & (!g3030) & (!g3579) & (g3580) & (!g3590)) + ((!g2779) & (!g3030) & (!g3579) & (g3580) & (g3590)) + ((!g2779) & (!g3030) & (g3579) & (!g3580) & (!g3590)) + ((!g2779) & (!g3030) & (g3579) & (!g3580) & (g3590)) + ((!g2779) & (!g3030) & (g3579) & (g3580) & (g3590)) + ((!g2779) & (g3030) & (!g3579) & (!g3580) & (!g3590)) + ((!g2779) & (g3030) & (!g3579) & (!g3580) & (g3590)) + ((!g2779) & (g3030) & (!g3579) & (g3580) & (!g3590)) + ((!g2779) & (g3030) & (!g3579) & (g3580) & (g3590)) + ((!g2779) & (g3030) & (g3579) & (!g3580) & (g3590)) + ((g2779) & (!g3030) & (!g3579) & (!g3580) & (!g3590)) + ((g2779) & (!g3030) & (!g3579) & (!g3580) & (g3590)) + ((g2779) & (!g3030) & (!g3579) & (g3580) & (g3590)) + ((g2779) & (g3030) & (!g3579) & (!g3580) & (g3590)));
	assign g3592 = (((!g2585) & (!g2825) & (!g3576) & (!g3577) & (!g3591)) + ((!g2585) & (!g2825) & (!g3576) & (!g3577) & (g3591)) + ((!g2585) & (!g2825) & (!g3576) & (g3577) & (!g3591)) + ((!g2585) & (!g2825) & (!g3576) & (g3577) & (g3591)) + ((!g2585) & (!g2825) & (g3576) & (!g3577) & (!g3591)) + ((!g2585) & (!g2825) & (g3576) & (!g3577) & (g3591)) + ((!g2585) & (!g2825) & (g3576) & (g3577) & (g3591)) + ((!g2585) & (g2825) & (!g3576) & (!g3577) & (!g3591)) + ((!g2585) & (g2825) & (!g3576) & (!g3577) & (g3591)) + ((!g2585) & (g2825) & (!g3576) & (g3577) & (!g3591)) + ((!g2585) & (g2825) & (!g3576) & (g3577) & (g3591)) + ((!g2585) & (g2825) & (g3576) & (!g3577) & (g3591)) + ((g2585) & (!g2825) & (!g3576) & (!g3577) & (!g3591)) + ((g2585) & (!g2825) & (!g3576) & (!g3577) & (g3591)) + ((g2585) & (!g2825) & (!g3576) & (g3577) & (g3591)) + ((g2585) & (g2825) & (!g3576) & (!g3577) & (g3591)));
	assign g3593 = (((!g2398) & (!g2627) & (!g3573) & (!g3574) & (!g3592)) + ((!g2398) & (!g2627) & (!g3573) & (!g3574) & (g3592)) + ((!g2398) & (!g2627) & (!g3573) & (g3574) & (!g3592)) + ((!g2398) & (!g2627) & (!g3573) & (g3574) & (g3592)) + ((!g2398) & (!g2627) & (g3573) & (!g3574) & (!g3592)) + ((!g2398) & (!g2627) & (g3573) & (!g3574) & (g3592)) + ((!g2398) & (!g2627) & (g3573) & (g3574) & (g3592)) + ((!g2398) & (g2627) & (!g3573) & (!g3574) & (!g3592)) + ((!g2398) & (g2627) & (!g3573) & (!g3574) & (g3592)) + ((!g2398) & (g2627) & (!g3573) & (g3574) & (!g3592)) + ((!g2398) & (g2627) & (!g3573) & (g3574) & (g3592)) + ((!g2398) & (g2627) & (g3573) & (!g3574) & (g3592)) + ((g2398) & (!g2627) & (!g3573) & (!g3574) & (!g3592)) + ((g2398) & (!g2627) & (!g3573) & (!g3574) & (g3592)) + ((g2398) & (!g2627) & (!g3573) & (g3574) & (g3592)) + ((g2398) & (g2627) & (!g3573) & (!g3574) & (g3592)));
	assign g3594 = (((!g2218) & (!g2436) & (!g3570) & (!g3571) & (!g3593)) + ((!g2218) & (!g2436) & (!g3570) & (!g3571) & (g3593)) + ((!g2218) & (!g2436) & (!g3570) & (g3571) & (!g3593)) + ((!g2218) & (!g2436) & (!g3570) & (g3571) & (g3593)) + ((!g2218) & (!g2436) & (g3570) & (!g3571) & (!g3593)) + ((!g2218) & (!g2436) & (g3570) & (!g3571) & (g3593)) + ((!g2218) & (!g2436) & (g3570) & (g3571) & (g3593)) + ((!g2218) & (g2436) & (!g3570) & (!g3571) & (!g3593)) + ((!g2218) & (g2436) & (!g3570) & (!g3571) & (g3593)) + ((!g2218) & (g2436) & (!g3570) & (g3571) & (!g3593)) + ((!g2218) & (g2436) & (!g3570) & (g3571) & (g3593)) + ((!g2218) & (g2436) & (g3570) & (!g3571) & (g3593)) + ((g2218) & (!g2436) & (!g3570) & (!g3571) & (!g3593)) + ((g2218) & (!g2436) & (!g3570) & (!g3571) & (g3593)) + ((g2218) & (!g2436) & (!g3570) & (g3571) & (g3593)) + ((g2218) & (g2436) & (!g3570) & (!g3571) & (g3593)));
	assign g3595 = (((!g2045) & (!g2252) & (!g3567) & (!g3568) & (!g3594)) + ((!g2045) & (!g2252) & (!g3567) & (!g3568) & (g3594)) + ((!g2045) & (!g2252) & (!g3567) & (g3568) & (!g3594)) + ((!g2045) & (!g2252) & (!g3567) & (g3568) & (g3594)) + ((!g2045) & (!g2252) & (g3567) & (!g3568) & (!g3594)) + ((!g2045) & (!g2252) & (g3567) & (!g3568) & (g3594)) + ((!g2045) & (!g2252) & (g3567) & (g3568) & (g3594)) + ((!g2045) & (g2252) & (!g3567) & (!g3568) & (!g3594)) + ((!g2045) & (g2252) & (!g3567) & (!g3568) & (g3594)) + ((!g2045) & (g2252) & (!g3567) & (g3568) & (!g3594)) + ((!g2045) & (g2252) & (!g3567) & (g3568) & (g3594)) + ((!g2045) & (g2252) & (g3567) & (!g3568) & (g3594)) + ((g2045) & (!g2252) & (!g3567) & (!g3568) & (!g3594)) + ((g2045) & (!g2252) & (!g3567) & (!g3568) & (g3594)) + ((g2045) & (!g2252) & (!g3567) & (g3568) & (g3594)) + ((g2045) & (g2252) & (!g3567) & (!g3568) & (g3594)));
	assign g3596 = (((!g1879) & (!g2075) & (!g3564) & (!g3565) & (!g3595)) + ((!g1879) & (!g2075) & (!g3564) & (!g3565) & (g3595)) + ((!g1879) & (!g2075) & (!g3564) & (g3565) & (!g3595)) + ((!g1879) & (!g2075) & (!g3564) & (g3565) & (g3595)) + ((!g1879) & (!g2075) & (g3564) & (!g3565) & (!g3595)) + ((!g1879) & (!g2075) & (g3564) & (!g3565) & (g3595)) + ((!g1879) & (!g2075) & (g3564) & (g3565) & (g3595)) + ((!g1879) & (g2075) & (!g3564) & (!g3565) & (!g3595)) + ((!g1879) & (g2075) & (!g3564) & (!g3565) & (g3595)) + ((!g1879) & (g2075) & (!g3564) & (g3565) & (!g3595)) + ((!g1879) & (g2075) & (!g3564) & (g3565) & (g3595)) + ((!g1879) & (g2075) & (g3564) & (!g3565) & (g3595)) + ((g1879) & (!g2075) & (!g3564) & (!g3565) & (!g3595)) + ((g1879) & (!g2075) & (!g3564) & (!g3565) & (g3595)) + ((g1879) & (!g2075) & (!g3564) & (g3565) & (g3595)) + ((g1879) & (g2075) & (!g3564) & (!g3565) & (g3595)));
	assign g3597 = (((!g1720) & (!g1905) & (!g3561) & (!g3562) & (!g3596)) + ((!g1720) & (!g1905) & (!g3561) & (!g3562) & (g3596)) + ((!g1720) & (!g1905) & (!g3561) & (g3562) & (!g3596)) + ((!g1720) & (!g1905) & (!g3561) & (g3562) & (g3596)) + ((!g1720) & (!g1905) & (g3561) & (!g3562) & (!g3596)) + ((!g1720) & (!g1905) & (g3561) & (!g3562) & (g3596)) + ((!g1720) & (!g1905) & (g3561) & (g3562) & (g3596)) + ((!g1720) & (g1905) & (!g3561) & (!g3562) & (!g3596)) + ((!g1720) & (g1905) & (!g3561) & (!g3562) & (g3596)) + ((!g1720) & (g1905) & (!g3561) & (g3562) & (!g3596)) + ((!g1720) & (g1905) & (!g3561) & (g3562) & (g3596)) + ((!g1720) & (g1905) & (g3561) & (!g3562) & (g3596)) + ((g1720) & (!g1905) & (!g3561) & (!g3562) & (!g3596)) + ((g1720) & (!g1905) & (!g3561) & (!g3562) & (g3596)) + ((g1720) & (!g1905) & (!g3561) & (g3562) & (g3596)) + ((g1720) & (g1905) & (!g3561) & (!g3562) & (g3596)));
	assign g3598 = (((!g1568) & (!g1742) & (!g3558) & (!g3559) & (!g3597)) + ((!g1568) & (!g1742) & (!g3558) & (!g3559) & (g3597)) + ((!g1568) & (!g1742) & (!g3558) & (g3559) & (!g3597)) + ((!g1568) & (!g1742) & (!g3558) & (g3559) & (g3597)) + ((!g1568) & (!g1742) & (g3558) & (!g3559) & (!g3597)) + ((!g1568) & (!g1742) & (g3558) & (!g3559) & (g3597)) + ((!g1568) & (!g1742) & (g3558) & (g3559) & (g3597)) + ((!g1568) & (g1742) & (!g3558) & (!g3559) & (!g3597)) + ((!g1568) & (g1742) & (!g3558) & (!g3559) & (g3597)) + ((!g1568) & (g1742) & (!g3558) & (g3559) & (!g3597)) + ((!g1568) & (g1742) & (!g3558) & (g3559) & (g3597)) + ((!g1568) & (g1742) & (g3558) & (!g3559) & (g3597)) + ((g1568) & (!g1742) & (!g3558) & (!g3559) & (!g3597)) + ((g1568) & (!g1742) & (!g3558) & (!g3559) & (g3597)) + ((g1568) & (!g1742) & (!g3558) & (g3559) & (g3597)) + ((g1568) & (g1742) & (!g3558) & (!g3559) & (g3597)));
	assign g3599 = (((!g1423) & (!g1586) & (!g3555) & (!g3556) & (!g3598)) + ((!g1423) & (!g1586) & (!g3555) & (!g3556) & (g3598)) + ((!g1423) & (!g1586) & (!g3555) & (g3556) & (!g3598)) + ((!g1423) & (!g1586) & (!g3555) & (g3556) & (g3598)) + ((!g1423) & (!g1586) & (g3555) & (!g3556) & (!g3598)) + ((!g1423) & (!g1586) & (g3555) & (!g3556) & (g3598)) + ((!g1423) & (!g1586) & (g3555) & (g3556) & (g3598)) + ((!g1423) & (g1586) & (!g3555) & (!g3556) & (!g3598)) + ((!g1423) & (g1586) & (!g3555) & (!g3556) & (g3598)) + ((!g1423) & (g1586) & (!g3555) & (g3556) & (!g3598)) + ((!g1423) & (g1586) & (!g3555) & (g3556) & (g3598)) + ((!g1423) & (g1586) & (g3555) & (!g3556) & (g3598)) + ((g1423) & (!g1586) & (!g3555) & (!g3556) & (!g3598)) + ((g1423) & (!g1586) & (!g3555) & (!g3556) & (g3598)) + ((g1423) & (!g1586) & (!g3555) & (g3556) & (g3598)) + ((g1423) & (g1586) & (!g3555) & (!g3556) & (g3598)));
	assign g3600 = (((!g1285) & (!g1437) & (!g3552) & (!g3553) & (!g3599)) + ((!g1285) & (!g1437) & (!g3552) & (!g3553) & (g3599)) + ((!g1285) & (!g1437) & (!g3552) & (g3553) & (!g3599)) + ((!g1285) & (!g1437) & (!g3552) & (g3553) & (g3599)) + ((!g1285) & (!g1437) & (g3552) & (!g3553) & (!g3599)) + ((!g1285) & (!g1437) & (g3552) & (!g3553) & (g3599)) + ((!g1285) & (!g1437) & (g3552) & (g3553) & (g3599)) + ((!g1285) & (g1437) & (!g3552) & (!g3553) & (!g3599)) + ((!g1285) & (g1437) & (!g3552) & (!g3553) & (g3599)) + ((!g1285) & (g1437) & (!g3552) & (g3553) & (!g3599)) + ((!g1285) & (g1437) & (!g3552) & (g3553) & (g3599)) + ((!g1285) & (g1437) & (g3552) & (!g3553) & (g3599)) + ((g1285) & (!g1437) & (!g3552) & (!g3553) & (!g3599)) + ((g1285) & (!g1437) & (!g3552) & (!g3553) & (g3599)) + ((g1285) & (!g1437) & (!g3552) & (g3553) & (g3599)) + ((g1285) & (g1437) & (!g3552) & (!g3553) & (g3599)));
	assign g3601 = (((!g1154) & (!g1295) & (!g3549) & (!g3550) & (!g3600)) + ((!g1154) & (!g1295) & (!g3549) & (!g3550) & (g3600)) + ((!g1154) & (!g1295) & (!g3549) & (g3550) & (!g3600)) + ((!g1154) & (!g1295) & (!g3549) & (g3550) & (g3600)) + ((!g1154) & (!g1295) & (g3549) & (!g3550) & (!g3600)) + ((!g1154) & (!g1295) & (g3549) & (!g3550) & (g3600)) + ((!g1154) & (!g1295) & (g3549) & (g3550) & (g3600)) + ((!g1154) & (g1295) & (!g3549) & (!g3550) & (!g3600)) + ((!g1154) & (g1295) & (!g3549) & (!g3550) & (g3600)) + ((!g1154) & (g1295) & (!g3549) & (g3550) & (!g3600)) + ((!g1154) & (g1295) & (!g3549) & (g3550) & (g3600)) + ((!g1154) & (g1295) & (g3549) & (!g3550) & (g3600)) + ((g1154) & (!g1295) & (!g3549) & (!g3550) & (!g3600)) + ((g1154) & (!g1295) & (!g3549) & (!g3550) & (g3600)) + ((g1154) & (!g1295) & (!g3549) & (g3550) & (g3600)) + ((g1154) & (g1295) & (!g3549) & (!g3550) & (g3600)));
	assign g3602 = (((!g1030) & (!g1160) & (!g3546) & (!g3547) & (!g3601)) + ((!g1030) & (!g1160) & (!g3546) & (!g3547) & (g3601)) + ((!g1030) & (!g1160) & (!g3546) & (g3547) & (!g3601)) + ((!g1030) & (!g1160) & (!g3546) & (g3547) & (g3601)) + ((!g1030) & (!g1160) & (g3546) & (!g3547) & (!g3601)) + ((!g1030) & (!g1160) & (g3546) & (!g3547) & (g3601)) + ((!g1030) & (!g1160) & (g3546) & (g3547) & (g3601)) + ((!g1030) & (g1160) & (!g3546) & (!g3547) & (!g3601)) + ((!g1030) & (g1160) & (!g3546) & (!g3547) & (g3601)) + ((!g1030) & (g1160) & (!g3546) & (g3547) & (!g3601)) + ((!g1030) & (g1160) & (!g3546) & (g3547) & (g3601)) + ((!g1030) & (g1160) & (g3546) & (!g3547) & (g3601)) + ((g1030) & (!g1160) & (!g3546) & (!g3547) & (!g3601)) + ((g1030) & (!g1160) & (!g3546) & (!g3547) & (g3601)) + ((g1030) & (!g1160) & (!g3546) & (g3547) & (g3601)) + ((g1030) & (g1160) & (!g3546) & (!g3547) & (g3601)));
	assign g3603 = (((!g914) & (!g1032) & (!g3543) & (!g3544) & (!g3602)) + ((!g914) & (!g1032) & (!g3543) & (!g3544) & (g3602)) + ((!g914) & (!g1032) & (!g3543) & (g3544) & (!g3602)) + ((!g914) & (!g1032) & (!g3543) & (g3544) & (g3602)) + ((!g914) & (!g1032) & (g3543) & (!g3544) & (!g3602)) + ((!g914) & (!g1032) & (g3543) & (!g3544) & (g3602)) + ((!g914) & (!g1032) & (g3543) & (g3544) & (g3602)) + ((!g914) & (g1032) & (!g3543) & (!g3544) & (!g3602)) + ((!g914) & (g1032) & (!g3543) & (!g3544) & (g3602)) + ((!g914) & (g1032) & (!g3543) & (g3544) & (!g3602)) + ((!g914) & (g1032) & (!g3543) & (g3544) & (g3602)) + ((!g914) & (g1032) & (g3543) & (!g3544) & (g3602)) + ((g914) & (!g1032) & (!g3543) & (!g3544) & (!g3602)) + ((g914) & (!g1032) & (!g3543) & (!g3544) & (g3602)) + ((g914) & (!g1032) & (!g3543) & (g3544) & (g3602)) + ((g914) & (g1032) & (!g3543) & (!g3544) & (g3602)));
	assign g3604 = (((!g803) & (!g851) & (!g3540) & (!g3541) & (!g3603)) + ((!g803) & (!g851) & (!g3540) & (!g3541) & (g3603)) + ((!g803) & (!g851) & (!g3540) & (g3541) & (!g3603)) + ((!g803) & (!g851) & (!g3540) & (g3541) & (g3603)) + ((!g803) & (!g851) & (g3540) & (!g3541) & (!g3603)) + ((!g803) & (!g851) & (g3540) & (!g3541) & (g3603)) + ((!g803) & (!g851) & (g3540) & (g3541) & (g3603)) + ((!g803) & (g851) & (!g3540) & (!g3541) & (!g3603)) + ((!g803) & (g851) & (!g3540) & (!g3541) & (g3603)) + ((!g803) & (g851) & (!g3540) & (g3541) & (!g3603)) + ((!g803) & (g851) & (!g3540) & (g3541) & (g3603)) + ((!g803) & (g851) & (g3540) & (!g3541) & (g3603)) + ((g803) & (!g851) & (!g3540) & (!g3541) & (!g3603)) + ((g803) & (!g851) & (!g3540) & (!g3541) & (g3603)) + ((g803) & (!g851) & (!g3540) & (g3541) & (g3603)) + ((g803) & (g851) & (!g3540) & (!g3541) & (g3603)));
	assign g3605 = (((!g700) & (!g744) & (!g3537) & (!g3538) & (!g3604)) + ((!g700) & (!g744) & (!g3537) & (!g3538) & (g3604)) + ((!g700) & (!g744) & (!g3537) & (g3538) & (!g3604)) + ((!g700) & (!g744) & (!g3537) & (g3538) & (g3604)) + ((!g700) & (!g744) & (g3537) & (!g3538) & (!g3604)) + ((!g700) & (!g744) & (g3537) & (!g3538) & (g3604)) + ((!g700) & (!g744) & (g3537) & (g3538) & (g3604)) + ((!g700) & (g744) & (!g3537) & (!g3538) & (!g3604)) + ((!g700) & (g744) & (!g3537) & (!g3538) & (g3604)) + ((!g700) & (g744) & (!g3537) & (g3538) & (!g3604)) + ((!g700) & (g744) & (!g3537) & (g3538) & (g3604)) + ((!g700) & (g744) & (g3537) & (!g3538) & (g3604)) + ((g700) & (!g744) & (!g3537) & (!g3538) & (!g3604)) + ((g700) & (!g744) & (!g3537) & (!g3538) & (g3604)) + ((g700) & (!g744) & (!g3537) & (g3538) & (g3604)) + ((g700) & (g744) & (!g3537) & (!g3538) & (g3604)));
	assign g3606 = (((!g604) & (!g645) & (!g3534) & (!g3535) & (!g3605)) + ((!g604) & (!g645) & (!g3534) & (!g3535) & (g3605)) + ((!g604) & (!g645) & (!g3534) & (g3535) & (!g3605)) + ((!g604) & (!g645) & (!g3534) & (g3535) & (g3605)) + ((!g604) & (!g645) & (g3534) & (!g3535) & (!g3605)) + ((!g604) & (!g645) & (g3534) & (!g3535) & (g3605)) + ((!g604) & (!g645) & (g3534) & (g3535) & (g3605)) + ((!g604) & (g645) & (!g3534) & (!g3535) & (!g3605)) + ((!g604) & (g645) & (!g3534) & (!g3535) & (g3605)) + ((!g604) & (g645) & (!g3534) & (g3535) & (!g3605)) + ((!g604) & (g645) & (!g3534) & (g3535) & (g3605)) + ((!g604) & (g645) & (g3534) & (!g3535) & (g3605)) + ((g604) & (!g645) & (!g3534) & (!g3535) & (!g3605)) + ((g604) & (!g645) & (!g3534) & (!g3535) & (g3605)) + ((g604) & (!g645) & (!g3534) & (g3535) & (g3605)) + ((g604) & (g645) & (!g3534) & (!g3535) & (g3605)));
	assign g3607 = (((!g515) & (!g553) & (!g3531) & (!g3532) & (!g3606)) + ((!g515) & (!g553) & (!g3531) & (!g3532) & (g3606)) + ((!g515) & (!g553) & (!g3531) & (g3532) & (!g3606)) + ((!g515) & (!g553) & (!g3531) & (g3532) & (g3606)) + ((!g515) & (!g553) & (g3531) & (!g3532) & (!g3606)) + ((!g515) & (!g553) & (g3531) & (!g3532) & (g3606)) + ((!g515) & (!g553) & (g3531) & (g3532) & (g3606)) + ((!g515) & (g553) & (!g3531) & (!g3532) & (!g3606)) + ((!g515) & (g553) & (!g3531) & (!g3532) & (g3606)) + ((!g515) & (g553) & (!g3531) & (g3532) & (!g3606)) + ((!g515) & (g553) & (!g3531) & (g3532) & (g3606)) + ((!g515) & (g553) & (g3531) & (!g3532) & (g3606)) + ((g515) & (!g553) & (!g3531) & (!g3532) & (!g3606)) + ((g515) & (!g553) & (!g3531) & (!g3532) & (g3606)) + ((g515) & (!g553) & (!g3531) & (g3532) & (g3606)) + ((g515) & (g553) & (!g3531) & (!g3532) & (g3606)));
	assign g3608 = (((!g433) & (!g468) & (!g3528) & (!g3529) & (!g3607)) + ((!g433) & (!g468) & (!g3528) & (!g3529) & (g3607)) + ((!g433) & (!g468) & (!g3528) & (g3529) & (!g3607)) + ((!g433) & (!g468) & (!g3528) & (g3529) & (g3607)) + ((!g433) & (!g468) & (g3528) & (!g3529) & (!g3607)) + ((!g433) & (!g468) & (g3528) & (!g3529) & (g3607)) + ((!g433) & (!g468) & (g3528) & (g3529) & (g3607)) + ((!g433) & (g468) & (!g3528) & (!g3529) & (!g3607)) + ((!g433) & (g468) & (!g3528) & (!g3529) & (g3607)) + ((!g433) & (g468) & (!g3528) & (g3529) & (!g3607)) + ((!g433) & (g468) & (!g3528) & (g3529) & (g3607)) + ((!g433) & (g468) & (g3528) & (!g3529) & (g3607)) + ((g433) & (!g468) & (!g3528) & (!g3529) & (!g3607)) + ((g433) & (!g468) & (!g3528) & (!g3529) & (g3607)) + ((g433) & (!g468) & (!g3528) & (g3529) & (g3607)) + ((g433) & (g468) & (!g3528) & (!g3529) & (g3607)));
	assign g3609 = (((!g358) & (!g390) & (!g3525) & (!g3526) & (!g3608)) + ((!g358) & (!g390) & (!g3525) & (!g3526) & (g3608)) + ((!g358) & (!g390) & (!g3525) & (g3526) & (!g3608)) + ((!g358) & (!g390) & (!g3525) & (g3526) & (g3608)) + ((!g358) & (!g390) & (g3525) & (!g3526) & (!g3608)) + ((!g358) & (!g390) & (g3525) & (!g3526) & (g3608)) + ((!g358) & (!g390) & (g3525) & (g3526) & (g3608)) + ((!g358) & (g390) & (!g3525) & (!g3526) & (!g3608)) + ((!g358) & (g390) & (!g3525) & (!g3526) & (g3608)) + ((!g358) & (g390) & (!g3525) & (g3526) & (!g3608)) + ((!g358) & (g390) & (!g3525) & (g3526) & (g3608)) + ((!g358) & (g390) & (g3525) & (!g3526) & (g3608)) + ((g358) & (!g390) & (!g3525) & (!g3526) & (!g3608)) + ((g358) & (!g390) & (!g3525) & (!g3526) & (g3608)) + ((g358) & (!g390) & (!g3525) & (g3526) & (g3608)) + ((g358) & (g390) & (!g3525) & (!g3526) & (g3608)));
	assign g3610 = (((!g290) & (!g319) & (!g3522) & (!g3523) & (!g3609)) + ((!g290) & (!g319) & (!g3522) & (!g3523) & (g3609)) + ((!g290) & (!g319) & (!g3522) & (g3523) & (!g3609)) + ((!g290) & (!g319) & (!g3522) & (g3523) & (g3609)) + ((!g290) & (!g319) & (g3522) & (!g3523) & (!g3609)) + ((!g290) & (!g319) & (g3522) & (!g3523) & (g3609)) + ((!g290) & (!g319) & (g3522) & (g3523) & (g3609)) + ((!g290) & (g319) & (!g3522) & (!g3523) & (!g3609)) + ((!g290) & (g319) & (!g3522) & (!g3523) & (g3609)) + ((!g290) & (g319) & (!g3522) & (g3523) & (!g3609)) + ((!g290) & (g319) & (!g3522) & (g3523) & (g3609)) + ((!g290) & (g319) & (g3522) & (!g3523) & (g3609)) + ((g290) & (!g319) & (!g3522) & (!g3523) & (!g3609)) + ((g290) & (!g319) & (!g3522) & (!g3523) & (g3609)) + ((g290) & (!g319) & (!g3522) & (g3523) & (g3609)) + ((g290) & (g319) & (!g3522) & (!g3523) & (g3609)));
	assign g3611 = (((!g229) & (!g255) & (!g3519) & (!g3520) & (!g3610)) + ((!g229) & (!g255) & (!g3519) & (!g3520) & (g3610)) + ((!g229) & (!g255) & (!g3519) & (g3520) & (!g3610)) + ((!g229) & (!g255) & (!g3519) & (g3520) & (g3610)) + ((!g229) & (!g255) & (g3519) & (!g3520) & (!g3610)) + ((!g229) & (!g255) & (g3519) & (!g3520) & (g3610)) + ((!g229) & (!g255) & (g3519) & (g3520) & (g3610)) + ((!g229) & (g255) & (!g3519) & (!g3520) & (!g3610)) + ((!g229) & (g255) & (!g3519) & (!g3520) & (g3610)) + ((!g229) & (g255) & (!g3519) & (g3520) & (!g3610)) + ((!g229) & (g255) & (!g3519) & (g3520) & (g3610)) + ((!g229) & (g255) & (g3519) & (!g3520) & (g3610)) + ((g229) & (!g255) & (!g3519) & (!g3520) & (!g3610)) + ((g229) & (!g255) & (!g3519) & (!g3520) & (g3610)) + ((g229) & (!g255) & (!g3519) & (g3520) & (g3610)) + ((g229) & (g255) & (!g3519) & (!g3520) & (g3610)));
	assign g3612 = (((!g174) & (!g198) & (!g3516) & (!g3517) & (!g3611)) + ((!g174) & (!g198) & (!g3516) & (!g3517) & (g3611)) + ((!g174) & (!g198) & (!g3516) & (g3517) & (!g3611)) + ((!g174) & (!g198) & (!g3516) & (g3517) & (g3611)) + ((!g174) & (!g198) & (g3516) & (!g3517) & (!g3611)) + ((!g174) & (!g198) & (g3516) & (!g3517) & (g3611)) + ((!g174) & (!g198) & (g3516) & (g3517) & (g3611)) + ((!g174) & (g198) & (!g3516) & (!g3517) & (!g3611)) + ((!g174) & (g198) & (!g3516) & (!g3517) & (g3611)) + ((!g174) & (g198) & (!g3516) & (g3517) & (!g3611)) + ((!g174) & (g198) & (!g3516) & (g3517) & (g3611)) + ((!g174) & (g198) & (g3516) & (!g3517) & (g3611)) + ((g174) & (!g198) & (!g3516) & (!g3517) & (!g3611)) + ((g174) & (!g198) & (!g3516) & (!g3517) & (g3611)) + ((g174) & (!g198) & (!g3516) & (g3517) & (g3611)) + ((g174) & (g198) & (!g3516) & (!g3517) & (g3611)));
	assign g3613 = (((!g127) & (!g147) & (!g3513) & (!g3514) & (!g3612)) + ((!g127) & (!g147) & (!g3513) & (!g3514) & (g3612)) + ((!g127) & (!g147) & (!g3513) & (g3514) & (!g3612)) + ((!g127) & (!g147) & (!g3513) & (g3514) & (g3612)) + ((!g127) & (!g147) & (g3513) & (!g3514) & (!g3612)) + ((!g127) & (!g147) & (g3513) & (!g3514) & (g3612)) + ((!g127) & (!g147) & (g3513) & (g3514) & (g3612)) + ((!g127) & (g147) & (!g3513) & (!g3514) & (!g3612)) + ((!g127) & (g147) & (!g3513) & (!g3514) & (g3612)) + ((!g127) & (g147) & (!g3513) & (g3514) & (!g3612)) + ((!g127) & (g147) & (!g3513) & (g3514) & (g3612)) + ((!g127) & (g147) & (g3513) & (!g3514) & (g3612)) + ((g127) & (!g147) & (!g3513) & (!g3514) & (!g3612)) + ((g127) & (!g147) & (!g3513) & (!g3514) & (g3612)) + ((g127) & (!g147) & (!g3513) & (g3514) & (g3612)) + ((g127) & (g147) & (!g3513) & (!g3514) & (g3612)));
	assign g3614 = (((!g87) & (!g104) & (!g3510) & (!g3511) & (!g3613)) + ((!g87) & (!g104) & (!g3510) & (!g3511) & (g3613)) + ((!g87) & (!g104) & (!g3510) & (g3511) & (!g3613)) + ((!g87) & (!g104) & (!g3510) & (g3511) & (g3613)) + ((!g87) & (!g104) & (g3510) & (!g3511) & (!g3613)) + ((!g87) & (!g104) & (g3510) & (!g3511) & (g3613)) + ((!g87) & (!g104) & (g3510) & (g3511) & (g3613)) + ((!g87) & (g104) & (!g3510) & (!g3511) & (!g3613)) + ((!g87) & (g104) & (!g3510) & (!g3511) & (g3613)) + ((!g87) & (g104) & (!g3510) & (g3511) & (!g3613)) + ((!g87) & (g104) & (!g3510) & (g3511) & (g3613)) + ((!g87) & (g104) & (g3510) & (!g3511) & (g3613)) + ((g87) & (!g104) & (!g3510) & (!g3511) & (!g3613)) + ((g87) & (!g104) & (!g3510) & (!g3511) & (g3613)) + ((g87) & (!g104) & (!g3510) & (g3511) & (g3613)) + ((g87) & (g104) & (!g3510) & (!g3511) & (g3613)));
	assign g3615 = (((!g54) & (!g68) & (!g3507) & (!g3508) & (!g3614)) + ((!g54) & (!g68) & (!g3507) & (!g3508) & (g3614)) + ((!g54) & (!g68) & (!g3507) & (g3508) & (!g3614)) + ((!g54) & (!g68) & (!g3507) & (g3508) & (g3614)) + ((!g54) & (!g68) & (g3507) & (!g3508) & (!g3614)) + ((!g54) & (!g68) & (g3507) & (!g3508) & (g3614)) + ((!g54) & (!g68) & (g3507) & (g3508) & (g3614)) + ((!g54) & (g68) & (!g3507) & (!g3508) & (!g3614)) + ((!g54) & (g68) & (!g3507) & (!g3508) & (g3614)) + ((!g54) & (g68) & (!g3507) & (g3508) & (!g3614)) + ((!g54) & (g68) & (!g3507) & (g3508) & (g3614)) + ((!g54) & (g68) & (g3507) & (!g3508) & (g3614)) + ((g54) & (!g68) & (!g3507) & (!g3508) & (!g3614)) + ((g54) & (!g68) & (!g3507) & (!g3508) & (g3614)) + ((g54) & (!g68) & (!g3507) & (g3508) & (g3614)) + ((g54) & (g68) & (!g3507) & (!g3508) & (g3614)));
	assign g3616 = (((!g27) & (!g39) & (!g3504) & (!g3505) & (!g3615)) + ((!g27) & (!g39) & (!g3504) & (!g3505) & (g3615)) + ((!g27) & (!g39) & (!g3504) & (g3505) & (!g3615)) + ((!g27) & (!g39) & (!g3504) & (g3505) & (g3615)) + ((!g27) & (!g39) & (g3504) & (!g3505) & (!g3615)) + ((!g27) & (!g39) & (g3504) & (!g3505) & (g3615)) + ((!g27) & (!g39) & (g3504) & (g3505) & (g3615)) + ((!g27) & (g39) & (!g3504) & (!g3505) & (!g3615)) + ((!g27) & (g39) & (!g3504) & (!g3505) & (g3615)) + ((!g27) & (g39) & (!g3504) & (g3505) & (!g3615)) + ((!g27) & (g39) & (!g3504) & (g3505) & (g3615)) + ((!g27) & (g39) & (g3504) & (!g3505) & (g3615)) + ((g27) & (!g39) & (!g3504) & (!g3505) & (!g3615)) + ((g27) & (!g39) & (!g3504) & (!g3505) & (g3615)) + ((g27) & (!g39) & (!g3504) & (g3505) & (g3615)) + ((g27) & (g39) & (!g3504) & (!g3505) & (g3615)));
	assign g3617 = (((!g8) & (!g18) & (!g3501) & (!g3502) & (!g3616)) + ((!g8) & (!g18) & (!g3501) & (!g3502) & (g3616)) + ((!g8) & (!g18) & (!g3501) & (g3502) & (!g3616)) + ((!g8) & (!g18) & (!g3501) & (g3502) & (g3616)) + ((!g8) & (!g18) & (g3501) & (!g3502) & (!g3616)) + ((!g8) & (!g18) & (g3501) & (!g3502) & (g3616)) + ((!g8) & (!g18) & (g3501) & (g3502) & (g3616)) + ((!g8) & (g18) & (!g3501) & (!g3502) & (!g3616)) + ((!g8) & (g18) & (!g3501) & (!g3502) & (g3616)) + ((!g8) & (g18) & (!g3501) & (g3502) & (!g3616)) + ((!g8) & (g18) & (!g3501) & (g3502) & (g3616)) + ((!g8) & (g18) & (g3501) & (!g3502) & (g3616)) + ((g8) & (!g18) & (!g3501) & (!g3502) & (!g3616)) + ((g8) & (!g18) & (!g3501) & (!g3502) & (g3616)) + ((g8) & (!g18) & (!g3501) & (g3502) & (g3616)) + ((g8) & (g18) & (!g3501) & (!g3502) & (g3616)));
	assign g3618 = (((!g4) & (!g2) & (!g3498) & (g3499) & (!g3617)) + ((!g4) & (!g2) & (g3498) & (!g3499) & (!g3617)) + ((!g4) & (!g2) & (g3498) & (!g3499) & (g3617)) + ((!g4) & (!g2) & (g3498) & (g3499) & (!g3617)) + ((!g4) & (!g2) & (g3498) & (g3499) & (g3617)) + ((!g4) & (g2) & (!g3498) & (!g3499) & (!g3617)) + ((!g4) & (g2) & (!g3498) & (g3499) & (!g3617)) + ((!g4) & (g2) & (!g3498) & (g3499) & (g3617)) + ((!g4) & (g2) & (g3498) & (!g3499) & (!g3617)) + ((!g4) & (g2) & (g3498) & (!g3499) & (g3617)) + ((!g4) & (g2) & (g3498) & (g3499) & (!g3617)) + ((!g4) & (g2) & (g3498) & (g3499) & (g3617)));
	assign g3619 = (((!g4) & (!g2) & (!g8) & (!g3403) & (!g3404) & (!g3490)) + ((!g4) & (!g2) & (!g8) & (!g3403) & (!g3404) & (g3490)) + ((!g4) & (!g2) & (!g8) & (!g3403) & (g3404) & (!g3490)) + ((!g4) & (!g2) & (!g8) & (!g3403) & (g3404) & (g3490)) + ((!g4) & (!g2) & (!g8) & (g3403) & (!g3404) & (!g3490)) + ((!g4) & (!g2) & (!g8) & (g3403) & (!g3404) & (g3490)) + ((!g4) & (!g2) & (!g8) & (g3403) & (g3404) & (!g3490)) + ((!g4) & (!g2) & (g8) & (!g3403) & (!g3404) & (!g3490)) + ((!g4) & (!g2) & (g8) & (!g3403) & (!g3404) & (g3490)) + ((!g4) & (!g2) & (g8) & (!g3403) & (g3404) & (!g3490)) + ((!g4) & (!g2) & (g8) & (!g3403) & (g3404) & (g3490)) + ((!g4) & (!g2) & (g8) & (g3403) & (!g3404) & (!g3490)) + ((!g4) & (g2) & (!g8) & (!g3403) & (!g3404) & (!g3490)) + ((!g4) & (g2) & (!g8) & (!g3403) & (!g3404) & (g3490)) + ((!g4) & (g2) & (!g8) & (!g3403) & (g3404) & (!g3490)) + ((!g4) & (g2) & (g8) & (!g3403) & (!g3404) & (!g3490)) + ((g4) & (!g2) & (!g8) & (g3403) & (g3404) & (g3490)) + ((g4) & (!g2) & (g8) & (g3403) & (!g3404) & (g3490)) + ((g4) & (!g2) & (g8) & (g3403) & (g3404) & (!g3490)) + ((g4) & (!g2) & (g8) & (g3403) & (g3404) & (g3490)) + ((g4) & (g2) & (!g8) & (!g3403) & (g3404) & (g3490)) + ((g4) & (g2) & (!g8) & (g3403) & (!g3404) & (!g3490)) + ((g4) & (g2) & (!g8) & (g3403) & (!g3404) & (g3490)) + ((g4) & (g2) & (!g8) & (g3403) & (g3404) & (!g3490)) + ((g4) & (g2) & (!g8) & (g3403) & (g3404) & (g3490)) + ((g4) & (g2) & (g8) & (!g3403) & (!g3404) & (g3490)) + ((g4) & (g2) & (g8) & (!g3403) & (g3404) & (!g3490)) + ((g4) & (g2) & (g8) & (!g3403) & (g3404) & (g3490)) + ((g4) & (g2) & (g8) & (g3403) & (!g3404) & (!g3490)) + ((g4) & (g2) & (g8) & (g3403) & (!g3404) & (g3490)) + ((g4) & (g2) & (g8) & (g3403) & (g3404) & (!g3490)) + ((g4) & (g2) & (g8) & (g3403) & (g3404) & (g3490)));
	assign g3620 = (((!g1) & (!g3403) & (!g3493) & (!g3495) & (g3497)) + ((!g1) & (!g3403) & (g3493) & (!g3495) & (g3497)) + ((!g1) & (!g3403) & (g3493) & (g3495) & (g3497)) + ((!g1) & (g3403) & (!g3493) & (!g3495) & (!g3497)) + ((!g1) & (g3403) & (!g3493) & (g3495) & (!g3497)) + ((!g1) & (g3403) & (!g3493) & (g3495) & (g3497)) + ((!g1) & (g3403) & (g3493) & (!g3495) & (!g3497)) + ((!g1) & (g3403) & (g3493) & (g3495) & (!g3497)));
	assign g3621 = (((!g3403) & (!g3401) & (!g3493) & (!g3495) & (g3497) & (g3619)) + ((!g3403) & (!g3401) & (g3493) & (!g3495) & (g3497) & (g3619)) + ((!g3403) & (!g3401) & (g3493) & (g3495) & (g3497) & (g3619)) + ((!g3403) & (g3401) & (!g3493) & (!g3495) & (g3497) & (!g3619)) + ((!g3403) & (g3401) & (g3493) & (!g3495) & (g3497) & (!g3619)) + ((!g3403) & (g3401) & (g3493) & (g3495) & (g3497) & (!g3619)) + ((g3403) & (!g3401) & (!g3493) & (!g3495) & (!g3497) & (g3619)) + ((g3403) & (!g3401) & (g3493) & (!g3495) & (!g3497) & (g3619)) + ((g3403) & (!g3401) & (g3493) & (g3495) & (!g3497) & (g3619)) + ((g3403) & (g3401) & (!g3493) & (!g3495) & (!g3497) & (!g3619)) + ((g3403) & (g3401) & (!g3493) & (g3495) & (!g3497) & (!g3619)) + ((g3403) & (g3401) & (!g3493) & (g3495) & (!g3497) & (g3619)) + ((g3403) & (g3401) & (!g3493) & (g3495) & (g3497) & (!g3619)) + ((g3403) & (g3401) & (!g3493) & (g3495) & (g3497) & (g3619)) + ((g3403) & (g3401) & (g3493) & (!g3495) & (!g3497) & (!g3619)) + ((g3403) & (g3401) & (g3493) & (g3495) & (!g3497) & (!g3619)));
	assign g3622 = (((!g4) & (!g1) & (!g3402) & (!g3491) & (!g3401) & (g3496)) + ((!g4) & (!g1) & (!g3402) & (!g3491) & (g3401) & (!g3496)) + ((!g4) & (!g1) & (!g3402) & (g3491) & (!g3401) & (!g3496)) + ((!g4) & (!g1) & (!g3402) & (g3491) & (!g3401) & (g3496)) + ((!g4) & (!g1) & (g3402) & (!g3491) & (!g3401) & (g3496)) + ((!g4) & (g1) & (!g3402) & (!g3491) & (!g3401) & (!g3496)) + ((!g4) & (g1) & (!g3402) & (!g3491) & (!g3401) & (g3496)) + ((!g4) & (g1) & (!g3402) & (!g3491) & (g3401) & (g3496)) + ((!g4) & (g1) & (!g3402) & (g3491) & (!g3401) & (g3496)) + ((!g4) & (g1) & (!g3402) & (g3491) & (g3401) & (g3496)) + ((!g4) & (g1) & (g3402) & (!g3491) & (g3401) & (!g3496)) + ((!g4) & (g1) & (g3402) & (!g3491) & (g3401) & (g3496)) + ((!g4) & (g1) & (g3402) & (g3491) & (!g3401) & (!g3496)) + ((!g4) & (g1) & (g3402) & (g3491) & (!g3401) & (g3496)) + ((!g4) & (g1) & (g3402) & (g3491) & (g3401) & (!g3496)) + ((!g4) & (g1) & (g3402) & (g3491) & (g3401) & (g3496)) + ((g4) & (!g1) & (!g3402) & (!g3491) & (!g3401) & (g3496)) + ((g4) & (!g1) & (!g3402) & (g3491) & (!g3401) & (g3496)) + ((g4) & (!g1) & (!g3402) & (g3491) & (g3401) & (!g3496)) + ((g4) & (!g1) & (g3402) & (!g3491) & (!g3401) & (!g3496)) + ((g4) & (!g1) & (g3402) & (!g3491) & (!g3401) & (g3496)) + ((g4) & (!g1) & (g3402) & (g3491) & (!g3401) & (g3496)) + ((g4) & (g1) & (!g3402) & (!g3491) & (!g3401) & (!g3496)) + ((g4) & (g1) & (!g3402) & (!g3491) & (!g3401) & (g3496)) + ((g4) & (g1) & (!g3402) & (!g3491) & (g3401) & (!g3496)) + ((g4) & (g1) & (!g3402) & (!g3491) & (g3401) & (g3496)) + ((g4) & (g1) & (!g3402) & (g3491) & (!g3401) & (!g3496)) + ((g4) & (g1) & (!g3402) & (g3491) & (!g3401) & (g3496)) + ((g4) & (g1) & (!g3402) & (g3491) & (g3401) & (g3496)) + ((g4) & (g1) & (g3402) & (g3491) & (g3401) & (!g3496)) + ((g4) & (g1) & (g3402) & (g3491) & (g3401) & (g3496)));
	assign g3623 = (((!g2) & (!g3499) & (!g3617) & (!g3620) & (!g3621) & (g3622)) + ((!g2) & (!g3499) & (!g3617) & (!g3620) & (g3621) & (g3622)) + ((!g2) & (!g3499) & (!g3617) & (g3620) & (!g3621) & (g3622)) + ((!g2) & (!g3499) & (!g3617) & (g3620) & (g3621) & (g3622)) + ((!g2) & (!g3499) & (g3617) & (!g3620) & (!g3621) & (g3622)) + ((!g2) & (!g3499) & (g3617) & (!g3620) & (g3621) & (g3622)) + ((!g2) & (!g3499) & (g3617) & (g3620) & (!g3621) & (g3622)) + ((!g2) & (!g3499) & (g3617) & (g3620) & (g3621) & (g3622)) + ((!g2) & (g3499) & (!g3617) & (!g3620) & (!g3621) & (g3622)) + ((!g2) & (g3499) & (g3617) & (!g3620) & (!g3621) & (g3622)) + ((!g2) & (g3499) & (g3617) & (!g3620) & (g3621) & (g3622)) + ((!g2) & (g3499) & (g3617) & (g3620) & (!g3621) & (g3622)) + ((!g2) & (g3499) & (g3617) & (g3620) & (g3621) & (g3622)) + ((g2) & (!g3499) & (!g3617) & (!g3620) & (!g3621) & (g3622)) + ((g2) & (!g3499) & (g3617) & (!g3620) & (!g3621) & (g3622)) + ((g2) & (!g3499) & (g3617) & (!g3620) & (g3621) & (g3622)) + ((g2) & (!g3499) & (g3617) & (g3620) & (!g3621) & (g3622)) + ((g2) & (!g3499) & (g3617) & (g3620) & (g3621) & (g3622)) + ((g2) & (g3499) & (!g3617) & (!g3620) & (!g3621) & (g3622)) + ((g2) & (g3499) & (g3617) & (!g3620) & (!g3621) & (g3622)));
	assign asqrtx0x = (((!g1) & (!g3401) & (!g3496) & (!g3618) & (!g3619) & (!g3623)) + ((!g1) & (!g3401) & (!g3496) & (!g3618) & (g3619) & (!g3623)) + ((!g1) & (!g3401) & (!g3496) & (g3618) & (!g3619) & (!g3623)) + ((!g1) & (!g3401) & (!g3496) & (g3618) & (!g3619) & (g3623)) + ((!g1) & (!g3401) & (!g3496) & (g3618) & (g3619) & (!g3623)) + ((!g1) & (!g3401) & (!g3496) & (g3618) & (g3619) & (g3623)) + ((!g1) & (!g3401) & (g3496) & (!g3618) & (!g3619) & (!g3623)) + ((!g1) & (!g3401) & (g3496) & (!g3618) & (g3619) & (!g3623)) + ((!g1) & (!g3401) & (g3496) & (g3618) & (!g3619) & (!g3623)) + ((!g1) & (!g3401) & (g3496) & (g3618) & (!g3619) & (g3623)) + ((!g1) & (!g3401) & (g3496) & (g3618) & (g3619) & (!g3623)) + ((!g1) & (!g3401) & (g3496) & (g3618) & (g3619) & (g3623)) + ((!g1) & (g3401) & (!g3496) & (!g3618) & (!g3619) & (!g3623)) + ((!g1) & (g3401) & (!g3496) & (!g3618) & (g3619) & (!g3623)) + ((!g1) & (g3401) & (!g3496) & (g3618) & (!g3619) & (!g3623)) + ((!g1) & (g3401) & (!g3496) & (g3618) & (!g3619) & (g3623)) + ((!g1) & (g3401) & (!g3496) & (g3618) & (g3619) & (!g3623)) + ((!g1) & (g3401) & (!g3496) & (g3618) & (g3619) & (g3623)) + ((!g1) & (g3401) & (g3496) & (!g3618) & (!g3619) & (!g3623)) + ((!g1) & (g3401) & (g3496) & (!g3618) & (g3619) & (!g3623)) + ((!g1) & (g3401) & (g3496) & (g3618) & (!g3619) & (!g3623)) + ((!g1) & (g3401) & (g3496) & (g3618) & (!g3619) & (g3623)) + ((!g1) & (g3401) & (g3496) & (g3618) & (g3619) & (!g3623)) + ((!g1) & (g3401) & (g3496) & (g3618) & (g3619) & (g3623)) + ((g1) & (!g3401) & (!g3496) & (!g3618) & (!g3619) & (!g3623)) + ((g1) & (!g3401) & (!g3496) & (!g3618) & (g3619) & (!g3623)) + ((g1) & (!g3401) & (!g3496) & (g3618) & (!g3619) & (!g3623)) + ((g1) & (!g3401) & (!g3496) & (g3618) & (g3619) & (!g3623)) + ((g1) & (!g3401) & (!g3496) & (g3618) & (g3619) & (g3623)) + ((g1) & (!g3401) & (g3496) & (!g3618) & (!g3619) & (!g3623)) + ((g1) & (!g3401) & (g3496) & (!g3618) & (g3619) & (!g3623)) + ((g1) & (!g3401) & (g3496) & (g3618) & (!g3619) & (!g3623)) + ((g1) & (!g3401) & (g3496) & (g3618) & (g3619) & (!g3623)) + ((g1) & (g3401) & (!g3496) & (!g3618) & (!g3619) & (!g3623)) + ((g1) & (g3401) & (!g3496) & (!g3618) & (g3619) & (!g3623)) + ((g1) & (g3401) & (!g3496) & (g3618) & (!g3619) & (!g3623)) + ((g1) & (g3401) & (!g3496) & (g3618) & (!g3619) & (g3623)) + ((g1) & (g3401) & (!g3496) & (g3618) & (g3619) & (!g3623)) + ((g1) & (g3401) & (g3496) & (!g3618) & (!g3619) & (!g3623)) + ((g1) & (g3401) & (g3496) & (!g3618) & (g3619) & (!g3623)) + ((g1) & (g3401) & (g3496) & (g3618) & (!g3619) & (!g3623)) + ((g1) & (g3401) & (g3496) & (g3618) & (!g3619) & (g3623)) + ((g1) & (g3401) & (g3496) & (g3618) & (g3619) & (!g3623)) + ((g1) & (g3401) & (g3496) & (g3618) & (g3619) & (g3623)));

endmodule