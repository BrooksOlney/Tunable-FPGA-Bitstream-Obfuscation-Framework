module apex4x6xv (i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_, o_1_, o_2_, o_12_, o_11_, o_14_, o_13_, o_16_, o_15_, o_18_, o_17_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

	input i_7_;
	input i_8_;
	input i_5_;
	input i_6_;
	input i_3_;
	input i_4_;
	input i_1_;
	input i_2_;
	input i_0_;
	output o_1_;
	output o_2_;
	output o_12_;
	output o_11_;
	output o_14_;
	output o_13_;
	output o_16_;
	output o_15_;
	output o_18_;
	output o_17_;
	output o_10_;
	output o_9_;
	output o_7_;
	output o_8_;
	output o_5_;
	output o_6_;
	output o_3_;
	output o_4_;

	wire [809 : 0] sk /* synthesis noprune */;

	lut_sub lut_3 ({sk[0], n_n110, x4863x, x4864x, x4865x, x4866x}, o_1_);
	defparam lut_3.LUT_SIZE = 6;
	defparam lut_3.mask = 64'h0f0f0f0f7fffffff;

	lut_sub lut_9 ({sk[1], x4991x, x4989x, x4990x}, o_2_);
	defparam lut_9.LUT_SIZE = 4;
	defparam lut_9.mask = 16'h037f;

	lut_sub lut_13 ({sk[2], x5048x, x5049x}, o_12_);
	defparam lut_13.LUT_SIZE = 3;
	defparam lut_13.mask = 8'h57;

	lut_sub lut_16 ({sk[3], x5110x, x5080x, x5081x, x5102x, x5103x, x5106x}, o_11_);
	defparam lut_16.LUT_SIZE = 7;
	defparam lut_16.mask = 128'h57ff57ff57ff5fff7fffffffffffffff;

	lut_sub lut_23 ({sk[4], x5169x, x5125x, x5123x, x5124x, x5162x, x5163x}, o_14_);
	defparam lut_23.LUT_SIZE = 7;
	defparam lut_23.mask = 128'h57ff57ff57ff5fff7fffffffffffffff;

	lut_sub lut_30 ({sk[5], x5220x, x5221x}, o_13_);
	defparam lut_30.LUT_SIZE = 3;
	defparam lut_30.mask = 8'h57;

	lut_sub lut_33 ({sk[6], x5232x, x178x, x258x, x310x, x5230x}, o_16_);
	defparam lut_33.LUT_SIZE = 6;
	defparam lut_33.mask = 64'h0f0f0f0f7fffffff;

	lut_sub lut_39 ({sk[7], x5249x, x5243x, x5244x, x5247x}, o_15_);
	defparam lut_39.LUT_SIZE = 5;
	defparam lut_39.mask = 32'h57577fff;

	lut_sub lut_44 ({sk[8], x5264x, x230x, x188x, x114x, x5259x, x6386x}, o_18_);
	defparam lut_44.LUT_SIZE = 7;
	defparam lut_44.mask = 128'h57ff57ff57ff5fffbfffffffffffffff;

	lut_sub lut_51 ({sk[9], x5271x, n_n91, x82x, n_n1259, n_n1176, x248x}, o_17_);
	defparam lut_51.LUT_SIZE = 7;
	defparam lut_51.mask = 128'h57ff57ff57ff5fff7f7f7fffffffffff;

	lut_sub lut_57 ({sk[10], x5373x, n_n655, x5372x}, o_10_);
	defparam lut_57.LUT_SIZE = 4;
	defparam lut_57.mask = 16'h037f;

	lut_sub lut_61 ({sk[11], x5403x, n_n324, n_n397, x5487x, x5488x, x5489x}, o_9_);
	defparam lut_61.LUT_SIZE = 7;
	defparam lut_61.mask = 128'h5f5fffff5f5fffff7fffffffffffffff;

	lut_sub lut_68 ({sk[12], x5539x, x5540x, x5589x, x5590x}, o_7_);
	defparam lut_68.LUT_SIZE = 5;
	defparam lut_68.mask = 32'h5f5f7fff;

	lut_sub lut_73 ({sk[13], x5685x, x5658x, x5648x, x5649x, x5650x, x5651x}, o_8_);
	defparam lut_73.LUT_SIZE = 7;
	defparam lut_73.mask = 128'h0000ffff0033ffff7fffffffffffffff;

	lut_sub lut_80 ({sk[14], x5732x, x5733x, x5779x, x5780x}, o_5_);
	defparam lut_80.LUT_SIZE = 5;
	defparam lut_80.mask = 32'h57577fff;

	lut_sub lut_85 ({sk[15], x5821x, x5822x, x5875x, x5876x}, o_6_);
	defparam lut_85.LUT_SIZE = 5;
	defparam lut_85.mask = 32'h57577fff;

	lut_sub lut_90 ({sk[16], n_n206, n_n208, n_n201, x5933x, x5939x, x5940x}, o_3_);
	defparam lut_90.LUT_SIZE = 7;
	defparam lut_90.mask = 128'h3fff7fff3fff7fff7fffffffffffffff;

	lut_sub lut_97 ({sk[17], x6028x, n_n243, x6019x, x6020x, x6021x, x6022x}, o_4_);
	defparam lut_97.LUT_SIZE = 7;
	defparam lut_97.mask = 128'h3fff7fff3fff7fff7fffffffffffffff;

	lut_sub lut_104 ({sk[18], n_n91, x4839x, n_n1120, n_n956, x128x, x355x}, n_n110);
	defparam lut_104.LUT_SIZE = 7;
	defparam lut_104.mask = 128'h3fff7fff3fff7fff5fffffff7fffffff;

	lut_sub lut_110 ({sk[19], x113x, x176x, x182x, x208x}, x4863x);
	defparam lut_110.LUT_SIZE = 5;
	defparam lut_110.mask = 32'h57577fff;

	lut_sub lut_115 ({sk[20], n_n86, n_n73, x27x, x252x, x329x, x6393x}, x4864x);
	defparam lut_115.LUT_SIZE = 7;
	defparam lut_115.mask = 128'h777f777fffffffff7f7f7f7f7f7f7fff;

	lut_sub lut_120 ({sk[21], x27x, x45x, x192x, x4847x, x4848x, x4850x}, x4865x);
	defparam lut_120.LUT_SIZE = 7;
	defparam lut_120.mask = 128'h777f777fffffffff7f7f7fff7fff7fff;

	lut_sub lut_126 ({sk[22], n_n58, x26x, x39x, x87x, x104x, x4861x}, x4866x);
	defparam lut_126.LUT_SIZE = 7;
	defparam lut_126.mask = 128'h777f777fffffffff7f7f7f7f7fffffff;

	lut_sub lut_132 ({sk[23], n_n136, n_n139, x4979x, x4980x, x4983x}, x4991x);
	defparam lut_132.LUT_SIZE = 6;
	defparam lut_132.mask = 64'h00ffffff7fffffff;

	lut_sub lut_138 ({sk[24], x4899x, x4897x, x4898x, x4981x, x4982x}, x4989x);
	defparam lut_138.LUT_SIZE = 6;
	defparam lut_138.mask = 64'h00ffffff7fffffff;

	lut_sub lut_144 ({sk[25], x4919x, n_n137, n_n135, x4917x, x4918x}, x4990x);
	defparam lut_144.LUT_SIZE = 6;
	defparam lut_144.mask = 64'h00ffffff7fffffff;

	lut_sub lut_150 ({sk[26], x179x, x181x, x222x, x255x, x5045x, x5046x}, x5048x);
	defparam lut_150.LUT_SIZE = 7;
	defparam lut_150.mask = 128'h3f3f3f3f7f7f7f7f7fffffffffffffff;

	lut_sub lut_157 ({sk[27], x5010x, x5029x, x5008x, x5009x, x5027x, x5028x}, x5049x);
	defparam lut_157.LUT_SIZE = 7;
	defparam lut_157.mask = 128'h3f3f3f3f7f7f7f7f7fffffffffffffff;

	lut_sub lut_164 ({sk[28], x5066x, x5064x, x5065x, x5104x, x5105x}, x5110x);
	defparam lut_164.LUT_SIZE = 6;
	defparam lut_164.mask = 64'h333333337fffffff;

	lut_sub lut_170 ({sk[29], x42x, n_n95, x297x, x147x, x202x, x6371x}, x5080x);
	defparam lut_170.LUT_SIZE = 7;
	defparam lut_170.mask = 128'h3f3f3f3f7f7f7f7fbfffbfffbfffffff;

	lut_sub lut_176 ({sk[30], x97x, x146x, x270x, x272x, x151x, x6350x}, x5081x);
	defparam lut_176.LUT_SIZE = 7;
	defparam lut_176.mask = 128'h3f3f3f3f7f7f7f7fbfffffffffffffff;

	lut_sub lut_183 ({sk[31], i_7_, i_6_, x39x, x93x, x197x, x5083x}, x5102x);
	defparam lut_183.LUT_SIZE = 7;
	defparam lut_183.mask = 128'h00ff00ff33ff33ff7f7f7f7f7f7f7fff;

	lut_sub lut_188 ({sk[32], x27x, n_n95, x117x, x133x, x148x, x323x}, x5103x);
	defparam lut_188.LUT_SIZE = 7;
	defparam lut_188.mask = 128'h00ff00ff33ff33ff7fff7fff7fffffff;

	lut_sub lut_194 ({sk[33], n_n1120, n_n1052, x233x, x5091x, x5092x}, x5106x);
	defparam lut_194.LUT_SIZE = 6;
	defparam lut_194.mask = 64'h7f7f7fff7fffffff;

	lut_sub lut_200 ({sk[34], x5139x, x5137x, x5138x, x5160x, x5161x, x5164x}, x5169x);
	defparam lut_200.LUT_SIZE = 7;
	defparam lut_200.mask = 128'h00ff00ff33ff33ff7fffffffffffffff;

	lut_sub lut_207 ({sk[35], n_n95, x41x, n_n949, n_n882, x296x, x5115x}, x5125x);
	defparam lut_207.LUT_SIZE = 7;
	defparam lut_207.mask = 128'h00ff00ff33ff33ff7fff7fff7fffffff;

	lut_sub lut_213 ({sk[36], n_n91, x29x, x271x, x145x, x146x, n_n939}, x5123x);
	defparam lut_213.LUT_SIZE = 7;
	defparam lut_213.mask = 128'h55ff55ff5fff5fff7fff7fff7fffffff;

	lut_sub lut_219 ({sk[37], n_n81, n_n91, n_n94, x270x, x272x, x6384x}, x5124x);
	defparam lut_219.LUT_SIZE = 7;
	defparam lut_219.mask = 128'h55ff55ff5fff5fffbfbfbfbfbfbfbfff;

	lut_sub lut_224 ({sk[38], x184x, x186x, x206x, x273x}, x5162x);
	defparam lut_224.LUT_SIZE = 5;
	defparam lut_224.mask = 32'h00ff7fff;

	lut_sub lut_229 ({sk[39], n_n58, n_n1259, x67x, n_n1330, n_n1267, x5156x}, x5163x);
	defparam lut_229.LUT_SIZE = 7;
	defparam lut_229.mask = 128'h55ff55ff5fff5fff7f7fffff7fffffff;

	lut_sub lut_235 ({sk[40], x89x, x183x, x184x, x186x, x5217x, x5218x}, x5220x);
	defparam lut_235.LUT_SIZE = 7;
	defparam lut_235.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_242 ({sk[41], x5185x, x5202x, x5183x, x5184x, x5200x, x5201x}, x5221x);
	defparam lut_242.LUT_SIZE = 7;
	defparam lut_242.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_249 ({sk[42], n_n1369, n_n1176, x187x, n_n1109, n_n1132, x294x}, x5232x);
	defparam lut_249.LUT_SIZE = 7;
	defparam lut_249.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_256 ({sk[43], i_7_, i_8_, i_6_, x76x, n_n74, n_n90}, x178x);
	defparam lut_256.LUT_SIZE = 7;
	defparam lut_256.mask = 128'h33ffffff33ffffff1100000f00000000;

	lut_sub lut_259 ({sk[44], i_7_, i_8_, i_6_, n_n74, x49x, n_n90}, x258x);
	defparam lut_259.LUT_SIZE = 7;
	defparam lut_259.mask = 128'h33ffffff33ffffff3300000500000000;

	lut_sub lut_262 ({sk[45], i_7_, i_8_, i_6_, n_n96, n_n90, x51x}, x310x);
	defparam lut_262.LUT_SIZE = 7;
	defparam lut_262.mask = 128'h33ffffff33ffffff0000000300570003;

	lut_sub lut_267 ({sk[46], i_7_, i_8_, i_6_, x43x, n_n1074, n_n1294}, x5230x);
	defparam lut_267.LUT_SIZE = 7;
	defparam lut_267.mask = 128'h33ffffff33ffffff777f77777f777f77;

	lut_sub lut_272 ({sk[47], x178x, x258x, x259x, x294x, x310x, x302x}, x5249x);
	defparam lut_272.LUT_SIZE = 7;
	defparam lut_272.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_279 ({sk[48], n_n93, n_n91, x43x, n_n1259, n_n1169, x86x}, x5243x);
	defparam lut_279.LUT_SIZE = 7;
	defparam lut_279.mask = 128'h33ffffff33ffffff3f3f7f7f3fff7fff;

	lut_sub lut_284 ({sk[49], i_7_, i_8_, i_6_, x73x, x67x, x51x}, x5244x);
	defparam lut_284.LUT_SIZE = 7;
	defparam lut_284.mask = 128'h33ffffff33ffffff3f0000000f000055;

	lut_sub lut_289 ({sk[50], n_n1324, n_n1369, x136x, x230x, x278x}, x5247x);
	defparam lut_289.LUT_SIZE = 6;
	defparam lut_289.mask = 64'h33ff33ff7fffffff;

	lut_sub lut_295 ({sk[51], n_n81, n_n82, n_n90, n_n1294, n_n1169, x6385x}, x5264x);
	defparam lut_295.LUT_SIZE = 7;
	defparam lut_295.mask = 128'h33ffffff33ffffffbfbfbfbfbfbfbfff;

	lut_sub lut_300 ({sk[52], i_7_, i_8_, i_6_, x49x, x86x}, x230x);
	defparam lut_300.LUT_SIZE = 6;
	defparam lut_300.mask = 64'h33ff33ff00003505;

	lut_sub lut_303 ({sk[53], i_7_, i_8_, i_6_, n_n81, n_n102, n_n90}, x188x);
	defparam lut_303.LUT_SIZE = 7;
	defparam lut_303.mask = 128'h33ffffff33ffffff0000050000110000;

	lut_sub lut_306 ({sk[54], i_5_, i_3_, i_4_, n_n93, n_n78, n_n94}, x114x);
	defparam lut_306.LUT_SIZE = 7;
	defparam lut_306.mask = 128'h33ffffff33ffffff0000001100000500;

	lut_sub lut_309 ({sk[55], i_7_, i_8_, i_1_, n_n1324, x72x, n_n1074}, x5259x);
	defparam lut_309.LUT_SIZE = 7;
	defparam lut_309.mask = 128'h33ffffff33ffffff7f5f5f5f5f5f5f5f;

	lut_sub lut_313 ({sk[56], n_n58, x39x, x136x, n_n937, x1315x, n_n941}, x6386x);
	defparam lut_313.LUT_SIZE = 7;
	defparam lut_313.mask = 128'h33ffffff33ffffff8000800080000000;

	lut_sub lut_316 ({sk[57], n_n58, x39x, x187x, x259x, x294x, n_n941}, x5271x);
	defparam lut_316.LUT_SIZE = 7;
	defparam lut_316.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_322 ({sk[58], i_7_, i_8_, i_6_}, n_n91);
	defparam lut_322.LUT_SIZE = 4;
	defparam lut_322.mask = 16'h7710;

	lut_sub lut_324 ({sk[59], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x82x);
	defparam lut_324.LUT_SIZE = 7;
	defparam lut_324.mask = 128'h33ffffff33ffffff0000000020000000;

	lut_sub lut_326 ({sk[60], i_7_, i_8_, i_6_, i_3_, x109x, n_n90}, n_n1259);
	defparam lut_326.LUT_SIZE = 7;
	defparam lut_326.mask = 128'h33ffffff33ffffff0000010000000000;

	lut_sub lut_328 ({sk[61], i_7_, i_8_, i_6_, n_n94, n_n74}, n_n1176);
	defparam lut_328.LUT_SIZE = 6;
	defparam lut_328.mask = 64'h33ff33ff00010000;

	lut_sub lut_330 ({sk[62], i_7_, i_8_, i_6_, n_n94, n_n77}, x248x);
	defparam lut_330.LUT_SIZE = 6;
	defparam lut_330.mask = 64'h33ff33ff00000001;

	lut_sub lut_332 ({sk[63], x5335x, x5333x, x5334x, x5367x, x5368x}, x5373x);
	defparam lut_332.LUT_SIZE = 6;
	defparam lut_332.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_338 ({sk[64], n_n663, x5308x, x5309x, x5310x, x5311x, x5312x}, n_n655);
	defparam lut_338.LUT_SIZE = 7;
	defparam lut_338.mask = 128'h0fffffff0fffffff7fffffffffffffff;

	lut_sub lut_345 ({sk[65], x137x, x90x, x298x, x5364x, x5365x, x5366x}, x5372x);
	defparam lut_345.LUT_SIZE = 7;
	defparam lut_345.mask = 128'h0fffffff0fffffff7fffffffffffffff;

	lut_sub lut_352 ({sk[66], n_n80, n_n86, n_n79, x168x, n_n652, x195x}, x5403x);
	defparam lut_352.LUT_SIZE = 7;
	defparam lut_352.mask = 128'h0fffffff0fffffff7f7f7f7f7f7f7fff;

	lut_sub lut_357 ({sk[67], n_n76, x297x, x129x, x193x, x5391x, n_n957}, n_n324);
	defparam lut_357.LUT_SIZE = 7;
	defparam lut_357.mask = 128'h0fffffff0fffffff7f7fffff7fffffff;

	lut_sub lut_363 ({sk[68], n_n91, x29x, x97x, n_n939, x125x, x5399x}, n_n397);
	defparam lut_363.LUT_SIZE = 7;
	defparam lut_363.mask = 128'h0fffffff0fffffff7fff7fff7fffffff;

	lut_sub lut_369 ({sk[69], x5388x, x5386x, x5387x, x5480x, x5481x}, x5487x);
	defparam lut_369.LUT_SIZE = 6;
	defparam lut_369.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_375 ({sk[70], x5421x, x5440x, x5419x, x5420x, x5438x, x5439x}, x5488x);
	defparam lut_375.LUT_SIZE = 7;
	defparam lut_375.mask = 128'h5555ffffffffffff7fffffffffffffff;

	lut_sub lut_382 ({sk[71], n_n593, n_n597, x5482x, x5483x}, x5489x);
	defparam lut_382.LUT_SIZE = 5;
	defparam lut_382.mask = 32'h0f0f7fff;

	lut_sub lut_387 ({sk[72], x278x, x159x, x300x, x5533x, x5536x}, x5539x);
	defparam lut_387.LUT_SIZE = 6;
	defparam lut_387.mask = 64'h33ff33ff7fffffff;

	lut_sub lut_393 ({sk[73], x5512x, x5510x, x5511x, x5534x, x5535x}, x5540x);
	defparam lut_393.LUT_SIZE = 6;
	defparam lut_393.mask = 64'h33ff33ff7fffffff;

	lut_sub lut_399 ({sk[74], x5580x, x5581x, x5582x, x5583x}, x5589x);
	defparam lut_399.LUT_SIZE = 5;
	defparam lut_399.mask = 32'h0f0f7fff;

	lut_sub lut_404 ({sk[75], x5556x, x5554x, x5555x, x5584x, x5585x}, x5590x);
	defparam lut_404.LUT_SIZE = 6;
	defparam lut_404.mask = 64'h33ff33ff7fffffff;

	lut_sub lut_410 ({sk[76], x5605x, x5606x, x5678x, x5679x, x5680x, x5681x}, x5685x);
	defparam lut_410.LUT_SIZE = 7;
	defparam lut_410.mask = 128'h5555ffffffffffff7fffffffffffffff;

	lut_sub lut_417 ({sk[77], x5622x, x5620x, x5621x, x5652x, x5653x}, x5658x);
	defparam lut_417.LUT_SIZE = 6;
	defparam lut_417.mask = 64'h33ff33ff7fffffff;

	lut_sub lut_423 ({sk[78], n_n91, x29x, n_n939, x162x, x91x, x266x}, x5648x);
	defparam lut_423.LUT_SIZE = 7;
	defparam lut_423.mask = 128'h5555ffffffffffff7fff7fff7fffffff;

	lut_sub lut_429 ({sk[79], x94x, x195x, x223x, x101x}, x5649x);
	defparam lut_429.LUT_SIZE = 5;
	defparam lut_429.mask = 32'h0f0f7fff;

	lut_sub lut_434 ({sk[80], n_n101, x115x, x236x, x128x, x283x, x218x}, x5650x);
	defparam lut_434.LUT_SIZE = 7;
	defparam lut_434.mask = 128'h000fffffffffffff77ffffff7fffffff;

	lut_sub lut_440 ({sk[81], n_n95, x21x, n_n1058, n_n977, n_n949, x6337x}, x5651x);
	defparam lut_440.LUT_SIZE = 7;
	defparam lut_440.mask = 128'h000fffffffffffffbfffbfffbfffffff;

	lut_sub lut_446 ({sk[82], x295x, x5716x, x5717x, x5718x, x5729x}, x5732x);
	defparam lut_446.LUT_SIZE = 6;
	defparam lut_446.mask = 64'h5f5f5f5f7fffffff;

	lut_sub lut_452 ({sk[83], x5707x, x5705x, x5706x, x5727x, x5728x}, x5733x);
	defparam lut_452.LUT_SIZE = 6;
	defparam lut_452.mask = 64'h5f5f5f5f7fffffff;

	lut_sub lut_458 ({sk[84], x5771x, x5772x, x5773x, x5774x}, x5779x);
	defparam lut_458.LUT_SIZE = 5;
	defparam lut_458.mask = 32'h0fff7fff;

	lut_sub lut_463 ({sk[85], x5748x, n_n324, x5746x, x5747x, x5775x}, x5780x);
	defparam lut_463.LUT_SIZE = 6;
	defparam lut_463.mask = 64'h5f5f5f5f7fffffff;

	lut_sub lut_469 ({sk[86], x5795x, x5793x, x5794x, x5813x, x5814x}, x5821x);
	defparam lut_469.LUT_SIZE = 6;
	defparam lut_469.mask = 64'h55ffffff7fffffff;

	lut_sub lut_475 ({sk[87], n_n397, x5815x, x5816x, x5817x}, x5822x);
	defparam lut_475.LUT_SIZE = 5;
	defparam lut_475.mask = 32'h5f5f7fff;

	lut_sub lut_480 ({sk[88], x176x, x88x, x301x, x5868x, x5869x, x5870x}, x5875x);
	defparam lut_480.LUT_SIZE = 7;
	defparam lut_480.mask = 128'h5555ffff55ffffff7fffffffffffffff;

	lut_sub lut_487 ({sk[89], n_n385, x5845x, x5843x, x5844x, x5871x}, x5876x);
	defparam lut_487.LUT_SIZE = 6;
	defparam lut_487.mask = 64'h55ffffff7fffffff;

	lut_sub lut_493 ({sk[90], n_n95, x44x, n_n980, n_n994, x149x, x6376x}, n_n206);
	defparam lut_493.LUT_SIZE = 7;
	defparam lut_493.mask = 128'h5555ffff55ffffffbfffbfffbfffffff;

	lut_sub lut_499 ({sk[91], n_n81, n_n85, n_n82, n_n241, x153x, x125x}, n_n208);
	defparam lut_499.LUT_SIZE = 7;
	defparam lut_499.mask = 128'h5555ffff55ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_504 ({sk[92], n_n93, n_n78, x57x, x86x, x100x, x6374x}, n_n201);
	defparam lut_504.LUT_SIZE = 7;
	defparam lut_504.mask = 128'h5555ffff55ffffff77777f7f77ff7fff;

	lut_sub lut_509 ({sk[93], n_n75, n_n85, x5338x, x5914x, x5916x, x6388x}, x5933x);
	defparam lut_509.LUT_SIZE = 7;
	defparam lut_509.mask = 128'h5555ffff55ffffffbfbfbfbfbfbfbfff;

	lut_sub lut_514 ({sk[94], x168x, n_n211, x5917x, x5918x, x5929x, x5930x}, x5939x);
	defparam lut_514.LUT_SIZE = 7;
	defparam lut_514.mask = 128'h5555ffff55ffffff7fffffffffffffff;

	lut_sub lut_521 ({sk[95], x5896x, x5894x, x5895x, x5931x, x5932x}, x5940x);
	defparam lut_521.LUT_SIZE = 6;
	defparam lut_521.mask = 64'h55ffffff7fffffff;

	lut_sub lut_527 ({sk[96], x5957x, n_n261, x5955x, x5956x, x6023x}, x6028x);
	defparam lut_527.LUT_SIZE = 6;
	defparam lut_527.mask = 64'h55ffffff7fffffff;

	lut_sub lut_533 ({sk[97], x5981x, x5982x, x5983x, x5984x, x5985x}, n_n243);
	defparam lut_533.LUT_SIZE = 6;
	defparam lut_533.mask = 64'h55ffffff7fffffff;

	lut_sub lut_539 ({sk[98], n_n1120, x197x, n_n944, n_n1122, n_n939, x94x}, x6019x);
	defparam lut_539.LUT_SIZE = 7;
	defparam lut_539.mask = 128'h5555ffff55ffffff7fffffffffffffff;

	lut_sub lut_546 ({sk[99], x251x, x321x, n_n1176, n_n974, x269x, x5996x}, x6020x);
	defparam lut_546.LUT_SIZE = 7;
	defparam lut_546.mask = 128'h5555ffff55ffffff7fffffffffffffff;

	lut_sub lut_553 ({sk[100], n_n91, x128x, n_n969, n_n1184, n_n1147, x6333x}, x6021x);
	defparam lut_553.LUT_SIZE = 7;
	defparam lut_553.mask = 128'h5555ffff55ffffffbfffbfffbfffffff;

	lut_sub lut_559 ({sk[101], i_2_, n_n78, n_n77, x107x, x6005x, x6015x}, x6022x);
	defparam lut_559.LUT_SIZE = 7;
	defparam lut_559.mask = 128'h5555ffff55ffffff777f777f777f77ff;

	lut_sub lut_564 ({sk[102], n_n38, n_n64, x239x, x308x, x121x, x304x}, n_n136);
	defparam lut_564.LUT_SIZE = 7;
	defparam lut_564.mask = 128'h5555ffff55ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_569 ({sk[103], n_n58, x81x, x44x, n_n1117, n_n1108, x6358x}, n_n139);
	defparam lut_569.LUT_SIZE = 7;
	defparam lut_569.mask = 128'h5555ffff55ffffffbfbfbfbfbfffffff;

	lut_sub lut_575 ({sk[104], x105x, x137x, x207x, x1442x, x1444x}, x4979x);
	defparam lut_575.LUT_SIZE = 6;
	defparam lut_575.mask = 64'h55ffffff7fffffff;

	lut_sub lut_581 ({sk[105], i_7_, i_8_, x254x, x53x, x63x, x4974x}, x4980x);
	defparam lut_581.LUT_SIZE = 7;
	defparam lut_581.mask = 128'h5555ffff55ffffff55ff77ff5fff55ff;

	lut_sub lut_586 ({sk[106], x232x, x136x, x4925x, x4926x, x4927x}, x4983x);
	defparam lut_586.LUT_SIZE = 6;
	defparam lut_586.mask = 64'h55ffffff7fffffff;

	lut_sub lut_592 ({sk[107], i_7_, i_8_, i_6_, n_n83, x64x, n_n77}, x179x);
	defparam lut_592.LUT_SIZE = 7;
	defparam lut_592.mask = 128'h5555ffff55ffffff0000000533000000;

	lut_sub lut_595 ({sk[108], i_7_, i_8_, i_6_, x26x, x23x}, x181x);
	defparam lut_595.LUT_SIZE = 6;
	defparam lut_595.mask = 64'h55ffffff00503000;

	lut_sub lut_598 ({sk[109], i_7_, i_8_, i_6_, x26x, n_n83, n_n77}, x222x);
	defparam lut_598.LUT_SIZE = 7;
	defparam lut_598.mask = 128'h5555ffff55ffffff00001100000f0000;

	lut_sub lut_601 ({sk[110], i_7_, i_8_, i_6_, n_n100, n_n84, n_n94}, x255x);
	defparam lut_601.LUT_SIZE = 7;
	defparam lut_601.mask = 128'h5555ffff55ffffff0300000000001100;

	lut_sub lut_604 ({sk[111], n_n78, x49x, n_n1369, x53x, x349x, x6354x}, x5045x);
	defparam lut_604.LUT_SIZE = 7;
	defparam lut_604.mask = 128'h5555ffff55ffffffbbffbbffbfffffff;

	lut_sub lut_610 ({sk[112], x87x, x61x, x88x, x178x, x231x, x301x}, x5046x);
	defparam lut_610.LUT_SIZE = 7;
	defparam lut_610.mask = 128'h5555ffff55ffffff7fffffffffffffff;

	lut_sub lut_617 ({sk[113], n_n73, x21x, x148x, x256x, x114x, x6353x}, x5010x);
	defparam lut_617.LUT_SIZE = 7;
	defparam lut_617.mask = 128'h5555ffff55ffffffbfffbfffbfffffff;

	lut_sub lut_623 ({sk[114], x135x, x291x, x204x, n_n978, x6372x}, x5029x);
	defparam lut_623.LUT_SIZE = 6;
	defparam lut_623.mask = 64'h55ffffffbfffffff;

	lut_sub lut_629 ({sk[115], n_n84, x32x, n_n1160, x265x, x283x, x196x}, x5008x);
	defparam lut_629.LUT_SIZE = 7;
	defparam lut_629.mask = 128'h5555ffff55ffffff7fff7fff7fffffff;

	lut_sub lut_635 ({sk[116], n_n95, x73x, n_n1022, n_n1093, n_n1128, x5005x}, x5009x);
	defparam lut_635.LUT_SIZE = 7;
	defparam lut_635.mask = 128'h5555ffff55ffffff7fff7fff7fffffff;

	lut_sub lut_641 ({sk[117], n_n95, x24x, x116x, x79x, x195x, n_n1014}, x5027x);
	defparam lut_641.LUT_SIZE = 7;
	defparam lut_641.mask = 128'h5555ffff55ffffff7fff7fff7fffffff;

	lut_sub lut_647 ({sk[118], n_n93, n_n100, n_n83, n_n77, x221x, x5024x}, x5028x);
	defparam lut_647.LUT_SIZE = 7;
	defparam lut_647.mask = 128'h5555ffff55ffffff77777777777f7f7f;

	lut_sub lut_652 ({sk[119], x87x, x61x, n_n554, x5055x, x5056x}, x5066x);
	defparam lut_652.LUT_SIZE = 6;
	defparam lut_652.mask = 64'h55ffffff7fffffff;

	lut_sub lut_658 ({sk[120], n_n91, n_n83, n_n77, x34x, x206x, x5059x}, x5064x);
	defparam lut_658.LUT_SIZE = 7;
	defparam lut_658.mask = 128'h5555ffff55ffffff777777777f7f7fff;

	lut_sub lut_663 ({sk[121], n_n73, n_n1153, x349x, n_n1267, x51x, x6352x}, x5065x);
	defparam lut_663.LUT_SIZE = 7;
	defparam lut_663.mask = 128'h5555ffff55ffffffafffffffbfffffff;

	lut_sub lut_669 ({sk[122], n_n83, x35x, x201x, x256x, x271x}, x5104x);
	defparam lut_669.LUT_SIZE = 6;
	defparam lut_669.mask = 64'h55ffffff7f7f7fff;

	lut_sub lut_674 ({sk[123], n_n86, n_n73, x39x, n_n1091, n_n1093, x6366x}, x5105x);
	defparam lut_674.LUT_SIZE = 7;
	defparam lut_674.mask = 128'h5555ffff55ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_679 ({sk[124], x106x, x197x, x5083x, x306x, x5130x}, x5139x);
	defparam lut_679.LUT_SIZE = 6;
	defparam lut_679.mask = 64'h55ffffff7fffffff;

	lut_sub lut_685 ({sk[125], i_8_, i_6_, x253x, x133x, x141x, x279x}, x5137x);
	defparam lut_685.LUT_SIZE = 7;
	defparam lut_685.mask = 128'h5555ffff55ffffff7f7f7f7f7fff7f7f;

	lut_sub lut_690 ({sk[126], n_n94, n_n74, n_n63, n_n1120, x267x, x6383x}, x5138x);
	defparam lut_690.LUT_SIZE = 7;
	defparam lut_690.mask = 128'h5555ffff55ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_695 ({sk[127], x113x, x182x, x105x, x93x}, x5160x);
	defparam lut_695.LUT_SIZE = 5;
	defparam lut_695.mask = 32'h5f5f7fff;

	lut_sub lut_700 ({sk[128], x117x, x89x, x123x, x183x}, x5161x);
	defparam lut_700.LUT_SIZE = 5;
	defparam lut_700.mask = 32'h5f5f7fff;

	lut_sub lut_705 ({sk[129], i_7_, i_6_, x233x, x51x, x5149x, x6378x}, x5164x);
	defparam lut_705.LUT_SIZE = 7;
	defparam lut_705.mask = 128'h5555ffff55ffffffbfffbbffbbffbbff;

	lut_sub lut_710 ({sk[130], i_5_, i_3_, i_4_, n_n101, n_n103, x20x}, x89x);
	defparam lut_710.LUT_SIZE = 7;
	defparam lut_710.mask = 128'h5555ffff55ffffff0000030000005500;

	lut_sub lut_713 ({sk[131], i_7_, i_8_, i_6_, x76x, n_n84, n_n90}, x183x);
	defparam lut_713.LUT_SIZE = 7;
	defparam lut_713.mask = 128'h5555ffff55ffffff00110f0000000000;

	lut_sub lut_716 ({sk[132], i_7_, i_8_, i_6_, n_n94, x40x, n_n77}, x184x);
	defparam lut_716.LUT_SIZE = 7;
	defparam lut_716.mask = 128'h5555ffff55ffffff3305000000000000;

	lut_sub lut_719 ({sk[133], i_7_, i_8_, i_6_, n_n100, n_n77, x128x}, x186x);
	defparam lut_719.LUT_SIZE = 7;
	defparam lut_719.mask = 128'h5555ffff55ffffff0300000000005500;

	lut_sub lut_722 ({sk[134], x323x, n_n1330, x185x, x258x, x5205x}, x5217x);
	defparam lut_722.LUT_SIZE = 6;
	defparam lut_722.mask = 64'h55ffffff7fffffff;

	lut_sub lut_728 ({sk[135], n_n91, x76x, n_n1279, x181x, x5206x, x6349x}, x5218x);
	defparam lut_728.LUT_SIZE = 7;
	defparam lut_728.mask = 128'h5555ffff55ffffffbfffbfffbfffffff;

	lut_sub lut_734 ({sk[136], i_7_, i_6_, x137x, x52x, x306x, x6348x}, x5185x);
	defparam lut_734.LUT_SIZE = 7;
	defparam lut_734.mask = 128'h5555ffff55ffffffbbffbbffbfffbbff;

	lut_sub lut_739 ({sk[137], n_n95, x52x, x128x, x125x, n_n1042, x6377x}, x5202x);
	defparam lut_739.LUT_SIZE = 7;
	defparam lut_739.mask = 128'h5555ffff55ffffffbfbfbfbfbfffffff;

	lut_sub lut_745 ({sk[138], n_n84, x32x, x254x, x88x, x273x, n_n1160}, x5183x);
	defparam lut_745.LUT_SIZE = 7;
	defparam lut_745.mask = 128'h5555ffff55ffffff7fff7fff7fffffff;

	lut_sub lut_751 ({sk[139], n_n91, x63x, n_n1132, n_n1130, x335x, x5179x}, x5184x);
	defparam lut_751.LUT_SIZE = 7;
	defparam lut_751.mask = 128'h5555ffff55ffffff7fff7fff7fffffff;

	lut_sub lut_757 ({sk[140], n_n93, x29x, x193x, n_n984, x195x, x274x}, x5200x);
	defparam lut_757.LUT_SIZE = 7;
	defparam lut_757.mask = 128'h5555ffff55ffffff7fff7fff7fffffff;

	lut_sub lut_763 ({sk[141], x64x, n_n95, n_n944, n_n1060, n_n1004, x6347x}, x5201x);
	defparam lut_763.LUT_SIZE = 7;
	defparam lut_763.mask = 128'h5555ffff55ffffffbfffbfffbfffffff;

	lut_sub lut_769 ({sk[142], i_8_, i_5_, i_3_, i_1_, i_0_, n_n73}, n_n1369);
	defparam lut_769.LUT_SIZE = 7;
	defparam lut_769.mask = 128'h5555ffff55ffffff0000000040000000;

	lut_sub lut_771 ({sk[143], n_n81, n_n93, n_n94, n_n95, n_n77, n_n90}, x187x);
	defparam lut_771.LUT_SIZE = 7;
	defparam lut_771.mask = 128'h5555ffff55ffffff01010101010101ff;

	lut_sub lut_774 ({sk[144], i_7_, i_8_, i_6_, n_n74, n_n90}, n_n1109);
	defparam lut_774.LUT_SIZE = 6;
	defparam lut_774.mask = 64'h55ffffff00000100;

	lut_sub lut_776 ({sk[145], i_5_, i_3_, i_4_, n_n93, n_n90}, n_n1132);
	defparam lut_776.LUT_SIZE = 6;
	defparam lut_776.mask = 64'h55ffffff00001000;

	lut_sub lut_778 ({sk[146], i_4_, i_1_, i_2_, i_0_, x28x, x5012x}, x294x);
	defparam lut_778.LUT_SIZE = 7;
	defparam lut_778.mask = 128'h5555ffff55fffffff0700000f0500000;

	lut_sub lut_782 ({sk[147], i_7_, i_8_, i_6_, n_n74, n_n96, n_n90}, x259x);
	defparam lut_782.LUT_SIZE = 7;
	defparam lut_782.mask = 128'h5555ffff55ffffff0011000000050000;

	lut_sub lut_785 ({sk[148], n_n81, n_n101, n_n102, n_n63, n_n90, x114x}, x302x);
	defparam lut_785.LUT_SIZE = 7;
	defparam lut_785.mask = 128'h5555ffff55ffffff5555557757575777;

	lut_sub lut_789 ({sk[149], i_5_, i_3_, i_4_}, n_n81);
	defparam lut_789.LUT_SIZE = 4;
	defparam lut_789.mask = 16'h7701;

	lut_sub lut_791 ({sk[150], i_7_, i_8_, i_6_}, n_n82);
	defparam lut_791.LUT_SIZE = 4;
	defparam lut_791.mask = 16'h7708;

	lut_sub lut_793 ({sk[151], i_1_, i_2_, i_0_}, n_n90);
	defparam lut_793.LUT_SIZE = 4;
	defparam lut_793.mask = 16'h7720;

	lut_sub lut_795 ({sk[152], i_7_, i_8_, i_6_, n_n84, n_n90}, n_n1294);
	defparam lut_795.LUT_SIZE = 6;
	defparam lut_795.mask = 64'h55ffffff10000000;

	lut_sub lut_797 ({sk[153], i_7_, i_8_, i_6_, n_n102, n_n90}, n_n1169);
	defparam lut_797.LUT_SIZE = 6;
	defparam lut_797.mask = 64'h55ffffff00010000;

	lut_sub lut_799 ({sk[154], n_n58, n_n91, n_n1109, x86x, n_n1125, n_n1128}, x6385x);
	defparam lut_799.LUT_SIZE = 7;
	defparam lut_799.mask = 128'h5555ffff55ffffff8800800080008000;

	lut_sub lut_802 ({sk[155], i_7_, i_8_, i_6_}, n_n58);
	defparam lut_802.LUT_SIZE = 4;
	defparam lut_802.mask = 16'h7702;

	lut_sub lut_804 ({sk[156], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x39x);
	defparam lut_804.LUT_SIZE = 7;
	defparam lut_804.mask = 128'h5555ffff55ffffff0000000800000000;

	lut_sub lut_806 ({sk[157], i_5_, i_3_, i_4_, n_n93, n_n94}, n_n941);
	defparam lut_806.LUT_SIZE = 6;
	defparam lut_806.mask = 64'h55ffffff00001000;

	lut_sub lut_808 ({sk[158], n_n52, n_n83, n_n96, x148x, x286x, x5331x}, x5335x);
	defparam lut_808.LUT_SIZE = 7;
	defparam lut_808.mask = 128'h5555ffff55ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_813 ({sk[159], x201x, x164x, x288x, x203x}, x5333x);
	defparam lut_813.LUT_SIZE = 5;
	defparam lut_813.mask = 32'h5f5f7fff;

	lut_sub lut_818 ({sk[160], x55x, n_n95, n_n1058, x156x, x5321x, x5323x}, x5334x);
	defparam lut_818.LUT_SIZE = 7;
	defparam lut_818.mask = 128'h5555ffff55ffffff7fff7fff7fffffff;

	lut_sub lut_824 ({sk[161], n_n70, x232x, n_n79, n_n53, x319x, x5352x}, x5367x);
	defparam lut_824.LUT_SIZE = 7;
	defparam lut_824.mask = 128'h5555ffff55ffffff7777ffff777fffff;

	lut_sub lut_829 ({sk[162], x197x, x5083x, x168x, x291x, x297x}, x5368x);
	defparam lut_829.LUT_SIZE = 6;
	defparam lut_829.mask = 64'h55ffffff7fffffff;

	lut_sub lut_835 ({sk[163], x310x, x5406x, x5407x, x5595x, x5596x}, x5605x);
	defparam lut_835.LUT_SIZE = 6;
	defparam lut_835.mask = 64'h55ffffff7fffffff;

	lut_sub lut_841 ({sk[164], x123x, x95x, x217x, x122x, x5597x, x5600x}, x5606x);
	defparam lut_841.LUT_SIZE = 7;
	defparam lut_841.mask = 128'h5555ffff55ffffff7fffffffffffffff;

	lut_sub lut_848 ({sk[165], n_n100, n_n96, n_n95, x81x, n_n211, x120x}, x5678x);
	defparam lut_848.LUT_SIZE = 7;
	defparam lut_848.mask = 128'h5555ffff55ffffff777f777f777f77ff;

	lut_sub lut_853 ({sk[166], n_n84, x32x, n_n1160, x191x, x264x, x265x}, x5679x);
	defparam lut_853.LUT_SIZE = 7;
	defparam lut_853.mask = 128'h5555ffff55ffffff7fff7fff7fffffff;

	lut_sub lut_859 ({sk[167], n_n95, x67x, n_n1169, n_n1145, x5664x, x6381x}, x5680x);
	defparam lut_859.LUT_SIZE = 7;
	defparam lut_859.mask = 128'h5555ffff55ffffffbfffbfffbfffffff;

	lut_sub lut_865 ({sk[168], n_n554, x5668x, x5669x, x5670x}, x5681x);
	defparam lut_865.LUT_SIZE = 5;
	defparam lut_865.mask = 32'h5f5f7fff;

	lut_sub lut_870 ({sk[169], n_n95, x34x, x167x, x287x, x6369x}, x5957x);
	defparam lut_870.LUT_SIZE = 6;
	defparam lut_870.mask = 64'h55ffffffbfbfbfff;

	lut_sub lut_875 ({sk[170], x64x, n_n95, x237x, x163x, n_n296, x284x}, n_n261);
	defparam lut_875.LUT_SIZE = 7;
	defparam lut_875.mask = 128'h5555ffff55ffffff7f7f7fff7f7fffff;

	lut_sub lut_881 ({sk[171], n_n95, x24x, x274x, n_n1014, x98x, x154x}, x5955x);
	defparam lut_881.LUT_SIZE = 7;
	defparam lut_881.mask = 128'h5555ffff55ffffff7fff7fff7fffffff;

	lut_sub lut_887 ({sk[172], n_n1057, n_n1087, x66x, x5442x, n_n1013, x5951x}, x5956x);
	defparam lut_887.LUT_SIZE = 7;
	defparam lut_887.mask = 128'h5555ffff55ffffff777fffffffffffff;

	lut_sub lut_893 ({sk[173], x150x, x153x, x125x, n_n652, x6007x}, x6023x);
	defparam lut_893.LUT_SIZE = 6;
	defparam lut_893.mask = 64'h55ffffff7fffffff;

	lut_sub lut_899 ({sk[174], i_3_, i_2_, i_0_}, n_n80);
	defparam lut_899.LUT_SIZE = 4;
	defparam lut_899.mask = 16'h7740;

	lut_sub lut_901 ({sk[175], i_7_, i_8_}, n_n75);
	defparam lut_901.LUT_SIZE = 3;
	defparam lut_901.mask = 8'h54;

	lut_sub lut_903 ({sk[176], i_7_, i_6_}, n_n38);
	defparam lut_903.LUT_SIZE = 3;
	defparam lut_903.mask = 8'h52;

	lut_sub lut_905 ({sk[177], i_7_, i_8_}, n_n64);
	defparam lut_905.LUT_SIZE = 3;
	defparam lut_905.mask = 8'h51;

	lut_sub lut_907 ({sk[178], i_7_, i_6_}, n_n52);
	defparam lut_907.LUT_SIZE = 3;
	defparam lut_907.mask = 8'h51;

	lut_sub lut_909 ({sk[179], i_8_, i_6_}, x77x);
	defparam lut_909.LUT_SIZE = 3;
	defparam lut_909.mask = 8'h54;

	lut_sub lut_911 ({sk[180], i_7_, i_8_, i_6_}, n_n101);
	defparam lut_911.LUT_SIZE = 4;
	defparam lut_911.mask = 16'h7704;

	lut_sub lut_913 ({sk[181], i_7_, i_8_}, n_n86);
	defparam lut_913.LUT_SIZE = 3;
	defparam lut_913.mask = 8'h58;

	lut_sub lut_915 ({sk[182], i_7_, i_8_, i_6_}, n_n93);
	defparam lut_915.LUT_SIZE = 4;
	defparam lut_915.mask = 16'h7740;

	lut_sub lut_917 ({sk[183], i_7_, i_6_}, n_n73);
	defparam lut_917.LUT_SIZE = 3;
	defparam lut_917.mask = 8'h58;

	lut_sub lut_919 ({sk[184], i_7_, i_8_, i_6_}, n_n78);
	defparam lut_919.LUT_SIZE = 4;
	defparam lut_919.mask = 16'h7780;

	lut_sub lut_921 ({sk[185], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x76x);
	defparam lut_921.LUT_SIZE = 7;
	defparam lut_921.mask = 128'h5555ffff55ffffff0200000000000000;

	lut_sub lut_923 ({sk[186], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x27x);
	defparam lut_923.LUT_SIZE = 7;
	defparam lut_923.mask = 128'h5555ffff55ffffff0000400000000000;

	lut_sub lut_925 ({sk[187], i_1_, i_2_, i_0_}, n_n100);
	defparam lut_925.LUT_SIZE = 4;
	defparam lut_925.mask = 16'h7740;

	lut_sub lut_927 ({sk[188], i_7_, i_8_, i_6_, n_n100, n_n74}, n_n1134);
	defparam lut_927.LUT_SIZE = 6;
	defparam lut_927.mask = 64'h55ffffff00000010;

	lut_sub lut_929 ({sk[189], i_7_, i_8_, i_3_, i_2_, i_0_, n_n87}, n_n1091);
	defparam lut_929.LUT_SIZE = 7;
	defparam lut_929.mask = 128'h5555ffff55ffffff0000000000000010;

	lut_sub lut_931 ({sk[190], i_7_, i_8_, i_5_, i_6_, i_4_}, x240x);
	defparam lut_931.LUT_SIZE = 6;
	defparam lut_931.mask = 64'h55ffffff00000800;

	lut_sub lut_933 ({sk[191], i_7_, i_8_, i_6_, x42x}, n_n1164);
	defparam lut_933.LUT_SIZE = 5;
	defparam lut_933.mask = 32'h5f5f1000;

	lut_sub lut_935 ({sk[192], i_5_, i_3_, i_4_, n_n85, n_n82}, n_n1021);
	defparam lut_935.LUT_SIZE = 6;
	defparam lut_935.mask = 64'h55ffffff00001000;

	lut_sub lut_937 ({sk[193], n_n100, n_n1134, n_n1091, x240x, n_n1164, n_n1021}, x4839x);
	defparam lut_937.LUT_SIZE = 7;
	defparam lut_937.mask = 128'h5555ffff55ffffff77ffffff7fffffff;

	lut_sub lut_943 ({sk[194], i_5_, i_3_, i_4_, n_n83, n_n95}, n_n1120);
	defparam lut_943.LUT_SIZE = 6;
	defparam lut_943.mask = 64'h55ffffff00000010;

	lut_sub lut_945 ({sk[195], i_7_, i_8_, i_6_, x42x}, n_n956);
	defparam lut_945.LUT_SIZE = 5;
	defparam lut_945.mask = 32'h5f5f4000;

	lut_sub lut_947 ({sk[196], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x128x);
	defparam lut_947.LUT_SIZE = 7;
	defparam lut_947.mask = 128'h03ff57ffffffffff0800000000000000;

	lut_sub lut_949 ({sk[197], i_7_, i_5_, i_6_, i_3_, i_4_, n_n83}, x355x);
	defparam lut_949.LUT_SIZE = 7;
	defparam lut_949.mask = 128'h03ff57ffffffffff0000010000000000;

	lut_sub lut_951 ({sk[198], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x57x);
	defparam lut_951.LUT_SIZE = 7;
	defparam lut_951.mask = 128'h03ff57ffffffffff0100000000000000;

	lut_sub lut_953 ({sk[199], i_1_, i_2_, i_0_}, n_n103);
	defparam lut_953.LUT_SIZE = 4;
	defparam lut_953.mask = 16'h7702;

	lut_sub lut_955 ({sk[200], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x26x);
	defparam lut_955.LUT_SIZE = 7;
	defparam lut_955.mask = 128'h03ff57ffffffffff0000000000000200;

	lut_sub lut_957 ({sk[201], i_5_, i_3_, i_4_}, n_n84);
	defparam lut_957.LUT_SIZE = 4;
	defparam lut_957.mask = 16'h7720;

	lut_sub lut_959 ({sk[202], i_1_, i_2_, i_0_}, n_n83);
	defparam lut_959.LUT_SIZE = 4;
	defparam lut_959.mask = 16'h7710;

	lut_sub lut_961 ({sk[203], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x32x);
	defparam lut_961.LUT_SIZE = 7;
	defparam lut_961.mask = 128'h03ff57ffffffffff0000001000000000;

	lut_sub lut_963 ({sk[204], i_5_, i_3_, i_4_}, n_n102);
	defparam lut_963.LUT_SIZE = 4;
	defparam lut_963.mask = 16'h7710;

	lut_sub lut_965 ({sk[205], i_1_, i_2_, i_0_}, n_n94);
	defparam lut_965.LUT_SIZE = 4;
	defparam lut_965.mask = 16'h7708;

	lut_sub lut_967 ({sk[206], i_5_, i_3_, i_4_}, n_n74);
	defparam lut_967.LUT_SIZE = 4;
	defparam lut_967.mask = 16'h7740;

	lut_sub lut_969 ({sk[207], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x40x);
	defparam lut_969.LUT_SIZE = 7;
	defparam lut_969.mask = 128'h03ff57ffffffffff0001000000000000;

	lut_sub lut_971 ({sk[208], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x45x);
	defparam lut_971.LUT_SIZE = 7;
	defparam lut_971.mask = 128'h03ff57ffffffffff0000000000004000;

	lut_sub lut_973 ({sk[209], i_5_, i_3_, i_4_}, n_n96);
	defparam lut_973.LUT_SIZE = 4;
	defparam lut_973.mask = 16'h7708;

	lut_sub lut_975 ({sk[210], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x55x);
	defparam lut_975.LUT_SIZE = 7;
	defparam lut_975.mask = 128'h03ff57ffffffffff0000000008000000;

	lut_sub lut_977 ({sk[211], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x58x);
	defparam lut_977.LUT_SIZE = 7;
	defparam lut_977.mask = 128'h03ff57ffffffffff0000001000000000;

	lut_sub lut_979 ({sk[212], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x64x);
	defparam lut_979.LUT_SIZE = 7;
	defparam lut_979.mask = 128'h03ff57ffffffffff0040000000000000;

	lut_sub lut_981 ({sk[213], i_1_, i_2_}, x75x);
	defparam lut_981.LUT_SIZE = 3;
	defparam lut_981.mask = 8'h54;

	lut_sub lut_983 ({sk[214], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x171x);
	defparam lut_983.LUT_SIZE = 7;
	defparam lut_983.mask = 128'h03ff57ffffffffff0000000000010000;

	lut_sub lut_985 ({sk[215], i_7_, i_8_, i_6_, n_n103, n_n74, x171x}, x87x);
	defparam lut_985.LUT_SIZE = 7;
	defparam lut_985.mask = 128'h03ff57ffffffffff5500550000030000;

	lut_sub lut_988 ({sk[216], i_5_, i_3_, i_4_}, n_n77);
	defparam lut_988.LUT_SIZE = 4;
	defparam lut_988.mask = 16'h7704;

	lut_sub lut_990 ({sk[217], i_7_, i_8_, i_6_, n_n100, x45x, n_n77}, x104x);
	defparam lut_990.LUT_SIZE = 7;
	defparam lut_990.mask = 128'h03ff57ffffffffff0000000500000033;

	lut_sub lut_993 ({sk[218], i_7_, i_8_, i_5_, i_6_, i_4_}, x318x);
	defparam lut_993.LUT_SIZE = 6;
	defparam lut_993.mask = 64'h11ffffff40000000;

	lut_sub lut_995 ({sk[219], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x63x);
	defparam lut_995.LUT_SIZE = 7;
	defparam lut_995.mask = 128'h03ff57ffffffffff0000000002000000;

	lut_sub lut_997 ({sk[220], i_3_, i_1_, i_0_, n_n101, x318x, x63x}, x113x);
	defparam lut_997.LUT_SIZE = 7;
	defparam lut_997.mask = 128'h03ff57ffffffffff0505050505370505;

	lut_sub lut_1000 ({sk[221], i_7_, i_8_}, n_n70);
	defparam lut_1000.LUT_SIZE = 3;
	defparam lut_1000.mask = 8'h52;

	lut_sub lut_1002 ({sk[222], i_7_, i_8_, i_6_}, n_n95);
	defparam lut_1002.LUT_SIZE = 4;
	defparam lut_1002.mask = 16'h7701;

	lut_sub lut_1004 ({sk[223], i_5_, i_4_}, x109x);
	defparam lut_1004.LUT_SIZE = 3;
	defparam lut_1004.mask = 8'h52;

	lut_sub lut_1006 ({sk[224], i_3_, n_n93, x57x, n_n83, n_n95, x109x}, x176x);
	defparam lut_1006.LUT_SIZE = 7;
	defparam lut_1006.mask = 128'h03ff57ffffffffff0033003300330537;

	lut_sub lut_1009 ({sk[225], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x34x);
	defparam lut_1009.LUT_SIZE = 7;
	defparam lut_1009.mask = 128'h03ff57ffffffffff0400000000000000;

	lut_sub lut_1011 ({sk[226], i_7_, i_8_, i_6_, n_n100, n_n84, x34x}, x182x);
	defparam lut_1011.LUT_SIZE = 7;
	defparam lut_1011.mask = 128'h03ff57ffffffffff0000550000000003;

	lut_sub lut_1014 ({sk[227], i_7_, i_8_, i_6_}, n_n63);
	defparam lut_1014.LUT_SIZE = 4;
	defparam lut_1014.mask = 16'h7720;

	lut_sub lut_1016 ({sk[228], i_7_, i_8_, i_6_}, x192x);
	defparam lut_1016.LUT_SIZE = 4;
	defparam lut_1016.mask = 16'h7724;

	lut_sub lut_1019 ({sk[229], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x74x);
	defparam lut_1019.LUT_SIZE = 7;
	defparam lut_1019.mask = 128'h03ff57ffffffffff0002000000000000;

	lut_sub lut_1021 ({sk[230], i_7_, i_8_, i_6_, n_n81, n_n94, x74x}, x208x);
	defparam lut_1021.LUT_SIZE = 7;
	defparam lut_1021.mask = 128'h03ff57ffffffffff0003000000000055;

	lut_sub lut_1024 ({sk[231], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x42x);
	defparam lut_1024.LUT_SIZE = 7;
	defparam lut_1024.mask = 128'h03ff57ffffffffff0000000001000000;

	lut_sub lut_1026 ({sk[232], i_7_, i_8_, i_6_, i_3_, n_n103, x109x}, x252x);
	defparam lut_1026.LUT_SIZE = 7;
	defparam lut_1026.mask = 128'h03ff57ffffffffff0001000000000000;

	lut_sub lut_1028 ({sk[233], i_1_, i_2_, i_0_}, n_n85);
	defparam lut_1028.LUT_SIZE = 4;
	defparam lut_1028.mask = 16'h7704;

	lut_sub lut_1030 ({sk[234], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x253x);
	defparam lut_1030.LUT_SIZE = 7;
	defparam lut_1030.mask = 128'h03ff57ffffffffff0000000000000004;

	lut_sub lut_1032 ({sk[235], i_6_, i_3_, i_1_, i_2_, i_0_}, x311x);
	defparam lut_1032.LUT_SIZE = 6;
	defparam lut_1032.mask = 64'h11ffffff00400000;

	lut_sub lut_1034 ({sk[236], i_7_, i_8_, i_6_, n_n81, n_n103}, x329x);
	defparam lut_1034.LUT_SIZE = 6;
	defparam lut_1034.mask = 64'h11ffffff00000100;

	lut_sub lut_1036 ({sk[237], i_7_, i_8_, i_5_, i_6_, i_4_}, x337x);
	defparam lut_1036.LUT_SIZE = 6;
	defparam lut_1036.mask = 64'h11ffffff00080000;

	lut_sub lut_1038 ({sk[238], i_7_, i_8_, i_6_, n_n100, n_n74}, n_n1077);
	defparam lut_1038.LUT_SIZE = 6;
	defparam lut_1038.mask = 64'h11ffffff00010000;

	lut_sub lut_1040 ({sk[239], i_7_, i_8_, i_6_, n_n71, x23x, n_n67}, x4888x);
	defparam lut_1040.LUT_SIZE = 7;
	defparam lut_1040.mask = 128'h03ff57ffffffffff0000000500330033;

	lut_sub lut_1043 ({sk[240], n_n38, x201x, x22x, x324x, x164x, x327x}, x4896x);
	defparam lut_1043.LUT_SIZE = 7;
	defparam lut_1043.mask = 128'h03ff57ffffffffff3737ffff37ffffff;

	lut_sub lut_1048 ({sk[241], n_n96, n_n85, n_n95, x34x, x4888x, x4896x}, x4899x);
	defparam lut_1048.LUT_SIZE = 7;
	defparam lut_1048.mask = 128'h03ff57ffffffffff777f777f777f77ff;

	lut_sub lut_1053 ({sk[242], i_7_, i_8_, i_5_, i_6_, i_4_}, x234x);
	defparam lut_1053.LUT_SIZE = 6;
	defparam lut_1053.mask = 64'h11ffffff00002000;

	lut_sub lut_1055 ({sk[243], i_7_, i_8_, n_n85, n_n76, x146x}, x298x);
	defparam lut_1055.LUT_SIZE = 6;
	defparam lut_1055.mask = 64'h11ffffff55575555;

	lut_sub lut_1058 ({sk[244], i_5_, i_3_, i_4_, n_n103, n_n82, x4901x}, x116x);
	defparam lut_1058.LUT_SIZE = 7;
	defparam lut_1058.mask = 128'h03ff57ffffffffff0003550000000000;

	lut_sub lut_1061 ({sk[245], i_7_, i_8_, i_6_, n_n100, n_n74, x221x}, n_n882);
	defparam lut_1061.LUT_SIZE = 7;
	defparam lut_1061.mask = 128'h03ff57ffffffffff5555555555555557;

	lut_sub lut_1064 ({sk[246], i_7_, i_0_, n_n80, n_n93, n_n77, x49x}, x4910x);
	defparam lut_1064.LUT_SIZE = 7;
	defparam lut_1064.mask = 128'h03ff57ffffffffff0505050505053705;

	lut_sub lut_1067 ({sk[247], n_n80, x234x, x298x, x116x, n_n882, x4910x}, x4919x);
	defparam lut_1067.LUT_SIZE = 7;
	defparam lut_1067.mask = 128'h03ff57ffffffffff7fff7fff7fffffff;

	lut_sub lut_1073 ({sk[248], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x73x);
	defparam lut_1073.LUT_SIZE = 7;
	defparam lut_1073.mask = 128'h03ff57ffffffffff0000000000000020;

	lut_sub lut_1075 ({sk[249], i_7_, i_8_, i_6_, n_n81, n_n90}, n_n1172);
	defparam lut_1075.LUT_SIZE = 6;
	defparam lut_1075.mask = 64'h11ffffff00000001;

	lut_sub lut_1077 ({sk[250], i_7_, i_8_, i_6_, x57x}, n_n1078);
	defparam lut_1077.LUT_SIZE = 5;
	defparam lut_1077.mask = 32'h0f0f4000;

	lut_sub lut_1079 ({sk[251], i_3_, i_2_, i_0_}, x245x);
	defparam lut_1079.LUT_SIZE = 4;
	defparam lut_1079.mask = 16'h7701;

	lut_sub lut_1081 ({sk[252], i_7_, i_8_, i_5_, i_6_, i_4_}, x38x);
	defparam lut_1081.LUT_SIZE = 6;
	defparam lut_1081.mask = 64'h11ffffff00000008;

	lut_sub lut_1083 ({sk[253], i_6_, i_3_, i_2_, i_0_, n_n64, x109x}, n_n1081);
	defparam lut_1083.LUT_SIZE = 7;
	defparam lut_1083.mask = 128'h03ff57ffffffffff0000000100000000;

	lut_sub lut_1085 ({sk[254], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x43x);
	defparam lut_1085.LUT_SIZE = 7;
	defparam lut_1085.mask = 128'h03ff57ffffffffff0020000000000000;

	lut_sub lut_1087 ({sk[255], i_7_, i_8_, i_6_, n_n74, n_n90}, n_n1279);
	defparam lut_1087.LUT_SIZE = 6;
	defparam lut_1087.mask = 64'h11ffffff10000000;

	lut_sub lut_1089 ({sk[256], i_7_, i_8_, i_6_, x29x, x23x}, x61x);
	defparam lut_1089.LUT_SIZE = 6;
	defparam lut_1089.mask = 64'h11ffffff00350000;

	lut_sub lut_1092 ({sk[257], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x22x);
	defparam lut_1092.LUT_SIZE = 7;
	defparam lut_1092.mask = 128'h03ff57ffffffffff0000020000000000;

	lut_sub lut_1094 ({sk[258], i_3_, i_1_, i_2_, n_n78, x52x, x339x}, x118x);
	defparam lut_1094.LUT_SIZE = 7;
	defparam lut_1094.mask = 128'h03ff57ffffffffff0303030303030357;

	lut_sub lut_1097 ({sk[259], i_7_, i_8_, i_6_, x39x, x239x, x81x}, x295x);
	defparam lut_1097.LUT_SIZE = 7;
	defparam lut_1097.mask = 128'h03ff57ffffffffff0000000f00000077;

	lut_sub lut_1101 ({sk[260], n_n78, x55x, x61x, x22x, x118x, x295x}, n_n137);
	defparam lut_1101.LUT_SIZE = 7;
	defparam lut_1101.mask = 128'h03ff57ffffffffff77ff77ff7fffffff;

	lut_sub lut_1107 ({sk[261], i_3_, i_1_, i_0_, x38x, x99x}, x231x);
	defparam lut_1107.LUT_SIZE = 6;
	defparam lut_1107.mask = 64'h11ffffff55575555;

	lut_sub lut_1110 ({sk[262], i_7_, i_8_, i_6_, i_4_, x311x, x46x}, x4933x);
	defparam lut_1110.LUT_SIZE = 7;
	defparam lut_1110.mask = 128'h03ff57ffffffffff0000035700000000;

	lut_sub lut_1113 ({sk[263], i_1_, i_0_, n_n93, n_n102, x354x, x62x}, x4934x);
	defparam lut_1113.LUT_SIZE = 7;
	defparam lut_1113.mask = 128'h03ff57ffffffffff11111111111f1111;

	lut_sub lut_1116 ({sk[264], i_7_, i_8_, i_6_, n_n81, n_n103, n_n77}, x4935x);
	defparam lut_1116.LUT_SIZE = 7;
	defparam lut_1116.mask = 128'h03ff57ffffffffff0011030300000000;

	lut_sub lut_1119 ({sk[265], x231x, x4933x, x4934x, x4935x}, n_n135);
	defparam lut_1119.LUT_SIZE = 5;
	defparam lut_1119.mask = 32'h0f0f7fff;

	lut_sub lut_1124 ({sk[266], i_5_, i_4_}, x325x);
	defparam lut_1124.LUT_SIZE = 3;
	defparam lut_1124.mask = 8'h54;

	lut_sub lut_1126 ({sk[267], i_7_, i_8_, i_6_, n_n102, n_n90}, n_n1153);
	defparam lut_1126.LUT_SIZE = 6;
	defparam lut_1126.mask = 64'h11ffffff00000010;

	lut_sub lut_1128 ({sk[268], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x239x);
	defparam lut_1128.LUT_SIZE = 7;
	defparam lut_1128.mask = 128'h03ff57ffffffffff0000000040000000;

	lut_sub lut_1130 ({sk[269], i_7_, i_8_, n_n84, n_n85, x46x, n_n87}, x308x);
	defparam lut_1130.LUT_SIZE = 7;
	defparam lut_1130.mask = 128'h03ff57ffffffffff000f050533330000;

	lut_sub lut_1134 ({sk[270], i_5_, i_3_, n_n75, n_n83, n_n66, x20x}, x121x);
	defparam lut_1134.LUT_SIZE = 7;
	defparam lut_1134.mask = 128'h03ff57ffffffffff0003000355570003;

	lut_sub lut_1137 ({sk[271], n_n101, x57x, n_n100, n_n77, x349x}, x304x);
	defparam lut_1137.LUT_SIZE = 6;
	defparam lut_1137.mask = 64'h11ffffff555557ff;

	lut_sub lut_1141 ({sk[272], i_5_, i_3_, i_4_, n_n95, n_n90}, n_n1297);
	defparam lut_1141.LUT_SIZE = 6;
	defparam lut_1141.mask = 64'h11ffffff00001000;

	lut_sub lut_1143 ({sk[273], i_7_, i_8_, i_6_, n_n102, n_n90}, n_n1324);
	defparam lut_1143.LUT_SIZE = 6;
	defparam lut_1143.mask = 64'h11ffffff01000000;

	lut_sub lut_1145 ({sk[274], i_7_, i_8_, i_6_, n_n100, n_n84}, n_n1092);
	defparam lut_1145.LUT_SIZE = 6;
	defparam lut_1145.mask = 64'h11ffffff00010000;

	lut_sub lut_1147 ({sk[275], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x81x);
	defparam lut_1147.LUT_SIZE = 7;
	defparam lut_1147.mask = 128'h03ff57ffffffffff0000000000000008;

	lut_sub lut_1149 ({sk[276], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x44x);
	defparam lut_1149.LUT_SIZE = 7;
	defparam lut_1149.mask = 128'h03ff57ffffffffff0000040000000000;

	lut_sub lut_1151 ({sk[277], i_7_, i_8_, i_1_, i_2_, i_0_, x354x}, n_n1117);
	defparam lut_1151.LUT_SIZE = 7;
	defparam lut_1151.mask = 128'h03ff57ffffffffff0000000000400000;

	lut_sub lut_1153 ({sk[278], i_7_, i_8_, i_6_, n_n81, n_n90}, n_n1108);
	defparam lut_1153.LUT_SIZE = 6;
	defparam lut_1153.mask = 64'h11ffffff01000000;

	lut_sub lut_1155 ({sk[279], x58x, n_n63, n_n95, x319x, x44x, x94x}, x6358x);
	defparam lut_1155.LUT_SIZE = 7;
	defparam lut_1155.mask = 128'h03ff57ffffffffffa0a08080a0008000;

	lut_sub lut_1160 ({sk[280], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x19x);
	defparam lut_1160.LUT_SIZE = 7;
	defparam lut_1160.mask = 128'h03ff57ffffffffff0000000000020000;

	lut_sub lut_1162 ({sk[281], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x29x);
	defparam lut_1162.LUT_SIZE = 7;
	defparam lut_1162.mask = 128'h03ff57ffffffffff0000000100000000;

	lut_sub lut_1164 ({sk[282], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x37x);
	defparam lut_1164.LUT_SIZE = 7;
	defparam lut_1164.mask = 128'h03ff57ffffffffff0000000008000000;

	lut_sub lut_1166 ({sk[283], i_1_, i_2_, i_0_, n_n81, n_n91, n_n74}, x105x);
	defparam lut_1166.LUT_SIZE = 7;
	defparam lut_1166.mask = 128'h03ff57ffffffffff0003001100000000;

	lut_sub lut_1169 ({sk[284], i_1_, i_0_}, x108x);
	defparam lut_1169.LUT_SIZE = 3;
	defparam lut_1169.mask = 8'h51;

	lut_sub lut_1171 ({sk[285], i_6_, i_3_, i_4_}, x127x);
	defparam lut_1171.LUT_SIZE = 4;
	defparam lut_1171.mask = 16'h7704;

	lut_sub lut_1173 ({sk[286], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x21x);
	defparam lut_1173.LUT_SIZE = 7;
	defparam lut_1173.mask = 128'h03ff57ffffffffff1000000000000000;

	lut_sub lut_1175 ({sk[287], i_7_, i_8_, i_6_, x40x, x21x}, x137x);
	defparam lut_1175.LUT_SIZE = 6;
	defparam lut_1175.mask = 64'h11ffffff50700000;

	lut_sub lut_1178 ({sk[288], i_7_, i_8_, i_6_, n_n84, x55x, n_n90}, x207x);
	defparam lut_1178.LUT_SIZE = 7;
	defparam lut_1178.mask = 128'h03ff57ffffffffff0000333305000500;

	lut_sub lut_1181 ({sk[289], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x35x);
	defparam lut_1181.LUT_SIZE = 7;
	defparam lut_1181.mask = 128'h03ff57ffffffffff0000500000800080;

	lut_sub lut_1184 ({sk[290], i_7_, i_6_, n_n103, n_n83, n_n102, x35x}, x106x);
	defparam lut_1184.LUT_SIZE = 7;
	defparam lut_1184.mask = 128'h03ff57ffffffffff0505050505370505;

	lut_sub lut_1187 ({sk[291], i_3_, i_1_, i_0_}, n_n67);
	defparam lut_1187.LUT_SIZE = 4;
	defparam lut_1187.mask = 16'h7740;

	lut_sub lut_1189 ({sk[292], i_7_, i_8_, i_6_, i_4_, x106x, n_n67}, x232x);
	defparam lut_1189.LUT_SIZE = 7;
	defparam lut_1189.mask = 128'h03ff57ffffffffff3373333333333333;

	lut_sub lut_1192 ({sk[293], i_7_, i_8_, i_6_, n_n103, n_n77}, x251x);
	defparam lut_1192.LUT_SIZE = 6;
	defparam lut_1192.mask = 64'h11ffffff00100000;

	lut_sub lut_1194 ({sk[294], i_5_, i_3_, i_4_, n_n93, n_n94}, n_n1070);
	defparam lut_1194.LUT_SIZE = 6;
	defparam lut_1194.mask = 64'h11ffffff10000000;

	lut_sub lut_1196 ({sk[295], i_5_, i_3_, i_4_, n_n93, n_n100, n_n94}, x254x);
	defparam lut_1196.LUT_SIZE = 7;
	defparam lut_1196.mask = 128'h03ff57ffffffffff0500000000000003;

	lut_sub lut_1199 ({sk[296], i_7_, i_8_, i_6_, x40x}, x321x);
	defparam lut_1199.LUT_SIZE = 5;
	defparam lut_1199.mask = 32'h0f0f0010;

	lut_sub lut_1201 ({sk[297], i_7_, i_8_, i_1_, i_2_, i_0_}, x328x);
	defparam lut_1201.LUT_SIZE = 6;
	defparam lut_1201.mask = 64'h11ffffff00000001;

	lut_sub lut_1203 ({sk[298], i_1_, i_2_}, x338x);
	defparam lut_1203.LUT_SIZE = 3;
	defparam lut_1203.mask = 8'h51;

	lut_sub lut_1205 ({sk[299], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x49x);
	defparam lut_1205.LUT_SIZE = 7;
	defparam lut_1205.mask = 128'h03ff57ffffffffff0000000000002000;

	lut_sub lut_1207 ({sk[300], i_5_, i_3_, i_4_, n_n100, n_n95}, n_n1204);
	defparam lut_1207.LUT_SIZE = 6;
	defparam lut_1207.mask = 64'h11ffffff00001000;

	lut_sub lut_1209 ({sk[301], i_7_, i_8_, i_6_, n_n96, n_n85, x43x}, x148x);
	defparam lut_1209.LUT_SIZE = 7;
	defparam lut_1209.mask = 128'h03ff57ffffffffff0055000000000003;

	lut_sub lut_1212 ({sk[302], i_7_, i_8_, i_6_, n_n102, n_n94, n_n96}, x256x);
	defparam lut_1212.LUT_SIZE = 7;
	defparam lut_1212.mask = 128'h03ff57ffffffffff0000030000001100;

	lut_sub lut_1215 ({sk[303], n_n91, x26x, n_n102, x83x, x20x, n_n1181}, x6353x);
	defparam lut_1215.LUT_SIZE = 7;
	defparam lut_1215.mask = 128'h03ff57ffffffffffaa88aa88a0800000;

	lut_sub lut_1220 ({sk[304], i_6_, i_3_, i_4_, i_1_, i_2_, i_0_}, x135x);
	defparam lut_1220.LUT_SIZE = 7;
	defparam lut_1220.mask = 128'h03ff57ffffffffffa080808080808080;

	lut_sub lut_1223 ({sk[305], i_7_, i_8_, i_6_, n_n84, n_n85, x97x}, x291x);
	defparam lut_1223.LUT_SIZE = 7;
	defparam lut_1223.mask = 128'h03ff57ffffffffff5555555555575555;

	lut_sub lut_1226 ({sk[306], i_5_, i_3_, i_4_, n_n103, n_n95, x317x}, x204x);
	defparam lut_1226.LUT_SIZE = 7;
	defparam lut_1226.mask = 128'h03ff57ffffffffff0000000300005500;

	lut_sub lut_1229 ({sk[307], i_5_, i_3_, i_4_, n_n83, n_n63}, n_n978);
	defparam lut_1229.LUT_SIZE = 6;
	defparam lut_1229.mask = 64'h11ffffff00000010;

	lut_sub lut_1231 ({sk[308], n_n81, n_n52, n_n103, n_n82, x23x, n_n1021}, x6372x);
	defparam lut_1231.LUT_SIZE = 7;
	defparam lut_1231.mask = 128'h03ff57ffffffffffaaaa8888aaa08880;

	lut_sub lut_1238 ({sk[309], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x23x);
	defparam lut_1238.LUT_SIZE = 7;
	defparam lut_1238.mask = 128'h03ff57ffffffffff0000000000000001;

	lut_sub lut_1240 ({sk[310], i_7_, i_8_, i_6_, n_n81, x40x, n_n90}, x88x);
	defparam lut_1240.LUT_SIZE = 7;
	defparam lut_1240.mask = 128'h03ff57ffffffffff0033000000000500;

	lut_sub lut_1243 ({sk[311], i_7_, i_8_, i_6_, n_n100, n_n77, x34x}, x99x);
	defparam lut_1243.LUT_SIZE = 7;
	defparam lut_1243.mask = 128'h03ff57ffffffffff0000000055000300;

	lut_sub lut_1246 ({sk[312], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x46x);
	defparam lut_1246.LUT_SIZE = 7;
	defparam lut_1246.mask = 128'h03ff57ffffffffff0000000000000400;

	lut_sub lut_1248 ({sk[313], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x41x);
	defparam lut_1248.LUT_SIZE = 7;
	defparam lut_1248.mask = 128'h03ff57ffffffffff0000004000000000;

	lut_sub lut_1250 ({sk[314], i_7_, i_8_, i_6_, x21x, x46x, x41x}, x301x);
	defparam lut_1250.LUT_SIZE = 7;
	defparam lut_1250.mask = 128'h03ff57ffffffffff0055000f00000033;

	lut_sub lut_1254 ({sk[315], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x53x);
	defparam lut_1254.LUT_SIZE = 7;
	defparam lut_1254.mask = 128'h03ff57ffffffffff0000000400000000;

	lut_sub lut_1256 ({sk[316], i_7_, i_8_, i_6_, n_n81, n_n103}, x349x);
	defparam lut_1256.LUT_SIZE = 6;
	defparam lut_1256.mask = 64'h11ffffff00000010;

	lut_sub lut_1258 ({sk[317], i_7_, i_8_, i_6_, n_n102, n_n85}, n_n1022);
	defparam lut_1258.LUT_SIZE = 6;
	defparam lut_1258.mask = 64'h11ffffff00000010;

	lut_sub lut_1260 ({sk[318], i_7_, i_8_, i_6_, n_n102, n_n94}, n_n1039);
	defparam lut_1260.LUT_SIZE = 6;
	defparam lut_1260.mask = 64'h11ffffff10000000;

	lut_sub lut_1262 ({sk[319], i_3_, i_2_, i_0_}, x241x);
	defparam lut_1262.LUT_SIZE = 4;
	defparam lut_1262.mask = 16'h7704;

	lut_sub lut_1264 ({sk[320], i_5_, i_6_, i_4_}, n_n87);
	defparam lut_1264.LUT_SIZE = 4;
	defparam lut_1264.mask = 16'h7704;

	lut_sub lut_1266 ({sk[321], i_8_, i_6_, n_n81, n_n85, x224x}, n_n554);
	defparam lut_1266.LUT_SIZE = 6;
	defparam lut_1266.mask = 64'h11ffffff55555755;

	lut_sub lut_1269 ({sk[322], i_7_, i_8_, i_6_, x26x, x45x}, x5055x);
	defparam lut_1269.LUT_SIZE = 6;
	defparam lut_1269.mask = 64'h11ffffff05000300;

	lut_sub lut_1272 ({sk[323], i_7_, i_8_, i_6_, n_n83, x34x, x354x}, x5056x);
	defparam lut_1272.LUT_SIZE = 7;
	defparam lut_1272.mask = 128'h03ff57ffffffffff0505000033000000;

	lut_sub lut_1275 ({sk[324], i_5_, i_3_, i_4_, n_n83, n_n82, x145x}, x297x);
	defparam lut_1275.LUT_SIZE = 7;
	defparam lut_1275.mask = 128'h03ff57ffffffffff5555555555555755;

	lut_sub lut_1278 ({sk[325], i_7_, i_8_, i_6_, n_n103, n_n102, x29x}, x147x);
	defparam lut_1278.LUT_SIZE = 7;
	defparam lut_1278.mask = 128'h03ff57ffffffffff0055030000000000;

	lut_sub lut_1281 ({sk[326], i_7_, i_8_, i_6_, n_n81, n_n103, n_n94}, x202x);
	defparam lut_1281.LUT_SIZE = 7;
	defparam lut_1281.mask = 128'h03ff57ffffffffff0000000503000000;

	lut_sub lut_1284 ({sk[327], i_7_, i_8_, i_6_, x63x, x347x, x23x}, x6371x);
	defparam lut_1284.LUT_SIZE = 7;
	defparam lut_1284.mask = 128'h03ff57fffffffffffff0ffffffaaff88;

	lut_sub lut_1293 ({sk[328], i_3_, i_1_, i_2_, i_0_, n_n93, x109x}, x97x);
	defparam lut_1293.LUT_SIZE = 7;
	defparam lut_1293.mask = 128'h03ff57ffffffffff0000100000100000;

	lut_sub lut_1296 ({sk[329], i_7_, i_8_, i_6_, x45x, x33x}, x146x);
	defparam lut_1296.LUT_SIZE = 6;
	defparam lut_1296.mask = 64'h11ffffff00070000;

	lut_sub lut_1299 ({sk[330], i_7_, i_8_, i_6_, x57x, x33x}, x270x);
	defparam lut_1299.LUT_SIZE = 6;
	defparam lut_1299.mask = 64'h11ffffff50300000;

	lut_sub lut_1302 ({sk[331], i_6_, i_3_, i_4_, n_n86, n_n100, n_n976}, x272x);
	defparam lut_1302.LUT_SIZE = 7;
	defparam lut_1302.mask = 128'h03ff57ffffffffff5755555555555555;

	lut_sub lut_1305 ({sk[332], i_7_, i_8_, i_6_, n_n81, n_n100, n_n77}, x151x);
	defparam lut_1305.LUT_SIZE = 7;
	defparam lut_1305.mask = 128'h03ff57ffffffffff0300000000000011;

	lut_sub lut_1308 ({sk[333], n_n84, n_n85, n_n95, x294x, n_n939, n_n978}, x6350x);
	defparam lut_1308.LUT_SIZE = 7;
	defparam lut_1308.mask = 128'h03ff57ffffffffff8080808080808000;

	lut_sub lut_1312 ({sk[334], i_6_, i_3_, i_2_, i_0_, n_n75, x109x}, n_n1093);
	defparam lut_1312.LUT_SIZE = 7;
	defparam lut_1312.mask = 128'h03ff57ffffffffff0010000000000000;

	lut_sub lut_1314 ({sk[335], i_7_, i_8_, i_6_, n_n94, n_n74}, n_n1052);
	defparam lut_1314.LUT_SIZE = 6;
	defparam lut_1314.mask = 64'h11ffffff00100000;

	lut_sub lut_1316 ({sk[336], i_5_, i_3_, i_4_, n_n101, n_n83, x37x}, x93x);
	defparam lut_1316.LUT_SIZE = 7;
	defparam lut_1316.mask = 128'h03ff57ffffffffff0055000300000000;

	lut_sub lut_1319 ({sk[337], i_5_, i_6_, i_4_}, n_n66);
	defparam lut_1319.LUT_SIZE = 4;
	defparam lut_1319.mask = 16'h7702;

	lut_sub lut_1321 ({sk[338], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x20x);
	defparam lut_1321.LUT_SIZE = 7;
	defparam lut_1321.mask = 128'h03ff57ffffffffff0004000000000000;

	lut_sub lut_1323 ({sk[339], i_3_, i_1_, i_2_}, x353x);
	defparam lut_1323.LUT_SIZE = 4;
	defparam lut_1323.mask = 16'h7740;

	lut_sub lut_1325 ({sk[340], i_7_, i_8_, n_n77, n_n66, x20x, x353x}, x117x);
	defparam lut_1325.LUT_SIZE = 7;
	defparam lut_1325.mask = 128'h03ff57ffffffffff0537003300330033;

	lut_sub lut_1328 ({sk[341], i_7_, i_8_, i_6_, n_n94, n_n74}, n_n1058);
	defparam lut_1328.LUT_SIZE = 6;
	defparam lut_1328.mask = 64'h11ffffff00000010;

	lut_sub lut_1330 ({sk[342], i_7_, i_6_, n_n103, n_n84, n_n1058}, x133x);
	defparam lut_1330.LUT_SIZE = 6;
	defparam lut_1330.mask = 64'h11ffffff55555755;

	lut_sub lut_1333 ({sk[343], i_5_, i_3_, i_4_, n_n94, n_n82}, x323x);
	defparam lut_1333.LUT_SIZE = 6;
	defparam lut_1333.mask = 64'h11ffffff10000000;

	lut_sub lut_1335 ({sk[344], i_7_, i_8_, i_6_, n_n103, n_n74, n_n85}, x201x);
	defparam lut_1335.LUT_SIZE = 7;
	defparam lut_1335.mask = 128'h03ff57ffffffffff0000000300110000;

	lut_sub lut_1338 ({sk[345], i_7_, i_8_, i_6_, n_n103, n_n77, n_n90}, x233x);
	defparam lut_1338.LUT_SIZE = 7;
	defparam lut_1338.mask = 128'h03ff57ffffffffff0000000300001300;

	lut_sub lut_1342 ({sk[346], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x347x);
	defparam lut_1342.LUT_SIZE = 7;
	defparam lut_1342.mask = 128'h03ff57ffffffffff4000000000000000;

	lut_sub lut_1344 ({sk[347], i_7_, i_8_, i_6_, n_n74, n_n90, x347x}, x197x);
	defparam lut_1344.LUT_SIZE = 7;
	defparam lut_1344.mask = 128'h03ff57ffffffffff5500550000030000;

	lut_sub lut_1347 ({sk[348], i_7_, i_8_, i_6_, x57x, x171x}, x5083x);
	defparam lut_1347.LUT_SIZE = 6;
	defparam lut_1347.mask = 64'h11ffffff30000505;

	lut_sub lut_1350 ({sk[349], i_7_, i_8_, i_6_, i_3_, i_4_}, x5085x);
	defparam lut_1350.LUT_SIZE = 6;
	defparam lut_1350.mask = 64'h11ffffff00000100;

	lut_sub lut_1352 ({sk[350], i_1_, i_2_, i_0_, x5085x}, n_n1020);
	defparam lut_1352.LUT_SIZE = 5;
	defparam lut_1352.mask = 32'h0f0f0040;

	lut_sub lut_1354 ({sk[351], i_1_, i_2_, i_0_, n_n74, n_n82, x5085x}, x271x);
	defparam lut_1354.LUT_SIZE = 7;
	defparam lut_1354.mask = 128'h03ff57ffffffffff0000000355000000;

	lut_sub lut_1357 ({sk[352], i_7_, i_8_, i_6_, n_n84, n_n85}, n_n949);
	defparam lut_1357.LUT_SIZE = 6;
	defparam lut_1357.mask = 64'h11ffffff00000100;

	lut_sub lut_1359 ({sk[353], i_7_, i_8_, i_6_, n_n84, n_n83, x144x}, x296x);
	defparam lut_1359.LUT_SIZE = 7;
	defparam lut_1359.mask = 128'h03ff57ffffffffff5555555557555555;

	lut_sub lut_1362 ({sk[354], i_7_, i_8_, i_6_, n_n83, n_n77, x29x}, x5115x);
	defparam lut_1362.LUT_SIZE = 7;
	defparam lut_1362.mask = 128'h03ff57ffffffffff0003000000550000;

	lut_sub lut_1365 ({sk[355], i_7_, i_8_, i_6_, x57x, x86x, x83x}, x306x);
	defparam lut_1365.LUT_SIZE = 7;
	defparam lut_1365.mask = 128'h03ff57ffffffffff330f550000000000;

	lut_sub lut_1369 ({sk[356], i_7_, i_8_, i_6_, n_n103, n_n96, x65x}, x5130x);
	defparam lut_1369.LUT_SIZE = 7;
	defparam lut_1369.mask = 128'h03ff57ffffffffff0355000000000000;

	lut_sub lut_1372 ({sk[357], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x67x);
	defparam lut_1372.LUT_SIZE = 7;
	defparam lut_1372.mask = 128'h03ff57ffffffffff0000080000000000;

	lut_sub lut_1374 ({sk[358], i_7_, i_8_, i_6_, n_n102, n_n90}, n_n1330);
	defparam lut_1374.LUT_SIZE = 6;
	defparam lut_1374.mask = 64'h11ffffff00000001;

	lut_sub lut_1376 ({sk[359], i_7_, i_8_, i_6_, n_n100, n_n84}, n_n1267);
	defparam lut_1376.LUT_SIZE = 6;
	defparam lut_1376.mask = 64'h11ffffff00000100;

	lut_sub lut_1378 ({sk[360], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x48x);
	defparam lut_1378.LUT_SIZE = 7;
	defparam lut_1378.mask = 128'h03ff57ffffffffff0000100000000000;

	lut_sub lut_1380 ({sk[361], i_7_, i_5_, i_3_, i_4_, i_0_}, x72x);
	defparam lut_1380.LUT_SIZE = 6;
	defparam lut_1380.mask = 64'h11ffffff80008080;

	lut_sub lut_1383 ({sk[362], i_3_, i_2_, i_0_, n_n93, x38x, x19x}, x123x);
	defparam lut_1383.LUT_SIZE = 7;
	defparam lut_1383.mask = 128'h03ff57ffffffffff0505053705050505;

	lut_sub lut_1386 ({sk[363], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x33x);
	defparam lut_1386.LUT_SIZE = 7;
	defparam lut_1386.mask = 128'h03ff57ffffffffff0000010000000000;

	lut_sub lut_1388 ({sk[364], i_7_, i_8_, i_6_, n_n85, n_n87, x33x}, x206x);
	defparam lut_1388.LUT_SIZE = 7;
	defparam lut_1388.mask = 128'h03ff57ffffffffff0000000000550303;

	lut_sub lut_1391 ({sk[365], i_5_, i_6_, i_3_}, n_n76);
	defparam lut_1391.LUT_SIZE = 4;
	defparam lut_1391.mask = 16'h7704;

	lut_sub lut_1393 ({sk[366], i_7_, i_8_, i_5_, i_6_, i_3_}, x244x);
	defparam lut_1393.LUT_SIZE = 6;
	defparam lut_1393.mask = 64'h11ffffff00000004;

	lut_sub lut_1395 ({sk[367], i_7_, i_8_, i_6_, n_n100, n_n96, x34x}, x273x);
	defparam lut_1395.LUT_SIZE = 7;
	defparam lut_1395.mask = 128'h03ff57ffffffffff0000000000550355;

	lut_sub lut_1398 ({sk[368], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x51x);
	defparam lut_1398.LUT_SIZE = 7;
	defparam lut_1398.mask = 128'h03ff57ffffffffff0000000000080000;

	lut_sub lut_1400 ({sk[369], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x52x);
	defparam lut_1400.LUT_SIZE = 7;
	defparam lut_1400.mask = 128'h03ff57ffffffffff0000000200000000;

	lut_sub lut_1402 ({sk[370], n_n101, x64x, x48x, n_n1088, n_n1181, x194x}, x6348x);
	defparam lut_1402.LUT_SIZE = 7;
	defparam lut_1402.mask = 128'h03ff57ffffffffffc080c080c0800000;

	lut_sub lut_1407 ({sk[371], i_7_, i_8_, i_6_, x42x, x86x, x52x}, x125x);
	defparam lut_1407.LUT_SIZE = 7;
	defparam lut_1407.mask = 128'h03ff57ffffffffff000000330055000f;

	lut_sub lut_1411 ({sk[372], i_5_, i_3_, i_4_, n_n93, n_n94}, n_n1042);
	defparam lut_1411.LUT_SIZE = 6;
	defparam lut_1411.mask = 64'h11ffffff00000010;

	lut_sub lut_1413 ({sk[373], n_n63, n_n85, x38x, x86x, x116x}, x6377x);
	defparam lut_1413.LUT_SIZE = 6;
	defparam lut_1413.mask = 64'h11ffffffaaa08880;

	lut_sub lut_1418 ({sk[374], i_5_, i_6_, i_4_}, n_n79);
	defparam lut_1418.LUT_SIZE = 4;
	defparam lut_1418.mask = 16'h7780;

	lut_sub lut_1420 ({sk[375], i_7_, i_8_, i_6_, n_n83, x34x, n_n79}, x185x);
	defparam lut_1420.LUT_SIZE = 7;
	defparam lut_1420.mask = 128'h03ff57ffffffffff0505003300000000;

	lut_sub lut_1423 ({sk[376], i_5_, i_6_, i_4_}, n_n40);
	defparam lut_1423.LUT_SIZE = 4;
	defparam lut_1423.mask = 16'h7740;

	lut_sub lut_1425 ({sk[377], i_7_, i_8_, i_6_, n_n94, n_n74}, n_n1074);
	defparam lut_1425.LUT_SIZE = 6;
	defparam lut_1425.mask = 64'h11ffffff00000100;

	lut_sub lut_1427 ({sk[378], i_6_, i_3_}, x28x);
	defparam lut_1427.LUT_SIZE = 3;
	defparam lut_1427.mask = 8'h58;

	lut_sub lut_1429 ({sk[379], i_5_, i_6_, i_3_, i_4_}, x5012x);
	defparam lut_1429.LUT_SIZE = 5;
	defparam lut_1429.mask = 32'h0f0f0800;

	lut_sub lut_1431 ({sk[380], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x86x);
	defparam lut_1431.LUT_SIZE = 7;
	defparam lut_1431.mask = 128'h03ff57ffffffffff0000000000000800;

	lut_sub lut_1433 ({sk[381], i_7_, i_8_, i_6_, n_n81, n_n90}, n_n1057);
	defparam lut_1433.LUT_SIZE = 6;
	defparam lut_1433.mask = 64'h11ffffff00001000;

	lut_sub lut_1435 ({sk[382], i_7_, i_8_, i_6_, n_n81, n_n90}, n_n1125);
	defparam lut_1435.LUT_SIZE = 6;
	defparam lut_1435.mask = 64'h11ffffff10000000;

	lut_sub lut_1437 ({sk[383], i_7_, i_8_, i_6_, n_n84, n_n94}, n_n1128);
	defparam lut_1437.LUT_SIZE = 6;
	defparam lut_1437.mask = 64'h11ffffff10000000;

	lut_sub lut_1439 ({sk[384], i_5_, i_3_, i_4_, n_n94, n_n82, n_n1330}, x136x);
	defparam lut_1439.LUT_SIZE = 7;
	defparam lut_1439.mask = 128'h03ff57ffffffffff5555555555555755;

	lut_sub lut_1442 ({sk[385], i_7_, i_5_, i_6_, i_3_, i_4_, n_n94}, x333x);
	defparam lut_1442.LUT_SIZE = 7;
	defparam lut_1442.mask = 128'h03ff57ffffffffff0000000000000004;

	lut_sub lut_1444 ({sk[386], i_7_, i_8_, i_6_, n_n74, n_n90, x86x}, x278x);
	defparam lut_1444.LUT_SIZE = 7;
	defparam lut_1444.mask = 128'h03ff57ffffffffff0000000003005700;

	lut_sub lut_1447 ({sk[387], i_1_, i_2_, i_0_}, n_n937);
	defparam lut_1447.LUT_SIZE = 4;
	defparam lut_1447.mask = 16'h7780;

	lut_sub lut_1449 ({sk[388], i_5_, i_6_, i_3_, i_4_, i_1_, i_0_}, x1315x);
	defparam lut_1449.LUT_SIZE = 7;
	defparam lut_1449.mask = 128'h03ff57ffffffffff8000000000000000;

	lut_sub lut_1451 ({sk[389], i_7_, i_8_, i_6_, n_n81, n_n94}, n_n1087);
	defparam lut_1451.LUT_SIZE = 6;
	defparam lut_1451.mask = 64'h11ffffff00100000;

	lut_sub lut_1453 ({sk[390], x241x, x93x, x318x, n_n1294, x290x, x217x}, n_n663);
	defparam lut_1453.LUT_SIZE = 7;
	defparam lut_1453.mask = 128'h03ff57ffffffffff7f7fffff7fffffff;

	lut_sub lut_1459 ({sk[391], x27x, n_n95, x323x, x191x, x71x, x118x}, x5308x);
	defparam lut_1459.LUT_SIZE = 7;
	defparam lut_1459.mask = 128'h03ff57ffffffffff7fff7fff7fffffff;

	lut_sub lut_1465 ({sk[392], n_n101, x74x, x174x, x339x, x5283x, x6346x}, x5309x);
	defparam lut_1465.LUT_SIZE = 7;
	defparam lut_1465.mask = 128'h03ff57ffffffffffbbbfbbbfbbbfffff;

	lut_sub lut_1470 ({sk[393], n_n95, x43x, x333x, x5288x, x5289x, x5290x}, x5310x);
	defparam lut_1470.LUT_SIZE = 7;
	defparam lut_1470.mask = 128'h03ff57ffffffffff7fff7fff7fffffff;

	lut_sub lut_1476 ({sk[394], x5291x, x5292x, x5293x, x5294x}, x5311x);
	defparam lut_1476.LUT_SIZE = 5;
	defparam lut_1476.mask = 32'h0f0f7fff;

	lut_sub lut_1481 ({sk[395], x207x, x61x, x308x, x5295x, x5296x}, x5312x);
	defparam lut_1481.LUT_SIZE = 6;
	defparam lut_1481.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1487 ({sk[396], i_7_, i_8_, i_6_, n_n85, n_n77}, n_n958);
	defparam lut_1487.LUT_SIZE = 6;
	defparam lut_1487.mask = 64'h11ffffff00000001;

	lut_sub lut_1489 ({sk[397], i_7_, i_8_, i_5_, i_6_, i_4_, n_n83}, n_n974);
	defparam lut_1489.LUT_SIZE = 7;
	defparam lut_1489.mask = 128'h03ff57ffffffffff0000000000040000;

	lut_sub lut_1491 ({sk[398], i_7_, i_8_, i_6_, n_n81, n_n94}, n_n989);
	defparam lut_1491.LUT_SIZE = 6;
	defparam lut_1491.mask = 64'h11ffffff00010000;

	lut_sub lut_1493 ({sk[399], i_7_, i_8_, i_6_, x29x}, n_n944);
	defparam lut_1493.LUT_SIZE = 5;
	defparam lut_1493.mask = 32'h0f0f0100;

	lut_sub lut_1495 ({sk[400], i_5_, i_3_, i_4_, n_n93, n_n83}, n_n982);
	defparam lut_1495.LUT_SIZE = 6;
	defparam lut_1495.mask = 64'h3333ffff00000001;

	lut_sub lut_1497 ({sk[401], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x24x);
	defparam lut_1497.LUT_SIZE = 7;
	defparam lut_1497.mask = 128'h0707ffff1717ffff0000000000400000;

	lut_sub lut_1499 ({sk[402], i_7_, i_8_, n_n103, x4871x, x59x}, x286x);
	defparam lut_1499.LUT_SIZE = 6;
	defparam lut_1499.mask = 64'h3333ffff55555557;

	lut_sub lut_1502 ({sk[403], x57x, n_n63, n_n95, x73x, x24x, x171x}, x5331x);
	defparam lut_1502.LUT_SIZE = 7;
	defparam lut_1502.mask = 128'h0707ffff1717ffff00335f7f0033ffff;

	lut_sub lut_1507 ({sk[404], i_7_, i_8_, i_5_, i_6_, i_4_, n_n90}, n_n1121);
	defparam lut_1507.LUT_SIZE = 7;
	defparam lut_1507.mask = 128'h0707ffff1717ffff0000000000010000;

	lut_sub lut_1509 ({sk[405], i_3_, i_1_, i_2_}, n_n53);
	defparam lut_1509.LUT_SIZE = 4;
	defparam lut_1509.mask = 16'h1f10;

	lut_sub lut_1511 ({sk[406], i_1_, i_2_}, x330x);
	defparam lut_1511.LUT_SIZE = 3;
	defparam lut_1511.mask = 8'h32;

	lut_sub lut_1513 ({sk[407], i_5_, i_3_, n_n80, n_n73, n_n40, x330x}, x70x);
	defparam lut_1513.LUT_SIZE = 7;
	defparam lut_1513.mask = 128'h0707ffff1717ffff0537003300330033;

	lut_sub lut_1516 ({sk[408], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x83x);
	defparam lut_1516.LUT_SIZE = 7;
	defparam lut_1516.mask = 128'h0707ffff1717ffff0000000000000100;

	lut_sub lut_1518 ({sk[409], i_7_, i_8_, i_6_, n_n94, n_n96, x73x}, x90x);
	defparam lut_1518.LUT_SIZE = 7;
	defparam lut_1518.mask = 128'h0707ffff1717ffff5700000003000000;

	lut_sub lut_1521 ({sk[410], i_7_, i_8_, i_6_, n_n83, n_n74, x128x}, x115x);
	defparam lut_1521.LUT_SIZE = 7;
	defparam lut_1521.mask = 128'h0707ffff1717ffff0300000000000055;

	lut_sub lut_1524 ({sk[411], i_7_, i_8_, i_6_, n_n100, n_n102, x115x}, x168x);
	defparam lut_1524.LUT_SIZE = 7;
	defparam lut_1524.mask = 128'h0707ffff1717ffff5555555555555557;

	lut_sub lut_1527 ({sk[412], i_7_, i_8_, i_5_, i_6_, i_4_, n_n67}, n_n977);
	defparam lut_1527.LUT_SIZE = 7;
	defparam lut_1527.mask = 128'h0707ffff1717ffff0000000000004000;

	lut_sub lut_1529 ({sk[413], i_5_, i_6_, i_4_}, x5338x);
	defparam lut_1529.LUT_SIZE = 4;
	defparam lut_1529.mask = 16'h1f01;

	lut_sub lut_1531 ({sk[414], i_7_, i_8_, n_n85, n_n79, x5338x, n_n67}, x215x);
	defparam lut_1531.LUT_SIZE = 7;
	defparam lut_1531.mask = 128'h0707ffff1717ffff0000003300000505;

	lut_sub lut_1534 ({sk[415], i_7_, i_8_, i_1_, i_2_, i_0_, n_n87}, x236x);
	defparam lut_1534.LUT_SIZE = 7;
	defparam lut_1534.mask = 128'h0707ffff1717ffff0000000000001000;

	lut_sub lut_1536 ({sk[416], i_7_, i_8_, i_6_, i_3_, i_4_, n_n90}, n_n1118);
	defparam lut_1536.LUT_SIZE = 7;
	defparam lut_1536.mask = 128'h0707ffff1717ffff0000001000000000;

	lut_sub lut_1538 ({sk[417], i_7_, i_8_, n_n84, n_n94, x127x, n_n90}, x262x);
	defparam lut_1538.LUT_SIZE = 7;
	defparam lut_1538.mask = 128'h0707ffff1717ffff00001111000f0000;

	lut_sub lut_1541 ({sk[418], i_7_, i_5_, i_6_, i_3_, i_4_, n_n103}, n_n993);
	defparam lut_1541.LUT_SIZE = 7;
	defparam lut_1541.mask = 128'h0707ffff1717ffff0000000100000000;

	lut_sub lut_1543 ({sk[419], i_7_, i_8_, i_6_, n_n83, n_n74, n_n993}, x275x);
	defparam lut_1543.LUT_SIZE = 7;
	defparam lut_1543.mask = 128'h0707ffff1717ffff5555555555555557;

	lut_sub lut_1546 ({sk[420], i_7_, i_8_, i_6_, n_n81, n_n94, n_n85}, x145x);
	defparam lut_1546.LUT_SIZE = 7;
	defparam lut_1546.mask = 128'h0707ffff1717ffff0300000005000000;

	lut_sub lut_1549 ({sk[421], i_7_, i_5_, i_6_, i_3_, i_4_, n_n90}, x319x);
	defparam lut_1549.LUT_SIZE = 7;
	defparam lut_1549.mask = 128'h0707ffff1717ffff0000100000000000;

	lut_sub lut_1551 ({sk[422], i_3_, n_n38, n_n64, n_n83, n_n74, n_n85}, x5379x);
	defparam lut_1551.LUT_SIZE = 7;
	defparam lut_1551.mask = 128'h0707ffff1717ffff001100110011001f;

	lut_sub lut_1554 ({sk[423], n_n80, x234x, x116x, n_n882, x296x, x5379x}, x5388x);
	defparam lut_1554.LUT_SIZE = 7;
	defparam lut_1554.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_1560 ({sk[424], i_1_, i_2_, i_0_, n_n102, n_n95, n_n949}, n_n652);
	defparam lut_1560.LUT_SIZE = 7;
	defparam lut_1560.mask = 128'h0707ffff1717ffff5555555555555757;

	lut_sub lut_1564 ({sk[425], i_7_, i_8_, i_6_, x42x, n_n90, x5012x}, x195x);
	defparam lut_1564.LUT_SIZE = 7;
	defparam lut_1564.mask = 128'h0707ffff1717ffff1f11111111111111;

	lut_sub lut_1567 ({sk[426], i_8_, i_5_, i_6_, i_3_, i_4_, n_n94}, n_n1045);
	defparam lut_1567.LUT_SIZE = 7;
	defparam lut_1567.mask = 128'h0707ffff1717ffff0000000004000000;

	lut_sub lut_1569 ({sk[427], i_7_, i_8_, i_6_, n_n102, n_n85}, n_n1043);
	defparam lut_1569.LUT_SIZE = 6;
	defparam lut_1569.mask = 64'h3333ffff00010000;

	lut_sub lut_1571 ({sk[428], i_5_, i_3_, i_4_, n_n93, n_n85, x95x}, x289x);
	defparam lut_1571.LUT_SIZE = 7;
	defparam lut_1571.mask = 128'h0707ffff1717ffff5555555555555557;

	lut_sub lut_1574 ({sk[429], i_7_, i_8_, i_6_, n_n100, n_n84, x96x}, x290x);
	defparam lut_1574.LUT_SIZE = 7;
	defparam lut_1574.mask = 128'h0707ffff1717ffff5555555557555555;

	lut_sub lut_1577 ({sk[430], i_7_, i_8_, i_6_, n_n96, n_n90, x74x}, x5406x);
	defparam lut_1577.LUT_SIZE = 7;
	defparam lut_1577.mask = 128'h0707ffff1717ffff0355000000000000;

	lut_sub lut_1580 ({sk[431], i_7_, i_8_, i_6_, n_n102, n_n77, n_n90}, x5407x);
	defparam lut_1580.LUT_SIZE = 7;
	defparam lut_1580.mask = 128'h0707ffff1717ffff0011050000000000;

	lut_sub lut_1583 ({sk[432], i_5_, i_3_, i_4_, n_n93, x32x, n_n94}, x5412x);
	defparam lut_1583.LUT_SIZE = 7;
	defparam lut_1583.mask = 128'h0707ffff1717ffff0000000000053300;

	lut_sub lut_1586 ({sk[433], x289x, x290x, x5406x, x5407x, x5412x}, x5421x);
	defparam lut_1586.LUT_SIZE = 6;
	defparam lut_1586.mask = 64'h3333ffff7fffffff;

	lut_sub lut_1592 ({sk[434], i_7_, i_8_, i_6_, x128x}, n_n1122);
	defparam lut_1592.LUT_SIZE = 5;
	defparam lut_1592.mask = 32'h0fff0010;

	lut_sub lut_1594 ({sk[435], i_5_, i_6_, i_3_, n_n91, x67x, x62x}, x158x);
	defparam lut_1594.LUT_SIZE = 7;
	defparam lut_1594.mask = 128'h0707ffff1717ffff0303030357030303;

	lut_sub lut_1597 ({sk[436], i_5_, i_3_, i_4_, x75x, x48x, x315x}, x5429x);
	defparam lut_1597.LUT_SIZE = 7;
	defparam lut_1597.mask = 128'h0707ffff1717ffff0505330005370000;

	lut_sub lut_1601 ({sk[437], i_7_, i_8_, i_6_, x23x, x33x}, x5430x);
	defparam lut_1601.LUT_SIZE = 6;
	defparam lut_1601.mask = 64'h3333ffff30000050;

	lut_sub lut_1604 ({sk[438], n_n101, x22x, x158x, x304x, x5429x, x5430x}, x5440x);
	defparam lut_1604.LUT_SIZE = 7;
	defparam lut_1604.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_1610 ({sk[439], i_7_, i_8_, i_1_, i_2_, i_0_}, x66x);
	defparam lut_1610.LUT_SIZE = 6;
	defparam lut_1610.mask = 64'h3333ffff00000002;

	lut_sub lut_1612 ({sk[440], i_6_, i_3_, i_4_}, x5442x);
	defparam lut_1612.LUT_SIZE = 4;
	defparam lut_1612.mask = 16'h1f02;

	lut_sub lut_1614 ({sk[441], i_6_, i_3_, i_2_, i_0_, n_n70, x109x}, n_n1101);
	defparam lut_1614.LUT_SIZE = 7;
	defparam lut_1614.mask = 128'h0707ffff1717ffff0010000000000000;

	lut_sub lut_1616 ({sk[442], i_7_, i_8_, i_6_, n_n84, n_n94, x23x}, x196x);
	defparam lut_1616.LUT_SIZE = 7;
	defparam lut_1616.mask = 128'h0707ffff1717ffff0003000055000000;

	lut_sub lut_1619 ({sk[443], i_7_, i_8_, i_5_, i_6_, x19x, n_n90}, x5446x);
	defparam lut_1619.LUT_SIZE = 7;
	defparam lut_1619.mask = 128'h0707ffff1717ffff0000353000000000;

	lut_sub lut_1622 ({sk[444], i_5_, n_n101, n_n91, x128x, x353x, x101x}, x6360x);
	defparam lut_1622.LUT_SIZE = 7;
	defparam lut_1622.mask = 128'h0707ffff1717ffffaaa08880aaa0aaa0;

	lut_sub lut_1629 ({sk[445], n_n86, n_n73, x67x, x196x, x5446x, x6360x}, n_n593);
	defparam lut_1629.LUT_SIZE = 7;
	defparam lut_1629.mask = 128'h0707ffff1717ffffbfbfbfbfbfbfbfff;

	lut_sub lut_1634 ({sk[446], i_7_, i_8_, i_3_, i_2_, i_0_, n_n71}, n_n1059);
	defparam lut_1634.LUT_SIZE = 7;
	defparam lut_1634.mask = 128'h0707ffff1717ffff0001000000000000;

	lut_sub lut_1636 ({sk[447], i_7_, i_8_, i_6_, n_n94, n_n74, n_n96}, x263x);
	defparam lut_1636.LUT_SIZE = 7;
	defparam lut_1636.mask = 128'h0707ffff1717ffff0000030000000500;

	lut_sub lut_1639 ({sk[448], i_7_, i_8_, i_6_, x73x, x325x, n_n53}, x91x);
	defparam lut_1639.LUT_SIZE = 7;
	defparam lut_1639.mask = 128'h0707ffff1717ffff000000000f001100;

	lut_sub lut_1642 ({sk[449], i_8_, i_3_, i_1_, i_0_, n_n40, n_n1060}, x156x);
	defparam lut_1642.LUT_SIZE = 7;
	defparam lut_1642.mask = 128'h0707ffff1717ffff5555555555555755;

	lut_sub lut_1645 ({sk[450], x133x, n_n1059, x263x, x91x, x156x}, n_n597);
	defparam lut_1645.LUT_SIZE = 6;
	defparam lut_1645.mask = 64'h3333ffff7fffffff;

	lut_sub lut_1651 ({sk[451], i_7_, i_6_, n_n102, n_n94, n_n1070}, x141x);
	defparam lut_1651.LUT_SIZE = 6;
	defparam lut_1651.mask = 64'h3333ffff55555557;

	lut_sub lut_1654 ({sk[452], i_7_, i_8_, i_6_, x76x, n_n79, n_n53}, x142x);
	defparam lut_1654.LUT_SIZE = 7;
	defparam lut_1654.mask = 128'h0707ffff1717ffff0f00000011110000;

	lut_sub lut_1657 ({sk[453], i_7_, i_8_, i_6_, n_n81, n_n94, x42x}, x150x);
	defparam lut_1657.LUT_SIZE = 7;
	defparam lut_1657.mask = 128'h0707ffff1717ffff0000550000000300;

	lut_sub lut_1660 ({sk[454], i_7_, i_8_, i_6_, n_n102, n_n90}, n_n1046);
	defparam lut_1660.LUT_SIZE = 6;
	defparam lut_1660.mask = 64'h3333ffff00000100;

	lut_sub lut_1662 ({sk[455], i_7_, i_8_, i_6_, n_n81, n_n90}, n_n1047);
	defparam lut_1662.LUT_SIZE = 6;
	defparam lut_1662.mask = 64'h3333ffff00100000;

	lut_sub lut_1664 ({sk[456], i_7_, i_8_, i_6_, x26x, n_n83, n_n102}, x279x);
	defparam lut_1664.LUT_SIZE = 7;
	defparam lut_1664.mask = 128'h0707ffff1717ffff0000000f00000011;

	lut_sub lut_1667 ({sk[457], i_5_, i_3_, i_4_, n_n94, n_n95}, n_n1048);
	defparam lut_1667.LUT_SIZE = 6;
	defparam lut_1667.mask = 64'h3333ffff00001000;

	lut_sub lut_1669 ({sk[458], i_5_, i_6_, i_4_}, n_n71);
	defparam lut_1669.LUT_SIZE = 4;
	defparam lut_1669.mask = 16'h1f20;

	lut_sub lut_1671 ({sk[459], i_7_, i_8_, i_3_, i_1_, i_0_}, x85x);
	defparam lut_1671.LUT_SIZE = 6;
	defparam lut_1671.mask = 64'h3333ffff00400000;

	lut_sub lut_1673 ({sk[460], i_3_, n_n94, n_n95, x109x, n_n71, x85x}, x282x);
	defparam lut_1673.LUT_SIZE = 7;
	defparam lut_1673.mask = 128'h0707ffff1717ffff1111111f11111111;

	lut_sub lut_1676 ({sk[461], i_7_, i_8_, i_6_, n_n100, n_n94, n_n74}, x285x);
	defparam lut_1676.LUT_SIZE = 7;
	defparam lut_1676.mask = 128'h0707ffff1717ffff0000000500110000;

	lut_sub lut_1679 ({sk[462], i_7_, i_8_, i_6_, n_n103, n_n74}, n_n1060);
	defparam lut_1679.LUT_SIZE = 6;
	defparam lut_1679.mask = 64'h3333ffff00100000;

	lut_sub lut_1681 ({sk[463], i_7_, i_8_, i_6_, n_n83, n_n77}, n_n969);
	defparam lut_1681.LUT_SIZE = 6;
	defparam lut_1681.mask = 64'h3333ffff01000000;

	lut_sub lut_1683 ({sk[464], i_8_, i_6_}, x331x);
	defparam lut_1683.LUT_SIZE = 3;
	defparam lut_1683.mask = 8'h38;

	lut_sub lut_1685 ({sk[465], i_8_, i_5_, i_6_, i_3_, i_4_, n_n100}, n_n939);
	defparam lut_1685.LUT_SIZE = 7;
	defparam lut_1685.mask = 128'h0707ffff1717ffff4000000000000000;

	lut_sub lut_1687 ({sk[466], i_6_, i_3_, i_4_}, x131x);
	defparam lut_1687.LUT_SIZE = 4;
	defparam lut_1687.mask = 16'h1f80;

	lut_sub lut_1689 ({sk[467], i_7_, i_8_, i_1_, i_2_, i_0_}, x5068x);
	defparam lut_1689.LUT_SIZE = 6;
	defparam lut_1689.mask = 64'h3333ffff40000000;

	lut_sub lut_1691 ({sk[468], i_7_, i_8_, i_6_, i_3_, i_4_, n_n100}, n_n971);
	defparam lut_1691.LUT_SIZE = 7;
	defparam lut_1691.mask = 128'h0707ffff1717ffff4000000000000000;

	lut_sub lut_1693 ({sk[469], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x107x);
	defparam lut_1693.LUT_SIZE = 7;
	defparam lut_1693.mask = 128'h0707ffff1717ffff0000000000040000;

	lut_sub lut_1695 ({sk[470], n_n78, x76x, n_n95, x21x, n_n40, x66x}, n_n421);
	defparam lut_1695.LUT_SIZE = 7;
	defparam lut_1695.mask = 128'h0707ffff1717ffff111f111f111fffff;

	lut_sub lut_1699 ({sk[471], i_3_, i_2_, i_0_, x329x, x38x}, x159x);
	defparam lut_1699.LUT_SIZE = 6;
	defparam lut_1699.mask = 64'h3333ffff33733333;

	lut_sub lut_1702 ({sk[472], n_n81, n_n101, n_n91, n_n83, x45x, x239x}, x300x);
	defparam lut_1702.LUT_SIZE = 7;
	defparam lut_1702.mask = 128'h0707ffff1717ffff00553377005f337f;

	lut_sub lut_1706 ({sk[473], x267x, x100x, x119x, x160x}, x5533x);
	defparam lut_1706.LUT_SIZE = 5;
	defparam lut_1706.mask = 32'h0fff7fff;

	lut_sub lut_1711 ({sk[474], n_n81, n_n84, x48x, x5519x, x5520x, x5522x}, x5536x);
	defparam lut_1711.LUT_SIZE = 7;
	defparam lut_1711.mask = 128'h0707ffff1717ffff7f7f7fff7fff7fff;

	lut_sub lut_1717 ({sk[475], n_n58, x262x, x44x, n_n1145, x265x, x6340x}, x5512x);
	defparam lut_1717.LUT_SIZE = 7;
	defparam lut_1717.mask = 128'h0707ffff1717ffffbfbfffffbfffffff;

	lut_sub lut_1723 ({sk[476], n_n91, x44x, x224x, n_n1108, x92x, x269x}, x5510x);
	defparam lut_1723.LUT_SIZE = 7;
	defparam lut_1723.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_1729 ({sk[477], n_n58, x64x, n_n1132, x101x, x102x, x5499x}, x5511x);
	defparam lut_1729.LUT_SIZE = 7;
	defparam lut_1729.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_1735 ({sk[478], n_n78, n_n1172, x216x, x23x, x166x, x220x}, x5534x);
	defparam lut_1735.LUT_SIZE = 7;
	defparam lut_1735.mask = 128'h0707ffff1717ffff77ffffff7fffffff;

	lut_sub lut_1741 ({sk[479], n_n78, n_n1259, x53x, n_n1176, n_n1184, x5529x}, x5535x);
	defparam lut_1741.LUT_SIZE = 7;
	defparam lut_1741.mask = 128'h0707ffff1717ffff7f7fffff7fffffff;

	lut_sub lut_1747 ({sk[480], i_7_, i_8_, i_3_, i_1_, i_0_, n_n87}, n_n947);
	defparam lut_1747.LUT_SIZE = 7;
	defparam lut_1747.mask = 128'h0707ffff1717ffff0400000000000000;

	lut_sub lut_1749 ({sk[481], i_7_, i_8_, i_6_, x29x, n_n947}, x162x);
	defparam lut_1749.LUT_SIZE = 6;
	defparam lut_1749.mask = 64'h3333ffff55555557;

	lut_sub lut_1752 ({sk[482], i_3_, i_4_}, x312x);
	defparam lut_1752.LUT_SIZE = 3;
	defparam lut_1752.mask = 8'h32;

	lut_sub lut_1754 ({sk[483], i_1_, i_2_, i_0_, x77x, x162x, x312x}, n_n241);
	defparam lut_1754.LUT_SIZE = 7;
	defparam lut_1754.mask = 128'h0707ffff1717ffff3333333333333337;

	lut_sub lut_1757 ({sk[484], i_7_, i_8_, n_n85, n_n76, n_n1026}, x5547x);
	defparam lut_1757.LUT_SIZE = 6;
	defparam lut_1757.mask = 64'h3333ffff57555555;

	lut_sub lut_1760 ({sk[485], n_n882, x147x, x202x, x286x, x5547x}, x5556x);
	defparam lut_1760.LUT_SIZE = 6;
	defparam lut_1760.mask = 64'h3333ffff7fffffff;

	lut_sub lut_1766 ({sk[486], i_1_, i_2_, i_0_, n_n70, x38x, n_n87}, x68x);
	defparam lut_1766.LUT_SIZE = 7;
	defparam lut_1766.mask = 128'h0707ffff1717ffff0000000000330005;

	lut_sub lut_1769 ({sk[487], i_3_, i_4_, n_n91, x108x, n_n87, x85x}, x138x);
	defparam lut_1769.LUT_SIZE = 7;
	defparam lut_1769.mask = 128'h0707ffff1717ffff1111111f11111111;

	lut_sub lut_1772 ({sk[488], n_n80, n_n86, n_n85, n_n95, n_n77, n_n79}, x153x);
	defparam lut_1772.LUT_SIZE = 7;
	defparam lut_1772.mask = 128'h0707ffff1717ffff0003000300035557;

	lut_sub lut_1775 ({sk[489], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x317x);
	defparam lut_1775.LUT_SIZE = 7;
	defparam lut_1775.mask = 128'h0707ffff1717ffff0000000010000000;

	lut_sub lut_1777 ({sk[490], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x4901x);
	defparam lut_1777.LUT_SIZE = 7;
	defparam lut_1777.mask = 128'h0707ffff1717ffff0000000000100000;

	lut_sub lut_1779 ({sk[491], i_7_, i_8_, i_6_, n_n84, n_n94}, n_n1184);
	defparam lut_1779.LUT_SIZE = 6;
	defparam lut_1779.mask = 64'h3333ffff00000001;

	lut_sub lut_1781 ({sk[492], i_7_, i_8_, i_6_, i_3_, i_4_, n_n94}, n_n1145);
	defparam lut_1781.LUT_SIZE = 7;
	defparam lut_1781.mask = 128'h0707ffff1717ffff0000000001000000;

	lut_sub lut_1783 ({sk[493], i_1_, i_0_}, x175x);
	defparam lut_1783.LUT_SIZE = 3;
	defparam lut_1783.mask = 8'h32;

	lut_sub lut_1785 ({sk[494], i_5_, i_3_, i_4_, n_n93, n_n94, n_n85}, x224x);
	defparam lut_1785.LUT_SIZE = 7;
	defparam lut_1785.mask = 128'h0707ffff1717ffff0000030500000000;

	lut_sub lut_1788 ({sk[495], i_7_, i_8_, i_1_, i_2_, i_0_, x130x}, x5595x);
	defparam lut_1788.LUT_SIZE = 7;
	defparam lut_1788.mask = 128'h0707ffff1717ffff0004004000000000;

	lut_sub lut_1791 ({sk[496], n_n100, n_n102, n_n70, n_n63, n_n71, x242x}, x5596x);
	defparam lut_1791.LUT_SIZE = 7;
	defparam lut_1791.mask = 128'h0707ffff1717ffff0011001100110f1f;

	lut_sub lut_1794 ({sk[497], i_5_, i_3_, i_4_, n_n91, n_n100, x20x}, x95x);
	defparam lut_1794.LUT_SIZE = 7;
	defparam lut_1794.mask = 128'h0707ffff1717ffff5500000300000000;

	lut_sub lut_1797 ({sk[498], i_7_, i_8_, i_6_, n_n81, n_n83, x43x}, x217x);
	defparam lut_1797.LUT_SIZE = 7;
	defparam lut_1797.mask = 128'h0707ffff1717ffff0000570000005500;

	lut_sub lut_1800 ({sk[499], i_5_, i_3_, i_4_, n_n100, x331x, x316x}, x122x);
	defparam lut_1800.LUT_SIZE = 7;
	defparam lut_1800.mask = 128'h0707ffff1717ffff5500000000000300;

	lut_sub lut_1803 ({sk[500], i_7_, i_8_, i_6_, x45x, x21x, x24x}, x5597x);
	defparam lut_1803.LUT_SIZE = 7;
	defparam lut_1803.mask = 128'h0707ffff1717ffff333300550000000f;

	lut_sub lut_1807 ({sk[501], n_n93, n_n78, x26x, x43x, x49x, x24x}, x5600x);
	defparam lut_1807.LUT_SIZE = 7;
	defparam lut_1807.mask = 128'h0707ffff1717ffff00007f7f00ff7fff;

	lut_sub lut_1812 ({sk[502], x148x, x114x, x296x, x167x, x5613x}, x5622x);
	defparam lut_1812.LUT_SIZE = 6;
	defparam lut_1812.mask = 64'h3333ffff7fffffff;

	lut_sub lut_1818 ({sk[503], n_n86, n_n73, x29x, x201x, x271x, x275x}, x5620x);
	defparam lut_1818.LUT_SIZE = 7;
	defparam lut_1818.mask = 128'h0707ffff1717ffff7f7f7f7f7f7f7fff;

	lut_sub lut_1823 ({sk[504], x57x, n_n63, n_n982, x152x, x5617x}, x5621x);
	defparam lut_1823.LUT_SIZE = 6;
	defparam lut_1823.mask = 64'h3333ffff7f7f7fff;

	lut_sub lut_1828 ({sk[505], n_n91, x45x, x97x, x125x, x33x, x5633x}, x5652x);
	defparam lut_1828.LUT_SIZE = 7;
	defparam lut_1828.mask = 128'h0707ffff1717ffff5fff5fff7fffffff;

	lut_sub lut_1834 ({sk[506], x279x, x153x, x204x, x287x, x6368x}, x5653x);
	defparam lut_1834.LUT_SIZE = 6;
	defparam lut_1834.mask = 64'h3333ffffbfffffff;

	lut_sub lut_1840 ({sk[507], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x65x);
	defparam lut_1840.LUT_SIZE = 7;
	defparam lut_1840.mask = 128'h0707ffff1717ffff0000000000000040;

	lut_sub lut_1842 ({sk[508], i_7_, i_8_, i_6_, n_n102, n_n90, x65x}, x216x);
	defparam lut_1842.LUT_SIZE = 7;
	defparam lut_1842.mask = 128'h0707ffff1717ffff0000000003000055;

	lut_sub lut_1845 ({sk[509], i_7_, i_8_, i_6_, x128x, x216x}, n_n211);
	defparam lut_1845.LUT_SIZE = 6;
	defparam lut_1845.mask = 64'h3333ffff55555575;

	lut_sub lut_1848 ({sk[510], i_4_, n_n70, n_n63, n_n85, x83x, x28x}, x120x);
	defparam lut_1848.LUT_SIZE = 7;
	defparam lut_1848.mask = 128'h0707ffff1717ffff0033003300330537;

	lut_sub lut_1851 ({sk[511], i_7_, i_8_, i_6_, n_n81, n_n83}, n_n1160);
	defparam lut_1851.LUT_SIZE = 6;
	defparam lut_1851.mask = 64'h3333ffff00000100;

	lut_sub lut_1853 ({sk[512], i_7_, i_8_, i_6_, n_n100, n_n84, x55x}, x191x);
	defparam lut_1853.LUT_SIZE = 7;
	defparam lut_1853.mask = 128'h0707ffff1717ffff0000000000550300;

	lut_sub lut_1856 ({sk[513], i_7_, i_8_, i_6_, n_n100, n_n74, x52x}, x264x);
	defparam lut_1856.LUT_SIZE = 7;
	defparam lut_1856.mask = 128'h0707ffff1717ffff5500000000030000;

	lut_sub lut_1859 ({sk[514], i_5_, i_3_, i_4_, n_n101, n_n85}, n_n1146);
	defparam lut_1859.LUT_SIZE = 6;
	defparam lut_1859.mask = 64'h3333ffff00001000;

	lut_sub lut_1861 ({sk[515], i_5_, i_3_, i_4_, n_n78, n_n103, x107x}, x265x);
	defparam lut_1861.LUT_SIZE = 7;
	defparam lut_1861.mask = 128'h0707ffff1717ffff0000000057000000;

	lut_sub lut_1864 ({sk[516], i_7_, i_8_, i_6_, n_n84, n_n83}, n_n980);
	defparam lut_1864.LUT_SIZE = 6;
	defparam lut_1864.mask = 64'h3333ffff00001000;

	lut_sub lut_1866 ({sk[517], i_7_, i_8_, i_6_, n_n84, n_n85}, n_n1130);
	defparam lut_1866.LUT_SIZE = 6;
	defparam lut_1866.mask = 64'h3333ffff00000010;

	lut_sub lut_1868 ({sk[518], i_3_, i_4_, i_1_, i_0_, n_n93, n_n1160}, x5716x);
	defparam lut_1868.LUT_SIZE = 7;
	defparam lut_1868.mask = 128'h0707ffff1717ffff5555555557555555;

	lut_sub lut_1871 ({sk[519], i_7_, i_8_, i_6_, n_n74, n_n85, x325x}, x5717x);
	defparam lut_1871.LUT_SIZE = 7;
	defparam lut_1871.mask = 128'h0707ffff1717ffff0000030011000000;

	lut_sub lut_1874 ({sk[520], i_5_, i_3_, i_4_, n_n93, n_n100, x37x}, x5718x);
	defparam lut_1874.LUT_SIZE = 7;
	defparam lut_1874.mask = 128'h0707ffff1717ffff0003000000000055;

	lut_sub lut_1877 ({sk[521], n_n91, x43x, n_n1134, x248x, n_n1147, x6336x}, x5729x);
	defparam lut_1877.LUT_SIZE = 7;
	defparam lut_1877.mask = 128'h0707ffff1717ffffbfffbfffbfffffff;

	lut_sub lut_1883 ({sk[522], x104x, x157x, x289x, x5696x, x5697x}, x5707x);
	defparam lut_1883.LUT_SIZE = 6;
	defparam lut_1883.mask = 64'h3333ffff7fffffff;

	lut_sub lut_1889 ({sk[523], n_n93, n_n103, n_n84, x213x, x96x, x6389x}, x5705x);
	defparam lut_1889.LUT_SIZE = 7;
	defparam lut_1889.mask = 128'h0707ffff1717ffffbfbfbfbfbfbfbfff;

	lut_sub lut_1894 ({sk[524], n_n38, n_n64, x239x, x5694x, x5695x, x6379x}, x5706x);
	defparam lut_1894.LUT_SIZE = 7;
	defparam lut_1894.mask = 128'h0707ffff1717ffffbfbfbfbfbfbfbfff;

	lut_sub lut_1899 ({sk[525], n_n101, x40x, x255x, x336x, x71x, x100x}, x5727x);
	defparam lut_1899.LUT_SIZE = 7;
	defparam lut_1899.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_1905 ({sk[526], n_n78, n_n1172, x23x, x160x, x166x, x121x}, x5728x);
	defparam lut_1905.LUT_SIZE = 7;
	defparam lut_1905.mask = 128'h0707ffff1717ffff7f7fffff7fffffff;

	lut_sub lut_1911 ({sk[527], i_5_, i_6_, i_3_}, x354x);
	defparam lut_1911.LUT_SIZE = 4;
	defparam lut_1911.mask = 16'h1f40;

	lut_sub lut_1913 ({sk[528], i_7_, i_8_, i_6_, n_n94, n_n74}, n_n1006);
	defparam lut_1913.LUT_SIZE = 6;
	defparam lut_1913.mask = 64'h3333ffff00000001;

	lut_sub lut_1915 ({sk[529], i_7_, i_8_, i_6_, n_n81, n_n90, x149x}, n_n296);
	defparam lut_1915.LUT_SIZE = 7;
	defparam lut_1915.mask = 128'h0707ffff1717ffff5555555555575555;

	lut_sub lut_1918 ({sk[530], i_3_, n_n58, n_n78, n_n83, x33x, n_n1002}, x6392x);
	defparam lut_1918.LUT_SIZE = 7;
	defparam lut_1918.mask = 128'h0707ffff1717ffffaa88aa88aa88a080;

	lut_sub lut_1925 ({sk[531], x188x, x114x, n_n1006, n_n296, x6392x}, x5748x);
	defparam lut_1925.LUT_SIZE = 6;
	defparam lut_1925.mask = 64'h3333ffffbfffffff;

	lut_sub lut_1931 ({sk[532], i_7_, i_8_, i_1_, i_2_, i_0_}, x129x);
	defparam lut_1931.LUT_SIZE = 6;
	defparam lut_1931.mask = 64'h3333ffff00040000;

	lut_sub lut_1933 ({sk[533], i_7_, i_8_, i_6_, n_n100, n_n77, x29x}, x193x);
	defparam lut_1933.LUT_SIZE = 7;
	defparam lut_1933.mask = 128'h0707ffff1717ffff0003000000550000;

	lut_sub lut_1936 ({sk[534], i_7_, i_8_, i_6_, n_n103, n_n77, x53x}, x5391x);
	defparam lut_1936.LUT_SIZE = 7;
	defparam lut_1936.mask = 128'h0707ffff1717ffff5500550300000003;

	lut_sub lut_1939 ({sk[535], i_7_, i_8_, i_6_, i_3_, n_n100, x109x}, n_n957);
	defparam lut_1939.LUT_SIZE = 7;
	defparam lut_1939.mask = 128'h0707ffff1717ffff0000000100000000;

	lut_sub lut_1941 ({sk[536], i_7_, i_8_, i_6_, n_n103, n_n102, x86x}, x79x);
	defparam lut_1941.LUT_SIZE = 7;
	defparam lut_1941.mask = 128'h0707ffff1717ffff0000005500030000;

	lut_sub lut_1944 ({sk[537], i_7_, i_8_, i_6_, n_n83, x109x, n_n67}, x103x);
	defparam lut_1944.LUT_SIZE = 7;
	defparam lut_1944.mask = 128'h0707ffff1717ffff0000000000130000;

	lut_sub lut_1947 ({sk[538], i_7_, i_8_, i_6_, n_n84, n_n85, x73x}, x161x);
	defparam lut_1947.LUT_SIZE = 7;
	defparam lut_1947.mask = 128'h0707ffff1717ffff0055000300000000;

	lut_sub lut_1950 ({sk[539], i_7_, i_8_, i_6_, x34x}, n_n1068);
	defparam lut_1950.LUT_SIZE = 5;
	defparam lut_1950.mask = 32'h0fff0001;

	lut_sub lut_1952 ({sk[540], i_7_, i_8_, i_6_, x34x, n_n87, n_n67}, x266x);
	defparam lut_1952.LUT_SIZE = 7;
	defparam lut_1952.mask = 128'h0707ffff1717ffff000011110000000f;

	lut_sub lut_1955 ({sk[541], x148x, x114x, n_n1026, x286x, x6370x}, x5795x);
	defparam lut_1955.LUT_SIZE = 6;
	defparam lut_1955.mask = 64'h3333ffffbfffffff;

	lut_sub lut_1961 ({sk[542], n_n95, x24x, x274x, n_n1014, x277x, x98x}, x5793x);
	defparam lut_1961.LUT_SIZE = 7;
	defparam lut_1961.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_1967 ({sk[543], n_n93, x76x, n_n1045, x154x, x212x, x280x}, x5794x);
	defparam lut_1967.LUT_SIZE = 7;
	defparam lut_1967.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_1973 ({sk[544], n_n91, x215x, x153x, x103x, x33x}, x5813x);
	defparam lut_1973.LUT_SIZE = 6;
	defparam lut_1973.mask = 64'h3333ffff3fff7fff;

	lut_sub lut_1978 ({sk[545], x145x, x131x, x5068x, x116x, n_n976, x147x}, x5814x);
	defparam lut_1978.LUT_SIZE = 7;
	defparam lut_1978.mask = 128'h0707ffff1717ffff7f7f7fffffffffff;

	lut_sub lut_1984 ({sk[546], n_n91, x81x, n_n956, x163x, x284x, x5798x}, x5815x);
	defparam lut_1984.LUT_SIZE = 7;
	defparam lut_1984.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_1990 ({sk[547], n_n95, x168x, n_n993, x237x, n_n1004, x6373x}, x5816x);
	defparam lut_1990.LUT_SIZE = 7;
	defparam lut_1990.mask = 128'h0707ffff1717ffffbbffffffbfffffff;

	lut_sub lut_1996 ({sk[548], x193x, x5391x, n_n652, x296x, x167x}, x5817x);
	defparam lut_1996.LUT_SIZE = 6;
	defparam lut_1996.mask = 64'h3333ffff7fffffff;

	lut_sub lut_2002 ({sk[549], i_7_, i_8_, i_6_, n_n103, n_n85, n_n77}, x71x);
	defparam lut_2002.LUT_SIZE = 7;
	defparam lut_2002.mask = 128'h0707ffff1717ffff0000000005110000;

	lut_sub lut_2005 ({sk[550], i_1_, i_2_, i_0_, n_n70, x127x, n_n1121}, x218x);
	defparam lut_2005.LUT_SIZE = 7;
	defparam lut_2005.mask = 128'h0707ffff1717ffff5555555555555557;

	lut_sub lut_2008 ({sk[551], i_6_, i_1_, i_0_, n_n58, x109x, x90x}, x5825x);
	defparam lut_2008.LUT_SIZE = 7;
	defparam lut_2008.mask = 128'h0707ffff1717ffff5557555555555555;

	lut_sub lut_2011 ({sk[552], n_n63, n_n1153, x19x, x71x, x218x, x5825x}, n_n385);
	defparam lut_2011.LUT_SIZE = 7;
	defparam lut_2011.mask = 128'h0707ffff1717ffff7f7fffff7fffffff;

	lut_sub lut_2017 ({sk[553], i_7_, i_8_, i_0_, n_n74, x63x, n_n67}, x5835x);
	defparam lut_2017.LUT_SIZE = 7;
	defparam lut_2017.mask = 128'h0707ffff1717ffff00003333000a0000;

	lut_sub lut_2020 ({sk[554], x150x, n_n1047, x285x, n_n421, n_n1068, x5835x}, x5845x);
	defparam lut_2020.LUT_SIZE = 7;
	defparam lut_2020.mask = 128'h0707ffff1717ffff7fffffffffffffff;

	lut_sub lut_2027 ({sk[555], i_7_, i_8_, i_6_, n_n74, n_n85, n_n1169}, x92x);
	defparam lut_2027.LUT_SIZE = 7;
	defparam lut_2027.mask = 128'h0707ffff1717ffff5555575555555555;

	lut_sub lut_2030 ({sk[556], i_7_, i_8_, i_1_, i_2_, i_0_}, x62x);
	defparam lut_2030.LUT_SIZE = 6;
	defparam lut_2030.mask = 64'h3333ffff10000000;

	lut_sub lut_2032 ({sk[557], i_7_, i_8_, i_1_, i_2_, i_0_}, x316x);
	defparam lut_2032.LUT_SIZE = 6;
	defparam lut_2032.mask = 64'h3333ffff00000020;

	lut_sub lut_2034 ({sk[558], i_7_, i_8_, i_6_, x23x}, x335x);
	defparam lut_2034.LUT_SIZE = 5;
	defparam lut_2034.mask = 32'h0fff0040;

	lut_sub lut_2036 ({sk[559], n_n73, x26x, n_n102, n_n94, n_n63, x20x}, x5886x);
	defparam lut_2036.LUT_SIZE = 7;
	defparam lut_2036.mask = 128'h0707ffff1717ffff005700570057ffff;

	lut_sub lut_2040 ({sk[560], n_n58, n_n78, x76x, n_n1020, x81x, n_n1108}, x6387x);
	defparam lut_2040.LUT_SIZE = 7;
	defparam lut_2040.mask = 128'h0707ffff1717ffff5f5f5fff7f7f7fff;

	lut_sub lut_2052 ({sk[561], n_n101, n_n1120, x128x, x138x, x5886x, x6387x}, x5896x);
	defparam lut_2052.LUT_SIZE = 7;
	defparam lut_2052.mask = 128'h0707ffff1717ffff7f7fffff7fffffff;

	lut_sub lut_2058 ({sk[562], i_7_, i_8_, i_6_, n_n103, n_n102}, n_n994);
	defparam lut_2058.LUT_SIZE = 6;
	defparam lut_2058.mask = 64'h3333ffff00010000;

	lut_sub lut_2060 ({sk[563], i_5_, n_n93, n_n73, n_n83, n_n76, x63x}, x149x);
	defparam lut_2060.LUT_SIZE = 7;
	defparam lut_2060.mask = 128'h0707ffff1717ffff00005555000c555d;

	lut_sub lut_2063 ({sk[564], n_n81, n_n103, n_n102, n_n63, n_n82, x103x}, x6376x);
	defparam lut_2063.LUT_SIZE = 7;
	defparam lut_2063.mask = 128'h0707ffff1717ffffaaaaaaa0aaaa8880;

	lut_sub lut_2069 ({sk[565], i_7_, i_8_, i_6_, n_n81, n_n103, x21x}, x100x);
	defparam lut_2069.LUT_SIZE = 7;
	defparam lut_2069.mask = 128'h0707ffff1717ffff0003000055000000;

	lut_sub lut_2072 ({sk[566], n_n52, n_n78, x27x, x34x, x264x, x22x}, x6374x);
	defparam lut_2072.LUT_SIZE = 7;
	defparam lut_2072.mask = 128'h0707ffff1717ffff333377ff3f3f7fff;

	lut_sub lut_2083 ({sk[567], i_7_, i_8_, n_n81, n_n100, n_n40, x107x}, x155x);
	defparam lut_2083.LUT_SIZE = 7;
	defparam lut_2083.mask = 128'h0707ffff1717ffff0055035700550055;

	lut_sub lut_2086 ({sk[568], i_3_, i_1_, i_2_, n_n95, x43x, x240x}, x157x);
	defparam lut_2086.LUT_SIZE = 7;
	defparam lut_2086.mask = 128'h0707ffff1717ffff0303035703030303;

	lut_sub lut_2089 ({sk[569], i_3_, i_1_, i_2_}, x174x);
	defparam lut_2089.LUT_SIZE = 4;
	defparam lut_2089.mask = 16'h1f04;

	lut_sub lut_2091 ({sk[570], i_7_, i_8_, i_6_, x26x, n_n83, n_n102}, x209x);
	defparam lut_2091.LUT_SIZE = 7;
	defparam lut_2091.mask = 128'h0707ffff1717ffff0000001100000f00;

	lut_sub lut_2094 ({sk[571], i_7_, i_8_, i_6_, n_n100, n_n84, x131x}, x210x);
	defparam lut_2094.LUT_SIZE = 7;
	defparam lut_2094.mask = 128'h0707ffff1717ffff0000000000030505;

	lut_sub lut_2097 ({sk[572], i_7_, i_8_, i_6_, n_n103, n_n77, x46x}, x213x);
	defparam lut_2097.LUT_SIZE = 7;
	defparam lut_2097.mask = 128'h0707ffff1717ffff5500000000030000;

	lut_sub lut_2100 ({sk[573], i_7_, i_8_, i_6_, x33x}, x336x);
	defparam lut_2100.LUT_SIZE = 5;
	defparam lut_2100.mask = 32'h0fff0001;

	lut_sub lut_2102 ({sk[574], i_7_, i_8_, i_6_, n_n103, x45x, n_n96}, x267x);
	defparam lut_2102.LUT_SIZE = 7;
	defparam lut_2102.mask = 128'h0707ffff1717ffff0033000500000000;

	lut_sub lut_2105 ({sk[575], i_5_, i_6_, i_3_}, x130x);
	defparam lut_2105.LUT_SIZE = 4;
	defparam lut_2105.mask = 16'h1f80;

	lut_sub lut_2107 ({sk[576], n_n58, n_n93, x58x, x66x, x23x, x130x}, x307x);
	defparam lut_2107.LUT_SIZE = 7;
	defparam lut_2107.mask = 128'h0707ffff1717ffff050505ff373737ff;

	lut_sub lut_2111 ({sk[577], i_7_, i_8_, i_5_, i_6_, i_4_}, x324x);
	defparam lut_2111.LUT_SIZE = 6;
	defparam lut_2111.mask = 64'h3333ffff00000080;

	lut_sub lut_2113 ({sk[578], i_7_, i_8_, i_3_, i_1_, i_2_, n_n87}, n_n1147);
	defparam lut_2113.LUT_SIZE = 7;
	defparam lut_2113.mask = 128'h0707ffff1717ffff0400000000000000;

	lut_sub lut_2115 ({sk[579], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x237x);
	defparam lut_2115.LUT_SIZE = 7;
	defparam lut_2115.mask = 128'h0707ffff1717ffff0010000000000000;

	lut_sub lut_2117 ({sk[580], i_7_, i_8_, n_n74, n_n85, n_n76, n_n1002}, x167x);
	defparam lut_2117.LUT_SIZE = 7;
	defparam lut_2117.mask = 128'h0707ffff1717ffff575755555555555f;

	lut_sub lut_2121 ({sk[581], i_8_, i_6_, x83x, x68x}, x287x);
	defparam lut_2121.LUT_SIZE = 5;
	defparam lut_2121.mask = 32'h0fff5755;

	lut_sub lut_2124 ({sk[582], i_7_, i_8_, i_6_, x39x, x282x, x65x}, x6369x);
	defparam lut_2124.LUT_SIZE = 7;
	defparam lut_2124.mask = 128'h0707ffff1717ffffcc88c0cccccccccc;

	lut_sub lut_2133 ({sk[583], i_7_, i_8_, i_6_, x83x}, n_n1088);
	defparam lut_2133.LUT_SIZE = 5;
	defparam lut_2133.mask = 32'h0fff0100;

	lut_sub lut_2135 ({sk[584], n_n81, n_n93, n_n85, x88x, x255x, x89x}, x5981x);
	defparam lut_2135.LUT_SIZE = 7;
	defparam lut_2135.mask = 128'h0707ffff1717ffff7f7f7f7f7f7f7fff;

	lut_sub lut_2140 ({sk[585], n_n78, n_n1297, x53x, x155x, x225x, x220x}, x5982x);
	defparam lut_2140.LUT_SIZE = 7;
	defparam lut_2140.mask = 128'h0707ffff1717ffff7f7fffff7fffffff;

	lut_sub lut_2146 ({sk[586], n_n78, n_n91, x82x, x22x, x6363x, x6364x}, x5983x);
	defparam lut_2146.LUT_SIZE = 7;
	defparam lut_2146.mask = 128'h0707ffff1717ffffeeeeeeffefefefff;

	lut_sub lut_2151 ({sk[587], x5965x, x5966x, x5967x, x5968x}, x5984x);
	defparam lut_2151.LUT_SIZE = 5;
	defparam lut_2151.mask = 32'h0fff7fff;

	lut_sub lut_2156 ({sk[588], x307x, x300x, x5969x, x5970x}, x5985x);
	defparam lut_2156.LUT_SIZE = 5;
	defparam lut_2156.mask = 32'h0fff7fff;

	lut_sub lut_2161 ({sk[589], i_7_, i_8_, i_6_, n_n84, n_n85, x33x}, x163x);
	defparam lut_2161.LUT_SIZE = 7;
	defparam lut_2161.mask = 128'h0707ffff1717ffff0000000055550003;

	lut_sub lut_2164 ({sk[590], i_7_, i_8_, i_6_, n_n103, n_n102, n_n978}, x284x);
	defparam lut_2164.LUT_SIZE = 7;
	defparam lut_2164.mask = 128'h0707ffff1717ffff5555555755555555;

	lut_sub lut_2167 ({sk[591], i_7_, i_8_, i_6_, n_n84, n_n83, x24x}, x94x);
	defparam lut_2167.LUT_SIZE = 7;
	defparam lut_2167.mask = 128'h0707ffff1717ffff0000000055000303;

	lut_sub lut_2170 ({sk[592], i_3_, i_2_, i_0_}, x242x);
	defparam lut_2170.LUT_SIZE = 4;
	defparam lut_2170.mask = 16'h1f02;

	lut_sub lut_2172 ({sk[593], i_7_, i_8_, i_6_, n_n84, n_n94, x171x}, x269x);
	defparam lut_2172.LUT_SIZE = 7;
	defparam lut_2172.mask = 128'h0707ffff1717ffff5755000000000000;

	lut_sub lut_2175 ({sk[594], i_7_, i_8_, i_6_, n_n81, x29x, n_n90}, x221x);
	defparam lut_2175.LUT_SIZE = 7;
	defparam lut_2175.mask = 128'h0707ffff1717ffff3300000000050000;

	lut_sub lut_2178 ({sk[595], i_7_, i_5_, i_6_, i_3_, i_4_, n_n85}, n_n976);
	defparam lut_2178.LUT_SIZE = 7;
	defparam lut_2178.mask = 128'h0707ffff1717ffff0010000000000000;

	lut_sub lut_2180 ({sk[596], i_7_, i_8_, i_6_, x86x, x347x}, x144x);
	defparam lut_2180.LUT_SIZE = 6;
	defparam lut_2180.mask = 64'h3333ffff00300005;

	lut_sub lut_2183 ({sk[597], i_5_, i_3_, i_4_, n_n93, n_n103}, n_n999);
	defparam lut_2183.LUT_SIZE = 6;
	defparam lut_2183.mask = 64'h3333ffff00001000;

	lut_sub lut_2185 ({sk[598], i_7_, i_8_, i_6_, x40x}, n_n1004);
	defparam lut_2185.LUT_SIZE = 5;
	defparam lut_2185.mask = 32'h0fff0100;

	lut_sub lut_2187 ({sk[599], i_7_, i_8_, i_6_, i_3_, n_n94, x109x}, n_n1181);
	defparam lut_2187.LUT_SIZE = 7;
	defparam lut_2187.mask = 128'h0707ffff1717ffff1000000000000000;

	lut_sub lut_2189 ({sk[600], i_5_, i_3_, i_4_}, x194x);
	defparam lut_2189.LUT_SIZE = 4;
	defparam lut_2189.mask = 16'h1f24;

	lut_sub lut_2192 ({sk[601], i_7_, i_8_, i_6_, x57x, x86x}, x205x);
	defparam lut_2192.LUT_SIZE = 6;
	defparam lut_2192.mask = 64'h3333ffff53000000;

	lut_sub lut_2195 ({sk[602], i_7_, i_8_, i_6_, n_n103, n_n102}, n_n984);
	defparam lut_2195.LUT_SIZE = 6;
	defparam lut_2195.mask = 64'h3333ffff00100000;

	lut_sub lut_2197 ({sk[603], i_5_, i_3_, i_4_, n_n83, n_n85, n_n82}, x274x);
	defparam lut_2197.LUT_SIZE = 7;
	defparam lut_2197.mask = 128'h0707ffff1717ffff0000000011000005;

	lut_sub lut_2200 ({sk[604], i_7_, i_8_, i_6_, n_n81, n_n103}, n_n1009);
	defparam lut_2200.LUT_SIZE = 6;
	defparam lut_2200.mask = 64'h3333ffff00000001;

	lut_sub lut_2202 ({sk[605], i_5_, i_6_, i_3_}, x4871x);
	defparam lut_2202.LUT_SIZE = 4;
	defparam lut_2202.mask = 16'h1f02;

	lut_sub lut_2204 ({sk[606], i_7_, i_8_, i_5_, i_6_, i_4_}, x339x);
	defparam lut_2204.LUT_SIZE = 6;
	defparam lut_2204.mask = 64'h3333ffff00800000;

	lut_sub lut_2206 ({sk[607], i_7_, i_8_, i_5_, i_6_, i_4_}, x315x);
	defparam lut_2206.LUT_SIZE = 6;
	defparam lut_2206.mask = 64'h3333ffff00000400;

	lut_sub lut_2208 ({sk[608], i_1_, i_2_, i_0_, n_n74, n_n95, x240x}, x59x);
	defparam lut_2208.LUT_SIZE = 7;
	defparam lut_2208.mask = 128'h0707ffff1717ffff0055000003000000;

	lut_sub lut_2211 ({sk[609], i_7_, i_5_, i_6_, i_4_, n_n982, n_n53}, x200x);
	defparam lut_2211.LUT_SIZE = 7;
	defparam lut_2211.mask = 128'h0707ffff1717ffff3333333333337333;

	lut_sub lut_2214 ({sk[610], i_7_, i_8_, i_6_, x109x, n_n969, n_n67}, x223x);
	defparam lut_2214.LUT_SIZE = 7;
	defparam lut_2214.mask = 128'h0707ffff1717ffff3333333333373333;

	lut_sub lut_2217 ({sk[611], i_1_, i_2_, i_0_, x77x, n_n947, x312x}, x5399x);
	defparam lut_2217.LUT_SIZE = 7;
	defparam lut_2217.mask = 128'h0707ffff1717ffff3333333333333337;

	lut_sub lut_2220 ({sk[612], i_7_, i_8_, i_6_, x76x}, n_n1013);
	defparam lut_2220.LUT_SIZE = 5;
	defparam lut_2220.mask = 32'h0fff1000;

	lut_sub lut_2222 ({sk[613], i_7_, i_8_, i_6_, n_n81, n_n100}, n_n1014);
	defparam lut_2222.LUT_SIZE = 6;
	defparam lut_2222.mask = 64'h3333ffff10000000;

	lut_sub lut_2224 ({sk[614], i_5_, i_6_, i_4_, n_n64, n_n85, x62x}, x152x);
	defparam lut_2224.LUT_SIZE = 7;
	defparam lut_2224.mask = 128'h0707ffff1717ffff0000000355000000;

	lut_sub lut_2227 ({sk[615], i_7_, i_8_, i_3_, i_2_, i_0_, n_n79}, n_n1002);
	defparam lut_2227.LUT_SIZE = 7;
	defparam lut_2227.mask = 128'h0707ffff1717ffff0000000100000000;

	lut_sub lut_2229 ({sk[616], i_7_, i_8_, i_6_, n_n96, n_n85, x171x}, x5613x);
	defparam lut_2229.LUT_SIZE = 7;
	defparam lut_2229.mask = 128'h0707ffff1717ffff0000550003000000;

	lut_sub lut_2232 ({sk[617], i_7_, i_8_, i_6_, i_3_, n_n83, x21x}, x164x);
	defparam lut_2232.LUT_SIZE = 7;
	defparam lut_2232.mask = 128'h0707ffff1717ffff0000000000003055;

	lut_sub lut_2235 ({sk[618], i_7_, i_8_, i_5_, i_6_, n_n83, n_n1046}, x277x);
	defparam lut_2235.LUT_SIZE = 7;
	defparam lut_2235.mask = 128'h0707ffff1717ffff5755555555555555;

	lut_sub lut_2238 ({sk[619], i_7_, i_8_, i_3_, i_1_, i_0_, n_n71}, n_n1026);
	defparam lut_2238.LUT_SIZE = 7;
	defparam lut_2238.mask = 128'h0707ffff1717ffff0000000004000000;

	lut_sub lut_2240 ({sk[620], i_7_, i_6_, i_3_, i_4_, n_n85}, x1581x);
	defparam lut_2240.LUT_SIZE = 6;
	defparam lut_2240.mask = 64'h3333ffff00001000;

	lut_sub lut_2242 ({sk[621], i_7_, i_8_, i_6_, i_3_, i_4_, i_0_}, x6359x);
	defparam lut_2242.LUT_SIZE = 7;
	defparam lut_2242.mask = 128'h0707ffff1717fffffffffffffbffffff;

	lut_sub lut_2257 ({sk[622], i_3_, i_1_, i_0_, x234x, x1581x, x6359x}, x288x);
	defparam lut_2257.LUT_SIZE = 7;
	defparam lut_2257.mask = 128'h0707ffff1717ffff3333bfbb3333bbbb;

	lut_sub lut_2261 ({sk[623], i_2_, i_0_}, x327x);
	defparam lut_2261.LUT_SIZE = 3;
	defparam lut_2261.mask = 8'h31;

	lut_sub lut_2263 ({sk[624], i_7_, i_1_, i_2_, i_0_, n_n76, n_n1004}, x203x);
	defparam lut_2263.LUT_SIZE = 7;
	defparam lut_2263.mask = 128'h0707ffff1717ffff5555555755555555;

	lut_sub lut_2266 ({sk[625], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x124x);
	defparam lut_2266.LUT_SIZE = 7;
	defparam lut_2266.mask = 128'h0707ffff1717ffff0000000000220000;

	lut_sub lut_2269 ({sk[626], i_1_, i_2_, i_0_, n_n91, n_n77, x34x}, x225x);
	defparam lut_2269.LUT_SIZE = 7;
	defparam lut_2269.mask = 128'h0707ffff1717ffff0505050705050505;

	lut_sub lut_2272 ({sk[627], n_n93, n_n78, n_n102, n_n94, n_n74, n_n90}, x96x);
	defparam lut_2272.LUT_SIZE = 7;
	defparam lut_2272.mask = 128'h0707ffff1717ffff0000005503030357;

	lut_sub lut_2275 ({sk[628], i_7_, i_6_, i_3_, n_n83, x109x, n_n1009}, x98x);
	defparam lut_2275.LUT_SIZE = 7;
	defparam lut_2275.mask = 128'h0707ffff1717ffff5555555555555755;

	lut_sub lut_2278 ({sk[629], i_7_, i_6_, i_3_, i_4_, n_n103, n_n1043}, x154x);
	defparam lut_2278.LUT_SIZE = 7;
	defparam lut_2278.mask = 128'h0707ffff1717ffff5555555575555555;

	lut_sub lut_2281 ({sk[630], i_7_, i_8_, i_6_, i_3_, n_n83, x53x}, x212x);
	defparam lut_2281.LUT_SIZE = 7;
	defparam lut_2281.mask = 128'h0707ffff1717ffff0000000000305500;

	lut_sub lut_2284 ({sk[631], i_7_, i_8_, i_6_, n_n102, n_n94, x171x}, x280x);
	defparam lut_2284.LUT_SIZE = 7;
	defparam lut_2284.mask = 128'h0707ffff1717ffff0003550000030000;

	lut_sub lut_2287 ({sk[632], i_7_, i_8_, i_6_, n_n1020, x23x, x33x}, x6370x);
	defparam lut_2287.LUT_SIZE = 7;
	defparam lut_2287.mask = 128'h0707ffff1717ffffa0f0f0f0f0c0f0c0;

	lut_sub lut_2298 ({sk[633], n_n91, n_n103, n_n84, n_n83, x90x, n_n1164}, x6340x);
	defparam lut_2298.LUT_SIZE = 7;
	defparam lut_2298.mask = 128'h0707ffff1717ffff8888888888808800;

	lut_sub lut_2302 ({sk[634], i_7_, i_8_, i_6_, x27x, n_n71, x242x}, x119x);
	defparam lut_2302.LUT_SIZE = 7;
	defparam lut_2302.mask = 128'h0707ffff1717ffff0000000000001f11;

	lut_sub lut_2305 ({sk[635], i_7_, i_8_, i_6_, n_n83, n_n74, x33x}, x160x);
	defparam lut_2305.LUT_SIZE = 7;
	defparam lut_2305.mask = 128'h0707ffff1717ffff0003000000035500;

	lut_sub lut_2308 ({sk[636], i_7_, i_8_, i_6_, n_n83, n_n77, n_n90}, x166x);
	defparam lut_2308.LUT_SIZE = 7;
	defparam lut_2308.mask = 128'h0707ffff1717ffff0000000003000011;

	lut_sub lut_2311 ({sk[637], i_7_, i_8_, i_6_, n_n74, n_n85, x65x}, x220x);
	defparam lut_2311.LUT_SIZE = 7;
	defparam lut_2311.mask = 128'h0707ffff1717ffff0003000055550000;

	lut_sub lut_2314 ({sk[638], i_7_, i_8_, i_6_, n_n81, n_n100, x33x}, x5696x);
	defparam lut_2314.LUT_SIZE = 7;
	defparam lut_2314.mask = 128'h0707ffff1717ffff0000000300550000;

	lut_sub lut_2317 ({sk[639], i_7_, i_8_, i_6_, n_n74, n_n85, x21x}, x5697x);
	defparam lut_2317.LUT_SIZE = 7;
	defparam lut_2317.mask = 128'h0707ffff1717ffff0003005500000000;

	lut_sub lut_2320 ({sk[640], i_7_, i_8_, i_6_, n_n83, n_n102, x44x}, x101x);
	defparam lut_2320.LUT_SIZE = 7;
	defparam lut_2320.mask = 128'h0707ffff1717ffff0000550003000000;

	lut_sub lut_2323 ({sk[641], i_5_, i_3_, i_1_, i_2_, i_0_, n_n93}, x899x);
	defparam lut_2323.LUT_SIZE = 7;
	defparam lut_2323.mask = 128'h0707ffff1717ffff0000000000000001;

	lut_sub lut_2325 ({sk[642], i_7_, i_8_, i_6_, n_n94, x109x, x899x}, x102x);
	defparam lut_2325.LUT_SIZE = 7;
	defparam lut_2325.mask = 128'h0707ffff1717ffff5555555555555557;

	lut_sub lut_2328 ({sk[643], i_7_, i_8_, i_6_, n_n100, n_n74, x82x}, x283x);
	defparam lut_2328.LUT_SIZE = 7;
	defparam lut_2328.mask = 128'h0707ffff1717ffff0055000000000300;

	lut_sub lut_2331 ({sk[644], i_7_, i_8_, i_3_, i_1_, i_2_, n_n40}, x1107x);
	defparam lut_2331.LUT_SIZE = 7;
	defparam lut_2331.mask = 128'h0707ffff1717ffff0000000000000001;

	lut_sub lut_2333 ({sk[645], i_8_, i_5_, i_3_, i_1_, i_0_, n_n52}, x1442x);
	defparam lut_2333.LUT_SIZE = 7;
	defparam lut_2333.mask = 128'h0707ffff1717ffff0000000000000001;

	lut_sub lut_2335 ({sk[646], i_7_, i_8_, i_5_, i_4_, n_n80}, x1444x);
	defparam lut_2335.LUT_SIZE = 6;
	defparam lut_2335.mask = 64'h3333ffff04000000;

	lut_sub lut_2337 ({sk[647], n_n80, n_n75, n_n81, x75x, x192x, x337x}, x4847x);
	defparam lut_2337.LUT_SIZE = 7;
	defparam lut_2337.mask = 128'h0707ffff1717ffff0000000c5555555d;

	lut_sub lut_2340 ({sk[648], i_7_, i_8_, i_6_, i_4_, x253x, x311x}, x4848x);
	defparam lut_2340.LUT_SIZE = 7;
	defparam lut_2340.mask = 128'h0707ffff1717ffff0000000005370033;

	lut_sub lut_2343 ({sk[649], i_7_, i_8_, i_6_, n_n81, n_n83, x64x}, x4850x);
	defparam lut_2343.LUT_SIZE = 7;
	defparam lut_2343.mask = 128'h0707ffff1717ffff0055000000030003;

	lut_sub lut_2346 ({sk[650], n_n101, n_n78, x32x, x40x, x55x, x58x}, x4861x);
	defparam lut_2346.LUT_SIZE = 7;
	defparam lut_2346.mask = 128'h0707ffff1717ffff00550f5f77777f7f;

	lut_sub lut_2351 ({sk[651], i_7_, i_8_, i_6_, x76x, x57x, x42x}, x6393x);
	defparam lut_2351.LUT_SIZE = 7;
	defparam lut_2351.mask = 128'h0707ffff1717ffff0033007f00550000;

	lut_sub lut_2359 ({sk[652], i_8_, n_n1022, n_n1052, x70x, x277x, x288x}, x4897x);
	defparam lut_2359.LUT_SIZE = 7;
	defparam lut_2359.mask = 128'h0707ffff1717ffff7fffffff77ffffff;

	lut_sub lut_2365 ({sk[653], n_n91, x53x, x66x, n_n1059, n_n1009, x4871x}, x6357x);
	defparam lut_2365.LUT_SIZE = 7;
	defparam lut_2365.mask = 128'h0707ffff1717ffffc080c080c0800000;

	lut_sub lut_2370 ({sk[654], n_n82, n_n1048, x237x, n_n1042, n_n1013, x6357x}, x4898x);
	defparam lut_2370.LUT_SIZE = 7;
	defparam lut_2370.mask = 128'h0707ffff1717ffffbfbfffffbfffffff;

	lut_sub lut_2376 ({sk[655], n_n93, n_n982, x24x, x204x, x202x, x203x}, x4917x);
	defparam lut_2376.LUT_SIZE = 7;
	defparam lut_2376.mask = 128'h0707ffff1717ffff7f7fffff7fffffff;

	lut_sub lut_2382 ({sk[656], n_n63, x42x, n_n95, x41x, x86x, n_n978}, x6355x);
	defparam lut_2382.LUT_SIZE = 7;
	defparam lut_2382.mask = 128'h0707ffff1717ffffaaa0aa0088808800;

	lut_sub lut_2387 ({sk[657], x253x, n_n82, n_n976, n_n984, n_n1006, x6355x}, x4918x);
	defparam lut_2387.LUT_SIZE = 7;
	defparam lut_2387.mask = 128'h0707ffff1717ffffbfffbfffbfffffff;

	lut_sub lut_2393 ({sk[658], i_7_, i_8_, i_6_, n_n100, n_n102, x49x}, x4925x);
	defparam lut_2393.LUT_SIZE = 7;
	defparam lut_2393.mask = 128'h0707ffff1717ffff0000035500000300;

	lut_sub lut_2396 ({sk[659], i_7_, i_8_, i_6_, x26x, n_n100, n_n84}, x4926x);
	defparam lut_2396.LUT_SIZE = 7;
	defparam lut_2396.mask = 128'h0707ffff1717ffff000011000f000000;

	lut_sub lut_2399 ({sk[660], i_7_, i_8_, i_6_, n_n81, n_n103, x21x}, x4927x);
	defparam lut_2399.LUT_SIZE = 7;
	defparam lut_2399.mask = 128'h0707ffff1717ffff0300000000550000;

	lut_sub lut_2402 ({sk[661], i_5_, n_n58, n_n78, n_n100, n_n102, x338x}, x4967x);
	defparam lut_2402.LUT_SIZE = 7;
	defparam lut_2402.mask = 128'h0707ffff1717ffff00001111000f111f;

	lut_sub lut_2405 ({sk[662], n_n81, n_n86, n_n1077, n_n1172, n_n1078, x108x}, x4974x);
	defparam lut_2405.LUT_SIZE = 7;
	defparam lut_2405.mask = 128'h0707ffff1717ffff3fff3fff3fff7fff;

	lut_sub lut_2410 ({sk[663], n_n73, x27x, x26x, n_n82, x19x, x29x}, x4978x);
	defparam lut_2410.LUT_SIZE = 7;
	defparam lut_2410.mask = 128'h0707ffff1717ffff07070f0f07ff0fff;

	lut_sub lut_2415 ({sk[664], n_n58, n_n102, n_n1081, n_n1279, n_n1297, n_n90}, x6356x);
	defparam lut_2415.LUT_SIZE = 7;
	defparam lut_2415.mask = 128'h0707ffff1717ffffc000c000c0008000;

	lut_sub lut_2419 ({sk[665], n_n91, x27x, n_n1324, x251x, x321x, x6356x}, x4981x);
	defparam lut_2419.LUT_SIZE = 7;
	defparam lut_2419.mask = 128'h0707ffff1717ffffbfffbfffbfffffff;

	lut_sub lut_2425 ({sk[666], n_n74, x37x, x127x, x328x, x4967x, x4978x}, x4982x);
	defparam lut_2425.LUT_SIZE = 7;
	defparam lut_2425.mask = 128'h0707ffff1717ffff777f777f777fffff;

	lut_sub lut_2430 ({sk[667], i_7_, i_8_, i_6_, n_n84, x42x, n_n85}, x4998x);
	defparam lut_2430.LUT_SIZE = 7;
	defparam lut_2430.mask = 128'h0707ffff1717ffff0033000000000500;

	lut_sub lut_2433 ({sk[668], i_7_, i_8_, i_6_, n_n103, n_n74, x4998x}, x5005x);
	defparam lut_2433.LUT_SIZE = 7;
	defparam lut_2433.mask = 128'h0707ffff1717ffff5555575755555555;

	lut_sub lut_2437 ({sk[669], n_n100, n_n102, n_n95, x128x, x44x, n_n1004}, x5024x);
	defparam lut_2437.LUT_SIZE = 7;
	defparam lut_2437.mask = 128'h0707ffff1717ffff557f557f557f55ff;

	lut_sub lut_2442 ({sk[670], n_n86, n_n63, x49x, n_n1204, x21x, x34x}, x6354x);
	defparam lut_2442.LUT_SIZE = 7;
	defparam lut_2442.mask = 128'h0707ffff1717fffff0f0a000c0c08000;

	lut_sub lut_2447 ({sk[671], i_7_, i_8_, i_6_, x27x, x73x, x124x}, x5059x);
	defparam lut_2447.LUT_SIZE = 7;
	defparam lut_2447.mask = 128'h0707ffff1717ffff0f55000000000033;

	lut_sub lut_2451 ({sk[672], n_n101, x64x, n_n95, x67x, n_n1146, n_n1164}, x6352x);
	defparam lut_2451.LUT_SIZE = 7;
	defparam lut_2451.mask = 128'h0707ffff1717ffff8880888088800000;

	lut_sub lut_2456 ({sk[673], i_7_, i_8_, i_6_, n_n74, x49x, n_n90}, x5091x);
	defparam lut_2456.LUT_SIZE = 7;
	defparam lut_2456.mask = 128'h0707ffff1717ffff0000003700330000;

	lut_sub lut_2460 ({sk[674], i_7_, i_8_, i_6_, x21x, x46x}, x5092x);
	defparam lut_2460.LUT_SIZE = 6;
	defparam lut_2460.mask = 64'h3333ffff03035000;

	lut_sub lut_2463 ({sk[675], x58x, n_n95, n_n1324, n_n1092, n_n1022, n_n1134}, x6366x);
	defparam lut_2463.LUT_SIZE = 7;
	defparam lut_2463.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_2477 ({sk[676], n_n81, n_n83, n_n82, n_n937, x1315x, n_n958}, x6384x);
	defparam lut_2477.LUT_SIZE = 7;
	defparam lut_2477.mask = 128'h0707ffff1717ffff8080808080808000;

	lut_sub lut_2481 ({sk[677], n_n74, x40x, n_n63, n_n1153, n_n1092, x107x}, x6383x);
	defparam lut_2481.LUT_SIZE = 7;
	defparam lut_2481.mask = 128'h0707ffff1717ffff3f3f3fff7f7f7fff;

	lut_sub lut_2493 ({sk[678], i_5_, i_3_, i_4_, n_n93, n_n90, x48x}, x5149x);
	defparam lut_2493.LUT_SIZE = 7;
	defparam lut_2493.mask = 128'h0707ffff1717ffff0000550000030000;

	lut_sub lut_2496 ({sk[679], i_7_, i_8_, i_1_, n_n1324, n_n1369, x72x}, x5156x);
	defparam lut_2496.LUT_SIZE = 7;
	defparam lut_2496.mask = 128'h0707ffff1717ffff7f3f3f3f3f3f3f3f;

	lut_sub lut_2500 ({sk[680], n_n101, x64x, n_n85, n_n82, x49x, x244x}, x6378x);
	defparam lut_2500.LUT_SIZE = 7;
	defparam lut_2500.mask = 128'h0707ffff1717ffffffaaf0a0cc88c080;

	lut_sub lut_2509 ({sk[681], n_n64, n_n100, n_n1204, n_n1128, n_n1184, n_n87}, x5179x);
	defparam lut_2509.LUT_SIZE = 7;
	defparam lut_2509.mask = 128'h0707ffff1717ffff3fff3fff3fff7fff;

	lut_sub lut_2514 ({sk[682], n_n84, n_n937, x1315x, n_n958, x317x, n_n999}, x6347x);
	defparam lut_2514.LUT_SIZE = 7;
	defparam lut_2514.mask = 128'h0707ffff1717ffffa000000080000000;

	lut_sub lut_2517 ({sk[683], i_7_, i_8_, i_6_, n_n103, n_n96, n_n90}, x5205x);
	defparam lut_2517.LUT_SIZE = 7;
	defparam lut_2517.mask = 128'h0707ffff1717ffff1100000000030000;

	lut_sub lut_2520 ({sk[684], i_7_, i_8_, i_6_, x325x, x49x, x241x}, x5206x);
	defparam lut_2520.LUT_SIZE = 7;
	defparam lut_2520.mask = 128'h0707ffff1717ffff0500003300000000;

	lut_sub lut_2523 ({sk[685], i_7_, i_8_, i_6_, x105x, x46x, x41x}, x6349x);
	defparam lut_2523.LUT_SIZE = 7;
	defparam lut_2523.mask = 128'h0707ffff1717fffff0a0f0f0c0f0f0c0;

	lut_sub lut_2534 ({sk[686], i_8_, i_5_, i_4_, n_n52, x75x, x252x}, x5283x);
	defparam lut_2534.LUT_SIZE = 7;
	defparam lut_2534.mask = 128'h0707ffff1717ffff5555555555555557;

	lut_sub lut_2537 ({sk[687], i_5_, i_6_, i_3_, n_n64, n_n90, x1107x}, x5288x);
	defparam lut_2537.LUT_SIZE = 7;
	defparam lut_2537.mask = 128'h0707ffff1717ffff5555555555555557;

	lut_sub lut_2540 ({sk[688], i_4_, n_n75, x75x, x311x, n_n77, x315x}, x5289x);
	defparam lut_2540.LUT_SIZE = 7;
	defparam lut_2540.mask = 128'h0707ffff1717ffff0011001100110f1f;

	lut_sub lut_2543 ({sk[689], i_1_, i_0_, n_n93, n_n102, x127x, x328x}, x5290x);
	defparam lut_2543.LUT_SIZE = 7;
	defparam lut_2543.mask = 128'h0707ffff1717ffff11111111111f1111;

	lut_sub lut_2546 ({sk[690], i_7_, i_8_, i_1_, i_2_, i_0_, n_n76}, x5291x);
	defparam lut_2546.LUT_SIZE = 7;
	defparam lut_2546.mask = 128'h0707ffff1717ffff0004000000001000;

	lut_sub lut_2549 ({sk[691], i_6_, i_3_, i_4_, x234x, x66x, x242x}, x5292x);
	defparam lut_2549.LUT_SIZE = 7;
	defparam lut_2549.mask = 128'h0707ffff1717ffff3705050505050505;

	lut_sub lut_2552 ({sk[692], i_5_, i_3_, i_4_, n_n93, n_n90, x85x}, x5293x);
	defparam lut_2552.LUT_SIZE = 7;
	defparam lut_2552.mask = 128'h0707ffff1717ffff0000030055005500;

	lut_sub lut_2555 ({sk[693], i_7_, i_8_, i_6_, n_n83, n_n102, x67x}, x5294x);
	defparam lut_2555.LUT_SIZE = 7;
	defparam lut_2555.mask = 128'h0707ffff1717ffff0000005503000000;

	lut_sub lut_2558 ({sk[694], i_5_, i_3_, i_4_, n_n93, n_n100, x32x}, x5295x);
	defparam lut_2558.LUT_SIZE = 7;
	defparam lut_2558.mask = 128'h0707ffff1717ffff0055030000000000;

	lut_sub lut_2561 ({sk[695], n_n101, n_n91, x57x, x42x, n_n77, x20x}, x5296x);
	defparam lut_2561.LUT_SIZE = 7;
	defparam lut_2561.mask = 128'h0707ffff1717ffff111111ff1f1f1fff;

	lut_sub lut_2565 ({sk[696], n_n78, n_n91, x82x, n_n1176, x22x, x336x}, x6346x);
	defparam lut_2565.LUT_SIZE = 7;
	defparam lut_2565.mask = 128'h0707ffff1717ffffa0a08080a0008000;

	lut_sub lut_2570 ({sk[697], i_8_, n_n81, n_n83, n_n85, n_n82, x28x}, x5321x);
	defparam lut_2570.LUT_SIZE = 7;
	defparam lut_2570.mask = 128'h0707ffff1717ffff0505053700000033;

	lut_sub lut_2573 ({sk[698], i_5_, i_3_, i_4_, n_n93, n_n103, n_n95}, x5323x);
	defparam lut_2573.LUT_SIZE = 7;
	defparam lut_2573.mask = 128'h0707ffff1717ffff0000000003000011;

	lut_sub lut_2576 ({sk[699], n_n64, n_n63, x42x, x109x, x338x, x83x}, x5352x);
	defparam lut_2576.LUT_SIZE = 7;
	defparam lut_2576.mask = 128'h0707ffff1717ffff555555ff575757ff;

	lut_sub lut_2580 ({sk[700], i_8_, x70x, x215x, x262x, x275x}, x5364x);
	defparam lut_2580.LUT_SIZE = 6;
	defparam lut_2580.mask = 64'h3333ffff7fff7f7f;

	lut_sub lut_2585 ({sk[701], n_n80, x245x, x38x, n_n1093, x234x, n_n958}, x6345x);
	defparam lut_2585.LUT_SIZE = 7;
	defparam lut_2585.mask = 128'h0707ffff1717ffffa0a0a00080808000;

	lut_sub lut_2590 ({sk[702], n_n82, n_n1074, n_n1087, n_n974, x74x, x6345x}, x5365x);
	defparam lut_2590.LUT_SIZE = 7;
	defparam lut_2590.mask = 128'h0707ffff1717ffffafffffffbfffffff;

	lut_sub lut_2596 ({sk[703], n_n101, n_n93, n_n989, x52x, x24x, n_n956}, x6344x);
	defparam lut_2596.LUT_SIZE = 7;
	defparam lut_2596.mask = 128'h0707ffff1717ffffaa008800a0008000;

	lut_sub lut_2601 ({sk[704], n_n91, x29x, n_n982, n_n1121, x236x, x6344x}, x5366x);
	defparam lut_2601.LUT_SIZE = 7;
	defparam lut_2601.mask = 128'h0707ffff1717ffffbfffbfffbfffffff;

	lut_sub lut_2607 ({sk[705], n_n93, n_n82, x29x, x237x, n_n976, n_n994}, x5383x);
	defparam lut_2607.LUT_SIZE = 7;
	defparam lut_2607.mask = 128'h0707ffff1717ffff77777f7f77ff7fff;

	lut_sub lut_2612 ({sk[706], n_n95, n_n993, x237x, x59x, x163x, x200x}, x5386x);
	defparam lut_2612.LUT_SIZE = 7;
	defparam lut_2612.mask = 128'h0707ffff1717ffff7f7fffff7fffffff;

	lut_sub lut_2618 ({sk[707], n_n91, x57x, x40x, n_n63, x223x, x5383x}, x5387x);
	defparam lut_2618.LUT_SIZE = 7;
	defparam lut_2618.mask = 128'h0707ffff1717ffff77777f7f77ff7fff;

	lut_sub lut_2623 ({sk[708], i_5_, i_3_, i_4_, n_n78, n_n85, x37x}, x5411x);
	defparam lut_2623.LUT_SIZE = 7;
	defparam lut_2623.mask = 128'h0707ffff1717ffff0000000000005700;

	lut_sub lut_2626 ({sk[709], n_n93, n_n100, n_n84, x208x, x209x, x210x}, x5419x);
	defparam lut_2626.LUT_SIZE = 7;
	defparam lut_2626.mask = 128'h0707ffff1717ffff7f7f7f7f7f7f7fff;

	lut_sub lut_2631 ({sk[710], i_7_, i_8_, i_6_, x57x, x51x, x63x}, x6343x);
	defparam lut_2631.LUT_SIZE = 7;
	defparam lut_2631.mask = 128'h0707ffff1717ffffffffffffff88ffc0;

	lut_sub lut_2637 ({sk[711], n_n91, x76x, x64x, n_n82, x5411x, x6343x}, x5420x);
	defparam lut_2637.LUT_SIZE = 7;
	defparam lut_2637.mask = 128'h0707ffff1717ffffbbbfbbbfbbbfffff;

	lut_sub lut_2642 ({sk[712], x99x, x205x, x119x, x122x}, x5438x);
	defparam lut_2642.LUT_SIZE = 5;
	defparam lut_2642.mask = 32'h0fff7fff;

	lut_sub lut_2647 ({sk[713], n_n93, x26x, x329x, n_n95, x43x, n_n1181}, x6342x);
	defparam lut_2647.LUT_SIZE = 7;
	defparam lut_2647.mask = 128'h0707ffff1717ffffa800a800a8000000;

	lut_sub lut_2652 ({sk[714], n_n93, n_n78, x45x, n_n1176, x22x, x6342x}, x5439x);
	defparam lut_2652.LUT_SIZE = 7;
	defparam lut_2652.mask = 128'h0707ffff1717ffffafafbfbfbfffbfff;

	lut_sub lut_2658 ({sk[715], i_7_, i_6_, i_3_, n_n1078, x325x, x330x}, x5460x);
	defparam lut_2658.LUT_SIZE = 7;
	defparam lut_2658.mask = 128'h0707ffff1717ffff0f0f0f0f0f1f0f0f;

	lut_sub lut_2661 ({sk[716], i_8_, i_5_, i_6_, i_4_, x241x, x355x}, x5467x);
	defparam lut_2661.LUT_SIZE = 7;
	defparam lut_2661.mask = 128'h0707ffff1717ffff5555555555557555;

	lut_sub lut_2664 ({sk[717], i_7_, i_8_, i_6_, n_n85, x127x, x21x}, x5468x);
	defparam lut_2664.LUT_SIZE = 7;
	defparam lut_2664.mask = 128'h0707ffff1717ffff0055035700000303;

	lut_sub lut_2667 ({sk[718], i_7_, i_8_, i_6_, n_n103, x325x, x44x}, x5469x);
	defparam lut_2667.LUT_SIZE = 7;
	defparam lut_2667.mask = 128'h0707ffff1717ffff0000005500000300;

	lut_sub lut_2670 ({sk[719], i_7_, i_8_, i_6_, x26x, x39x, x58x}, x5472x);
	defparam lut_2670.LUT_SIZE = 7;
	defparam lut_2670.mask = 128'h0707ffff1717ffff0f003f0f00000055;

	lut_sub lut_2675 ({sk[720], n_n91, x40x, n_n63, x53x, x319x, n_n1045}, x5475x);
	defparam lut_2675.LUT_SIZE = 7;
	defparam lut_2675.mask = 128'h0707ffff1717ffff777777ff7f7f7fff;

	lut_sub lut_2680 ({sk[721], n_n91, n_n100, n_n74, n_n1074, x282x, x5472x}, x5480x);
	defparam lut_2680.LUT_SIZE = 7;
	defparam lut_2680.mask = 128'h0707ffff1717ffff7f7f7f7f7f7f7fff;

	lut_sub lut_2685 ({sk[722], n_n93, n_n74, n_n90, n_n1125, x5460x, x5475x}, x5481x);
	defparam lut_2685.LUT_SIZE = 7;
	defparam lut_2685.mask = 128'h0707ffff1717ffff7f7f7f7f7f7f7fff;

	lut_sub lut_2690 ({sk[723], n_n91, x74x, n_n1122, x66x, x5442x, n_n1101}, x6341x);
	defparam lut_2690.LUT_SIZE = 7;
	defparam lut_2690.mask = 128'h0707ffff1717ffffa800a800a8000000;

	lut_sub lut_2695 ({sk[724], n_n81, n_n83, n_n82, n_n1118, x5467x, x6341x}, x5482x);
	defparam lut_2695.LUT_SIZE = 7;
	defparam lut_2695.mask = 128'h0707ffff1717ffffbfbfbfbfbfbfbfff;

	lut_sub lut_2700 ({sk[725], x188x, x141x, x142x, x150x, x5468x, x5469x}, x5483x);
	defparam lut_2700.LUT_SIZE = 7;
	defparam lut_2700.mask = 128'h0707ffff1717ffff7fffffffffffffff;

	lut_sub lut_2707 ({sk[726], i_8_, i_5_, i_4_, n_n38, n_n1153, x175x}, x5499x);
	defparam lut_2707.LUT_SIZE = 7;
	defparam lut_2707.mask = 128'h0707ffff1717ffff3733333333333333;

	lut_sub lut_2710 ({sk[727], i_7_, i_8_, n_n96, n_n85, n_n87, x174x}, x5519x);
	defparam lut_2710.LUT_SIZE = 7;
	defparam lut_2710.mask = 128'h0707ffff1717ffff0000000f00001111;

	lut_sub lut_2713 ({sk[728], i_7_, i_8_, i_6_, n_n81, n_n94, x49x}, x5520x);
	defparam lut_2713.LUT_SIZE = 7;
	defparam lut_2713.mask = 128'h0707ffff1717ffff0000000000550003;

	lut_sub lut_2716 ({sk[729], i_7_, i_8_, i_6_, n_n100, n_n102, n_n77}, x5522x);
	defparam lut_2716.LUT_SIZE = 7;
	defparam lut_2716.mask = 128'h0707ffff1717ffff0000030000000500;

	lut_sub lut_2719 ({sk[730], n_n101, n_n91, x64x, x46x, x51x, x74x}, x5529x);
	defparam lut_2719.LUT_SIZE = 7;
	defparam lut_2719.mask = 128'h0707ffff1717ffff00000f0f77ff7fff;

	lut_sub lut_2724 ({sk[731], n_n75, n_n71, x270x, n_n67, x200x, x152x}, x5554x);
	defparam lut_2724.LUT_SIZE = 7;
	defparam lut_2724.mask = 128'h0707ffff1717ffff77ff77ff77ff7fff;

	lut_sub lut_2729 ({sk[732], n_n82, x237x, x144x, n_n1013, x212x, x284x}, x5555x);
	defparam lut_2729.LUT_SIZE = 7;
	defparam lut_2729.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_2735 ({sk[733], i_8_, i_6_, n_n103, n_n77, n_n1059}, x5568x);
	defparam lut_2735.LUT_SIZE = 6;
	defparam lut_2735.mask = 64'h3333ffff55555557;

	lut_sub lut_2738 ({sk[734], n_n91, x64x, x254x, n_n1074, x68x, x138x}, x5580x);
	defparam lut_2738.LUT_SIZE = 7;
	defparam lut_2738.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_2744 ({sk[735], n_n82, x29x, n_n1087, x153x, x204x, x263x}, x5581x);
	defparam lut_2744.LUT_SIZE = 7;
	defparam lut_2744.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_2750 ({sk[736], i_8_, i_6_, n_n1093, x67x, n_n1057, n_n956}, x6339x);
	defparam lut_2750.LUT_SIZE = 7;
	defparam lut_2750.mask = 128'h0707ffff1717ffff8800880080008800;

	lut_sub lut_2754 ({sk[737], n_n82, x24x, n_n1043, n_n1101, n_n1060, x6339x}, x5582x);
	defparam lut_2754.LUT_SIZE = 7;
	defparam lut_2754.mask = 128'h0707ffff1717ffffbfffbfffbfffffff;

	lut_sub lut_2760 ({sk[738], x77x, n_n78, x39x, n_n1058, x81x, n_n939}, x6338x);
	defparam lut_2760.LUT_SIZE = 7;
	defparam lut_2760.mask = 128'h0707ffff1717ffffa0a08080a0008000;

	lut_sub lut_2765 ({sk[739], n_n74, n_n1046, n_n969, n_n971, x107x, x6338x}, x5583x);
	defparam lut_2765.LUT_SIZE = 7;
	defparam lut_2765.mask = 128'h0707ffff1717ffffafffffffbfffffff;

	lut_sub lut_2771 ({sk[740], n_n95, x41x, x115x, x97x, x125x, x5568x}, x5584x);
	defparam lut_2771.LUT_SIZE = 7;
	defparam lut_2771.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_2777 ({sk[741], n_n80, x234x, x298x, n_n421, n_n241, x116x}, x5585x);
	defparam lut_2777.LUT_SIZE = 7;
	defparam lut_2777.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_2783 ({sk[742], n_n81, n_n103, n_n82, n_n1047, n_n1013, n_n1014}, x5617x);
	defparam lut_2783.LUT_SIZE = 7;
	defparam lut_2783.mask = 128'h0707ffff1717ffff7f7f7f7f7f7f7fff;

	lut_sub lut_2788 ({sk[743], i_1_, n_n64, n_n91, n_n94, n_n77, n_n66}, x5633x);
	defparam lut_2788.LUT_SIZE = 7;
	defparam lut_2788.mask = 128'h0707ffff1717ffff0000050500330537;

	lut_sub lut_2791 ({sk[744], n_n93, n_n78, x81x, n_n1101, x65x, n_n978}, x6337x);
	defparam lut_2791.LUT_SIZE = 7;
	defparam lut_2791.mask = 128'h0707ffff1717ffffa0a0a00080808000;

	lut_sub lut_2796 ({sk[745], i_7_, i_8_, i_6_, x53x, x63x, x33x}, x6368x);
	defparam lut_2796.LUT_SIZE = 7;
	defparam lut_2796.mask = 128'h0707ffff1717fffff0ffc0cca0a0ffff;

	lut_sub lut_2807 ({sk[746], i_5_, i_3_, n_n38, n_n91, n_n94, x42x}, x5664x);
	defparam lut_2807.LUT_SIZE = 7;
	defparam lut_2807.mask = 128'h0707ffff1717ffff0505050505370505;

	lut_sub lut_2810 ({sk[747], i_5_, i_3_, i_4_, n_n91, n_n94}, x5668x);
	defparam lut_2810.LUT_SIZE = 6;
	defparam lut_2810.mask = 64'h3333ffff10110000;

	lut_sub lut_2813 ({sk[748], i_3_, n_n93, n_n83, x109x, x66x, n_n71}, x5669x);
	defparam lut_2813.LUT_SIZE = 7;
	defparam lut_2813.mask = 128'h0707ffff1717ffff111111111111111f;

	lut_sub lut_2816 ({sk[749], i_7_, i_8_, i_6_, x57x, n_n77, n_n90}, x5670x);
	defparam lut_2816.LUT_SIZE = 7;
	defparam lut_2816.mask = 128'h0707ffff1717ffff00000000000f1100;

	lut_sub lut_2819 ({sk[750], i_7_, i_8_, i_6_, x73x, x67x, x51x}, x6381x);
	defparam lut_2819.LUT_SIZE = 7;
	defparam lut_2819.mask = 128'h0707ffff1717ffffaaffaaffffffc0ff;

	lut_sub lut_2826 ({sk[751], i_7_, i_8_, n_n94, x38x, x174x, x130x}, x5694x);
	defparam lut_2826.LUT_SIZE = 7;
	defparam lut_2826.mask = 128'h0707ffff1717ffff0303035703030303;

	lut_sub lut_2829 ({sk[752], i_5_, i_6_, i_3_, i_4_, x66x, x107x}, x5695x);
	defparam lut_2829.LUT_SIZE = 7;
	defparam lut_2829.mask = 128'h0707ffff1717ffff3000000030050005;

	lut_sub lut_2832 ({sk[753], i_7_, i_8_, i_6_, x42x, x82x, x49x}, x6389x);
	defparam lut_2832.LUT_SIZE = 7;
	defparam lut_2832.mask = 128'h0707ffff1717ffffffffaaf0ffccffff;

	lut_sub lut_2846 ({sk[754], i_5_, n_n101, x26x, x328x, x24x, x28x}, x6379x);
	defparam lut_2846.LUT_SIZE = 7;
	defparam lut_2846.mask = 128'h0707ffff1717ffffffffcc00fafac800;

	lut_sub lut_2853 ({sk[755], n_n91, x333x, x22x, x174x, n_n1181, x339x}, x6336x);
	defparam lut_2853.LUT_SIZE = 7;
	defparam lut_2853.mask = 128'h0707ffff1717ffffc8c80000c8000000;

	lut_sub lut_2858 ({sk[756], i_7_, i_8_, i_6_, n_n83, n_n74, n_n1021}, x5738x);
	defparam lut_2858.LUT_SIZE = 7;
	defparam lut_2858.mask = 128'h0707ffff1717ffff5555555555555557;

	lut_sub lut_2861 ({sk[757], n_n93, x29x, n_n984, x152x, x151x, x202x}, x5746x);
	defparam lut_2861.LUT_SIZE = 7;
	defparam lut_2861.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_2867 ({sk[758], n_n58, x53x, n_n994, x98x, x280x, x5738x}, x5747x);
	defparam lut_2867.LUT_SIZE = 7;
	defparam lut_2867.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_2873 ({sk[759], i_7_, i_8_, i_6_, x245x, x109x, x67x}, x5758x);
	defparam lut_2873.LUT_SIZE = 7;
	defparam lut_2873.mask = 128'h0707ffff1717ffff0003000355550000;

	lut_sub lut_2876 ({sk[760], i_7_, i_8_, i_6_, x44x, x347x, n_n1117}, x5768x);
	defparam lut_2876.LUT_SIZE = 7;
	defparam lut_2876.mask = 128'h0707ffff1717ffff5555555555555f7f;

	lut_sub lut_2881 ({sk[761], n_n82, x29x, n_n1087, x79x, x91x, x103x}, x5771x);
	defparam lut_2881.LUT_SIZE = 7;
	defparam lut_2881.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_2887 ({sk[762], n_n91, x29x, n_n939, x162x, x161x, x266x}, x5772x);
	defparam lut_2887.LUT_SIZE = 7;
	defparam lut_2887.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_2893 ({sk[763], n_n1077, n_n1081, n_n1120, n_n1122, x66x, x5442x}, x6391x);
	defparam lut_2893.LUT_SIZE = 7;
	defparam lut_2893.mask = 128'h0707ffff1717ffff1fffffffffffffff;

	lut_sub lut_2907 ({sk[764], n_n64, n_n100, x241x, n_n982, n_n87, x6391x}, x5773x);
	defparam lut_2907.LUT_SIZE = 7;
	defparam lut_2907.mask = 128'h0707ffff1717ffff5f5f5f5f5f7f7f7f;

	lut_sub lut_2912 ({sk[765], x55x, n_n95, n_n1132, n_n971, n_n980, x5768x}, x5774x);
	defparam lut_2912.LUT_SIZE = 7;
	defparam lut_2912.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_2918 ({sk[766], x256x, x215x, x291x, x141x, x142x, x5758x}, x5775x);
	defparam lut_2918.LUT_SIZE = 7;
	defparam lut_2918.mask = 128'h0707ffff1717ffff7fffffffffffffff;

	lut_sub lut_2925 ({sk[767], i_5_, i_4_, i_1_, n_n80, n_n58, x234x}, x5798x);
	defparam lut_2925.LUT_SIZE = 7;
	defparam lut_2925.mask = 128'h0707ffff1717ffff0537050505050505;

	lut_sub lut_2928 ({sk[768], n_n93, n_n83, x64x, n_n95, n_n77, x63x}, x6373x);
	defparam lut_2928.LUT_SIZE = 7;
	defparam lut_2928.mask = 128'h0707ffff1717fffffff0fff0aaa08880;

	lut_sub lut_2935 ({sk[769], n_n82, x29x, n_n1087, x263x, x161x, x102x}, x5843x);
	defparam lut_2935.LUT_SIZE = 7;
	defparam lut_2935.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_2941 ({sk[770], n_n91, x26x, n_n100, n_n84, n_n1091, x83x}, x6335x);
	defparam lut_2941.LUT_SIZE = 7;
	defparam lut_2941.mask = 128'h0707ffff1717ffffcccccccc88800000;

	lut_sub lut_2945 ({sk[771], n_n82, n_n1109, x24x, x355x, n_n1117, x6335x}, x5844x);
	defparam lut_2945.LUT_SIZE = 7;
	defparam lut_2945.mask = 128'h0707ffff1717ffffbfbfffffbfffffff;

	lut_sub lut_2951 ({sk[772], i_5_, i_6_, i_3_, n_n93, x22x, x316x}, x5852x);
	defparam lut_2951.LUT_SIZE = 7;
	defparam lut_2951.mask = 128'h0707ffff1717ffff0303030303030357;

	lut_sub lut_2954 ({sk[773], i_7_, i_8_, i_1_, i_2_, i_0_, n_n76}, x5853x);
	defparam lut_2954.LUT_SIZE = 7;
	defparam lut_2954.mask = 128'h0707ffff1717ffff0004000000000010;

	lut_sub lut_2957 ({sk[774], i_7_, i_8_, i_6_, n_n100, n_n102, n_n96}, x5854x);
	defparam lut_2957.LUT_SIZE = 7;
	defparam lut_2957.mask = 128'h0707ffff1717ffff0000030500030000;

	lut_sub lut_2961 ({sk[775], i_7_, i_8_, i_6_, x45x, x49x}, x5855x);
	defparam lut_2961.LUT_SIZE = 6;
	defparam lut_2961.mask = 64'h3333ffff00305000;

	lut_sub lut_2964 ({sk[776], i_7_, i_8_, i_6_, n_n103, n_n84, x21x}, x5857x);
	defparam lut_2964.LUT_SIZE = 7;
	defparam lut_2964.mask = 128'h0707ffff1717ffff0000000055030003;

	lut_sub lut_2967 ({sk[777], x222x, x185x, x120x, x92x}, x5868x);
	defparam lut_2967.LUT_SIZE = 5;
	defparam lut_2967.mask = 32'h0fff7fff;

	lut_sub lut_2972 ({sk[778], i_7_, i_8_, i_6_, x82x, x49x, x86x}, x6380x);
	defparam lut_2972.LUT_SIZE = 7;
	defparam lut_2972.mask = 128'h0707ffff1717ffffccfffff0ffffaaff;

	lut_sub lut_2987 ({sk[779], n_n78, n_n84, n_n90, x158x, x159x, x6380x}, x5869x);
	defparam lut_2987.LUT_SIZE = 7;
	defparam lut_2987.mask = 128'h0707ffff1717ffffbfbfbfbfbfbfbfff;

	lut_sub lut_2992 ({sk[780], i_7_, i_8_, i_6_, x46x, x86x, x128x}, x6375x);
	defparam lut_2992.LUT_SIZE = 7;
	defparam lut_2992.mask = 128'h0707ffff1717ffffccffffa0ffffffff;

	lut_sub lut_3001 ({sk[781], n_n82, x23x, x5852x, x5853x, x6375x}, x5870x);
	defparam lut_3001.LUT_SIZE = 6;
	defparam lut_3001.mask = 64'h3333ffffbfbfbfff;

	lut_sub lut_3006 ({sk[782], n_n91, x39x, x24x, x5854x, x5855x, x5857x}, x5871x);
	defparam lut_3006.LUT_SIZE = 7;
	defparam lut_3006.mask = 128'h0707ffff1717ffff7f7f7f7f7fffffff;

	lut_sub lut_3012 ({sk[783], n_n1092, n_n1074, n_n1045, n_n1060, x152x, x151x}, x5894x);
	defparam lut_3012.LUT_SIZE = 7;
	defparam lut_3012.mask = 128'h0707ffff1717ffff7fffffffffffffff;

	lut_sub lut_3019 ({sk[784], n_n78, x55x, n_n95, n_n1145, n_n1146, x33x}, x6334x);
	defparam lut_3019.LUT_SIZE = 7;
	defparam lut_3019.mask = 128'h0707ffff1717ffffc0c0c00080808000;

	lut_sub lut_3024 ({sk[785], x174x, n_n1147, n_n1009, x339x, n_n1013, x6334x}, x5895x);
	defparam lut_3024.LUT_SIZE = 7;
	defparam lut_3024.mask = 128'h0707ffff1717ffffbbffffffbfffffff;

	lut_sub lut_3030 ({sk[786], i_3_, i_1_, i_2_, n_n64, n_n79, n_n87}, x5914x);
	defparam lut_3030.LUT_SIZE = 7;
	defparam lut_3030.mask = 128'h0707ffff1717ffff0000000300050000;

	lut_sub lut_3033 ({sk[787], i_7_, i_8_, i_6_, n_n81, n_n103, x45x}, x5916x);
	defparam lut_3033.LUT_SIZE = 7;
	defparam lut_3033.mask = 128'h0707ffff1717ffff0000030300000055;

	lut_sub lut_3036 ({sk[788], i_7_, i_8_, i_6_, n_n103, n_n84, x21x}, x5917x);
	defparam lut_3036.LUT_SIZE = 7;
	defparam lut_3036.mask = 128'h0707ffff1717ffff0000000000570003;

	lut_sub lut_3039 ({sk[789], i_5_, i_3_, i_4_, n_n58, n_n103, x20x}, x5918x);
	defparam lut_3039.LUT_SIZE = 7;
	defparam lut_3039.mask = 128'h0707ffff1717ffff0000000000035500;

	lut_sub lut_3042 ({sk[790], n_n101, n_n93, x29x, x24x, x5391x, x307x}, x5929x);
	defparam lut_3042.LUT_SIZE = 7;
	defparam lut_3042.mask = 128'h0707ffff1717ffff77777f7f77ff7fff;

	lut_sub lut_3047 ({sk[791], n_n84, x32x, x179x, n_n1160, x92x, x155x}, x5930x);
	defparam lut_3047.LUT_SIZE = 7;
	defparam lut_3047.mask = 128'h0707ffff1717ffff7fff7fff7fffffff;

	lut_sub lut_3053 ({sk[792], x157x, x209x, x210x, x213x}, x5931x);
	defparam lut_3053.LUT_SIZE = 5;
	defparam lut_3053.mask = 32'h0fff7fff;

	lut_sub lut_3058 ({sk[793], i_7_, i_8_, i_6_, x42x, x63x, x86x}, x6382x);
	defparam lut_3058.LUT_SIZE = 7;
	defparam lut_3058.mask = 128'h0707ffff1717ffffccfffff0ffffaaff;

	lut_sub lut_3073 ({sk[794], x321x, x131x, x5068x, x336x, x267x, x6382x}, x5932x);
	defparam lut_3073.LUT_SIZE = 7;
	defparam lut_3073.mask = 128'h0707ffff1717ffffbfbfbfffffffffff;

	lut_sub lut_3079 ({sk[795], n_n101, n_n93, x38x, x82x, x74x, x174x}, x6388x);
	defparam lut_3079.LUT_SIZE = 7;
	defparam lut_3079.mask = 128'h0707ffff1717ffffffaacc88f0a0c080;

	lut_sub lut_3088 ({sk[796], i_5_, i_4_, n_n58, n_n1039, x327x, x280x}, x5951x);
	defparam lut_3088.LUT_SIZE = 7;
	defparam lut_3088.mask = 128'h0707ffff1717ffff5f7f5f5f5f5f5f5f;

	lut_sub lut_3092 ({sk[797], i_7_, i_8_, n_n80, n_n103, x337x, x130x}, x5965x);
	defparam lut_3092.LUT_SIZE = 7;
	defparam lut_3092.mask = 128'h0707ffff1717ffff0537003300330033;

	lut_sub lut_3095 ({sk[798], i_7_, i_8_, n_n81, n_n103, n_n100, n_n76}, x5966x);
	defparam lut_3095.LUT_SIZE = 7;
	defparam lut_3095.mask = 128'h0707ffff1717ffff000f000000001111;

	lut_sub lut_3098 ({sk[799], i_7_, i_8_, i_6_, n_n96, n_n85, x19x}, x5967x);
	defparam lut_3098.LUT_SIZE = 7;
	defparam lut_3098.mask = 128'h0707ffff1717ffff0000035700550000;

	lut_sub lut_3102 ({sk[800], i_7_, i_8_, i_6_, x76x, n_n103, n_n71}, x5968x);
	defparam lut_3102.LUT_SIZE = 7;
	defparam lut_3102.mask = 128'h0707ffff1717ffff00000f0000001111;

	lut_sub lut_3105 ({sk[801], i_7_, i_8_, i_6_, n_n100, n_n102, n_n90}, x5969x);
	defparam lut_3105.LUT_SIZE = 7;
	defparam lut_3105.mask = 128'h0707ffff1717ffff0000110000030000;

	lut_sub lut_3108 ({sk[802], i_5_, i_3_, i_4_, n_n91, n_n83, x37x}, x5970x);
	defparam lut_3108.LUT_SIZE = 7;
	defparam lut_3108.mask = 128'h0707ffff1717ffff0000000000000355;

	lut_sub lut_3111 ({sk[803], n_n58, n_n78, n_n84, x239x, n_n90, x323x}, x6363x);
	defparam lut_3111.LUT_SIZE = 7;
	defparam lut_3111.mask = 128'h0707ffff1717ffffaaaaaa88a0a0a080;

	lut_sub lut_3118 ({sk[804], i_7_, i_8_, i_6_, n_n85, x325x, x24x}, x6364x);
	defparam lut_3118.LUT_SIZE = 7;
	defparam lut_3118.mask = 128'h0707ffff1717ffffaafffffffcaaffff;

	lut_sub lut_3127 ({sk[805], i_7_, i_8_, i_6_, i_4_, x27x, x242x}, x5996x);
	defparam lut_3127.LUT_SIZE = 7;
	defparam lut_3127.mask = 128'h0707ffff1717ffff0000003350000000;

	lut_sub lut_3130 ({sk[806], i_7_, i_8_, i_6_, x21x, x33x}, x6005x);
	defparam lut_3130.LUT_SIZE = 6;
	defparam lut_3130.mask = 64'h3333ffff03030005;

	lut_sub lut_3133 ({sk[807], i_7_, i_8_, n_n102, n_n85, n_n977, x5338x}, x6007x);
	defparam lut_3133.LUT_SIZE = 7;
	defparam lut_3133.mask = 128'h0707ffff1717ffff33333737333f3333;

	lut_sub lut_3137 ({sk[808], n_n101, n_n91, x29x, x63x, x83x, x22x}, x6015x);
	defparam lut_3137.LUT_SIZE = 7;
	defparam lut_3137.mask = 128'h0707ffff1717ffff00007f7f00ff7fff;

	lut_sub lut_3142 ({sk[809], n_n78, n_n84, n_n941, x237x, n_n1164, x4901x}, x6333x);
	defparam lut_3142.LUT_SIZE = 7;
	defparam lut_3142.mask = 128'h0707ffff1717ffffcc008800c0008000;


endmodule