module ks_seq_qmap_map (sk, i_37_, i_7_, i_5_, i_36_, i_34_, i_35_, i_33_, i_32_, i_31_, i_16_, i_9_, i_40_, i_38_, i_39_, i_11_, i_12_, i_15_, i_24_, i_17_, i_22_, i_2_, i_1_, i_3_, i_4_, i_13_, i_0_, i_10_, i_27_, i_25_, i_26_, i_18_, i_19_, i_30_, i_28_, i_29_, i_21_, i_23_, i_14_, i_20_, i_8_, i_6_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_);

	input i_37_;
	input i_7_;
	input i_5_;
	input i_36_;
	input i_34_;
	input i_35_;
	input i_33_;
	input i_32_;
	input i_31_;
	input i_16_;
	input i_9_;
	input i_40_;
	input i_38_;
	input i_39_;
	input i_11_;
	input i_12_;
	input i_15_;
	input i_24_;
	input i_17_;
	input i_22_;
	input i_2_;
	input i_1_;
	input i_3_;
	input i_4_;
	input i_13_;
	input i_0_;
	input i_10_;
	input i_27_;
	input i_25_;
	input i_26_;
	input i_18_;
	input i_19_;
	input i_30_;
	input i_28_;
	input i_29_;
	input i_21_;
	input i_23_;
	input i_14_;
	input i_20_;
	input i_8_;
	input i_6_;
	output o_0_;
	output o_1_;
	output o_2_;
	output o_3_;
	output o_4_;
	output o_5_;
	output o_6_;
	output o_7_;
	output o_8_;
	output o_9_;
	output o_10_;
	output o_11_;
	output o_12_;
	output o_13_;
	output o_14_;
	output o_15_;
	output o_16_;
	output o_17_;
	output o_18_;
	output o_19_;
	output o_20_;
	output o_21_;
	output o_22_;
	output o_23_;
	output o_24_;
	output o_25_;
	output o_26_;
	output o_27_;
	output o_28_;
	output o_29_;
	output o_30_;
	output o_31_;
	output o_32_;
	output o_33_;
	output o_34_;

	input [127 : 0] sk /* synthesis noprune */;


	wire g159, g207, g230, g287, g328, g421, g439, g440, g441, g453, g458, g459, g184, g469, g519, g526, g554, g565, g597, g613, g616;
	wire g617, g607, g615, g619, g610, g660, g689, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14;
	wire g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35;
	wire g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56;
	wire g57, g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77;
	wire g78, g79, g80, g81, g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98;
	wire g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g692, g111, g112, g113, g114, g115, g116, g117, g118;
	wire g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g136, g137, g138, g139;
	wire g140, g141, g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g747, g158, g160;
	wire g161, g162, g163, g164, g165, g166, g167, g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178, g691, g179, g180;
	wire g181, g182, g183, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195, g196, g197, g198, g199, g200, g201, g202;
	wire g203, g204, g205, g206, g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219, g220, g221, g222, g223, g224;
	wire g225, g226, g227, g228, g229, g231, g232, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242, g243, g244, g245, g246;
	wire g247, g248, g249, g250, g251, g252, g253, g254, g255, g256, g257, g258, g259, g260, g261, g262, g740, g263, g264, g265, g266;
	wire g267, g268, g269, g270, g729, g271, g272, g273, g274, g275, g276, g277, g278, g279, g280, g281, g282, g283, g284, g285, g286;
	wire g288, g289, g290, g291, g292, g293, g294, g295, g296, g297, g298, g299, g300, g301, g302, g303, g304, g305, g306, g307, g308;
	wire g309, g310, g311, g312, g313, g314, g315, g316, g317, g318, g319, g320, g321, g322, g323, g324, g325, g326, g327, g329, g330;
	wire g331, g332, g333, g334, g335, g336, g337, g338, g339, g340, g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351;
	wire g352, g353, g354, g355, g356, g357, g723, g358, g359, g360, g361, g362, g363, g364, g365, g366, g367, g368, g369, g370, g371;
	wire g372, g373, g374, g375, g376, g377, g378, g379, g381, g382, g383, g384, g385, g386, g387, g388, g389, g390, g391, g392, g393;
	wire g394, g395, g396, g397, g398, g399, g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410, g411, g412, g413, g414;
	wire g415, g416, g417, g418, g419, g420, g422, g423, g424, g425, g426, g427, g428, g429, g430, g431, g432, g433, g434, g435, g436;
	wire g437, g438, g442, g443, g444, g445, g446, g447, g449, g450, g451, g452, g454, g455, g457, g460, g461, g462, g463, g464, g465;
	wire g466, g467, g468, g470, g471, g472, g473, g474, g475, g476, g477, g478, g479, g480, g481, g482, g483, g484, g485, g486, g487;
	wire g488, g489, g491, g492, g493, g494, g495, g496, g497, g498, g499, g500, g501, g502, g503, g504, g505, g506, g507, g508, g509;
	wire g510, g511, g512, g513, g514, g515, g516, g517, g518, g520, g521, g522, g523, g524, g525, g712, g527, g528, g529, g530, g531;
	wire g532, g533, g534, g535, g536, g537, g538, g539, g540, g541, g542, g543, g544, g545, g546, g547, g548, g549, g550, g551, g552;
	wire g553, g555, g556, g557, g558, g559, g560, g561, g562, g563, g564, g566, g567, g568, g569, g570, g571, g572, g573, g574, g576;
	wire g577, g578, g704, g579, g580, g581, g582, g583, g584, g585, g586, g587, g588, g589, g590, g591, g592, g593, g594, g595, g693;
	wire g596, g598, g599, g600, g601, g602, g603, g604, g605, g606, g608, g609, g611, g612, g614, g618, g620, g621, g622, g623, g624;
	wire g626, g627, g629, g630, g631, g632, g633, g634, g635, g636, g637, g638, g639, g640, g641, g642, g643, g644, g645, g646, g647;
	wire g648, g649, g650, g651, g652, g653, g654, g655, g656, g657, g658, g659, g661, g662, g663, g664, g665, g666, g667, g668, g669;
	wire g670, g671, g672, g673, g674, g675, g676, g677, g678, g679, g680, g681, g682, g683, g684, g685, g686, g687, g688, g690, g694;
	wire g695, g696, g699, g697, g698, g702, g703, g700, g701, g705, g706, g707, g709, g708, g711, g710, g713, g714, g715, g717, g716;
	wire g720, g718, g719, g721, g722, g724, g725, g726, g727, g728, g730, g731, g732, g735, g733, g734, g737, g738, g736, g739, g741;
	wire g742, g743, g744, g745, g746, g748, g749, g750, g753, g751, g752, g756, g757, g754, g755, g758, g759;

	assign o_0_ = (((sk[0]) & (!g159)));
	assign o_1_ = (((sk[1]) & (!g207)));
	assign o_2_ = (((sk[2]) & (!g230)));
	assign o_3_ = (((sk[3]) & (!g287)));
	assign o_4_ = (((sk[4]) & (!g328)));
	assign o_6_ = (((sk[5]) & (!g421)));
	assign o_7_ = (((sk[6]) & (!g439)));
	assign o_8_ = (((sk[7]) & (!g440)));
	assign o_9_ = (((sk[8]) & (!g441)));
	assign o_11_ = (((sk[9]) & (!g453)));
	assign o_13_ = (((sk[10]) & (!g458)));
	assign o_14_ = (((sk[11]) & (!g459)));
	assign o_15_ = (((sk[12]) & (!g184)));
	assign o_16_ = (((sk[13]) & (!g469)));
	assign o_18_ = (((sk[14]) & (!g519)));
	assign o_19_ = (((sk[15]) & (!g526)));
	assign o_20_ = (((sk[16]) & (!g554)));
	assign o_21_ = (((sk[17]) & (!g565)));
	assign o_23_ = (((sk[18]) & (!g597)));
	assign o_24_ = (((sk[19]) & (!g613)));
	assign o_25_ = (((sk[20]) & (!g616)));
	assign o_26_ = (((sk[21]) & (!g617)));
	assign o_27_ = (((sk[22]) & (!g607)));
	assign o_28_ = (((sk[23]) & (!g615)));
	assign o_29_ = (((sk[24]) & (!g619)));
	assign o_32_ = (((sk[25]) & (!g610)));
	assign o_33_ = (((sk[26]) & (!g660)));
	assign o_34_ = (((sk[27]) & (!g689)));
	assign g1 = (((i_7_) & (!sk[28]) & (!i_5_)) + ((!i_7_) & (sk[28]) & (i_5_)));
	assign g2 = (((i_36_) & (!sk[29]) & (!i_34_) & (!i_35_)) + ((!i_36_) & (!sk[29]) & (i_34_) & (!i_35_)) + ((!i_36_) & (sk[29]) & (!i_34_) & (!i_35_)));
	assign g3 = (((!sk[30]) & (i_33_) & (!i_32_) & (!i_31_)) + ((!sk[30]) & (!i_33_) & (i_32_) & (!i_31_)) + ((!sk[30]) & (i_33_) & (!i_32_) & (!i_31_)));
	assign g4 = (((!g1) & (!sk[31]) & (g2) & (!g3) & (!i_16_) & (!i_9_)) + ((g1) & (!sk[31]) & (!g2) & (g3) & (!i_16_) & (!i_9_)) + ((!g1) & (!sk[31]) & (!g2) & (!g3) & (i_16_) & (i_9_)) + ((!g1) & (!sk[31]) & (g2) & (g3) & (!i_16_) & (!i_9_)));
	assign g5 = (((!sk[32]) & (i_34_) & (!i_35_)) + ((sk[32]) & (!i_34_) & (i_35_)));
	assign g6 = (((!sk[33]) & (i_7_) & (!i_33_) & (!i_32_)) + ((!sk[33]) & (!i_7_) & (i_33_) & (!i_32_)) + ((!sk[33]) & (!i_7_) & (i_33_) & (!i_32_)));
	assign g7 = (((!sk[34]) & (i_36_) & (!g5) & (!g6)) + ((!sk[34]) & (!i_36_) & (g5) & (!g6)) + ((!sk[34]) & (i_36_) & (g5) & (g6)));
	assign g8 = (((i_37_) & (!i_38_) & (!sk[35]) & (!i_39_)) + ((!i_37_) & (i_38_) & (!sk[35]) & (!i_39_)) + ((i_37_) & (!i_38_) & (!sk[35]) & (i_39_)));
	assign g9 = (((i_40_) & (!sk[36]) & (!g7) & (!g8)) + ((!i_40_) & (!sk[36]) & (g7) & (!g8)) + ((!i_40_) & (!sk[36]) & (g7) & (g8)));
	assign g10 = (((!sk[37]) & (!i_33_) & (i_34_) & (!i_35_)) + ((!sk[37]) & (i_33_) & (!i_34_) & (!i_35_)) + ((sk[37]) & (!i_33_) & (!i_34_) & (!i_35_)) + ((!sk[37]) & (i_33_) & (!i_34_) & (!i_35_)));
	assign g11 = (((i_32_) & (!sk[38]) & (!i_15_)) + ((!i_32_) & (sk[38]) & (i_15_)));
	assign g12 = (((g10) & (!sk[39]) & (!g11) & (!i_24_)) + ((!g10) & (!sk[39]) & (g11) & (!i_24_)) + ((!g10) & (!sk[39]) & (g11) & (!i_24_)));
	assign g13 = (((!i_36_) & (!sk[40]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((i_36_) & (!sk[40]) & (!i_37_) & (i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (!sk[40]) & (!i_37_) & (!i_38_) & (i_39_) & (i_40_)) + ((!i_36_) & (sk[40]) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (!sk[40]) & (i_37_) & (!i_38_) & (!i_39_) & (i_40_)));
	assign g14 = (((!sk[41]) & (i_38_) & (!i_39_)) + ((sk[41]) & (!i_38_) & (!i_39_)));
	assign g15 = (((i_36_) & (!i_37_) & (!i_38_) & (!sk[42]) & (!i_39_)) + ((!i_36_) & (!i_37_) & (i_38_) & (!sk[42]) & (!i_39_)) + ((!i_36_) & (!i_37_) & (i_38_) & (!sk[42]) & (i_39_)) + ((!i_36_) & (!i_37_) & (!i_38_) & (sk[42]) & (!i_39_)));
	assign g16 = (((!i_36_) & (i_40_) & (!sk[43]) & (!g14) & (!g15)) + ((i_36_) & (!i_40_) & (!sk[43]) & (g14) & (!g15)) + ((!i_36_) & (!i_40_) & (sk[43]) & (!g14) & (!g15)) + ((i_36_) & (!i_40_) & (sk[43]) & (!g14) & (!g15)) + ((!i_36_) & (!i_40_) & (sk[43]) & (!g14) & (!g15)));
	assign g17 = (((!i_11_) & (!g1) & (i_12_) & (g12) & (g13) & (!g16)) + ((i_11_) & (!g1) & (!i_12_) & (g12) & (!g13) & (!g16)));
	assign g18 = (((!sk[45]) & (!i_11_) & (i_12_) & (!i_15_)) + ((!sk[45]) & (!i_11_) & (!i_12_) & (i_15_)) + ((!sk[45]) & (i_11_) & (!i_12_) & (i_15_)) + ((!sk[45]) & (!i_11_) & (i_12_) & (i_15_)));
	assign g19 = (((!sk[46]) & (!i_38_) & (i_40_) & (!g18)) + ((!sk[46]) & (!i_38_) & (!i_40_) & (g18)) + ((!sk[46]) & (i_38_) & (!i_40_) & (g18)));
	assign g20 = (((i_37_) & (!g4) & (!g9) & (!sk[47]) & (!g17) & (!g19)) + ((!i_37_) & (g4) & (!g9) & (!sk[47]) & (!g17) & (!g19)) + ((i_37_) & (!g4) & (!g9) & (!sk[47]) & (!g17) & (!g19)) + ((!i_37_) & (!g4) & (g9) & (!sk[47]) & (!g17) & (g19)) + ((!i_37_) & (!g4) & (!g9) & (sk[47]) & (!g17) & (!g19)) + ((!i_37_) & (!g4) & (!g9) & (sk[47]) & (!g17) & (!g19)));
	assign g21 = (((!sk[48]) & (!i_37_) & (i_38_) & (!i_39_)) + ((!sk[48]) & (!i_37_) & (!i_38_) & (i_39_)) + ((sk[48]) & (i_37_) & (!i_38_) & (!i_39_)));
	assign g22 = (((!sk[49]) & (!i_11_) & (i_12_)) + ((sk[49]) & (!i_11_) & (!i_12_)));
	assign g23 = (((!g1) & (!sk[50]) & (g22) & (!i_15_)) + ((!g1) & (!sk[50]) & (!g22) & (i_15_)) + ((!g1) & (!sk[50]) & (!g22) & (i_15_)));
	assign g24 = (((!i_16_) & (!sk[51]) & (i_17_)) + ((!i_16_) & (sk[51]) & (!i_17_)));
	assign g25 = (((!g3) & (g23) & (!sk[52]) & (!g24)) + ((!g3) & (!g23) & (!sk[52]) & (g24)) + ((g3) & (g23) & (!sk[52]) & (g24)));
	assign g26 = (((!sk[53]) & (!i_11_) & (i_15_)) + ((!sk[53]) & (i_11_) & (i_15_)));
	assign g27 = (((!i_36_) & (!sk[54]) & (i_37_) & (!i_38_)) + ((!i_36_) & (!sk[54]) & (!i_37_) & (i_38_)) + ((!i_36_) & (!sk[54]) & (!i_37_) & (i_38_)));
	assign g28 = (((i_39_) & (!sk[55]) & (g27)) + ((!i_39_) & (!sk[55]) & (g27)));
	assign g29 = (((!sk[56]) & (!g1) & (i_12_) & (!g28) & (!g12)) + ((!sk[56]) & (g1) & (!i_12_) & (g28) & (!g12)) + ((!sk[56]) & (!g1) & (i_12_) & (g28) & (g12)));
	assign g30 = (((!sk[57]) & (!i_38_) & (i_40_)) + ((sk[57]) & (!i_38_) & (!i_40_)) + ((!sk[57]) & (i_38_) & (i_40_)));
	assign g31 = (((!g1) & (g2) & (!sk[58]) & (!g3)) + ((!g1) & (!g2) & (!sk[58]) & (g3)) + ((!g1) & (g2) & (!sk[58]) & (g3)));
	assign g32 = (((!i_38_) & (!sk[59]) & (i_39_) & (!i_17_)) + ((!i_38_) & (!sk[59]) & (!i_39_) & (i_17_)) + ((i_38_) & (!sk[59]) & (i_39_) & (!i_17_)));
	assign g33 = (((g30) & (!g31) & (!sk[60]) & (!i_9_) & (!g4) & (!g32)) + ((!g30) & (g31) & (!sk[60]) & (!i_9_) & (!g4) & (!g32)) + ((!g30) & (!g31) & (sk[60]) & (!i_9_) & (g4) & (!g32)) + ((!g30) & (!g31) & (!sk[60]) & (i_9_) & (!g4) & (g32)) + ((!g30) & (g31) & (!sk[60]) & (!i_9_) & (!g4) & (g32)));
	assign g34 = (((!g1) & (!sk[61]) & (i_9_)) + ((!g1) & (sk[61]) & (!i_9_)));
	assign g35 = (((!g2) & (g21) & (!sk[62]) & (!g18)) + ((!g2) & (!g21) & (!sk[62]) & (g18)) + ((g2) & (g21) & (!sk[62]) & (g18)));
	assign g36 = (((!sk[63]) & (g3) & (!i_16_) & (!i_17_) & (!g34) & (!g35)) + ((!sk[63]) & (!g3) & (i_16_) & (!i_17_) & (!g34) & (!g35)) + ((!sk[63]) & (!g3) & (!i_16_) & (i_17_) & (!g34) & (g35)) + ((!sk[63]) & (g3) & (!i_16_) & (!i_17_) & (g34) & (g35)) + ((!sk[63]) & (g3) & (!i_16_) & (!i_17_) & (g34) & (g35)));
	assign g37 = (((!sk[64]) & (!i_12_) & (i_15_)) + ((!sk[64]) & (i_12_) & (i_15_)));
	assign g38 = (((!i_37_) & (!i_39_) & (!g30) & (!g26) & (g4) & (g37)) + ((!i_37_) & (i_39_) & (!g30) & (g26) & (g4) & (!g37)) + ((!i_37_) & (i_39_) & (!g30) & (!g26) & (g4) & (g37)));
	assign g39 = (((!i_37_) & (!sk[66]) & (i_38_) & (!i_39_) & (!i_40_)) + ((i_37_) & (!sk[66]) & (!i_38_) & (i_39_) & (!i_40_)) + ((i_37_) & (!sk[66]) & (i_38_) & (i_39_) & (!i_40_)) + ((!i_37_) & (!sk[66]) & (i_38_) & (i_39_) & (!i_40_)));
	assign g40 = (((g31) & (!i_9_) & (!g32) & (!g37) & (!sk[67]) & (!g39)) + ((!g31) & (i_9_) & (!g32) & (!g37) & (!sk[67]) & (!g39)) + ((g31) & (!i_9_) & (!g32) & (!g37) & (!sk[67]) & (g39)) + ((!g31) & (!i_9_) & (g32) & (!g37) & (!sk[67]) & (g39)) + ((g31) & (!i_9_) & (g32) & (g37) & (!sk[67]) & (!g39)));
	assign g41 = (((!g26) & (!g29) & (!g33) & (!g36) & (!g38) & (!g40)) + ((!g26) & (!g29) & (!g33) & (!g36) & (!g38) & (!g40)));
	assign g42 = (((!sk[69]) & (!i_22_) & (g10) & (!g11)) + ((!sk[69]) & (!i_22_) & (!g10) & (g11)) + ((!sk[69]) & (!i_22_) & (!g10) & (g11)));
	assign g43 = (((!g1) & (!sk[70]) & (g22)) + ((!g1) & (sk[70]) & (!g22)));
	assign g44 = (((g42) & (!sk[71]) & (g43)) + ((!g42) & (!sk[71]) & (g43)));
	assign g45 = (((!i_36_) & (!sk[72]) & (i_37_) & (!i_38_)) + ((!i_36_) & (!sk[72]) & (!i_37_) & (i_38_)) + ((!i_36_) & (!sk[72]) & (i_37_) & (!i_38_)));
	assign g46 = (((!i_39_) & (!sk[73]) & (g45)) + ((!i_39_) & (!sk[73]) & (g45)));
	assign g47 = (((!i_2_) & (i_1_) & (!sk[74]) & (!i_3_) & (!i_4_)) + ((i_2_) & (!i_1_) & (!sk[74]) & (i_3_) & (!i_4_)) + ((!i_2_) & (!i_1_) & (sk[74]) & (!i_3_) & (!i_4_)));
	assign g48 = (((!sk[75]) & (!i_7_) & (i_32_)) + ((sk[75]) & (!i_7_) & (!i_32_)));
	assign g49 = (((!sk[76]) & (!i_33_) & (!i_34_) & (i_35_)) + ((!sk[76]) & (!i_33_) & (i_34_) & (!i_35_)) + ((sk[76]) & (!i_33_) & (!i_34_) & (!i_35_)) + ((!sk[76]) & (!i_33_) & (i_34_) & (!i_35_)));
	assign g50 = (((!sk[77]) & (g28) & (!g46) & (!g47) & (!g48) & (!g49)) + ((!sk[77]) & (!g28) & (g46) & (!g47) & (!g48) & (!g49)) + ((!sk[77]) & (!g28) & (!g46) & (g47) & (!g48) & (g49)) + ((!sk[77]) & (g28) & (!g46) & (!g47) & (g48) & (!g49)) + ((!sk[77]) & (!g28) & (g46) & (!g47) & (g48) & (!g49)));
	assign g51 = (((!sk[78]) & (!i_36_) & (i_35_)) + ((sk[78]) & (!i_36_) & (!i_35_)));
	assign g52 = (((i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (!sk[79]) & (!g51)) + ((!i_37_) & (i_38_) & (!i_39_) & (!i_40_) & (!sk[79]) & (!g51)) + ((!i_37_) & (!i_38_) & (i_39_) & (!i_40_) & (!sk[79]) & (g51)) + ((i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (!sk[79]) & (g51)) + ((!i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (sk[79]) & (g51)));
	assign g53 = (((!i_33_) & (i_34_) & (!i_32_) & (!sk[80]) & (!i_31_)) + ((i_33_) & (!i_34_) & (i_32_) & (!sk[80]) & (!i_31_)) + ((i_33_) & (!i_34_) & (!i_32_) & (sk[80]) & (!i_31_)));
	assign g54 = (((!i_7_) & (i_11_) & (!sk[81]) & (!i_5_) & (!i_12_)) + ((i_7_) & (!i_11_) & (!sk[81]) & (i_5_) & (!i_12_)) + ((!i_7_) & (!i_11_) & (sk[81]) & (!i_5_) & (!i_12_)));
	assign g55 = (((!sk[82]) & (g53) & (!g54) & (!i_13_)) + ((!sk[82]) & (!g53) & (!g54) & (i_13_)) + ((!sk[82]) & (g53) & (g54) & (i_13_)));
	assign g56 = (((i_33_) & (!sk[83]) & (!i_34_) & (!i_35_)) + ((!i_33_) & (!sk[83]) & (!i_34_) & (i_35_)) + ((i_33_) & (!sk[83]) & (!i_34_) & (!i_35_)));
	assign g57 = (((i_7_) & (!i_5_) & (!i_13_) & (!sk[84]) & (!i_15_)) + ((!i_7_) & (i_5_) & (!i_13_) & (!sk[84]) & (!i_15_)) + ((!i_7_) & (!i_5_) & (i_13_) & (sk[84]) & (!i_15_)));
	assign g58 = (((g56) & (!i_32_) & (!sk[85]) & (!i_31_) & (!g57)) + ((!g56) & (i_32_) & (!sk[85]) & (!i_31_) & (!g57)) + ((g56) & (!i_32_) & (!sk[85]) & (!i_31_) & (g57)));
	assign g59 = (((!sk[86]) & (i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!sk[86]) & (!i_36_) & (!i_37_) & (i_38_) & (!i_39_) & (!i_40_)) + ((sk[86]) & (!i_36_) & (!i_37_) & (!i_38_) & (i_39_) & (!i_40_)) + ((sk[86]) & (!i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (i_40_)) + ((sk[86]) & (!i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_)));
	assign g60 = (((!sk[87]) & (g52) & (!g55) & (!g58) & (!g59)) + ((!sk[87]) & (!g52) & (g55) & (!g58) & (!g59)) + ((!sk[87]) & (g52) & (g55) & (!g58) & (!g59)) + ((sk[87]) & (!g52) & (!g55) & (g58) & (g59)));
	assign g61 = (((i_37_) & (!sk[88]) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_37_) & (!sk[88]) & (i_38_) & (!i_39_) & (!i_40_)) + ((!i_37_) & (!sk[88]) & (i_38_) & (i_39_) & (!i_40_)));
	assign g62 = (((!i_11_) & (!g1) & (!i_12_) & (!i_15_) & (g31) & (g61)) + ((!i_11_) & (!g1) & (!i_12_) & (!i_15_) & (g31) & (g61)) + ((!i_11_) & (!g1) & (!i_12_) & (!i_15_) & (g31) & (g61)));
	assign g63 = (((g28) & (!g44) & (!g50) & (!g60) & (!sk[90]) & (!g62)) + ((!g28) & (!g44) & (g50) & (!g60) & (!sk[90]) & (!g62)) + ((!g28) & (!g44) & (!g50) & (!g60) & (sk[90]) & (!g62)) + ((!g28) & (!g44) & (!g50) & (!g60) & (sk[90]) & (!g62)));
	assign g64 = (((g2) & (!g21) & (!g25) & (!g41) & (!sk[91]) & (!g63)) + ((!g2) & (g21) & (!g25) & (!g41) & (!sk[91]) & (!g63)) + ((!g2) & (!g21) & (!g25) & (g41) & (sk[91]) & (g63)) + ((!g2) & (!g21) & (!g25) & (g41) & (sk[91]) & (g63)) + ((!g2) & (!g21) & (!g25) & (g41) & (sk[91]) & (g63)));
	assign g65 = (((!i_33_) & (!sk[92]) & (i_34_) & (!i_32_)) + ((i_33_) & (!sk[92]) & (!i_34_) & (i_32_)) + ((i_33_) & (sk[92]) & (!i_34_) & (!i_32_)));
	assign g66 = (((!sk[93]) & (!i_36_) & (i_37_) & (!i_35_) & (!g65)) + ((!sk[93]) & (!i_36_) & (!i_37_) & (i_35_) & (!g65)) + ((!sk[93]) & (i_36_) & (i_37_) & (i_35_) & (g65)));
	assign g67 = (((!i_3_) & (!sk[94]) & (i_4_)) + ((!i_3_) & (!sk[94]) & (i_4_)));
	assign g68 = (((i_7_) & (!i_2_) & (!i_1_) & (!sk[95]) & (!i_0_) & (!g67)) + ((!i_7_) & (i_2_) & (!i_1_) & (!sk[95]) & (!i_0_) & (!g67)) + ((!i_7_) & (i_2_) & (!i_1_) & (!sk[95]) & (i_0_) & (!g67)) + ((!i_7_) & (!i_2_) & (!i_1_) & (sk[95]) & (i_0_) & (!g67)) + ((!i_7_) & (!i_2_) & (!i_1_) & (sk[95]) & (i_0_) & (!g67)));
	assign g69 = (((!i_38_) & (!sk[96]) & (i_40_)) + ((!i_38_) & (sk[96]) & (!i_40_)));
	assign g70 = (((!sk[97]) & (!i_7_) & (g65)) + ((!sk[97]) & (!i_7_) & (g65)));
	assign g71 = (((!i_36_) & (i_37_) & (!sk[98]) & (!i_35_)) + ((i_36_) & (!i_37_) & (!sk[98]) & (i_35_)) + ((i_36_) & (!i_37_) & (sk[98]) & (!i_35_)));
	assign g72 = (((!g70) & (!sk[99]) & (i_10_) & (!i_27_) & (!g71)) + ((!g70) & (!sk[99]) & (!i_10_) & (i_27_) & (!g71)) + ((g70) & (!sk[99]) & (i_10_) & (i_27_) & (g71)));
	assign g73 = (((!sk[100]) & (!i_39_) & (i_40_)) + ((sk[100]) & (!i_39_) & (!i_40_)));
	assign g74 = (((!i_38_) & (g72) & (!sk[101]) & (!g73)) + ((i_38_) & (g72) & (!sk[101]) & (g73)) + ((i_38_) & (!g72) & (!sk[101]) & (g73)));
	assign g75 = (((!i_1_) & (!sk[102]) & (i_3_) & (!i_4_)) + ((i_1_) & (!sk[102]) & (!i_3_) & (i_4_)) + ((!i_1_) & (sk[102]) & (!i_3_) & (!i_4_)));
	assign g76 = (((!sk[103]) & (!i_39_) & (i_40_)) + ((!sk[103]) & (!i_39_) & (i_40_)));
	assign g77 = (((!sk[104]) & (!i_38_) & (g76)) + ((!sk[104]) & (i_38_) & (g76)));
	assign g78 = (((!i_36_) & (!sk[105]) & (i_35_)) + ((i_36_) & (sk[105]) & (!i_35_)));
	assign g79 = (((!i_38_) & (!sk[106]) & (i_39_) & (!i_40_)) + ((i_38_) & (!sk[106]) & (!i_39_) & (i_40_)) + ((i_38_) & (!sk[106]) & (i_39_) & (i_40_)));
	assign g80 = (((!i_37_) & (g77) & (!g78) & (!sk[107]) & (!g79)) + ((!i_37_) & (!g77) & (g78) & (!sk[107]) & (!g79)) + ((i_37_) & (g77) & (g78) & (!sk[107]) & (!g79)) + ((!i_37_) & (!g77) & (g78) & (!sk[107]) & (g79)));
	assign g81 = (((i_2_) & (!g75) & (!g70) & (!sk[108]) & (!i_0_) & (!g80)) + ((!i_2_) & (g75) & (!g70) & (!sk[108]) & (!i_0_) & (!g80)) + ((i_2_) & (!g75) & (g70) & (!sk[108]) & (i_0_) & (g80)) + ((!i_2_) & (!g75) & (g70) & (sk[108]) & (i_0_) & (g80)));
	assign g82 = (((g66) & (!g68) & (!g69) & (!g74) & (!sk[109]) & (!g81)) + ((!g66) & (g68) & (!g69) & (!g74) & (!sk[109]) & (!g81)) + ((!g66) & (!g68) & (!g69) & (!g74) & (sk[109]) & (!g81)) + ((!g66) & (!g68) & (!g69) & (!g74) & (sk[109]) & (!g81)) + ((!g66) & (!g68) & (!g69) & (!g74) & (sk[109]) & (!g81)));
	assign g83 = (((!i_36_) & (!sk[110]) & (i_37_) & (!i_35_)) + ((i_36_) & (!sk[110]) & (!i_37_) & (i_35_)) + ((!i_36_) & (!sk[110]) & (i_37_) & (i_35_)));
	assign g84 = (((!sk[111]) & (!i_38_) & (g65) & (!g76) & (!g83)) + ((!sk[111]) & (!i_38_) & (!g65) & (g76) & (!g83)) + ((!sk[111]) & (!i_38_) & (g65) & (g76) & (g83)));
	assign g85 = (((!sk[112]) & (!i_22_) & (g23) & (!i_24_) & (!g84)) + ((!sk[112]) & (!i_22_) & (!g23) & (i_24_) & (!g84)) + ((!sk[112]) & (!i_22_) & (g23) & (i_24_) & (g84)));
	assign g86 = (((i_36_) & (!i_37_) & (!sk[113]) & (!i_38_) & (!g10) & (!g49)) + ((!i_36_) & (i_37_) & (!sk[113]) & (!i_38_) & (!g10) & (!g49)) + ((i_36_) & (i_37_) & (!sk[113]) & (i_38_) & (!g10) & (!g49)) + ((!i_36_) & (!i_37_) & (sk[113]) & (!i_38_) & (!g10) & (!g49)));
	assign g87 = (((!sk[114]) & (!i_2_) & (i_1_) & (!i_3_) & (!i_0_)) + ((!sk[114]) & (!i_2_) & (!i_1_) & (i_3_) & (!i_0_)) + ((sk[114]) & (i_2_) & (!i_1_) & (!i_3_) & (i_0_)));
	assign g88 = (((!i_36_) & (!sk[115]) & (i_37_) & (!i_35_)) + ((i_36_) & (!sk[115]) & (!i_37_) & (i_35_)));
	assign g89 = (((g14) & (!sk[116]) & (!g70) & (!g88) & (!i_25_) & (!i_26_)) + ((!g14) & (!sk[116]) & (g70) & (!g88) & (!i_25_) & (!i_26_)) + ((g14) & (!sk[116]) & (g70) & (g88) & (!i_25_) & (!i_26_)));
	assign g90 = (((!g48) & (!sk[117]) & (g86) & (!g87) & (!g89)) + ((!g48) & (!sk[117]) & (!g86) & (g87) & (!g89)) + ((!g48) & (sk[117]) & (!g86) & (!g87) & (!g89)) + ((!g48) & (sk[117]) & (!g86) & (!g87) & (!g89)) + ((!g48) & (sk[117]) & (!g86) & (!g87) & (!g89)));
	assign g91 = (((g23) & (!g34) & (!g18) & (!i_18_) & (!sk[118]) & (!i_19_)) + ((!g23) & (g34) & (!g18) & (!i_18_) & (!sk[118]) & (!i_19_)) + ((!g23) & (g34) & (g18) & (!i_18_) & (!sk[118]) & (!i_19_)) + ((g23) & (!g34) & (!g18) & (!i_18_) & (!sk[118]) & (!i_19_)));
	assign g92 = (((!i_1_) & (i_4_) & (!sk[119]) & (!i_0_)) + ((i_1_) & (!i_4_) & (!sk[119]) & (i_0_)) + ((!i_1_) & (!i_4_) & (sk[119]) & (i_0_)));
	assign g93 = (((!sk[120]) & (!g92) & (g7)) + ((!sk[120]) & (g92) & (g7)));
	assign g94 = (((!sk[121]) & (!i_36_) & (i_34_) & (!i_35_)) + ((sk[121]) & (!i_36_) & (!i_34_) & (!i_35_)) + ((!sk[121]) & (i_36_) & (!i_34_) & (i_35_)) + ((!sk[121]) & (i_36_) & (i_34_) & (!i_35_)) + ((!sk[121]) & (!i_36_) & (i_34_) & (i_35_)));
	assign g95 = (((!sk[122]) & (!g6) & (g94)) + ((sk[122]) & (g6) & (!g94)));
	assign g96 = (((g92) & (!sk[123]) & (g95)) + ((!g92) & (!sk[123]) & (g95)));
	assign g97 = (((!sk[124]) & (!i_37_) & (i_38_) & (!g93) & (!g96)) + ((!sk[124]) & (!i_37_) & (!i_38_) & (g93) & (!g96)) + ((!sk[124]) & (i_37_) & (i_38_) & (g93) & (!g96)) + ((sk[124]) & (!i_37_) & (!i_38_) & (!g93) & (g96)));
	assign g98 = (((!i_37_) & (!sk[125]) & (i_38_) & (!i_39_)) + ((i_37_) & (!sk[125]) & (!i_38_) & (i_39_)) + ((!i_37_) & (sk[125]) & (!i_38_) & (i_39_)));
	assign g99 = (((!i_40_) & (!sk[126]) & (g95) & (!g77) & (!g98)) + ((!i_40_) & (!sk[126]) & (!g95) & (g77) & (!g98)) + ((!i_40_) & (!sk[126]) & (g95) & (g77) & (!g98)) + ((i_40_) & (!sk[126]) & (g95) & (!g77) & (g98)));
	assign g100 = (((!i_37_) & (!sk[127]) & (i_38_)) + ((!i_37_) & (sk[127]) & (!i_38_)));
	assign g101 = (((i_39_) & (!sk[0]) & (i_40_)) + ((!i_39_) & (!sk[0]) & (i_40_)));
	assign g102 = (((!sk[1]) & (!g56) & (i_32_)) + ((sk[1]) & (g56) & (!i_32_)));
	assign g103 = (((!sk[2]) & (!i_36_) & (g100) & (!g101) & (!g102)) + ((!sk[2]) & (!i_36_) & (!g100) & (g101) & (!g102)) + ((!sk[2]) & (i_36_) & (g100) & (g101) & (g102)));
	assign g104 = (((!sk[3]) & (!i_38_) & (i_39_)) + ((sk[3]) & (i_38_) & (!i_39_)));
	assign g105 = (((!i_36_) & (!sk[4]) & (i_40_) & (!g104)) + ((i_36_) & (!sk[4]) & (!i_40_) & (g104)) + ((!i_36_) & (!sk[4]) & (i_40_) & (g104)));
	assign g106 = (((!i_33_) & (i_35_) & (!sk[5]) & (!i_32_)) + ((i_33_) & (!i_35_) & (!sk[5]) & (i_32_)) + ((i_33_) & (!i_35_) & (sk[5]) & (!i_32_)));
	assign g107 = (((!g1) & (i_30_) & (!i_28_) & (!sk[6]) & (!i_29_)) + ((!g1) & (!i_30_) & (i_28_) & (!sk[6]) & (!i_29_)) + ((!g1) & (i_30_) & (!i_28_) & (!sk[6]) & (i_29_)));
	assign g108 = (((!sk[7]) & (!g1) & (i_30_) & (!i_28_) & (!i_29_)) + ((!sk[7]) & (!g1) & (!i_30_) & (i_28_) & (!i_29_)) + ((!sk[7]) & (!g1) & (!i_30_) & (i_28_) & (!i_29_)));
	assign g109 = (((i_31_) & (!g105) & (!sk[8]) & (!g106) & (!g107) & (!g108)) + ((!i_31_) & (g105) & (!sk[8]) & (!g106) & (!g107) & (!g108)) + ((!i_31_) & (g105) & (!sk[8]) & (g106) & (g107) & (!g108)) + ((!i_31_) & (g105) & (!sk[8]) & (g106) & (!g107) & (g108)));
	assign g110 = (((i_7_) & (!i_11_) & (!sk[9]) & (!g99) & (!g103) & (!g109)) + ((!i_7_) & (i_11_) & (!sk[9]) & (!g99) & (!g103) & (!g109)) + ((i_7_) & (!i_11_) & (!sk[9]) & (!g99) & (!g103) & (!g109)) + ((!i_7_) & (!i_11_) & (sk[9]) & (!g99) & (!g103) & (!g109)) + ((!i_7_) & (!i_11_) & (sk[9]) & (!g99) & (!g103) & (!g109)));
	assign g111 = (((!sk[10]) & (g85) & (!g90) & (!g692) & (!g97) & (!g110)) + ((!sk[10]) & (!g85) & (g90) & (!g692) & (!g97) & (!g110)) + ((!sk[10]) & (!g85) & (g90) & (!g692) & (!g97) & (g110)));
	assign g112 = (((!i_37_) & (i_38_) & (!sk[11]) & (!i_39_)) + ((!i_37_) & (i_38_) & (!sk[11]) & (i_39_)) + ((i_37_) & (!i_38_) & (!sk[11]) & (i_39_)));
	assign g113 = (((i_40_) & (!sk[12]) & (g112)) + ((!i_40_) & (!sk[12]) & (g112)));
	assign g114 = (((!g24) & (g31) & (!g37) & (!sk[13]) & (!g113)) + ((!g24) & (!g31) & (g37) & (!sk[13]) & (!g113)) + ((g24) & (g31) & (g37) & (!sk[13]) & (g113)));
	assign g115 = (((!sk[14]) & (!i_39_) & (i_40_)) + ((sk[14]) & (i_39_) & (!i_40_)));
	assign g116 = (((!sk[15]) & (!i_37_) & (i_38_)) + ((!sk[15]) & (i_37_) & (i_38_)));
	assign g117 = (((i_36_) & (!g10) & (!g48) & (!sk[16]) & (!g116) & (!i_0_)) + ((!i_36_) & (g10) & (!g48) & (!sk[16]) & (!g116) & (!i_0_)) + ((!i_36_) & (!g10) & (g48) & (sk[16]) & (g116) & (i_0_)));
	assign g118 = (((!i_38_) & (!sk[17]) & (g115)) + ((!i_38_) & (!sk[17]) & (g115)));
	assign g119 = (((!i_37_) & (g51) & (!sk[18]) & (!g118)) + ((i_37_) & (g51) & (!sk[18]) & (g118)) + ((i_37_) & (!g51) & (!sk[18]) & (g118)));
	assign g120 = (((!g53) & (g115) & (g117) & (!g107) & (!g108) & (!g119)) + ((g53) & (!g115) & (!g117) & (g107) & (!g108) & (g119)) + ((g53) & (!g115) & (!g117) & (!g107) & (g108) & (g119)));
	assign g121 = (((!i_36_) & (i_34_) & (!sk[20]) & (!i_35_)) + ((i_36_) & (!i_34_) & (!sk[20]) & (i_35_)) + ((!i_36_) & (!i_34_) & (sk[20]) & (i_35_)));
	assign g122 = (((!i_33_) & (!sk[21]) & (i_32_)) + ((!i_33_) & (sk[21]) & (!i_32_)));
	assign g123 = (((g122) & (!sk[22]) & (!i_22_) & (!g23) & (!i_24_) & (!i_21_)) + ((!g122) & (!sk[22]) & (i_22_) & (!g23) & (!i_24_) & (!i_21_)) + ((!g122) & (!sk[22]) & (i_22_) & (g23) & (i_24_) & (i_21_)));
	assign g124 = (((!sk[23]) & (!i_40_) & (g21)) + ((!sk[23]) & (i_40_) & (g21)));
	assign g125 = (((!sk[24]) & (!g122) & (g121)) + ((!sk[24]) & (!g122) & (g121)));
	assign g126 = (((!sk[25]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (!g125)) + ((!sk[25]) & (!i_37_) & (i_38_) & (!i_39_) & (!i_40_) & (!g125)) + ((!sk[25]) & (!i_37_) & (i_38_) & (i_39_) & (!i_40_) & (g125)) + ((sk[25]) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (g125)));
	assign g127 = (((g23) & (!g121) & (!g123) & (!sk[26]) & (!g124) & (!g126)) + ((!g23) & (g121) & (!g123) & (!sk[26]) & (!g124) & (!g126)) + ((g23) & (!g121) & (!g123) & (!sk[26]) & (!g124) & (g126)) + ((!g23) & (g121) & (g123) & (!sk[26]) & (g124) & (!g126)));
	assign g128 = (((!sk[27]) & (!i_32_) & (g54) & (!i_13_) & (!g10)) + ((!sk[27]) & (!i_32_) & (!g54) & (i_13_) & (!g10)) + ((!sk[27]) & (!i_32_) & (g54) & (i_13_) & (!g10)));
	assign g129 = (((!sk[28]) & (!i_36_) & (i_40_) & (!g14)) + ((!sk[28]) & (i_36_) & (!i_40_) & (g14)) + ((!sk[28]) & (!i_36_) & (i_40_) & (g14)));
	assign g130 = (((!g122) & (!sk[29]) & (g94)) + ((!g122) & (sk[29]) & (!g94)));
	assign g131 = (((!i_38_) & (!sk[30]) & (i_39_) & (!i_40_)) + ((i_38_) & (!sk[30]) & (!i_39_) & (i_40_)) + ((!i_38_) & (!sk[30]) & (i_39_) & (i_40_)));
	assign g132 = (((!sk[31]) & (!g130) & (g131)) + ((!sk[31]) & (g130) & (g131)));
	assign g133 = (((!g23) & (g128) & (!sk[32]) & (!g129) & (!g132)) + ((!g23) & (g128) & (!sk[32]) & (g129) & (!g132)) + ((!g23) & (!g128) & (!sk[32]) & (g129) & (!g132)) + ((g23) & (!g128) & (sk[32]) & (!g129) & (g132)));
	assign g134 = (((!sk[33]) & (!i_34_) & (g51) & (!g122)) + ((!sk[33]) & (i_34_) & (!g51) & (g122)) + ((!sk[33]) & (i_34_) & (g51) & (!g122)));
	assign g135 = (((!i_38_) & (!sk[34]) & (g101) & (!g134)) + ((i_38_) & (!sk[34]) & (!g101) & (g134)) + ((!i_38_) & (!sk[34]) & (g101) & (g134)));
	assign g136 = (((!sk[35]) & (!i_36_) & (i_37_) & (!i_35_)) + ((!sk[35]) & (i_36_) & (!i_37_) & (i_35_)) + ((sk[35]) & (!i_36_) & (!i_37_) & (!i_35_)));
	assign g137 = (((!i_38_) & (i_40_) & (!sk[36]) & (!g55) & (!g136)) + ((!i_38_) & (!i_40_) & (!sk[36]) & (g55) & (!g136)) + ((i_38_) & (!i_40_) & (!sk[36]) & (g55) & (g136)));
	assign g138 = (((!g56) & (i_32_) & (!sk[37]) & (!i_31_)) + ((g56) & (!i_32_) & (!sk[37]) & (i_31_)) + ((g56) & (!i_32_) & (sk[37]) & (!i_31_)));
	assign g139 = (((!sk[38]) & (!i_38_) & (g76)) + ((!sk[38]) & (!i_38_) & (g76)));
	assign g140 = (((!i_40_) & (!g27) & (!g138) & (g57) & (g139) & (g125)) + ((!i_40_) & (g27) & (g138) & (g57) & (!g139) & (!g125)));
	assign g141 = (((g1) & (!i_13_) & (!sk[40]) & (!g135) & (!g137) & (!g140)) + ((!g1) & (i_13_) & (!sk[40]) & (!g135) & (!g137) & (!g140)) + ((g1) & (!i_13_) & (!sk[40]) & (!g135) & (!g137) & (!g140)) + ((!g1) & (!i_13_) & (sk[40]) & (!g135) & (!g137) & (!g140)) + ((!g1) & (!i_13_) & (sk[40]) & (!g135) & (!g137) & (!g140)));
	assign g142 = (((g114) & (!sk[41]) & (!g120) & (!g127) & (!g133) & (!g141)) + ((!g114) & (!sk[41]) & (g120) & (!g127) & (!g133) & (!g141)) + ((!g114) & (sk[41]) & (!g120) & (!g127) & (!g133) & (g141)));
	assign g143 = (((!g10) & (!sk[42]) & (g11)) + ((!g10) & (!sk[42]) & (g11)));
	assign g144 = (((g143) & (!sk[43]) & (g43)) + ((!g143) & (!sk[43]) & (g43)));
	assign g145 = (((!i_11_) & (g1) & (!i_12_) & (!sk[44]) & (!g24)) + ((!i_11_) & (!g1) & (i_12_) & (!sk[44]) & (!g24)) + ((i_11_) & (!g1) & (!i_12_) & (sk[44]) & (g24)));
	assign g146 = (((!g56) & (i_31_) & (!g11) & (!sk[45]) & (!g145)) + ((!g56) & (!i_31_) & (g11) & (!sk[45]) & (!g145)) + ((g56) & (!i_31_) & (g11) & (!sk[45]) & (g145)));
	assign g147 = (((!sk[46]) & (i_37_) & (!i_38_) & (!i_39_) & (!g57) & (!g125)) + ((!sk[46]) & (!i_37_) & (i_38_) & (!i_39_) & (!g57) & (!g125)) + ((!sk[46]) & (!i_37_) & (i_38_) & (i_39_) & (g57) & (g125)) + ((sk[46]) & (!i_37_) & (!i_38_) & (!i_39_) & (g57) & (g125)));
	assign g148 = (((!sk[47]) & (!i_34_) & (g6) & (!g78)) + ((!sk[47]) & (i_34_) & (!g6) & (g78)) + ((!sk[47]) & (!i_34_) & (g6) & (g78)));
	assign g149 = (((i_37_) & (!i_38_) & (!sk[48]) & (!i_39_) & (!i_40_) & (!g148)) + ((!i_37_) & (i_38_) & (!sk[48]) & (!i_39_) & (!i_40_) & (!g148)) + ((i_37_) & (i_38_) & (!sk[48]) & (i_39_) & (!i_40_) & (g148)));
	assign g150 = (((!g128) & (!sk[49]) & (g147) & (!g15) & (!g149)) + ((!g128) & (!sk[49]) & (!g147) & (g15) & (!g149)) + ((!g128) & (sk[49]) & (!g147) & (!g15) & (!g149)) + ((!g128) & (!sk[49]) & (!g147) & (g15) & (!g149)));
	assign g151 = (((!i_36_) & (i_37_) & (!sk[50]) & (!i_35_)) + ((i_36_) & (!i_37_) & (!sk[50]) & (i_35_)) + ((!i_36_) & (!i_37_) & (sk[50]) & (i_35_)));
	assign g152 = (((sk[51]) & (!i_38_) & (!i_39_) & (!g65) & (!g151)) + ((!sk[51]) & (!i_38_) & (i_39_) & (!g65) & (!g151)) + ((!sk[51]) & (!i_38_) & (!i_39_) & (g65) & (!g151)) + ((sk[51]) & (!i_38_) & (!i_39_) & (!g65) & (!g151)) + ((!sk[51]) & (!i_38_) & (!i_39_) & (g65) & (!g151)));
	assign g153 = (((!sk[52]) & (!i_22_) & (i_24_) & (!i_21_)) + ((!sk[52]) & (i_22_) & (!i_24_) & (i_21_)) + ((!sk[52]) & (i_22_) & (i_24_) & (!i_21_)));
	assign g154 = (((!sk[53]) & (!g18) & (i_23_) & (!g153)) + ((!sk[53]) & (g18) & (!i_23_) & (g153)));
	assign g155 = (((!g1) & (!sk[54]) & (i_9_)) + ((!g1) & (!sk[54]) & (i_9_)));
	assign g156 = (((g125) & (!i_18_) & (!sk[55]) & (!g124) & (!g155) & (!i_19_)) + ((!g125) & (i_18_) & (!sk[55]) & (!g124) & (!g155) & (!i_19_)) + ((g125) & (i_18_) & (!sk[55]) & (g124) & (g155) & (!i_19_)) + ((g125) & (!i_18_) & (!sk[55]) & (g124) & (g155) & (i_19_)));
	assign g157 = (((!i_32_) & (g10) & (!g45) & (!sk[56]) & (!g76)) + ((!i_32_) & (!g10) & (g45) & (!sk[56]) & (!g76)) + ((!i_32_) & (!g10) & (g45) & (!sk[56]) & (g76)));
	assign g158 = (((!g28) & (!i_21_) & (!g144) & (!g146) & (g150) & (g747)) + ((!g28) & (!i_21_) & (!g144) & (!g146) & (g150) & (g747)) + ((!g28) & (!i_21_) & (!g144) & (!g146) & (g150) & (g747)));
	assign g159 = (((g20) & (g64) & (g82) & (g111) & (g142) & (g158)));
	assign g160 = (((!sk[59]) & (!i_36_) & (g5)) + ((!sk[59]) & (i_36_) & (g5)));
	assign g161 = (((g100) & (!g122) & (!i_25_) & (!i_26_) & (!sk[60]) & (!g160)) + ((!g100) & (g122) & (!i_25_) & (!i_26_) & (!sk[60]) & (!g160)) + ((g100) & (!g122) & (i_25_) & (!i_26_) & (!sk[60]) & (g160)) + ((g100) & (!g122) & (!i_25_) & (i_26_) & (!sk[60]) & (g160)));
	assign g162 = (((!i_33_) & (!sk[61]) & (i_34_)) + ((!i_33_) & (sk[61]) & (!i_34_)));
	assign g163 = (((!i_11_) & (!sk[62]) & (i_36_) & (!i_12_)) + ((i_11_) & (!sk[62]) & (!i_36_) & (i_12_)) + ((!i_11_) & (!sk[62]) & (i_36_) & (i_12_)));
	assign g164 = (((i_40_) & (!g162) & (!i_32_) & (!sk[63]) & (!g98) & (!g163)) + ((!i_40_) & (g162) & (!i_32_) & (!sk[63]) & (!g98) & (!g163)) + ((i_40_) & (!g162) & (!i_32_) & (!sk[63]) & (g98) & (g163)));
	assign g165 = (((g101) & (!sk[64]) & (g27)) + ((!g101) & (!sk[64]) & (g27)));
	assign g166 = (((i_5_) & (!i_16_) & (!i_17_) & (!sk[65]) & (!i_9_) & (!g18)) + ((!i_5_) & (i_16_) & (!i_17_) & (!sk[65]) & (!i_9_) & (!g18)) + ((!i_5_) & (i_16_) & (i_17_) & (!sk[65]) & (!i_9_) & (g18)) + ((!i_5_) & (i_16_) & (!i_17_) & (!sk[65]) & (i_9_) & (g18)) + ((!i_5_) & (!i_16_) & (i_17_) & (sk[65]) & (i_9_) & (g18)));
	assign g167 = (((!g102) & (g165) & (!sk[66]) & (!g166)) + ((g102) & (g165) & (!sk[66]) & (g166)) + ((g102) & (!g165) & (!sk[66]) & (g166)));
	assign g168 = (((!sk[67]) & (!i_37_) & (g51) & (!g14)) + ((!sk[67]) & (i_37_) & (!g51) & (g14)) + ((!sk[67]) & (i_37_) & (g51) & (g14)));
	assign g169 = (((i_5_) & (!sk[68]) & (!i_15_) & (!i_16_) & (!i_17_) & (!i_9_)) + ((!i_5_) & (!sk[68]) & (i_15_) & (!i_16_) & (!i_17_) & (!i_9_)) + ((!i_5_) & (!sk[68]) & (i_15_) & (i_16_) & (i_17_) & (!i_9_)) + ((!i_5_) & (!sk[68]) & (i_15_) & (i_16_) & (!i_17_) & (i_9_)) + ((!i_5_) & (!sk[68]) & (i_15_) & (!i_16_) & (i_17_) & (i_9_)));
	assign g170 = (((!i_12_) & (!sk[69]) & (i_14_) & (!g169)) + ((i_12_) & (!sk[69]) & (!i_14_) & (g169)));
	assign g171 = (((!sk[70]) & (!i_16_) & (i_17_)) + ((!sk[70]) & (i_16_) & (i_17_)));
	assign g172 = (((!sk[71]) & (!i_5_) & (i_13_) & (!i_15_)) + ((!sk[71]) & (i_5_) & (!i_13_) & (i_15_)) + ((sk[71]) & (!i_5_) & (!i_13_) & (!i_15_)));
	assign g173 = (((!i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (i_35_)) + ((!i_36_) & (!i_37_) & (!i_38_) & (i_39_) & (!i_40_) & (!i_35_)) + ((!i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (!i_35_)) + ((!i_36_) & (!i_37_) & (!i_38_) & (i_39_) & (i_40_) & (!i_35_)) + ((!i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (!i_35_)));
	assign g174 = (((!g51) & (i_31_) & (!sk[73]) & (!i_5_) & (!g37)) + ((!g51) & (!i_31_) & (!sk[73]) & (i_5_) & (!g37)) + ((g51) & (i_31_) & (!sk[73]) & (!i_5_) & (!g37)));
	assign g175 = (((!i_38_) & (i_39_) & (!sk[74]) & (!g83) & (!g174)) + ((!i_38_) & (!i_39_) & (!sk[74]) & (g83) & (!g174)) + ((i_38_) & (!i_39_) & (sk[74]) & (!g83) & (!g174)) + ((!i_38_) & (!i_39_) & (sk[74]) & (!g83) & (!g174)) + ((!i_38_) & (!i_39_) & (sk[74]) & (!g83) & (!g174)));
	assign g176 = (((i_36_) & (!i_37_) & (!i_38_) & (i_39_) & (!i_40_) & (i_35_)) + ((!i_36_) & (i_37_) & (!i_38_) & (i_39_) & (i_40_) & (i_35_)) + ((!i_36_) & (!i_37_) & (i_38_) & (!i_39_) & (i_40_) & (i_35_)) + ((i_36_) & (!i_37_) & (!i_38_) & (i_39_) & (!i_40_) & (i_35_)) + ((!i_36_) & (i_37_) & (i_38_) & (!i_39_) & (!i_40_) & (i_35_)) + ((i_36_) & (i_37_) & (i_38_) & (i_39_) & (i_40_) & (!i_35_)));
	assign g177 = (((!sk[76]) & (!g172) & (g173) & (!g175) & (!g176)) + ((!sk[76]) & (!g172) & (!g173) & (g175) & (!g176)) + ((!sk[76]) & (!g172) & (!g173) & (g175) & (!g176)) + ((!sk[76]) & (!g172) & (!g173) & (g175) & (!g176)));
	assign g178 = (((i_34_) & (!g51) & (!sk[77]) & (!g122) & (!g47) & (!g113)) + ((!i_34_) & (g51) & (!sk[77]) & (!g122) & (!g47) & (!g113)) + ((!i_34_) & (!g51) & (sk[77]) & (!g122) & (!g47) & (!g113)) + ((!i_34_) & (g51) & (!sk[77]) & (!g122) & (g47) & (g113)));
	assign g179 = (((i_34_) & (!g168) & (!g170) & (!g691) & (!g177) & (g178)) + ((!i_34_) & (!g168) & (!g170) & (!g691) & (!g177) & (g178)) + ((!i_34_) & (g168) & (g170) & (!g691) & (!g177) & (g178)) + ((!i_34_) & (g168) & (!g170) & (g691) & (!g177) & (g178)));
	assign g180 = (((!sk[79]) & (!g27) & (g106) & (!g73)) + ((!sk[79]) & (g27) & (!g106) & (g73)) + ((!sk[79]) & (g27) & (g106) & (g73)));
	assign g181 = (((!g101) & (!sk[80]) & (g45) & (!g152) & (!g106)) + ((!g101) & (!sk[80]) & (!g45) & (g152) & (!g106)) + ((!g101) & (!sk[80]) & (!g45) & (g152) & (!g106)) + ((!g101) & (!sk[80]) & (!g45) & (g152) & (!g106)));
	assign g182 = (((!g30) & (!sk[81]) & (g65) & (!g83)) + ((g30) & (!sk[81]) & (!g65) & (g83)) + ((!g30) & (!sk[81]) & (g65) & (g83)));
	assign g183 = (((!sk[82]) & (i_36_) & (!i_32_) & (!i_31_) & (!i_5_) & (!g21)) + ((!sk[82]) & (!i_36_) & (i_32_) & (!i_31_) & (!i_5_) & (!g21)) + ((sk[82]) & (!i_36_) & (!i_32_) & (i_31_) & (!i_5_) & (!g21)));
	assign g184 = (((!sk[83]) & (!i_7_) & (i_33_)) + ((sk[83]) & (!i_7_) & (!i_33_)) + ((!sk[83]) & (!i_7_) & (i_33_)));
	assign g185 = (((!g122) & (i_5_) & (!sk[84]) & (!g22) & (!i_13_)) + ((!g122) & (!i_5_) & (!sk[84]) & (g22) & (!i_13_)) + ((!g122) & (!i_5_) & (!sk[84]) & (g22) & (!i_13_)));
	assign g186 = (((!i_37_) & (!sk[85]) & (g51) & (!g131) & (!g185)) + ((!i_37_) & (!sk[85]) & (!g51) & (g131) & (!g185)) + ((i_37_) & (!sk[85]) & (g51) & (g131) & (g185)));
	assign g187 = (((!i_38_) & (i_39_) & (!sk[86]) & (!i_40_)) + ((i_38_) & (!i_39_) & (!sk[86]) & (i_40_)) + ((!i_38_) & (!i_39_) & (sk[86]) & (!i_40_)));
	assign g188 = (((!i_34_) & (!sk[87]) & (g122) & (!g71) & (!g187)) + ((!i_34_) & (!sk[87]) & (!g122) & (g71) & (!g187)) + ((i_34_) & (!sk[87]) & (!g122) & (g71) & (g187)));
	assign g189 = (((!i_38_) & (!sk[88]) & (g136) & (!g73)) + ((i_38_) & (!sk[88]) & (!g136) & (g73)) + ((i_38_) & (!sk[88]) & (g136) & (g73)));
	assign g190 = (((!i_37_) & (!sk[89]) & (i_38_) & (!i_39_) & (!i_40_)) + ((!i_37_) & (!sk[89]) & (!i_38_) & (i_39_) & (!i_40_)) + ((!i_37_) & (!sk[89]) & (!i_38_) & (i_39_) & (!i_40_)) + ((!i_37_) & (!sk[89]) & (!i_38_) & (i_39_) & (i_40_)) + ((i_37_) & (sk[89]) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_37_) & (sk[89]) & (!i_38_) & (!i_39_) & (i_40_)));
	assign g191 = (((g2) & (!g188) & (!sk[90]) & (!g185) & (!g189) & (!g190)) + ((!g2) & (g188) & (!sk[90]) & (!g185) & (!g189) & (!g190)) + ((!g2) & (!g188) & (sk[90]) & (!g185) & (!g189) & (!g190)) + ((!g2) & (!g188) & (sk[90]) & (!g185) & (!g189) & (!g190)) + ((!g2) & (!g188) & (sk[90]) & (!g185) & (!g189) & (!g190)));
	assign g192 = (((!sk[91]) & (g56) & (!g183) & (!g184) & (!g186) & (!g191)) + ((!sk[91]) & (!g56) & (g183) & (!g184) & (!g186) & (!g191)) + ((sk[91]) & (!g56) & (!g183) & (g184) & (!g186) & (g191)) + ((sk[91]) & (!g56) & (!g183) & (g184) & (!g186) & (g191)));
	assign g193 = (((g180) & (!g172) & (!g181) & (!g182) & (!sk[92]) & (!g192)) + ((!g180) & (g172) & (!g181) & (!g182) & (!sk[92]) & (!g192)) + ((!g180) & (!g172) & (!g181) & (!g182) & (sk[92]) & (g192)) + ((!g180) & (!g172) & (g181) & (!g182) & (sk[92]) & (g192)));
	assign g194 = (((!sk[93]) & (!i_31_) & (g122) & (!g2)) + ((!sk[93]) & (i_31_) & (!g122) & (g2)));
	assign g195 = (((!i_16_) & (i_17_) & (!sk[94]) & (!i_9_)) + ((!i_16_) & (!i_17_) & (sk[94]) & (!i_9_)) + ((i_16_) & (!i_17_) & (!sk[94]) & (i_9_)) + ((!i_16_) & (!i_17_) & (sk[94]) & (!i_9_)) + ((!i_16_) & (!i_17_) & (sk[94]) & (!i_9_)));
	assign g196 = (((g194) & (!sk[95]) & (g195)) + ((!g194) & (!sk[95]) & (g195)));
	assign g197 = (((!i_34_) & (!sk[96]) & (g122)) + ((i_34_) & (sk[96]) & (!g122)));
	assign g198 = (((!i_5_) & (!sk[97]) & (g18)) + ((!i_5_) & (!sk[97]) & (g18)));
	assign g199 = (((!sk[98]) & (!i_37_) & (g76)) + ((!sk[98]) & (!i_37_) & (g76)));
	assign g200 = (((!i_24_) & (!g125) & (g197) & (g189) & (!g198) & (!g199)) + ((i_24_) & (g125) & (!g197) & (!g189) & (g198) & (g199)));
	assign g201 = (((!i_11_) & (i_12_) & (!sk[100]) & (!i_14_)) + ((i_11_) & (i_12_) & (!sk[100]) & (i_14_)) + ((i_11_) & (!i_12_) & (!sk[100]) & (i_14_)));
	assign g202 = (((i_15_) & (!i_16_) & (!i_17_) & (!sk[101]) & (!i_9_) & (!g201)) + ((!i_15_) & (i_16_) & (!i_17_) & (!sk[101]) & (!i_9_) & (!g201)) + ((i_15_) & (i_16_) & (i_17_) & (!sk[101]) & (!i_9_) & (g201)) + ((i_15_) & (i_16_) & (!i_17_) & (!sk[101]) & (i_9_) & (g201)) + ((i_15_) & (!i_16_) & (i_17_) & (!sk[101]) & (i_9_) & (g201)));
	assign g203 = (((!g65) & (!sk[102]) & (g136) & (!g79) & (!g202)) + ((!g65) & (!sk[102]) & (!g136) & (g79) & (!g202)) + ((g65) & (!sk[102]) & (g136) & (g79) & (g202)));
	assign g204 = (((!i_5_) & (g22) & (!i_13_) & (!sk[103]) & (!g125)) + ((!i_5_) & (!g22) & (i_13_) & (!sk[103]) & (!g125)) + ((!i_5_) & (g22) & (!i_13_) & (!sk[103]) & (g125)));
	assign g205 = (((!sk[104]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (!g204)) + ((!sk[104]) & (!i_37_) & (i_38_) & (!i_39_) & (!i_40_) & (!g204)) + ((!sk[104]) & (!i_37_) & (i_38_) & (i_39_) & (!i_40_) & (g204)) + ((!sk[104]) & (i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (g204)) + ((sk[104]) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (g204)));
	assign g206 = (((i_5_) & (!g196) & (!g200) & (!g203) & (!sk[105]) & (!g205)) + ((!i_5_) & (g196) & (!g200) & (!g203) & (!sk[105]) & (!g205)) + ((i_5_) & (!g196) & (!g200) & (!g203) & (!sk[105]) & (!g205)) + ((!i_5_) & (!g196) & (!g200) & (!g203) & (sk[105]) & (!g205)));
	assign g207 = (((!g161) & (!g164) & (!g167) & (!g179) & (g193) & (g206)));
	assign g208 = (((!g2) & (!g21) & (!g3) & (!g113) & (g184) & (!g691)) + ((!g2) & (!g21) & (!g3) & (!g113) & (g184) & (!g691)) + ((!g2) & (!g21) & (!g3) & (!g113) & (g184) & (!g691)) + ((!g2) & (!g21) & (!g3) & (!g113) & (g184) & (!g691)));
	assign g209 = (((i_5_) & (!g3) & (!sk[108]) & (!i_30_) & (!i_28_) & (!i_29_)) + ((!i_5_) & (g3) & (!sk[108]) & (!i_30_) & (!i_28_) & (!i_29_)) + ((!i_5_) & (g3) & (!sk[108]) & (!i_30_) & (!i_28_) & (!i_29_)) + ((!i_5_) & (g3) & (!sk[108]) & (!i_30_) & (i_28_) & (i_29_)) + ((!i_5_) & (g3) & (!sk[108]) & (i_30_) & (!i_28_) & (!i_29_)));
	assign g210 = (((!g2) & (g77) & (!g119) & (!sk[109]) & (!g209)) + ((!g2) & (!g77) & (g119) & (!sk[109]) & (!g209)) + ((!g2) & (!g77) & (g119) & (!sk[109]) & (g209)) + ((g2) & (g77) & (!g119) & (!sk[109]) & (g209)));
	assign g211 = (((!g14) & (g65) & (!sk[110]) & (!g83)) + ((g14) & (g65) & (!sk[110]) & (g83)) + ((g14) & (!g65) & (!sk[110]) & (g83)));
	assign g212 = (((i_5_) & (!sk[111]) & (!i_9_) & (!g18) & (!i_18_) & (!i_19_)) + ((!i_5_) & (!sk[111]) & (i_9_) & (!g18) & (!i_18_) & (!i_19_)) + ((!i_5_) & (!sk[111]) & (i_9_) & (g18) & (i_18_) & (!i_19_)) + ((!i_5_) & (!sk[111]) & (i_9_) & (g18) & (!i_18_) & (i_19_)) + ((!i_5_) & (sk[111]) & (!i_9_) & (g18) & (i_18_) & (i_19_)));
	assign g213 = (((!i_23_) & (g153) & (!sk[112]) & (!g212)) + ((i_23_) & (g153) & (!sk[112]) & (g212)) + ((i_23_) & (!g153) & (!sk[112]) & (g212)));
	assign g214 = (((!sk[113]) & (!i_34_) & (g122) & (!g78)) + ((!sk[113]) & (i_34_) & (!g122) & (g78)) + ((sk[113]) & (!i_34_) & (!g122) & (g78)));
	assign g215 = (((!i_37_) & (!sk[114]) & (g104)) + ((!i_37_) & (!sk[114]) & (g104)));
	assign g216 = (((!i_36_) & (i_37_) & (!sk[115]) & (!i_38_)) + ((i_36_) & (!i_37_) & (!sk[115]) & (i_38_)));
	assign g217 = (((!sk[116]) & (!g65) & (g76) & (!g216)) + ((!sk[116]) & (g65) & (!g76) & (g216)) + ((!sk[116]) & (g65) & (g76) & (g216)));
	assign g218 = (((!sk[117]) & (i_10_) & (!i_27_) & (!g214) & (!g215) & (!g217)) + ((!sk[117]) & (!i_10_) & (i_27_) & (!g214) & (!g215) & (!g217)) + ((!sk[117]) & (i_10_) & (i_27_) & (!g214) & (!g215) & (!g217)) + ((sk[117]) & (!i_10_) & (!i_27_) & (!g214) & (!g215) & (!g217)) + ((sk[117]) & (!i_10_) & (!i_27_) & (!g214) & (!g215) & (!g217)));
	assign g219 = (((!sk[118]) & (!i_37_) & (g51) & (!g197)) + ((!sk[118]) & (i_37_) & (!g51) & (g197)) + ((!sk[118]) & (i_37_) & (g51) & (g197)));
	assign g220 = (((!g112) & (!sk[119]) & (g124)) + ((!g112) & (sk[119]) & (!g124)));
	assign g221 = (((!sk[120]) & (g47) & (!g130) & (!g118) & (!g219) & (!g220)) + ((!sk[120]) & (!g47) & (g130) & (!g118) & (!g219) & (!g220)) + ((sk[120]) & (!g47) & (!g130) & (g118) & (g219) & (!g220)) + ((!sk[120]) & (g47) & (g130) & (!g118) & (!g219) & (!g220)));
	assign g222 = (((!i_5_) & (!sk[121]) & (i_9_) & (!g18) & (!i_18_)) + ((!i_5_) & (!sk[121]) & (!i_9_) & (g18) & (!i_18_)) + ((!i_5_) & (!sk[121]) & (i_9_) & (g18) & (!i_18_)) + ((!i_5_) & (!sk[121]) & (!i_9_) & (g18) & (i_18_)));
	assign g223 = (((!g125) & (!g153) & (!g79) & (g204) & (g199) & (!g222)) + ((g125) & (g153) & (g79) & (!g204) & (!g199) & (g222)));
	assign g224 = (((g211) & (!sk[123]) & (!g213) & (!g218) & (!g221) & (!g223)) + ((!g211) & (!sk[123]) & (g213) & (!g218) & (!g221) & (!g223)) + ((!g211) & (sk[123]) & (!g213) & (g218) & (!g221) & (!g223)) + ((!g211) & (sk[123]) & (!g213) & (g218) & (!g221) & (!g223)));
	assign g225 = (((!i_37_) & (!sk[124]) & (g14)) + ((!i_37_) & (!sk[124]) & (g14)));
	assign g226 = (((!g122) & (!sk[125]) & (g160) & (!g225)) + ((g122) & (!sk[125]) & (!g160) & (g225)) + ((!g122) & (!sk[125]) & (g160) & (g225)));
	assign g227 = (((!i_36_) & (!i_37_) & (i_38_) & (!i_39_) & (i_40_) & (i_35_)) + ((i_36_) & (i_37_) & (!i_38_) & (i_39_) & (!i_40_) & (!i_35_)) + ((i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (!i_35_)) + ((!i_36_) & (i_37_) & (i_38_) & (i_39_) & (i_40_) & (i_35_)) + ((i_36_) & (!i_37_) & (i_38_) & (i_39_) & (!i_40_) & (i_35_)) + ((!i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (i_35_)));
	assign g228 = (((!sk[127]) & (!g76) & (g151) & (!g172) & (!g227)) + ((!sk[127]) & (!g76) & (!g151) & (g172) & (!g227)) + ((sk[127]) & (!g76) & (!g151) & (!g172) & (!g227)) + ((sk[127]) & (!g76) & (!g151) & (!g172) & (!g227)) + ((sk[127]) & (!g76) & (!g151) & (!g172) & (!g227)));
	assign g229 = (((g65) & (!i_25_) & (!sk[0]) & (!i_26_) & (!g226) & (!g228)) + ((!g65) & (i_25_) & (!sk[0]) & (!i_26_) & (!g226) & (!g228)) + ((!g65) & (!i_25_) & (sk[0]) & (!i_26_) & (!g226) & (!g228)) + ((!g65) & (!i_25_) & (sk[0]) & (!i_26_) & (!g226) & (!g228)) + ((!g65) & (!i_25_) & (sk[0]) & (!i_26_) & (!g226) & (g228)) + ((!g65) & (!i_25_) & (sk[0]) & (!i_26_) & (!g226) & (g228)));
	assign g230 = (((g200) & (!sk[1]) & (!g208) & (!g210) & (!g224) & (!g229)) + ((!g200) & (!sk[1]) & (g208) & (!g210) & (!g224) & (!g229)) + ((!g200) & (!sk[1]) & (g208) & (!g210) & (g224) & (g229)));
	assign g231 = (((!i_22_) & (g112) & (!g125) & (!sk[2]) & (!g198)) + ((!i_22_) & (!g112) & (g125) & (!sk[2]) & (!g198)) + ((!i_22_) & (g112) & (g125) & (!sk[2]) & (g198)));
	assign g232 = (((!sk[3]) & (!i_5_) & (i_9_)) + ((sk[3]) & (!i_5_) & (!i_9_)));
	assign g233 = (((!i_11_) & (!sk[4]) & (i_38_) & (!i_39_) & (!g232)) + ((!i_11_) & (!sk[4]) & (!i_38_) & (i_39_) & (!g232)) + ((i_11_) & (!sk[4]) & (!i_38_) & (i_39_) & (g232)));
	assign g234 = (((i_36_) & (i_37_) & (!sk[5]) & (!i_38_) & (!i_39_)) + ((!i_36_) & (i_37_) & (!sk[5]) & (!i_38_) & (!i_39_)) + ((!i_36_) & (!i_37_) & (!sk[5]) & (i_38_) & (!i_39_)) + ((i_36_) & (!i_37_) & (!sk[5]) & (i_38_) & (i_39_)));
	assign g235 = (((i_40_) & (!sk[6]) & (!i_32_) & (!g47) & (!i_0_) & (!g234)) + ((!i_40_) & (!sk[6]) & (i_32_) & (!g47) & (!i_0_) & (!g234)) + ((i_40_) & (!sk[6]) & (!i_32_) & (!g47) & (i_0_) & (g234)));
	assign g236 = (((i_36_) & (!g11) & (!i_16_) & (!g233) & (!sk[7]) & (!g235)) + ((!i_36_) & (g11) & (!i_16_) & (!g233) & (!sk[7]) & (!g235)) + ((i_36_) & (!g11) & (!i_16_) & (!g233) & (!sk[7]) & (!g235)) + ((!i_36_) & (!g11) & (!i_16_) & (!g233) & (sk[7]) & (!g235)) + ((!i_36_) & (!g11) & (i_16_) & (!g233) & (sk[7]) & (!g235)) + ((!i_36_) & (!g11) & (!i_16_) & (!g233) & (sk[7]) & (!g235)));
	assign g237 = (((!sk[8]) & (i_11_) & (!i_36_) & (!g30) & (!i_12_) & (!g232)) + ((!sk[8]) & (!i_11_) & (i_36_) & (!g30) & (!i_12_) & (!g232)) + ((sk[8]) & (!i_11_) & (!i_36_) & (!g30) & (i_12_) & (g232)) + ((!sk[8]) & (i_11_) & (!i_36_) & (!g30) & (!i_12_) & (g232)));
	assign g238 = (((i_39_) & (!g30) & (!g22) & (!g45) & (!sk[9]) & (!g232)) + ((!i_39_) & (g30) & (!g22) & (!g45) & (!sk[9]) & (!g232)) + ((!i_39_) & (g30) & (!g22) & (!g45) & (!sk[9]) & (!g232)) + ((!i_39_) & (!g30) & (g22) & (!g45) & (sk[9]) & (!g232)) + ((!i_39_) & (!g30) & (!g22) & (!g45) & (sk[9]) & (!g232)));
	assign g239 = (((i_36_) & (!g11) & (!i_16_) & (!sk[10]) & (!g237) & (!g238)) + ((!i_36_) & (g11) & (!i_16_) & (!sk[10]) & (!g237) & (!g238)) + ((!i_36_) & (g11) & (!i_16_) & (!sk[10]) & (g237) & (!g238)));
	assign g240 = (((g56) & (!g183) & (!sk[11]) & (!g231) & (!g236) & (!g239)) + ((!g56) & (g183) & (!sk[11]) & (!g231) & (!g236) & (!g239)) + ((!g56) & (!g183) & (sk[11]) & (!g231) & (!g236) & (!g239)) + ((!g56) & (!g183) & (sk[11]) & (!g231) & (g236) & (!g239)));
	assign g241 = (((g10) & (!i_2_) & (!i_1_) & (!i_0_) & (!sk[12]) & (!g67)) + ((!g10) & (i_2_) & (!i_1_) & (!i_0_) & (!sk[12]) & (!g67)) + ((!g10) & (i_2_) & (!i_1_) & (i_0_) & (!sk[12]) & (!g67)) + ((!g10) & (!i_2_) & (!i_1_) & (i_0_) & (sk[12]) & (!g67)) + ((!g10) & (!i_2_) & (!i_1_) & (i_0_) & (sk[12]) & (!g67)));
	assign g242 = (((!i_37_) & (!i_32_) & (!i_25_) & (!g69) & (g226) & (!g241)) + ((i_37_) & (!i_32_) & (!i_25_) & (g69) & (!g226) & (g241)));
	assign g243 = (((!i_22_) & (g125) & (!sk[14]) & (!i_21_) & (!g198)) + ((!i_22_) & (!g125) & (!sk[14]) & (i_21_) & (!g198)) + ((!i_22_) & (g125) & (!sk[14]) & (!i_21_) & (g198)) + ((!i_22_) & (g125) & (!sk[14]) & (!i_21_) & (g198)));
	assign g244 = (((!i_37_) & (i_38_) & (!g187) & (!sk[15]) & (!g243)) + ((!i_37_) & (!i_38_) & (g187) & (!sk[15]) & (!g243)) + ((!i_37_) & (!i_38_) & (g187) & (!sk[15]) & (g243)) + ((i_37_) & (!i_38_) & (!g187) & (sk[15]) & (g243)));
	assign g245 = (((i_37_) & (!i_38_) & (!sk[16]) & (!i_39_) & (!i_40_) & (!g92)) + ((!i_37_) & (i_38_) & (!sk[16]) & (!i_39_) & (!i_40_) & (!g92)) + ((!i_37_) & (i_38_) & (!sk[16]) & (i_39_) & (!i_40_) & (!g92)) + ((!i_37_) & (i_38_) & (!sk[16]) & (!i_39_) & (!i_40_) & (!g92)) + ((i_37_) & (!i_38_) & (!sk[16]) & (!i_39_) & (i_40_) & (!g92)) + ((!i_37_) & (!i_38_) & (sk[16]) & (!i_39_) & (!i_40_) & (g92)));
	assign g246 = (((!sk[17]) & (!g27) & (g115)) + ((!sk[17]) & (g27) & (g115)));
	assign g247 = (((!i_13_) & (!sk[18]) & (g45) & (!g76) & (!g246)) + ((!i_13_) & (!sk[18]) & (!g45) & (g76) & (!g246)) + ((i_13_) & (sk[18]) & (!g45) & (!g76) & (!g246)) + ((!i_13_) & (sk[18]) & (!g45) & (!g76) & (!g246)) + ((!i_13_) & (sk[18]) & (!g45) & (!g76) & (!g246)));
	assign g248 = (((!sk[19]) & (!i_5_) & (i_12_) & (!i_13_) & (!i_15_)) + ((!sk[19]) & (!i_5_) & (!i_12_) & (i_13_) & (!i_15_)) + ((sk[19]) & (!i_5_) & (!i_12_) & (!i_13_) & (i_15_)) + ((sk[19]) & (!i_5_) & (!i_12_) & (!i_13_) & (!i_15_)));
	assign g249 = (((!sk[20]) & (g106) & (!g202) & (!g165) & (!g247) & (!g248)) + ((!sk[20]) & (!g106) & (g202) & (!g165) & (!g247) & (!g248)) + ((!sk[20]) & (g106) & (g202) & (g165) & (!g247) & (!g248)) + ((!sk[20]) & (g106) & (!g202) & (!g165) & (!g247) & (g248)));
	assign g250 = (((i_37_) & (!i_38_) & (!i_39_) & (!i_34_) & (!sk[21]) & (!g51)) + ((!i_37_) & (i_38_) & (!i_39_) & (!i_34_) & (!sk[21]) & (!g51)) + ((!i_37_) & (i_38_) & (i_39_) & (!i_34_) & (!sk[21]) & (g51)) + ((i_37_) & (!i_38_) & (!i_39_) & (!i_34_) & (!sk[21]) & (g51)));
	assign g251 = (((!sk[22]) & (!i_2_) & (i_1_) & (!g49) & (!i_0_)) + ((!sk[22]) & (!i_2_) & (!i_1_) & (g49) & (!i_0_)) + ((sk[22]) & (i_2_) & (!i_1_) & (!g49) & (i_0_)));
	assign g252 = (((i_11_) & (!g122) & (!sk[23]) & (!i_5_) & (!i_12_) & (!i_15_)) + ((!i_11_) & (g122) & (!sk[23]) & (!i_5_) & (!i_12_) & (!i_15_)) + ((i_11_) & (!g122) & (!sk[23]) & (!i_5_) & (!i_12_) & (i_15_)) + ((!i_11_) & (!g122) & (sk[23]) & (!i_5_) & (i_12_) & (i_15_)));
	assign g253 = (((i_36_) & (!i_37_) & (!sk[24]) & (!i_40_) & (!i_32_) & (!g67)) + ((!i_36_) & (i_37_) & (!sk[24]) & (!i_40_) & (!i_32_) & (!g67)) + ((!i_36_) & (!i_37_) & (sk[24]) & (!i_40_) & (!i_32_) & (g67)));
	assign g254 = (((!g250) & (g251) & (!sk[25]) & (!g252) & (!g253)) + ((g250) & (!g251) & (!sk[25]) & (g252) & (!g253)) + ((!g250) & (!g251) & (!sk[25]) & (g252) & (!g253)) + ((!g250) & (g251) & (!sk[25]) & (!g252) & (g253)));
	assign g255 = (((!i_33_) & (!sk[26]) & (g51)) + ((!i_33_) & (sk[26]) & (!g51)) + ((!i_33_) & (!sk[26]) & (g51)));
	assign g256 = (((!i_12_) & (g11) & (!sk[27]) & (!i_17_) & (!g232)) + ((!i_12_) & (!g11) & (!sk[27]) & (i_17_) & (!g232)) + ((i_12_) & (g11) & (!sk[27]) & (!i_17_) & (g232)));
	assign g257 = (((!i_32_) & (i_5_) & (!g24) & (!sk[28]) & (!g37)) + ((!i_32_) & (!i_5_) & (g24) & (!sk[28]) & (!g37)) + ((!i_32_) & (!i_5_) & (g24) & (!sk[28]) & (g37)));
	assign g258 = (((g56) & (g46) & (!g113) & (!g255) & (g256) & (!g257)) + ((g56) & (g46) & (!g113) & (!g255) & (!g256) & (g257)) + ((!g56) & (!g46) & (g113) & (!g255) & (!g256) & (g257)));
	assign g259 = (((!g134) & (!g244) & (!g245) & (!g249) & (!g254) & (!g258)) + ((!g134) & (!g244) & (!g245) & (!g249) & (!g254) & (!g258)));
	assign g260 = (((!i_38_) & (!sk[31]) & (i_39_) & (!i_40_)) + ((i_38_) & (!sk[31]) & (!i_39_) & (i_40_)) + ((i_38_) & (!sk[31]) & (i_39_) & (!i_40_)));
	assign g261 = (((g51) & (!i_31_) & (!i_5_) & (!i_9_) & (g260) & (!i_14_)) + ((g51) & (i_31_) & (!i_5_) & (!i_9_) & (!g260) & (!i_14_)));
	assign g262 = (((i_36_) & (i_37_) & (!i_38_) & (i_39_) & (!i_40_) & (!i_35_)) + ((!i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (i_35_)) + ((i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (!i_35_)) + ((i_36_) & (!i_37_) & (i_38_) & (!i_39_) & (i_40_) & (i_35_)) + ((i_36_) & (!i_37_) & (i_38_) & (i_39_) & (!i_40_) & (i_35_)) + ((!i_36_) & (i_37_) & (!i_38_) & (i_39_) & (!i_40_) & (i_35_)));
	assign g263 = (((!sk[34]) & (!g65) & (g175) & (!g740) & (!g261) & (!g262)) + ((!sk[34]) & (g65) & (!g175) & (!g740) & (!g261) & (!g262)) + ((!sk[34]) & (g65) & (!g175) & (!g740) & (!g261) & (!g262)) + ((!sk[34]) & (g65) & (!g175) & (!g740) & (g261) & (!g262)) + ((!sk[34]) & (g65) & (!g175) & (!g740) & (!g261) & (g262)));
	assign g264 = (((!sk[35]) & (!i_37_) & (i_38_) & (!g65) & (!i_5_)) + ((!sk[35]) & (!i_37_) & (!i_38_) & (g65) & (!i_5_)) + ((!sk[35]) & (i_37_) & (!i_38_) & (g65) & (!i_5_)));
	assign g265 = (((i_37_) & (!sk[36]) & (!g115) & (!g125) & (!i_0_) & (!g264)) + ((!i_37_) & (!sk[36]) & (g115) & (!g125) & (!i_0_) & (!g264)) + ((!i_37_) & (!sk[36]) & (g115) & (!g125) & (!i_0_) & (g264)) + ((i_37_) & (!sk[36]) & (g115) & (g125) & (i_0_) & (!g264)));
	assign g266 = (((!g260) & (!sk[37]) & (i_21_) & (!i_23_)) + ((g260) & (!sk[37]) & (!i_21_) & (i_23_)) + ((g260) & (sk[37]) & (!i_21_) & (!i_23_)));
	assign g267 = (((!g122) & (!sk[38]) & (i_22_) & (!i_21_)) + ((!g122) & (sk[38]) & (!i_22_) & (!i_21_)) + ((g122) & (!sk[38]) & (!i_22_) & (i_21_)) + ((!g122) & (!sk[38]) & (i_22_) & (!i_21_)));
	assign g268 = (((i_40_) & (!sk[39]) & (!i_32_) & (!i_16_) & (!g215) & (!g255)) + ((!i_40_) & (!sk[39]) & (i_32_) & (!i_16_) & (!g215) & (!g255)) + ((!i_40_) & (sk[39]) & (!i_32_) & (!i_16_) & (g215) & (!g255)));
	assign g269 = (((!g22) & (i_15_) & (!sk[40]) & (!g232)) + ((!g22) & (i_15_) & (!sk[40]) & (g232)) + ((g22) & (!i_15_) & (!sk[40]) & (g232)));
	assign g270 = (((i_18_) & (!g152) & (!i_21_) & (!g268) & (!sk[41]) & (!g269)) + ((!i_18_) & (g152) & (!i_21_) & (!g268) & (!sk[41]) & (!g269)) + ((!i_18_) & (!g152) & (!i_21_) & (g268) & (sk[41]) & (g269)) + ((!i_18_) & (!g152) & (!i_21_) & (!g268) & (sk[41]) & (g269)));
	assign g271 = (((!sk[42]) & (g198) & (!g263) & (!g265) & (!g729) & (!g270)) + ((!sk[42]) & (!g198) & (g263) & (!g265) & (!g729) & (!g270)) + ((sk[42]) & (!g198) & (!g263) & (!g265) & (!g729) & (!g270)) + ((!sk[42]) & (g198) & (!g263) & (!g265) & (g729) & (!g270)));
	assign g272 = (((!i_24_) & (!sk[43]) & (g125) & (!g198)) + ((i_24_) & (!sk[43]) & (!g125) & (g198)) + ((!i_24_) & (!sk[43]) & (g125) & (g198)));
	assign g273 = (((!i_30_) & (i_28_) & (!sk[44]) & (!i_29_)) + ((i_30_) & (!i_28_) & (!sk[44]) & (i_29_)) + ((!i_30_) & (!i_28_) & (sk[44]) & (!i_29_)));
	assign g274 = (((!sk[45]) & (!i_37_) & (i_38_) & (!i_39_) & (!g232)) + ((!sk[45]) & (!i_37_) & (!i_38_) & (i_39_) & (!g232)) + ((!sk[45]) & (i_37_) & (i_38_) & (i_39_) & (g232)));
	assign g275 = (((!i_36_) & (i_38_) & (!sk[46]) & (!i_39_)) + ((!i_36_) & (i_38_) & (!sk[46]) & (i_39_)) + ((i_36_) & (!i_38_) & (!sk[46]) & (i_39_)));
	assign g276 = (((i_12_) & (!i_15_) & (!i_17_) & (!g232) & (!sk[47]) & (!g275)) + ((!i_12_) & (i_15_) & (!i_17_) & (!g232) & (!sk[47]) & (!g275)) + ((i_12_) & (i_15_) & (!i_17_) & (g232) & (!sk[47]) & (g275)));
	assign g277 = (((!sk[48]) & (!g131) & (g163) & (!g274) & (!g276)) + ((!sk[48]) & (!g131) & (!g163) & (g274) & (!g276)) + ((sk[48]) & (!g131) & (!g163) & (!g274) & (!g276)) + ((!sk[48]) & (!g131) & (g163) & (!g274) & (!g276)));
	assign g278 = (((!sk[49]) & (!i_5_) & (g105) & (!g273) & (!g277)) + ((!sk[49]) & (!i_5_) & (!g105) & (g273) & (!g277)) + ((!sk[49]) & (!i_5_) & (!g105) & (g273) & (g277)) + ((sk[49]) & (!i_5_) & (!g105) & (!g273) & (g277)) + ((!sk[49]) & (i_5_) & (g105) & (!g273) & (g277)));
	assign g279 = (((g102) & (!i_10_) & (!i_27_) & (!sk[50]) & (!g73) & (!g216)) + ((!g102) & (i_10_) & (!i_27_) & (!sk[50]) & (!g73) & (!g216)) + ((g102) & (i_10_) & (i_27_) & (!sk[50]) & (g73) & (g216)));
	assign g280 = (((!sk[51]) & (!i_36_) & (g10) & (!g116)) + ((!sk[51]) & (i_36_) & (!g10) & (g116)));
	assign g281 = (((!i_36_) & (!sk[52]) & (g14)) + ((!i_36_) & (!sk[52]) & (g14)));
	assign g282 = (((i_32_) & (!i_2_) & (!i_1_) & (!i_0_) & (!sk[53]) & (!g67)) + ((!i_32_) & (i_2_) & (!i_1_) & (!i_0_) & (!sk[53]) & (!g67)) + ((!i_32_) & (i_2_) & (!i_1_) & (i_0_) & (!sk[53]) & (g67)));
	assign g283 = (((!g49) & (g280) & (!sk[54]) & (!g281) & (!g282)) + ((!g49) & (!g280) & (!sk[54]) & (g281) & (!g282)) + ((!g49) & (g280) & (!sk[54]) & (!g281) & (g282)) + ((!g49) & (!g280) & (!sk[54]) & (g281) & (g282)));
	assign g284 = (((!g21) & (!sk[55]) & (g47) & (!g130) & (!g184)) + ((!g21) & (!sk[55]) & (!g47) & (g130) & (!g184)) + ((!g21) & (!sk[55]) & (g47) & (!g130) & (g184)) + ((!g21) & (sk[55]) & (!g47) & (!g130) & (g184)) + ((!g21) & (!sk[55]) & (!g47) & (g130) & (g184)));
	assign g285 = (((g112) & (!g272) & (!g279) & (!g283) & (!sk[56]) & (!g284)) + ((!g112) & (g272) & (!g279) & (!g283) & (!sk[56]) & (!g284)) + ((!g112) & (!g272) & (!g279) & (!g283) & (sk[56]) & (g284)) + ((!g112) & (!g272) & (!g279) & (!g283) & (sk[56]) & (g284)));
	assign g286 = (((g102) & (!sk[57]) & (!g14) & (!g272) & (!g278) & (!g285)) + ((!g102) & (!sk[57]) & (g14) & (!g272) & (!g278) & (!g285)) + ((!g102) & (sk[57]) & (!g14) & (!g272) & (!g278) & (g285)) + ((!g102) & (!sk[57]) & (g14) & (!g272) & (!g278) & (g285)) + ((!g102) & (sk[57]) & (!g14) & (!g272) & (g278) & (g285)) + ((!g102) & (!sk[57]) & (g14) & (!g272) & (g278) & (g285)));
	assign g287 = (((g240) & (!sk[58]) & (!g242) & (!g259) & (!g271) & (!g286)) + ((!g240) & (!sk[58]) & (g242) & (!g259) & (!g271) & (!g286)) + ((g240) & (!sk[58]) & (!g242) & (g259) & (g271) & (g286)));
	assign g288 = (((i_7_) & (!sk[59]) & (!i_5_) & (!i_30_) & (!i_28_) & (!i_29_)) + ((!i_7_) & (!sk[59]) & (i_5_) & (!i_30_) & (!i_28_) & (!i_29_)) + ((!i_7_) & (sk[59]) & (!i_5_) & (!i_30_) & (i_28_) & (i_29_)) + ((!i_7_) & (sk[59]) & (!i_5_) & (!i_30_) & (!i_28_) & (!i_29_)) + ((!i_7_) & (sk[59]) & (!i_5_) & (i_30_) & (!i_28_) & (!i_29_)));
	assign g289 = (((!sk[60]) & (!g1) & (i_30_) & (!i_29_) & (!g288)) + ((!sk[60]) & (!g1) & (!i_30_) & (i_29_) & (!g288)) + ((!sk[60]) & (!g1) & (i_30_) & (!i_29_) & (!g288)) + ((sk[60]) & (!g1) & (!i_30_) & (!i_29_) & (!g288)) + ((!sk[60]) & (g1) & (!i_30_) & (i_29_) & (!g288)));
	assign g290 = (((g65) & (!g1) & (!i_15_) & (!sk[61]) & (!i_24_) & (!g151)) + ((!g65) & (g1) & (!i_15_) & (!sk[61]) & (!i_24_) & (!g151)) + ((g65) & (!g1) & (!i_15_) & (!sk[61]) & (!i_24_) & (g151)) + ((g65) & (!g1) & (!i_15_) & (!sk[61]) & (i_24_) & (g151)));
	assign g291 = (((g122) & (!g139) & (!sk[62]) & (!g119) & (!g289) & (!g290)) + ((!g122) & (g139) & (!sk[62]) & (!g119) & (!g289) & (!g290)) + ((!g122) & (g139) & (!sk[62]) & (!g119) & (!g289) & (g290)) + ((!g122) & (!g139) & (sk[62]) & (g119) & (!g289) & (!g290)));
	assign g292 = (((i_9_) & (!i_18_) & (!g153) & (!sk[63]) & (!g144) & (!g165)) + ((!i_9_) & (i_18_) & (!g153) & (!sk[63]) & (!g144) & (!g165)) + ((i_9_) & (!i_18_) & (g153) & (!sk[63]) & (g144) & (g165)) + ((!i_9_) & (i_18_) & (g153) & (!sk[63]) & (g144) & (g165)));
	assign g293 = (((!i_36_) & (!sk[64]) & (g56) & (!g48)) + ((i_36_) & (!sk[64]) & (!g56) & (g48)) + ((!i_36_) & (!sk[64]) & (g56) & (g48)));
	assign g294 = (((!sk[65]) & (!g102) & (g1) & (!g105) & (!g273)) + ((!sk[65]) & (!g102) & (!g1) & (g105) & (!g273)) + ((!sk[65]) & (g102) & (!g1) & (g105) & (g273)));
	assign g295 = (((i_31_) & (!i_5_) & (!sk[66]) & (!g24) & (!g293) & (!g294)) + ((!i_31_) & (i_5_) & (!sk[66]) & (!g24) & (!g293) & (!g294)) + ((!i_31_) & (i_5_) & (!sk[66]) & (!g24) & (!g293) & (!g294)) + ((!i_31_) & (!i_5_) & (sk[66]) & (!g24) & (!g293) & (!g294)) + ((!i_31_) & (!i_5_) & (sk[66]) & (!g24) & (!g293) & (!g294)) + ((!i_31_) & (!i_5_) & (sk[66]) & (!g24) & (!g293) & (!g294)));
	assign g296 = (((i_40_) & (!sk[67]) & (!g117) & (!g95) & (!g8) & (!g215)) + ((!i_40_) & (!sk[67]) & (g117) & (!g95) & (!g8) & (!g215)) + ((!i_40_) & (sk[67]) & (!g117) & (g95) & (g8) & (!g215)) + ((!i_40_) & (sk[67]) & (!g117) & (g95) & (!g8) & (g215)));
	assign g297 = (((!g1) & (i_12_) & (!i_15_) & (!sk[68]) & (!g194)) + ((!g1) & (!i_12_) & (i_15_) & (!sk[68]) & (!g194)) + ((!g1) & (!i_12_) & (!i_15_) & (sk[68]) & (g194)) + ((!g1) & (!i_12_) & (!i_15_) & (sk[68]) & (g194)));
	assign g298 = (((!g57) & (g130) & (!g8) & (!sk[69]) & (!g297)) + ((!g57) & (!g130) & (g8) & (!sk[69]) & (!g297)) + ((!g57) & (!g130) & (!g8) & (sk[69]) & (!g297)) + ((!g57) & (!g130) & (!g8) & (sk[69]) & (!g297)) + ((!g57) & (!g130) & (!g8) & (sk[69]) & (!g297)));
	assign g299 = (((!i_37_) & (i_38_) & (!i_39_) & (i_40_) & (g93) & (!g96)) + ((!i_37_) & (!i_38_) & (i_39_) & (!i_40_) & (!g93) & (g96)) + ((!i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (!g93) & (g96)));
	assign g300 = (((g292) & (!sk[71]) & (!g295) & (!g296) & (!g298) & (!g299)) + ((!g292) & (!sk[71]) & (g295) & (!g296) & (!g298) & (!g299)) + ((!g292) & (!sk[71]) & (g295) & (!g296) & (g298) & (!g299)));
	assign g301 = (((!g122) & (g1) & (!i_13_) & (!sk[72]) & (!i_15_)) + ((!g122) & (!g1) & (i_13_) & (!sk[72]) & (!i_15_)) + ((!g122) & (!g1) & (!i_13_) & (sk[72]) & (!i_15_)));
	assign g302 = (((!g2) & (g45) & (g128) & (!sk[73]) & (!g98) & (!g301)) + ((g2) & (!g45) & (!g128) & (!sk[73]) & (!g98) & (!g301)) + ((!g2) & (g45) & (!g128) & (!sk[73]) & (!g98) & (!g301)) + ((g2) & (!g45) & (!g128) & (!sk[73]) & (g98) & (g301)));
	assign g303 = (((i_36_) & (g100) & (!g10) & (g48) & (i_25_) & (!i_26_)) + ((i_36_) & (g100) & (!g10) & (g48) & (!i_25_) & (!i_26_)));
	assign g304 = (((!sk[75]) & (i_7_) & (!g102) & (!i_10_) & (!i_27_) & (!g216)) + ((!sk[75]) & (!i_7_) & (g102) & (!i_10_) & (!i_27_) & (!g216)) + ((!sk[75]) & (!i_7_) & (g102) & (!i_10_) & (!i_27_) & (g216)) + ((!sk[75]) & (!i_7_) & (g102) & (!i_10_) & (!i_27_) & (g216)));
	assign g305 = (((!sk[76]) & (i_40_) & (!i_34_) & (!g6) & (!g78) & (!g225)) + ((!sk[76]) & (!i_40_) & (i_34_) & (!g6) & (!g78) & (!g225)) + ((!sk[76]) & (!i_40_) & (i_34_) & (g6) & (g78) & (g225)));
	assign g306 = (((i_38_) & (!g101) & (!i_35_) & (!sk[77]) & (!g70) & (!g163)) + ((!i_38_) & (g101) & (!i_35_) & (!sk[77]) & (!g70) & (!g163)) + ((!i_38_) & (g101) & (!i_35_) & (!sk[77]) & (g70) & (g163)));
	assign g307 = (((!i_7_) & (i_33_) & (!sk[78]) & (!g11)) + ((!i_7_) & (i_33_) & (!sk[78]) & (g11)) + ((i_7_) & (!i_33_) & (!sk[78]) & (g11)));
	assign g308 = (((i_5_) & (!g22) & (!i_16_) & (!i_17_) & (!sk[79]) & (!i_9_)) + ((!i_5_) & (g22) & (!i_16_) & (!i_17_) & (!sk[79]) & (!i_9_)) + ((!i_5_) & (!g22) & (i_16_) & (i_17_) & (sk[79]) & (!i_9_)) + ((!i_5_) & (!g22) & (i_16_) & (!i_17_) & (sk[79]) & (i_9_)) + ((!i_5_) & (!g22) & (!i_16_) & (i_17_) & (sk[79]) & (i_9_)));
	assign g309 = (((!sk[80]) & (g2) & (!g21) & (!g113) & (!g307) & (!g308)) + ((!sk[80]) & (!g2) & (g21) & (!g113) & (!g307) & (!g308)) + ((!sk[80]) & (g2) & (g21) & (!g113) & (g307) & (g308)) + ((!sk[80]) & (g2) & (!g21) & (g113) & (g307) & (g308)));
	assign g310 = (((!sk[81]) & (i_37_) & (!i_35_) & (!g65) & (!g21) & (!g79)) + ((!sk[81]) & (!i_37_) & (i_35_) & (!g65) & (!g21) & (!g79)) + ((!sk[81]) & (i_37_) & (!i_35_) & (g65) & (!g21) & (!g79)) + ((sk[81]) & (!i_37_) & (!i_35_) & (g65) & (!g21) & (!g79)));
	assign g311 = (((!i_36_) & (i_31_) & (!sk[82]) & (!g1)) + ((i_36_) & (!i_31_) & (!sk[82]) & (g1)) + ((!i_36_) & (i_31_) & (!sk[82]) & (!g1)));
	assign g312 = (((g102) & (!sk[83]) & (!i_9_) & (!g171) & (!g310) & (!g311)) + ((!g102) & (!sk[83]) & (i_9_) & (!g171) & (!g310) & (!g311)) + ((!g102) & (sk[83]) & (!i_9_) & (!g171) & (g310) & (g311)) + ((g102) & (!sk[83]) & (!i_9_) & (!g171) & (!g310) & (g311)));
	assign g313 = (((g201) & (!g305) & (!sk[84]) & (!g306) & (!g309) & (!g312)) + ((!g201) & (g305) & (!sk[84]) & (!g306) & (!g309) & (!g312)) + ((g201) & (!g305) & (!sk[84]) & (!g306) & (!g309) & (!g312)) + ((!g201) & (!g305) & (sk[84]) & (!g306) & (!g309) & (!g312)));
	assign g314 = (((i_39_) & (!i_40_) & (!g302) & (!g303) & (!g304) & (g313)) + ((i_39_) & (!i_40_) & (!g302) & (!g303) & (!g304) & (g313)) + ((!i_39_) & (!i_40_) & (!g302) & (!g303) & (!g304) & (g313)) + ((!i_39_) & (!i_40_) & (!g302) & (!g303) & (!g304) & (g313)));
	assign g315 = (((!sk[86]) & (!i_40_) & (g8)) + ((!sk[86]) & (i_40_) & (g8)));
	assign g316 = (((!sk[87]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (!g121)) + ((!sk[87]) & (!i_37_) & (i_38_) & (!i_39_) & (!i_40_) & (!g121)) + ((!sk[87]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (g121)) + ((!sk[87]) & (i_37_) & (!i_38_) & (i_39_) & (i_40_) & (g121)));
	assign g317 = (((i_36_) & (!i_37_) & (!i_34_) & (!g77) & (!sk[88]) & (!g316)) + ((!i_36_) & (i_37_) & (!i_34_) & (!g77) & (!sk[88]) & (!g316)) + ((!i_36_) & (i_37_) & (!i_34_) & (!g77) & (!sk[88]) & (!g316)) + ((!i_36_) & (!i_37_) & (!i_34_) & (!g77) & (sk[88]) & (!g316)) + ((!i_36_) & (!i_37_) & (i_34_) & (!g77) & (sk[88]) & (!g316)) + ((!i_36_) & (!i_37_) & (!i_34_) & (!g77) & (sk[88]) & (!g316)));
	assign g318 = (((!i_37_) & (g260) & (!sk[89]) & (!g5)) + ((i_37_) & (g260) & (!sk[89]) & (g5)) + ((i_37_) & (!g260) & (!sk[89]) & (g5)));
	assign g319 = (((g61) & (!g92) & (g160) & (!sk[90]) & (!g318)) + ((!g61) & (g92) & (!g160) & (!sk[90]) & (!g318)) + ((!g61) & (!g92) & (g160) & (!sk[90]) & (!g318)) + ((!g61) & (g92) & (!g160) & (!sk[90]) & (g318)));
	assign g320 = (((!sk[91]) & (i_34_) & (!g78) & (!g315) & (!g317) & (!g319)) + ((!sk[91]) & (!i_34_) & (g78) & (!g315) & (!g317) & (!g319)) + ((!sk[91]) & (i_34_) & (!g78) & (!g315) & (g317) & (!g319)) + ((sk[91]) & (!i_34_) & (!g78) & (!g315) & (g317) & (!g319)) + ((!sk[91]) & (!i_34_) & (g78) & (!g315) & (g317) & (!g319)));
	assign g321 = (((i_7_) & (!i_33_) & (!i_32_) & (!sk[92]) & (!g150) & (!g320)) + ((!i_7_) & (i_33_) & (!i_32_) & (!sk[92]) & (!g150) & (!g320)) + ((i_7_) & (!i_33_) & (!i_32_) & (!sk[92]) & (g150) & (!g320)) + ((!i_7_) & (!i_33_) & (!i_32_) & (sk[92]) & (g150) & (!g320)) + ((!i_7_) & (!i_33_) & (i_32_) & (sk[92]) & (g150) & (!g320)) + ((!i_7_) & (!i_33_) & (!i_32_) & (sk[92]) & (g150) & (g320)));
	assign g322 = (((i_36_) & (!sk[93]) & (!g100) & (!g101) & (!g102) & (!i_13_)) + ((!i_36_) & (!sk[93]) & (g100) & (!g101) & (!g102) & (!i_13_)) + ((!i_36_) & (!sk[93]) & (g100) & (g101) & (g102) & (!i_13_)));
	assign g323 = (((i_39_) & (!i_32_) & (!i_13_) & (!g45) & (!sk[94]) & (!g49)) + ((!i_39_) & (i_32_) & (!i_13_) & (!g45) & (!sk[94]) & (!g49)) + ((i_39_) & (!i_32_) & (i_13_) & (g45) & (!sk[94]) & (!g49)));
	assign g324 = (((!sk[95]) & (i_40_) & (!g125) & (!g225) & (!g322) & (!g323)) + ((!sk[95]) & (!i_40_) & (g125) & (!g225) & (!g322) & (!g323)) + ((sk[95]) & (!i_40_) & (!g125) & (!g225) & (!g322) & (!g323)) + ((sk[95]) & (!i_40_) & (!g125) & (!g225) & (!g322) & (!g323)) + ((!sk[95]) & (!i_40_) & (g125) & (!g225) & (!g322) & (!g323)));
	assign g325 = (((!sk[96]) & (g23) & (!g18) & (!i_18_) & (!g155) & (!i_19_)) + ((!sk[96]) & (!g23) & (g18) & (!i_18_) & (!g155) & (!i_19_)) + ((!sk[96]) & (!g23) & (g18) & (i_18_) & (g155) & (!i_19_)) + ((!sk[96]) & (g23) & (!g18) & (i_18_) & (!g155) & (i_19_)) + ((!sk[96]) & (!g23) & (g18) & (!i_18_) & (g155) & (i_19_)));
	assign g326 = (((!sk[97]) & (g57) & (!g125) & (!i_23_) & (!g153) & (!g325)) + ((!sk[97]) & (!g57) & (g125) & (!i_23_) & (!g153) & (!g325)) + ((!sk[97]) & (g57) & (g125) & (!i_23_) & (!g153) & (!g325)) + ((!sk[97]) & (!g57) & (g125) & (i_23_) & (g153) & (g325)));
	assign g327 = (((!sk[98]) & (i_37_) & (!g30) & (!g54) & (!g324) & (!g326)) + ((!sk[98]) & (!i_37_) & (g30) & (!g54) & (!g324) & (!g326)) + ((sk[98]) & (!i_37_) & (!g30) & (g54) & (!g324) & (!g326)) + ((!sk[98]) & (i_37_) & (!g30) & (!g54) & (!g324) & (g326)));
	assign g328 = (((g291) & (!sk[99]) & (!g300) & (!g314) & (!g321) & (!g327)) + ((!g291) & (!sk[99]) & (g300) & (!g314) & (!g321) & (!g327)) + ((!g291) & (!sk[99]) & (g300) & (g314) & (g321) & (!g327)));
	assign g329 = (((!sk[100]) & (!g25) & (g136) & (!g79)) + ((!sk[100]) & (g25) & (!g136) & (g79)) + ((!sk[100]) & (g25) & (g136) & (g79)));
	assign g330 = (((!sk[101]) & (i_7_) & (!i_2_) & (!i_1_) & (!i_0_) & (!g67)) + ((!sk[101]) & (!i_7_) & (i_2_) & (!i_1_) & (!i_0_) & (!g67)) + ((!sk[101]) & (!i_7_) & (i_2_) & (!i_1_) & (i_0_) & (g67)));
	assign g331 = (((!i_38_) & (g66) & (!sk[102]) & (!g330)) + ((i_38_) & (g66) & (!sk[102]) & (g330)) + ((i_38_) & (!g66) & (!sk[102]) & (g330)));
	assign g332 = (((!g124) & (!sk[103]) & (g148) & (!g331)) + ((g124) & (!sk[103]) & (!g148) & (g331)) + ((!g124) & (sk[103]) & (!g148) & (!g331)) + ((!g124) & (!sk[103]) & (g148) & (!g331)));
	assign g333 = (((!i_32_) & (!sk[104]) & (g54) & (!i_13_) & (!g10)) + ((!i_32_) & (!sk[104]) & (!g54) & (i_13_) & (!g10)) + ((!i_32_) & (!sk[104]) & (g54) & (!i_13_) & (!g10)));
	assign g334 = (((!i_36_) & (g100) & (!g76) & (!sk[105]) & (!g333)) + ((!i_36_) & (!g100) & (g76) & (!sk[105]) & (!g333)) + ((!i_36_) & (g100) & (g76) & (!sk[105]) & (g333)));
	assign g335 = (((i_31_) & (!sk[106]) & (!g54) & (!i_13_) & (!g180) & (!g334)) + ((!i_31_) & (!sk[106]) & (g54) & (!i_13_) & (!g180) & (!g334)) + ((i_31_) & (!sk[106]) & (!g54) & (!i_13_) & (!g180) & (!g334)) + ((!i_31_) & (sk[106]) & (!g54) & (!i_13_) & (!g180) & (!g334)) + ((!i_31_) & (!sk[106]) & (g54) & (!i_13_) & (!g180) & (!g334)) + ((!i_31_) & (!sk[106]) & (g54) & (!i_13_) & (!g180) & (!g334)));
	assign g336 = (((!g138) & (!sk[107]) & (i_30_) & (!i_29_)) + ((g138) & (!sk[107]) & (!i_30_) & (i_29_)) + ((g138) & (sk[107]) & (!i_30_) & (!i_29_)));
	assign g337 = (((!g1) & (g44) & (g46) & (!sk[108]) & (!g105) & (!g336)) + ((g1) & (!g44) & (!g46) & (!sk[108]) & (!g105) & (!g336)) + ((!g1) & (g44) & (!g46) & (!sk[108]) & (!g105) & (!g336)) + ((!g1) & (!g44) & (!g46) & (sk[108]) & (g105) & (g336)));
	assign g338 = (((!i_38_) & (!sk[109]) & (g51) & (!g76)) + ((i_38_) & (!sk[109]) & (!g51) & (g76)) + ((i_38_) & (!sk[109]) & (g51) & (g76)));
	assign g339 = (((!g53) & (!sk[110]) & (g107) & (!g338)) + ((g53) & (!sk[110]) & (!g107) & (g338)) + ((g53) & (!sk[110]) & (g107) & (g338)));
	assign g340 = (((!i_36_) & (i_38_) & (!i_39_) & (!sk[111]) & (!g92)) + ((!i_36_) & (!i_38_) & (i_39_) & (!sk[111]) & (!g92)) + ((!i_36_) & (i_38_) & (!i_39_) & (!sk[111]) & (!g92)) + ((i_36_) & (!i_38_) & (!i_39_) & (sk[111]) & (!g92)));
	assign g341 = (((!i_36_) & (i_37_) & (!i_38_) & (!sk[112]) & (!i_35_)) + ((!i_36_) & (!i_37_) & (i_38_) & (!sk[112]) & (!i_35_)) + ((!i_36_) & (i_37_) & (!i_38_) & (!sk[112]) & (i_35_)) + ((i_36_) & (i_37_) & (!i_38_) & (!sk[112]) & (!i_35_)) + ((i_36_) & (!i_37_) & (!i_38_) & (sk[112]) & (i_35_)));
	assign g342 = (((i_37_) & (!i_40_) & (!sk[113]) & (!i_34_) & (!g6) & (!g341)) + ((!i_37_) & (i_40_) & (!sk[113]) & (!i_34_) & (!g6) & (!g341)) + ((!i_37_) & (!i_40_) & (sk[113]) & (!i_34_) & (g6) & (g341)) + ((!i_37_) & (!i_40_) & (sk[113]) & (!i_34_) & (g6) & (g341)));
	assign g343 = (((i_37_) & (!i_39_) & (!i_40_) & (!g7) & (!sk[114]) & (!g95)) + ((!i_37_) & (i_39_) & (!i_40_) & (!g7) & (!sk[114]) & (!g95)) + ((!i_37_) & (i_39_) & (!i_40_) & (g7) & (!sk[114]) & (!g95)) + ((!i_37_) & (i_39_) & (i_40_) & (!g7) & (!sk[114]) & (g95)));
	assign g344 = (((g303) & (!sk[115]) & (!g339) & (!g340) & (!g342) & (!g343)) + ((!g303) & (!sk[115]) & (g339) & (!g340) & (!g342) & (!g343)) + ((!g303) & (sk[115]) & (!g339) & (g340) & (!g342) & (!g343)) + ((!g303) & (sk[115]) & (!g339) & (!g340) & (!g342) & (!g343)));
	assign g345 = (((g329) & (!sk[116]) & (!g332) & (!g335) & (!g337) & (!g344)) + ((!g329) & (!sk[116]) & (g332) & (!g335) & (!g337) & (!g344)) + ((!g329) & (!sk[116]) & (g332) & (g335) & (!g337) & (g344)));
	assign g346 = (((!sk[117]) & (!i_37_) & (g104)) + ((!sk[117]) & (i_37_) & (g104)));
	assign g347 = (((!i_38_) & (g70) & (!sk[118]) & (!g78)) + ((i_38_) & (g70) & (!sk[118]) & (g78)) + ((i_38_) & (!g70) & (!sk[118]) & (g78)));
	assign g348 = (((!sk[119]) & (g47) & (!i_0_) & (!g93) & (!g346) & (!g347)) + ((!sk[119]) & (!g47) & (i_0_) & (!g93) & (!g346) & (!g347)) + ((sk[119]) & (!g47) & (!i_0_) & (g93) & (g346) & (!g347)) + ((!sk[119]) & (!g47) & (i_0_) & (!g93) & (!g346) & (g347)));
	assign g349 = (((!i_37_) & (!i_38_) & (i_39_) & (!g121) & (!g148) & (!g301)) + ((i_37_) & (!i_38_) & (!i_39_) & (!g121) & (!g148) & (!g301)) + ((!i_37_) & (!i_38_) & (!i_39_) & (!g121) & (!g148) & (!g301)) + ((!i_37_) & (i_38_) & (!i_39_) & (!g121) & (!g148) & (!g301)) + ((!i_37_) & (!i_38_) & (!i_39_) & (!g121) & (!g148) & (!g301)) + ((!i_37_) & (!i_38_) & (i_39_) & (!g121) & (!g148) & (!g301)));
	assign g350 = (((!sk[121]) & (!i_33_) & (i_32_) & (!g51) & (!i_31_)) + ((!sk[121]) & (!i_33_) & (!i_32_) & (g51) & (!i_31_)) + ((!sk[121]) & (i_33_) & (!i_32_) & (g51) & (!i_31_)));
	assign g351 = (((!i_36_) & (g162) & (!sk[122]) & (!g48) & (!g98)) + ((!i_36_) & (!g162) & (!sk[122]) & (g48) & (!g98)) + ((i_36_) & (!g162) & (!sk[122]) & (g48) & (g98)));
	assign g352 = (((i_40_) & (!g44) & (!sk[123]) & (!g281) & (!g95) & (!g215)) + ((!i_40_) & (g44) & (!sk[123]) & (!g281) & (!g95) & (!g215)) + ((!i_40_) & (!g44) & (sk[123]) & (!g281) & (!g95) & (!g215)) + ((!i_40_) & (!g44) & (sk[123]) & (!g281) & (!g95) & (!g215)) + ((!i_40_) & (!g44) & (sk[123]) & (!g281) & (!g95) & (!g215)) + ((!i_40_) & (!g44) & (sk[123]) & (!g281) & (!g95) & (!g215)));
	assign g353 = (((!i_37_) & (!sk[124]) & (i_38_) & (!i_35_) & (!g65)) + ((!i_37_) & (!sk[124]) & (!i_38_) & (i_35_) & (!g65)) + ((i_37_) & (!sk[124]) & (!i_38_) & (i_35_) & (g65)));
	assign g354 = (((g57) & (!g68) & (!g215) & (!sk[125]) & (!g350) & (!g353)) + ((!g57) & (g68) & (!g215) & (!sk[125]) & (!g350) & (!g353)) + ((!g57) & (g68) & (!g215) & (!sk[125]) & (!g350) & (g353)) + ((g57) & (!g68) & (g215) & (!sk[125]) & (g350) & (!g353)));
	assign g355 = (((!g10) & (!sk[126]) & (g11) & (!i_21_)) + ((g10) & (!sk[126]) & (!g11) & (i_21_)) + ((!g10) & (!sk[126]) & (g11) & (!i_21_)));
	assign g356 = (((!sk[127]) & (!i_11_) & (g1) & (!i_12_) & (!g355)) + ((!sk[127]) & (!i_11_) & (!g1) & (i_12_) & (!g355)) + ((!sk[127]) & (!i_11_) & (!g1) & (i_12_) & (g355)) + ((sk[127]) & (i_11_) & (!g1) & (!i_12_) & (g355)));
	assign g357 = (((i_11_) & (!g1) & (!sk[0]) & (!g28) & (!g12) & (!g356)) + ((!i_11_) & (g1) & (!sk[0]) & (!g28) & (!g12) & (!g356)) + ((!i_11_) & (!g1) & (sk[0]) & (g28) & (!g12) & (g356)) + ((i_11_) & (!g1) & (!sk[0]) & (g28) & (g12) & (!g356)));
	assign g358 = (((g348) & (!g723) & (!sk[1]) & (!g352) & (!g354) & (!g357)) + ((!g348) & (g723) & (!sk[1]) & (!g352) & (!g354) & (!g357)) + ((!g348) & (g723) & (!sk[1]) & (!g352) & (!g354) & (!g357)) + ((!g348) & (!g723) & (sk[1]) & (g352) & (!g354) & (!g357)));
	assign g359 = (((!i_11_) & (g1) & (!g37) & (!sk[2]) & (!i_14_)) + ((!i_11_) & (!g1) & (g37) & (!sk[2]) & (!i_14_)) + ((i_11_) & (!g1) & (g37) & (!sk[2]) & (!i_14_)));
	assign g360 = (((g2) & (!g21) & (!sk[3]) & (!g136) & (!g79) & (!g359)) + ((!g2) & (g21) & (!sk[3]) & (!g136) & (!g79) & (!g359)) + ((g2) & (g21) & (!sk[3]) & (!g136) & (!g79) & (g359)) + ((!g2) & (!g21) & (sk[3]) & (g136) & (g79) & (g359)));
	assign g361 = (((!sk[4]) & (!g1) & (i_30_) & (!i_28_) & (!i_29_)) + ((!sk[4]) & (!g1) & (!i_30_) & (i_28_) & (!i_29_)) + ((sk[4]) & (!g1) & (!i_30_) & (!i_28_) & (!i_29_)) + ((!sk[4]) & (g1) & (!i_30_) & (i_28_) & (!i_29_)));
	assign g362 = (((i_37_) & (!i_38_) & (!i_34_) & (!g1) & (!sk[5]) & (!g361)) + ((!i_37_) & (i_38_) & (!i_34_) & (!g1) & (!sk[5]) & (!g361)) + ((i_37_) & (!i_38_) & (!i_34_) & (!g1) & (!sk[5]) & (!g361)));
	assign g363 = (((g100) & (!sk[6]) & (!g104) & (!g72) & (!g73) & (!g96)) + ((!g100) & (!sk[6]) & (g104) & (!g72) & (!g73) & (!g96)) + ((!g100) & (!sk[6]) & (g104) & (g72) & (!g73) & (!g96)) + ((g100) & (!sk[6]) & (!g104) & (!g72) & (!g73) & (g96)));
	assign g364 = (((g3) & (!g115) & (!g360) & (!sk[7]) & (!g362) & (!g363)) + ((!g3) & (g115) & (!g360) & (!sk[7]) & (!g362) & (!g363)) + ((!g3) & (!g115) & (!g360) & (sk[7]) & (!g362) & (!g363)) + ((!g3) & (!g115) & (!g360) & (sk[7]) & (!g362) & (!g363)) + ((!g3) & (!g115) & (!g360) & (sk[7]) & (!g362) & (!g363)));
	assign g365 = (((g122) & (!g1) & (!i_9_) & (!i_18_) & (!sk[8]) & (!i_21_)) + ((!g122) & (g1) & (!i_9_) & (!i_18_) & (!sk[8]) & (!i_21_)) + ((!g122) & (!g1) & (!i_9_) & (!i_18_) & (sk[8]) & (!i_21_)));
	assign g366 = (((!sk[9]) & (!g26) & (g37) & (!g365)) + ((!sk[9]) & (g26) & (!g37) & (g365)) + ((!sk[9]) & (!g26) & (g37) & (g365)));
	assign g367 = (((g122) & (!g121) & (!sk[10]) & (!i_21_) & (!g91) & (!g366)) + ((!g122) & (g121) & (!sk[10]) & (!i_21_) & (!g91) & (!g366)) + ((!g122) & (g121) & (!sk[10]) & (!i_21_) & (!g91) & (g366)) + ((!g122) & (g121) & (!sk[10]) & (!i_21_) & (g91) & (!g366)));
	assign g368 = (((i_37_) & (!g10) & (!sk[11]) & (!g48) & (!g115) & (!i_0_)) + ((!i_37_) & (g10) & (!sk[11]) & (!g48) & (!g115) & (!i_0_)) + ((i_37_) & (!g10) & (!sk[11]) & (g48) & (g115) & (i_0_)));
	assign g369 = (((!i_11_) & (!sk[12]) & (g1) & (!i_12_) & (!g12)) + ((!i_11_) & (!sk[12]) & (!g1) & (i_12_) & (!g12)) + ((!i_11_) & (!sk[12]) & (!g1) & (i_12_) & (g12)) + ((i_11_) & (sk[12]) & (!g1) & (!i_12_) & (g12)));
	assign g370 = (((i_40_) & (!sk[13]) & (!g14) & (!g356) & (!g368) & (!g369)) + ((!i_40_) & (!sk[13]) & (g14) & (!g356) & (!g368) & (!g369)) + ((!i_40_) & (sk[13]) & (!g14) & (!g356) & (!g368) & (!g369)) + ((i_40_) & (!sk[13]) & (!g14) & (!g356) & (!g368) & (!g369)) + ((!i_40_) & (!sk[13]) & (g14) & (!g356) & (!g368) & (!g369)));
	assign g371 = (((i_38_) & (g3) & (!i_16_) & (g34) & (g18) & (g73)));
	assign g372 = (((!g1) & (i_15_) & (!g3) & (!sk[15]) & (!g131)) + ((!g1) & (!i_15_) & (g3) & (!sk[15]) & (!g131)) + ((!g1) & (!i_15_) & (g3) & (!sk[15]) & (g131)));
	assign g373 = (((!i_38_) & (!sk[16]) & (g197) & (!g330) & (!g372)) + ((!i_38_) & (!sk[16]) & (!g197) & (g330) & (!g372)) + ((i_38_) & (sk[16]) & (!g197) & (!g330) & (!g372)) + ((!i_38_) & (sk[16]) & (!g197) & (!g330) & (!g372)) + ((!i_38_) & (sk[16]) & (!g197) & (!g330) & (!g372)));
	assign g374 = (((!i_15_) & (!sk[17]) & (i_21_) & (!i_23_) & (!g211)) + ((!i_15_) & (!sk[17]) & (!i_21_) & (i_23_) & (!g211)) + ((i_15_) & (sk[17]) & (!i_21_) & (!i_23_) & (g211)));
	assign g375 = (((!i_22_) & (!sk[18]) & (g11) & (!i_21_)) + ((!i_22_) & (!sk[18]) & (g11) & (!i_21_)) + ((i_22_) & (!sk[18]) & (!g11) & (i_21_)));
	assign g376 = (((!i_36_) & (g49) & (!sk[19]) & (!g131)) + ((i_36_) & (!g49) & (!sk[19]) & (g131)) + ((!i_36_) & (!g49) & (sk[19]) & (g131)));
	assign g377 = (((g143) & (!sk[20]) & (!g61) & (!i_23_) & (!g375) & (!g376)) + ((!g143) & (!sk[20]) & (g61) & (!i_23_) & (!g375) & (!g376)) + ((g143) & (!sk[20]) & (g61) & (!i_23_) & (!g375) & (!g376)) + ((!g143) & (sk[20]) & (!g61) & (!i_23_) & (g375) & (g376)));
	assign g378 = (((!g43) & (!g136) & (!g371) & (!g373) & (!g374) & (!g377)) + ((!g43) & (!g136) & (!g371) & (g373) & (!g374) & (!g377)) + ((!g43) & (!g136) & (!g371) & (!g373) & (!g374) & (!g377)) + ((!g43) & (!g136) & (!g371) & (g373) & (!g374) & (!g377)));
	assign g379 = (((i_36_) & (!sk[22]) & (!g21) & (!g367) & (!g370) & (!g378)) + ((!i_36_) & (!sk[22]) & (g21) & (!g367) & (!g370) & (!g378)) + ((i_36_) & (!sk[22]) & (!g21) & (!g367) & (!g370) & (g378)) + ((i_36_) & (!sk[22]) & (!g21) & (!g367) & (!g370) & (g378)) + ((!i_36_) & (sk[22]) & (!g21) & (!g367) & (g370) & (g378)) + ((!i_36_) & (!sk[22]) & (g21) & (!g367) & (g370) & (g378)));
	assign o_5_ = (((!g64) & (sk[23]) & (!g345) & (!g358) & (!g364) & (!g379)) + ((!g64) & (!sk[23]) & (g345) & (!g358) & (!g364) & (!g379)) + ((g64) & (!sk[23]) & (!g345) & (!g358) & (!g364) & (!g379)) + ((!g64) & (!sk[23]) & (g345) & (!g358) & (!g364) & (!g379)) + ((!g64) & (!sk[23]) & (g345) & (!g358) & (!g364) & (!g379)) + ((!g64) & (!sk[23]) & (g345) & (!g358) & (!g364) & (!g379)));
	assign g381 = (((!i_15_) & (g31) & (!sk[24]) & (!g98)) + ((!i_15_) & (g31) & (!sk[24]) & (g98)) + ((i_15_) & (!g31) & (!sk[24]) & (g98)));
	assign g382 = (((!i_11_) & (g95) & (!sk[25]) & (!g346) & (!g351)) + ((!i_11_) & (g95) & (!sk[25]) & (g346) & (!g351)) + ((!i_11_) & (!g95) & (!sk[25]) & (g346) & (!g351)) + ((i_11_) & (!g95) & (sk[25]) & (!g346) & (g351)));
	assign g383 = (((i_40_) & (!g45) & (!g333) & (!sk[26]) & (!g381) & (!g382)) + ((!i_40_) & (g45) & (!g333) & (!sk[26]) & (!g381) & (!g382)) + ((i_40_) & (!g45) & (!g333) & (!sk[26]) & (g381) & (!g382)) + ((i_40_) & (!g45) & (!g333) & (!sk[26]) & (!g381) & (g382)) + ((i_40_) & (g45) & (g333) & (!sk[26]) & (!g381) & (!g382)));
	assign g384 = (((!sk[27]) & (!i_40_) & (g105) & (!g8)) + ((sk[27]) & (!i_40_) & (!g105) & (!g8)) + ((!sk[27]) & (i_40_) & (!g105) & (g8)));
	assign g385 = (((i_11_) & (!sk[28]) & (i_12_)) + ((!i_11_) & (!sk[28]) & (i_12_)));
	assign g386 = (((i_36_) & (!sk[29]) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (!sk[29]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (!sk[29]) & (i_37_) & (!i_38_) & (!i_39_) & (i_40_)) + ((!i_36_) & (sk[29]) & (!i_37_) & (!i_38_) & (i_39_) & (i_40_)));
	assign g387 = (((g54) & (!g155) & (!sk[30]) & (!g385) & (!g246) & (!g386)) + ((!g54) & (g155) & (!sk[30]) & (!g385) & (!g246) & (!g386)) + ((g54) & (!g155) & (!sk[30]) & (!g385) & (!g246) & (g386)) + ((!g54) & (g155) & (!sk[30]) & (!g385) & (g246) & (!g386)));
	assign g388 = (((g102) & (!i_31_) & (!sk[31]) & (!g288) & (!g384) & (!g387)) + ((!g102) & (i_31_) & (!sk[31]) & (!g288) & (!g384) & (!g387)) + ((g102) & (!i_31_) & (!sk[31]) & (!g288) & (!g384) & (g387)) + ((g102) & (!i_31_) & (!sk[31]) & (g288) & (!g384) & (!g387)));
	assign g389 = (((i_22_) & (!i_24_) & (!sk[32]) & (!i_23_) & (!g182) & (!g325)) + ((!i_22_) & (i_24_) & (!sk[32]) & (!i_23_) & (!g182) & (!g325)) + ((i_22_) & (i_24_) & (!sk[32]) & (i_23_) & (g182) & (g325)));
	assign g390 = (((!i_22_) & (!sk[33]) & (g23) & (!i_21_)) + ((i_22_) & (!sk[33]) & (!g23) & (i_21_)) + ((i_22_) & (!sk[33]) & (g23) & (i_21_)));
	assign g391 = (((!sk[34]) & (!i_37_) & (g5) & (!g6) & (!g77)) + ((!sk[34]) & (!i_37_) & (!g5) & (g6) & (!g77)) + ((!sk[34]) & (!i_37_) & (g5) & (g6) & (g77)));
	assign g392 = (((i_32_) & (!g28) & (!g10) & (!i_24_) & (!sk[35]) & (!i_23_)) + ((!i_32_) & (g28) & (!g10) & (!i_24_) & (!sk[35]) & (!i_23_)) + ((!i_32_) & (g28) & (!g10) & (i_24_) & (!sk[35]) & (i_23_)));
	assign g393 = (((!i_38_) & (g5) & (!sk[36]) & (!g6)) + ((!i_38_) & (g5) & (!sk[36]) & (g6)) + ((i_38_) & (!g5) & (!sk[36]) & (g6)));
	assign g394 = (((i_36_) & (!i_37_) & (!i_39_) & (!i_40_) & (!g7) & (g393)) + ((!i_36_) & (!i_37_) & (i_39_) & (!i_40_) & (g7) & (!g393)) + ((!i_36_) & (i_37_) & (i_39_) & (!i_40_) & (!g7) & (g393)));
	assign g395 = (((!sk[38]) & (!i_37_) & (g14) & (!g5)) + ((!sk[38]) & (i_37_) & (!g14) & (g5)) + ((!sk[38]) & (!i_37_) & (g14) & (g5)));
	assign g396 = (((i_24_) & (!g123) & (!g144) & (!g199) & (!sk[39]) & (!g395)) + ((!i_24_) & (g123) & (!g144) & (!g199) & (!sk[39]) & (!g395)) + ((!i_24_) & (g123) & (!g144) & (!g199) & (!sk[39]) & (g395)) + ((i_24_) & (!g123) & (g144) & (g199) & (!sk[39]) & (!g395)));
	assign g397 = (((g390) & (!g391) & (!g392) & (!g394) & (!sk[40]) & (!g396)) + ((!g390) & (g391) & (!g392) & (!g394) & (!sk[40]) & (!g396)) + ((!g390) & (!g391) & (!g392) & (!g394) & (sk[40]) & (!g396)) + ((!g390) & (!g391) & (!g392) & (!g394) & (sk[40]) & (!g396)));
	assign g398 = (((!i_37_) & (i_38_) & (!sk[41]) & (!i_39_) & (!i_40_)) + ((!i_37_) & (!i_38_) & (!sk[41]) & (i_39_) & (!i_40_)) + ((!i_37_) & (i_38_) & (!sk[41]) & (!i_39_) & (i_40_)) + ((!i_37_) & (i_38_) & (!sk[41]) & (i_39_) & (!i_40_)) + ((i_37_) & (i_38_) & (!sk[41]) & (!i_39_) & (!i_40_)));
	assign g399 = (((!g101) & (g45) & (!sk[42]) & (!g49)) + ((g101) & (!g45) & (!sk[42]) & (g49)) + ((g101) & (g45) & (!sk[42]) & (!g49)));
	assign g400 = (((!i_32_) & (!sk[43]) & (g54) & (!i_13_) & (!g399)) + ((!i_32_) & (!sk[43]) & (!g54) & (i_13_) & (!g399)) + ((!i_32_) & (!sk[43]) & (g54) & (!i_13_) & (g399)));
	assign g401 = (((i_37_) & (!i_38_) & (!i_39_) & (!sk[44]) & (!i_40_) & (!g51)) + ((!i_37_) & (i_38_) & (!i_39_) & (!sk[44]) & (!i_40_) & (!g51)) + ((i_37_) & (!i_38_) & (!i_39_) & (!sk[44]) & (!i_40_) & (g51)) + ((!i_37_) & (!i_38_) & (!i_39_) & (sk[44]) & (i_40_) & (g51)) + ((!i_37_) & (!i_38_) & (i_39_) & (sk[44]) & (!i_40_) & (g51)) + ((!i_37_) & (!i_38_) & (i_39_) & (sk[44]) & (i_40_) & (g51)));
	assign g402 = (((!i_40_) & (g55) & (!g148) & (!g8) & (g189) & (!g401)) + ((!i_40_) & (g55) & (!g148) & (!g8) & (!g189) & (g401)) + ((!i_40_) & (!g55) & (g148) & (g8) & (!g189) & (!g401)));
	assign g403 = (((!sk[46]) & (!i_15_) & (g138) & (!g155) & (!g246)) + ((!sk[46]) & (!i_15_) & (!g138) & (g155) & (!g246)) + ((!sk[46]) & (!i_15_) & (g138) & (g155) & (g246)));
	assign g404 = (((i_37_) & (!g122) & (!g57) & (!g76) & (!sk[47]) & (!g5)) + ((!i_37_) & (g122) & (!g57) & (!g76) & (!sk[47]) & (!g5)) + ((!i_37_) & (!g122) & (g57) & (g76) & (sk[47]) & (g5)));
	assign g405 = (((g1) & (!g22) & (!i_9_) & (!sk[48]) & (!i_18_) & (!i_21_)) + ((!g1) & (g22) & (!i_9_) & (!sk[48]) & (!i_18_) & (!i_21_)) + ((!g1) & (!g22) & (i_9_) & (sk[48]) & (!i_18_) & (!i_21_)) + ((!g1) & (!g22) & (!i_9_) & (sk[48]) & (i_18_) & (!i_21_)) + ((!g1) & (!g22) & (!i_9_) & (sk[48]) & (!i_18_) & (i_21_)));
	assign g406 = (((!i_37_) & (i_38_) & (!i_40_) & (!sk[49]) & (!i_15_)) + ((!i_37_) & (!i_38_) & (i_40_) & (!sk[49]) & (!i_15_)) + ((!i_37_) & (i_38_) & (i_40_) & (!sk[49]) & (i_15_)));
	assign g407 = (((i_22_) & (!i_24_) & (!g125) & (!sk[50]) & (!g405) & (!g406)) + ((!i_22_) & (i_24_) & (!g125) & (!sk[50]) & (!g405) & (!g406)) + ((i_22_) & (i_24_) & (g125) & (!sk[50]) & (g405) & (g406)));
	assign g408 = (((!g47) & (g48) & (!sk[51]) & (!g49)) + ((g47) & (!g48) & (!sk[51]) & (g49)) + ((g47) & (g48) & (!sk[51]) & (!g49)));
	assign g409 = (((i_36_) & (!sk[52]) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (!sk[52]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (!sk[52]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (sk[52]) & (!i_37_) & (!i_38_) & (!i_39_) & (i_40_)) + ((!i_36_) & (sk[52]) & (!i_37_) & (!i_38_) & (i_39_) & (!i_40_)) + ((!i_36_) & (sk[52]) & (!i_37_) & (!i_38_) & (i_39_) & (i_40_)) + ((!i_36_) & (sk[52]) & (!i_37_) & (i_38_) & (!i_39_) & (!i_40_)));
	assign g410 = (((!g58) & (!sk[53]) & (g165) & (!g408) & (!g409)) + ((!g58) & (!sk[53]) & (!g165) & (g408) & (!g409)) + ((!g58) & (!sk[53]) & (g165) & (g408) & (!g409)) + ((g58) & (sk[53]) & (!g165) & (!g408) & (g409)));
	assign g411 = (((!i_40_) & (!g28) & (g128) & (g199) & (!g225) & (!g333)) + ((!i_40_) & (g28) & (!g128) & (!g199) & (!g225) & (g333)) + ((!i_40_) & (!g28) & (!g128) & (!g199) & (g225) & (g333)));
	assign g412 = (((g403) & (!sk[55]) & (!g404) & (!g407) & (!g410) & (!g411)) + ((!g403) & (!sk[55]) & (g404) & (!g407) & (!g410) & (!g411)) + ((!g403) & (sk[55]) & (!g404) & (!g407) & (!g410) & (!g411)));
	assign g413 = (((g93) & (!g398) & (!g400) & (!g402) & (!sk[56]) & (!g412)) + ((!g93) & (g398) & (!g400) & (!g402) & (!sk[56]) & (!g412)) + ((!g93) & (!g398) & (!g400) & (!g402) & (sk[56]) & (g412)) + ((!g93) & (!g398) & (!g400) & (!g402) & (sk[56]) & (g412)));
	assign g414 = (((!i_15_) & (g31) & (!sk[57]) & (!g124)) + ((!i_15_) & (g31) & (!sk[57]) & (g124)) + ((i_15_) & (!g31) & (!sk[57]) & (g124)));
	assign g415 = (((!sk[58]) & (!g131) & (g219) & (!g390)) + ((!sk[58]) & (g131) & (!g219) & (g390)) + ((!sk[58]) & (g131) & (g219) & (g390)));
	assign g416 = (((g1) & (!g138) & (!i_30_) & (!sk[59]) & (!i_29_) & (!g384)) + ((!g1) & (g138) & (!i_30_) & (!sk[59]) & (!i_29_) & (!g384)) + ((!g1) & (g138) & (!i_30_) & (!sk[59]) & (i_29_) & (!g384)));
	assign g417 = (((!i_36_) & (!i_37_) & (i_38_) & (i_39_) & (!i_40_) & (g5)) + ((!i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (g5)) + ((!i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (g5)));
	assign g418 = (((!sk[61]) & (!g94) & (g315) & (!g301) & (!g417)) + ((!sk[61]) & (!g94) & (!g315) & (g301) & (!g417)) + ((!sk[61]) & (!g94) & (!g315) & (g301) & (g417)) + ((!sk[61]) & (!g94) & (g315) & (g301) & (!g417)));
	assign g419 = (((i_37_) & (!g30) & (!g121) & (!sk[62]) & (!g123) & (!g418)) + ((!i_37_) & (g30) & (!g121) & (!sk[62]) & (!g123) & (!g418)) + ((!i_37_) & (g30) & (!g121) & (!sk[62]) & (!g123) & (!g418)) + ((!i_37_) & (!g30) & (!g121) & (sk[62]) & (!g123) & (!g418)) + ((!i_37_) & (!g30) & (!g121) & (sk[62]) & (!g123) & (!g418)) + ((!i_37_) & (!g30) & (!g121) & (sk[62]) & (!g123) & (!g418)));
	assign g420 = (((!g73) & (!g304) & (!g414) & (!g415) & (!g416) & (g419)) + ((!g73) & (!g304) & (!g414) & (!g415) & (!g416) & (g419)));
	assign g421 = (((!g383) & (!g388) & (!g389) & (g397) & (g413) & (g420)));
	assign g422 = (((!sk[65]) & (!i_11_) & (i_12_) & (!g103)) + ((!sk[65]) & (i_11_) & (!i_12_) & (g103)) + ((!sk[65]) & (!i_11_) & (i_12_) & (g103)));
	assign g423 = (((g65) & (!i_22_) & (!i_24_) & (!i_21_) & (!sk[66]) & (!g198)) + ((!g65) & (i_22_) & (!i_24_) & (!i_21_) & (!sk[66]) & (!g198)) + ((g65) & (i_22_) & (i_24_) & (i_21_) & (!sk[66]) & (g198)));
	assign g424 = (((!g151) & (g79) & (!g187) & (!sk[67]) & (!g423)) + ((!g151) & (!g79) & (g187) & (!sk[67]) & (!g423)) + ((g151) & (g79) & (!g187) & (!sk[67]) & (g423)) + ((g151) & (!g79) & (g187) & (!sk[67]) & (g423)));
	assign g425 = (((!sk[68]) & (i_5_) & (!i_9_) & (!g18) & (!i_18_) & (!i_19_)) + ((!sk[68]) & (!i_5_) & (i_9_) & (!g18) & (!i_18_) & (!i_19_)) + ((!sk[68]) & (!i_5_) & (i_9_) & (g18) & (!i_18_) & (!i_19_)) + ((sk[68]) & (!i_5_) & (!i_9_) & (g18) & (i_18_) & (i_19_)));
	assign g426 = (((!sk[69]) & (!i_24_) & (i_18_) & (!i_23_) & (!i_19_)) + ((!sk[69]) & (!i_24_) & (!i_18_) & (i_23_) & (!i_19_)) + ((!sk[69]) & (i_24_) & (i_18_) & (i_23_) & (!i_19_)) + ((!sk[69]) & (i_24_) & (!i_18_) & (i_23_) & (i_19_)));
	assign g427 = (((g112) & (i_24_) & (g125) & (i_21_) & (i_23_) & (g198)));
	assign g428 = (((!sk[71]) & (!i_32_) & (i_21_) & (!g198) & (!g376)) + ((!sk[71]) & (!i_32_) & (!i_21_) & (g198) & (!g376)) + ((!sk[71]) & (!i_32_) & (i_21_) & (g198) & (g376)));
	assign g429 = (((g157) & (!sk[72]) & (!g425) & (!g426) & (!g427) & (!g428)) + ((!g157) & (!sk[72]) & (g425) & (!g426) & (!g427) & (!g428)) + ((!g157) & (sk[72]) & (!g425) & (!g426) & (!g427) & (!g428)) + ((!g157) & (sk[72]) & (!g425) & (!g426) & (!g427) & (!g428)) + ((!g157) & (!sk[72]) & (g425) & (!g426) & (!g427) & (!g428)));
	assign g430 = (((i_5_) & (!g45) & (!g115) & (!sk[73]) & (!i_28_) & (!g336)) + ((!i_5_) & (g45) & (!g115) & (!sk[73]) & (!i_28_) & (!g336)) + ((!i_5_) & (g45) & (g115) & (!sk[73]) & (!i_28_) & (g336)));
	assign g431 = (((!i_5_) & (g77) & (!g273) & (!sk[74]) & (!g350)) + ((!i_5_) & (!g77) & (g273) & (!sk[74]) & (!g350)) + ((!i_5_) & (g77) & (g273) & (!sk[74]) & (g350)));
	assign g432 = (((!sk[75]) & (!g139) & (g83)) + ((!sk[75]) & (g139) & (g83)));
	assign g433 = (((!g136) & (!sk[76]) & (g131) & (!g104) & (!g338)) + ((!g136) & (!sk[76]) & (!g131) & (g104) & (!g338)) + ((!g136) & (sk[76]) & (!g131) & (!g104) & (!g338)) + ((!g136) & (sk[76]) & (!g131) & (!g104) & (!g338)));
	assign g434 = (((!g197) & (g423) & (!sk[77]) & (!g432) & (!g433)) + ((!g197) & (g423) & (!sk[77]) & (g432) & (!g433)) + ((!g197) & (!g423) & (!sk[77]) & (g432) & (!g433)) + ((g197) & (!g423) & (sk[77]) & (!g432) & (!g433)));
	assign g435 = (((i_22_) & (!g429) & (!sk[78]) & (!g430) & (!g431) & (!g434)) + ((!i_22_) & (g429) & (!sk[78]) & (!g430) & (!g431) & (!g434)) + ((!i_22_) & (g429) & (!sk[78]) & (!g430) & (!g431) & (!g434)) + ((!i_22_) & (!g429) & (sk[78]) & (!g430) & (!g431) & (!g434)));
	assign g436 = (((!i_22_) & (!sk[79]) & (i_24_) & (!g222)) + ((i_22_) & (!sk[79]) & (!i_24_) & (g222)) + ((i_22_) & (!sk[79]) & (i_24_) & (g222)));
	assign g437 = (((i_38_) & (!i_39_) & (!sk[80]) & (!i_40_) & (!g65) & (!g88)) + ((!i_38_) & (i_39_) & (!sk[80]) & (!i_40_) & (!g65) & (!g88)) + ((i_38_) & (!i_39_) & (!sk[80]) & (i_40_) & (g65) & (g88)) + ((i_38_) & (i_39_) & (!sk[80]) & (!i_40_) & (g65) & (g88)));
	assign g438 = (((g65) & (!g151) & (!g79) & (!g436) & (!sk[81]) & (!g437)) + ((!g65) & (g151) & (!g79) & (!g436) & (!sk[81]) & (!g437)) + ((!g65) & (!g151) & (!g79) & (!g436) & (sk[81]) & (!g437)) + ((!g65) & (!g151) & (!g79) & (!g436) & (sk[81]) & (!g437)) + ((!g65) & (!g151) & (!g79) & (!g436) & (sk[81]) & (!g437)) + ((!g65) & (!g151) & (!g79) & (!g436) & (sk[81]) & (!g437)));
	assign g439 = (((g422) & (!g424) & (!g208) & (!g435) & (!sk[82]) & (!g438)) + ((!g422) & (g424) & (!g208) & (!g435) & (!sk[82]) & (!g438)) + ((!g422) & (!g424) & (g208) & (g435) & (sk[82]) & (g438)));
	assign g440 = (((!g77) & (g184) & (!g219) & (!sk[83]) & (!g422)) + ((!g77) & (!g184) & (g219) & (!sk[83]) & (!g422)) + ((!g77) & (g184) & (!g219) & (!sk[83]) & (!g422)) + ((!g77) & (g184) & (!g219) & (!sk[83]) & (!g422)));
	assign g441 = (((!g84) & (g213) & (!sk[84]) & (!g208) & (!g430)) + ((!g84) & (!g213) & (!sk[84]) & (g208) & (!g430)) + ((!g84) & (!g213) & (!sk[84]) & (g208) & (!g430)) + ((!g84) & (!g213) & (!sk[84]) & (g208) & (!g430)));
	assign g442 = (((!i_36_) & (!sk[85]) & (g100) & (!g73)) + ((i_36_) & (!sk[85]) & (!g100) & (g73)) + ((!i_36_) & (!sk[85]) & (g100) & (g73)));
	assign g443 = (((g10) & (!g45) & (!g76) & (!g165) & (!sk[86]) & (!g442)) + ((!g10) & (g45) & (!g76) & (!g165) & (!sk[86]) & (!g442)) + ((!g10) & (g45) & (g76) & (!g165) & (!sk[86]) & (!g442)) + ((!g10) & (!g45) & (!g76) & (g165) & (sk[86]) & (!g442)) + ((!g10) & (!g45) & (!g76) & (!g165) & (sk[86]) & (g442)));
	assign g444 = (((g11) & (!g43) & (!i_25_) & (!i_20_) & (!sk[87]) & (!g443)) + ((!g11) & (g43) & (!i_25_) & (!i_20_) & (!sk[87]) & (!g443)) + ((g11) & (g43) & (i_25_) & (!i_20_) & (!sk[87]) & (g443)) + ((g11) & (g43) & (!i_25_) & (i_20_) & (!sk[87]) & (g443)));
	assign g445 = (((!i_24_) & (g152) & (!g132) & (!sk[88]) & (!i_23_)) + ((!i_24_) & (!g152) & (g132) & (!sk[88]) & (!i_23_)) + ((!i_24_) & (!g152) & (!g132) & (sk[88]) & (!i_23_)) + ((!i_24_) & (!g152) & (!g132) & (sk[88]) & (!i_23_)));
	assign g446 = (((!i_40_) & (!sk[89]) & (g95) & (!g98) & (!g215)) + ((!i_40_) & (!sk[89]) & (!g95) & (g98) & (!g215)) + ((!i_40_) & (!sk[89]) & (g95) & (!g98) & (g215)) + ((i_40_) & (!sk[89]) & (g95) & (g98) & (!g215)));
	assign g447 = (((!sk[90]) & (i_25_) & (!g390) & (!i_20_) & (!g445) & (!g446)) + ((!sk[90]) & (!i_25_) & (g390) & (!i_20_) & (!g445) & (!g446)) + ((sk[90]) & (!i_25_) & (!g390) & (!i_20_) & (!g445) & (!g446)) + ((!sk[90]) & (!i_25_) & (g390) & (!i_20_) & (g445) & (!g446)) + ((!sk[90]) & (!i_25_) & (g390) & (!i_20_) & (!g445) & (!g446)));
	assign o_10_ = (((i_22_) & (!i_24_) & (!i_21_) & (!g444) & (!sk[91]) & (!g447)) + ((!i_22_) & (i_24_) & (!i_21_) & (!g444) & (!sk[91]) & (!g447)) + ((!i_22_) & (!i_24_) & (!i_21_) & (!g444) & (sk[91]) & (!g447)) + ((i_22_) & (i_24_) & (i_21_) & (g444) & (!sk[91]) & (!g447)));
	assign g449 = (((!sk[92]) & (i_31_) & (!g1) & (!g105) & (!g106) & (!g273)) + ((!sk[92]) & (!i_31_) & (g1) & (!g105) & (!g106) & (!g273)) + ((sk[92]) & (!i_31_) & (!g1) & (g105) & (g106) & (g273)));
	assign g450 = (((g56) & (!sk[93]) & (g46) & (!g165)) + ((!g56) & (!sk[93]) & (g46) & (!g165)) + ((g56) & (!sk[93]) & (!g46) & (g165)));
	assign g451 = (((i_11_) & (!i_31_) & (!i_12_) & (!sk[94]) & (!g11) & (!g450)) + ((!i_11_) & (i_31_) & (!i_12_) & (!sk[94]) & (!g11) & (!g450)) + ((i_11_) & (!i_31_) & (!i_12_) & (!sk[94]) & (g11) & (g450)) + ((!i_11_) & (!i_31_) & (i_12_) & (sk[94]) & (g11) & (g450)));
	assign g452 = (((g1) & (!i_16_) & (!i_17_) & (!i_9_) & (!sk[95]) & (!g451)) + ((!g1) & (i_16_) & (!i_17_) & (!i_9_) & (!sk[95]) & (!g451)) + ((!g1) & (i_16_) & (i_17_) & (!i_9_) & (!sk[95]) & (g451)) + ((!g1) & (i_16_) & (!i_17_) & (i_9_) & (!sk[95]) & (g451)) + ((!g1) & (!i_16_) & (i_17_) & (i_9_) & (sk[95]) & (g451)));
	assign g453 = (((!g95) & (!g99) & (!g215) & (!g292) & (!g449) & (!g452)) + ((!g95) & (!g99) & (!g215) & (!g292) & (!g449) & (!g452)));
	assign g454 = (((!sk[97]) & (!i_7_) & (i_5_) & (!i_0_)) + ((!sk[97]) & (i_7_) & (!i_5_) & (i_0_)) + ((!sk[97]) & (!i_7_) & (i_5_) & (!i_0_)));
	assign g455 = (((!sk[98]) & (i_37_) & (!i_38_) & (!i_40_) & (!g160) & (!g94)) + ((!sk[98]) & (!i_37_) & (i_38_) & (!i_40_) & (!g160) & (!g94)) + ((!sk[98]) & (i_37_) & (i_38_) & (!i_40_) & (g160) & (!g94)) + ((sk[98]) & (!i_37_) & (!i_38_) & (!i_40_) & (!g160) & (!g94)));
	assign o_12_ = (((!g122) & (g454) & (!sk[99]) & (!i_8_) & (!g455)) + ((!g122) & (!g454) & (!sk[99]) & (i_8_) & (!g455)) + ((!g122) & (g454) & (!sk[99]) & (i_8_) & (g455)));
	assign g457 = (((!i_38_) & (!i_39_) & (!i_40_) & (!g65) & (!g151) & (g184)) + ((!i_38_) & (!i_39_) & (!i_40_) & (!g65) & (!g151) & (g184)) + ((i_38_) & (i_39_) & (!i_40_) & (!g65) & (!g151) & (g184)) + ((!i_38_) & (!i_39_) & (i_40_) & (!g65) & (!g151) & (g184)) + ((!i_38_) & (!i_39_) & (!i_40_) & (!g65) & (!g151) & (g184)));
	assign g458 = (((!g14) & (g65) & (!sk[101]) & (!g88) & (!g457)) + ((!g14) & (!g65) & (!sk[101]) & (g88) & (!g457)) + ((!g14) & (!g65) & (sk[101]) & (!g88) & (g457)) + ((!g14) & (!g65) & (sk[101]) & (!g88) & (g457)) + ((!g14) & (!g65) & (sk[101]) & (!g88) & (g457)));
	assign g459 = (((!i_13_) & (!sk[102]) & (g226) & (!g457)) + ((!i_13_) & (sk[102]) & (!g226) & (g457)) + ((i_13_) & (!sk[102]) & (!g226) & (g457)));
	assign g460 = (((!sk[103]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (!g95)) + ((!sk[103]) & (!i_37_) & (i_38_) & (!i_39_) & (!i_40_) & (!g95)) + ((!sk[103]) & (i_37_) & (i_38_) & (i_39_) & (!i_40_) & (g95)));
	assign g461 = (((!i_2_) & (i_1_) & (!sk[104]) & (!i_0_)) + ((i_2_) & (!i_1_) & (!sk[104]) & (i_0_)) + ((!i_2_) & (!i_1_) & (sk[104]) & (i_0_)));
	assign g462 = (((!i_3_) & (i_4_) & (!sk[105]) & (!g461)) + ((i_3_) & (!i_4_) & (!sk[105]) & (g461)) + ((!i_3_) & (!i_4_) & (sk[105]) & (g461)));
	assign g463 = (((i_37_) & (!sk[106]) & (!g104) & (!g78) & (!g79) & (!g462)) + ((!i_37_) & (!sk[106]) & (g104) & (!g78) & (!g79) & (!g462)) + ((i_37_) & (!sk[106]) & (g104) & (g78) & (!g79) & (g462)) + ((!i_37_) & (sk[106]) & (!g104) & (g78) & (g79) & (g462)));
	assign g464 = (((g30) & (!g22) & (!sk[107]) & (!g70) & (!g71) & (!g463)) + ((!g30) & (g22) & (!sk[107]) & (!g70) & (!g71) & (!g463)) + ((!g30) & (!g22) & (sk[107]) & (g70) & (!g71) & (g463)) + ((!g30) & (g22) & (!sk[107]) & (g70) & (g71) & (!g463)));
	assign g465 = (((!i_2_) & (i_1_) & (!sk[108]) & (!i_0_)) + ((!i_2_) & (i_1_) & (!sk[108]) & (i_0_)) + ((i_2_) & (!i_1_) & (!sk[108]) & (i_0_)));
	assign g466 = (((!sk[109]) & (!i_7_) & (g67) & (!g465)) + ((!sk[109]) & (i_7_) & (!g67) & (g465)) + ((!sk[109]) & (!i_7_) & (g67) & (g465)));
	assign g467 = (((i_36_) & (!i_40_) & (!i_34_) & (!i_35_) & (!sk[110]) & (!g6)) + ((!i_36_) & (i_40_) & (!i_34_) & (!i_35_) & (!sk[110]) & (!g6)) + ((!i_36_) & (i_40_) & (!i_34_) & (i_35_) & (!sk[110]) & (g6)) + ((i_36_) & (!i_40_) & (!i_34_) & (!i_35_) & (!sk[110]) & (g6)));
	assign g468 = (((g66) & (!g187) & (!sk[111]) & (!g346) & (!g466) & (!g467)) + ((!g66) & (g187) & (!sk[111]) & (!g346) & (!g466) & (!g467)) + ((g66) & (g187) & (!sk[111]) & (!g346) & (g466) & (!g467)) + ((!g66) & (!g187) & (sk[111]) & (g346) & (!g466) & (g467)));
	assign g469 = (((g148) & (!sk[112]) & (!g225) & (!g460) & (!g464) & (!g468)) + ((!g148) & (!sk[112]) & (g225) & (!g460) & (!g464) & (!g468)) + ((!g148) & (sk[112]) & (!g225) & (!g460) & (!g464) & (!g468)) + ((!g148) & (sk[112]) & (!g225) & (!g460) & (!g464) & (!g468)));
	assign g470 = (((!i_37_) & (!sk[113]) & (i_38_) & (!i_39_) & (!g51)) + ((!i_37_) & (!sk[113]) & (!i_38_) & (i_39_) & (!g51)) + ((i_37_) & (!sk[113]) & (i_38_) & (i_39_) & (g51)));
	assign g471 = (((i_38_) & (!g51) & (!g115) & (!sk[114]) & (!g232) & (!g470)) + ((!i_38_) & (g51) & (!g115) & (!sk[114]) & (!g232) & (!g470)) + ((!i_38_) & (!g51) & (!g115) & (sk[114]) & (g232) & (g470)) + ((i_38_) & (g51) & (g115) & (!sk[114]) & (g232) & (!g470)));
	assign g472 = (((i_37_) & (!i_38_) & (!i_39_) & (!g51) & (!sk[115]) & (!i_17_)) + ((!i_37_) & (i_38_) & (!i_39_) & (!g51) & (!sk[115]) & (!i_17_)) + ((!i_37_) & (i_38_) & (i_39_) & (g51) & (!sk[115]) & (!i_17_)) + ((i_37_) & (!i_38_) & (!i_39_) & (g51) & (!sk[115]) & (!i_17_)));
	assign g473 = (((i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (!sk[116]) & (!g51)) + ((!i_37_) & (i_38_) & (!i_39_) & (!i_40_) & (!sk[116]) & (!g51)) + ((!i_37_) & (i_38_) & (i_39_) & (!i_40_) & (!sk[116]) & (g51)) + ((i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (!sk[116]) & (g51)) + ((!i_37_) & (i_38_) & (!i_39_) & (!i_40_) & (!sk[116]) & (g51)) + ((!i_37_) & (!i_38_) & (i_39_) & (!i_40_) & (sk[116]) & (g51)) + ((!i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (sk[116]) & (g51)));
	assign g474 = (((!sk[117]) & (i_16_) & (!g269) & (!g471) & (!g472) & (!g473)) + ((!sk[117]) & (!i_16_) & (g269) & (!g471) & (!g472) & (!g473)) + ((sk[117]) & (!i_16_) & (!g269) & (!g471) & (!g472) & (!g473)) + ((!sk[117]) & (i_16_) & (!g269) & (!g471) & (!g472) & (!g473)) + ((!sk[117]) & (!i_16_) & (g269) & (!g471) & (!g472) & (!g473)));
	assign g475 = (((i_36_) & (i_37_) & (!i_38_) & (!g67) & (g241) & (!g251)) + ((!i_36_) & (!i_37_) & (!i_38_) & (g67) & (!g241) & (g251)));
	assign g476 = (((!i_40_) & (i_32_) & (!sk[119]) & (!g475)) + ((i_40_) & (!i_32_) & (!sk[119]) & (g475)) + ((!i_40_) & (!i_32_) & (sk[119]) & (g475)));
	assign g477 = (((!sk[120]) & (!g94) & (g267) & (!g315)) + ((!sk[120]) & (g94) & (!g267) & (g315)) + ((!sk[120]) & (!g94) & (g267) & (g315)));
	assign g478 = (((!sk[121]) & (!g168) & (g136) & (!g79)) + ((sk[121]) & (!g168) & (!g136) & (!g79)) + ((!sk[121]) & (g168) & (!g136) & (g79)) + ((!sk[121]) & (!g168) & (g136) & (!g79)));
	assign g479 = (((g53) & (!g24) & (!g198) & (!sk[122]) & (!g477) & (!g478)) + ((!g53) & (g24) & (!g198) & (!sk[122]) & (!g477) & (!g478)) + ((!g53) & (!g24) & (g198) & (sk[122]) & (g477) & (!g478)) + ((g53) & (g24) & (g198) & (!sk[122]) & (!g477) & (!g478)));
	assign g480 = (((!g139) & (g225) & (!sk[123]) & (!g272)) + ((g139) & (!g225) & (!sk[123]) & (g272)) + ((!g139) & (g225) & (!sk[123]) & (g272)));
	assign g481 = (((!i_40_) & (!sk[124]) & (g121) & (!i_23_) & (!g198)) + ((!i_40_) & (!sk[124]) & (!g121) & (i_23_) & (!g198)) + ((!i_40_) & (!sk[124]) & (g121) & (!i_23_) & (g198)));
	assign g482 = (((g122) & (!g112) & (!g47) & (!g94) & (!sk[125]) & (!g481)) + ((!g122) & (g112) & (!g47) & (!g94) & (!sk[125]) & (!g481)) + ((!g122) & (g112) & (!g47) & (!g94) & (!sk[125]) & (g481)) + ((!g122) & (g112) & (!g47) & (!g94) & (!sk[125]) & (!g481)));
	assign g483 = (((g56) & (!i_32_) & (!i_31_) & (i_30_) & (!i_28_) & (i_29_)) + ((g56) & (!i_32_) & (!i_31_) & (!i_30_) & (i_28_) & (!i_29_)));
	assign g484 = (((i_5_) & (!sk[127]) & (!g45) & (!g115) & (!g105) & (!g483)) + ((!i_5_) & (!sk[127]) & (g45) & (!g115) & (!g105) & (!g483)) + ((!i_5_) & (!sk[127]) & (g45) & (g115) & (!g105) & (g483)) + ((!i_5_) & (sk[127]) & (!g45) & (!g115) & (g105) & (g483)));
	assign g485 = (((!i_32_) & (g47) & (!sk[0]) & (!i_0_)) + ((i_32_) & (!g47) & (!sk[0]) & (i_0_)) + ((!i_32_) & (!g47) & (sk[0]) & (i_0_)));
	assign g486 = (((i_36_) & (!sk[1]) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (!sk[1]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((i_36_) & (!sk[1]) & (!i_37_) & (i_38_) & (i_39_) & (i_40_)) + ((i_36_) & (!sk[1]) & (i_37_) & (i_38_) & (!i_39_) & (i_40_)));
	assign g487 = (((!sk[2]) & (g56) & (!g118) & (!g66) & (!g485) & (!g486)) + ((!sk[2]) & (!g56) & (g118) & (!g66) & (!g485) & (!g486)) + ((!sk[2]) & (!g56) & (g118) & (g66) & (!g485) & (!g486)) + ((!sk[2]) & (g56) & (!g118) & (!g66) & (g485) & (g486)));
	assign g488 = (((i_40_) & (!g220) & (!g225) & (!g243) & (!sk[3]) & (!g487)) + ((!i_40_) & (g220) & (!g225) & (!g243) & (!sk[3]) & (!g487)) + ((i_40_) & (g220) & (!g225) & (!g243) & (!sk[3]) & (!g487)) + ((!i_40_) & (g220) & (!g225) & (!g243) & (!sk[3]) & (!g487)) + ((!i_40_) & (!g220) & (!g225) & (!g243) & (sk[3]) & (!g487)));
	assign g489 = (((!sk[4]) & (g479) & (!g480) & (!g482) & (!g484) & (!g488)) + ((!sk[4]) & (!g479) & (g480) & (!g482) & (!g484) & (!g488)) + ((sk[4]) & (!g479) & (!g480) & (!g482) & (!g484) & (g488)));
	assign o_17_ = (((!sk[5]) & (!g53) & (g474) & (!g476) & (!g285) & (!g489)) + ((!sk[5]) & (g53) & (!g474) & (!g476) & (!g285) & (!g489)) + ((sk[5]) & (!g53) & (!g474) & (g476) & (!g285) & (!g489)) + ((sk[5]) & (!g53) & (!g474) & (!g476) & (!g285) & (!g489)) + ((sk[5]) & (!g53) & (!g474) & (!g476) & (!g285) & (!g489)));
	assign g491 = (((!i_37_) & (!sk[6]) & (i_38_) & (!i_31_) & (!g1)) + ((!i_37_) & (!sk[6]) & (!i_38_) & (i_31_) & (!g1)) + ((i_37_) & (!sk[6]) & (i_38_) & (!i_31_) & (!g1)) + ((!i_37_) & (sk[6]) & (!i_38_) & (!i_31_) & (!g1)));
	assign g492 = (((i_36_) & (!g56) & (!sk[7]) & (!g353) & (!g466) & (!g491)) + ((!i_36_) & (g56) & (!sk[7]) & (!g353) & (!g466) & (!g491)) + ((!i_36_) & (!g56) & (sk[7]) & (g353) & (g466) & (!g491)) + ((!i_36_) & (g56) & (!sk[7]) & (!g353) & (!g466) & (g491)));
	assign g493 = (((!sk[8]) & (!g24) & (i_9_)) + ((!sk[8]) & (!g24) & (i_9_)));
	assign g494 = (((!sk[9]) & (i_11_) & (!i_12_) & (!i_15_) & (!g171) & (!g493)) + ((!sk[9]) & (!i_11_) & (i_12_) & (!i_15_) & (!g171) & (!g493)) + ((!sk[9]) & (i_11_) & (i_12_) & (i_15_) & (g171) & (!g493)) + ((!sk[9]) & (i_11_) & (i_12_) & (i_15_) & (!g171) & (g493)));
	assign g495 = (((i_7_) & (!g162) & (!i_14_) & (!g478) & (!sk[10]) & (!g494)) + ((!i_7_) & (g162) & (!i_14_) & (!g478) & (!sk[10]) & (!g494)) + ((!i_7_) & (!g162) & (i_14_) & (!g478) & (sk[10]) & (g494)));
	assign g496 = (((i_36_) & (!sk[11]) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (!sk[11]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (sk[11]) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (!sk[11]) & (i_37_) & (!i_38_) & (i_39_) & (i_40_)) + ((!i_36_) & (sk[11]) & (!i_37_) & (i_38_) & (!i_39_) & (!i_40_)));
	assign g497 = (((!sk[12]) & (!i_31_) & (g1) & (!i_16_) & (!i_9_)) + ((!sk[12]) & (!i_31_) & (!g1) & (i_16_) & (!i_9_)) + ((!sk[12]) & (!i_31_) & (!g1) & (i_16_) & (!i_9_)) + ((sk[12]) & (!i_31_) & (!g1) & (!i_16_) & (i_9_)));
	assign g498 = (((!sk[13]) & (!g56) & (g18) & (!g496) & (!g497)) + ((!sk[13]) & (!g56) & (!g18) & (g496) & (!g497)) + ((!sk[13]) & (g56) & (g18) & (g496) & (g497)));
	assign g499 = (((i_40_) & (!g95) & (!sk[14]) & (!g104) & (!g347) & (!g462)) + ((!i_40_) & (g95) & (!sk[14]) & (!g104) & (!g347) & (!g462)) + ((!i_40_) & (g95) & (!sk[14]) & (g104) & (!g347) & (!g462)) + ((i_40_) & (!g95) & (!sk[14]) & (!g104) & (g347) & (g462)));
	assign g500 = (((!sk[15]) & (g5) & (!g116) & (!g92) & (!g71) & (!g187)) + ((!sk[15]) & (!g5) & (g116) & (!g92) & (!g71) & (!g187)) + ((!sk[15]) & (g5) & (g116) & (g92) & (!g71) & (!g187)) + ((sk[15]) & (!g5) & (!g116) & (!g92) & (g71) & (g187)));
	assign g501 = (((!g116) & (g6) & (!sk[16]) & (!g467) & (!g500)) + ((g116) & (!g6) & (!sk[16]) & (g467) & (!g500)) + ((!g116) & (!g6) & (!sk[16]) & (g467) & (!g500)) + ((!g116) & (g6) & (!sk[16]) & (!g467) & (g500)));
	assign g502 = (((i_37_) & (!i_38_) & (!i_39_) & (!sk[17]) & (!i_40_) & (!g148)) + ((!i_37_) & (i_38_) & (!i_39_) & (!sk[17]) & (!i_40_) & (!g148)) + ((i_37_) & (!i_38_) & (i_39_) & (!sk[17]) & (!i_40_) & (g148)) + ((!i_37_) & (i_38_) & (i_39_) & (!sk[17]) & (!i_40_) & (g148)) + ((!i_37_) & (!i_38_) & (!i_39_) & (sk[17]) & (i_40_) & (g148)) + ((!i_37_) & (!i_38_) & (!i_39_) & (sk[17]) & (i_40_) & (g148)));
	assign g503 = (((!sk[18]) & (!i_7_) & (i_33_) & (!i_32_) & (!g2)) + ((!sk[18]) & (!i_7_) & (!i_33_) & (i_32_) & (!g2)) + ((!sk[18]) & (!i_7_) & (i_33_) & (i_32_) & (g2)));
	assign g504 = (((i_37_) & (!g76) & (!sk[19]) & (!g5) & (!g301) & (!g503)) + ((!i_37_) & (g76) & (!sk[19]) & (!g5) & (!g301) & (!g503)) + ((i_37_) & (!g76) & (!sk[19]) & (!g5) & (!g301) & (!g503)) + ((!i_37_) & (!g76) & (sk[19]) & (!g5) & (!g301) & (!g503)) + ((!i_37_) & (!g76) & (sk[19]) & (!g5) & (!g301) & (!g503)) + ((!i_37_) & (!g76) & (sk[19]) & (!g5) & (!g301) & (!g503)));
	assign g505 = (((i_37_) & (!i_38_) & (i_39_) & (!i_40_) & (g95) & (!g333)) + ((!i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (!g95) & (g333)) + ((!i_37_) & (!i_38_) & (i_39_) & (i_40_) & (g95) & (!g333)));
	assign g506 = (((!sk[21]) & (!i_33_) & (i_31_) & (!g2)) + ((!sk[21]) & (i_33_) & (!i_31_) & (g2)));
	assign g507 = (((i_40_) & (!g77) & (!g8) & (!sk[22]) & (!g289) & (!g506)) + ((!i_40_) & (g77) & (!g8) & (!sk[22]) & (!g289) & (!g506)) + ((!i_40_) & (g77) & (!g8) & (!sk[22]) & (!g289) & (g506)) + ((!i_40_) & (!g77) & (g8) & (sk[22]) & (!g289) & (g506)));
	assign g508 = (((!sk[23]) & (g117) & (!g502) & (!g504) & (!g505) & (!g507)) + ((!sk[23]) & (!g117) & (g502) & (!g504) & (!g505) & (!g507)) + ((sk[23]) & (!g117) & (!g502) & (g504) & (!g505) & (!g507)));
	assign g509 = (((g495) & (!sk[24]) & (!g498) & (!g499) & (!g501) & (!g508)) + ((!g495) & (!sk[24]) & (g498) & (!g499) & (!g501) & (!g508)) + ((!g495) & (sk[24]) & (!g498) & (!g499) & (!g501) & (g508)));
	assign g510 = (((!i_37_) & (i_39_) & (!sk[25]) & (!g118) & (!g96)) + ((!i_37_) & (!i_39_) & (!sk[25]) & (g118) & (!g96)) + ((!i_37_) & (!i_39_) & (!sk[25]) & (g118) & (g96)) + ((!i_37_) & (!i_39_) & (sk[25]) & (!g118) & (g96)));
	assign g511 = (((i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (g123) & (!g6)) + ((!i_37_) & (i_38_) & (!i_39_) & (i_40_) & (g123) & (!g6)) + ((i_37_) & (i_38_) & (!i_39_) & (!i_40_) & (!g123) & (g6)) + ((i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (!g123) & (g6)));
	assign g512 = (((!i_7_) & (!i_11_) & (!i_38_) & (i_40_) & (!i_10_) & (!i_27_)) + ((!i_7_) & (!i_11_) & (i_38_) & (!i_40_) & (!i_10_) & (!i_27_)) + ((!i_7_) & (!i_11_) & (i_38_) & (!i_40_) & (!i_10_) & (!i_27_)));
	assign g513 = (((!i_37_) & (!sk[28]) & (i_38_) & (!i_39_) & (!i_40_)) + ((!i_37_) & (!sk[28]) & (!i_38_) & (i_39_) & (!i_40_)) + ((i_37_) & (!sk[28]) & (!i_38_) & (i_39_) & (i_40_)) + ((!i_37_) & (sk[28]) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_37_) & (sk[28]) & (!i_38_) & (!i_39_) & (i_40_)));
	assign g514 = (((i_36_) & (!g102) & (!g408) & (!g512) & (!sk[29]) & (!g513)) + ((!i_36_) & (g102) & (!g408) & (!g512) & (!sk[29]) & (!g513)) + ((i_36_) & (g102) & (!g408) & (g512) & (!sk[29]) & (!g513)) + ((!i_36_) & (!g102) & (g408) & (!g512) & (sk[29]) & (!g513)));
	assign g515 = (((i_38_) & (!i_40_) & (!g51) & (!sk[30]) & (!i_15_) & (!g385)) + ((!i_38_) & (i_40_) & (!g51) & (!sk[30]) & (!i_15_) & (!g385)) + ((i_38_) & (!i_40_) & (g51) & (!sk[30]) & (i_15_) & (g385)));
	assign g516 = (((!g162) & (i_31_) & (!sk[31]) & (!g155)) + ((g162) & (!i_31_) & (!sk[31]) & (g155)) + ((!g162) & (!i_31_) & (sk[31]) & (g155)));
	assign g517 = (((g135) & (!g390) & (!g470) & (!g515) & (!sk[32]) & (!g516)) + ((!g135) & (g390) & (!g470) & (!g515) & (!sk[32]) & (!g516)) + ((!g135) & (!g390) & (!g470) & (!g515) & (sk[32]) & (!g516)) + ((!g135) & (!g390) & (!g470) & (!g515) & (sk[32]) & (!g516)) + ((!g135) & (!g390) & (!g470) & (!g515) & (sk[32]) & (!g516)) + ((!g135) & (!g390) & (!g470) & (!g515) & (sk[32]) & (!g516)));
	assign g518 = (((g121) & (!g510) & (!g511) & (!sk[33]) & (!g514) & (!g517)) + ((!g121) & (g510) & (!g511) & (!sk[33]) & (!g514) & (!g517)) + ((!g121) & (!g510) & (!g511) & (sk[33]) & (!g514) & (g517)) + ((!g121) & (!g510) & (!g511) & (sk[33]) & (!g514) & (g517)));
	assign g519 = (((g73) & (!sk[34]) & (!g492) & (!g397) & (!g509) & (!g518)) + ((!g73) & (!sk[34]) & (g492) & (!g397) & (!g509) & (!g518)) + ((!g73) & (sk[34]) & (!g492) & (g397) & (g509) & (g518)) + ((!g73) & (sk[34]) & (!g492) & (g397) & (g509) & (g518)));
	assign g520 = (((!sk[35]) & (!i_7_) & (g67) & (!g461)) + ((!sk[35]) & (i_7_) & (!g67) & (g461)) + ((!sk[35]) & (!i_7_) & (g67) & (g461)));
	assign g521 = (((i_38_) & (!g101) & (!g197) & (!g136) & (g66) & (g520)) + ((!i_38_) & (!g101) & (g197) & (g136) & (!g66) & (g520)));
	assign g522 = (((!sk[37]) & (!g45) & (g73) & (!g408)) + ((!sk[37]) & (g45) & (!g73) & (g408)) + ((!sk[37]) & (g45) & (g73) & (g408)));
	assign g523 = (((!i_38_) & (i_39_) & (!i_40_) & (!sk[38]) & (!g121)) + ((!i_38_) & (!i_39_) & (i_40_) & (!sk[38]) & (!g121)) + ((!i_38_) & (i_39_) & (i_40_) & (!sk[38]) & (g121)) + ((i_38_) & (!i_39_) & (!i_40_) & (sk[38]) & (g121)));
	assign g524 = (((!sk[39]) & (i_40_) & (!g21) & (!g7) & (!g148) & (!g8)) + ((!sk[39]) & (!i_40_) & (g21) & (!g7) & (!g148) & (!g8)) + ((!sk[39]) & (!i_40_) & (g21) & (!g7) & (g148) & (!g8)) + ((!sk[39]) & (i_40_) & (!g21) & (g7) & (!g148) & (g8)));
	assign g525 = (((i_37_) & (!g6) & (!sk[40]) & (!g522) & (!g523) & (!g524)) + ((!i_37_) & (g6) & (!sk[40]) & (!g522) & (!g523) & (!g524)) + ((i_37_) & (!g6) & (!sk[40]) & (!g522) & (!g523) & (!g524)) + ((!i_37_) & (!g6) & (sk[40]) & (!g522) & (!g523) & (!g524)) + ((!i_37_) & (!g6) & (sk[40]) & (!g522) & (!g523) & (!g524)));
	assign g526 = (((g48) & (!i_6_) & (!g712) & (!g521) & (!sk[41]) & (!g525)) + ((!g48) & (i_6_) & (!g712) & (!g521) & (!sk[41]) & (!g525)) + ((!g48) & (!i_6_) & (!g712) & (!g521) & (sk[41]) & (g525)) + ((!g48) & (!i_6_) & (!g712) & (!g521) & (sk[41]) & (g525)) + ((!g48) & (!i_6_) & (g712) & (!g521) & (sk[41]) & (g525)));
	assign g527 = (((g122) & (!g2) & (!g21) & (!g24) & (!sk[42]) & (!g112)) + ((!g122) & (g2) & (!g21) & (!g24) & (!sk[42]) & (!g112)) + ((!g122) & (g2) & (g21) & (!g24) & (!sk[42]) & (!g112)) + ((!g122) & (g2) & (!g21) & (!g24) & (!sk[42]) & (g112)));
	assign g528 = (((g65) & (!i_9_) & (!g260) & (!sk[43]) & (!g136) & (!g527)) + ((!g65) & (i_9_) & (!g260) & (!sk[43]) & (!g136) & (!g527)) + ((!g65) & (i_9_) & (!g260) & (!sk[43]) & (!g136) & (g527)) + ((g65) & (i_9_) & (g260) & (!sk[43]) & (g136) & (!g527)));
	assign g529 = (((!sk[44]) & (i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!sk[44]) & (!i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!sk[44]) & (i_36_) & (i_37_) & (i_38_) & (!i_39_) & (i_40_)) + ((sk[44]) & (!i_36_) & (!i_37_) & (i_38_) & (i_39_) & (!i_40_)));
	assign g530 = (((!i_37_) & (i_35_) & (!sk[45]) & (!i_13_)) + ((i_37_) & (!i_35_) & (!sk[45]) & (i_13_)) + ((!i_37_) & (i_35_) & (!sk[45]) & (!i_13_)));
	assign g531 = (((!i_36_) & (!i_38_) & (!i_39_) & (i_40_) & (!g136) & (!g530)) + ((!i_36_) & (!i_38_) & (i_39_) & (!i_40_) & (g136) & (!g530)));
	assign g532 = (((!g168) & (!g151) & (!g187) & (!g189) & (!g165) & (!g531)) + ((!g168) & (!g151) & (!g187) & (!g189) & (!g165) & (!g531)));
	assign g533 = (((g65) & (!sk[48]) & (!g22) & (!g454) & (!g529) & (!g532)) + ((!g65) & (!sk[48]) & (g22) & (!g454) & (!g529) & (!g532)) + ((g65) & (!sk[48]) & (!g22) & (g454) & (g529) & (!g532)) + ((g65) & (!sk[48]) & (g22) & (!g454) & (!g529) & (!g532)));
	assign g534 = (((!g122) & (g2) & (!sk[49]) & (!g21) & (!g113)) + ((!g122) & (!g2) & (!sk[49]) & (g21) & (!g113)) + ((!g122) & (g2) & (!sk[49]) & (g21) & (!g113)) + ((!g122) & (g2) & (!sk[49]) & (!g21) & (g113)));
	assign g535 = (((!sk[50]) & (g171) & (!g493) & (!i_14_) & (!g385) & (!g534)) + ((!sk[50]) & (!g171) & (g493) & (!i_14_) & (!g385) & (!g534)) + ((!sk[50]) & (g171) & (!g493) & (!i_14_) & (!g385) & (g534)) + ((!sk[50]) & (!g171) & (g493) & (!i_14_) & (!g385) & (g534)) + ((!sk[50]) & (g171) & (!g493) & (!i_14_) & (!g385) & (g534)));
	assign g536 = (((i_12_) & (!g196) & (!sk[51]) & (!g528) & (!g533) & (!g535)) + ((!i_12_) & (g196) & (!sk[51]) & (!g528) & (!g533) & (!g535)) + ((i_12_) & (!g196) & (!sk[51]) & (!g528) & (!g533) & (!g535)) + ((!i_12_) & (!g196) & (sk[51]) & (!g528) & (!g533) & (!g535)));
	assign g537 = (((!sk[52]) & (!g28) & (g10) & (!g255) & (!g315)) + ((!sk[52]) & (!g28) & (!g10) & (g255) & (!g315)) + ((sk[52]) & (g28) & (!g10) & (!g255) & (!g315)) + ((sk[52]) & (!g28) & (!g10) & (!g255) & (g315)));
	assign g538 = (((i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (!sk[53]) & (!i_40_)) + ((!i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (!sk[53]) & (!i_40_)) + ((!i_36_) & (!i_37_) & (!i_38_) & (i_39_) & (sk[53]) & (!i_40_)) + ((!i_36_) & (!i_37_) & (i_38_) & (!i_39_) & (sk[53]) & (!i_40_)) + ((!i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (sk[53]) & (i_40_)));
	assign g539 = (((g162) & (!i_35_) & (!g46) & (!g442) & (!sk[54]) & (!g538)) + ((!g162) & (i_35_) & (!g46) & (!g442) & (!sk[54]) & (!g538)) + ((!g162) & (i_35_) & (!g46) & (g442) & (!sk[54]) & (!g538)) + ((!g162) & (!i_35_) & (g46) & (!g442) & (sk[54]) & (!g538)) + ((!g162) & (!i_35_) & (!g46) & (!g442) & (sk[54]) & (g538)));
	assign g540 = (((!i_37_) & (i_38_) & (!i_39_) & (!sk[55]) & (!i_40_)) + ((!i_37_) & (!i_38_) & (i_39_) & (!sk[55]) & (!i_40_)) + ((!i_37_) & (i_38_) & (i_39_) & (!sk[55]) & (i_40_)) + ((i_37_) & (!i_38_) & (!i_39_) & (sk[55]) & (i_40_)));
	assign g541 = (((!sk[56]) & (!i_13_) & (g28) & (!i_9_) & (!g129)) + ((!sk[56]) & (!i_13_) & (!g28) & (i_9_) & (!g129)) + ((!sk[56]) & (!i_13_) & (g28) & (i_9_) & (!g129)) + ((sk[56]) & (i_13_) & (!g28) & (!i_9_) & (g129)));
	assign g542 = (((!sk[57]) & (i_36_) & (!g162) & (!g70) & (!g540) & (!g541)) + ((!sk[57]) & (!i_36_) & (g162) & (!g70) & (!g540) & (!g541)) + ((sk[57]) & (!i_36_) & (!g162) & (g70) & (!g540) & (g541)) + ((sk[57]) & (!i_36_) & (!g162) & (!g70) & (g540) & (!g541)));
	assign g543 = (((!sk[58]) & (i_15_) & (!g48) & (!g537) & (!g539) & (!g542)) + ((!sk[58]) & (!i_15_) & (g48) & (!g537) & (!g539) & (!g542)) + ((!sk[58]) & (!i_15_) & (g48) & (g537) & (!g539) & (!g542)) + ((!sk[58]) & (!i_15_) & (g48) & (!g537) & (g539) & (!g542)) + ((!sk[58]) & (!i_15_) & (g48) & (!g537) & (!g539) & (g542)));
	assign g544 = (((i_37_) & (!sk[59]) & (!i_40_) & (!g162) & (!i_35_) & (!g281)) + ((!i_37_) & (!sk[59]) & (i_40_) & (!g162) & (!i_35_) & (!g281)) + ((!i_37_) & (sk[59]) & (!i_40_) & (!g162) & (!i_35_) & (g281)) + ((!i_37_) & (!sk[59]) & (i_40_) & (!g162) & (i_35_) & (g281)));
	assign g545 = (((!i_36_) & (!i_37_) & (i_38_) & (!g101) & (!g106) & (g66)) + ((!i_36_) & (!i_37_) & (!i_38_) & (!g101) & (g106) & (!g66)));
	assign g546 = (((!sk[61]) & (g65) & (!g71) & (!g79) & (!g454) & (!g545)) + ((!sk[61]) & (!g65) & (g71) & (!g79) & (!g454) & (!g545)) + ((sk[61]) & (!g65) & (!g71) & (!g79) & (g454) & (g545)) + ((!sk[61]) & (g65) & (g71) & (g79) & (g454) & (!g545)));
	assign g547 = (((i_5_) & (!sk[62]) & (!g48) & (!g537) & (!g544) & (!g546)) + ((!i_5_) & (!sk[62]) & (g48) & (!g537) & (!g544) & (!g546)) + ((!i_5_) & (sk[62]) & (!g48) & (!g537) & (!g544) & (!g546)) + ((!i_5_) & (sk[62]) & (!g48) & (!g537) & (!g544) & (!g546)) + ((!i_5_) & (!sk[62]) & (g48) & (!g537) & (!g544) & (!g546)));
	assign g548 = (((!sk[63]) & (i_7_) & (!g122) & (!i_5_) & (!g2) & (!g195)) + ((!sk[63]) & (!i_7_) & (g122) & (!i_5_) & (!g2) & (!g195)) + ((sk[63]) & (!i_7_) & (!g122) & (i_5_) & (g2) & (g195)));
	assign g549 = (((i_36_) & (!g162) & (!i_5_) & (!g61) & (!sk[64]) & (!g48)) + ((!i_36_) & (g162) & (!i_5_) & (!g61) & (!sk[64]) & (!g48)) + ((!i_36_) & (!g162) & (i_5_) & (g61) & (sk[64]) & (g48)));
	assign g550 = (((i_37_) & (!sk[65]) & (!i_38_) & (!i_39_) & (!i_40_) & (!i_31_)) + ((!i_37_) & (!sk[65]) & (i_38_) & (!i_39_) & (!i_40_) & (!i_31_)) + ((i_37_) & (!sk[65]) & (!i_38_) & (!i_39_) & (!i_40_) & (!i_31_)) + ((!i_37_) & (!sk[65]) & (i_38_) & (i_39_) & (i_40_) & (!i_31_)) + ((!i_37_) & (!sk[65]) & (i_38_) & (i_39_) & (!i_40_) & (!i_31_)));
	assign g551 = (((i_31_) & (!i_5_) & (!g293) & (!sk[66]) & (!g549) & (!g550)) + ((!i_31_) & (i_5_) & (!g293) & (!sk[66]) & (!g549) & (!g550)) + ((!i_31_) & (!i_5_) & (!g293) & (sk[66]) & (!g549) & (!g550)) + ((!i_31_) & (!i_5_) & (!g293) & (sk[66]) & (!g549) & (!g550)) + ((!i_31_) & (!i_5_) & (!g293) & (sk[66]) & (!g549) & (g550)));
	assign g552 = (((i_7_) & (!sk[67]) & (!g22) & (!g181) & (!g548) & (!g551)) + ((!i_7_) & (!sk[67]) & (g22) & (!g181) & (!g548) & (!g551)) + ((i_7_) & (!sk[67]) & (!g22) & (!g181) & (!g548) & (g551)) + ((!i_7_) & (sk[67]) & (!g22) & (!g181) & (!g548) & (g551)) + ((!i_7_) & (!sk[67]) & (g22) & (g181) & (!g548) & (g551)));
	assign g553 = (((i_7_) & (!i_11_) & (!sk[68]) & (!g103) & (!g528) & (!g552)) + ((!i_7_) & (i_11_) & (!sk[68]) & (!g103) & (!g528) & (!g552)) + ((i_7_) & (!i_11_) & (!sk[68]) & (!g103) & (!g528) & (g552)) + ((!i_7_) & (i_11_) & (!sk[68]) & (!g103) & (!g528) & (g552)) + ((!i_7_) & (!i_11_) & (sk[68]) & (!g103) & (!g528) & (g552)));
	assign g554 = (((i_7_) & (!g536) & (!sk[69]) & (!g543) & (!g547) & (!g553)) + ((!i_7_) & (g536) & (!sk[69]) & (!g543) & (!g547) & (!g553)) + ((i_7_) & (!g536) & (!sk[69]) & (!g543) & (g547) & (g553)) + ((!i_7_) & (g536) & (!sk[69]) & (!g543) & (g547) & (g553)));
	assign g555 = (((i_36_) & (!i_38_) & (!i_39_) & (i_40_) & (!g88) & (!i_6_)) + ((i_36_) & (i_38_) & (i_39_) & (i_40_) & (g88) & (!i_6_)));
	assign g556 = (((!sk[71]) & (i_36_) & (!i_37_) & (!i_0_) & (!g187) & (!g555)) + ((!sk[71]) & (!i_36_) & (i_37_) & (!i_0_) & (!g187) & (!g555)) + ((sk[71]) & (!i_36_) & (!i_37_) & (!i_0_) & (!g187) & (!g555)) + ((sk[71]) & (!i_36_) & (!i_37_) & (!i_0_) & (!g187) & (!g555)) + ((!sk[71]) & (!i_36_) & (i_37_) & (i_0_) & (!g187) & (!g555)) + ((!sk[71]) & (!i_36_) & (i_37_) & (!i_0_) & (!g187) & (!g555)));
	assign g557 = (((!i_36_) & (!sk[72]) & (i_37_) & (!g5) & (!g79)) + ((!i_36_) & (!sk[72]) & (!i_37_) & (g5) & (!g79)) + ((!i_36_) & (!sk[72]) & (!i_37_) & (g5) & (g79)) + ((i_36_) & (!sk[72]) & (i_37_) & (g5) & (!g79)));
	assign g558 = (((!i_36_) & (g100) & (!sk[73]) & (!i_35_) & (!g73)) + ((!i_36_) & (!g100) & (!sk[73]) & (i_35_) & (!g73)) + ((i_36_) & (g100) & (!sk[73]) & (!i_35_) & (g73)));
	assign g559 = (((!sk[74]) & (i_37_) & (!i_34_) & (!g51) & (!g79) & (!i_6_)) + ((!sk[74]) & (!i_37_) & (i_34_) & (!g51) & (!g79) & (!i_6_)) + ((!sk[74]) & (i_37_) & (i_34_) & (g51) & (g79) & (!i_6_)));
	assign g560 = (((i_34_) & (!i_32_) & (!g51) & (!sk[75]) & (!g558) & (!g559)) + ((!i_34_) & (i_32_) & (!g51) & (!sk[75]) & (!g558) & (!g559)) + ((!i_34_) & (!i_32_) & (!g51) & (sk[75]) & (!g558) & (!g559)) + ((i_34_) & (!i_32_) & (!g51) & (!sk[75]) & (!g558) & (!g559)) + ((!i_34_) & (!i_32_) & (g51) & (sk[75]) & (!g558) & (!g559)));
	assign g561 = (((!sk[76]) & (!i_34_) & (g113) & (!g78)) + ((!sk[76]) & (i_34_) & (!g113) & (g78)) + ((!sk[76]) & (!i_34_) & (g113) & (g78)));
	assign g562 = (((!i_37_) & (i_38_) & (!g101) & (!g160) & (!g94) & (!g318)) + ((i_37_) & (!i_38_) & (!g101) & (!g160) & (!g94) & (!g318)) + ((!i_37_) & (!i_38_) & (g101) & (!g160) & (!g94) & (!g318)) + ((!i_37_) & (i_38_) & (!g101) & (!g160) & (!g94) & (!g318)) + ((!i_37_) & (!i_38_) & (!g101) & (!g160) & (g94) & (!g318)));
	assign g563 = (((i_36_) & (!i_37_) & (!sk[78]) & (!i_34_) & (!g77) & (!g562)) + ((!i_36_) & (i_37_) & (!sk[78]) & (!i_34_) & (!g77) & (!g562)) + ((!i_36_) & (!i_37_) & (sk[78]) & (!i_34_) & (!g77) & (g562)) + ((!i_36_) & (!i_37_) & (sk[78]) & (!i_34_) & (!g77) & (g562)) + ((!i_36_) & (!i_37_) & (sk[78]) & (i_34_) & (!g77) & (g562)) + ((!i_36_) & (!i_37_) & (sk[78]) & (!i_34_) & (!g77) & (g562)));
	assign g564 = (((i_33_) & (g1) & (!i_0_) & (!sk[79]) & (!g561) & (!g563)) + ((i_33_) & (!g1) & (i_0_) & (!sk[79]) & (!g561) & (!g563)) + ((i_33_) & (!g1) & (!i_0_) & (!sk[79]) & (!g561) & (!g563)) + ((!i_33_) & (g1) & (!i_0_) & (!sk[79]) & (!g561) & (!g563)) + ((i_33_) & (!g1) & (!i_0_) & (!sk[79]) & (!g561) & (g563)));
	assign g565 = (((i_7_) & (!g556) & (!g557) & (!sk[80]) & (!g560) & (!g564)) + ((!i_7_) & (g556) & (!g557) & (!sk[80]) & (!g560) & (!g564)) + ((i_7_) & (!g556) & (!g557) & (!sk[80]) & (!g560) & (g564)) + ((!i_7_) & (g556) & (!g557) & (!sk[80]) & (g560) & (g564)) + ((!i_7_) & (!g556) & (!g557) & (sk[80]) & (g560) & (g564)));
	assign g566 = (((!i_37_) & (i_40_) & (!i_31_) & (!sk[81]) & (!i_9_)) + ((!i_37_) & (!i_40_) & (i_31_) & (!sk[81]) & (!i_9_)) + ((!i_37_) & (!i_40_) & (!i_31_) & (sk[81]) & (i_9_)));
	assign g567 = (((!i_11_) & (!i_5_) & (!i_12_) & (!i_15_) & (!i_14_) & (!g566)) + ((!i_11_) & (!i_5_) & (!i_12_) & (!i_15_) & (!i_14_) & (!g566)) + ((!i_11_) & (!i_5_) & (!i_12_) & (!i_15_) & (!i_14_) & (!g566)) + ((!i_11_) & (!i_5_) & (!i_12_) & (!i_15_) & (!i_14_) & (!g566)) + ((i_11_) & (!i_5_) & (i_12_) & (i_15_) & (i_14_) & (!g566)));
	assign g568 = (((!i_37_) & (!sk[83]) & (i_38_) & (!i_39_) & (!i_40_)) + ((!i_37_) & (!sk[83]) & (!i_38_) & (i_39_) & (!i_40_)) + ((!i_37_) & (sk[83]) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_37_) & (!sk[83]) & (i_38_) & (i_39_) & (i_40_)));
	assign g569 = (((!i_16_) & (!sk[84]) & (i_17_) & (!i_9_) & (!g568)) + ((!i_16_) & (!sk[84]) & (!i_17_) & (i_9_) & (!g568)) + ((i_16_) & (!sk[84]) & (i_17_) & (!i_9_) & (g568)) + ((i_16_) & (!sk[84]) & (!i_17_) & (i_9_) & (g568)) + ((!i_16_) & (!sk[84]) & (i_17_) & (i_9_) & (g568)));
	assign g570 = (((!i_33_) & (!sk[85]) & (i_5_) & (!g2) & (!g569)) + ((!i_33_) & (!sk[85]) & (!i_5_) & (g2) & (!g569)) + ((i_33_) & (!sk[85]) & (i_5_) & (g2) & (!g569)));
	assign g571 = (((!i_16_) & (!sk[86]) & (i_9_) & (!g18)) + ((i_16_) & (!sk[86]) & (!i_9_) & (g18)) + ((!i_16_) & (!sk[86]) & (i_9_) & (g18)));
	assign g572 = (((!i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (g506) & (g571)) + ((i_37_) & (i_38_) & (!i_39_) & (!i_40_) & (g506) & (!g571)) + ((!i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (g506) & (!g571)) + ((!i_37_) & (!i_38_) & (i_39_) & (i_40_) & (g506) & (g571)) + ((!i_37_) & (i_38_) & (!i_39_) & (!i_40_) & (g506) & (g571)));
	assign g573 = (((i_36_) & (!g56) & (!sk[88]) & (!g567) & (!g570) & (!g572)) + ((!i_36_) & (g56) & (!sk[88]) & (!g567) & (!g570) & (!g572)) + ((i_36_) & (!g56) & (!sk[88]) & (!g567) & (!g570) & (!g572)) + ((!i_36_) & (!g56) & (sk[88]) & (!g567) & (!g570) & (!g572)) + ((!i_36_) & (!g56) & (sk[88]) & (g567) & (!g570) & (!g572)));
	assign g574 = (((i_39_) & (!i_40_) & (i_35_) & (g65) & (g116) & (g454)) + ((!i_39_) & (i_40_) & (!i_35_) & (g65) & (g116) & (g454)));
	assign o_22_ = (((i_7_) & (!sk[90]) & (!g573) & (!g503) & (!g547) & (!g574)) + ((!i_7_) & (!sk[90]) & (g573) & (!g503) & (!g547) & (!g574)) + ((!i_7_) & (sk[90]) & (!g573) & (!g503) & (!g547) & (!g574)) + ((!i_7_) & (sk[90]) & (!g573) & (g503) & (!g547) & (!g574)) + ((!i_7_) & (sk[90]) & (!g573) & (!g503) & (!g547) & (!g574)) + ((!i_7_) & (sk[90]) & (!g573) & (!g503) & (!g547) & (g574)));
	assign g576 = (((!sk[91]) & (!i_36_) & (g100) & (!g106) & (!g73)) + ((!sk[91]) & (!i_36_) & (!g100) & (g106) & (!g73)) + ((!sk[91]) & (i_36_) & (g100) & (g106) & (g73)));
	assign g577 = (((i_38_) & (!i_39_) & (!sk[92]) & (!g122) & (!g136) & (!g385)) + ((!i_38_) & (i_39_) & (!sk[92]) & (!g122) & (!g136) & (!g385)) + ((i_38_) & (i_39_) & (!sk[92]) & (!g122) & (g136) & (!g385)));
	assign g578 = (((!sk[93]) & (i_37_) & (!g122) & (!g5) & (!i_0_) & (!g69)) + ((!sk[93]) & (!i_37_) & (g122) & (!g5) & (!i_0_) & (!g69)) + ((!sk[93]) & (i_37_) & (!g122) & (g5) & (i_0_) & (g69)));
	assign g579 = (((!i_38_) & (g73) & (!g219) & (!sk[94]) & (!g704)) + ((!i_38_) & (!g73) & (g219) & (!sk[94]) & (!g704)) + ((!i_38_) & (g73) & (!g219) & (!sk[94]) & (g704)) + ((!i_38_) & (!g73) & (!g219) & (sk[94]) & (g704)) + ((i_38_) & (!g73) & (!g219) & (sk[94]) & (g704)));
	assign g580 = (((i_37_) & (!i_38_) & (!g47) & (!g87) & (!sk[95]) & (!g130)) + ((!i_37_) & (i_38_) & (!g47) & (!g87) & (!sk[95]) & (!g130)) + ((i_37_) & (!i_38_) & (!g47) & (!g87) & (!sk[95]) & (g130)) + ((!i_37_) & (!i_38_) & (!g47) & (g87) & (sk[95]) & (g130)));
	assign g581 = (((i_31_) & (!g122) & (!i_5_) & (!sk[96]) & (!g2) & (!g580)) + ((!i_31_) & (g122) & (!i_5_) & (!sk[96]) & (!g2) & (!g580)) + ((!i_31_) & (g122) & (!i_5_) & (!sk[96]) & (!g2) & (!g580)) + ((!i_31_) & (!g122) & (!i_5_) & (sk[96]) & (!g2) & (!g580)) + ((!i_31_) & (!g122) & (!i_5_) & (sk[96]) & (!g2) & (!g580)));
	assign g582 = (((!i_34_) & (g30) & (!sk[97]) & (!i_15_) & (!g106)) + ((!i_34_) & (!g30) & (!sk[97]) & (i_15_) & (!g106)) + ((!i_34_) & (!g30) & (sk[97]) & (!i_15_) & (g106)));
	assign g583 = (((!sk[98]) & (i_40_) & (!g27) & (!g105) & (!g106) & (!g582)) + ((!sk[98]) & (!i_40_) & (g27) & (!g105) & (!g106) & (!g582)) + ((sk[98]) & (!i_40_) & (!g27) & (!g105) & (!g106) & (!g582)) + ((sk[98]) & (!i_40_) & (!g27) & (!g105) & (!g106) & (!g582)) + ((sk[98]) & (!i_40_) & (!g27) & (!g105) & (!g106) & (!g582)));
	assign g584 = (((!i_38_) & (g101) & (!g134) & (!sk[99]) & (!g152)) + ((!i_38_) & (!g101) & (g134) & (!sk[99]) & (!g152)) + ((i_38_) & (g101) & (!g134) & (!sk[99]) & (g152)) + ((!i_38_) & (!g101) & (!g134) & (sk[99]) & (g152)) + ((!i_38_) & (!g101) & (!g134) & (sk[99]) & (g152)));
	assign g585 = (((!sk[100]) & (i_38_) & (!i_39_) & (!g122) & (!i_15_) & (!g2)) + ((!sk[100]) & (!i_38_) & (i_39_) & (!g122) & (!i_15_) & (!g2)) + ((!sk[100]) & (i_38_) & (i_39_) & (!g122) & (!i_15_) & (g2)) + ((!sk[100]) & (!i_38_) & (i_39_) & (!g122) & (!i_15_) & (g2)));
	assign g586 = (((i_37_) & (!i_38_) & (!g134) & (!sk[101]) & (!g92) & (!g585)) + ((!i_37_) & (i_38_) & (!g134) & (!sk[101]) & (!g92) & (!g585)) + ((!i_37_) & (!i_38_) & (!g134) & (sk[101]) & (!g92) & (g585)) + ((!i_37_) & (!i_38_) & (g134) & (sk[101]) & (g92) & (!g585)));
	assign g587 = (((g184) & (!g581) & (!g583) & (!g584) & (!sk[102]) & (!g586)) + ((!g184) & (g581) & (!g583) & (!g584) & (!sk[102]) & (!g586)) + ((g184) & (g581) & (g583) & (g584) & (!sk[102]) & (!g586)));
	assign g588 = (((!g22) & (i_16_) & (!sk[103]) & (!i_9_) & (!g255)) + ((!g22) & (i_16_) & (!sk[103]) & (!i_9_) & (!g255)) + ((!g22) & (!i_16_) & (!sk[103]) & (i_9_) & (!g255)) + ((!g22) & (!i_16_) & (!sk[103]) & (i_9_) & (!g255)) + ((!g22) & (!i_16_) & (sk[103]) & (!i_9_) & (g255)));
	assign g589 = (((!i_37_) & (g51) & (!g122) & (!i_15_) & (!g5) & (!g87)) + ((i_37_) & (!g51) & (!g122) & (!i_15_) & (g5) & (g87)));
	assign g590 = (((i_34_) & (!i_5_) & (!i_0_) & (!g106) & (!g214) & (!g589)) + ((!i_34_) & (!i_5_) & (!i_0_) & (!g106) & (!g214) & (!g589)) + ((!i_34_) & (!i_5_) & (!i_0_) & (!g106) & (!g214) & (!g589)) + ((i_34_) & (!i_5_) & (!i_0_) & (!g106) & (!g214) & (!g589)) + ((!i_34_) & (!i_5_) & (!i_0_) & (!g106) & (!g214) & (!g589)) + ((!i_34_) & (!i_5_) & (!i_0_) & (!g106) & (!g214) & (!g589)));
	assign g591 = (((i_37_) & (!i_38_) & (!sk[106]) & (!i_39_) & (!i_40_) & (!g92)) + ((!i_37_) & (i_38_) & (!sk[106]) & (!i_39_) & (!i_40_) & (!g92)) + ((i_37_) & (i_38_) & (!sk[106]) & (!i_39_) & (!i_40_) & (g92)) + ((!i_37_) & (!i_38_) & (sk[106]) & (!i_39_) & (!i_40_) & (!g92)) + ((!i_37_) & (i_38_) & (!sk[106]) & (i_39_) & (!i_40_) & (!g92)) + ((i_37_) & (!i_38_) & (!sk[106]) & (i_39_) & (!i_40_) & (!g92)) + ((!i_37_) & (!i_38_) & (sk[106]) & (!i_39_) & (i_40_) & (!g92)));
	assign g592 = (((i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (i_35_)) + ((!i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (i_35_)) + ((!i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (i_35_)) + ((i_36_) & (i_37_) & (!i_38_) & (i_39_) & (!i_40_) & (!i_35_)) + ((i_36_) & (!i_37_) & (i_38_) & (!i_39_) & (!i_40_) & (!i_35_)) + ((!i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (!i_35_)) + ((i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (!i_35_)) + ((i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (!i_35_)) + ((!i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (!i_35_)));
	assign g593 = (((!i_38_) & (!i_39_) & (!i_40_) & (!g22) & (!i_16_) & (!i_9_)) + ((!i_38_) & (i_39_) & (!i_40_) & (g22) & (!i_16_) & (!i_9_)) + ((!i_38_) & (!i_39_) & (i_40_) & (g22) & (!i_16_) & (!i_9_)));
	assign g594 = (((i_36_) & (!sk[109]) & (!i_39_) & (!g102) & (!g30) & (!g593)) + ((!i_36_) & (!sk[109]) & (i_39_) & (!g102) & (!g30) & (!g593)) + ((!i_36_) & (!sk[109]) & (i_39_) & (g102) & (!g30) & (g593)) + ((!i_36_) & (sk[109]) & (!i_39_) & (g102) & (!g30) & (g593)));
	assign g595 = (((i_35_) & (!g65) & (!sk[110]) & (!g591) & (!g592) & (!g594)) + ((!i_35_) & (g65) & (!sk[110]) & (!g591) & (!g592) & (!g594)) + ((!i_35_) & (!g65) & (sk[110]) & (!g591) & (!g592) & (!g594)) + ((!i_35_) & (!g65) & (sk[110]) & (!g591) & (!g592) & (!g594)) + ((!i_35_) & (!g65) & (sk[110]) & (!g591) & (!g592) & (!g594)));
	assign g596 = (((i_38_) & (!i_9_) & (!sk[111]) & (!g585) & (!g693) & (!g595)) + ((!i_38_) & (i_9_) & (!sk[111]) & (!g585) & (!g693) & (!g595)) + ((!i_38_) & (i_9_) & (!sk[111]) & (!g585) & (!g693) & (g595)) + ((!i_38_) & (i_9_) & (!sk[111]) & (!g585) & (g693) & (g595)) + ((!i_38_) & (!i_9_) & (sk[111]) & (!g585) & (!g693) & (g595)) + ((!i_38_) & (!i_9_) & (sk[111]) & (!g585) & (g693) & (g595)));
	assign g597 = (((!g576) & (!g577) & (!g578) & (g579) & (g587) & (g596)));
	assign g598 = (((!g112) & (!sk[113]) & (g18) & (!g121) & (!g365)) + ((!g112) & (!sk[113]) & (!g18) & (g121) & (!g365)) + ((g112) & (!sk[113]) & (g18) & (g121) & (g365)));
	assign g599 = (((!sk[114]) & (!g23) & (g84) & (!i_21_) & (!i_23_)) + ((!sk[114]) & (!g23) & (!g84) & (i_21_) & (!i_23_)) + ((!sk[114]) & (g23) & (g84) & (!i_21_) & (!i_23_)));
	assign g600 = (((!sk[115]) & (!g43) & (g375) & (!g399)) + ((!sk[115]) & (g43) & (!g375) & (g399)) + ((!sk[115]) & (g43) & (g375) & (g399)));
	assign g601 = (((!g143) & (!sk[116]) & (g43) & (!i_23_) & (!g246)) + ((!g143) & (!sk[116]) & (!g43) & (i_23_) & (!g246)) + ((g143) & (!sk[116]) & (g43) & (!i_23_) & (g246)));
	assign g602 = (((i_36_) & (!sk[117]) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (!sk[117]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_)) + ((!i_36_) & (!sk[117]) & (i_37_) & (!i_38_) & (!i_39_) & (i_40_)) + ((!i_36_) & (sk[117]) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_40_)));
	assign g603 = (((i_11_) & (!g1) & (!i_12_) & (g28) & (g42) & (!g602)) + ((!i_11_) & (!g1) & (i_12_) & (g28) & (g42) & (!g602)) + ((i_11_) & (!g1) & (!i_12_) & (!g28) & (g42) & (g602)) + ((!i_11_) & (!g1) & (i_12_) & (!g28) & (g42) & (g602)));
	assign g604 = (((i_11_) & (!g1) & (!i_12_) & (g246) & (g355) & (!g442)) + ((!i_11_) & (!g1) & (i_12_) & (g246) & (g355) & (!g442)) + ((i_11_) & (!g1) & (!i_12_) & (!g246) & (g355) & (g442)) + ((!i_11_) & (!g1) & (i_12_) & (!g246) & (g355) & (g442)));
	assign g605 = (((g2) & (g21) & (g3) & (g23) & (g24) & (!g113)) + ((g2) & (!g21) & (g3) & (g23) & (g24) & (g113)));
	assign g606 = (((!g599) & (!g600) & (!g601) & (!g603) & (!g604) & (!g605)));
	assign g607 = (((!g124) & (!g367) & (g41) & (g20) & (!g598) & (g606)) + ((!g124) & (!g367) & (g41) & (g20) & (!g598) & (g606)));
	assign g608 = (((g53) & (!sk[123]) & (!g107) & (!g108) & (!g119) & (!g338)) + ((!g53) & (!sk[123]) & (g107) & (!g108) & (!g119) & (!g338)) + ((g53) & (!sk[123]) & (g107) & (!g108) & (g119) & (!g338)) + ((g53) & (!sk[123]) & (!g107) & (g108) & (g119) & (!g338)) + ((g53) & (!sk[123]) & (g107) & (!g108) & (!g119) & (g338)) + ((g53) & (!sk[123]) & (!g107) & (g108) & (!g119) & (g338)));
	assign g609 = (((!g197) & (g136) & (!g69) & (!sk[124]) & (!g330)) + ((!g197) & (!g136) & (g69) & (!sk[124]) & (!g330)) + ((g197) & (g136) & (g69) & (!sk[124]) & (g330)));
	assign g610 = (((!i_40_) & (!sk[125]) & (g121) & (!g6) & (!g346)) + ((i_40_) & (!sk[125]) & (!g121) & (g6) & (!g346)) + ((!i_40_) & (!sk[125]) & (!g121) & (g6) & (!g346)) + ((!i_40_) & (sk[125]) & (!g121) & (!g6) & (!g346)) + ((!i_40_) & (!sk[125]) & (!g121) & (g6) & (!g346)));
	assign g611 = (((!g331) & (!sk[126]) & (g609) & (!g50) & (!g610)) + ((!g331) & (!sk[126]) & (!g609) & (g50) & (!g610)) + ((!g331) & (sk[126]) & (!g609) & (!g50) & (g610)));
	assign g612 = (((!g14) & (!sk[127]) & (g134) & (!g330) & (!g611)) + ((!g14) & (!sk[127]) & (!g134) & (g330) & (!g611)) + ((!g14) & (sk[127]) & (!g134) & (!g330) & (g611)) + ((!g14) & (sk[127]) & (!g134) & (!g330) & (g611)) + ((!g14) & (sk[127]) & (!g134) & (!g330) & (g611)));
	assign g613 = (((g607) & (!sk[0]) & (!g305) & (!g608) & (!g82) & (!g612)) + ((!g607) & (!sk[0]) & (g305) & (!g608) & (!g82) & (!g612)) + ((g607) & (!sk[0]) & (!g305) & (!g608) & (g82) & (g612)));
	assign g614 = (((!g14) & (g197) & (!sk[1]) & (!g136) & (!g330)) + ((!g14) & (!g197) & (!sk[1]) & (g136) & (!g330)) + ((g14) & (g197) & (!sk[1]) & (g136) & (g330)));
	assign g615 = (((!g74) & (g331) & (!g609) & (!sk[2]) & (!g614)) + ((!g74) & (!g331) & (g609) & (!sk[2]) & (!g614)) + ((!g74) & (!g331) & (!g609) & (sk[2]) & (!g614)));
	assign g616 = (((!g607) & (g305) & (!sk[3]) & (!g608) & (!g615)) + ((!g607) & (!g305) & (!sk[3]) & (g608) & (!g615)) + ((g607) & (!g305) & (sk[3]) & (!g608) & (g615)));
	assign g617 = (((!g66) & (!g68) & (!g81) & (!g187) & (!g305) & (!g50)) + ((!g66) & (!g68) & (!g81) & (!g187) & (!g305) & (!g50)) + ((!g66) & (!g68) & (!g81) & (!g187) & (!g305) & (!g50)));
	assign g618 = (((g23) & (!i_24_) & (!g131) & (!g126) & (!sk[5]) & (!g219)) + ((!g23) & (i_24_) & (!g131) & (!g126) & (!sk[5]) & (!g219)) + ((g23) & (i_24_) & (!g131) & (g126) & (!sk[5]) & (!g219)) + ((g23) & (!i_24_) & (g131) & (!g126) & (!sk[5]) & (g219)));
	assign g619 = (((i_22_) & (!i_21_) & (!g9) & (!sk[6]) & (!g608) & (!g618)) + ((!i_22_) & (i_21_) & (!g9) & (!sk[6]) & (!g608) & (!g618)) + ((!i_22_) & (i_21_) & (!g9) & (!sk[6]) & (!g608) & (!g618)) + ((!i_22_) & (!i_21_) & (!g9) & (sk[6]) & (!g608) & (!g618)) + ((!i_22_) & (!i_21_) & (!g9) & (sk[6]) & (!g608) & (!g618)));
	assign g620 = (((i_38_) & (!sk[7]) & (i_39_) & (!i_40_)) + ((!i_38_) & (!sk[7]) & (i_39_) & (!i_40_)) + ((i_38_) & (!sk[7]) & (!i_39_) & (i_40_)) + ((!i_38_) & (sk[7]) & (!i_39_) & (!i_40_)));
	assign g621 = (((i_22_) & (!sk[8]) & (!g151) & (!g266) & (!g432) & (!g620)) + ((!i_22_) & (!sk[8]) & (g151) & (!g266) & (!g432) & (!g620)) + ((!i_22_) & (!sk[8]) & (g151) & (g266) & (!g432) & (!g620)) + ((!i_22_) & (sk[8]) & (!g151) & (!g266) & (g432) & (!g620)) + ((!i_22_) & (!sk[8]) & (g151) & (!g266) & (!g432) & (g620)));
	assign g622 = (((!sk[9]) & (!g151) & (i_21_) & (!g187) & (!g621)) + ((!sk[9]) & (!g151) & (!i_21_) & (g187) & (!g621)) + ((!sk[9]) & (!g151) & (i_21_) & (!g187) & (!g621)) + ((sk[9]) & (!g151) & (!i_21_) & (!g187) & (!g621)) + ((!sk[9]) & (!g151) & (!i_21_) & (g187) & (!g621)));
	assign g623 = (((!sk[10]) & (!i_24_) & (g84) & (!i_21_) & (!i_23_)) + ((!sk[10]) & (!i_24_) & (!g84) & (i_21_) & (!i_23_)) + ((!sk[10]) & (i_24_) & (g84) & (!i_21_) & (!i_23_)));
	assign g624 = (((!g74) & (g325) & (!sk[11]) & (!g600) & (!g623)) + ((!g74) & (!g325) & (!sk[11]) & (g600) & (!g623)) + ((!g74) & (!g325) & (sk[11]) & (!g600) & (!g623)) + ((!g74) & (!g325) & (sk[11]) & (!g600) & (!g623)));
	assign o_30_ = (((g65) & (!g23) & (!i_24_) & (!sk[12]) & (!g622) & (!g624)) + ((!g65) & (g23) & (!i_24_) & (!sk[12]) & (!g622) & (!g624)) + ((!g65) & (!g23) & (!i_24_) & (sk[12]) & (!g622) & (!g624)) + ((g65) & (g23) & (i_24_) & (!sk[12]) & (!g622) & (!g624)));
	assign g626 = (((!i_22_) & (g84) & (!sk[13]) & (!i_21_) & (!g325)) + ((!i_22_) & (!g84) & (!sk[13]) & (i_21_) & (!g325)) + ((i_22_) & (g84) & (!sk[13]) & (!i_21_) & (g325)));
	assign g627 = (((!g61) & (g125) & (!g390) & (!sk[14]) & (!g626)) + ((!g61) & (!g125) & (g390) & (!sk[14]) & (!g626)) + ((!g61) & (!g125) & (!g390) & (sk[14]) & (!g626)) + ((!g61) & (!g125) & (!g390) & (sk[14]) & (!g626)) + ((!g61) & (!g125) & (!g390) & (sk[14]) & (!g626)));
	assign o_31_ = (((g29) & (!sk[15]) & (!i_23_) & (!g17) & (!g615) & (!g627)) + ((!g29) & (!sk[15]) & (i_23_) & (!g17) & (!g615) & (!g627)) + ((!g29) & (sk[15]) & (!i_23_) & (g17) & (!g615) & (!g627)) + ((!g29) & (sk[15]) & (!i_23_) & (!g17) & (!g615) & (!g627)) + ((!g29) & (sk[15]) & (!i_23_) & (!g17) & (!g615) & (!g627)));
	assign g629 = (((!sk[16]) & (!i_31_) & (i_5_) & (!i_15_) & (!g401)) + ((!sk[16]) & (!i_31_) & (!i_5_) & (i_15_) & (!g401)) + ((sk[16]) & (!i_31_) & (!i_5_) & (!i_15_) & (g401)));
	assign g630 = (((!g100) & (i_35_) & (!sk[17]) & (!g73) & (!g172)) + ((!g100) & (!i_35_) & (!sk[17]) & (g73) & (!g172)) + ((g100) & (i_35_) & (!sk[17]) & (g73) & (g172)));
	assign g631 = (((i_36_) & (!i_37_) & (i_38_) & (i_39_) & (!i_40_) & (!i_35_)) + ((i_36_) & (i_37_) & (!i_38_) & (i_39_) & (i_40_) & (i_35_)) + ((i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (!i_35_)));
	assign g632 = (((g101) & (!sk[19]) & (!g151) & (!g204) & (!g220) & (!g436)) + ((!g101) & (!sk[19]) & (g151) & (!g204) & (!g220) & (!g436)) + ((!g101) & (sk[19]) & (!g151) & (g204) & (!g220) & (!g436)) + ((g101) & (!sk[19]) & (g151) & (!g204) & (!g220) & (g436)));
	assign g633 = (((g65) & (g629) & (!sk[20]) & (!g630) & (!g631) & (!g632)) + ((g65) & (!g629) & (!sk[20]) & (!g630) & (!g631) & (!g632)) + ((!g65) & (g629) & (!sk[20]) & (!g630) & (!g631) & (!g632)) + ((g65) & (!g629) & (!sk[20]) & (g630) & (!g631) & (!g632)) + ((g65) & (!g629) & (!sk[20]) & (!g630) & (g631) & (!g632)) + ((g65) & (!g629) & (!sk[20]) & (!g630) & (!g631) & (g632)));
	assign g634 = (((!sk[21]) & (i_37_) & (!i_34_) & (!i_35_) & (!g3) & (!g260)) + ((!sk[21]) & (!i_37_) & (i_34_) & (!i_35_) & (!g3) & (!g260)) + ((sk[21]) & (!i_37_) & (!i_34_) & (!i_35_) & (g3) & (g260)));
	assign g635 = (((!sk[22]) & (g56) & (!i_32_) & (!i_31_) & (!g24) & (!g46)) + ((!sk[22]) & (!g56) & (i_32_) & (!i_31_) & (!g24) & (!g46)) + ((!sk[22]) & (g56) & (!i_32_) & (!i_31_) & (!g24) & (g46)));
	assign g636 = (((g24) & (!g138) & (!sk[23]) & (!g275) & (!g634) & (!g635)) + ((!g24) & (g138) & (!sk[23]) & (!g275) & (!g634) & (!g635)) + ((g24) & (!g138) & (!sk[23]) & (!g275) & (!g634) & (!g635)) + ((!g24) & (!g138) & (sk[23]) & (!g275) & (!g634) & (!g635)) + ((!g24) & (!g138) & (sk[23]) & (!g275) & (!g634) & (!g635)));
	assign g637 = (((!i_31_) & (i_5_) & (!i_15_) & (!sk[24]) & (!g180)) + ((!i_31_) & (!i_5_) & (i_15_) & (!sk[24]) & (!g180)) + ((!i_31_) & (!i_5_) & (!i_15_) & (sk[24]) & (g180)));
	assign g638 = (((!i_5_) & (i_9_) & (!sk[25]) & (!g637)) + ((i_5_) & (!i_9_) & (!sk[25]) & (g637)) + ((!i_5_) & (!i_9_) & (sk[25]) & (!g637)) + ((i_5_) & (!i_9_) & (sk[25]) & (!g637)));
	assign g639 = (((!sk[26]) & (!i_40_) & (g56) & (!g46) & (!g275)) + ((!sk[26]) & (!i_40_) & (!g56) & (g46) & (!g275)) + ((!sk[26]) & (!i_40_) & (g56) & (g46) & (!g275)) + ((sk[26]) & (i_40_) & (!g56) & (!g46) & (g275)));
	assign g640 = (((!sk[27]) & (!g24) & (g138) & (!i_14_)) + ((!sk[27]) & (g24) & (!g138) & (i_14_)) + ((!sk[27]) & (!g24) & (g138) & (!i_14_)));
	assign g641 = (((!sk[28]) & (g53) & (!g470) & (!g637) & (!g639) & (!g640)) + ((!sk[28]) & (!g53) & (g470) & (!g637) & (!g639) & (!g640)) + ((sk[28]) & (!g53) & (!g470) & (!g637) & (!g639) & (!g640)) + ((sk[28]) & (!g53) & (!g470) & (!g637) & (!g639) & (!g640)) + ((sk[28]) & (!g53) & (!g470) & (!g637) & (!g639) & (!g640)) + ((sk[28]) & (!g53) & (!g470) & (!g637) & (!g639) & (!g640)));
	assign g642 = (((!i_12_) & (!i_15_) & (!g634) & (!g636) & (!g638) & (!g641)) + ((!i_12_) & (!i_15_) & (g634) & (!g636) & (!g638) & (!g641)) + ((!i_12_) & (!i_15_) & (!g634) & (!g636) & (!g638) & (!g641)));
	assign g643 = (((!g100) & (i_40_) & (!sk[30]) & (!g122) & (!i_6_)) + ((!g100) & (!i_40_) & (!sk[30]) & (g122) & (!i_6_)) + ((!g100) & (i_40_) & (!sk[30]) & (!g122) & (i_6_)));
	assign g644 = (((!g116) & (g160) & (!sk[31]) & (!g94) & (!g643)) + ((!g116) & (!g160) & (!sk[31]) & (g94) & (!g643)) + ((!g116) & (g160) & (!sk[31]) & (!g94) & (g643)) + ((g116) & (!g160) & (sk[31]) & (!g94) & (g643)));
	assign g645 = (((!sk[32]) & (!i_37_) & (i_38_) & (!i_39_) & (!i_40_)) + ((!sk[32]) & (!i_37_) & (!i_38_) & (i_39_) & (!i_40_)) + ((!sk[32]) & (!i_37_) & (!i_38_) & (i_39_) & (!i_40_)) + ((sk[32]) & (!i_37_) & (!i_38_) & (!i_39_) & (i_40_)) + ((!sk[32]) & (!i_37_) & (!i_38_) & (i_39_) & (i_40_)) + ((sk[32]) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_)));
	assign g646 = (((i_37_) & (!sk[33]) & (!g122) & (!i_13_) & (!g5) & (!g187)) + ((!i_37_) & (!sk[33]) & (g122) & (!i_13_) & (!g5) & (!g187)) + ((!i_37_) & (sk[33]) & (!g122) & (!i_13_) & (g5) & (g187)));
	assign g647 = (((g2) & (!g3) & (!sk[34]) & (!g189) & (!g645) & (!g646)) + ((!g2) & (g3) & (!sk[34]) & (!g189) & (!g645) & (!g646)) + ((!g2) & (!g3) & (sk[34]) & (!g189) & (!g645) & (!g646)) + ((!g2) & (!g3) & (sk[34]) & (!g189) & (!g645) & (!g646)) + ((!g2) & (!g3) & (sk[34]) & (!g189) & (!g645) & (!g646)));
	assign g648 = (((i_5_) & (!g22) & (!i_13_) & (!g132) & (!g644) & (!g647)) + ((!i_5_) & (!g22) & (!i_13_) & (!g132) & (!g644) & (!g647)) + ((!i_5_) & (!g22) & (i_13_) & (!g132) & (!g644) & (g647)) + ((!i_5_) & (!g22) & (!i_13_) & (!g132) & (!g644) & (g647)));
	assign g649 = (((i_32_) & (!i_31_) & (!i_5_) & (!sk[36]) & (!g171) & (!g201)) + ((!i_32_) & (i_31_) & (!i_5_) & (!sk[36]) & (!g171) & (!g201)) + ((!i_32_) & (!i_31_) & (!i_5_) & (sk[36]) & (g171) & (!g201)));
	assign g650 = (((!sk[37]) & (g100) & (!i_39_) & (!i_40_) & (!i_35_) & (!g151)) + ((!sk[37]) & (!g100) & (i_39_) & (!i_40_) & (!i_35_) & (!g151)) + ((!sk[37]) & (!g100) & (i_39_) & (i_40_) & (!i_35_) & (g151)) + ((!sk[37]) & (g100) & (!i_39_) & (!i_40_) & (i_35_) & (!g151)));
	assign g651 = (((i_36_) & (!sk[38]) & (!i_32_) & (!g10) & (!g67) & (!g187)) + ((!i_36_) & (!sk[38]) & (i_32_) & (!g10) & (!g67) & (!g187)) + ((i_36_) & (!sk[38]) & (!i_32_) & (!g10) & (g67) & (g187)));
	assign g652 = (((!g423) & (!sk[39]) & (g465) & (!g650) & (!g651)) + ((g423) & (!sk[39]) & (!g465) & (g650) & (!g651)) + ((!g423) & (!sk[39]) & (!g465) & (g650) & (!g651)) + ((!g423) & (!sk[39]) & (g465) & (!g650) & (g651)));
	assign g653 = (((!sk[40]) & (!i_40_) & (g98) & (!g214)) + ((!sk[40]) & (i_40_) & (!g98) & (g214)) + ((!sk[40]) & (i_40_) & (g98) & (g214)));
	assign g654 = (((i_40_) & (!g122) & (!sk[41]) & (!g21) & (!g47) & (!g94)) + ((!i_40_) & (g122) & (!sk[41]) & (!g21) & (!g47) & (!g94)) + ((!i_40_) & (!g122) & (sk[41]) & (g21) & (g47) & (!g94)));
	assign g655 = (((i_33_) & (i_32_) & (!g86) & (!g67) & (!g461) & (!g654)) + ((!i_33_) & (!i_32_) & (!g86) & (!g67) & (!g461) & (!g654)) + ((!i_33_) & (!i_32_) & (!g86) & (!g67) & (!g461) & (!g654)) + ((!i_33_) & (!i_32_) & (!g86) & (!g67) & (!g461) & (!g654)));
	assign g656 = (((!g22) & (g218) & (!g653) & (!sk[43]) & (!g655)) + ((!g22) & (!g218) & (g653) & (!sk[43]) & (!g655)) + ((g22) & (g218) & (!g653) & (!sk[43]) & (g655)) + ((!g22) & (g218) & (!g653) & (!sk[43]) & (g655)));
	assign g657 = (((!sk[44]) & (g450) & (!g458) & (!g649) & (!g652) & (!g656)) + ((!sk[44]) & (!g450) & (g458) & (!g649) & (!g652) & (!g656)) + ((!sk[44]) & (!g450) & (g458) & (!g649) & (!g652) & (g656)) + ((!sk[44]) & (!g450) & (g458) & (!g649) & (!g652) & (g656)));
	assign g658 = (((!sk[45]) & (!g135) & (g84) & (!g152) & (!g172)) + ((!sk[45]) & (!g135) & (!g84) & (g152) & (!g172)) + ((!sk[45]) & (!g135) & (g84) & (!g152) & (g172)) + ((sk[45]) & (!g135) & (!g84) & (!g152) & (g172)) + ((!sk[45]) & (g135) & (!g84) & (g152) & (g172)));
	assign g659 = (((i_11_) & (!sk[46]) & (!i_5_) & (!i_9_) & (!g636) & (!g658)) + ((!i_11_) & (!sk[46]) & (i_5_) & (!i_9_) & (!g636) & (!g658)) + ((i_11_) & (!sk[46]) & (!i_5_) & (!i_9_) & (!g636) & (!g658)) + ((!i_11_) & (!sk[46]) & (i_5_) & (!i_9_) & (!g636) & (!g658)) + ((!i_11_) & (sk[46]) & (!i_5_) & (!i_9_) & (!g636) & (!g658)) + ((!i_11_) & (sk[46]) & (!i_5_) & (!i_9_) & (g636) & (!g658)));
	assign g660 = (((!g633) & (!g642) & (g648) & (g435) & (g657) & (g659)));
	assign g661 = (((i_36_) & (!i_37_) & (i_38_) & (i_39_) & (!i_40_) & (g462)) + ((i_36_) & (i_37_) & (i_38_) & (!i_39_) & (i_40_) & (g462)));
	assign g662 = (((!sk[49]) & (i_36_) & (!i_5_) & (!i_15_) & (!g201) & (!g661)) + ((!sk[49]) & (!i_36_) & (i_5_) & (!i_15_) & (!g201) & (!g661)) + ((!sk[49]) & (i_36_) & (!i_5_) & (!i_15_) & (!g201) & (!g661)) + ((sk[49]) & (!i_36_) & (!i_5_) & (!i_15_) & (!g201) & (!g661)) + ((!sk[49]) & (!i_36_) & (i_5_) & (i_15_) & (g201) & (!g661)));
	assign g663 = (((i_36_) & (!sk[50]) & (!g162) & (!i_35_) & (!g112) & (!g260)) + ((!i_36_) & (!sk[50]) & (g162) & (!i_35_) & (!g112) & (!g260)) + ((!i_36_) & (sk[50]) & (!g162) & (!i_35_) & (g112) & (!g260)) + ((!i_36_) & (sk[50]) & (!g162) & (!i_35_) & (!g112) & (g260)));
	assign g664 = (((g100) & (!g101) & (!g280) & (!g255) & (!sk[51]) & (!g663)) + ((!g100) & (g101) & (!g280) & (!g255) & (!sk[51]) & (!g663)) + ((!g100) & (g101) & (!g280) & (!g255) & (!sk[51]) & (!g663)) + ((!g100) & (!g101) & (!g280) & (!g255) & (sk[51]) & (!g663)) + ((!g100) & (!g101) & (!g280) & (g255) & (sk[51]) & (!g663)));
	assign g665 = (((i_36_) & (!i_40_) & (!g162) & (!sk[52]) & (!g346) & (!g664)) + ((!i_36_) & (i_40_) & (!g162) & (!sk[52]) & (!g346) & (!g664)) + ((!i_36_) & (!i_40_) & (!g162) & (sk[52]) & (!g346) & (g664)) + ((!i_36_) & (!i_40_) & (!g162) & (sk[52]) & (!g346) & (g664)) + ((!i_36_) & (!i_40_) & (g162) & (sk[52]) & (!g346) & (g664)) + ((!i_36_) & (!i_40_) & (!g162) & (sk[52]) & (!g346) & (g664)));
	assign g666 = (((i_36_) & (!i_40_) & (!sk[53]) & (!g162) & (!g21) & (!g465)) + ((!i_36_) & (i_40_) & (!sk[53]) & (!g162) & (!g21) & (!g465)) + ((i_36_) & (!i_40_) & (!sk[53]) & (!g162) & (g21) & (g465)));
	assign g667 = (((!i_36_) & (g100) & (!sk[54]) & (!g101) & (!g49)) + ((!i_36_) & (!g100) & (!sk[54]) & (g101) & (!g49)) + ((!i_36_) & (g100) & (!sk[54]) & (!g101) & (!g49)));
	assign g668 = (((!sk[55]) & (g280) & (!g67) & (!g461) & (!g666) & (!g667)) + ((!sk[55]) & (!g280) & (g67) & (!g461) & (!g666) & (!g667)) + ((!sk[55]) & (!g280) & (g67) & (!g461) & (g666) & (!g667)) + ((!sk[55]) & (g280) & (g67) & (g461) & (!g666) & (!g667)) + ((!sk[55]) & (!g280) & (g67) & (g461) & (!g666) & (g667)));
	assign g669 = (((!sk[56]) & (i_32_) & (!i_5_) & (!i_0_) & (!g665) & (!g668)) + ((!sk[56]) & (!i_32_) & (i_5_) & (!i_0_) & (!g665) & (!g668)) + ((sk[56]) & (!i_32_) & (!i_5_) & (!i_0_) & (!g665) & (g668)) + ((!sk[56]) & (!i_32_) & (i_5_) & (!i_0_) & (!g665) & (!g668)));
	assign g670 = (((i_37_) & (!i_35_) & (!g53) & (!sk[57]) & (!i_9_) & (!g260)) + ((!i_37_) & (i_35_) & (!g53) & (!sk[57]) & (!i_9_) & (!g260)) + ((!i_37_) & (!i_35_) & (g53) & (sk[57]) & (i_9_) & (g260)));
	assign g671 = (((i_11_) & (!i_38_) & (!sk[58]) & (!g73) & (!g219) & (!g653)) + ((!i_11_) & (i_38_) & (!sk[58]) & (!g73) & (!g219) & (!g653)) + ((i_11_) & (!i_38_) & (!sk[58]) & (!g73) & (!g219) & (g653)) + ((!i_11_) & (i_38_) & (!sk[58]) & (g73) & (g219) & (!g653)));
	assign g672 = (((!g2) & (g21) & (!g3) & (!sk[59]) & (!g201)) + ((!g2) & (!g21) & (g3) & (!sk[59]) & (!g201)) + ((g2) & (g21) & (g3) & (!sk[59]) & (!g201)));
	assign g673 = (((!sk[60]) & (!g53) & (g136) & (!g79) & (!g672)) + ((!sk[60]) & (!g53) & (!g136) & (g79) & (!g672)) + ((sk[60]) & (!g53) & (!g136) & (!g79) & (!g672)) + ((sk[60]) & (!g53) & (!g136) & (!g79) & (!g672)) + ((sk[60]) & (!g53) & (!g136) & (!g79) & (!g672)));
	assign g674 = (((i_39_) & (!sk[61]) & (!g53) & (!i_15_) & (!i_9_) & (!g136)) + ((!i_39_) & (!sk[61]) & (g53) & (!i_15_) & (!i_9_) & (!g136)) + ((i_39_) & (!sk[61]) & (g53) & (!i_15_) & (i_9_) & (g136)));
	assign g675 = (((g171) & (!g493) & (!g673) & (!g203) & (!sk[62]) & (!g674)) + ((!g171) & (g493) & (!g673) & (!g203) & (!sk[62]) & (!g674)) + ((!g171) & (!g493) & (!g673) & (!g203) & (sk[62]) & (!g674)) + ((!g171) & (!g493) & (g673) & (!g203) & (sk[62]) & (!g674)));
	assign g676 = (((g385) & (!g457) & (!g670) & (!sk[63]) & (!g671) & (!g675)) + ((!g385) & (g457) & (!g670) & (!sk[63]) & (!g671) & (!g675)) + ((g385) & (g457) & (!g670) & (!sk[63]) & (!g671) & (g675)) + ((!g385) & (g457) & (!g670) & (!sk[63]) & (!g671) & (g675)));
	assign g677 = (((!i_37_) & (i_38_) & (i_39_) & (i_40_) & (g160) & (!g94)) + ((i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (g160) & (!g94)) + ((i_37_) & (i_38_) & (i_39_) & (i_40_) & (!g160) & (!g94)));
	assign g678 = (((i_36_) & (!i_37_) & (!i_40_) & (!g162) & (!sk[65]) & (!g104)) + ((!i_36_) & (i_37_) & (!i_40_) & (!g162) & (!sk[65]) & (!g104)) + ((!i_36_) & (!i_37_) & (!i_40_) & (!g162) & (sk[65]) & (g104)));
	assign g679 = (((!i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (i_40_) & (g56)) + ((!i_36_) & (!i_37_) & (!i_38_) & (i_39_) & (!i_40_) & (g56)) + ((!i_36_) & (i_37_) & (!i_38_) & (!i_39_) & (!i_40_) & (g56)) + ((!i_36_) & (!i_37_) & (!i_38_) & (i_39_) & (i_40_) & (g56)));
	assign g680 = (((i_32_) & (!i_31_) & (!sk[67]) & (!i_15_) & (!g678) & (!g679)) + ((!i_32_) & (i_31_) & (!sk[67]) & (!i_15_) & (!g678) & (!g679)) + ((!i_32_) & (!i_31_) & (sk[67]) & (!i_15_) & (g678) & (!g679)) + ((!i_32_) & (!i_31_) & (sk[67]) & (!i_15_) & (!g678) & (g679)));
	assign g681 = (((i_31_) & (!g22) & (!sk[68]) & (!g27) & (!g73) & (!g401)) + ((!i_31_) & (g22) & (!sk[68]) & (!g27) & (!g73) & (!g401)) + ((!i_31_) & (g22) & (!sk[68]) & (!g27) & (!g73) & (g401)) + ((!i_31_) & (g22) & (!sk[68]) & (g27) & (g73) & (!g401)));
	assign g682 = (((!i_37_) & (g260) & (!sk[69]) & (!g78) & (!g187)) + ((!i_37_) & (!g260) & (!sk[69]) & (g78) & (!g187)) + ((!i_37_) & (g260) & (!sk[69]) & (g78) & (!g187)) + ((i_37_) & (!g260) & (!sk[69]) & (g78) & (g187)));
	assign g683 = (((!g51) & (i_5_) & (!g195) & (!sk[70]) & (!g682)) + ((!g51) & (!i_5_) & (g195) & (!sk[70]) & (!g682)) + ((!g51) & (!i_5_) & (!g195) & (sk[70]) & (!g682)) + ((!g51) & (!i_5_) & (!g195) & (sk[70]) & (!g682)) + ((!g51) & (!i_5_) & (!g195) & (sk[70]) & (!g682)));
	assign g684 = (((!i_36_) & (!i_37_) & (i_38_) & (!i_39_) & (!i_34_) & (!i_35_)) + ((!i_36_) & (!i_37_) & (!i_38_) & (i_39_) & (!i_34_) & (!i_35_)) + ((!i_36_) & (!i_37_) & (i_38_) & (i_39_) & (!i_34_) & (!i_35_)) + ((!i_36_) & (!i_37_) & (!i_38_) & (!i_39_) & (!i_34_) & (!i_35_)));
	assign g685 = (((!i_37_) & (g51) & (!sk[72]) & (!g131) & (!g684)) + ((!i_37_) & (!g51) & (!sk[72]) & (g131) & (!g684)) + ((!i_37_) & (!g51) & (sk[72]) & (!g131) & (!g684)) + ((!i_37_) & (!g51) & (sk[72]) & (!g131) & (!g684)) + ((!i_37_) & (!g51) & (sk[72]) & (!g131) & (!g684)));
	assign g686 = (((!sk[73]) & (g122) & (!i_5_) & (!g139) & (!g121) & (!g685)) + ((!sk[73]) & (!g122) & (i_5_) & (!g139) & (!g121) & (!g685)) + ((!sk[73]) & (!g122) & (i_5_) & (!g139) & (!g121) & (!g685)) + ((!sk[73]) & (!g122) & (i_5_) & (g139) & (g121) & (!g685)));
	assign g687 = (((!g65) & (g681) & (!g683) & (!sk[74]) & (!g686)) + ((!g65) & (!g681) & (g683) & (!sk[74]) & (!g686)) + ((!g65) & (!g681) & (g683) & (!sk[74]) & (!g686)) + ((!g65) & (!g681) & (!g683) & (sk[74]) & (!g686)));
	assign g688 = (((!sk[75]) & (g122) & (!i_6_) & (!g677) & (!g680) & (!g687)) + ((!sk[75]) & (!g122) & (i_6_) & (!g677) & (!g680) & (!g687)) + ((!sk[75]) & (g122) & (!i_6_) & (!g677) & (!g680) & (g687)) + ((sk[75]) & (!g122) & (!i_6_) & (!g677) & (!g680) & (g687)) + ((!sk[75]) & (!g122) & (i_6_) & (!g677) & (!g680) & (g687)));
	assign g689 = (((g102) & (!g662) & (!g669) & (!g676) & (!sk[76]) & (!g688)) + ((!g102) & (g662) & (!g669) & (!g676) & (!sk[76]) & (!g688)) + ((!g102) & (g662) & (!g669) & (g676) & (!sk[76]) & (g688)) + ((!g102) & (!g662) & (!g669) & (g676) & (sk[76]) & (g688)));
	assign g690 = (((i_17_) & (i_16_) & (i_15_) & (!i_12_) & (i_11_) & (!i_9_)) + ((i_17_) & (i_16_) & (i_15_) & (i_12_) & (!i_11_) & (!i_9_)) + ((i_17_) & (!i_16_) & (i_15_) & (!i_12_) & (i_11_) & (i_9_)) + ((!i_17_) & (i_16_) & (i_15_) & (!i_12_) & (i_11_) & (i_9_)) + ((i_17_) & (!i_16_) & (i_15_) & (i_12_) & (!i_11_) & (i_9_)) + ((!i_17_) & (i_16_) & (i_15_) & (i_12_) & (!i_11_) & (i_9_)));
	assign g691 = (((!sk[78]) & (!g690) & (i_5_)) + ((sk[78]) & (g690) & (!i_5_)));
	assign g692 = (((!i_19_) & (g23) & (!i_18_) & (!g18) & (!g34) & (g84)) + ((!i_19_) & (!g23) & (!i_18_) & (g18) & (g34) & (g84)) + ((!i_19_) & (!g23) & (!i_18_) & (g18) & (g34) & (g84)));
	assign g693 = (((!sk[80]) & (!g694) & (g695)) + ((sk[80]) & (!g694) & (!g695)));
	assign g694 = (((!i_32_) & (!sk[81]) & (g696)) + ((!i_32_) & (!sk[81]) & (g696)));
	assign g695 = (((!sk[82]) & (!i_32_) & (g699)) + ((!sk[82]) & (i_32_) & (g699)));
	assign g696 = (((!sk[83]) & (!g697) & (g698)) + ((sk[83]) & (!g697) & (!g698)));
	assign g697 = (((!sk[84]) & (!i_37_) & (g702)) + ((!sk[84]) & (!i_37_) & (g702)));
	assign g698 = (((i_37_) & (!sk[85]) & (g703)) + ((!i_37_) & (!sk[85]) & (g703)));
	assign g699 = (((!sk[86]) & (!g700) & (g701)) + ((sk[86]) & (!g700) & (!g701)));
	assign g700 = (((!i_37_) & (!sk[87]) & (g590)) + ((!i_37_) & (!sk[87]) & (g590)));
	assign g701 = (((!sk[88]) & (!i_37_) & (g590)) + ((!sk[88]) & (i_37_) & (g590)));
	assign g702 = (((g588) & (!sk[89]) & (g590)) + ((!g588) & (!sk[89]) & (g590)));
	assign g703 = (((!sk[90]) & (!i_5_) & (g162) & (!i_0_) & (!g590)) + ((!sk[90]) & (!i_5_) & (!g162) & (i_0_) & (!g590)) + ((!sk[90]) & (!i_5_) & (g162) & (!i_0_) & (g590)) + ((!sk[90]) & (!i_5_) & (!g162) & (i_0_) & (g590)) + ((sk[90]) & (!i_5_) & (!g162) & (!i_0_) & (g590)));
	assign g704 = (((!sk[91]) & (!g705) & (g706)) + ((sk[91]) & (!g705) & (!g706)));
	assign g705 = (((!i_37_) & (!sk[92]) & (g707)) + ((!i_37_) & (!sk[92]) & (g707)));
	assign g706 = (((i_37_) & (!sk[93]) & (g709)) + ((!i_37_) & (!sk[93]) & (g709)));
	assign g707 = (((!i_0_) & (!sk[94]) & (g708)) + ((!i_0_) & (sk[94]) & (!g708)));
	assign g708 = (((!i_0_) & (!sk[95]) & (g711)) + ((!i_0_) & (!sk[95]) & (g711)));
	assign g709 = (((!i_0_) & (!sk[96]) & (g710)) + ((i_0_) & (sk[96]) & (!g710)));
	assign g710 = (((!i_0_) & (!sk[97]) & (g125)) + ((i_0_) & (sk[97]) & (!g125)));
	assign g711 = (((!i_38_) & (g255) & (!sk[98]) & (!i_32_) & (!i_5_)) + ((!i_38_) & (!g255) & (!sk[98]) & (i_32_) & (!i_5_)) + ((i_38_) & (!g255) & (sk[98]) & (!i_32_) & (!i_5_)) + ((!i_38_) & (!g255) & (sk[98]) & (!i_32_) & (!i_5_)));
	assign g712 = (((!sk[99]) & (!g713) & (g714)) + ((sk[99]) & (!g713) & (!g714)));
	assign g713 = (((!i_37_) & (!sk[100]) & (g715)) + ((!i_37_) & (!sk[100]) & (g715)));
	assign g714 = (((!sk[101]) & (!i_37_) & (g717)) + ((!sk[101]) & (i_37_) & (g717)));
	assign g715 = (((!i_36_) & (!sk[102]) & (g716)) + ((i_36_) & (sk[102]) & (!g716)));
	assign g716 = (((!sk[103]) & (!i_36_) & (g720)) + ((!sk[103]) & (i_36_) & (g720)));
	assign g717 = (((!g718) & (!sk[104]) & (g719)) + ((!g718) & (sk[104]) & (!g719)));
	assign g718 = (((!sk[105]) & (!i_36_) & (g721)) + ((!sk[105]) & (!i_36_) & (g721)));
	assign g719 = (((!sk[106]) & (!i_36_) & (g722)) + ((!sk[106]) & (i_36_) & (g722)));
	assign g720 = (((!sk[107]) & (!i_40_) & (!i_39_) & (g10) & (!i_38_)) + ((!sk[107]) & (!i_40_) & (i_39_) & (!g10) & (!i_38_)) + ((sk[107]) & (!i_40_) & (!i_39_) & (!g10) & (!i_38_)) + ((!sk[107]) & (!i_40_) & (i_39_) & (!g10) & (!i_38_)) + ((!sk[107]) & (!i_40_) & (i_39_) & (!g10) & (!i_38_)));
	assign g721 = (((!i_40_) & (!i_39_) & (!sk[108]) & (g49) & (!i_38_)) + ((!i_40_) & (!i_39_) & (sk[108]) & (!g49) & (!i_38_)) + ((!i_40_) & (i_39_) & (!sk[108]) & (!g49) & (!i_38_)) + ((!i_40_) & (!i_39_) & (sk[108]) & (!g49) & (!i_38_)) + ((!i_40_) & (!i_39_) & (sk[108]) & (!g49) & (!i_38_)));
	assign g722 = (((!sk[109]) & (!i_40_) & (g10) & (!i_38_)) + ((sk[109]) & (!i_40_) & (!g10) & (!i_38_)) + ((!sk[109]) & (i_40_) & (!g10) & (i_38_)));
	assign g723 = (((!sk[110]) & (!i_40_) & (g724)) + ((!sk[110]) & (i_40_) & (g724)));
	assign g724 = (((!g725) & (!sk[111]) & (g726)) + ((!g725) & (sk[111]) & (!g726)));
	assign g725 = (((!g22) & (!sk[112]) & (g727)) + ((!g22) & (!sk[112]) & (g727)));
	assign g726 = (((!sk[113]) & (!g22) & (g728)) + ((!sk[113]) & (g22) & (g728)));
	assign g727 = (((!sk[114]) & (!g351) & (g349)) + ((!sk[114]) & (!g351) & (g349)));
	assign g728 = (((!g350) & (!sk[115]) & (g98) & (!g1) & (!g349)) + ((!g350) & (!sk[115]) & (!g98) & (g1) & (!g349)) + ((!g350) & (!sk[115]) & (!g98) & (g1) & (g349)) + ((!g350) & (sk[115]) & (!g98) & (!g1) & (g349)) + ((!g350) & (!sk[115]) & (g98) & (!g1) & (g349)));
	assign g729 = (((!sk[116]) & (!g730) & (g731)) + ((sk[116]) & (!g730) & (!g731)));
	assign g730 = (((!sk[117]) & (!g30) & (g732)) + ((!sk[117]) & (!g30) & (g732)));
	assign g731 = (((!sk[118]) & (!g30) & (g735)) + ((!sk[118]) & (g30) & (g735)));
	assign g732 = (((!sk[119]) & (!g733) & (g734)) + ((sk[119]) & (!g733) & (!g734)));
	assign g733 = (((!sk[120]) & (!i_37_) & (g737)) + ((!sk[120]) & (!i_37_) & (g737)));
	assign g734 = (((!sk[121]) & (!i_37_) & (g738)) + ((!sk[121]) & (i_37_) & (g738)));
	assign g735 = (((!sk[122]) & (!i_37_) & (g736)) + ((sk[122]) & (!i_37_) & (!g736)));
	assign g736 = (((!sk[123]) & (!i_37_) & (g739)) + ((!sk[123]) & (!i_37_) & (g739)));
	assign g737 = (((!g5) & (g122) & (!sk[124]) & (!g266)) + ((!g5) & (!g122) & (sk[124]) & (!g266)) + ((!g5) & (!g122) & (sk[124]) & (!g266)) + ((g5) & (!g122) & (!sk[124]) & (g266)));
	assign g738 = (((!sk[125]) & (!g267) & (g94)) + ((sk[125]) & (!g267) & (!g94)));
	assign g739 = (((!g5) & (g122) & (!sk[126]) & (!g266)) + ((!g5) & (!g122) & (sk[126]) & (!g266)) + ((!g5) & (!g122) & (sk[126]) & (!g266)) + ((g5) & (!g122) & (!sk[126]) & (g266)));
	assign g740 = (((!sk[127]) & (!i_36_) & (g741)) + ((sk[127]) & (i_36_) & (!g741)));
	assign g741 = (((!sk[0]) & (!i_36_) & (g742)) + ((!sk[0]) & (i_36_) & (g742)));
	assign g742 = (((!sk[1]) & (!g743) & (g744)) + ((sk[1]) & (!g743) & (!g744)));
	assign g743 = (((!sk[2]) & (!i_40_) & (g745)) + ((!sk[2]) & (!i_40_) & (g745)));
	assign g744 = (((!sk[3]) & (!i_40_) & (g746)) + ((!sk[3]) & (i_40_) & (g746)));
	assign g745 = (((!i_37_) & (!sk[4]) & (i_39_) & (!i_35_) & (!g92)) + ((!i_37_) & (!sk[4]) & (!i_39_) & (i_35_) & (!g92)) + ((!i_37_) & (sk[4]) & (!i_39_) & (!i_35_) & (!g92)) + ((!i_37_) & (!sk[4]) & (!i_39_) & (i_35_) & (!g92)) + ((!i_37_) & (!sk[4]) & (!i_39_) & (i_35_) & (!g92)));
	assign g746 = (((!i_37_) & (!i_39_) & (sk[5]) & (!i_38_) & (!g92)) + ((!i_37_) & (!i_39_) & (!sk[5]) & (i_38_) & (!g92)) + ((!i_37_) & (!i_39_) & (!sk[5]) & (i_38_) & (!g92)) + ((!i_37_) & (i_39_) & (!sk[5]) & (!i_38_) & (!g92)) + ((!i_37_) & (!i_39_) & (!sk[5]) & (i_38_) & (!g92)));
	assign g747 = (((!g748) & (!sk[6]) & (g749)) + ((!g748) & (sk[6]) & (!g749)));
	assign g748 = (((!sk[7]) & (!g152) & (g750)) + ((!sk[7]) & (!g152) & (g750)));
	assign g749 = (((!sk[8]) & (!g152) & (g753)) + ((!sk[8]) & (g152) & (g753)));
	assign g750 = (((!g751) & (!sk[9]) & (g752)) + ((!g751) & (sk[9]) & (!g752)));
	assign g751 = (((!sk[10]) & (!i_18_) & (g756)) + ((!sk[10]) & (!i_18_) & (g756)));
	assign g752 = (((!sk[11]) & (!i_18_) & (g757)) + ((!sk[11]) & (i_18_) & (g757)));
	assign g753 = (((!sk[12]) & (!g754) & (g755)) + ((sk[12]) & (!g754) & (!g755)));
	assign g754 = (((!i_18_) & (!sk[13]) & (g758)) + ((!i_18_) & (!sk[13]) & (g758)));
	assign g755 = (((!sk[14]) & (!i_18_) & (g759)) + ((!sk[14]) & (i_18_) & (g759)));
	assign g756 = (((!g34) & (!sk[15]) & (g156) & (!g18) & (!g154)) + ((!g34) & (!sk[15]) & (!g156) & (g18) & (!g154)) + ((!g34) & (sk[15]) & (!g156) & (!g18) & (!g154)) + ((!g34) & (!sk[15]) & (!g156) & (g18) & (!g154)) + ((!g34) & (!sk[15]) & (g156) & (!g18) & (!g154)) + ((!g34) & (!sk[15]) & (g156) & (!g18) & (!g154)));
	assign g757 = (((!g34) & (!sk[16]) & (g156) & (!g157) & (!g154)) + ((!g34) & (!sk[16]) & (!g156) & (g157) & (!g154)) + ((!g34) & (sk[16]) & (!g156) & (!g157) & (!g154)) + ((!g34) & (sk[16]) & (!g156) & (!g157) & (!g154)) + ((!g34) & (!sk[16]) & (!g156) & (g157) & (!g154)));
	assign g758 = (((!sk[17]) & (!g156) & (g154)) + ((sk[17]) & (!g156) & (!g154)) + ((!sk[17]) & (!g156) & (g154)));
	assign g759 = (((!g34) & (g156) & (!g157) & (!sk[18]) & (!g154)) + ((!g34) & (!g156) & (g157) & (!sk[18]) & (!g154)) + ((!g34) & (!g156) & (!g157) & (sk[18]) & (!g154)) + ((!g34) & (!g156) & (!g157) & (sk[18]) & (!g154)) + ((!g34) & (!g156) & (!g157) & (sk[18]) & (!g154)));

endmodule