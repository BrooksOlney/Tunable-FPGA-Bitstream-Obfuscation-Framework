module ks__altor32_qmap_map (sk, dmem_ack_i, clk_i, rst_i, dmem_stall_i, nmi_i, intr_i, dmem_dat_ix28x, dmem_dat_ix27x, dmem_dat_ix31x, dmem_dat_ix30x, dmem_dat_ix29x, dmem_dat_ix26x, dmem_dat_ix7x, dmem_dat_ix6x, dmem_dat_ix2x, dmem_dat_ix1x, dmem_dat_ix0x, dmem_dat_ix3x, dmem_dat_ix9x, dmem_dat_ix8x, dmem_dat_ix25x, dmem_dat_ix23x, dmem_dat_ix22x, dmem_dat_ix24x, dmem_dat_ix20x, dmem_dat_ix16x, dmem_dat_ix19x, dmem_dat_ix18x, dmem_dat_ix17x, dmem_dat_ix10x, dmem_dat_ix11x, dmem_dat_ix4x, dmem_dat_ix12x, dmem_dat_ix5x, dmem_dat_ix13x, dmem_dat_ix21x, dmem_dat_ix14x, dmem_dat_ix15x, fault_o, break_o, imem_addr_ox0x, imem_addr_ox1x, imem_addr_ox2x, imem_addr_ox3x, imem_addr_ox4x, imem_addr_ox5x, imem_addr_ox6x, imem_addr_ox7x, imem_addr_ox8x, imem_addr_ox9x, imem_addr_ox10x, imem_addr_ox11x, imem_addr_ox12x, imem_addr_ox13x, imem_addr_ox14x, imem_addr_ox15x, imem_addr_ox16x, imem_addr_ox17x, imem_addr_ox18x, imem_addr_ox19x, imem_addr_ox20x, imem_addr_ox21x, imem_addr_ox22x, imem_addr_ox23x, imem_addr_ox24x, imem_addr_ox25x, imem_addr_ox26x, imem_addr_ox27x, imem_addr_ox28x, imem_addr_ox29x, imem_addr_ox30x, imem_addr_ox31x, imem_cti_ox0x, imem_cti_ox1x, imem_cti_ox2x, imem_cyc_o, imem_stb_o, dmem_addr_ox0x, dmem_addr_ox1x, dmem_addr_ox2x, dmem_addr_ox3x, dmem_addr_ox4x, dmem_addr_ox5x, dmem_addr_ox6x, dmem_addr_ox7x, dmem_addr_ox8x, dmem_addr_ox9x, dmem_addr_ox10x, dmem_addr_ox11x, dmem_addr_ox12x, dmem_addr_ox13x, dmem_addr_ox14x, dmem_addr_ox15x, dmem_addr_ox16x, dmem_addr_ox17x, dmem_addr_ox18x, dmem_addr_ox19x, dmem_addr_ox20x, dmem_addr_ox21x, dmem_addr_ox22x, dmem_addr_ox23x, dmem_addr_ox24x, dmem_addr_ox25x, dmem_addr_ox26x, dmem_addr_ox27x, dmem_addr_ox28x, dmem_addr_ox29x, dmem_addr_ox30x, dmem_addr_ox31x, dmem_dat_ox0x, dmem_dat_ox1x, dmem_dat_ox2x, dmem_dat_ox3x, dmem_dat_ox4x, dmem_dat_ox5x, dmem_dat_ox6x, dmem_dat_ox7x, dmem_dat_ox8x, dmem_dat_ox9x, dmem_dat_ox10x, dmem_dat_ox11x, dmem_dat_ox12x, dmem_dat_ox13x, dmem_dat_ox14x, dmem_dat_ox15x, dmem_dat_ox16x, dmem_dat_ox17x, dmem_dat_ox18x, dmem_dat_ox19x, dmem_dat_ox20x, dmem_dat_ox21x, dmem_dat_ox22x, dmem_dat_ox23x, dmem_dat_ox24x, dmem_dat_ox25x, dmem_dat_ox26x, dmem_dat_ox27x, dmem_dat_ox28x, dmem_dat_ox29x, dmem_dat_ox30x, dmem_dat_ox31x, dmem_cti_ox0x, dmem_cti_ox1x, dmem_cti_ox2x, dmem_cyc_o, dmem_stb_o, dmem_we_o, dmem_sel_ox0x, dmem_sel_ox1x, dmem_sel_ox2x, dmem_sel_ox3x);

	input dmem_ack_i;
	input clk_i;
	input rst_i;
	input dmem_stall_i;
	input nmi_i;
	input intr_i;
	input dmem_dat_ix28x;
	input dmem_dat_ix27x;
	input dmem_dat_ix31x;
	input dmem_dat_ix30x;
	input dmem_dat_ix29x;
	input dmem_dat_ix26x;
	input dmem_dat_ix7x;
	input dmem_dat_ix6x;
	input dmem_dat_ix2x;
	input dmem_dat_ix1x;
	input dmem_dat_ix0x;
	input dmem_dat_ix3x;
	input dmem_dat_ix9x;
	input dmem_dat_ix8x;
	input dmem_dat_ix25x;
	input dmem_dat_ix23x;
	input dmem_dat_ix22x;
	input dmem_dat_ix24x;
	input dmem_dat_ix20x;
	input dmem_dat_ix16x;
	input dmem_dat_ix19x;
	input dmem_dat_ix18x;
	input dmem_dat_ix17x;
	input dmem_dat_ix10x;
	input dmem_dat_ix11x;
	input dmem_dat_ix4x;
	input dmem_dat_ix12x;
	input dmem_dat_ix5x;
	input dmem_dat_ix13x;
	input dmem_dat_ix21x;
	input dmem_dat_ix14x;
	input dmem_dat_ix15x;
	output fault_o;
	output break_o;
	output imem_addr_ox0x;
	output imem_addr_ox1x;
	output imem_addr_ox2x;
	output imem_addr_ox3x;
	output imem_addr_ox4x;
	output imem_addr_ox5x;
	output imem_addr_ox6x;
	output imem_addr_ox7x;
	output imem_addr_ox8x;
	output imem_addr_ox9x;
	output imem_addr_ox10x;
	output imem_addr_ox11x;
	output imem_addr_ox12x;
	output imem_addr_ox13x;
	output imem_addr_ox14x;
	output imem_addr_ox15x;
	output imem_addr_ox16x;
	output imem_addr_ox17x;
	output imem_addr_ox18x;
	output imem_addr_ox19x;
	output imem_addr_ox20x;
	output imem_addr_ox21x;
	output imem_addr_ox22x;
	output imem_addr_ox23x;
	output imem_addr_ox24x;
	output imem_addr_ox25x;
	output imem_addr_ox26x;
	output imem_addr_ox27x;
	output imem_addr_ox28x;
	output imem_addr_ox29x;
	output imem_addr_ox30x;
	output imem_addr_ox31x;
	output imem_cti_ox0x;
	output imem_cti_ox1x;
	output imem_cti_ox2x;
	output imem_cyc_o;
	output imem_stb_o;
	output dmem_addr_ox0x;
	output dmem_addr_ox1x;
	output dmem_addr_ox2x;
	output dmem_addr_ox3x;
	output dmem_addr_ox4x;
	output dmem_addr_ox5x;
	output dmem_addr_ox6x;
	output dmem_addr_ox7x;
	output dmem_addr_ox8x;
	output dmem_addr_ox9x;
	output dmem_addr_ox10x;
	output dmem_addr_ox11x;
	output dmem_addr_ox12x;
	output dmem_addr_ox13x;
	output dmem_addr_ox14x;
	output dmem_addr_ox15x;
	output dmem_addr_ox16x;
	output dmem_addr_ox17x;
	output dmem_addr_ox18x;
	output dmem_addr_ox19x;
	output dmem_addr_ox20x;
	output dmem_addr_ox21x;
	output dmem_addr_ox22x;
	output dmem_addr_ox23x;
	output dmem_addr_ox24x;
	output dmem_addr_ox25x;
	output dmem_addr_ox26x;
	output dmem_addr_ox27x;
	output dmem_addr_ox28x;
	output dmem_addr_ox29x;
	output dmem_addr_ox30x;
	output dmem_addr_ox31x;
	output dmem_dat_ox0x;
	output dmem_dat_ox1x;
	output dmem_dat_ox2x;
	output dmem_dat_ox3x;
	output dmem_dat_ox4x;
	output dmem_dat_ox5x;
	output dmem_dat_ox6x;
	output dmem_dat_ox7x;
	output dmem_dat_ox8x;
	output dmem_dat_ox9x;
	output dmem_dat_ox10x;
	output dmem_dat_ox11x;
	output dmem_dat_ox12x;
	output dmem_dat_ox13x;
	output dmem_dat_ox14x;
	output dmem_dat_ox15x;
	output dmem_dat_ox16x;
	output dmem_dat_ox17x;
	output dmem_dat_ox18x;
	output dmem_dat_ox19x;
	output dmem_dat_ox20x;
	output dmem_dat_ox21x;
	output dmem_dat_ox22x;
	output dmem_dat_ox23x;
	output dmem_dat_ox24x;
	output dmem_dat_ox25x;
	output dmem_dat_ox26x;
	output dmem_dat_ox27x;
	output dmem_dat_ox28x;
	output dmem_dat_ox29x;
	output dmem_dat_ox30x;
	output dmem_dat_ox31x;
	output dmem_cti_ox0x;
	output dmem_cti_ox1x;
	output dmem_cti_ox2x;
	output dmem_cyc_o;
	output dmem_stb_o;
	output dmem_we_o;
	output dmem_sel_ox0x;
	output dmem_sel_ox1x;
	output dmem_sel_ox2x;
	output dmem_sel_ox3x;

	input [127 : 0] sk /* synthesis noprune */;


	wire gnd, vcc, g139, g127, g3893, g140, g3894, g274, g3895, g3882, g3896;
	wire g363, g3897, g3871, g3898, g452, g3899, g3860, g3900, g540, g3901, g585;
	wire g3902, g3849, g3903, g681, g3904, g728, g3905, g775, g3906, g822, g3907;
	wire g869, g3908, g917, g3909, g962, g3910, g1007, g3911, g1052, g3912, g1097;
	wire g3913, g1142, g3914, g1187, g3915, g1232, g3916, g1277, g3917, g1322, g3918;
	wire g1367, g3919, g1412, g3920, g1457, g3921, g1501, g3922, g1546, g3923, g1591;
	wire g3924, g1609, g1608, g3925, g1621, g3926, g1633, g3927, g1645, g3928, g1657;
	wire g3929, g1669, g3930, g1681, g3931, g1693, g3932, g1708, g3933, g1721, g3934;
	wire g1734, g3935, g1747, g3936, g1760, g3937, g1773, g3938, g1786, g3939, g1799;
	wire g3940, g1813, g3941, g1826, g3942, g1839, g3943, g1852, g3944, g1865, g3945;
	wire g1878, g3946, g1891, g3947, g1904, g3948, g1918, g3949, g1931, g3950, g1944;
	wire g3951, g1957, g3952, g1970, g3953, g1983, g3954, g1996, g3955, g2009, g3956;
	wire g2015, g2014, g3957, g2016, g3958, g2017, g3959, g2018, g3960, g2059, g2058;
	wire g3961, g2063, g3962, g2064, g3963, g3964, g3965, g3966, g3967, g3968, g84;
	wire g3969, g3970, g3971, g3972, g3973, g3974, g3975, g3976, g93, g94, g95;
	wire g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106;
	wire g3977, g3978, g3979, g3980, g111, g112, g113, g114, g115, g116, g117;
	wire g118, g119, g120, g121, g122, g123, g124, g125, g130, g131, g132;
	wire g133, g134, g135, g136, g137, g138, g2069, g3981, g3982, g2140, g3777;
	wire g3983, g2142, g3984, g2144, g3985, g2145, g3986, g3987, g3988, g149, g2146;
	wire g3989, g2148, g3990, g2150, g3991, g2151, g3992, g154, g2152, g3993, g2153;
	wire g3994, g2155, g3995, g2157, g3996, g159, g2158, g3997, g2159, g3998, g2160;
	wire g3999, g2161, g4000, g164, g4001, g4002, g167, g2162, g4003, g2164, g4004;
	wire g2166, g4005, g2168, g4006, g172, g2169, g4007, g2170, g4008, g2171, g4009;
	wire g2172, g4010, g177, g2173, g4011, g2174, g4012, g2175, g4013, g2176, g4014;
	wire g182, g2177, g4015, g2178, g4016, g2179, g4017, g186, g187, g188, g2210;
	wire g4018, g4019, g4020, g4021, g193, g4022, g4023, g4024, g4025, g198, g4026;
	wire g4027, g4028, g4029, g203, g4030, g4031, g4032, g4033, g208, g209, g4034;
	wire g4035, g4036, g4037, g214, g4038, g4039, g4040, g4041, g219, g4042, g4043;
	wire g4044, g4045, g224, g4046, g4047, g4048, g228, g229, g230, g231, g2229;
	wire g4049, g4050, g4051, g4052, g236, g4053, g4054, g4055, g4056, g241, g4057;
	wire g4058, g4059, g4060, g246, g4061, g4062, g4063, g4064, g251, g252, g4065;
	wire g4066, g4067, g4068, g257, g4069, g4070, g4071, g261, g4072, g4073, g4074;
	wire g4075, g266, g4076, g4077, g4078, g4079, g271, g272, g273, g2235, g4080;
	wire g2256, g4081, g4082, g4083, g4084, g280, g4085, g4086, g4087, g4088, g285;
	wire g4089, g4090, g4091, g4092, g290, g4093, g4094, g4095, g4096, g295, g296;
	wire g4097, g4098, g4099, g4100, g301, g4101, g4102, g4103, g305, g4104, g4105;
	wire g4106, g4107, g310, g4108, g4109, g4110, g4111, g315, g316, g317, g4112;
	wire g2263, g4113, g320, g2282, g4114, g4115, g4116, g4117, g325, g4118, g4119;
	wire g4120, g4121, g330, g4122, g4123, g4124, g4125, g335, g4126, g4127, g4128;
	wire g4129, g340, g341, g4130, g4131, g4132, g4133, g346, g4134, g4135, g4136;
	wire g350, g4137, g4138, g4139, g4140, g355, g4141, g4142, g4143, g4144, g360;
	wire g361, g362, g4145, g2288, g4146, g2304, g4147, g4148, g4149, g4150, g370;
	wire g4151, g4152, g4153, g4154, g375, g4155, g4156, g4157, g4158, g380, g4159;
	wire g4160, g4161, g4162, g385, g386, g4163, g4164, g4165, g4166, g391, g4167;
	wire g4168, g4169, g395, g4170, g4171, g4172, g4173, g400, g4174, g4175, g4176;
	wire g4177, g405, g406, g407, g2311, g4178, g409, g2328, g4179, g4180, g4181;
	wire g4182, g414, g4183, g4184, g4185, g4186, g419, g4187, g4188, g4189, g4190;
	wire g424, g4191, g4192, g4193, g4194, g429, g430, g4195, g4196, g4197, g4198;
	wire g435, g4199, g4200, g4201, g439, g4202, g4203, g4204, g4205, g444, g4206;
	wire g4207, g4208, g4209, g449, g450, g451, g2337, g4210, g3676, g4211, g4212;
	wire g4213, g4214, g458, g4215, g4216, g4217, g4218, g463, g4219, g4220, g4221;
	wire g4222, g468, g4223, g4224, g4225, g4226, g473, g474, g4227, g4228, g4229;
	wire g4230, g479, g4231, g4232, g4233, g483, g4234, g4235, g4236, g4237, g488;
	wire g4238, g4239, g4240, g4241, g493, g494, g495, g2361, g4242, g4243, g497;
	wire g2378, g4244, g4245, g4246, g4247, g502, g4248, g4249, g4250, g4251, g507;
	wire g4252, g4253, g4254, g4255, g512, g4256, g4257, g4258, g4259, g517, g518;
	wire g4260, g4261, g4262, g4263, g523, g4264, g4265, g4266, g527, g4267, g4268;
	wire g4269, g4270, g532, g4271, g4272, g4273, g4274, g537, g538, g539, g2388;
	wire g4275, g542, g2407, g4276, g4277, g4278, g4279, g547, g4280, g4281, g4282;
	wire g4283, g552, g4284, g4285, g4286, g4287, g557, g4288, g4289, g4290, g4291;
	wire g562, g563, g4292, g4293, g4294, g4295, g568, g4296, g4297, g4298, g572;
	wire g4299, g4300, g4301, g4302, g577, g4303, g4304, g4305, g4306, g582, g583;
	wire g584, g4307, g2415, g4308, g2431, g4309, g4310, g4311, g4312, g592, g4313;
	wire g4314, g4315, g4316, g597, g4317, g4318, g4319, g4320, g602, g4321, g4322;
	wire g4323, g4324, g607, g608, g4325, g4326, g4327, g4328, g613, g4329, g4330;
	wire g4331, g617, g4332, g4333, g4334, g4335, g622, g4336, g4337, g4338, g4339;
	wire g627, g628, g629, g3627, g4340, g2454, g4341, g4342, g4343, g4344, g635;
	wire g4345, g4346, g4347, g4348, g640, g4349, g4350, g4351, g4352, g645, g4353;
	wire g4354, g4355, g4356, g650, g651, g4357, g4358, g4359, g4360, g656, g4361;
	wire g4362, g4363, g660, g4364, g4365, g4366, g4367, g665, g4368, g4369, g4370;
	wire g4371, g670, g671, g672, g673, g674, g675, g676, g4372, g4373, g679;
	wire g680, g2473, g4374, g4375, g4376, g4377, g686, g4378, g4379, g4380, g4381;
	wire g691, g4382, g4383, g4384, g4385, g696, g4386, g4387, g4388, g4389, g701;
	wire g702, g4390, g4391, g4392, g4393, g707, g4394, g4395, g4396, g711, g4397;
	wire g4398, g4399, g4400, g716, g4401, g4402, g4403, g4404, g721, g722, g723;
	wire g2479, g4405, g725, g4406, g727, g2495, g4407, g4408, g4409, g4410, g733;
	wire g4411, g4412, g4413, g4414, g738, g4415, g4416, g4417, g4418, g743, g4419;
	wire g4420, g4421, g4422, g748, g749, g4423, g4424, g4425, g4426, g754, g4427;
	wire g4428, g4429, g758, g4430, g4431, g4432, g4433, g763, g4434, g4435, g4436;
	wire g4437, g768, g769, g770, g2504, g4438, g772, g4439, g774, g2520, g4440;
	wire g4441, g4442, g4443, g780, g4444, g4445, g4446, g4447, g785, g4448, g4449;
	wire g4450, g4451, g790, g4452, g4453, g4454, g4455, g795, g796, g4456, g4457;
	wire g4458, g4459, g801, g4460, g4461, g4462, g805, g4463, g4464, g4465, g4466;
	wire g810, g4467, g4468, g4469, g4470, g815, g816, g817, g2526, g4471, g819;
	wire g4472, g821, g2542, g4473, g4474, g4475, g4476, g827, g4477, g4478, g4479;
	wire g4480, g832, g4481, g4482, g4483, g4484, g837, g4485, g4486, g4487, g4488;
	wire g842, g843, g4489, g4490, g4491, g4492, g848, g4493, g4494, g4495, g852;
	wire g4496, g4497, g4498, g4499, g857, g4500, g4501, g4502, g4503, g862, g863;
	wire g864, g2548, g4504, g866, g4505, g868, g3539, g4506, g4507, g4508, g4509;
	wire g874, g4510, g4511, g4512, g4513, g879, g4514, g4515, g4516, g4517, g884;
	wire g4518, g4519, g4520, g4521, g889, g890, g4522, g4523, g4524, g4525, g895;
	wire g4526, g4527, g4528, g899, g4529, g4530, g4531, g4532, g904, g4533, g4534;
	wire g4535, g4536, g909, g910, g911, g2569, g4537, g3134, g3135, g913, g914;
	wire g915, g916, g3515, g4538, g4539, g4540, g4541, g922, g4542, g4543, g4544;
	wire g4545, g927, g4546, g4547, g4548, g4549, g932, g4550, g4551, g4552, g4553;
	wire g937, g938, g4554, g4555, g4556, g4557, g943, g4558, g4559, g4560, g947;
	wire g4561, g4562, g4563, g4564, g952, g4565, g4566, g4567, g4568, g957, g958;
	wire g959, g2589, g4569, g961, g3491, g4570, g4571, g4572, g4573, g967, g4574;
	wire g4575, g4576, g4577, g972, g4578, g4579, g4580, g4581, g977, g4582, g4583;
	wire g4584, g4585, g982, g983, g4586, g4587, g4588, g4589, g988, g4590, g4591;
	wire g4592, g992, g4593, g4594, g4595, g4596, g997, g4597, g4598, g4599, g4600;
	wire g1002, g1003, g1004, g2607, g4601, g1006, g3468, g4602, g4603, g4604, g4605;
	wire g1012, g4606, g4607, g4608, g4609, g1017, g4610, g4611, g4612, g4613, g1022;
	wire g4614, g4615, g4616, g4617, g1027, g1028, g4618, g4619, g4620, g4621, g1033;
	wire g4622, g4623, g4624, g1037, g4625, g4626, g4627, g4628, g1042, g4629, g4630;
	wire g4631, g4632, g1047, g1048, g1049, g2624, g4633, g1051, g3444, g4634, g4635;
	wire g4636, g4637, g1057, g4638, g4639, g4640, g4641, g1062, g4642, g4643, g4644;
	wire g4645, g1067, g4646, g4647, g4648, g4649, g1072, g1073, g4650, g4651, g4652;
	wire g4653, g1078, g4654, g4655, g4656, g1082, g4657, g4658, g4659, g4660, g1087;
	wire g4661, g4662, g4663, g4664, g1092, g1093, g1094, g2641, g4665, g1096, g3420;
	wire g4666, g4667, g4668, g4669, g1102, g4670, g4671, g4672, g4673, g1107, g4674;
	wire g4675, g4676, g4677, g1112, g4678, g4679, g4680, g4681, g1117, g1118, g4682;
	wire g4683, g4684, g4685, g1123, g4686, g4687, g4688, g1127, g4689, g4690, g4691;
	wire g4692, g1132, g4693, g4694, g4695, g4696, g1137, g1138, g1139, g2659, g4697;
	wire g1141, g3836, g3397, g4698, g4699, g4700, g4701, g1147, g4702, g4703, g4704;
	wire g4705, g1152, g4706, g4707, g4708, g4709, g1157, g4710, g4711, g4712, g4713;
	wire g1162, g1163, g4714, g4715, g4716, g4717, g1168, g4718, g4719, g4720, g1172;
	wire g4721, g4722, g4723, g4724, g1177, g4725, g4726, g4727, g4728, g1182, g1183;
	wire g1184, g2679, g4729, g1186, g3373, g4730, g4731, g4732, g4733, g1192, g4734;
	wire g4735, g4736, g4737, g1197, g4738, g4739, g4740, g4741, g1202, g4742, g4743;
	wire g4744, g4745, g1207, g1208, g4746, g4747, g4748, g4749, g1213, g4750, g4751;
	wire g4752, g1217, g4753, g4754, g4755, g4756, g1222, g4757, g4758, g4759, g4760;
	wire g1227, g1228, g1229, g2698, g4761, g1231, g3349, g4762, g4763, g4764, g4765;
	wire g1237, g4766, g4767, g4768, g4769, g1242, g4770, g4771, g4772, g4773, g1247;
	wire g4774, g4775, g4776, g4777, g1252, g1253, g4778, g4779, g4780, g4781, g1258;
	wire g4782, g4783, g4784, g1262, g4785, g4786, g4787, g4788, g1267, g4789, g4790;
	wire g4791, g4792, g1272, g1273, g1274, g2714, g4793, g1276, g3325, g4794, g4795;
	wire g4796, g4797, g1282, g4798, g4799, g4800, g4801, g1287, g4802, g4803, g4804;
	wire g4805, g1292, g4806, g4807, g4808, g4809, g1297, g1298, g4810, g4811, g4812;
	wire g4813, g1303, g4814, g4815, g4816, g1307, g4817, g4818, g4819, g4820, g1312;
	wire g4821, g4822, g4823, g4824, g1317, g1318, g1319, g2733, g4825, g1321, g3302;
	wire g4826, g4827, g4828, g4829, g1327, g4830, g4831, g4832, g4833, g1332, g4834;
	wire g4835, g4836, g4837, g1337, g4838, g4839, g4840, g4841, g1342, g1343, g4842;
	wire g4843, g4844, g4845, g1348, g4846, g4847, g4848, g1352, g4849, g4850, g4851;
	wire g4852, g1357, g4853, g4854, g4855, g4856, g1362, g1363, g1364, g2750, g4857;
	wire g1366, g3823, g3278, g4858, g4859, g4860, g4861, g1372, g4862, g4863, g4864;
	wire g4865, g1377, g4866, g4867, g4868, g4869, g1382, g4870, g4871, g4872, g4873;
	wire g1387, g1388, g4874, g4875, g4876, g4877, g1393, g4878, g4879, g4880, g1397;
	wire g4881, g4882, g4883, g4884, g1402, g4885, g4886, g4887, g4888, g1407, g1408;
	wire g1409, g2769, g4889, g1411, g2787, g4890, g4891, g4892, g4893, g1417, g4894;
	wire g4895, g4896, g4897, g1422, g4898, g4899, g4900, g4901, g1427, g4902, g4903;
	wire g4904, g4905, g1432, g1433, g4906, g4907, g4908, g4909, g1438, g4910, g4911;
	wire g4912, g1442, g4913, g4914, g4915, g4916, g1447, g4917, g4918, g4919, g4920;
	wire g1452, g1453, g1454, g2793, g4921, g1456, g2805, g4922, g4923, g4924, g4925;
	wire g1462, g4926, g4927, g4928, g4929, g1467, g4930, g4931, g4932, g4933, g1472;
	wire g4934, g4935, g4936, g4937, g1477, g1478, g4938, g4939, g4940, g4941, g1483;
	wire g4942, g4943, g4944, g1487, g4945, g4946, g4947, g4948, g1492, g4949, g4950;
	wire g4951, g4952, g1497, g1498, g1499, g2810, g4953, g3118, g2821, g4954, g4955;
	wire g4956, g4957, g1506, g4958, g4959, g4960, g4961, g1511, g4962, g4963, g4964;
	wire g4965, g1516, g4966, g4967, g4968, g4969, g1521, g1522, g4970, g4971, g4972;
	wire g4973, g1527, g4974, g4975, g4976, g1531, g4977, g4978, g4979, g4980, g1536;
	wire g4981, g4982, g4983, g4984, g1541, g1542, g1543, g2825, g4985, g1545, g2830;
	wire g4986, g2841, g4987, g4988, g4989, g4990, g1552, g4991, g4992, g4993, g4994;
	wire g1557, g4995, g4996, g4997, g4998, g1562, g4999, g5000, g5001, g5002, g1567;
	wire g1568, g5003, g5004, g5005, g5006, g1573, g5007, g5008, g5009, g1577, g5010;
	wire g5011, g5012, g5013, g1582, g5014, g5015, g5016, g5017, g1587, g1588, g1589;
	wire g1590, g1592, g1593, g1594, g1595, g1596, g1597, g1598, g1599, g1600, g1601;
	wire g1602, g1603, g1604, g1605, g1606, g1607, g1610, g1611, g1612, g1613, g1614;
	wire g1615, g1616, g1617, g1618, g1619, g1620, g1622, g1623, g1624, g1625, g1626;
	wire g1627, g1628, g1629, g1630, g1631, g1632, g1634, g1635, g1636, g1637, g1638;
	wire g1639, g1640, g1641, g1642, g1643, g1644, g1646, g1647, g1648, g1649, g1650;
	wire g1651, g1652, g1653, g1654, g1655, g1656, g1658, g1659, g1660, g1661, g1662;
	wire g1663, g1664, g1665, g1666, g1667, g1668, g1670, g1671, g1672, g1673, g1674;
	wire g1675, g1676, g1677, g1678, g1679, g1680, g1682, g1683, g1684, g1685, g1686;
	wire g1687, g1688, g1689, g1690, g1691, g1692, g1694, g1695, g1696, g1697, g1698;
	wire g1699, g1700, g1701, g1702, g1703, g1704, g1705, g1706, g1707, g1709, g1710;
	wire g1711, g1712, g1713, g1714, g1715, g1716, g1717, g1718, g1719, g1720, g1722;
	wire g1723, g1724, g1725, g1726, g1727, g1728, g1729, g1730, g1731, g1732, g1733;
	wire g1735, g1736, g1737, g1738, g1739, g1740, g1741, g1742, g1743, g1744, g1745;
	wire g1746, g1748, g1749, g1750, g1751, g1752, g1753, g1754, g1755, g1756, g1757;
	wire g1758, g1759, g1761, g1762, g1763, g1764, g1765, g1766, g1767, g1768, g1769;
	wire g1770, g1771, g1772, g1774, g1775, g1776, g1777, g1778, g1779, g1780, g1781;
	wire g1782, g1783, g1784, g1785, g1787, g1788, g1789, g1790, g1791, g1792, g1793;
	wire g1794, g1795, g1796, g1797, g1798, g1800, g1801, g1802, g1803, g1804, g1805;
	wire g1806, g1807, g1808, g1809, g1810, g1811, g1812, g1814, g1815, g1816, g1817;
	wire g1818, g1819, g1820, g1821, g1822, g1823, g1824, g1825, g1827, g1828, g1829;
	wire g1830, g1831, g1832, g1833, g1834, g1835, g1836, g1837, g1838, g1840, g1841;
	wire g1842, g1843, g1844, g1845, g1846, g1847, g1848, g1849, g1850, g1851, g1853;
	wire g1854, g1855, g1856, g1857, g1858, g1859, g1860, g1861, g1862, g1863, g1864;
	wire g1866, g1867, g1868, g1869, g1870, g1871, g1872, g1873, g1874, g1875, g1876;
	wire g1877, g1879, g1880, g1881, g1882, g1883, g1884, g1885, g1886, g1887, g1888;
	wire g1889, g1890, g1892, g1893, g1894, g1895, g1896, g1897, g1898, g1899, g1900;
	wire g1901, g1902, g1903, g1905, g1906, g1907, g1908, g1909, g1910, g1911, g1912;
	wire g1913, g1914, g1915, g1916, g1917, g1919, g1920, g1921, g1922, g1923, g1924;
	wire g1925, g1926, g1927, g1928, g1929, g1930, g1932, g1933, g1934, g1935, g1936;
	wire g1937, g1938, g1939, g1940, g1941, g1942, g1943, g1945, g1946, g1947, g1948;
	wire g1949, g1950, g1951, g1952, g1953, g1954, g1955, g1956, g1958, g1959, g1960;
	wire g1961, g1962, g1963, g1964, g1965, g1966, g1967, g1968, g1969, g1971, g1972;
	wire g1973, g1974, g1975, g1976, g1977, g1978, g1979, g1980, g1981, g1982, g1984;
	wire g1985, g1986, g1987, g1988, g1989, g1990, g1991, g1992, g1993, g1994, g1995;
	wire g1997, g1998, g1999, g2000, g2001, g2002, g2003, g2004, g2005, g2006, g2007;
	wire g2008, g2010, g2011, g2012, g2013, g2020, g2021, g2022, g2024, g2025, g2917;
	wire g5018, g2027, g2028, g2029, g2030, g2031, g2032, g2033, g2034, g2921, g2918;
	wire g5019, g2036, g2037, g2924, g2922, g5020, g2039, g2040, g2041, g2042, g2043;
	wire g2044, g2045, g2046, g2047, g2048, g2049, g2050, g2051, g2052, g2053, g2054;
	wire g2925, g5021, g2056, g2057, g2926, g5022, g2061, g2062, g2065, g2927, g5023;
	wire g2067, g2068, g2072, g2075, g2078, g2973, g5024, g2082, g2087, g2092, g2097;
	wire g2102, g2103, g2107, g2112, g2117, g2122, g2123, g3801, g3788, g2126, g2127;
	wire g5025, g5026, g2130, g2131, g2132, g2133, g2139, g2141, g2143, g2147, g2149;
	wire g2154, g2156, g2163, g2165, g2167, g2180, g2181, g2182, g2183, g2184, g2185;
	wire g2186, g2187, g2188, g2189, g2190, g2191, g2192, g2193, g2194, g2195, g2196;
	wire g2197, g2198, g2199, g2200, g2201, g2202, g2203, g3147, g2204, g2205, g2206;
	wire g2207, g2208, g2209, g2211, g2212, g2213, g2214, g2215, g2216, g2217, g2218;
	wire g2219, g2220, g2221, g2222, g2223, g2224, g3764, g2225, g2226, g2227, g2228;
	wire g2230, g3056, g5027, g2232, g2233, g2234, g2236, g2237, g2238, g2239, g2240;
	wire g2241, g2242, g2243, g2244, g2245, g2246, g2247, g2248, g2249, g2250, g2251;
	wire g3751, g2252, g2253, g2254, g2255, g2257, g3057, g5028, g2259, g2260, g2261;
	wire g2262, g2264, g2265, g2266, g2267, g3125, g2268, g2269, g2270, g2271, g2272;
	wire g2273, g2274, g2275, g2276, g3738, g2277, g2278, g2279, g2280, g2281, g2283;
	wire g3058, g5029, g2285, g2286, g2287, g2290, g2291, g2292, g2293, g2294, g2295;
	wire g2296, g2297, g2298, g2299, g2300, g3725, g2301, g2302, g2303, g2305, g3060;
	wire g5030, g2307, g2308, g2309, g2310, g2313, g2314, g2315, g2316, g2317, g2318;
	wire g2319, g2320, g2321, g2322, g2323, g2324, g3712, g2325, g2326, g2327, g2329;
	wire g2330, g2331, g2332, g3066, g5031, g2334, g2335, g2336, g2338, g2339, g2341;
	wire g2342, g2343, g2344, g2345, g2346, g2347, g2348, g2349, g2350, g2351, g2352;
	wire g2353, g2354, g2355, g2356, g3068, g5032, g2358, g2359, g2360, g2362, g2363;
	wire g2364, g2366, g2367, g2368, g2369, g2370, g2371, g2372, g2373, g2374, g2375;
	wire g2376, g3663, g2377, g2379, g2380, g2381, g2382, g3070, g5033, g2384, g2385;
	wire g2386, g2387, g2389, g2390, g2392, g2393, g2394, g2395, g2396, g2397, g2398;
	wire g2399, g2400, g2401, g2402, g2403, g2404, g2405, g3650, g2406, g2408, g2409;
	wire g2410, g2411, g2412, g3073, g5034, g2414, g2416, g2417, g2419, g2420, g2421;
	wire g2422, g2423, g2424, g2425, g2426, g2427, g2428, g2429, g3638, g2430, g3075;
	wire g5035, g2433, g2434, g2435, g2436, g2437, g2438, g2440, g2441, g2442, g2443;
	wire g2444, g2445, g2446, g2447, g2448, g2449, g2450, g2451, g2452, g3614, g2453;
	wire g2455, g2456, g2458, g2459, g2460, g2461, g2462, g2463, g2464, g2465, g2466;
	wire g2467, g2468, g2469, g2470, g2471, g3601, g2472, g2474, g2475, g3239, g5036;
	wire g2477, g2478, g2480, g2481, g2483, g2484, g2485, g2486, g2487, g2488, g2489;
	wire g2490, g2491, g2492, g2493, g3588, g2494, g2496, g2497, g2498, g3080, g5037;
	wire g2500, g2501, g2502, g2503, g2505, g2506, g2508, g2509, g2510, g2511, g2512;
	wire g2513, g2514, g2515, g2516, g2517, g2518, g3575, g2519, g2521, g2522, g3226;
	wire g5038, g2524, g2525, g2527, g2528, g3119, g2530, g2531, g2532, g2533, g2534;
	wire g2535, g2536, g2537, g2538, g2539, g2540, g3562, g2541, g2543, g3083, g5039;
	wire g2545, g2546, g2547, g2549, g2550, g3137, g3138, g2552, g2553, g2554, g2555;
	wire g2556, g2557, g2558, g2559, g2560, g2561, g3550, g2562, g2563, g2564, g2565;
	wire g3087, g5040, g2567, g2568, g2571, g2572, g2573, g2574, g2575, g2576, g2577;
	wire g2578, g2579, g2580, g2581, g2582, g3526, g2583, g2584, g2585, g2586, g3213;
	wire g5041, g2588, g2591, g2592, g2593, g2594, g2595, g2596, g2597, g3502, g2598;
	wire g2599, g2600, g2601, g2602, g2603, g2604, g3200, g5042, g2606, g2609, g2610;
	wire g2611, g2612, g2613, g2614, g2615, g2616, g2617, g3479, g2618, g2619, g2620;
	wire g2621, g3091, g5043, g2623, g3127, g2626, g2627, g2628, g2629, g2630, g2631;
	wire g2632, g2633, g2634, g3455, g2635, g2636, g2637, g2638, g3093, g5044, g2640;
	wire g2643, g2644, g2645, g2646, g2647, g2648, g2649, g2650, g2651, g2652, g3431;
	wire g2653, g2654, g2655, g2656, g3187, g5045, g2658, g2661, g3126, g2662, g2663;
	wire g2664, g2665, g2666, g2667, g2668, g2669, g2670, g2671, g3408, g2672, g2673;
	wire g2674, g2675, g2676, g3098, g5046, g2678, g2681, g2682, g2683, g2684, g2685;
	wire g2686, g2687, g2688, g2689, g3384, g2690, g2691, g2692, g2693, g2694, g2695;
	wire g3174, g5047, g2697, g2700, g2701, g2702, g2703, g2704, g2705, g2706, g2707;
	wire g2708, g3360, g2709, g2710, g2711, g3101, g5048, g2713, g2716, g2717, g2718;
	wire g2719, g2720, g2721, g2722, g2723, g2724, g2725, g3336, g2726, g2727, g2728;
	wire g2729, g2730, g3103, g5049, g2732, g2735, g2736, g2737, g2738, g2739, g2740;
	wire g2741, g2742, g2743, g2744, g3313, g2745, g2746, g2747, g3161, g5050, g2749;
	wire g2752, g2753, g2754, g2755, g2756, g2757, g2758, g2759, g2760, g2761, g2762;
	wire g3289, g2763, g2764, g2765, g2766, g3148, g5051, g2768, g2770, g2772, g2773;
	wire g2774, g2775, g2776, g2777, g2778, g2779, g2780, g3265, g2781, g2782, g2783;
	wire g2784, g2785, g2786, g2788, g2789, g2790, g3107, g5052, g2792, g2795, g2796;
	wire g2797, g2798, g2799, g3116, g2800, g2801, g2802, g2803, g2804, g2806, g2807;
	wire g3109, g5053, g2809, g2812, g2813, g2814, g2815, g3131, g3132, g2816, g2817;
	wire g2818, g2819, g2820, g2822, g2823, g3111, g5054, g3252, g2826, g3112, g5055;
	wire g2828, g2829, g2832, g2833, g2834, g2835, g2836, g2837, g2838, g2839, g3140;
	wire g2840, g2842, g2843, g2844, g2845, g2846, g2847, g2848, g2849, g2850, g2851;
	wire g2852, g2853, g2854, g2855, g2856, g2857, g2858, g2859, g2860, g2861, g2862;
	wire g2863, g2864, g2865, g2866, g2867, g2868, g2869, g2870, g2871, g2872, g2873;
	wire g2874, g2875, g2876, g2877, g2878, g2879, g2880, g2881, g2882, g2883, g2884;
	wire g2885, g2886, g2887, g2888, g2889, g2890, g2891, g2892, g2893, g2894, g2895;
	wire g2896, g2897, g2898, g2899, g2900, g2901, g2902, g2903, g2904, g2905, g2906;
	wire g2907, g2908, g2909, g2910, g2911, g2912, g2913, g3114, g5056, g2915, g2916;
	wire g2919, g2920, g2923, g2928, g2929, g2930, g2931, g3139, g2932, g2933, g2934;
	wire g2935, g2936, g2937, g2938, g2939, g2940, g2941, g2942, g2943, g2944, g2945;
	wire g2946, g2947, g2948, g2949, g2950, g2951, g2952, g2953, g2954, g2955, g2956;
	wire g2957, g2958, g2959, g2960, g2961, g2962, g2963, g2964, g2965, g2966, g2967;
	wire g2968, g3115, g5057, g3120, g3121, g2970, g2971, g3122, g2972, g2974, g2975;
	wire g2976, g2977, g2978, g2979, g2980, g2981, g2982, g2983, g2984, g2985, g2986;
	wire g2987, g2988, g2989, g2990, g2991, g2992, g2993, g2994, g2995, g2996, g2997;
	wire g2998, g2999, g3000, g3001, g3002, g3003, g3004, g3005, g3006, g3007, g3008;
	wire g3009, g3010, g3011, g3012, g3013, g3014, g3015, g3016, g3017, g3018, g3019;
	wire g3020, g3021, g3022, g3023, g3024, g3124, g3025, g3026, g3027, g3028, g3029;
	wire g3030, g3031, g3032, g3033, g3034, g3035, g3036, g3037, g3038, g3039, g3040;
	wire g3041, g3042, g3043, g3044, g3045, g3046, g3047, g3048, g3049, g3050, g3051;
	wire g3052, g3053, g3054, g3055, g3059, g3061, g3062, g3063, g3064, g3065, g3067;
	wire g3069, g3071, g3072, g3074, g3076, g3077, g3078, g3079, g3081, g3082, g3084;
	wire g3085, g3086, g3088, g3089, g3090, g3092, g3094, g3095, g3096, g3097, g3099;
	wire g3100, g3102, g3104, g3105, g3106, g3108, g3110, g3113, g3117, g3123, g3128;
	wire g3129, g3130, g3133, g3136, g3141, g3142, g3143, g3144, g3145, g3146, g3149;
	wire g3150, g3151, g3154, g3152, g3153, g3157, g3158, g3155, g3156, g3159, g3160;
	wire g3162, g3163, g3164, g3167, g3165, g3166, g3170, g3171, g3168, g3169, g3172;
	wire g3173, g3175, g3176, g3177, g3180, g3178, g3179, g3183, g3184, g3181, g3182;
	wire g3185, g3186, g3188, g3189, g3190, g3193, g3191, g3192, g3196, g3197, g3194;
	wire g3195, g3198, g3199, g3201, g3202, g3203, g3206, g3204, g3205, g3209, g3210;
	wire g3207, g3208, g3211, g3212, g3214, g3215, g3216, g3219, g3217, g3218, g3222;
	wire g3223, g3220, g3221, g3224, g3225, g3227, g3228, g3229, g3232, g3230, g3231;
	wire g3235, g3236, g3233, g3234, g3237, g3238, g3240, g3241, g3242, g3245, g3243;
	wire g3244, g3248, g3249, g3246, g3247, g3250, g3251, g3253, g3254, g3255, g3258;
	wire g3256, g3257, g3261, g3262, g3259, g3260, g3263, g3264, g3266, g3267, g3268;
	wire g3271, g3269, g3270, g3274, g3275, g3272, g3273, g3276, g3277, g3279, g3280;
	wire g3281, g3284, g3282, g3283, g3285, g3286, g3287, g3288, g3290, g3291, g3292;
	wire g3295, g3293, g3294, g3298, g3299, g3296, g3297, g3300, g3301, g3303, g3304;
	wire g3305, g3308, g3306, g3307, g3309, g3310, g3311, g3312, g3314, g3315, g3316;
	wire g3319, g3317, g3318, g3322, g3320, g3321, g3323, g3324, g3326, g3327, g3328;
	wire g3331, g3329, g3330, g3332, g3333, g3334, g3335, g3337, g3338, g3339, g3342;
	wire g3340, g3341, g3345, g3346, g3343, g3344, g3347, g3348, g3350, g3351, g3352;
	wire g3355, g3353, g3354, g3356, g3357, g3358, g3359, g3361, g3362, g3363, g3366;
	wire g3364, g3365, g3369, g3370, g3367, g3368, g3371, g3372, g3374, g3375, g3376;
	wire g3379, g3377, g3378, g3380, g3381, g3382, g3383, g3385, g3386, g3387, g3390;
	wire g3388, g3389, g3393, g3394, g3391, g3392, g3395, g3396, g3398, g3399, g3400;
	wire g3403, g3401, g3402, g3404, g3405, g3406, g3407, g3409, g3410, g3411, g3414;
	wire g3412, g3413, g3417, g3415, g3416, g3418, g3419, g3421, g3422, g3423, g3426;
	wire g3424, g3425, g3427, g3428, g3429, g3430, g3432, g3433, g3434, g3437, g3435;
	wire g3436, g3440, g3441, g3438, g3439, g3442, g3443, g3445, g3446, g3447, g3450;
	wire g3448, g3449, g3451, g3452, g3453, g3454, g3456, g3457, g3458, g3461, g3459;
	wire g3460, g3464, g3465, g3462, g3463, g3466, g3467, g3469, g3470, g3471, g3474;
	wire g3472, g3473, g3475, g3476, g3477, g3478, g3480, g3481, g3482, g3485, g3483;
	wire g3484, g3488, g3486, g3487, g3489, g3490, g3492, g3493, g3494, g3497, g3495;
	wire g3496, g3498, g3499, g3500, g3501, g3503, g3504, g3505, g3508, g3506, g3507;
	wire g3511, g3512, g3509, g3510, g3513, g3514, g3516, g3517, g3518, g3521, g3519;
	wire g3520, g3522, g3523, g3524, g3525, g3527, g3528, g3529, g3532, g3530, g3531;
	wire g3535, g3536, g3533, g3534, g3537, g3538, g3540, g3541, g3542, g3545, g3543;
	wire g3544, g3546, g3547, g3548, g3549, g3551, g3552, g3553, g3556, g3554, g3555;
	wire g3559, g3557, g3558, g3560, g3561, g3563, g3564, g3565, g3568, g3566, g3567;
	wire g3571, g3572, g3569, g3570, g3573, g3574, g3576, g3577, g3578, g3581, g3579;
	wire g3580, g3584, g3585, g3582, g3583, g3586, g3587, g3589, g3590, g3591, g3594;
	wire g3592, g3593, g3597, g3598, g3595, g3596, g3599, g3600, g3602, g3603, g3604;
	wire g3607, g3605, g3606, g3610, g3611, g3608, g3609, g3612, g3613, g3615, g3616;
	wire g3617, g3620, g3618, g3619, g3623, g3624, g3621, g3622, g3625, g3626, g3628;
	wire g3629, g3630, g3633, g3631, g3632, g3636, g3634, g3635, g3637, g3639, g3640;
	wire g3641, g3644, g3642, g3643, g3647, g3645, g3646, g3648, g3649, g3651, g3652;
	wire g3653, g3656, g3654, g3655, g3659, g3660, g3657, g3658, g3661, g3662, g3664;
	wire g3665, g3666, g3669, g3667, g3668, g3672, g3673, g3670, g3671, g3674, g3675;
	wire g3677, g3678, g3679, g3682, g3680, g3681, g3687, g3685, g3683, g3684, g3686;
	wire g3688, g3689, g3690, g3693, g3691, g3692, g3696, g3697, g3694, g3695, g3698;
	wire g3699, g3700, g3701, g3702, g3703, g3706, g3704, g3705, g3709, g3707, g3708;
	wire g3710, g3711, g3713, g3714, g3715, g3718, g3716, g3717, g3721, g3722, g3719;
	wire g3720, g3723, g3724, g3726, g3727, g3728, g3731, g3729, g3730, g3734, g3735;
	wire g3732, g3733, g3736, g3737, g3739, g3740, g3741, g3744, g3742, g3743, g3747;
	wire g3748, g3745, g3746, g3749, g3750, g3752, g3753, g3754, g3757, g3755, g3756;
	wire g3760, g3761, g3758, g3759, g3762, g3763, g3765, g3766, g3767, g3770, g3768;
	wire g3769, g3773, g3774, g3771, g3772, g3775, g3776, g3778, g3779, g3780, g3783;
	wire g3781, g3782, g3786, g3784, g3785, g3787, g3789, g3790, g3791, g3794, g3792;
	wire g3793, g3797, g3798, g3795, g3796, g3799, g3800, g3802, g3803, g3804, g3807;
	wire g3805, g3806, g3810, g3811, g3808, g3809, g3812, g3813, g3815, g3816, g3814;
	wire g3817, g3820, g3818, g3819, g3821, g3822, g3824, g3825, g3826, g3829, g3827;
	wire g3828, g3832, g3833, g3830, g3831, g3834, g3835, g3837, g3838, g3839, g3842;
	wire g3840, g3841, g3845, g3846, g3843, g3844, g3847, g3848, g3850, g3851, g3852;
	wire g3855, g3853, g3854, g3858, g3856, g3857, g3859, g3861, g3862, g3863, g3866;
	wire g3864, g3865, g3869, g3867, g3868, g3870, g3872, g3873, g3874, g3877, g3875;
	wire g3876, g3880, g3878, g3879, g3881, g3883, g3884, g3885, g3888, g3886, g3887;
	wire g3891, g3889, g3890, g3892;


	reg g1, break_o, dmem_addr_ox0x, dmem_addr_ox1x, dmem_addr_ox2x, dmem_addr_ox3x, dmem_addr_ox4x, dmem_addr_ox5x, dmem_addr_ox6x;
	reg dmem_addr_ox7x, dmem_addr_ox8x, dmem_addr_ox9x, dmem_addr_ox10x, dmem_addr_ox11x, dmem_addr_ox12x, dmem_addr_ox13x, dmem_addr_ox14x, dmem_addr_ox15x;
	reg dmem_addr_ox16x, dmem_addr_ox17x, dmem_addr_ox18x, dmem_addr_ox19x, dmem_addr_ox20x, dmem_addr_ox21x, dmem_addr_ox22x, dmem_addr_ox23x, dmem_addr_ox24x;
	reg dmem_addr_ox25x, dmem_addr_ox26x, dmem_addr_ox27x, dmem_addr_ox28x, dmem_addr_ox29x, dmem_addr_ox30x, dmem_addr_ox31x, g35, g36;
	reg g37, g38, g39, g40, g41, g42, g43, g44, g45;
	reg g46, g47, g48, g49, g50, g51, g52, g53, g54;
	reg g55, g56, g57, g58, g59, g60, g61, g62, g63;
	reg g64, g65, g66, g67, g68, g69, dmem_sel_ox0x, dmem_sel_ox1x, dmem_sel_ox2x;
	reg dmem_sel_ox3x, g74, g75, g76, g77, g78, g79, g80, g81;
	reg g82, g83, g85, g86, g87, g88, g89, g90, g91;
	reg g92, g107, g108, g109, g110, g126, g128, g129, g141;
	reg g142, g143, g144, g145, g146, g147, g148, g150, g151;
	reg g152, g153, g155, g156, g157, g158, g160, g161, g162;
	reg g163, g165, g166, g168, g169, g170, g171, g173, g174;
	reg g175, g176, g178, g179, g180, g181, g183, g184, g185;
	reg g189, g190, g191, g192, g194, g195, g196, g197, g199;
	reg g200, g201, g202, g204, g205, g206, g207, g210, g211;
	reg g212, g213, g215, g216, g217, g218, g220, g221, g222;
	reg g223, g225, g226, g227, g232, g233, g234, g235, g237;
	reg g238, g239, g240, g242, g243, g244, g245, g247, g248;
	reg g249, g250, g253, g254, g255, g256, g258, g259, g260;
	reg g262, g263, g264, g265, g267, g268, g269, g270, g275;
	reg g276, g277, g278, g279, g281, g282, g283, g284, g286;
	reg g287, g288, g289, g291, g292, g293, g294, g297, g298;
	reg g299, g300, g302, g303, g304, g306, g307, g308, g309;
	reg g311, g312, g313, g314, g318, g319, g321, g322, g323;
	reg g324, g326, g327, g328, g329, g331, g332, g333, g334;
	reg g336, g337, g338, g339, g342, g343, g344, g345, g347;
	reg g348, g349, g351, g352, g353, g354, g356, g357, g358;
	reg g359, g364, g365, g366, g367, g368, g369, g371, g372;
	reg g373, g374, g376, g377, g378, g379, g381, g382, g383;
	reg g384, g387, g388, g389, g390, g392, g393, g394, g396;
	reg g397, g398, g399, g401, g402, g403, g404, g408, g410;
	reg g411, g412, g413, g415, g416, g417, g418, g420, g421;
	reg g422, g423, g425, g426, g427, g428, g431, g432, g433;
	reg g434, g436, g437, g438, g440, g441, g442, g443, g445;
	reg g446, g447, g448, g453, g454, g455, g456, g457, g459;
	reg g460, g461, g462, g464, g465, g466, g467, g469, g470;
	reg g471, g472, g475, g476, g477, g478, g480, g481, g482;
	reg g484, g485, g486, g487, g489, g490, g491, g492, g496;
	reg g498, g499, g500, g501, g503, g504, g505, g506, g508;
	reg g509, g510, g511, g513, g514, g515, g516, g519, g520;
	reg g521, g522, g524, g525, g526, g528, g529, g530, g531;
	reg g533, g534, g535, g536, g541, g543, g544, g545, g546;
	reg g548, g549, g550, g551, g553, g554, g555, g556, g558;
	reg g559, g560, g561, g564, g565, g566, g567, g569, g570;
	reg g571, g573, g574, g575, g576, g578, g579, g580, g581;
	reg g586, g587, g588, g589, g590, g591, g593, g594, g595;
	reg g596, g598, g599, g600, g601, g603, g604, g605, g606;
	reg g609, g610, g611, g612, g614, g615, g616, g618, g619;
	reg g620, g621, g623, g624, g625, g626, g630, g631, g632;
	reg g633, g634, g636, g637, g638, g639, g641, g642, g643;
	reg g644, g646, g647, g648, g649, g652, g653, g654, g655;
	reg g657, g658, g659, g661, g662, g663, g664, g666, g667;
	reg g668, g669, g677, g678, g682, g683, g684, g685, g687;
	reg g688, g689, g690, g692, g693, g694, g695, g697, g698;
	reg g699, g700, g703, g704, g705, g706, g708, g709, g710;
	reg g712, g713, g714, g715, g717, g718, g719, g720, g724;
	reg g726, g729, g730, g731, g732, g734, g735, g736, g737;
	reg g739, g740, g741, g742, g744, g745, g746, g747, g750;
	reg g751, g752, g753, g755, g756, g757, g759, g760, g761;
	reg g762, g764, g765, g766, g767, g771, g773, g776, g777;
	reg g778, g779, g781, g782, g783, g784, g786, g787, g788;
	reg g789, g791, g792, g793, g794, g797, g798, g799, g800;
	reg g802, g803, g804, g806, g807, g808, g809, g811, g812;
	reg g813, g814, g818, g820, g823, g824, g825, g826, g828;
	reg g829, g830, g831, g833, g834, g835, g836, g838, g839;
	reg g840, g841, g844, g845, g846, g847, g849, g850, g851;
	reg g853, g854, g855, g856, g858, g859, g860, g861, g865;
	reg g867, g870, g871, g872, g873, g875, g876, g877, g878;
	reg g880, g881, g882, g883, g885, g886, g887, g888, g891;
	reg g892, g893, g894, g896, g897, g898, g900, g901, g902;
	reg g903, g905, g906, g907, g908, g912, g918, g919, g920;
	reg g921, g923, g924, g925, g926, g928, g929, g930, g931;
	reg g933, g934, g935, g936, g939, g940, g941, g942, g944;
	reg g945, g946, g948, g949, g950, g951, g953, g954, g955;
	reg g956, g960, g963, g964, g965, g966, g968, g969, g970;
	reg g971, g973, g974, g975, g976, g978, g979, g980, g981;
	reg g984, g985, g986, g987, g989, g990, g991, g993, g994;
	reg g995, g996, g998, g999, g1000, g1001, g1005, g1008, g1009;
	reg g1010, g1011, g1013, g1014, g1015, g1016, g1018, g1019, g1020;
	reg g1021, g1023, g1024, g1025, g1026, g1029, g1030, g1031, g1032;
	reg g1034, g1035, g1036, g1038, g1039, g1040, g1041, g1043, g1044;
	reg g1045, g1046, g1050, g1053, g1054, g1055, g1056, g1058, g1059;
	reg g1060, g1061, g1063, g1064, g1065, g1066, g1068, g1069, g1070;
	reg g1071, g1074, g1075, g1076, g1077, g1079, g1080, g1081, g1083;
	reg g1084, g1085, g1086, g1088, g1089, g1090, g1091, g1095, g1098;
	reg g1099, g1100, g1101, g1103, g1104, g1105, g1106, g1108, g1109;
	reg g1110, g1111, g1113, g1114, g1115, g1116, g1119, g1120, g1121;
	reg g1122, g1124, g1125, g1126, g1128, g1129, g1130, g1131, g1133;
	reg g1134, g1135, g1136, g1140, g1143, g1144, g1145, g1146, g1148;
	reg g1149, g1150, g1151, g1153, g1154, g1155, g1156, g1158, g1159;
	reg g1160, g1161, g1164, g1165, g1166, g1167, g1169, g1170, g1171;
	reg g1173, g1174, g1175, g1176, g1178, g1179, g1180, g1181, g1185;
	reg g1188, g1189, g1190, g1191, g1193, g1194, g1195, g1196, g1198;
	reg g1199, g1200, g1201, g1203, g1204, g1205, g1206, g1209, g1210;
	reg g1211, g1212, g1214, g1215, g1216, g1218, g1219, g1220, g1221;
	reg g1223, g1224, g1225, g1226, g1230, g1233, g1234, g1235, g1236;
	reg g1238, g1239, g1240, g1241, g1243, g1244, g1245, g1246, g1248;
	reg g1249, g1250, g1251, g1254, g1255, g1256, g1257, g1259, g1260;
	reg g1261, g1263, g1264, g1265, g1266, g1268, g1269, g1270, g1271;
	reg g1275, g1278, g1279, g1280, g1281, g1283, g1284, g1285, g1286;
	reg g1288, g1289, g1290, g1291, g1293, g1294, g1295, g1296, g1299;
	reg g1300, g1301, g1302, g1304, g1305, g1306, g1308, g1309, g1310;
	reg g1311, g1313, g1314, g1315, g1316, g1320, g1323, g1324, g1325;
	reg g1326, g1328, g1329, g1330, g1331, g1333, g1334, g1335, g1336;
	reg g1338, g1339, g1340, g1341, g1344, g1345, g1346, g1347, g1349;
	reg g1350, g1351, g1353, g1354, g1355, g1356, g1358, g1359, g1360;
	reg g1361, g1365, g1368, g1369, g1370, g1371, g1373, g1374, g1375;
	reg g1376, g1378, g1379, g1380, g1381, g1383, g1384, g1385, g1386;
	reg g1389, g1390, g1391, g1392, g1394, g1395, g1396, g1398, g1399;
	reg g1400, g1401, g1403, g1404, g1405, g1406, g1410, g1413, g1414;
	reg g1415, g1416, g1418, g1419, g1420, g1421, g1423, g1424, g1425;
	reg g1426, g1428, g1429, g1430, g1431, g1434, g1435, g1436, g1437;
	reg g1439, g1440, g1441, g1443, g1444, g1445, g1446, g1448, g1449;
	reg g1450, g1451, g1455, g1458, g1459, g1460, g1461, g1463, g1464;
	reg g1465, g1466, g1468, g1469, g1470, g1471, g1473, g1474, g1475;
	reg g1476, g1479, g1480, g1481, g1482, g1484, g1485, g1486, g1488;
	reg g1489, g1490, g1491, g1493, g1494, g1495, g1496, g1500, g1502;
	reg g1503, g1504, g1505, g1507, g1508, g1509, g1510, g1512, g1513;
	reg g1514, g1515, g1517, g1518, g1519, g1520, g1523, g1524, g1525;
	reg g1526, g1528, g1529, g1530, g1532, g1533, g1534, g1535, g1537;
	reg g1538, g1539, g1540, g1544, g1547, g1548, g1549, g1550, g1551;
	reg g1553, g1554, g1555, g1556, g1558, g1559, g1560, g1561, g1563;
	reg g1564, g1565, g1566, g1569, g1570, g1571, g1572, g1574, g1575;
	reg g1576, g1578, g1579, g1580, g1581, g1583, g1584, g1585, g1586;
	reg g2019, g2023, g2026, g2035, g2038, g2055, g2060, g2066, g2070;
	reg g2071, g2073, g2074, g2076, g2077, g2079, g2080, g2081, g2083;
	reg g2084, g2085, g2086, g2088, g2089, g2090, g2091, g2093, g2094;
	reg g2095, g2096, g2098, g2099, g2100, g2101, g2104, g2105, g2106;
	reg g2108, g2109, g2110, g2111, g2113, g2114, g2115, g2116, g2118;
	reg g2119, g2120, g2121, g2124, g2125, g2128, g2129, g2134, g2135;
	reg g2136, g2137, g2138, g2231, g2258, g2284, g2289, g2306, g2312;
	reg g2333, g2340, g2357, g2365, g2383, g2391, g2413, g2418, g2432;
	reg g2439, g2457, g2476, g2482, g2499, g2507, g2523, g2529, g2544;
	reg g2551, g2566, g2570, g2587, g2590, g2605, g2608, g2622, g2625;
	reg g2639, g2642, g2657, g2660, g2677, g2680, g2696, g2699, g2712;
	reg g2715, g2731, g2734, g2748, g2751, g2767, g2771, g2791, g2794;
	reg g2808, g2811, g2824, g2827, g2831, g2914, g2969;

	always @ (posedge clk_i) begin g1 <= g124; end
	always @ (posedge clk_i) begin break_o <= g125; end
	always @ (posedge clk_i) begin dmem_addr_ox0x <= g3893; end
	always @ (posedge clk_i) begin dmem_addr_ox1x <= g3894; end
	always @ (posedge clk_i) begin dmem_addr_ox2x <= g3895; end
	always @ (posedge clk_i) begin dmem_addr_ox3x <= g3896; end
	always @ (posedge clk_i) begin dmem_addr_ox4x <= g3897; end
	always @ (posedge clk_i) begin dmem_addr_ox5x <= g3898; end
	always @ (posedge clk_i) begin dmem_addr_ox6x <= g3899; end
	always @ (posedge clk_i) begin dmem_addr_ox7x <= g3900; end
	always @ (posedge clk_i) begin dmem_addr_ox8x <= g3901; end
	always @ (posedge clk_i) begin dmem_addr_ox9x <= g3902; end
	always @ (posedge clk_i) begin dmem_addr_ox10x <= g3903; end
	always @ (posedge clk_i) begin dmem_addr_ox11x <= g3904; end
	always @ (posedge clk_i) begin dmem_addr_ox12x <= g3905; end
	always @ (posedge clk_i) begin dmem_addr_ox13x <= g3906; end
	always @ (posedge clk_i) begin dmem_addr_ox14x <= g3907; end
	always @ (posedge clk_i) begin dmem_addr_ox15x <= g3908; end
	always @ (posedge clk_i) begin dmem_addr_ox16x <= g3909; end
	always @ (posedge clk_i) begin dmem_addr_ox17x <= g3910; end
	always @ (posedge clk_i) begin dmem_addr_ox18x <= g3911; end
	always @ (posedge clk_i) begin dmem_addr_ox19x <= g3912; end
	always @ (posedge clk_i) begin dmem_addr_ox20x <= g3913; end
	always @ (posedge clk_i) begin dmem_addr_ox21x <= g3914; end
	always @ (posedge clk_i) begin dmem_addr_ox22x <= g3915; end
	always @ (posedge clk_i) begin dmem_addr_ox23x <= g3916; end
	always @ (posedge clk_i) begin dmem_addr_ox24x <= g3917; end
	always @ (posedge clk_i) begin dmem_addr_ox25x <= g3918; end
	always @ (posedge clk_i) begin dmem_addr_ox26x <= g3919; end
	always @ (posedge clk_i) begin dmem_addr_ox27x <= g3920; end
	always @ (posedge clk_i) begin dmem_addr_ox28x <= g3921; end
	always @ (posedge clk_i) begin dmem_addr_ox29x <= g3922; end
	always @ (posedge clk_i) begin dmem_addr_ox30x <= g3923; end
	always @ (posedge clk_i) begin dmem_addr_ox31x <= g3924; end
	always @ (posedge clk_i) begin g35 <= g3925; end
	always @ (posedge clk_i) begin g36 <= g3926; end
	always @ (posedge clk_i) begin g37 <= g3927; end
	always @ (posedge clk_i) begin g38 <= g3928; end
	always @ (posedge clk_i) begin g39 <= g3929; end
	always @ (posedge clk_i) begin g40 <= g3930; end
	always @ (posedge clk_i) begin g41 <= g3931; end
	always @ (posedge clk_i) begin g42 <= g3932; end
	always @ (posedge clk_i) begin g43 <= g3933; end
	always @ (posedge clk_i) begin g44 <= g3934; end
	always @ (posedge clk_i) begin g45 <= g3935; end
	always @ (posedge clk_i) begin g46 <= g3936; end
	always @ (posedge clk_i) begin g47 <= g3937; end
	always @ (posedge clk_i) begin g48 <= g3938; end
	always @ (posedge clk_i) begin g49 <= g3939; end
	always @ (posedge clk_i) begin g50 <= g3940; end
	always @ (posedge clk_i) begin g51 <= g3941; end
	always @ (posedge clk_i) begin g52 <= g3942; end
	always @ (posedge clk_i) begin g53 <= g3943; end
	always @ (posedge clk_i) begin g54 <= g3944; end
	always @ (posedge clk_i) begin g55 <= g3945; end
	always @ (posedge clk_i) begin g56 <= g3946; end
	always @ (posedge clk_i) begin g57 <= g3947; end
	always @ (posedge clk_i) begin g58 <= g3948; end
	always @ (posedge clk_i) begin g59 <= g3949; end
	always @ (posedge clk_i) begin g60 <= g3950; end
	always @ (posedge clk_i) begin g61 <= g3951; end
	always @ (posedge clk_i) begin g62 <= g3952; end
	always @ (posedge clk_i) begin g63 <= g3953; end
	always @ (posedge clk_i) begin g64 <= g3954; end
	always @ (posedge clk_i) begin g65 <= g3955; end
	always @ (posedge clk_i) begin g66 <= g3956; end
	always @ (posedge clk_i) begin g67 <= g3814; end
	always @ (posedge clk_i) begin g68 <= g2011; end
	always @ (posedge clk_i) begin g69 <= g2013; end
	always @ (posedge clk_i) begin dmem_sel_ox0x <= g3957; end
	always @ (posedge clk_i) begin dmem_sel_ox1x <= g3958; end
	always @ (posedge clk_i) begin dmem_sel_ox2x <= g3959; end
	always @ (posedge clk_i) begin dmem_sel_ox3x <= g3960; end
	always @ (posedge clk_i) begin g74 <= g138; end
	always @ (posedge clk_i) begin g75 <= g2021; end
	always @ (posedge clk_i) begin g76 <= g3961; end
	always @ (posedge clk_i) begin g77 <= g3962; end
	always @ (posedge clk_i) begin g78 <= g3963; end
	always @ (posedge clk_i) begin g79 <= g3964; end
	always @ (posedge clk_i) begin g80 <= g3965; end
	always @ (posedge clk_i) begin g81 <= g3966; end
	always @ (posedge clk_i) begin g82 <= g3967; end
	always @ (posedge clk_i) begin g83 <= g3968; end
	always @ (posedge clk_i) begin g85 <= g3969; end
	always @ (posedge clk_i) begin g86 <= g3970; end
	always @ (posedge clk_i) begin g87 <= g3971; end
	always @ (posedge clk_i) begin g88 <= g3972; end
	always @ (posedge clk_i) begin g89 <= g3973; end
	always @ (posedge clk_i) begin g90 <= g3974; end
	always @ (posedge clk_i) begin g91 <= g3975; end
	always @ (posedge clk_i) begin g92 <= g3976; end
	always @ (posedge clk_i) begin g107 <= g3977; end
	always @ (posedge clk_i) begin g108 <= g3978; end
	always @ (posedge clk_i) begin g109 <= g3979; end
	always @ (posedge clk_i) begin g110 <= g3980; end
	always @ (posedge clk_i) begin g126 <= g2064; end
	always @ (posedge clk_i) begin g128 <= vcc; end
	always @ (posedge clk_i) begin g129 <= g2065; end
	always @ (posedge clk_i) begin g141 <= g3981; end
	always @ (posedge clk_i) begin g142 <= g3982; end
	always @ (posedge clk_i) begin g143 <= g3983; end
	always @ (posedge clk_i) begin g144 <= g3984; end
	always @ (posedge clk_i) begin g145 <= g3985; end
	always @ (posedge clk_i) begin g146 <= g3986; end
	always @ (posedge clk_i) begin g147 <= g3987; end
	always @ (posedge clk_i) begin g148 <= g3988; end
	always @ (posedge clk_i) begin g150 <= g3989; end
	always @ (posedge clk_i) begin g151 <= g3990; end
	always @ (posedge clk_i) begin g152 <= g3991; end
	always @ (posedge clk_i) begin g153 <= g3992; end
	always @ (posedge clk_i) begin g155 <= g3993; end
	always @ (posedge clk_i) begin g156 <= g3994; end
	always @ (posedge clk_i) begin g157 <= g3995; end
	always @ (posedge clk_i) begin g158 <= g3996; end
	always @ (posedge clk_i) begin g160 <= g3997; end
	always @ (posedge clk_i) begin g161 <= g3998; end
	always @ (posedge clk_i) begin g162 <= g3999; end
	always @ (posedge clk_i) begin g163 <= g4000; end
	always @ (posedge clk_i) begin g165 <= g4001; end
	always @ (posedge clk_i) begin g166 <= g4002; end
	always @ (posedge clk_i) begin g168 <= g4003; end
	always @ (posedge clk_i) begin g169 <= g4004; end
	always @ (posedge clk_i) begin g170 <= g4005; end
	always @ (posedge clk_i) begin g171 <= g4006; end
	always @ (posedge clk_i) begin g173 <= g4007; end
	always @ (posedge clk_i) begin g174 <= g4008; end
	always @ (posedge clk_i) begin g175 <= g4009; end
	always @ (posedge clk_i) begin g176 <= g4010; end
	always @ (posedge clk_i) begin g178 <= g4011; end
	always @ (posedge clk_i) begin g179 <= g4012; end
	always @ (posedge clk_i) begin g180 <= g4013; end
	always @ (posedge clk_i) begin g181 <= g4014; end
	always @ (posedge clk_i) begin g183 <= g4015; end
	always @ (posedge clk_i) begin g184 <= g4016; end
	always @ (posedge clk_i) begin g185 <= g4017; end
	always @ (posedge clk_i) begin g189 <= g4018; end
	always @ (posedge clk_i) begin g190 <= g4019; end
	always @ (posedge clk_i) begin g191 <= g4020; end
	always @ (posedge clk_i) begin g192 <= g4021; end
	always @ (posedge clk_i) begin g194 <= g4022; end
	always @ (posedge clk_i) begin g195 <= g4023; end
	always @ (posedge clk_i) begin g196 <= g4024; end
	always @ (posedge clk_i) begin g197 <= g4025; end
	always @ (posedge clk_i) begin g199 <= g4026; end
	always @ (posedge clk_i) begin g200 <= g4027; end
	always @ (posedge clk_i) begin g201 <= g4028; end
	always @ (posedge clk_i) begin g202 <= g4029; end
	always @ (posedge clk_i) begin g204 <= g4030; end
	always @ (posedge clk_i) begin g205 <= g4031; end
	always @ (posedge clk_i) begin g206 <= g4032; end
	always @ (posedge clk_i) begin g207 <= g4033; end
	always @ (posedge clk_i) begin g210 <= g4034; end
	always @ (posedge clk_i) begin g211 <= g4035; end
	always @ (posedge clk_i) begin g212 <= g4036; end
	always @ (posedge clk_i) begin g213 <= g4037; end
	always @ (posedge clk_i) begin g215 <= g4038; end
	always @ (posedge clk_i) begin g216 <= g4039; end
	always @ (posedge clk_i) begin g217 <= g4040; end
	always @ (posedge clk_i) begin g218 <= g4041; end
	always @ (posedge clk_i) begin g220 <= g4042; end
	always @ (posedge clk_i) begin g221 <= g4043; end
	always @ (posedge clk_i) begin g222 <= g4044; end
	always @ (posedge clk_i) begin g223 <= g4045; end
	always @ (posedge clk_i) begin g225 <= g4046; end
	always @ (posedge clk_i) begin g226 <= g4047; end
	always @ (posedge clk_i) begin g227 <= g4048; end
	always @ (posedge clk_i) begin g232 <= g4049; end
	always @ (posedge clk_i) begin g233 <= g4050; end
	always @ (posedge clk_i) begin g234 <= g4051; end
	always @ (posedge clk_i) begin g235 <= g4052; end
	always @ (posedge clk_i) begin g237 <= g4053; end
	always @ (posedge clk_i) begin g238 <= g4054; end
	always @ (posedge clk_i) begin g239 <= g4055; end
	always @ (posedge clk_i) begin g240 <= g4056; end
	always @ (posedge clk_i) begin g242 <= g4057; end
	always @ (posedge clk_i) begin g243 <= g4058; end
	always @ (posedge clk_i) begin g244 <= g4059; end
	always @ (posedge clk_i) begin g245 <= g4060; end
	always @ (posedge clk_i) begin g247 <= g4061; end
	always @ (posedge clk_i) begin g248 <= g4062; end
	always @ (posedge clk_i) begin g249 <= g4063; end
	always @ (posedge clk_i) begin g250 <= g4064; end
	always @ (posedge clk_i) begin g253 <= g4065; end
	always @ (posedge clk_i) begin g254 <= g4066; end
	always @ (posedge clk_i) begin g255 <= g4067; end
	always @ (posedge clk_i) begin g256 <= g4068; end
	always @ (posedge clk_i) begin g258 <= g4069; end
	always @ (posedge clk_i) begin g259 <= g4070; end
	always @ (posedge clk_i) begin g260 <= g4071; end
	always @ (posedge clk_i) begin g262 <= g4072; end
	always @ (posedge clk_i) begin g263 <= g4073; end
	always @ (posedge clk_i) begin g264 <= g4074; end
	always @ (posedge clk_i) begin g265 <= g4075; end
	always @ (posedge clk_i) begin g267 <= g4076; end
	always @ (posedge clk_i) begin g268 <= g4077; end
	always @ (posedge clk_i) begin g269 <= g4078; end
	always @ (posedge clk_i) begin g270 <= g4079; end
	always @ (posedge clk_i) begin g275 <= g4080; end
	always @ (posedge clk_i) begin g276 <= g4081; end
	always @ (posedge clk_i) begin g277 <= g4082; end
	always @ (posedge clk_i) begin g278 <= g4083; end
	always @ (posedge clk_i) begin g279 <= g4084; end
	always @ (posedge clk_i) begin g281 <= g4085; end
	always @ (posedge clk_i) begin g282 <= g4086; end
	always @ (posedge clk_i) begin g283 <= g4087; end
	always @ (posedge clk_i) begin g284 <= g4088; end
	always @ (posedge clk_i) begin g286 <= g4089; end
	always @ (posedge clk_i) begin g287 <= g4090; end
	always @ (posedge clk_i) begin g288 <= g4091; end
	always @ (posedge clk_i) begin g289 <= g4092; end
	always @ (posedge clk_i) begin g291 <= g4093; end
	always @ (posedge clk_i) begin g292 <= g4094; end
	always @ (posedge clk_i) begin g293 <= g4095; end
	always @ (posedge clk_i) begin g294 <= g4096; end
	always @ (posedge clk_i) begin g297 <= g4097; end
	always @ (posedge clk_i) begin g298 <= g4098; end
	always @ (posedge clk_i) begin g299 <= g4099; end
	always @ (posedge clk_i) begin g300 <= g4100; end
	always @ (posedge clk_i) begin g302 <= g4101; end
	always @ (posedge clk_i) begin g303 <= g4102; end
	always @ (posedge clk_i) begin g304 <= g4103; end
	always @ (posedge clk_i) begin g306 <= g4104; end
	always @ (posedge clk_i) begin g307 <= g4105; end
	always @ (posedge clk_i) begin g308 <= g4106; end
	always @ (posedge clk_i) begin g309 <= g4107; end
	always @ (posedge clk_i) begin g311 <= g4108; end
	always @ (posedge clk_i) begin g312 <= g4109; end
	always @ (posedge clk_i) begin g313 <= g4110; end
	always @ (posedge clk_i) begin g314 <= g4111; end
	always @ (posedge clk_i) begin g318 <= g4112; end
	always @ (posedge clk_i) begin g319 <= g4113; end
	always @ (posedge clk_i) begin g321 <= g4114; end
	always @ (posedge clk_i) begin g322 <= g4115; end
	always @ (posedge clk_i) begin g323 <= g4116; end
	always @ (posedge clk_i) begin g324 <= g4117; end
	always @ (posedge clk_i) begin g326 <= g4118; end
	always @ (posedge clk_i) begin g327 <= g4119; end
	always @ (posedge clk_i) begin g328 <= g4120; end
	always @ (posedge clk_i) begin g329 <= g4121; end
	always @ (posedge clk_i) begin g331 <= g4122; end
	always @ (posedge clk_i) begin g332 <= g4123; end
	always @ (posedge clk_i) begin g333 <= g4124; end
	always @ (posedge clk_i) begin g334 <= g4125; end
	always @ (posedge clk_i) begin g336 <= g4126; end
	always @ (posedge clk_i) begin g337 <= g4127; end
	always @ (posedge clk_i) begin g338 <= g4128; end
	always @ (posedge clk_i) begin g339 <= g4129; end
	always @ (posedge clk_i) begin g342 <= g4130; end
	always @ (posedge clk_i) begin g343 <= g4131; end
	always @ (posedge clk_i) begin g344 <= g4132; end
	always @ (posedge clk_i) begin g345 <= g4133; end
	always @ (posedge clk_i) begin g347 <= g4134; end
	always @ (posedge clk_i) begin g348 <= g4135; end
	always @ (posedge clk_i) begin g349 <= g4136; end
	always @ (posedge clk_i) begin g351 <= g4137; end
	always @ (posedge clk_i) begin g352 <= g4138; end
	always @ (posedge clk_i) begin g353 <= g4139; end
	always @ (posedge clk_i) begin g354 <= g4140; end
	always @ (posedge clk_i) begin g356 <= g4141; end
	always @ (posedge clk_i) begin g357 <= g4142; end
	always @ (posedge clk_i) begin g358 <= g4143; end
	always @ (posedge clk_i) begin g359 <= g4144; end
	always @ (posedge clk_i) begin g364 <= g4145; end
	always @ (posedge clk_i) begin g365 <= g4146; end
	always @ (posedge clk_i) begin g366 <= g4147; end
	always @ (posedge clk_i) begin g367 <= g4148; end
	always @ (posedge clk_i) begin g368 <= g4149; end
	always @ (posedge clk_i) begin g369 <= g4150; end
	always @ (posedge clk_i) begin g371 <= g4151; end
	always @ (posedge clk_i) begin g372 <= g4152; end
	always @ (posedge clk_i) begin g373 <= g4153; end
	always @ (posedge clk_i) begin g374 <= g4154; end
	always @ (posedge clk_i) begin g376 <= g4155; end
	always @ (posedge clk_i) begin g377 <= g4156; end
	always @ (posedge clk_i) begin g378 <= g4157; end
	always @ (posedge clk_i) begin g379 <= g4158; end
	always @ (posedge clk_i) begin g381 <= g4159; end
	always @ (posedge clk_i) begin g382 <= g4160; end
	always @ (posedge clk_i) begin g383 <= g4161; end
	always @ (posedge clk_i) begin g384 <= g4162; end
	always @ (posedge clk_i) begin g387 <= g4163; end
	always @ (posedge clk_i) begin g388 <= g4164; end
	always @ (posedge clk_i) begin g389 <= g4165; end
	always @ (posedge clk_i) begin g390 <= g4166; end
	always @ (posedge clk_i) begin g392 <= g4167; end
	always @ (posedge clk_i) begin g393 <= g4168; end
	always @ (posedge clk_i) begin g394 <= g4169; end
	always @ (posedge clk_i) begin g396 <= g4170; end
	always @ (posedge clk_i) begin g397 <= g4171; end
	always @ (posedge clk_i) begin g398 <= g4172; end
	always @ (posedge clk_i) begin g399 <= g4173; end
	always @ (posedge clk_i) begin g401 <= g4174; end
	always @ (posedge clk_i) begin g402 <= g4175; end
	always @ (posedge clk_i) begin g403 <= g4176; end
	always @ (posedge clk_i) begin g404 <= g4177; end
	always @ (posedge clk_i) begin g408 <= g4178; end
	always @ (posedge clk_i) begin g410 <= g4179; end
	always @ (posedge clk_i) begin g411 <= g4180; end
	always @ (posedge clk_i) begin g412 <= g4181; end
	always @ (posedge clk_i) begin g413 <= g4182; end
	always @ (posedge clk_i) begin g415 <= g4183; end
	always @ (posedge clk_i) begin g416 <= g4184; end
	always @ (posedge clk_i) begin g417 <= g4185; end
	always @ (posedge clk_i) begin g418 <= g4186; end
	always @ (posedge clk_i) begin g420 <= g4187; end
	always @ (posedge clk_i) begin g421 <= g4188; end
	always @ (posedge clk_i) begin g422 <= g4189; end
	always @ (posedge clk_i) begin g423 <= g4190; end
	always @ (posedge clk_i) begin g425 <= g4191; end
	always @ (posedge clk_i) begin g426 <= g4192; end
	always @ (posedge clk_i) begin g427 <= g4193; end
	always @ (posedge clk_i) begin g428 <= g4194; end
	always @ (posedge clk_i) begin g431 <= g4195; end
	always @ (posedge clk_i) begin g432 <= g4196; end
	always @ (posedge clk_i) begin g433 <= g4197; end
	always @ (posedge clk_i) begin g434 <= g4198; end
	always @ (posedge clk_i) begin g436 <= g4199; end
	always @ (posedge clk_i) begin g437 <= g4200; end
	always @ (posedge clk_i) begin g438 <= g4201; end
	always @ (posedge clk_i) begin g440 <= g4202; end
	always @ (posedge clk_i) begin g441 <= g4203; end
	always @ (posedge clk_i) begin g442 <= g4204; end
	always @ (posedge clk_i) begin g443 <= g4205; end
	always @ (posedge clk_i) begin g445 <= g4206; end
	always @ (posedge clk_i) begin g446 <= g4207; end
	always @ (posedge clk_i) begin g447 <= g4208; end
	always @ (posedge clk_i) begin g448 <= g4209; end
	always @ (posedge clk_i) begin g453 <= g4210; end
	always @ (posedge clk_i) begin g454 <= g4211; end
	always @ (posedge clk_i) begin g455 <= g4212; end
	always @ (posedge clk_i) begin g456 <= g4213; end
	always @ (posedge clk_i) begin g457 <= g4214; end
	always @ (posedge clk_i) begin g459 <= g4215; end
	always @ (posedge clk_i) begin g460 <= g4216; end
	always @ (posedge clk_i) begin g461 <= g4217; end
	always @ (posedge clk_i) begin g462 <= g4218; end
	always @ (posedge clk_i) begin g464 <= g4219; end
	always @ (posedge clk_i) begin g465 <= g4220; end
	always @ (posedge clk_i) begin g466 <= g4221; end
	always @ (posedge clk_i) begin g467 <= g4222; end
	always @ (posedge clk_i) begin g469 <= g4223; end
	always @ (posedge clk_i) begin g470 <= g4224; end
	always @ (posedge clk_i) begin g471 <= g4225; end
	always @ (posedge clk_i) begin g472 <= g4226; end
	always @ (posedge clk_i) begin g475 <= g4227; end
	always @ (posedge clk_i) begin g476 <= g4228; end
	always @ (posedge clk_i) begin g477 <= g4229; end
	always @ (posedge clk_i) begin g478 <= g4230; end
	always @ (posedge clk_i) begin g480 <= g4231; end
	always @ (posedge clk_i) begin g481 <= g4232; end
	always @ (posedge clk_i) begin g482 <= g4233; end
	always @ (posedge clk_i) begin g484 <= g4234; end
	always @ (posedge clk_i) begin g485 <= g4235; end
	always @ (posedge clk_i) begin g486 <= g4236; end
	always @ (posedge clk_i) begin g487 <= g4237; end
	always @ (posedge clk_i) begin g489 <= g4238; end
	always @ (posedge clk_i) begin g490 <= g4239; end
	always @ (posedge clk_i) begin g491 <= g4240; end
	always @ (posedge clk_i) begin g492 <= g4241; end
	always @ (posedge clk_i) begin g496 <= g4243; end
	always @ (posedge clk_i) begin g498 <= g4244; end
	always @ (posedge clk_i) begin g499 <= g4245; end
	always @ (posedge clk_i) begin g500 <= g4246; end
	always @ (posedge clk_i) begin g501 <= g4247; end
	always @ (posedge clk_i) begin g503 <= g4248; end
	always @ (posedge clk_i) begin g504 <= g4249; end
	always @ (posedge clk_i) begin g505 <= g4250; end
	always @ (posedge clk_i) begin g506 <= g4251; end
	always @ (posedge clk_i) begin g508 <= g4252; end
	always @ (posedge clk_i) begin g509 <= g4253; end
	always @ (posedge clk_i) begin g510 <= g4254; end
	always @ (posedge clk_i) begin g511 <= g4255; end
	always @ (posedge clk_i) begin g513 <= g4256; end
	always @ (posedge clk_i) begin g514 <= g4257; end
	always @ (posedge clk_i) begin g515 <= g4258; end
	always @ (posedge clk_i) begin g516 <= g4259; end
	always @ (posedge clk_i) begin g519 <= g4260; end
	always @ (posedge clk_i) begin g520 <= g4261; end
	always @ (posedge clk_i) begin g521 <= g4262; end
	always @ (posedge clk_i) begin g522 <= g4263; end
	always @ (posedge clk_i) begin g524 <= g4264; end
	always @ (posedge clk_i) begin g525 <= g4265; end
	always @ (posedge clk_i) begin g526 <= g4266; end
	always @ (posedge clk_i) begin g528 <= g4267; end
	always @ (posedge clk_i) begin g529 <= g4268; end
	always @ (posedge clk_i) begin g530 <= g4269; end
	always @ (posedge clk_i) begin g531 <= g4270; end
	always @ (posedge clk_i) begin g533 <= g4271; end
	always @ (posedge clk_i) begin g534 <= g4272; end
	always @ (posedge clk_i) begin g535 <= g4273; end
	always @ (posedge clk_i) begin g536 <= g4274; end
	always @ (posedge clk_i) begin g541 <= g4275; end
	always @ (posedge clk_i) begin g543 <= g4276; end
	always @ (posedge clk_i) begin g544 <= g4277; end
	always @ (posedge clk_i) begin g545 <= g4278; end
	always @ (posedge clk_i) begin g546 <= g4279; end
	always @ (posedge clk_i) begin g548 <= g4280; end
	always @ (posedge clk_i) begin g549 <= g4281; end
	always @ (posedge clk_i) begin g550 <= g4282; end
	always @ (posedge clk_i) begin g551 <= g4283; end
	always @ (posedge clk_i) begin g553 <= g4284; end
	always @ (posedge clk_i) begin g554 <= g4285; end
	always @ (posedge clk_i) begin g555 <= g4286; end
	always @ (posedge clk_i) begin g556 <= g4287; end
	always @ (posedge clk_i) begin g558 <= g4288; end
	always @ (posedge clk_i) begin g559 <= g4289; end
	always @ (posedge clk_i) begin g560 <= g4290; end
	always @ (posedge clk_i) begin g561 <= g4291; end
	always @ (posedge clk_i) begin g564 <= g4292; end
	always @ (posedge clk_i) begin g565 <= g4293; end
	always @ (posedge clk_i) begin g566 <= g4294; end
	always @ (posedge clk_i) begin g567 <= g4295; end
	always @ (posedge clk_i) begin g569 <= g4296; end
	always @ (posedge clk_i) begin g570 <= g4297; end
	always @ (posedge clk_i) begin g571 <= g4298; end
	always @ (posedge clk_i) begin g573 <= g4299; end
	always @ (posedge clk_i) begin g574 <= g4300; end
	always @ (posedge clk_i) begin g575 <= g4301; end
	always @ (posedge clk_i) begin g576 <= g4302; end
	always @ (posedge clk_i) begin g578 <= g4303; end
	always @ (posedge clk_i) begin g579 <= g4304; end
	always @ (posedge clk_i) begin g580 <= g4305; end
	always @ (posedge clk_i) begin g581 <= g4306; end
	always @ (posedge clk_i) begin g586 <= g4307; end
	always @ (posedge clk_i) begin g587 <= g4308; end
	always @ (posedge clk_i) begin g588 <= g4309; end
	always @ (posedge clk_i) begin g589 <= g4310; end
	always @ (posedge clk_i) begin g590 <= g4311; end
	always @ (posedge clk_i) begin g591 <= g4312; end
	always @ (posedge clk_i) begin g593 <= g4313; end
	always @ (posedge clk_i) begin g594 <= g4314; end
	always @ (posedge clk_i) begin g595 <= g4315; end
	always @ (posedge clk_i) begin g596 <= g4316; end
	always @ (posedge clk_i) begin g598 <= g4317; end
	always @ (posedge clk_i) begin g599 <= g4318; end
	always @ (posedge clk_i) begin g600 <= g4319; end
	always @ (posedge clk_i) begin g601 <= g4320; end
	always @ (posedge clk_i) begin g603 <= g4321; end
	always @ (posedge clk_i) begin g604 <= g4322; end
	always @ (posedge clk_i) begin g605 <= g4323; end
	always @ (posedge clk_i) begin g606 <= g4324; end
	always @ (posedge clk_i) begin g609 <= g4325; end
	always @ (posedge clk_i) begin g610 <= g4326; end
	always @ (posedge clk_i) begin g611 <= g4327; end
	always @ (posedge clk_i) begin g612 <= g4328; end
	always @ (posedge clk_i) begin g614 <= g4329; end
	always @ (posedge clk_i) begin g615 <= g4330; end
	always @ (posedge clk_i) begin g616 <= g4331; end
	always @ (posedge clk_i) begin g618 <= g4332; end
	always @ (posedge clk_i) begin g619 <= g4333; end
	always @ (posedge clk_i) begin g620 <= g4334; end
	always @ (posedge clk_i) begin g621 <= g4335; end
	always @ (posedge clk_i) begin g623 <= g4336; end
	always @ (posedge clk_i) begin g624 <= g4337; end
	always @ (posedge clk_i) begin g625 <= g4338; end
	always @ (posedge clk_i) begin g626 <= g4339; end
	always @ (posedge clk_i) begin g630 <= g4340; end
	always @ (posedge clk_i) begin g631 <= g4341; end
	always @ (posedge clk_i) begin g632 <= g4342; end
	always @ (posedge clk_i) begin g633 <= g4343; end
	always @ (posedge clk_i) begin g634 <= g4344; end
	always @ (posedge clk_i) begin g636 <= g4345; end
	always @ (posedge clk_i) begin g637 <= g4346; end
	always @ (posedge clk_i) begin g638 <= g4347; end
	always @ (posedge clk_i) begin g639 <= g4348; end
	always @ (posedge clk_i) begin g641 <= g4349; end
	always @ (posedge clk_i) begin g642 <= g4350; end
	always @ (posedge clk_i) begin g643 <= g4351; end
	always @ (posedge clk_i) begin g644 <= g4352; end
	always @ (posedge clk_i) begin g646 <= g4353; end
	always @ (posedge clk_i) begin g647 <= g4354; end
	always @ (posedge clk_i) begin g648 <= g4355; end
	always @ (posedge clk_i) begin g649 <= g4356; end
	always @ (posedge clk_i) begin g652 <= g4357; end
	always @ (posedge clk_i) begin g653 <= g4358; end
	always @ (posedge clk_i) begin g654 <= g4359; end
	always @ (posedge clk_i) begin g655 <= g4360; end
	always @ (posedge clk_i) begin g657 <= g4361; end
	always @ (posedge clk_i) begin g658 <= g4362; end
	always @ (posedge clk_i) begin g659 <= g4363; end
	always @ (posedge clk_i) begin g661 <= g4364; end
	always @ (posedge clk_i) begin g662 <= g4365; end
	always @ (posedge clk_i) begin g663 <= g4366; end
	always @ (posedge clk_i) begin g664 <= g4367; end
	always @ (posedge clk_i) begin g666 <= g4368; end
	always @ (posedge clk_i) begin g667 <= g4369; end
	always @ (posedge clk_i) begin g668 <= g4370; end
	always @ (posedge clk_i) begin g669 <= g4371; end
	always @ (posedge clk_i) begin g677 <= g4372; end
	always @ (posedge clk_i) begin g678 <= g4373; end
	always @ (posedge clk_i) begin g682 <= g4374; end
	always @ (posedge clk_i) begin g683 <= g4375; end
	always @ (posedge clk_i) begin g684 <= g4376; end
	always @ (posedge clk_i) begin g685 <= g4377; end
	always @ (posedge clk_i) begin g687 <= g4378; end
	always @ (posedge clk_i) begin g688 <= g4379; end
	always @ (posedge clk_i) begin g689 <= g4380; end
	always @ (posedge clk_i) begin g690 <= g4381; end
	always @ (posedge clk_i) begin g692 <= g4382; end
	always @ (posedge clk_i) begin g693 <= g4383; end
	always @ (posedge clk_i) begin g694 <= g4384; end
	always @ (posedge clk_i) begin g695 <= g4385; end
	always @ (posedge clk_i) begin g697 <= g4386; end
	always @ (posedge clk_i) begin g698 <= g4387; end
	always @ (posedge clk_i) begin g699 <= g4388; end
	always @ (posedge clk_i) begin g700 <= g4389; end
	always @ (posedge clk_i) begin g703 <= g4390; end
	always @ (posedge clk_i) begin g704 <= g4391; end
	always @ (posedge clk_i) begin g705 <= g4392; end
	always @ (posedge clk_i) begin g706 <= g4393; end
	always @ (posedge clk_i) begin g708 <= g4394; end
	always @ (posedge clk_i) begin g709 <= g4395; end
	always @ (posedge clk_i) begin g710 <= g4396; end
	always @ (posedge clk_i) begin g712 <= g4397; end
	always @ (posedge clk_i) begin g713 <= g4398; end
	always @ (posedge clk_i) begin g714 <= g4399; end
	always @ (posedge clk_i) begin g715 <= g4400; end
	always @ (posedge clk_i) begin g717 <= g4401; end
	always @ (posedge clk_i) begin g718 <= g4402; end
	always @ (posedge clk_i) begin g719 <= g4403; end
	always @ (posedge clk_i) begin g720 <= g4404; end
	always @ (posedge clk_i) begin g724 <= g4405; end
	always @ (posedge clk_i) begin g726 <= g4406; end
	always @ (posedge clk_i) begin g729 <= g4407; end
	always @ (posedge clk_i) begin g730 <= g4408; end
	always @ (posedge clk_i) begin g731 <= g4409; end
	always @ (posedge clk_i) begin g732 <= g4410; end
	always @ (posedge clk_i) begin g734 <= g4411; end
	always @ (posedge clk_i) begin g735 <= g4412; end
	always @ (posedge clk_i) begin g736 <= g4413; end
	always @ (posedge clk_i) begin g737 <= g4414; end
	always @ (posedge clk_i) begin g739 <= g4415; end
	always @ (posedge clk_i) begin g740 <= g4416; end
	always @ (posedge clk_i) begin g741 <= g4417; end
	always @ (posedge clk_i) begin g742 <= g4418; end
	always @ (posedge clk_i) begin g744 <= g4419; end
	always @ (posedge clk_i) begin g745 <= g4420; end
	always @ (posedge clk_i) begin g746 <= g4421; end
	always @ (posedge clk_i) begin g747 <= g4422; end
	always @ (posedge clk_i) begin g750 <= g4423; end
	always @ (posedge clk_i) begin g751 <= g4424; end
	always @ (posedge clk_i) begin g752 <= g4425; end
	always @ (posedge clk_i) begin g753 <= g4426; end
	always @ (posedge clk_i) begin g755 <= g4427; end
	always @ (posedge clk_i) begin g756 <= g4428; end
	always @ (posedge clk_i) begin g757 <= g4429; end
	always @ (posedge clk_i) begin g759 <= g4430; end
	always @ (posedge clk_i) begin g760 <= g4431; end
	always @ (posedge clk_i) begin g761 <= g4432; end
	always @ (posedge clk_i) begin g762 <= g4433; end
	always @ (posedge clk_i) begin g764 <= g4434; end
	always @ (posedge clk_i) begin g765 <= g4435; end
	always @ (posedge clk_i) begin g766 <= g4436; end
	always @ (posedge clk_i) begin g767 <= g4437; end
	always @ (posedge clk_i) begin g771 <= g4438; end
	always @ (posedge clk_i) begin g773 <= g4439; end
	always @ (posedge clk_i) begin g776 <= g4440; end
	always @ (posedge clk_i) begin g777 <= g4441; end
	always @ (posedge clk_i) begin g778 <= g4442; end
	always @ (posedge clk_i) begin g779 <= g4443; end
	always @ (posedge clk_i) begin g781 <= g4444; end
	always @ (posedge clk_i) begin g782 <= g4445; end
	always @ (posedge clk_i) begin g783 <= g4446; end
	always @ (posedge clk_i) begin g784 <= g4447; end
	always @ (posedge clk_i) begin g786 <= g4448; end
	always @ (posedge clk_i) begin g787 <= g4449; end
	always @ (posedge clk_i) begin g788 <= g4450; end
	always @ (posedge clk_i) begin g789 <= g4451; end
	always @ (posedge clk_i) begin g791 <= g4452; end
	always @ (posedge clk_i) begin g792 <= g4453; end
	always @ (posedge clk_i) begin g793 <= g4454; end
	always @ (posedge clk_i) begin g794 <= g4455; end
	always @ (posedge clk_i) begin g797 <= g4456; end
	always @ (posedge clk_i) begin g798 <= g4457; end
	always @ (posedge clk_i) begin g799 <= g4458; end
	always @ (posedge clk_i) begin g800 <= g4459; end
	always @ (posedge clk_i) begin g802 <= g4460; end
	always @ (posedge clk_i) begin g803 <= g4461; end
	always @ (posedge clk_i) begin g804 <= g4462; end
	always @ (posedge clk_i) begin g806 <= g4463; end
	always @ (posedge clk_i) begin g807 <= g4464; end
	always @ (posedge clk_i) begin g808 <= g4465; end
	always @ (posedge clk_i) begin g809 <= g4466; end
	always @ (posedge clk_i) begin g811 <= g4467; end
	always @ (posedge clk_i) begin g812 <= g4468; end
	always @ (posedge clk_i) begin g813 <= g4469; end
	always @ (posedge clk_i) begin g814 <= g4470; end
	always @ (posedge clk_i) begin g818 <= g4471; end
	always @ (posedge clk_i) begin g820 <= g4472; end
	always @ (posedge clk_i) begin g823 <= g4473; end
	always @ (posedge clk_i) begin g824 <= g4474; end
	always @ (posedge clk_i) begin g825 <= g4475; end
	always @ (posedge clk_i) begin g826 <= g4476; end
	always @ (posedge clk_i) begin g828 <= g4477; end
	always @ (posedge clk_i) begin g829 <= g4478; end
	always @ (posedge clk_i) begin g830 <= g4479; end
	always @ (posedge clk_i) begin g831 <= g4480; end
	always @ (posedge clk_i) begin g833 <= g4481; end
	always @ (posedge clk_i) begin g834 <= g4482; end
	always @ (posedge clk_i) begin g835 <= g4483; end
	always @ (posedge clk_i) begin g836 <= g4484; end
	always @ (posedge clk_i) begin g838 <= g4485; end
	always @ (posedge clk_i) begin g839 <= g4486; end
	always @ (posedge clk_i) begin g840 <= g4487; end
	always @ (posedge clk_i) begin g841 <= g4488; end
	always @ (posedge clk_i) begin g844 <= g4489; end
	always @ (posedge clk_i) begin g845 <= g4490; end
	always @ (posedge clk_i) begin g846 <= g4491; end
	always @ (posedge clk_i) begin g847 <= g4492; end
	always @ (posedge clk_i) begin g849 <= g4493; end
	always @ (posedge clk_i) begin g850 <= g4494; end
	always @ (posedge clk_i) begin g851 <= g4495; end
	always @ (posedge clk_i) begin g853 <= g4496; end
	always @ (posedge clk_i) begin g854 <= g4497; end
	always @ (posedge clk_i) begin g855 <= g4498; end
	always @ (posedge clk_i) begin g856 <= g4499; end
	always @ (posedge clk_i) begin g858 <= g4500; end
	always @ (posedge clk_i) begin g859 <= g4501; end
	always @ (posedge clk_i) begin g860 <= g4502; end
	always @ (posedge clk_i) begin g861 <= g4503; end
	always @ (posedge clk_i) begin g865 <= g4504; end
	always @ (posedge clk_i) begin g867 <= g4505; end
	always @ (posedge clk_i) begin g870 <= g4506; end
	always @ (posedge clk_i) begin g871 <= g4507; end
	always @ (posedge clk_i) begin g872 <= g4508; end
	always @ (posedge clk_i) begin g873 <= g4509; end
	always @ (posedge clk_i) begin g875 <= g4510; end
	always @ (posedge clk_i) begin g876 <= g4511; end
	always @ (posedge clk_i) begin g877 <= g4512; end
	always @ (posedge clk_i) begin g878 <= g4513; end
	always @ (posedge clk_i) begin g880 <= g4514; end
	always @ (posedge clk_i) begin g881 <= g4515; end
	always @ (posedge clk_i) begin g882 <= g4516; end
	always @ (posedge clk_i) begin g883 <= g4517; end
	always @ (posedge clk_i) begin g885 <= g4518; end
	always @ (posedge clk_i) begin g886 <= g4519; end
	always @ (posedge clk_i) begin g887 <= g4520; end
	always @ (posedge clk_i) begin g888 <= g4521; end
	always @ (posedge clk_i) begin g891 <= g4522; end
	always @ (posedge clk_i) begin g892 <= g4523; end
	always @ (posedge clk_i) begin g893 <= g4524; end
	always @ (posedge clk_i) begin g894 <= g4525; end
	always @ (posedge clk_i) begin g896 <= g4526; end
	always @ (posedge clk_i) begin g897 <= g4527; end
	always @ (posedge clk_i) begin g898 <= g4528; end
	always @ (posedge clk_i) begin g900 <= g4529; end
	always @ (posedge clk_i) begin g901 <= g4530; end
	always @ (posedge clk_i) begin g902 <= g4531; end
	always @ (posedge clk_i) begin g903 <= g4532; end
	always @ (posedge clk_i) begin g905 <= g4533; end
	always @ (posedge clk_i) begin g906 <= g4534; end
	always @ (posedge clk_i) begin g907 <= g4535; end
	always @ (posedge clk_i) begin g908 <= g4536; end
	always @ (posedge clk_i) begin g912 <= g4537; end
	always @ (posedge clk_i) begin g918 <= g4538; end
	always @ (posedge clk_i) begin g919 <= g4539; end
	always @ (posedge clk_i) begin g920 <= g4540; end
	always @ (posedge clk_i) begin g921 <= g4541; end
	always @ (posedge clk_i) begin g923 <= g4542; end
	always @ (posedge clk_i) begin g924 <= g4543; end
	always @ (posedge clk_i) begin g925 <= g4544; end
	always @ (posedge clk_i) begin g926 <= g4545; end
	always @ (posedge clk_i) begin g928 <= g4546; end
	always @ (posedge clk_i) begin g929 <= g4547; end
	always @ (posedge clk_i) begin g930 <= g4548; end
	always @ (posedge clk_i) begin g931 <= g4549; end
	always @ (posedge clk_i) begin g933 <= g4550; end
	always @ (posedge clk_i) begin g934 <= g4551; end
	always @ (posedge clk_i) begin g935 <= g4552; end
	always @ (posedge clk_i) begin g936 <= g4553; end
	always @ (posedge clk_i) begin g939 <= g4554; end
	always @ (posedge clk_i) begin g940 <= g4555; end
	always @ (posedge clk_i) begin g941 <= g4556; end
	always @ (posedge clk_i) begin g942 <= g4557; end
	always @ (posedge clk_i) begin g944 <= g4558; end
	always @ (posedge clk_i) begin g945 <= g4559; end
	always @ (posedge clk_i) begin g946 <= g4560; end
	always @ (posedge clk_i) begin g948 <= g4561; end
	always @ (posedge clk_i) begin g949 <= g4562; end
	always @ (posedge clk_i) begin g950 <= g4563; end
	always @ (posedge clk_i) begin g951 <= g4564; end
	always @ (posedge clk_i) begin g953 <= g4565; end
	always @ (posedge clk_i) begin g954 <= g4566; end
	always @ (posedge clk_i) begin g955 <= g4567; end
	always @ (posedge clk_i) begin g956 <= g4568; end
	always @ (posedge clk_i) begin g960 <= g4569; end
	always @ (posedge clk_i) begin g963 <= g4570; end
	always @ (posedge clk_i) begin g964 <= g4571; end
	always @ (posedge clk_i) begin g965 <= g4572; end
	always @ (posedge clk_i) begin g966 <= g4573; end
	always @ (posedge clk_i) begin g968 <= g4574; end
	always @ (posedge clk_i) begin g969 <= g4575; end
	always @ (posedge clk_i) begin g970 <= g4576; end
	always @ (posedge clk_i) begin g971 <= g4577; end
	always @ (posedge clk_i) begin g973 <= g4578; end
	always @ (posedge clk_i) begin g974 <= g4579; end
	always @ (posedge clk_i) begin g975 <= g4580; end
	always @ (posedge clk_i) begin g976 <= g4581; end
	always @ (posedge clk_i) begin g978 <= g4582; end
	always @ (posedge clk_i) begin g979 <= g4583; end
	always @ (posedge clk_i) begin g980 <= g4584; end
	always @ (posedge clk_i) begin g981 <= g4585; end
	always @ (posedge clk_i) begin g984 <= g4586; end
	always @ (posedge clk_i) begin g985 <= g4587; end
	always @ (posedge clk_i) begin g986 <= g4588; end
	always @ (posedge clk_i) begin g987 <= g4589; end
	always @ (posedge clk_i) begin g989 <= g4590; end
	always @ (posedge clk_i) begin g990 <= g4591; end
	always @ (posedge clk_i) begin g991 <= g4592; end
	always @ (posedge clk_i) begin g993 <= g4593; end
	always @ (posedge clk_i) begin g994 <= g4594; end
	always @ (posedge clk_i) begin g995 <= g4595; end
	always @ (posedge clk_i) begin g996 <= g4596; end
	always @ (posedge clk_i) begin g998 <= g4597; end
	always @ (posedge clk_i) begin g999 <= g4598; end
	always @ (posedge clk_i) begin g1000 <= g4599; end
	always @ (posedge clk_i) begin g1001 <= g4600; end
	always @ (posedge clk_i) begin g1005 <= g4601; end
	always @ (posedge clk_i) begin g1008 <= g4602; end
	always @ (posedge clk_i) begin g1009 <= g4603; end
	always @ (posedge clk_i) begin g1010 <= g4604; end
	always @ (posedge clk_i) begin g1011 <= g4605; end
	always @ (posedge clk_i) begin g1013 <= g4606; end
	always @ (posedge clk_i) begin g1014 <= g4607; end
	always @ (posedge clk_i) begin g1015 <= g4608; end
	always @ (posedge clk_i) begin g1016 <= g4609; end
	always @ (posedge clk_i) begin g1018 <= g4610; end
	always @ (posedge clk_i) begin g1019 <= g4611; end
	always @ (posedge clk_i) begin g1020 <= g4612; end
	always @ (posedge clk_i) begin g1021 <= g4613; end
	always @ (posedge clk_i) begin g1023 <= g4614; end
	always @ (posedge clk_i) begin g1024 <= g4615; end
	always @ (posedge clk_i) begin g1025 <= g4616; end
	always @ (posedge clk_i) begin g1026 <= g4617; end
	always @ (posedge clk_i) begin g1029 <= g4618; end
	always @ (posedge clk_i) begin g1030 <= g4619; end
	always @ (posedge clk_i) begin g1031 <= g4620; end
	always @ (posedge clk_i) begin g1032 <= g4621; end
	always @ (posedge clk_i) begin g1034 <= g4622; end
	always @ (posedge clk_i) begin g1035 <= g4623; end
	always @ (posedge clk_i) begin g1036 <= g4624; end
	always @ (posedge clk_i) begin g1038 <= g4625; end
	always @ (posedge clk_i) begin g1039 <= g4626; end
	always @ (posedge clk_i) begin g1040 <= g4627; end
	always @ (posedge clk_i) begin g1041 <= g4628; end
	always @ (posedge clk_i) begin g1043 <= g4629; end
	always @ (posedge clk_i) begin g1044 <= g4630; end
	always @ (posedge clk_i) begin g1045 <= g4631; end
	always @ (posedge clk_i) begin g1046 <= g4632; end
	always @ (posedge clk_i) begin g1050 <= g4633; end
	always @ (posedge clk_i) begin g1053 <= g4634; end
	always @ (posedge clk_i) begin g1054 <= g4635; end
	always @ (posedge clk_i) begin g1055 <= g4636; end
	always @ (posedge clk_i) begin g1056 <= g4637; end
	always @ (posedge clk_i) begin g1058 <= g4638; end
	always @ (posedge clk_i) begin g1059 <= g4639; end
	always @ (posedge clk_i) begin g1060 <= g4640; end
	always @ (posedge clk_i) begin g1061 <= g4641; end
	always @ (posedge clk_i) begin g1063 <= g4642; end
	always @ (posedge clk_i) begin g1064 <= g4643; end
	always @ (posedge clk_i) begin g1065 <= g4644; end
	always @ (posedge clk_i) begin g1066 <= g4645; end
	always @ (posedge clk_i) begin g1068 <= g4646; end
	always @ (posedge clk_i) begin g1069 <= g4647; end
	always @ (posedge clk_i) begin g1070 <= g4648; end
	always @ (posedge clk_i) begin g1071 <= g4649; end
	always @ (posedge clk_i) begin g1074 <= g4650; end
	always @ (posedge clk_i) begin g1075 <= g4651; end
	always @ (posedge clk_i) begin g1076 <= g4652; end
	always @ (posedge clk_i) begin g1077 <= g4653; end
	always @ (posedge clk_i) begin g1079 <= g4654; end
	always @ (posedge clk_i) begin g1080 <= g4655; end
	always @ (posedge clk_i) begin g1081 <= g4656; end
	always @ (posedge clk_i) begin g1083 <= g4657; end
	always @ (posedge clk_i) begin g1084 <= g4658; end
	always @ (posedge clk_i) begin g1085 <= g4659; end
	always @ (posedge clk_i) begin g1086 <= g4660; end
	always @ (posedge clk_i) begin g1088 <= g4661; end
	always @ (posedge clk_i) begin g1089 <= g4662; end
	always @ (posedge clk_i) begin g1090 <= g4663; end
	always @ (posedge clk_i) begin g1091 <= g4664; end
	always @ (posedge clk_i) begin g1095 <= g4665; end
	always @ (posedge clk_i) begin g1098 <= g4666; end
	always @ (posedge clk_i) begin g1099 <= g4667; end
	always @ (posedge clk_i) begin g1100 <= g4668; end
	always @ (posedge clk_i) begin g1101 <= g4669; end
	always @ (posedge clk_i) begin g1103 <= g4670; end
	always @ (posedge clk_i) begin g1104 <= g4671; end
	always @ (posedge clk_i) begin g1105 <= g4672; end
	always @ (posedge clk_i) begin g1106 <= g4673; end
	always @ (posedge clk_i) begin g1108 <= g4674; end
	always @ (posedge clk_i) begin g1109 <= g4675; end
	always @ (posedge clk_i) begin g1110 <= g4676; end
	always @ (posedge clk_i) begin g1111 <= g4677; end
	always @ (posedge clk_i) begin g1113 <= g4678; end
	always @ (posedge clk_i) begin g1114 <= g4679; end
	always @ (posedge clk_i) begin g1115 <= g4680; end
	always @ (posedge clk_i) begin g1116 <= g4681; end
	always @ (posedge clk_i) begin g1119 <= g4682; end
	always @ (posedge clk_i) begin g1120 <= g4683; end
	always @ (posedge clk_i) begin g1121 <= g4684; end
	always @ (posedge clk_i) begin g1122 <= g4685; end
	always @ (posedge clk_i) begin g1124 <= g4686; end
	always @ (posedge clk_i) begin g1125 <= g4687; end
	always @ (posedge clk_i) begin g1126 <= g4688; end
	always @ (posedge clk_i) begin g1128 <= g4689; end
	always @ (posedge clk_i) begin g1129 <= g4690; end
	always @ (posedge clk_i) begin g1130 <= g4691; end
	always @ (posedge clk_i) begin g1131 <= g4692; end
	always @ (posedge clk_i) begin g1133 <= g4693; end
	always @ (posedge clk_i) begin g1134 <= g4694; end
	always @ (posedge clk_i) begin g1135 <= g4695; end
	always @ (posedge clk_i) begin g1136 <= g4696; end
	always @ (posedge clk_i) begin g1140 <= g4697; end
	always @ (posedge clk_i) begin g1143 <= g4698; end
	always @ (posedge clk_i) begin g1144 <= g4699; end
	always @ (posedge clk_i) begin g1145 <= g4700; end
	always @ (posedge clk_i) begin g1146 <= g4701; end
	always @ (posedge clk_i) begin g1148 <= g4702; end
	always @ (posedge clk_i) begin g1149 <= g4703; end
	always @ (posedge clk_i) begin g1150 <= g4704; end
	always @ (posedge clk_i) begin g1151 <= g4705; end
	always @ (posedge clk_i) begin g1153 <= g4706; end
	always @ (posedge clk_i) begin g1154 <= g4707; end
	always @ (posedge clk_i) begin g1155 <= g4708; end
	always @ (posedge clk_i) begin g1156 <= g4709; end
	always @ (posedge clk_i) begin g1158 <= g4710; end
	always @ (posedge clk_i) begin g1159 <= g4711; end
	always @ (posedge clk_i) begin g1160 <= g4712; end
	always @ (posedge clk_i) begin g1161 <= g4713; end
	always @ (posedge clk_i) begin g1164 <= g4714; end
	always @ (posedge clk_i) begin g1165 <= g4715; end
	always @ (posedge clk_i) begin g1166 <= g4716; end
	always @ (posedge clk_i) begin g1167 <= g4717; end
	always @ (posedge clk_i) begin g1169 <= g4718; end
	always @ (posedge clk_i) begin g1170 <= g4719; end
	always @ (posedge clk_i) begin g1171 <= g4720; end
	always @ (posedge clk_i) begin g1173 <= g4721; end
	always @ (posedge clk_i) begin g1174 <= g4722; end
	always @ (posedge clk_i) begin g1175 <= g4723; end
	always @ (posedge clk_i) begin g1176 <= g4724; end
	always @ (posedge clk_i) begin g1178 <= g4725; end
	always @ (posedge clk_i) begin g1179 <= g4726; end
	always @ (posedge clk_i) begin g1180 <= g4727; end
	always @ (posedge clk_i) begin g1181 <= g4728; end
	always @ (posedge clk_i) begin g1185 <= g4729; end
	always @ (posedge clk_i) begin g1188 <= g4730; end
	always @ (posedge clk_i) begin g1189 <= g4731; end
	always @ (posedge clk_i) begin g1190 <= g4732; end
	always @ (posedge clk_i) begin g1191 <= g4733; end
	always @ (posedge clk_i) begin g1193 <= g4734; end
	always @ (posedge clk_i) begin g1194 <= g4735; end
	always @ (posedge clk_i) begin g1195 <= g4736; end
	always @ (posedge clk_i) begin g1196 <= g4737; end
	always @ (posedge clk_i) begin g1198 <= g4738; end
	always @ (posedge clk_i) begin g1199 <= g4739; end
	always @ (posedge clk_i) begin g1200 <= g4740; end
	always @ (posedge clk_i) begin g1201 <= g4741; end
	always @ (posedge clk_i) begin g1203 <= g4742; end
	always @ (posedge clk_i) begin g1204 <= g4743; end
	always @ (posedge clk_i) begin g1205 <= g4744; end
	always @ (posedge clk_i) begin g1206 <= g4745; end
	always @ (posedge clk_i) begin g1209 <= g4746; end
	always @ (posedge clk_i) begin g1210 <= g4747; end
	always @ (posedge clk_i) begin g1211 <= g4748; end
	always @ (posedge clk_i) begin g1212 <= g4749; end
	always @ (posedge clk_i) begin g1214 <= g4750; end
	always @ (posedge clk_i) begin g1215 <= g4751; end
	always @ (posedge clk_i) begin g1216 <= g4752; end
	always @ (posedge clk_i) begin g1218 <= g4753; end
	always @ (posedge clk_i) begin g1219 <= g4754; end
	always @ (posedge clk_i) begin g1220 <= g4755; end
	always @ (posedge clk_i) begin g1221 <= g4756; end
	always @ (posedge clk_i) begin g1223 <= g4757; end
	always @ (posedge clk_i) begin g1224 <= g4758; end
	always @ (posedge clk_i) begin g1225 <= g4759; end
	always @ (posedge clk_i) begin g1226 <= g4760; end
	always @ (posedge clk_i) begin g1230 <= g4761; end
	always @ (posedge clk_i) begin g1233 <= g4762; end
	always @ (posedge clk_i) begin g1234 <= g4763; end
	always @ (posedge clk_i) begin g1235 <= g4764; end
	always @ (posedge clk_i) begin g1236 <= g4765; end
	always @ (posedge clk_i) begin g1238 <= g4766; end
	always @ (posedge clk_i) begin g1239 <= g4767; end
	always @ (posedge clk_i) begin g1240 <= g4768; end
	always @ (posedge clk_i) begin g1241 <= g4769; end
	always @ (posedge clk_i) begin g1243 <= g4770; end
	always @ (posedge clk_i) begin g1244 <= g4771; end
	always @ (posedge clk_i) begin g1245 <= g4772; end
	always @ (posedge clk_i) begin g1246 <= g4773; end
	always @ (posedge clk_i) begin g1248 <= g4774; end
	always @ (posedge clk_i) begin g1249 <= g4775; end
	always @ (posedge clk_i) begin g1250 <= g4776; end
	always @ (posedge clk_i) begin g1251 <= g4777; end
	always @ (posedge clk_i) begin g1254 <= g4778; end
	always @ (posedge clk_i) begin g1255 <= g4779; end
	always @ (posedge clk_i) begin g1256 <= g4780; end
	always @ (posedge clk_i) begin g1257 <= g4781; end
	always @ (posedge clk_i) begin g1259 <= g4782; end
	always @ (posedge clk_i) begin g1260 <= g4783; end
	always @ (posedge clk_i) begin g1261 <= g4784; end
	always @ (posedge clk_i) begin g1263 <= g4785; end
	always @ (posedge clk_i) begin g1264 <= g4786; end
	always @ (posedge clk_i) begin g1265 <= g4787; end
	always @ (posedge clk_i) begin g1266 <= g4788; end
	always @ (posedge clk_i) begin g1268 <= g4789; end
	always @ (posedge clk_i) begin g1269 <= g4790; end
	always @ (posedge clk_i) begin g1270 <= g4791; end
	always @ (posedge clk_i) begin g1271 <= g4792; end
	always @ (posedge clk_i) begin g1275 <= g4793; end
	always @ (posedge clk_i) begin g1278 <= g4794; end
	always @ (posedge clk_i) begin g1279 <= g4795; end
	always @ (posedge clk_i) begin g1280 <= g4796; end
	always @ (posedge clk_i) begin g1281 <= g4797; end
	always @ (posedge clk_i) begin g1283 <= g4798; end
	always @ (posedge clk_i) begin g1284 <= g4799; end
	always @ (posedge clk_i) begin g1285 <= g4800; end
	always @ (posedge clk_i) begin g1286 <= g4801; end
	always @ (posedge clk_i) begin g1288 <= g4802; end
	always @ (posedge clk_i) begin g1289 <= g4803; end
	always @ (posedge clk_i) begin g1290 <= g4804; end
	always @ (posedge clk_i) begin g1291 <= g4805; end
	always @ (posedge clk_i) begin g1293 <= g4806; end
	always @ (posedge clk_i) begin g1294 <= g4807; end
	always @ (posedge clk_i) begin g1295 <= g4808; end
	always @ (posedge clk_i) begin g1296 <= g4809; end
	always @ (posedge clk_i) begin g1299 <= g4810; end
	always @ (posedge clk_i) begin g1300 <= g4811; end
	always @ (posedge clk_i) begin g1301 <= g4812; end
	always @ (posedge clk_i) begin g1302 <= g4813; end
	always @ (posedge clk_i) begin g1304 <= g4814; end
	always @ (posedge clk_i) begin g1305 <= g4815; end
	always @ (posedge clk_i) begin g1306 <= g4816; end
	always @ (posedge clk_i) begin g1308 <= g4817; end
	always @ (posedge clk_i) begin g1309 <= g4818; end
	always @ (posedge clk_i) begin g1310 <= g4819; end
	always @ (posedge clk_i) begin g1311 <= g4820; end
	always @ (posedge clk_i) begin g1313 <= g4821; end
	always @ (posedge clk_i) begin g1314 <= g4822; end
	always @ (posedge clk_i) begin g1315 <= g4823; end
	always @ (posedge clk_i) begin g1316 <= g4824; end
	always @ (posedge clk_i) begin g1320 <= g4825; end
	always @ (posedge clk_i) begin g1323 <= g4826; end
	always @ (posedge clk_i) begin g1324 <= g4827; end
	always @ (posedge clk_i) begin g1325 <= g4828; end
	always @ (posedge clk_i) begin g1326 <= g4829; end
	always @ (posedge clk_i) begin g1328 <= g4830; end
	always @ (posedge clk_i) begin g1329 <= g4831; end
	always @ (posedge clk_i) begin g1330 <= g4832; end
	always @ (posedge clk_i) begin g1331 <= g4833; end
	always @ (posedge clk_i) begin g1333 <= g4834; end
	always @ (posedge clk_i) begin g1334 <= g4835; end
	always @ (posedge clk_i) begin g1335 <= g4836; end
	always @ (posedge clk_i) begin g1336 <= g4837; end
	always @ (posedge clk_i) begin g1338 <= g4838; end
	always @ (posedge clk_i) begin g1339 <= g4839; end
	always @ (posedge clk_i) begin g1340 <= g4840; end
	always @ (posedge clk_i) begin g1341 <= g4841; end
	always @ (posedge clk_i) begin g1344 <= g4842; end
	always @ (posedge clk_i) begin g1345 <= g4843; end
	always @ (posedge clk_i) begin g1346 <= g4844; end
	always @ (posedge clk_i) begin g1347 <= g4845; end
	always @ (posedge clk_i) begin g1349 <= g4846; end
	always @ (posedge clk_i) begin g1350 <= g4847; end
	always @ (posedge clk_i) begin g1351 <= g4848; end
	always @ (posedge clk_i) begin g1353 <= g4849; end
	always @ (posedge clk_i) begin g1354 <= g4850; end
	always @ (posedge clk_i) begin g1355 <= g4851; end
	always @ (posedge clk_i) begin g1356 <= g4852; end
	always @ (posedge clk_i) begin g1358 <= g4853; end
	always @ (posedge clk_i) begin g1359 <= g4854; end
	always @ (posedge clk_i) begin g1360 <= g4855; end
	always @ (posedge clk_i) begin g1361 <= g4856; end
	always @ (posedge clk_i) begin g1365 <= g4857; end
	always @ (posedge clk_i) begin g1368 <= g4858; end
	always @ (posedge clk_i) begin g1369 <= g4859; end
	always @ (posedge clk_i) begin g1370 <= g4860; end
	always @ (posedge clk_i) begin g1371 <= g4861; end
	always @ (posedge clk_i) begin g1373 <= g4862; end
	always @ (posedge clk_i) begin g1374 <= g4863; end
	always @ (posedge clk_i) begin g1375 <= g4864; end
	always @ (posedge clk_i) begin g1376 <= g4865; end
	always @ (posedge clk_i) begin g1378 <= g4866; end
	always @ (posedge clk_i) begin g1379 <= g4867; end
	always @ (posedge clk_i) begin g1380 <= g4868; end
	always @ (posedge clk_i) begin g1381 <= g4869; end
	always @ (posedge clk_i) begin g1383 <= g4870; end
	always @ (posedge clk_i) begin g1384 <= g4871; end
	always @ (posedge clk_i) begin g1385 <= g4872; end
	always @ (posedge clk_i) begin g1386 <= g4873; end
	always @ (posedge clk_i) begin g1389 <= g4874; end
	always @ (posedge clk_i) begin g1390 <= g4875; end
	always @ (posedge clk_i) begin g1391 <= g4876; end
	always @ (posedge clk_i) begin g1392 <= g4877; end
	always @ (posedge clk_i) begin g1394 <= g4878; end
	always @ (posedge clk_i) begin g1395 <= g4879; end
	always @ (posedge clk_i) begin g1396 <= g4880; end
	always @ (posedge clk_i) begin g1398 <= g4881; end
	always @ (posedge clk_i) begin g1399 <= g4882; end
	always @ (posedge clk_i) begin g1400 <= g4883; end
	always @ (posedge clk_i) begin g1401 <= g4884; end
	always @ (posedge clk_i) begin g1403 <= g4885; end
	always @ (posedge clk_i) begin g1404 <= g4886; end
	always @ (posedge clk_i) begin g1405 <= g4887; end
	always @ (posedge clk_i) begin g1406 <= g4888; end
	always @ (posedge clk_i) begin g1410 <= g4889; end
	always @ (posedge clk_i) begin g1413 <= g4890; end
	always @ (posedge clk_i) begin g1414 <= g4891; end
	always @ (posedge clk_i) begin g1415 <= g4892; end
	always @ (posedge clk_i) begin g1416 <= g4893; end
	always @ (posedge clk_i) begin g1418 <= g4894; end
	always @ (posedge clk_i) begin g1419 <= g4895; end
	always @ (posedge clk_i) begin g1420 <= g4896; end
	always @ (posedge clk_i) begin g1421 <= g4897; end
	always @ (posedge clk_i) begin g1423 <= g4898; end
	always @ (posedge clk_i) begin g1424 <= g4899; end
	always @ (posedge clk_i) begin g1425 <= g4900; end
	always @ (posedge clk_i) begin g1426 <= g4901; end
	always @ (posedge clk_i) begin g1428 <= g4902; end
	always @ (posedge clk_i) begin g1429 <= g4903; end
	always @ (posedge clk_i) begin g1430 <= g4904; end
	always @ (posedge clk_i) begin g1431 <= g4905; end
	always @ (posedge clk_i) begin g1434 <= g4906; end
	always @ (posedge clk_i) begin g1435 <= g4907; end
	always @ (posedge clk_i) begin g1436 <= g4908; end
	always @ (posedge clk_i) begin g1437 <= g4909; end
	always @ (posedge clk_i) begin g1439 <= g4910; end
	always @ (posedge clk_i) begin g1440 <= g4911; end
	always @ (posedge clk_i) begin g1441 <= g4912; end
	always @ (posedge clk_i) begin g1443 <= g4913; end
	always @ (posedge clk_i) begin g1444 <= g4914; end
	always @ (posedge clk_i) begin g1445 <= g4915; end
	always @ (posedge clk_i) begin g1446 <= g4916; end
	always @ (posedge clk_i) begin g1448 <= g4917; end
	always @ (posedge clk_i) begin g1449 <= g4918; end
	always @ (posedge clk_i) begin g1450 <= g4919; end
	always @ (posedge clk_i) begin g1451 <= g4920; end
	always @ (posedge clk_i) begin g1455 <= g4921; end
	always @ (posedge clk_i) begin g1458 <= g4922; end
	always @ (posedge clk_i) begin g1459 <= g4923; end
	always @ (posedge clk_i) begin g1460 <= g4924; end
	always @ (posedge clk_i) begin g1461 <= g4925; end
	always @ (posedge clk_i) begin g1463 <= g4926; end
	always @ (posedge clk_i) begin g1464 <= g4927; end
	always @ (posedge clk_i) begin g1465 <= g4928; end
	always @ (posedge clk_i) begin g1466 <= g4929; end
	always @ (posedge clk_i) begin g1468 <= g4930; end
	always @ (posedge clk_i) begin g1469 <= g4931; end
	always @ (posedge clk_i) begin g1470 <= g4932; end
	always @ (posedge clk_i) begin g1471 <= g4933; end
	always @ (posedge clk_i) begin g1473 <= g4934; end
	always @ (posedge clk_i) begin g1474 <= g4935; end
	always @ (posedge clk_i) begin g1475 <= g4936; end
	always @ (posedge clk_i) begin g1476 <= g4937; end
	always @ (posedge clk_i) begin g1479 <= g4938; end
	always @ (posedge clk_i) begin g1480 <= g4939; end
	always @ (posedge clk_i) begin g1481 <= g4940; end
	always @ (posedge clk_i) begin g1482 <= g4941; end
	always @ (posedge clk_i) begin g1484 <= g4942; end
	always @ (posedge clk_i) begin g1485 <= g4943; end
	always @ (posedge clk_i) begin g1486 <= g4944; end
	always @ (posedge clk_i) begin g1488 <= g4945; end
	always @ (posedge clk_i) begin g1489 <= g4946; end
	always @ (posedge clk_i) begin g1490 <= g4947; end
	always @ (posedge clk_i) begin g1491 <= g4948; end
	always @ (posedge clk_i) begin g1493 <= g4949; end
	always @ (posedge clk_i) begin g1494 <= g4950; end
	always @ (posedge clk_i) begin g1495 <= g4951; end
	always @ (posedge clk_i) begin g1496 <= g4952; end
	always @ (posedge clk_i) begin g1500 <= g4953; end
	always @ (posedge clk_i) begin g1502 <= g4954; end
	always @ (posedge clk_i) begin g1503 <= g4955; end
	always @ (posedge clk_i) begin g1504 <= g4956; end
	always @ (posedge clk_i) begin g1505 <= g4957; end
	always @ (posedge clk_i) begin g1507 <= g4958; end
	always @ (posedge clk_i) begin g1508 <= g4959; end
	always @ (posedge clk_i) begin g1509 <= g4960; end
	always @ (posedge clk_i) begin g1510 <= g4961; end
	always @ (posedge clk_i) begin g1512 <= g4962; end
	always @ (posedge clk_i) begin g1513 <= g4963; end
	always @ (posedge clk_i) begin g1514 <= g4964; end
	always @ (posedge clk_i) begin g1515 <= g4965; end
	always @ (posedge clk_i) begin g1517 <= g4966; end
	always @ (posedge clk_i) begin g1518 <= g4967; end
	always @ (posedge clk_i) begin g1519 <= g4968; end
	always @ (posedge clk_i) begin g1520 <= g4969; end
	always @ (posedge clk_i) begin g1523 <= g4970; end
	always @ (posedge clk_i) begin g1524 <= g4971; end
	always @ (posedge clk_i) begin g1525 <= g4972; end
	always @ (posedge clk_i) begin g1526 <= g4973; end
	always @ (posedge clk_i) begin g1528 <= g4974; end
	always @ (posedge clk_i) begin g1529 <= g4975; end
	always @ (posedge clk_i) begin g1530 <= g4976; end
	always @ (posedge clk_i) begin g1532 <= g4977; end
	always @ (posedge clk_i) begin g1533 <= g4978; end
	always @ (posedge clk_i) begin g1534 <= g4979; end
	always @ (posedge clk_i) begin g1535 <= g4980; end
	always @ (posedge clk_i) begin g1537 <= g4981; end
	always @ (posedge clk_i) begin g1538 <= g4982; end
	always @ (posedge clk_i) begin g1539 <= g4983; end
	always @ (posedge clk_i) begin g1540 <= g4984; end
	always @ (posedge clk_i) begin g1544 <= g4985; end
	always @ (posedge clk_i) begin g1547 <= g4986; end
	always @ (posedge clk_i) begin g1548 <= g4987; end
	always @ (posedge clk_i) begin g1549 <= g4988; end
	always @ (posedge clk_i) begin g1550 <= g4989; end
	always @ (posedge clk_i) begin g1551 <= g4990; end
	always @ (posedge clk_i) begin g1553 <= g4991; end
	always @ (posedge clk_i) begin g1554 <= g4992; end
	always @ (posedge clk_i) begin g1555 <= g4993; end
	always @ (posedge clk_i) begin g1556 <= g4994; end
	always @ (posedge clk_i) begin g1558 <= g4995; end
	always @ (posedge clk_i) begin g1559 <= g4996; end
	always @ (posedge clk_i) begin g1560 <= g4997; end
	always @ (posedge clk_i) begin g1561 <= g4998; end
	always @ (posedge clk_i) begin g1563 <= g4999; end
	always @ (posedge clk_i) begin g1564 <= g5000; end
	always @ (posedge clk_i) begin g1565 <= g5001; end
	always @ (posedge clk_i) begin g1566 <= g5002; end
	always @ (posedge clk_i) begin g1569 <= g5003; end
	always @ (posedge clk_i) begin g1570 <= g5004; end
	always @ (posedge clk_i) begin g1571 <= g5005; end
	always @ (posedge clk_i) begin g1572 <= g5006; end
	always @ (posedge clk_i) begin g1574 <= g5007; end
	always @ (posedge clk_i) begin g1575 <= g5008; end
	always @ (posedge clk_i) begin g1576 <= g5009; end
	always @ (posedge clk_i) begin g1578 <= g5010; end
	always @ (posedge clk_i) begin g1579 <= g5011; end
	always @ (posedge clk_i) begin g1580 <= g5012; end
	always @ (posedge clk_i) begin g1581 <= g5013; end
	always @ (posedge clk_i) begin g1583 <= g5014; end
	always @ (posedge clk_i) begin g1584 <= g5015; end
	always @ (posedge clk_i) begin g1585 <= g5016; end
	always @ (posedge clk_i) begin g1586 <= g5017; end
	always @ (posedge clk_i) begin g2019 <= g2842; end
	always @ (posedge clk_i) begin g2023 <= g2844; end
	always @ (posedge clk_i) begin g2026 <= g5018; end
	always @ (posedge clk_i) begin g2035 <= g5019; end
	always @ (posedge clk_i) begin g2038 <= g5020; end
	always @ (posedge clk_i) begin g2055 <= g5021; end
	always @ (posedge clk_i) begin g2060 <= g5022; end
	always @ (posedge clk_i) begin g2066 <= g5023; end
	always @ (posedge clk_i) begin g2070 <= g2953; end
	always @ (posedge clk_i) begin g2071 <= g2964; end
	always @ (posedge clk_i) begin g2073 <= g2965; end
	always @ (posedge clk_i) begin g2074 <= g2966; end
	always @ (posedge clk_i) begin g2076 <= g2967; end
	always @ (posedge clk_i) begin g2077 <= g2968; end
	always @ (posedge clk_i) begin g2079 <= g5024; end
	always @ (posedge clk_i) begin g2080 <= g2975; end
	always @ (posedge clk_i) begin g2081 <= g2976; end
	always @ (posedge clk_i) begin g2083 <= g2982; end
	always @ (posedge clk_i) begin g2084 <= g2984; end
	always @ (posedge clk_i) begin g2085 <= g2986; end
	always @ (posedge clk_i) begin g2086 <= g2988; end
	always @ (posedge clk_i) begin g2088 <= g2990; end
	always @ (posedge clk_i) begin g2089 <= g2992; end
	always @ (posedge clk_i) begin g2090 <= g2994; end
	always @ (posedge clk_i) begin g2091 <= g2996; end
	always @ (posedge clk_i) begin g2093 <= g2998; end
	always @ (posedge clk_i) begin g2094 <= g3000; end
	always @ (posedge clk_i) begin g2095 <= g3002; end
	always @ (posedge clk_i) begin g2096 <= g3004; end
	always @ (posedge clk_i) begin g2098 <= g3006; end
	always @ (posedge clk_i) begin g2099 <= g3008; end
	always @ (posedge clk_i) begin g2100 <= g3010; end
	always @ (posedge clk_i) begin g2101 <= g3012; end
	always @ (posedge clk_i) begin g2104 <= g3014; end
	always @ (posedge clk_i) begin g2105 <= g3020; end
	always @ (posedge clk_i) begin g2106 <= g3022; end
	always @ (posedge clk_i) begin g2108 <= g3024; end
	always @ (posedge clk_i) begin g2109 <= g3025; end
	always @ (posedge clk_i) begin g2110 <= g3029; end
	always @ (posedge clk_i) begin g2111 <= g3030; end
	always @ (posedge clk_i) begin g2113 <= g3032; end
	always @ (posedge clk_i) begin g2114 <= g3034; end
	always @ (posedge clk_i) begin g2115 <= g3036; end
	always @ (posedge clk_i) begin g2116 <= g3038; end
	always @ (posedge clk_i) begin g2118 <= g3039; end
	always @ (posedge clk_i) begin g2119 <= g3040; end
	always @ (posedge clk_i) begin g2120 <= g3041; end
	always @ (posedge clk_i) begin g2121 <= g3042; end
	always @ (posedge clk_i) begin g2124 <= g3044; end
	always @ (posedge clk_i) begin g2125 <= g3047; end
	always @ (posedge clk_i) begin g2128 <= g5025; end
	always @ (posedge clk_i) begin g2129 <= g5026; end
	always @ (posedge clk_i) begin g2134 <= g3051; end
	always @ (posedge clk_i) begin g2135 <= g3052; end
	always @ (posedge clk_i) begin g2136 <= g3053; end
	always @ (posedge clk_i) begin g2137 <= g3054; end
	always @ (posedge clk_i) begin g2138 <= g3055; end
	always @ (posedge clk_i) begin g2231 <= g5027; end
	always @ (posedge clk_i) begin g2258 <= g5028; end
	always @ (posedge clk_i) begin g2284 <= g5029; end
	always @ (posedge clk_i) begin g2289 <= g3059; end
	always @ (posedge clk_i) begin g2306 <= g5030; end
	always @ (posedge clk_i) begin g2312 <= g3065; end
	always @ (posedge clk_i) begin g2333 <= g5031; end
	always @ (posedge clk_i) begin g2340 <= g3067; end
	always @ (posedge clk_i) begin g2357 <= g5032; end
	always @ (posedge clk_i) begin g2365 <= g3069; end
	always @ (posedge clk_i) begin g2383 <= g5033; end
	always @ (posedge clk_i) begin g2391 <= g3071; end
	always @ (posedge clk_i) begin g2413 <= g5034; end
	always @ (posedge clk_i) begin g2418 <= g3074; end
	always @ (posedge clk_i) begin g2432 <= g5035; end
	always @ (posedge clk_i) begin g2439 <= g3076; end
	always @ (posedge clk_i) begin g2457 <= g3077; end
	always @ (posedge clk_i) begin g2476 <= g5036; end
	always @ (posedge clk_i) begin g2482 <= g3078; end
	always @ (posedge clk_i) begin g2499 <= g5037; end
	always @ (posedge clk_i) begin g2507 <= g3081; end
	always @ (posedge clk_i) begin g2523 <= g5038; end
	always @ (posedge clk_i) begin g2529 <= g3082; end
	always @ (posedge clk_i) begin g2544 <= g5039; end
	always @ (posedge clk_i) begin g2551 <= g3085; end
	always @ (posedge clk_i) begin g2566 <= g5040; end
	always @ (posedge clk_i) begin g2570 <= g3088; end
	always @ (posedge clk_i) begin g2587 <= g5041; end
	always @ (posedge clk_i) begin g2590 <= g3089; end
	always @ (posedge clk_i) begin g2605 <= g5042; end
	always @ (posedge clk_i) begin g2608 <= g3090; end
	always @ (posedge clk_i) begin g2622 <= g5043; end
	always @ (posedge clk_i) begin g2625 <= g3092; end
	always @ (posedge clk_i) begin g2639 <= g5044; end
	always @ (posedge clk_i) begin g2642 <= g3094; end
	always @ (posedge clk_i) begin g2657 <= g5045; end
	always @ (posedge clk_i) begin g2660 <= g3095; end
	always @ (posedge clk_i) begin g2677 <= g5046; end
	always @ (posedge clk_i) begin g2680 <= g3099; end
	always @ (posedge clk_i) begin g2696 <= g5047; end
	always @ (posedge clk_i) begin g2699 <= g3100; end
	always @ (posedge clk_i) begin g2712 <= g5048; end
	always @ (posedge clk_i) begin g2715 <= g3102; end
	always @ (posedge clk_i) begin g2731 <= g5049; end
	always @ (posedge clk_i) begin g2734 <= g3104; end
	always @ (posedge clk_i) begin g2748 <= g5050; end
	always @ (posedge clk_i) begin g2751 <= g3105; end
	always @ (posedge clk_i) begin g2767 <= g5051; end
	always @ (posedge clk_i) begin g2771 <= g3106; end
	always @ (posedge clk_i) begin g2791 <= g5052; end
	always @ (posedge clk_i) begin g2794 <= g3108; end
	always @ (posedge clk_i) begin g2808 <= g5053; end
	always @ (posedge clk_i) begin g2811 <= g3110; end
	always @ (posedge clk_i) begin g2824 <= g5054; end
	always @ (posedge clk_i) begin g2827 <= g5055; end
	always @ (posedge clk_i) begin g2831 <= g3113; end
	always @ (posedge clk_i) begin g2914 <= g5056; end
	always @ (posedge clk_i) begin g2969 <= g5057; end

	assign fault_o = (((sk[0]) & (g1)));
	assign imem_addr_ox0x = (((sk[1]) & (gnd)));
	assign imem_addr_ox1x = (((sk[2]) & (gnd)));
	assign imem_addr_ox2x = (((sk[3]) & (gnd)));
	assign imem_addr_ox3x = (((sk[4]) & (gnd)));
	assign imem_addr_ox4x = (((sk[5]) & (gnd)));
	assign imem_addr_ox5x = (((sk[6]) & (gnd)));
	assign imem_addr_ox6x = (((sk[7]) & (gnd)));
	assign imem_addr_ox7x = (((sk[8]) & (gnd)));
	assign imem_addr_ox8x = (((sk[9]) & (gnd)));
	assign imem_addr_ox9x = (((sk[10]) & (gnd)));
	assign imem_addr_ox10x = (((sk[11]) & (gnd)));
	assign imem_addr_ox11x = (((sk[12]) & (gnd)));
	assign imem_addr_ox12x = (((sk[13]) & (gnd)));
	assign imem_addr_ox13x = (((sk[14]) & (gnd)));
	assign imem_addr_ox14x = (((sk[15]) & (gnd)));
	assign imem_addr_ox15x = (((sk[16]) & (gnd)));
	assign imem_addr_ox16x = (((sk[17]) & (gnd)));
	assign imem_addr_ox17x = (((sk[18]) & (gnd)));
	assign imem_addr_ox18x = (((sk[19]) & (gnd)));
	assign imem_addr_ox19x = (((sk[20]) & (gnd)));
	assign imem_addr_ox20x = (((sk[21]) & (gnd)));
	assign imem_addr_ox21x = (((sk[22]) & (gnd)));
	assign imem_addr_ox22x = (((sk[23]) & (gnd)));
	assign imem_addr_ox23x = (((sk[24]) & (gnd)));
	assign imem_addr_ox24x = (((sk[25]) & (gnd)));
	assign imem_addr_ox25x = (((sk[26]) & (gnd)));
	assign imem_addr_ox26x = (((sk[27]) & (gnd)));
	assign imem_addr_ox27x = (((sk[28]) & (gnd)));
	assign imem_addr_ox28x = (((sk[29]) & (gnd)));
	assign imem_addr_ox29x = (((sk[30]) & (gnd)));
	assign imem_addr_ox30x = (((sk[31]) & (gnd)));
	assign imem_addr_ox31x = (((sk[32]) & (gnd)));
	assign imem_cti_ox0x = (((sk[33]) & (gnd)));
	assign imem_cti_ox1x = (((sk[34]) & (gnd)));
	assign imem_cti_ox2x = (((sk[35]) & (gnd)));
	assign imem_cyc_o = (((sk[36]) & (gnd)));
	assign imem_stb_o = (((sk[37]) & (gnd)));
	assign dmem_dat_ox0x = (((sk[38]) & (g35)));
	assign dmem_dat_ox1x = (((sk[39]) & (g36)));
	assign dmem_dat_ox2x = (((sk[40]) & (g37)));
	assign dmem_dat_ox3x = (((sk[41]) & (g38)));
	assign dmem_dat_ox4x = (((sk[42]) & (g39)));
	assign dmem_dat_ox5x = (((sk[43]) & (g40)));
	assign dmem_dat_ox6x = (((sk[44]) & (g41)));
	assign dmem_dat_ox7x = (((sk[45]) & (g42)));
	assign dmem_dat_ox8x = (((sk[46]) & (g43)));
	assign dmem_dat_ox9x = (((sk[47]) & (g44)));
	assign dmem_dat_ox10x = (((sk[48]) & (g45)));
	assign dmem_dat_ox11x = (((sk[49]) & (g46)));
	assign dmem_dat_ox12x = (((sk[50]) & (g47)));
	assign dmem_dat_ox13x = (((sk[51]) & (g48)));
	assign dmem_dat_ox14x = (((sk[52]) & (g49)));
	assign dmem_dat_ox15x = (((sk[53]) & (g50)));
	assign dmem_dat_ox16x = (((sk[54]) & (g51)));
	assign dmem_dat_ox17x = (((sk[55]) & (g52)));
	assign dmem_dat_ox18x = (((sk[56]) & (g53)));
	assign dmem_dat_ox19x = (((sk[57]) & (g54)));
	assign dmem_dat_ox20x = (((sk[58]) & (g55)));
	assign dmem_dat_ox21x = (((sk[59]) & (g56)));
	assign dmem_dat_ox22x = (((sk[60]) & (g57)));
	assign dmem_dat_ox23x = (((sk[61]) & (g58)));
	assign dmem_dat_ox24x = (((sk[62]) & (g59)));
	assign dmem_dat_ox25x = (((sk[63]) & (g60)));
	assign dmem_dat_ox26x = (((sk[64]) & (g61)));
	assign dmem_dat_ox27x = (((sk[65]) & (g62)));
	assign dmem_dat_ox28x = (((sk[66]) & (g63)));
	assign dmem_dat_ox29x = (((sk[67]) & (g64)));
	assign dmem_dat_ox30x = (((sk[68]) & (g65)));
	assign dmem_dat_ox31x = (((sk[69]) & (g66)));
	assign dmem_cti_ox0x = (((sk[70]) & (vcc)));
	assign dmem_cti_ox1x = (((sk[71]) & (vcc)));
	assign dmem_cti_ox2x = (((sk[72]) & (vcc)));
	assign dmem_cyc_o = (((sk[73]) & (g67)));
	assign dmem_stb_o = (((sk[74]) & (g68)));
	assign dmem_we_o = (((sk[75]) & (g69)));
	assign g3893 = (((!g139) & (sk[76]) & (g127) & (!dmem_addr_ox0x)) + ((!g139) & (sk[76]) & (g127) & (dmem_addr_ox0x)) + ((g139) & (!sk[76]) & (!g127) & (!dmem_addr_ox0x)) + ((g139) & (!sk[76]) & (!g127) & (dmem_addr_ox0x)) + ((g139) & (!sk[76]) & (g127) & (!dmem_addr_ox0x)) + ((g139) & (!sk[76]) & (g127) & (dmem_addr_ox0x)) + ((g139) & (sk[76]) & (!g127) & (dmem_addr_ox0x)) + ((g139) & (sk[76]) & (g127) & (dmem_addr_ox0x)));
	assign g3894 = (((!g139) & (!sk[77]) & (!g140) & (dmem_addr_ox1x)) + ((!g139) & (!sk[77]) & (g140) & (!dmem_addr_ox1x)) + ((!g139) & (!sk[77]) & (g140) & (dmem_addr_ox1x)) + ((!g139) & (sk[77]) & (g140) & (!dmem_addr_ox1x)) + ((!g139) & (sk[77]) & (g140) & (dmem_addr_ox1x)) + ((g139) & (!sk[77]) & (!g140) & (dmem_addr_ox1x)) + ((g139) & (!sk[77]) & (g140) & (!dmem_addr_ox1x)) + ((g139) & (!sk[77]) & (g140) & (dmem_addr_ox1x)) + ((g139) & (sk[77]) & (!g140) & (dmem_addr_ox1x)) + ((g139) & (sk[77]) & (g140) & (dmem_addr_ox1x)));
	assign g3895 = (((!sk[78]) & (!g139) & (!g274) & (dmem_addr_ox2x)) + ((!sk[78]) & (!g139) & (g274) & (!dmem_addr_ox2x)) + ((!sk[78]) & (!g139) & (g274) & (dmem_addr_ox2x)) + ((!sk[78]) & (g139) & (!g274) & (dmem_addr_ox2x)) + ((!sk[78]) & (g139) & (g274) & (!dmem_addr_ox2x)) + ((!sk[78]) & (g139) & (g274) & (dmem_addr_ox2x)) + ((sk[78]) & (!g139) & (g274) & (!dmem_addr_ox2x)) + ((sk[78]) & (!g139) & (g274) & (dmem_addr_ox2x)) + ((sk[78]) & (g139) & (!g274) & (dmem_addr_ox2x)) + ((sk[78]) & (g139) & (g274) & (dmem_addr_ox2x)));
	assign g3896 = (((!g139) & (!sk[79]) & (!g3882) & (dmem_addr_ox3x)) + ((!g139) & (!sk[79]) & (g3882) & (!dmem_addr_ox3x)) + ((!g139) & (!sk[79]) & (g3882) & (dmem_addr_ox3x)) + ((!g139) & (sk[79]) & (g3882) & (!dmem_addr_ox3x)) + ((!g139) & (sk[79]) & (g3882) & (dmem_addr_ox3x)) + ((g139) & (!sk[79]) & (!g3882) & (dmem_addr_ox3x)) + ((g139) & (!sk[79]) & (g3882) & (!dmem_addr_ox3x)) + ((g139) & (!sk[79]) & (g3882) & (dmem_addr_ox3x)) + ((g139) & (sk[79]) & (!g3882) & (dmem_addr_ox3x)) + ((g139) & (sk[79]) & (g3882) & (dmem_addr_ox3x)));
	assign g3897 = (((!sk[80]) & (!g139) & (!g363) & (dmem_addr_ox4x)) + ((!sk[80]) & (!g139) & (g363) & (!dmem_addr_ox4x)) + ((!sk[80]) & (!g139) & (g363) & (dmem_addr_ox4x)) + ((!sk[80]) & (g139) & (!g363) & (dmem_addr_ox4x)) + ((!sk[80]) & (g139) & (g363) & (!dmem_addr_ox4x)) + ((!sk[80]) & (g139) & (g363) & (dmem_addr_ox4x)) + ((sk[80]) & (!g139) & (g363) & (!dmem_addr_ox4x)) + ((sk[80]) & (!g139) & (g363) & (dmem_addr_ox4x)) + ((sk[80]) & (g139) & (!g363) & (dmem_addr_ox4x)) + ((sk[80]) & (g139) & (g363) & (dmem_addr_ox4x)));
	assign g3898 = (((!sk[81]) & (!g139) & (!g3871) & (dmem_addr_ox5x)) + ((!sk[81]) & (!g139) & (g3871) & (!dmem_addr_ox5x)) + ((!sk[81]) & (!g139) & (g3871) & (dmem_addr_ox5x)) + ((!sk[81]) & (g139) & (!g3871) & (dmem_addr_ox5x)) + ((!sk[81]) & (g139) & (g3871) & (!dmem_addr_ox5x)) + ((!sk[81]) & (g139) & (g3871) & (dmem_addr_ox5x)) + ((sk[81]) & (!g139) & (g3871) & (!dmem_addr_ox5x)) + ((sk[81]) & (!g139) & (g3871) & (dmem_addr_ox5x)) + ((sk[81]) & (g139) & (!g3871) & (dmem_addr_ox5x)) + ((sk[81]) & (g139) & (g3871) & (dmem_addr_ox5x)));
	assign g3899 = (((!g139) & (!sk[82]) & (!g452) & (dmem_addr_ox6x)) + ((!g139) & (!sk[82]) & (g452) & (!dmem_addr_ox6x)) + ((!g139) & (!sk[82]) & (g452) & (dmem_addr_ox6x)) + ((!g139) & (sk[82]) & (g452) & (!dmem_addr_ox6x)) + ((!g139) & (sk[82]) & (g452) & (dmem_addr_ox6x)) + ((g139) & (!sk[82]) & (!g452) & (dmem_addr_ox6x)) + ((g139) & (!sk[82]) & (g452) & (!dmem_addr_ox6x)) + ((g139) & (!sk[82]) & (g452) & (dmem_addr_ox6x)) + ((g139) & (sk[82]) & (!g452) & (dmem_addr_ox6x)) + ((g139) & (sk[82]) & (g452) & (dmem_addr_ox6x)));
	assign g3900 = (((!sk[83]) & (!g139) & (!g3860) & (dmem_addr_ox7x)) + ((!sk[83]) & (!g139) & (g3860) & (!dmem_addr_ox7x)) + ((!sk[83]) & (!g139) & (g3860) & (dmem_addr_ox7x)) + ((!sk[83]) & (g139) & (!g3860) & (dmem_addr_ox7x)) + ((!sk[83]) & (g139) & (g3860) & (!dmem_addr_ox7x)) + ((!sk[83]) & (g139) & (g3860) & (dmem_addr_ox7x)) + ((sk[83]) & (!g139) & (g3860) & (!dmem_addr_ox7x)) + ((sk[83]) & (!g139) & (g3860) & (dmem_addr_ox7x)) + ((sk[83]) & (g139) & (!g3860) & (dmem_addr_ox7x)) + ((sk[83]) & (g139) & (g3860) & (dmem_addr_ox7x)));
	assign g3901 = (((!g139) & (!sk[84]) & (!g540) & (dmem_addr_ox8x)) + ((!g139) & (!sk[84]) & (g540) & (!dmem_addr_ox8x)) + ((!g139) & (!sk[84]) & (g540) & (dmem_addr_ox8x)) + ((!g139) & (sk[84]) & (g540) & (!dmem_addr_ox8x)) + ((!g139) & (sk[84]) & (g540) & (dmem_addr_ox8x)) + ((g139) & (!sk[84]) & (!g540) & (dmem_addr_ox8x)) + ((g139) & (!sk[84]) & (g540) & (!dmem_addr_ox8x)) + ((g139) & (!sk[84]) & (g540) & (dmem_addr_ox8x)) + ((g139) & (sk[84]) & (!g540) & (dmem_addr_ox8x)) + ((g139) & (sk[84]) & (g540) & (dmem_addr_ox8x)));
	assign g3902 = (((!sk[85]) & (!g139) & (!g585) & (dmem_addr_ox9x)) + ((!sk[85]) & (!g139) & (g585) & (!dmem_addr_ox9x)) + ((!sk[85]) & (!g139) & (g585) & (dmem_addr_ox9x)) + ((!sk[85]) & (g139) & (!g585) & (dmem_addr_ox9x)) + ((!sk[85]) & (g139) & (g585) & (!dmem_addr_ox9x)) + ((!sk[85]) & (g139) & (g585) & (dmem_addr_ox9x)) + ((sk[85]) & (!g139) & (g585) & (!dmem_addr_ox9x)) + ((sk[85]) & (!g139) & (g585) & (dmem_addr_ox9x)) + ((sk[85]) & (g139) & (!g585) & (dmem_addr_ox9x)) + ((sk[85]) & (g139) & (g585) & (dmem_addr_ox9x)));
	assign g3903 = (((!sk[86]) & (!g139) & (!g3849) & (dmem_addr_ox10x)) + ((!sk[86]) & (!g139) & (g3849) & (!dmem_addr_ox10x)) + ((!sk[86]) & (!g139) & (g3849) & (dmem_addr_ox10x)) + ((!sk[86]) & (g139) & (!g3849) & (dmem_addr_ox10x)) + ((!sk[86]) & (g139) & (g3849) & (!dmem_addr_ox10x)) + ((!sk[86]) & (g139) & (g3849) & (dmem_addr_ox10x)) + ((sk[86]) & (!g139) & (g3849) & (!dmem_addr_ox10x)) + ((sk[86]) & (!g139) & (g3849) & (dmem_addr_ox10x)) + ((sk[86]) & (g139) & (!g3849) & (dmem_addr_ox10x)) + ((sk[86]) & (g139) & (g3849) & (dmem_addr_ox10x)));
	assign g3904 = (((!g139) & (!g681) & (!sk[87]) & (dmem_addr_ox11x)) + ((!g139) & (g681) & (!sk[87]) & (!dmem_addr_ox11x)) + ((!g139) & (g681) & (!sk[87]) & (dmem_addr_ox11x)) + ((!g139) & (g681) & (sk[87]) & (!dmem_addr_ox11x)) + ((!g139) & (g681) & (sk[87]) & (dmem_addr_ox11x)) + ((g139) & (!g681) & (!sk[87]) & (dmem_addr_ox11x)) + ((g139) & (!g681) & (sk[87]) & (dmem_addr_ox11x)) + ((g139) & (g681) & (!sk[87]) & (!dmem_addr_ox11x)) + ((g139) & (g681) & (!sk[87]) & (dmem_addr_ox11x)) + ((g139) & (g681) & (sk[87]) & (dmem_addr_ox11x)));
	assign g3905 = (((!g139) & (!g728) & (!sk[88]) & (dmem_addr_ox12x)) + ((!g139) & (g728) & (!sk[88]) & (!dmem_addr_ox12x)) + ((!g139) & (g728) & (!sk[88]) & (dmem_addr_ox12x)) + ((!g139) & (g728) & (sk[88]) & (!dmem_addr_ox12x)) + ((!g139) & (g728) & (sk[88]) & (dmem_addr_ox12x)) + ((g139) & (!g728) & (!sk[88]) & (dmem_addr_ox12x)) + ((g139) & (!g728) & (sk[88]) & (dmem_addr_ox12x)) + ((g139) & (g728) & (!sk[88]) & (!dmem_addr_ox12x)) + ((g139) & (g728) & (!sk[88]) & (dmem_addr_ox12x)) + ((g139) & (g728) & (sk[88]) & (dmem_addr_ox12x)));
	assign g3906 = (((!sk[89]) & (!g139) & (!g775) & (dmem_addr_ox13x)) + ((!sk[89]) & (!g139) & (g775) & (!dmem_addr_ox13x)) + ((!sk[89]) & (!g139) & (g775) & (dmem_addr_ox13x)) + ((!sk[89]) & (g139) & (!g775) & (dmem_addr_ox13x)) + ((!sk[89]) & (g139) & (g775) & (!dmem_addr_ox13x)) + ((!sk[89]) & (g139) & (g775) & (dmem_addr_ox13x)) + ((sk[89]) & (!g139) & (g775) & (!dmem_addr_ox13x)) + ((sk[89]) & (!g139) & (g775) & (dmem_addr_ox13x)) + ((sk[89]) & (g139) & (!g775) & (dmem_addr_ox13x)) + ((sk[89]) & (g139) & (g775) & (dmem_addr_ox13x)));
	assign g3907 = (((!g139) & (!g822) & (!sk[90]) & (dmem_addr_ox14x)) + ((!g139) & (g822) & (!sk[90]) & (!dmem_addr_ox14x)) + ((!g139) & (g822) & (!sk[90]) & (dmem_addr_ox14x)) + ((!g139) & (g822) & (sk[90]) & (!dmem_addr_ox14x)) + ((!g139) & (g822) & (sk[90]) & (dmem_addr_ox14x)) + ((g139) & (!g822) & (!sk[90]) & (dmem_addr_ox14x)) + ((g139) & (!g822) & (sk[90]) & (dmem_addr_ox14x)) + ((g139) & (g822) & (!sk[90]) & (!dmem_addr_ox14x)) + ((g139) & (g822) & (!sk[90]) & (dmem_addr_ox14x)) + ((g139) & (g822) & (sk[90]) & (dmem_addr_ox14x)));
	assign g3908 = (((!g139) & (!g869) & (!sk[91]) & (dmem_addr_ox15x)) + ((!g139) & (g869) & (!sk[91]) & (!dmem_addr_ox15x)) + ((!g139) & (g869) & (!sk[91]) & (dmem_addr_ox15x)) + ((!g139) & (g869) & (sk[91]) & (!dmem_addr_ox15x)) + ((!g139) & (g869) & (sk[91]) & (dmem_addr_ox15x)) + ((g139) & (!g869) & (!sk[91]) & (dmem_addr_ox15x)) + ((g139) & (!g869) & (sk[91]) & (dmem_addr_ox15x)) + ((g139) & (g869) & (!sk[91]) & (!dmem_addr_ox15x)) + ((g139) & (g869) & (!sk[91]) & (dmem_addr_ox15x)) + ((g139) & (g869) & (sk[91]) & (dmem_addr_ox15x)));
	assign g3909 = (((!g139) & (!g917) & (!sk[92]) & (dmem_addr_ox16x)) + ((!g139) & (g917) & (!sk[92]) & (!dmem_addr_ox16x)) + ((!g139) & (g917) & (!sk[92]) & (dmem_addr_ox16x)) + ((!g139) & (g917) & (sk[92]) & (!dmem_addr_ox16x)) + ((!g139) & (g917) & (sk[92]) & (dmem_addr_ox16x)) + ((g139) & (!g917) & (!sk[92]) & (dmem_addr_ox16x)) + ((g139) & (!g917) & (sk[92]) & (dmem_addr_ox16x)) + ((g139) & (g917) & (!sk[92]) & (!dmem_addr_ox16x)) + ((g139) & (g917) & (!sk[92]) & (dmem_addr_ox16x)) + ((g139) & (g917) & (sk[92]) & (dmem_addr_ox16x)));
	assign g3910 = (((!g139) & (!g962) & (!sk[93]) & (dmem_addr_ox17x)) + ((!g139) & (g962) & (!sk[93]) & (!dmem_addr_ox17x)) + ((!g139) & (g962) & (!sk[93]) & (dmem_addr_ox17x)) + ((!g139) & (g962) & (sk[93]) & (!dmem_addr_ox17x)) + ((!g139) & (g962) & (sk[93]) & (dmem_addr_ox17x)) + ((g139) & (!g962) & (!sk[93]) & (dmem_addr_ox17x)) + ((g139) & (!g962) & (sk[93]) & (dmem_addr_ox17x)) + ((g139) & (g962) & (!sk[93]) & (!dmem_addr_ox17x)) + ((g139) & (g962) & (!sk[93]) & (dmem_addr_ox17x)) + ((g139) & (g962) & (sk[93]) & (dmem_addr_ox17x)));
	assign g3911 = (((!sk[94]) & (!g139) & (!g1007) & (dmem_addr_ox18x)) + ((!sk[94]) & (!g139) & (g1007) & (!dmem_addr_ox18x)) + ((!sk[94]) & (!g139) & (g1007) & (dmem_addr_ox18x)) + ((!sk[94]) & (g139) & (!g1007) & (dmem_addr_ox18x)) + ((!sk[94]) & (g139) & (g1007) & (!dmem_addr_ox18x)) + ((!sk[94]) & (g139) & (g1007) & (dmem_addr_ox18x)) + ((sk[94]) & (!g139) & (g1007) & (!dmem_addr_ox18x)) + ((sk[94]) & (!g139) & (g1007) & (dmem_addr_ox18x)) + ((sk[94]) & (g139) & (!g1007) & (dmem_addr_ox18x)) + ((sk[94]) & (g139) & (g1007) & (dmem_addr_ox18x)));
	assign g3912 = (((!g139) & (!g1052) & (!sk[95]) & (dmem_addr_ox19x)) + ((!g139) & (g1052) & (!sk[95]) & (!dmem_addr_ox19x)) + ((!g139) & (g1052) & (!sk[95]) & (dmem_addr_ox19x)) + ((!g139) & (g1052) & (sk[95]) & (!dmem_addr_ox19x)) + ((!g139) & (g1052) & (sk[95]) & (dmem_addr_ox19x)) + ((g139) & (!g1052) & (!sk[95]) & (dmem_addr_ox19x)) + ((g139) & (!g1052) & (sk[95]) & (dmem_addr_ox19x)) + ((g139) & (g1052) & (!sk[95]) & (!dmem_addr_ox19x)) + ((g139) & (g1052) & (!sk[95]) & (dmem_addr_ox19x)) + ((g139) & (g1052) & (sk[95]) & (dmem_addr_ox19x)));
	assign g3913 = (((!sk[96]) & (!g139) & (!g1097) & (dmem_addr_ox20x)) + ((!sk[96]) & (!g139) & (g1097) & (!dmem_addr_ox20x)) + ((!sk[96]) & (!g139) & (g1097) & (dmem_addr_ox20x)) + ((!sk[96]) & (g139) & (!g1097) & (dmem_addr_ox20x)) + ((!sk[96]) & (g139) & (g1097) & (!dmem_addr_ox20x)) + ((!sk[96]) & (g139) & (g1097) & (dmem_addr_ox20x)) + ((sk[96]) & (!g139) & (g1097) & (!dmem_addr_ox20x)) + ((sk[96]) & (!g139) & (g1097) & (dmem_addr_ox20x)) + ((sk[96]) & (g139) & (!g1097) & (dmem_addr_ox20x)) + ((sk[96]) & (g139) & (g1097) & (dmem_addr_ox20x)));
	assign g3914 = (((!g139) & (!g1142) & (!sk[97]) & (dmem_addr_ox21x)) + ((!g139) & (g1142) & (!sk[97]) & (!dmem_addr_ox21x)) + ((!g139) & (g1142) & (!sk[97]) & (dmem_addr_ox21x)) + ((!g139) & (g1142) & (sk[97]) & (!dmem_addr_ox21x)) + ((!g139) & (g1142) & (sk[97]) & (dmem_addr_ox21x)) + ((g139) & (!g1142) & (!sk[97]) & (dmem_addr_ox21x)) + ((g139) & (!g1142) & (sk[97]) & (dmem_addr_ox21x)) + ((g139) & (g1142) & (!sk[97]) & (!dmem_addr_ox21x)) + ((g139) & (g1142) & (!sk[97]) & (dmem_addr_ox21x)) + ((g139) & (g1142) & (sk[97]) & (dmem_addr_ox21x)));
	assign g3915 = (((!g139) & (!sk[98]) & (!g1187) & (dmem_addr_ox22x)) + ((!g139) & (!sk[98]) & (g1187) & (!dmem_addr_ox22x)) + ((!g139) & (!sk[98]) & (g1187) & (dmem_addr_ox22x)) + ((!g139) & (sk[98]) & (g1187) & (!dmem_addr_ox22x)) + ((!g139) & (sk[98]) & (g1187) & (dmem_addr_ox22x)) + ((g139) & (!sk[98]) & (!g1187) & (dmem_addr_ox22x)) + ((g139) & (!sk[98]) & (g1187) & (!dmem_addr_ox22x)) + ((g139) & (!sk[98]) & (g1187) & (dmem_addr_ox22x)) + ((g139) & (sk[98]) & (!g1187) & (dmem_addr_ox22x)) + ((g139) & (sk[98]) & (g1187) & (dmem_addr_ox22x)));
	assign g3916 = (((!g139) & (!g1232) & (!sk[99]) & (dmem_addr_ox23x)) + ((!g139) & (g1232) & (!sk[99]) & (!dmem_addr_ox23x)) + ((!g139) & (g1232) & (!sk[99]) & (dmem_addr_ox23x)) + ((!g139) & (g1232) & (sk[99]) & (!dmem_addr_ox23x)) + ((!g139) & (g1232) & (sk[99]) & (dmem_addr_ox23x)) + ((g139) & (!g1232) & (!sk[99]) & (dmem_addr_ox23x)) + ((g139) & (!g1232) & (sk[99]) & (dmem_addr_ox23x)) + ((g139) & (g1232) & (!sk[99]) & (!dmem_addr_ox23x)) + ((g139) & (g1232) & (!sk[99]) & (dmem_addr_ox23x)) + ((g139) & (g1232) & (sk[99]) & (dmem_addr_ox23x)));
	assign g3917 = (((!sk[100]) & (!g139) & (!g1277) & (dmem_addr_ox24x)) + ((!sk[100]) & (!g139) & (g1277) & (!dmem_addr_ox24x)) + ((!sk[100]) & (!g139) & (g1277) & (dmem_addr_ox24x)) + ((!sk[100]) & (g139) & (!g1277) & (dmem_addr_ox24x)) + ((!sk[100]) & (g139) & (g1277) & (!dmem_addr_ox24x)) + ((!sk[100]) & (g139) & (g1277) & (dmem_addr_ox24x)) + ((sk[100]) & (!g139) & (g1277) & (!dmem_addr_ox24x)) + ((sk[100]) & (!g139) & (g1277) & (dmem_addr_ox24x)) + ((sk[100]) & (g139) & (!g1277) & (dmem_addr_ox24x)) + ((sk[100]) & (g139) & (g1277) & (dmem_addr_ox24x)));
	assign g3918 = (((!g139) & (!g1322) & (!sk[101]) & (dmem_addr_ox25x)) + ((!g139) & (g1322) & (!sk[101]) & (!dmem_addr_ox25x)) + ((!g139) & (g1322) & (!sk[101]) & (dmem_addr_ox25x)) + ((!g139) & (g1322) & (sk[101]) & (!dmem_addr_ox25x)) + ((!g139) & (g1322) & (sk[101]) & (dmem_addr_ox25x)) + ((g139) & (!g1322) & (!sk[101]) & (dmem_addr_ox25x)) + ((g139) & (!g1322) & (sk[101]) & (dmem_addr_ox25x)) + ((g139) & (g1322) & (!sk[101]) & (!dmem_addr_ox25x)) + ((g139) & (g1322) & (!sk[101]) & (dmem_addr_ox25x)) + ((g139) & (g1322) & (sk[101]) & (dmem_addr_ox25x)));
	assign g3919 = (((!sk[102]) & (!g139) & (!g1367) & (dmem_addr_ox26x)) + ((!sk[102]) & (!g139) & (g1367) & (!dmem_addr_ox26x)) + ((!sk[102]) & (!g139) & (g1367) & (dmem_addr_ox26x)) + ((!sk[102]) & (g139) & (!g1367) & (dmem_addr_ox26x)) + ((!sk[102]) & (g139) & (g1367) & (!dmem_addr_ox26x)) + ((!sk[102]) & (g139) & (g1367) & (dmem_addr_ox26x)) + ((sk[102]) & (!g139) & (g1367) & (!dmem_addr_ox26x)) + ((sk[102]) & (!g139) & (g1367) & (dmem_addr_ox26x)) + ((sk[102]) & (g139) & (!g1367) & (dmem_addr_ox26x)) + ((sk[102]) & (g139) & (g1367) & (dmem_addr_ox26x)));
	assign g3920 = (((!g139) & (!sk[103]) & (!g1412) & (dmem_addr_ox27x)) + ((!g139) & (!sk[103]) & (g1412) & (!dmem_addr_ox27x)) + ((!g139) & (!sk[103]) & (g1412) & (dmem_addr_ox27x)) + ((!g139) & (sk[103]) & (g1412) & (!dmem_addr_ox27x)) + ((!g139) & (sk[103]) & (g1412) & (dmem_addr_ox27x)) + ((g139) & (!sk[103]) & (!g1412) & (dmem_addr_ox27x)) + ((g139) & (!sk[103]) & (g1412) & (!dmem_addr_ox27x)) + ((g139) & (!sk[103]) & (g1412) & (dmem_addr_ox27x)) + ((g139) & (sk[103]) & (!g1412) & (dmem_addr_ox27x)) + ((g139) & (sk[103]) & (g1412) & (dmem_addr_ox27x)));
	assign g3921 = (((!g139) & (!sk[104]) & (!g1457) & (dmem_addr_ox28x)) + ((!g139) & (!sk[104]) & (g1457) & (!dmem_addr_ox28x)) + ((!g139) & (!sk[104]) & (g1457) & (dmem_addr_ox28x)) + ((!g139) & (sk[104]) & (g1457) & (!dmem_addr_ox28x)) + ((!g139) & (sk[104]) & (g1457) & (dmem_addr_ox28x)) + ((g139) & (!sk[104]) & (!g1457) & (dmem_addr_ox28x)) + ((g139) & (!sk[104]) & (g1457) & (!dmem_addr_ox28x)) + ((g139) & (!sk[104]) & (g1457) & (dmem_addr_ox28x)) + ((g139) & (sk[104]) & (!g1457) & (dmem_addr_ox28x)) + ((g139) & (sk[104]) & (g1457) & (dmem_addr_ox28x)));
	assign g3922 = (((!g139) & (!sk[105]) & (!g1501) & (dmem_addr_ox29x)) + ((!g139) & (!sk[105]) & (g1501) & (!dmem_addr_ox29x)) + ((!g139) & (!sk[105]) & (g1501) & (dmem_addr_ox29x)) + ((!g139) & (sk[105]) & (g1501) & (!dmem_addr_ox29x)) + ((!g139) & (sk[105]) & (g1501) & (dmem_addr_ox29x)) + ((g139) & (!sk[105]) & (!g1501) & (dmem_addr_ox29x)) + ((g139) & (!sk[105]) & (g1501) & (!dmem_addr_ox29x)) + ((g139) & (!sk[105]) & (g1501) & (dmem_addr_ox29x)) + ((g139) & (sk[105]) & (!g1501) & (dmem_addr_ox29x)) + ((g139) & (sk[105]) & (g1501) & (dmem_addr_ox29x)));
	assign g3923 = (((!g139) & (!sk[106]) & (!g1546) & (dmem_addr_ox30x)) + ((!g139) & (!sk[106]) & (g1546) & (!dmem_addr_ox30x)) + ((!g139) & (!sk[106]) & (g1546) & (dmem_addr_ox30x)) + ((!g139) & (sk[106]) & (g1546) & (!dmem_addr_ox30x)) + ((!g139) & (sk[106]) & (g1546) & (dmem_addr_ox30x)) + ((g139) & (!sk[106]) & (!g1546) & (dmem_addr_ox30x)) + ((g139) & (!sk[106]) & (g1546) & (!dmem_addr_ox30x)) + ((g139) & (!sk[106]) & (g1546) & (dmem_addr_ox30x)) + ((g139) & (sk[106]) & (!g1546) & (dmem_addr_ox30x)) + ((g139) & (sk[106]) & (g1546) & (dmem_addr_ox30x)));
	assign g3924 = (((!g139) & (!sk[107]) & (!g1591) & (dmem_addr_ox31x)) + ((!g139) & (!sk[107]) & (g1591) & (!dmem_addr_ox31x)) + ((!g139) & (!sk[107]) & (g1591) & (dmem_addr_ox31x)) + ((!g139) & (sk[107]) & (g1591) & (!dmem_addr_ox31x)) + ((!g139) & (sk[107]) & (g1591) & (dmem_addr_ox31x)) + ((g139) & (!sk[107]) & (!g1591) & (dmem_addr_ox31x)) + ((g139) & (!sk[107]) & (g1591) & (!dmem_addr_ox31x)) + ((g139) & (!sk[107]) & (g1591) & (dmem_addr_ox31x)) + ((g139) & (sk[107]) & (!g1591) & (dmem_addr_ox31x)) + ((g139) & (sk[107]) & (g1591) & (dmem_addr_ox31x)));
	assign g3925 = (((!g1609) & (!g1608) & (!sk[108]) & (g35)) + ((!g1609) & (!g1608) & (sk[108]) & (g35)) + ((!g1609) & (g1608) & (!sk[108]) & (!g35)) + ((!g1609) & (g1608) & (!sk[108]) & (g35)) + ((!g1609) & (g1608) & (sk[108]) & (g35)) + ((g1609) & (!g1608) & (!sk[108]) & (g35)) + ((g1609) & (g1608) & (!sk[108]) & (!g35)) + ((g1609) & (g1608) & (!sk[108]) & (g35)) + ((g1609) & (g1608) & (sk[108]) & (!g35)) + ((g1609) & (g1608) & (sk[108]) & (g35)));
	assign g3926 = (((!sk[109]) & (!g1609) & (!g1621) & (g36)) + ((!sk[109]) & (!g1609) & (g1621) & (!g36)) + ((!sk[109]) & (!g1609) & (g1621) & (g36)) + ((!sk[109]) & (g1609) & (!g1621) & (g36)) + ((!sk[109]) & (g1609) & (g1621) & (!g36)) + ((!sk[109]) & (g1609) & (g1621) & (g36)) + ((sk[109]) & (!g1609) & (!g1621) & (g36)) + ((sk[109]) & (!g1609) & (g1621) & (g36)) + ((sk[109]) & (g1609) & (g1621) & (!g36)) + ((sk[109]) & (g1609) & (g1621) & (g36)));
	assign g3927 = (((!g1609) & (!sk[110]) & (!g1633) & (g37)) + ((!g1609) & (!sk[110]) & (g1633) & (!g37)) + ((!g1609) & (!sk[110]) & (g1633) & (g37)) + ((!g1609) & (sk[110]) & (!g1633) & (g37)) + ((!g1609) & (sk[110]) & (g1633) & (g37)) + ((g1609) & (!sk[110]) & (!g1633) & (g37)) + ((g1609) & (!sk[110]) & (g1633) & (!g37)) + ((g1609) & (!sk[110]) & (g1633) & (g37)) + ((g1609) & (sk[110]) & (g1633) & (!g37)) + ((g1609) & (sk[110]) & (g1633) & (g37)));
	assign g3928 = (((!g1609) & (!sk[111]) & (!g1645) & (g38)) + ((!g1609) & (!sk[111]) & (g1645) & (!g38)) + ((!g1609) & (!sk[111]) & (g1645) & (g38)) + ((!g1609) & (sk[111]) & (!g1645) & (g38)) + ((!g1609) & (sk[111]) & (g1645) & (g38)) + ((g1609) & (!sk[111]) & (!g1645) & (g38)) + ((g1609) & (!sk[111]) & (g1645) & (!g38)) + ((g1609) & (!sk[111]) & (g1645) & (g38)) + ((g1609) & (sk[111]) & (g1645) & (!g38)) + ((g1609) & (sk[111]) & (g1645) & (g38)));
	assign g3929 = (((!g1609) & (!g1657) & (!sk[112]) & (g39)) + ((!g1609) & (!g1657) & (sk[112]) & (g39)) + ((!g1609) & (g1657) & (!sk[112]) & (!g39)) + ((!g1609) & (g1657) & (!sk[112]) & (g39)) + ((!g1609) & (g1657) & (sk[112]) & (g39)) + ((g1609) & (!g1657) & (!sk[112]) & (g39)) + ((g1609) & (g1657) & (!sk[112]) & (!g39)) + ((g1609) & (g1657) & (!sk[112]) & (g39)) + ((g1609) & (g1657) & (sk[112]) & (!g39)) + ((g1609) & (g1657) & (sk[112]) & (g39)));
	assign g3930 = (((!g1609) & (!sk[113]) & (!g1669) & (g40)) + ((!g1609) & (!sk[113]) & (g1669) & (!g40)) + ((!g1609) & (!sk[113]) & (g1669) & (g40)) + ((!g1609) & (sk[113]) & (!g1669) & (g40)) + ((!g1609) & (sk[113]) & (g1669) & (g40)) + ((g1609) & (!sk[113]) & (!g1669) & (g40)) + ((g1609) & (!sk[113]) & (g1669) & (!g40)) + ((g1609) & (!sk[113]) & (g1669) & (g40)) + ((g1609) & (sk[113]) & (g1669) & (!g40)) + ((g1609) & (sk[113]) & (g1669) & (g40)));
	assign g3931 = (((!g1609) & (!g1681) & (!sk[114]) & (g41)) + ((!g1609) & (!g1681) & (sk[114]) & (g41)) + ((!g1609) & (g1681) & (!sk[114]) & (!g41)) + ((!g1609) & (g1681) & (!sk[114]) & (g41)) + ((!g1609) & (g1681) & (sk[114]) & (g41)) + ((g1609) & (!g1681) & (!sk[114]) & (g41)) + ((g1609) & (g1681) & (!sk[114]) & (!g41)) + ((g1609) & (g1681) & (!sk[114]) & (g41)) + ((g1609) & (g1681) & (sk[114]) & (!g41)) + ((g1609) & (g1681) & (sk[114]) & (g41)));
	assign g3932 = (((!sk[115]) & (!g1609) & (!g1693) & (g42)) + ((!sk[115]) & (!g1609) & (g1693) & (!g42)) + ((!sk[115]) & (!g1609) & (g1693) & (g42)) + ((!sk[115]) & (g1609) & (!g1693) & (g42)) + ((!sk[115]) & (g1609) & (g1693) & (!g42)) + ((!sk[115]) & (g1609) & (g1693) & (g42)) + ((sk[115]) & (!g1609) & (!g1693) & (g42)) + ((sk[115]) & (!g1609) & (g1693) & (g42)) + ((sk[115]) & (g1609) & (g1693) & (!g42)) + ((sk[115]) & (g1609) & (g1693) & (g42)));
	assign g3933 = (((!sk[116]) & (!g1609) & (!g1708) & (g43)) + ((!sk[116]) & (!g1609) & (g1708) & (!g43)) + ((!sk[116]) & (!g1609) & (g1708) & (g43)) + ((!sk[116]) & (g1609) & (!g1708) & (g43)) + ((!sk[116]) & (g1609) & (g1708) & (!g43)) + ((!sk[116]) & (g1609) & (g1708) & (g43)) + ((sk[116]) & (!g1609) & (!g1708) & (g43)) + ((sk[116]) & (!g1609) & (g1708) & (g43)) + ((sk[116]) & (g1609) & (g1708) & (!g43)) + ((sk[116]) & (g1609) & (g1708) & (g43)));
	assign g3934 = (((!g1609) & (!sk[117]) & (!g1721) & (g44)) + ((!g1609) & (!sk[117]) & (g1721) & (!g44)) + ((!g1609) & (!sk[117]) & (g1721) & (g44)) + ((!g1609) & (sk[117]) & (!g1721) & (g44)) + ((!g1609) & (sk[117]) & (g1721) & (g44)) + ((g1609) & (!sk[117]) & (!g1721) & (g44)) + ((g1609) & (!sk[117]) & (g1721) & (!g44)) + ((g1609) & (!sk[117]) & (g1721) & (g44)) + ((g1609) & (sk[117]) & (g1721) & (!g44)) + ((g1609) & (sk[117]) & (g1721) & (g44)));
	assign g3935 = (((!sk[118]) & (!g1609) & (!g1734) & (g45)) + ((!sk[118]) & (!g1609) & (g1734) & (!g45)) + ((!sk[118]) & (!g1609) & (g1734) & (g45)) + ((!sk[118]) & (g1609) & (!g1734) & (g45)) + ((!sk[118]) & (g1609) & (g1734) & (!g45)) + ((!sk[118]) & (g1609) & (g1734) & (g45)) + ((sk[118]) & (!g1609) & (!g1734) & (g45)) + ((sk[118]) & (!g1609) & (g1734) & (g45)) + ((sk[118]) & (g1609) & (g1734) & (!g45)) + ((sk[118]) & (g1609) & (g1734) & (g45)));
	assign g3936 = (((!g1609) & (!g1747) & (!sk[119]) & (g46)) + ((!g1609) & (!g1747) & (sk[119]) & (g46)) + ((!g1609) & (g1747) & (!sk[119]) & (!g46)) + ((!g1609) & (g1747) & (!sk[119]) & (g46)) + ((!g1609) & (g1747) & (sk[119]) & (g46)) + ((g1609) & (!g1747) & (!sk[119]) & (g46)) + ((g1609) & (g1747) & (!sk[119]) & (!g46)) + ((g1609) & (g1747) & (!sk[119]) & (g46)) + ((g1609) & (g1747) & (sk[119]) & (!g46)) + ((g1609) & (g1747) & (sk[119]) & (g46)));
	assign g3937 = (((!g1609) & (!sk[120]) & (!g1760) & (g47)) + ((!g1609) & (!sk[120]) & (g1760) & (!g47)) + ((!g1609) & (!sk[120]) & (g1760) & (g47)) + ((!g1609) & (sk[120]) & (!g1760) & (g47)) + ((!g1609) & (sk[120]) & (g1760) & (g47)) + ((g1609) & (!sk[120]) & (!g1760) & (g47)) + ((g1609) & (!sk[120]) & (g1760) & (!g47)) + ((g1609) & (!sk[120]) & (g1760) & (g47)) + ((g1609) & (sk[120]) & (g1760) & (!g47)) + ((g1609) & (sk[120]) & (g1760) & (g47)));
	assign g3938 = (((!sk[121]) & (!g1609) & (!g1773) & (g48)) + ((!sk[121]) & (!g1609) & (g1773) & (!g48)) + ((!sk[121]) & (!g1609) & (g1773) & (g48)) + ((!sk[121]) & (g1609) & (!g1773) & (g48)) + ((!sk[121]) & (g1609) & (g1773) & (!g48)) + ((!sk[121]) & (g1609) & (g1773) & (g48)) + ((sk[121]) & (!g1609) & (!g1773) & (g48)) + ((sk[121]) & (!g1609) & (g1773) & (g48)) + ((sk[121]) & (g1609) & (g1773) & (!g48)) + ((sk[121]) & (g1609) & (g1773) & (g48)));
	assign g3939 = (((!g1609) & (!sk[122]) & (!g1786) & (g49)) + ((!g1609) & (!sk[122]) & (g1786) & (!g49)) + ((!g1609) & (!sk[122]) & (g1786) & (g49)) + ((!g1609) & (sk[122]) & (!g1786) & (g49)) + ((!g1609) & (sk[122]) & (g1786) & (g49)) + ((g1609) & (!sk[122]) & (!g1786) & (g49)) + ((g1609) & (!sk[122]) & (g1786) & (!g49)) + ((g1609) & (!sk[122]) & (g1786) & (g49)) + ((g1609) & (sk[122]) & (g1786) & (!g49)) + ((g1609) & (sk[122]) & (g1786) & (g49)));
	assign g3940 = (((!g1609) & (!g1799) & (!sk[123]) & (g50)) + ((!g1609) & (!g1799) & (sk[123]) & (g50)) + ((!g1609) & (g1799) & (!sk[123]) & (!g50)) + ((!g1609) & (g1799) & (!sk[123]) & (g50)) + ((!g1609) & (g1799) & (sk[123]) & (g50)) + ((g1609) & (!g1799) & (!sk[123]) & (g50)) + ((g1609) & (g1799) & (!sk[123]) & (!g50)) + ((g1609) & (g1799) & (!sk[123]) & (g50)) + ((g1609) & (g1799) & (sk[123]) & (!g50)) + ((g1609) & (g1799) & (sk[123]) & (g50)));
	assign g3941 = (((!g1609) & (!g1813) & (!sk[124]) & (g51)) + ((!g1609) & (!g1813) & (sk[124]) & (g51)) + ((!g1609) & (g1813) & (!sk[124]) & (!g51)) + ((!g1609) & (g1813) & (!sk[124]) & (g51)) + ((!g1609) & (g1813) & (sk[124]) & (g51)) + ((g1609) & (!g1813) & (!sk[124]) & (g51)) + ((g1609) & (g1813) & (!sk[124]) & (!g51)) + ((g1609) & (g1813) & (!sk[124]) & (g51)) + ((g1609) & (g1813) & (sk[124]) & (!g51)) + ((g1609) & (g1813) & (sk[124]) & (g51)));
	assign g3942 = (((!sk[125]) & (!g1609) & (!g1826) & (g52)) + ((!sk[125]) & (!g1609) & (g1826) & (!g52)) + ((!sk[125]) & (!g1609) & (g1826) & (g52)) + ((!sk[125]) & (g1609) & (!g1826) & (g52)) + ((!sk[125]) & (g1609) & (g1826) & (!g52)) + ((!sk[125]) & (g1609) & (g1826) & (g52)) + ((sk[125]) & (!g1609) & (!g1826) & (g52)) + ((sk[125]) & (!g1609) & (g1826) & (g52)) + ((sk[125]) & (g1609) & (g1826) & (!g52)) + ((sk[125]) & (g1609) & (g1826) & (g52)));
	assign g3943 = (((!g1609) & (!g1839) & (!sk[126]) & (g53)) + ((!g1609) & (!g1839) & (sk[126]) & (g53)) + ((!g1609) & (g1839) & (!sk[126]) & (!g53)) + ((!g1609) & (g1839) & (!sk[126]) & (g53)) + ((!g1609) & (g1839) & (sk[126]) & (g53)) + ((g1609) & (!g1839) & (!sk[126]) & (g53)) + ((g1609) & (g1839) & (!sk[126]) & (!g53)) + ((g1609) & (g1839) & (!sk[126]) & (g53)) + ((g1609) & (g1839) & (sk[126]) & (!g53)) + ((g1609) & (g1839) & (sk[126]) & (g53)));
	assign g3944 = (((!g1609) & (!g1852) & (!sk[127]) & (g54)) + ((!g1609) & (!g1852) & (sk[127]) & (g54)) + ((!g1609) & (g1852) & (!sk[127]) & (!g54)) + ((!g1609) & (g1852) & (!sk[127]) & (g54)) + ((!g1609) & (g1852) & (sk[127]) & (g54)) + ((g1609) & (!g1852) & (!sk[127]) & (g54)) + ((g1609) & (g1852) & (!sk[127]) & (!g54)) + ((g1609) & (g1852) & (!sk[127]) & (g54)) + ((g1609) & (g1852) & (sk[127]) & (!g54)) + ((g1609) & (g1852) & (sk[127]) & (g54)));
	assign g3945 = (((!sk[0]) & (!g1609) & (!g1865) & (g55)) + ((!sk[0]) & (!g1609) & (g1865) & (!g55)) + ((!sk[0]) & (!g1609) & (g1865) & (g55)) + ((!sk[0]) & (g1609) & (!g1865) & (g55)) + ((!sk[0]) & (g1609) & (g1865) & (!g55)) + ((!sk[0]) & (g1609) & (g1865) & (g55)) + ((sk[0]) & (!g1609) & (!g1865) & (g55)) + ((sk[0]) & (!g1609) & (g1865) & (g55)) + ((sk[0]) & (g1609) & (g1865) & (!g55)) + ((sk[0]) & (g1609) & (g1865) & (g55)));
	assign g3946 = (((!g1609) & (!g1878) & (!sk[1]) & (g56)) + ((!g1609) & (!g1878) & (sk[1]) & (g56)) + ((!g1609) & (g1878) & (!sk[1]) & (!g56)) + ((!g1609) & (g1878) & (!sk[1]) & (g56)) + ((!g1609) & (g1878) & (sk[1]) & (g56)) + ((g1609) & (!g1878) & (!sk[1]) & (g56)) + ((g1609) & (g1878) & (!sk[1]) & (!g56)) + ((g1609) & (g1878) & (!sk[1]) & (g56)) + ((g1609) & (g1878) & (sk[1]) & (!g56)) + ((g1609) & (g1878) & (sk[1]) & (g56)));
	assign g3947 = (((!g1609) & (!g1891) & (!sk[2]) & (g57)) + ((!g1609) & (!g1891) & (sk[2]) & (g57)) + ((!g1609) & (g1891) & (!sk[2]) & (!g57)) + ((!g1609) & (g1891) & (!sk[2]) & (g57)) + ((!g1609) & (g1891) & (sk[2]) & (g57)) + ((g1609) & (!g1891) & (!sk[2]) & (g57)) + ((g1609) & (g1891) & (!sk[2]) & (!g57)) + ((g1609) & (g1891) & (!sk[2]) & (g57)) + ((g1609) & (g1891) & (sk[2]) & (!g57)) + ((g1609) & (g1891) & (sk[2]) & (g57)));
	assign g3948 = (((!g1609) & (!sk[3]) & (!g1904) & (g58)) + ((!g1609) & (!sk[3]) & (g1904) & (!g58)) + ((!g1609) & (!sk[3]) & (g1904) & (g58)) + ((!g1609) & (sk[3]) & (!g1904) & (g58)) + ((!g1609) & (sk[3]) & (g1904) & (g58)) + ((g1609) & (!sk[3]) & (!g1904) & (g58)) + ((g1609) & (!sk[3]) & (g1904) & (!g58)) + ((g1609) & (!sk[3]) & (g1904) & (g58)) + ((g1609) & (sk[3]) & (g1904) & (!g58)) + ((g1609) & (sk[3]) & (g1904) & (g58)));
	assign g3949 = (((!sk[4]) & (!g1609) & (!g1918) & (g59)) + ((!sk[4]) & (!g1609) & (g1918) & (!g59)) + ((!sk[4]) & (!g1609) & (g1918) & (g59)) + ((!sk[4]) & (g1609) & (!g1918) & (g59)) + ((!sk[4]) & (g1609) & (g1918) & (!g59)) + ((!sk[4]) & (g1609) & (g1918) & (g59)) + ((sk[4]) & (!g1609) & (!g1918) & (g59)) + ((sk[4]) & (!g1609) & (g1918) & (g59)) + ((sk[4]) & (g1609) & (g1918) & (!g59)) + ((sk[4]) & (g1609) & (g1918) & (g59)));
	assign g3950 = (((!g1609) & (!sk[5]) & (!g1931) & (g60)) + ((!g1609) & (!sk[5]) & (g1931) & (!g60)) + ((!g1609) & (!sk[5]) & (g1931) & (g60)) + ((!g1609) & (sk[5]) & (!g1931) & (g60)) + ((!g1609) & (sk[5]) & (g1931) & (g60)) + ((g1609) & (!sk[5]) & (!g1931) & (g60)) + ((g1609) & (!sk[5]) & (g1931) & (!g60)) + ((g1609) & (!sk[5]) & (g1931) & (g60)) + ((g1609) & (sk[5]) & (g1931) & (!g60)) + ((g1609) & (sk[5]) & (g1931) & (g60)));
	assign g3951 = (((!g1609) & (!sk[6]) & (!g1944) & (g61)) + ((!g1609) & (!sk[6]) & (g1944) & (!g61)) + ((!g1609) & (!sk[6]) & (g1944) & (g61)) + ((!g1609) & (sk[6]) & (!g1944) & (g61)) + ((!g1609) & (sk[6]) & (g1944) & (g61)) + ((g1609) & (!sk[6]) & (!g1944) & (g61)) + ((g1609) & (!sk[6]) & (g1944) & (!g61)) + ((g1609) & (!sk[6]) & (g1944) & (g61)) + ((g1609) & (sk[6]) & (g1944) & (!g61)) + ((g1609) & (sk[6]) & (g1944) & (g61)));
	assign g3952 = (((!g1609) & (!sk[7]) & (!g1957) & (g62)) + ((!g1609) & (!sk[7]) & (g1957) & (!g62)) + ((!g1609) & (!sk[7]) & (g1957) & (g62)) + ((!g1609) & (sk[7]) & (!g1957) & (g62)) + ((!g1609) & (sk[7]) & (g1957) & (g62)) + ((g1609) & (!sk[7]) & (!g1957) & (g62)) + ((g1609) & (!sk[7]) & (g1957) & (!g62)) + ((g1609) & (!sk[7]) & (g1957) & (g62)) + ((g1609) & (sk[7]) & (g1957) & (!g62)) + ((g1609) & (sk[7]) & (g1957) & (g62)));
	assign g3953 = (((!sk[8]) & (!g1609) & (!g1970) & (g63)) + ((!sk[8]) & (!g1609) & (g1970) & (!g63)) + ((!sk[8]) & (!g1609) & (g1970) & (g63)) + ((!sk[8]) & (g1609) & (!g1970) & (g63)) + ((!sk[8]) & (g1609) & (g1970) & (!g63)) + ((!sk[8]) & (g1609) & (g1970) & (g63)) + ((sk[8]) & (!g1609) & (!g1970) & (g63)) + ((sk[8]) & (!g1609) & (g1970) & (g63)) + ((sk[8]) & (g1609) & (g1970) & (!g63)) + ((sk[8]) & (g1609) & (g1970) & (g63)));
	assign g3954 = (((!g1609) & (!g1983) & (!sk[9]) & (g64)) + ((!g1609) & (!g1983) & (sk[9]) & (g64)) + ((!g1609) & (g1983) & (!sk[9]) & (!g64)) + ((!g1609) & (g1983) & (!sk[9]) & (g64)) + ((!g1609) & (g1983) & (sk[9]) & (g64)) + ((g1609) & (!g1983) & (!sk[9]) & (g64)) + ((g1609) & (g1983) & (!sk[9]) & (!g64)) + ((g1609) & (g1983) & (!sk[9]) & (g64)) + ((g1609) & (g1983) & (sk[9]) & (!g64)) + ((g1609) & (g1983) & (sk[9]) & (g64)));
	assign g3955 = (((!g1609) & (!sk[10]) & (!g1996) & (g65)) + ((!g1609) & (!sk[10]) & (g1996) & (!g65)) + ((!g1609) & (!sk[10]) & (g1996) & (g65)) + ((!g1609) & (sk[10]) & (!g1996) & (g65)) + ((!g1609) & (sk[10]) & (g1996) & (g65)) + ((g1609) & (!sk[10]) & (!g1996) & (g65)) + ((g1609) & (!sk[10]) & (g1996) & (!g65)) + ((g1609) & (!sk[10]) & (g1996) & (g65)) + ((g1609) & (sk[10]) & (g1996) & (!g65)) + ((g1609) & (sk[10]) & (g1996) & (g65)));
	assign g3956 = (((!sk[11]) & (!g1609) & (!g2009) & (g66)) + ((!sk[11]) & (!g1609) & (g2009) & (!g66)) + ((!sk[11]) & (!g1609) & (g2009) & (g66)) + ((!sk[11]) & (g1609) & (!g2009) & (g66)) + ((!sk[11]) & (g1609) & (g2009) & (!g66)) + ((!sk[11]) & (g1609) & (g2009) & (g66)) + ((sk[11]) & (!g1609) & (!g2009) & (g66)) + ((sk[11]) & (!g1609) & (g2009) & (g66)) + ((sk[11]) & (g1609) & (g2009) & (!g66)) + ((sk[11]) & (g1609) & (g2009) & (g66)));
	assign g3957 = (((!g2015) & (!sk[12]) & (!g2014) & (dmem_sel_ox0x)) + ((!g2015) & (!sk[12]) & (g2014) & (!dmem_sel_ox0x)) + ((!g2015) & (!sk[12]) & (g2014) & (dmem_sel_ox0x)) + ((!g2015) & (sk[12]) & (!g2014) & (dmem_sel_ox0x)) + ((!g2015) & (sk[12]) & (g2014) & (dmem_sel_ox0x)) + ((g2015) & (!sk[12]) & (!g2014) & (dmem_sel_ox0x)) + ((g2015) & (!sk[12]) & (g2014) & (!dmem_sel_ox0x)) + ((g2015) & (!sk[12]) & (g2014) & (dmem_sel_ox0x)) + ((g2015) & (sk[12]) & (g2014) & (!dmem_sel_ox0x)) + ((g2015) & (sk[12]) & (g2014) & (dmem_sel_ox0x)));
	assign g3958 = (((!g2015) & (!sk[13]) & (!g2016) & (dmem_sel_ox1x)) + ((!g2015) & (!sk[13]) & (g2016) & (!dmem_sel_ox1x)) + ((!g2015) & (!sk[13]) & (g2016) & (dmem_sel_ox1x)) + ((!g2015) & (sk[13]) & (!g2016) & (dmem_sel_ox1x)) + ((!g2015) & (sk[13]) & (g2016) & (dmem_sel_ox1x)) + ((g2015) & (!sk[13]) & (!g2016) & (dmem_sel_ox1x)) + ((g2015) & (!sk[13]) & (g2016) & (!dmem_sel_ox1x)) + ((g2015) & (!sk[13]) & (g2016) & (dmem_sel_ox1x)) + ((g2015) & (sk[13]) & (g2016) & (!dmem_sel_ox1x)) + ((g2015) & (sk[13]) & (g2016) & (dmem_sel_ox1x)));
	assign g3959 = (((!sk[14]) & (!g2015) & (!g2017) & (dmem_sel_ox2x)) + ((!sk[14]) & (!g2015) & (g2017) & (!dmem_sel_ox2x)) + ((!sk[14]) & (!g2015) & (g2017) & (dmem_sel_ox2x)) + ((!sk[14]) & (g2015) & (!g2017) & (dmem_sel_ox2x)) + ((!sk[14]) & (g2015) & (g2017) & (!dmem_sel_ox2x)) + ((!sk[14]) & (g2015) & (g2017) & (dmem_sel_ox2x)) + ((sk[14]) & (!g2015) & (!g2017) & (dmem_sel_ox2x)) + ((sk[14]) & (!g2015) & (g2017) & (dmem_sel_ox2x)) + ((sk[14]) & (g2015) & (g2017) & (!dmem_sel_ox2x)) + ((sk[14]) & (g2015) & (g2017) & (dmem_sel_ox2x)));
	assign g3960 = (((!g2015) & (!g2018) & (!sk[15]) & (dmem_sel_ox3x)) + ((!g2015) & (!g2018) & (sk[15]) & (dmem_sel_ox3x)) + ((!g2015) & (g2018) & (!sk[15]) & (!dmem_sel_ox3x)) + ((!g2015) & (g2018) & (!sk[15]) & (dmem_sel_ox3x)) + ((!g2015) & (g2018) & (sk[15]) & (dmem_sel_ox3x)) + ((g2015) & (!g2018) & (!sk[15]) & (dmem_sel_ox3x)) + ((g2015) & (g2018) & (!sk[15]) & (!dmem_sel_ox3x)) + ((g2015) & (g2018) & (!sk[15]) & (dmem_sel_ox3x)) + ((g2015) & (g2018) & (sk[15]) & (!dmem_sel_ox3x)) + ((g2015) & (g2018) & (sk[15]) & (dmem_sel_ox3x)));
	assign g3961 = (((!g2059) & (!g2058) & (!sk[16]) & (g76)) + ((!g2059) & (!g2058) & (sk[16]) & (g76)) + ((!g2059) & (g2058) & (!sk[16]) & (!g76)) + ((!g2059) & (g2058) & (!sk[16]) & (g76)) + ((!g2059) & (g2058) & (sk[16]) & (g76)) + ((g2059) & (!g2058) & (!sk[16]) & (g76)) + ((g2059) & (g2058) & (!sk[16]) & (!g76)) + ((g2059) & (g2058) & (!sk[16]) & (g76)) + ((g2059) & (g2058) & (sk[16]) & (!g76)) + ((g2059) & (g2058) & (sk[16]) & (g76)));
	assign g3962 = (((!sk[17]) & (!g2059) & (!g2063) & (g77)) + ((!sk[17]) & (!g2059) & (g2063) & (!g77)) + ((!sk[17]) & (!g2059) & (g2063) & (g77)) + ((!sk[17]) & (g2059) & (!g2063) & (g77)) + ((!sk[17]) & (g2059) & (g2063) & (!g77)) + ((!sk[17]) & (g2059) & (g2063) & (g77)) + ((sk[17]) & (!g2059) & (!g2063) & (g77)) + ((sk[17]) & (!g2059) & (g2063) & (g77)) + ((sk[17]) & (g2059) & (g2063) & (!g77)) + ((sk[17]) & (g2059) & (g2063) & (g77)));
	assign g3963 = (((!g2064) & (!dmem_dat_ix28x) & (!sk[18]) & (g78)) + ((!g2064) & (!dmem_dat_ix28x) & (sk[18]) & (g78)) + ((!g2064) & (dmem_dat_ix28x) & (!sk[18]) & (!g78)) + ((!g2064) & (dmem_dat_ix28x) & (!sk[18]) & (g78)) + ((!g2064) & (dmem_dat_ix28x) & (sk[18]) & (g78)) + ((g2064) & (!dmem_dat_ix28x) & (!sk[18]) & (g78)) + ((g2064) & (dmem_dat_ix28x) & (!sk[18]) & (!g78)) + ((g2064) & (dmem_dat_ix28x) & (!sk[18]) & (g78)) + ((g2064) & (dmem_dat_ix28x) & (sk[18]) & (!g78)) + ((g2064) & (dmem_dat_ix28x) & (sk[18]) & (g78)));
	assign g3964 = (((!g2064) & (!sk[19]) & (!dmem_dat_ix27x) & (g79)) + ((!g2064) & (!sk[19]) & (dmem_dat_ix27x) & (!g79)) + ((!g2064) & (!sk[19]) & (dmem_dat_ix27x) & (g79)) + ((!g2064) & (sk[19]) & (!dmem_dat_ix27x) & (g79)) + ((!g2064) & (sk[19]) & (dmem_dat_ix27x) & (g79)) + ((g2064) & (!sk[19]) & (!dmem_dat_ix27x) & (g79)) + ((g2064) & (!sk[19]) & (dmem_dat_ix27x) & (!g79)) + ((g2064) & (!sk[19]) & (dmem_dat_ix27x) & (g79)) + ((g2064) & (sk[19]) & (dmem_dat_ix27x) & (!g79)) + ((g2064) & (sk[19]) & (dmem_dat_ix27x) & (g79)));
	assign g3965 = (((!sk[20]) & (!g2064) & (!dmem_dat_ix31x) & (g80)) + ((!sk[20]) & (!g2064) & (dmem_dat_ix31x) & (!g80)) + ((!sk[20]) & (!g2064) & (dmem_dat_ix31x) & (g80)) + ((!sk[20]) & (g2064) & (!dmem_dat_ix31x) & (g80)) + ((!sk[20]) & (g2064) & (dmem_dat_ix31x) & (!g80)) + ((!sk[20]) & (g2064) & (dmem_dat_ix31x) & (g80)) + ((sk[20]) & (!g2064) & (!dmem_dat_ix31x) & (g80)) + ((sk[20]) & (!g2064) & (dmem_dat_ix31x) & (g80)) + ((sk[20]) & (g2064) & (dmem_dat_ix31x) & (!g80)) + ((sk[20]) & (g2064) & (dmem_dat_ix31x) & (g80)));
	assign g3966 = (((!g2064) & (!dmem_dat_ix30x) & (!sk[21]) & (g81)) + ((!g2064) & (!dmem_dat_ix30x) & (sk[21]) & (g81)) + ((!g2064) & (dmem_dat_ix30x) & (!sk[21]) & (!g81)) + ((!g2064) & (dmem_dat_ix30x) & (!sk[21]) & (g81)) + ((!g2064) & (dmem_dat_ix30x) & (sk[21]) & (g81)) + ((g2064) & (!dmem_dat_ix30x) & (!sk[21]) & (g81)) + ((g2064) & (dmem_dat_ix30x) & (!sk[21]) & (!g81)) + ((g2064) & (dmem_dat_ix30x) & (!sk[21]) & (g81)) + ((g2064) & (dmem_dat_ix30x) & (sk[21]) & (!g81)) + ((g2064) & (dmem_dat_ix30x) & (sk[21]) & (g81)));
	assign g3967 = (((!g2064) & (!dmem_dat_ix29x) & (!sk[22]) & (g82)) + ((!g2064) & (!dmem_dat_ix29x) & (sk[22]) & (g82)) + ((!g2064) & (dmem_dat_ix29x) & (!sk[22]) & (!g82)) + ((!g2064) & (dmem_dat_ix29x) & (!sk[22]) & (g82)) + ((!g2064) & (dmem_dat_ix29x) & (sk[22]) & (g82)) + ((g2064) & (!dmem_dat_ix29x) & (!sk[22]) & (g82)) + ((g2064) & (dmem_dat_ix29x) & (!sk[22]) & (!g82)) + ((g2064) & (dmem_dat_ix29x) & (!sk[22]) & (g82)) + ((g2064) & (dmem_dat_ix29x) & (sk[22]) & (!g82)) + ((g2064) & (dmem_dat_ix29x) & (sk[22]) & (g82)));
	assign g3968 = (((!g2064) & (!dmem_dat_ix26x) & (!sk[23]) & (g83)) + ((!g2064) & (!dmem_dat_ix26x) & (sk[23]) & (g83)) + ((!g2064) & (dmem_dat_ix26x) & (!sk[23]) & (!g83)) + ((!g2064) & (dmem_dat_ix26x) & (!sk[23]) & (g83)) + ((!g2064) & (dmem_dat_ix26x) & (sk[23]) & (g83)) + ((g2064) & (!dmem_dat_ix26x) & (!sk[23]) & (g83)) + ((g2064) & (dmem_dat_ix26x) & (!sk[23]) & (!g83)) + ((g2064) & (dmem_dat_ix26x) & (!sk[23]) & (g83)) + ((g2064) & (dmem_dat_ix26x) & (sk[23]) & (!g83)) + ((g2064) & (dmem_dat_ix26x) & (sk[23]) & (g83)));
	assign g84 = (((!g78) & (!g79) & (g80) & (g81) & (g82) & (!g83)));
	assign g3969 = (((!g2064) & (!dmem_dat_ix7x) & (!sk[25]) & (g85)) + ((!g2064) & (!dmem_dat_ix7x) & (sk[25]) & (g85)) + ((!g2064) & (dmem_dat_ix7x) & (!sk[25]) & (!g85)) + ((!g2064) & (dmem_dat_ix7x) & (!sk[25]) & (g85)) + ((!g2064) & (dmem_dat_ix7x) & (sk[25]) & (g85)) + ((g2064) & (!dmem_dat_ix7x) & (!sk[25]) & (g85)) + ((g2064) & (dmem_dat_ix7x) & (!sk[25]) & (!g85)) + ((g2064) & (dmem_dat_ix7x) & (!sk[25]) & (g85)) + ((g2064) & (dmem_dat_ix7x) & (sk[25]) & (!g85)) + ((g2064) & (dmem_dat_ix7x) & (sk[25]) & (g85)));
	assign g3970 = (((!g2064) & (!dmem_dat_ix6x) & (!sk[26]) & (g86)) + ((!g2064) & (!dmem_dat_ix6x) & (sk[26]) & (g86)) + ((!g2064) & (dmem_dat_ix6x) & (!sk[26]) & (!g86)) + ((!g2064) & (dmem_dat_ix6x) & (!sk[26]) & (g86)) + ((!g2064) & (dmem_dat_ix6x) & (sk[26]) & (g86)) + ((g2064) & (!dmem_dat_ix6x) & (!sk[26]) & (g86)) + ((g2064) & (dmem_dat_ix6x) & (!sk[26]) & (!g86)) + ((g2064) & (dmem_dat_ix6x) & (!sk[26]) & (g86)) + ((g2064) & (dmem_dat_ix6x) & (sk[26]) & (!g86)) + ((g2064) & (dmem_dat_ix6x) & (sk[26]) & (g86)));
	assign g3971 = (((!sk[27]) & (!g2064) & (!dmem_dat_ix2x) & (g87)) + ((!sk[27]) & (!g2064) & (dmem_dat_ix2x) & (!g87)) + ((!sk[27]) & (!g2064) & (dmem_dat_ix2x) & (g87)) + ((!sk[27]) & (g2064) & (!dmem_dat_ix2x) & (g87)) + ((!sk[27]) & (g2064) & (dmem_dat_ix2x) & (!g87)) + ((!sk[27]) & (g2064) & (dmem_dat_ix2x) & (g87)) + ((sk[27]) & (!g2064) & (!dmem_dat_ix2x) & (g87)) + ((sk[27]) & (!g2064) & (dmem_dat_ix2x) & (g87)) + ((sk[27]) & (g2064) & (dmem_dat_ix2x) & (!g87)) + ((sk[27]) & (g2064) & (dmem_dat_ix2x) & (g87)));
	assign g3972 = (((!g2064) & (!dmem_dat_ix1x) & (!sk[28]) & (g88)) + ((!g2064) & (!dmem_dat_ix1x) & (sk[28]) & (g88)) + ((!g2064) & (dmem_dat_ix1x) & (!sk[28]) & (!g88)) + ((!g2064) & (dmem_dat_ix1x) & (!sk[28]) & (g88)) + ((!g2064) & (dmem_dat_ix1x) & (sk[28]) & (g88)) + ((g2064) & (!dmem_dat_ix1x) & (!sk[28]) & (g88)) + ((g2064) & (dmem_dat_ix1x) & (!sk[28]) & (!g88)) + ((g2064) & (dmem_dat_ix1x) & (!sk[28]) & (g88)) + ((g2064) & (dmem_dat_ix1x) & (sk[28]) & (!g88)) + ((g2064) & (dmem_dat_ix1x) & (sk[28]) & (g88)));
	assign g3973 = (((!g2064) & (!sk[29]) & (!dmem_dat_ix0x) & (g89)) + ((!g2064) & (!sk[29]) & (dmem_dat_ix0x) & (!g89)) + ((!g2064) & (!sk[29]) & (dmem_dat_ix0x) & (g89)) + ((!g2064) & (sk[29]) & (!dmem_dat_ix0x) & (g89)) + ((!g2064) & (sk[29]) & (dmem_dat_ix0x) & (g89)) + ((g2064) & (!sk[29]) & (!dmem_dat_ix0x) & (g89)) + ((g2064) & (!sk[29]) & (dmem_dat_ix0x) & (!g89)) + ((g2064) & (!sk[29]) & (dmem_dat_ix0x) & (g89)) + ((g2064) & (sk[29]) & (dmem_dat_ix0x) & (!g89)) + ((g2064) & (sk[29]) & (dmem_dat_ix0x) & (g89)));
	assign g3974 = (((!sk[30]) & (!g2064) & (!dmem_dat_ix3x) & (g90)) + ((!sk[30]) & (!g2064) & (dmem_dat_ix3x) & (!g90)) + ((!sk[30]) & (!g2064) & (dmem_dat_ix3x) & (g90)) + ((!sk[30]) & (g2064) & (!dmem_dat_ix3x) & (g90)) + ((!sk[30]) & (g2064) & (dmem_dat_ix3x) & (!g90)) + ((!sk[30]) & (g2064) & (dmem_dat_ix3x) & (g90)) + ((sk[30]) & (!g2064) & (!dmem_dat_ix3x) & (g90)) + ((sk[30]) & (!g2064) & (dmem_dat_ix3x) & (g90)) + ((sk[30]) & (g2064) & (dmem_dat_ix3x) & (!g90)) + ((sk[30]) & (g2064) & (dmem_dat_ix3x) & (g90)));
	assign g3975 = (((!g2064) & (!dmem_dat_ix9x) & (!sk[31]) & (g91)) + ((!g2064) & (!dmem_dat_ix9x) & (sk[31]) & (g91)) + ((!g2064) & (dmem_dat_ix9x) & (!sk[31]) & (!g91)) + ((!g2064) & (dmem_dat_ix9x) & (!sk[31]) & (g91)) + ((!g2064) & (dmem_dat_ix9x) & (sk[31]) & (g91)) + ((g2064) & (!dmem_dat_ix9x) & (!sk[31]) & (g91)) + ((g2064) & (dmem_dat_ix9x) & (!sk[31]) & (!g91)) + ((g2064) & (dmem_dat_ix9x) & (!sk[31]) & (g91)) + ((g2064) & (dmem_dat_ix9x) & (sk[31]) & (!g91)) + ((g2064) & (dmem_dat_ix9x) & (sk[31]) & (g91)));
	assign g3976 = (((!sk[32]) & (!g2064) & (!dmem_dat_ix8x) & (g92)) + ((!sk[32]) & (!g2064) & (dmem_dat_ix8x) & (!g92)) + ((!sk[32]) & (!g2064) & (dmem_dat_ix8x) & (g92)) + ((!sk[32]) & (g2064) & (!dmem_dat_ix8x) & (g92)) + ((!sk[32]) & (g2064) & (dmem_dat_ix8x) & (!g92)) + ((!sk[32]) & (g2064) & (dmem_dat_ix8x) & (g92)) + ((sk[32]) & (!g2064) & (!dmem_dat_ix8x) & (g92)) + ((sk[32]) & (!g2064) & (dmem_dat_ix8x) & (g92)) + ((sk[32]) & (g2064) & (dmem_dat_ix8x) & (!g92)) + ((sk[32]) & (g2064) & (dmem_dat_ix8x) & (g92)));
	assign g93 = (((!g87) & (!g88) & (!g89) & (g90) & (!g91) & (!g92)));
	assign g94 = (((!g85) & (!g86) & (!sk[34]) & (!g84) & (g93)) + ((!g85) & (!g86) & (!sk[34]) & (g84) & (!g93)) + ((!g85) & (!g86) & (!sk[34]) & (g84) & (g93)) + ((!g85) & (g86) & (!sk[34]) & (!g84) & (!g93)) + ((!g85) & (g86) & (!sk[34]) & (!g84) & (g93)) + ((!g85) & (g86) & (!sk[34]) & (g84) & (!g93)) + ((!g85) & (g86) & (!sk[34]) & (g84) & (g93)) + ((!g85) & (g86) & (sk[34]) & (g84) & (g93)) + ((g85) & (!g86) & (!sk[34]) & (!g84) & (g93)) + ((g85) & (!g86) & (!sk[34]) & (g84) & (!g93)) + ((g85) & (!g86) & (!sk[34]) & (g84) & (g93)) + ((g85) & (g86) & (!sk[34]) & (!g84) & (!g93)) + ((g85) & (g86) & (!sk[34]) & (!g84) & (g93)) + ((g85) & (g86) & (!sk[34]) & (g84) & (!g93)) + ((g85) & (g86) & (!sk[34]) & (g84) & (g93)));
	assign g95 = (((!g85) & (!g86) & (!sk[35]) & (g93)) + ((!g85) & (!g86) & (sk[35]) & (g93)) + ((!g85) & (g86) & (!sk[35]) & (!g93)) + ((!g85) & (g86) & (!sk[35]) & (g93)) + ((g85) & (!g86) & (!sk[35]) & (g93)) + ((g85) & (g86) & (!sk[35]) & (!g93)) + ((g85) & (g86) & (!sk[35]) & (g93)));
	assign g96 = (((g85) & (!sk[36]) & (!g86)) + ((g85) & (!sk[36]) & (g86)) + ((g85) & (sk[36]) & (!g86)));
	assign g97 = (((!g85) & (!g86) & (g89) & (!g90) & (!g91) & (!g92)));
	assign g98 = (((!g87) & (sk[38]) & (g88)) + ((g87) & (!sk[38]) & (!g88)) + ((g87) & (!sk[38]) & (g88)));
	assign g99 = (((!g78) & (!g79) & (g80) & (!g81) & (g82) & (g83)));
	assign g100 = (((!g96) & (!g84) & (!g93) & (!g97) & (!g98) & (!g99)) + ((!g96) & (!g84) & (!g93) & (!g97) & (g98) & (!g99)) + ((!g96) & (!g84) & (!g93) & (g97) & (!g98) & (!g99)) + ((!g96) & (!g84) & (!g93) & (g97) & (g98) & (!g99)) + ((!g96) & (!g84) & (g93) & (!g97) & (!g98) & (!g99)) + ((!g96) & (!g84) & (g93) & (!g97) & (g98) & (!g99)) + ((!g96) & (!g84) & (g93) & (g97) & (!g98) & (!g99)) + ((!g96) & (!g84) & (g93) & (g97) & (g98) & (!g99)) + ((!g96) & (g84) & (!g93) & (!g97) & (!g98) & (!g99)) + ((!g96) & (g84) & (!g93) & (!g97) & (g98) & (!g99)) + ((!g96) & (g84) & (!g93) & (g97) & (!g98) & (!g99)) + ((!g96) & (g84) & (g93) & (!g97) & (!g98) & (!g99)) + ((!g96) & (g84) & (g93) & (!g97) & (g98) & (!g99)) + ((!g96) & (g84) & (g93) & (g97) & (!g98) & (!g99)) + ((g96) & (!g84) & (!g93) & (!g97) & (!g98) & (!g99)) + ((g96) & (!g84) & (!g93) & (!g97) & (g98) & (!g99)) + ((g96) & (!g84) & (!g93) & (g97) & (!g98) & (!g99)) + ((g96) & (!g84) & (!g93) & (g97) & (g98) & (!g99)) + ((g96) & (!g84) & (g93) & (!g97) & (!g98) & (!g99)) + ((g96) & (!g84) & (g93) & (!g97) & (g98) & (!g99)) + ((g96) & (!g84) & (g93) & (g97) & (!g98) & (!g99)) + ((g96) & (!g84) & (g93) & (g97) & (g98) & (!g99)) + ((g96) & (g84) & (!g93) & (!g97) & (!g98) & (!g99)) + ((g96) & (g84) & (!g93) & (!g97) & (g98) & (!g99)) + ((g96) & (g84) & (!g93) & (g97) & (!g98) & (!g99)));
	assign g101 = (((!sk[41]) & (!g84) & (!g88) & (g97)) + ((!sk[41]) & (!g84) & (g88) & (!g97)) + ((!sk[41]) & (!g84) & (g88) & (g97)) + ((!sk[41]) & (g84) & (!g88) & (g97)) + ((!sk[41]) & (g84) & (g88) & (!g97)) + ((!sk[41]) & (g84) & (g88) & (g97)) + ((sk[41]) & (g84) & (!g88) & (g97)));
	assign g102 = (((!g85) & (!g86) & (!g90) & (!g91) & (sk[42]) & (!g92)) + ((!g85) & (!g86) & (!g90) & (g91) & (!sk[42]) & (!g92)) + ((!g85) & (!g86) & (!g90) & (g91) & (!sk[42]) & (g92)) + ((!g85) & (!g86) & (g90) & (!g91) & (!sk[42]) & (!g92)) + ((!g85) & (!g86) & (g90) & (!g91) & (!sk[42]) & (g92)) + ((!g85) & (!g86) & (g90) & (g91) & (!sk[42]) & (!g92)) + ((!g85) & (!g86) & (g90) & (g91) & (!sk[42]) & (g92)) + ((!g85) & (g86) & (!g90) & (!g91) & (!sk[42]) & (!g92)) + ((!g85) & (g86) & (!g90) & (!g91) & (!sk[42]) & (g92)) + ((!g85) & (g86) & (!g90) & (g91) & (!sk[42]) & (!g92)) + ((!g85) & (g86) & (!g90) & (g91) & (!sk[42]) & (g92)) + ((!g85) & (g86) & (g90) & (!g91) & (!sk[42]) & (!g92)) + ((!g85) & (g86) & (g90) & (!g91) & (!sk[42]) & (g92)) + ((!g85) & (g86) & (g90) & (g91) & (!sk[42]) & (!g92)) + ((!g85) & (g86) & (g90) & (g91) & (!sk[42]) & (g92)) + ((g85) & (!g86) & (!g90) & (g91) & (!sk[42]) & (!g92)) + ((g85) & (!g86) & (!g90) & (g91) & (!sk[42]) & (g92)) + ((g85) & (!g86) & (g90) & (!g91) & (!sk[42]) & (!g92)) + ((g85) & (!g86) & (g90) & (!g91) & (!sk[42]) & (g92)) + ((g85) & (!g86) & (g90) & (g91) & (!sk[42]) & (!g92)) + ((g85) & (!g86) & (g90) & (g91) & (!sk[42]) & (g92)) + ((g85) & (g86) & (!g90) & (!g91) & (!sk[42]) & (!g92)) + ((g85) & (g86) & (!g90) & (!g91) & (!sk[42]) & (g92)) + ((g85) & (g86) & (!g90) & (g91) & (!sk[42]) & (!g92)) + ((g85) & (g86) & (!g90) & (g91) & (!sk[42]) & (g92)) + ((g85) & (g86) & (g90) & (!g91) & (!sk[42]) & (!g92)) + ((g85) & (g86) & (g90) & (!g91) & (!sk[42]) & (g92)) + ((g85) & (g86) & (g90) & (g91) & (!sk[42]) & (!g92)) + ((g85) & (g86) & (g90) & (g91) & (!sk[42]) & (g92)));
	assign g103 = (((!g84) & (!sk[43]) & (!g88) & (!g89) & (g102)) + ((!g84) & (!sk[43]) & (!g88) & (g89) & (!g102)) + ((!g84) & (!sk[43]) & (!g88) & (g89) & (g102)) + ((!g84) & (!sk[43]) & (g88) & (!g89) & (!g102)) + ((!g84) & (!sk[43]) & (g88) & (!g89) & (g102)) + ((!g84) & (!sk[43]) & (g88) & (g89) & (!g102)) + ((!g84) & (!sk[43]) & (g88) & (g89) & (g102)) + ((g84) & (!sk[43]) & (!g88) & (!g89) & (g102)) + ((g84) & (!sk[43]) & (!g88) & (g89) & (!g102)) + ((g84) & (!sk[43]) & (!g88) & (g89) & (g102)) + ((g84) & (!sk[43]) & (g88) & (!g89) & (!g102)) + ((g84) & (!sk[43]) & (g88) & (!g89) & (g102)) + ((g84) & (!sk[43]) & (g88) & (g89) & (!g102)) + ((g84) & (!sk[43]) & (g88) & (g89) & (g102)) + ((g84) & (sk[43]) & (!g88) & (!g89) & (g102)));
	assign g104 = (((!g84) & (!g94) & (!g95) & (g100) & (!g101) & (!g103)) + ((!g84) & (!g94) & (g95) & (g100) & (!g101) & (!g103)) + ((g84) & (!g94) & (!g95) & (g100) & (!g101) & (!g103)));
	assign g105 = (((!g78) & (!sk[45]) & (!g79) & (!g80) & (g81) & (!g82)) + ((!g78) & (!sk[45]) & (!g79) & (!g80) & (g81) & (g82)) + ((!g78) & (!sk[45]) & (!g79) & (g80) & (!g81) & (!g82)) + ((!g78) & (!sk[45]) & (!g79) & (g80) & (!g81) & (g82)) + ((!g78) & (!sk[45]) & (!g79) & (g80) & (g81) & (!g82)) + ((!g78) & (!sk[45]) & (!g79) & (g80) & (g81) & (g82)) + ((!g78) & (!sk[45]) & (g79) & (!g80) & (!g81) & (!g82)) + ((!g78) & (!sk[45]) & (g79) & (!g80) & (!g81) & (g82)) + ((!g78) & (!sk[45]) & (g79) & (!g80) & (g81) & (!g82)) + ((!g78) & (!sk[45]) & (g79) & (!g80) & (g81) & (g82)) + ((!g78) & (!sk[45]) & (g79) & (g80) & (!g81) & (!g82)) + ((!g78) & (!sk[45]) & (g79) & (g80) & (!g81) & (g82)) + ((!g78) & (!sk[45]) & (g79) & (g80) & (g81) & (!g82)) + ((!g78) & (!sk[45]) & (g79) & (g80) & (g81) & (g82)) + ((g78) & (!sk[45]) & (!g79) & (!g80) & (g81) & (!g82)) + ((g78) & (!sk[45]) & (!g79) & (!g80) & (g81) & (g82)) + ((g78) & (!sk[45]) & (!g79) & (g80) & (!g81) & (!g82)) + ((g78) & (!sk[45]) & (!g79) & (g80) & (!g81) & (g82)) + ((g78) & (!sk[45]) & (!g79) & (g80) & (g81) & (!g82)) + ((g78) & (!sk[45]) & (!g79) & (g80) & (g81) & (g82)) + ((g78) & (!sk[45]) & (g79) & (!g80) & (!g81) & (!g82)) + ((g78) & (!sk[45]) & (g79) & (!g80) & (!g81) & (g82)) + ((g78) & (!sk[45]) & (g79) & (!g80) & (g81) & (!g82)) + ((g78) & (!sk[45]) & (g79) & (!g80) & (g81) & (g82)) + ((g78) & (!sk[45]) & (g79) & (g80) & (!g81) & (!g82)) + ((g78) & (!sk[45]) & (g79) & (g80) & (!g81) & (g82)) + ((g78) & (!sk[45]) & (g79) & (g80) & (g81) & (!g82)) + ((g78) & (!sk[45]) & (g79) & (g80) & (g81) & (g82)) + ((g78) & (sk[45]) & (!g79) & (!g80) & (!g81) & (!g82)));
	assign g106 = (((!g78) & (!g79) & (g80) & (g81) & (g82) & (g83)) + ((g78) & (g79) & (g80) & (!g81) & (g82) & (g83)));
	assign g3977 = (((!sk[47]) & (!g2064) & (!dmem_dat_ix25x) & (g107)) + ((!sk[47]) & (!g2064) & (dmem_dat_ix25x) & (!g107)) + ((!sk[47]) & (!g2064) & (dmem_dat_ix25x) & (g107)) + ((!sk[47]) & (g2064) & (!dmem_dat_ix25x) & (g107)) + ((!sk[47]) & (g2064) & (dmem_dat_ix25x) & (!g107)) + ((!sk[47]) & (g2064) & (dmem_dat_ix25x) & (g107)) + ((sk[47]) & (!g2064) & (!dmem_dat_ix25x) & (g107)) + ((sk[47]) & (!g2064) & (dmem_dat_ix25x) & (g107)) + ((sk[47]) & (g2064) & (dmem_dat_ix25x) & (!g107)) + ((sk[47]) & (g2064) & (dmem_dat_ix25x) & (g107)));
	assign g3978 = (((!sk[48]) & (!g2064) & (!dmem_dat_ix23x) & (g108)) + ((!sk[48]) & (!g2064) & (dmem_dat_ix23x) & (!g108)) + ((!sk[48]) & (!g2064) & (dmem_dat_ix23x) & (g108)) + ((!sk[48]) & (g2064) & (!dmem_dat_ix23x) & (g108)) + ((!sk[48]) & (g2064) & (dmem_dat_ix23x) & (!g108)) + ((!sk[48]) & (g2064) & (dmem_dat_ix23x) & (g108)) + ((sk[48]) & (!g2064) & (!dmem_dat_ix23x) & (g108)) + ((sk[48]) & (!g2064) & (dmem_dat_ix23x) & (g108)) + ((sk[48]) & (g2064) & (dmem_dat_ix23x) & (!g108)) + ((sk[48]) & (g2064) & (dmem_dat_ix23x) & (g108)));
	assign g3979 = (((!sk[49]) & (!g2064) & (!dmem_dat_ix22x) & (g109)) + ((!sk[49]) & (!g2064) & (dmem_dat_ix22x) & (!g109)) + ((!sk[49]) & (!g2064) & (dmem_dat_ix22x) & (g109)) + ((!sk[49]) & (g2064) & (!dmem_dat_ix22x) & (g109)) + ((!sk[49]) & (g2064) & (dmem_dat_ix22x) & (!g109)) + ((!sk[49]) & (g2064) & (dmem_dat_ix22x) & (g109)) + ((sk[49]) & (!g2064) & (!dmem_dat_ix22x) & (g109)) + ((sk[49]) & (!g2064) & (dmem_dat_ix22x) & (g109)) + ((sk[49]) & (g2064) & (dmem_dat_ix22x) & (!g109)) + ((sk[49]) & (g2064) & (dmem_dat_ix22x) & (g109)));
	assign g3980 = (((!sk[50]) & (!g2064) & (!dmem_dat_ix24x) & (g110)) + ((!sk[50]) & (!g2064) & (dmem_dat_ix24x) & (!g110)) + ((!sk[50]) & (!g2064) & (dmem_dat_ix24x) & (g110)) + ((!sk[50]) & (g2064) & (!dmem_dat_ix24x) & (g110)) + ((!sk[50]) & (g2064) & (dmem_dat_ix24x) & (!g110)) + ((!sk[50]) & (g2064) & (dmem_dat_ix24x) & (g110)) + ((sk[50]) & (!g2064) & (!dmem_dat_ix24x) & (g110)) + ((sk[50]) & (!g2064) & (dmem_dat_ix24x) & (g110)) + ((sk[50]) & (g2064) & (dmem_dat_ix24x) & (!g110)) + ((sk[50]) & (g2064) & (dmem_dat_ix24x) & (g110)));
	assign g111 = (((g80) & (g82) & (!g107) & (!g108) & (!g109) & (!g110)) + ((g80) & (g82) & (!g107) & (!g108) & (g109) & (!g110)) + ((g80) & (g82) & (!g107) & (!g108) & (g109) & (g110)) + ((g80) & (g82) & (!g107) & (g108) & (!g109) & (!g110)) + ((g80) & (g82) & (!g107) & (g108) & (!g109) & (g110)));
	assign g112 = (((!g83) & (!g105) & (!g106) & (!sk[52]) & (g111)) + ((!g83) & (!g105) & (g106) & (!sk[52]) & (!g111)) + ((!g83) & (!g105) & (g106) & (!sk[52]) & (g111)) + ((!g83) & (g105) & (!g106) & (!sk[52]) & (!g111)) + ((!g83) & (g105) & (!g106) & (!sk[52]) & (g111)) + ((!g83) & (g105) & (g106) & (!sk[52]) & (!g111)) + ((!g83) & (g105) & (g106) & (!sk[52]) & (g111)) + ((g83) & (!g105) & (!g106) & (!sk[52]) & (g111)) + ((g83) & (!g105) & (g106) & (!sk[52]) & (!g111)) + ((g83) & (!g105) & (g106) & (!sk[52]) & (g111)) + ((g83) & (!g105) & (g106) & (sk[52]) & (g111)) + ((g83) & (g105) & (!g106) & (!sk[52]) & (!g111)) + ((g83) & (g105) & (!g106) & (!sk[52]) & (g111)) + ((g83) & (g105) & (!g106) & (sk[52]) & (!g111)) + ((g83) & (g105) & (!g106) & (sk[52]) & (g111)) + ((g83) & (g105) & (g106) & (!sk[52]) & (!g111)) + ((g83) & (g105) & (g106) & (!sk[52]) & (g111)) + ((g83) & (g105) & (g106) & (sk[52]) & (!g111)) + ((g83) & (g105) & (g106) & (sk[52]) & (g111)));
	assign g113 = (((!sk[53]) & (!g84) & (!g89) & (!g102) & (g98)) + ((!sk[53]) & (!g84) & (!g89) & (g102) & (!g98)) + ((!sk[53]) & (!g84) & (!g89) & (g102) & (g98)) + ((!sk[53]) & (!g84) & (g89) & (!g102) & (!g98)) + ((!sk[53]) & (!g84) & (g89) & (!g102) & (g98)) + ((!sk[53]) & (!g84) & (g89) & (g102) & (!g98)) + ((!sk[53]) & (!g84) & (g89) & (g102) & (g98)) + ((!sk[53]) & (g84) & (!g89) & (!g102) & (g98)) + ((!sk[53]) & (g84) & (!g89) & (g102) & (!g98)) + ((!sk[53]) & (g84) & (!g89) & (g102) & (g98)) + ((!sk[53]) & (g84) & (g89) & (!g102) & (!g98)) + ((!sk[53]) & (g84) & (g89) & (!g102) & (g98)) + ((!sk[53]) & (g84) & (g89) & (g102) & (!g98)) + ((!sk[53]) & (g84) & (g89) & (g102) & (g98)) + ((sk[53]) & (g84) & (!g89) & (g102) & (g98)));
	assign g114 = (((!sk[54]) & (!g78) & (!g79) & (!g80) & (g81)) + ((!sk[54]) & (!g78) & (!g79) & (g80) & (!g81)) + ((!sk[54]) & (!g78) & (!g79) & (g80) & (g81)) + ((!sk[54]) & (!g78) & (g79) & (!g80) & (!g81)) + ((!sk[54]) & (!g78) & (g79) & (!g80) & (g81)) + ((!sk[54]) & (!g78) & (g79) & (g80) & (!g81)) + ((!sk[54]) & (!g78) & (g79) & (g80) & (g81)) + ((!sk[54]) & (g78) & (!g79) & (!g80) & (g81)) + ((!sk[54]) & (g78) & (!g79) & (g80) & (!g81)) + ((!sk[54]) & (g78) & (!g79) & (g80) & (g81)) + ((!sk[54]) & (g78) & (g79) & (!g80) & (!g81)) + ((!sk[54]) & (g78) & (g79) & (!g80) & (g81)) + ((!sk[54]) & (g78) & (g79) & (g80) & (!g81)) + ((!sk[54]) & (g78) & (g79) & (g80) & (g81)) + ((sk[54]) & (!g78) & (!g79) & (!g80) & (!g81)));
	assign g115 = (((!g82) & (!g83) & (!sk[55]) & (g107)) + ((!g82) & (g83) & (!sk[55]) & (!g107)) + ((!g82) & (g83) & (!sk[55]) & (g107)) + ((g82) & (!g83) & (!sk[55]) & (g107)) + ((g82) & (!g83) & (sk[55]) & (!g107)) + ((g82) & (g83) & (!sk[55]) & (!g107)) + ((g82) & (g83) & (!sk[55]) & (g107)));
	assign g116 = (((!g78) & (!g79) & (!g80) & (!g81) & (!g82) & (!g83)) + ((!g78) & (!g79) & (!g80) & (!g81) & (g82) & (g83)) + ((!g78) & (!g79) & (!g80) & (g81) & (!g82) & (g83)));
	assign g117 = (((!sk[57]) & (!g114) & (!g115) & (g116)) + ((!sk[57]) & (!g114) & (g115) & (!g116)) + ((!sk[57]) & (!g114) & (g115) & (g116)) + ((!sk[57]) & (g114) & (!g115) & (g116)) + ((!sk[57]) & (g114) & (g115) & (!g116)) + ((!sk[57]) & (g114) & (g115) & (g116)) + ((sk[57]) & (!g114) & (!g115) & (!g116)) + ((sk[57]) & (!g114) & (g115) & (!g116)) + ((sk[57]) & (g114) & (!g115) & (!g116)));
	assign g118 = (((g78) & (g79) & (g80) & (!g81) & (g82) & (!g83)));
	assign g119 = (((!g78) & (!g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((!g78) & (g79) & (!g80) & (g81) & (!g82) & (!g83)) + ((!g78) & (g79) & (g80) & (!g81) & (g82) & (!g83)) + ((g78) & (!g79) & (g80) & (!g81) & (g82) & (g83)) + ((g78) & (g79) & (!g80) & (!g81) & (!g82) & (!g83)));
	assign g120 = (((!g78) & (!g79) & (g80) & (!g81) & (!g82) & (g83)) + ((!g78) & (!g79) & (g80) & (g81) & (!g82) & (!g83)) + ((!g78) & (g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((!g78) & (g79) & (g80) & (!g81) & (!g82) & (!g83)) + ((!g78) & (g79) & (g80) & (!g81) & (!g82) & (g83)) + ((!g78) & (g79) & (g80) & (!g81) & (g82) & (g83)) + ((g78) & (!g79) & (!g80) & (!g81) & (!g82) & (!g83)) + ((g78) & (!g79) & (g80) & (!g81) & (!g82) & (!g83)) + ((g78) & (!g79) & (g80) & (!g81) & (!g82) & (g83)) + ((g78) & (!g79) & (g80) & (g81) & (!g82) & (g83)) + ((g78) & (g79) & (g80) & (!g81) & (!g82) & (!g83)) + ((g78) & (g79) & (g80) & (!g81) & (!g82) & (g83)) + ((g78) & (g79) & (g80) & (g81) & (!g82) & (!g83)) + ((g78) & (g79) & (g80) & (g81) & (!g82) & (g83)));
	assign g121 = (((!g118) & (!g85) & (!sk[61]) & (!g86) & (g119) & (!g120)) + ((!g118) & (!g85) & (!sk[61]) & (!g86) & (g119) & (g120)) + ((!g118) & (!g85) & (!sk[61]) & (g86) & (!g119) & (!g120)) + ((!g118) & (!g85) & (!sk[61]) & (g86) & (!g119) & (g120)) + ((!g118) & (!g85) & (!sk[61]) & (g86) & (g119) & (!g120)) + ((!g118) & (!g85) & (!sk[61]) & (g86) & (g119) & (g120)) + ((!g118) & (!g85) & (sk[61]) & (!g86) & (!g119) & (!g120)) + ((!g118) & (!g85) & (sk[61]) & (g86) & (!g119) & (!g120)) + ((!g118) & (g85) & (!sk[61]) & (!g86) & (!g119) & (!g120)) + ((!g118) & (g85) & (!sk[61]) & (!g86) & (!g119) & (g120)) + ((!g118) & (g85) & (!sk[61]) & (!g86) & (g119) & (!g120)) + ((!g118) & (g85) & (!sk[61]) & (!g86) & (g119) & (g120)) + ((!g118) & (g85) & (!sk[61]) & (g86) & (!g119) & (!g120)) + ((!g118) & (g85) & (!sk[61]) & (g86) & (!g119) & (g120)) + ((!g118) & (g85) & (!sk[61]) & (g86) & (g119) & (!g120)) + ((!g118) & (g85) & (!sk[61]) & (g86) & (g119) & (g120)) + ((!g118) & (g85) & (sk[61]) & (!g86) & (!g119) & (!g120)) + ((!g118) & (g85) & (sk[61]) & (g86) & (!g119) & (!g120)) + ((g118) & (!g85) & (!sk[61]) & (!g86) & (g119) & (!g120)) + ((g118) & (!g85) & (!sk[61]) & (!g86) & (g119) & (g120)) + ((g118) & (!g85) & (!sk[61]) & (g86) & (!g119) & (!g120)) + ((g118) & (!g85) & (!sk[61]) & (g86) & (!g119) & (g120)) + ((g118) & (!g85) & (!sk[61]) & (g86) & (g119) & (!g120)) + ((g118) & (!g85) & (!sk[61]) & (g86) & (g119) & (g120)) + ((g118) & (g85) & (!sk[61]) & (!g86) & (!g119) & (!g120)) + ((g118) & (g85) & (!sk[61]) & (!g86) & (!g119) & (g120)) + ((g118) & (g85) & (!sk[61]) & (!g86) & (g119) & (!g120)) + ((g118) & (g85) & (!sk[61]) & (!g86) & (g119) & (g120)) + ((g118) & (g85) & (!sk[61]) & (g86) & (!g119) & (!g120)) + ((g118) & (g85) & (!sk[61]) & (g86) & (!g119) & (g120)) + ((g118) & (g85) & (!sk[61]) & (g86) & (g119) & (!g120)) + ((g118) & (g85) & (!sk[61]) & (g86) & (g119) & (g120)) + ((g118) & (g85) & (sk[61]) & (g86) & (!g119) & (!g120)));
	assign g122 = (((!g112) & (!g113) & (!g117) & (!sk[62]) & (g121)) + ((!g112) & (!g113) & (g117) & (!sk[62]) & (!g121)) + ((!g112) & (!g113) & (g117) & (!sk[62]) & (g121)) + ((!g112) & (!g113) & (g117) & (sk[62]) & (g121)) + ((!g112) & (g113) & (!g117) & (!sk[62]) & (!g121)) + ((!g112) & (g113) & (!g117) & (!sk[62]) & (g121)) + ((!g112) & (g113) & (g117) & (!sk[62]) & (!g121)) + ((!g112) & (g113) & (g117) & (!sk[62]) & (g121)) + ((g112) & (!g113) & (!g117) & (!sk[62]) & (g121)) + ((g112) & (!g113) & (g117) & (!sk[62]) & (!g121)) + ((g112) & (!g113) & (g117) & (!sk[62]) & (g121)) + ((g112) & (g113) & (!g117) & (!sk[62]) & (!g121)) + ((g112) & (g113) & (!g117) & (!sk[62]) & (g121)) + ((g112) & (g113) & (g117) & (!sk[62]) & (!g121)) + ((g112) & (g113) & (g117) & (!sk[62]) & (g121)));
	assign g123 = (((!g76) & (!g77) & (!sk[63]) & (!g104) & (g122)) + ((!g76) & (!g77) & (!sk[63]) & (g104) & (!g122)) + ((!g76) & (!g77) & (!sk[63]) & (g104) & (g122)) + ((!g76) & (!g77) & (sk[63]) & (g104) & (g122)) + ((!g76) & (g77) & (!sk[63]) & (!g104) & (!g122)) + ((!g76) & (g77) & (!sk[63]) & (!g104) & (g122)) + ((!g76) & (g77) & (!sk[63]) & (g104) & (!g122)) + ((!g76) & (g77) & (!sk[63]) & (g104) & (g122)) + ((!g76) & (g77) & (sk[63]) & (!g104) & (!g122)) + ((!g76) & (g77) & (sk[63]) & (!g104) & (g122)) + ((!g76) & (g77) & (sk[63]) & (g104) & (!g122)) + ((!g76) & (g77) & (sk[63]) & (g104) & (g122)) + ((g76) & (!g77) & (!sk[63]) & (!g104) & (g122)) + ((g76) & (!g77) & (!sk[63]) & (g104) & (!g122)) + ((g76) & (!g77) & (!sk[63]) & (g104) & (g122)) + ((g76) & (!g77) & (sk[63]) & (!g104) & (!g122)) + ((g76) & (!g77) & (sk[63]) & (!g104) & (g122)) + ((g76) & (!g77) & (sk[63]) & (g104) & (!g122)) + ((g76) & (!g77) & (sk[63]) & (g104) & (g122)) + ((g76) & (g77) & (!sk[63]) & (!g104) & (!g122)) + ((g76) & (g77) & (!sk[63]) & (!g104) & (g122)) + ((g76) & (g77) & (!sk[63]) & (g104) & (!g122)) + ((g76) & (g77) & (!sk[63]) & (g104) & (g122)) + ((g76) & (g77) & (sk[63]) & (!g104) & (!g122)) + ((g76) & (g77) & (sk[63]) & (!g104) & (g122)) + ((g76) & (g77) & (sk[63]) & (g104) & (!g122)) + ((g76) & (g77) & (sk[63]) & (g104) & (g122)));
	assign g124 = (((!g1) & (!sk[64]) & (!g74) & (!dmem_ack_i) & (g75) & (!g123)) + ((!g1) & (!sk[64]) & (!g74) & (!dmem_ack_i) & (g75) & (g123)) + ((!g1) & (!sk[64]) & (!g74) & (dmem_ack_i) & (!g75) & (!g123)) + ((!g1) & (!sk[64]) & (!g74) & (dmem_ack_i) & (!g75) & (g123)) + ((!g1) & (!sk[64]) & (!g74) & (dmem_ack_i) & (g75) & (!g123)) + ((!g1) & (!sk[64]) & (!g74) & (dmem_ack_i) & (g75) & (g123)) + ((!g1) & (!sk[64]) & (g74) & (!dmem_ack_i) & (!g75) & (!g123)) + ((!g1) & (!sk[64]) & (g74) & (!dmem_ack_i) & (!g75) & (g123)) + ((!g1) & (!sk[64]) & (g74) & (!dmem_ack_i) & (g75) & (!g123)) + ((!g1) & (!sk[64]) & (g74) & (!dmem_ack_i) & (g75) & (g123)) + ((!g1) & (!sk[64]) & (g74) & (dmem_ack_i) & (!g75) & (!g123)) + ((!g1) & (!sk[64]) & (g74) & (dmem_ack_i) & (!g75) & (g123)) + ((!g1) & (!sk[64]) & (g74) & (dmem_ack_i) & (g75) & (!g123)) + ((!g1) & (!sk[64]) & (g74) & (dmem_ack_i) & (g75) & (g123)) + ((!g1) & (sk[64]) & (!g74) & (dmem_ack_i) & (g75) & (g123)) + ((!g1) & (sk[64]) & (g74) & (!dmem_ack_i) & (!g75) & (g123)) + ((!g1) & (sk[64]) & (g74) & (!dmem_ack_i) & (g75) & (g123)) + ((!g1) & (sk[64]) & (g74) & (dmem_ack_i) & (!g75) & (g123)) + ((!g1) & (sk[64]) & (g74) & (dmem_ack_i) & (g75) & (g123)) + ((g1) & (!sk[64]) & (!g74) & (!dmem_ack_i) & (g75) & (!g123)) + ((g1) & (!sk[64]) & (!g74) & (!dmem_ack_i) & (g75) & (g123)) + ((g1) & (!sk[64]) & (!g74) & (dmem_ack_i) & (!g75) & (!g123)) + ((g1) & (!sk[64]) & (!g74) & (dmem_ack_i) & (!g75) & (g123)) + ((g1) & (!sk[64]) & (!g74) & (dmem_ack_i) & (g75) & (!g123)) + ((g1) & (!sk[64]) & (!g74) & (dmem_ack_i) & (g75) & (g123)) + ((g1) & (!sk[64]) & (g74) & (!dmem_ack_i) & (!g75) & (!g123)) + ((g1) & (!sk[64]) & (g74) & (!dmem_ack_i) & (!g75) & (g123)) + ((g1) & (!sk[64]) & (g74) & (!dmem_ack_i) & (g75) & (!g123)) + ((g1) & (!sk[64]) & (g74) & (!dmem_ack_i) & (g75) & (g123)) + ((g1) & (!sk[64]) & (g74) & (dmem_ack_i) & (!g75) & (!g123)) + ((g1) & (!sk[64]) & (g74) & (dmem_ack_i) & (!g75) & (g123)) + ((g1) & (!sk[64]) & (g74) & (dmem_ack_i) & (g75) & (!g123)) + ((g1) & (!sk[64]) & (g74) & (dmem_ack_i) & (g75) & (g123)) + ((g1) & (sk[64]) & (!g74) & (!dmem_ack_i) & (!g75) & (!g123)) + ((g1) & (sk[64]) & (!g74) & (!dmem_ack_i) & (!g75) & (g123)) + ((g1) & (sk[64]) & (!g74) & (!dmem_ack_i) & (g75) & (!g123)) + ((g1) & (sk[64]) & (!g74) & (!dmem_ack_i) & (g75) & (g123)) + ((g1) & (sk[64]) & (!g74) & (dmem_ack_i) & (!g75) & (!g123)) + ((g1) & (sk[64]) & (!g74) & (dmem_ack_i) & (!g75) & (g123)) + ((g1) & (sk[64]) & (!g74) & (dmem_ack_i) & (g75) & (!g123)) + ((g1) & (sk[64]) & (!g74) & (dmem_ack_i) & (g75) & (g123)) + ((g1) & (sk[64]) & (g74) & (!dmem_ack_i) & (!g75) & (!g123)) + ((g1) & (sk[64]) & (g74) & (!dmem_ack_i) & (!g75) & (g123)) + ((g1) & (sk[64]) & (g74) & (!dmem_ack_i) & (g75) & (!g123)) + ((g1) & (sk[64]) & (g74) & (!dmem_ack_i) & (g75) & (g123)) + ((g1) & (sk[64]) & (g74) & (dmem_ack_i) & (!g75) & (!g123)) + ((g1) & (sk[64]) & (g74) & (dmem_ack_i) & (!g75) & (g123)) + ((g1) & (sk[64]) & (g74) & (dmem_ack_i) & (g75) & (!g123)) + ((g1) & (sk[64]) & (g74) & (dmem_ack_i) & (g75) & (g123)));
	assign g125 = (((!g110) & (!sk[65]) & (!g114) & (g115)) + ((!g110) & (!sk[65]) & (g114) & (!g115)) + ((!g110) & (!sk[65]) & (g114) & (g115)) + ((g110) & (!sk[65]) & (!g114) & (g115)) + ((g110) & (!sk[65]) & (g114) & (!g115)) + ((g110) & (!sk[65]) & (g114) & (g115)) + ((g110) & (sk[65]) & (g114) & (g115)));
	assign g127 = (((g77) & (!sk[66]) & (!g126)) + ((g77) & (!sk[66]) & (g126)) + ((g77) & (sk[66]) & (!g126)));
	assign g130 = (((!sk[67]) & (!g74) & (!g75) & (!g128) & (g129)) + ((!sk[67]) & (!g74) & (!g75) & (g128) & (!g129)) + ((!sk[67]) & (!g74) & (!g75) & (g128) & (g129)) + ((!sk[67]) & (!g74) & (g75) & (!g128) & (!g129)) + ((!sk[67]) & (!g74) & (g75) & (!g128) & (g129)) + ((!sk[67]) & (!g74) & (g75) & (g128) & (!g129)) + ((!sk[67]) & (!g74) & (g75) & (g128) & (g129)) + ((!sk[67]) & (g74) & (!g75) & (!g128) & (g129)) + ((!sk[67]) & (g74) & (!g75) & (g128) & (!g129)) + ((!sk[67]) & (g74) & (!g75) & (g128) & (g129)) + ((!sk[67]) & (g74) & (g75) & (!g128) & (!g129)) + ((!sk[67]) & (g74) & (g75) & (!g128) & (g129)) + ((!sk[67]) & (g74) & (g75) & (g128) & (!g129)) + ((!sk[67]) & (g74) & (g75) & (g128) & (g129)) + ((sk[67]) & (!g74) & (!g75) & (g128) & (!g129)));
	assign g131 = (((!g78) & (!g82) & (!sk[68]) & (g83)) + ((!g78) & (g82) & (!sk[68]) & (!g83)) + ((!g78) & (g82) & (!sk[68]) & (g83)) + ((g78) & (!g82) & (!sk[68]) & (g83)) + ((g78) & (!g82) & (sk[68]) & (g83)) + ((g78) & (g82) & (!sk[68]) & (!g83)) + ((g78) & (g82) & (!sk[68]) & (g83)));
	assign g132 = (((!g79) & (!sk[69]) & (!g80) & (!g81) & (g131)) + ((!g79) & (!sk[69]) & (!g80) & (g81) & (!g131)) + ((!g79) & (!sk[69]) & (!g80) & (g81) & (g131)) + ((!g79) & (!sk[69]) & (g80) & (!g81) & (!g131)) + ((!g79) & (!sk[69]) & (g80) & (!g81) & (g131)) + ((!g79) & (!sk[69]) & (g80) & (g81) & (!g131)) + ((!g79) & (!sk[69]) & (g80) & (g81) & (g131)) + ((!g79) & (sk[69]) & (g80) & (g81) & (g131)) + ((g79) & (!sk[69]) & (!g80) & (!g81) & (g131)) + ((g79) & (!sk[69]) & (!g80) & (g81) & (!g131)) + ((g79) & (!sk[69]) & (!g80) & (g81) & (g131)) + ((g79) & (!sk[69]) & (g80) & (!g81) & (!g131)) + ((g79) & (!sk[69]) & (g80) & (!g81) & (g131)) + ((g79) & (!sk[69]) & (g80) & (g81) & (!g131)) + ((g79) & (!sk[69]) & (g80) & (g81) & (g131)));
	assign g133 = (((!g78) & (!sk[70]) & (!g82) & (g83)) + ((!g78) & (!sk[70]) & (g82) & (!g83)) + ((!g78) & (!sk[70]) & (g82) & (g83)) + ((g78) & (!sk[70]) & (!g82) & (g83)) + ((g78) & (!sk[70]) & (g82) & (!g83)) + ((g78) & (!sk[70]) & (g82) & (g83)) + ((g78) & (sk[70]) & (!g82) & (!g83)));
	assign g134 = (((!g79) & (!g80) & (!sk[71]) & (!g81) & (g131) & (!g133)) + ((!g79) & (!g80) & (!sk[71]) & (!g81) & (g131) & (g133)) + ((!g79) & (!g80) & (!sk[71]) & (g81) & (!g131) & (!g133)) + ((!g79) & (!g80) & (!sk[71]) & (g81) & (!g131) & (g133)) + ((!g79) & (!g80) & (!sk[71]) & (g81) & (g131) & (!g133)) + ((!g79) & (!g80) & (!sk[71]) & (g81) & (g131) & (g133)) + ((!g79) & (g80) & (!sk[71]) & (!g81) & (!g131) & (!g133)) + ((!g79) & (g80) & (!sk[71]) & (!g81) & (!g131) & (g133)) + ((!g79) & (g80) & (!sk[71]) & (!g81) & (g131) & (!g133)) + ((!g79) & (g80) & (!sk[71]) & (!g81) & (g131) & (g133)) + ((!g79) & (g80) & (!sk[71]) & (g81) & (!g131) & (!g133)) + ((!g79) & (g80) & (!sk[71]) & (g81) & (!g131) & (g133)) + ((!g79) & (g80) & (!sk[71]) & (g81) & (g131) & (!g133)) + ((!g79) & (g80) & (!sk[71]) & (g81) & (g131) & (g133)) + ((g79) & (!g80) & (!sk[71]) & (!g81) & (g131) & (!g133)) + ((g79) & (!g80) & (!sk[71]) & (!g81) & (g131) & (g133)) + ((g79) & (!g80) & (!sk[71]) & (g81) & (!g131) & (!g133)) + ((g79) & (!g80) & (!sk[71]) & (g81) & (!g131) & (g133)) + ((g79) & (!g80) & (!sk[71]) & (g81) & (g131) & (!g133)) + ((g79) & (!g80) & (!sk[71]) & (g81) & (g131) & (g133)) + ((g79) & (g80) & (!sk[71]) & (!g81) & (!g131) & (!g133)) + ((g79) & (g80) & (!sk[71]) & (!g81) & (!g131) & (g133)) + ((g79) & (g80) & (!sk[71]) & (!g81) & (g131) & (!g133)) + ((g79) & (g80) & (!sk[71]) & (!g81) & (g131) & (g133)) + ((g79) & (g80) & (!sk[71]) & (g81) & (!g131) & (!g133)) + ((g79) & (g80) & (!sk[71]) & (g81) & (!g131) & (g133)) + ((g79) & (g80) & (!sk[71]) & (g81) & (g131) & (!g133)) + ((g79) & (g80) & (!sk[71]) & (g81) & (g131) & (g133)) + ((g79) & (g80) & (sk[71]) & (g81) & (!g131) & (g133)) + ((g79) & (g80) & (sk[71]) & (g81) & (g131) & (!g133)) + ((g79) & (g80) & (sk[71]) & (g81) & (g131) & (g133)));
	assign g135 = (((!sk[72]) & (g80) & (!g81)) + ((!sk[72]) & (g80) & (g81)) + ((sk[72]) & (g80) & (!g81)));
	assign g136 = (((!g78) & (!g79) & (!g135) & (!sk[73]) & (g82) & (!g83)) + ((!g78) & (!g79) & (!g135) & (!sk[73]) & (g82) & (g83)) + ((!g78) & (!g79) & (g135) & (!sk[73]) & (!g82) & (!g83)) + ((!g78) & (!g79) & (g135) & (!sk[73]) & (!g82) & (g83)) + ((!g78) & (!g79) & (g135) & (!sk[73]) & (g82) & (!g83)) + ((!g78) & (!g79) & (g135) & (!sk[73]) & (g82) & (g83)) + ((!g78) & (!g79) & (g135) & (sk[73]) & (!g82) & (g83)) + ((!g78) & (g79) & (!g135) & (!sk[73]) & (!g82) & (!g83)) + ((!g78) & (g79) & (!g135) & (!sk[73]) & (!g82) & (g83)) + ((!g78) & (g79) & (!g135) & (!sk[73]) & (g82) & (!g83)) + ((!g78) & (g79) & (!g135) & (!sk[73]) & (g82) & (g83)) + ((!g78) & (g79) & (g135) & (!sk[73]) & (!g82) & (!g83)) + ((!g78) & (g79) & (g135) & (!sk[73]) & (!g82) & (g83)) + ((!g78) & (g79) & (g135) & (!sk[73]) & (g82) & (!g83)) + ((!g78) & (g79) & (g135) & (!sk[73]) & (g82) & (g83)) + ((!g78) & (g79) & (g135) & (sk[73]) & (!g82) & (!g83)) + ((!g78) & (g79) & (g135) & (sk[73]) & (!g82) & (g83)) + ((g78) & (!g79) & (!g135) & (!sk[73]) & (g82) & (!g83)) + ((g78) & (!g79) & (!g135) & (!sk[73]) & (g82) & (g83)) + ((g78) & (!g79) & (g135) & (!sk[73]) & (!g82) & (!g83)) + ((g78) & (!g79) & (g135) & (!sk[73]) & (!g82) & (g83)) + ((g78) & (!g79) & (g135) & (!sk[73]) & (g82) & (!g83)) + ((g78) & (!g79) & (g135) & (!sk[73]) & (g82) & (g83)) + ((g78) & (!g79) & (g135) & (sk[73]) & (!g82) & (!g83)) + ((g78) & (!g79) & (g135) & (sk[73]) & (!g82) & (g83)) + ((g78) & (g79) & (!g135) & (!sk[73]) & (!g82) & (!g83)) + ((g78) & (g79) & (!g135) & (!sk[73]) & (!g82) & (g83)) + ((g78) & (g79) & (!g135) & (!sk[73]) & (g82) & (!g83)) + ((g78) & (g79) & (!g135) & (!sk[73]) & (g82) & (g83)) + ((g78) & (g79) & (g135) & (!sk[73]) & (!g82) & (!g83)) + ((g78) & (g79) & (g135) & (!sk[73]) & (!g82) & (g83)) + ((g78) & (g79) & (g135) & (!sk[73]) & (g82) & (!g83)) + ((g78) & (g79) & (g135) & (!sk[73]) & (g82) & (g83)) + ((g78) & (g79) & (g135) & (sk[73]) & (!g82) & (!g83)));
	assign g137 = (((!g132) & (!g134) & (!sk[74]) & (g136)) + ((!g132) & (!g134) & (sk[74]) & (!g136)) + ((!g132) & (g134) & (!sk[74]) & (!g136)) + ((!g132) & (g134) & (!sk[74]) & (g136)) + ((g132) & (!g134) & (!sk[74]) & (g136)) + ((g132) & (g134) & (!sk[74]) & (!g136)) + ((g132) & (g134) & (!sk[74]) & (g136)));
	assign g138 = (((g137) & (!sk[75]) & (!g126)) + ((g137) & (!sk[75]) & (g126)) + ((g137) & (sk[75]) & (g126)));
	assign g139 = (((!sk[76]) & (g130) & (!g138)) + ((!sk[76]) & (g130) & (g138)) + ((sk[76]) & (!g130) & (!g138)) + ((sk[76]) & (!g130) & (g138)) + ((sk[76]) & (g130) & (g138)));
	assign g140 = (((!sk[77]) & (g76) & (!g126)) + ((!sk[77]) & (g76) & (g126)) + ((sk[77]) & (g76) & (!g126)));
	assign g3981 = (((!g2059) & (!sk[78]) & (!g2069) & (g141)) + ((!g2059) & (!sk[78]) & (g2069) & (!g141)) + ((!g2059) & (!sk[78]) & (g2069) & (g141)) + ((!g2059) & (sk[78]) & (!g2069) & (g141)) + ((!g2059) & (sk[78]) & (g2069) & (g141)) + ((g2059) & (!sk[78]) & (!g2069) & (g141)) + ((g2059) & (!sk[78]) & (g2069) & (!g141)) + ((g2059) & (!sk[78]) & (g2069) & (g141)) + ((g2059) & (sk[78]) & (g2069) & (!g141)) + ((g2059) & (sk[78]) & (g2069) & (g141)));
	assign g3982 = (((!g2064) & (!dmem_dat_ix20x) & (!sk[79]) & (g142)) + ((!g2064) & (!dmem_dat_ix20x) & (sk[79]) & (g142)) + ((!g2064) & (dmem_dat_ix20x) & (!sk[79]) & (!g142)) + ((!g2064) & (dmem_dat_ix20x) & (!sk[79]) & (g142)) + ((!g2064) & (dmem_dat_ix20x) & (sk[79]) & (g142)) + ((g2064) & (!dmem_dat_ix20x) & (!sk[79]) & (g142)) + ((g2064) & (dmem_dat_ix20x) & (!sk[79]) & (!g142)) + ((g2064) & (dmem_dat_ix20x) & (!sk[79]) & (g142)) + ((g2064) & (dmem_dat_ix20x) & (sk[79]) & (!g142)) + ((g2064) & (dmem_dat_ix20x) & (sk[79]) & (g142)));
	assign g3983 = (((!sk[80]) & (!g2140) & (!g3777) & (g143)) + ((!sk[80]) & (!g2140) & (g3777) & (!g143)) + ((!sk[80]) & (!g2140) & (g3777) & (g143)) + ((!sk[80]) & (g2140) & (!g3777) & (g143)) + ((!sk[80]) & (g2140) & (g3777) & (!g143)) + ((!sk[80]) & (g2140) & (g3777) & (g143)) + ((sk[80]) & (!g2140) & (!g3777) & (g143)) + ((sk[80]) & (!g2140) & (g3777) & (g143)) + ((sk[80]) & (g2140) & (g3777) & (!g143)) + ((sk[80]) & (g2140) & (g3777) & (g143)));
	assign g3984 = (((!sk[81]) & (!g2142) & (!g3777) & (g144)) + ((!sk[81]) & (!g2142) & (g3777) & (!g144)) + ((!sk[81]) & (!g2142) & (g3777) & (g144)) + ((!sk[81]) & (g2142) & (!g3777) & (g144)) + ((!sk[81]) & (g2142) & (g3777) & (!g144)) + ((!sk[81]) & (g2142) & (g3777) & (g144)) + ((sk[81]) & (!g2142) & (!g3777) & (g144)) + ((sk[81]) & (!g2142) & (g3777) & (g144)) + ((sk[81]) & (g2142) & (g3777) & (!g144)) + ((sk[81]) & (g2142) & (g3777) & (g144)));
	assign g3985 = (((!g2144) & (!sk[82]) & (!g3777) & (g145)) + ((!g2144) & (!sk[82]) & (g3777) & (!g145)) + ((!g2144) & (!sk[82]) & (g3777) & (g145)) + ((!g2144) & (sk[82]) & (!g3777) & (g145)) + ((!g2144) & (sk[82]) & (g3777) & (g145)) + ((g2144) & (!sk[82]) & (!g3777) & (g145)) + ((g2144) & (!sk[82]) & (g3777) & (!g145)) + ((g2144) & (!sk[82]) & (g3777) & (g145)) + ((g2144) & (sk[82]) & (g3777) & (!g145)) + ((g2144) & (sk[82]) & (g3777) & (g145)));
	assign g3986 = (((!g2145) & (!g3777) & (!sk[83]) & (g146)) + ((!g2145) & (!g3777) & (sk[83]) & (g146)) + ((!g2145) & (g3777) & (!sk[83]) & (!g146)) + ((!g2145) & (g3777) & (!sk[83]) & (g146)) + ((!g2145) & (g3777) & (sk[83]) & (g146)) + ((g2145) & (!g3777) & (!sk[83]) & (g146)) + ((g2145) & (g3777) & (!sk[83]) & (!g146)) + ((g2145) & (g3777) & (!sk[83]) & (g146)) + ((g2145) & (g3777) & (sk[83]) & (!g146)) + ((g2145) & (g3777) & (sk[83]) & (g146)));
	assign g3987 = (((!g2064) & (!dmem_dat_ix19x) & (!sk[84]) & (g147)) + ((!g2064) & (!dmem_dat_ix19x) & (sk[84]) & (g147)) + ((!g2064) & (dmem_dat_ix19x) & (!sk[84]) & (!g147)) + ((!g2064) & (dmem_dat_ix19x) & (!sk[84]) & (g147)) + ((!g2064) & (dmem_dat_ix19x) & (sk[84]) & (g147)) + ((g2064) & (!dmem_dat_ix19x) & (!sk[84]) & (g147)) + ((g2064) & (dmem_dat_ix19x) & (!sk[84]) & (!g147)) + ((g2064) & (dmem_dat_ix19x) & (!sk[84]) & (g147)) + ((g2064) & (dmem_dat_ix19x) & (sk[84]) & (!g147)) + ((g2064) & (dmem_dat_ix19x) & (sk[84]) & (g147)));
	assign g3988 = (((!g2064) & (!dmem_dat_ix18x) & (!sk[85]) & (g148)) + ((!g2064) & (!dmem_dat_ix18x) & (sk[85]) & (g148)) + ((!g2064) & (dmem_dat_ix18x) & (!sk[85]) & (!g148)) + ((!g2064) & (dmem_dat_ix18x) & (!sk[85]) & (g148)) + ((!g2064) & (dmem_dat_ix18x) & (sk[85]) & (g148)) + ((g2064) & (!dmem_dat_ix18x) & (!sk[85]) & (g148)) + ((g2064) & (dmem_dat_ix18x) & (!sk[85]) & (!g148)) + ((g2064) & (dmem_dat_ix18x) & (!sk[85]) & (g148)) + ((g2064) & (dmem_dat_ix18x) & (sk[85]) & (!g148)) + ((g2064) & (dmem_dat_ix18x) & (sk[85]) & (g148)));
	assign g149 = (((!g143) & (!g144) & (!g145) & (g146) & (g147) & (g148)) + ((!g143) & (!g144) & (g145) & (!g146) & (!g147) & (g148)) + ((!g143) & (!g144) & (g145) & (g146) & (!g147) & (g148)) + ((!g143) & (!g144) & (g145) & (g146) & (g147) & (g148)) + ((!g143) & (g144) & (!g145) & (!g146) & (g147) & (!g148)) + ((!g143) & (g144) & (!g145) & (g146) & (g147) & (!g148)) + ((!g143) & (g144) & (!g145) & (g146) & (g147) & (g148)) + ((!g143) & (g144) & (g145) & (!g146) & (!g147) & (g148)) + ((!g143) & (g144) & (g145) & (!g146) & (g147) & (!g148)) + ((!g143) & (g144) & (g145) & (g146) & (!g147) & (g148)) + ((!g143) & (g144) & (g145) & (g146) & (g147) & (!g148)) + ((!g143) & (g144) & (g145) & (g146) & (g147) & (g148)) + ((g143) & (!g144) & (!g145) & (!g146) & (!g147) & (!g148)) + ((g143) & (!g144) & (!g145) & (g146) & (!g147) & (!g148)) + ((g143) & (!g144) & (!g145) & (g146) & (g147) & (g148)) + ((g143) & (!g144) & (g145) & (!g146) & (!g147) & (!g148)) + ((g143) & (!g144) & (g145) & (!g146) & (!g147) & (g148)) + ((g143) & (!g144) & (g145) & (g146) & (!g147) & (!g148)) + ((g143) & (!g144) & (g145) & (g146) & (!g147) & (g148)) + ((g143) & (!g144) & (g145) & (g146) & (g147) & (g148)) + ((g143) & (g144) & (!g145) & (!g146) & (!g147) & (!g148)) + ((g143) & (g144) & (!g145) & (!g146) & (g147) & (!g148)) + ((g143) & (g144) & (!g145) & (g146) & (!g147) & (!g148)) + ((g143) & (g144) & (!g145) & (g146) & (g147) & (!g148)) + ((g143) & (g144) & (!g145) & (g146) & (g147) & (g148)) + ((g143) & (g144) & (g145) & (!g146) & (!g147) & (!g148)) + ((g143) & (g144) & (g145) & (!g146) & (!g147) & (g148)) + ((g143) & (g144) & (g145) & (!g146) & (g147) & (!g148)) + ((g143) & (g144) & (g145) & (g146) & (!g147) & (!g148)) + ((g143) & (g144) & (g145) & (g146) & (!g147) & (g148)) + ((g143) & (g144) & (g145) & (g146) & (g147) & (!g148)) + ((g143) & (g144) & (g145) & (g146) & (g147) & (g148)));
	assign g3989 = (((!sk[87]) & (!g2146) & (!g3777) & (g150)) + ((!sk[87]) & (!g2146) & (g3777) & (!g150)) + ((!sk[87]) & (!g2146) & (g3777) & (g150)) + ((!sk[87]) & (g2146) & (!g3777) & (g150)) + ((!sk[87]) & (g2146) & (g3777) & (!g150)) + ((!sk[87]) & (g2146) & (g3777) & (g150)) + ((sk[87]) & (!g2146) & (!g3777) & (g150)) + ((sk[87]) & (!g2146) & (g3777) & (g150)) + ((sk[87]) & (g2146) & (g3777) & (!g150)) + ((sk[87]) & (g2146) & (g3777) & (g150)));
	assign g3990 = (((!g2148) & (!g3777) & (!sk[88]) & (g151)) + ((!g2148) & (!g3777) & (sk[88]) & (g151)) + ((!g2148) & (g3777) & (!sk[88]) & (!g151)) + ((!g2148) & (g3777) & (!sk[88]) & (g151)) + ((!g2148) & (g3777) & (sk[88]) & (g151)) + ((g2148) & (!g3777) & (!sk[88]) & (g151)) + ((g2148) & (g3777) & (!sk[88]) & (!g151)) + ((g2148) & (g3777) & (!sk[88]) & (g151)) + ((g2148) & (g3777) & (sk[88]) & (!g151)) + ((g2148) & (g3777) & (sk[88]) & (g151)));
	assign g3991 = (((!g2150) & (!g3777) & (!sk[89]) & (g152)) + ((!g2150) & (!g3777) & (sk[89]) & (g152)) + ((!g2150) & (g3777) & (!sk[89]) & (!g152)) + ((!g2150) & (g3777) & (!sk[89]) & (g152)) + ((!g2150) & (g3777) & (sk[89]) & (g152)) + ((g2150) & (!g3777) & (!sk[89]) & (g152)) + ((g2150) & (g3777) & (!sk[89]) & (!g152)) + ((g2150) & (g3777) & (!sk[89]) & (g152)) + ((g2150) & (g3777) & (sk[89]) & (!g152)) + ((g2150) & (g3777) & (sk[89]) & (g152)));
	assign g3992 = (((!g2151) & (!g3777) & (!sk[90]) & (g153)) + ((!g2151) & (!g3777) & (sk[90]) & (g153)) + ((!g2151) & (g3777) & (!sk[90]) & (!g153)) + ((!g2151) & (g3777) & (!sk[90]) & (g153)) + ((!g2151) & (g3777) & (sk[90]) & (g153)) + ((g2151) & (!g3777) & (!sk[90]) & (g153)) + ((g2151) & (g3777) & (!sk[90]) & (!g153)) + ((g2151) & (g3777) & (!sk[90]) & (g153)) + ((g2151) & (g3777) & (sk[90]) & (!g153)) + ((g2151) & (g3777) & (sk[90]) & (g153)));
	assign g154 = (((!g150) & (!g151) & (!g152) & (g153) & (g147) & (g148)) + ((!g150) & (!g151) & (g152) & (!g153) & (!g147) & (g148)) + ((!g150) & (!g151) & (g152) & (g153) & (!g147) & (g148)) + ((!g150) & (!g151) & (g152) & (g153) & (g147) & (g148)) + ((!g150) & (g151) & (!g152) & (!g153) & (g147) & (!g148)) + ((!g150) & (g151) & (!g152) & (g153) & (g147) & (!g148)) + ((!g150) & (g151) & (!g152) & (g153) & (g147) & (g148)) + ((!g150) & (g151) & (g152) & (!g153) & (!g147) & (g148)) + ((!g150) & (g151) & (g152) & (!g153) & (g147) & (!g148)) + ((!g150) & (g151) & (g152) & (g153) & (!g147) & (g148)) + ((!g150) & (g151) & (g152) & (g153) & (g147) & (!g148)) + ((!g150) & (g151) & (g152) & (g153) & (g147) & (g148)) + ((g150) & (!g151) & (!g152) & (!g153) & (!g147) & (!g148)) + ((g150) & (!g151) & (!g152) & (g153) & (!g147) & (!g148)) + ((g150) & (!g151) & (!g152) & (g153) & (g147) & (g148)) + ((g150) & (!g151) & (g152) & (!g153) & (!g147) & (!g148)) + ((g150) & (!g151) & (g152) & (!g153) & (!g147) & (g148)) + ((g150) & (!g151) & (g152) & (g153) & (!g147) & (!g148)) + ((g150) & (!g151) & (g152) & (g153) & (!g147) & (g148)) + ((g150) & (!g151) & (g152) & (g153) & (g147) & (g148)) + ((g150) & (g151) & (!g152) & (!g153) & (!g147) & (!g148)) + ((g150) & (g151) & (!g152) & (!g153) & (g147) & (!g148)) + ((g150) & (g151) & (!g152) & (g153) & (!g147) & (!g148)) + ((g150) & (g151) & (!g152) & (g153) & (g147) & (!g148)) + ((g150) & (g151) & (!g152) & (g153) & (g147) & (g148)) + ((g150) & (g151) & (g152) & (!g153) & (!g147) & (!g148)) + ((g150) & (g151) & (g152) & (!g153) & (!g147) & (g148)) + ((g150) & (g151) & (g152) & (!g153) & (g147) & (!g148)) + ((g150) & (g151) & (g152) & (g153) & (!g147) & (!g148)) + ((g150) & (g151) & (g152) & (g153) & (!g147) & (g148)) + ((g150) & (g151) & (g152) & (g153) & (g147) & (!g148)) + ((g150) & (g151) & (g152) & (g153) & (g147) & (g148)));
	assign g3993 = (((!g2152) & (!g3777) & (!sk[92]) & (g155)) + ((!g2152) & (!g3777) & (sk[92]) & (g155)) + ((!g2152) & (g3777) & (!sk[92]) & (!g155)) + ((!g2152) & (g3777) & (!sk[92]) & (g155)) + ((!g2152) & (g3777) & (sk[92]) & (g155)) + ((g2152) & (!g3777) & (!sk[92]) & (g155)) + ((g2152) & (g3777) & (!sk[92]) & (!g155)) + ((g2152) & (g3777) & (!sk[92]) & (g155)) + ((g2152) & (g3777) & (sk[92]) & (!g155)) + ((g2152) & (g3777) & (sk[92]) & (g155)));
	assign g3994 = (((!g2153) & (!g3777) & (!sk[93]) & (g156)) + ((!g2153) & (!g3777) & (sk[93]) & (g156)) + ((!g2153) & (g3777) & (!sk[93]) & (!g156)) + ((!g2153) & (g3777) & (!sk[93]) & (g156)) + ((!g2153) & (g3777) & (sk[93]) & (g156)) + ((g2153) & (!g3777) & (!sk[93]) & (g156)) + ((g2153) & (g3777) & (!sk[93]) & (!g156)) + ((g2153) & (g3777) & (!sk[93]) & (g156)) + ((g2153) & (g3777) & (sk[93]) & (!g156)) + ((g2153) & (g3777) & (sk[93]) & (g156)));
	assign g3995 = (((!g2155) & (!sk[94]) & (!g3777) & (g157)) + ((!g2155) & (!sk[94]) & (g3777) & (!g157)) + ((!g2155) & (!sk[94]) & (g3777) & (g157)) + ((!g2155) & (sk[94]) & (!g3777) & (g157)) + ((!g2155) & (sk[94]) & (g3777) & (g157)) + ((g2155) & (!sk[94]) & (!g3777) & (g157)) + ((g2155) & (!sk[94]) & (g3777) & (!g157)) + ((g2155) & (!sk[94]) & (g3777) & (g157)) + ((g2155) & (sk[94]) & (g3777) & (!g157)) + ((g2155) & (sk[94]) & (g3777) & (g157)));
	assign g3996 = (((!sk[95]) & (!g2157) & (!g3777) & (g158)) + ((!sk[95]) & (!g2157) & (g3777) & (!g158)) + ((!sk[95]) & (!g2157) & (g3777) & (g158)) + ((!sk[95]) & (g2157) & (!g3777) & (g158)) + ((!sk[95]) & (g2157) & (g3777) & (!g158)) + ((!sk[95]) & (g2157) & (g3777) & (g158)) + ((sk[95]) & (!g2157) & (!g3777) & (g158)) + ((sk[95]) & (!g2157) & (g3777) & (g158)) + ((sk[95]) & (g2157) & (g3777) & (!g158)) + ((sk[95]) & (g2157) & (g3777) & (g158)));
	assign g159 = (((!g155) & (!g156) & (!g157) & (g158) & (g147) & (g148)) + ((!g155) & (!g156) & (g157) & (!g158) & (!g147) & (g148)) + ((!g155) & (!g156) & (g157) & (g158) & (!g147) & (g148)) + ((!g155) & (!g156) & (g157) & (g158) & (g147) & (g148)) + ((!g155) & (g156) & (!g157) & (!g158) & (g147) & (!g148)) + ((!g155) & (g156) & (!g157) & (g158) & (g147) & (!g148)) + ((!g155) & (g156) & (!g157) & (g158) & (g147) & (g148)) + ((!g155) & (g156) & (g157) & (!g158) & (!g147) & (g148)) + ((!g155) & (g156) & (g157) & (!g158) & (g147) & (!g148)) + ((!g155) & (g156) & (g157) & (g158) & (!g147) & (g148)) + ((!g155) & (g156) & (g157) & (g158) & (g147) & (!g148)) + ((!g155) & (g156) & (g157) & (g158) & (g147) & (g148)) + ((g155) & (!g156) & (!g157) & (!g158) & (!g147) & (!g148)) + ((g155) & (!g156) & (!g157) & (g158) & (!g147) & (!g148)) + ((g155) & (!g156) & (!g157) & (g158) & (g147) & (g148)) + ((g155) & (!g156) & (g157) & (!g158) & (!g147) & (!g148)) + ((g155) & (!g156) & (g157) & (!g158) & (!g147) & (g148)) + ((g155) & (!g156) & (g157) & (g158) & (!g147) & (!g148)) + ((g155) & (!g156) & (g157) & (g158) & (!g147) & (g148)) + ((g155) & (!g156) & (g157) & (g158) & (g147) & (g148)) + ((g155) & (g156) & (!g157) & (!g158) & (!g147) & (!g148)) + ((g155) & (g156) & (!g157) & (!g158) & (g147) & (!g148)) + ((g155) & (g156) & (!g157) & (g158) & (!g147) & (!g148)) + ((g155) & (g156) & (!g157) & (g158) & (g147) & (!g148)) + ((g155) & (g156) & (!g157) & (g158) & (g147) & (g148)) + ((g155) & (g156) & (g157) & (!g158) & (!g147) & (!g148)) + ((g155) & (g156) & (g157) & (!g158) & (!g147) & (g148)) + ((g155) & (g156) & (g157) & (!g158) & (g147) & (!g148)) + ((g155) & (g156) & (g157) & (g158) & (!g147) & (!g148)) + ((g155) & (g156) & (g157) & (g158) & (!g147) & (g148)) + ((g155) & (g156) & (g157) & (g158) & (g147) & (!g148)) + ((g155) & (g156) & (g157) & (g158) & (g147) & (g148)));
	assign g3997 = (((!g2158) & (!g3777) & (!sk[97]) & (g160)) + ((!g2158) & (!g3777) & (sk[97]) & (g160)) + ((!g2158) & (g3777) & (!sk[97]) & (!g160)) + ((!g2158) & (g3777) & (!sk[97]) & (g160)) + ((!g2158) & (g3777) & (sk[97]) & (g160)) + ((g2158) & (!g3777) & (!sk[97]) & (g160)) + ((g2158) & (g3777) & (!sk[97]) & (!g160)) + ((g2158) & (g3777) & (!sk[97]) & (g160)) + ((g2158) & (g3777) & (sk[97]) & (!g160)) + ((g2158) & (g3777) & (sk[97]) & (g160)));
	assign g3998 = (((!g2159) & (!g3777) & (!sk[98]) & (g161)) + ((!g2159) & (!g3777) & (sk[98]) & (g161)) + ((!g2159) & (g3777) & (!sk[98]) & (!g161)) + ((!g2159) & (g3777) & (!sk[98]) & (g161)) + ((!g2159) & (g3777) & (sk[98]) & (g161)) + ((g2159) & (!g3777) & (!sk[98]) & (g161)) + ((g2159) & (g3777) & (!sk[98]) & (!g161)) + ((g2159) & (g3777) & (!sk[98]) & (g161)) + ((g2159) & (g3777) & (sk[98]) & (!g161)) + ((g2159) & (g3777) & (sk[98]) & (g161)));
	assign g3999 = (((!g2160) & (!sk[99]) & (!g3777) & (g162)) + ((!g2160) & (!sk[99]) & (g3777) & (!g162)) + ((!g2160) & (!sk[99]) & (g3777) & (g162)) + ((!g2160) & (sk[99]) & (!g3777) & (g162)) + ((!g2160) & (sk[99]) & (g3777) & (g162)) + ((g2160) & (!sk[99]) & (!g3777) & (g162)) + ((g2160) & (!sk[99]) & (g3777) & (!g162)) + ((g2160) & (!sk[99]) & (g3777) & (g162)) + ((g2160) & (sk[99]) & (g3777) & (!g162)) + ((g2160) & (sk[99]) & (g3777) & (g162)));
	assign g4000 = (((!sk[100]) & (!g2161) & (!g3777) & (g163)) + ((!sk[100]) & (!g2161) & (g3777) & (!g163)) + ((!sk[100]) & (!g2161) & (g3777) & (g163)) + ((!sk[100]) & (g2161) & (!g3777) & (g163)) + ((!sk[100]) & (g2161) & (g3777) & (!g163)) + ((!sk[100]) & (g2161) & (g3777) & (g163)) + ((sk[100]) & (!g2161) & (!g3777) & (g163)) + ((sk[100]) & (!g2161) & (g3777) & (g163)) + ((sk[100]) & (g2161) & (g3777) & (!g163)) + ((sk[100]) & (g2161) & (g3777) & (g163)));
	assign g164 = (((!g160) & (!g161) & (!g162) & (g163) & (g147) & (g148)) + ((!g160) & (!g161) & (g162) & (!g163) & (!g147) & (g148)) + ((!g160) & (!g161) & (g162) & (g163) & (!g147) & (g148)) + ((!g160) & (!g161) & (g162) & (g163) & (g147) & (g148)) + ((!g160) & (g161) & (!g162) & (!g163) & (g147) & (!g148)) + ((!g160) & (g161) & (!g162) & (g163) & (g147) & (!g148)) + ((!g160) & (g161) & (!g162) & (g163) & (g147) & (g148)) + ((!g160) & (g161) & (g162) & (!g163) & (!g147) & (g148)) + ((!g160) & (g161) & (g162) & (!g163) & (g147) & (!g148)) + ((!g160) & (g161) & (g162) & (g163) & (!g147) & (g148)) + ((!g160) & (g161) & (g162) & (g163) & (g147) & (!g148)) + ((!g160) & (g161) & (g162) & (g163) & (g147) & (g148)) + ((g160) & (!g161) & (!g162) & (!g163) & (!g147) & (!g148)) + ((g160) & (!g161) & (!g162) & (g163) & (!g147) & (!g148)) + ((g160) & (!g161) & (!g162) & (g163) & (g147) & (g148)) + ((g160) & (!g161) & (g162) & (!g163) & (!g147) & (!g148)) + ((g160) & (!g161) & (g162) & (!g163) & (!g147) & (g148)) + ((g160) & (!g161) & (g162) & (g163) & (!g147) & (!g148)) + ((g160) & (!g161) & (g162) & (g163) & (!g147) & (g148)) + ((g160) & (!g161) & (g162) & (g163) & (g147) & (g148)) + ((g160) & (g161) & (!g162) & (!g163) & (!g147) & (!g148)) + ((g160) & (g161) & (!g162) & (!g163) & (g147) & (!g148)) + ((g160) & (g161) & (!g162) & (g163) & (!g147) & (!g148)) + ((g160) & (g161) & (!g162) & (g163) & (g147) & (!g148)) + ((g160) & (g161) & (!g162) & (g163) & (g147) & (g148)) + ((g160) & (g161) & (g162) & (!g163) & (!g147) & (!g148)) + ((g160) & (g161) & (g162) & (!g163) & (!g147) & (g148)) + ((g160) & (g161) & (g162) & (!g163) & (g147) & (!g148)) + ((g160) & (g161) & (g162) & (g163) & (!g147) & (!g148)) + ((g160) & (g161) & (g162) & (g163) & (!g147) & (g148)) + ((g160) & (g161) & (g162) & (g163) & (g147) & (!g148)) + ((g160) & (g161) & (g162) & (g163) & (g147) & (g148)));
	assign g4001 = (((!sk[102]) & (!g2064) & (!dmem_dat_ix16x) & (g165)) + ((!sk[102]) & (!g2064) & (dmem_dat_ix16x) & (!g165)) + ((!sk[102]) & (!g2064) & (dmem_dat_ix16x) & (g165)) + ((!sk[102]) & (g2064) & (!dmem_dat_ix16x) & (g165)) + ((!sk[102]) & (g2064) & (dmem_dat_ix16x) & (!g165)) + ((!sk[102]) & (g2064) & (dmem_dat_ix16x) & (g165)) + ((sk[102]) & (!g2064) & (!dmem_dat_ix16x) & (g165)) + ((sk[102]) & (!g2064) & (dmem_dat_ix16x) & (g165)) + ((sk[102]) & (g2064) & (dmem_dat_ix16x) & (!g165)) + ((sk[102]) & (g2064) & (dmem_dat_ix16x) & (g165)));
	assign g4002 = (((!sk[103]) & (!g2064) & (!dmem_dat_ix17x) & (g166)) + ((!sk[103]) & (!g2064) & (dmem_dat_ix17x) & (!g166)) + ((!sk[103]) & (!g2064) & (dmem_dat_ix17x) & (g166)) + ((!sk[103]) & (g2064) & (!dmem_dat_ix17x) & (g166)) + ((!sk[103]) & (g2064) & (dmem_dat_ix17x) & (!g166)) + ((!sk[103]) & (g2064) & (dmem_dat_ix17x) & (g166)) + ((sk[103]) & (!g2064) & (!dmem_dat_ix17x) & (g166)) + ((sk[103]) & (!g2064) & (dmem_dat_ix17x) & (g166)) + ((sk[103]) & (g2064) & (dmem_dat_ix17x) & (!g166)) + ((sk[103]) & (g2064) & (dmem_dat_ix17x) & (g166)));
	assign g167 = (((!g149) & (!g154) & (!g159) & (g164) & (g165) & (g166)) + ((!g149) & (!g154) & (g159) & (!g164) & (!g165) & (g166)) + ((!g149) & (!g154) & (g159) & (g164) & (!g165) & (g166)) + ((!g149) & (!g154) & (g159) & (g164) & (g165) & (g166)) + ((!g149) & (g154) & (!g159) & (!g164) & (g165) & (!g166)) + ((!g149) & (g154) & (!g159) & (g164) & (g165) & (!g166)) + ((!g149) & (g154) & (!g159) & (g164) & (g165) & (g166)) + ((!g149) & (g154) & (g159) & (!g164) & (!g165) & (g166)) + ((!g149) & (g154) & (g159) & (!g164) & (g165) & (!g166)) + ((!g149) & (g154) & (g159) & (g164) & (!g165) & (g166)) + ((!g149) & (g154) & (g159) & (g164) & (g165) & (!g166)) + ((!g149) & (g154) & (g159) & (g164) & (g165) & (g166)) + ((g149) & (!g154) & (!g159) & (!g164) & (!g165) & (!g166)) + ((g149) & (!g154) & (!g159) & (g164) & (!g165) & (!g166)) + ((g149) & (!g154) & (!g159) & (g164) & (g165) & (g166)) + ((g149) & (!g154) & (g159) & (!g164) & (!g165) & (!g166)) + ((g149) & (!g154) & (g159) & (!g164) & (!g165) & (g166)) + ((g149) & (!g154) & (g159) & (g164) & (!g165) & (!g166)) + ((g149) & (!g154) & (g159) & (g164) & (!g165) & (g166)) + ((g149) & (!g154) & (g159) & (g164) & (g165) & (g166)) + ((g149) & (g154) & (!g159) & (!g164) & (!g165) & (!g166)) + ((g149) & (g154) & (!g159) & (!g164) & (g165) & (!g166)) + ((g149) & (g154) & (!g159) & (g164) & (!g165) & (!g166)) + ((g149) & (g154) & (!g159) & (g164) & (g165) & (!g166)) + ((g149) & (g154) & (!g159) & (g164) & (g165) & (g166)) + ((g149) & (g154) & (g159) & (!g164) & (!g165) & (!g166)) + ((g149) & (g154) & (g159) & (!g164) & (!g165) & (g166)) + ((g149) & (g154) & (g159) & (!g164) & (g165) & (!g166)) + ((g149) & (g154) & (g159) & (g164) & (!g165) & (!g166)) + ((g149) & (g154) & (g159) & (g164) & (!g165) & (g166)) + ((g149) & (g154) & (g159) & (g164) & (g165) & (!g166)) + ((g149) & (g154) & (g159) & (g164) & (g165) & (g166)));
	assign g4003 = (((!g2162) & (!g3777) & (!sk[105]) & (g168)) + ((!g2162) & (!g3777) & (sk[105]) & (g168)) + ((!g2162) & (g3777) & (!sk[105]) & (!g168)) + ((!g2162) & (g3777) & (!sk[105]) & (g168)) + ((!g2162) & (g3777) & (sk[105]) & (g168)) + ((g2162) & (!g3777) & (!sk[105]) & (g168)) + ((g2162) & (g3777) & (!sk[105]) & (!g168)) + ((g2162) & (g3777) & (!sk[105]) & (g168)) + ((g2162) & (g3777) & (sk[105]) & (!g168)) + ((g2162) & (g3777) & (sk[105]) & (g168)));
	assign g4004 = (((!g2164) & (!sk[106]) & (!g3777) & (g169)) + ((!g2164) & (!sk[106]) & (g3777) & (!g169)) + ((!g2164) & (!sk[106]) & (g3777) & (g169)) + ((!g2164) & (sk[106]) & (!g3777) & (g169)) + ((!g2164) & (sk[106]) & (g3777) & (g169)) + ((g2164) & (!sk[106]) & (!g3777) & (g169)) + ((g2164) & (!sk[106]) & (g3777) & (!g169)) + ((g2164) & (!sk[106]) & (g3777) & (g169)) + ((g2164) & (sk[106]) & (g3777) & (!g169)) + ((g2164) & (sk[106]) & (g3777) & (g169)));
	assign g4005 = (((!g2166) & (!g3777) & (!sk[107]) & (g170)) + ((!g2166) & (!g3777) & (sk[107]) & (g170)) + ((!g2166) & (g3777) & (!sk[107]) & (!g170)) + ((!g2166) & (g3777) & (!sk[107]) & (g170)) + ((!g2166) & (g3777) & (sk[107]) & (g170)) + ((g2166) & (!g3777) & (!sk[107]) & (g170)) + ((g2166) & (g3777) & (!sk[107]) & (!g170)) + ((g2166) & (g3777) & (!sk[107]) & (g170)) + ((g2166) & (g3777) & (sk[107]) & (!g170)) + ((g2166) & (g3777) & (sk[107]) & (g170)));
	assign g4006 = (((!g2168) & (!g3777) & (!sk[108]) & (g171)) + ((!g2168) & (!g3777) & (sk[108]) & (g171)) + ((!g2168) & (g3777) & (!sk[108]) & (!g171)) + ((!g2168) & (g3777) & (!sk[108]) & (g171)) + ((!g2168) & (g3777) & (sk[108]) & (g171)) + ((g2168) & (!g3777) & (!sk[108]) & (g171)) + ((g2168) & (g3777) & (!sk[108]) & (!g171)) + ((g2168) & (g3777) & (!sk[108]) & (g171)) + ((g2168) & (g3777) & (sk[108]) & (!g171)) + ((g2168) & (g3777) & (sk[108]) & (g171)));
	assign g172 = (((!g168) & (!g169) & (!g170) & (g171) & (g165) & (g166)) + ((!g168) & (!g169) & (g170) & (!g171) & (!g165) & (g166)) + ((!g168) & (!g169) & (g170) & (g171) & (!g165) & (g166)) + ((!g168) & (!g169) & (g170) & (g171) & (g165) & (g166)) + ((!g168) & (g169) & (!g170) & (!g171) & (g165) & (!g166)) + ((!g168) & (g169) & (!g170) & (g171) & (g165) & (!g166)) + ((!g168) & (g169) & (!g170) & (g171) & (g165) & (g166)) + ((!g168) & (g169) & (g170) & (!g171) & (!g165) & (g166)) + ((!g168) & (g169) & (g170) & (!g171) & (g165) & (!g166)) + ((!g168) & (g169) & (g170) & (g171) & (!g165) & (g166)) + ((!g168) & (g169) & (g170) & (g171) & (g165) & (!g166)) + ((!g168) & (g169) & (g170) & (g171) & (g165) & (g166)) + ((g168) & (!g169) & (!g170) & (!g171) & (!g165) & (!g166)) + ((g168) & (!g169) & (!g170) & (g171) & (!g165) & (!g166)) + ((g168) & (!g169) & (!g170) & (g171) & (g165) & (g166)) + ((g168) & (!g169) & (g170) & (!g171) & (!g165) & (!g166)) + ((g168) & (!g169) & (g170) & (!g171) & (!g165) & (g166)) + ((g168) & (!g169) & (g170) & (g171) & (!g165) & (!g166)) + ((g168) & (!g169) & (g170) & (g171) & (!g165) & (g166)) + ((g168) & (!g169) & (g170) & (g171) & (g165) & (g166)) + ((g168) & (g169) & (!g170) & (!g171) & (!g165) & (!g166)) + ((g168) & (g169) & (!g170) & (!g171) & (g165) & (!g166)) + ((g168) & (g169) & (!g170) & (g171) & (!g165) & (!g166)) + ((g168) & (g169) & (!g170) & (g171) & (g165) & (!g166)) + ((g168) & (g169) & (!g170) & (g171) & (g165) & (g166)) + ((g168) & (g169) & (g170) & (!g171) & (!g165) & (!g166)) + ((g168) & (g169) & (g170) & (!g171) & (!g165) & (g166)) + ((g168) & (g169) & (g170) & (!g171) & (g165) & (!g166)) + ((g168) & (g169) & (g170) & (g171) & (!g165) & (!g166)) + ((g168) & (g169) & (g170) & (g171) & (!g165) & (g166)) + ((g168) & (g169) & (g170) & (g171) & (g165) & (!g166)) + ((g168) & (g169) & (g170) & (g171) & (g165) & (g166)));
	assign g4007 = (((!sk[110]) & (!g2169) & (!g3777) & (g173)) + ((!sk[110]) & (!g2169) & (g3777) & (!g173)) + ((!sk[110]) & (!g2169) & (g3777) & (g173)) + ((!sk[110]) & (g2169) & (!g3777) & (g173)) + ((!sk[110]) & (g2169) & (g3777) & (!g173)) + ((!sk[110]) & (g2169) & (g3777) & (g173)) + ((sk[110]) & (!g2169) & (!g3777) & (g173)) + ((sk[110]) & (!g2169) & (g3777) & (g173)) + ((sk[110]) & (g2169) & (g3777) & (!g173)) + ((sk[110]) & (g2169) & (g3777) & (g173)));
	assign g4008 = (((!g2170) & (!g3777) & (!sk[111]) & (g174)) + ((!g2170) & (!g3777) & (sk[111]) & (g174)) + ((!g2170) & (g3777) & (!sk[111]) & (!g174)) + ((!g2170) & (g3777) & (!sk[111]) & (g174)) + ((!g2170) & (g3777) & (sk[111]) & (g174)) + ((g2170) & (!g3777) & (!sk[111]) & (g174)) + ((g2170) & (g3777) & (!sk[111]) & (!g174)) + ((g2170) & (g3777) & (!sk[111]) & (g174)) + ((g2170) & (g3777) & (sk[111]) & (!g174)) + ((g2170) & (g3777) & (sk[111]) & (g174)));
	assign g4009 = (((!sk[112]) & (!g2171) & (!g3777) & (g175)) + ((!sk[112]) & (!g2171) & (g3777) & (!g175)) + ((!sk[112]) & (!g2171) & (g3777) & (g175)) + ((!sk[112]) & (g2171) & (!g3777) & (g175)) + ((!sk[112]) & (g2171) & (g3777) & (!g175)) + ((!sk[112]) & (g2171) & (g3777) & (g175)) + ((sk[112]) & (!g2171) & (!g3777) & (g175)) + ((sk[112]) & (!g2171) & (g3777) & (g175)) + ((sk[112]) & (g2171) & (g3777) & (!g175)) + ((sk[112]) & (g2171) & (g3777) & (g175)));
	assign g4010 = (((!g2172) & (!sk[113]) & (!g3777) & (g176)) + ((!g2172) & (!sk[113]) & (g3777) & (!g176)) + ((!g2172) & (!sk[113]) & (g3777) & (g176)) + ((!g2172) & (sk[113]) & (!g3777) & (g176)) + ((!g2172) & (sk[113]) & (g3777) & (g176)) + ((g2172) & (!sk[113]) & (!g3777) & (g176)) + ((g2172) & (!sk[113]) & (g3777) & (!g176)) + ((g2172) & (!sk[113]) & (g3777) & (g176)) + ((g2172) & (sk[113]) & (g3777) & (!g176)) + ((g2172) & (sk[113]) & (g3777) & (g176)));
	assign g177 = (((!g173) & (!g174) & (!g175) & (g176) & (g165) & (g166)) + ((!g173) & (!g174) & (g175) & (!g176) & (!g165) & (g166)) + ((!g173) & (!g174) & (g175) & (g176) & (!g165) & (g166)) + ((!g173) & (!g174) & (g175) & (g176) & (g165) & (g166)) + ((!g173) & (g174) & (!g175) & (!g176) & (g165) & (!g166)) + ((!g173) & (g174) & (!g175) & (g176) & (g165) & (!g166)) + ((!g173) & (g174) & (!g175) & (g176) & (g165) & (g166)) + ((!g173) & (g174) & (g175) & (!g176) & (!g165) & (g166)) + ((!g173) & (g174) & (g175) & (!g176) & (g165) & (!g166)) + ((!g173) & (g174) & (g175) & (g176) & (!g165) & (g166)) + ((!g173) & (g174) & (g175) & (g176) & (g165) & (!g166)) + ((!g173) & (g174) & (g175) & (g176) & (g165) & (g166)) + ((g173) & (!g174) & (!g175) & (!g176) & (!g165) & (!g166)) + ((g173) & (!g174) & (!g175) & (g176) & (!g165) & (!g166)) + ((g173) & (!g174) & (!g175) & (g176) & (g165) & (g166)) + ((g173) & (!g174) & (g175) & (!g176) & (!g165) & (!g166)) + ((g173) & (!g174) & (g175) & (!g176) & (!g165) & (g166)) + ((g173) & (!g174) & (g175) & (g176) & (!g165) & (!g166)) + ((g173) & (!g174) & (g175) & (g176) & (!g165) & (g166)) + ((g173) & (!g174) & (g175) & (g176) & (g165) & (g166)) + ((g173) & (g174) & (!g175) & (!g176) & (!g165) & (!g166)) + ((g173) & (g174) & (!g175) & (!g176) & (g165) & (!g166)) + ((g173) & (g174) & (!g175) & (g176) & (!g165) & (!g166)) + ((g173) & (g174) & (!g175) & (g176) & (g165) & (!g166)) + ((g173) & (g174) & (!g175) & (g176) & (g165) & (g166)) + ((g173) & (g174) & (g175) & (!g176) & (!g165) & (!g166)) + ((g173) & (g174) & (g175) & (!g176) & (!g165) & (g166)) + ((g173) & (g174) & (g175) & (!g176) & (g165) & (!g166)) + ((g173) & (g174) & (g175) & (g176) & (!g165) & (!g166)) + ((g173) & (g174) & (g175) & (g176) & (!g165) & (g166)) + ((g173) & (g174) & (g175) & (g176) & (g165) & (!g166)) + ((g173) & (g174) & (g175) & (g176) & (g165) & (g166)));
	assign g4011 = (((!sk[115]) & (!g2173) & (!g3777) & (g178)) + ((!sk[115]) & (!g2173) & (g3777) & (!g178)) + ((!sk[115]) & (!g2173) & (g3777) & (g178)) + ((!sk[115]) & (g2173) & (!g3777) & (g178)) + ((!sk[115]) & (g2173) & (g3777) & (!g178)) + ((!sk[115]) & (g2173) & (g3777) & (g178)) + ((sk[115]) & (!g2173) & (!g3777) & (g178)) + ((sk[115]) & (!g2173) & (g3777) & (g178)) + ((sk[115]) & (g2173) & (g3777) & (!g178)) + ((sk[115]) & (g2173) & (g3777) & (g178)));
	assign g4012 = (((!g2174) & (!sk[116]) & (!g3777) & (g179)) + ((!g2174) & (!sk[116]) & (g3777) & (!g179)) + ((!g2174) & (!sk[116]) & (g3777) & (g179)) + ((!g2174) & (sk[116]) & (!g3777) & (g179)) + ((!g2174) & (sk[116]) & (g3777) & (g179)) + ((g2174) & (!sk[116]) & (!g3777) & (g179)) + ((g2174) & (!sk[116]) & (g3777) & (!g179)) + ((g2174) & (!sk[116]) & (g3777) & (g179)) + ((g2174) & (sk[116]) & (g3777) & (!g179)) + ((g2174) & (sk[116]) & (g3777) & (g179)));
	assign g4013 = (((!g2175) & (!g3777) & (!sk[117]) & (g180)) + ((!g2175) & (!g3777) & (sk[117]) & (g180)) + ((!g2175) & (g3777) & (!sk[117]) & (!g180)) + ((!g2175) & (g3777) & (!sk[117]) & (g180)) + ((!g2175) & (g3777) & (sk[117]) & (g180)) + ((g2175) & (!g3777) & (!sk[117]) & (g180)) + ((g2175) & (g3777) & (!sk[117]) & (!g180)) + ((g2175) & (g3777) & (!sk[117]) & (g180)) + ((g2175) & (g3777) & (sk[117]) & (!g180)) + ((g2175) & (g3777) & (sk[117]) & (g180)));
	assign g4014 = (((!g2176) & (!g3777) & (!sk[118]) & (g181)) + ((!g2176) & (!g3777) & (sk[118]) & (g181)) + ((!g2176) & (g3777) & (!sk[118]) & (!g181)) + ((!g2176) & (g3777) & (!sk[118]) & (g181)) + ((!g2176) & (g3777) & (sk[118]) & (g181)) + ((g2176) & (!g3777) & (!sk[118]) & (g181)) + ((g2176) & (g3777) & (!sk[118]) & (!g181)) + ((g2176) & (g3777) & (!sk[118]) & (g181)) + ((g2176) & (g3777) & (sk[118]) & (!g181)) + ((g2176) & (g3777) & (sk[118]) & (g181)));
	assign g182 = (((!g178) & (!g179) & (!g180) & (g181) & (g165) & (g166)) + ((!g178) & (!g179) & (g180) & (!g181) & (!g165) & (g166)) + ((!g178) & (!g179) & (g180) & (g181) & (!g165) & (g166)) + ((!g178) & (!g179) & (g180) & (g181) & (g165) & (g166)) + ((!g178) & (g179) & (!g180) & (!g181) & (g165) & (!g166)) + ((!g178) & (g179) & (!g180) & (g181) & (g165) & (!g166)) + ((!g178) & (g179) & (!g180) & (g181) & (g165) & (g166)) + ((!g178) & (g179) & (g180) & (!g181) & (!g165) & (g166)) + ((!g178) & (g179) & (g180) & (!g181) & (g165) & (!g166)) + ((!g178) & (g179) & (g180) & (g181) & (!g165) & (g166)) + ((!g178) & (g179) & (g180) & (g181) & (g165) & (!g166)) + ((!g178) & (g179) & (g180) & (g181) & (g165) & (g166)) + ((g178) & (!g179) & (!g180) & (!g181) & (!g165) & (!g166)) + ((g178) & (!g179) & (!g180) & (g181) & (!g165) & (!g166)) + ((g178) & (!g179) & (!g180) & (g181) & (g165) & (g166)) + ((g178) & (!g179) & (g180) & (!g181) & (!g165) & (!g166)) + ((g178) & (!g179) & (g180) & (!g181) & (!g165) & (g166)) + ((g178) & (!g179) & (g180) & (g181) & (!g165) & (!g166)) + ((g178) & (!g179) & (g180) & (g181) & (!g165) & (g166)) + ((g178) & (!g179) & (g180) & (g181) & (g165) & (g166)) + ((g178) & (g179) & (!g180) & (!g181) & (!g165) & (!g166)) + ((g178) & (g179) & (!g180) & (!g181) & (g165) & (!g166)) + ((g178) & (g179) & (!g180) & (g181) & (!g165) & (!g166)) + ((g178) & (g179) & (!g180) & (g181) & (g165) & (!g166)) + ((g178) & (g179) & (!g180) & (g181) & (g165) & (g166)) + ((g178) & (g179) & (g180) & (!g181) & (!g165) & (!g166)) + ((g178) & (g179) & (g180) & (!g181) & (!g165) & (g166)) + ((g178) & (g179) & (g180) & (!g181) & (g165) & (!g166)) + ((g178) & (g179) & (g180) & (g181) & (!g165) & (!g166)) + ((g178) & (g179) & (g180) & (g181) & (!g165) & (g166)) + ((g178) & (g179) & (g180) & (g181) & (g165) & (!g166)) + ((g178) & (g179) & (g180) & (g181) & (g165) & (g166)));
	assign g4015 = (((!g2177) & (!sk[120]) & (!g3777) & (g183)) + ((!g2177) & (!sk[120]) & (g3777) & (!g183)) + ((!g2177) & (!sk[120]) & (g3777) & (g183)) + ((!g2177) & (sk[120]) & (!g3777) & (g183)) + ((!g2177) & (sk[120]) & (g3777) & (g183)) + ((g2177) & (!sk[120]) & (!g3777) & (g183)) + ((g2177) & (!sk[120]) & (g3777) & (!g183)) + ((g2177) & (!sk[120]) & (g3777) & (g183)) + ((g2177) & (sk[120]) & (g3777) & (!g183)) + ((g2177) & (sk[120]) & (g3777) & (g183)));
	assign g4016 = (((!g2178) & (!sk[121]) & (!g3777) & (g184)) + ((!g2178) & (!sk[121]) & (g3777) & (!g184)) + ((!g2178) & (!sk[121]) & (g3777) & (g184)) + ((!g2178) & (sk[121]) & (!g3777) & (g184)) + ((!g2178) & (sk[121]) & (g3777) & (g184)) + ((g2178) & (!sk[121]) & (!g3777) & (g184)) + ((g2178) & (!sk[121]) & (g3777) & (!g184)) + ((g2178) & (!sk[121]) & (g3777) & (g184)) + ((g2178) & (sk[121]) & (g3777) & (!g184)) + ((g2178) & (sk[121]) & (g3777) & (g184)));
	assign g4017 = (((!g2179) & (!g3777) & (!sk[122]) & (g185)) + ((!g2179) & (!g3777) & (sk[122]) & (g185)) + ((!g2179) & (g3777) & (!sk[122]) & (!g185)) + ((!g2179) & (g3777) & (!sk[122]) & (g185)) + ((!g2179) & (g3777) & (sk[122]) & (g185)) + ((g2179) & (!g3777) & (!sk[122]) & (g185)) + ((g2179) & (g3777) & (!sk[122]) & (!g185)) + ((g2179) & (g3777) & (!sk[122]) & (g185)) + ((g2179) & (g3777) & (sk[122]) & (!g185)) + ((g2179) & (g3777) & (sk[122]) & (g185)));
	assign g186 = (((!g165) & (!g166) & (!g183) & (g184) & (!sk[123]) & (!g185)) + ((!g165) & (!g166) & (!g183) & (g184) & (!sk[123]) & (g185)) + ((!g165) & (!g166) & (g183) & (!g184) & (!sk[123]) & (!g185)) + ((!g165) & (!g166) & (g183) & (!g184) & (!sk[123]) & (g185)) + ((!g165) & (!g166) & (g183) & (g184) & (!sk[123]) & (!g185)) + ((!g165) & (!g166) & (g183) & (g184) & (!sk[123]) & (g185)) + ((!g165) & (g166) & (!g183) & (!g184) & (!sk[123]) & (!g185)) + ((!g165) & (g166) & (!g183) & (!g184) & (!sk[123]) & (g185)) + ((!g165) & (g166) & (!g183) & (!g184) & (sk[123]) & (g185)) + ((!g165) & (g166) & (!g183) & (g184) & (!sk[123]) & (!g185)) + ((!g165) & (g166) & (!g183) & (g184) & (!sk[123]) & (g185)) + ((!g165) & (g166) & (!g183) & (g184) & (sk[123]) & (g185)) + ((!g165) & (g166) & (g183) & (!g184) & (!sk[123]) & (!g185)) + ((!g165) & (g166) & (g183) & (!g184) & (!sk[123]) & (g185)) + ((!g165) & (g166) & (g183) & (!g184) & (sk[123]) & (g185)) + ((!g165) & (g166) & (g183) & (g184) & (!sk[123]) & (!g185)) + ((!g165) & (g166) & (g183) & (g184) & (!sk[123]) & (g185)) + ((!g165) & (g166) & (g183) & (g184) & (sk[123]) & (g185)) + ((g165) & (!g166) & (!g183) & (g184) & (!sk[123]) & (!g185)) + ((g165) & (!g166) & (!g183) & (g184) & (!sk[123]) & (g185)) + ((g165) & (!g166) & (g183) & (!g184) & (!sk[123]) & (!g185)) + ((g165) & (!g166) & (g183) & (!g184) & (!sk[123]) & (g185)) + ((g165) & (!g166) & (g183) & (!g184) & (sk[123]) & (!g185)) + ((g165) & (!g166) & (g183) & (!g184) & (sk[123]) & (g185)) + ((g165) & (!g166) & (g183) & (g184) & (!sk[123]) & (!g185)) + ((g165) & (!g166) & (g183) & (g184) & (!sk[123]) & (g185)) + ((g165) & (!g166) & (g183) & (g184) & (sk[123]) & (!g185)) + ((g165) & (!g166) & (g183) & (g184) & (sk[123]) & (g185)) + ((g165) & (g166) & (!g183) & (!g184) & (!sk[123]) & (!g185)) + ((g165) & (g166) & (!g183) & (!g184) & (!sk[123]) & (g185)) + ((g165) & (g166) & (!g183) & (g184) & (!sk[123]) & (!g185)) + ((g165) & (g166) & (!g183) & (g184) & (!sk[123]) & (g185)) + ((g165) & (g166) & (!g183) & (g184) & (sk[123]) & (!g185)) + ((g165) & (g166) & (!g183) & (g184) & (sk[123]) & (g185)) + ((g165) & (g166) & (g183) & (!g184) & (!sk[123]) & (!g185)) + ((g165) & (g166) & (g183) & (!g184) & (!sk[123]) & (g185)) + ((g165) & (g166) & (g183) & (g184) & (!sk[123]) & (!g185)) + ((g165) & (g166) & (g183) & (g184) & (!sk[123]) & (g185)) + ((g165) & (g166) & (g183) & (g184) & (sk[123]) & (!g185)) + ((g165) & (g166) & (g183) & (g184) & (sk[123]) & (g185)));
	assign g187 = (((!g147) & (!g148) & (!g172) & (!g177) & (!g182) & (g186)) + ((!g147) & (!g148) & (!g172) & (!g177) & (g182) & (g186)) + ((!g147) & (!g148) & (!g172) & (g177) & (!g182) & (g186)) + ((!g147) & (!g148) & (!g172) & (g177) & (g182) & (g186)) + ((!g147) & (!g148) & (g172) & (!g177) & (!g182) & (g186)) + ((!g147) & (!g148) & (g172) & (!g177) & (g182) & (g186)) + ((!g147) & (!g148) & (g172) & (g177) & (!g182) & (g186)) + ((!g147) & (!g148) & (g172) & (g177) & (g182) & (g186)) + ((!g147) & (g148) & (!g172) & (g177) & (!g182) & (!g186)) + ((!g147) & (g148) & (!g172) & (g177) & (!g182) & (g186)) + ((!g147) & (g148) & (!g172) & (g177) & (g182) & (!g186)) + ((!g147) & (g148) & (!g172) & (g177) & (g182) & (g186)) + ((!g147) & (g148) & (g172) & (g177) & (!g182) & (!g186)) + ((!g147) & (g148) & (g172) & (g177) & (!g182) & (g186)) + ((!g147) & (g148) & (g172) & (g177) & (g182) & (!g186)) + ((!g147) & (g148) & (g172) & (g177) & (g182) & (g186)) + ((g147) & (!g148) & (!g172) & (!g177) & (g182) & (!g186)) + ((g147) & (!g148) & (!g172) & (!g177) & (g182) & (g186)) + ((g147) & (!g148) & (!g172) & (g177) & (g182) & (!g186)) + ((g147) & (!g148) & (!g172) & (g177) & (g182) & (g186)) + ((g147) & (!g148) & (g172) & (!g177) & (g182) & (!g186)) + ((g147) & (!g148) & (g172) & (!g177) & (g182) & (g186)) + ((g147) & (!g148) & (g172) & (g177) & (g182) & (!g186)) + ((g147) & (!g148) & (g172) & (g177) & (g182) & (g186)) + ((g147) & (g148) & (g172) & (!g177) & (!g182) & (!g186)) + ((g147) & (g148) & (g172) & (!g177) & (!g182) & (g186)) + ((g147) & (g148) & (g172) & (!g177) & (g182) & (!g186)) + ((g147) & (g148) & (g172) & (!g177) & (g182) & (g186)) + ((g147) & (g148) & (g172) & (g177) & (!g182) & (!g186)) + ((g147) & (g148) & (g172) & (g177) & (!g182) & (g186)) + ((g147) & (g148) & (g172) & (g177) & (g182) & (!g186)) + ((g147) & (g148) & (g172) & (g177) & (g182) & (g186)));
	assign g188 = (((!g142) & (!g167) & (!sk[125]) & (g187)) + ((!g142) & (!g167) & (sk[125]) & (g187)) + ((!g142) & (g167) & (!sk[125]) & (!g187)) + ((!g142) & (g167) & (!sk[125]) & (g187)) + ((!g142) & (g167) & (sk[125]) & (g187)) + ((g142) & (!g167) & (!sk[125]) & (g187)) + ((g142) & (g167) & (!sk[125]) & (!g187)) + ((g142) & (g167) & (!sk[125]) & (g187)) + ((g142) & (g167) & (sk[125]) & (!g187)) + ((g142) & (g167) & (sk[125]) & (g187)));
	assign g4018 = (((!g2140) & (!g2210) & (!sk[126]) & (g189)) + ((!g2140) & (!g2210) & (sk[126]) & (g189)) + ((!g2140) & (g2210) & (!sk[126]) & (!g189)) + ((!g2140) & (g2210) & (!sk[126]) & (g189)) + ((!g2140) & (g2210) & (sk[126]) & (g189)) + ((g2140) & (!g2210) & (!sk[126]) & (g189)) + ((g2140) & (g2210) & (!sk[126]) & (!g189)) + ((g2140) & (g2210) & (!sk[126]) & (g189)) + ((g2140) & (g2210) & (sk[126]) & (!g189)) + ((g2140) & (g2210) & (sk[126]) & (g189)));
	assign g4019 = (((!g2146) & (!sk[127]) & (!g2210) & (g190)) + ((!g2146) & (!sk[127]) & (g2210) & (!g190)) + ((!g2146) & (!sk[127]) & (g2210) & (g190)) + ((!g2146) & (sk[127]) & (!g2210) & (g190)) + ((!g2146) & (sk[127]) & (g2210) & (g190)) + ((g2146) & (!sk[127]) & (!g2210) & (g190)) + ((g2146) & (!sk[127]) & (g2210) & (!g190)) + ((g2146) & (!sk[127]) & (g2210) & (g190)) + ((g2146) & (sk[127]) & (g2210) & (!g190)) + ((g2146) & (sk[127]) & (g2210) & (g190)));
	assign g4020 = (((!g2152) & (!sk[0]) & (!g2210) & (g191)) + ((!g2152) & (!sk[0]) & (g2210) & (!g191)) + ((!g2152) & (!sk[0]) & (g2210) & (g191)) + ((!g2152) & (sk[0]) & (!g2210) & (g191)) + ((!g2152) & (sk[0]) & (g2210) & (g191)) + ((g2152) & (!sk[0]) & (!g2210) & (g191)) + ((g2152) & (!sk[0]) & (g2210) & (!g191)) + ((g2152) & (!sk[0]) & (g2210) & (g191)) + ((g2152) & (sk[0]) & (g2210) & (!g191)) + ((g2152) & (sk[0]) & (g2210) & (g191)));
	assign g4021 = (((!sk[1]) & (!g2158) & (!g2210) & (g192)) + ((!sk[1]) & (!g2158) & (g2210) & (!g192)) + ((!sk[1]) & (!g2158) & (g2210) & (g192)) + ((!sk[1]) & (g2158) & (!g2210) & (g192)) + ((!sk[1]) & (g2158) & (g2210) & (!g192)) + ((!sk[1]) & (g2158) & (g2210) & (g192)) + ((sk[1]) & (!g2158) & (!g2210) & (g192)) + ((sk[1]) & (!g2158) & (g2210) & (g192)) + ((sk[1]) & (g2158) & (g2210) & (!g192)) + ((sk[1]) & (g2158) & (g2210) & (g192)));
	assign g193 = (((!g189) & (!g190) & (!g191) & (g192) & (g165) & (g166)) + ((!g189) & (!g190) & (g191) & (!g192) & (!g165) & (g166)) + ((!g189) & (!g190) & (g191) & (g192) & (!g165) & (g166)) + ((!g189) & (!g190) & (g191) & (g192) & (g165) & (g166)) + ((!g189) & (g190) & (!g191) & (!g192) & (g165) & (!g166)) + ((!g189) & (g190) & (!g191) & (g192) & (g165) & (!g166)) + ((!g189) & (g190) & (!g191) & (g192) & (g165) & (g166)) + ((!g189) & (g190) & (g191) & (!g192) & (!g165) & (g166)) + ((!g189) & (g190) & (g191) & (!g192) & (g165) & (!g166)) + ((!g189) & (g190) & (g191) & (g192) & (!g165) & (g166)) + ((!g189) & (g190) & (g191) & (g192) & (g165) & (!g166)) + ((!g189) & (g190) & (g191) & (g192) & (g165) & (g166)) + ((g189) & (!g190) & (!g191) & (!g192) & (!g165) & (!g166)) + ((g189) & (!g190) & (!g191) & (g192) & (!g165) & (!g166)) + ((g189) & (!g190) & (!g191) & (g192) & (g165) & (g166)) + ((g189) & (!g190) & (g191) & (!g192) & (!g165) & (!g166)) + ((g189) & (!g190) & (g191) & (!g192) & (!g165) & (g166)) + ((g189) & (!g190) & (g191) & (g192) & (!g165) & (!g166)) + ((g189) & (!g190) & (g191) & (g192) & (!g165) & (g166)) + ((g189) & (!g190) & (g191) & (g192) & (g165) & (g166)) + ((g189) & (g190) & (!g191) & (!g192) & (!g165) & (!g166)) + ((g189) & (g190) & (!g191) & (!g192) & (g165) & (!g166)) + ((g189) & (g190) & (!g191) & (g192) & (!g165) & (!g166)) + ((g189) & (g190) & (!g191) & (g192) & (g165) & (!g166)) + ((g189) & (g190) & (!g191) & (g192) & (g165) & (g166)) + ((g189) & (g190) & (g191) & (!g192) & (!g165) & (!g166)) + ((g189) & (g190) & (g191) & (!g192) & (!g165) & (g166)) + ((g189) & (g190) & (g191) & (!g192) & (g165) & (!g166)) + ((g189) & (g190) & (g191) & (g192) & (!g165) & (!g166)) + ((g189) & (g190) & (g191) & (g192) & (!g165) & (g166)) + ((g189) & (g190) & (g191) & (g192) & (g165) & (!g166)) + ((g189) & (g190) & (g191) & (g192) & (g165) & (g166)));
	assign g4022 = (((!sk[3]) & (!g2142) & (!g2210) & (g194)) + ((!sk[3]) & (!g2142) & (g2210) & (!g194)) + ((!sk[3]) & (!g2142) & (g2210) & (g194)) + ((!sk[3]) & (g2142) & (!g2210) & (g194)) + ((!sk[3]) & (g2142) & (g2210) & (!g194)) + ((!sk[3]) & (g2142) & (g2210) & (g194)) + ((sk[3]) & (!g2142) & (!g2210) & (g194)) + ((sk[3]) & (!g2142) & (g2210) & (g194)) + ((sk[3]) & (g2142) & (g2210) & (!g194)) + ((sk[3]) & (g2142) & (g2210) & (g194)));
	assign g4023 = (((!sk[4]) & (!g2148) & (!g2210) & (g195)) + ((!sk[4]) & (!g2148) & (g2210) & (!g195)) + ((!sk[4]) & (!g2148) & (g2210) & (g195)) + ((!sk[4]) & (g2148) & (!g2210) & (g195)) + ((!sk[4]) & (g2148) & (g2210) & (!g195)) + ((!sk[4]) & (g2148) & (g2210) & (g195)) + ((sk[4]) & (!g2148) & (!g2210) & (g195)) + ((sk[4]) & (!g2148) & (g2210) & (g195)) + ((sk[4]) & (g2148) & (g2210) & (!g195)) + ((sk[4]) & (g2148) & (g2210) & (g195)));
	assign g4024 = (((!sk[5]) & (!g2153) & (!g2210) & (g196)) + ((!sk[5]) & (!g2153) & (g2210) & (!g196)) + ((!sk[5]) & (!g2153) & (g2210) & (g196)) + ((!sk[5]) & (g2153) & (!g2210) & (g196)) + ((!sk[5]) & (g2153) & (g2210) & (!g196)) + ((!sk[5]) & (g2153) & (g2210) & (g196)) + ((sk[5]) & (!g2153) & (!g2210) & (g196)) + ((sk[5]) & (!g2153) & (g2210) & (g196)) + ((sk[5]) & (g2153) & (g2210) & (!g196)) + ((sk[5]) & (g2153) & (g2210) & (g196)));
	assign g4025 = (((!g2159) & (!sk[6]) & (!g2210) & (g197)) + ((!g2159) & (!sk[6]) & (g2210) & (!g197)) + ((!g2159) & (!sk[6]) & (g2210) & (g197)) + ((!g2159) & (sk[6]) & (!g2210) & (g197)) + ((!g2159) & (sk[6]) & (g2210) & (g197)) + ((g2159) & (!sk[6]) & (!g2210) & (g197)) + ((g2159) & (!sk[6]) & (g2210) & (!g197)) + ((g2159) & (!sk[6]) & (g2210) & (g197)) + ((g2159) & (sk[6]) & (g2210) & (!g197)) + ((g2159) & (sk[6]) & (g2210) & (g197)));
	assign g198 = (((!g194) & (!g195) & (!g196) & (g197) & (g165) & (g166)) + ((!g194) & (!g195) & (g196) & (!g197) & (!g165) & (g166)) + ((!g194) & (!g195) & (g196) & (g197) & (!g165) & (g166)) + ((!g194) & (!g195) & (g196) & (g197) & (g165) & (g166)) + ((!g194) & (g195) & (!g196) & (!g197) & (g165) & (!g166)) + ((!g194) & (g195) & (!g196) & (g197) & (g165) & (!g166)) + ((!g194) & (g195) & (!g196) & (g197) & (g165) & (g166)) + ((!g194) & (g195) & (g196) & (!g197) & (!g165) & (g166)) + ((!g194) & (g195) & (g196) & (!g197) & (g165) & (!g166)) + ((!g194) & (g195) & (g196) & (g197) & (!g165) & (g166)) + ((!g194) & (g195) & (g196) & (g197) & (g165) & (!g166)) + ((!g194) & (g195) & (g196) & (g197) & (g165) & (g166)) + ((g194) & (!g195) & (!g196) & (!g197) & (!g165) & (!g166)) + ((g194) & (!g195) & (!g196) & (g197) & (!g165) & (!g166)) + ((g194) & (!g195) & (!g196) & (g197) & (g165) & (g166)) + ((g194) & (!g195) & (g196) & (!g197) & (!g165) & (!g166)) + ((g194) & (!g195) & (g196) & (!g197) & (!g165) & (g166)) + ((g194) & (!g195) & (g196) & (g197) & (!g165) & (!g166)) + ((g194) & (!g195) & (g196) & (g197) & (!g165) & (g166)) + ((g194) & (!g195) & (g196) & (g197) & (g165) & (g166)) + ((g194) & (g195) & (!g196) & (!g197) & (!g165) & (!g166)) + ((g194) & (g195) & (!g196) & (!g197) & (g165) & (!g166)) + ((g194) & (g195) & (!g196) & (g197) & (!g165) & (!g166)) + ((g194) & (g195) & (!g196) & (g197) & (g165) & (!g166)) + ((g194) & (g195) & (!g196) & (g197) & (g165) & (g166)) + ((g194) & (g195) & (g196) & (!g197) & (!g165) & (!g166)) + ((g194) & (g195) & (g196) & (!g197) & (!g165) & (g166)) + ((g194) & (g195) & (g196) & (!g197) & (g165) & (!g166)) + ((g194) & (g195) & (g196) & (g197) & (!g165) & (!g166)) + ((g194) & (g195) & (g196) & (g197) & (!g165) & (g166)) + ((g194) & (g195) & (g196) & (g197) & (g165) & (!g166)) + ((g194) & (g195) & (g196) & (g197) & (g165) & (g166)));
	assign g4026 = (((!g2144) & (!g2210) & (!sk[8]) & (g199)) + ((!g2144) & (!g2210) & (sk[8]) & (g199)) + ((!g2144) & (g2210) & (!sk[8]) & (!g199)) + ((!g2144) & (g2210) & (!sk[8]) & (g199)) + ((!g2144) & (g2210) & (sk[8]) & (g199)) + ((g2144) & (!g2210) & (!sk[8]) & (g199)) + ((g2144) & (g2210) & (!sk[8]) & (!g199)) + ((g2144) & (g2210) & (!sk[8]) & (g199)) + ((g2144) & (g2210) & (sk[8]) & (!g199)) + ((g2144) & (g2210) & (sk[8]) & (g199)));
	assign g4027 = (((!sk[9]) & (!g2150) & (!g2210) & (g200)) + ((!sk[9]) & (!g2150) & (g2210) & (!g200)) + ((!sk[9]) & (!g2150) & (g2210) & (g200)) + ((!sk[9]) & (g2150) & (!g2210) & (g200)) + ((!sk[9]) & (g2150) & (g2210) & (!g200)) + ((!sk[9]) & (g2150) & (g2210) & (g200)) + ((sk[9]) & (!g2150) & (!g2210) & (g200)) + ((sk[9]) & (!g2150) & (g2210) & (g200)) + ((sk[9]) & (g2150) & (g2210) & (!g200)) + ((sk[9]) & (g2150) & (g2210) & (g200)));
	assign g4028 = (((!g2155) & (!g2210) & (!sk[10]) & (g201)) + ((!g2155) & (!g2210) & (sk[10]) & (g201)) + ((!g2155) & (g2210) & (!sk[10]) & (!g201)) + ((!g2155) & (g2210) & (!sk[10]) & (g201)) + ((!g2155) & (g2210) & (sk[10]) & (g201)) + ((g2155) & (!g2210) & (!sk[10]) & (g201)) + ((g2155) & (g2210) & (!sk[10]) & (!g201)) + ((g2155) & (g2210) & (!sk[10]) & (g201)) + ((g2155) & (g2210) & (sk[10]) & (!g201)) + ((g2155) & (g2210) & (sk[10]) & (g201)));
	assign g4029 = (((!g2160) & (!g2210) & (!sk[11]) & (g202)) + ((!g2160) & (!g2210) & (sk[11]) & (g202)) + ((!g2160) & (g2210) & (!sk[11]) & (!g202)) + ((!g2160) & (g2210) & (!sk[11]) & (g202)) + ((!g2160) & (g2210) & (sk[11]) & (g202)) + ((g2160) & (!g2210) & (!sk[11]) & (g202)) + ((g2160) & (g2210) & (!sk[11]) & (!g202)) + ((g2160) & (g2210) & (!sk[11]) & (g202)) + ((g2160) & (g2210) & (sk[11]) & (!g202)) + ((g2160) & (g2210) & (sk[11]) & (g202)));
	assign g203 = (((!g199) & (!g200) & (!g201) & (g202) & (g165) & (g166)) + ((!g199) & (!g200) & (g201) & (!g202) & (!g165) & (g166)) + ((!g199) & (!g200) & (g201) & (g202) & (!g165) & (g166)) + ((!g199) & (!g200) & (g201) & (g202) & (g165) & (g166)) + ((!g199) & (g200) & (!g201) & (!g202) & (g165) & (!g166)) + ((!g199) & (g200) & (!g201) & (g202) & (g165) & (!g166)) + ((!g199) & (g200) & (!g201) & (g202) & (g165) & (g166)) + ((!g199) & (g200) & (g201) & (!g202) & (!g165) & (g166)) + ((!g199) & (g200) & (g201) & (!g202) & (g165) & (!g166)) + ((!g199) & (g200) & (g201) & (g202) & (!g165) & (g166)) + ((!g199) & (g200) & (g201) & (g202) & (g165) & (!g166)) + ((!g199) & (g200) & (g201) & (g202) & (g165) & (g166)) + ((g199) & (!g200) & (!g201) & (!g202) & (!g165) & (!g166)) + ((g199) & (!g200) & (!g201) & (g202) & (!g165) & (!g166)) + ((g199) & (!g200) & (!g201) & (g202) & (g165) & (g166)) + ((g199) & (!g200) & (g201) & (!g202) & (!g165) & (!g166)) + ((g199) & (!g200) & (g201) & (!g202) & (!g165) & (g166)) + ((g199) & (!g200) & (g201) & (g202) & (!g165) & (!g166)) + ((g199) & (!g200) & (g201) & (g202) & (!g165) & (g166)) + ((g199) & (!g200) & (g201) & (g202) & (g165) & (g166)) + ((g199) & (g200) & (!g201) & (!g202) & (!g165) & (!g166)) + ((g199) & (g200) & (!g201) & (!g202) & (g165) & (!g166)) + ((g199) & (g200) & (!g201) & (g202) & (!g165) & (!g166)) + ((g199) & (g200) & (!g201) & (g202) & (g165) & (!g166)) + ((g199) & (g200) & (!g201) & (g202) & (g165) & (g166)) + ((g199) & (g200) & (g201) & (!g202) & (!g165) & (!g166)) + ((g199) & (g200) & (g201) & (!g202) & (!g165) & (g166)) + ((g199) & (g200) & (g201) & (!g202) & (g165) & (!g166)) + ((g199) & (g200) & (g201) & (g202) & (!g165) & (!g166)) + ((g199) & (g200) & (g201) & (g202) & (!g165) & (g166)) + ((g199) & (g200) & (g201) & (g202) & (g165) & (!g166)) + ((g199) & (g200) & (g201) & (g202) & (g165) & (g166)));
	assign g4030 = (((!sk[13]) & (!g2145) & (!g2210) & (g204)) + ((!sk[13]) & (!g2145) & (g2210) & (!g204)) + ((!sk[13]) & (!g2145) & (g2210) & (g204)) + ((!sk[13]) & (g2145) & (!g2210) & (g204)) + ((!sk[13]) & (g2145) & (g2210) & (!g204)) + ((!sk[13]) & (g2145) & (g2210) & (g204)) + ((sk[13]) & (!g2145) & (!g2210) & (g204)) + ((sk[13]) & (!g2145) & (g2210) & (g204)) + ((sk[13]) & (g2145) & (g2210) & (!g204)) + ((sk[13]) & (g2145) & (g2210) & (g204)));
	assign g4031 = (((!g2151) & (!sk[14]) & (!g2210) & (g205)) + ((!g2151) & (!sk[14]) & (g2210) & (!g205)) + ((!g2151) & (!sk[14]) & (g2210) & (g205)) + ((!g2151) & (sk[14]) & (!g2210) & (g205)) + ((!g2151) & (sk[14]) & (g2210) & (g205)) + ((g2151) & (!sk[14]) & (!g2210) & (g205)) + ((g2151) & (!sk[14]) & (g2210) & (!g205)) + ((g2151) & (!sk[14]) & (g2210) & (g205)) + ((g2151) & (sk[14]) & (g2210) & (!g205)) + ((g2151) & (sk[14]) & (g2210) & (g205)));
	assign g4032 = (((!g2157) & (!g2210) & (!sk[15]) & (g206)) + ((!g2157) & (!g2210) & (sk[15]) & (g206)) + ((!g2157) & (g2210) & (!sk[15]) & (!g206)) + ((!g2157) & (g2210) & (!sk[15]) & (g206)) + ((!g2157) & (g2210) & (sk[15]) & (g206)) + ((g2157) & (!g2210) & (!sk[15]) & (g206)) + ((g2157) & (g2210) & (!sk[15]) & (!g206)) + ((g2157) & (g2210) & (!sk[15]) & (g206)) + ((g2157) & (g2210) & (sk[15]) & (!g206)) + ((g2157) & (g2210) & (sk[15]) & (g206)));
	assign g4033 = (((!sk[16]) & (!g2161) & (!g2210) & (g207)) + ((!sk[16]) & (!g2161) & (g2210) & (!g207)) + ((!sk[16]) & (!g2161) & (g2210) & (g207)) + ((!sk[16]) & (g2161) & (!g2210) & (g207)) + ((!sk[16]) & (g2161) & (g2210) & (!g207)) + ((!sk[16]) & (g2161) & (g2210) & (g207)) + ((sk[16]) & (!g2161) & (!g2210) & (g207)) + ((sk[16]) & (!g2161) & (g2210) & (g207)) + ((sk[16]) & (g2161) & (g2210) & (!g207)) + ((sk[16]) & (g2161) & (g2210) & (g207)));
	assign g208 = (((!g204) & (!g205) & (!g206) & (g207) & (g165) & (g166)) + ((!g204) & (!g205) & (g206) & (!g207) & (!g165) & (g166)) + ((!g204) & (!g205) & (g206) & (g207) & (!g165) & (g166)) + ((!g204) & (!g205) & (g206) & (g207) & (g165) & (g166)) + ((!g204) & (g205) & (!g206) & (!g207) & (g165) & (!g166)) + ((!g204) & (g205) & (!g206) & (g207) & (g165) & (!g166)) + ((!g204) & (g205) & (!g206) & (g207) & (g165) & (g166)) + ((!g204) & (g205) & (g206) & (!g207) & (!g165) & (g166)) + ((!g204) & (g205) & (g206) & (!g207) & (g165) & (!g166)) + ((!g204) & (g205) & (g206) & (g207) & (!g165) & (g166)) + ((!g204) & (g205) & (g206) & (g207) & (g165) & (!g166)) + ((!g204) & (g205) & (g206) & (g207) & (g165) & (g166)) + ((g204) & (!g205) & (!g206) & (!g207) & (!g165) & (!g166)) + ((g204) & (!g205) & (!g206) & (g207) & (!g165) & (!g166)) + ((g204) & (!g205) & (!g206) & (g207) & (g165) & (g166)) + ((g204) & (!g205) & (g206) & (!g207) & (!g165) & (!g166)) + ((g204) & (!g205) & (g206) & (!g207) & (!g165) & (g166)) + ((g204) & (!g205) & (g206) & (g207) & (!g165) & (!g166)) + ((g204) & (!g205) & (g206) & (g207) & (!g165) & (g166)) + ((g204) & (!g205) & (g206) & (g207) & (g165) & (g166)) + ((g204) & (g205) & (!g206) & (!g207) & (!g165) & (!g166)) + ((g204) & (g205) & (!g206) & (!g207) & (g165) & (!g166)) + ((g204) & (g205) & (!g206) & (g207) & (!g165) & (!g166)) + ((g204) & (g205) & (!g206) & (g207) & (g165) & (!g166)) + ((g204) & (g205) & (!g206) & (g207) & (g165) & (g166)) + ((g204) & (g205) & (g206) & (!g207) & (!g165) & (!g166)) + ((g204) & (g205) & (g206) & (!g207) & (!g165) & (g166)) + ((g204) & (g205) & (g206) & (!g207) & (g165) & (!g166)) + ((g204) & (g205) & (g206) & (g207) & (!g165) & (!g166)) + ((g204) & (g205) & (g206) & (g207) & (!g165) & (g166)) + ((g204) & (g205) & (g206) & (g207) & (g165) & (!g166)) + ((g204) & (g205) & (g206) & (g207) & (g165) & (g166)));
	assign g209 = (((!g193) & (!g198) & (!g203) & (g208) & (g147) & (g148)) + ((!g193) & (!g198) & (g203) & (!g208) & (!g147) & (g148)) + ((!g193) & (!g198) & (g203) & (g208) & (!g147) & (g148)) + ((!g193) & (!g198) & (g203) & (g208) & (g147) & (g148)) + ((!g193) & (g198) & (!g203) & (!g208) & (g147) & (!g148)) + ((!g193) & (g198) & (!g203) & (g208) & (g147) & (!g148)) + ((!g193) & (g198) & (!g203) & (g208) & (g147) & (g148)) + ((!g193) & (g198) & (g203) & (!g208) & (!g147) & (g148)) + ((!g193) & (g198) & (g203) & (!g208) & (g147) & (!g148)) + ((!g193) & (g198) & (g203) & (g208) & (!g147) & (g148)) + ((!g193) & (g198) & (g203) & (g208) & (g147) & (!g148)) + ((!g193) & (g198) & (g203) & (g208) & (g147) & (g148)) + ((g193) & (!g198) & (!g203) & (!g208) & (!g147) & (!g148)) + ((g193) & (!g198) & (!g203) & (g208) & (!g147) & (!g148)) + ((g193) & (!g198) & (!g203) & (g208) & (g147) & (g148)) + ((g193) & (!g198) & (g203) & (!g208) & (!g147) & (!g148)) + ((g193) & (!g198) & (g203) & (!g208) & (!g147) & (g148)) + ((g193) & (!g198) & (g203) & (g208) & (!g147) & (!g148)) + ((g193) & (!g198) & (g203) & (g208) & (!g147) & (g148)) + ((g193) & (!g198) & (g203) & (g208) & (g147) & (g148)) + ((g193) & (g198) & (!g203) & (!g208) & (!g147) & (!g148)) + ((g193) & (g198) & (!g203) & (!g208) & (g147) & (!g148)) + ((g193) & (g198) & (!g203) & (g208) & (!g147) & (!g148)) + ((g193) & (g198) & (!g203) & (g208) & (g147) & (!g148)) + ((g193) & (g198) & (!g203) & (g208) & (g147) & (g148)) + ((g193) & (g198) & (g203) & (!g208) & (!g147) & (!g148)) + ((g193) & (g198) & (g203) & (!g208) & (!g147) & (g148)) + ((g193) & (g198) & (g203) & (!g208) & (g147) & (!g148)) + ((g193) & (g198) & (g203) & (g208) & (!g147) & (!g148)) + ((g193) & (g198) & (g203) & (g208) & (!g147) & (g148)) + ((g193) & (g198) & (g203) & (g208) & (g147) & (!g148)) + ((g193) & (g198) & (g203) & (g208) & (g147) & (g148)));
	assign g4034 = (((!g2162) & (!sk[19]) & (!g2210) & (g210)) + ((!g2162) & (!sk[19]) & (g2210) & (!g210)) + ((!g2162) & (!sk[19]) & (g2210) & (g210)) + ((!g2162) & (sk[19]) & (!g2210) & (g210)) + ((!g2162) & (sk[19]) & (g2210) & (g210)) + ((g2162) & (!sk[19]) & (!g2210) & (g210)) + ((g2162) & (!sk[19]) & (g2210) & (!g210)) + ((g2162) & (!sk[19]) & (g2210) & (g210)) + ((g2162) & (sk[19]) & (g2210) & (!g210)) + ((g2162) & (sk[19]) & (g2210) & (g210)));
	assign g4035 = (((!g2164) & (!g2210) & (!sk[20]) & (g211)) + ((!g2164) & (!g2210) & (sk[20]) & (g211)) + ((!g2164) & (g2210) & (!sk[20]) & (!g211)) + ((!g2164) & (g2210) & (!sk[20]) & (g211)) + ((!g2164) & (g2210) & (sk[20]) & (g211)) + ((g2164) & (!g2210) & (!sk[20]) & (g211)) + ((g2164) & (g2210) & (!sk[20]) & (!g211)) + ((g2164) & (g2210) & (!sk[20]) & (g211)) + ((g2164) & (g2210) & (sk[20]) & (!g211)) + ((g2164) & (g2210) & (sk[20]) & (g211)));
	assign g4036 = (((!g2166) & (!sk[21]) & (!g2210) & (g212)) + ((!g2166) & (!sk[21]) & (g2210) & (!g212)) + ((!g2166) & (!sk[21]) & (g2210) & (g212)) + ((!g2166) & (sk[21]) & (!g2210) & (g212)) + ((!g2166) & (sk[21]) & (g2210) & (g212)) + ((g2166) & (!sk[21]) & (!g2210) & (g212)) + ((g2166) & (!sk[21]) & (g2210) & (!g212)) + ((g2166) & (!sk[21]) & (g2210) & (g212)) + ((g2166) & (sk[21]) & (g2210) & (!g212)) + ((g2166) & (sk[21]) & (g2210) & (g212)));
	assign g4037 = (((!g2168) & (!sk[22]) & (!g2210) & (g213)) + ((!g2168) & (!sk[22]) & (g2210) & (!g213)) + ((!g2168) & (!sk[22]) & (g2210) & (g213)) + ((!g2168) & (sk[22]) & (!g2210) & (g213)) + ((!g2168) & (sk[22]) & (g2210) & (g213)) + ((g2168) & (!sk[22]) & (!g2210) & (g213)) + ((g2168) & (!sk[22]) & (g2210) & (!g213)) + ((g2168) & (!sk[22]) & (g2210) & (g213)) + ((g2168) & (sk[22]) & (g2210) & (!g213)) + ((g2168) & (sk[22]) & (g2210) & (g213)));
	assign g214 = (((!g210) & (!g211) & (!g212) & (g213) & (g165) & (g166)) + ((!g210) & (!g211) & (g212) & (!g213) & (!g165) & (g166)) + ((!g210) & (!g211) & (g212) & (g213) & (!g165) & (g166)) + ((!g210) & (!g211) & (g212) & (g213) & (g165) & (g166)) + ((!g210) & (g211) & (!g212) & (!g213) & (g165) & (!g166)) + ((!g210) & (g211) & (!g212) & (g213) & (g165) & (!g166)) + ((!g210) & (g211) & (!g212) & (g213) & (g165) & (g166)) + ((!g210) & (g211) & (g212) & (!g213) & (!g165) & (g166)) + ((!g210) & (g211) & (g212) & (!g213) & (g165) & (!g166)) + ((!g210) & (g211) & (g212) & (g213) & (!g165) & (g166)) + ((!g210) & (g211) & (g212) & (g213) & (g165) & (!g166)) + ((!g210) & (g211) & (g212) & (g213) & (g165) & (g166)) + ((g210) & (!g211) & (!g212) & (!g213) & (!g165) & (!g166)) + ((g210) & (!g211) & (!g212) & (g213) & (!g165) & (!g166)) + ((g210) & (!g211) & (!g212) & (g213) & (g165) & (g166)) + ((g210) & (!g211) & (g212) & (!g213) & (!g165) & (!g166)) + ((g210) & (!g211) & (g212) & (!g213) & (!g165) & (g166)) + ((g210) & (!g211) & (g212) & (g213) & (!g165) & (!g166)) + ((g210) & (!g211) & (g212) & (g213) & (!g165) & (g166)) + ((g210) & (!g211) & (g212) & (g213) & (g165) & (g166)) + ((g210) & (g211) & (!g212) & (!g213) & (!g165) & (!g166)) + ((g210) & (g211) & (!g212) & (!g213) & (g165) & (!g166)) + ((g210) & (g211) & (!g212) & (g213) & (!g165) & (!g166)) + ((g210) & (g211) & (!g212) & (g213) & (g165) & (!g166)) + ((g210) & (g211) & (!g212) & (g213) & (g165) & (g166)) + ((g210) & (g211) & (g212) & (!g213) & (!g165) & (!g166)) + ((g210) & (g211) & (g212) & (!g213) & (!g165) & (g166)) + ((g210) & (g211) & (g212) & (!g213) & (g165) & (!g166)) + ((g210) & (g211) & (g212) & (g213) & (!g165) & (!g166)) + ((g210) & (g211) & (g212) & (g213) & (!g165) & (g166)) + ((g210) & (g211) & (g212) & (g213) & (g165) & (!g166)) + ((g210) & (g211) & (g212) & (g213) & (g165) & (g166)));
	assign g4038 = (((!g2169) & (!g2210) & (!sk[24]) & (g215)) + ((!g2169) & (!g2210) & (sk[24]) & (g215)) + ((!g2169) & (g2210) & (!sk[24]) & (!g215)) + ((!g2169) & (g2210) & (!sk[24]) & (g215)) + ((!g2169) & (g2210) & (sk[24]) & (g215)) + ((g2169) & (!g2210) & (!sk[24]) & (g215)) + ((g2169) & (g2210) & (!sk[24]) & (!g215)) + ((g2169) & (g2210) & (!sk[24]) & (g215)) + ((g2169) & (g2210) & (sk[24]) & (!g215)) + ((g2169) & (g2210) & (sk[24]) & (g215)));
	assign g4039 = (((!g2170) & (!sk[25]) & (!g2210) & (g216)) + ((!g2170) & (!sk[25]) & (g2210) & (!g216)) + ((!g2170) & (!sk[25]) & (g2210) & (g216)) + ((!g2170) & (sk[25]) & (!g2210) & (g216)) + ((!g2170) & (sk[25]) & (g2210) & (g216)) + ((g2170) & (!sk[25]) & (!g2210) & (g216)) + ((g2170) & (!sk[25]) & (g2210) & (!g216)) + ((g2170) & (!sk[25]) & (g2210) & (g216)) + ((g2170) & (sk[25]) & (g2210) & (!g216)) + ((g2170) & (sk[25]) & (g2210) & (g216)));
	assign g4040 = (((!sk[26]) & (!g2171) & (!g2210) & (g217)) + ((!sk[26]) & (!g2171) & (g2210) & (!g217)) + ((!sk[26]) & (!g2171) & (g2210) & (g217)) + ((!sk[26]) & (g2171) & (!g2210) & (g217)) + ((!sk[26]) & (g2171) & (g2210) & (!g217)) + ((!sk[26]) & (g2171) & (g2210) & (g217)) + ((sk[26]) & (!g2171) & (!g2210) & (g217)) + ((sk[26]) & (!g2171) & (g2210) & (g217)) + ((sk[26]) & (g2171) & (g2210) & (!g217)) + ((sk[26]) & (g2171) & (g2210) & (g217)));
	assign g4041 = (((!g2172) & (!sk[27]) & (!g2210) & (g218)) + ((!g2172) & (!sk[27]) & (g2210) & (!g218)) + ((!g2172) & (!sk[27]) & (g2210) & (g218)) + ((!g2172) & (sk[27]) & (!g2210) & (g218)) + ((!g2172) & (sk[27]) & (g2210) & (g218)) + ((g2172) & (!sk[27]) & (!g2210) & (g218)) + ((g2172) & (!sk[27]) & (g2210) & (!g218)) + ((g2172) & (!sk[27]) & (g2210) & (g218)) + ((g2172) & (sk[27]) & (g2210) & (!g218)) + ((g2172) & (sk[27]) & (g2210) & (g218)));
	assign g219 = (((!g215) & (!g216) & (!g217) & (g218) & (g165) & (g166)) + ((!g215) & (!g216) & (g217) & (!g218) & (!g165) & (g166)) + ((!g215) & (!g216) & (g217) & (g218) & (!g165) & (g166)) + ((!g215) & (!g216) & (g217) & (g218) & (g165) & (g166)) + ((!g215) & (g216) & (!g217) & (!g218) & (g165) & (!g166)) + ((!g215) & (g216) & (!g217) & (g218) & (g165) & (!g166)) + ((!g215) & (g216) & (!g217) & (g218) & (g165) & (g166)) + ((!g215) & (g216) & (g217) & (!g218) & (!g165) & (g166)) + ((!g215) & (g216) & (g217) & (!g218) & (g165) & (!g166)) + ((!g215) & (g216) & (g217) & (g218) & (!g165) & (g166)) + ((!g215) & (g216) & (g217) & (g218) & (g165) & (!g166)) + ((!g215) & (g216) & (g217) & (g218) & (g165) & (g166)) + ((g215) & (!g216) & (!g217) & (!g218) & (!g165) & (!g166)) + ((g215) & (!g216) & (!g217) & (g218) & (!g165) & (!g166)) + ((g215) & (!g216) & (!g217) & (g218) & (g165) & (g166)) + ((g215) & (!g216) & (g217) & (!g218) & (!g165) & (!g166)) + ((g215) & (!g216) & (g217) & (!g218) & (!g165) & (g166)) + ((g215) & (!g216) & (g217) & (g218) & (!g165) & (!g166)) + ((g215) & (!g216) & (g217) & (g218) & (!g165) & (g166)) + ((g215) & (!g216) & (g217) & (g218) & (g165) & (g166)) + ((g215) & (g216) & (!g217) & (!g218) & (!g165) & (!g166)) + ((g215) & (g216) & (!g217) & (!g218) & (g165) & (!g166)) + ((g215) & (g216) & (!g217) & (g218) & (!g165) & (!g166)) + ((g215) & (g216) & (!g217) & (g218) & (g165) & (!g166)) + ((g215) & (g216) & (!g217) & (g218) & (g165) & (g166)) + ((g215) & (g216) & (g217) & (!g218) & (!g165) & (!g166)) + ((g215) & (g216) & (g217) & (!g218) & (!g165) & (g166)) + ((g215) & (g216) & (g217) & (!g218) & (g165) & (!g166)) + ((g215) & (g216) & (g217) & (g218) & (!g165) & (!g166)) + ((g215) & (g216) & (g217) & (g218) & (!g165) & (g166)) + ((g215) & (g216) & (g217) & (g218) & (g165) & (!g166)) + ((g215) & (g216) & (g217) & (g218) & (g165) & (g166)));
	assign g4042 = (((!g2173) & (!g2210) & (!sk[29]) & (g220)) + ((!g2173) & (!g2210) & (sk[29]) & (g220)) + ((!g2173) & (g2210) & (!sk[29]) & (!g220)) + ((!g2173) & (g2210) & (!sk[29]) & (g220)) + ((!g2173) & (g2210) & (sk[29]) & (g220)) + ((g2173) & (!g2210) & (!sk[29]) & (g220)) + ((g2173) & (g2210) & (!sk[29]) & (!g220)) + ((g2173) & (g2210) & (!sk[29]) & (g220)) + ((g2173) & (g2210) & (sk[29]) & (!g220)) + ((g2173) & (g2210) & (sk[29]) & (g220)));
	assign g4043 = (((!g2174) & (!sk[30]) & (!g2210) & (g221)) + ((!g2174) & (!sk[30]) & (g2210) & (!g221)) + ((!g2174) & (!sk[30]) & (g2210) & (g221)) + ((!g2174) & (sk[30]) & (!g2210) & (g221)) + ((!g2174) & (sk[30]) & (g2210) & (g221)) + ((g2174) & (!sk[30]) & (!g2210) & (g221)) + ((g2174) & (!sk[30]) & (g2210) & (!g221)) + ((g2174) & (!sk[30]) & (g2210) & (g221)) + ((g2174) & (sk[30]) & (g2210) & (!g221)) + ((g2174) & (sk[30]) & (g2210) & (g221)));
	assign g4044 = (((!g2175) & (!sk[31]) & (!g2210) & (g222)) + ((!g2175) & (!sk[31]) & (g2210) & (!g222)) + ((!g2175) & (!sk[31]) & (g2210) & (g222)) + ((!g2175) & (sk[31]) & (!g2210) & (g222)) + ((!g2175) & (sk[31]) & (g2210) & (g222)) + ((g2175) & (!sk[31]) & (!g2210) & (g222)) + ((g2175) & (!sk[31]) & (g2210) & (!g222)) + ((g2175) & (!sk[31]) & (g2210) & (g222)) + ((g2175) & (sk[31]) & (g2210) & (!g222)) + ((g2175) & (sk[31]) & (g2210) & (g222)));
	assign g4045 = (((!sk[32]) & (!g2176) & (!g2210) & (g223)) + ((!sk[32]) & (!g2176) & (g2210) & (!g223)) + ((!sk[32]) & (!g2176) & (g2210) & (g223)) + ((!sk[32]) & (g2176) & (!g2210) & (g223)) + ((!sk[32]) & (g2176) & (g2210) & (!g223)) + ((!sk[32]) & (g2176) & (g2210) & (g223)) + ((sk[32]) & (!g2176) & (!g2210) & (g223)) + ((sk[32]) & (!g2176) & (g2210) & (g223)) + ((sk[32]) & (g2176) & (g2210) & (!g223)) + ((sk[32]) & (g2176) & (g2210) & (g223)));
	assign g224 = (((!g220) & (!g221) & (!g222) & (g223) & (g165) & (g166)) + ((!g220) & (!g221) & (g222) & (!g223) & (!g165) & (g166)) + ((!g220) & (!g221) & (g222) & (g223) & (!g165) & (g166)) + ((!g220) & (!g221) & (g222) & (g223) & (g165) & (g166)) + ((!g220) & (g221) & (!g222) & (!g223) & (g165) & (!g166)) + ((!g220) & (g221) & (!g222) & (g223) & (g165) & (!g166)) + ((!g220) & (g221) & (!g222) & (g223) & (g165) & (g166)) + ((!g220) & (g221) & (g222) & (!g223) & (!g165) & (g166)) + ((!g220) & (g221) & (g222) & (!g223) & (g165) & (!g166)) + ((!g220) & (g221) & (g222) & (g223) & (!g165) & (g166)) + ((!g220) & (g221) & (g222) & (g223) & (g165) & (!g166)) + ((!g220) & (g221) & (g222) & (g223) & (g165) & (g166)) + ((g220) & (!g221) & (!g222) & (!g223) & (!g165) & (!g166)) + ((g220) & (!g221) & (!g222) & (g223) & (!g165) & (!g166)) + ((g220) & (!g221) & (!g222) & (g223) & (g165) & (g166)) + ((g220) & (!g221) & (g222) & (!g223) & (!g165) & (!g166)) + ((g220) & (!g221) & (g222) & (!g223) & (!g165) & (g166)) + ((g220) & (!g221) & (g222) & (g223) & (!g165) & (!g166)) + ((g220) & (!g221) & (g222) & (g223) & (!g165) & (g166)) + ((g220) & (!g221) & (g222) & (g223) & (g165) & (g166)) + ((g220) & (g221) & (!g222) & (!g223) & (!g165) & (!g166)) + ((g220) & (g221) & (!g222) & (!g223) & (g165) & (!g166)) + ((g220) & (g221) & (!g222) & (g223) & (!g165) & (!g166)) + ((g220) & (g221) & (!g222) & (g223) & (g165) & (!g166)) + ((g220) & (g221) & (!g222) & (g223) & (g165) & (g166)) + ((g220) & (g221) & (g222) & (!g223) & (!g165) & (!g166)) + ((g220) & (g221) & (g222) & (!g223) & (!g165) & (g166)) + ((g220) & (g221) & (g222) & (!g223) & (g165) & (!g166)) + ((g220) & (g221) & (g222) & (g223) & (!g165) & (!g166)) + ((g220) & (g221) & (g222) & (g223) & (!g165) & (g166)) + ((g220) & (g221) & (g222) & (g223) & (g165) & (!g166)) + ((g220) & (g221) & (g222) & (g223) & (g165) & (g166)));
	assign g4046 = (((!g2177) & (!g2210) & (!sk[34]) & (g225)) + ((!g2177) & (!g2210) & (sk[34]) & (g225)) + ((!g2177) & (g2210) & (!sk[34]) & (!g225)) + ((!g2177) & (g2210) & (!sk[34]) & (g225)) + ((!g2177) & (g2210) & (sk[34]) & (g225)) + ((g2177) & (!g2210) & (!sk[34]) & (g225)) + ((g2177) & (g2210) & (!sk[34]) & (!g225)) + ((g2177) & (g2210) & (!sk[34]) & (g225)) + ((g2177) & (g2210) & (sk[34]) & (!g225)) + ((g2177) & (g2210) & (sk[34]) & (g225)));
	assign g4047 = (((!sk[35]) & (!g2178) & (!g2210) & (g226)) + ((!sk[35]) & (!g2178) & (g2210) & (!g226)) + ((!sk[35]) & (!g2178) & (g2210) & (g226)) + ((!sk[35]) & (g2178) & (!g2210) & (g226)) + ((!sk[35]) & (g2178) & (g2210) & (!g226)) + ((!sk[35]) & (g2178) & (g2210) & (g226)) + ((sk[35]) & (!g2178) & (!g2210) & (g226)) + ((sk[35]) & (!g2178) & (g2210) & (g226)) + ((sk[35]) & (g2178) & (g2210) & (!g226)) + ((sk[35]) & (g2178) & (g2210) & (g226)));
	assign g4048 = (((!sk[36]) & (!g2179) & (!g2210) & (g227)) + ((!sk[36]) & (!g2179) & (g2210) & (!g227)) + ((!sk[36]) & (!g2179) & (g2210) & (g227)) + ((!sk[36]) & (g2179) & (!g2210) & (g227)) + ((!sk[36]) & (g2179) & (g2210) & (!g227)) + ((!sk[36]) & (g2179) & (g2210) & (g227)) + ((sk[36]) & (!g2179) & (!g2210) & (g227)) + ((sk[36]) & (!g2179) & (g2210) & (g227)) + ((sk[36]) & (g2179) & (g2210) & (!g227)) + ((sk[36]) & (g2179) & (g2210) & (g227)));
	assign g228 = (((!g165) & (!sk[37]) & (!g166) & (!g225) & (g226) & (!g227)) + ((!g165) & (!sk[37]) & (!g166) & (!g225) & (g226) & (g227)) + ((!g165) & (!sk[37]) & (!g166) & (g225) & (!g226) & (!g227)) + ((!g165) & (!sk[37]) & (!g166) & (g225) & (!g226) & (g227)) + ((!g165) & (!sk[37]) & (!g166) & (g225) & (g226) & (!g227)) + ((!g165) & (!sk[37]) & (!g166) & (g225) & (g226) & (g227)) + ((!g165) & (!sk[37]) & (g166) & (!g225) & (!g226) & (!g227)) + ((!g165) & (!sk[37]) & (g166) & (!g225) & (!g226) & (g227)) + ((!g165) & (!sk[37]) & (g166) & (!g225) & (g226) & (!g227)) + ((!g165) & (!sk[37]) & (g166) & (!g225) & (g226) & (g227)) + ((!g165) & (!sk[37]) & (g166) & (g225) & (!g226) & (!g227)) + ((!g165) & (!sk[37]) & (g166) & (g225) & (!g226) & (g227)) + ((!g165) & (!sk[37]) & (g166) & (g225) & (g226) & (!g227)) + ((!g165) & (!sk[37]) & (g166) & (g225) & (g226) & (g227)) + ((!g165) & (sk[37]) & (g166) & (!g225) & (!g226) & (g227)) + ((!g165) & (sk[37]) & (g166) & (!g225) & (g226) & (g227)) + ((!g165) & (sk[37]) & (g166) & (g225) & (!g226) & (g227)) + ((!g165) & (sk[37]) & (g166) & (g225) & (g226) & (g227)) + ((g165) & (!sk[37]) & (!g166) & (!g225) & (g226) & (!g227)) + ((g165) & (!sk[37]) & (!g166) & (!g225) & (g226) & (g227)) + ((g165) & (!sk[37]) & (!g166) & (g225) & (!g226) & (!g227)) + ((g165) & (!sk[37]) & (!g166) & (g225) & (!g226) & (g227)) + ((g165) & (!sk[37]) & (!g166) & (g225) & (g226) & (!g227)) + ((g165) & (!sk[37]) & (!g166) & (g225) & (g226) & (g227)) + ((g165) & (!sk[37]) & (g166) & (!g225) & (!g226) & (!g227)) + ((g165) & (!sk[37]) & (g166) & (!g225) & (!g226) & (g227)) + ((g165) & (!sk[37]) & (g166) & (!g225) & (g226) & (!g227)) + ((g165) & (!sk[37]) & (g166) & (!g225) & (g226) & (g227)) + ((g165) & (!sk[37]) & (g166) & (g225) & (!g226) & (!g227)) + ((g165) & (!sk[37]) & (g166) & (g225) & (!g226) & (g227)) + ((g165) & (!sk[37]) & (g166) & (g225) & (g226) & (!g227)) + ((g165) & (!sk[37]) & (g166) & (g225) & (g226) & (g227)) + ((g165) & (sk[37]) & (!g166) & (g225) & (!g226) & (!g227)) + ((g165) & (sk[37]) & (!g166) & (g225) & (!g226) & (g227)) + ((g165) & (sk[37]) & (!g166) & (g225) & (g226) & (!g227)) + ((g165) & (sk[37]) & (!g166) & (g225) & (g226) & (g227)) + ((g165) & (sk[37]) & (g166) & (!g225) & (g226) & (!g227)) + ((g165) & (sk[37]) & (g166) & (!g225) & (g226) & (g227)) + ((g165) & (sk[37]) & (g166) & (g225) & (g226) & (!g227)) + ((g165) & (sk[37]) & (g166) & (g225) & (g226) & (g227)));
	assign g229 = (((!g147) & (!g148) & (!g214) & (!g219) & (!g224) & (g228)) + ((!g147) & (!g148) & (!g214) & (!g219) & (g224) & (g228)) + ((!g147) & (!g148) & (!g214) & (g219) & (!g224) & (g228)) + ((!g147) & (!g148) & (!g214) & (g219) & (g224) & (g228)) + ((!g147) & (!g148) & (g214) & (!g219) & (!g224) & (g228)) + ((!g147) & (!g148) & (g214) & (!g219) & (g224) & (g228)) + ((!g147) & (!g148) & (g214) & (g219) & (!g224) & (g228)) + ((!g147) & (!g148) & (g214) & (g219) & (g224) & (g228)) + ((!g147) & (g148) & (!g214) & (g219) & (!g224) & (!g228)) + ((!g147) & (g148) & (!g214) & (g219) & (!g224) & (g228)) + ((!g147) & (g148) & (!g214) & (g219) & (g224) & (!g228)) + ((!g147) & (g148) & (!g214) & (g219) & (g224) & (g228)) + ((!g147) & (g148) & (g214) & (g219) & (!g224) & (!g228)) + ((!g147) & (g148) & (g214) & (g219) & (!g224) & (g228)) + ((!g147) & (g148) & (g214) & (g219) & (g224) & (!g228)) + ((!g147) & (g148) & (g214) & (g219) & (g224) & (g228)) + ((g147) & (!g148) & (!g214) & (!g219) & (g224) & (!g228)) + ((g147) & (!g148) & (!g214) & (!g219) & (g224) & (g228)) + ((g147) & (!g148) & (!g214) & (g219) & (g224) & (!g228)) + ((g147) & (!g148) & (!g214) & (g219) & (g224) & (g228)) + ((g147) & (!g148) & (g214) & (!g219) & (g224) & (!g228)) + ((g147) & (!g148) & (g214) & (!g219) & (g224) & (g228)) + ((g147) & (!g148) & (g214) & (g219) & (g224) & (!g228)) + ((g147) & (!g148) & (g214) & (g219) & (g224) & (g228)) + ((g147) & (g148) & (g214) & (!g219) & (!g224) & (!g228)) + ((g147) & (g148) & (g214) & (!g219) & (!g224) & (g228)) + ((g147) & (g148) & (g214) & (!g219) & (g224) & (!g228)) + ((g147) & (g148) & (g214) & (!g219) & (g224) & (g228)) + ((g147) & (g148) & (g214) & (g219) & (!g224) & (!g228)) + ((g147) & (g148) & (g214) & (g219) & (!g224) & (g228)) + ((g147) & (g148) & (g214) & (g219) & (g224) & (!g228)) + ((g147) & (g148) & (g214) & (g219) & (g224) & (g228)));
	assign g230 = (((!sk[39]) & (!g142) & (!g209) & (g229)) + ((!sk[39]) & (!g142) & (g209) & (!g229)) + ((!sk[39]) & (!g142) & (g209) & (g229)) + ((!sk[39]) & (g142) & (!g209) & (g229)) + ((!sk[39]) & (g142) & (g209) & (!g229)) + ((!sk[39]) & (g142) & (g209) & (g229)) + ((sk[39]) & (!g142) & (!g209) & (g229)) + ((sk[39]) & (!g142) & (g209) & (g229)) + ((sk[39]) & (g142) & (g209) & (!g229)) + ((sk[39]) & (g142) & (g209) & (g229)));
	assign g231 = (((!g88) & (!g89) & (!g188) & (!sk[40]) & (g230)) + ((!g88) & (!g89) & (g188) & (!sk[40]) & (!g230)) + ((!g88) & (!g89) & (g188) & (!sk[40]) & (g230)) + ((!g88) & (g89) & (!g188) & (!sk[40]) & (!g230)) + ((!g88) & (g89) & (!g188) & (!sk[40]) & (g230)) + ((!g88) & (g89) & (g188) & (!sk[40]) & (!g230)) + ((!g88) & (g89) & (g188) & (!sk[40]) & (g230)) + ((!g88) & (g89) & (g188) & (sk[40]) & (g230)) + ((g88) & (!g89) & (!g188) & (!sk[40]) & (g230)) + ((g88) & (!g89) & (!g188) & (sk[40]) & (g230)) + ((g88) & (!g89) & (g188) & (!sk[40]) & (!g230)) + ((g88) & (!g89) & (g188) & (!sk[40]) & (g230)) + ((g88) & (!g89) & (g188) & (sk[40]) & (g230)) + ((g88) & (g89) & (!g188) & (!sk[40]) & (!g230)) + ((g88) & (g89) & (!g188) & (!sk[40]) & (g230)) + ((g88) & (g89) & (!g188) & (sk[40]) & (g230)) + ((g88) & (g89) & (g188) & (!sk[40]) & (!g230)) + ((g88) & (g89) & (g188) & (!sk[40]) & (g230)) + ((g88) & (g89) & (g188) & (sk[40]) & (!g230)) + ((g88) & (g89) & (g188) & (sk[40]) & (g230)));
	assign g4049 = (((!g2140) & (!sk[41]) & (!g2229) & (g232)) + ((!g2140) & (!sk[41]) & (g2229) & (!g232)) + ((!g2140) & (!sk[41]) & (g2229) & (g232)) + ((!g2140) & (sk[41]) & (!g2229) & (g232)) + ((!g2140) & (sk[41]) & (g2229) & (g232)) + ((g2140) & (!sk[41]) & (!g2229) & (g232)) + ((g2140) & (!sk[41]) & (g2229) & (!g232)) + ((g2140) & (!sk[41]) & (g2229) & (g232)) + ((g2140) & (sk[41]) & (g2229) & (!g232)) + ((g2140) & (sk[41]) & (g2229) & (g232)));
	assign g4050 = (((!g2142) & (!sk[42]) & (!g2229) & (g233)) + ((!g2142) & (!sk[42]) & (g2229) & (!g233)) + ((!g2142) & (!sk[42]) & (g2229) & (g233)) + ((!g2142) & (sk[42]) & (!g2229) & (g233)) + ((!g2142) & (sk[42]) & (g2229) & (g233)) + ((g2142) & (!sk[42]) & (!g2229) & (g233)) + ((g2142) & (!sk[42]) & (g2229) & (!g233)) + ((g2142) & (!sk[42]) & (g2229) & (g233)) + ((g2142) & (sk[42]) & (g2229) & (!g233)) + ((g2142) & (sk[42]) & (g2229) & (g233)));
	assign g4051 = (((!g2144) & (!sk[43]) & (!g2229) & (g234)) + ((!g2144) & (!sk[43]) & (g2229) & (!g234)) + ((!g2144) & (!sk[43]) & (g2229) & (g234)) + ((!g2144) & (sk[43]) & (!g2229) & (g234)) + ((!g2144) & (sk[43]) & (g2229) & (g234)) + ((g2144) & (!sk[43]) & (!g2229) & (g234)) + ((g2144) & (!sk[43]) & (g2229) & (!g234)) + ((g2144) & (!sk[43]) & (g2229) & (g234)) + ((g2144) & (sk[43]) & (g2229) & (!g234)) + ((g2144) & (sk[43]) & (g2229) & (g234)));
	assign g4052 = (((!g2145) & (!g2229) & (!sk[44]) & (g235)) + ((!g2145) & (!g2229) & (sk[44]) & (g235)) + ((!g2145) & (g2229) & (!sk[44]) & (!g235)) + ((!g2145) & (g2229) & (!sk[44]) & (g235)) + ((!g2145) & (g2229) & (sk[44]) & (g235)) + ((g2145) & (!g2229) & (!sk[44]) & (g235)) + ((g2145) & (g2229) & (!sk[44]) & (!g235)) + ((g2145) & (g2229) & (!sk[44]) & (g235)) + ((g2145) & (g2229) & (sk[44]) & (!g235)) + ((g2145) & (g2229) & (sk[44]) & (g235)));
	assign g236 = (((!g232) & (!g233) & (!g234) & (g235) & (g147) & (g148)) + ((!g232) & (!g233) & (g234) & (!g235) & (!g147) & (g148)) + ((!g232) & (!g233) & (g234) & (g235) & (!g147) & (g148)) + ((!g232) & (!g233) & (g234) & (g235) & (g147) & (g148)) + ((!g232) & (g233) & (!g234) & (!g235) & (g147) & (!g148)) + ((!g232) & (g233) & (!g234) & (g235) & (g147) & (!g148)) + ((!g232) & (g233) & (!g234) & (g235) & (g147) & (g148)) + ((!g232) & (g233) & (g234) & (!g235) & (!g147) & (g148)) + ((!g232) & (g233) & (g234) & (!g235) & (g147) & (!g148)) + ((!g232) & (g233) & (g234) & (g235) & (!g147) & (g148)) + ((!g232) & (g233) & (g234) & (g235) & (g147) & (!g148)) + ((!g232) & (g233) & (g234) & (g235) & (g147) & (g148)) + ((g232) & (!g233) & (!g234) & (!g235) & (!g147) & (!g148)) + ((g232) & (!g233) & (!g234) & (g235) & (!g147) & (!g148)) + ((g232) & (!g233) & (!g234) & (g235) & (g147) & (g148)) + ((g232) & (!g233) & (g234) & (!g235) & (!g147) & (!g148)) + ((g232) & (!g233) & (g234) & (!g235) & (!g147) & (g148)) + ((g232) & (!g233) & (g234) & (g235) & (!g147) & (!g148)) + ((g232) & (!g233) & (g234) & (g235) & (!g147) & (g148)) + ((g232) & (!g233) & (g234) & (g235) & (g147) & (g148)) + ((g232) & (g233) & (!g234) & (!g235) & (!g147) & (!g148)) + ((g232) & (g233) & (!g234) & (!g235) & (g147) & (!g148)) + ((g232) & (g233) & (!g234) & (g235) & (!g147) & (!g148)) + ((g232) & (g233) & (!g234) & (g235) & (g147) & (!g148)) + ((g232) & (g233) & (!g234) & (g235) & (g147) & (g148)) + ((g232) & (g233) & (g234) & (!g235) & (!g147) & (!g148)) + ((g232) & (g233) & (g234) & (!g235) & (!g147) & (g148)) + ((g232) & (g233) & (g234) & (!g235) & (g147) & (!g148)) + ((g232) & (g233) & (g234) & (g235) & (!g147) & (!g148)) + ((g232) & (g233) & (g234) & (g235) & (!g147) & (g148)) + ((g232) & (g233) & (g234) & (g235) & (g147) & (!g148)) + ((g232) & (g233) & (g234) & (g235) & (g147) & (g148)));
	assign g4053 = (((!g2146) & (!g2229) & (!sk[46]) & (g237)) + ((!g2146) & (!g2229) & (sk[46]) & (g237)) + ((!g2146) & (g2229) & (!sk[46]) & (!g237)) + ((!g2146) & (g2229) & (!sk[46]) & (g237)) + ((!g2146) & (g2229) & (sk[46]) & (g237)) + ((g2146) & (!g2229) & (!sk[46]) & (g237)) + ((g2146) & (g2229) & (!sk[46]) & (!g237)) + ((g2146) & (g2229) & (!sk[46]) & (g237)) + ((g2146) & (g2229) & (sk[46]) & (!g237)) + ((g2146) & (g2229) & (sk[46]) & (g237)));
	assign g4054 = (((!g2148) & (!sk[47]) & (!g2229) & (g238)) + ((!g2148) & (!sk[47]) & (g2229) & (!g238)) + ((!g2148) & (!sk[47]) & (g2229) & (g238)) + ((!g2148) & (sk[47]) & (!g2229) & (g238)) + ((!g2148) & (sk[47]) & (g2229) & (g238)) + ((g2148) & (!sk[47]) & (!g2229) & (g238)) + ((g2148) & (!sk[47]) & (g2229) & (!g238)) + ((g2148) & (!sk[47]) & (g2229) & (g238)) + ((g2148) & (sk[47]) & (g2229) & (!g238)) + ((g2148) & (sk[47]) & (g2229) & (g238)));
	assign g4055 = (((!g2150) & (!g2229) & (!sk[48]) & (g239)) + ((!g2150) & (!g2229) & (sk[48]) & (g239)) + ((!g2150) & (g2229) & (!sk[48]) & (!g239)) + ((!g2150) & (g2229) & (!sk[48]) & (g239)) + ((!g2150) & (g2229) & (sk[48]) & (g239)) + ((g2150) & (!g2229) & (!sk[48]) & (g239)) + ((g2150) & (g2229) & (!sk[48]) & (!g239)) + ((g2150) & (g2229) & (!sk[48]) & (g239)) + ((g2150) & (g2229) & (sk[48]) & (!g239)) + ((g2150) & (g2229) & (sk[48]) & (g239)));
	assign g4056 = (((!sk[49]) & (!g2151) & (!g2229) & (g240)) + ((!sk[49]) & (!g2151) & (g2229) & (!g240)) + ((!sk[49]) & (!g2151) & (g2229) & (g240)) + ((!sk[49]) & (g2151) & (!g2229) & (g240)) + ((!sk[49]) & (g2151) & (g2229) & (!g240)) + ((!sk[49]) & (g2151) & (g2229) & (g240)) + ((sk[49]) & (!g2151) & (!g2229) & (g240)) + ((sk[49]) & (!g2151) & (g2229) & (g240)) + ((sk[49]) & (g2151) & (g2229) & (!g240)) + ((sk[49]) & (g2151) & (g2229) & (g240)));
	assign g241 = (((!g237) & (!g238) & (!g239) & (g240) & (g147) & (g148)) + ((!g237) & (!g238) & (g239) & (!g240) & (!g147) & (g148)) + ((!g237) & (!g238) & (g239) & (g240) & (!g147) & (g148)) + ((!g237) & (!g238) & (g239) & (g240) & (g147) & (g148)) + ((!g237) & (g238) & (!g239) & (!g240) & (g147) & (!g148)) + ((!g237) & (g238) & (!g239) & (g240) & (g147) & (!g148)) + ((!g237) & (g238) & (!g239) & (g240) & (g147) & (g148)) + ((!g237) & (g238) & (g239) & (!g240) & (!g147) & (g148)) + ((!g237) & (g238) & (g239) & (!g240) & (g147) & (!g148)) + ((!g237) & (g238) & (g239) & (g240) & (!g147) & (g148)) + ((!g237) & (g238) & (g239) & (g240) & (g147) & (!g148)) + ((!g237) & (g238) & (g239) & (g240) & (g147) & (g148)) + ((g237) & (!g238) & (!g239) & (!g240) & (!g147) & (!g148)) + ((g237) & (!g238) & (!g239) & (g240) & (!g147) & (!g148)) + ((g237) & (!g238) & (!g239) & (g240) & (g147) & (g148)) + ((g237) & (!g238) & (g239) & (!g240) & (!g147) & (!g148)) + ((g237) & (!g238) & (g239) & (!g240) & (!g147) & (g148)) + ((g237) & (!g238) & (g239) & (g240) & (!g147) & (!g148)) + ((g237) & (!g238) & (g239) & (g240) & (!g147) & (g148)) + ((g237) & (!g238) & (g239) & (g240) & (g147) & (g148)) + ((g237) & (g238) & (!g239) & (!g240) & (!g147) & (!g148)) + ((g237) & (g238) & (!g239) & (!g240) & (g147) & (!g148)) + ((g237) & (g238) & (!g239) & (g240) & (!g147) & (!g148)) + ((g237) & (g238) & (!g239) & (g240) & (g147) & (!g148)) + ((g237) & (g238) & (!g239) & (g240) & (g147) & (g148)) + ((g237) & (g238) & (g239) & (!g240) & (!g147) & (!g148)) + ((g237) & (g238) & (g239) & (!g240) & (!g147) & (g148)) + ((g237) & (g238) & (g239) & (!g240) & (g147) & (!g148)) + ((g237) & (g238) & (g239) & (g240) & (!g147) & (!g148)) + ((g237) & (g238) & (g239) & (g240) & (!g147) & (g148)) + ((g237) & (g238) & (g239) & (g240) & (g147) & (!g148)) + ((g237) & (g238) & (g239) & (g240) & (g147) & (g148)));
	assign g4057 = (((!g2152) & (!sk[51]) & (!g2229) & (g242)) + ((!g2152) & (!sk[51]) & (g2229) & (!g242)) + ((!g2152) & (!sk[51]) & (g2229) & (g242)) + ((!g2152) & (sk[51]) & (!g2229) & (g242)) + ((!g2152) & (sk[51]) & (g2229) & (g242)) + ((g2152) & (!sk[51]) & (!g2229) & (g242)) + ((g2152) & (!sk[51]) & (g2229) & (!g242)) + ((g2152) & (!sk[51]) & (g2229) & (g242)) + ((g2152) & (sk[51]) & (g2229) & (!g242)) + ((g2152) & (sk[51]) & (g2229) & (g242)));
	assign g4058 = (((!g2153) & (!g2229) & (!sk[52]) & (g243)) + ((!g2153) & (!g2229) & (sk[52]) & (g243)) + ((!g2153) & (g2229) & (!sk[52]) & (!g243)) + ((!g2153) & (g2229) & (!sk[52]) & (g243)) + ((!g2153) & (g2229) & (sk[52]) & (g243)) + ((g2153) & (!g2229) & (!sk[52]) & (g243)) + ((g2153) & (g2229) & (!sk[52]) & (!g243)) + ((g2153) & (g2229) & (!sk[52]) & (g243)) + ((g2153) & (g2229) & (sk[52]) & (!g243)) + ((g2153) & (g2229) & (sk[52]) & (g243)));
	assign g4059 = (((!sk[53]) & (!g2155) & (!g2229) & (g244)) + ((!sk[53]) & (!g2155) & (g2229) & (!g244)) + ((!sk[53]) & (!g2155) & (g2229) & (g244)) + ((!sk[53]) & (g2155) & (!g2229) & (g244)) + ((!sk[53]) & (g2155) & (g2229) & (!g244)) + ((!sk[53]) & (g2155) & (g2229) & (g244)) + ((sk[53]) & (!g2155) & (!g2229) & (g244)) + ((sk[53]) & (!g2155) & (g2229) & (g244)) + ((sk[53]) & (g2155) & (g2229) & (!g244)) + ((sk[53]) & (g2155) & (g2229) & (g244)));
	assign g4060 = (((!g2157) & (!g2229) & (!sk[54]) & (g245)) + ((!g2157) & (!g2229) & (sk[54]) & (g245)) + ((!g2157) & (g2229) & (!sk[54]) & (!g245)) + ((!g2157) & (g2229) & (!sk[54]) & (g245)) + ((!g2157) & (g2229) & (sk[54]) & (g245)) + ((g2157) & (!g2229) & (!sk[54]) & (g245)) + ((g2157) & (g2229) & (!sk[54]) & (!g245)) + ((g2157) & (g2229) & (!sk[54]) & (g245)) + ((g2157) & (g2229) & (sk[54]) & (!g245)) + ((g2157) & (g2229) & (sk[54]) & (g245)));
	assign g246 = (((!g242) & (!g243) & (!g244) & (g245) & (g147) & (g148)) + ((!g242) & (!g243) & (g244) & (!g245) & (!g147) & (g148)) + ((!g242) & (!g243) & (g244) & (g245) & (!g147) & (g148)) + ((!g242) & (!g243) & (g244) & (g245) & (g147) & (g148)) + ((!g242) & (g243) & (!g244) & (!g245) & (g147) & (!g148)) + ((!g242) & (g243) & (!g244) & (g245) & (g147) & (!g148)) + ((!g242) & (g243) & (!g244) & (g245) & (g147) & (g148)) + ((!g242) & (g243) & (g244) & (!g245) & (!g147) & (g148)) + ((!g242) & (g243) & (g244) & (!g245) & (g147) & (!g148)) + ((!g242) & (g243) & (g244) & (g245) & (!g147) & (g148)) + ((!g242) & (g243) & (g244) & (g245) & (g147) & (!g148)) + ((!g242) & (g243) & (g244) & (g245) & (g147) & (g148)) + ((g242) & (!g243) & (!g244) & (!g245) & (!g147) & (!g148)) + ((g242) & (!g243) & (!g244) & (g245) & (!g147) & (!g148)) + ((g242) & (!g243) & (!g244) & (g245) & (g147) & (g148)) + ((g242) & (!g243) & (g244) & (!g245) & (!g147) & (!g148)) + ((g242) & (!g243) & (g244) & (!g245) & (!g147) & (g148)) + ((g242) & (!g243) & (g244) & (g245) & (!g147) & (!g148)) + ((g242) & (!g243) & (g244) & (g245) & (!g147) & (g148)) + ((g242) & (!g243) & (g244) & (g245) & (g147) & (g148)) + ((g242) & (g243) & (!g244) & (!g245) & (!g147) & (!g148)) + ((g242) & (g243) & (!g244) & (!g245) & (g147) & (!g148)) + ((g242) & (g243) & (!g244) & (g245) & (!g147) & (!g148)) + ((g242) & (g243) & (!g244) & (g245) & (g147) & (!g148)) + ((g242) & (g243) & (!g244) & (g245) & (g147) & (g148)) + ((g242) & (g243) & (g244) & (!g245) & (!g147) & (!g148)) + ((g242) & (g243) & (g244) & (!g245) & (!g147) & (g148)) + ((g242) & (g243) & (g244) & (!g245) & (g147) & (!g148)) + ((g242) & (g243) & (g244) & (g245) & (!g147) & (!g148)) + ((g242) & (g243) & (g244) & (g245) & (!g147) & (g148)) + ((g242) & (g243) & (g244) & (g245) & (g147) & (!g148)) + ((g242) & (g243) & (g244) & (g245) & (g147) & (g148)));
	assign g4061 = (((!sk[56]) & (!g2158) & (!g2229) & (g247)) + ((!sk[56]) & (!g2158) & (g2229) & (!g247)) + ((!sk[56]) & (!g2158) & (g2229) & (g247)) + ((!sk[56]) & (g2158) & (!g2229) & (g247)) + ((!sk[56]) & (g2158) & (g2229) & (!g247)) + ((!sk[56]) & (g2158) & (g2229) & (g247)) + ((sk[56]) & (!g2158) & (!g2229) & (g247)) + ((sk[56]) & (!g2158) & (g2229) & (g247)) + ((sk[56]) & (g2158) & (g2229) & (!g247)) + ((sk[56]) & (g2158) & (g2229) & (g247)));
	assign g4062 = (((!g2159) & (!g2229) & (!sk[57]) & (g248)) + ((!g2159) & (!g2229) & (sk[57]) & (g248)) + ((!g2159) & (g2229) & (!sk[57]) & (!g248)) + ((!g2159) & (g2229) & (!sk[57]) & (g248)) + ((!g2159) & (g2229) & (sk[57]) & (g248)) + ((g2159) & (!g2229) & (!sk[57]) & (g248)) + ((g2159) & (g2229) & (!sk[57]) & (!g248)) + ((g2159) & (g2229) & (!sk[57]) & (g248)) + ((g2159) & (g2229) & (sk[57]) & (!g248)) + ((g2159) & (g2229) & (sk[57]) & (g248)));
	assign g4063 = (((!g2160) & (!g2229) & (!sk[58]) & (g249)) + ((!g2160) & (!g2229) & (sk[58]) & (g249)) + ((!g2160) & (g2229) & (!sk[58]) & (!g249)) + ((!g2160) & (g2229) & (!sk[58]) & (g249)) + ((!g2160) & (g2229) & (sk[58]) & (g249)) + ((g2160) & (!g2229) & (!sk[58]) & (g249)) + ((g2160) & (g2229) & (!sk[58]) & (!g249)) + ((g2160) & (g2229) & (!sk[58]) & (g249)) + ((g2160) & (g2229) & (sk[58]) & (!g249)) + ((g2160) & (g2229) & (sk[58]) & (g249)));
	assign g4064 = (((!g2161) & (!g2229) & (!sk[59]) & (g250)) + ((!g2161) & (!g2229) & (sk[59]) & (g250)) + ((!g2161) & (g2229) & (!sk[59]) & (!g250)) + ((!g2161) & (g2229) & (!sk[59]) & (g250)) + ((!g2161) & (g2229) & (sk[59]) & (g250)) + ((g2161) & (!g2229) & (!sk[59]) & (g250)) + ((g2161) & (g2229) & (!sk[59]) & (!g250)) + ((g2161) & (g2229) & (!sk[59]) & (g250)) + ((g2161) & (g2229) & (sk[59]) & (!g250)) + ((g2161) & (g2229) & (sk[59]) & (g250)));
	assign g251 = (((!g247) & (!g248) & (!g249) & (g250) & (g147) & (g148)) + ((!g247) & (!g248) & (g249) & (!g250) & (!g147) & (g148)) + ((!g247) & (!g248) & (g249) & (g250) & (!g147) & (g148)) + ((!g247) & (!g248) & (g249) & (g250) & (g147) & (g148)) + ((!g247) & (g248) & (!g249) & (!g250) & (g147) & (!g148)) + ((!g247) & (g248) & (!g249) & (g250) & (g147) & (!g148)) + ((!g247) & (g248) & (!g249) & (g250) & (g147) & (g148)) + ((!g247) & (g248) & (g249) & (!g250) & (!g147) & (g148)) + ((!g247) & (g248) & (g249) & (!g250) & (g147) & (!g148)) + ((!g247) & (g248) & (g249) & (g250) & (!g147) & (g148)) + ((!g247) & (g248) & (g249) & (g250) & (g147) & (!g148)) + ((!g247) & (g248) & (g249) & (g250) & (g147) & (g148)) + ((g247) & (!g248) & (!g249) & (!g250) & (!g147) & (!g148)) + ((g247) & (!g248) & (!g249) & (g250) & (!g147) & (!g148)) + ((g247) & (!g248) & (!g249) & (g250) & (g147) & (g148)) + ((g247) & (!g248) & (g249) & (!g250) & (!g147) & (!g148)) + ((g247) & (!g248) & (g249) & (!g250) & (!g147) & (g148)) + ((g247) & (!g248) & (g249) & (g250) & (!g147) & (!g148)) + ((g247) & (!g248) & (g249) & (g250) & (!g147) & (g148)) + ((g247) & (!g248) & (g249) & (g250) & (g147) & (g148)) + ((g247) & (g248) & (!g249) & (!g250) & (!g147) & (!g148)) + ((g247) & (g248) & (!g249) & (!g250) & (g147) & (!g148)) + ((g247) & (g248) & (!g249) & (g250) & (!g147) & (!g148)) + ((g247) & (g248) & (!g249) & (g250) & (g147) & (!g148)) + ((g247) & (g248) & (!g249) & (g250) & (g147) & (g148)) + ((g247) & (g248) & (g249) & (!g250) & (!g147) & (!g148)) + ((g247) & (g248) & (g249) & (!g250) & (!g147) & (g148)) + ((g247) & (g248) & (g249) & (!g250) & (g147) & (!g148)) + ((g247) & (g248) & (g249) & (g250) & (!g147) & (!g148)) + ((g247) & (g248) & (g249) & (g250) & (!g147) & (g148)) + ((g247) & (g248) & (g249) & (g250) & (g147) & (!g148)) + ((g247) & (g248) & (g249) & (g250) & (g147) & (g148)));
	assign g252 = (((!g236) & (!g241) & (!g246) & (g251) & (g165) & (g166)) + ((!g236) & (!g241) & (g246) & (!g251) & (!g165) & (g166)) + ((!g236) & (!g241) & (g246) & (g251) & (!g165) & (g166)) + ((!g236) & (!g241) & (g246) & (g251) & (g165) & (g166)) + ((!g236) & (g241) & (!g246) & (!g251) & (g165) & (!g166)) + ((!g236) & (g241) & (!g246) & (g251) & (g165) & (!g166)) + ((!g236) & (g241) & (!g246) & (g251) & (g165) & (g166)) + ((!g236) & (g241) & (g246) & (!g251) & (!g165) & (g166)) + ((!g236) & (g241) & (g246) & (!g251) & (g165) & (!g166)) + ((!g236) & (g241) & (g246) & (g251) & (!g165) & (g166)) + ((!g236) & (g241) & (g246) & (g251) & (g165) & (!g166)) + ((!g236) & (g241) & (g246) & (g251) & (g165) & (g166)) + ((g236) & (!g241) & (!g246) & (!g251) & (!g165) & (!g166)) + ((g236) & (!g241) & (!g246) & (g251) & (!g165) & (!g166)) + ((g236) & (!g241) & (!g246) & (g251) & (g165) & (g166)) + ((g236) & (!g241) & (g246) & (!g251) & (!g165) & (!g166)) + ((g236) & (!g241) & (g246) & (!g251) & (!g165) & (g166)) + ((g236) & (!g241) & (g246) & (g251) & (!g165) & (!g166)) + ((g236) & (!g241) & (g246) & (g251) & (!g165) & (g166)) + ((g236) & (!g241) & (g246) & (g251) & (g165) & (g166)) + ((g236) & (g241) & (!g246) & (!g251) & (!g165) & (!g166)) + ((g236) & (g241) & (!g246) & (!g251) & (g165) & (!g166)) + ((g236) & (g241) & (!g246) & (g251) & (!g165) & (!g166)) + ((g236) & (g241) & (!g246) & (g251) & (g165) & (!g166)) + ((g236) & (g241) & (!g246) & (g251) & (g165) & (g166)) + ((g236) & (g241) & (g246) & (!g251) & (!g165) & (!g166)) + ((g236) & (g241) & (g246) & (!g251) & (!g165) & (g166)) + ((g236) & (g241) & (g246) & (!g251) & (g165) & (!g166)) + ((g236) & (g241) & (g246) & (g251) & (!g165) & (!g166)) + ((g236) & (g241) & (g246) & (g251) & (!g165) & (g166)) + ((g236) & (g241) & (g246) & (g251) & (g165) & (!g166)) + ((g236) & (g241) & (g246) & (g251) & (g165) & (g166)));
	assign g4065 = (((!g2173) & (!g2229) & (!sk[62]) & (g253)) + ((!g2173) & (!g2229) & (sk[62]) & (g253)) + ((!g2173) & (g2229) & (!sk[62]) & (!g253)) + ((!g2173) & (g2229) & (!sk[62]) & (g253)) + ((!g2173) & (g2229) & (sk[62]) & (g253)) + ((g2173) & (!g2229) & (!sk[62]) & (g253)) + ((g2173) & (g2229) & (!sk[62]) & (!g253)) + ((g2173) & (g2229) & (!sk[62]) & (g253)) + ((g2173) & (g2229) & (sk[62]) & (!g253)) + ((g2173) & (g2229) & (sk[62]) & (g253)));
	assign g4066 = (((!g2174) & (!sk[63]) & (!g2229) & (g254)) + ((!g2174) & (!sk[63]) & (g2229) & (!g254)) + ((!g2174) & (!sk[63]) & (g2229) & (g254)) + ((!g2174) & (sk[63]) & (!g2229) & (g254)) + ((!g2174) & (sk[63]) & (g2229) & (g254)) + ((g2174) & (!sk[63]) & (!g2229) & (g254)) + ((g2174) & (!sk[63]) & (g2229) & (!g254)) + ((g2174) & (!sk[63]) & (g2229) & (g254)) + ((g2174) & (sk[63]) & (g2229) & (!g254)) + ((g2174) & (sk[63]) & (g2229) & (g254)));
	assign g4067 = (((!g2175) & (!sk[64]) & (!g2229) & (g255)) + ((!g2175) & (!sk[64]) & (g2229) & (!g255)) + ((!g2175) & (!sk[64]) & (g2229) & (g255)) + ((!g2175) & (sk[64]) & (!g2229) & (g255)) + ((!g2175) & (sk[64]) & (g2229) & (g255)) + ((g2175) & (!sk[64]) & (!g2229) & (g255)) + ((g2175) & (!sk[64]) & (g2229) & (!g255)) + ((g2175) & (!sk[64]) & (g2229) & (g255)) + ((g2175) & (sk[64]) & (g2229) & (!g255)) + ((g2175) & (sk[64]) & (g2229) & (g255)));
	assign g4068 = (((!g2176) & (!sk[65]) & (!g2229) & (g256)) + ((!g2176) & (!sk[65]) & (g2229) & (!g256)) + ((!g2176) & (!sk[65]) & (g2229) & (g256)) + ((!g2176) & (sk[65]) & (!g2229) & (g256)) + ((!g2176) & (sk[65]) & (g2229) & (g256)) + ((g2176) & (!sk[65]) & (!g2229) & (g256)) + ((g2176) & (!sk[65]) & (g2229) & (!g256)) + ((g2176) & (!sk[65]) & (g2229) & (g256)) + ((g2176) & (sk[65]) & (g2229) & (!g256)) + ((g2176) & (sk[65]) & (g2229) & (g256)));
	assign g257 = (((!g253) & (!g254) & (!g255) & (g256) & (g165) & (g166)) + ((!g253) & (!g254) & (g255) & (!g256) & (!g165) & (g166)) + ((!g253) & (!g254) & (g255) & (g256) & (!g165) & (g166)) + ((!g253) & (!g254) & (g255) & (g256) & (g165) & (g166)) + ((!g253) & (g254) & (!g255) & (!g256) & (g165) & (!g166)) + ((!g253) & (g254) & (!g255) & (g256) & (g165) & (!g166)) + ((!g253) & (g254) & (!g255) & (g256) & (g165) & (g166)) + ((!g253) & (g254) & (g255) & (!g256) & (!g165) & (g166)) + ((!g253) & (g254) & (g255) & (!g256) & (g165) & (!g166)) + ((!g253) & (g254) & (g255) & (g256) & (!g165) & (g166)) + ((!g253) & (g254) & (g255) & (g256) & (g165) & (!g166)) + ((!g253) & (g254) & (g255) & (g256) & (g165) & (g166)) + ((g253) & (!g254) & (!g255) & (!g256) & (!g165) & (!g166)) + ((g253) & (!g254) & (!g255) & (g256) & (!g165) & (!g166)) + ((g253) & (!g254) & (!g255) & (g256) & (g165) & (g166)) + ((g253) & (!g254) & (g255) & (!g256) & (!g165) & (!g166)) + ((g253) & (!g254) & (g255) & (!g256) & (!g165) & (g166)) + ((g253) & (!g254) & (g255) & (g256) & (!g165) & (!g166)) + ((g253) & (!g254) & (g255) & (g256) & (!g165) & (g166)) + ((g253) & (!g254) & (g255) & (g256) & (g165) & (g166)) + ((g253) & (g254) & (!g255) & (!g256) & (!g165) & (!g166)) + ((g253) & (g254) & (!g255) & (!g256) & (g165) & (!g166)) + ((g253) & (g254) & (!g255) & (g256) & (!g165) & (!g166)) + ((g253) & (g254) & (!g255) & (g256) & (g165) & (!g166)) + ((g253) & (g254) & (!g255) & (g256) & (g165) & (g166)) + ((g253) & (g254) & (g255) & (!g256) & (!g165) & (!g166)) + ((g253) & (g254) & (g255) & (!g256) & (!g165) & (g166)) + ((g253) & (g254) & (g255) & (!g256) & (g165) & (!g166)) + ((g253) & (g254) & (g255) & (g256) & (!g165) & (!g166)) + ((g253) & (g254) & (g255) & (g256) & (!g165) & (g166)) + ((g253) & (g254) & (g255) & (g256) & (g165) & (!g166)) + ((g253) & (g254) & (g255) & (g256) & (g165) & (g166)));
	assign g4069 = (((!sk[67]) & (!g2177) & (!g2229) & (g258)) + ((!sk[67]) & (!g2177) & (g2229) & (!g258)) + ((!sk[67]) & (!g2177) & (g2229) & (g258)) + ((!sk[67]) & (g2177) & (!g2229) & (g258)) + ((!sk[67]) & (g2177) & (g2229) & (!g258)) + ((!sk[67]) & (g2177) & (g2229) & (g258)) + ((sk[67]) & (!g2177) & (!g2229) & (g258)) + ((sk[67]) & (!g2177) & (g2229) & (g258)) + ((sk[67]) & (g2177) & (g2229) & (!g258)) + ((sk[67]) & (g2177) & (g2229) & (g258)));
	assign g4070 = (((!g2178) & (!sk[68]) & (!g2229) & (g259)) + ((!g2178) & (!sk[68]) & (g2229) & (!g259)) + ((!g2178) & (!sk[68]) & (g2229) & (g259)) + ((!g2178) & (sk[68]) & (!g2229) & (g259)) + ((!g2178) & (sk[68]) & (g2229) & (g259)) + ((g2178) & (!sk[68]) & (!g2229) & (g259)) + ((g2178) & (!sk[68]) & (g2229) & (!g259)) + ((g2178) & (!sk[68]) & (g2229) & (g259)) + ((g2178) & (sk[68]) & (g2229) & (!g259)) + ((g2178) & (sk[68]) & (g2229) & (g259)));
	assign g4071 = (((!g2179) & (!sk[69]) & (!g2229) & (g260)) + ((!g2179) & (!sk[69]) & (g2229) & (!g260)) + ((!g2179) & (!sk[69]) & (g2229) & (g260)) + ((!g2179) & (sk[69]) & (!g2229) & (g260)) + ((!g2179) & (sk[69]) & (g2229) & (g260)) + ((g2179) & (!sk[69]) & (!g2229) & (g260)) + ((g2179) & (!sk[69]) & (g2229) & (!g260)) + ((g2179) & (!sk[69]) & (g2229) & (g260)) + ((g2179) & (sk[69]) & (g2229) & (!g260)) + ((g2179) & (sk[69]) & (g2229) & (g260)));
	assign g261 = (((!sk[70]) & (!g165) & (!g166) & (!g258) & (g259) & (!g260)) + ((!sk[70]) & (!g165) & (!g166) & (!g258) & (g259) & (g260)) + ((!sk[70]) & (!g165) & (!g166) & (g258) & (!g259) & (!g260)) + ((!sk[70]) & (!g165) & (!g166) & (g258) & (!g259) & (g260)) + ((!sk[70]) & (!g165) & (!g166) & (g258) & (g259) & (!g260)) + ((!sk[70]) & (!g165) & (!g166) & (g258) & (g259) & (g260)) + ((!sk[70]) & (!g165) & (g166) & (!g258) & (!g259) & (!g260)) + ((!sk[70]) & (!g165) & (g166) & (!g258) & (!g259) & (g260)) + ((!sk[70]) & (!g165) & (g166) & (!g258) & (g259) & (!g260)) + ((!sk[70]) & (!g165) & (g166) & (!g258) & (g259) & (g260)) + ((!sk[70]) & (!g165) & (g166) & (g258) & (!g259) & (!g260)) + ((!sk[70]) & (!g165) & (g166) & (g258) & (!g259) & (g260)) + ((!sk[70]) & (!g165) & (g166) & (g258) & (g259) & (!g260)) + ((!sk[70]) & (!g165) & (g166) & (g258) & (g259) & (g260)) + ((!sk[70]) & (g165) & (!g166) & (!g258) & (g259) & (!g260)) + ((!sk[70]) & (g165) & (!g166) & (!g258) & (g259) & (g260)) + ((!sk[70]) & (g165) & (!g166) & (g258) & (!g259) & (!g260)) + ((!sk[70]) & (g165) & (!g166) & (g258) & (!g259) & (g260)) + ((!sk[70]) & (g165) & (!g166) & (g258) & (g259) & (!g260)) + ((!sk[70]) & (g165) & (!g166) & (g258) & (g259) & (g260)) + ((!sk[70]) & (g165) & (g166) & (!g258) & (!g259) & (!g260)) + ((!sk[70]) & (g165) & (g166) & (!g258) & (!g259) & (g260)) + ((!sk[70]) & (g165) & (g166) & (!g258) & (g259) & (!g260)) + ((!sk[70]) & (g165) & (g166) & (!g258) & (g259) & (g260)) + ((!sk[70]) & (g165) & (g166) & (g258) & (!g259) & (!g260)) + ((!sk[70]) & (g165) & (g166) & (g258) & (!g259) & (g260)) + ((!sk[70]) & (g165) & (g166) & (g258) & (g259) & (!g260)) + ((!sk[70]) & (g165) & (g166) & (g258) & (g259) & (g260)) + ((sk[70]) & (!g165) & (g166) & (!g258) & (!g259) & (g260)) + ((sk[70]) & (!g165) & (g166) & (!g258) & (g259) & (g260)) + ((sk[70]) & (!g165) & (g166) & (g258) & (!g259) & (g260)) + ((sk[70]) & (!g165) & (g166) & (g258) & (g259) & (g260)) + ((sk[70]) & (g165) & (!g166) & (g258) & (!g259) & (!g260)) + ((sk[70]) & (g165) & (!g166) & (g258) & (!g259) & (g260)) + ((sk[70]) & (g165) & (!g166) & (g258) & (g259) & (!g260)) + ((sk[70]) & (g165) & (!g166) & (g258) & (g259) & (g260)) + ((sk[70]) & (g165) & (g166) & (!g258) & (g259) & (!g260)) + ((sk[70]) & (g165) & (g166) & (!g258) & (g259) & (g260)) + ((sk[70]) & (g165) & (g166) & (g258) & (g259) & (!g260)) + ((sk[70]) & (g165) & (g166) & (g258) & (g259) & (g260)));
	assign g4072 = (((!g2162) & (!sk[71]) & (!g2229) & (g262)) + ((!g2162) & (!sk[71]) & (g2229) & (!g262)) + ((!g2162) & (!sk[71]) & (g2229) & (g262)) + ((!g2162) & (sk[71]) & (!g2229) & (g262)) + ((!g2162) & (sk[71]) & (g2229) & (g262)) + ((g2162) & (!sk[71]) & (!g2229) & (g262)) + ((g2162) & (!sk[71]) & (g2229) & (!g262)) + ((g2162) & (!sk[71]) & (g2229) & (g262)) + ((g2162) & (sk[71]) & (g2229) & (!g262)) + ((g2162) & (sk[71]) & (g2229) & (g262)));
	assign g4073 = (((!g2164) & (!sk[72]) & (!g2229) & (g263)) + ((!g2164) & (!sk[72]) & (g2229) & (!g263)) + ((!g2164) & (!sk[72]) & (g2229) & (g263)) + ((!g2164) & (sk[72]) & (!g2229) & (g263)) + ((!g2164) & (sk[72]) & (g2229) & (g263)) + ((g2164) & (!sk[72]) & (!g2229) & (g263)) + ((g2164) & (!sk[72]) & (g2229) & (!g263)) + ((g2164) & (!sk[72]) & (g2229) & (g263)) + ((g2164) & (sk[72]) & (g2229) & (!g263)) + ((g2164) & (sk[72]) & (g2229) & (g263)));
	assign g4074 = (((!g2166) & (!sk[73]) & (!g2229) & (g264)) + ((!g2166) & (!sk[73]) & (g2229) & (!g264)) + ((!g2166) & (!sk[73]) & (g2229) & (g264)) + ((!g2166) & (sk[73]) & (!g2229) & (g264)) + ((!g2166) & (sk[73]) & (g2229) & (g264)) + ((g2166) & (!sk[73]) & (!g2229) & (g264)) + ((g2166) & (!sk[73]) & (g2229) & (!g264)) + ((g2166) & (!sk[73]) & (g2229) & (g264)) + ((g2166) & (sk[73]) & (g2229) & (!g264)) + ((g2166) & (sk[73]) & (g2229) & (g264)));
	assign g4075 = (((!sk[74]) & (!g2168) & (!g2229) & (g265)) + ((!sk[74]) & (!g2168) & (g2229) & (!g265)) + ((!sk[74]) & (!g2168) & (g2229) & (g265)) + ((!sk[74]) & (g2168) & (!g2229) & (g265)) + ((!sk[74]) & (g2168) & (g2229) & (!g265)) + ((!sk[74]) & (g2168) & (g2229) & (g265)) + ((sk[74]) & (!g2168) & (!g2229) & (g265)) + ((sk[74]) & (!g2168) & (g2229) & (g265)) + ((sk[74]) & (g2168) & (g2229) & (!g265)) + ((sk[74]) & (g2168) & (g2229) & (g265)));
	assign g266 = (((!g262) & (!g263) & (!g264) & (g265) & (g165) & (g166)) + ((!g262) & (!g263) & (g264) & (!g265) & (!g165) & (g166)) + ((!g262) & (!g263) & (g264) & (g265) & (!g165) & (g166)) + ((!g262) & (!g263) & (g264) & (g265) & (g165) & (g166)) + ((!g262) & (g263) & (!g264) & (!g265) & (g165) & (!g166)) + ((!g262) & (g263) & (!g264) & (g265) & (g165) & (!g166)) + ((!g262) & (g263) & (!g264) & (g265) & (g165) & (g166)) + ((!g262) & (g263) & (g264) & (!g265) & (!g165) & (g166)) + ((!g262) & (g263) & (g264) & (!g265) & (g165) & (!g166)) + ((!g262) & (g263) & (g264) & (g265) & (!g165) & (g166)) + ((!g262) & (g263) & (g264) & (g265) & (g165) & (!g166)) + ((!g262) & (g263) & (g264) & (g265) & (g165) & (g166)) + ((g262) & (!g263) & (!g264) & (!g265) & (!g165) & (!g166)) + ((g262) & (!g263) & (!g264) & (g265) & (!g165) & (!g166)) + ((g262) & (!g263) & (!g264) & (g265) & (g165) & (g166)) + ((g262) & (!g263) & (g264) & (!g265) & (!g165) & (!g166)) + ((g262) & (!g263) & (g264) & (!g265) & (!g165) & (g166)) + ((g262) & (!g263) & (g264) & (g265) & (!g165) & (!g166)) + ((g262) & (!g263) & (g264) & (g265) & (!g165) & (g166)) + ((g262) & (!g263) & (g264) & (g265) & (g165) & (g166)) + ((g262) & (g263) & (!g264) & (!g265) & (!g165) & (!g166)) + ((g262) & (g263) & (!g264) & (!g265) & (g165) & (!g166)) + ((g262) & (g263) & (!g264) & (g265) & (!g165) & (!g166)) + ((g262) & (g263) & (!g264) & (g265) & (g165) & (!g166)) + ((g262) & (g263) & (!g264) & (g265) & (g165) & (g166)) + ((g262) & (g263) & (g264) & (!g265) & (!g165) & (!g166)) + ((g262) & (g263) & (g264) & (!g265) & (!g165) & (g166)) + ((g262) & (g263) & (g264) & (!g265) & (g165) & (!g166)) + ((g262) & (g263) & (g264) & (g265) & (!g165) & (!g166)) + ((g262) & (g263) & (g264) & (g265) & (!g165) & (g166)) + ((g262) & (g263) & (g264) & (g265) & (g165) & (!g166)) + ((g262) & (g263) & (g264) & (g265) & (g165) & (g166)));
	assign g4076 = (((!g2169) & (!g2229) & (!sk[76]) & (g267)) + ((!g2169) & (!g2229) & (sk[76]) & (g267)) + ((!g2169) & (g2229) & (!sk[76]) & (!g267)) + ((!g2169) & (g2229) & (!sk[76]) & (g267)) + ((!g2169) & (g2229) & (sk[76]) & (g267)) + ((g2169) & (!g2229) & (!sk[76]) & (g267)) + ((g2169) & (g2229) & (!sk[76]) & (!g267)) + ((g2169) & (g2229) & (!sk[76]) & (g267)) + ((g2169) & (g2229) & (sk[76]) & (!g267)) + ((g2169) & (g2229) & (sk[76]) & (g267)));
	assign g4077 = (((!g2170) & (!sk[77]) & (!g2229) & (g268)) + ((!g2170) & (!sk[77]) & (g2229) & (!g268)) + ((!g2170) & (!sk[77]) & (g2229) & (g268)) + ((!g2170) & (sk[77]) & (!g2229) & (g268)) + ((!g2170) & (sk[77]) & (g2229) & (g268)) + ((g2170) & (!sk[77]) & (!g2229) & (g268)) + ((g2170) & (!sk[77]) & (g2229) & (!g268)) + ((g2170) & (!sk[77]) & (g2229) & (g268)) + ((g2170) & (sk[77]) & (g2229) & (!g268)) + ((g2170) & (sk[77]) & (g2229) & (g268)));
	assign g4078 = (((!g2171) & (!g2229) & (!sk[78]) & (g269)) + ((!g2171) & (!g2229) & (sk[78]) & (g269)) + ((!g2171) & (g2229) & (!sk[78]) & (!g269)) + ((!g2171) & (g2229) & (!sk[78]) & (g269)) + ((!g2171) & (g2229) & (sk[78]) & (g269)) + ((g2171) & (!g2229) & (!sk[78]) & (g269)) + ((g2171) & (g2229) & (!sk[78]) & (!g269)) + ((g2171) & (g2229) & (!sk[78]) & (g269)) + ((g2171) & (g2229) & (sk[78]) & (!g269)) + ((g2171) & (g2229) & (sk[78]) & (g269)));
	assign g4079 = (((!g2172) & (!sk[79]) & (!g2229) & (g270)) + ((!g2172) & (!sk[79]) & (g2229) & (!g270)) + ((!g2172) & (!sk[79]) & (g2229) & (g270)) + ((!g2172) & (sk[79]) & (!g2229) & (g270)) + ((!g2172) & (sk[79]) & (g2229) & (g270)) + ((g2172) & (!sk[79]) & (!g2229) & (g270)) + ((g2172) & (!sk[79]) & (g2229) & (!g270)) + ((g2172) & (!sk[79]) & (g2229) & (g270)) + ((g2172) & (sk[79]) & (g2229) & (!g270)) + ((g2172) & (sk[79]) & (g2229) & (g270)));
	assign g271 = (((!g267) & (!g268) & (!g269) & (g270) & (g165) & (g166)) + ((!g267) & (!g268) & (g269) & (!g270) & (!g165) & (g166)) + ((!g267) & (!g268) & (g269) & (g270) & (!g165) & (g166)) + ((!g267) & (!g268) & (g269) & (g270) & (g165) & (g166)) + ((!g267) & (g268) & (!g269) & (!g270) & (g165) & (!g166)) + ((!g267) & (g268) & (!g269) & (g270) & (g165) & (!g166)) + ((!g267) & (g268) & (!g269) & (g270) & (g165) & (g166)) + ((!g267) & (g268) & (g269) & (!g270) & (!g165) & (g166)) + ((!g267) & (g268) & (g269) & (!g270) & (g165) & (!g166)) + ((!g267) & (g268) & (g269) & (g270) & (!g165) & (g166)) + ((!g267) & (g268) & (g269) & (g270) & (g165) & (!g166)) + ((!g267) & (g268) & (g269) & (g270) & (g165) & (g166)) + ((g267) & (!g268) & (!g269) & (!g270) & (!g165) & (!g166)) + ((g267) & (!g268) & (!g269) & (g270) & (!g165) & (!g166)) + ((g267) & (!g268) & (!g269) & (g270) & (g165) & (g166)) + ((g267) & (!g268) & (g269) & (!g270) & (!g165) & (!g166)) + ((g267) & (!g268) & (g269) & (!g270) & (!g165) & (g166)) + ((g267) & (!g268) & (g269) & (g270) & (!g165) & (!g166)) + ((g267) & (!g268) & (g269) & (g270) & (!g165) & (g166)) + ((g267) & (!g268) & (g269) & (g270) & (g165) & (g166)) + ((g267) & (g268) & (!g269) & (!g270) & (!g165) & (!g166)) + ((g267) & (g268) & (!g269) & (!g270) & (g165) & (!g166)) + ((g267) & (g268) & (!g269) & (g270) & (!g165) & (!g166)) + ((g267) & (g268) & (!g269) & (g270) & (g165) & (!g166)) + ((g267) & (g268) & (!g269) & (g270) & (g165) & (g166)) + ((g267) & (g268) & (g269) & (!g270) & (!g165) & (!g166)) + ((g267) & (g268) & (g269) & (!g270) & (!g165) & (g166)) + ((g267) & (g268) & (g269) & (!g270) & (g165) & (!g166)) + ((g267) & (g268) & (g269) & (g270) & (!g165) & (!g166)) + ((g267) & (g268) & (g269) & (g270) & (!g165) & (g166)) + ((g267) & (g268) & (g269) & (g270) & (g165) & (!g166)) + ((g267) & (g268) & (g269) & (g270) & (g165) & (g166)));
	assign g272 = (((!g147) & (!g148) & (!g257) & (g261) & (!g266) & (!g271)) + ((!g147) & (!g148) & (!g257) & (g261) & (!g266) & (g271)) + ((!g147) & (!g148) & (!g257) & (g261) & (g266) & (!g271)) + ((!g147) & (!g148) & (!g257) & (g261) & (g266) & (g271)) + ((!g147) & (!g148) & (g257) & (g261) & (!g266) & (!g271)) + ((!g147) & (!g148) & (g257) & (g261) & (!g266) & (g271)) + ((!g147) & (!g148) & (g257) & (g261) & (g266) & (!g271)) + ((!g147) & (!g148) & (g257) & (g261) & (g266) & (g271)) + ((!g147) & (g148) & (!g257) & (!g261) & (!g266) & (g271)) + ((!g147) & (g148) & (!g257) & (!g261) & (g266) & (g271)) + ((!g147) & (g148) & (!g257) & (g261) & (!g266) & (g271)) + ((!g147) & (g148) & (!g257) & (g261) & (g266) & (g271)) + ((!g147) & (g148) & (g257) & (!g261) & (!g266) & (g271)) + ((!g147) & (g148) & (g257) & (!g261) & (g266) & (g271)) + ((!g147) & (g148) & (g257) & (g261) & (!g266) & (g271)) + ((!g147) & (g148) & (g257) & (g261) & (g266) & (g271)) + ((g147) & (!g148) & (g257) & (!g261) & (!g266) & (!g271)) + ((g147) & (!g148) & (g257) & (!g261) & (!g266) & (g271)) + ((g147) & (!g148) & (g257) & (!g261) & (g266) & (!g271)) + ((g147) & (!g148) & (g257) & (!g261) & (g266) & (g271)) + ((g147) & (!g148) & (g257) & (g261) & (!g266) & (!g271)) + ((g147) & (!g148) & (g257) & (g261) & (!g266) & (g271)) + ((g147) & (!g148) & (g257) & (g261) & (g266) & (!g271)) + ((g147) & (!g148) & (g257) & (g261) & (g266) & (g271)) + ((g147) & (g148) & (!g257) & (!g261) & (g266) & (!g271)) + ((g147) & (g148) & (!g257) & (!g261) & (g266) & (g271)) + ((g147) & (g148) & (!g257) & (g261) & (g266) & (!g271)) + ((g147) & (g148) & (!g257) & (g261) & (g266) & (g271)) + ((g147) & (g148) & (g257) & (!g261) & (g266) & (!g271)) + ((g147) & (g148) & (g257) & (!g261) & (g266) & (g271)) + ((g147) & (g148) & (g257) & (g261) & (g266) & (!g271)) + ((g147) & (g148) & (g257) & (g261) & (g266) & (g271)));
	assign g273 = (((!g142) & (!g252) & (!sk[82]) & (g272)) + ((!g142) & (!g252) & (sk[82]) & (g272)) + ((!g142) & (g252) & (!sk[82]) & (!g272)) + ((!g142) & (g252) & (!sk[82]) & (g272)) + ((!g142) & (g252) & (sk[82]) & (g272)) + ((g142) & (!g252) & (!sk[82]) & (g272)) + ((g142) & (g252) & (!sk[82]) & (!g272)) + ((g142) & (g252) & (!sk[82]) & (g272)) + ((g142) & (g252) & (sk[82]) & (!g272)) + ((g142) & (g252) & (sk[82]) & (g272)));
	assign g274 = (((!sk[83]) & (!g87) & (!g126) & (!g141) & (g231) & (!g273)) + ((!sk[83]) & (!g87) & (!g126) & (!g141) & (g231) & (g273)) + ((!sk[83]) & (!g87) & (!g126) & (g141) & (!g231) & (!g273)) + ((!sk[83]) & (!g87) & (!g126) & (g141) & (!g231) & (g273)) + ((!sk[83]) & (!g87) & (!g126) & (g141) & (g231) & (!g273)) + ((!sk[83]) & (!g87) & (!g126) & (g141) & (g231) & (g273)) + ((!sk[83]) & (!g87) & (g126) & (!g141) & (!g231) & (!g273)) + ((!sk[83]) & (!g87) & (g126) & (!g141) & (!g231) & (g273)) + ((!sk[83]) & (!g87) & (g126) & (!g141) & (g231) & (!g273)) + ((!sk[83]) & (!g87) & (g126) & (!g141) & (g231) & (g273)) + ((!sk[83]) & (!g87) & (g126) & (g141) & (!g231) & (!g273)) + ((!sk[83]) & (!g87) & (g126) & (g141) & (!g231) & (g273)) + ((!sk[83]) & (!g87) & (g126) & (g141) & (g231) & (!g273)) + ((!sk[83]) & (!g87) & (g126) & (g141) & (g231) & (g273)) + ((!sk[83]) & (g87) & (!g126) & (!g141) & (g231) & (!g273)) + ((!sk[83]) & (g87) & (!g126) & (!g141) & (g231) & (g273)) + ((!sk[83]) & (g87) & (!g126) & (g141) & (!g231) & (!g273)) + ((!sk[83]) & (g87) & (!g126) & (g141) & (!g231) & (g273)) + ((!sk[83]) & (g87) & (!g126) & (g141) & (g231) & (!g273)) + ((!sk[83]) & (g87) & (!g126) & (g141) & (g231) & (g273)) + ((!sk[83]) & (g87) & (g126) & (!g141) & (!g231) & (!g273)) + ((!sk[83]) & (g87) & (g126) & (!g141) & (!g231) & (g273)) + ((!sk[83]) & (g87) & (g126) & (!g141) & (g231) & (!g273)) + ((!sk[83]) & (g87) & (g126) & (!g141) & (g231) & (g273)) + ((!sk[83]) & (g87) & (g126) & (g141) & (!g231) & (!g273)) + ((!sk[83]) & (g87) & (g126) & (g141) & (!g231) & (g273)) + ((!sk[83]) & (g87) & (g126) & (g141) & (g231) & (!g273)) + ((!sk[83]) & (g87) & (g126) & (g141) & (g231) & (g273)) + ((sk[83]) & (!g87) & (!g126) & (g141) & (!g231) & (!g273)) + ((sk[83]) & (!g87) & (!g126) & (g141) & (!g231) & (g273)) + ((sk[83]) & (!g87) & (!g126) & (g141) & (g231) & (!g273)) + ((sk[83]) & (!g87) & (!g126) & (g141) & (g231) & (g273)) + ((sk[83]) & (!g87) & (g126) & (!g141) & (!g231) & (g273)) + ((sk[83]) & (!g87) & (g126) & (!g141) & (g231) & (!g273)) + ((sk[83]) & (!g87) & (g126) & (g141) & (!g231) & (g273)) + ((sk[83]) & (!g87) & (g126) & (g141) & (g231) & (!g273)) + ((sk[83]) & (g87) & (!g126) & (g141) & (!g231) & (!g273)) + ((sk[83]) & (g87) & (!g126) & (g141) & (!g231) & (g273)) + ((sk[83]) & (g87) & (!g126) & (g141) & (g231) & (!g273)) + ((sk[83]) & (g87) & (!g126) & (g141) & (g231) & (g273)) + ((sk[83]) & (g87) & (g126) & (!g141) & (!g231) & (!g273)) + ((sk[83]) & (g87) & (g126) & (!g141) & (g231) & (g273)) + ((sk[83]) & (g87) & (g126) & (g141) & (!g231) & (!g273)) + ((sk[83]) & (g87) & (g126) & (g141) & (g231) & (g273)));
	assign g4080 = (((!g2059) & (!g2235) & (!sk[84]) & (g275)) + ((!g2059) & (!g2235) & (sk[84]) & (g275)) + ((!g2059) & (g2235) & (!sk[84]) & (!g275)) + ((!g2059) & (g2235) & (!sk[84]) & (g275)) + ((!g2059) & (g2235) & (sk[84]) & (g275)) + ((g2059) & (!g2235) & (!sk[84]) & (g275)) + ((g2059) & (g2235) & (!sk[84]) & (!g275)) + ((g2059) & (g2235) & (!sk[84]) & (g275)) + ((g2059) & (g2235) & (sk[84]) & (!g275)) + ((g2059) & (g2235) & (sk[84]) & (g275)));
	assign g4081 = (((!g2140) & (!sk[85]) & (!g2256) & (g276)) + ((!g2140) & (!sk[85]) & (g2256) & (!g276)) + ((!g2140) & (!sk[85]) & (g2256) & (g276)) + ((!g2140) & (sk[85]) & (!g2256) & (g276)) + ((!g2140) & (sk[85]) & (g2256) & (g276)) + ((g2140) & (!sk[85]) & (!g2256) & (g276)) + ((g2140) & (!sk[85]) & (g2256) & (!g276)) + ((g2140) & (!sk[85]) & (g2256) & (g276)) + ((g2140) & (sk[85]) & (g2256) & (!g276)) + ((g2140) & (sk[85]) & (g2256) & (g276)));
	assign g4082 = (((!g2146) & (!sk[86]) & (!g2256) & (g277)) + ((!g2146) & (!sk[86]) & (g2256) & (!g277)) + ((!g2146) & (!sk[86]) & (g2256) & (g277)) + ((!g2146) & (sk[86]) & (!g2256) & (g277)) + ((!g2146) & (sk[86]) & (g2256) & (g277)) + ((g2146) & (!sk[86]) & (!g2256) & (g277)) + ((g2146) & (!sk[86]) & (g2256) & (!g277)) + ((g2146) & (!sk[86]) & (g2256) & (g277)) + ((g2146) & (sk[86]) & (g2256) & (!g277)) + ((g2146) & (sk[86]) & (g2256) & (g277)));
	assign g4083 = (((!g2152) & (!sk[87]) & (!g2256) & (g278)) + ((!g2152) & (!sk[87]) & (g2256) & (!g278)) + ((!g2152) & (!sk[87]) & (g2256) & (g278)) + ((!g2152) & (sk[87]) & (!g2256) & (g278)) + ((!g2152) & (sk[87]) & (g2256) & (g278)) + ((g2152) & (!sk[87]) & (!g2256) & (g278)) + ((g2152) & (!sk[87]) & (g2256) & (!g278)) + ((g2152) & (!sk[87]) & (g2256) & (g278)) + ((g2152) & (sk[87]) & (g2256) & (!g278)) + ((g2152) & (sk[87]) & (g2256) & (g278)));
	assign g4084 = (((!sk[88]) & (!g2158) & (!g2256) & (g279)) + ((!sk[88]) & (!g2158) & (g2256) & (!g279)) + ((!sk[88]) & (!g2158) & (g2256) & (g279)) + ((!sk[88]) & (g2158) & (!g2256) & (g279)) + ((!sk[88]) & (g2158) & (g2256) & (!g279)) + ((!sk[88]) & (g2158) & (g2256) & (g279)) + ((sk[88]) & (!g2158) & (!g2256) & (g279)) + ((sk[88]) & (!g2158) & (g2256) & (g279)) + ((sk[88]) & (g2158) & (g2256) & (!g279)) + ((sk[88]) & (g2158) & (g2256) & (g279)));
	assign g280 = (((!g276) & (!g277) & (!g278) & (g279) & (g165) & (g166)) + ((!g276) & (!g277) & (g278) & (!g279) & (!g165) & (g166)) + ((!g276) & (!g277) & (g278) & (g279) & (!g165) & (g166)) + ((!g276) & (!g277) & (g278) & (g279) & (g165) & (g166)) + ((!g276) & (g277) & (!g278) & (!g279) & (g165) & (!g166)) + ((!g276) & (g277) & (!g278) & (g279) & (g165) & (!g166)) + ((!g276) & (g277) & (!g278) & (g279) & (g165) & (g166)) + ((!g276) & (g277) & (g278) & (!g279) & (!g165) & (g166)) + ((!g276) & (g277) & (g278) & (!g279) & (g165) & (!g166)) + ((!g276) & (g277) & (g278) & (g279) & (!g165) & (g166)) + ((!g276) & (g277) & (g278) & (g279) & (g165) & (!g166)) + ((!g276) & (g277) & (g278) & (g279) & (g165) & (g166)) + ((g276) & (!g277) & (!g278) & (!g279) & (!g165) & (!g166)) + ((g276) & (!g277) & (!g278) & (g279) & (!g165) & (!g166)) + ((g276) & (!g277) & (!g278) & (g279) & (g165) & (g166)) + ((g276) & (!g277) & (g278) & (!g279) & (!g165) & (!g166)) + ((g276) & (!g277) & (g278) & (!g279) & (!g165) & (g166)) + ((g276) & (!g277) & (g278) & (g279) & (!g165) & (!g166)) + ((g276) & (!g277) & (g278) & (g279) & (!g165) & (g166)) + ((g276) & (!g277) & (g278) & (g279) & (g165) & (g166)) + ((g276) & (g277) & (!g278) & (!g279) & (!g165) & (!g166)) + ((g276) & (g277) & (!g278) & (!g279) & (g165) & (!g166)) + ((g276) & (g277) & (!g278) & (g279) & (!g165) & (!g166)) + ((g276) & (g277) & (!g278) & (g279) & (g165) & (!g166)) + ((g276) & (g277) & (!g278) & (g279) & (g165) & (g166)) + ((g276) & (g277) & (g278) & (!g279) & (!g165) & (!g166)) + ((g276) & (g277) & (g278) & (!g279) & (!g165) & (g166)) + ((g276) & (g277) & (g278) & (!g279) & (g165) & (!g166)) + ((g276) & (g277) & (g278) & (g279) & (!g165) & (!g166)) + ((g276) & (g277) & (g278) & (g279) & (!g165) & (g166)) + ((g276) & (g277) & (g278) & (g279) & (g165) & (!g166)) + ((g276) & (g277) & (g278) & (g279) & (g165) & (g166)));
	assign g4085 = (((!sk[90]) & (!g2142) & (!g2256) & (g281)) + ((!sk[90]) & (!g2142) & (g2256) & (!g281)) + ((!sk[90]) & (!g2142) & (g2256) & (g281)) + ((!sk[90]) & (g2142) & (!g2256) & (g281)) + ((!sk[90]) & (g2142) & (g2256) & (!g281)) + ((!sk[90]) & (g2142) & (g2256) & (g281)) + ((sk[90]) & (!g2142) & (!g2256) & (g281)) + ((sk[90]) & (!g2142) & (g2256) & (g281)) + ((sk[90]) & (g2142) & (g2256) & (!g281)) + ((sk[90]) & (g2142) & (g2256) & (g281)));
	assign g4086 = (((!g2148) & (!sk[91]) & (!g2256) & (g282)) + ((!g2148) & (!sk[91]) & (g2256) & (!g282)) + ((!g2148) & (!sk[91]) & (g2256) & (g282)) + ((!g2148) & (sk[91]) & (!g2256) & (g282)) + ((!g2148) & (sk[91]) & (g2256) & (g282)) + ((g2148) & (!sk[91]) & (!g2256) & (g282)) + ((g2148) & (!sk[91]) & (g2256) & (!g282)) + ((g2148) & (!sk[91]) & (g2256) & (g282)) + ((g2148) & (sk[91]) & (g2256) & (!g282)) + ((g2148) & (sk[91]) & (g2256) & (g282)));
	assign g4087 = (((!g2153) & (!sk[92]) & (!g2256) & (g283)) + ((!g2153) & (!sk[92]) & (g2256) & (!g283)) + ((!g2153) & (!sk[92]) & (g2256) & (g283)) + ((!g2153) & (sk[92]) & (!g2256) & (g283)) + ((!g2153) & (sk[92]) & (g2256) & (g283)) + ((g2153) & (!sk[92]) & (!g2256) & (g283)) + ((g2153) & (!sk[92]) & (g2256) & (!g283)) + ((g2153) & (!sk[92]) & (g2256) & (g283)) + ((g2153) & (sk[92]) & (g2256) & (!g283)) + ((g2153) & (sk[92]) & (g2256) & (g283)));
	assign g4088 = (((!sk[93]) & (!g2159) & (!g2256) & (g284)) + ((!sk[93]) & (!g2159) & (g2256) & (!g284)) + ((!sk[93]) & (!g2159) & (g2256) & (g284)) + ((!sk[93]) & (g2159) & (!g2256) & (g284)) + ((!sk[93]) & (g2159) & (g2256) & (!g284)) + ((!sk[93]) & (g2159) & (g2256) & (g284)) + ((sk[93]) & (!g2159) & (!g2256) & (g284)) + ((sk[93]) & (!g2159) & (g2256) & (g284)) + ((sk[93]) & (g2159) & (g2256) & (!g284)) + ((sk[93]) & (g2159) & (g2256) & (g284)));
	assign g285 = (((!g281) & (!g282) & (!g283) & (g284) & (g165) & (g166)) + ((!g281) & (!g282) & (g283) & (!g284) & (!g165) & (g166)) + ((!g281) & (!g282) & (g283) & (g284) & (!g165) & (g166)) + ((!g281) & (!g282) & (g283) & (g284) & (g165) & (g166)) + ((!g281) & (g282) & (!g283) & (!g284) & (g165) & (!g166)) + ((!g281) & (g282) & (!g283) & (g284) & (g165) & (!g166)) + ((!g281) & (g282) & (!g283) & (g284) & (g165) & (g166)) + ((!g281) & (g282) & (g283) & (!g284) & (!g165) & (g166)) + ((!g281) & (g282) & (g283) & (!g284) & (g165) & (!g166)) + ((!g281) & (g282) & (g283) & (g284) & (!g165) & (g166)) + ((!g281) & (g282) & (g283) & (g284) & (g165) & (!g166)) + ((!g281) & (g282) & (g283) & (g284) & (g165) & (g166)) + ((g281) & (!g282) & (!g283) & (!g284) & (!g165) & (!g166)) + ((g281) & (!g282) & (!g283) & (g284) & (!g165) & (!g166)) + ((g281) & (!g282) & (!g283) & (g284) & (g165) & (g166)) + ((g281) & (!g282) & (g283) & (!g284) & (!g165) & (!g166)) + ((g281) & (!g282) & (g283) & (!g284) & (!g165) & (g166)) + ((g281) & (!g282) & (g283) & (g284) & (!g165) & (!g166)) + ((g281) & (!g282) & (g283) & (g284) & (!g165) & (g166)) + ((g281) & (!g282) & (g283) & (g284) & (g165) & (g166)) + ((g281) & (g282) & (!g283) & (!g284) & (!g165) & (!g166)) + ((g281) & (g282) & (!g283) & (!g284) & (g165) & (!g166)) + ((g281) & (g282) & (!g283) & (g284) & (!g165) & (!g166)) + ((g281) & (g282) & (!g283) & (g284) & (g165) & (!g166)) + ((g281) & (g282) & (!g283) & (g284) & (g165) & (g166)) + ((g281) & (g282) & (g283) & (!g284) & (!g165) & (!g166)) + ((g281) & (g282) & (g283) & (!g284) & (!g165) & (g166)) + ((g281) & (g282) & (g283) & (!g284) & (g165) & (!g166)) + ((g281) & (g282) & (g283) & (g284) & (!g165) & (!g166)) + ((g281) & (g282) & (g283) & (g284) & (!g165) & (g166)) + ((g281) & (g282) & (g283) & (g284) & (g165) & (!g166)) + ((g281) & (g282) & (g283) & (g284) & (g165) & (g166)));
	assign g4089 = (((!sk[95]) & (!g2144) & (!g2256) & (g286)) + ((!sk[95]) & (!g2144) & (g2256) & (!g286)) + ((!sk[95]) & (!g2144) & (g2256) & (g286)) + ((!sk[95]) & (g2144) & (!g2256) & (g286)) + ((!sk[95]) & (g2144) & (g2256) & (!g286)) + ((!sk[95]) & (g2144) & (g2256) & (g286)) + ((sk[95]) & (!g2144) & (!g2256) & (g286)) + ((sk[95]) & (!g2144) & (g2256) & (g286)) + ((sk[95]) & (g2144) & (g2256) & (!g286)) + ((sk[95]) & (g2144) & (g2256) & (g286)));
	assign g4090 = (((!sk[96]) & (!g2150) & (!g2256) & (g287)) + ((!sk[96]) & (!g2150) & (g2256) & (!g287)) + ((!sk[96]) & (!g2150) & (g2256) & (g287)) + ((!sk[96]) & (g2150) & (!g2256) & (g287)) + ((!sk[96]) & (g2150) & (g2256) & (!g287)) + ((!sk[96]) & (g2150) & (g2256) & (g287)) + ((sk[96]) & (!g2150) & (!g2256) & (g287)) + ((sk[96]) & (!g2150) & (g2256) & (g287)) + ((sk[96]) & (g2150) & (g2256) & (!g287)) + ((sk[96]) & (g2150) & (g2256) & (g287)));
	assign g4091 = (((!sk[97]) & (!g2155) & (!g2256) & (g288)) + ((!sk[97]) & (!g2155) & (g2256) & (!g288)) + ((!sk[97]) & (!g2155) & (g2256) & (g288)) + ((!sk[97]) & (g2155) & (!g2256) & (g288)) + ((!sk[97]) & (g2155) & (g2256) & (!g288)) + ((!sk[97]) & (g2155) & (g2256) & (g288)) + ((sk[97]) & (!g2155) & (!g2256) & (g288)) + ((sk[97]) & (!g2155) & (g2256) & (g288)) + ((sk[97]) & (g2155) & (g2256) & (!g288)) + ((sk[97]) & (g2155) & (g2256) & (g288)));
	assign g4092 = (((!g2160) & (!sk[98]) & (!g2256) & (g289)) + ((!g2160) & (!sk[98]) & (g2256) & (!g289)) + ((!g2160) & (!sk[98]) & (g2256) & (g289)) + ((!g2160) & (sk[98]) & (!g2256) & (g289)) + ((!g2160) & (sk[98]) & (g2256) & (g289)) + ((g2160) & (!sk[98]) & (!g2256) & (g289)) + ((g2160) & (!sk[98]) & (g2256) & (!g289)) + ((g2160) & (!sk[98]) & (g2256) & (g289)) + ((g2160) & (sk[98]) & (g2256) & (!g289)) + ((g2160) & (sk[98]) & (g2256) & (g289)));
	assign g290 = (((!g286) & (!g287) & (!g288) & (g289) & (g165) & (g166)) + ((!g286) & (!g287) & (g288) & (!g289) & (!g165) & (g166)) + ((!g286) & (!g287) & (g288) & (g289) & (!g165) & (g166)) + ((!g286) & (!g287) & (g288) & (g289) & (g165) & (g166)) + ((!g286) & (g287) & (!g288) & (!g289) & (g165) & (!g166)) + ((!g286) & (g287) & (!g288) & (g289) & (g165) & (!g166)) + ((!g286) & (g287) & (!g288) & (g289) & (g165) & (g166)) + ((!g286) & (g287) & (g288) & (!g289) & (!g165) & (g166)) + ((!g286) & (g287) & (g288) & (!g289) & (g165) & (!g166)) + ((!g286) & (g287) & (g288) & (g289) & (!g165) & (g166)) + ((!g286) & (g287) & (g288) & (g289) & (g165) & (!g166)) + ((!g286) & (g287) & (g288) & (g289) & (g165) & (g166)) + ((g286) & (!g287) & (!g288) & (!g289) & (!g165) & (!g166)) + ((g286) & (!g287) & (!g288) & (g289) & (!g165) & (!g166)) + ((g286) & (!g287) & (!g288) & (g289) & (g165) & (g166)) + ((g286) & (!g287) & (g288) & (!g289) & (!g165) & (!g166)) + ((g286) & (!g287) & (g288) & (!g289) & (!g165) & (g166)) + ((g286) & (!g287) & (g288) & (g289) & (!g165) & (!g166)) + ((g286) & (!g287) & (g288) & (g289) & (!g165) & (g166)) + ((g286) & (!g287) & (g288) & (g289) & (g165) & (g166)) + ((g286) & (g287) & (!g288) & (!g289) & (!g165) & (!g166)) + ((g286) & (g287) & (!g288) & (!g289) & (g165) & (!g166)) + ((g286) & (g287) & (!g288) & (g289) & (!g165) & (!g166)) + ((g286) & (g287) & (!g288) & (g289) & (g165) & (!g166)) + ((g286) & (g287) & (!g288) & (g289) & (g165) & (g166)) + ((g286) & (g287) & (g288) & (!g289) & (!g165) & (!g166)) + ((g286) & (g287) & (g288) & (!g289) & (!g165) & (g166)) + ((g286) & (g287) & (g288) & (!g289) & (g165) & (!g166)) + ((g286) & (g287) & (g288) & (g289) & (!g165) & (!g166)) + ((g286) & (g287) & (g288) & (g289) & (!g165) & (g166)) + ((g286) & (g287) & (g288) & (g289) & (g165) & (!g166)) + ((g286) & (g287) & (g288) & (g289) & (g165) & (g166)));
	assign g4093 = (((!g2145) & (!sk[100]) & (!g2256) & (g291)) + ((!g2145) & (!sk[100]) & (g2256) & (!g291)) + ((!g2145) & (!sk[100]) & (g2256) & (g291)) + ((!g2145) & (sk[100]) & (!g2256) & (g291)) + ((!g2145) & (sk[100]) & (g2256) & (g291)) + ((g2145) & (!sk[100]) & (!g2256) & (g291)) + ((g2145) & (!sk[100]) & (g2256) & (!g291)) + ((g2145) & (!sk[100]) & (g2256) & (g291)) + ((g2145) & (sk[100]) & (g2256) & (!g291)) + ((g2145) & (sk[100]) & (g2256) & (g291)));
	assign g4094 = (((!sk[101]) & (!g2151) & (!g2256) & (g292)) + ((!sk[101]) & (!g2151) & (g2256) & (!g292)) + ((!sk[101]) & (!g2151) & (g2256) & (g292)) + ((!sk[101]) & (g2151) & (!g2256) & (g292)) + ((!sk[101]) & (g2151) & (g2256) & (!g292)) + ((!sk[101]) & (g2151) & (g2256) & (g292)) + ((sk[101]) & (!g2151) & (!g2256) & (g292)) + ((sk[101]) & (!g2151) & (g2256) & (g292)) + ((sk[101]) & (g2151) & (g2256) & (!g292)) + ((sk[101]) & (g2151) & (g2256) & (g292)));
	assign g4095 = (((!sk[102]) & (!g2157) & (!g2256) & (g293)) + ((!sk[102]) & (!g2157) & (g2256) & (!g293)) + ((!sk[102]) & (!g2157) & (g2256) & (g293)) + ((!sk[102]) & (g2157) & (!g2256) & (g293)) + ((!sk[102]) & (g2157) & (g2256) & (!g293)) + ((!sk[102]) & (g2157) & (g2256) & (g293)) + ((sk[102]) & (!g2157) & (!g2256) & (g293)) + ((sk[102]) & (!g2157) & (g2256) & (g293)) + ((sk[102]) & (g2157) & (g2256) & (!g293)) + ((sk[102]) & (g2157) & (g2256) & (g293)));
	assign g4096 = (((!g2161) & (!sk[103]) & (!g2256) & (g294)) + ((!g2161) & (!sk[103]) & (g2256) & (!g294)) + ((!g2161) & (!sk[103]) & (g2256) & (g294)) + ((!g2161) & (sk[103]) & (!g2256) & (g294)) + ((!g2161) & (sk[103]) & (g2256) & (g294)) + ((g2161) & (!sk[103]) & (!g2256) & (g294)) + ((g2161) & (!sk[103]) & (g2256) & (!g294)) + ((g2161) & (!sk[103]) & (g2256) & (g294)) + ((g2161) & (sk[103]) & (g2256) & (!g294)) + ((g2161) & (sk[103]) & (g2256) & (g294)));
	assign g295 = (((!g291) & (!g292) & (!g293) & (g294) & (g165) & (g166)) + ((!g291) & (!g292) & (g293) & (!g294) & (!g165) & (g166)) + ((!g291) & (!g292) & (g293) & (g294) & (!g165) & (g166)) + ((!g291) & (!g292) & (g293) & (g294) & (g165) & (g166)) + ((!g291) & (g292) & (!g293) & (!g294) & (g165) & (!g166)) + ((!g291) & (g292) & (!g293) & (g294) & (g165) & (!g166)) + ((!g291) & (g292) & (!g293) & (g294) & (g165) & (g166)) + ((!g291) & (g292) & (g293) & (!g294) & (!g165) & (g166)) + ((!g291) & (g292) & (g293) & (!g294) & (g165) & (!g166)) + ((!g291) & (g292) & (g293) & (g294) & (!g165) & (g166)) + ((!g291) & (g292) & (g293) & (g294) & (g165) & (!g166)) + ((!g291) & (g292) & (g293) & (g294) & (g165) & (g166)) + ((g291) & (!g292) & (!g293) & (!g294) & (!g165) & (!g166)) + ((g291) & (!g292) & (!g293) & (g294) & (!g165) & (!g166)) + ((g291) & (!g292) & (!g293) & (g294) & (g165) & (g166)) + ((g291) & (!g292) & (g293) & (!g294) & (!g165) & (!g166)) + ((g291) & (!g292) & (g293) & (!g294) & (!g165) & (g166)) + ((g291) & (!g292) & (g293) & (g294) & (!g165) & (!g166)) + ((g291) & (!g292) & (g293) & (g294) & (!g165) & (g166)) + ((g291) & (!g292) & (g293) & (g294) & (g165) & (g166)) + ((g291) & (g292) & (!g293) & (!g294) & (!g165) & (!g166)) + ((g291) & (g292) & (!g293) & (!g294) & (g165) & (!g166)) + ((g291) & (g292) & (!g293) & (g294) & (!g165) & (!g166)) + ((g291) & (g292) & (!g293) & (g294) & (g165) & (!g166)) + ((g291) & (g292) & (!g293) & (g294) & (g165) & (g166)) + ((g291) & (g292) & (g293) & (!g294) & (!g165) & (!g166)) + ((g291) & (g292) & (g293) & (!g294) & (!g165) & (g166)) + ((g291) & (g292) & (g293) & (!g294) & (g165) & (!g166)) + ((g291) & (g292) & (g293) & (g294) & (!g165) & (!g166)) + ((g291) & (g292) & (g293) & (g294) & (!g165) & (g166)) + ((g291) & (g292) & (g293) & (g294) & (g165) & (!g166)) + ((g291) & (g292) & (g293) & (g294) & (g165) & (g166)));
	assign g296 = (((!g280) & (!g285) & (!g290) & (g295) & (g147) & (g148)) + ((!g280) & (!g285) & (g290) & (!g295) & (!g147) & (g148)) + ((!g280) & (!g285) & (g290) & (g295) & (!g147) & (g148)) + ((!g280) & (!g285) & (g290) & (g295) & (g147) & (g148)) + ((!g280) & (g285) & (!g290) & (!g295) & (g147) & (!g148)) + ((!g280) & (g285) & (!g290) & (g295) & (g147) & (!g148)) + ((!g280) & (g285) & (!g290) & (g295) & (g147) & (g148)) + ((!g280) & (g285) & (g290) & (!g295) & (!g147) & (g148)) + ((!g280) & (g285) & (g290) & (!g295) & (g147) & (!g148)) + ((!g280) & (g285) & (g290) & (g295) & (!g147) & (g148)) + ((!g280) & (g285) & (g290) & (g295) & (g147) & (!g148)) + ((!g280) & (g285) & (g290) & (g295) & (g147) & (g148)) + ((g280) & (!g285) & (!g290) & (!g295) & (!g147) & (!g148)) + ((g280) & (!g285) & (!g290) & (g295) & (!g147) & (!g148)) + ((g280) & (!g285) & (!g290) & (g295) & (g147) & (g148)) + ((g280) & (!g285) & (g290) & (!g295) & (!g147) & (!g148)) + ((g280) & (!g285) & (g290) & (!g295) & (!g147) & (g148)) + ((g280) & (!g285) & (g290) & (g295) & (!g147) & (!g148)) + ((g280) & (!g285) & (g290) & (g295) & (!g147) & (g148)) + ((g280) & (!g285) & (g290) & (g295) & (g147) & (g148)) + ((g280) & (g285) & (!g290) & (!g295) & (!g147) & (!g148)) + ((g280) & (g285) & (!g290) & (!g295) & (g147) & (!g148)) + ((g280) & (g285) & (!g290) & (g295) & (!g147) & (!g148)) + ((g280) & (g285) & (!g290) & (g295) & (g147) & (!g148)) + ((g280) & (g285) & (!g290) & (g295) & (g147) & (g148)) + ((g280) & (g285) & (g290) & (!g295) & (!g147) & (!g148)) + ((g280) & (g285) & (g290) & (!g295) & (!g147) & (g148)) + ((g280) & (g285) & (g290) & (!g295) & (g147) & (!g148)) + ((g280) & (g285) & (g290) & (g295) & (!g147) & (!g148)) + ((g280) & (g285) & (g290) & (g295) & (!g147) & (g148)) + ((g280) & (g285) & (g290) & (g295) & (g147) & (!g148)) + ((g280) & (g285) & (g290) & (g295) & (g147) & (g148)));
	assign g4097 = (((!g2173) & (!sk[106]) & (!g2256) & (g297)) + ((!g2173) & (!sk[106]) & (g2256) & (!g297)) + ((!g2173) & (!sk[106]) & (g2256) & (g297)) + ((!g2173) & (sk[106]) & (!g2256) & (g297)) + ((!g2173) & (sk[106]) & (g2256) & (g297)) + ((g2173) & (!sk[106]) & (!g2256) & (g297)) + ((g2173) & (!sk[106]) & (g2256) & (!g297)) + ((g2173) & (!sk[106]) & (g2256) & (g297)) + ((g2173) & (sk[106]) & (g2256) & (!g297)) + ((g2173) & (sk[106]) & (g2256) & (g297)));
	assign g4098 = (((!g2174) & (!g2256) & (!sk[107]) & (g298)) + ((!g2174) & (!g2256) & (sk[107]) & (g298)) + ((!g2174) & (g2256) & (!sk[107]) & (!g298)) + ((!g2174) & (g2256) & (!sk[107]) & (g298)) + ((!g2174) & (g2256) & (sk[107]) & (g298)) + ((g2174) & (!g2256) & (!sk[107]) & (g298)) + ((g2174) & (g2256) & (!sk[107]) & (!g298)) + ((g2174) & (g2256) & (!sk[107]) & (g298)) + ((g2174) & (g2256) & (sk[107]) & (!g298)) + ((g2174) & (g2256) & (sk[107]) & (g298)));
	assign g4099 = (((!g2175) & (!sk[108]) & (!g2256) & (g299)) + ((!g2175) & (!sk[108]) & (g2256) & (!g299)) + ((!g2175) & (!sk[108]) & (g2256) & (g299)) + ((!g2175) & (sk[108]) & (!g2256) & (g299)) + ((!g2175) & (sk[108]) & (g2256) & (g299)) + ((g2175) & (!sk[108]) & (!g2256) & (g299)) + ((g2175) & (!sk[108]) & (g2256) & (!g299)) + ((g2175) & (!sk[108]) & (g2256) & (g299)) + ((g2175) & (sk[108]) & (g2256) & (!g299)) + ((g2175) & (sk[108]) & (g2256) & (g299)));
	assign g4100 = (((!g2176) & (!g2256) & (!sk[109]) & (g300)) + ((!g2176) & (!g2256) & (sk[109]) & (g300)) + ((!g2176) & (g2256) & (!sk[109]) & (!g300)) + ((!g2176) & (g2256) & (!sk[109]) & (g300)) + ((!g2176) & (g2256) & (sk[109]) & (g300)) + ((g2176) & (!g2256) & (!sk[109]) & (g300)) + ((g2176) & (g2256) & (!sk[109]) & (!g300)) + ((g2176) & (g2256) & (!sk[109]) & (g300)) + ((g2176) & (g2256) & (sk[109]) & (!g300)) + ((g2176) & (g2256) & (sk[109]) & (g300)));
	assign g301 = (((!g297) & (!g298) & (!g299) & (g300) & (g165) & (g166)) + ((!g297) & (!g298) & (g299) & (!g300) & (!g165) & (g166)) + ((!g297) & (!g298) & (g299) & (g300) & (!g165) & (g166)) + ((!g297) & (!g298) & (g299) & (g300) & (g165) & (g166)) + ((!g297) & (g298) & (!g299) & (!g300) & (g165) & (!g166)) + ((!g297) & (g298) & (!g299) & (g300) & (g165) & (!g166)) + ((!g297) & (g298) & (!g299) & (g300) & (g165) & (g166)) + ((!g297) & (g298) & (g299) & (!g300) & (!g165) & (g166)) + ((!g297) & (g298) & (g299) & (!g300) & (g165) & (!g166)) + ((!g297) & (g298) & (g299) & (g300) & (!g165) & (g166)) + ((!g297) & (g298) & (g299) & (g300) & (g165) & (!g166)) + ((!g297) & (g298) & (g299) & (g300) & (g165) & (g166)) + ((g297) & (!g298) & (!g299) & (!g300) & (!g165) & (!g166)) + ((g297) & (!g298) & (!g299) & (g300) & (!g165) & (!g166)) + ((g297) & (!g298) & (!g299) & (g300) & (g165) & (g166)) + ((g297) & (!g298) & (g299) & (!g300) & (!g165) & (!g166)) + ((g297) & (!g298) & (g299) & (!g300) & (!g165) & (g166)) + ((g297) & (!g298) & (g299) & (g300) & (!g165) & (!g166)) + ((g297) & (!g298) & (g299) & (g300) & (!g165) & (g166)) + ((g297) & (!g298) & (g299) & (g300) & (g165) & (g166)) + ((g297) & (g298) & (!g299) & (!g300) & (!g165) & (!g166)) + ((g297) & (g298) & (!g299) & (!g300) & (g165) & (!g166)) + ((g297) & (g298) & (!g299) & (g300) & (!g165) & (!g166)) + ((g297) & (g298) & (!g299) & (g300) & (g165) & (!g166)) + ((g297) & (g298) & (!g299) & (g300) & (g165) & (g166)) + ((g297) & (g298) & (g299) & (!g300) & (!g165) & (!g166)) + ((g297) & (g298) & (g299) & (!g300) & (!g165) & (g166)) + ((g297) & (g298) & (g299) & (!g300) & (g165) & (!g166)) + ((g297) & (g298) & (g299) & (g300) & (!g165) & (!g166)) + ((g297) & (g298) & (g299) & (g300) & (!g165) & (g166)) + ((g297) & (g298) & (g299) & (g300) & (g165) & (!g166)) + ((g297) & (g298) & (g299) & (g300) & (g165) & (g166)));
	assign g4101 = (((!sk[111]) & (!g2177) & (!g2256) & (g302)) + ((!sk[111]) & (!g2177) & (g2256) & (!g302)) + ((!sk[111]) & (!g2177) & (g2256) & (g302)) + ((!sk[111]) & (g2177) & (!g2256) & (g302)) + ((!sk[111]) & (g2177) & (g2256) & (!g302)) + ((!sk[111]) & (g2177) & (g2256) & (g302)) + ((sk[111]) & (!g2177) & (!g2256) & (g302)) + ((sk[111]) & (!g2177) & (g2256) & (g302)) + ((sk[111]) & (g2177) & (g2256) & (!g302)) + ((sk[111]) & (g2177) & (g2256) & (g302)));
	assign g4102 = (((!sk[112]) & (!g2178) & (!g2256) & (g303)) + ((!sk[112]) & (!g2178) & (g2256) & (!g303)) + ((!sk[112]) & (!g2178) & (g2256) & (g303)) + ((!sk[112]) & (g2178) & (!g2256) & (g303)) + ((!sk[112]) & (g2178) & (g2256) & (!g303)) + ((!sk[112]) & (g2178) & (g2256) & (g303)) + ((sk[112]) & (!g2178) & (!g2256) & (g303)) + ((sk[112]) & (!g2178) & (g2256) & (g303)) + ((sk[112]) & (g2178) & (g2256) & (!g303)) + ((sk[112]) & (g2178) & (g2256) & (g303)));
	assign g4103 = (((!sk[113]) & (!g2179) & (!g2256) & (g304)) + ((!sk[113]) & (!g2179) & (g2256) & (!g304)) + ((!sk[113]) & (!g2179) & (g2256) & (g304)) + ((!sk[113]) & (g2179) & (!g2256) & (g304)) + ((!sk[113]) & (g2179) & (g2256) & (!g304)) + ((!sk[113]) & (g2179) & (g2256) & (g304)) + ((sk[113]) & (!g2179) & (!g2256) & (g304)) + ((sk[113]) & (!g2179) & (g2256) & (g304)) + ((sk[113]) & (g2179) & (g2256) & (!g304)) + ((sk[113]) & (g2179) & (g2256) & (g304)));
	assign g305 = (((!g165) & (!g166) & (!sk[114]) & (!g302) & (g303) & (!g304)) + ((!g165) & (!g166) & (!sk[114]) & (!g302) & (g303) & (g304)) + ((!g165) & (!g166) & (!sk[114]) & (g302) & (!g303) & (!g304)) + ((!g165) & (!g166) & (!sk[114]) & (g302) & (!g303) & (g304)) + ((!g165) & (!g166) & (!sk[114]) & (g302) & (g303) & (!g304)) + ((!g165) & (!g166) & (!sk[114]) & (g302) & (g303) & (g304)) + ((!g165) & (g166) & (!sk[114]) & (!g302) & (!g303) & (!g304)) + ((!g165) & (g166) & (!sk[114]) & (!g302) & (!g303) & (g304)) + ((!g165) & (g166) & (!sk[114]) & (!g302) & (g303) & (!g304)) + ((!g165) & (g166) & (!sk[114]) & (!g302) & (g303) & (g304)) + ((!g165) & (g166) & (!sk[114]) & (g302) & (!g303) & (!g304)) + ((!g165) & (g166) & (!sk[114]) & (g302) & (!g303) & (g304)) + ((!g165) & (g166) & (!sk[114]) & (g302) & (g303) & (!g304)) + ((!g165) & (g166) & (!sk[114]) & (g302) & (g303) & (g304)) + ((!g165) & (g166) & (sk[114]) & (!g302) & (!g303) & (g304)) + ((!g165) & (g166) & (sk[114]) & (!g302) & (g303) & (g304)) + ((!g165) & (g166) & (sk[114]) & (g302) & (!g303) & (g304)) + ((!g165) & (g166) & (sk[114]) & (g302) & (g303) & (g304)) + ((g165) & (!g166) & (!sk[114]) & (!g302) & (g303) & (!g304)) + ((g165) & (!g166) & (!sk[114]) & (!g302) & (g303) & (g304)) + ((g165) & (!g166) & (!sk[114]) & (g302) & (!g303) & (!g304)) + ((g165) & (!g166) & (!sk[114]) & (g302) & (!g303) & (g304)) + ((g165) & (!g166) & (!sk[114]) & (g302) & (g303) & (!g304)) + ((g165) & (!g166) & (!sk[114]) & (g302) & (g303) & (g304)) + ((g165) & (!g166) & (sk[114]) & (g302) & (!g303) & (!g304)) + ((g165) & (!g166) & (sk[114]) & (g302) & (!g303) & (g304)) + ((g165) & (!g166) & (sk[114]) & (g302) & (g303) & (!g304)) + ((g165) & (!g166) & (sk[114]) & (g302) & (g303) & (g304)) + ((g165) & (g166) & (!sk[114]) & (!g302) & (!g303) & (!g304)) + ((g165) & (g166) & (!sk[114]) & (!g302) & (!g303) & (g304)) + ((g165) & (g166) & (!sk[114]) & (!g302) & (g303) & (!g304)) + ((g165) & (g166) & (!sk[114]) & (!g302) & (g303) & (g304)) + ((g165) & (g166) & (!sk[114]) & (g302) & (!g303) & (!g304)) + ((g165) & (g166) & (!sk[114]) & (g302) & (!g303) & (g304)) + ((g165) & (g166) & (!sk[114]) & (g302) & (g303) & (!g304)) + ((g165) & (g166) & (!sk[114]) & (g302) & (g303) & (g304)) + ((g165) & (g166) & (sk[114]) & (!g302) & (g303) & (!g304)) + ((g165) & (g166) & (sk[114]) & (!g302) & (g303) & (g304)) + ((g165) & (g166) & (sk[114]) & (g302) & (g303) & (!g304)) + ((g165) & (g166) & (sk[114]) & (g302) & (g303) & (g304)));
	assign g4104 = (((!sk[115]) & (!g2162) & (!g2256) & (g306)) + ((!sk[115]) & (!g2162) & (g2256) & (!g306)) + ((!sk[115]) & (!g2162) & (g2256) & (g306)) + ((!sk[115]) & (g2162) & (!g2256) & (g306)) + ((!sk[115]) & (g2162) & (g2256) & (!g306)) + ((!sk[115]) & (g2162) & (g2256) & (g306)) + ((sk[115]) & (!g2162) & (!g2256) & (g306)) + ((sk[115]) & (!g2162) & (g2256) & (g306)) + ((sk[115]) & (g2162) & (g2256) & (!g306)) + ((sk[115]) & (g2162) & (g2256) & (g306)));
	assign g4105 = (((!g2164) & (!g2256) & (!sk[116]) & (g307)) + ((!g2164) & (!g2256) & (sk[116]) & (g307)) + ((!g2164) & (g2256) & (!sk[116]) & (!g307)) + ((!g2164) & (g2256) & (!sk[116]) & (g307)) + ((!g2164) & (g2256) & (sk[116]) & (g307)) + ((g2164) & (!g2256) & (!sk[116]) & (g307)) + ((g2164) & (g2256) & (!sk[116]) & (!g307)) + ((g2164) & (g2256) & (!sk[116]) & (g307)) + ((g2164) & (g2256) & (sk[116]) & (!g307)) + ((g2164) & (g2256) & (sk[116]) & (g307)));
	assign g4106 = (((!g2166) & (!sk[117]) & (!g2256) & (g308)) + ((!g2166) & (!sk[117]) & (g2256) & (!g308)) + ((!g2166) & (!sk[117]) & (g2256) & (g308)) + ((!g2166) & (sk[117]) & (!g2256) & (g308)) + ((!g2166) & (sk[117]) & (g2256) & (g308)) + ((g2166) & (!sk[117]) & (!g2256) & (g308)) + ((g2166) & (!sk[117]) & (g2256) & (!g308)) + ((g2166) & (!sk[117]) & (g2256) & (g308)) + ((g2166) & (sk[117]) & (g2256) & (!g308)) + ((g2166) & (sk[117]) & (g2256) & (g308)));
	assign g4107 = (((!g2168) & (!sk[118]) & (!g2256) & (g309)) + ((!g2168) & (!sk[118]) & (g2256) & (!g309)) + ((!g2168) & (!sk[118]) & (g2256) & (g309)) + ((!g2168) & (sk[118]) & (!g2256) & (g309)) + ((!g2168) & (sk[118]) & (g2256) & (g309)) + ((g2168) & (!sk[118]) & (!g2256) & (g309)) + ((g2168) & (!sk[118]) & (g2256) & (!g309)) + ((g2168) & (!sk[118]) & (g2256) & (g309)) + ((g2168) & (sk[118]) & (g2256) & (!g309)) + ((g2168) & (sk[118]) & (g2256) & (g309)));
	assign g310 = (((!g306) & (!g307) & (!g308) & (g309) & (g165) & (g166)) + ((!g306) & (!g307) & (g308) & (!g309) & (!g165) & (g166)) + ((!g306) & (!g307) & (g308) & (g309) & (!g165) & (g166)) + ((!g306) & (!g307) & (g308) & (g309) & (g165) & (g166)) + ((!g306) & (g307) & (!g308) & (!g309) & (g165) & (!g166)) + ((!g306) & (g307) & (!g308) & (g309) & (g165) & (!g166)) + ((!g306) & (g307) & (!g308) & (g309) & (g165) & (g166)) + ((!g306) & (g307) & (g308) & (!g309) & (!g165) & (g166)) + ((!g306) & (g307) & (g308) & (!g309) & (g165) & (!g166)) + ((!g306) & (g307) & (g308) & (g309) & (!g165) & (g166)) + ((!g306) & (g307) & (g308) & (g309) & (g165) & (!g166)) + ((!g306) & (g307) & (g308) & (g309) & (g165) & (g166)) + ((g306) & (!g307) & (!g308) & (!g309) & (!g165) & (!g166)) + ((g306) & (!g307) & (!g308) & (g309) & (!g165) & (!g166)) + ((g306) & (!g307) & (!g308) & (g309) & (g165) & (g166)) + ((g306) & (!g307) & (g308) & (!g309) & (!g165) & (!g166)) + ((g306) & (!g307) & (g308) & (!g309) & (!g165) & (g166)) + ((g306) & (!g307) & (g308) & (g309) & (!g165) & (!g166)) + ((g306) & (!g307) & (g308) & (g309) & (!g165) & (g166)) + ((g306) & (!g307) & (g308) & (g309) & (g165) & (g166)) + ((g306) & (g307) & (!g308) & (!g309) & (!g165) & (!g166)) + ((g306) & (g307) & (!g308) & (!g309) & (g165) & (!g166)) + ((g306) & (g307) & (!g308) & (g309) & (!g165) & (!g166)) + ((g306) & (g307) & (!g308) & (g309) & (g165) & (!g166)) + ((g306) & (g307) & (!g308) & (g309) & (g165) & (g166)) + ((g306) & (g307) & (g308) & (!g309) & (!g165) & (!g166)) + ((g306) & (g307) & (g308) & (!g309) & (!g165) & (g166)) + ((g306) & (g307) & (g308) & (!g309) & (g165) & (!g166)) + ((g306) & (g307) & (g308) & (g309) & (!g165) & (!g166)) + ((g306) & (g307) & (g308) & (g309) & (!g165) & (g166)) + ((g306) & (g307) & (g308) & (g309) & (g165) & (!g166)) + ((g306) & (g307) & (g308) & (g309) & (g165) & (g166)));
	assign g4108 = (((!g2169) & (!g2256) & (!sk[120]) & (g311)) + ((!g2169) & (!g2256) & (sk[120]) & (g311)) + ((!g2169) & (g2256) & (!sk[120]) & (!g311)) + ((!g2169) & (g2256) & (!sk[120]) & (g311)) + ((!g2169) & (g2256) & (sk[120]) & (g311)) + ((g2169) & (!g2256) & (!sk[120]) & (g311)) + ((g2169) & (g2256) & (!sk[120]) & (!g311)) + ((g2169) & (g2256) & (!sk[120]) & (g311)) + ((g2169) & (g2256) & (sk[120]) & (!g311)) + ((g2169) & (g2256) & (sk[120]) & (g311)));
	assign g4109 = (((!g2170) & (!g2256) & (!sk[121]) & (g312)) + ((!g2170) & (!g2256) & (sk[121]) & (g312)) + ((!g2170) & (g2256) & (!sk[121]) & (!g312)) + ((!g2170) & (g2256) & (!sk[121]) & (g312)) + ((!g2170) & (g2256) & (sk[121]) & (g312)) + ((g2170) & (!g2256) & (!sk[121]) & (g312)) + ((g2170) & (g2256) & (!sk[121]) & (!g312)) + ((g2170) & (g2256) & (!sk[121]) & (g312)) + ((g2170) & (g2256) & (sk[121]) & (!g312)) + ((g2170) & (g2256) & (sk[121]) & (g312)));
	assign g4110 = (((!g2171) & (!g2256) & (!sk[122]) & (g313)) + ((!g2171) & (!g2256) & (sk[122]) & (g313)) + ((!g2171) & (g2256) & (!sk[122]) & (!g313)) + ((!g2171) & (g2256) & (!sk[122]) & (g313)) + ((!g2171) & (g2256) & (sk[122]) & (g313)) + ((g2171) & (!g2256) & (!sk[122]) & (g313)) + ((g2171) & (g2256) & (!sk[122]) & (!g313)) + ((g2171) & (g2256) & (!sk[122]) & (g313)) + ((g2171) & (g2256) & (sk[122]) & (!g313)) + ((g2171) & (g2256) & (sk[122]) & (g313)));
	assign g4111 = (((!g2172) & (!g2256) & (!sk[123]) & (g314)) + ((!g2172) & (!g2256) & (sk[123]) & (g314)) + ((!g2172) & (g2256) & (!sk[123]) & (!g314)) + ((!g2172) & (g2256) & (!sk[123]) & (g314)) + ((!g2172) & (g2256) & (sk[123]) & (g314)) + ((g2172) & (!g2256) & (!sk[123]) & (g314)) + ((g2172) & (g2256) & (!sk[123]) & (!g314)) + ((g2172) & (g2256) & (!sk[123]) & (g314)) + ((g2172) & (g2256) & (sk[123]) & (!g314)) + ((g2172) & (g2256) & (sk[123]) & (g314)));
	assign g315 = (((!g311) & (!g312) & (!g313) & (g314) & (g165) & (g166)) + ((!g311) & (!g312) & (g313) & (!g314) & (!g165) & (g166)) + ((!g311) & (!g312) & (g313) & (g314) & (!g165) & (g166)) + ((!g311) & (!g312) & (g313) & (g314) & (g165) & (g166)) + ((!g311) & (g312) & (!g313) & (!g314) & (g165) & (!g166)) + ((!g311) & (g312) & (!g313) & (g314) & (g165) & (!g166)) + ((!g311) & (g312) & (!g313) & (g314) & (g165) & (g166)) + ((!g311) & (g312) & (g313) & (!g314) & (!g165) & (g166)) + ((!g311) & (g312) & (g313) & (!g314) & (g165) & (!g166)) + ((!g311) & (g312) & (g313) & (g314) & (!g165) & (g166)) + ((!g311) & (g312) & (g313) & (g314) & (g165) & (!g166)) + ((!g311) & (g312) & (g313) & (g314) & (g165) & (g166)) + ((g311) & (!g312) & (!g313) & (!g314) & (!g165) & (!g166)) + ((g311) & (!g312) & (!g313) & (g314) & (!g165) & (!g166)) + ((g311) & (!g312) & (!g313) & (g314) & (g165) & (g166)) + ((g311) & (!g312) & (g313) & (!g314) & (!g165) & (!g166)) + ((g311) & (!g312) & (g313) & (!g314) & (!g165) & (g166)) + ((g311) & (!g312) & (g313) & (g314) & (!g165) & (!g166)) + ((g311) & (!g312) & (g313) & (g314) & (!g165) & (g166)) + ((g311) & (!g312) & (g313) & (g314) & (g165) & (g166)) + ((g311) & (g312) & (!g313) & (!g314) & (!g165) & (!g166)) + ((g311) & (g312) & (!g313) & (!g314) & (g165) & (!g166)) + ((g311) & (g312) & (!g313) & (g314) & (!g165) & (!g166)) + ((g311) & (g312) & (!g313) & (g314) & (g165) & (!g166)) + ((g311) & (g312) & (!g313) & (g314) & (g165) & (g166)) + ((g311) & (g312) & (g313) & (!g314) & (!g165) & (!g166)) + ((g311) & (g312) & (g313) & (!g314) & (!g165) & (g166)) + ((g311) & (g312) & (g313) & (!g314) & (g165) & (!g166)) + ((g311) & (g312) & (g313) & (g314) & (!g165) & (!g166)) + ((g311) & (g312) & (g313) & (g314) & (!g165) & (g166)) + ((g311) & (g312) & (g313) & (g314) & (g165) & (!g166)) + ((g311) & (g312) & (g313) & (g314) & (g165) & (g166)));
	assign g316 = (((!g147) & (!g148) & (!g301) & (g305) & (!g310) & (!g315)) + ((!g147) & (!g148) & (!g301) & (g305) & (!g310) & (g315)) + ((!g147) & (!g148) & (!g301) & (g305) & (g310) & (!g315)) + ((!g147) & (!g148) & (!g301) & (g305) & (g310) & (g315)) + ((!g147) & (!g148) & (g301) & (g305) & (!g310) & (!g315)) + ((!g147) & (!g148) & (g301) & (g305) & (!g310) & (g315)) + ((!g147) & (!g148) & (g301) & (g305) & (g310) & (!g315)) + ((!g147) & (!g148) & (g301) & (g305) & (g310) & (g315)) + ((!g147) & (g148) & (!g301) & (!g305) & (!g310) & (g315)) + ((!g147) & (g148) & (!g301) & (!g305) & (g310) & (g315)) + ((!g147) & (g148) & (!g301) & (g305) & (!g310) & (g315)) + ((!g147) & (g148) & (!g301) & (g305) & (g310) & (g315)) + ((!g147) & (g148) & (g301) & (!g305) & (!g310) & (g315)) + ((!g147) & (g148) & (g301) & (!g305) & (g310) & (g315)) + ((!g147) & (g148) & (g301) & (g305) & (!g310) & (g315)) + ((!g147) & (g148) & (g301) & (g305) & (g310) & (g315)) + ((g147) & (!g148) & (g301) & (!g305) & (!g310) & (!g315)) + ((g147) & (!g148) & (g301) & (!g305) & (!g310) & (g315)) + ((g147) & (!g148) & (g301) & (!g305) & (g310) & (!g315)) + ((g147) & (!g148) & (g301) & (!g305) & (g310) & (g315)) + ((g147) & (!g148) & (g301) & (g305) & (!g310) & (!g315)) + ((g147) & (!g148) & (g301) & (g305) & (!g310) & (g315)) + ((g147) & (!g148) & (g301) & (g305) & (g310) & (!g315)) + ((g147) & (!g148) & (g301) & (g305) & (g310) & (g315)) + ((g147) & (g148) & (!g301) & (!g305) & (g310) & (!g315)) + ((g147) & (g148) & (!g301) & (!g305) & (g310) & (g315)) + ((g147) & (g148) & (!g301) & (g305) & (g310) & (!g315)) + ((g147) & (g148) & (!g301) & (g305) & (g310) & (g315)) + ((g147) & (g148) & (g301) & (!g305) & (g310) & (!g315)) + ((g147) & (g148) & (g301) & (!g305) & (g310) & (g315)) + ((g147) & (g148) & (g301) & (g305) & (g310) & (!g315)) + ((g147) & (g148) & (g301) & (g305) & (g310) & (g315)));
	assign g317 = (((!sk[126]) & (!g142) & (!g296) & (g316)) + ((!sk[126]) & (!g142) & (g296) & (!g316)) + ((!sk[126]) & (!g142) & (g296) & (g316)) + ((!sk[126]) & (g142) & (!g296) & (g316)) + ((!sk[126]) & (g142) & (g296) & (!g316)) + ((!sk[126]) & (g142) & (g296) & (g316)) + ((sk[126]) & (!g142) & (!g296) & (g316)) + ((sk[126]) & (!g142) & (g296) & (g316)) + ((sk[126]) & (g142) & (g296) & (!g316)) + ((sk[126]) & (g142) & (g296) & (g316)));
	assign g4112 = (((!g2064) & (!dmem_dat_ix4x) & (!sk[127]) & (g318)) + ((!g2064) & (!dmem_dat_ix4x) & (sk[127]) & (g318)) + ((!g2064) & (dmem_dat_ix4x) & (!sk[127]) & (!g318)) + ((!g2064) & (dmem_dat_ix4x) & (!sk[127]) & (g318)) + ((!g2064) & (dmem_dat_ix4x) & (sk[127]) & (g318)) + ((g2064) & (!dmem_dat_ix4x) & (!sk[127]) & (g318)) + ((g2064) & (dmem_dat_ix4x) & (!sk[127]) & (!g318)) + ((g2064) & (dmem_dat_ix4x) & (!sk[127]) & (g318)) + ((g2064) & (dmem_dat_ix4x) & (sk[127]) & (!g318)) + ((g2064) & (dmem_dat_ix4x) & (sk[127]) & (g318)));
	assign g4113 = (((!g2059) & (!sk[0]) & (!g2263) & (g319)) + ((!g2059) & (!sk[0]) & (g2263) & (!g319)) + ((!g2059) & (!sk[0]) & (g2263) & (g319)) + ((!g2059) & (sk[0]) & (!g2263) & (g319)) + ((!g2059) & (sk[0]) & (g2263) & (g319)) + ((g2059) & (!sk[0]) & (!g2263) & (g319)) + ((g2059) & (!sk[0]) & (g2263) & (!g319)) + ((g2059) & (!sk[0]) & (g2263) & (g319)) + ((g2059) & (sk[0]) & (g2263) & (!g319)) + ((g2059) & (sk[0]) & (g2263) & (g319)));
	assign g320 = (((!g87) & (!sk[1]) & (!g90) & (!g231) & (g273) & (!g317)) + ((!g87) & (!sk[1]) & (!g90) & (!g231) & (g273) & (g317)) + ((!g87) & (!sk[1]) & (!g90) & (g231) & (!g273) & (!g317)) + ((!g87) & (!sk[1]) & (!g90) & (g231) & (!g273) & (g317)) + ((!g87) & (!sk[1]) & (!g90) & (g231) & (g273) & (!g317)) + ((!g87) & (!sk[1]) & (!g90) & (g231) & (g273) & (g317)) + ((!g87) & (!sk[1]) & (g90) & (!g231) & (!g273) & (!g317)) + ((!g87) & (!sk[1]) & (g90) & (!g231) & (!g273) & (g317)) + ((!g87) & (!sk[1]) & (g90) & (!g231) & (g273) & (!g317)) + ((!g87) & (!sk[1]) & (g90) & (!g231) & (g273) & (g317)) + ((!g87) & (!sk[1]) & (g90) & (g231) & (!g273) & (!g317)) + ((!g87) & (!sk[1]) & (g90) & (g231) & (!g273) & (g317)) + ((!g87) & (!sk[1]) & (g90) & (g231) & (g273) & (!g317)) + ((!g87) & (!sk[1]) & (g90) & (g231) & (g273) & (g317)) + ((!g87) & (sk[1]) & (!g90) & (g231) & (g273) & (g317)) + ((!g87) & (sk[1]) & (g90) & (!g231) & (!g273) & (g317)) + ((!g87) & (sk[1]) & (g90) & (!g231) & (g273) & (g317)) + ((!g87) & (sk[1]) & (g90) & (g231) & (!g273) & (g317)) + ((!g87) & (sk[1]) & (g90) & (g231) & (g273) & (!g317)) + ((!g87) & (sk[1]) & (g90) & (g231) & (g273) & (g317)) + ((g87) & (!sk[1]) & (!g90) & (!g231) & (g273) & (!g317)) + ((g87) & (!sk[1]) & (!g90) & (!g231) & (g273) & (g317)) + ((g87) & (!sk[1]) & (!g90) & (g231) & (!g273) & (!g317)) + ((g87) & (!sk[1]) & (!g90) & (g231) & (!g273) & (g317)) + ((g87) & (!sk[1]) & (!g90) & (g231) & (g273) & (!g317)) + ((g87) & (!sk[1]) & (!g90) & (g231) & (g273) & (g317)) + ((g87) & (!sk[1]) & (g90) & (!g231) & (!g273) & (!g317)) + ((g87) & (!sk[1]) & (g90) & (!g231) & (!g273) & (g317)) + ((g87) & (!sk[1]) & (g90) & (!g231) & (g273) & (!g317)) + ((g87) & (!sk[1]) & (g90) & (!g231) & (g273) & (g317)) + ((g87) & (!sk[1]) & (g90) & (g231) & (!g273) & (!g317)) + ((g87) & (!sk[1]) & (g90) & (g231) & (!g273) & (g317)) + ((g87) & (!sk[1]) & (g90) & (g231) & (g273) & (!g317)) + ((g87) & (!sk[1]) & (g90) & (g231) & (g273) & (g317)) + ((g87) & (sk[1]) & (!g90) & (!g231) & (g273) & (g317)) + ((g87) & (sk[1]) & (!g90) & (g231) & (!g273) & (g317)) + ((g87) & (sk[1]) & (!g90) & (g231) & (g273) & (g317)) + ((g87) & (sk[1]) & (g90) & (!g231) & (!g273) & (g317)) + ((g87) & (sk[1]) & (g90) & (!g231) & (g273) & (!g317)) + ((g87) & (sk[1]) & (g90) & (!g231) & (g273) & (g317)) + ((g87) & (sk[1]) & (g90) & (g231) & (!g273) & (!g317)) + ((g87) & (sk[1]) & (g90) & (g231) & (!g273) & (g317)) + ((g87) & (sk[1]) & (g90) & (g231) & (g273) & (!g317)) + ((g87) & (sk[1]) & (g90) & (g231) & (g273) & (g317)));
	assign g4114 = (((!g2140) & (!sk[2]) & (!g2282) & (g321)) + ((!g2140) & (!sk[2]) & (g2282) & (!g321)) + ((!g2140) & (!sk[2]) & (g2282) & (g321)) + ((!g2140) & (sk[2]) & (!g2282) & (g321)) + ((!g2140) & (sk[2]) & (g2282) & (g321)) + ((g2140) & (!sk[2]) & (!g2282) & (g321)) + ((g2140) & (!sk[2]) & (g2282) & (!g321)) + ((g2140) & (!sk[2]) & (g2282) & (g321)) + ((g2140) & (sk[2]) & (g2282) & (!g321)) + ((g2140) & (sk[2]) & (g2282) & (g321)));
	assign g4115 = (((!sk[3]) & (!g2142) & (!g2282) & (g322)) + ((!sk[3]) & (!g2142) & (g2282) & (!g322)) + ((!sk[3]) & (!g2142) & (g2282) & (g322)) + ((!sk[3]) & (g2142) & (!g2282) & (g322)) + ((!sk[3]) & (g2142) & (g2282) & (!g322)) + ((!sk[3]) & (g2142) & (g2282) & (g322)) + ((sk[3]) & (!g2142) & (!g2282) & (g322)) + ((sk[3]) & (!g2142) & (g2282) & (g322)) + ((sk[3]) & (g2142) & (g2282) & (!g322)) + ((sk[3]) & (g2142) & (g2282) & (g322)));
	assign g4116 = (((!sk[4]) & (!g2144) & (!g2282) & (g323)) + ((!sk[4]) & (!g2144) & (g2282) & (!g323)) + ((!sk[4]) & (!g2144) & (g2282) & (g323)) + ((!sk[4]) & (g2144) & (!g2282) & (g323)) + ((!sk[4]) & (g2144) & (g2282) & (!g323)) + ((!sk[4]) & (g2144) & (g2282) & (g323)) + ((sk[4]) & (!g2144) & (!g2282) & (g323)) + ((sk[4]) & (!g2144) & (g2282) & (g323)) + ((sk[4]) & (g2144) & (g2282) & (!g323)) + ((sk[4]) & (g2144) & (g2282) & (g323)));
	assign g4117 = (((!g2145) & (!g2282) & (!sk[5]) & (g324)) + ((!g2145) & (!g2282) & (sk[5]) & (g324)) + ((!g2145) & (g2282) & (!sk[5]) & (!g324)) + ((!g2145) & (g2282) & (!sk[5]) & (g324)) + ((!g2145) & (g2282) & (sk[5]) & (g324)) + ((g2145) & (!g2282) & (!sk[5]) & (g324)) + ((g2145) & (g2282) & (!sk[5]) & (!g324)) + ((g2145) & (g2282) & (!sk[5]) & (g324)) + ((g2145) & (g2282) & (sk[5]) & (!g324)) + ((g2145) & (g2282) & (sk[5]) & (g324)));
	assign g325 = (((!g321) & (!g322) & (!g323) & (g324) & (g147) & (g148)) + ((!g321) & (!g322) & (g323) & (!g324) & (!g147) & (g148)) + ((!g321) & (!g322) & (g323) & (g324) & (!g147) & (g148)) + ((!g321) & (!g322) & (g323) & (g324) & (g147) & (g148)) + ((!g321) & (g322) & (!g323) & (!g324) & (g147) & (!g148)) + ((!g321) & (g322) & (!g323) & (g324) & (g147) & (!g148)) + ((!g321) & (g322) & (!g323) & (g324) & (g147) & (g148)) + ((!g321) & (g322) & (g323) & (!g324) & (!g147) & (g148)) + ((!g321) & (g322) & (g323) & (!g324) & (g147) & (!g148)) + ((!g321) & (g322) & (g323) & (g324) & (!g147) & (g148)) + ((!g321) & (g322) & (g323) & (g324) & (g147) & (!g148)) + ((!g321) & (g322) & (g323) & (g324) & (g147) & (g148)) + ((g321) & (!g322) & (!g323) & (!g324) & (!g147) & (!g148)) + ((g321) & (!g322) & (!g323) & (g324) & (!g147) & (!g148)) + ((g321) & (!g322) & (!g323) & (g324) & (g147) & (g148)) + ((g321) & (!g322) & (g323) & (!g324) & (!g147) & (!g148)) + ((g321) & (!g322) & (g323) & (!g324) & (!g147) & (g148)) + ((g321) & (!g322) & (g323) & (g324) & (!g147) & (!g148)) + ((g321) & (!g322) & (g323) & (g324) & (!g147) & (g148)) + ((g321) & (!g322) & (g323) & (g324) & (g147) & (g148)) + ((g321) & (g322) & (!g323) & (!g324) & (!g147) & (!g148)) + ((g321) & (g322) & (!g323) & (!g324) & (g147) & (!g148)) + ((g321) & (g322) & (!g323) & (g324) & (!g147) & (!g148)) + ((g321) & (g322) & (!g323) & (g324) & (g147) & (!g148)) + ((g321) & (g322) & (!g323) & (g324) & (g147) & (g148)) + ((g321) & (g322) & (g323) & (!g324) & (!g147) & (!g148)) + ((g321) & (g322) & (g323) & (!g324) & (!g147) & (g148)) + ((g321) & (g322) & (g323) & (!g324) & (g147) & (!g148)) + ((g321) & (g322) & (g323) & (g324) & (!g147) & (!g148)) + ((g321) & (g322) & (g323) & (g324) & (!g147) & (g148)) + ((g321) & (g322) & (g323) & (g324) & (g147) & (!g148)) + ((g321) & (g322) & (g323) & (g324) & (g147) & (g148)));
	assign g4118 = (((!g2146) & (!sk[7]) & (!g2282) & (g326)) + ((!g2146) & (!sk[7]) & (g2282) & (!g326)) + ((!g2146) & (!sk[7]) & (g2282) & (g326)) + ((!g2146) & (sk[7]) & (!g2282) & (g326)) + ((!g2146) & (sk[7]) & (g2282) & (g326)) + ((g2146) & (!sk[7]) & (!g2282) & (g326)) + ((g2146) & (!sk[7]) & (g2282) & (!g326)) + ((g2146) & (!sk[7]) & (g2282) & (g326)) + ((g2146) & (sk[7]) & (g2282) & (!g326)) + ((g2146) & (sk[7]) & (g2282) & (g326)));
	assign g4119 = (((!sk[8]) & (!g2148) & (!g2282) & (g327)) + ((!sk[8]) & (!g2148) & (g2282) & (!g327)) + ((!sk[8]) & (!g2148) & (g2282) & (g327)) + ((!sk[8]) & (g2148) & (!g2282) & (g327)) + ((!sk[8]) & (g2148) & (g2282) & (!g327)) + ((!sk[8]) & (g2148) & (g2282) & (g327)) + ((sk[8]) & (!g2148) & (!g2282) & (g327)) + ((sk[8]) & (!g2148) & (g2282) & (g327)) + ((sk[8]) & (g2148) & (g2282) & (!g327)) + ((sk[8]) & (g2148) & (g2282) & (g327)));
	assign g4120 = (((!sk[9]) & (!g2150) & (!g2282) & (g328)) + ((!sk[9]) & (!g2150) & (g2282) & (!g328)) + ((!sk[9]) & (!g2150) & (g2282) & (g328)) + ((!sk[9]) & (g2150) & (!g2282) & (g328)) + ((!sk[9]) & (g2150) & (g2282) & (!g328)) + ((!sk[9]) & (g2150) & (g2282) & (g328)) + ((sk[9]) & (!g2150) & (!g2282) & (g328)) + ((sk[9]) & (!g2150) & (g2282) & (g328)) + ((sk[9]) & (g2150) & (g2282) & (!g328)) + ((sk[9]) & (g2150) & (g2282) & (g328)));
	assign g4121 = (((!g2151) & (!g2282) & (!sk[10]) & (g329)) + ((!g2151) & (!g2282) & (sk[10]) & (g329)) + ((!g2151) & (g2282) & (!sk[10]) & (!g329)) + ((!g2151) & (g2282) & (!sk[10]) & (g329)) + ((!g2151) & (g2282) & (sk[10]) & (g329)) + ((g2151) & (!g2282) & (!sk[10]) & (g329)) + ((g2151) & (g2282) & (!sk[10]) & (!g329)) + ((g2151) & (g2282) & (!sk[10]) & (g329)) + ((g2151) & (g2282) & (sk[10]) & (!g329)) + ((g2151) & (g2282) & (sk[10]) & (g329)));
	assign g330 = (((!g326) & (!g327) & (!g328) & (g329) & (g147) & (g148)) + ((!g326) & (!g327) & (g328) & (!g329) & (!g147) & (g148)) + ((!g326) & (!g327) & (g328) & (g329) & (!g147) & (g148)) + ((!g326) & (!g327) & (g328) & (g329) & (g147) & (g148)) + ((!g326) & (g327) & (!g328) & (!g329) & (g147) & (!g148)) + ((!g326) & (g327) & (!g328) & (g329) & (g147) & (!g148)) + ((!g326) & (g327) & (!g328) & (g329) & (g147) & (g148)) + ((!g326) & (g327) & (g328) & (!g329) & (!g147) & (g148)) + ((!g326) & (g327) & (g328) & (!g329) & (g147) & (!g148)) + ((!g326) & (g327) & (g328) & (g329) & (!g147) & (g148)) + ((!g326) & (g327) & (g328) & (g329) & (g147) & (!g148)) + ((!g326) & (g327) & (g328) & (g329) & (g147) & (g148)) + ((g326) & (!g327) & (!g328) & (!g329) & (!g147) & (!g148)) + ((g326) & (!g327) & (!g328) & (g329) & (!g147) & (!g148)) + ((g326) & (!g327) & (!g328) & (g329) & (g147) & (g148)) + ((g326) & (!g327) & (g328) & (!g329) & (!g147) & (!g148)) + ((g326) & (!g327) & (g328) & (!g329) & (!g147) & (g148)) + ((g326) & (!g327) & (g328) & (g329) & (!g147) & (!g148)) + ((g326) & (!g327) & (g328) & (g329) & (!g147) & (g148)) + ((g326) & (!g327) & (g328) & (g329) & (g147) & (g148)) + ((g326) & (g327) & (!g328) & (!g329) & (!g147) & (!g148)) + ((g326) & (g327) & (!g328) & (!g329) & (g147) & (!g148)) + ((g326) & (g327) & (!g328) & (g329) & (!g147) & (!g148)) + ((g326) & (g327) & (!g328) & (g329) & (g147) & (!g148)) + ((g326) & (g327) & (!g328) & (g329) & (g147) & (g148)) + ((g326) & (g327) & (g328) & (!g329) & (!g147) & (!g148)) + ((g326) & (g327) & (g328) & (!g329) & (!g147) & (g148)) + ((g326) & (g327) & (g328) & (!g329) & (g147) & (!g148)) + ((g326) & (g327) & (g328) & (g329) & (!g147) & (!g148)) + ((g326) & (g327) & (g328) & (g329) & (!g147) & (g148)) + ((g326) & (g327) & (g328) & (g329) & (g147) & (!g148)) + ((g326) & (g327) & (g328) & (g329) & (g147) & (g148)));
	assign g4122 = (((!g2152) & (!sk[12]) & (!g2282) & (g331)) + ((!g2152) & (!sk[12]) & (g2282) & (!g331)) + ((!g2152) & (!sk[12]) & (g2282) & (g331)) + ((!g2152) & (sk[12]) & (!g2282) & (g331)) + ((!g2152) & (sk[12]) & (g2282) & (g331)) + ((g2152) & (!sk[12]) & (!g2282) & (g331)) + ((g2152) & (!sk[12]) & (g2282) & (!g331)) + ((g2152) & (!sk[12]) & (g2282) & (g331)) + ((g2152) & (sk[12]) & (g2282) & (!g331)) + ((g2152) & (sk[12]) & (g2282) & (g331)));
	assign g4123 = (((!sk[13]) & (!g2153) & (!g2282) & (g332)) + ((!sk[13]) & (!g2153) & (g2282) & (!g332)) + ((!sk[13]) & (!g2153) & (g2282) & (g332)) + ((!sk[13]) & (g2153) & (!g2282) & (g332)) + ((!sk[13]) & (g2153) & (g2282) & (!g332)) + ((!sk[13]) & (g2153) & (g2282) & (g332)) + ((sk[13]) & (!g2153) & (!g2282) & (g332)) + ((sk[13]) & (!g2153) & (g2282) & (g332)) + ((sk[13]) & (g2153) & (g2282) & (!g332)) + ((sk[13]) & (g2153) & (g2282) & (g332)));
	assign g4124 = (((!sk[14]) & (!g2155) & (!g2282) & (g333)) + ((!sk[14]) & (!g2155) & (g2282) & (!g333)) + ((!sk[14]) & (!g2155) & (g2282) & (g333)) + ((!sk[14]) & (g2155) & (!g2282) & (g333)) + ((!sk[14]) & (g2155) & (g2282) & (!g333)) + ((!sk[14]) & (g2155) & (g2282) & (g333)) + ((sk[14]) & (!g2155) & (!g2282) & (g333)) + ((sk[14]) & (!g2155) & (g2282) & (g333)) + ((sk[14]) & (g2155) & (g2282) & (!g333)) + ((sk[14]) & (g2155) & (g2282) & (g333)));
	assign g4125 = (((!g2157) & (!g2282) & (!sk[15]) & (g334)) + ((!g2157) & (!g2282) & (sk[15]) & (g334)) + ((!g2157) & (g2282) & (!sk[15]) & (!g334)) + ((!g2157) & (g2282) & (!sk[15]) & (g334)) + ((!g2157) & (g2282) & (sk[15]) & (g334)) + ((g2157) & (!g2282) & (!sk[15]) & (g334)) + ((g2157) & (g2282) & (!sk[15]) & (!g334)) + ((g2157) & (g2282) & (!sk[15]) & (g334)) + ((g2157) & (g2282) & (sk[15]) & (!g334)) + ((g2157) & (g2282) & (sk[15]) & (g334)));
	assign g335 = (((!g331) & (!g332) & (!g333) & (g334) & (g147) & (g148)) + ((!g331) & (!g332) & (g333) & (!g334) & (!g147) & (g148)) + ((!g331) & (!g332) & (g333) & (g334) & (!g147) & (g148)) + ((!g331) & (!g332) & (g333) & (g334) & (g147) & (g148)) + ((!g331) & (g332) & (!g333) & (!g334) & (g147) & (!g148)) + ((!g331) & (g332) & (!g333) & (g334) & (g147) & (!g148)) + ((!g331) & (g332) & (!g333) & (g334) & (g147) & (g148)) + ((!g331) & (g332) & (g333) & (!g334) & (!g147) & (g148)) + ((!g331) & (g332) & (g333) & (!g334) & (g147) & (!g148)) + ((!g331) & (g332) & (g333) & (g334) & (!g147) & (g148)) + ((!g331) & (g332) & (g333) & (g334) & (g147) & (!g148)) + ((!g331) & (g332) & (g333) & (g334) & (g147) & (g148)) + ((g331) & (!g332) & (!g333) & (!g334) & (!g147) & (!g148)) + ((g331) & (!g332) & (!g333) & (g334) & (!g147) & (!g148)) + ((g331) & (!g332) & (!g333) & (g334) & (g147) & (g148)) + ((g331) & (!g332) & (g333) & (!g334) & (!g147) & (!g148)) + ((g331) & (!g332) & (g333) & (!g334) & (!g147) & (g148)) + ((g331) & (!g332) & (g333) & (g334) & (!g147) & (!g148)) + ((g331) & (!g332) & (g333) & (g334) & (!g147) & (g148)) + ((g331) & (!g332) & (g333) & (g334) & (g147) & (g148)) + ((g331) & (g332) & (!g333) & (!g334) & (!g147) & (!g148)) + ((g331) & (g332) & (!g333) & (!g334) & (g147) & (!g148)) + ((g331) & (g332) & (!g333) & (g334) & (!g147) & (!g148)) + ((g331) & (g332) & (!g333) & (g334) & (g147) & (!g148)) + ((g331) & (g332) & (!g333) & (g334) & (g147) & (g148)) + ((g331) & (g332) & (g333) & (!g334) & (!g147) & (!g148)) + ((g331) & (g332) & (g333) & (!g334) & (!g147) & (g148)) + ((g331) & (g332) & (g333) & (!g334) & (g147) & (!g148)) + ((g331) & (g332) & (g333) & (g334) & (!g147) & (!g148)) + ((g331) & (g332) & (g333) & (g334) & (!g147) & (g148)) + ((g331) & (g332) & (g333) & (g334) & (g147) & (!g148)) + ((g331) & (g332) & (g333) & (g334) & (g147) & (g148)));
	assign g4126 = (((!g2158) & (!g2282) & (!sk[17]) & (g336)) + ((!g2158) & (!g2282) & (sk[17]) & (g336)) + ((!g2158) & (g2282) & (!sk[17]) & (!g336)) + ((!g2158) & (g2282) & (!sk[17]) & (g336)) + ((!g2158) & (g2282) & (sk[17]) & (g336)) + ((g2158) & (!g2282) & (!sk[17]) & (g336)) + ((g2158) & (g2282) & (!sk[17]) & (!g336)) + ((g2158) & (g2282) & (!sk[17]) & (g336)) + ((g2158) & (g2282) & (sk[17]) & (!g336)) + ((g2158) & (g2282) & (sk[17]) & (g336)));
	assign g4127 = (((!sk[18]) & (!g2159) & (!g2282) & (g337)) + ((!sk[18]) & (!g2159) & (g2282) & (!g337)) + ((!sk[18]) & (!g2159) & (g2282) & (g337)) + ((!sk[18]) & (g2159) & (!g2282) & (g337)) + ((!sk[18]) & (g2159) & (g2282) & (!g337)) + ((!sk[18]) & (g2159) & (g2282) & (g337)) + ((sk[18]) & (!g2159) & (!g2282) & (g337)) + ((sk[18]) & (!g2159) & (g2282) & (g337)) + ((sk[18]) & (g2159) & (g2282) & (!g337)) + ((sk[18]) & (g2159) & (g2282) & (g337)));
	assign g4128 = (((!g2160) & (!sk[19]) & (!g2282) & (g338)) + ((!g2160) & (!sk[19]) & (g2282) & (!g338)) + ((!g2160) & (!sk[19]) & (g2282) & (g338)) + ((!g2160) & (sk[19]) & (!g2282) & (g338)) + ((!g2160) & (sk[19]) & (g2282) & (g338)) + ((g2160) & (!sk[19]) & (!g2282) & (g338)) + ((g2160) & (!sk[19]) & (g2282) & (!g338)) + ((g2160) & (!sk[19]) & (g2282) & (g338)) + ((g2160) & (sk[19]) & (g2282) & (!g338)) + ((g2160) & (sk[19]) & (g2282) & (g338)));
	assign g4129 = (((!g2161) & (!sk[20]) & (!g2282) & (g339)) + ((!g2161) & (!sk[20]) & (g2282) & (!g339)) + ((!g2161) & (!sk[20]) & (g2282) & (g339)) + ((!g2161) & (sk[20]) & (!g2282) & (g339)) + ((!g2161) & (sk[20]) & (g2282) & (g339)) + ((g2161) & (!sk[20]) & (!g2282) & (g339)) + ((g2161) & (!sk[20]) & (g2282) & (!g339)) + ((g2161) & (!sk[20]) & (g2282) & (g339)) + ((g2161) & (sk[20]) & (g2282) & (!g339)) + ((g2161) & (sk[20]) & (g2282) & (g339)));
	assign g340 = (((!g336) & (!g337) & (!g338) & (g339) & (g147) & (g148)) + ((!g336) & (!g337) & (g338) & (!g339) & (!g147) & (g148)) + ((!g336) & (!g337) & (g338) & (g339) & (!g147) & (g148)) + ((!g336) & (!g337) & (g338) & (g339) & (g147) & (g148)) + ((!g336) & (g337) & (!g338) & (!g339) & (g147) & (!g148)) + ((!g336) & (g337) & (!g338) & (g339) & (g147) & (!g148)) + ((!g336) & (g337) & (!g338) & (g339) & (g147) & (g148)) + ((!g336) & (g337) & (g338) & (!g339) & (!g147) & (g148)) + ((!g336) & (g337) & (g338) & (!g339) & (g147) & (!g148)) + ((!g336) & (g337) & (g338) & (g339) & (!g147) & (g148)) + ((!g336) & (g337) & (g338) & (g339) & (g147) & (!g148)) + ((!g336) & (g337) & (g338) & (g339) & (g147) & (g148)) + ((g336) & (!g337) & (!g338) & (!g339) & (!g147) & (!g148)) + ((g336) & (!g337) & (!g338) & (g339) & (!g147) & (!g148)) + ((g336) & (!g337) & (!g338) & (g339) & (g147) & (g148)) + ((g336) & (!g337) & (g338) & (!g339) & (!g147) & (!g148)) + ((g336) & (!g337) & (g338) & (!g339) & (!g147) & (g148)) + ((g336) & (!g337) & (g338) & (g339) & (!g147) & (!g148)) + ((g336) & (!g337) & (g338) & (g339) & (!g147) & (g148)) + ((g336) & (!g337) & (g338) & (g339) & (g147) & (g148)) + ((g336) & (g337) & (!g338) & (!g339) & (!g147) & (!g148)) + ((g336) & (g337) & (!g338) & (!g339) & (g147) & (!g148)) + ((g336) & (g337) & (!g338) & (g339) & (!g147) & (!g148)) + ((g336) & (g337) & (!g338) & (g339) & (g147) & (!g148)) + ((g336) & (g337) & (!g338) & (g339) & (g147) & (g148)) + ((g336) & (g337) & (g338) & (!g339) & (!g147) & (!g148)) + ((g336) & (g337) & (g338) & (!g339) & (!g147) & (g148)) + ((g336) & (g337) & (g338) & (!g339) & (g147) & (!g148)) + ((g336) & (g337) & (g338) & (g339) & (!g147) & (!g148)) + ((g336) & (g337) & (g338) & (g339) & (!g147) & (g148)) + ((g336) & (g337) & (g338) & (g339) & (g147) & (!g148)) + ((g336) & (g337) & (g338) & (g339) & (g147) & (g148)));
	assign g341 = (((!g325) & (!g330) & (!g335) & (g340) & (g165) & (g166)) + ((!g325) & (!g330) & (g335) & (!g340) & (!g165) & (g166)) + ((!g325) & (!g330) & (g335) & (g340) & (!g165) & (g166)) + ((!g325) & (!g330) & (g335) & (g340) & (g165) & (g166)) + ((!g325) & (g330) & (!g335) & (!g340) & (g165) & (!g166)) + ((!g325) & (g330) & (!g335) & (g340) & (g165) & (!g166)) + ((!g325) & (g330) & (!g335) & (g340) & (g165) & (g166)) + ((!g325) & (g330) & (g335) & (!g340) & (!g165) & (g166)) + ((!g325) & (g330) & (g335) & (!g340) & (g165) & (!g166)) + ((!g325) & (g330) & (g335) & (g340) & (!g165) & (g166)) + ((!g325) & (g330) & (g335) & (g340) & (g165) & (!g166)) + ((!g325) & (g330) & (g335) & (g340) & (g165) & (g166)) + ((g325) & (!g330) & (!g335) & (!g340) & (!g165) & (!g166)) + ((g325) & (!g330) & (!g335) & (g340) & (!g165) & (!g166)) + ((g325) & (!g330) & (!g335) & (g340) & (g165) & (g166)) + ((g325) & (!g330) & (g335) & (!g340) & (!g165) & (!g166)) + ((g325) & (!g330) & (g335) & (!g340) & (!g165) & (g166)) + ((g325) & (!g330) & (g335) & (g340) & (!g165) & (!g166)) + ((g325) & (!g330) & (g335) & (g340) & (!g165) & (g166)) + ((g325) & (!g330) & (g335) & (g340) & (g165) & (g166)) + ((g325) & (g330) & (!g335) & (!g340) & (!g165) & (!g166)) + ((g325) & (g330) & (!g335) & (!g340) & (g165) & (!g166)) + ((g325) & (g330) & (!g335) & (g340) & (!g165) & (!g166)) + ((g325) & (g330) & (!g335) & (g340) & (g165) & (!g166)) + ((g325) & (g330) & (!g335) & (g340) & (g165) & (g166)) + ((g325) & (g330) & (g335) & (!g340) & (!g165) & (!g166)) + ((g325) & (g330) & (g335) & (!g340) & (!g165) & (g166)) + ((g325) & (g330) & (g335) & (!g340) & (g165) & (!g166)) + ((g325) & (g330) & (g335) & (g340) & (!g165) & (!g166)) + ((g325) & (g330) & (g335) & (g340) & (!g165) & (g166)) + ((g325) & (g330) & (g335) & (g340) & (g165) & (!g166)) + ((g325) & (g330) & (g335) & (g340) & (g165) & (g166)));
	assign g4130 = (((!sk[23]) & (!g2173) & (!g2282) & (g342)) + ((!sk[23]) & (!g2173) & (g2282) & (!g342)) + ((!sk[23]) & (!g2173) & (g2282) & (g342)) + ((!sk[23]) & (g2173) & (!g2282) & (g342)) + ((!sk[23]) & (g2173) & (g2282) & (!g342)) + ((!sk[23]) & (g2173) & (g2282) & (g342)) + ((sk[23]) & (!g2173) & (!g2282) & (g342)) + ((sk[23]) & (!g2173) & (g2282) & (g342)) + ((sk[23]) & (g2173) & (g2282) & (!g342)) + ((sk[23]) & (g2173) & (g2282) & (g342)));
	assign g4131 = (((!sk[24]) & (!g2174) & (!g2282) & (g343)) + ((!sk[24]) & (!g2174) & (g2282) & (!g343)) + ((!sk[24]) & (!g2174) & (g2282) & (g343)) + ((!sk[24]) & (g2174) & (!g2282) & (g343)) + ((!sk[24]) & (g2174) & (g2282) & (!g343)) + ((!sk[24]) & (g2174) & (g2282) & (g343)) + ((sk[24]) & (!g2174) & (!g2282) & (g343)) + ((sk[24]) & (!g2174) & (g2282) & (g343)) + ((sk[24]) & (g2174) & (g2282) & (!g343)) + ((sk[24]) & (g2174) & (g2282) & (g343)));
	assign g4132 = (((!g2175) & (!g2282) & (!sk[25]) & (g344)) + ((!g2175) & (!g2282) & (sk[25]) & (g344)) + ((!g2175) & (g2282) & (!sk[25]) & (!g344)) + ((!g2175) & (g2282) & (!sk[25]) & (g344)) + ((!g2175) & (g2282) & (sk[25]) & (g344)) + ((g2175) & (!g2282) & (!sk[25]) & (g344)) + ((g2175) & (g2282) & (!sk[25]) & (!g344)) + ((g2175) & (g2282) & (!sk[25]) & (g344)) + ((g2175) & (g2282) & (sk[25]) & (!g344)) + ((g2175) & (g2282) & (sk[25]) & (g344)));
	assign g4133 = (((!sk[26]) & (!g2176) & (!g2282) & (g345)) + ((!sk[26]) & (!g2176) & (g2282) & (!g345)) + ((!sk[26]) & (!g2176) & (g2282) & (g345)) + ((!sk[26]) & (g2176) & (!g2282) & (g345)) + ((!sk[26]) & (g2176) & (g2282) & (!g345)) + ((!sk[26]) & (g2176) & (g2282) & (g345)) + ((sk[26]) & (!g2176) & (!g2282) & (g345)) + ((sk[26]) & (!g2176) & (g2282) & (g345)) + ((sk[26]) & (g2176) & (g2282) & (!g345)) + ((sk[26]) & (g2176) & (g2282) & (g345)));
	assign g346 = (((!g342) & (!g343) & (!g344) & (g345) & (g165) & (g166)) + ((!g342) & (!g343) & (g344) & (!g345) & (!g165) & (g166)) + ((!g342) & (!g343) & (g344) & (g345) & (!g165) & (g166)) + ((!g342) & (!g343) & (g344) & (g345) & (g165) & (g166)) + ((!g342) & (g343) & (!g344) & (!g345) & (g165) & (!g166)) + ((!g342) & (g343) & (!g344) & (g345) & (g165) & (!g166)) + ((!g342) & (g343) & (!g344) & (g345) & (g165) & (g166)) + ((!g342) & (g343) & (g344) & (!g345) & (!g165) & (g166)) + ((!g342) & (g343) & (g344) & (!g345) & (g165) & (!g166)) + ((!g342) & (g343) & (g344) & (g345) & (!g165) & (g166)) + ((!g342) & (g343) & (g344) & (g345) & (g165) & (!g166)) + ((!g342) & (g343) & (g344) & (g345) & (g165) & (g166)) + ((g342) & (!g343) & (!g344) & (!g345) & (!g165) & (!g166)) + ((g342) & (!g343) & (!g344) & (g345) & (!g165) & (!g166)) + ((g342) & (!g343) & (!g344) & (g345) & (g165) & (g166)) + ((g342) & (!g343) & (g344) & (!g345) & (!g165) & (!g166)) + ((g342) & (!g343) & (g344) & (!g345) & (!g165) & (g166)) + ((g342) & (!g343) & (g344) & (g345) & (!g165) & (!g166)) + ((g342) & (!g343) & (g344) & (g345) & (!g165) & (g166)) + ((g342) & (!g343) & (g344) & (g345) & (g165) & (g166)) + ((g342) & (g343) & (!g344) & (!g345) & (!g165) & (!g166)) + ((g342) & (g343) & (!g344) & (!g345) & (g165) & (!g166)) + ((g342) & (g343) & (!g344) & (g345) & (!g165) & (!g166)) + ((g342) & (g343) & (!g344) & (g345) & (g165) & (!g166)) + ((g342) & (g343) & (!g344) & (g345) & (g165) & (g166)) + ((g342) & (g343) & (g344) & (!g345) & (!g165) & (!g166)) + ((g342) & (g343) & (g344) & (!g345) & (!g165) & (g166)) + ((g342) & (g343) & (g344) & (!g345) & (g165) & (!g166)) + ((g342) & (g343) & (g344) & (g345) & (!g165) & (!g166)) + ((g342) & (g343) & (g344) & (g345) & (!g165) & (g166)) + ((g342) & (g343) & (g344) & (g345) & (g165) & (!g166)) + ((g342) & (g343) & (g344) & (g345) & (g165) & (g166)));
	assign g4134 = (((!sk[28]) & (!g2177) & (!g2282) & (g347)) + ((!sk[28]) & (!g2177) & (g2282) & (!g347)) + ((!sk[28]) & (!g2177) & (g2282) & (g347)) + ((!sk[28]) & (g2177) & (!g2282) & (g347)) + ((!sk[28]) & (g2177) & (g2282) & (!g347)) + ((!sk[28]) & (g2177) & (g2282) & (g347)) + ((sk[28]) & (!g2177) & (!g2282) & (g347)) + ((sk[28]) & (!g2177) & (g2282) & (g347)) + ((sk[28]) & (g2177) & (g2282) & (!g347)) + ((sk[28]) & (g2177) & (g2282) & (g347)));
	assign g4135 = (((!sk[29]) & (!g2178) & (!g2282) & (g348)) + ((!sk[29]) & (!g2178) & (g2282) & (!g348)) + ((!sk[29]) & (!g2178) & (g2282) & (g348)) + ((!sk[29]) & (g2178) & (!g2282) & (g348)) + ((!sk[29]) & (g2178) & (g2282) & (!g348)) + ((!sk[29]) & (g2178) & (g2282) & (g348)) + ((sk[29]) & (!g2178) & (!g2282) & (g348)) + ((sk[29]) & (!g2178) & (g2282) & (g348)) + ((sk[29]) & (g2178) & (g2282) & (!g348)) + ((sk[29]) & (g2178) & (g2282) & (g348)));
	assign g4136 = (((!g2179) & (!g2282) & (!sk[30]) & (g349)) + ((!g2179) & (!g2282) & (sk[30]) & (g349)) + ((!g2179) & (g2282) & (!sk[30]) & (!g349)) + ((!g2179) & (g2282) & (!sk[30]) & (g349)) + ((!g2179) & (g2282) & (sk[30]) & (g349)) + ((g2179) & (!g2282) & (!sk[30]) & (g349)) + ((g2179) & (g2282) & (!sk[30]) & (!g349)) + ((g2179) & (g2282) & (!sk[30]) & (g349)) + ((g2179) & (g2282) & (sk[30]) & (!g349)) + ((g2179) & (g2282) & (sk[30]) & (g349)));
	assign g350 = (((!g165) & (!sk[31]) & (!g166) & (!g347) & (g348) & (!g349)) + ((!g165) & (!sk[31]) & (!g166) & (!g347) & (g348) & (g349)) + ((!g165) & (!sk[31]) & (!g166) & (g347) & (!g348) & (!g349)) + ((!g165) & (!sk[31]) & (!g166) & (g347) & (!g348) & (g349)) + ((!g165) & (!sk[31]) & (!g166) & (g347) & (g348) & (!g349)) + ((!g165) & (!sk[31]) & (!g166) & (g347) & (g348) & (g349)) + ((!g165) & (!sk[31]) & (g166) & (!g347) & (!g348) & (!g349)) + ((!g165) & (!sk[31]) & (g166) & (!g347) & (!g348) & (g349)) + ((!g165) & (!sk[31]) & (g166) & (!g347) & (g348) & (!g349)) + ((!g165) & (!sk[31]) & (g166) & (!g347) & (g348) & (g349)) + ((!g165) & (!sk[31]) & (g166) & (g347) & (!g348) & (!g349)) + ((!g165) & (!sk[31]) & (g166) & (g347) & (!g348) & (g349)) + ((!g165) & (!sk[31]) & (g166) & (g347) & (g348) & (!g349)) + ((!g165) & (!sk[31]) & (g166) & (g347) & (g348) & (g349)) + ((!g165) & (sk[31]) & (g166) & (!g347) & (!g348) & (g349)) + ((!g165) & (sk[31]) & (g166) & (!g347) & (g348) & (g349)) + ((!g165) & (sk[31]) & (g166) & (g347) & (!g348) & (g349)) + ((!g165) & (sk[31]) & (g166) & (g347) & (g348) & (g349)) + ((g165) & (!sk[31]) & (!g166) & (!g347) & (g348) & (!g349)) + ((g165) & (!sk[31]) & (!g166) & (!g347) & (g348) & (g349)) + ((g165) & (!sk[31]) & (!g166) & (g347) & (!g348) & (!g349)) + ((g165) & (!sk[31]) & (!g166) & (g347) & (!g348) & (g349)) + ((g165) & (!sk[31]) & (!g166) & (g347) & (g348) & (!g349)) + ((g165) & (!sk[31]) & (!g166) & (g347) & (g348) & (g349)) + ((g165) & (!sk[31]) & (g166) & (!g347) & (!g348) & (!g349)) + ((g165) & (!sk[31]) & (g166) & (!g347) & (!g348) & (g349)) + ((g165) & (!sk[31]) & (g166) & (!g347) & (g348) & (!g349)) + ((g165) & (!sk[31]) & (g166) & (!g347) & (g348) & (g349)) + ((g165) & (!sk[31]) & (g166) & (g347) & (!g348) & (!g349)) + ((g165) & (!sk[31]) & (g166) & (g347) & (!g348) & (g349)) + ((g165) & (!sk[31]) & (g166) & (g347) & (g348) & (!g349)) + ((g165) & (!sk[31]) & (g166) & (g347) & (g348) & (g349)) + ((g165) & (sk[31]) & (!g166) & (g347) & (!g348) & (!g349)) + ((g165) & (sk[31]) & (!g166) & (g347) & (!g348) & (g349)) + ((g165) & (sk[31]) & (!g166) & (g347) & (g348) & (!g349)) + ((g165) & (sk[31]) & (!g166) & (g347) & (g348) & (g349)) + ((g165) & (sk[31]) & (g166) & (!g347) & (g348) & (!g349)) + ((g165) & (sk[31]) & (g166) & (!g347) & (g348) & (g349)) + ((g165) & (sk[31]) & (g166) & (g347) & (g348) & (!g349)) + ((g165) & (sk[31]) & (g166) & (g347) & (g348) & (g349)));
	assign g4137 = (((!sk[32]) & (!g2162) & (!g2282) & (g351)) + ((!sk[32]) & (!g2162) & (g2282) & (!g351)) + ((!sk[32]) & (!g2162) & (g2282) & (g351)) + ((!sk[32]) & (g2162) & (!g2282) & (g351)) + ((!sk[32]) & (g2162) & (g2282) & (!g351)) + ((!sk[32]) & (g2162) & (g2282) & (g351)) + ((sk[32]) & (!g2162) & (!g2282) & (g351)) + ((sk[32]) & (!g2162) & (g2282) & (g351)) + ((sk[32]) & (g2162) & (g2282) & (!g351)) + ((sk[32]) & (g2162) & (g2282) & (g351)));
	assign g4138 = (((!g2164) & (!g2282) & (!sk[33]) & (g352)) + ((!g2164) & (!g2282) & (sk[33]) & (g352)) + ((!g2164) & (g2282) & (!sk[33]) & (!g352)) + ((!g2164) & (g2282) & (!sk[33]) & (g352)) + ((!g2164) & (g2282) & (sk[33]) & (g352)) + ((g2164) & (!g2282) & (!sk[33]) & (g352)) + ((g2164) & (g2282) & (!sk[33]) & (!g352)) + ((g2164) & (g2282) & (!sk[33]) & (g352)) + ((g2164) & (g2282) & (sk[33]) & (!g352)) + ((g2164) & (g2282) & (sk[33]) & (g352)));
	assign g4139 = (((!g2166) & (!sk[34]) & (!g2282) & (g353)) + ((!g2166) & (!sk[34]) & (g2282) & (!g353)) + ((!g2166) & (!sk[34]) & (g2282) & (g353)) + ((!g2166) & (sk[34]) & (!g2282) & (g353)) + ((!g2166) & (sk[34]) & (g2282) & (g353)) + ((g2166) & (!sk[34]) & (!g2282) & (g353)) + ((g2166) & (!sk[34]) & (g2282) & (!g353)) + ((g2166) & (!sk[34]) & (g2282) & (g353)) + ((g2166) & (sk[34]) & (g2282) & (!g353)) + ((g2166) & (sk[34]) & (g2282) & (g353)));
	assign g4140 = (((!g2168) & (!sk[35]) & (!g2282) & (g354)) + ((!g2168) & (!sk[35]) & (g2282) & (!g354)) + ((!g2168) & (!sk[35]) & (g2282) & (g354)) + ((!g2168) & (sk[35]) & (!g2282) & (g354)) + ((!g2168) & (sk[35]) & (g2282) & (g354)) + ((g2168) & (!sk[35]) & (!g2282) & (g354)) + ((g2168) & (!sk[35]) & (g2282) & (!g354)) + ((g2168) & (!sk[35]) & (g2282) & (g354)) + ((g2168) & (sk[35]) & (g2282) & (!g354)) + ((g2168) & (sk[35]) & (g2282) & (g354)));
	assign g355 = (((!g351) & (!g352) & (!g353) & (g354) & (g165) & (g166)) + ((!g351) & (!g352) & (g353) & (!g354) & (!g165) & (g166)) + ((!g351) & (!g352) & (g353) & (g354) & (!g165) & (g166)) + ((!g351) & (!g352) & (g353) & (g354) & (g165) & (g166)) + ((!g351) & (g352) & (!g353) & (!g354) & (g165) & (!g166)) + ((!g351) & (g352) & (!g353) & (g354) & (g165) & (!g166)) + ((!g351) & (g352) & (!g353) & (g354) & (g165) & (g166)) + ((!g351) & (g352) & (g353) & (!g354) & (!g165) & (g166)) + ((!g351) & (g352) & (g353) & (!g354) & (g165) & (!g166)) + ((!g351) & (g352) & (g353) & (g354) & (!g165) & (g166)) + ((!g351) & (g352) & (g353) & (g354) & (g165) & (!g166)) + ((!g351) & (g352) & (g353) & (g354) & (g165) & (g166)) + ((g351) & (!g352) & (!g353) & (!g354) & (!g165) & (!g166)) + ((g351) & (!g352) & (!g353) & (g354) & (!g165) & (!g166)) + ((g351) & (!g352) & (!g353) & (g354) & (g165) & (g166)) + ((g351) & (!g352) & (g353) & (!g354) & (!g165) & (!g166)) + ((g351) & (!g352) & (g353) & (!g354) & (!g165) & (g166)) + ((g351) & (!g352) & (g353) & (g354) & (!g165) & (!g166)) + ((g351) & (!g352) & (g353) & (g354) & (!g165) & (g166)) + ((g351) & (!g352) & (g353) & (g354) & (g165) & (g166)) + ((g351) & (g352) & (!g353) & (!g354) & (!g165) & (!g166)) + ((g351) & (g352) & (!g353) & (!g354) & (g165) & (!g166)) + ((g351) & (g352) & (!g353) & (g354) & (!g165) & (!g166)) + ((g351) & (g352) & (!g353) & (g354) & (g165) & (!g166)) + ((g351) & (g352) & (!g353) & (g354) & (g165) & (g166)) + ((g351) & (g352) & (g353) & (!g354) & (!g165) & (!g166)) + ((g351) & (g352) & (g353) & (!g354) & (!g165) & (g166)) + ((g351) & (g352) & (g353) & (!g354) & (g165) & (!g166)) + ((g351) & (g352) & (g353) & (g354) & (!g165) & (!g166)) + ((g351) & (g352) & (g353) & (g354) & (!g165) & (g166)) + ((g351) & (g352) & (g353) & (g354) & (g165) & (!g166)) + ((g351) & (g352) & (g353) & (g354) & (g165) & (g166)));
	assign g4141 = (((!g2169) & (!sk[37]) & (!g2282) & (g356)) + ((!g2169) & (!sk[37]) & (g2282) & (!g356)) + ((!g2169) & (!sk[37]) & (g2282) & (g356)) + ((!g2169) & (sk[37]) & (!g2282) & (g356)) + ((!g2169) & (sk[37]) & (g2282) & (g356)) + ((g2169) & (!sk[37]) & (!g2282) & (g356)) + ((g2169) & (!sk[37]) & (g2282) & (!g356)) + ((g2169) & (!sk[37]) & (g2282) & (g356)) + ((g2169) & (sk[37]) & (g2282) & (!g356)) + ((g2169) & (sk[37]) & (g2282) & (g356)));
	assign g4142 = (((!sk[38]) & (!g2170) & (!g2282) & (g357)) + ((!sk[38]) & (!g2170) & (g2282) & (!g357)) + ((!sk[38]) & (!g2170) & (g2282) & (g357)) + ((!sk[38]) & (g2170) & (!g2282) & (g357)) + ((!sk[38]) & (g2170) & (g2282) & (!g357)) + ((!sk[38]) & (g2170) & (g2282) & (g357)) + ((sk[38]) & (!g2170) & (!g2282) & (g357)) + ((sk[38]) & (!g2170) & (g2282) & (g357)) + ((sk[38]) & (g2170) & (g2282) & (!g357)) + ((sk[38]) & (g2170) & (g2282) & (g357)));
	assign g4143 = (((!sk[39]) & (!g2171) & (!g2282) & (g358)) + ((!sk[39]) & (!g2171) & (g2282) & (!g358)) + ((!sk[39]) & (!g2171) & (g2282) & (g358)) + ((!sk[39]) & (g2171) & (!g2282) & (g358)) + ((!sk[39]) & (g2171) & (g2282) & (!g358)) + ((!sk[39]) & (g2171) & (g2282) & (g358)) + ((sk[39]) & (!g2171) & (!g2282) & (g358)) + ((sk[39]) & (!g2171) & (g2282) & (g358)) + ((sk[39]) & (g2171) & (g2282) & (!g358)) + ((sk[39]) & (g2171) & (g2282) & (g358)));
	assign g4144 = (((!g2172) & (!sk[40]) & (!g2282) & (g359)) + ((!g2172) & (!sk[40]) & (g2282) & (!g359)) + ((!g2172) & (!sk[40]) & (g2282) & (g359)) + ((!g2172) & (sk[40]) & (!g2282) & (g359)) + ((!g2172) & (sk[40]) & (g2282) & (g359)) + ((g2172) & (!sk[40]) & (!g2282) & (g359)) + ((g2172) & (!sk[40]) & (g2282) & (!g359)) + ((g2172) & (!sk[40]) & (g2282) & (g359)) + ((g2172) & (sk[40]) & (g2282) & (!g359)) + ((g2172) & (sk[40]) & (g2282) & (g359)));
	assign g360 = (((!g356) & (!g357) & (!g358) & (g359) & (g165) & (g166)) + ((!g356) & (!g357) & (g358) & (!g359) & (!g165) & (g166)) + ((!g356) & (!g357) & (g358) & (g359) & (!g165) & (g166)) + ((!g356) & (!g357) & (g358) & (g359) & (g165) & (g166)) + ((!g356) & (g357) & (!g358) & (!g359) & (g165) & (!g166)) + ((!g356) & (g357) & (!g358) & (g359) & (g165) & (!g166)) + ((!g356) & (g357) & (!g358) & (g359) & (g165) & (g166)) + ((!g356) & (g357) & (g358) & (!g359) & (!g165) & (g166)) + ((!g356) & (g357) & (g358) & (!g359) & (g165) & (!g166)) + ((!g356) & (g357) & (g358) & (g359) & (!g165) & (g166)) + ((!g356) & (g357) & (g358) & (g359) & (g165) & (!g166)) + ((!g356) & (g357) & (g358) & (g359) & (g165) & (g166)) + ((g356) & (!g357) & (!g358) & (!g359) & (!g165) & (!g166)) + ((g356) & (!g357) & (!g358) & (g359) & (!g165) & (!g166)) + ((g356) & (!g357) & (!g358) & (g359) & (g165) & (g166)) + ((g356) & (!g357) & (g358) & (!g359) & (!g165) & (!g166)) + ((g356) & (!g357) & (g358) & (!g359) & (!g165) & (g166)) + ((g356) & (!g357) & (g358) & (g359) & (!g165) & (!g166)) + ((g356) & (!g357) & (g358) & (g359) & (!g165) & (g166)) + ((g356) & (!g357) & (g358) & (g359) & (g165) & (g166)) + ((g356) & (g357) & (!g358) & (!g359) & (!g165) & (!g166)) + ((g356) & (g357) & (!g358) & (!g359) & (g165) & (!g166)) + ((g356) & (g357) & (!g358) & (g359) & (!g165) & (!g166)) + ((g356) & (g357) & (!g358) & (g359) & (g165) & (!g166)) + ((g356) & (g357) & (!g358) & (g359) & (g165) & (g166)) + ((g356) & (g357) & (g358) & (!g359) & (!g165) & (!g166)) + ((g356) & (g357) & (g358) & (!g359) & (!g165) & (g166)) + ((g356) & (g357) & (g358) & (!g359) & (g165) & (!g166)) + ((g356) & (g357) & (g358) & (g359) & (!g165) & (!g166)) + ((g356) & (g357) & (g358) & (g359) & (!g165) & (g166)) + ((g356) & (g357) & (g358) & (g359) & (g165) & (!g166)) + ((g356) & (g357) & (g358) & (g359) & (g165) & (g166)));
	assign g361 = (((!g147) & (!g148) & (!g346) & (g350) & (!g355) & (!g360)) + ((!g147) & (!g148) & (!g346) & (g350) & (!g355) & (g360)) + ((!g147) & (!g148) & (!g346) & (g350) & (g355) & (!g360)) + ((!g147) & (!g148) & (!g346) & (g350) & (g355) & (g360)) + ((!g147) & (!g148) & (g346) & (g350) & (!g355) & (!g360)) + ((!g147) & (!g148) & (g346) & (g350) & (!g355) & (g360)) + ((!g147) & (!g148) & (g346) & (g350) & (g355) & (!g360)) + ((!g147) & (!g148) & (g346) & (g350) & (g355) & (g360)) + ((!g147) & (g148) & (!g346) & (!g350) & (!g355) & (g360)) + ((!g147) & (g148) & (!g346) & (!g350) & (g355) & (g360)) + ((!g147) & (g148) & (!g346) & (g350) & (!g355) & (g360)) + ((!g147) & (g148) & (!g346) & (g350) & (g355) & (g360)) + ((!g147) & (g148) & (g346) & (!g350) & (!g355) & (g360)) + ((!g147) & (g148) & (g346) & (!g350) & (g355) & (g360)) + ((!g147) & (g148) & (g346) & (g350) & (!g355) & (g360)) + ((!g147) & (g148) & (g346) & (g350) & (g355) & (g360)) + ((g147) & (!g148) & (g346) & (!g350) & (!g355) & (!g360)) + ((g147) & (!g148) & (g346) & (!g350) & (!g355) & (g360)) + ((g147) & (!g148) & (g346) & (!g350) & (g355) & (!g360)) + ((g147) & (!g148) & (g346) & (!g350) & (g355) & (g360)) + ((g147) & (!g148) & (g346) & (g350) & (!g355) & (!g360)) + ((g147) & (!g148) & (g346) & (g350) & (!g355) & (g360)) + ((g147) & (!g148) & (g346) & (g350) & (g355) & (!g360)) + ((g147) & (!g148) & (g346) & (g350) & (g355) & (g360)) + ((g147) & (g148) & (!g346) & (!g350) & (g355) & (!g360)) + ((g147) & (g148) & (!g346) & (!g350) & (g355) & (g360)) + ((g147) & (g148) & (!g346) & (g350) & (g355) & (!g360)) + ((g147) & (g148) & (!g346) & (g350) & (g355) & (g360)) + ((g147) & (g148) & (g346) & (!g350) & (g355) & (!g360)) + ((g147) & (g148) & (g346) & (!g350) & (g355) & (g360)) + ((g147) & (g148) & (g346) & (g350) & (g355) & (!g360)) + ((g147) & (g148) & (g346) & (g350) & (g355) & (g360)));
	assign g362 = (((!g142) & (!g341) & (!sk[43]) & (g361)) + ((!g142) & (!g341) & (sk[43]) & (g361)) + ((!g142) & (g341) & (!sk[43]) & (!g361)) + ((!g142) & (g341) & (!sk[43]) & (g361)) + ((!g142) & (g341) & (sk[43]) & (g361)) + ((g142) & (!g341) & (!sk[43]) & (g361)) + ((g142) & (g341) & (!sk[43]) & (!g361)) + ((g142) & (g341) & (!sk[43]) & (g361)) + ((g142) & (g341) & (sk[43]) & (!g361)) + ((g142) & (g341) & (sk[43]) & (g361)));
	assign g363 = (((!g126) & (!g318) & (!g319) & (!sk[44]) & (g320) & (!g362)) + ((!g126) & (!g318) & (!g319) & (!sk[44]) & (g320) & (g362)) + ((!g126) & (!g318) & (g319) & (!sk[44]) & (!g320) & (!g362)) + ((!g126) & (!g318) & (g319) & (!sk[44]) & (!g320) & (g362)) + ((!g126) & (!g318) & (g319) & (!sk[44]) & (g320) & (!g362)) + ((!g126) & (!g318) & (g319) & (!sk[44]) & (g320) & (g362)) + ((!g126) & (!g318) & (g319) & (sk[44]) & (!g320) & (!g362)) + ((!g126) & (!g318) & (g319) & (sk[44]) & (!g320) & (g362)) + ((!g126) & (!g318) & (g319) & (sk[44]) & (g320) & (!g362)) + ((!g126) & (!g318) & (g319) & (sk[44]) & (g320) & (g362)) + ((!g126) & (g318) & (!g319) & (!sk[44]) & (!g320) & (!g362)) + ((!g126) & (g318) & (!g319) & (!sk[44]) & (!g320) & (g362)) + ((!g126) & (g318) & (!g319) & (!sk[44]) & (g320) & (!g362)) + ((!g126) & (g318) & (!g319) & (!sk[44]) & (g320) & (g362)) + ((!g126) & (g318) & (g319) & (!sk[44]) & (!g320) & (!g362)) + ((!g126) & (g318) & (g319) & (!sk[44]) & (!g320) & (g362)) + ((!g126) & (g318) & (g319) & (!sk[44]) & (g320) & (!g362)) + ((!g126) & (g318) & (g319) & (!sk[44]) & (g320) & (g362)) + ((!g126) & (g318) & (g319) & (sk[44]) & (!g320) & (!g362)) + ((!g126) & (g318) & (g319) & (sk[44]) & (!g320) & (g362)) + ((!g126) & (g318) & (g319) & (sk[44]) & (g320) & (!g362)) + ((!g126) & (g318) & (g319) & (sk[44]) & (g320) & (g362)) + ((g126) & (!g318) & (!g319) & (!sk[44]) & (g320) & (!g362)) + ((g126) & (!g318) & (!g319) & (!sk[44]) & (g320) & (g362)) + ((g126) & (!g318) & (!g319) & (sk[44]) & (!g320) & (g362)) + ((g126) & (!g318) & (!g319) & (sk[44]) & (g320) & (!g362)) + ((g126) & (!g318) & (g319) & (!sk[44]) & (!g320) & (!g362)) + ((g126) & (!g318) & (g319) & (!sk[44]) & (!g320) & (g362)) + ((g126) & (!g318) & (g319) & (!sk[44]) & (g320) & (!g362)) + ((g126) & (!g318) & (g319) & (!sk[44]) & (g320) & (g362)) + ((g126) & (!g318) & (g319) & (sk[44]) & (!g320) & (g362)) + ((g126) & (!g318) & (g319) & (sk[44]) & (g320) & (!g362)) + ((g126) & (g318) & (!g319) & (!sk[44]) & (!g320) & (!g362)) + ((g126) & (g318) & (!g319) & (!sk[44]) & (!g320) & (g362)) + ((g126) & (g318) & (!g319) & (!sk[44]) & (g320) & (!g362)) + ((g126) & (g318) & (!g319) & (!sk[44]) & (g320) & (g362)) + ((g126) & (g318) & (!g319) & (sk[44]) & (!g320) & (!g362)) + ((g126) & (g318) & (!g319) & (sk[44]) & (g320) & (g362)) + ((g126) & (g318) & (g319) & (!sk[44]) & (!g320) & (!g362)) + ((g126) & (g318) & (g319) & (!sk[44]) & (!g320) & (g362)) + ((g126) & (g318) & (g319) & (!sk[44]) & (g320) & (!g362)) + ((g126) & (g318) & (g319) & (!sk[44]) & (g320) & (g362)) + ((g126) & (g318) & (g319) & (sk[44]) & (!g320) & (!g362)) + ((g126) & (g318) & (g319) & (sk[44]) & (g320) & (g362)));
	assign g4145 = (((!g2064) & (!dmem_dat_ix5x) & (!sk[45]) & (g364)) + ((!g2064) & (!dmem_dat_ix5x) & (sk[45]) & (g364)) + ((!g2064) & (dmem_dat_ix5x) & (!sk[45]) & (!g364)) + ((!g2064) & (dmem_dat_ix5x) & (!sk[45]) & (g364)) + ((!g2064) & (dmem_dat_ix5x) & (sk[45]) & (g364)) + ((g2064) & (!dmem_dat_ix5x) & (!sk[45]) & (g364)) + ((g2064) & (dmem_dat_ix5x) & (!sk[45]) & (!g364)) + ((g2064) & (dmem_dat_ix5x) & (!sk[45]) & (g364)) + ((g2064) & (dmem_dat_ix5x) & (sk[45]) & (!g364)) + ((g2064) & (dmem_dat_ix5x) & (sk[45]) & (g364)));
	assign g4146 = (((!sk[46]) & (!g2059) & (!g2288) & (g365)) + ((!sk[46]) & (!g2059) & (g2288) & (!g365)) + ((!sk[46]) & (!g2059) & (g2288) & (g365)) + ((!sk[46]) & (g2059) & (!g2288) & (g365)) + ((!sk[46]) & (g2059) & (g2288) & (!g365)) + ((!sk[46]) & (g2059) & (g2288) & (g365)) + ((sk[46]) & (!g2059) & (!g2288) & (g365)) + ((sk[46]) & (!g2059) & (g2288) & (g365)) + ((sk[46]) & (g2059) & (g2288) & (!g365)) + ((sk[46]) & (g2059) & (g2288) & (g365)));
	assign g4147 = (((!g2140) & (!sk[47]) & (!g2304) & (g366)) + ((!g2140) & (!sk[47]) & (g2304) & (!g366)) + ((!g2140) & (!sk[47]) & (g2304) & (g366)) + ((!g2140) & (sk[47]) & (!g2304) & (g366)) + ((!g2140) & (sk[47]) & (g2304) & (g366)) + ((g2140) & (!sk[47]) & (!g2304) & (g366)) + ((g2140) & (!sk[47]) & (g2304) & (!g366)) + ((g2140) & (!sk[47]) & (g2304) & (g366)) + ((g2140) & (sk[47]) & (g2304) & (!g366)) + ((g2140) & (sk[47]) & (g2304) & (g366)));
	assign g4148 = (((!g2146) & (!g2304) & (!sk[48]) & (g367)) + ((!g2146) & (!g2304) & (sk[48]) & (g367)) + ((!g2146) & (g2304) & (!sk[48]) & (!g367)) + ((!g2146) & (g2304) & (!sk[48]) & (g367)) + ((!g2146) & (g2304) & (sk[48]) & (g367)) + ((g2146) & (!g2304) & (!sk[48]) & (g367)) + ((g2146) & (g2304) & (!sk[48]) & (!g367)) + ((g2146) & (g2304) & (!sk[48]) & (g367)) + ((g2146) & (g2304) & (sk[48]) & (!g367)) + ((g2146) & (g2304) & (sk[48]) & (g367)));
	assign g4149 = (((!sk[49]) & (!g2152) & (!g2304) & (g368)) + ((!sk[49]) & (!g2152) & (g2304) & (!g368)) + ((!sk[49]) & (!g2152) & (g2304) & (g368)) + ((!sk[49]) & (g2152) & (!g2304) & (g368)) + ((!sk[49]) & (g2152) & (g2304) & (!g368)) + ((!sk[49]) & (g2152) & (g2304) & (g368)) + ((sk[49]) & (!g2152) & (!g2304) & (g368)) + ((sk[49]) & (!g2152) & (g2304) & (g368)) + ((sk[49]) & (g2152) & (g2304) & (!g368)) + ((sk[49]) & (g2152) & (g2304) & (g368)));
	assign g4150 = (((!sk[50]) & (!g2158) & (!g2304) & (g369)) + ((!sk[50]) & (!g2158) & (g2304) & (!g369)) + ((!sk[50]) & (!g2158) & (g2304) & (g369)) + ((!sk[50]) & (g2158) & (!g2304) & (g369)) + ((!sk[50]) & (g2158) & (g2304) & (!g369)) + ((!sk[50]) & (g2158) & (g2304) & (g369)) + ((sk[50]) & (!g2158) & (!g2304) & (g369)) + ((sk[50]) & (!g2158) & (g2304) & (g369)) + ((sk[50]) & (g2158) & (g2304) & (!g369)) + ((sk[50]) & (g2158) & (g2304) & (g369)));
	assign g370 = (((!g366) & (!g367) & (!g368) & (g369) & (g165) & (g166)) + ((!g366) & (!g367) & (g368) & (!g369) & (!g165) & (g166)) + ((!g366) & (!g367) & (g368) & (g369) & (!g165) & (g166)) + ((!g366) & (!g367) & (g368) & (g369) & (g165) & (g166)) + ((!g366) & (g367) & (!g368) & (!g369) & (g165) & (!g166)) + ((!g366) & (g367) & (!g368) & (g369) & (g165) & (!g166)) + ((!g366) & (g367) & (!g368) & (g369) & (g165) & (g166)) + ((!g366) & (g367) & (g368) & (!g369) & (!g165) & (g166)) + ((!g366) & (g367) & (g368) & (!g369) & (g165) & (!g166)) + ((!g366) & (g367) & (g368) & (g369) & (!g165) & (g166)) + ((!g366) & (g367) & (g368) & (g369) & (g165) & (!g166)) + ((!g366) & (g367) & (g368) & (g369) & (g165) & (g166)) + ((g366) & (!g367) & (!g368) & (!g369) & (!g165) & (!g166)) + ((g366) & (!g367) & (!g368) & (g369) & (!g165) & (!g166)) + ((g366) & (!g367) & (!g368) & (g369) & (g165) & (g166)) + ((g366) & (!g367) & (g368) & (!g369) & (!g165) & (!g166)) + ((g366) & (!g367) & (g368) & (!g369) & (!g165) & (g166)) + ((g366) & (!g367) & (g368) & (g369) & (!g165) & (!g166)) + ((g366) & (!g367) & (g368) & (g369) & (!g165) & (g166)) + ((g366) & (!g367) & (g368) & (g369) & (g165) & (g166)) + ((g366) & (g367) & (!g368) & (!g369) & (!g165) & (!g166)) + ((g366) & (g367) & (!g368) & (!g369) & (g165) & (!g166)) + ((g366) & (g367) & (!g368) & (g369) & (!g165) & (!g166)) + ((g366) & (g367) & (!g368) & (g369) & (g165) & (!g166)) + ((g366) & (g367) & (!g368) & (g369) & (g165) & (g166)) + ((g366) & (g367) & (g368) & (!g369) & (!g165) & (!g166)) + ((g366) & (g367) & (g368) & (!g369) & (!g165) & (g166)) + ((g366) & (g367) & (g368) & (!g369) & (g165) & (!g166)) + ((g366) & (g367) & (g368) & (g369) & (!g165) & (!g166)) + ((g366) & (g367) & (g368) & (g369) & (!g165) & (g166)) + ((g366) & (g367) & (g368) & (g369) & (g165) & (!g166)) + ((g366) & (g367) & (g368) & (g369) & (g165) & (g166)));
	assign g4151 = (((!g2142) & (!g2304) & (!sk[52]) & (g371)) + ((!g2142) & (!g2304) & (sk[52]) & (g371)) + ((!g2142) & (g2304) & (!sk[52]) & (!g371)) + ((!g2142) & (g2304) & (!sk[52]) & (g371)) + ((!g2142) & (g2304) & (sk[52]) & (g371)) + ((g2142) & (!g2304) & (!sk[52]) & (g371)) + ((g2142) & (g2304) & (!sk[52]) & (!g371)) + ((g2142) & (g2304) & (!sk[52]) & (g371)) + ((g2142) & (g2304) & (sk[52]) & (!g371)) + ((g2142) & (g2304) & (sk[52]) & (g371)));
	assign g4152 = (((!g2148) & (!sk[53]) & (!g2304) & (g372)) + ((!g2148) & (!sk[53]) & (g2304) & (!g372)) + ((!g2148) & (!sk[53]) & (g2304) & (g372)) + ((!g2148) & (sk[53]) & (!g2304) & (g372)) + ((!g2148) & (sk[53]) & (g2304) & (g372)) + ((g2148) & (!sk[53]) & (!g2304) & (g372)) + ((g2148) & (!sk[53]) & (g2304) & (!g372)) + ((g2148) & (!sk[53]) & (g2304) & (g372)) + ((g2148) & (sk[53]) & (g2304) & (!g372)) + ((g2148) & (sk[53]) & (g2304) & (g372)));
	assign g4153 = (((!sk[54]) & (!g2153) & (!g2304) & (g373)) + ((!sk[54]) & (!g2153) & (g2304) & (!g373)) + ((!sk[54]) & (!g2153) & (g2304) & (g373)) + ((!sk[54]) & (g2153) & (!g2304) & (g373)) + ((!sk[54]) & (g2153) & (g2304) & (!g373)) + ((!sk[54]) & (g2153) & (g2304) & (g373)) + ((sk[54]) & (!g2153) & (!g2304) & (g373)) + ((sk[54]) & (!g2153) & (g2304) & (g373)) + ((sk[54]) & (g2153) & (g2304) & (!g373)) + ((sk[54]) & (g2153) & (g2304) & (g373)));
	assign g4154 = (((!sk[55]) & (!g2159) & (!g2304) & (g374)) + ((!sk[55]) & (!g2159) & (g2304) & (!g374)) + ((!sk[55]) & (!g2159) & (g2304) & (g374)) + ((!sk[55]) & (g2159) & (!g2304) & (g374)) + ((!sk[55]) & (g2159) & (g2304) & (!g374)) + ((!sk[55]) & (g2159) & (g2304) & (g374)) + ((sk[55]) & (!g2159) & (!g2304) & (g374)) + ((sk[55]) & (!g2159) & (g2304) & (g374)) + ((sk[55]) & (g2159) & (g2304) & (!g374)) + ((sk[55]) & (g2159) & (g2304) & (g374)));
	assign g375 = (((!g371) & (!g372) & (!g373) & (g374) & (g165) & (g166)) + ((!g371) & (!g372) & (g373) & (!g374) & (!g165) & (g166)) + ((!g371) & (!g372) & (g373) & (g374) & (!g165) & (g166)) + ((!g371) & (!g372) & (g373) & (g374) & (g165) & (g166)) + ((!g371) & (g372) & (!g373) & (!g374) & (g165) & (!g166)) + ((!g371) & (g372) & (!g373) & (g374) & (g165) & (!g166)) + ((!g371) & (g372) & (!g373) & (g374) & (g165) & (g166)) + ((!g371) & (g372) & (g373) & (!g374) & (!g165) & (g166)) + ((!g371) & (g372) & (g373) & (!g374) & (g165) & (!g166)) + ((!g371) & (g372) & (g373) & (g374) & (!g165) & (g166)) + ((!g371) & (g372) & (g373) & (g374) & (g165) & (!g166)) + ((!g371) & (g372) & (g373) & (g374) & (g165) & (g166)) + ((g371) & (!g372) & (!g373) & (!g374) & (!g165) & (!g166)) + ((g371) & (!g372) & (!g373) & (g374) & (!g165) & (!g166)) + ((g371) & (!g372) & (!g373) & (g374) & (g165) & (g166)) + ((g371) & (!g372) & (g373) & (!g374) & (!g165) & (!g166)) + ((g371) & (!g372) & (g373) & (!g374) & (!g165) & (g166)) + ((g371) & (!g372) & (g373) & (g374) & (!g165) & (!g166)) + ((g371) & (!g372) & (g373) & (g374) & (!g165) & (g166)) + ((g371) & (!g372) & (g373) & (g374) & (g165) & (g166)) + ((g371) & (g372) & (!g373) & (!g374) & (!g165) & (!g166)) + ((g371) & (g372) & (!g373) & (!g374) & (g165) & (!g166)) + ((g371) & (g372) & (!g373) & (g374) & (!g165) & (!g166)) + ((g371) & (g372) & (!g373) & (g374) & (g165) & (!g166)) + ((g371) & (g372) & (!g373) & (g374) & (g165) & (g166)) + ((g371) & (g372) & (g373) & (!g374) & (!g165) & (!g166)) + ((g371) & (g372) & (g373) & (!g374) & (!g165) & (g166)) + ((g371) & (g372) & (g373) & (!g374) & (g165) & (!g166)) + ((g371) & (g372) & (g373) & (g374) & (!g165) & (!g166)) + ((g371) & (g372) & (g373) & (g374) & (!g165) & (g166)) + ((g371) & (g372) & (g373) & (g374) & (g165) & (!g166)) + ((g371) & (g372) & (g373) & (g374) & (g165) & (g166)));
	assign g4155 = (((!g2144) & (!g2304) & (!sk[57]) & (g376)) + ((!g2144) & (!g2304) & (sk[57]) & (g376)) + ((!g2144) & (g2304) & (!sk[57]) & (!g376)) + ((!g2144) & (g2304) & (!sk[57]) & (g376)) + ((!g2144) & (g2304) & (sk[57]) & (g376)) + ((g2144) & (!g2304) & (!sk[57]) & (g376)) + ((g2144) & (g2304) & (!sk[57]) & (!g376)) + ((g2144) & (g2304) & (!sk[57]) & (g376)) + ((g2144) & (g2304) & (sk[57]) & (!g376)) + ((g2144) & (g2304) & (sk[57]) & (g376)));
	assign g4156 = (((!g2150) & (!g2304) & (!sk[58]) & (g377)) + ((!g2150) & (!g2304) & (sk[58]) & (g377)) + ((!g2150) & (g2304) & (!sk[58]) & (!g377)) + ((!g2150) & (g2304) & (!sk[58]) & (g377)) + ((!g2150) & (g2304) & (sk[58]) & (g377)) + ((g2150) & (!g2304) & (!sk[58]) & (g377)) + ((g2150) & (g2304) & (!sk[58]) & (!g377)) + ((g2150) & (g2304) & (!sk[58]) & (g377)) + ((g2150) & (g2304) & (sk[58]) & (!g377)) + ((g2150) & (g2304) & (sk[58]) & (g377)));
	assign g4157 = (((!g2155) & (!g2304) & (!sk[59]) & (g378)) + ((!g2155) & (!g2304) & (sk[59]) & (g378)) + ((!g2155) & (g2304) & (!sk[59]) & (!g378)) + ((!g2155) & (g2304) & (!sk[59]) & (g378)) + ((!g2155) & (g2304) & (sk[59]) & (g378)) + ((g2155) & (!g2304) & (!sk[59]) & (g378)) + ((g2155) & (g2304) & (!sk[59]) & (!g378)) + ((g2155) & (g2304) & (!sk[59]) & (g378)) + ((g2155) & (g2304) & (sk[59]) & (!g378)) + ((g2155) & (g2304) & (sk[59]) & (g378)));
	assign g4158 = (((!g2160) & (!sk[60]) & (!g2304) & (g379)) + ((!g2160) & (!sk[60]) & (g2304) & (!g379)) + ((!g2160) & (!sk[60]) & (g2304) & (g379)) + ((!g2160) & (sk[60]) & (!g2304) & (g379)) + ((!g2160) & (sk[60]) & (g2304) & (g379)) + ((g2160) & (!sk[60]) & (!g2304) & (g379)) + ((g2160) & (!sk[60]) & (g2304) & (!g379)) + ((g2160) & (!sk[60]) & (g2304) & (g379)) + ((g2160) & (sk[60]) & (g2304) & (!g379)) + ((g2160) & (sk[60]) & (g2304) & (g379)));
	assign g380 = (((!g376) & (!g377) & (!g378) & (g379) & (g165) & (g166)) + ((!g376) & (!g377) & (g378) & (!g379) & (!g165) & (g166)) + ((!g376) & (!g377) & (g378) & (g379) & (!g165) & (g166)) + ((!g376) & (!g377) & (g378) & (g379) & (g165) & (g166)) + ((!g376) & (g377) & (!g378) & (!g379) & (g165) & (!g166)) + ((!g376) & (g377) & (!g378) & (g379) & (g165) & (!g166)) + ((!g376) & (g377) & (!g378) & (g379) & (g165) & (g166)) + ((!g376) & (g377) & (g378) & (!g379) & (!g165) & (g166)) + ((!g376) & (g377) & (g378) & (!g379) & (g165) & (!g166)) + ((!g376) & (g377) & (g378) & (g379) & (!g165) & (g166)) + ((!g376) & (g377) & (g378) & (g379) & (g165) & (!g166)) + ((!g376) & (g377) & (g378) & (g379) & (g165) & (g166)) + ((g376) & (!g377) & (!g378) & (!g379) & (!g165) & (!g166)) + ((g376) & (!g377) & (!g378) & (g379) & (!g165) & (!g166)) + ((g376) & (!g377) & (!g378) & (g379) & (g165) & (g166)) + ((g376) & (!g377) & (g378) & (!g379) & (!g165) & (!g166)) + ((g376) & (!g377) & (g378) & (!g379) & (!g165) & (g166)) + ((g376) & (!g377) & (g378) & (g379) & (!g165) & (!g166)) + ((g376) & (!g377) & (g378) & (g379) & (!g165) & (g166)) + ((g376) & (!g377) & (g378) & (g379) & (g165) & (g166)) + ((g376) & (g377) & (!g378) & (!g379) & (!g165) & (!g166)) + ((g376) & (g377) & (!g378) & (!g379) & (g165) & (!g166)) + ((g376) & (g377) & (!g378) & (g379) & (!g165) & (!g166)) + ((g376) & (g377) & (!g378) & (g379) & (g165) & (!g166)) + ((g376) & (g377) & (!g378) & (g379) & (g165) & (g166)) + ((g376) & (g377) & (g378) & (!g379) & (!g165) & (!g166)) + ((g376) & (g377) & (g378) & (!g379) & (!g165) & (g166)) + ((g376) & (g377) & (g378) & (!g379) & (g165) & (!g166)) + ((g376) & (g377) & (g378) & (g379) & (!g165) & (!g166)) + ((g376) & (g377) & (g378) & (g379) & (!g165) & (g166)) + ((g376) & (g377) & (g378) & (g379) & (g165) & (!g166)) + ((g376) & (g377) & (g378) & (g379) & (g165) & (g166)));
	assign g4159 = (((!g2145) & (!sk[62]) & (!g2304) & (g381)) + ((!g2145) & (!sk[62]) & (g2304) & (!g381)) + ((!g2145) & (!sk[62]) & (g2304) & (g381)) + ((!g2145) & (sk[62]) & (!g2304) & (g381)) + ((!g2145) & (sk[62]) & (g2304) & (g381)) + ((g2145) & (!sk[62]) & (!g2304) & (g381)) + ((g2145) & (!sk[62]) & (g2304) & (!g381)) + ((g2145) & (!sk[62]) & (g2304) & (g381)) + ((g2145) & (sk[62]) & (g2304) & (!g381)) + ((g2145) & (sk[62]) & (g2304) & (g381)));
	assign g4160 = (((!sk[63]) & (!g2151) & (!g2304) & (g382)) + ((!sk[63]) & (!g2151) & (g2304) & (!g382)) + ((!sk[63]) & (!g2151) & (g2304) & (g382)) + ((!sk[63]) & (g2151) & (!g2304) & (g382)) + ((!sk[63]) & (g2151) & (g2304) & (!g382)) + ((!sk[63]) & (g2151) & (g2304) & (g382)) + ((sk[63]) & (!g2151) & (!g2304) & (g382)) + ((sk[63]) & (!g2151) & (g2304) & (g382)) + ((sk[63]) & (g2151) & (g2304) & (!g382)) + ((sk[63]) & (g2151) & (g2304) & (g382)));
	assign g4161 = (((!g2157) & (!g2304) & (!sk[64]) & (g383)) + ((!g2157) & (!g2304) & (sk[64]) & (g383)) + ((!g2157) & (g2304) & (!sk[64]) & (!g383)) + ((!g2157) & (g2304) & (!sk[64]) & (g383)) + ((!g2157) & (g2304) & (sk[64]) & (g383)) + ((g2157) & (!g2304) & (!sk[64]) & (g383)) + ((g2157) & (g2304) & (!sk[64]) & (!g383)) + ((g2157) & (g2304) & (!sk[64]) & (g383)) + ((g2157) & (g2304) & (sk[64]) & (!g383)) + ((g2157) & (g2304) & (sk[64]) & (g383)));
	assign g4162 = (((!g2161) & (!g2304) & (!sk[65]) & (g384)) + ((!g2161) & (!g2304) & (sk[65]) & (g384)) + ((!g2161) & (g2304) & (!sk[65]) & (!g384)) + ((!g2161) & (g2304) & (!sk[65]) & (g384)) + ((!g2161) & (g2304) & (sk[65]) & (g384)) + ((g2161) & (!g2304) & (!sk[65]) & (g384)) + ((g2161) & (g2304) & (!sk[65]) & (!g384)) + ((g2161) & (g2304) & (!sk[65]) & (g384)) + ((g2161) & (g2304) & (sk[65]) & (!g384)) + ((g2161) & (g2304) & (sk[65]) & (g384)));
	assign g385 = (((!g381) & (!g382) & (!g383) & (g384) & (g165) & (g166)) + ((!g381) & (!g382) & (g383) & (!g384) & (!g165) & (g166)) + ((!g381) & (!g382) & (g383) & (g384) & (!g165) & (g166)) + ((!g381) & (!g382) & (g383) & (g384) & (g165) & (g166)) + ((!g381) & (g382) & (!g383) & (!g384) & (g165) & (!g166)) + ((!g381) & (g382) & (!g383) & (g384) & (g165) & (!g166)) + ((!g381) & (g382) & (!g383) & (g384) & (g165) & (g166)) + ((!g381) & (g382) & (g383) & (!g384) & (!g165) & (g166)) + ((!g381) & (g382) & (g383) & (!g384) & (g165) & (!g166)) + ((!g381) & (g382) & (g383) & (g384) & (!g165) & (g166)) + ((!g381) & (g382) & (g383) & (g384) & (g165) & (!g166)) + ((!g381) & (g382) & (g383) & (g384) & (g165) & (g166)) + ((g381) & (!g382) & (!g383) & (!g384) & (!g165) & (!g166)) + ((g381) & (!g382) & (!g383) & (g384) & (!g165) & (!g166)) + ((g381) & (!g382) & (!g383) & (g384) & (g165) & (g166)) + ((g381) & (!g382) & (g383) & (!g384) & (!g165) & (!g166)) + ((g381) & (!g382) & (g383) & (!g384) & (!g165) & (g166)) + ((g381) & (!g382) & (g383) & (g384) & (!g165) & (!g166)) + ((g381) & (!g382) & (g383) & (g384) & (!g165) & (g166)) + ((g381) & (!g382) & (g383) & (g384) & (g165) & (g166)) + ((g381) & (g382) & (!g383) & (!g384) & (!g165) & (!g166)) + ((g381) & (g382) & (!g383) & (!g384) & (g165) & (!g166)) + ((g381) & (g382) & (!g383) & (g384) & (!g165) & (!g166)) + ((g381) & (g382) & (!g383) & (g384) & (g165) & (!g166)) + ((g381) & (g382) & (!g383) & (g384) & (g165) & (g166)) + ((g381) & (g382) & (g383) & (!g384) & (!g165) & (!g166)) + ((g381) & (g382) & (g383) & (!g384) & (!g165) & (g166)) + ((g381) & (g382) & (g383) & (!g384) & (g165) & (!g166)) + ((g381) & (g382) & (g383) & (g384) & (!g165) & (!g166)) + ((g381) & (g382) & (g383) & (g384) & (!g165) & (g166)) + ((g381) & (g382) & (g383) & (g384) & (g165) & (!g166)) + ((g381) & (g382) & (g383) & (g384) & (g165) & (g166)));
	assign g386 = (((!g370) & (!g375) & (!g380) & (g385) & (g147) & (g148)) + ((!g370) & (!g375) & (g380) & (!g385) & (!g147) & (g148)) + ((!g370) & (!g375) & (g380) & (g385) & (!g147) & (g148)) + ((!g370) & (!g375) & (g380) & (g385) & (g147) & (g148)) + ((!g370) & (g375) & (!g380) & (!g385) & (g147) & (!g148)) + ((!g370) & (g375) & (!g380) & (g385) & (g147) & (!g148)) + ((!g370) & (g375) & (!g380) & (g385) & (g147) & (g148)) + ((!g370) & (g375) & (g380) & (!g385) & (!g147) & (g148)) + ((!g370) & (g375) & (g380) & (!g385) & (g147) & (!g148)) + ((!g370) & (g375) & (g380) & (g385) & (!g147) & (g148)) + ((!g370) & (g375) & (g380) & (g385) & (g147) & (!g148)) + ((!g370) & (g375) & (g380) & (g385) & (g147) & (g148)) + ((g370) & (!g375) & (!g380) & (!g385) & (!g147) & (!g148)) + ((g370) & (!g375) & (!g380) & (g385) & (!g147) & (!g148)) + ((g370) & (!g375) & (!g380) & (g385) & (g147) & (g148)) + ((g370) & (!g375) & (g380) & (!g385) & (!g147) & (!g148)) + ((g370) & (!g375) & (g380) & (!g385) & (!g147) & (g148)) + ((g370) & (!g375) & (g380) & (g385) & (!g147) & (!g148)) + ((g370) & (!g375) & (g380) & (g385) & (!g147) & (g148)) + ((g370) & (!g375) & (g380) & (g385) & (g147) & (g148)) + ((g370) & (g375) & (!g380) & (!g385) & (!g147) & (!g148)) + ((g370) & (g375) & (!g380) & (!g385) & (g147) & (!g148)) + ((g370) & (g375) & (!g380) & (g385) & (!g147) & (!g148)) + ((g370) & (g375) & (!g380) & (g385) & (g147) & (!g148)) + ((g370) & (g375) & (!g380) & (g385) & (g147) & (g148)) + ((g370) & (g375) & (g380) & (!g385) & (!g147) & (!g148)) + ((g370) & (g375) & (g380) & (!g385) & (!g147) & (g148)) + ((g370) & (g375) & (g380) & (!g385) & (g147) & (!g148)) + ((g370) & (g375) & (g380) & (g385) & (!g147) & (!g148)) + ((g370) & (g375) & (g380) & (g385) & (!g147) & (g148)) + ((g370) & (g375) & (g380) & (g385) & (g147) & (!g148)) + ((g370) & (g375) & (g380) & (g385) & (g147) & (g148)));
	assign g4163 = (((!sk[68]) & (!g2173) & (!g2304) & (g387)) + ((!sk[68]) & (!g2173) & (g2304) & (!g387)) + ((!sk[68]) & (!g2173) & (g2304) & (g387)) + ((!sk[68]) & (g2173) & (!g2304) & (g387)) + ((!sk[68]) & (g2173) & (g2304) & (!g387)) + ((!sk[68]) & (g2173) & (g2304) & (g387)) + ((sk[68]) & (!g2173) & (!g2304) & (g387)) + ((sk[68]) & (!g2173) & (g2304) & (g387)) + ((sk[68]) & (g2173) & (g2304) & (!g387)) + ((sk[68]) & (g2173) & (g2304) & (g387)));
	assign g4164 = (((!sk[69]) & (!g2174) & (!g2304) & (g388)) + ((!sk[69]) & (!g2174) & (g2304) & (!g388)) + ((!sk[69]) & (!g2174) & (g2304) & (g388)) + ((!sk[69]) & (g2174) & (!g2304) & (g388)) + ((!sk[69]) & (g2174) & (g2304) & (!g388)) + ((!sk[69]) & (g2174) & (g2304) & (g388)) + ((sk[69]) & (!g2174) & (!g2304) & (g388)) + ((sk[69]) & (!g2174) & (g2304) & (g388)) + ((sk[69]) & (g2174) & (g2304) & (!g388)) + ((sk[69]) & (g2174) & (g2304) & (g388)));
	assign g4165 = (((!g2175) & (!g2304) & (!sk[70]) & (g389)) + ((!g2175) & (!g2304) & (sk[70]) & (g389)) + ((!g2175) & (g2304) & (!sk[70]) & (!g389)) + ((!g2175) & (g2304) & (!sk[70]) & (g389)) + ((!g2175) & (g2304) & (sk[70]) & (g389)) + ((g2175) & (!g2304) & (!sk[70]) & (g389)) + ((g2175) & (g2304) & (!sk[70]) & (!g389)) + ((g2175) & (g2304) & (!sk[70]) & (g389)) + ((g2175) & (g2304) & (sk[70]) & (!g389)) + ((g2175) & (g2304) & (sk[70]) & (g389)));
	assign g4166 = (((!sk[71]) & (!g2176) & (!g2304) & (g390)) + ((!sk[71]) & (!g2176) & (g2304) & (!g390)) + ((!sk[71]) & (!g2176) & (g2304) & (g390)) + ((!sk[71]) & (g2176) & (!g2304) & (g390)) + ((!sk[71]) & (g2176) & (g2304) & (!g390)) + ((!sk[71]) & (g2176) & (g2304) & (g390)) + ((sk[71]) & (!g2176) & (!g2304) & (g390)) + ((sk[71]) & (!g2176) & (g2304) & (g390)) + ((sk[71]) & (g2176) & (g2304) & (!g390)) + ((sk[71]) & (g2176) & (g2304) & (g390)));
	assign g391 = (((!g387) & (!g388) & (!g389) & (g390) & (g165) & (g166)) + ((!g387) & (!g388) & (g389) & (!g390) & (!g165) & (g166)) + ((!g387) & (!g388) & (g389) & (g390) & (!g165) & (g166)) + ((!g387) & (!g388) & (g389) & (g390) & (g165) & (g166)) + ((!g387) & (g388) & (!g389) & (!g390) & (g165) & (!g166)) + ((!g387) & (g388) & (!g389) & (g390) & (g165) & (!g166)) + ((!g387) & (g388) & (!g389) & (g390) & (g165) & (g166)) + ((!g387) & (g388) & (g389) & (!g390) & (!g165) & (g166)) + ((!g387) & (g388) & (g389) & (!g390) & (g165) & (!g166)) + ((!g387) & (g388) & (g389) & (g390) & (!g165) & (g166)) + ((!g387) & (g388) & (g389) & (g390) & (g165) & (!g166)) + ((!g387) & (g388) & (g389) & (g390) & (g165) & (g166)) + ((g387) & (!g388) & (!g389) & (!g390) & (!g165) & (!g166)) + ((g387) & (!g388) & (!g389) & (g390) & (!g165) & (!g166)) + ((g387) & (!g388) & (!g389) & (g390) & (g165) & (g166)) + ((g387) & (!g388) & (g389) & (!g390) & (!g165) & (!g166)) + ((g387) & (!g388) & (g389) & (!g390) & (!g165) & (g166)) + ((g387) & (!g388) & (g389) & (g390) & (!g165) & (!g166)) + ((g387) & (!g388) & (g389) & (g390) & (!g165) & (g166)) + ((g387) & (!g388) & (g389) & (g390) & (g165) & (g166)) + ((g387) & (g388) & (!g389) & (!g390) & (!g165) & (!g166)) + ((g387) & (g388) & (!g389) & (!g390) & (g165) & (!g166)) + ((g387) & (g388) & (!g389) & (g390) & (!g165) & (!g166)) + ((g387) & (g388) & (!g389) & (g390) & (g165) & (!g166)) + ((g387) & (g388) & (!g389) & (g390) & (g165) & (g166)) + ((g387) & (g388) & (g389) & (!g390) & (!g165) & (!g166)) + ((g387) & (g388) & (g389) & (!g390) & (!g165) & (g166)) + ((g387) & (g388) & (g389) & (!g390) & (g165) & (!g166)) + ((g387) & (g388) & (g389) & (g390) & (!g165) & (!g166)) + ((g387) & (g388) & (g389) & (g390) & (!g165) & (g166)) + ((g387) & (g388) & (g389) & (g390) & (g165) & (!g166)) + ((g387) & (g388) & (g389) & (g390) & (g165) & (g166)));
	assign g4167 = (((!g2177) & (!sk[73]) & (!g2304) & (g392)) + ((!g2177) & (!sk[73]) & (g2304) & (!g392)) + ((!g2177) & (!sk[73]) & (g2304) & (g392)) + ((!g2177) & (sk[73]) & (!g2304) & (g392)) + ((!g2177) & (sk[73]) & (g2304) & (g392)) + ((g2177) & (!sk[73]) & (!g2304) & (g392)) + ((g2177) & (!sk[73]) & (g2304) & (!g392)) + ((g2177) & (!sk[73]) & (g2304) & (g392)) + ((g2177) & (sk[73]) & (g2304) & (!g392)) + ((g2177) & (sk[73]) & (g2304) & (g392)));
	assign g4168 = (((!g2178) & (!g2304) & (!sk[74]) & (g393)) + ((!g2178) & (!g2304) & (sk[74]) & (g393)) + ((!g2178) & (g2304) & (!sk[74]) & (!g393)) + ((!g2178) & (g2304) & (!sk[74]) & (g393)) + ((!g2178) & (g2304) & (sk[74]) & (g393)) + ((g2178) & (!g2304) & (!sk[74]) & (g393)) + ((g2178) & (g2304) & (!sk[74]) & (!g393)) + ((g2178) & (g2304) & (!sk[74]) & (g393)) + ((g2178) & (g2304) & (sk[74]) & (!g393)) + ((g2178) & (g2304) & (sk[74]) & (g393)));
	assign g4169 = (((!g2179) & (!g2304) & (!sk[75]) & (g394)) + ((!g2179) & (!g2304) & (sk[75]) & (g394)) + ((!g2179) & (g2304) & (!sk[75]) & (!g394)) + ((!g2179) & (g2304) & (!sk[75]) & (g394)) + ((!g2179) & (g2304) & (sk[75]) & (g394)) + ((g2179) & (!g2304) & (!sk[75]) & (g394)) + ((g2179) & (g2304) & (!sk[75]) & (!g394)) + ((g2179) & (g2304) & (!sk[75]) & (g394)) + ((g2179) & (g2304) & (sk[75]) & (!g394)) + ((g2179) & (g2304) & (sk[75]) & (g394)));
	assign g395 = (((!g165) & (!g166) & (!g392) & (!sk[76]) & (g393) & (!g394)) + ((!g165) & (!g166) & (!g392) & (!sk[76]) & (g393) & (g394)) + ((!g165) & (!g166) & (g392) & (!sk[76]) & (!g393) & (!g394)) + ((!g165) & (!g166) & (g392) & (!sk[76]) & (!g393) & (g394)) + ((!g165) & (!g166) & (g392) & (!sk[76]) & (g393) & (!g394)) + ((!g165) & (!g166) & (g392) & (!sk[76]) & (g393) & (g394)) + ((!g165) & (g166) & (!g392) & (!sk[76]) & (!g393) & (!g394)) + ((!g165) & (g166) & (!g392) & (!sk[76]) & (!g393) & (g394)) + ((!g165) & (g166) & (!g392) & (!sk[76]) & (g393) & (!g394)) + ((!g165) & (g166) & (!g392) & (!sk[76]) & (g393) & (g394)) + ((!g165) & (g166) & (!g392) & (sk[76]) & (!g393) & (g394)) + ((!g165) & (g166) & (!g392) & (sk[76]) & (g393) & (g394)) + ((!g165) & (g166) & (g392) & (!sk[76]) & (!g393) & (!g394)) + ((!g165) & (g166) & (g392) & (!sk[76]) & (!g393) & (g394)) + ((!g165) & (g166) & (g392) & (!sk[76]) & (g393) & (!g394)) + ((!g165) & (g166) & (g392) & (!sk[76]) & (g393) & (g394)) + ((!g165) & (g166) & (g392) & (sk[76]) & (!g393) & (g394)) + ((!g165) & (g166) & (g392) & (sk[76]) & (g393) & (g394)) + ((g165) & (!g166) & (!g392) & (!sk[76]) & (g393) & (!g394)) + ((g165) & (!g166) & (!g392) & (!sk[76]) & (g393) & (g394)) + ((g165) & (!g166) & (g392) & (!sk[76]) & (!g393) & (!g394)) + ((g165) & (!g166) & (g392) & (!sk[76]) & (!g393) & (g394)) + ((g165) & (!g166) & (g392) & (!sk[76]) & (g393) & (!g394)) + ((g165) & (!g166) & (g392) & (!sk[76]) & (g393) & (g394)) + ((g165) & (!g166) & (g392) & (sk[76]) & (!g393) & (!g394)) + ((g165) & (!g166) & (g392) & (sk[76]) & (!g393) & (g394)) + ((g165) & (!g166) & (g392) & (sk[76]) & (g393) & (!g394)) + ((g165) & (!g166) & (g392) & (sk[76]) & (g393) & (g394)) + ((g165) & (g166) & (!g392) & (!sk[76]) & (!g393) & (!g394)) + ((g165) & (g166) & (!g392) & (!sk[76]) & (!g393) & (g394)) + ((g165) & (g166) & (!g392) & (!sk[76]) & (g393) & (!g394)) + ((g165) & (g166) & (!g392) & (!sk[76]) & (g393) & (g394)) + ((g165) & (g166) & (!g392) & (sk[76]) & (g393) & (!g394)) + ((g165) & (g166) & (!g392) & (sk[76]) & (g393) & (g394)) + ((g165) & (g166) & (g392) & (!sk[76]) & (!g393) & (!g394)) + ((g165) & (g166) & (g392) & (!sk[76]) & (!g393) & (g394)) + ((g165) & (g166) & (g392) & (!sk[76]) & (g393) & (!g394)) + ((g165) & (g166) & (g392) & (!sk[76]) & (g393) & (g394)) + ((g165) & (g166) & (g392) & (sk[76]) & (g393) & (!g394)) + ((g165) & (g166) & (g392) & (sk[76]) & (g393) & (g394)));
	assign g4170 = (((!g2162) & (!sk[77]) & (!g2304) & (g396)) + ((!g2162) & (!sk[77]) & (g2304) & (!g396)) + ((!g2162) & (!sk[77]) & (g2304) & (g396)) + ((!g2162) & (sk[77]) & (!g2304) & (g396)) + ((!g2162) & (sk[77]) & (g2304) & (g396)) + ((g2162) & (!sk[77]) & (!g2304) & (g396)) + ((g2162) & (!sk[77]) & (g2304) & (!g396)) + ((g2162) & (!sk[77]) & (g2304) & (g396)) + ((g2162) & (sk[77]) & (g2304) & (!g396)) + ((g2162) & (sk[77]) & (g2304) & (g396)));
	assign g4171 = (((!g2164) & (!g2304) & (!sk[78]) & (g397)) + ((!g2164) & (!g2304) & (sk[78]) & (g397)) + ((!g2164) & (g2304) & (!sk[78]) & (!g397)) + ((!g2164) & (g2304) & (!sk[78]) & (g397)) + ((!g2164) & (g2304) & (sk[78]) & (g397)) + ((g2164) & (!g2304) & (!sk[78]) & (g397)) + ((g2164) & (g2304) & (!sk[78]) & (!g397)) + ((g2164) & (g2304) & (!sk[78]) & (g397)) + ((g2164) & (g2304) & (sk[78]) & (!g397)) + ((g2164) & (g2304) & (sk[78]) & (g397)));
	assign g4172 = (((!sk[79]) & (!g2166) & (!g2304) & (g398)) + ((!sk[79]) & (!g2166) & (g2304) & (!g398)) + ((!sk[79]) & (!g2166) & (g2304) & (g398)) + ((!sk[79]) & (g2166) & (!g2304) & (g398)) + ((!sk[79]) & (g2166) & (g2304) & (!g398)) + ((!sk[79]) & (g2166) & (g2304) & (g398)) + ((sk[79]) & (!g2166) & (!g2304) & (g398)) + ((sk[79]) & (!g2166) & (g2304) & (g398)) + ((sk[79]) & (g2166) & (g2304) & (!g398)) + ((sk[79]) & (g2166) & (g2304) & (g398)));
	assign g4173 = (((!sk[80]) & (!g2168) & (!g2304) & (g399)) + ((!sk[80]) & (!g2168) & (g2304) & (!g399)) + ((!sk[80]) & (!g2168) & (g2304) & (g399)) + ((!sk[80]) & (g2168) & (!g2304) & (g399)) + ((!sk[80]) & (g2168) & (g2304) & (!g399)) + ((!sk[80]) & (g2168) & (g2304) & (g399)) + ((sk[80]) & (!g2168) & (!g2304) & (g399)) + ((sk[80]) & (!g2168) & (g2304) & (g399)) + ((sk[80]) & (g2168) & (g2304) & (!g399)) + ((sk[80]) & (g2168) & (g2304) & (g399)));
	assign g400 = (((!g396) & (!g397) & (!g398) & (g399) & (g165) & (g166)) + ((!g396) & (!g397) & (g398) & (!g399) & (!g165) & (g166)) + ((!g396) & (!g397) & (g398) & (g399) & (!g165) & (g166)) + ((!g396) & (!g397) & (g398) & (g399) & (g165) & (g166)) + ((!g396) & (g397) & (!g398) & (!g399) & (g165) & (!g166)) + ((!g396) & (g397) & (!g398) & (g399) & (g165) & (!g166)) + ((!g396) & (g397) & (!g398) & (g399) & (g165) & (g166)) + ((!g396) & (g397) & (g398) & (!g399) & (!g165) & (g166)) + ((!g396) & (g397) & (g398) & (!g399) & (g165) & (!g166)) + ((!g396) & (g397) & (g398) & (g399) & (!g165) & (g166)) + ((!g396) & (g397) & (g398) & (g399) & (g165) & (!g166)) + ((!g396) & (g397) & (g398) & (g399) & (g165) & (g166)) + ((g396) & (!g397) & (!g398) & (!g399) & (!g165) & (!g166)) + ((g396) & (!g397) & (!g398) & (g399) & (!g165) & (!g166)) + ((g396) & (!g397) & (!g398) & (g399) & (g165) & (g166)) + ((g396) & (!g397) & (g398) & (!g399) & (!g165) & (!g166)) + ((g396) & (!g397) & (g398) & (!g399) & (!g165) & (g166)) + ((g396) & (!g397) & (g398) & (g399) & (!g165) & (!g166)) + ((g396) & (!g397) & (g398) & (g399) & (!g165) & (g166)) + ((g396) & (!g397) & (g398) & (g399) & (g165) & (g166)) + ((g396) & (g397) & (!g398) & (!g399) & (!g165) & (!g166)) + ((g396) & (g397) & (!g398) & (!g399) & (g165) & (!g166)) + ((g396) & (g397) & (!g398) & (g399) & (!g165) & (!g166)) + ((g396) & (g397) & (!g398) & (g399) & (g165) & (!g166)) + ((g396) & (g397) & (!g398) & (g399) & (g165) & (g166)) + ((g396) & (g397) & (g398) & (!g399) & (!g165) & (!g166)) + ((g396) & (g397) & (g398) & (!g399) & (!g165) & (g166)) + ((g396) & (g397) & (g398) & (!g399) & (g165) & (!g166)) + ((g396) & (g397) & (g398) & (g399) & (!g165) & (!g166)) + ((g396) & (g397) & (g398) & (g399) & (!g165) & (g166)) + ((g396) & (g397) & (g398) & (g399) & (g165) & (!g166)) + ((g396) & (g397) & (g398) & (g399) & (g165) & (g166)));
	assign g4174 = (((!g2169) & (!g2304) & (!sk[82]) & (g401)) + ((!g2169) & (!g2304) & (sk[82]) & (g401)) + ((!g2169) & (g2304) & (!sk[82]) & (!g401)) + ((!g2169) & (g2304) & (!sk[82]) & (g401)) + ((!g2169) & (g2304) & (sk[82]) & (g401)) + ((g2169) & (!g2304) & (!sk[82]) & (g401)) + ((g2169) & (g2304) & (!sk[82]) & (!g401)) + ((g2169) & (g2304) & (!sk[82]) & (g401)) + ((g2169) & (g2304) & (sk[82]) & (!g401)) + ((g2169) & (g2304) & (sk[82]) & (g401)));
	assign g4175 = (((!g2170) & (!sk[83]) & (!g2304) & (g402)) + ((!g2170) & (!sk[83]) & (g2304) & (!g402)) + ((!g2170) & (!sk[83]) & (g2304) & (g402)) + ((!g2170) & (sk[83]) & (!g2304) & (g402)) + ((!g2170) & (sk[83]) & (g2304) & (g402)) + ((g2170) & (!sk[83]) & (!g2304) & (g402)) + ((g2170) & (!sk[83]) & (g2304) & (!g402)) + ((g2170) & (!sk[83]) & (g2304) & (g402)) + ((g2170) & (sk[83]) & (g2304) & (!g402)) + ((g2170) & (sk[83]) & (g2304) & (g402)));
	assign g4176 = (((!sk[84]) & (!g2171) & (!g2304) & (g403)) + ((!sk[84]) & (!g2171) & (g2304) & (!g403)) + ((!sk[84]) & (!g2171) & (g2304) & (g403)) + ((!sk[84]) & (g2171) & (!g2304) & (g403)) + ((!sk[84]) & (g2171) & (g2304) & (!g403)) + ((!sk[84]) & (g2171) & (g2304) & (g403)) + ((sk[84]) & (!g2171) & (!g2304) & (g403)) + ((sk[84]) & (!g2171) & (g2304) & (g403)) + ((sk[84]) & (g2171) & (g2304) & (!g403)) + ((sk[84]) & (g2171) & (g2304) & (g403)));
	assign g4177 = (((!g2172) & (!g2304) & (!sk[85]) & (g404)) + ((!g2172) & (!g2304) & (sk[85]) & (g404)) + ((!g2172) & (g2304) & (!sk[85]) & (!g404)) + ((!g2172) & (g2304) & (!sk[85]) & (g404)) + ((!g2172) & (g2304) & (sk[85]) & (g404)) + ((g2172) & (!g2304) & (!sk[85]) & (g404)) + ((g2172) & (g2304) & (!sk[85]) & (!g404)) + ((g2172) & (g2304) & (!sk[85]) & (g404)) + ((g2172) & (g2304) & (sk[85]) & (!g404)) + ((g2172) & (g2304) & (sk[85]) & (g404)));
	assign g405 = (((!g401) & (!g402) & (!g403) & (g404) & (g165) & (g166)) + ((!g401) & (!g402) & (g403) & (!g404) & (!g165) & (g166)) + ((!g401) & (!g402) & (g403) & (g404) & (!g165) & (g166)) + ((!g401) & (!g402) & (g403) & (g404) & (g165) & (g166)) + ((!g401) & (g402) & (!g403) & (!g404) & (g165) & (!g166)) + ((!g401) & (g402) & (!g403) & (g404) & (g165) & (!g166)) + ((!g401) & (g402) & (!g403) & (g404) & (g165) & (g166)) + ((!g401) & (g402) & (g403) & (!g404) & (!g165) & (g166)) + ((!g401) & (g402) & (g403) & (!g404) & (g165) & (!g166)) + ((!g401) & (g402) & (g403) & (g404) & (!g165) & (g166)) + ((!g401) & (g402) & (g403) & (g404) & (g165) & (!g166)) + ((!g401) & (g402) & (g403) & (g404) & (g165) & (g166)) + ((g401) & (!g402) & (!g403) & (!g404) & (!g165) & (!g166)) + ((g401) & (!g402) & (!g403) & (g404) & (!g165) & (!g166)) + ((g401) & (!g402) & (!g403) & (g404) & (g165) & (g166)) + ((g401) & (!g402) & (g403) & (!g404) & (!g165) & (!g166)) + ((g401) & (!g402) & (g403) & (!g404) & (!g165) & (g166)) + ((g401) & (!g402) & (g403) & (g404) & (!g165) & (!g166)) + ((g401) & (!g402) & (g403) & (g404) & (!g165) & (g166)) + ((g401) & (!g402) & (g403) & (g404) & (g165) & (g166)) + ((g401) & (g402) & (!g403) & (!g404) & (!g165) & (!g166)) + ((g401) & (g402) & (!g403) & (!g404) & (g165) & (!g166)) + ((g401) & (g402) & (!g403) & (g404) & (!g165) & (!g166)) + ((g401) & (g402) & (!g403) & (g404) & (g165) & (!g166)) + ((g401) & (g402) & (!g403) & (g404) & (g165) & (g166)) + ((g401) & (g402) & (g403) & (!g404) & (!g165) & (!g166)) + ((g401) & (g402) & (g403) & (!g404) & (!g165) & (g166)) + ((g401) & (g402) & (g403) & (!g404) & (g165) & (!g166)) + ((g401) & (g402) & (g403) & (g404) & (!g165) & (!g166)) + ((g401) & (g402) & (g403) & (g404) & (!g165) & (g166)) + ((g401) & (g402) & (g403) & (g404) & (g165) & (!g166)) + ((g401) & (g402) & (g403) & (g404) & (g165) & (g166)));
	assign g406 = (((!g147) & (!g148) & (!g391) & (g395) & (!g400) & (!g405)) + ((!g147) & (!g148) & (!g391) & (g395) & (!g400) & (g405)) + ((!g147) & (!g148) & (!g391) & (g395) & (g400) & (!g405)) + ((!g147) & (!g148) & (!g391) & (g395) & (g400) & (g405)) + ((!g147) & (!g148) & (g391) & (g395) & (!g400) & (!g405)) + ((!g147) & (!g148) & (g391) & (g395) & (!g400) & (g405)) + ((!g147) & (!g148) & (g391) & (g395) & (g400) & (!g405)) + ((!g147) & (!g148) & (g391) & (g395) & (g400) & (g405)) + ((!g147) & (g148) & (!g391) & (!g395) & (!g400) & (g405)) + ((!g147) & (g148) & (!g391) & (!g395) & (g400) & (g405)) + ((!g147) & (g148) & (!g391) & (g395) & (!g400) & (g405)) + ((!g147) & (g148) & (!g391) & (g395) & (g400) & (g405)) + ((!g147) & (g148) & (g391) & (!g395) & (!g400) & (g405)) + ((!g147) & (g148) & (g391) & (!g395) & (g400) & (g405)) + ((!g147) & (g148) & (g391) & (g395) & (!g400) & (g405)) + ((!g147) & (g148) & (g391) & (g395) & (g400) & (g405)) + ((g147) & (!g148) & (g391) & (!g395) & (!g400) & (!g405)) + ((g147) & (!g148) & (g391) & (!g395) & (!g400) & (g405)) + ((g147) & (!g148) & (g391) & (!g395) & (g400) & (!g405)) + ((g147) & (!g148) & (g391) & (!g395) & (g400) & (g405)) + ((g147) & (!g148) & (g391) & (g395) & (!g400) & (!g405)) + ((g147) & (!g148) & (g391) & (g395) & (!g400) & (g405)) + ((g147) & (!g148) & (g391) & (g395) & (g400) & (!g405)) + ((g147) & (!g148) & (g391) & (g395) & (g400) & (g405)) + ((g147) & (g148) & (!g391) & (!g395) & (g400) & (!g405)) + ((g147) & (g148) & (!g391) & (!g395) & (g400) & (g405)) + ((g147) & (g148) & (!g391) & (g395) & (g400) & (!g405)) + ((g147) & (g148) & (!g391) & (g395) & (g400) & (g405)) + ((g147) & (g148) & (g391) & (!g395) & (g400) & (!g405)) + ((g147) & (g148) & (g391) & (!g395) & (g400) & (g405)) + ((g147) & (g148) & (g391) & (g395) & (g400) & (!g405)) + ((g147) & (g148) & (g391) & (g395) & (g400) & (g405)));
	assign g407 = (((!sk[88]) & (!g142) & (!g386) & (g406)) + ((!sk[88]) & (!g142) & (g386) & (!g406)) + ((!sk[88]) & (!g142) & (g386) & (g406)) + ((!sk[88]) & (g142) & (!g386) & (g406)) + ((!sk[88]) & (g142) & (g386) & (!g406)) + ((!sk[88]) & (g142) & (g386) & (g406)) + ((sk[88]) & (!g142) & (!g386) & (g406)) + ((sk[88]) & (!g142) & (g386) & (g406)) + ((sk[88]) & (g142) & (g386) & (!g406)) + ((sk[88]) & (g142) & (g386) & (g406)));
	assign g4178 = (((!sk[89]) & (!g2059) & (!g2311) & (g408)) + ((!sk[89]) & (!g2059) & (g2311) & (!g408)) + ((!sk[89]) & (!g2059) & (g2311) & (g408)) + ((!sk[89]) & (g2059) & (!g2311) & (g408)) + ((!sk[89]) & (g2059) & (g2311) & (!g408)) + ((!sk[89]) & (g2059) & (g2311) & (g408)) + ((sk[89]) & (!g2059) & (!g2311) & (g408)) + ((sk[89]) & (!g2059) & (g2311) & (g408)) + ((sk[89]) & (g2059) & (g2311) & (!g408)) + ((sk[89]) & (g2059) & (g2311) & (g408)));
	assign g409 = (((!sk[90]) & (!g318) & (!g364) & (!g320) & (g362) & (!g407)) + ((!sk[90]) & (!g318) & (!g364) & (!g320) & (g362) & (g407)) + ((!sk[90]) & (!g318) & (!g364) & (g320) & (!g362) & (!g407)) + ((!sk[90]) & (!g318) & (!g364) & (g320) & (!g362) & (g407)) + ((!sk[90]) & (!g318) & (!g364) & (g320) & (g362) & (!g407)) + ((!sk[90]) & (!g318) & (!g364) & (g320) & (g362) & (g407)) + ((!sk[90]) & (!g318) & (g364) & (!g320) & (!g362) & (!g407)) + ((!sk[90]) & (!g318) & (g364) & (!g320) & (!g362) & (g407)) + ((!sk[90]) & (!g318) & (g364) & (!g320) & (g362) & (!g407)) + ((!sk[90]) & (!g318) & (g364) & (!g320) & (g362) & (g407)) + ((!sk[90]) & (!g318) & (g364) & (g320) & (!g362) & (!g407)) + ((!sk[90]) & (!g318) & (g364) & (g320) & (!g362) & (g407)) + ((!sk[90]) & (!g318) & (g364) & (g320) & (g362) & (!g407)) + ((!sk[90]) & (!g318) & (g364) & (g320) & (g362) & (g407)) + ((!sk[90]) & (g318) & (!g364) & (!g320) & (g362) & (!g407)) + ((!sk[90]) & (g318) & (!g364) & (!g320) & (g362) & (g407)) + ((!sk[90]) & (g318) & (!g364) & (g320) & (!g362) & (!g407)) + ((!sk[90]) & (g318) & (!g364) & (g320) & (!g362) & (g407)) + ((!sk[90]) & (g318) & (!g364) & (g320) & (g362) & (!g407)) + ((!sk[90]) & (g318) & (!g364) & (g320) & (g362) & (g407)) + ((!sk[90]) & (g318) & (g364) & (!g320) & (!g362) & (!g407)) + ((!sk[90]) & (g318) & (g364) & (!g320) & (!g362) & (g407)) + ((!sk[90]) & (g318) & (g364) & (!g320) & (g362) & (!g407)) + ((!sk[90]) & (g318) & (g364) & (!g320) & (g362) & (g407)) + ((!sk[90]) & (g318) & (g364) & (g320) & (!g362) & (!g407)) + ((!sk[90]) & (g318) & (g364) & (g320) & (!g362) & (g407)) + ((!sk[90]) & (g318) & (g364) & (g320) & (g362) & (!g407)) + ((!sk[90]) & (g318) & (g364) & (g320) & (g362) & (g407)) + ((sk[90]) & (!g318) & (!g364) & (g320) & (g362) & (g407)) + ((sk[90]) & (!g318) & (g364) & (!g320) & (!g362) & (g407)) + ((sk[90]) & (!g318) & (g364) & (!g320) & (g362) & (g407)) + ((sk[90]) & (!g318) & (g364) & (g320) & (!g362) & (g407)) + ((sk[90]) & (!g318) & (g364) & (g320) & (g362) & (!g407)) + ((sk[90]) & (!g318) & (g364) & (g320) & (g362) & (g407)) + ((sk[90]) & (g318) & (!g364) & (!g320) & (g362) & (g407)) + ((sk[90]) & (g318) & (!g364) & (g320) & (!g362) & (g407)) + ((sk[90]) & (g318) & (!g364) & (g320) & (g362) & (g407)) + ((sk[90]) & (g318) & (g364) & (!g320) & (!g362) & (g407)) + ((sk[90]) & (g318) & (g364) & (!g320) & (g362) & (!g407)) + ((sk[90]) & (g318) & (g364) & (!g320) & (g362) & (g407)) + ((sk[90]) & (g318) & (g364) & (g320) & (!g362) & (!g407)) + ((sk[90]) & (g318) & (g364) & (g320) & (!g362) & (g407)) + ((sk[90]) & (g318) & (g364) & (g320) & (g362) & (!g407)) + ((sk[90]) & (g318) & (g364) & (g320) & (g362) & (g407)));
	assign g4179 = (((!g2140) & (!sk[91]) & (!g2328) & (g410)) + ((!g2140) & (!sk[91]) & (g2328) & (!g410)) + ((!g2140) & (!sk[91]) & (g2328) & (g410)) + ((!g2140) & (sk[91]) & (!g2328) & (g410)) + ((!g2140) & (sk[91]) & (g2328) & (g410)) + ((g2140) & (!sk[91]) & (!g2328) & (g410)) + ((g2140) & (!sk[91]) & (g2328) & (!g410)) + ((g2140) & (!sk[91]) & (g2328) & (g410)) + ((g2140) & (sk[91]) & (g2328) & (!g410)) + ((g2140) & (sk[91]) & (g2328) & (g410)));
	assign g4180 = (((!sk[92]) & (!g2142) & (!g2328) & (g411)) + ((!sk[92]) & (!g2142) & (g2328) & (!g411)) + ((!sk[92]) & (!g2142) & (g2328) & (g411)) + ((!sk[92]) & (g2142) & (!g2328) & (g411)) + ((!sk[92]) & (g2142) & (g2328) & (!g411)) + ((!sk[92]) & (g2142) & (g2328) & (g411)) + ((sk[92]) & (!g2142) & (!g2328) & (g411)) + ((sk[92]) & (!g2142) & (g2328) & (g411)) + ((sk[92]) & (g2142) & (g2328) & (!g411)) + ((sk[92]) & (g2142) & (g2328) & (g411)));
	assign g4181 = (((!g2144) & (!g2328) & (!sk[93]) & (g412)) + ((!g2144) & (!g2328) & (sk[93]) & (g412)) + ((!g2144) & (g2328) & (!sk[93]) & (!g412)) + ((!g2144) & (g2328) & (!sk[93]) & (g412)) + ((!g2144) & (g2328) & (sk[93]) & (g412)) + ((g2144) & (!g2328) & (!sk[93]) & (g412)) + ((g2144) & (g2328) & (!sk[93]) & (!g412)) + ((g2144) & (g2328) & (!sk[93]) & (g412)) + ((g2144) & (g2328) & (sk[93]) & (!g412)) + ((g2144) & (g2328) & (sk[93]) & (g412)));
	assign g4182 = (((!g2145) & (!sk[94]) & (!g2328) & (g413)) + ((!g2145) & (!sk[94]) & (g2328) & (!g413)) + ((!g2145) & (!sk[94]) & (g2328) & (g413)) + ((!g2145) & (sk[94]) & (!g2328) & (g413)) + ((!g2145) & (sk[94]) & (g2328) & (g413)) + ((g2145) & (!sk[94]) & (!g2328) & (g413)) + ((g2145) & (!sk[94]) & (g2328) & (!g413)) + ((g2145) & (!sk[94]) & (g2328) & (g413)) + ((g2145) & (sk[94]) & (g2328) & (!g413)) + ((g2145) & (sk[94]) & (g2328) & (g413)));
	assign g414 = (((!g410) & (!g411) & (!g412) & (g413) & (g147) & (g148)) + ((!g410) & (!g411) & (g412) & (!g413) & (!g147) & (g148)) + ((!g410) & (!g411) & (g412) & (g413) & (!g147) & (g148)) + ((!g410) & (!g411) & (g412) & (g413) & (g147) & (g148)) + ((!g410) & (g411) & (!g412) & (!g413) & (g147) & (!g148)) + ((!g410) & (g411) & (!g412) & (g413) & (g147) & (!g148)) + ((!g410) & (g411) & (!g412) & (g413) & (g147) & (g148)) + ((!g410) & (g411) & (g412) & (!g413) & (!g147) & (g148)) + ((!g410) & (g411) & (g412) & (!g413) & (g147) & (!g148)) + ((!g410) & (g411) & (g412) & (g413) & (!g147) & (g148)) + ((!g410) & (g411) & (g412) & (g413) & (g147) & (!g148)) + ((!g410) & (g411) & (g412) & (g413) & (g147) & (g148)) + ((g410) & (!g411) & (!g412) & (!g413) & (!g147) & (!g148)) + ((g410) & (!g411) & (!g412) & (g413) & (!g147) & (!g148)) + ((g410) & (!g411) & (!g412) & (g413) & (g147) & (g148)) + ((g410) & (!g411) & (g412) & (!g413) & (!g147) & (!g148)) + ((g410) & (!g411) & (g412) & (!g413) & (!g147) & (g148)) + ((g410) & (!g411) & (g412) & (g413) & (!g147) & (!g148)) + ((g410) & (!g411) & (g412) & (g413) & (!g147) & (g148)) + ((g410) & (!g411) & (g412) & (g413) & (g147) & (g148)) + ((g410) & (g411) & (!g412) & (!g413) & (!g147) & (!g148)) + ((g410) & (g411) & (!g412) & (!g413) & (g147) & (!g148)) + ((g410) & (g411) & (!g412) & (g413) & (!g147) & (!g148)) + ((g410) & (g411) & (!g412) & (g413) & (g147) & (!g148)) + ((g410) & (g411) & (!g412) & (g413) & (g147) & (g148)) + ((g410) & (g411) & (g412) & (!g413) & (!g147) & (!g148)) + ((g410) & (g411) & (g412) & (!g413) & (!g147) & (g148)) + ((g410) & (g411) & (g412) & (!g413) & (g147) & (!g148)) + ((g410) & (g411) & (g412) & (g413) & (!g147) & (!g148)) + ((g410) & (g411) & (g412) & (g413) & (!g147) & (g148)) + ((g410) & (g411) & (g412) & (g413) & (g147) & (!g148)) + ((g410) & (g411) & (g412) & (g413) & (g147) & (g148)));
	assign g4183 = (((!g2146) & (!g2328) & (!sk[96]) & (g415)) + ((!g2146) & (!g2328) & (sk[96]) & (g415)) + ((!g2146) & (g2328) & (!sk[96]) & (!g415)) + ((!g2146) & (g2328) & (!sk[96]) & (g415)) + ((!g2146) & (g2328) & (sk[96]) & (g415)) + ((g2146) & (!g2328) & (!sk[96]) & (g415)) + ((g2146) & (g2328) & (!sk[96]) & (!g415)) + ((g2146) & (g2328) & (!sk[96]) & (g415)) + ((g2146) & (g2328) & (sk[96]) & (!g415)) + ((g2146) & (g2328) & (sk[96]) & (g415)));
	assign g4184 = (((!g2148) & (!g2328) & (!sk[97]) & (g416)) + ((!g2148) & (!g2328) & (sk[97]) & (g416)) + ((!g2148) & (g2328) & (!sk[97]) & (!g416)) + ((!g2148) & (g2328) & (!sk[97]) & (g416)) + ((!g2148) & (g2328) & (sk[97]) & (g416)) + ((g2148) & (!g2328) & (!sk[97]) & (g416)) + ((g2148) & (g2328) & (!sk[97]) & (!g416)) + ((g2148) & (g2328) & (!sk[97]) & (g416)) + ((g2148) & (g2328) & (sk[97]) & (!g416)) + ((g2148) & (g2328) & (sk[97]) & (g416)));
	assign g4185 = (((!g2150) & (!g2328) & (!sk[98]) & (g417)) + ((!g2150) & (!g2328) & (sk[98]) & (g417)) + ((!g2150) & (g2328) & (!sk[98]) & (!g417)) + ((!g2150) & (g2328) & (!sk[98]) & (g417)) + ((!g2150) & (g2328) & (sk[98]) & (g417)) + ((g2150) & (!g2328) & (!sk[98]) & (g417)) + ((g2150) & (g2328) & (!sk[98]) & (!g417)) + ((g2150) & (g2328) & (!sk[98]) & (g417)) + ((g2150) & (g2328) & (sk[98]) & (!g417)) + ((g2150) & (g2328) & (sk[98]) & (g417)));
	assign g4186 = (((!g2151) & (!g2328) & (!sk[99]) & (g418)) + ((!g2151) & (!g2328) & (sk[99]) & (g418)) + ((!g2151) & (g2328) & (!sk[99]) & (!g418)) + ((!g2151) & (g2328) & (!sk[99]) & (g418)) + ((!g2151) & (g2328) & (sk[99]) & (g418)) + ((g2151) & (!g2328) & (!sk[99]) & (g418)) + ((g2151) & (g2328) & (!sk[99]) & (!g418)) + ((g2151) & (g2328) & (!sk[99]) & (g418)) + ((g2151) & (g2328) & (sk[99]) & (!g418)) + ((g2151) & (g2328) & (sk[99]) & (g418)));
	assign g419 = (((!g415) & (!g416) & (!g417) & (g418) & (g147) & (g148)) + ((!g415) & (!g416) & (g417) & (!g418) & (!g147) & (g148)) + ((!g415) & (!g416) & (g417) & (g418) & (!g147) & (g148)) + ((!g415) & (!g416) & (g417) & (g418) & (g147) & (g148)) + ((!g415) & (g416) & (!g417) & (!g418) & (g147) & (!g148)) + ((!g415) & (g416) & (!g417) & (g418) & (g147) & (!g148)) + ((!g415) & (g416) & (!g417) & (g418) & (g147) & (g148)) + ((!g415) & (g416) & (g417) & (!g418) & (!g147) & (g148)) + ((!g415) & (g416) & (g417) & (!g418) & (g147) & (!g148)) + ((!g415) & (g416) & (g417) & (g418) & (!g147) & (g148)) + ((!g415) & (g416) & (g417) & (g418) & (g147) & (!g148)) + ((!g415) & (g416) & (g417) & (g418) & (g147) & (g148)) + ((g415) & (!g416) & (!g417) & (!g418) & (!g147) & (!g148)) + ((g415) & (!g416) & (!g417) & (g418) & (!g147) & (!g148)) + ((g415) & (!g416) & (!g417) & (g418) & (g147) & (g148)) + ((g415) & (!g416) & (g417) & (!g418) & (!g147) & (!g148)) + ((g415) & (!g416) & (g417) & (!g418) & (!g147) & (g148)) + ((g415) & (!g416) & (g417) & (g418) & (!g147) & (!g148)) + ((g415) & (!g416) & (g417) & (g418) & (!g147) & (g148)) + ((g415) & (!g416) & (g417) & (g418) & (g147) & (g148)) + ((g415) & (g416) & (!g417) & (!g418) & (!g147) & (!g148)) + ((g415) & (g416) & (!g417) & (!g418) & (g147) & (!g148)) + ((g415) & (g416) & (!g417) & (g418) & (!g147) & (!g148)) + ((g415) & (g416) & (!g417) & (g418) & (g147) & (!g148)) + ((g415) & (g416) & (!g417) & (g418) & (g147) & (g148)) + ((g415) & (g416) & (g417) & (!g418) & (!g147) & (!g148)) + ((g415) & (g416) & (g417) & (!g418) & (!g147) & (g148)) + ((g415) & (g416) & (g417) & (!g418) & (g147) & (!g148)) + ((g415) & (g416) & (g417) & (g418) & (!g147) & (!g148)) + ((g415) & (g416) & (g417) & (g418) & (!g147) & (g148)) + ((g415) & (g416) & (g417) & (g418) & (g147) & (!g148)) + ((g415) & (g416) & (g417) & (g418) & (g147) & (g148)));
	assign g4187 = (((!g2152) & (!sk[101]) & (!g2328) & (g420)) + ((!g2152) & (!sk[101]) & (g2328) & (!g420)) + ((!g2152) & (!sk[101]) & (g2328) & (g420)) + ((!g2152) & (sk[101]) & (!g2328) & (g420)) + ((!g2152) & (sk[101]) & (g2328) & (g420)) + ((g2152) & (!sk[101]) & (!g2328) & (g420)) + ((g2152) & (!sk[101]) & (g2328) & (!g420)) + ((g2152) & (!sk[101]) & (g2328) & (g420)) + ((g2152) & (sk[101]) & (g2328) & (!g420)) + ((g2152) & (sk[101]) & (g2328) & (g420)));
	assign g4188 = (((!sk[102]) & (!g2153) & (!g2328) & (g421)) + ((!sk[102]) & (!g2153) & (g2328) & (!g421)) + ((!sk[102]) & (!g2153) & (g2328) & (g421)) + ((!sk[102]) & (g2153) & (!g2328) & (g421)) + ((!sk[102]) & (g2153) & (g2328) & (!g421)) + ((!sk[102]) & (g2153) & (g2328) & (g421)) + ((sk[102]) & (!g2153) & (!g2328) & (g421)) + ((sk[102]) & (!g2153) & (g2328) & (g421)) + ((sk[102]) & (g2153) & (g2328) & (!g421)) + ((sk[102]) & (g2153) & (g2328) & (g421)));
	assign g4189 = (((!g2155) & (!g2328) & (!sk[103]) & (g422)) + ((!g2155) & (!g2328) & (sk[103]) & (g422)) + ((!g2155) & (g2328) & (!sk[103]) & (!g422)) + ((!g2155) & (g2328) & (!sk[103]) & (g422)) + ((!g2155) & (g2328) & (sk[103]) & (g422)) + ((g2155) & (!g2328) & (!sk[103]) & (g422)) + ((g2155) & (g2328) & (!sk[103]) & (!g422)) + ((g2155) & (g2328) & (!sk[103]) & (g422)) + ((g2155) & (g2328) & (sk[103]) & (!g422)) + ((g2155) & (g2328) & (sk[103]) & (g422)));
	assign g4190 = (((!sk[104]) & (!g2157) & (!g2328) & (g423)) + ((!sk[104]) & (!g2157) & (g2328) & (!g423)) + ((!sk[104]) & (!g2157) & (g2328) & (g423)) + ((!sk[104]) & (g2157) & (!g2328) & (g423)) + ((!sk[104]) & (g2157) & (g2328) & (!g423)) + ((!sk[104]) & (g2157) & (g2328) & (g423)) + ((sk[104]) & (!g2157) & (!g2328) & (g423)) + ((sk[104]) & (!g2157) & (g2328) & (g423)) + ((sk[104]) & (g2157) & (g2328) & (!g423)) + ((sk[104]) & (g2157) & (g2328) & (g423)));
	assign g424 = (((!g420) & (!g421) & (!g422) & (g423) & (g147) & (g148)) + ((!g420) & (!g421) & (g422) & (!g423) & (!g147) & (g148)) + ((!g420) & (!g421) & (g422) & (g423) & (!g147) & (g148)) + ((!g420) & (!g421) & (g422) & (g423) & (g147) & (g148)) + ((!g420) & (g421) & (!g422) & (!g423) & (g147) & (!g148)) + ((!g420) & (g421) & (!g422) & (g423) & (g147) & (!g148)) + ((!g420) & (g421) & (!g422) & (g423) & (g147) & (g148)) + ((!g420) & (g421) & (g422) & (!g423) & (!g147) & (g148)) + ((!g420) & (g421) & (g422) & (!g423) & (g147) & (!g148)) + ((!g420) & (g421) & (g422) & (g423) & (!g147) & (g148)) + ((!g420) & (g421) & (g422) & (g423) & (g147) & (!g148)) + ((!g420) & (g421) & (g422) & (g423) & (g147) & (g148)) + ((g420) & (!g421) & (!g422) & (!g423) & (!g147) & (!g148)) + ((g420) & (!g421) & (!g422) & (g423) & (!g147) & (!g148)) + ((g420) & (!g421) & (!g422) & (g423) & (g147) & (g148)) + ((g420) & (!g421) & (g422) & (!g423) & (!g147) & (!g148)) + ((g420) & (!g421) & (g422) & (!g423) & (!g147) & (g148)) + ((g420) & (!g421) & (g422) & (g423) & (!g147) & (!g148)) + ((g420) & (!g421) & (g422) & (g423) & (!g147) & (g148)) + ((g420) & (!g421) & (g422) & (g423) & (g147) & (g148)) + ((g420) & (g421) & (!g422) & (!g423) & (!g147) & (!g148)) + ((g420) & (g421) & (!g422) & (!g423) & (g147) & (!g148)) + ((g420) & (g421) & (!g422) & (g423) & (!g147) & (!g148)) + ((g420) & (g421) & (!g422) & (g423) & (g147) & (!g148)) + ((g420) & (g421) & (!g422) & (g423) & (g147) & (g148)) + ((g420) & (g421) & (g422) & (!g423) & (!g147) & (!g148)) + ((g420) & (g421) & (g422) & (!g423) & (!g147) & (g148)) + ((g420) & (g421) & (g422) & (!g423) & (g147) & (!g148)) + ((g420) & (g421) & (g422) & (g423) & (!g147) & (!g148)) + ((g420) & (g421) & (g422) & (g423) & (!g147) & (g148)) + ((g420) & (g421) & (g422) & (g423) & (g147) & (!g148)) + ((g420) & (g421) & (g422) & (g423) & (g147) & (g148)));
	assign g4191 = (((!g2158) & (!sk[106]) & (!g2328) & (g425)) + ((!g2158) & (!sk[106]) & (g2328) & (!g425)) + ((!g2158) & (!sk[106]) & (g2328) & (g425)) + ((!g2158) & (sk[106]) & (!g2328) & (g425)) + ((!g2158) & (sk[106]) & (g2328) & (g425)) + ((g2158) & (!sk[106]) & (!g2328) & (g425)) + ((g2158) & (!sk[106]) & (g2328) & (!g425)) + ((g2158) & (!sk[106]) & (g2328) & (g425)) + ((g2158) & (sk[106]) & (g2328) & (!g425)) + ((g2158) & (sk[106]) & (g2328) & (g425)));
	assign g4192 = (((!sk[107]) & (!g2159) & (!g2328) & (g426)) + ((!sk[107]) & (!g2159) & (g2328) & (!g426)) + ((!sk[107]) & (!g2159) & (g2328) & (g426)) + ((!sk[107]) & (g2159) & (!g2328) & (g426)) + ((!sk[107]) & (g2159) & (g2328) & (!g426)) + ((!sk[107]) & (g2159) & (g2328) & (g426)) + ((sk[107]) & (!g2159) & (!g2328) & (g426)) + ((sk[107]) & (!g2159) & (g2328) & (g426)) + ((sk[107]) & (g2159) & (g2328) & (!g426)) + ((sk[107]) & (g2159) & (g2328) & (g426)));
	assign g4193 = (((!g2160) & (!sk[108]) & (!g2328) & (g427)) + ((!g2160) & (!sk[108]) & (g2328) & (!g427)) + ((!g2160) & (!sk[108]) & (g2328) & (g427)) + ((!g2160) & (sk[108]) & (!g2328) & (g427)) + ((!g2160) & (sk[108]) & (g2328) & (g427)) + ((g2160) & (!sk[108]) & (!g2328) & (g427)) + ((g2160) & (!sk[108]) & (g2328) & (!g427)) + ((g2160) & (!sk[108]) & (g2328) & (g427)) + ((g2160) & (sk[108]) & (g2328) & (!g427)) + ((g2160) & (sk[108]) & (g2328) & (g427)));
	assign g4194 = (((!g2161) & (!sk[109]) & (!g2328) & (g428)) + ((!g2161) & (!sk[109]) & (g2328) & (!g428)) + ((!g2161) & (!sk[109]) & (g2328) & (g428)) + ((!g2161) & (sk[109]) & (!g2328) & (g428)) + ((!g2161) & (sk[109]) & (g2328) & (g428)) + ((g2161) & (!sk[109]) & (!g2328) & (g428)) + ((g2161) & (!sk[109]) & (g2328) & (!g428)) + ((g2161) & (!sk[109]) & (g2328) & (g428)) + ((g2161) & (sk[109]) & (g2328) & (!g428)) + ((g2161) & (sk[109]) & (g2328) & (g428)));
	assign g429 = (((!g425) & (!g426) & (!g427) & (g428) & (g147) & (g148)) + ((!g425) & (!g426) & (g427) & (!g428) & (!g147) & (g148)) + ((!g425) & (!g426) & (g427) & (g428) & (!g147) & (g148)) + ((!g425) & (!g426) & (g427) & (g428) & (g147) & (g148)) + ((!g425) & (g426) & (!g427) & (!g428) & (g147) & (!g148)) + ((!g425) & (g426) & (!g427) & (g428) & (g147) & (!g148)) + ((!g425) & (g426) & (!g427) & (g428) & (g147) & (g148)) + ((!g425) & (g426) & (g427) & (!g428) & (!g147) & (g148)) + ((!g425) & (g426) & (g427) & (!g428) & (g147) & (!g148)) + ((!g425) & (g426) & (g427) & (g428) & (!g147) & (g148)) + ((!g425) & (g426) & (g427) & (g428) & (g147) & (!g148)) + ((!g425) & (g426) & (g427) & (g428) & (g147) & (g148)) + ((g425) & (!g426) & (!g427) & (!g428) & (!g147) & (!g148)) + ((g425) & (!g426) & (!g427) & (g428) & (!g147) & (!g148)) + ((g425) & (!g426) & (!g427) & (g428) & (g147) & (g148)) + ((g425) & (!g426) & (g427) & (!g428) & (!g147) & (!g148)) + ((g425) & (!g426) & (g427) & (!g428) & (!g147) & (g148)) + ((g425) & (!g426) & (g427) & (g428) & (!g147) & (!g148)) + ((g425) & (!g426) & (g427) & (g428) & (!g147) & (g148)) + ((g425) & (!g426) & (g427) & (g428) & (g147) & (g148)) + ((g425) & (g426) & (!g427) & (!g428) & (!g147) & (!g148)) + ((g425) & (g426) & (!g427) & (!g428) & (g147) & (!g148)) + ((g425) & (g426) & (!g427) & (g428) & (!g147) & (!g148)) + ((g425) & (g426) & (!g427) & (g428) & (g147) & (!g148)) + ((g425) & (g426) & (!g427) & (g428) & (g147) & (g148)) + ((g425) & (g426) & (g427) & (!g428) & (!g147) & (!g148)) + ((g425) & (g426) & (g427) & (!g428) & (!g147) & (g148)) + ((g425) & (g426) & (g427) & (!g428) & (g147) & (!g148)) + ((g425) & (g426) & (g427) & (g428) & (!g147) & (!g148)) + ((g425) & (g426) & (g427) & (g428) & (!g147) & (g148)) + ((g425) & (g426) & (g427) & (g428) & (g147) & (!g148)) + ((g425) & (g426) & (g427) & (g428) & (g147) & (g148)));
	assign g430 = (((!g414) & (!g419) & (!g424) & (g429) & (g165) & (g166)) + ((!g414) & (!g419) & (g424) & (!g429) & (!g165) & (g166)) + ((!g414) & (!g419) & (g424) & (g429) & (!g165) & (g166)) + ((!g414) & (!g419) & (g424) & (g429) & (g165) & (g166)) + ((!g414) & (g419) & (!g424) & (!g429) & (g165) & (!g166)) + ((!g414) & (g419) & (!g424) & (g429) & (g165) & (!g166)) + ((!g414) & (g419) & (!g424) & (g429) & (g165) & (g166)) + ((!g414) & (g419) & (g424) & (!g429) & (!g165) & (g166)) + ((!g414) & (g419) & (g424) & (!g429) & (g165) & (!g166)) + ((!g414) & (g419) & (g424) & (g429) & (!g165) & (g166)) + ((!g414) & (g419) & (g424) & (g429) & (g165) & (!g166)) + ((!g414) & (g419) & (g424) & (g429) & (g165) & (g166)) + ((g414) & (!g419) & (!g424) & (!g429) & (!g165) & (!g166)) + ((g414) & (!g419) & (!g424) & (g429) & (!g165) & (!g166)) + ((g414) & (!g419) & (!g424) & (g429) & (g165) & (g166)) + ((g414) & (!g419) & (g424) & (!g429) & (!g165) & (!g166)) + ((g414) & (!g419) & (g424) & (!g429) & (!g165) & (g166)) + ((g414) & (!g419) & (g424) & (g429) & (!g165) & (!g166)) + ((g414) & (!g419) & (g424) & (g429) & (!g165) & (g166)) + ((g414) & (!g419) & (g424) & (g429) & (g165) & (g166)) + ((g414) & (g419) & (!g424) & (!g429) & (!g165) & (!g166)) + ((g414) & (g419) & (!g424) & (!g429) & (g165) & (!g166)) + ((g414) & (g419) & (!g424) & (g429) & (!g165) & (!g166)) + ((g414) & (g419) & (!g424) & (g429) & (g165) & (!g166)) + ((g414) & (g419) & (!g424) & (g429) & (g165) & (g166)) + ((g414) & (g419) & (g424) & (!g429) & (!g165) & (!g166)) + ((g414) & (g419) & (g424) & (!g429) & (!g165) & (g166)) + ((g414) & (g419) & (g424) & (!g429) & (g165) & (!g166)) + ((g414) & (g419) & (g424) & (g429) & (!g165) & (!g166)) + ((g414) & (g419) & (g424) & (g429) & (!g165) & (g166)) + ((g414) & (g419) & (g424) & (g429) & (g165) & (!g166)) + ((g414) & (g419) & (g424) & (g429) & (g165) & (g166)));
	assign g4195 = (((!g2173) & (!sk[112]) & (!g2328) & (g431)) + ((!g2173) & (!sk[112]) & (g2328) & (!g431)) + ((!g2173) & (!sk[112]) & (g2328) & (g431)) + ((!g2173) & (sk[112]) & (!g2328) & (g431)) + ((!g2173) & (sk[112]) & (g2328) & (g431)) + ((g2173) & (!sk[112]) & (!g2328) & (g431)) + ((g2173) & (!sk[112]) & (g2328) & (!g431)) + ((g2173) & (!sk[112]) & (g2328) & (g431)) + ((g2173) & (sk[112]) & (g2328) & (!g431)) + ((g2173) & (sk[112]) & (g2328) & (g431)));
	assign g4196 = (((!g2174) & (!g2328) & (!sk[113]) & (g432)) + ((!g2174) & (!g2328) & (sk[113]) & (g432)) + ((!g2174) & (g2328) & (!sk[113]) & (!g432)) + ((!g2174) & (g2328) & (!sk[113]) & (g432)) + ((!g2174) & (g2328) & (sk[113]) & (g432)) + ((g2174) & (!g2328) & (!sk[113]) & (g432)) + ((g2174) & (g2328) & (!sk[113]) & (!g432)) + ((g2174) & (g2328) & (!sk[113]) & (g432)) + ((g2174) & (g2328) & (sk[113]) & (!g432)) + ((g2174) & (g2328) & (sk[113]) & (g432)));
	assign g4197 = (((!g2175) & (!sk[114]) & (!g2328) & (g433)) + ((!g2175) & (!sk[114]) & (g2328) & (!g433)) + ((!g2175) & (!sk[114]) & (g2328) & (g433)) + ((!g2175) & (sk[114]) & (!g2328) & (g433)) + ((!g2175) & (sk[114]) & (g2328) & (g433)) + ((g2175) & (!sk[114]) & (!g2328) & (g433)) + ((g2175) & (!sk[114]) & (g2328) & (!g433)) + ((g2175) & (!sk[114]) & (g2328) & (g433)) + ((g2175) & (sk[114]) & (g2328) & (!g433)) + ((g2175) & (sk[114]) & (g2328) & (g433)));
	assign g4198 = (((!g2176) & (!g2328) & (!sk[115]) & (g434)) + ((!g2176) & (!g2328) & (sk[115]) & (g434)) + ((!g2176) & (g2328) & (!sk[115]) & (!g434)) + ((!g2176) & (g2328) & (!sk[115]) & (g434)) + ((!g2176) & (g2328) & (sk[115]) & (g434)) + ((g2176) & (!g2328) & (!sk[115]) & (g434)) + ((g2176) & (g2328) & (!sk[115]) & (!g434)) + ((g2176) & (g2328) & (!sk[115]) & (g434)) + ((g2176) & (g2328) & (sk[115]) & (!g434)) + ((g2176) & (g2328) & (sk[115]) & (g434)));
	assign g435 = (((!g431) & (!g432) & (!g433) & (g434) & (g165) & (g166)) + ((!g431) & (!g432) & (g433) & (!g434) & (!g165) & (g166)) + ((!g431) & (!g432) & (g433) & (g434) & (!g165) & (g166)) + ((!g431) & (!g432) & (g433) & (g434) & (g165) & (g166)) + ((!g431) & (g432) & (!g433) & (!g434) & (g165) & (!g166)) + ((!g431) & (g432) & (!g433) & (g434) & (g165) & (!g166)) + ((!g431) & (g432) & (!g433) & (g434) & (g165) & (g166)) + ((!g431) & (g432) & (g433) & (!g434) & (!g165) & (g166)) + ((!g431) & (g432) & (g433) & (!g434) & (g165) & (!g166)) + ((!g431) & (g432) & (g433) & (g434) & (!g165) & (g166)) + ((!g431) & (g432) & (g433) & (g434) & (g165) & (!g166)) + ((!g431) & (g432) & (g433) & (g434) & (g165) & (g166)) + ((g431) & (!g432) & (!g433) & (!g434) & (!g165) & (!g166)) + ((g431) & (!g432) & (!g433) & (g434) & (!g165) & (!g166)) + ((g431) & (!g432) & (!g433) & (g434) & (g165) & (g166)) + ((g431) & (!g432) & (g433) & (!g434) & (!g165) & (!g166)) + ((g431) & (!g432) & (g433) & (!g434) & (!g165) & (g166)) + ((g431) & (!g432) & (g433) & (g434) & (!g165) & (!g166)) + ((g431) & (!g432) & (g433) & (g434) & (!g165) & (g166)) + ((g431) & (!g432) & (g433) & (g434) & (g165) & (g166)) + ((g431) & (g432) & (!g433) & (!g434) & (!g165) & (!g166)) + ((g431) & (g432) & (!g433) & (!g434) & (g165) & (!g166)) + ((g431) & (g432) & (!g433) & (g434) & (!g165) & (!g166)) + ((g431) & (g432) & (!g433) & (g434) & (g165) & (!g166)) + ((g431) & (g432) & (!g433) & (g434) & (g165) & (g166)) + ((g431) & (g432) & (g433) & (!g434) & (!g165) & (!g166)) + ((g431) & (g432) & (g433) & (!g434) & (!g165) & (g166)) + ((g431) & (g432) & (g433) & (!g434) & (g165) & (!g166)) + ((g431) & (g432) & (g433) & (g434) & (!g165) & (!g166)) + ((g431) & (g432) & (g433) & (g434) & (!g165) & (g166)) + ((g431) & (g432) & (g433) & (g434) & (g165) & (!g166)) + ((g431) & (g432) & (g433) & (g434) & (g165) & (g166)));
	assign g4199 = (((!g2177) & (!g2328) & (!sk[117]) & (g436)) + ((!g2177) & (!g2328) & (sk[117]) & (g436)) + ((!g2177) & (g2328) & (!sk[117]) & (!g436)) + ((!g2177) & (g2328) & (!sk[117]) & (g436)) + ((!g2177) & (g2328) & (sk[117]) & (g436)) + ((g2177) & (!g2328) & (!sk[117]) & (g436)) + ((g2177) & (g2328) & (!sk[117]) & (!g436)) + ((g2177) & (g2328) & (!sk[117]) & (g436)) + ((g2177) & (g2328) & (sk[117]) & (!g436)) + ((g2177) & (g2328) & (sk[117]) & (g436)));
	assign g4200 = (((!g2178) & (!g2328) & (!sk[118]) & (g437)) + ((!g2178) & (!g2328) & (sk[118]) & (g437)) + ((!g2178) & (g2328) & (!sk[118]) & (!g437)) + ((!g2178) & (g2328) & (!sk[118]) & (g437)) + ((!g2178) & (g2328) & (sk[118]) & (g437)) + ((g2178) & (!g2328) & (!sk[118]) & (g437)) + ((g2178) & (g2328) & (!sk[118]) & (!g437)) + ((g2178) & (g2328) & (!sk[118]) & (g437)) + ((g2178) & (g2328) & (sk[118]) & (!g437)) + ((g2178) & (g2328) & (sk[118]) & (g437)));
	assign g4201 = (((!g2179) & (!sk[119]) & (!g2328) & (g438)) + ((!g2179) & (!sk[119]) & (g2328) & (!g438)) + ((!g2179) & (!sk[119]) & (g2328) & (g438)) + ((!g2179) & (sk[119]) & (!g2328) & (g438)) + ((!g2179) & (sk[119]) & (g2328) & (g438)) + ((g2179) & (!sk[119]) & (!g2328) & (g438)) + ((g2179) & (!sk[119]) & (g2328) & (!g438)) + ((g2179) & (!sk[119]) & (g2328) & (g438)) + ((g2179) & (sk[119]) & (g2328) & (!g438)) + ((g2179) & (sk[119]) & (g2328) & (g438)));
	assign g439 = (((!g165) & (!g166) & (!sk[120]) & (!g436) & (g437) & (!g438)) + ((!g165) & (!g166) & (!sk[120]) & (!g436) & (g437) & (g438)) + ((!g165) & (!g166) & (!sk[120]) & (g436) & (!g437) & (!g438)) + ((!g165) & (!g166) & (!sk[120]) & (g436) & (!g437) & (g438)) + ((!g165) & (!g166) & (!sk[120]) & (g436) & (g437) & (!g438)) + ((!g165) & (!g166) & (!sk[120]) & (g436) & (g437) & (g438)) + ((!g165) & (g166) & (!sk[120]) & (!g436) & (!g437) & (!g438)) + ((!g165) & (g166) & (!sk[120]) & (!g436) & (!g437) & (g438)) + ((!g165) & (g166) & (!sk[120]) & (!g436) & (g437) & (!g438)) + ((!g165) & (g166) & (!sk[120]) & (!g436) & (g437) & (g438)) + ((!g165) & (g166) & (!sk[120]) & (g436) & (!g437) & (!g438)) + ((!g165) & (g166) & (!sk[120]) & (g436) & (!g437) & (g438)) + ((!g165) & (g166) & (!sk[120]) & (g436) & (g437) & (!g438)) + ((!g165) & (g166) & (!sk[120]) & (g436) & (g437) & (g438)) + ((!g165) & (g166) & (sk[120]) & (!g436) & (!g437) & (g438)) + ((!g165) & (g166) & (sk[120]) & (!g436) & (g437) & (g438)) + ((!g165) & (g166) & (sk[120]) & (g436) & (!g437) & (g438)) + ((!g165) & (g166) & (sk[120]) & (g436) & (g437) & (g438)) + ((g165) & (!g166) & (!sk[120]) & (!g436) & (g437) & (!g438)) + ((g165) & (!g166) & (!sk[120]) & (!g436) & (g437) & (g438)) + ((g165) & (!g166) & (!sk[120]) & (g436) & (!g437) & (!g438)) + ((g165) & (!g166) & (!sk[120]) & (g436) & (!g437) & (g438)) + ((g165) & (!g166) & (!sk[120]) & (g436) & (g437) & (!g438)) + ((g165) & (!g166) & (!sk[120]) & (g436) & (g437) & (g438)) + ((g165) & (!g166) & (sk[120]) & (g436) & (!g437) & (!g438)) + ((g165) & (!g166) & (sk[120]) & (g436) & (!g437) & (g438)) + ((g165) & (!g166) & (sk[120]) & (g436) & (g437) & (!g438)) + ((g165) & (!g166) & (sk[120]) & (g436) & (g437) & (g438)) + ((g165) & (g166) & (!sk[120]) & (!g436) & (!g437) & (!g438)) + ((g165) & (g166) & (!sk[120]) & (!g436) & (!g437) & (g438)) + ((g165) & (g166) & (!sk[120]) & (!g436) & (g437) & (!g438)) + ((g165) & (g166) & (!sk[120]) & (!g436) & (g437) & (g438)) + ((g165) & (g166) & (!sk[120]) & (g436) & (!g437) & (!g438)) + ((g165) & (g166) & (!sk[120]) & (g436) & (!g437) & (g438)) + ((g165) & (g166) & (!sk[120]) & (g436) & (g437) & (!g438)) + ((g165) & (g166) & (!sk[120]) & (g436) & (g437) & (g438)) + ((g165) & (g166) & (sk[120]) & (!g436) & (g437) & (!g438)) + ((g165) & (g166) & (sk[120]) & (!g436) & (g437) & (g438)) + ((g165) & (g166) & (sk[120]) & (g436) & (g437) & (!g438)) + ((g165) & (g166) & (sk[120]) & (g436) & (g437) & (g438)));
	assign g4202 = (((!g2162) & (!g2328) & (!sk[121]) & (g440)) + ((!g2162) & (!g2328) & (sk[121]) & (g440)) + ((!g2162) & (g2328) & (!sk[121]) & (!g440)) + ((!g2162) & (g2328) & (!sk[121]) & (g440)) + ((!g2162) & (g2328) & (sk[121]) & (g440)) + ((g2162) & (!g2328) & (!sk[121]) & (g440)) + ((g2162) & (g2328) & (!sk[121]) & (!g440)) + ((g2162) & (g2328) & (!sk[121]) & (g440)) + ((g2162) & (g2328) & (sk[121]) & (!g440)) + ((g2162) & (g2328) & (sk[121]) & (g440)));
	assign g4203 = (((!sk[122]) & (!g2164) & (!g2328) & (g441)) + ((!sk[122]) & (!g2164) & (g2328) & (!g441)) + ((!sk[122]) & (!g2164) & (g2328) & (g441)) + ((!sk[122]) & (g2164) & (!g2328) & (g441)) + ((!sk[122]) & (g2164) & (g2328) & (!g441)) + ((!sk[122]) & (g2164) & (g2328) & (g441)) + ((sk[122]) & (!g2164) & (!g2328) & (g441)) + ((sk[122]) & (!g2164) & (g2328) & (g441)) + ((sk[122]) & (g2164) & (g2328) & (!g441)) + ((sk[122]) & (g2164) & (g2328) & (g441)));
	assign g4204 = (((!g2166) & (!g2328) & (!sk[123]) & (g442)) + ((!g2166) & (!g2328) & (sk[123]) & (g442)) + ((!g2166) & (g2328) & (!sk[123]) & (!g442)) + ((!g2166) & (g2328) & (!sk[123]) & (g442)) + ((!g2166) & (g2328) & (sk[123]) & (g442)) + ((g2166) & (!g2328) & (!sk[123]) & (g442)) + ((g2166) & (g2328) & (!sk[123]) & (!g442)) + ((g2166) & (g2328) & (!sk[123]) & (g442)) + ((g2166) & (g2328) & (sk[123]) & (!g442)) + ((g2166) & (g2328) & (sk[123]) & (g442)));
	assign g4205 = (((!sk[124]) & (!g2168) & (!g2328) & (g443)) + ((!sk[124]) & (!g2168) & (g2328) & (!g443)) + ((!sk[124]) & (!g2168) & (g2328) & (g443)) + ((!sk[124]) & (g2168) & (!g2328) & (g443)) + ((!sk[124]) & (g2168) & (g2328) & (!g443)) + ((!sk[124]) & (g2168) & (g2328) & (g443)) + ((sk[124]) & (!g2168) & (!g2328) & (g443)) + ((sk[124]) & (!g2168) & (g2328) & (g443)) + ((sk[124]) & (g2168) & (g2328) & (!g443)) + ((sk[124]) & (g2168) & (g2328) & (g443)));
	assign g444 = (((!g440) & (!g441) & (!g442) & (g443) & (g165) & (g166)) + ((!g440) & (!g441) & (g442) & (!g443) & (!g165) & (g166)) + ((!g440) & (!g441) & (g442) & (g443) & (!g165) & (g166)) + ((!g440) & (!g441) & (g442) & (g443) & (g165) & (g166)) + ((!g440) & (g441) & (!g442) & (!g443) & (g165) & (!g166)) + ((!g440) & (g441) & (!g442) & (g443) & (g165) & (!g166)) + ((!g440) & (g441) & (!g442) & (g443) & (g165) & (g166)) + ((!g440) & (g441) & (g442) & (!g443) & (!g165) & (g166)) + ((!g440) & (g441) & (g442) & (!g443) & (g165) & (!g166)) + ((!g440) & (g441) & (g442) & (g443) & (!g165) & (g166)) + ((!g440) & (g441) & (g442) & (g443) & (g165) & (!g166)) + ((!g440) & (g441) & (g442) & (g443) & (g165) & (g166)) + ((g440) & (!g441) & (!g442) & (!g443) & (!g165) & (!g166)) + ((g440) & (!g441) & (!g442) & (g443) & (!g165) & (!g166)) + ((g440) & (!g441) & (!g442) & (g443) & (g165) & (g166)) + ((g440) & (!g441) & (g442) & (!g443) & (!g165) & (!g166)) + ((g440) & (!g441) & (g442) & (!g443) & (!g165) & (g166)) + ((g440) & (!g441) & (g442) & (g443) & (!g165) & (!g166)) + ((g440) & (!g441) & (g442) & (g443) & (!g165) & (g166)) + ((g440) & (!g441) & (g442) & (g443) & (g165) & (g166)) + ((g440) & (g441) & (!g442) & (!g443) & (!g165) & (!g166)) + ((g440) & (g441) & (!g442) & (!g443) & (g165) & (!g166)) + ((g440) & (g441) & (!g442) & (g443) & (!g165) & (!g166)) + ((g440) & (g441) & (!g442) & (g443) & (g165) & (!g166)) + ((g440) & (g441) & (!g442) & (g443) & (g165) & (g166)) + ((g440) & (g441) & (g442) & (!g443) & (!g165) & (!g166)) + ((g440) & (g441) & (g442) & (!g443) & (!g165) & (g166)) + ((g440) & (g441) & (g442) & (!g443) & (g165) & (!g166)) + ((g440) & (g441) & (g442) & (g443) & (!g165) & (!g166)) + ((g440) & (g441) & (g442) & (g443) & (!g165) & (g166)) + ((g440) & (g441) & (g442) & (g443) & (g165) & (!g166)) + ((g440) & (g441) & (g442) & (g443) & (g165) & (g166)));
	assign g4206 = (((!sk[126]) & (!g2169) & (!g2328) & (g445)) + ((!sk[126]) & (!g2169) & (g2328) & (!g445)) + ((!sk[126]) & (!g2169) & (g2328) & (g445)) + ((!sk[126]) & (g2169) & (!g2328) & (g445)) + ((!sk[126]) & (g2169) & (g2328) & (!g445)) + ((!sk[126]) & (g2169) & (g2328) & (g445)) + ((sk[126]) & (!g2169) & (!g2328) & (g445)) + ((sk[126]) & (!g2169) & (g2328) & (g445)) + ((sk[126]) & (g2169) & (g2328) & (!g445)) + ((sk[126]) & (g2169) & (g2328) & (g445)));
	assign g4207 = (((!g2170) & (!sk[127]) & (!g2328) & (g446)) + ((!g2170) & (!sk[127]) & (g2328) & (!g446)) + ((!g2170) & (!sk[127]) & (g2328) & (g446)) + ((!g2170) & (sk[127]) & (!g2328) & (g446)) + ((!g2170) & (sk[127]) & (g2328) & (g446)) + ((g2170) & (!sk[127]) & (!g2328) & (g446)) + ((g2170) & (!sk[127]) & (g2328) & (!g446)) + ((g2170) & (!sk[127]) & (g2328) & (g446)) + ((g2170) & (sk[127]) & (g2328) & (!g446)) + ((g2170) & (sk[127]) & (g2328) & (g446)));
	assign g4208 = (((!g2171) & (!g2328) & (!sk[0]) & (g447)) + ((!g2171) & (!g2328) & (sk[0]) & (g447)) + ((!g2171) & (g2328) & (!sk[0]) & (!g447)) + ((!g2171) & (g2328) & (!sk[0]) & (g447)) + ((!g2171) & (g2328) & (sk[0]) & (g447)) + ((g2171) & (!g2328) & (!sk[0]) & (g447)) + ((g2171) & (g2328) & (!sk[0]) & (!g447)) + ((g2171) & (g2328) & (!sk[0]) & (g447)) + ((g2171) & (g2328) & (sk[0]) & (!g447)) + ((g2171) & (g2328) & (sk[0]) & (g447)));
	assign g4209 = (((!g2172) & (!sk[1]) & (!g2328) & (g448)) + ((!g2172) & (!sk[1]) & (g2328) & (!g448)) + ((!g2172) & (!sk[1]) & (g2328) & (g448)) + ((!g2172) & (sk[1]) & (!g2328) & (g448)) + ((!g2172) & (sk[1]) & (g2328) & (g448)) + ((g2172) & (!sk[1]) & (!g2328) & (g448)) + ((g2172) & (!sk[1]) & (g2328) & (!g448)) + ((g2172) & (!sk[1]) & (g2328) & (g448)) + ((g2172) & (sk[1]) & (g2328) & (!g448)) + ((g2172) & (sk[1]) & (g2328) & (g448)));
	assign g449 = (((!g445) & (!g446) & (!g447) & (g448) & (g165) & (g166)) + ((!g445) & (!g446) & (g447) & (!g448) & (!g165) & (g166)) + ((!g445) & (!g446) & (g447) & (g448) & (!g165) & (g166)) + ((!g445) & (!g446) & (g447) & (g448) & (g165) & (g166)) + ((!g445) & (g446) & (!g447) & (!g448) & (g165) & (!g166)) + ((!g445) & (g446) & (!g447) & (g448) & (g165) & (!g166)) + ((!g445) & (g446) & (!g447) & (g448) & (g165) & (g166)) + ((!g445) & (g446) & (g447) & (!g448) & (!g165) & (g166)) + ((!g445) & (g446) & (g447) & (!g448) & (g165) & (!g166)) + ((!g445) & (g446) & (g447) & (g448) & (!g165) & (g166)) + ((!g445) & (g446) & (g447) & (g448) & (g165) & (!g166)) + ((!g445) & (g446) & (g447) & (g448) & (g165) & (g166)) + ((g445) & (!g446) & (!g447) & (!g448) & (!g165) & (!g166)) + ((g445) & (!g446) & (!g447) & (g448) & (!g165) & (!g166)) + ((g445) & (!g446) & (!g447) & (g448) & (g165) & (g166)) + ((g445) & (!g446) & (g447) & (!g448) & (!g165) & (!g166)) + ((g445) & (!g446) & (g447) & (!g448) & (!g165) & (g166)) + ((g445) & (!g446) & (g447) & (g448) & (!g165) & (!g166)) + ((g445) & (!g446) & (g447) & (g448) & (!g165) & (g166)) + ((g445) & (!g446) & (g447) & (g448) & (g165) & (g166)) + ((g445) & (g446) & (!g447) & (!g448) & (!g165) & (!g166)) + ((g445) & (g446) & (!g447) & (!g448) & (g165) & (!g166)) + ((g445) & (g446) & (!g447) & (g448) & (!g165) & (!g166)) + ((g445) & (g446) & (!g447) & (g448) & (g165) & (!g166)) + ((g445) & (g446) & (!g447) & (g448) & (g165) & (g166)) + ((g445) & (g446) & (g447) & (!g448) & (!g165) & (!g166)) + ((g445) & (g446) & (g447) & (!g448) & (!g165) & (g166)) + ((g445) & (g446) & (g447) & (!g448) & (g165) & (!g166)) + ((g445) & (g446) & (g447) & (g448) & (!g165) & (!g166)) + ((g445) & (g446) & (g447) & (g448) & (!g165) & (g166)) + ((g445) & (g446) & (g447) & (g448) & (g165) & (!g166)) + ((g445) & (g446) & (g447) & (g448) & (g165) & (g166)));
	assign g450 = (((!g147) & (!g148) & (!g435) & (g439) & (!g444) & (!g449)) + ((!g147) & (!g148) & (!g435) & (g439) & (!g444) & (g449)) + ((!g147) & (!g148) & (!g435) & (g439) & (g444) & (!g449)) + ((!g147) & (!g148) & (!g435) & (g439) & (g444) & (g449)) + ((!g147) & (!g148) & (g435) & (g439) & (!g444) & (!g449)) + ((!g147) & (!g148) & (g435) & (g439) & (!g444) & (g449)) + ((!g147) & (!g148) & (g435) & (g439) & (g444) & (!g449)) + ((!g147) & (!g148) & (g435) & (g439) & (g444) & (g449)) + ((!g147) & (g148) & (!g435) & (!g439) & (!g444) & (g449)) + ((!g147) & (g148) & (!g435) & (!g439) & (g444) & (g449)) + ((!g147) & (g148) & (!g435) & (g439) & (!g444) & (g449)) + ((!g147) & (g148) & (!g435) & (g439) & (g444) & (g449)) + ((!g147) & (g148) & (g435) & (!g439) & (!g444) & (g449)) + ((!g147) & (g148) & (g435) & (!g439) & (g444) & (g449)) + ((!g147) & (g148) & (g435) & (g439) & (!g444) & (g449)) + ((!g147) & (g148) & (g435) & (g439) & (g444) & (g449)) + ((g147) & (!g148) & (g435) & (!g439) & (!g444) & (!g449)) + ((g147) & (!g148) & (g435) & (!g439) & (!g444) & (g449)) + ((g147) & (!g148) & (g435) & (!g439) & (g444) & (!g449)) + ((g147) & (!g148) & (g435) & (!g439) & (g444) & (g449)) + ((g147) & (!g148) & (g435) & (g439) & (!g444) & (!g449)) + ((g147) & (!g148) & (g435) & (g439) & (!g444) & (g449)) + ((g147) & (!g148) & (g435) & (g439) & (g444) & (!g449)) + ((g147) & (!g148) & (g435) & (g439) & (g444) & (g449)) + ((g147) & (g148) & (!g435) & (!g439) & (g444) & (!g449)) + ((g147) & (g148) & (!g435) & (!g439) & (g444) & (g449)) + ((g147) & (g148) & (!g435) & (g439) & (g444) & (!g449)) + ((g147) & (g148) & (!g435) & (g439) & (g444) & (g449)) + ((g147) & (g148) & (g435) & (!g439) & (g444) & (!g449)) + ((g147) & (g148) & (g435) & (!g439) & (g444) & (g449)) + ((g147) & (g148) & (g435) & (g439) & (g444) & (!g449)) + ((g147) & (g148) & (g435) & (g439) & (g444) & (g449)));
	assign g451 = (((!sk[4]) & (!g142) & (!g430) & (g450)) + ((!sk[4]) & (!g142) & (g430) & (!g450)) + ((!sk[4]) & (!g142) & (g430) & (g450)) + ((!sk[4]) & (g142) & (!g430) & (g450)) + ((!sk[4]) & (g142) & (g430) & (!g450)) + ((!sk[4]) & (g142) & (g430) & (g450)) + ((sk[4]) & (!g142) & (!g430) & (g450)) + ((sk[4]) & (!g142) & (g430) & (g450)) + ((sk[4]) & (g142) & (g430) & (!g450)) + ((sk[4]) & (g142) & (g430) & (g450)));
	assign g452 = (((!sk[5]) & (!g86) & (!g126) & (!g408) & (g409) & (!g451)) + ((!sk[5]) & (!g86) & (!g126) & (!g408) & (g409) & (g451)) + ((!sk[5]) & (!g86) & (!g126) & (g408) & (!g409) & (!g451)) + ((!sk[5]) & (!g86) & (!g126) & (g408) & (!g409) & (g451)) + ((!sk[5]) & (!g86) & (!g126) & (g408) & (g409) & (!g451)) + ((!sk[5]) & (!g86) & (!g126) & (g408) & (g409) & (g451)) + ((!sk[5]) & (!g86) & (g126) & (!g408) & (!g409) & (!g451)) + ((!sk[5]) & (!g86) & (g126) & (!g408) & (!g409) & (g451)) + ((!sk[5]) & (!g86) & (g126) & (!g408) & (g409) & (!g451)) + ((!sk[5]) & (!g86) & (g126) & (!g408) & (g409) & (g451)) + ((!sk[5]) & (!g86) & (g126) & (g408) & (!g409) & (!g451)) + ((!sk[5]) & (!g86) & (g126) & (g408) & (!g409) & (g451)) + ((!sk[5]) & (!g86) & (g126) & (g408) & (g409) & (!g451)) + ((!sk[5]) & (!g86) & (g126) & (g408) & (g409) & (g451)) + ((!sk[5]) & (g86) & (!g126) & (!g408) & (g409) & (!g451)) + ((!sk[5]) & (g86) & (!g126) & (!g408) & (g409) & (g451)) + ((!sk[5]) & (g86) & (!g126) & (g408) & (!g409) & (!g451)) + ((!sk[5]) & (g86) & (!g126) & (g408) & (!g409) & (g451)) + ((!sk[5]) & (g86) & (!g126) & (g408) & (g409) & (!g451)) + ((!sk[5]) & (g86) & (!g126) & (g408) & (g409) & (g451)) + ((!sk[5]) & (g86) & (g126) & (!g408) & (!g409) & (!g451)) + ((!sk[5]) & (g86) & (g126) & (!g408) & (!g409) & (g451)) + ((!sk[5]) & (g86) & (g126) & (!g408) & (g409) & (!g451)) + ((!sk[5]) & (g86) & (g126) & (!g408) & (g409) & (g451)) + ((!sk[5]) & (g86) & (g126) & (g408) & (!g409) & (!g451)) + ((!sk[5]) & (g86) & (g126) & (g408) & (!g409) & (g451)) + ((!sk[5]) & (g86) & (g126) & (g408) & (g409) & (!g451)) + ((!sk[5]) & (g86) & (g126) & (g408) & (g409) & (g451)) + ((sk[5]) & (!g86) & (!g126) & (g408) & (!g409) & (!g451)) + ((sk[5]) & (!g86) & (!g126) & (g408) & (!g409) & (g451)) + ((sk[5]) & (!g86) & (!g126) & (g408) & (g409) & (!g451)) + ((sk[5]) & (!g86) & (!g126) & (g408) & (g409) & (g451)) + ((sk[5]) & (!g86) & (g126) & (!g408) & (!g409) & (g451)) + ((sk[5]) & (!g86) & (g126) & (!g408) & (g409) & (!g451)) + ((sk[5]) & (!g86) & (g126) & (g408) & (!g409) & (g451)) + ((sk[5]) & (!g86) & (g126) & (g408) & (g409) & (!g451)) + ((sk[5]) & (g86) & (!g126) & (g408) & (!g409) & (!g451)) + ((sk[5]) & (g86) & (!g126) & (g408) & (!g409) & (g451)) + ((sk[5]) & (g86) & (!g126) & (g408) & (g409) & (!g451)) + ((sk[5]) & (g86) & (!g126) & (g408) & (g409) & (g451)) + ((sk[5]) & (g86) & (g126) & (!g408) & (!g409) & (!g451)) + ((sk[5]) & (g86) & (g126) & (!g408) & (g409) & (g451)) + ((sk[5]) & (g86) & (g126) & (g408) & (!g409) & (!g451)) + ((sk[5]) & (g86) & (g126) & (g408) & (g409) & (g451)));
	assign g4210 = (((!sk[6]) & (!g2059) & (!g2337) & (g453)) + ((!sk[6]) & (!g2059) & (g2337) & (!g453)) + ((!sk[6]) & (!g2059) & (g2337) & (g453)) + ((!sk[6]) & (g2059) & (!g2337) & (g453)) + ((!sk[6]) & (g2059) & (g2337) & (!g453)) + ((!sk[6]) & (g2059) & (g2337) & (g453)) + ((sk[6]) & (!g2059) & (!g2337) & (g453)) + ((sk[6]) & (!g2059) & (g2337) & (g453)) + ((sk[6]) & (g2059) & (g2337) & (!g453)) + ((sk[6]) & (g2059) & (g2337) & (g453)));
	assign g4211 = (((!g2140) & (!sk[7]) & (!g3676) & (g454)) + ((!g2140) & (!sk[7]) & (g3676) & (!g454)) + ((!g2140) & (!sk[7]) & (g3676) & (g454)) + ((!g2140) & (sk[7]) & (!g3676) & (g454)) + ((!g2140) & (sk[7]) & (g3676) & (g454)) + ((g2140) & (!sk[7]) & (!g3676) & (g454)) + ((g2140) & (!sk[7]) & (g3676) & (!g454)) + ((g2140) & (!sk[7]) & (g3676) & (g454)) + ((g2140) & (sk[7]) & (g3676) & (!g454)) + ((g2140) & (sk[7]) & (g3676) & (g454)));
	assign g4212 = (((!sk[8]) & (!g2146) & (!g3676) & (g455)) + ((!sk[8]) & (!g2146) & (g3676) & (!g455)) + ((!sk[8]) & (!g2146) & (g3676) & (g455)) + ((!sk[8]) & (g2146) & (!g3676) & (g455)) + ((!sk[8]) & (g2146) & (g3676) & (!g455)) + ((!sk[8]) & (g2146) & (g3676) & (g455)) + ((sk[8]) & (!g2146) & (!g3676) & (g455)) + ((sk[8]) & (!g2146) & (g3676) & (g455)) + ((sk[8]) & (g2146) & (g3676) & (!g455)) + ((sk[8]) & (g2146) & (g3676) & (g455)));
	assign g4213 = (((!g2152) & (!sk[9]) & (!g3676) & (g456)) + ((!g2152) & (!sk[9]) & (g3676) & (!g456)) + ((!g2152) & (!sk[9]) & (g3676) & (g456)) + ((!g2152) & (sk[9]) & (!g3676) & (g456)) + ((!g2152) & (sk[9]) & (g3676) & (g456)) + ((g2152) & (!sk[9]) & (!g3676) & (g456)) + ((g2152) & (!sk[9]) & (g3676) & (!g456)) + ((g2152) & (!sk[9]) & (g3676) & (g456)) + ((g2152) & (sk[9]) & (g3676) & (!g456)) + ((g2152) & (sk[9]) & (g3676) & (g456)));
	assign g4214 = (((!sk[10]) & (!g2158) & (!g3676) & (g457)) + ((!sk[10]) & (!g2158) & (g3676) & (!g457)) + ((!sk[10]) & (!g2158) & (g3676) & (g457)) + ((!sk[10]) & (g2158) & (!g3676) & (g457)) + ((!sk[10]) & (g2158) & (g3676) & (!g457)) + ((!sk[10]) & (g2158) & (g3676) & (g457)) + ((sk[10]) & (!g2158) & (!g3676) & (g457)) + ((sk[10]) & (!g2158) & (g3676) & (g457)) + ((sk[10]) & (g2158) & (g3676) & (!g457)) + ((sk[10]) & (g2158) & (g3676) & (g457)));
	assign g458 = (((!g454) & (!g455) & (!g456) & (g457) & (g165) & (g166)) + ((!g454) & (!g455) & (g456) & (!g457) & (!g165) & (g166)) + ((!g454) & (!g455) & (g456) & (g457) & (!g165) & (g166)) + ((!g454) & (!g455) & (g456) & (g457) & (g165) & (g166)) + ((!g454) & (g455) & (!g456) & (!g457) & (g165) & (!g166)) + ((!g454) & (g455) & (!g456) & (g457) & (g165) & (!g166)) + ((!g454) & (g455) & (!g456) & (g457) & (g165) & (g166)) + ((!g454) & (g455) & (g456) & (!g457) & (!g165) & (g166)) + ((!g454) & (g455) & (g456) & (!g457) & (g165) & (!g166)) + ((!g454) & (g455) & (g456) & (g457) & (!g165) & (g166)) + ((!g454) & (g455) & (g456) & (g457) & (g165) & (!g166)) + ((!g454) & (g455) & (g456) & (g457) & (g165) & (g166)) + ((g454) & (!g455) & (!g456) & (!g457) & (!g165) & (!g166)) + ((g454) & (!g455) & (!g456) & (g457) & (!g165) & (!g166)) + ((g454) & (!g455) & (!g456) & (g457) & (g165) & (g166)) + ((g454) & (!g455) & (g456) & (!g457) & (!g165) & (!g166)) + ((g454) & (!g455) & (g456) & (!g457) & (!g165) & (g166)) + ((g454) & (!g455) & (g456) & (g457) & (!g165) & (!g166)) + ((g454) & (!g455) & (g456) & (g457) & (!g165) & (g166)) + ((g454) & (!g455) & (g456) & (g457) & (g165) & (g166)) + ((g454) & (g455) & (!g456) & (!g457) & (!g165) & (!g166)) + ((g454) & (g455) & (!g456) & (!g457) & (g165) & (!g166)) + ((g454) & (g455) & (!g456) & (g457) & (!g165) & (!g166)) + ((g454) & (g455) & (!g456) & (g457) & (g165) & (!g166)) + ((g454) & (g455) & (!g456) & (g457) & (g165) & (g166)) + ((g454) & (g455) & (g456) & (!g457) & (!g165) & (!g166)) + ((g454) & (g455) & (g456) & (!g457) & (!g165) & (g166)) + ((g454) & (g455) & (g456) & (!g457) & (g165) & (!g166)) + ((g454) & (g455) & (g456) & (g457) & (!g165) & (!g166)) + ((g454) & (g455) & (g456) & (g457) & (!g165) & (g166)) + ((g454) & (g455) & (g456) & (g457) & (g165) & (!g166)) + ((g454) & (g455) & (g456) & (g457) & (g165) & (g166)));
	assign g4215 = (((!g2142) & (!sk[12]) & (!g3676) & (g459)) + ((!g2142) & (!sk[12]) & (g3676) & (!g459)) + ((!g2142) & (!sk[12]) & (g3676) & (g459)) + ((!g2142) & (sk[12]) & (!g3676) & (g459)) + ((!g2142) & (sk[12]) & (g3676) & (g459)) + ((g2142) & (!sk[12]) & (!g3676) & (g459)) + ((g2142) & (!sk[12]) & (g3676) & (!g459)) + ((g2142) & (!sk[12]) & (g3676) & (g459)) + ((g2142) & (sk[12]) & (g3676) & (!g459)) + ((g2142) & (sk[12]) & (g3676) & (g459)));
	assign g4216 = (((!g2148) & (!g3676) & (!sk[13]) & (g460)) + ((!g2148) & (!g3676) & (sk[13]) & (g460)) + ((!g2148) & (g3676) & (!sk[13]) & (!g460)) + ((!g2148) & (g3676) & (!sk[13]) & (g460)) + ((!g2148) & (g3676) & (sk[13]) & (g460)) + ((g2148) & (!g3676) & (!sk[13]) & (g460)) + ((g2148) & (g3676) & (!sk[13]) & (!g460)) + ((g2148) & (g3676) & (!sk[13]) & (g460)) + ((g2148) & (g3676) & (sk[13]) & (!g460)) + ((g2148) & (g3676) & (sk[13]) & (g460)));
	assign g4217 = (((!sk[14]) & (!g2153) & (!g3676) & (g461)) + ((!sk[14]) & (!g2153) & (g3676) & (!g461)) + ((!sk[14]) & (!g2153) & (g3676) & (g461)) + ((!sk[14]) & (g2153) & (!g3676) & (g461)) + ((!sk[14]) & (g2153) & (g3676) & (!g461)) + ((!sk[14]) & (g2153) & (g3676) & (g461)) + ((sk[14]) & (!g2153) & (!g3676) & (g461)) + ((sk[14]) & (!g2153) & (g3676) & (g461)) + ((sk[14]) & (g2153) & (g3676) & (!g461)) + ((sk[14]) & (g2153) & (g3676) & (g461)));
	assign g4218 = (((!g2159) & (!sk[15]) & (!g3676) & (g462)) + ((!g2159) & (!sk[15]) & (g3676) & (!g462)) + ((!g2159) & (!sk[15]) & (g3676) & (g462)) + ((!g2159) & (sk[15]) & (!g3676) & (g462)) + ((!g2159) & (sk[15]) & (g3676) & (g462)) + ((g2159) & (!sk[15]) & (!g3676) & (g462)) + ((g2159) & (!sk[15]) & (g3676) & (!g462)) + ((g2159) & (!sk[15]) & (g3676) & (g462)) + ((g2159) & (sk[15]) & (g3676) & (!g462)) + ((g2159) & (sk[15]) & (g3676) & (g462)));
	assign g463 = (((!g459) & (!g460) & (!g461) & (g462) & (g165) & (g166)) + ((!g459) & (!g460) & (g461) & (!g462) & (!g165) & (g166)) + ((!g459) & (!g460) & (g461) & (g462) & (!g165) & (g166)) + ((!g459) & (!g460) & (g461) & (g462) & (g165) & (g166)) + ((!g459) & (g460) & (!g461) & (!g462) & (g165) & (!g166)) + ((!g459) & (g460) & (!g461) & (g462) & (g165) & (!g166)) + ((!g459) & (g460) & (!g461) & (g462) & (g165) & (g166)) + ((!g459) & (g460) & (g461) & (!g462) & (!g165) & (g166)) + ((!g459) & (g460) & (g461) & (!g462) & (g165) & (!g166)) + ((!g459) & (g460) & (g461) & (g462) & (!g165) & (g166)) + ((!g459) & (g460) & (g461) & (g462) & (g165) & (!g166)) + ((!g459) & (g460) & (g461) & (g462) & (g165) & (g166)) + ((g459) & (!g460) & (!g461) & (!g462) & (!g165) & (!g166)) + ((g459) & (!g460) & (!g461) & (g462) & (!g165) & (!g166)) + ((g459) & (!g460) & (!g461) & (g462) & (g165) & (g166)) + ((g459) & (!g460) & (g461) & (!g462) & (!g165) & (!g166)) + ((g459) & (!g460) & (g461) & (!g462) & (!g165) & (g166)) + ((g459) & (!g460) & (g461) & (g462) & (!g165) & (!g166)) + ((g459) & (!g460) & (g461) & (g462) & (!g165) & (g166)) + ((g459) & (!g460) & (g461) & (g462) & (g165) & (g166)) + ((g459) & (g460) & (!g461) & (!g462) & (!g165) & (!g166)) + ((g459) & (g460) & (!g461) & (!g462) & (g165) & (!g166)) + ((g459) & (g460) & (!g461) & (g462) & (!g165) & (!g166)) + ((g459) & (g460) & (!g461) & (g462) & (g165) & (!g166)) + ((g459) & (g460) & (!g461) & (g462) & (g165) & (g166)) + ((g459) & (g460) & (g461) & (!g462) & (!g165) & (!g166)) + ((g459) & (g460) & (g461) & (!g462) & (!g165) & (g166)) + ((g459) & (g460) & (g461) & (!g462) & (g165) & (!g166)) + ((g459) & (g460) & (g461) & (g462) & (!g165) & (!g166)) + ((g459) & (g460) & (g461) & (g462) & (!g165) & (g166)) + ((g459) & (g460) & (g461) & (g462) & (g165) & (!g166)) + ((g459) & (g460) & (g461) & (g462) & (g165) & (g166)));
	assign g4219 = (((!g2144) & (!sk[17]) & (!g3676) & (g464)) + ((!g2144) & (!sk[17]) & (g3676) & (!g464)) + ((!g2144) & (!sk[17]) & (g3676) & (g464)) + ((!g2144) & (sk[17]) & (!g3676) & (g464)) + ((!g2144) & (sk[17]) & (g3676) & (g464)) + ((g2144) & (!sk[17]) & (!g3676) & (g464)) + ((g2144) & (!sk[17]) & (g3676) & (!g464)) + ((g2144) & (!sk[17]) & (g3676) & (g464)) + ((g2144) & (sk[17]) & (g3676) & (!g464)) + ((g2144) & (sk[17]) & (g3676) & (g464)));
	assign g4220 = (((!g2150) & (!sk[18]) & (!g3676) & (g465)) + ((!g2150) & (!sk[18]) & (g3676) & (!g465)) + ((!g2150) & (!sk[18]) & (g3676) & (g465)) + ((!g2150) & (sk[18]) & (!g3676) & (g465)) + ((!g2150) & (sk[18]) & (g3676) & (g465)) + ((g2150) & (!sk[18]) & (!g3676) & (g465)) + ((g2150) & (!sk[18]) & (g3676) & (!g465)) + ((g2150) & (!sk[18]) & (g3676) & (g465)) + ((g2150) & (sk[18]) & (g3676) & (!g465)) + ((g2150) & (sk[18]) & (g3676) & (g465)));
	assign g4221 = (((!g2155) & (!g3676) & (!sk[19]) & (g466)) + ((!g2155) & (!g3676) & (sk[19]) & (g466)) + ((!g2155) & (g3676) & (!sk[19]) & (!g466)) + ((!g2155) & (g3676) & (!sk[19]) & (g466)) + ((!g2155) & (g3676) & (sk[19]) & (g466)) + ((g2155) & (!g3676) & (!sk[19]) & (g466)) + ((g2155) & (g3676) & (!sk[19]) & (!g466)) + ((g2155) & (g3676) & (!sk[19]) & (g466)) + ((g2155) & (g3676) & (sk[19]) & (!g466)) + ((g2155) & (g3676) & (sk[19]) & (g466)));
	assign g4222 = (((!g2160) & (!sk[20]) & (!g3676) & (g467)) + ((!g2160) & (!sk[20]) & (g3676) & (!g467)) + ((!g2160) & (!sk[20]) & (g3676) & (g467)) + ((!g2160) & (sk[20]) & (!g3676) & (g467)) + ((!g2160) & (sk[20]) & (g3676) & (g467)) + ((g2160) & (!sk[20]) & (!g3676) & (g467)) + ((g2160) & (!sk[20]) & (g3676) & (!g467)) + ((g2160) & (!sk[20]) & (g3676) & (g467)) + ((g2160) & (sk[20]) & (g3676) & (!g467)) + ((g2160) & (sk[20]) & (g3676) & (g467)));
	assign g468 = (((!g464) & (!g465) & (!g466) & (g467) & (g165) & (g166)) + ((!g464) & (!g465) & (g466) & (!g467) & (!g165) & (g166)) + ((!g464) & (!g465) & (g466) & (g467) & (!g165) & (g166)) + ((!g464) & (!g465) & (g466) & (g467) & (g165) & (g166)) + ((!g464) & (g465) & (!g466) & (!g467) & (g165) & (!g166)) + ((!g464) & (g465) & (!g466) & (g467) & (g165) & (!g166)) + ((!g464) & (g465) & (!g466) & (g467) & (g165) & (g166)) + ((!g464) & (g465) & (g466) & (!g467) & (!g165) & (g166)) + ((!g464) & (g465) & (g466) & (!g467) & (g165) & (!g166)) + ((!g464) & (g465) & (g466) & (g467) & (!g165) & (g166)) + ((!g464) & (g465) & (g466) & (g467) & (g165) & (!g166)) + ((!g464) & (g465) & (g466) & (g467) & (g165) & (g166)) + ((g464) & (!g465) & (!g466) & (!g467) & (!g165) & (!g166)) + ((g464) & (!g465) & (!g466) & (g467) & (!g165) & (!g166)) + ((g464) & (!g465) & (!g466) & (g467) & (g165) & (g166)) + ((g464) & (!g465) & (g466) & (!g467) & (!g165) & (!g166)) + ((g464) & (!g465) & (g466) & (!g467) & (!g165) & (g166)) + ((g464) & (!g465) & (g466) & (g467) & (!g165) & (!g166)) + ((g464) & (!g465) & (g466) & (g467) & (!g165) & (g166)) + ((g464) & (!g465) & (g466) & (g467) & (g165) & (g166)) + ((g464) & (g465) & (!g466) & (!g467) & (!g165) & (!g166)) + ((g464) & (g465) & (!g466) & (!g467) & (g165) & (!g166)) + ((g464) & (g465) & (!g466) & (g467) & (!g165) & (!g166)) + ((g464) & (g465) & (!g466) & (g467) & (g165) & (!g166)) + ((g464) & (g465) & (!g466) & (g467) & (g165) & (g166)) + ((g464) & (g465) & (g466) & (!g467) & (!g165) & (!g166)) + ((g464) & (g465) & (g466) & (!g467) & (!g165) & (g166)) + ((g464) & (g465) & (g466) & (!g467) & (g165) & (!g166)) + ((g464) & (g465) & (g466) & (g467) & (!g165) & (!g166)) + ((g464) & (g465) & (g466) & (g467) & (!g165) & (g166)) + ((g464) & (g465) & (g466) & (g467) & (g165) & (!g166)) + ((g464) & (g465) & (g466) & (g467) & (g165) & (g166)));
	assign g4223 = (((!g2145) & (!g3676) & (!sk[22]) & (g469)) + ((!g2145) & (!g3676) & (sk[22]) & (g469)) + ((!g2145) & (g3676) & (!sk[22]) & (!g469)) + ((!g2145) & (g3676) & (!sk[22]) & (g469)) + ((!g2145) & (g3676) & (sk[22]) & (g469)) + ((g2145) & (!g3676) & (!sk[22]) & (g469)) + ((g2145) & (g3676) & (!sk[22]) & (!g469)) + ((g2145) & (g3676) & (!sk[22]) & (g469)) + ((g2145) & (g3676) & (sk[22]) & (!g469)) + ((g2145) & (g3676) & (sk[22]) & (g469)));
	assign g4224 = (((!sk[23]) & (!g2151) & (!g3676) & (g470)) + ((!sk[23]) & (!g2151) & (g3676) & (!g470)) + ((!sk[23]) & (!g2151) & (g3676) & (g470)) + ((!sk[23]) & (g2151) & (!g3676) & (g470)) + ((!sk[23]) & (g2151) & (g3676) & (!g470)) + ((!sk[23]) & (g2151) & (g3676) & (g470)) + ((sk[23]) & (!g2151) & (!g3676) & (g470)) + ((sk[23]) & (!g2151) & (g3676) & (g470)) + ((sk[23]) & (g2151) & (g3676) & (!g470)) + ((sk[23]) & (g2151) & (g3676) & (g470)));
	assign g4225 = (((!g2157) & (!g3676) & (!sk[24]) & (g471)) + ((!g2157) & (!g3676) & (sk[24]) & (g471)) + ((!g2157) & (g3676) & (!sk[24]) & (!g471)) + ((!g2157) & (g3676) & (!sk[24]) & (g471)) + ((!g2157) & (g3676) & (sk[24]) & (g471)) + ((g2157) & (!g3676) & (!sk[24]) & (g471)) + ((g2157) & (g3676) & (!sk[24]) & (!g471)) + ((g2157) & (g3676) & (!sk[24]) & (g471)) + ((g2157) & (g3676) & (sk[24]) & (!g471)) + ((g2157) & (g3676) & (sk[24]) & (g471)));
	assign g4226 = (((!g2161) & (!sk[25]) & (!g3676) & (g472)) + ((!g2161) & (!sk[25]) & (g3676) & (!g472)) + ((!g2161) & (!sk[25]) & (g3676) & (g472)) + ((!g2161) & (sk[25]) & (!g3676) & (g472)) + ((!g2161) & (sk[25]) & (g3676) & (g472)) + ((g2161) & (!sk[25]) & (!g3676) & (g472)) + ((g2161) & (!sk[25]) & (g3676) & (!g472)) + ((g2161) & (!sk[25]) & (g3676) & (g472)) + ((g2161) & (sk[25]) & (g3676) & (!g472)) + ((g2161) & (sk[25]) & (g3676) & (g472)));
	assign g473 = (((!g469) & (!g470) & (!g471) & (g472) & (g165) & (g166)) + ((!g469) & (!g470) & (g471) & (!g472) & (!g165) & (g166)) + ((!g469) & (!g470) & (g471) & (g472) & (!g165) & (g166)) + ((!g469) & (!g470) & (g471) & (g472) & (g165) & (g166)) + ((!g469) & (g470) & (!g471) & (!g472) & (g165) & (!g166)) + ((!g469) & (g470) & (!g471) & (g472) & (g165) & (!g166)) + ((!g469) & (g470) & (!g471) & (g472) & (g165) & (g166)) + ((!g469) & (g470) & (g471) & (!g472) & (!g165) & (g166)) + ((!g469) & (g470) & (g471) & (!g472) & (g165) & (!g166)) + ((!g469) & (g470) & (g471) & (g472) & (!g165) & (g166)) + ((!g469) & (g470) & (g471) & (g472) & (g165) & (!g166)) + ((!g469) & (g470) & (g471) & (g472) & (g165) & (g166)) + ((g469) & (!g470) & (!g471) & (!g472) & (!g165) & (!g166)) + ((g469) & (!g470) & (!g471) & (g472) & (!g165) & (!g166)) + ((g469) & (!g470) & (!g471) & (g472) & (g165) & (g166)) + ((g469) & (!g470) & (g471) & (!g472) & (!g165) & (!g166)) + ((g469) & (!g470) & (g471) & (!g472) & (!g165) & (g166)) + ((g469) & (!g470) & (g471) & (g472) & (!g165) & (!g166)) + ((g469) & (!g470) & (g471) & (g472) & (!g165) & (g166)) + ((g469) & (!g470) & (g471) & (g472) & (g165) & (g166)) + ((g469) & (g470) & (!g471) & (!g472) & (!g165) & (!g166)) + ((g469) & (g470) & (!g471) & (!g472) & (g165) & (!g166)) + ((g469) & (g470) & (!g471) & (g472) & (!g165) & (!g166)) + ((g469) & (g470) & (!g471) & (g472) & (g165) & (!g166)) + ((g469) & (g470) & (!g471) & (g472) & (g165) & (g166)) + ((g469) & (g470) & (g471) & (!g472) & (!g165) & (!g166)) + ((g469) & (g470) & (g471) & (!g472) & (!g165) & (g166)) + ((g469) & (g470) & (g471) & (!g472) & (g165) & (!g166)) + ((g469) & (g470) & (g471) & (g472) & (!g165) & (!g166)) + ((g469) & (g470) & (g471) & (g472) & (!g165) & (g166)) + ((g469) & (g470) & (g471) & (g472) & (g165) & (!g166)) + ((g469) & (g470) & (g471) & (g472) & (g165) & (g166)));
	assign g474 = (((!g458) & (!g463) & (!g468) & (g473) & (g147) & (g148)) + ((!g458) & (!g463) & (g468) & (!g473) & (!g147) & (g148)) + ((!g458) & (!g463) & (g468) & (g473) & (!g147) & (g148)) + ((!g458) & (!g463) & (g468) & (g473) & (g147) & (g148)) + ((!g458) & (g463) & (!g468) & (!g473) & (g147) & (!g148)) + ((!g458) & (g463) & (!g468) & (g473) & (g147) & (!g148)) + ((!g458) & (g463) & (!g468) & (g473) & (g147) & (g148)) + ((!g458) & (g463) & (g468) & (!g473) & (!g147) & (g148)) + ((!g458) & (g463) & (g468) & (!g473) & (g147) & (!g148)) + ((!g458) & (g463) & (g468) & (g473) & (!g147) & (g148)) + ((!g458) & (g463) & (g468) & (g473) & (g147) & (!g148)) + ((!g458) & (g463) & (g468) & (g473) & (g147) & (g148)) + ((g458) & (!g463) & (!g468) & (!g473) & (!g147) & (!g148)) + ((g458) & (!g463) & (!g468) & (g473) & (!g147) & (!g148)) + ((g458) & (!g463) & (!g468) & (g473) & (g147) & (g148)) + ((g458) & (!g463) & (g468) & (!g473) & (!g147) & (!g148)) + ((g458) & (!g463) & (g468) & (!g473) & (!g147) & (g148)) + ((g458) & (!g463) & (g468) & (g473) & (!g147) & (!g148)) + ((g458) & (!g463) & (g468) & (g473) & (!g147) & (g148)) + ((g458) & (!g463) & (g468) & (g473) & (g147) & (g148)) + ((g458) & (g463) & (!g468) & (!g473) & (!g147) & (!g148)) + ((g458) & (g463) & (!g468) & (!g473) & (g147) & (!g148)) + ((g458) & (g463) & (!g468) & (g473) & (!g147) & (!g148)) + ((g458) & (g463) & (!g468) & (g473) & (g147) & (!g148)) + ((g458) & (g463) & (!g468) & (g473) & (g147) & (g148)) + ((g458) & (g463) & (g468) & (!g473) & (!g147) & (!g148)) + ((g458) & (g463) & (g468) & (!g473) & (!g147) & (g148)) + ((g458) & (g463) & (g468) & (!g473) & (g147) & (!g148)) + ((g458) & (g463) & (g468) & (g473) & (!g147) & (!g148)) + ((g458) & (g463) & (g468) & (g473) & (!g147) & (g148)) + ((g458) & (g463) & (g468) & (g473) & (g147) & (!g148)) + ((g458) & (g463) & (g468) & (g473) & (g147) & (g148)));
	assign g4227 = (((!sk[28]) & (!g2173) & (!g3676) & (g475)) + ((!sk[28]) & (!g2173) & (g3676) & (!g475)) + ((!sk[28]) & (!g2173) & (g3676) & (g475)) + ((!sk[28]) & (g2173) & (!g3676) & (g475)) + ((!sk[28]) & (g2173) & (g3676) & (!g475)) + ((!sk[28]) & (g2173) & (g3676) & (g475)) + ((sk[28]) & (!g2173) & (!g3676) & (g475)) + ((sk[28]) & (!g2173) & (g3676) & (g475)) + ((sk[28]) & (g2173) & (g3676) & (!g475)) + ((sk[28]) & (g2173) & (g3676) & (g475)));
	assign g4228 = (((!g2174) & (!sk[29]) & (!g3676) & (g476)) + ((!g2174) & (!sk[29]) & (g3676) & (!g476)) + ((!g2174) & (!sk[29]) & (g3676) & (g476)) + ((!g2174) & (sk[29]) & (!g3676) & (g476)) + ((!g2174) & (sk[29]) & (g3676) & (g476)) + ((g2174) & (!sk[29]) & (!g3676) & (g476)) + ((g2174) & (!sk[29]) & (g3676) & (!g476)) + ((g2174) & (!sk[29]) & (g3676) & (g476)) + ((g2174) & (sk[29]) & (g3676) & (!g476)) + ((g2174) & (sk[29]) & (g3676) & (g476)));
	assign g4229 = (((!g2175) & (!sk[30]) & (!g3676) & (g477)) + ((!g2175) & (!sk[30]) & (g3676) & (!g477)) + ((!g2175) & (!sk[30]) & (g3676) & (g477)) + ((!g2175) & (sk[30]) & (!g3676) & (g477)) + ((!g2175) & (sk[30]) & (g3676) & (g477)) + ((g2175) & (!sk[30]) & (!g3676) & (g477)) + ((g2175) & (!sk[30]) & (g3676) & (!g477)) + ((g2175) & (!sk[30]) & (g3676) & (g477)) + ((g2175) & (sk[30]) & (g3676) & (!g477)) + ((g2175) & (sk[30]) & (g3676) & (g477)));
	assign g4230 = (((!sk[31]) & (!g2176) & (!g3676) & (g478)) + ((!sk[31]) & (!g2176) & (g3676) & (!g478)) + ((!sk[31]) & (!g2176) & (g3676) & (g478)) + ((!sk[31]) & (g2176) & (!g3676) & (g478)) + ((!sk[31]) & (g2176) & (g3676) & (!g478)) + ((!sk[31]) & (g2176) & (g3676) & (g478)) + ((sk[31]) & (!g2176) & (!g3676) & (g478)) + ((sk[31]) & (!g2176) & (g3676) & (g478)) + ((sk[31]) & (g2176) & (g3676) & (!g478)) + ((sk[31]) & (g2176) & (g3676) & (g478)));
	assign g479 = (((!g475) & (!g476) & (!g477) & (g478) & (g165) & (g166)) + ((!g475) & (!g476) & (g477) & (!g478) & (!g165) & (g166)) + ((!g475) & (!g476) & (g477) & (g478) & (!g165) & (g166)) + ((!g475) & (!g476) & (g477) & (g478) & (g165) & (g166)) + ((!g475) & (g476) & (!g477) & (!g478) & (g165) & (!g166)) + ((!g475) & (g476) & (!g477) & (g478) & (g165) & (!g166)) + ((!g475) & (g476) & (!g477) & (g478) & (g165) & (g166)) + ((!g475) & (g476) & (g477) & (!g478) & (!g165) & (g166)) + ((!g475) & (g476) & (g477) & (!g478) & (g165) & (!g166)) + ((!g475) & (g476) & (g477) & (g478) & (!g165) & (g166)) + ((!g475) & (g476) & (g477) & (g478) & (g165) & (!g166)) + ((!g475) & (g476) & (g477) & (g478) & (g165) & (g166)) + ((g475) & (!g476) & (!g477) & (!g478) & (!g165) & (!g166)) + ((g475) & (!g476) & (!g477) & (g478) & (!g165) & (!g166)) + ((g475) & (!g476) & (!g477) & (g478) & (g165) & (g166)) + ((g475) & (!g476) & (g477) & (!g478) & (!g165) & (!g166)) + ((g475) & (!g476) & (g477) & (!g478) & (!g165) & (g166)) + ((g475) & (!g476) & (g477) & (g478) & (!g165) & (!g166)) + ((g475) & (!g476) & (g477) & (g478) & (!g165) & (g166)) + ((g475) & (!g476) & (g477) & (g478) & (g165) & (g166)) + ((g475) & (g476) & (!g477) & (!g478) & (!g165) & (!g166)) + ((g475) & (g476) & (!g477) & (!g478) & (g165) & (!g166)) + ((g475) & (g476) & (!g477) & (g478) & (!g165) & (!g166)) + ((g475) & (g476) & (!g477) & (g478) & (g165) & (!g166)) + ((g475) & (g476) & (!g477) & (g478) & (g165) & (g166)) + ((g475) & (g476) & (g477) & (!g478) & (!g165) & (!g166)) + ((g475) & (g476) & (g477) & (!g478) & (!g165) & (g166)) + ((g475) & (g476) & (g477) & (!g478) & (g165) & (!g166)) + ((g475) & (g476) & (g477) & (g478) & (!g165) & (!g166)) + ((g475) & (g476) & (g477) & (g478) & (!g165) & (g166)) + ((g475) & (g476) & (g477) & (g478) & (g165) & (!g166)) + ((g475) & (g476) & (g477) & (g478) & (g165) & (g166)));
	assign g4231 = (((!g2177) & (!sk[33]) & (!g3676) & (g480)) + ((!g2177) & (!sk[33]) & (g3676) & (!g480)) + ((!g2177) & (!sk[33]) & (g3676) & (g480)) + ((!g2177) & (sk[33]) & (!g3676) & (g480)) + ((!g2177) & (sk[33]) & (g3676) & (g480)) + ((g2177) & (!sk[33]) & (!g3676) & (g480)) + ((g2177) & (!sk[33]) & (g3676) & (!g480)) + ((g2177) & (!sk[33]) & (g3676) & (g480)) + ((g2177) & (sk[33]) & (g3676) & (!g480)) + ((g2177) & (sk[33]) & (g3676) & (g480)));
	assign g4232 = (((!g2178) & (!sk[34]) & (!g3676) & (g481)) + ((!g2178) & (!sk[34]) & (g3676) & (!g481)) + ((!g2178) & (!sk[34]) & (g3676) & (g481)) + ((!g2178) & (sk[34]) & (!g3676) & (g481)) + ((!g2178) & (sk[34]) & (g3676) & (g481)) + ((g2178) & (!sk[34]) & (!g3676) & (g481)) + ((g2178) & (!sk[34]) & (g3676) & (!g481)) + ((g2178) & (!sk[34]) & (g3676) & (g481)) + ((g2178) & (sk[34]) & (g3676) & (!g481)) + ((g2178) & (sk[34]) & (g3676) & (g481)));
	assign g4233 = (((!g2179) & (!sk[35]) & (!g3676) & (g482)) + ((!g2179) & (!sk[35]) & (g3676) & (!g482)) + ((!g2179) & (!sk[35]) & (g3676) & (g482)) + ((!g2179) & (sk[35]) & (!g3676) & (g482)) + ((!g2179) & (sk[35]) & (g3676) & (g482)) + ((g2179) & (!sk[35]) & (!g3676) & (g482)) + ((g2179) & (!sk[35]) & (g3676) & (!g482)) + ((g2179) & (!sk[35]) & (g3676) & (g482)) + ((g2179) & (sk[35]) & (g3676) & (!g482)) + ((g2179) & (sk[35]) & (g3676) & (g482)));
	assign g483 = (((!g165) & (!g166) & (!g480) & (!sk[36]) & (g481) & (!g482)) + ((!g165) & (!g166) & (!g480) & (!sk[36]) & (g481) & (g482)) + ((!g165) & (!g166) & (g480) & (!sk[36]) & (!g481) & (!g482)) + ((!g165) & (!g166) & (g480) & (!sk[36]) & (!g481) & (g482)) + ((!g165) & (!g166) & (g480) & (!sk[36]) & (g481) & (!g482)) + ((!g165) & (!g166) & (g480) & (!sk[36]) & (g481) & (g482)) + ((!g165) & (g166) & (!g480) & (!sk[36]) & (!g481) & (!g482)) + ((!g165) & (g166) & (!g480) & (!sk[36]) & (!g481) & (g482)) + ((!g165) & (g166) & (!g480) & (!sk[36]) & (g481) & (!g482)) + ((!g165) & (g166) & (!g480) & (!sk[36]) & (g481) & (g482)) + ((!g165) & (g166) & (!g480) & (sk[36]) & (!g481) & (g482)) + ((!g165) & (g166) & (!g480) & (sk[36]) & (g481) & (g482)) + ((!g165) & (g166) & (g480) & (!sk[36]) & (!g481) & (!g482)) + ((!g165) & (g166) & (g480) & (!sk[36]) & (!g481) & (g482)) + ((!g165) & (g166) & (g480) & (!sk[36]) & (g481) & (!g482)) + ((!g165) & (g166) & (g480) & (!sk[36]) & (g481) & (g482)) + ((!g165) & (g166) & (g480) & (sk[36]) & (!g481) & (g482)) + ((!g165) & (g166) & (g480) & (sk[36]) & (g481) & (g482)) + ((g165) & (!g166) & (!g480) & (!sk[36]) & (g481) & (!g482)) + ((g165) & (!g166) & (!g480) & (!sk[36]) & (g481) & (g482)) + ((g165) & (!g166) & (g480) & (!sk[36]) & (!g481) & (!g482)) + ((g165) & (!g166) & (g480) & (!sk[36]) & (!g481) & (g482)) + ((g165) & (!g166) & (g480) & (!sk[36]) & (g481) & (!g482)) + ((g165) & (!g166) & (g480) & (!sk[36]) & (g481) & (g482)) + ((g165) & (!g166) & (g480) & (sk[36]) & (!g481) & (!g482)) + ((g165) & (!g166) & (g480) & (sk[36]) & (!g481) & (g482)) + ((g165) & (!g166) & (g480) & (sk[36]) & (g481) & (!g482)) + ((g165) & (!g166) & (g480) & (sk[36]) & (g481) & (g482)) + ((g165) & (g166) & (!g480) & (!sk[36]) & (!g481) & (!g482)) + ((g165) & (g166) & (!g480) & (!sk[36]) & (!g481) & (g482)) + ((g165) & (g166) & (!g480) & (!sk[36]) & (g481) & (!g482)) + ((g165) & (g166) & (!g480) & (!sk[36]) & (g481) & (g482)) + ((g165) & (g166) & (!g480) & (sk[36]) & (g481) & (!g482)) + ((g165) & (g166) & (!g480) & (sk[36]) & (g481) & (g482)) + ((g165) & (g166) & (g480) & (!sk[36]) & (!g481) & (!g482)) + ((g165) & (g166) & (g480) & (!sk[36]) & (!g481) & (g482)) + ((g165) & (g166) & (g480) & (!sk[36]) & (g481) & (!g482)) + ((g165) & (g166) & (g480) & (!sk[36]) & (g481) & (g482)) + ((g165) & (g166) & (g480) & (sk[36]) & (g481) & (!g482)) + ((g165) & (g166) & (g480) & (sk[36]) & (g481) & (g482)));
	assign g4234 = (((!g2162) & (!sk[37]) & (!g3676) & (g484)) + ((!g2162) & (!sk[37]) & (g3676) & (!g484)) + ((!g2162) & (!sk[37]) & (g3676) & (g484)) + ((!g2162) & (sk[37]) & (!g3676) & (g484)) + ((!g2162) & (sk[37]) & (g3676) & (g484)) + ((g2162) & (!sk[37]) & (!g3676) & (g484)) + ((g2162) & (!sk[37]) & (g3676) & (!g484)) + ((g2162) & (!sk[37]) & (g3676) & (g484)) + ((g2162) & (sk[37]) & (g3676) & (!g484)) + ((g2162) & (sk[37]) & (g3676) & (g484)));
	assign g4235 = (((!sk[38]) & (!g2164) & (!g3676) & (g485)) + ((!sk[38]) & (!g2164) & (g3676) & (!g485)) + ((!sk[38]) & (!g2164) & (g3676) & (g485)) + ((!sk[38]) & (g2164) & (!g3676) & (g485)) + ((!sk[38]) & (g2164) & (g3676) & (!g485)) + ((!sk[38]) & (g2164) & (g3676) & (g485)) + ((sk[38]) & (!g2164) & (!g3676) & (g485)) + ((sk[38]) & (!g2164) & (g3676) & (g485)) + ((sk[38]) & (g2164) & (g3676) & (!g485)) + ((sk[38]) & (g2164) & (g3676) & (g485)));
	assign g4236 = (((!g2166) & (!sk[39]) & (!g3676) & (g486)) + ((!g2166) & (!sk[39]) & (g3676) & (!g486)) + ((!g2166) & (!sk[39]) & (g3676) & (g486)) + ((!g2166) & (sk[39]) & (!g3676) & (g486)) + ((!g2166) & (sk[39]) & (g3676) & (g486)) + ((g2166) & (!sk[39]) & (!g3676) & (g486)) + ((g2166) & (!sk[39]) & (g3676) & (!g486)) + ((g2166) & (!sk[39]) & (g3676) & (g486)) + ((g2166) & (sk[39]) & (g3676) & (!g486)) + ((g2166) & (sk[39]) & (g3676) & (g486)));
	assign g4237 = (((!g2168) & (!sk[40]) & (!g3676) & (g487)) + ((!g2168) & (!sk[40]) & (g3676) & (!g487)) + ((!g2168) & (!sk[40]) & (g3676) & (g487)) + ((!g2168) & (sk[40]) & (!g3676) & (g487)) + ((!g2168) & (sk[40]) & (g3676) & (g487)) + ((g2168) & (!sk[40]) & (!g3676) & (g487)) + ((g2168) & (!sk[40]) & (g3676) & (!g487)) + ((g2168) & (!sk[40]) & (g3676) & (g487)) + ((g2168) & (sk[40]) & (g3676) & (!g487)) + ((g2168) & (sk[40]) & (g3676) & (g487)));
	assign g488 = (((!g484) & (!g485) & (!g486) & (g487) & (g165) & (g166)) + ((!g484) & (!g485) & (g486) & (!g487) & (!g165) & (g166)) + ((!g484) & (!g485) & (g486) & (g487) & (!g165) & (g166)) + ((!g484) & (!g485) & (g486) & (g487) & (g165) & (g166)) + ((!g484) & (g485) & (!g486) & (!g487) & (g165) & (!g166)) + ((!g484) & (g485) & (!g486) & (g487) & (g165) & (!g166)) + ((!g484) & (g485) & (!g486) & (g487) & (g165) & (g166)) + ((!g484) & (g485) & (g486) & (!g487) & (!g165) & (g166)) + ((!g484) & (g485) & (g486) & (!g487) & (g165) & (!g166)) + ((!g484) & (g485) & (g486) & (g487) & (!g165) & (g166)) + ((!g484) & (g485) & (g486) & (g487) & (g165) & (!g166)) + ((!g484) & (g485) & (g486) & (g487) & (g165) & (g166)) + ((g484) & (!g485) & (!g486) & (!g487) & (!g165) & (!g166)) + ((g484) & (!g485) & (!g486) & (g487) & (!g165) & (!g166)) + ((g484) & (!g485) & (!g486) & (g487) & (g165) & (g166)) + ((g484) & (!g485) & (g486) & (!g487) & (!g165) & (!g166)) + ((g484) & (!g485) & (g486) & (!g487) & (!g165) & (g166)) + ((g484) & (!g485) & (g486) & (g487) & (!g165) & (!g166)) + ((g484) & (!g485) & (g486) & (g487) & (!g165) & (g166)) + ((g484) & (!g485) & (g486) & (g487) & (g165) & (g166)) + ((g484) & (g485) & (!g486) & (!g487) & (!g165) & (!g166)) + ((g484) & (g485) & (!g486) & (!g487) & (g165) & (!g166)) + ((g484) & (g485) & (!g486) & (g487) & (!g165) & (!g166)) + ((g484) & (g485) & (!g486) & (g487) & (g165) & (!g166)) + ((g484) & (g485) & (!g486) & (g487) & (g165) & (g166)) + ((g484) & (g485) & (g486) & (!g487) & (!g165) & (!g166)) + ((g484) & (g485) & (g486) & (!g487) & (!g165) & (g166)) + ((g484) & (g485) & (g486) & (!g487) & (g165) & (!g166)) + ((g484) & (g485) & (g486) & (g487) & (!g165) & (!g166)) + ((g484) & (g485) & (g486) & (g487) & (!g165) & (g166)) + ((g484) & (g485) & (g486) & (g487) & (g165) & (!g166)) + ((g484) & (g485) & (g486) & (g487) & (g165) & (g166)));
	assign g4238 = (((!g2169) & (!g3676) & (!sk[42]) & (g489)) + ((!g2169) & (!g3676) & (sk[42]) & (g489)) + ((!g2169) & (g3676) & (!sk[42]) & (!g489)) + ((!g2169) & (g3676) & (!sk[42]) & (g489)) + ((!g2169) & (g3676) & (sk[42]) & (g489)) + ((g2169) & (!g3676) & (!sk[42]) & (g489)) + ((g2169) & (g3676) & (!sk[42]) & (!g489)) + ((g2169) & (g3676) & (!sk[42]) & (g489)) + ((g2169) & (g3676) & (sk[42]) & (!g489)) + ((g2169) & (g3676) & (sk[42]) & (g489)));
	assign g4239 = (((!g2170) & (!sk[43]) & (!g3676) & (g490)) + ((!g2170) & (!sk[43]) & (g3676) & (!g490)) + ((!g2170) & (!sk[43]) & (g3676) & (g490)) + ((!g2170) & (sk[43]) & (!g3676) & (g490)) + ((!g2170) & (sk[43]) & (g3676) & (g490)) + ((g2170) & (!sk[43]) & (!g3676) & (g490)) + ((g2170) & (!sk[43]) & (g3676) & (!g490)) + ((g2170) & (!sk[43]) & (g3676) & (g490)) + ((g2170) & (sk[43]) & (g3676) & (!g490)) + ((g2170) & (sk[43]) & (g3676) & (g490)));
	assign g4240 = (((!g2171) & (!sk[44]) & (!g3676) & (g491)) + ((!g2171) & (!sk[44]) & (g3676) & (!g491)) + ((!g2171) & (!sk[44]) & (g3676) & (g491)) + ((!g2171) & (sk[44]) & (!g3676) & (g491)) + ((!g2171) & (sk[44]) & (g3676) & (g491)) + ((g2171) & (!sk[44]) & (!g3676) & (g491)) + ((g2171) & (!sk[44]) & (g3676) & (!g491)) + ((g2171) & (!sk[44]) & (g3676) & (g491)) + ((g2171) & (sk[44]) & (g3676) & (!g491)) + ((g2171) & (sk[44]) & (g3676) & (g491)));
	assign g4241 = (((!g2172) & (!g3676) & (!sk[45]) & (g492)) + ((!g2172) & (!g3676) & (sk[45]) & (g492)) + ((!g2172) & (g3676) & (!sk[45]) & (!g492)) + ((!g2172) & (g3676) & (!sk[45]) & (g492)) + ((!g2172) & (g3676) & (sk[45]) & (g492)) + ((g2172) & (!g3676) & (!sk[45]) & (g492)) + ((g2172) & (g3676) & (!sk[45]) & (!g492)) + ((g2172) & (g3676) & (!sk[45]) & (g492)) + ((g2172) & (g3676) & (sk[45]) & (!g492)) + ((g2172) & (g3676) & (sk[45]) & (g492)));
	assign g493 = (((!g489) & (!g490) & (!g491) & (g492) & (g165) & (g166)) + ((!g489) & (!g490) & (g491) & (!g492) & (!g165) & (g166)) + ((!g489) & (!g490) & (g491) & (g492) & (!g165) & (g166)) + ((!g489) & (!g490) & (g491) & (g492) & (g165) & (g166)) + ((!g489) & (g490) & (!g491) & (!g492) & (g165) & (!g166)) + ((!g489) & (g490) & (!g491) & (g492) & (g165) & (!g166)) + ((!g489) & (g490) & (!g491) & (g492) & (g165) & (g166)) + ((!g489) & (g490) & (g491) & (!g492) & (!g165) & (g166)) + ((!g489) & (g490) & (g491) & (!g492) & (g165) & (!g166)) + ((!g489) & (g490) & (g491) & (g492) & (!g165) & (g166)) + ((!g489) & (g490) & (g491) & (g492) & (g165) & (!g166)) + ((!g489) & (g490) & (g491) & (g492) & (g165) & (g166)) + ((g489) & (!g490) & (!g491) & (!g492) & (!g165) & (!g166)) + ((g489) & (!g490) & (!g491) & (g492) & (!g165) & (!g166)) + ((g489) & (!g490) & (!g491) & (g492) & (g165) & (g166)) + ((g489) & (!g490) & (g491) & (!g492) & (!g165) & (!g166)) + ((g489) & (!g490) & (g491) & (!g492) & (!g165) & (g166)) + ((g489) & (!g490) & (g491) & (g492) & (!g165) & (!g166)) + ((g489) & (!g490) & (g491) & (g492) & (!g165) & (g166)) + ((g489) & (!g490) & (g491) & (g492) & (g165) & (g166)) + ((g489) & (g490) & (!g491) & (!g492) & (!g165) & (!g166)) + ((g489) & (g490) & (!g491) & (!g492) & (g165) & (!g166)) + ((g489) & (g490) & (!g491) & (g492) & (!g165) & (!g166)) + ((g489) & (g490) & (!g491) & (g492) & (g165) & (!g166)) + ((g489) & (g490) & (!g491) & (g492) & (g165) & (g166)) + ((g489) & (g490) & (g491) & (!g492) & (!g165) & (!g166)) + ((g489) & (g490) & (g491) & (!g492) & (!g165) & (g166)) + ((g489) & (g490) & (g491) & (!g492) & (g165) & (!g166)) + ((g489) & (g490) & (g491) & (g492) & (!g165) & (!g166)) + ((g489) & (g490) & (g491) & (g492) & (!g165) & (g166)) + ((g489) & (g490) & (g491) & (g492) & (g165) & (!g166)) + ((g489) & (g490) & (g491) & (g492) & (g165) & (g166)));
	assign g494 = (((!g147) & (!g148) & (!g479) & (g483) & (!g488) & (!g493)) + ((!g147) & (!g148) & (!g479) & (g483) & (!g488) & (g493)) + ((!g147) & (!g148) & (!g479) & (g483) & (g488) & (!g493)) + ((!g147) & (!g148) & (!g479) & (g483) & (g488) & (g493)) + ((!g147) & (!g148) & (g479) & (g483) & (!g488) & (!g493)) + ((!g147) & (!g148) & (g479) & (g483) & (!g488) & (g493)) + ((!g147) & (!g148) & (g479) & (g483) & (g488) & (!g493)) + ((!g147) & (!g148) & (g479) & (g483) & (g488) & (g493)) + ((!g147) & (g148) & (!g479) & (!g483) & (!g488) & (g493)) + ((!g147) & (g148) & (!g479) & (!g483) & (g488) & (g493)) + ((!g147) & (g148) & (!g479) & (g483) & (!g488) & (g493)) + ((!g147) & (g148) & (!g479) & (g483) & (g488) & (g493)) + ((!g147) & (g148) & (g479) & (!g483) & (!g488) & (g493)) + ((!g147) & (g148) & (g479) & (!g483) & (g488) & (g493)) + ((!g147) & (g148) & (g479) & (g483) & (!g488) & (g493)) + ((!g147) & (g148) & (g479) & (g483) & (g488) & (g493)) + ((g147) & (!g148) & (g479) & (!g483) & (!g488) & (!g493)) + ((g147) & (!g148) & (g479) & (!g483) & (!g488) & (g493)) + ((g147) & (!g148) & (g479) & (!g483) & (g488) & (!g493)) + ((g147) & (!g148) & (g479) & (!g483) & (g488) & (g493)) + ((g147) & (!g148) & (g479) & (g483) & (!g488) & (!g493)) + ((g147) & (!g148) & (g479) & (g483) & (!g488) & (g493)) + ((g147) & (!g148) & (g479) & (g483) & (g488) & (!g493)) + ((g147) & (!g148) & (g479) & (g483) & (g488) & (g493)) + ((g147) & (g148) & (!g479) & (!g483) & (g488) & (!g493)) + ((g147) & (g148) & (!g479) & (!g483) & (g488) & (g493)) + ((g147) & (g148) & (!g479) & (g483) & (g488) & (!g493)) + ((g147) & (g148) & (!g479) & (g483) & (g488) & (g493)) + ((g147) & (g148) & (g479) & (!g483) & (g488) & (!g493)) + ((g147) & (g148) & (g479) & (!g483) & (g488) & (g493)) + ((g147) & (g148) & (g479) & (g483) & (g488) & (!g493)) + ((g147) & (g148) & (g479) & (g483) & (g488) & (g493)));
	assign g495 = (((!g142) & (!sk[48]) & (!g474) & (g494)) + ((!g142) & (!sk[48]) & (g474) & (!g494)) + ((!g142) & (!sk[48]) & (g474) & (g494)) + ((!g142) & (sk[48]) & (!g474) & (g494)) + ((!g142) & (sk[48]) & (g474) & (g494)) + ((g142) & (!sk[48]) & (!g474) & (g494)) + ((g142) & (!sk[48]) & (g474) & (!g494)) + ((g142) & (!sk[48]) & (g474) & (g494)) + ((g142) & (sk[48]) & (g474) & (!g494)) + ((g142) & (sk[48]) & (g474) & (g494)));
	assign g4242 = (((sk[49]) & (!g2361)));
	assign g4243 = (((!g2059) & (!g4242) & (!sk[50]) & (g496)) + ((!g2059) & (!g4242) & (sk[50]) & (g496)) + ((!g2059) & (g4242) & (!sk[50]) & (!g496)) + ((!g2059) & (g4242) & (!sk[50]) & (g496)) + ((!g2059) & (g4242) & (sk[50]) & (g496)) + ((g2059) & (!g4242) & (!sk[50]) & (g496)) + ((g2059) & (g4242) & (!sk[50]) & (!g496)) + ((g2059) & (g4242) & (!sk[50]) & (g496)) + ((g2059) & (g4242) & (sk[50]) & (!g496)) + ((g2059) & (g4242) & (sk[50]) & (g496)));
	assign g497 = (((!g85) & (!sk[51]) & (!g86) & (!g409) & (g451) & (!g495)) + ((!g85) & (!sk[51]) & (!g86) & (!g409) & (g451) & (g495)) + ((!g85) & (!sk[51]) & (!g86) & (g409) & (!g451) & (!g495)) + ((!g85) & (!sk[51]) & (!g86) & (g409) & (!g451) & (g495)) + ((!g85) & (!sk[51]) & (!g86) & (g409) & (g451) & (!g495)) + ((!g85) & (!sk[51]) & (!g86) & (g409) & (g451) & (g495)) + ((!g85) & (!sk[51]) & (g86) & (!g409) & (!g451) & (!g495)) + ((!g85) & (!sk[51]) & (g86) & (!g409) & (!g451) & (g495)) + ((!g85) & (!sk[51]) & (g86) & (!g409) & (g451) & (!g495)) + ((!g85) & (!sk[51]) & (g86) & (!g409) & (g451) & (g495)) + ((!g85) & (!sk[51]) & (g86) & (g409) & (!g451) & (!g495)) + ((!g85) & (!sk[51]) & (g86) & (g409) & (!g451) & (g495)) + ((!g85) & (!sk[51]) & (g86) & (g409) & (g451) & (!g495)) + ((!g85) & (!sk[51]) & (g86) & (g409) & (g451) & (g495)) + ((!g85) & (sk[51]) & (!g86) & (g409) & (g451) & (g495)) + ((!g85) & (sk[51]) & (g86) & (!g409) & (g451) & (g495)) + ((!g85) & (sk[51]) & (g86) & (g409) & (!g451) & (g495)) + ((!g85) & (sk[51]) & (g86) & (g409) & (g451) & (g495)) + ((g85) & (!sk[51]) & (!g86) & (!g409) & (g451) & (!g495)) + ((g85) & (!sk[51]) & (!g86) & (!g409) & (g451) & (g495)) + ((g85) & (!sk[51]) & (!g86) & (g409) & (!g451) & (!g495)) + ((g85) & (!sk[51]) & (!g86) & (g409) & (!g451) & (g495)) + ((g85) & (!sk[51]) & (!g86) & (g409) & (g451) & (!g495)) + ((g85) & (!sk[51]) & (!g86) & (g409) & (g451) & (g495)) + ((g85) & (!sk[51]) & (g86) & (!g409) & (!g451) & (!g495)) + ((g85) & (!sk[51]) & (g86) & (!g409) & (!g451) & (g495)) + ((g85) & (!sk[51]) & (g86) & (!g409) & (g451) & (!g495)) + ((g85) & (!sk[51]) & (g86) & (!g409) & (g451) & (g495)) + ((g85) & (!sk[51]) & (g86) & (g409) & (!g451) & (!g495)) + ((g85) & (!sk[51]) & (g86) & (g409) & (!g451) & (g495)) + ((g85) & (!sk[51]) & (g86) & (g409) & (g451) & (!g495)) + ((g85) & (!sk[51]) & (g86) & (g409) & (g451) & (g495)) + ((g85) & (sk[51]) & (!g86) & (!g409) & (!g451) & (g495)) + ((g85) & (sk[51]) & (!g86) & (!g409) & (g451) & (g495)) + ((g85) & (sk[51]) & (!g86) & (g409) & (!g451) & (g495)) + ((g85) & (sk[51]) & (!g86) & (g409) & (g451) & (!g495)) + ((g85) & (sk[51]) & (!g86) & (g409) & (g451) & (g495)) + ((g85) & (sk[51]) & (g86) & (!g409) & (!g451) & (g495)) + ((g85) & (sk[51]) & (g86) & (!g409) & (g451) & (!g495)) + ((g85) & (sk[51]) & (g86) & (!g409) & (g451) & (g495)) + ((g85) & (sk[51]) & (g86) & (g409) & (!g451) & (!g495)) + ((g85) & (sk[51]) & (g86) & (g409) & (!g451) & (g495)) + ((g85) & (sk[51]) & (g86) & (g409) & (g451) & (!g495)) + ((g85) & (sk[51]) & (g86) & (g409) & (g451) & (g495)));
	assign g4244 = (((!g2140) & (!g2378) & (!sk[52]) & (g498)) + ((!g2140) & (!g2378) & (sk[52]) & (g498)) + ((!g2140) & (g2378) & (!sk[52]) & (!g498)) + ((!g2140) & (g2378) & (!sk[52]) & (g498)) + ((!g2140) & (g2378) & (sk[52]) & (g498)) + ((g2140) & (!g2378) & (!sk[52]) & (g498)) + ((g2140) & (g2378) & (!sk[52]) & (!g498)) + ((g2140) & (g2378) & (!sk[52]) & (g498)) + ((g2140) & (g2378) & (sk[52]) & (!g498)) + ((g2140) & (g2378) & (sk[52]) & (g498)));
	assign g4245 = (((!g2142) & (!g2378) & (!sk[53]) & (g499)) + ((!g2142) & (!g2378) & (sk[53]) & (g499)) + ((!g2142) & (g2378) & (!sk[53]) & (!g499)) + ((!g2142) & (g2378) & (!sk[53]) & (g499)) + ((!g2142) & (g2378) & (sk[53]) & (g499)) + ((g2142) & (!g2378) & (!sk[53]) & (g499)) + ((g2142) & (g2378) & (!sk[53]) & (!g499)) + ((g2142) & (g2378) & (!sk[53]) & (g499)) + ((g2142) & (g2378) & (sk[53]) & (!g499)) + ((g2142) & (g2378) & (sk[53]) & (g499)));
	assign g4246 = (((!sk[54]) & (!g2144) & (!g2378) & (g500)) + ((!sk[54]) & (!g2144) & (g2378) & (!g500)) + ((!sk[54]) & (!g2144) & (g2378) & (g500)) + ((!sk[54]) & (g2144) & (!g2378) & (g500)) + ((!sk[54]) & (g2144) & (g2378) & (!g500)) + ((!sk[54]) & (g2144) & (g2378) & (g500)) + ((sk[54]) & (!g2144) & (!g2378) & (g500)) + ((sk[54]) & (!g2144) & (g2378) & (g500)) + ((sk[54]) & (g2144) & (g2378) & (!g500)) + ((sk[54]) & (g2144) & (g2378) & (g500)));
	assign g4247 = (((!sk[55]) & (!g2145) & (!g2378) & (g501)) + ((!sk[55]) & (!g2145) & (g2378) & (!g501)) + ((!sk[55]) & (!g2145) & (g2378) & (g501)) + ((!sk[55]) & (g2145) & (!g2378) & (g501)) + ((!sk[55]) & (g2145) & (g2378) & (!g501)) + ((!sk[55]) & (g2145) & (g2378) & (g501)) + ((sk[55]) & (!g2145) & (!g2378) & (g501)) + ((sk[55]) & (!g2145) & (g2378) & (g501)) + ((sk[55]) & (g2145) & (g2378) & (!g501)) + ((sk[55]) & (g2145) & (g2378) & (g501)));
	assign g502 = (((!g498) & (!g499) & (!g500) & (g501) & (g147) & (g148)) + ((!g498) & (!g499) & (g500) & (!g501) & (!g147) & (g148)) + ((!g498) & (!g499) & (g500) & (g501) & (!g147) & (g148)) + ((!g498) & (!g499) & (g500) & (g501) & (g147) & (g148)) + ((!g498) & (g499) & (!g500) & (!g501) & (g147) & (!g148)) + ((!g498) & (g499) & (!g500) & (g501) & (g147) & (!g148)) + ((!g498) & (g499) & (!g500) & (g501) & (g147) & (g148)) + ((!g498) & (g499) & (g500) & (!g501) & (!g147) & (g148)) + ((!g498) & (g499) & (g500) & (!g501) & (g147) & (!g148)) + ((!g498) & (g499) & (g500) & (g501) & (!g147) & (g148)) + ((!g498) & (g499) & (g500) & (g501) & (g147) & (!g148)) + ((!g498) & (g499) & (g500) & (g501) & (g147) & (g148)) + ((g498) & (!g499) & (!g500) & (!g501) & (!g147) & (!g148)) + ((g498) & (!g499) & (!g500) & (g501) & (!g147) & (!g148)) + ((g498) & (!g499) & (!g500) & (g501) & (g147) & (g148)) + ((g498) & (!g499) & (g500) & (!g501) & (!g147) & (!g148)) + ((g498) & (!g499) & (g500) & (!g501) & (!g147) & (g148)) + ((g498) & (!g499) & (g500) & (g501) & (!g147) & (!g148)) + ((g498) & (!g499) & (g500) & (g501) & (!g147) & (g148)) + ((g498) & (!g499) & (g500) & (g501) & (g147) & (g148)) + ((g498) & (g499) & (!g500) & (!g501) & (!g147) & (!g148)) + ((g498) & (g499) & (!g500) & (!g501) & (g147) & (!g148)) + ((g498) & (g499) & (!g500) & (g501) & (!g147) & (!g148)) + ((g498) & (g499) & (!g500) & (g501) & (g147) & (!g148)) + ((g498) & (g499) & (!g500) & (g501) & (g147) & (g148)) + ((g498) & (g499) & (g500) & (!g501) & (!g147) & (!g148)) + ((g498) & (g499) & (g500) & (!g501) & (!g147) & (g148)) + ((g498) & (g499) & (g500) & (!g501) & (g147) & (!g148)) + ((g498) & (g499) & (g500) & (g501) & (!g147) & (!g148)) + ((g498) & (g499) & (g500) & (g501) & (!g147) & (g148)) + ((g498) & (g499) & (g500) & (g501) & (g147) & (!g148)) + ((g498) & (g499) & (g500) & (g501) & (g147) & (g148)));
	assign g4248 = (((!g2146) & (!sk[57]) & (!g2378) & (g503)) + ((!g2146) & (!sk[57]) & (g2378) & (!g503)) + ((!g2146) & (!sk[57]) & (g2378) & (g503)) + ((!g2146) & (sk[57]) & (!g2378) & (g503)) + ((!g2146) & (sk[57]) & (g2378) & (g503)) + ((g2146) & (!sk[57]) & (!g2378) & (g503)) + ((g2146) & (!sk[57]) & (g2378) & (!g503)) + ((g2146) & (!sk[57]) & (g2378) & (g503)) + ((g2146) & (sk[57]) & (g2378) & (!g503)) + ((g2146) & (sk[57]) & (g2378) & (g503)));
	assign g4249 = (((!g2148) & (!sk[58]) & (!g2378) & (g504)) + ((!g2148) & (!sk[58]) & (g2378) & (!g504)) + ((!g2148) & (!sk[58]) & (g2378) & (g504)) + ((!g2148) & (sk[58]) & (!g2378) & (g504)) + ((!g2148) & (sk[58]) & (g2378) & (g504)) + ((g2148) & (!sk[58]) & (!g2378) & (g504)) + ((g2148) & (!sk[58]) & (g2378) & (!g504)) + ((g2148) & (!sk[58]) & (g2378) & (g504)) + ((g2148) & (sk[58]) & (g2378) & (!g504)) + ((g2148) & (sk[58]) & (g2378) & (g504)));
	assign g4250 = (((!sk[59]) & (!g2150) & (!g2378) & (g505)) + ((!sk[59]) & (!g2150) & (g2378) & (!g505)) + ((!sk[59]) & (!g2150) & (g2378) & (g505)) + ((!sk[59]) & (g2150) & (!g2378) & (g505)) + ((!sk[59]) & (g2150) & (g2378) & (!g505)) + ((!sk[59]) & (g2150) & (g2378) & (g505)) + ((sk[59]) & (!g2150) & (!g2378) & (g505)) + ((sk[59]) & (!g2150) & (g2378) & (g505)) + ((sk[59]) & (g2150) & (g2378) & (!g505)) + ((sk[59]) & (g2150) & (g2378) & (g505)));
	assign g4251 = (((!g2151) & (!g2378) & (!sk[60]) & (g506)) + ((!g2151) & (!g2378) & (sk[60]) & (g506)) + ((!g2151) & (g2378) & (!sk[60]) & (!g506)) + ((!g2151) & (g2378) & (!sk[60]) & (g506)) + ((!g2151) & (g2378) & (sk[60]) & (g506)) + ((g2151) & (!g2378) & (!sk[60]) & (g506)) + ((g2151) & (g2378) & (!sk[60]) & (!g506)) + ((g2151) & (g2378) & (!sk[60]) & (g506)) + ((g2151) & (g2378) & (sk[60]) & (!g506)) + ((g2151) & (g2378) & (sk[60]) & (g506)));
	assign g507 = (((!g503) & (!g504) & (!g505) & (g506) & (g147) & (g148)) + ((!g503) & (!g504) & (g505) & (!g506) & (!g147) & (g148)) + ((!g503) & (!g504) & (g505) & (g506) & (!g147) & (g148)) + ((!g503) & (!g504) & (g505) & (g506) & (g147) & (g148)) + ((!g503) & (g504) & (!g505) & (!g506) & (g147) & (!g148)) + ((!g503) & (g504) & (!g505) & (g506) & (g147) & (!g148)) + ((!g503) & (g504) & (!g505) & (g506) & (g147) & (g148)) + ((!g503) & (g504) & (g505) & (!g506) & (!g147) & (g148)) + ((!g503) & (g504) & (g505) & (!g506) & (g147) & (!g148)) + ((!g503) & (g504) & (g505) & (g506) & (!g147) & (g148)) + ((!g503) & (g504) & (g505) & (g506) & (g147) & (!g148)) + ((!g503) & (g504) & (g505) & (g506) & (g147) & (g148)) + ((g503) & (!g504) & (!g505) & (!g506) & (!g147) & (!g148)) + ((g503) & (!g504) & (!g505) & (g506) & (!g147) & (!g148)) + ((g503) & (!g504) & (!g505) & (g506) & (g147) & (g148)) + ((g503) & (!g504) & (g505) & (!g506) & (!g147) & (!g148)) + ((g503) & (!g504) & (g505) & (!g506) & (!g147) & (g148)) + ((g503) & (!g504) & (g505) & (g506) & (!g147) & (!g148)) + ((g503) & (!g504) & (g505) & (g506) & (!g147) & (g148)) + ((g503) & (!g504) & (g505) & (g506) & (g147) & (g148)) + ((g503) & (g504) & (!g505) & (!g506) & (!g147) & (!g148)) + ((g503) & (g504) & (!g505) & (!g506) & (g147) & (!g148)) + ((g503) & (g504) & (!g505) & (g506) & (!g147) & (!g148)) + ((g503) & (g504) & (!g505) & (g506) & (g147) & (!g148)) + ((g503) & (g504) & (!g505) & (g506) & (g147) & (g148)) + ((g503) & (g504) & (g505) & (!g506) & (!g147) & (!g148)) + ((g503) & (g504) & (g505) & (!g506) & (!g147) & (g148)) + ((g503) & (g504) & (g505) & (!g506) & (g147) & (!g148)) + ((g503) & (g504) & (g505) & (g506) & (!g147) & (!g148)) + ((g503) & (g504) & (g505) & (g506) & (!g147) & (g148)) + ((g503) & (g504) & (g505) & (g506) & (g147) & (!g148)) + ((g503) & (g504) & (g505) & (g506) & (g147) & (g148)));
	assign g4252 = (((!sk[62]) & (!g2152) & (!g2378) & (g508)) + ((!sk[62]) & (!g2152) & (g2378) & (!g508)) + ((!sk[62]) & (!g2152) & (g2378) & (g508)) + ((!sk[62]) & (g2152) & (!g2378) & (g508)) + ((!sk[62]) & (g2152) & (g2378) & (!g508)) + ((!sk[62]) & (g2152) & (g2378) & (g508)) + ((sk[62]) & (!g2152) & (!g2378) & (g508)) + ((sk[62]) & (!g2152) & (g2378) & (g508)) + ((sk[62]) & (g2152) & (g2378) & (!g508)) + ((sk[62]) & (g2152) & (g2378) & (g508)));
	assign g4253 = (((!g2153) & (!sk[63]) & (!g2378) & (g509)) + ((!g2153) & (!sk[63]) & (g2378) & (!g509)) + ((!g2153) & (!sk[63]) & (g2378) & (g509)) + ((!g2153) & (sk[63]) & (!g2378) & (g509)) + ((!g2153) & (sk[63]) & (g2378) & (g509)) + ((g2153) & (!sk[63]) & (!g2378) & (g509)) + ((g2153) & (!sk[63]) & (g2378) & (!g509)) + ((g2153) & (!sk[63]) & (g2378) & (g509)) + ((g2153) & (sk[63]) & (g2378) & (!g509)) + ((g2153) & (sk[63]) & (g2378) & (g509)));
	assign g4254 = (((!g2155) & (!g2378) & (!sk[64]) & (g510)) + ((!g2155) & (!g2378) & (sk[64]) & (g510)) + ((!g2155) & (g2378) & (!sk[64]) & (!g510)) + ((!g2155) & (g2378) & (!sk[64]) & (g510)) + ((!g2155) & (g2378) & (sk[64]) & (g510)) + ((g2155) & (!g2378) & (!sk[64]) & (g510)) + ((g2155) & (g2378) & (!sk[64]) & (!g510)) + ((g2155) & (g2378) & (!sk[64]) & (g510)) + ((g2155) & (g2378) & (sk[64]) & (!g510)) + ((g2155) & (g2378) & (sk[64]) & (g510)));
	assign g4255 = (((!sk[65]) & (!g2157) & (!g2378) & (g511)) + ((!sk[65]) & (!g2157) & (g2378) & (!g511)) + ((!sk[65]) & (!g2157) & (g2378) & (g511)) + ((!sk[65]) & (g2157) & (!g2378) & (g511)) + ((!sk[65]) & (g2157) & (g2378) & (!g511)) + ((!sk[65]) & (g2157) & (g2378) & (g511)) + ((sk[65]) & (!g2157) & (!g2378) & (g511)) + ((sk[65]) & (!g2157) & (g2378) & (g511)) + ((sk[65]) & (g2157) & (g2378) & (!g511)) + ((sk[65]) & (g2157) & (g2378) & (g511)));
	assign g512 = (((!g508) & (!g509) & (!g510) & (g511) & (g147) & (g148)) + ((!g508) & (!g509) & (g510) & (!g511) & (!g147) & (g148)) + ((!g508) & (!g509) & (g510) & (g511) & (!g147) & (g148)) + ((!g508) & (!g509) & (g510) & (g511) & (g147) & (g148)) + ((!g508) & (g509) & (!g510) & (!g511) & (g147) & (!g148)) + ((!g508) & (g509) & (!g510) & (g511) & (g147) & (!g148)) + ((!g508) & (g509) & (!g510) & (g511) & (g147) & (g148)) + ((!g508) & (g509) & (g510) & (!g511) & (!g147) & (g148)) + ((!g508) & (g509) & (g510) & (!g511) & (g147) & (!g148)) + ((!g508) & (g509) & (g510) & (g511) & (!g147) & (g148)) + ((!g508) & (g509) & (g510) & (g511) & (g147) & (!g148)) + ((!g508) & (g509) & (g510) & (g511) & (g147) & (g148)) + ((g508) & (!g509) & (!g510) & (!g511) & (!g147) & (!g148)) + ((g508) & (!g509) & (!g510) & (g511) & (!g147) & (!g148)) + ((g508) & (!g509) & (!g510) & (g511) & (g147) & (g148)) + ((g508) & (!g509) & (g510) & (!g511) & (!g147) & (!g148)) + ((g508) & (!g509) & (g510) & (!g511) & (!g147) & (g148)) + ((g508) & (!g509) & (g510) & (g511) & (!g147) & (!g148)) + ((g508) & (!g509) & (g510) & (g511) & (!g147) & (g148)) + ((g508) & (!g509) & (g510) & (g511) & (g147) & (g148)) + ((g508) & (g509) & (!g510) & (!g511) & (!g147) & (!g148)) + ((g508) & (g509) & (!g510) & (!g511) & (g147) & (!g148)) + ((g508) & (g509) & (!g510) & (g511) & (!g147) & (!g148)) + ((g508) & (g509) & (!g510) & (g511) & (g147) & (!g148)) + ((g508) & (g509) & (!g510) & (g511) & (g147) & (g148)) + ((g508) & (g509) & (g510) & (!g511) & (!g147) & (!g148)) + ((g508) & (g509) & (g510) & (!g511) & (!g147) & (g148)) + ((g508) & (g509) & (g510) & (!g511) & (g147) & (!g148)) + ((g508) & (g509) & (g510) & (g511) & (!g147) & (!g148)) + ((g508) & (g509) & (g510) & (g511) & (!g147) & (g148)) + ((g508) & (g509) & (g510) & (g511) & (g147) & (!g148)) + ((g508) & (g509) & (g510) & (g511) & (g147) & (g148)));
	assign g4256 = (((!sk[67]) & (!g2158) & (!g2378) & (g513)) + ((!sk[67]) & (!g2158) & (g2378) & (!g513)) + ((!sk[67]) & (!g2158) & (g2378) & (g513)) + ((!sk[67]) & (g2158) & (!g2378) & (g513)) + ((!sk[67]) & (g2158) & (g2378) & (!g513)) + ((!sk[67]) & (g2158) & (g2378) & (g513)) + ((sk[67]) & (!g2158) & (!g2378) & (g513)) + ((sk[67]) & (!g2158) & (g2378) & (g513)) + ((sk[67]) & (g2158) & (g2378) & (!g513)) + ((sk[67]) & (g2158) & (g2378) & (g513)));
	assign g4257 = (((!g2159) & (!g2378) & (!sk[68]) & (g514)) + ((!g2159) & (!g2378) & (sk[68]) & (g514)) + ((!g2159) & (g2378) & (!sk[68]) & (!g514)) + ((!g2159) & (g2378) & (!sk[68]) & (g514)) + ((!g2159) & (g2378) & (sk[68]) & (g514)) + ((g2159) & (!g2378) & (!sk[68]) & (g514)) + ((g2159) & (g2378) & (!sk[68]) & (!g514)) + ((g2159) & (g2378) & (!sk[68]) & (g514)) + ((g2159) & (g2378) & (sk[68]) & (!g514)) + ((g2159) & (g2378) & (sk[68]) & (g514)));
	assign g4258 = (((!g2160) & (!g2378) & (!sk[69]) & (g515)) + ((!g2160) & (!g2378) & (sk[69]) & (g515)) + ((!g2160) & (g2378) & (!sk[69]) & (!g515)) + ((!g2160) & (g2378) & (!sk[69]) & (g515)) + ((!g2160) & (g2378) & (sk[69]) & (g515)) + ((g2160) & (!g2378) & (!sk[69]) & (g515)) + ((g2160) & (g2378) & (!sk[69]) & (!g515)) + ((g2160) & (g2378) & (!sk[69]) & (g515)) + ((g2160) & (g2378) & (sk[69]) & (!g515)) + ((g2160) & (g2378) & (sk[69]) & (g515)));
	assign g4259 = (((!g2161) & (!g2378) & (!sk[70]) & (g516)) + ((!g2161) & (!g2378) & (sk[70]) & (g516)) + ((!g2161) & (g2378) & (!sk[70]) & (!g516)) + ((!g2161) & (g2378) & (!sk[70]) & (g516)) + ((!g2161) & (g2378) & (sk[70]) & (g516)) + ((g2161) & (!g2378) & (!sk[70]) & (g516)) + ((g2161) & (g2378) & (!sk[70]) & (!g516)) + ((g2161) & (g2378) & (!sk[70]) & (g516)) + ((g2161) & (g2378) & (sk[70]) & (!g516)) + ((g2161) & (g2378) & (sk[70]) & (g516)));
	assign g517 = (((!g513) & (!g514) & (!g515) & (g516) & (g147) & (g148)) + ((!g513) & (!g514) & (g515) & (!g516) & (!g147) & (g148)) + ((!g513) & (!g514) & (g515) & (g516) & (!g147) & (g148)) + ((!g513) & (!g514) & (g515) & (g516) & (g147) & (g148)) + ((!g513) & (g514) & (!g515) & (!g516) & (g147) & (!g148)) + ((!g513) & (g514) & (!g515) & (g516) & (g147) & (!g148)) + ((!g513) & (g514) & (!g515) & (g516) & (g147) & (g148)) + ((!g513) & (g514) & (g515) & (!g516) & (!g147) & (g148)) + ((!g513) & (g514) & (g515) & (!g516) & (g147) & (!g148)) + ((!g513) & (g514) & (g515) & (g516) & (!g147) & (g148)) + ((!g513) & (g514) & (g515) & (g516) & (g147) & (!g148)) + ((!g513) & (g514) & (g515) & (g516) & (g147) & (g148)) + ((g513) & (!g514) & (!g515) & (!g516) & (!g147) & (!g148)) + ((g513) & (!g514) & (!g515) & (g516) & (!g147) & (!g148)) + ((g513) & (!g514) & (!g515) & (g516) & (g147) & (g148)) + ((g513) & (!g514) & (g515) & (!g516) & (!g147) & (!g148)) + ((g513) & (!g514) & (g515) & (!g516) & (!g147) & (g148)) + ((g513) & (!g514) & (g515) & (g516) & (!g147) & (!g148)) + ((g513) & (!g514) & (g515) & (g516) & (!g147) & (g148)) + ((g513) & (!g514) & (g515) & (g516) & (g147) & (g148)) + ((g513) & (g514) & (!g515) & (!g516) & (!g147) & (!g148)) + ((g513) & (g514) & (!g515) & (!g516) & (g147) & (!g148)) + ((g513) & (g514) & (!g515) & (g516) & (!g147) & (!g148)) + ((g513) & (g514) & (!g515) & (g516) & (g147) & (!g148)) + ((g513) & (g514) & (!g515) & (g516) & (g147) & (g148)) + ((g513) & (g514) & (g515) & (!g516) & (!g147) & (!g148)) + ((g513) & (g514) & (g515) & (!g516) & (!g147) & (g148)) + ((g513) & (g514) & (g515) & (!g516) & (g147) & (!g148)) + ((g513) & (g514) & (g515) & (g516) & (!g147) & (!g148)) + ((g513) & (g514) & (g515) & (g516) & (!g147) & (g148)) + ((g513) & (g514) & (g515) & (g516) & (g147) & (!g148)) + ((g513) & (g514) & (g515) & (g516) & (g147) & (g148)));
	assign g518 = (((!g502) & (!g507) & (!g512) & (g517) & (g165) & (g166)) + ((!g502) & (!g507) & (g512) & (!g517) & (!g165) & (g166)) + ((!g502) & (!g507) & (g512) & (g517) & (!g165) & (g166)) + ((!g502) & (!g507) & (g512) & (g517) & (g165) & (g166)) + ((!g502) & (g507) & (!g512) & (!g517) & (g165) & (!g166)) + ((!g502) & (g507) & (!g512) & (g517) & (g165) & (!g166)) + ((!g502) & (g507) & (!g512) & (g517) & (g165) & (g166)) + ((!g502) & (g507) & (g512) & (!g517) & (!g165) & (g166)) + ((!g502) & (g507) & (g512) & (!g517) & (g165) & (!g166)) + ((!g502) & (g507) & (g512) & (g517) & (!g165) & (g166)) + ((!g502) & (g507) & (g512) & (g517) & (g165) & (!g166)) + ((!g502) & (g507) & (g512) & (g517) & (g165) & (g166)) + ((g502) & (!g507) & (!g512) & (!g517) & (!g165) & (!g166)) + ((g502) & (!g507) & (!g512) & (g517) & (!g165) & (!g166)) + ((g502) & (!g507) & (!g512) & (g517) & (g165) & (g166)) + ((g502) & (!g507) & (g512) & (!g517) & (!g165) & (!g166)) + ((g502) & (!g507) & (g512) & (!g517) & (!g165) & (g166)) + ((g502) & (!g507) & (g512) & (g517) & (!g165) & (!g166)) + ((g502) & (!g507) & (g512) & (g517) & (!g165) & (g166)) + ((g502) & (!g507) & (g512) & (g517) & (g165) & (g166)) + ((g502) & (g507) & (!g512) & (!g517) & (!g165) & (!g166)) + ((g502) & (g507) & (!g512) & (!g517) & (g165) & (!g166)) + ((g502) & (g507) & (!g512) & (g517) & (!g165) & (!g166)) + ((g502) & (g507) & (!g512) & (g517) & (g165) & (!g166)) + ((g502) & (g507) & (!g512) & (g517) & (g165) & (g166)) + ((g502) & (g507) & (g512) & (!g517) & (!g165) & (!g166)) + ((g502) & (g507) & (g512) & (!g517) & (!g165) & (g166)) + ((g502) & (g507) & (g512) & (!g517) & (g165) & (!g166)) + ((g502) & (g507) & (g512) & (g517) & (!g165) & (!g166)) + ((g502) & (g507) & (g512) & (g517) & (!g165) & (g166)) + ((g502) & (g507) & (g512) & (g517) & (g165) & (!g166)) + ((g502) & (g507) & (g512) & (g517) & (g165) & (g166)));
	assign g4260 = (((!g2173) & (!g2378) & (!sk[73]) & (g519)) + ((!g2173) & (!g2378) & (sk[73]) & (g519)) + ((!g2173) & (g2378) & (!sk[73]) & (!g519)) + ((!g2173) & (g2378) & (!sk[73]) & (g519)) + ((!g2173) & (g2378) & (sk[73]) & (g519)) + ((g2173) & (!g2378) & (!sk[73]) & (g519)) + ((g2173) & (g2378) & (!sk[73]) & (!g519)) + ((g2173) & (g2378) & (!sk[73]) & (g519)) + ((g2173) & (g2378) & (sk[73]) & (!g519)) + ((g2173) & (g2378) & (sk[73]) & (g519)));
	assign g4261 = (((!g2174) & (!g2378) & (!sk[74]) & (g520)) + ((!g2174) & (!g2378) & (sk[74]) & (g520)) + ((!g2174) & (g2378) & (!sk[74]) & (!g520)) + ((!g2174) & (g2378) & (!sk[74]) & (g520)) + ((!g2174) & (g2378) & (sk[74]) & (g520)) + ((g2174) & (!g2378) & (!sk[74]) & (g520)) + ((g2174) & (g2378) & (!sk[74]) & (!g520)) + ((g2174) & (g2378) & (!sk[74]) & (g520)) + ((g2174) & (g2378) & (sk[74]) & (!g520)) + ((g2174) & (g2378) & (sk[74]) & (g520)));
	assign g4262 = (((!g2175) & (!g2378) & (!sk[75]) & (g521)) + ((!g2175) & (!g2378) & (sk[75]) & (g521)) + ((!g2175) & (g2378) & (!sk[75]) & (!g521)) + ((!g2175) & (g2378) & (!sk[75]) & (g521)) + ((!g2175) & (g2378) & (sk[75]) & (g521)) + ((g2175) & (!g2378) & (!sk[75]) & (g521)) + ((g2175) & (g2378) & (!sk[75]) & (!g521)) + ((g2175) & (g2378) & (!sk[75]) & (g521)) + ((g2175) & (g2378) & (sk[75]) & (!g521)) + ((g2175) & (g2378) & (sk[75]) & (g521)));
	assign g4263 = (((!g2176) & (!g2378) & (!sk[76]) & (g522)) + ((!g2176) & (!g2378) & (sk[76]) & (g522)) + ((!g2176) & (g2378) & (!sk[76]) & (!g522)) + ((!g2176) & (g2378) & (!sk[76]) & (g522)) + ((!g2176) & (g2378) & (sk[76]) & (g522)) + ((g2176) & (!g2378) & (!sk[76]) & (g522)) + ((g2176) & (g2378) & (!sk[76]) & (!g522)) + ((g2176) & (g2378) & (!sk[76]) & (g522)) + ((g2176) & (g2378) & (sk[76]) & (!g522)) + ((g2176) & (g2378) & (sk[76]) & (g522)));
	assign g523 = (((!g519) & (!g520) & (!g521) & (g522) & (g165) & (g166)) + ((!g519) & (!g520) & (g521) & (!g522) & (!g165) & (g166)) + ((!g519) & (!g520) & (g521) & (g522) & (!g165) & (g166)) + ((!g519) & (!g520) & (g521) & (g522) & (g165) & (g166)) + ((!g519) & (g520) & (!g521) & (!g522) & (g165) & (!g166)) + ((!g519) & (g520) & (!g521) & (g522) & (g165) & (!g166)) + ((!g519) & (g520) & (!g521) & (g522) & (g165) & (g166)) + ((!g519) & (g520) & (g521) & (!g522) & (!g165) & (g166)) + ((!g519) & (g520) & (g521) & (!g522) & (g165) & (!g166)) + ((!g519) & (g520) & (g521) & (g522) & (!g165) & (g166)) + ((!g519) & (g520) & (g521) & (g522) & (g165) & (!g166)) + ((!g519) & (g520) & (g521) & (g522) & (g165) & (g166)) + ((g519) & (!g520) & (!g521) & (!g522) & (!g165) & (!g166)) + ((g519) & (!g520) & (!g521) & (g522) & (!g165) & (!g166)) + ((g519) & (!g520) & (!g521) & (g522) & (g165) & (g166)) + ((g519) & (!g520) & (g521) & (!g522) & (!g165) & (!g166)) + ((g519) & (!g520) & (g521) & (!g522) & (!g165) & (g166)) + ((g519) & (!g520) & (g521) & (g522) & (!g165) & (!g166)) + ((g519) & (!g520) & (g521) & (g522) & (!g165) & (g166)) + ((g519) & (!g520) & (g521) & (g522) & (g165) & (g166)) + ((g519) & (g520) & (!g521) & (!g522) & (!g165) & (!g166)) + ((g519) & (g520) & (!g521) & (!g522) & (g165) & (!g166)) + ((g519) & (g520) & (!g521) & (g522) & (!g165) & (!g166)) + ((g519) & (g520) & (!g521) & (g522) & (g165) & (!g166)) + ((g519) & (g520) & (!g521) & (g522) & (g165) & (g166)) + ((g519) & (g520) & (g521) & (!g522) & (!g165) & (!g166)) + ((g519) & (g520) & (g521) & (!g522) & (!g165) & (g166)) + ((g519) & (g520) & (g521) & (!g522) & (g165) & (!g166)) + ((g519) & (g520) & (g521) & (g522) & (!g165) & (!g166)) + ((g519) & (g520) & (g521) & (g522) & (!g165) & (g166)) + ((g519) & (g520) & (g521) & (g522) & (g165) & (!g166)) + ((g519) & (g520) & (g521) & (g522) & (g165) & (g166)));
	assign g4264 = (((!g2177) & (!g2378) & (!sk[78]) & (g524)) + ((!g2177) & (!g2378) & (sk[78]) & (g524)) + ((!g2177) & (g2378) & (!sk[78]) & (!g524)) + ((!g2177) & (g2378) & (!sk[78]) & (g524)) + ((!g2177) & (g2378) & (sk[78]) & (g524)) + ((g2177) & (!g2378) & (!sk[78]) & (g524)) + ((g2177) & (g2378) & (!sk[78]) & (!g524)) + ((g2177) & (g2378) & (!sk[78]) & (g524)) + ((g2177) & (g2378) & (sk[78]) & (!g524)) + ((g2177) & (g2378) & (sk[78]) & (g524)));
	assign g4265 = (((!g2178) & (!g2378) & (!sk[79]) & (g525)) + ((!g2178) & (!g2378) & (sk[79]) & (g525)) + ((!g2178) & (g2378) & (!sk[79]) & (!g525)) + ((!g2178) & (g2378) & (!sk[79]) & (g525)) + ((!g2178) & (g2378) & (sk[79]) & (g525)) + ((g2178) & (!g2378) & (!sk[79]) & (g525)) + ((g2178) & (g2378) & (!sk[79]) & (!g525)) + ((g2178) & (g2378) & (!sk[79]) & (g525)) + ((g2178) & (g2378) & (sk[79]) & (!g525)) + ((g2178) & (g2378) & (sk[79]) & (g525)));
	assign g4266 = (((!g2179) & (!sk[80]) & (!g2378) & (g526)) + ((!g2179) & (!sk[80]) & (g2378) & (!g526)) + ((!g2179) & (!sk[80]) & (g2378) & (g526)) + ((!g2179) & (sk[80]) & (!g2378) & (g526)) + ((!g2179) & (sk[80]) & (g2378) & (g526)) + ((g2179) & (!sk[80]) & (!g2378) & (g526)) + ((g2179) & (!sk[80]) & (g2378) & (!g526)) + ((g2179) & (!sk[80]) & (g2378) & (g526)) + ((g2179) & (sk[80]) & (g2378) & (!g526)) + ((g2179) & (sk[80]) & (g2378) & (g526)));
	assign g527 = (((!g165) & (!sk[81]) & (!g166) & (!g524) & (g525) & (!g526)) + ((!g165) & (!sk[81]) & (!g166) & (!g524) & (g525) & (g526)) + ((!g165) & (!sk[81]) & (!g166) & (g524) & (!g525) & (!g526)) + ((!g165) & (!sk[81]) & (!g166) & (g524) & (!g525) & (g526)) + ((!g165) & (!sk[81]) & (!g166) & (g524) & (g525) & (!g526)) + ((!g165) & (!sk[81]) & (!g166) & (g524) & (g525) & (g526)) + ((!g165) & (!sk[81]) & (g166) & (!g524) & (!g525) & (!g526)) + ((!g165) & (!sk[81]) & (g166) & (!g524) & (!g525) & (g526)) + ((!g165) & (!sk[81]) & (g166) & (!g524) & (g525) & (!g526)) + ((!g165) & (!sk[81]) & (g166) & (!g524) & (g525) & (g526)) + ((!g165) & (!sk[81]) & (g166) & (g524) & (!g525) & (!g526)) + ((!g165) & (!sk[81]) & (g166) & (g524) & (!g525) & (g526)) + ((!g165) & (!sk[81]) & (g166) & (g524) & (g525) & (!g526)) + ((!g165) & (!sk[81]) & (g166) & (g524) & (g525) & (g526)) + ((!g165) & (sk[81]) & (g166) & (!g524) & (!g525) & (g526)) + ((!g165) & (sk[81]) & (g166) & (!g524) & (g525) & (g526)) + ((!g165) & (sk[81]) & (g166) & (g524) & (!g525) & (g526)) + ((!g165) & (sk[81]) & (g166) & (g524) & (g525) & (g526)) + ((g165) & (!sk[81]) & (!g166) & (!g524) & (g525) & (!g526)) + ((g165) & (!sk[81]) & (!g166) & (!g524) & (g525) & (g526)) + ((g165) & (!sk[81]) & (!g166) & (g524) & (!g525) & (!g526)) + ((g165) & (!sk[81]) & (!g166) & (g524) & (!g525) & (g526)) + ((g165) & (!sk[81]) & (!g166) & (g524) & (g525) & (!g526)) + ((g165) & (!sk[81]) & (!g166) & (g524) & (g525) & (g526)) + ((g165) & (!sk[81]) & (g166) & (!g524) & (!g525) & (!g526)) + ((g165) & (!sk[81]) & (g166) & (!g524) & (!g525) & (g526)) + ((g165) & (!sk[81]) & (g166) & (!g524) & (g525) & (!g526)) + ((g165) & (!sk[81]) & (g166) & (!g524) & (g525) & (g526)) + ((g165) & (!sk[81]) & (g166) & (g524) & (!g525) & (!g526)) + ((g165) & (!sk[81]) & (g166) & (g524) & (!g525) & (g526)) + ((g165) & (!sk[81]) & (g166) & (g524) & (g525) & (!g526)) + ((g165) & (!sk[81]) & (g166) & (g524) & (g525) & (g526)) + ((g165) & (sk[81]) & (!g166) & (g524) & (!g525) & (!g526)) + ((g165) & (sk[81]) & (!g166) & (g524) & (!g525) & (g526)) + ((g165) & (sk[81]) & (!g166) & (g524) & (g525) & (!g526)) + ((g165) & (sk[81]) & (!g166) & (g524) & (g525) & (g526)) + ((g165) & (sk[81]) & (g166) & (!g524) & (g525) & (!g526)) + ((g165) & (sk[81]) & (g166) & (!g524) & (g525) & (g526)) + ((g165) & (sk[81]) & (g166) & (g524) & (g525) & (!g526)) + ((g165) & (sk[81]) & (g166) & (g524) & (g525) & (g526)));
	assign g4267 = (((!sk[82]) & (!g2162) & (!g2378) & (g528)) + ((!sk[82]) & (!g2162) & (g2378) & (!g528)) + ((!sk[82]) & (!g2162) & (g2378) & (g528)) + ((!sk[82]) & (g2162) & (!g2378) & (g528)) + ((!sk[82]) & (g2162) & (g2378) & (!g528)) + ((!sk[82]) & (g2162) & (g2378) & (g528)) + ((sk[82]) & (!g2162) & (!g2378) & (g528)) + ((sk[82]) & (!g2162) & (g2378) & (g528)) + ((sk[82]) & (g2162) & (g2378) & (!g528)) + ((sk[82]) & (g2162) & (g2378) & (g528)));
	assign g4268 = (((!g2164) & (!g2378) & (!sk[83]) & (g529)) + ((!g2164) & (!g2378) & (sk[83]) & (g529)) + ((!g2164) & (g2378) & (!sk[83]) & (!g529)) + ((!g2164) & (g2378) & (!sk[83]) & (g529)) + ((!g2164) & (g2378) & (sk[83]) & (g529)) + ((g2164) & (!g2378) & (!sk[83]) & (g529)) + ((g2164) & (g2378) & (!sk[83]) & (!g529)) + ((g2164) & (g2378) & (!sk[83]) & (g529)) + ((g2164) & (g2378) & (sk[83]) & (!g529)) + ((g2164) & (g2378) & (sk[83]) & (g529)));
	assign g4269 = (((!g2166) & (!sk[84]) & (!g2378) & (g530)) + ((!g2166) & (!sk[84]) & (g2378) & (!g530)) + ((!g2166) & (!sk[84]) & (g2378) & (g530)) + ((!g2166) & (sk[84]) & (!g2378) & (g530)) + ((!g2166) & (sk[84]) & (g2378) & (g530)) + ((g2166) & (!sk[84]) & (!g2378) & (g530)) + ((g2166) & (!sk[84]) & (g2378) & (!g530)) + ((g2166) & (!sk[84]) & (g2378) & (g530)) + ((g2166) & (sk[84]) & (g2378) & (!g530)) + ((g2166) & (sk[84]) & (g2378) & (g530)));
	assign g4270 = (((!sk[85]) & (!g2168) & (!g2378) & (g531)) + ((!sk[85]) & (!g2168) & (g2378) & (!g531)) + ((!sk[85]) & (!g2168) & (g2378) & (g531)) + ((!sk[85]) & (g2168) & (!g2378) & (g531)) + ((!sk[85]) & (g2168) & (g2378) & (!g531)) + ((!sk[85]) & (g2168) & (g2378) & (g531)) + ((sk[85]) & (!g2168) & (!g2378) & (g531)) + ((sk[85]) & (!g2168) & (g2378) & (g531)) + ((sk[85]) & (g2168) & (g2378) & (!g531)) + ((sk[85]) & (g2168) & (g2378) & (g531)));
	assign g532 = (((!g528) & (!g529) & (!g530) & (g531) & (g165) & (g166)) + ((!g528) & (!g529) & (g530) & (!g531) & (!g165) & (g166)) + ((!g528) & (!g529) & (g530) & (g531) & (!g165) & (g166)) + ((!g528) & (!g529) & (g530) & (g531) & (g165) & (g166)) + ((!g528) & (g529) & (!g530) & (!g531) & (g165) & (!g166)) + ((!g528) & (g529) & (!g530) & (g531) & (g165) & (!g166)) + ((!g528) & (g529) & (!g530) & (g531) & (g165) & (g166)) + ((!g528) & (g529) & (g530) & (!g531) & (!g165) & (g166)) + ((!g528) & (g529) & (g530) & (!g531) & (g165) & (!g166)) + ((!g528) & (g529) & (g530) & (g531) & (!g165) & (g166)) + ((!g528) & (g529) & (g530) & (g531) & (g165) & (!g166)) + ((!g528) & (g529) & (g530) & (g531) & (g165) & (g166)) + ((g528) & (!g529) & (!g530) & (!g531) & (!g165) & (!g166)) + ((g528) & (!g529) & (!g530) & (g531) & (!g165) & (!g166)) + ((g528) & (!g529) & (!g530) & (g531) & (g165) & (g166)) + ((g528) & (!g529) & (g530) & (!g531) & (!g165) & (!g166)) + ((g528) & (!g529) & (g530) & (!g531) & (!g165) & (g166)) + ((g528) & (!g529) & (g530) & (g531) & (!g165) & (!g166)) + ((g528) & (!g529) & (g530) & (g531) & (!g165) & (g166)) + ((g528) & (!g529) & (g530) & (g531) & (g165) & (g166)) + ((g528) & (g529) & (!g530) & (!g531) & (!g165) & (!g166)) + ((g528) & (g529) & (!g530) & (!g531) & (g165) & (!g166)) + ((g528) & (g529) & (!g530) & (g531) & (!g165) & (!g166)) + ((g528) & (g529) & (!g530) & (g531) & (g165) & (!g166)) + ((g528) & (g529) & (!g530) & (g531) & (g165) & (g166)) + ((g528) & (g529) & (g530) & (!g531) & (!g165) & (!g166)) + ((g528) & (g529) & (g530) & (!g531) & (!g165) & (g166)) + ((g528) & (g529) & (g530) & (!g531) & (g165) & (!g166)) + ((g528) & (g529) & (g530) & (g531) & (!g165) & (!g166)) + ((g528) & (g529) & (g530) & (g531) & (!g165) & (g166)) + ((g528) & (g529) & (g530) & (g531) & (g165) & (!g166)) + ((g528) & (g529) & (g530) & (g531) & (g165) & (g166)));
	assign g4271 = (((!sk[87]) & (!g2169) & (!g2378) & (g533)) + ((!sk[87]) & (!g2169) & (g2378) & (!g533)) + ((!sk[87]) & (!g2169) & (g2378) & (g533)) + ((!sk[87]) & (g2169) & (!g2378) & (g533)) + ((!sk[87]) & (g2169) & (g2378) & (!g533)) + ((!sk[87]) & (g2169) & (g2378) & (g533)) + ((sk[87]) & (!g2169) & (!g2378) & (g533)) + ((sk[87]) & (!g2169) & (g2378) & (g533)) + ((sk[87]) & (g2169) & (g2378) & (!g533)) + ((sk[87]) & (g2169) & (g2378) & (g533)));
	assign g4272 = (((!g2170) & (!g2378) & (!sk[88]) & (g534)) + ((!g2170) & (!g2378) & (sk[88]) & (g534)) + ((!g2170) & (g2378) & (!sk[88]) & (!g534)) + ((!g2170) & (g2378) & (!sk[88]) & (g534)) + ((!g2170) & (g2378) & (sk[88]) & (g534)) + ((g2170) & (!g2378) & (!sk[88]) & (g534)) + ((g2170) & (g2378) & (!sk[88]) & (!g534)) + ((g2170) & (g2378) & (!sk[88]) & (g534)) + ((g2170) & (g2378) & (sk[88]) & (!g534)) + ((g2170) & (g2378) & (sk[88]) & (g534)));
	assign g4273 = (((!sk[89]) & (!g2171) & (!g2378) & (g535)) + ((!sk[89]) & (!g2171) & (g2378) & (!g535)) + ((!sk[89]) & (!g2171) & (g2378) & (g535)) + ((!sk[89]) & (g2171) & (!g2378) & (g535)) + ((!sk[89]) & (g2171) & (g2378) & (!g535)) + ((!sk[89]) & (g2171) & (g2378) & (g535)) + ((sk[89]) & (!g2171) & (!g2378) & (g535)) + ((sk[89]) & (!g2171) & (g2378) & (g535)) + ((sk[89]) & (g2171) & (g2378) & (!g535)) + ((sk[89]) & (g2171) & (g2378) & (g535)));
	assign g4274 = (((!g2172) & (!g2378) & (!sk[90]) & (g536)) + ((!g2172) & (!g2378) & (sk[90]) & (g536)) + ((!g2172) & (g2378) & (!sk[90]) & (!g536)) + ((!g2172) & (g2378) & (!sk[90]) & (g536)) + ((!g2172) & (g2378) & (sk[90]) & (g536)) + ((g2172) & (!g2378) & (!sk[90]) & (g536)) + ((g2172) & (g2378) & (!sk[90]) & (!g536)) + ((g2172) & (g2378) & (!sk[90]) & (g536)) + ((g2172) & (g2378) & (sk[90]) & (!g536)) + ((g2172) & (g2378) & (sk[90]) & (g536)));
	assign g537 = (((!g533) & (!g534) & (!g535) & (g536) & (g165) & (g166)) + ((!g533) & (!g534) & (g535) & (!g536) & (!g165) & (g166)) + ((!g533) & (!g534) & (g535) & (g536) & (!g165) & (g166)) + ((!g533) & (!g534) & (g535) & (g536) & (g165) & (g166)) + ((!g533) & (g534) & (!g535) & (!g536) & (g165) & (!g166)) + ((!g533) & (g534) & (!g535) & (g536) & (g165) & (!g166)) + ((!g533) & (g534) & (!g535) & (g536) & (g165) & (g166)) + ((!g533) & (g534) & (g535) & (!g536) & (!g165) & (g166)) + ((!g533) & (g534) & (g535) & (!g536) & (g165) & (!g166)) + ((!g533) & (g534) & (g535) & (g536) & (!g165) & (g166)) + ((!g533) & (g534) & (g535) & (g536) & (g165) & (!g166)) + ((!g533) & (g534) & (g535) & (g536) & (g165) & (g166)) + ((g533) & (!g534) & (!g535) & (!g536) & (!g165) & (!g166)) + ((g533) & (!g534) & (!g535) & (g536) & (!g165) & (!g166)) + ((g533) & (!g534) & (!g535) & (g536) & (g165) & (g166)) + ((g533) & (!g534) & (g535) & (!g536) & (!g165) & (!g166)) + ((g533) & (!g534) & (g535) & (!g536) & (!g165) & (g166)) + ((g533) & (!g534) & (g535) & (g536) & (!g165) & (!g166)) + ((g533) & (!g534) & (g535) & (g536) & (!g165) & (g166)) + ((g533) & (!g534) & (g535) & (g536) & (g165) & (g166)) + ((g533) & (g534) & (!g535) & (!g536) & (!g165) & (!g166)) + ((g533) & (g534) & (!g535) & (!g536) & (g165) & (!g166)) + ((g533) & (g534) & (!g535) & (g536) & (!g165) & (!g166)) + ((g533) & (g534) & (!g535) & (g536) & (g165) & (!g166)) + ((g533) & (g534) & (!g535) & (g536) & (g165) & (g166)) + ((g533) & (g534) & (g535) & (!g536) & (!g165) & (!g166)) + ((g533) & (g534) & (g535) & (!g536) & (!g165) & (g166)) + ((g533) & (g534) & (g535) & (!g536) & (g165) & (!g166)) + ((g533) & (g534) & (g535) & (g536) & (!g165) & (!g166)) + ((g533) & (g534) & (g535) & (g536) & (!g165) & (g166)) + ((g533) & (g534) & (g535) & (g536) & (g165) & (!g166)) + ((g533) & (g534) & (g535) & (g536) & (g165) & (g166)));
	assign g538 = (((!g147) & (!g148) & (!g523) & (g527) & (!g532) & (!g537)) + ((!g147) & (!g148) & (!g523) & (g527) & (!g532) & (g537)) + ((!g147) & (!g148) & (!g523) & (g527) & (g532) & (!g537)) + ((!g147) & (!g148) & (!g523) & (g527) & (g532) & (g537)) + ((!g147) & (!g148) & (g523) & (g527) & (!g532) & (!g537)) + ((!g147) & (!g148) & (g523) & (g527) & (!g532) & (g537)) + ((!g147) & (!g148) & (g523) & (g527) & (g532) & (!g537)) + ((!g147) & (!g148) & (g523) & (g527) & (g532) & (g537)) + ((!g147) & (g148) & (!g523) & (!g527) & (!g532) & (g537)) + ((!g147) & (g148) & (!g523) & (!g527) & (g532) & (g537)) + ((!g147) & (g148) & (!g523) & (g527) & (!g532) & (g537)) + ((!g147) & (g148) & (!g523) & (g527) & (g532) & (g537)) + ((!g147) & (g148) & (g523) & (!g527) & (!g532) & (g537)) + ((!g147) & (g148) & (g523) & (!g527) & (g532) & (g537)) + ((!g147) & (g148) & (g523) & (g527) & (!g532) & (g537)) + ((!g147) & (g148) & (g523) & (g527) & (g532) & (g537)) + ((g147) & (!g148) & (g523) & (!g527) & (!g532) & (!g537)) + ((g147) & (!g148) & (g523) & (!g527) & (!g532) & (g537)) + ((g147) & (!g148) & (g523) & (!g527) & (g532) & (!g537)) + ((g147) & (!g148) & (g523) & (!g527) & (g532) & (g537)) + ((g147) & (!g148) & (g523) & (g527) & (!g532) & (!g537)) + ((g147) & (!g148) & (g523) & (g527) & (!g532) & (g537)) + ((g147) & (!g148) & (g523) & (g527) & (g532) & (!g537)) + ((g147) & (!g148) & (g523) & (g527) & (g532) & (g537)) + ((g147) & (g148) & (!g523) & (!g527) & (g532) & (!g537)) + ((g147) & (g148) & (!g523) & (!g527) & (g532) & (g537)) + ((g147) & (g148) & (!g523) & (g527) & (g532) & (!g537)) + ((g147) & (g148) & (!g523) & (g527) & (g532) & (g537)) + ((g147) & (g148) & (g523) & (!g527) & (g532) & (!g537)) + ((g147) & (g148) & (g523) & (!g527) & (g532) & (g537)) + ((g147) & (g148) & (g523) & (g527) & (g532) & (!g537)) + ((g147) & (g148) & (g523) & (g527) & (g532) & (g537)));
	assign g539 = (((!sk[93]) & (!g142) & (!g518) & (g538)) + ((!sk[93]) & (!g142) & (g518) & (!g538)) + ((!sk[93]) & (!g142) & (g518) & (g538)) + ((!sk[93]) & (g142) & (!g518) & (g538)) + ((!sk[93]) & (g142) & (g518) & (!g538)) + ((!sk[93]) & (g142) & (g518) & (g538)) + ((sk[93]) & (!g142) & (!g518) & (g538)) + ((sk[93]) & (!g142) & (g518) & (g538)) + ((sk[93]) & (g142) & (g518) & (!g538)) + ((sk[93]) & (g142) & (g518) & (g538)));
	assign g540 = (((!g92) & (!g126) & (!g496) & (!sk[94]) & (g497) & (!g539)) + ((!g92) & (!g126) & (!g496) & (!sk[94]) & (g497) & (g539)) + ((!g92) & (!g126) & (!g496) & (sk[94]) & (!g497) & (!g539)) + ((!g92) & (!g126) & (!g496) & (sk[94]) & (!g497) & (g539)) + ((!g92) & (!g126) & (!g496) & (sk[94]) & (g497) & (!g539)) + ((!g92) & (!g126) & (!g496) & (sk[94]) & (g497) & (g539)) + ((!g92) & (!g126) & (g496) & (!sk[94]) & (!g497) & (!g539)) + ((!g92) & (!g126) & (g496) & (!sk[94]) & (!g497) & (g539)) + ((!g92) & (!g126) & (g496) & (!sk[94]) & (g497) & (!g539)) + ((!g92) & (!g126) & (g496) & (!sk[94]) & (g497) & (g539)) + ((!g92) & (g126) & (!g496) & (!sk[94]) & (!g497) & (!g539)) + ((!g92) & (g126) & (!g496) & (!sk[94]) & (!g497) & (g539)) + ((!g92) & (g126) & (!g496) & (!sk[94]) & (g497) & (!g539)) + ((!g92) & (g126) & (!g496) & (!sk[94]) & (g497) & (g539)) + ((!g92) & (g126) & (!g496) & (sk[94]) & (!g497) & (g539)) + ((!g92) & (g126) & (!g496) & (sk[94]) & (g497) & (!g539)) + ((!g92) & (g126) & (g496) & (!sk[94]) & (!g497) & (!g539)) + ((!g92) & (g126) & (g496) & (!sk[94]) & (!g497) & (g539)) + ((!g92) & (g126) & (g496) & (!sk[94]) & (g497) & (!g539)) + ((!g92) & (g126) & (g496) & (!sk[94]) & (g497) & (g539)) + ((!g92) & (g126) & (g496) & (sk[94]) & (!g497) & (g539)) + ((!g92) & (g126) & (g496) & (sk[94]) & (g497) & (!g539)) + ((g92) & (!g126) & (!g496) & (!sk[94]) & (g497) & (!g539)) + ((g92) & (!g126) & (!g496) & (!sk[94]) & (g497) & (g539)) + ((g92) & (!g126) & (!g496) & (sk[94]) & (!g497) & (!g539)) + ((g92) & (!g126) & (!g496) & (sk[94]) & (!g497) & (g539)) + ((g92) & (!g126) & (!g496) & (sk[94]) & (g497) & (!g539)) + ((g92) & (!g126) & (!g496) & (sk[94]) & (g497) & (g539)) + ((g92) & (!g126) & (g496) & (!sk[94]) & (!g497) & (!g539)) + ((g92) & (!g126) & (g496) & (!sk[94]) & (!g497) & (g539)) + ((g92) & (!g126) & (g496) & (!sk[94]) & (g497) & (!g539)) + ((g92) & (!g126) & (g496) & (!sk[94]) & (g497) & (g539)) + ((g92) & (g126) & (!g496) & (!sk[94]) & (!g497) & (!g539)) + ((g92) & (g126) & (!g496) & (!sk[94]) & (!g497) & (g539)) + ((g92) & (g126) & (!g496) & (!sk[94]) & (g497) & (!g539)) + ((g92) & (g126) & (!g496) & (!sk[94]) & (g497) & (g539)) + ((g92) & (g126) & (!g496) & (sk[94]) & (!g497) & (!g539)) + ((g92) & (g126) & (!g496) & (sk[94]) & (g497) & (g539)) + ((g92) & (g126) & (g496) & (!sk[94]) & (!g497) & (!g539)) + ((g92) & (g126) & (g496) & (!sk[94]) & (!g497) & (g539)) + ((g92) & (g126) & (g496) & (!sk[94]) & (g497) & (!g539)) + ((g92) & (g126) & (g496) & (!sk[94]) & (g497) & (g539)) + ((g92) & (g126) & (g496) & (sk[94]) & (!g497) & (!g539)) + ((g92) & (g126) & (g496) & (sk[94]) & (g497) & (g539)));
	assign g4275 = (((!g2059) & (!sk[95]) & (!g2388) & (g541)) + ((!g2059) & (!sk[95]) & (g2388) & (!g541)) + ((!g2059) & (!sk[95]) & (g2388) & (g541)) + ((!g2059) & (sk[95]) & (!g2388) & (g541)) + ((!g2059) & (sk[95]) & (g2388) & (g541)) + ((g2059) & (!sk[95]) & (!g2388) & (g541)) + ((g2059) & (!sk[95]) & (g2388) & (!g541)) + ((g2059) & (!sk[95]) & (g2388) & (g541)) + ((g2059) & (sk[95]) & (g2388) & (!g541)) + ((g2059) & (sk[95]) & (g2388) & (g541)));
	assign g542 = (((!sk[96]) & (!g92) & (!g497) & (g539)) + ((!sk[96]) & (!g92) & (g497) & (!g539)) + ((!sk[96]) & (!g92) & (g497) & (g539)) + ((!sk[96]) & (g92) & (!g497) & (g539)) + ((!sk[96]) & (g92) & (g497) & (!g539)) + ((!sk[96]) & (g92) & (g497) & (g539)) + ((sk[96]) & (!g92) & (g497) & (g539)) + ((sk[96]) & (g92) & (!g497) & (g539)) + ((sk[96]) & (g92) & (g497) & (!g539)) + ((sk[96]) & (g92) & (g497) & (g539)));
	assign g4276 = (((!sk[97]) & (!g2140) & (!g2407) & (g543)) + ((!sk[97]) & (!g2140) & (g2407) & (!g543)) + ((!sk[97]) & (!g2140) & (g2407) & (g543)) + ((!sk[97]) & (g2140) & (!g2407) & (g543)) + ((!sk[97]) & (g2140) & (g2407) & (!g543)) + ((!sk[97]) & (g2140) & (g2407) & (g543)) + ((sk[97]) & (!g2140) & (!g2407) & (g543)) + ((sk[97]) & (!g2140) & (g2407) & (g543)) + ((sk[97]) & (g2140) & (g2407) & (!g543)) + ((sk[97]) & (g2140) & (g2407) & (g543)));
	assign g4277 = (((!sk[98]) & (!g2146) & (!g2407) & (g544)) + ((!sk[98]) & (!g2146) & (g2407) & (!g544)) + ((!sk[98]) & (!g2146) & (g2407) & (g544)) + ((!sk[98]) & (g2146) & (!g2407) & (g544)) + ((!sk[98]) & (g2146) & (g2407) & (!g544)) + ((!sk[98]) & (g2146) & (g2407) & (g544)) + ((sk[98]) & (!g2146) & (!g2407) & (g544)) + ((sk[98]) & (!g2146) & (g2407) & (g544)) + ((sk[98]) & (g2146) & (g2407) & (!g544)) + ((sk[98]) & (g2146) & (g2407) & (g544)));
	assign g4278 = (((!g2152) & (!g2407) & (!sk[99]) & (g545)) + ((!g2152) & (!g2407) & (sk[99]) & (g545)) + ((!g2152) & (g2407) & (!sk[99]) & (!g545)) + ((!g2152) & (g2407) & (!sk[99]) & (g545)) + ((!g2152) & (g2407) & (sk[99]) & (g545)) + ((g2152) & (!g2407) & (!sk[99]) & (g545)) + ((g2152) & (g2407) & (!sk[99]) & (!g545)) + ((g2152) & (g2407) & (!sk[99]) & (g545)) + ((g2152) & (g2407) & (sk[99]) & (!g545)) + ((g2152) & (g2407) & (sk[99]) & (g545)));
	assign g4279 = (((!sk[100]) & (!g2158) & (!g2407) & (g546)) + ((!sk[100]) & (!g2158) & (g2407) & (!g546)) + ((!sk[100]) & (!g2158) & (g2407) & (g546)) + ((!sk[100]) & (g2158) & (!g2407) & (g546)) + ((!sk[100]) & (g2158) & (g2407) & (!g546)) + ((!sk[100]) & (g2158) & (g2407) & (g546)) + ((sk[100]) & (!g2158) & (!g2407) & (g546)) + ((sk[100]) & (!g2158) & (g2407) & (g546)) + ((sk[100]) & (g2158) & (g2407) & (!g546)) + ((sk[100]) & (g2158) & (g2407) & (g546)));
	assign g547 = (((!g543) & (!g544) & (!g545) & (g546) & (g165) & (g166)) + ((!g543) & (!g544) & (g545) & (!g546) & (!g165) & (g166)) + ((!g543) & (!g544) & (g545) & (g546) & (!g165) & (g166)) + ((!g543) & (!g544) & (g545) & (g546) & (g165) & (g166)) + ((!g543) & (g544) & (!g545) & (!g546) & (g165) & (!g166)) + ((!g543) & (g544) & (!g545) & (g546) & (g165) & (!g166)) + ((!g543) & (g544) & (!g545) & (g546) & (g165) & (g166)) + ((!g543) & (g544) & (g545) & (!g546) & (!g165) & (g166)) + ((!g543) & (g544) & (g545) & (!g546) & (g165) & (!g166)) + ((!g543) & (g544) & (g545) & (g546) & (!g165) & (g166)) + ((!g543) & (g544) & (g545) & (g546) & (g165) & (!g166)) + ((!g543) & (g544) & (g545) & (g546) & (g165) & (g166)) + ((g543) & (!g544) & (!g545) & (!g546) & (!g165) & (!g166)) + ((g543) & (!g544) & (!g545) & (g546) & (!g165) & (!g166)) + ((g543) & (!g544) & (!g545) & (g546) & (g165) & (g166)) + ((g543) & (!g544) & (g545) & (!g546) & (!g165) & (!g166)) + ((g543) & (!g544) & (g545) & (!g546) & (!g165) & (g166)) + ((g543) & (!g544) & (g545) & (g546) & (!g165) & (!g166)) + ((g543) & (!g544) & (g545) & (g546) & (!g165) & (g166)) + ((g543) & (!g544) & (g545) & (g546) & (g165) & (g166)) + ((g543) & (g544) & (!g545) & (!g546) & (!g165) & (!g166)) + ((g543) & (g544) & (!g545) & (!g546) & (g165) & (!g166)) + ((g543) & (g544) & (!g545) & (g546) & (!g165) & (!g166)) + ((g543) & (g544) & (!g545) & (g546) & (g165) & (!g166)) + ((g543) & (g544) & (!g545) & (g546) & (g165) & (g166)) + ((g543) & (g544) & (g545) & (!g546) & (!g165) & (!g166)) + ((g543) & (g544) & (g545) & (!g546) & (!g165) & (g166)) + ((g543) & (g544) & (g545) & (!g546) & (g165) & (!g166)) + ((g543) & (g544) & (g545) & (g546) & (!g165) & (!g166)) + ((g543) & (g544) & (g545) & (g546) & (!g165) & (g166)) + ((g543) & (g544) & (g545) & (g546) & (g165) & (!g166)) + ((g543) & (g544) & (g545) & (g546) & (g165) & (g166)));
	assign g4280 = (((!g2142) & (!sk[102]) & (!g2407) & (g548)) + ((!g2142) & (!sk[102]) & (g2407) & (!g548)) + ((!g2142) & (!sk[102]) & (g2407) & (g548)) + ((!g2142) & (sk[102]) & (!g2407) & (g548)) + ((!g2142) & (sk[102]) & (g2407) & (g548)) + ((g2142) & (!sk[102]) & (!g2407) & (g548)) + ((g2142) & (!sk[102]) & (g2407) & (!g548)) + ((g2142) & (!sk[102]) & (g2407) & (g548)) + ((g2142) & (sk[102]) & (g2407) & (!g548)) + ((g2142) & (sk[102]) & (g2407) & (g548)));
	assign g4281 = (((!g2148) & (!sk[103]) & (!g2407) & (g549)) + ((!g2148) & (!sk[103]) & (g2407) & (!g549)) + ((!g2148) & (!sk[103]) & (g2407) & (g549)) + ((!g2148) & (sk[103]) & (!g2407) & (g549)) + ((!g2148) & (sk[103]) & (g2407) & (g549)) + ((g2148) & (!sk[103]) & (!g2407) & (g549)) + ((g2148) & (!sk[103]) & (g2407) & (!g549)) + ((g2148) & (!sk[103]) & (g2407) & (g549)) + ((g2148) & (sk[103]) & (g2407) & (!g549)) + ((g2148) & (sk[103]) & (g2407) & (g549)));
	assign g4282 = (((!g2153) & (!sk[104]) & (!g2407) & (g550)) + ((!g2153) & (!sk[104]) & (g2407) & (!g550)) + ((!g2153) & (!sk[104]) & (g2407) & (g550)) + ((!g2153) & (sk[104]) & (!g2407) & (g550)) + ((!g2153) & (sk[104]) & (g2407) & (g550)) + ((g2153) & (!sk[104]) & (!g2407) & (g550)) + ((g2153) & (!sk[104]) & (g2407) & (!g550)) + ((g2153) & (!sk[104]) & (g2407) & (g550)) + ((g2153) & (sk[104]) & (g2407) & (!g550)) + ((g2153) & (sk[104]) & (g2407) & (g550)));
	assign g4283 = (((!g2159) & (!g2407) & (!sk[105]) & (g551)) + ((!g2159) & (!g2407) & (sk[105]) & (g551)) + ((!g2159) & (g2407) & (!sk[105]) & (!g551)) + ((!g2159) & (g2407) & (!sk[105]) & (g551)) + ((!g2159) & (g2407) & (sk[105]) & (g551)) + ((g2159) & (!g2407) & (!sk[105]) & (g551)) + ((g2159) & (g2407) & (!sk[105]) & (!g551)) + ((g2159) & (g2407) & (!sk[105]) & (g551)) + ((g2159) & (g2407) & (sk[105]) & (!g551)) + ((g2159) & (g2407) & (sk[105]) & (g551)));
	assign g552 = (((!g548) & (!g549) & (!g550) & (g551) & (g165) & (g166)) + ((!g548) & (!g549) & (g550) & (!g551) & (!g165) & (g166)) + ((!g548) & (!g549) & (g550) & (g551) & (!g165) & (g166)) + ((!g548) & (!g549) & (g550) & (g551) & (g165) & (g166)) + ((!g548) & (g549) & (!g550) & (!g551) & (g165) & (!g166)) + ((!g548) & (g549) & (!g550) & (g551) & (g165) & (!g166)) + ((!g548) & (g549) & (!g550) & (g551) & (g165) & (g166)) + ((!g548) & (g549) & (g550) & (!g551) & (!g165) & (g166)) + ((!g548) & (g549) & (g550) & (!g551) & (g165) & (!g166)) + ((!g548) & (g549) & (g550) & (g551) & (!g165) & (g166)) + ((!g548) & (g549) & (g550) & (g551) & (g165) & (!g166)) + ((!g548) & (g549) & (g550) & (g551) & (g165) & (g166)) + ((g548) & (!g549) & (!g550) & (!g551) & (!g165) & (!g166)) + ((g548) & (!g549) & (!g550) & (g551) & (!g165) & (!g166)) + ((g548) & (!g549) & (!g550) & (g551) & (g165) & (g166)) + ((g548) & (!g549) & (g550) & (!g551) & (!g165) & (!g166)) + ((g548) & (!g549) & (g550) & (!g551) & (!g165) & (g166)) + ((g548) & (!g549) & (g550) & (g551) & (!g165) & (!g166)) + ((g548) & (!g549) & (g550) & (g551) & (!g165) & (g166)) + ((g548) & (!g549) & (g550) & (g551) & (g165) & (g166)) + ((g548) & (g549) & (!g550) & (!g551) & (!g165) & (!g166)) + ((g548) & (g549) & (!g550) & (!g551) & (g165) & (!g166)) + ((g548) & (g549) & (!g550) & (g551) & (!g165) & (!g166)) + ((g548) & (g549) & (!g550) & (g551) & (g165) & (!g166)) + ((g548) & (g549) & (!g550) & (g551) & (g165) & (g166)) + ((g548) & (g549) & (g550) & (!g551) & (!g165) & (!g166)) + ((g548) & (g549) & (g550) & (!g551) & (!g165) & (g166)) + ((g548) & (g549) & (g550) & (!g551) & (g165) & (!g166)) + ((g548) & (g549) & (g550) & (g551) & (!g165) & (!g166)) + ((g548) & (g549) & (g550) & (g551) & (!g165) & (g166)) + ((g548) & (g549) & (g550) & (g551) & (g165) & (!g166)) + ((g548) & (g549) & (g550) & (g551) & (g165) & (g166)));
	assign g4284 = (((!sk[107]) & (!g2144) & (!g2407) & (g553)) + ((!sk[107]) & (!g2144) & (g2407) & (!g553)) + ((!sk[107]) & (!g2144) & (g2407) & (g553)) + ((!sk[107]) & (g2144) & (!g2407) & (g553)) + ((!sk[107]) & (g2144) & (g2407) & (!g553)) + ((!sk[107]) & (g2144) & (g2407) & (g553)) + ((sk[107]) & (!g2144) & (!g2407) & (g553)) + ((sk[107]) & (!g2144) & (g2407) & (g553)) + ((sk[107]) & (g2144) & (g2407) & (!g553)) + ((sk[107]) & (g2144) & (g2407) & (g553)));
	assign g4285 = (((!g2150) & (!sk[108]) & (!g2407) & (g554)) + ((!g2150) & (!sk[108]) & (g2407) & (!g554)) + ((!g2150) & (!sk[108]) & (g2407) & (g554)) + ((!g2150) & (sk[108]) & (!g2407) & (g554)) + ((!g2150) & (sk[108]) & (g2407) & (g554)) + ((g2150) & (!sk[108]) & (!g2407) & (g554)) + ((g2150) & (!sk[108]) & (g2407) & (!g554)) + ((g2150) & (!sk[108]) & (g2407) & (g554)) + ((g2150) & (sk[108]) & (g2407) & (!g554)) + ((g2150) & (sk[108]) & (g2407) & (g554)));
	assign g4286 = (((!sk[109]) & (!g2155) & (!g2407) & (g555)) + ((!sk[109]) & (!g2155) & (g2407) & (!g555)) + ((!sk[109]) & (!g2155) & (g2407) & (g555)) + ((!sk[109]) & (g2155) & (!g2407) & (g555)) + ((!sk[109]) & (g2155) & (g2407) & (!g555)) + ((!sk[109]) & (g2155) & (g2407) & (g555)) + ((sk[109]) & (!g2155) & (!g2407) & (g555)) + ((sk[109]) & (!g2155) & (g2407) & (g555)) + ((sk[109]) & (g2155) & (g2407) & (!g555)) + ((sk[109]) & (g2155) & (g2407) & (g555)));
	assign g4287 = (((!g2160) & (!g2407) & (!sk[110]) & (g556)) + ((!g2160) & (!g2407) & (sk[110]) & (g556)) + ((!g2160) & (g2407) & (!sk[110]) & (!g556)) + ((!g2160) & (g2407) & (!sk[110]) & (g556)) + ((!g2160) & (g2407) & (sk[110]) & (g556)) + ((g2160) & (!g2407) & (!sk[110]) & (g556)) + ((g2160) & (g2407) & (!sk[110]) & (!g556)) + ((g2160) & (g2407) & (!sk[110]) & (g556)) + ((g2160) & (g2407) & (sk[110]) & (!g556)) + ((g2160) & (g2407) & (sk[110]) & (g556)));
	assign g557 = (((!g553) & (!g554) & (!g555) & (g556) & (g165) & (g166)) + ((!g553) & (!g554) & (g555) & (!g556) & (!g165) & (g166)) + ((!g553) & (!g554) & (g555) & (g556) & (!g165) & (g166)) + ((!g553) & (!g554) & (g555) & (g556) & (g165) & (g166)) + ((!g553) & (g554) & (!g555) & (!g556) & (g165) & (!g166)) + ((!g553) & (g554) & (!g555) & (g556) & (g165) & (!g166)) + ((!g553) & (g554) & (!g555) & (g556) & (g165) & (g166)) + ((!g553) & (g554) & (g555) & (!g556) & (!g165) & (g166)) + ((!g553) & (g554) & (g555) & (!g556) & (g165) & (!g166)) + ((!g553) & (g554) & (g555) & (g556) & (!g165) & (g166)) + ((!g553) & (g554) & (g555) & (g556) & (g165) & (!g166)) + ((!g553) & (g554) & (g555) & (g556) & (g165) & (g166)) + ((g553) & (!g554) & (!g555) & (!g556) & (!g165) & (!g166)) + ((g553) & (!g554) & (!g555) & (g556) & (!g165) & (!g166)) + ((g553) & (!g554) & (!g555) & (g556) & (g165) & (g166)) + ((g553) & (!g554) & (g555) & (!g556) & (!g165) & (!g166)) + ((g553) & (!g554) & (g555) & (!g556) & (!g165) & (g166)) + ((g553) & (!g554) & (g555) & (g556) & (!g165) & (!g166)) + ((g553) & (!g554) & (g555) & (g556) & (!g165) & (g166)) + ((g553) & (!g554) & (g555) & (g556) & (g165) & (g166)) + ((g553) & (g554) & (!g555) & (!g556) & (!g165) & (!g166)) + ((g553) & (g554) & (!g555) & (!g556) & (g165) & (!g166)) + ((g553) & (g554) & (!g555) & (g556) & (!g165) & (!g166)) + ((g553) & (g554) & (!g555) & (g556) & (g165) & (!g166)) + ((g553) & (g554) & (!g555) & (g556) & (g165) & (g166)) + ((g553) & (g554) & (g555) & (!g556) & (!g165) & (!g166)) + ((g553) & (g554) & (g555) & (!g556) & (!g165) & (g166)) + ((g553) & (g554) & (g555) & (!g556) & (g165) & (!g166)) + ((g553) & (g554) & (g555) & (g556) & (!g165) & (!g166)) + ((g553) & (g554) & (g555) & (g556) & (!g165) & (g166)) + ((g553) & (g554) & (g555) & (g556) & (g165) & (!g166)) + ((g553) & (g554) & (g555) & (g556) & (g165) & (g166)));
	assign g4288 = (((!g2145) & (!g2407) & (!sk[112]) & (g558)) + ((!g2145) & (!g2407) & (sk[112]) & (g558)) + ((!g2145) & (g2407) & (!sk[112]) & (!g558)) + ((!g2145) & (g2407) & (!sk[112]) & (g558)) + ((!g2145) & (g2407) & (sk[112]) & (g558)) + ((g2145) & (!g2407) & (!sk[112]) & (g558)) + ((g2145) & (g2407) & (!sk[112]) & (!g558)) + ((g2145) & (g2407) & (!sk[112]) & (g558)) + ((g2145) & (g2407) & (sk[112]) & (!g558)) + ((g2145) & (g2407) & (sk[112]) & (g558)));
	assign g4289 = (((!g2151) & (!g2407) & (!sk[113]) & (g559)) + ((!g2151) & (!g2407) & (sk[113]) & (g559)) + ((!g2151) & (g2407) & (!sk[113]) & (!g559)) + ((!g2151) & (g2407) & (!sk[113]) & (g559)) + ((!g2151) & (g2407) & (sk[113]) & (g559)) + ((g2151) & (!g2407) & (!sk[113]) & (g559)) + ((g2151) & (g2407) & (!sk[113]) & (!g559)) + ((g2151) & (g2407) & (!sk[113]) & (g559)) + ((g2151) & (g2407) & (sk[113]) & (!g559)) + ((g2151) & (g2407) & (sk[113]) & (g559)));
	assign g4290 = (((!g2157) & (!g2407) & (!sk[114]) & (g560)) + ((!g2157) & (!g2407) & (sk[114]) & (g560)) + ((!g2157) & (g2407) & (!sk[114]) & (!g560)) + ((!g2157) & (g2407) & (!sk[114]) & (g560)) + ((!g2157) & (g2407) & (sk[114]) & (g560)) + ((g2157) & (!g2407) & (!sk[114]) & (g560)) + ((g2157) & (g2407) & (!sk[114]) & (!g560)) + ((g2157) & (g2407) & (!sk[114]) & (g560)) + ((g2157) & (g2407) & (sk[114]) & (!g560)) + ((g2157) & (g2407) & (sk[114]) & (g560)));
	assign g4291 = (((!g2161) & (!g2407) & (!sk[115]) & (g561)) + ((!g2161) & (!g2407) & (sk[115]) & (g561)) + ((!g2161) & (g2407) & (!sk[115]) & (!g561)) + ((!g2161) & (g2407) & (!sk[115]) & (g561)) + ((!g2161) & (g2407) & (sk[115]) & (g561)) + ((g2161) & (!g2407) & (!sk[115]) & (g561)) + ((g2161) & (g2407) & (!sk[115]) & (!g561)) + ((g2161) & (g2407) & (!sk[115]) & (g561)) + ((g2161) & (g2407) & (sk[115]) & (!g561)) + ((g2161) & (g2407) & (sk[115]) & (g561)));
	assign g562 = (((!g558) & (!g559) & (!g560) & (g561) & (g165) & (g166)) + ((!g558) & (!g559) & (g560) & (!g561) & (!g165) & (g166)) + ((!g558) & (!g559) & (g560) & (g561) & (!g165) & (g166)) + ((!g558) & (!g559) & (g560) & (g561) & (g165) & (g166)) + ((!g558) & (g559) & (!g560) & (!g561) & (g165) & (!g166)) + ((!g558) & (g559) & (!g560) & (g561) & (g165) & (!g166)) + ((!g558) & (g559) & (!g560) & (g561) & (g165) & (g166)) + ((!g558) & (g559) & (g560) & (!g561) & (!g165) & (g166)) + ((!g558) & (g559) & (g560) & (!g561) & (g165) & (!g166)) + ((!g558) & (g559) & (g560) & (g561) & (!g165) & (g166)) + ((!g558) & (g559) & (g560) & (g561) & (g165) & (!g166)) + ((!g558) & (g559) & (g560) & (g561) & (g165) & (g166)) + ((g558) & (!g559) & (!g560) & (!g561) & (!g165) & (!g166)) + ((g558) & (!g559) & (!g560) & (g561) & (!g165) & (!g166)) + ((g558) & (!g559) & (!g560) & (g561) & (g165) & (g166)) + ((g558) & (!g559) & (g560) & (!g561) & (!g165) & (!g166)) + ((g558) & (!g559) & (g560) & (!g561) & (!g165) & (g166)) + ((g558) & (!g559) & (g560) & (g561) & (!g165) & (!g166)) + ((g558) & (!g559) & (g560) & (g561) & (!g165) & (g166)) + ((g558) & (!g559) & (g560) & (g561) & (g165) & (g166)) + ((g558) & (g559) & (!g560) & (!g561) & (!g165) & (!g166)) + ((g558) & (g559) & (!g560) & (!g561) & (g165) & (!g166)) + ((g558) & (g559) & (!g560) & (g561) & (!g165) & (!g166)) + ((g558) & (g559) & (!g560) & (g561) & (g165) & (!g166)) + ((g558) & (g559) & (!g560) & (g561) & (g165) & (g166)) + ((g558) & (g559) & (g560) & (!g561) & (!g165) & (!g166)) + ((g558) & (g559) & (g560) & (!g561) & (!g165) & (g166)) + ((g558) & (g559) & (g560) & (!g561) & (g165) & (!g166)) + ((g558) & (g559) & (g560) & (g561) & (!g165) & (!g166)) + ((g558) & (g559) & (g560) & (g561) & (!g165) & (g166)) + ((g558) & (g559) & (g560) & (g561) & (g165) & (!g166)) + ((g558) & (g559) & (g560) & (g561) & (g165) & (g166)));
	assign g563 = (((!g547) & (!g552) & (!g557) & (g562) & (g147) & (g148)) + ((!g547) & (!g552) & (g557) & (!g562) & (!g147) & (g148)) + ((!g547) & (!g552) & (g557) & (g562) & (!g147) & (g148)) + ((!g547) & (!g552) & (g557) & (g562) & (g147) & (g148)) + ((!g547) & (g552) & (!g557) & (!g562) & (g147) & (!g148)) + ((!g547) & (g552) & (!g557) & (g562) & (g147) & (!g148)) + ((!g547) & (g552) & (!g557) & (g562) & (g147) & (g148)) + ((!g547) & (g552) & (g557) & (!g562) & (!g147) & (g148)) + ((!g547) & (g552) & (g557) & (!g562) & (g147) & (!g148)) + ((!g547) & (g552) & (g557) & (g562) & (!g147) & (g148)) + ((!g547) & (g552) & (g557) & (g562) & (g147) & (!g148)) + ((!g547) & (g552) & (g557) & (g562) & (g147) & (g148)) + ((g547) & (!g552) & (!g557) & (!g562) & (!g147) & (!g148)) + ((g547) & (!g552) & (!g557) & (g562) & (!g147) & (!g148)) + ((g547) & (!g552) & (!g557) & (g562) & (g147) & (g148)) + ((g547) & (!g552) & (g557) & (!g562) & (!g147) & (!g148)) + ((g547) & (!g552) & (g557) & (!g562) & (!g147) & (g148)) + ((g547) & (!g552) & (g557) & (g562) & (!g147) & (!g148)) + ((g547) & (!g552) & (g557) & (g562) & (!g147) & (g148)) + ((g547) & (!g552) & (g557) & (g562) & (g147) & (g148)) + ((g547) & (g552) & (!g557) & (!g562) & (!g147) & (!g148)) + ((g547) & (g552) & (!g557) & (!g562) & (g147) & (!g148)) + ((g547) & (g552) & (!g557) & (g562) & (!g147) & (!g148)) + ((g547) & (g552) & (!g557) & (g562) & (g147) & (!g148)) + ((g547) & (g552) & (!g557) & (g562) & (g147) & (g148)) + ((g547) & (g552) & (g557) & (!g562) & (!g147) & (!g148)) + ((g547) & (g552) & (g557) & (!g562) & (!g147) & (g148)) + ((g547) & (g552) & (g557) & (!g562) & (g147) & (!g148)) + ((g547) & (g552) & (g557) & (g562) & (!g147) & (!g148)) + ((g547) & (g552) & (g557) & (g562) & (!g147) & (g148)) + ((g547) & (g552) & (g557) & (g562) & (g147) & (!g148)) + ((g547) & (g552) & (g557) & (g562) & (g147) & (g148)));
	assign g4292 = (((!sk[118]) & (!g2173) & (!g2407) & (g564)) + ((!sk[118]) & (!g2173) & (g2407) & (!g564)) + ((!sk[118]) & (!g2173) & (g2407) & (g564)) + ((!sk[118]) & (g2173) & (!g2407) & (g564)) + ((!sk[118]) & (g2173) & (g2407) & (!g564)) + ((!sk[118]) & (g2173) & (g2407) & (g564)) + ((sk[118]) & (!g2173) & (!g2407) & (g564)) + ((sk[118]) & (!g2173) & (g2407) & (g564)) + ((sk[118]) & (g2173) & (g2407) & (!g564)) + ((sk[118]) & (g2173) & (g2407) & (g564)));
	assign g4293 = (((!sk[119]) & (!g2174) & (!g2407) & (g565)) + ((!sk[119]) & (!g2174) & (g2407) & (!g565)) + ((!sk[119]) & (!g2174) & (g2407) & (g565)) + ((!sk[119]) & (g2174) & (!g2407) & (g565)) + ((!sk[119]) & (g2174) & (g2407) & (!g565)) + ((!sk[119]) & (g2174) & (g2407) & (g565)) + ((sk[119]) & (!g2174) & (!g2407) & (g565)) + ((sk[119]) & (!g2174) & (g2407) & (g565)) + ((sk[119]) & (g2174) & (g2407) & (!g565)) + ((sk[119]) & (g2174) & (g2407) & (g565)));
	assign g4294 = (((!g2175) & (!sk[120]) & (!g2407) & (g566)) + ((!g2175) & (!sk[120]) & (g2407) & (!g566)) + ((!g2175) & (!sk[120]) & (g2407) & (g566)) + ((!g2175) & (sk[120]) & (!g2407) & (g566)) + ((!g2175) & (sk[120]) & (g2407) & (g566)) + ((g2175) & (!sk[120]) & (!g2407) & (g566)) + ((g2175) & (!sk[120]) & (g2407) & (!g566)) + ((g2175) & (!sk[120]) & (g2407) & (g566)) + ((g2175) & (sk[120]) & (g2407) & (!g566)) + ((g2175) & (sk[120]) & (g2407) & (g566)));
	assign g4295 = (((!g2176) & (!g2407) & (!sk[121]) & (g567)) + ((!g2176) & (!g2407) & (sk[121]) & (g567)) + ((!g2176) & (g2407) & (!sk[121]) & (!g567)) + ((!g2176) & (g2407) & (!sk[121]) & (g567)) + ((!g2176) & (g2407) & (sk[121]) & (g567)) + ((g2176) & (!g2407) & (!sk[121]) & (g567)) + ((g2176) & (g2407) & (!sk[121]) & (!g567)) + ((g2176) & (g2407) & (!sk[121]) & (g567)) + ((g2176) & (g2407) & (sk[121]) & (!g567)) + ((g2176) & (g2407) & (sk[121]) & (g567)));
	assign g568 = (((!g564) & (!g565) & (!g566) & (g567) & (g165) & (g166)) + ((!g564) & (!g565) & (g566) & (!g567) & (!g165) & (g166)) + ((!g564) & (!g565) & (g566) & (g567) & (!g165) & (g166)) + ((!g564) & (!g565) & (g566) & (g567) & (g165) & (g166)) + ((!g564) & (g565) & (!g566) & (!g567) & (g165) & (!g166)) + ((!g564) & (g565) & (!g566) & (g567) & (g165) & (!g166)) + ((!g564) & (g565) & (!g566) & (g567) & (g165) & (g166)) + ((!g564) & (g565) & (g566) & (!g567) & (!g165) & (g166)) + ((!g564) & (g565) & (g566) & (!g567) & (g165) & (!g166)) + ((!g564) & (g565) & (g566) & (g567) & (!g165) & (g166)) + ((!g564) & (g565) & (g566) & (g567) & (g165) & (!g166)) + ((!g564) & (g565) & (g566) & (g567) & (g165) & (g166)) + ((g564) & (!g565) & (!g566) & (!g567) & (!g165) & (!g166)) + ((g564) & (!g565) & (!g566) & (g567) & (!g165) & (!g166)) + ((g564) & (!g565) & (!g566) & (g567) & (g165) & (g166)) + ((g564) & (!g565) & (g566) & (!g567) & (!g165) & (!g166)) + ((g564) & (!g565) & (g566) & (!g567) & (!g165) & (g166)) + ((g564) & (!g565) & (g566) & (g567) & (!g165) & (!g166)) + ((g564) & (!g565) & (g566) & (g567) & (!g165) & (g166)) + ((g564) & (!g565) & (g566) & (g567) & (g165) & (g166)) + ((g564) & (g565) & (!g566) & (!g567) & (!g165) & (!g166)) + ((g564) & (g565) & (!g566) & (!g567) & (g165) & (!g166)) + ((g564) & (g565) & (!g566) & (g567) & (!g165) & (!g166)) + ((g564) & (g565) & (!g566) & (g567) & (g165) & (!g166)) + ((g564) & (g565) & (!g566) & (g567) & (g165) & (g166)) + ((g564) & (g565) & (g566) & (!g567) & (!g165) & (!g166)) + ((g564) & (g565) & (g566) & (!g567) & (!g165) & (g166)) + ((g564) & (g565) & (g566) & (!g567) & (g165) & (!g166)) + ((g564) & (g565) & (g566) & (g567) & (!g165) & (!g166)) + ((g564) & (g565) & (g566) & (g567) & (!g165) & (g166)) + ((g564) & (g565) & (g566) & (g567) & (g165) & (!g166)) + ((g564) & (g565) & (g566) & (g567) & (g165) & (g166)));
	assign g4296 = (((!sk[123]) & (!g2177) & (!g2407) & (g569)) + ((!sk[123]) & (!g2177) & (g2407) & (!g569)) + ((!sk[123]) & (!g2177) & (g2407) & (g569)) + ((!sk[123]) & (g2177) & (!g2407) & (g569)) + ((!sk[123]) & (g2177) & (g2407) & (!g569)) + ((!sk[123]) & (g2177) & (g2407) & (g569)) + ((sk[123]) & (!g2177) & (!g2407) & (g569)) + ((sk[123]) & (!g2177) & (g2407) & (g569)) + ((sk[123]) & (g2177) & (g2407) & (!g569)) + ((sk[123]) & (g2177) & (g2407) & (g569)));
	assign g4297 = (((!sk[124]) & (!g2178) & (!g2407) & (g570)) + ((!sk[124]) & (!g2178) & (g2407) & (!g570)) + ((!sk[124]) & (!g2178) & (g2407) & (g570)) + ((!sk[124]) & (g2178) & (!g2407) & (g570)) + ((!sk[124]) & (g2178) & (g2407) & (!g570)) + ((!sk[124]) & (g2178) & (g2407) & (g570)) + ((sk[124]) & (!g2178) & (!g2407) & (g570)) + ((sk[124]) & (!g2178) & (g2407) & (g570)) + ((sk[124]) & (g2178) & (g2407) & (!g570)) + ((sk[124]) & (g2178) & (g2407) & (g570)));
	assign g4298 = (((!g2179) & (!g2407) & (!sk[125]) & (g571)) + ((!g2179) & (!g2407) & (sk[125]) & (g571)) + ((!g2179) & (g2407) & (!sk[125]) & (!g571)) + ((!g2179) & (g2407) & (!sk[125]) & (g571)) + ((!g2179) & (g2407) & (sk[125]) & (g571)) + ((g2179) & (!g2407) & (!sk[125]) & (g571)) + ((g2179) & (g2407) & (!sk[125]) & (!g571)) + ((g2179) & (g2407) & (!sk[125]) & (g571)) + ((g2179) & (g2407) & (sk[125]) & (!g571)) + ((g2179) & (g2407) & (sk[125]) & (g571)));
	assign g572 = (((!g165) & (!g166) & (!g569) & (!sk[126]) & (g570) & (!g571)) + ((!g165) & (!g166) & (!g569) & (!sk[126]) & (g570) & (g571)) + ((!g165) & (!g166) & (g569) & (!sk[126]) & (!g570) & (!g571)) + ((!g165) & (!g166) & (g569) & (!sk[126]) & (!g570) & (g571)) + ((!g165) & (!g166) & (g569) & (!sk[126]) & (g570) & (!g571)) + ((!g165) & (!g166) & (g569) & (!sk[126]) & (g570) & (g571)) + ((!g165) & (g166) & (!g569) & (!sk[126]) & (!g570) & (!g571)) + ((!g165) & (g166) & (!g569) & (!sk[126]) & (!g570) & (g571)) + ((!g165) & (g166) & (!g569) & (!sk[126]) & (g570) & (!g571)) + ((!g165) & (g166) & (!g569) & (!sk[126]) & (g570) & (g571)) + ((!g165) & (g166) & (!g569) & (sk[126]) & (!g570) & (g571)) + ((!g165) & (g166) & (!g569) & (sk[126]) & (g570) & (g571)) + ((!g165) & (g166) & (g569) & (!sk[126]) & (!g570) & (!g571)) + ((!g165) & (g166) & (g569) & (!sk[126]) & (!g570) & (g571)) + ((!g165) & (g166) & (g569) & (!sk[126]) & (g570) & (!g571)) + ((!g165) & (g166) & (g569) & (!sk[126]) & (g570) & (g571)) + ((!g165) & (g166) & (g569) & (sk[126]) & (!g570) & (g571)) + ((!g165) & (g166) & (g569) & (sk[126]) & (g570) & (g571)) + ((g165) & (!g166) & (!g569) & (!sk[126]) & (g570) & (!g571)) + ((g165) & (!g166) & (!g569) & (!sk[126]) & (g570) & (g571)) + ((g165) & (!g166) & (g569) & (!sk[126]) & (!g570) & (!g571)) + ((g165) & (!g166) & (g569) & (!sk[126]) & (!g570) & (g571)) + ((g165) & (!g166) & (g569) & (!sk[126]) & (g570) & (!g571)) + ((g165) & (!g166) & (g569) & (!sk[126]) & (g570) & (g571)) + ((g165) & (!g166) & (g569) & (sk[126]) & (!g570) & (!g571)) + ((g165) & (!g166) & (g569) & (sk[126]) & (!g570) & (g571)) + ((g165) & (!g166) & (g569) & (sk[126]) & (g570) & (!g571)) + ((g165) & (!g166) & (g569) & (sk[126]) & (g570) & (g571)) + ((g165) & (g166) & (!g569) & (!sk[126]) & (!g570) & (!g571)) + ((g165) & (g166) & (!g569) & (!sk[126]) & (!g570) & (g571)) + ((g165) & (g166) & (!g569) & (!sk[126]) & (g570) & (!g571)) + ((g165) & (g166) & (!g569) & (!sk[126]) & (g570) & (g571)) + ((g165) & (g166) & (!g569) & (sk[126]) & (g570) & (!g571)) + ((g165) & (g166) & (!g569) & (sk[126]) & (g570) & (g571)) + ((g165) & (g166) & (g569) & (!sk[126]) & (!g570) & (!g571)) + ((g165) & (g166) & (g569) & (!sk[126]) & (!g570) & (g571)) + ((g165) & (g166) & (g569) & (!sk[126]) & (g570) & (!g571)) + ((g165) & (g166) & (g569) & (!sk[126]) & (g570) & (g571)) + ((g165) & (g166) & (g569) & (sk[126]) & (g570) & (!g571)) + ((g165) & (g166) & (g569) & (sk[126]) & (g570) & (g571)));
	assign g4299 = (((!g2162) & (!g2407) & (!sk[127]) & (g573)) + ((!g2162) & (!g2407) & (sk[127]) & (g573)) + ((!g2162) & (g2407) & (!sk[127]) & (!g573)) + ((!g2162) & (g2407) & (!sk[127]) & (g573)) + ((!g2162) & (g2407) & (sk[127]) & (g573)) + ((g2162) & (!g2407) & (!sk[127]) & (g573)) + ((g2162) & (g2407) & (!sk[127]) & (!g573)) + ((g2162) & (g2407) & (!sk[127]) & (g573)) + ((g2162) & (g2407) & (sk[127]) & (!g573)) + ((g2162) & (g2407) & (sk[127]) & (g573)));
	assign g4300 = (((!sk[0]) & (!g2164) & (!g2407) & (g574)) + ((!sk[0]) & (!g2164) & (g2407) & (!g574)) + ((!sk[0]) & (!g2164) & (g2407) & (g574)) + ((!sk[0]) & (g2164) & (!g2407) & (g574)) + ((!sk[0]) & (g2164) & (g2407) & (!g574)) + ((!sk[0]) & (g2164) & (g2407) & (g574)) + ((sk[0]) & (!g2164) & (!g2407) & (g574)) + ((sk[0]) & (!g2164) & (g2407) & (g574)) + ((sk[0]) & (g2164) & (g2407) & (!g574)) + ((sk[0]) & (g2164) & (g2407) & (g574)));
	assign g4301 = (((!g2166) & (!g2407) & (!sk[1]) & (g575)) + ((!g2166) & (!g2407) & (sk[1]) & (g575)) + ((!g2166) & (g2407) & (!sk[1]) & (!g575)) + ((!g2166) & (g2407) & (!sk[1]) & (g575)) + ((!g2166) & (g2407) & (sk[1]) & (g575)) + ((g2166) & (!g2407) & (!sk[1]) & (g575)) + ((g2166) & (g2407) & (!sk[1]) & (!g575)) + ((g2166) & (g2407) & (!sk[1]) & (g575)) + ((g2166) & (g2407) & (sk[1]) & (!g575)) + ((g2166) & (g2407) & (sk[1]) & (g575)));
	assign g4302 = (((!sk[2]) & (!g2168) & (!g2407) & (g576)) + ((!sk[2]) & (!g2168) & (g2407) & (!g576)) + ((!sk[2]) & (!g2168) & (g2407) & (g576)) + ((!sk[2]) & (g2168) & (!g2407) & (g576)) + ((!sk[2]) & (g2168) & (g2407) & (!g576)) + ((!sk[2]) & (g2168) & (g2407) & (g576)) + ((sk[2]) & (!g2168) & (!g2407) & (g576)) + ((sk[2]) & (!g2168) & (g2407) & (g576)) + ((sk[2]) & (g2168) & (g2407) & (!g576)) + ((sk[2]) & (g2168) & (g2407) & (g576)));
	assign g577 = (((!g573) & (!g574) & (!g575) & (g576) & (g165) & (g166)) + ((!g573) & (!g574) & (g575) & (!g576) & (!g165) & (g166)) + ((!g573) & (!g574) & (g575) & (g576) & (!g165) & (g166)) + ((!g573) & (!g574) & (g575) & (g576) & (g165) & (g166)) + ((!g573) & (g574) & (!g575) & (!g576) & (g165) & (!g166)) + ((!g573) & (g574) & (!g575) & (g576) & (g165) & (!g166)) + ((!g573) & (g574) & (!g575) & (g576) & (g165) & (g166)) + ((!g573) & (g574) & (g575) & (!g576) & (!g165) & (g166)) + ((!g573) & (g574) & (g575) & (!g576) & (g165) & (!g166)) + ((!g573) & (g574) & (g575) & (g576) & (!g165) & (g166)) + ((!g573) & (g574) & (g575) & (g576) & (g165) & (!g166)) + ((!g573) & (g574) & (g575) & (g576) & (g165) & (g166)) + ((g573) & (!g574) & (!g575) & (!g576) & (!g165) & (!g166)) + ((g573) & (!g574) & (!g575) & (g576) & (!g165) & (!g166)) + ((g573) & (!g574) & (!g575) & (g576) & (g165) & (g166)) + ((g573) & (!g574) & (g575) & (!g576) & (!g165) & (!g166)) + ((g573) & (!g574) & (g575) & (!g576) & (!g165) & (g166)) + ((g573) & (!g574) & (g575) & (g576) & (!g165) & (!g166)) + ((g573) & (!g574) & (g575) & (g576) & (!g165) & (g166)) + ((g573) & (!g574) & (g575) & (g576) & (g165) & (g166)) + ((g573) & (g574) & (!g575) & (!g576) & (!g165) & (!g166)) + ((g573) & (g574) & (!g575) & (!g576) & (g165) & (!g166)) + ((g573) & (g574) & (!g575) & (g576) & (!g165) & (!g166)) + ((g573) & (g574) & (!g575) & (g576) & (g165) & (!g166)) + ((g573) & (g574) & (!g575) & (g576) & (g165) & (g166)) + ((g573) & (g574) & (g575) & (!g576) & (!g165) & (!g166)) + ((g573) & (g574) & (g575) & (!g576) & (!g165) & (g166)) + ((g573) & (g574) & (g575) & (!g576) & (g165) & (!g166)) + ((g573) & (g574) & (g575) & (g576) & (!g165) & (!g166)) + ((g573) & (g574) & (g575) & (g576) & (!g165) & (g166)) + ((g573) & (g574) & (g575) & (g576) & (g165) & (!g166)) + ((g573) & (g574) & (g575) & (g576) & (g165) & (g166)));
	assign g4303 = (((!g2169) & (!sk[4]) & (!g2407) & (g578)) + ((!g2169) & (!sk[4]) & (g2407) & (!g578)) + ((!g2169) & (!sk[4]) & (g2407) & (g578)) + ((!g2169) & (sk[4]) & (!g2407) & (g578)) + ((!g2169) & (sk[4]) & (g2407) & (g578)) + ((g2169) & (!sk[4]) & (!g2407) & (g578)) + ((g2169) & (!sk[4]) & (g2407) & (!g578)) + ((g2169) & (!sk[4]) & (g2407) & (g578)) + ((g2169) & (sk[4]) & (g2407) & (!g578)) + ((g2169) & (sk[4]) & (g2407) & (g578)));
	assign g4304 = (((!g2170) & (!g2407) & (!sk[5]) & (g579)) + ((!g2170) & (!g2407) & (sk[5]) & (g579)) + ((!g2170) & (g2407) & (!sk[5]) & (!g579)) + ((!g2170) & (g2407) & (!sk[5]) & (g579)) + ((!g2170) & (g2407) & (sk[5]) & (g579)) + ((g2170) & (!g2407) & (!sk[5]) & (g579)) + ((g2170) & (g2407) & (!sk[5]) & (!g579)) + ((g2170) & (g2407) & (!sk[5]) & (g579)) + ((g2170) & (g2407) & (sk[5]) & (!g579)) + ((g2170) & (g2407) & (sk[5]) & (g579)));
	assign g4305 = (((!g2171) & (!g2407) & (!sk[6]) & (g580)) + ((!g2171) & (!g2407) & (sk[6]) & (g580)) + ((!g2171) & (g2407) & (!sk[6]) & (!g580)) + ((!g2171) & (g2407) & (!sk[6]) & (g580)) + ((!g2171) & (g2407) & (sk[6]) & (g580)) + ((g2171) & (!g2407) & (!sk[6]) & (g580)) + ((g2171) & (g2407) & (!sk[6]) & (!g580)) + ((g2171) & (g2407) & (!sk[6]) & (g580)) + ((g2171) & (g2407) & (sk[6]) & (!g580)) + ((g2171) & (g2407) & (sk[6]) & (g580)));
	assign g4306 = (((!g2172) & (!g2407) & (!sk[7]) & (g581)) + ((!g2172) & (!g2407) & (sk[7]) & (g581)) + ((!g2172) & (g2407) & (!sk[7]) & (!g581)) + ((!g2172) & (g2407) & (!sk[7]) & (g581)) + ((!g2172) & (g2407) & (sk[7]) & (g581)) + ((g2172) & (!g2407) & (!sk[7]) & (g581)) + ((g2172) & (g2407) & (!sk[7]) & (!g581)) + ((g2172) & (g2407) & (!sk[7]) & (g581)) + ((g2172) & (g2407) & (sk[7]) & (!g581)) + ((g2172) & (g2407) & (sk[7]) & (g581)));
	assign g582 = (((!g578) & (!g579) & (!g580) & (g581) & (g165) & (g166)) + ((!g578) & (!g579) & (g580) & (!g581) & (!g165) & (g166)) + ((!g578) & (!g579) & (g580) & (g581) & (!g165) & (g166)) + ((!g578) & (!g579) & (g580) & (g581) & (g165) & (g166)) + ((!g578) & (g579) & (!g580) & (!g581) & (g165) & (!g166)) + ((!g578) & (g579) & (!g580) & (g581) & (g165) & (!g166)) + ((!g578) & (g579) & (!g580) & (g581) & (g165) & (g166)) + ((!g578) & (g579) & (g580) & (!g581) & (!g165) & (g166)) + ((!g578) & (g579) & (g580) & (!g581) & (g165) & (!g166)) + ((!g578) & (g579) & (g580) & (g581) & (!g165) & (g166)) + ((!g578) & (g579) & (g580) & (g581) & (g165) & (!g166)) + ((!g578) & (g579) & (g580) & (g581) & (g165) & (g166)) + ((g578) & (!g579) & (!g580) & (!g581) & (!g165) & (!g166)) + ((g578) & (!g579) & (!g580) & (g581) & (!g165) & (!g166)) + ((g578) & (!g579) & (!g580) & (g581) & (g165) & (g166)) + ((g578) & (!g579) & (g580) & (!g581) & (!g165) & (!g166)) + ((g578) & (!g579) & (g580) & (!g581) & (!g165) & (g166)) + ((g578) & (!g579) & (g580) & (g581) & (!g165) & (!g166)) + ((g578) & (!g579) & (g580) & (g581) & (!g165) & (g166)) + ((g578) & (!g579) & (g580) & (g581) & (g165) & (g166)) + ((g578) & (g579) & (!g580) & (!g581) & (!g165) & (!g166)) + ((g578) & (g579) & (!g580) & (!g581) & (g165) & (!g166)) + ((g578) & (g579) & (!g580) & (g581) & (!g165) & (!g166)) + ((g578) & (g579) & (!g580) & (g581) & (g165) & (!g166)) + ((g578) & (g579) & (!g580) & (g581) & (g165) & (g166)) + ((g578) & (g579) & (g580) & (!g581) & (!g165) & (!g166)) + ((g578) & (g579) & (g580) & (!g581) & (!g165) & (g166)) + ((g578) & (g579) & (g580) & (!g581) & (g165) & (!g166)) + ((g578) & (g579) & (g580) & (g581) & (!g165) & (!g166)) + ((g578) & (g579) & (g580) & (g581) & (!g165) & (g166)) + ((g578) & (g579) & (g580) & (g581) & (g165) & (!g166)) + ((g578) & (g579) & (g580) & (g581) & (g165) & (g166)));
	assign g583 = (((!g147) & (!g148) & (!g568) & (g572) & (!g577) & (!g582)) + ((!g147) & (!g148) & (!g568) & (g572) & (!g577) & (g582)) + ((!g147) & (!g148) & (!g568) & (g572) & (g577) & (!g582)) + ((!g147) & (!g148) & (!g568) & (g572) & (g577) & (g582)) + ((!g147) & (!g148) & (g568) & (g572) & (!g577) & (!g582)) + ((!g147) & (!g148) & (g568) & (g572) & (!g577) & (g582)) + ((!g147) & (!g148) & (g568) & (g572) & (g577) & (!g582)) + ((!g147) & (!g148) & (g568) & (g572) & (g577) & (g582)) + ((!g147) & (g148) & (!g568) & (!g572) & (!g577) & (g582)) + ((!g147) & (g148) & (!g568) & (!g572) & (g577) & (g582)) + ((!g147) & (g148) & (!g568) & (g572) & (!g577) & (g582)) + ((!g147) & (g148) & (!g568) & (g572) & (g577) & (g582)) + ((!g147) & (g148) & (g568) & (!g572) & (!g577) & (g582)) + ((!g147) & (g148) & (g568) & (!g572) & (g577) & (g582)) + ((!g147) & (g148) & (g568) & (g572) & (!g577) & (g582)) + ((!g147) & (g148) & (g568) & (g572) & (g577) & (g582)) + ((g147) & (!g148) & (g568) & (!g572) & (!g577) & (!g582)) + ((g147) & (!g148) & (g568) & (!g572) & (!g577) & (g582)) + ((g147) & (!g148) & (g568) & (!g572) & (g577) & (!g582)) + ((g147) & (!g148) & (g568) & (!g572) & (g577) & (g582)) + ((g147) & (!g148) & (g568) & (g572) & (!g577) & (!g582)) + ((g147) & (!g148) & (g568) & (g572) & (!g577) & (g582)) + ((g147) & (!g148) & (g568) & (g572) & (g577) & (!g582)) + ((g147) & (!g148) & (g568) & (g572) & (g577) & (g582)) + ((g147) & (g148) & (!g568) & (!g572) & (g577) & (!g582)) + ((g147) & (g148) & (!g568) & (!g572) & (g577) & (g582)) + ((g147) & (g148) & (!g568) & (g572) & (g577) & (!g582)) + ((g147) & (g148) & (!g568) & (g572) & (g577) & (g582)) + ((g147) & (g148) & (g568) & (!g572) & (g577) & (!g582)) + ((g147) & (g148) & (g568) & (!g572) & (g577) & (g582)) + ((g147) & (g148) & (g568) & (g572) & (g577) & (!g582)) + ((g147) & (g148) & (g568) & (g572) & (g577) & (g582)));
	assign g584 = (((!sk[10]) & (!g142) & (!g563) & (g583)) + ((!sk[10]) & (!g142) & (g563) & (!g583)) + ((!sk[10]) & (!g142) & (g563) & (g583)) + ((!sk[10]) & (g142) & (!g563) & (g583)) + ((!sk[10]) & (g142) & (g563) & (!g583)) + ((!sk[10]) & (g142) & (g563) & (g583)) + ((sk[10]) & (!g142) & (!g563) & (g583)) + ((sk[10]) & (!g142) & (g563) & (g583)) + ((sk[10]) & (g142) & (g563) & (!g583)) + ((sk[10]) & (g142) & (g563) & (g583)));
	assign g585 = (((!g91) & (!g126) & (!sk[11]) & (!g541) & (g542) & (!g584)) + ((!g91) & (!g126) & (!sk[11]) & (!g541) & (g542) & (g584)) + ((!g91) & (!g126) & (!sk[11]) & (g541) & (!g542) & (!g584)) + ((!g91) & (!g126) & (!sk[11]) & (g541) & (!g542) & (g584)) + ((!g91) & (!g126) & (!sk[11]) & (g541) & (g542) & (!g584)) + ((!g91) & (!g126) & (!sk[11]) & (g541) & (g542) & (g584)) + ((!g91) & (!g126) & (sk[11]) & (g541) & (!g542) & (!g584)) + ((!g91) & (!g126) & (sk[11]) & (g541) & (!g542) & (g584)) + ((!g91) & (!g126) & (sk[11]) & (g541) & (g542) & (!g584)) + ((!g91) & (!g126) & (sk[11]) & (g541) & (g542) & (g584)) + ((!g91) & (g126) & (!sk[11]) & (!g541) & (!g542) & (!g584)) + ((!g91) & (g126) & (!sk[11]) & (!g541) & (!g542) & (g584)) + ((!g91) & (g126) & (!sk[11]) & (!g541) & (g542) & (!g584)) + ((!g91) & (g126) & (!sk[11]) & (!g541) & (g542) & (g584)) + ((!g91) & (g126) & (!sk[11]) & (g541) & (!g542) & (!g584)) + ((!g91) & (g126) & (!sk[11]) & (g541) & (!g542) & (g584)) + ((!g91) & (g126) & (!sk[11]) & (g541) & (g542) & (!g584)) + ((!g91) & (g126) & (!sk[11]) & (g541) & (g542) & (g584)) + ((!g91) & (g126) & (sk[11]) & (!g541) & (!g542) & (g584)) + ((!g91) & (g126) & (sk[11]) & (!g541) & (g542) & (!g584)) + ((!g91) & (g126) & (sk[11]) & (g541) & (!g542) & (g584)) + ((!g91) & (g126) & (sk[11]) & (g541) & (g542) & (!g584)) + ((g91) & (!g126) & (!sk[11]) & (!g541) & (g542) & (!g584)) + ((g91) & (!g126) & (!sk[11]) & (!g541) & (g542) & (g584)) + ((g91) & (!g126) & (!sk[11]) & (g541) & (!g542) & (!g584)) + ((g91) & (!g126) & (!sk[11]) & (g541) & (!g542) & (g584)) + ((g91) & (!g126) & (!sk[11]) & (g541) & (g542) & (!g584)) + ((g91) & (!g126) & (!sk[11]) & (g541) & (g542) & (g584)) + ((g91) & (!g126) & (sk[11]) & (g541) & (!g542) & (!g584)) + ((g91) & (!g126) & (sk[11]) & (g541) & (!g542) & (g584)) + ((g91) & (!g126) & (sk[11]) & (g541) & (g542) & (!g584)) + ((g91) & (!g126) & (sk[11]) & (g541) & (g542) & (g584)) + ((g91) & (g126) & (!sk[11]) & (!g541) & (!g542) & (!g584)) + ((g91) & (g126) & (!sk[11]) & (!g541) & (!g542) & (g584)) + ((g91) & (g126) & (!sk[11]) & (!g541) & (g542) & (!g584)) + ((g91) & (g126) & (!sk[11]) & (!g541) & (g542) & (g584)) + ((g91) & (g126) & (!sk[11]) & (g541) & (!g542) & (!g584)) + ((g91) & (g126) & (!sk[11]) & (g541) & (!g542) & (g584)) + ((g91) & (g126) & (!sk[11]) & (g541) & (g542) & (!g584)) + ((g91) & (g126) & (!sk[11]) & (g541) & (g542) & (g584)) + ((g91) & (g126) & (sk[11]) & (!g541) & (!g542) & (!g584)) + ((g91) & (g126) & (sk[11]) & (!g541) & (g542) & (g584)) + ((g91) & (g126) & (sk[11]) & (g541) & (!g542) & (!g584)) + ((g91) & (g126) & (sk[11]) & (g541) & (g542) & (g584)));
	assign g4307 = (((!g2064) & (!sk[12]) & (!dmem_dat_ix10x) & (g586)) + ((!g2064) & (!sk[12]) & (dmem_dat_ix10x) & (!g586)) + ((!g2064) & (!sk[12]) & (dmem_dat_ix10x) & (g586)) + ((!g2064) & (sk[12]) & (!dmem_dat_ix10x) & (g586)) + ((!g2064) & (sk[12]) & (dmem_dat_ix10x) & (g586)) + ((g2064) & (!sk[12]) & (!dmem_dat_ix10x) & (g586)) + ((g2064) & (!sk[12]) & (dmem_dat_ix10x) & (!g586)) + ((g2064) & (!sk[12]) & (dmem_dat_ix10x) & (g586)) + ((g2064) & (sk[12]) & (dmem_dat_ix10x) & (!g586)) + ((g2064) & (sk[12]) & (dmem_dat_ix10x) & (g586)));
	assign g4308 = (((!g2059) & (!sk[13]) & (!g2415) & (g587)) + ((!g2059) & (!sk[13]) & (g2415) & (!g587)) + ((!g2059) & (!sk[13]) & (g2415) & (g587)) + ((!g2059) & (sk[13]) & (!g2415) & (g587)) + ((!g2059) & (sk[13]) & (g2415) & (g587)) + ((g2059) & (!sk[13]) & (!g2415) & (g587)) + ((g2059) & (!sk[13]) & (g2415) & (!g587)) + ((g2059) & (!sk[13]) & (g2415) & (g587)) + ((g2059) & (sk[13]) & (g2415) & (!g587)) + ((g2059) & (sk[13]) & (g2415) & (g587)));
	assign g4309 = (((!g2140) & (!g2431) & (!sk[14]) & (g588)) + ((!g2140) & (!g2431) & (sk[14]) & (g588)) + ((!g2140) & (g2431) & (!sk[14]) & (!g588)) + ((!g2140) & (g2431) & (!sk[14]) & (g588)) + ((!g2140) & (g2431) & (sk[14]) & (g588)) + ((g2140) & (!g2431) & (!sk[14]) & (g588)) + ((g2140) & (g2431) & (!sk[14]) & (!g588)) + ((g2140) & (g2431) & (!sk[14]) & (g588)) + ((g2140) & (g2431) & (sk[14]) & (!g588)) + ((g2140) & (g2431) & (sk[14]) & (g588)));
	assign g4310 = (((!g2142) & (!g2431) & (!sk[15]) & (g589)) + ((!g2142) & (!g2431) & (sk[15]) & (g589)) + ((!g2142) & (g2431) & (!sk[15]) & (!g589)) + ((!g2142) & (g2431) & (!sk[15]) & (g589)) + ((!g2142) & (g2431) & (sk[15]) & (g589)) + ((g2142) & (!g2431) & (!sk[15]) & (g589)) + ((g2142) & (g2431) & (!sk[15]) & (!g589)) + ((g2142) & (g2431) & (!sk[15]) & (g589)) + ((g2142) & (g2431) & (sk[15]) & (!g589)) + ((g2142) & (g2431) & (sk[15]) & (g589)));
	assign g4311 = (((!g2144) & (!sk[16]) & (!g2431) & (g590)) + ((!g2144) & (!sk[16]) & (g2431) & (!g590)) + ((!g2144) & (!sk[16]) & (g2431) & (g590)) + ((!g2144) & (sk[16]) & (!g2431) & (g590)) + ((!g2144) & (sk[16]) & (g2431) & (g590)) + ((g2144) & (!sk[16]) & (!g2431) & (g590)) + ((g2144) & (!sk[16]) & (g2431) & (!g590)) + ((g2144) & (!sk[16]) & (g2431) & (g590)) + ((g2144) & (sk[16]) & (g2431) & (!g590)) + ((g2144) & (sk[16]) & (g2431) & (g590)));
	assign g4312 = (((!sk[17]) & (!g2145) & (!g2431) & (g591)) + ((!sk[17]) & (!g2145) & (g2431) & (!g591)) + ((!sk[17]) & (!g2145) & (g2431) & (g591)) + ((!sk[17]) & (g2145) & (!g2431) & (g591)) + ((!sk[17]) & (g2145) & (g2431) & (!g591)) + ((!sk[17]) & (g2145) & (g2431) & (g591)) + ((sk[17]) & (!g2145) & (!g2431) & (g591)) + ((sk[17]) & (!g2145) & (g2431) & (g591)) + ((sk[17]) & (g2145) & (g2431) & (!g591)) + ((sk[17]) & (g2145) & (g2431) & (g591)));
	assign g592 = (((!g588) & (!g589) & (!g590) & (g591) & (g147) & (g148)) + ((!g588) & (!g589) & (g590) & (!g591) & (!g147) & (g148)) + ((!g588) & (!g589) & (g590) & (g591) & (!g147) & (g148)) + ((!g588) & (!g589) & (g590) & (g591) & (g147) & (g148)) + ((!g588) & (g589) & (!g590) & (!g591) & (g147) & (!g148)) + ((!g588) & (g589) & (!g590) & (g591) & (g147) & (!g148)) + ((!g588) & (g589) & (!g590) & (g591) & (g147) & (g148)) + ((!g588) & (g589) & (g590) & (!g591) & (!g147) & (g148)) + ((!g588) & (g589) & (g590) & (!g591) & (g147) & (!g148)) + ((!g588) & (g589) & (g590) & (g591) & (!g147) & (g148)) + ((!g588) & (g589) & (g590) & (g591) & (g147) & (!g148)) + ((!g588) & (g589) & (g590) & (g591) & (g147) & (g148)) + ((g588) & (!g589) & (!g590) & (!g591) & (!g147) & (!g148)) + ((g588) & (!g589) & (!g590) & (g591) & (!g147) & (!g148)) + ((g588) & (!g589) & (!g590) & (g591) & (g147) & (g148)) + ((g588) & (!g589) & (g590) & (!g591) & (!g147) & (!g148)) + ((g588) & (!g589) & (g590) & (!g591) & (!g147) & (g148)) + ((g588) & (!g589) & (g590) & (g591) & (!g147) & (!g148)) + ((g588) & (!g589) & (g590) & (g591) & (!g147) & (g148)) + ((g588) & (!g589) & (g590) & (g591) & (g147) & (g148)) + ((g588) & (g589) & (!g590) & (!g591) & (!g147) & (!g148)) + ((g588) & (g589) & (!g590) & (!g591) & (g147) & (!g148)) + ((g588) & (g589) & (!g590) & (g591) & (!g147) & (!g148)) + ((g588) & (g589) & (!g590) & (g591) & (g147) & (!g148)) + ((g588) & (g589) & (!g590) & (g591) & (g147) & (g148)) + ((g588) & (g589) & (g590) & (!g591) & (!g147) & (!g148)) + ((g588) & (g589) & (g590) & (!g591) & (!g147) & (g148)) + ((g588) & (g589) & (g590) & (!g591) & (g147) & (!g148)) + ((g588) & (g589) & (g590) & (g591) & (!g147) & (!g148)) + ((g588) & (g589) & (g590) & (g591) & (!g147) & (g148)) + ((g588) & (g589) & (g590) & (g591) & (g147) & (!g148)) + ((g588) & (g589) & (g590) & (g591) & (g147) & (g148)));
	assign g4313 = (((!g2146) & (!sk[19]) & (!g2431) & (g593)) + ((!g2146) & (!sk[19]) & (g2431) & (!g593)) + ((!g2146) & (!sk[19]) & (g2431) & (g593)) + ((!g2146) & (sk[19]) & (!g2431) & (g593)) + ((!g2146) & (sk[19]) & (g2431) & (g593)) + ((g2146) & (!sk[19]) & (!g2431) & (g593)) + ((g2146) & (!sk[19]) & (g2431) & (!g593)) + ((g2146) & (!sk[19]) & (g2431) & (g593)) + ((g2146) & (sk[19]) & (g2431) & (!g593)) + ((g2146) & (sk[19]) & (g2431) & (g593)));
	assign g4314 = (((!g2148) & (!g2431) & (!sk[20]) & (g594)) + ((!g2148) & (!g2431) & (sk[20]) & (g594)) + ((!g2148) & (g2431) & (!sk[20]) & (!g594)) + ((!g2148) & (g2431) & (!sk[20]) & (g594)) + ((!g2148) & (g2431) & (sk[20]) & (g594)) + ((g2148) & (!g2431) & (!sk[20]) & (g594)) + ((g2148) & (g2431) & (!sk[20]) & (!g594)) + ((g2148) & (g2431) & (!sk[20]) & (g594)) + ((g2148) & (g2431) & (sk[20]) & (!g594)) + ((g2148) & (g2431) & (sk[20]) & (g594)));
	assign g4315 = (((!sk[21]) & (!g2150) & (!g2431) & (g595)) + ((!sk[21]) & (!g2150) & (g2431) & (!g595)) + ((!sk[21]) & (!g2150) & (g2431) & (g595)) + ((!sk[21]) & (g2150) & (!g2431) & (g595)) + ((!sk[21]) & (g2150) & (g2431) & (!g595)) + ((!sk[21]) & (g2150) & (g2431) & (g595)) + ((sk[21]) & (!g2150) & (!g2431) & (g595)) + ((sk[21]) & (!g2150) & (g2431) & (g595)) + ((sk[21]) & (g2150) & (g2431) & (!g595)) + ((sk[21]) & (g2150) & (g2431) & (g595)));
	assign g4316 = (((!g2151) & (!g2431) & (!sk[22]) & (g596)) + ((!g2151) & (!g2431) & (sk[22]) & (g596)) + ((!g2151) & (g2431) & (!sk[22]) & (!g596)) + ((!g2151) & (g2431) & (!sk[22]) & (g596)) + ((!g2151) & (g2431) & (sk[22]) & (g596)) + ((g2151) & (!g2431) & (!sk[22]) & (g596)) + ((g2151) & (g2431) & (!sk[22]) & (!g596)) + ((g2151) & (g2431) & (!sk[22]) & (g596)) + ((g2151) & (g2431) & (sk[22]) & (!g596)) + ((g2151) & (g2431) & (sk[22]) & (g596)));
	assign g597 = (((!g593) & (!g594) & (!g595) & (g596) & (g147) & (g148)) + ((!g593) & (!g594) & (g595) & (!g596) & (!g147) & (g148)) + ((!g593) & (!g594) & (g595) & (g596) & (!g147) & (g148)) + ((!g593) & (!g594) & (g595) & (g596) & (g147) & (g148)) + ((!g593) & (g594) & (!g595) & (!g596) & (g147) & (!g148)) + ((!g593) & (g594) & (!g595) & (g596) & (g147) & (!g148)) + ((!g593) & (g594) & (!g595) & (g596) & (g147) & (g148)) + ((!g593) & (g594) & (g595) & (!g596) & (!g147) & (g148)) + ((!g593) & (g594) & (g595) & (!g596) & (g147) & (!g148)) + ((!g593) & (g594) & (g595) & (g596) & (!g147) & (g148)) + ((!g593) & (g594) & (g595) & (g596) & (g147) & (!g148)) + ((!g593) & (g594) & (g595) & (g596) & (g147) & (g148)) + ((g593) & (!g594) & (!g595) & (!g596) & (!g147) & (!g148)) + ((g593) & (!g594) & (!g595) & (g596) & (!g147) & (!g148)) + ((g593) & (!g594) & (!g595) & (g596) & (g147) & (g148)) + ((g593) & (!g594) & (g595) & (!g596) & (!g147) & (!g148)) + ((g593) & (!g594) & (g595) & (!g596) & (!g147) & (g148)) + ((g593) & (!g594) & (g595) & (g596) & (!g147) & (!g148)) + ((g593) & (!g594) & (g595) & (g596) & (!g147) & (g148)) + ((g593) & (!g594) & (g595) & (g596) & (g147) & (g148)) + ((g593) & (g594) & (!g595) & (!g596) & (!g147) & (!g148)) + ((g593) & (g594) & (!g595) & (!g596) & (g147) & (!g148)) + ((g593) & (g594) & (!g595) & (g596) & (!g147) & (!g148)) + ((g593) & (g594) & (!g595) & (g596) & (g147) & (!g148)) + ((g593) & (g594) & (!g595) & (g596) & (g147) & (g148)) + ((g593) & (g594) & (g595) & (!g596) & (!g147) & (!g148)) + ((g593) & (g594) & (g595) & (!g596) & (!g147) & (g148)) + ((g593) & (g594) & (g595) & (!g596) & (g147) & (!g148)) + ((g593) & (g594) & (g595) & (g596) & (!g147) & (!g148)) + ((g593) & (g594) & (g595) & (g596) & (!g147) & (g148)) + ((g593) & (g594) & (g595) & (g596) & (g147) & (!g148)) + ((g593) & (g594) & (g595) & (g596) & (g147) & (g148)));
	assign g4317 = (((!g2152) & (!sk[24]) & (!g2431) & (g598)) + ((!g2152) & (!sk[24]) & (g2431) & (!g598)) + ((!g2152) & (!sk[24]) & (g2431) & (g598)) + ((!g2152) & (sk[24]) & (!g2431) & (g598)) + ((!g2152) & (sk[24]) & (g2431) & (g598)) + ((g2152) & (!sk[24]) & (!g2431) & (g598)) + ((g2152) & (!sk[24]) & (g2431) & (!g598)) + ((g2152) & (!sk[24]) & (g2431) & (g598)) + ((g2152) & (sk[24]) & (g2431) & (!g598)) + ((g2152) & (sk[24]) & (g2431) & (g598)));
	assign g4318 = (((!g2153) & (!sk[25]) & (!g2431) & (g599)) + ((!g2153) & (!sk[25]) & (g2431) & (!g599)) + ((!g2153) & (!sk[25]) & (g2431) & (g599)) + ((!g2153) & (sk[25]) & (!g2431) & (g599)) + ((!g2153) & (sk[25]) & (g2431) & (g599)) + ((g2153) & (!sk[25]) & (!g2431) & (g599)) + ((g2153) & (!sk[25]) & (g2431) & (!g599)) + ((g2153) & (!sk[25]) & (g2431) & (g599)) + ((g2153) & (sk[25]) & (g2431) & (!g599)) + ((g2153) & (sk[25]) & (g2431) & (g599)));
	assign g4319 = (((!g2155) & (!sk[26]) & (!g2431) & (g600)) + ((!g2155) & (!sk[26]) & (g2431) & (!g600)) + ((!g2155) & (!sk[26]) & (g2431) & (g600)) + ((!g2155) & (sk[26]) & (!g2431) & (g600)) + ((!g2155) & (sk[26]) & (g2431) & (g600)) + ((g2155) & (!sk[26]) & (!g2431) & (g600)) + ((g2155) & (!sk[26]) & (g2431) & (!g600)) + ((g2155) & (!sk[26]) & (g2431) & (g600)) + ((g2155) & (sk[26]) & (g2431) & (!g600)) + ((g2155) & (sk[26]) & (g2431) & (g600)));
	assign g4320 = (((!sk[27]) & (!g2157) & (!g2431) & (g601)) + ((!sk[27]) & (!g2157) & (g2431) & (!g601)) + ((!sk[27]) & (!g2157) & (g2431) & (g601)) + ((!sk[27]) & (g2157) & (!g2431) & (g601)) + ((!sk[27]) & (g2157) & (g2431) & (!g601)) + ((!sk[27]) & (g2157) & (g2431) & (g601)) + ((sk[27]) & (!g2157) & (!g2431) & (g601)) + ((sk[27]) & (!g2157) & (g2431) & (g601)) + ((sk[27]) & (g2157) & (g2431) & (!g601)) + ((sk[27]) & (g2157) & (g2431) & (g601)));
	assign g602 = (((!g598) & (!g599) & (!g600) & (g601) & (g147) & (g148)) + ((!g598) & (!g599) & (g600) & (!g601) & (!g147) & (g148)) + ((!g598) & (!g599) & (g600) & (g601) & (!g147) & (g148)) + ((!g598) & (!g599) & (g600) & (g601) & (g147) & (g148)) + ((!g598) & (g599) & (!g600) & (!g601) & (g147) & (!g148)) + ((!g598) & (g599) & (!g600) & (g601) & (g147) & (!g148)) + ((!g598) & (g599) & (!g600) & (g601) & (g147) & (g148)) + ((!g598) & (g599) & (g600) & (!g601) & (!g147) & (g148)) + ((!g598) & (g599) & (g600) & (!g601) & (g147) & (!g148)) + ((!g598) & (g599) & (g600) & (g601) & (!g147) & (g148)) + ((!g598) & (g599) & (g600) & (g601) & (g147) & (!g148)) + ((!g598) & (g599) & (g600) & (g601) & (g147) & (g148)) + ((g598) & (!g599) & (!g600) & (!g601) & (!g147) & (!g148)) + ((g598) & (!g599) & (!g600) & (g601) & (!g147) & (!g148)) + ((g598) & (!g599) & (!g600) & (g601) & (g147) & (g148)) + ((g598) & (!g599) & (g600) & (!g601) & (!g147) & (!g148)) + ((g598) & (!g599) & (g600) & (!g601) & (!g147) & (g148)) + ((g598) & (!g599) & (g600) & (g601) & (!g147) & (!g148)) + ((g598) & (!g599) & (g600) & (g601) & (!g147) & (g148)) + ((g598) & (!g599) & (g600) & (g601) & (g147) & (g148)) + ((g598) & (g599) & (!g600) & (!g601) & (!g147) & (!g148)) + ((g598) & (g599) & (!g600) & (!g601) & (g147) & (!g148)) + ((g598) & (g599) & (!g600) & (g601) & (!g147) & (!g148)) + ((g598) & (g599) & (!g600) & (g601) & (g147) & (!g148)) + ((g598) & (g599) & (!g600) & (g601) & (g147) & (g148)) + ((g598) & (g599) & (g600) & (!g601) & (!g147) & (!g148)) + ((g598) & (g599) & (g600) & (!g601) & (!g147) & (g148)) + ((g598) & (g599) & (g600) & (!g601) & (g147) & (!g148)) + ((g598) & (g599) & (g600) & (g601) & (!g147) & (!g148)) + ((g598) & (g599) & (g600) & (g601) & (!g147) & (g148)) + ((g598) & (g599) & (g600) & (g601) & (g147) & (!g148)) + ((g598) & (g599) & (g600) & (g601) & (g147) & (g148)));
	assign g4321 = (((!g2158) & (!g2431) & (!sk[29]) & (g603)) + ((!g2158) & (!g2431) & (sk[29]) & (g603)) + ((!g2158) & (g2431) & (!sk[29]) & (!g603)) + ((!g2158) & (g2431) & (!sk[29]) & (g603)) + ((!g2158) & (g2431) & (sk[29]) & (g603)) + ((g2158) & (!g2431) & (!sk[29]) & (g603)) + ((g2158) & (g2431) & (!sk[29]) & (!g603)) + ((g2158) & (g2431) & (!sk[29]) & (g603)) + ((g2158) & (g2431) & (sk[29]) & (!g603)) + ((g2158) & (g2431) & (sk[29]) & (g603)));
	assign g4322 = (((!g2159) & (!sk[30]) & (!g2431) & (g604)) + ((!g2159) & (!sk[30]) & (g2431) & (!g604)) + ((!g2159) & (!sk[30]) & (g2431) & (g604)) + ((!g2159) & (sk[30]) & (!g2431) & (g604)) + ((!g2159) & (sk[30]) & (g2431) & (g604)) + ((g2159) & (!sk[30]) & (!g2431) & (g604)) + ((g2159) & (!sk[30]) & (g2431) & (!g604)) + ((g2159) & (!sk[30]) & (g2431) & (g604)) + ((g2159) & (sk[30]) & (g2431) & (!g604)) + ((g2159) & (sk[30]) & (g2431) & (g604)));
	assign g4323 = (((!g2160) & (!g2431) & (!sk[31]) & (g605)) + ((!g2160) & (!g2431) & (sk[31]) & (g605)) + ((!g2160) & (g2431) & (!sk[31]) & (!g605)) + ((!g2160) & (g2431) & (!sk[31]) & (g605)) + ((!g2160) & (g2431) & (sk[31]) & (g605)) + ((g2160) & (!g2431) & (!sk[31]) & (g605)) + ((g2160) & (g2431) & (!sk[31]) & (!g605)) + ((g2160) & (g2431) & (!sk[31]) & (g605)) + ((g2160) & (g2431) & (sk[31]) & (!g605)) + ((g2160) & (g2431) & (sk[31]) & (g605)));
	assign g4324 = (((!sk[32]) & (!g2161) & (!g2431) & (g606)) + ((!sk[32]) & (!g2161) & (g2431) & (!g606)) + ((!sk[32]) & (!g2161) & (g2431) & (g606)) + ((!sk[32]) & (g2161) & (!g2431) & (g606)) + ((!sk[32]) & (g2161) & (g2431) & (!g606)) + ((!sk[32]) & (g2161) & (g2431) & (g606)) + ((sk[32]) & (!g2161) & (!g2431) & (g606)) + ((sk[32]) & (!g2161) & (g2431) & (g606)) + ((sk[32]) & (g2161) & (g2431) & (!g606)) + ((sk[32]) & (g2161) & (g2431) & (g606)));
	assign g607 = (((!g603) & (!g604) & (!g605) & (g606) & (g147) & (g148)) + ((!g603) & (!g604) & (g605) & (!g606) & (!g147) & (g148)) + ((!g603) & (!g604) & (g605) & (g606) & (!g147) & (g148)) + ((!g603) & (!g604) & (g605) & (g606) & (g147) & (g148)) + ((!g603) & (g604) & (!g605) & (!g606) & (g147) & (!g148)) + ((!g603) & (g604) & (!g605) & (g606) & (g147) & (!g148)) + ((!g603) & (g604) & (!g605) & (g606) & (g147) & (g148)) + ((!g603) & (g604) & (g605) & (!g606) & (!g147) & (g148)) + ((!g603) & (g604) & (g605) & (!g606) & (g147) & (!g148)) + ((!g603) & (g604) & (g605) & (g606) & (!g147) & (g148)) + ((!g603) & (g604) & (g605) & (g606) & (g147) & (!g148)) + ((!g603) & (g604) & (g605) & (g606) & (g147) & (g148)) + ((g603) & (!g604) & (!g605) & (!g606) & (!g147) & (!g148)) + ((g603) & (!g604) & (!g605) & (g606) & (!g147) & (!g148)) + ((g603) & (!g604) & (!g605) & (g606) & (g147) & (g148)) + ((g603) & (!g604) & (g605) & (!g606) & (!g147) & (!g148)) + ((g603) & (!g604) & (g605) & (!g606) & (!g147) & (g148)) + ((g603) & (!g604) & (g605) & (g606) & (!g147) & (!g148)) + ((g603) & (!g604) & (g605) & (g606) & (!g147) & (g148)) + ((g603) & (!g604) & (g605) & (g606) & (g147) & (g148)) + ((g603) & (g604) & (!g605) & (!g606) & (!g147) & (!g148)) + ((g603) & (g604) & (!g605) & (!g606) & (g147) & (!g148)) + ((g603) & (g604) & (!g605) & (g606) & (!g147) & (!g148)) + ((g603) & (g604) & (!g605) & (g606) & (g147) & (!g148)) + ((g603) & (g604) & (!g605) & (g606) & (g147) & (g148)) + ((g603) & (g604) & (g605) & (!g606) & (!g147) & (!g148)) + ((g603) & (g604) & (g605) & (!g606) & (!g147) & (g148)) + ((g603) & (g604) & (g605) & (!g606) & (g147) & (!g148)) + ((g603) & (g604) & (g605) & (g606) & (!g147) & (!g148)) + ((g603) & (g604) & (g605) & (g606) & (!g147) & (g148)) + ((g603) & (g604) & (g605) & (g606) & (g147) & (!g148)) + ((g603) & (g604) & (g605) & (g606) & (g147) & (g148)));
	assign g608 = (((!g592) & (!g597) & (!g602) & (g607) & (g165) & (g166)) + ((!g592) & (!g597) & (g602) & (!g607) & (!g165) & (g166)) + ((!g592) & (!g597) & (g602) & (g607) & (!g165) & (g166)) + ((!g592) & (!g597) & (g602) & (g607) & (g165) & (g166)) + ((!g592) & (g597) & (!g602) & (!g607) & (g165) & (!g166)) + ((!g592) & (g597) & (!g602) & (g607) & (g165) & (!g166)) + ((!g592) & (g597) & (!g602) & (g607) & (g165) & (g166)) + ((!g592) & (g597) & (g602) & (!g607) & (!g165) & (g166)) + ((!g592) & (g597) & (g602) & (!g607) & (g165) & (!g166)) + ((!g592) & (g597) & (g602) & (g607) & (!g165) & (g166)) + ((!g592) & (g597) & (g602) & (g607) & (g165) & (!g166)) + ((!g592) & (g597) & (g602) & (g607) & (g165) & (g166)) + ((g592) & (!g597) & (!g602) & (!g607) & (!g165) & (!g166)) + ((g592) & (!g597) & (!g602) & (g607) & (!g165) & (!g166)) + ((g592) & (!g597) & (!g602) & (g607) & (g165) & (g166)) + ((g592) & (!g597) & (g602) & (!g607) & (!g165) & (!g166)) + ((g592) & (!g597) & (g602) & (!g607) & (!g165) & (g166)) + ((g592) & (!g597) & (g602) & (g607) & (!g165) & (!g166)) + ((g592) & (!g597) & (g602) & (g607) & (!g165) & (g166)) + ((g592) & (!g597) & (g602) & (g607) & (g165) & (g166)) + ((g592) & (g597) & (!g602) & (!g607) & (!g165) & (!g166)) + ((g592) & (g597) & (!g602) & (!g607) & (g165) & (!g166)) + ((g592) & (g597) & (!g602) & (g607) & (!g165) & (!g166)) + ((g592) & (g597) & (!g602) & (g607) & (g165) & (!g166)) + ((g592) & (g597) & (!g602) & (g607) & (g165) & (g166)) + ((g592) & (g597) & (g602) & (!g607) & (!g165) & (!g166)) + ((g592) & (g597) & (g602) & (!g607) & (!g165) & (g166)) + ((g592) & (g597) & (g602) & (!g607) & (g165) & (!g166)) + ((g592) & (g597) & (g602) & (g607) & (!g165) & (!g166)) + ((g592) & (g597) & (g602) & (g607) & (!g165) & (g166)) + ((g592) & (g597) & (g602) & (g607) & (g165) & (!g166)) + ((g592) & (g597) & (g602) & (g607) & (g165) & (g166)));
	assign g4325 = (((!sk[35]) & (!g2173) & (!g2431) & (g609)) + ((!sk[35]) & (!g2173) & (g2431) & (!g609)) + ((!sk[35]) & (!g2173) & (g2431) & (g609)) + ((!sk[35]) & (g2173) & (!g2431) & (g609)) + ((!sk[35]) & (g2173) & (g2431) & (!g609)) + ((!sk[35]) & (g2173) & (g2431) & (g609)) + ((sk[35]) & (!g2173) & (!g2431) & (g609)) + ((sk[35]) & (!g2173) & (g2431) & (g609)) + ((sk[35]) & (g2173) & (g2431) & (!g609)) + ((sk[35]) & (g2173) & (g2431) & (g609)));
	assign g4326 = (((!g2174) & (!g2431) & (!sk[36]) & (g610)) + ((!g2174) & (!g2431) & (sk[36]) & (g610)) + ((!g2174) & (g2431) & (!sk[36]) & (!g610)) + ((!g2174) & (g2431) & (!sk[36]) & (g610)) + ((!g2174) & (g2431) & (sk[36]) & (g610)) + ((g2174) & (!g2431) & (!sk[36]) & (g610)) + ((g2174) & (g2431) & (!sk[36]) & (!g610)) + ((g2174) & (g2431) & (!sk[36]) & (g610)) + ((g2174) & (g2431) & (sk[36]) & (!g610)) + ((g2174) & (g2431) & (sk[36]) & (g610)));
	assign g4327 = (((!sk[37]) & (!g2175) & (!g2431) & (g611)) + ((!sk[37]) & (!g2175) & (g2431) & (!g611)) + ((!sk[37]) & (!g2175) & (g2431) & (g611)) + ((!sk[37]) & (g2175) & (!g2431) & (g611)) + ((!sk[37]) & (g2175) & (g2431) & (!g611)) + ((!sk[37]) & (g2175) & (g2431) & (g611)) + ((sk[37]) & (!g2175) & (!g2431) & (g611)) + ((sk[37]) & (!g2175) & (g2431) & (g611)) + ((sk[37]) & (g2175) & (g2431) & (!g611)) + ((sk[37]) & (g2175) & (g2431) & (g611)));
	assign g4328 = (((!sk[38]) & (!g2176) & (!g2431) & (g612)) + ((!sk[38]) & (!g2176) & (g2431) & (!g612)) + ((!sk[38]) & (!g2176) & (g2431) & (g612)) + ((!sk[38]) & (g2176) & (!g2431) & (g612)) + ((!sk[38]) & (g2176) & (g2431) & (!g612)) + ((!sk[38]) & (g2176) & (g2431) & (g612)) + ((sk[38]) & (!g2176) & (!g2431) & (g612)) + ((sk[38]) & (!g2176) & (g2431) & (g612)) + ((sk[38]) & (g2176) & (g2431) & (!g612)) + ((sk[38]) & (g2176) & (g2431) & (g612)));
	assign g613 = (((!g609) & (!g610) & (!g611) & (g612) & (g165) & (g166)) + ((!g609) & (!g610) & (g611) & (!g612) & (!g165) & (g166)) + ((!g609) & (!g610) & (g611) & (g612) & (!g165) & (g166)) + ((!g609) & (!g610) & (g611) & (g612) & (g165) & (g166)) + ((!g609) & (g610) & (!g611) & (!g612) & (g165) & (!g166)) + ((!g609) & (g610) & (!g611) & (g612) & (g165) & (!g166)) + ((!g609) & (g610) & (!g611) & (g612) & (g165) & (g166)) + ((!g609) & (g610) & (g611) & (!g612) & (!g165) & (g166)) + ((!g609) & (g610) & (g611) & (!g612) & (g165) & (!g166)) + ((!g609) & (g610) & (g611) & (g612) & (!g165) & (g166)) + ((!g609) & (g610) & (g611) & (g612) & (g165) & (!g166)) + ((!g609) & (g610) & (g611) & (g612) & (g165) & (g166)) + ((g609) & (!g610) & (!g611) & (!g612) & (!g165) & (!g166)) + ((g609) & (!g610) & (!g611) & (g612) & (!g165) & (!g166)) + ((g609) & (!g610) & (!g611) & (g612) & (g165) & (g166)) + ((g609) & (!g610) & (g611) & (!g612) & (!g165) & (!g166)) + ((g609) & (!g610) & (g611) & (!g612) & (!g165) & (g166)) + ((g609) & (!g610) & (g611) & (g612) & (!g165) & (!g166)) + ((g609) & (!g610) & (g611) & (g612) & (!g165) & (g166)) + ((g609) & (!g610) & (g611) & (g612) & (g165) & (g166)) + ((g609) & (g610) & (!g611) & (!g612) & (!g165) & (!g166)) + ((g609) & (g610) & (!g611) & (!g612) & (g165) & (!g166)) + ((g609) & (g610) & (!g611) & (g612) & (!g165) & (!g166)) + ((g609) & (g610) & (!g611) & (g612) & (g165) & (!g166)) + ((g609) & (g610) & (!g611) & (g612) & (g165) & (g166)) + ((g609) & (g610) & (g611) & (!g612) & (!g165) & (!g166)) + ((g609) & (g610) & (g611) & (!g612) & (!g165) & (g166)) + ((g609) & (g610) & (g611) & (!g612) & (g165) & (!g166)) + ((g609) & (g610) & (g611) & (g612) & (!g165) & (!g166)) + ((g609) & (g610) & (g611) & (g612) & (!g165) & (g166)) + ((g609) & (g610) & (g611) & (g612) & (g165) & (!g166)) + ((g609) & (g610) & (g611) & (g612) & (g165) & (g166)));
	assign g4329 = (((!g2177) & (!sk[40]) & (!g2431) & (g614)) + ((!g2177) & (!sk[40]) & (g2431) & (!g614)) + ((!g2177) & (!sk[40]) & (g2431) & (g614)) + ((!g2177) & (sk[40]) & (!g2431) & (g614)) + ((!g2177) & (sk[40]) & (g2431) & (g614)) + ((g2177) & (!sk[40]) & (!g2431) & (g614)) + ((g2177) & (!sk[40]) & (g2431) & (!g614)) + ((g2177) & (!sk[40]) & (g2431) & (g614)) + ((g2177) & (sk[40]) & (g2431) & (!g614)) + ((g2177) & (sk[40]) & (g2431) & (g614)));
	assign g4330 = (((!sk[41]) & (!g2178) & (!g2431) & (g615)) + ((!sk[41]) & (!g2178) & (g2431) & (!g615)) + ((!sk[41]) & (!g2178) & (g2431) & (g615)) + ((!sk[41]) & (g2178) & (!g2431) & (g615)) + ((!sk[41]) & (g2178) & (g2431) & (!g615)) + ((!sk[41]) & (g2178) & (g2431) & (g615)) + ((sk[41]) & (!g2178) & (!g2431) & (g615)) + ((sk[41]) & (!g2178) & (g2431) & (g615)) + ((sk[41]) & (g2178) & (g2431) & (!g615)) + ((sk[41]) & (g2178) & (g2431) & (g615)));
	assign g4331 = (((!sk[42]) & (!g2179) & (!g2431) & (g616)) + ((!sk[42]) & (!g2179) & (g2431) & (!g616)) + ((!sk[42]) & (!g2179) & (g2431) & (g616)) + ((!sk[42]) & (g2179) & (!g2431) & (g616)) + ((!sk[42]) & (g2179) & (g2431) & (!g616)) + ((!sk[42]) & (g2179) & (g2431) & (g616)) + ((sk[42]) & (!g2179) & (!g2431) & (g616)) + ((sk[42]) & (!g2179) & (g2431) & (g616)) + ((sk[42]) & (g2179) & (g2431) & (!g616)) + ((sk[42]) & (g2179) & (g2431) & (g616)));
	assign g617 = (((!g165) & (!g166) & (!sk[43]) & (!g614) & (g615) & (!g616)) + ((!g165) & (!g166) & (!sk[43]) & (!g614) & (g615) & (g616)) + ((!g165) & (!g166) & (!sk[43]) & (g614) & (!g615) & (!g616)) + ((!g165) & (!g166) & (!sk[43]) & (g614) & (!g615) & (g616)) + ((!g165) & (!g166) & (!sk[43]) & (g614) & (g615) & (!g616)) + ((!g165) & (!g166) & (!sk[43]) & (g614) & (g615) & (g616)) + ((!g165) & (g166) & (!sk[43]) & (!g614) & (!g615) & (!g616)) + ((!g165) & (g166) & (!sk[43]) & (!g614) & (!g615) & (g616)) + ((!g165) & (g166) & (!sk[43]) & (!g614) & (g615) & (!g616)) + ((!g165) & (g166) & (!sk[43]) & (!g614) & (g615) & (g616)) + ((!g165) & (g166) & (!sk[43]) & (g614) & (!g615) & (!g616)) + ((!g165) & (g166) & (!sk[43]) & (g614) & (!g615) & (g616)) + ((!g165) & (g166) & (!sk[43]) & (g614) & (g615) & (!g616)) + ((!g165) & (g166) & (!sk[43]) & (g614) & (g615) & (g616)) + ((!g165) & (g166) & (sk[43]) & (!g614) & (!g615) & (g616)) + ((!g165) & (g166) & (sk[43]) & (!g614) & (g615) & (g616)) + ((!g165) & (g166) & (sk[43]) & (g614) & (!g615) & (g616)) + ((!g165) & (g166) & (sk[43]) & (g614) & (g615) & (g616)) + ((g165) & (!g166) & (!sk[43]) & (!g614) & (g615) & (!g616)) + ((g165) & (!g166) & (!sk[43]) & (!g614) & (g615) & (g616)) + ((g165) & (!g166) & (!sk[43]) & (g614) & (!g615) & (!g616)) + ((g165) & (!g166) & (!sk[43]) & (g614) & (!g615) & (g616)) + ((g165) & (!g166) & (!sk[43]) & (g614) & (g615) & (!g616)) + ((g165) & (!g166) & (!sk[43]) & (g614) & (g615) & (g616)) + ((g165) & (!g166) & (sk[43]) & (g614) & (!g615) & (!g616)) + ((g165) & (!g166) & (sk[43]) & (g614) & (!g615) & (g616)) + ((g165) & (!g166) & (sk[43]) & (g614) & (g615) & (!g616)) + ((g165) & (!g166) & (sk[43]) & (g614) & (g615) & (g616)) + ((g165) & (g166) & (!sk[43]) & (!g614) & (!g615) & (!g616)) + ((g165) & (g166) & (!sk[43]) & (!g614) & (!g615) & (g616)) + ((g165) & (g166) & (!sk[43]) & (!g614) & (g615) & (!g616)) + ((g165) & (g166) & (!sk[43]) & (!g614) & (g615) & (g616)) + ((g165) & (g166) & (!sk[43]) & (g614) & (!g615) & (!g616)) + ((g165) & (g166) & (!sk[43]) & (g614) & (!g615) & (g616)) + ((g165) & (g166) & (!sk[43]) & (g614) & (g615) & (!g616)) + ((g165) & (g166) & (!sk[43]) & (g614) & (g615) & (g616)) + ((g165) & (g166) & (sk[43]) & (!g614) & (g615) & (!g616)) + ((g165) & (g166) & (sk[43]) & (!g614) & (g615) & (g616)) + ((g165) & (g166) & (sk[43]) & (g614) & (g615) & (!g616)) + ((g165) & (g166) & (sk[43]) & (g614) & (g615) & (g616)));
	assign g4332 = (((!g2162) & (!g2431) & (!sk[44]) & (g618)) + ((!g2162) & (!g2431) & (sk[44]) & (g618)) + ((!g2162) & (g2431) & (!sk[44]) & (!g618)) + ((!g2162) & (g2431) & (!sk[44]) & (g618)) + ((!g2162) & (g2431) & (sk[44]) & (g618)) + ((g2162) & (!g2431) & (!sk[44]) & (g618)) + ((g2162) & (g2431) & (!sk[44]) & (!g618)) + ((g2162) & (g2431) & (!sk[44]) & (g618)) + ((g2162) & (g2431) & (sk[44]) & (!g618)) + ((g2162) & (g2431) & (sk[44]) & (g618)));
	assign g4333 = (((!sk[45]) & (!g2164) & (!g2431) & (g619)) + ((!sk[45]) & (!g2164) & (g2431) & (!g619)) + ((!sk[45]) & (!g2164) & (g2431) & (g619)) + ((!sk[45]) & (g2164) & (!g2431) & (g619)) + ((!sk[45]) & (g2164) & (g2431) & (!g619)) + ((!sk[45]) & (g2164) & (g2431) & (g619)) + ((sk[45]) & (!g2164) & (!g2431) & (g619)) + ((sk[45]) & (!g2164) & (g2431) & (g619)) + ((sk[45]) & (g2164) & (g2431) & (!g619)) + ((sk[45]) & (g2164) & (g2431) & (g619)));
	assign g4334 = (((!g2166) & (!sk[46]) & (!g2431) & (g620)) + ((!g2166) & (!sk[46]) & (g2431) & (!g620)) + ((!g2166) & (!sk[46]) & (g2431) & (g620)) + ((!g2166) & (sk[46]) & (!g2431) & (g620)) + ((!g2166) & (sk[46]) & (g2431) & (g620)) + ((g2166) & (!sk[46]) & (!g2431) & (g620)) + ((g2166) & (!sk[46]) & (g2431) & (!g620)) + ((g2166) & (!sk[46]) & (g2431) & (g620)) + ((g2166) & (sk[46]) & (g2431) & (!g620)) + ((g2166) & (sk[46]) & (g2431) & (g620)));
	assign g4335 = (((!sk[47]) & (!g2168) & (!g2431) & (g621)) + ((!sk[47]) & (!g2168) & (g2431) & (!g621)) + ((!sk[47]) & (!g2168) & (g2431) & (g621)) + ((!sk[47]) & (g2168) & (!g2431) & (g621)) + ((!sk[47]) & (g2168) & (g2431) & (!g621)) + ((!sk[47]) & (g2168) & (g2431) & (g621)) + ((sk[47]) & (!g2168) & (!g2431) & (g621)) + ((sk[47]) & (!g2168) & (g2431) & (g621)) + ((sk[47]) & (g2168) & (g2431) & (!g621)) + ((sk[47]) & (g2168) & (g2431) & (g621)));
	assign g622 = (((!g618) & (!g619) & (!g620) & (g621) & (g165) & (g166)) + ((!g618) & (!g619) & (g620) & (!g621) & (!g165) & (g166)) + ((!g618) & (!g619) & (g620) & (g621) & (!g165) & (g166)) + ((!g618) & (!g619) & (g620) & (g621) & (g165) & (g166)) + ((!g618) & (g619) & (!g620) & (!g621) & (g165) & (!g166)) + ((!g618) & (g619) & (!g620) & (g621) & (g165) & (!g166)) + ((!g618) & (g619) & (!g620) & (g621) & (g165) & (g166)) + ((!g618) & (g619) & (g620) & (!g621) & (!g165) & (g166)) + ((!g618) & (g619) & (g620) & (!g621) & (g165) & (!g166)) + ((!g618) & (g619) & (g620) & (g621) & (!g165) & (g166)) + ((!g618) & (g619) & (g620) & (g621) & (g165) & (!g166)) + ((!g618) & (g619) & (g620) & (g621) & (g165) & (g166)) + ((g618) & (!g619) & (!g620) & (!g621) & (!g165) & (!g166)) + ((g618) & (!g619) & (!g620) & (g621) & (!g165) & (!g166)) + ((g618) & (!g619) & (!g620) & (g621) & (g165) & (g166)) + ((g618) & (!g619) & (g620) & (!g621) & (!g165) & (!g166)) + ((g618) & (!g619) & (g620) & (!g621) & (!g165) & (g166)) + ((g618) & (!g619) & (g620) & (g621) & (!g165) & (!g166)) + ((g618) & (!g619) & (g620) & (g621) & (!g165) & (g166)) + ((g618) & (!g619) & (g620) & (g621) & (g165) & (g166)) + ((g618) & (g619) & (!g620) & (!g621) & (!g165) & (!g166)) + ((g618) & (g619) & (!g620) & (!g621) & (g165) & (!g166)) + ((g618) & (g619) & (!g620) & (g621) & (!g165) & (!g166)) + ((g618) & (g619) & (!g620) & (g621) & (g165) & (!g166)) + ((g618) & (g619) & (!g620) & (g621) & (g165) & (g166)) + ((g618) & (g619) & (g620) & (!g621) & (!g165) & (!g166)) + ((g618) & (g619) & (g620) & (!g621) & (!g165) & (g166)) + ((g618) & (g619) & (g620) & (!g621) & (g165) & (!g166)) + ((g618) & (g619) & (g620) & (g621) & (!g165) & (!g166)) + ((g618) & (g619) & (g620) & (g621) & (!g165) & (g166)) + ((g618) & (g619) & (g620) & (g621) & (g165) & (!g166)) + ((g618) & (g619) & (g620) & (g621) & (g165) & (g166)));
	assign g4336 = (((!g2169) & (!sk[49]) & (!g2431) & (g623)) + ((!g2169) & (!sk[49]) & (g2431) & (!g623)) + ((!g2169) & (!sk[49]) & (g2431) & (g623)) + ((!g2169) & (sk[49]) & (!g2431) & (g623)) + ((!g2169) & (sk[49]) & (g2431) & (g623)) + ((g2169) & (!sk[49]) & (!g2431) & (g623)) + ((g2169) & (!sk[49]) & (g2431) & (!g623)) + ((g2169) & (!sk[49]) & (g2431) & (g623)) + ((g2169) & (sk[49]) & (g2431) & (!g623)) + ((g2169) & (sk[49]) & (g2431) & (g623)));
	assign g4337 = (((!g2170) & (!sk[50]) & (!g2431) & (g624)) + ((!g2170) & (!sk[50]) & (g2431) & (!g624)) + ((!g2170) & (!sk[50]) & (g2431) & (g624)) + ((!g2170) & (sk[50]) & (!g2431) & (g624)) + ((!g2170) & (sk[50]) & (g2431) & (g624)) + ((g2170) & (!sk[50]) & (!g2431) & (g624)) + ((g2170) & (!sk[50]) & (g2431) & (!g624)) + ((g2170) & (!sk[50]) & (g2431) & (g624)) + ((g2170) & (sk[50]) & (g2431) & (!g624)) + ((g2170) & (sk[50]) & (g2431) & (g624)));
	assign g4338 = (((!g2171) & (!g2431) & (!sk[51]) & (g625)) + ((!g2171) & (!g2431) & (sk[51]) & (g625)) + ((!g2171) & (g2431) & (!sk[51]) & (!g625)) + ((!g2171) & (g2431) & (!sk[51]) & (g625)) + ((!g2171) & (g2431) & (sk[51]) & (g625)) + ((g2171) & (!g2431) & (!sk[51]) & (g625)) + ((g2171) & (g2431) & (!sk[51]) & (!g625)) + ((g2171) & (g2431) & (!sk[51]) & (g625)) + ((g2171) & (g2431) & (sk[51]) & (!g625)) + ((g2171) & (g2431) & (sk[51]) & (g625)));
	assign g4339 = (((!sk[52]) & (!g2172) & (!g2431) & (g626)) + ((!sk[52]) & (!g2172) & (g2431) & (!g626)) + ((!sk[52]) & (!g2172) & (g2431) & (g626)) + ((!sk[52]) & (g2172) & (!g2431) & (g626)) + ((!sk[52]) & (g2172) & (g2431) & (!g626)) + ((!sk[52]) & (g2172) & (g2431) & (g626)) + ((sk[52]) & (!g2172) & (!g2431) & (g626)) + ((sk[52]) & (!g2172) & (g2431) & (g626)) + ((sk[52]) & (g2172) & (g2431) & (!g626)) + ((sk[52]) & (g2172) & (g2431) & (g626)));
	assign g627 = (((!g623) & (!g624) & (!g625) & (g626) & (g165) & (g166)) + ((!g623) & (!g624) & (g625) & (!g626) & (!g165) & (g166)) + ((!g623) & (!g624) & (g625) & (g626) & (!g165) & (g166)) + ((!g623) & (!g624) & (g625) & (g626) & (g165) & (g166)) + ((!g623) & (g624) & (!g625) & (!g626) & (g165) & (!g166)) + ((!g623) & (g624) & (!g625) & (g626) & (g165) & (!g166)) + ((!g623) & (g624) & (!g625) & (g626) & (g165) & (g166)) + ((!g623) & (g624) & (g625) & (!g626) & (!g165) & (g166)) + ((!g623) & (g624) & (g625) & (!g626) & (g165) & (!g166)) + ((!g623) & (g624) & (g625) & (g626) & (!g165) & (g166)) + ((!g623) & (g624) & (g625) & (g626) & (g165) & (!g166)) + ((!g623) & (g624) & (g625) & (g626) & (g165) & (g166)) + ((g623) & (!g624) & (!g625) & (!g626) & (!g165) & (!g166)) + ((g623) & (!g624) & (!g625) & (g626) & (!g165) & (!g166)) + ((g623) & (!g624) & (!g625) & (g626) & (g165) & (g166)) + ((g623) & (!g624) & (g625) & (!g626) & (!g165) & (!g166)) + ((g623) & (!g624) & (g625) & (!g626) & (!g165) & (g166)) + ((g623) & (!g624) & (g625) & (g626) & (!g165) & (!g166)) + ((g623) & (!g624) & (g625) & (g626) & (!g165) & (g166)) + ((g623) & (!g624) & (g625) & (g626) & (g165) & (g166)) + ((g623) & (g624) & (!g625) & (!g626) & (!g165) & (!g166)) + ((g623) & (g624) & (!g625) & (!g626) & (g165) & (!g166)) + ((g623) & (g624) & (!g625) & (g626) & (!g165) & (!g166)) + ((g623) & (g624) & (!g625) & (g626) & (g165) & (!g166)) + ((g623) & (g624) & (!g625) & (g626) & (g165) & (g166)) + ((g623) & (g624) & (g625) & (!g626) & (!g165) & (!g166)) + ((g623) & (g624) & (g625) & (!g626) & (!g165) & (g166)) + ((g623) & (g624) & (g625) & (!g626) & (g165) & (!g166)) + ((g623) & (g624) & (g625) & (g626) & (!g165) & (!g166)) + ((g623) & (g624) & (g625) & (g626) & (!g165) & (g166)) + ((g623) & (g624) & (g625) & (g626) & (g165) & (!g166)) + ((g623) & (g624) & (g625) & (g626) & (g165) & (g166)));
	assign g628 = (((!g147) & (!g148) & (!g613) & (g617) & (!g622) & (!g627)) + ((!g147) & (!g148) & (!g613) & (g617) & (!g622) & (g627)) + ((!g147) & (!g148) & (!g613) & (g617) & (g622) & (!g627)) + ((!g147) & (!g148) & (!g613) & (g617) & (g622) & (g627)) + ((!g147) & (!g148) & (g613) & (g617) & (!g622) & (!g627)) + ((!g147) & (!g148) & (g613) & (g617) & (!g622) & (g627)) + ((!g147) & (!g148) & (g613) & (g617) & (g622) & (!g627)) + ((!g147) & (!g148) & (g613) & (g617) & (g622) & (g627)) + ((!g147) & (g148) & (!g613) & (!g617) & (!g622) & (g627)) + ((!g147) & (g148) & (!g613) & (!g617) & (g622) & (g627)) + ((!g147) & (g148) & (!g613) & (g617) & (!g622) & (g627)) + ((!g147) & (g148) & (!g613) & (g617) & (g622) & (g627)) + ((!g147) & (g148) & (g613) & (!g617) & (!g622) & (g627)) + ((!g147) & (g148) & (g613) & (!g617) & (g622) & (g627)) + ((!g147) & (g148) & (g613) & (g617) & (!g622) & (g627)) + ((!g147) & (g148) & (g613) & (g617) & (g622) & (g627)) + ((g147) & (!g148) & (g613) & (!g617) & (!g622) & (!g627)) + ((g147) & (!g148) & (g613) & (!g617) & (!g622) & (g627)) + ((g147) & (!g148) & (g613) & (!g617) & (g622) & (!g627)) + ((g147) & (!g148) & (g613) & (!g617) & (g622) & (g627)) + ((g147) & (!g148) & (g613) & (g617) & (!g622) & (!g627)) + ((g147) & (!g148) & (g613) & (g617) & (!g622) & (g627)) + ((g147) & (!g148) & (g613) & (g617) & (g622) & (!g627)) + ((g147) & (!g148) & (g613) & (g617) & (g622) & (g627)) + ((g147) & (g148) & (!g613) & (!g617) & (g622) & (!g627)) + ((g147) & (g148) & (!g613) & (!g617) & (g622) & (g627)) + ((g147) & (g148) & (!g613) & (g617) & (g622) & (!g627)) + ((g147) & (g148) & (!g613) & (g617) & (g622) & (g627)) + ((g147) & (g148) & (g613) & (!g617) & (g622) & (!g627)) + ((g147) & (g148) & (g613) & (!g617) & (g622) & (g627)) + ((g147) & (g148) & (g613) & (g617) & (g622) & (!g627)) + ((g147) & (g148) & (g613) & (g617) & (g622) & (g627)));
	assign g629 = (((!g142) & (!sk[55]) & (!g608) & (g628)) + ((!g142) & (!sk[55]) & (g608) & (!g628)) + ((!g142) & (!sk[55]) & (g608) & (g628)) + ((!g142) & (sk[55]) & (!g608) & (g628)) + ((!g142) & (sk[55]) & (g608) & (g628)) + ((g142) & (!sk[55]) & (!g608) & (g628)) + ((g142) & (!sk[55]) & (g608) & (!g628)) + ((g142) & (!sk[55]) & (g608) & (g628)) + ((g142) & (sk[55]) & (g608) & (!g628)) + ((g142) & (sk[55]) & (g608) & (g628)));
	assign g4340 = (((!g2059) & (!sk[56]) & (!g3627) & (g630)) + ((!g2059) & (!sk[56]) & (g3627) & (!g630)) + ((!g2059) & (!sk[56]) & (g3627) & (g630)) + ((!g2059) & (sk[56]) & (!g3627) & (g630)) + ((!g2059) & (sk[56]) & (g3627) & (g630)) + ((g2059) & (!sk[56]) & (!g3627) & (g630)) + ((g2059) & (!sk[56]) & (g3627) & (!g630)) + ((g2059) & (!sk[56]) & (g3627) & (g630)) + ((g2059) & (sk[56]) & (g3627) & (!g630)) + ((g2059) & (sk[56]) & (g3627) & (g630)));
	assign g4341 = (((!g2140) & (!g2454) & (!sk[57]) & (g631)) + ((!g2140) & (!g2454) & (sk[57]) & (g631)) + ((!g2140) & (g2454) & (!sk[57]) & (!g631)) + ((!g2140) & (g2454) & (!sk[57]) & (g631)) + ((!g2140) & (g2454) & (sk[57]) & (g631)) + ((g2140) & (!g2454) & (!sk[57]) & (g631)) + ((g2140) & (g2454) & (!sk[57]) & (!g631)) + ((g2140) & (g2454) & (!sk[57]) & (g631)) + ((g2140) & (g2454) & (sk[57]) & (!g631)) + ((g2140) & (g2454) & (sk[57]) & (g631)));
	assign g4342 = (((!g2142) & (!sk[58]) & (!g2454) & (g632)) + ((!g2142) & (!sk[58]) & (g2454) & (!g632)) + ((!g2142) & (!sk[58]) & (g2454) & (g632)) + ((!g2142) & (sk[58]) & (!g2454) & (g632)) + ((!g2142) & (sk[58]) & (g2454) & (g632)) + ((g2142) & (!sk[58]) & (!g2454) & (g632)) + ((g2142) & (!sk[58]) & (g2454) & (!g632)) + ((g2142) & (!sk[58]) & (g2454) & (g632)) + ((g2142) & (sk[58]) & (g2454) & (!g632)) + ((g2142) & (sk[58]) & (g2454) & (g632)));
	assign g4343 = (((!g2144) & (!sk[59]) & (!g2454) & (g633)) + ((!g2144) & (!sk[59]) & (g2454) & (!g633)) + ((!g2144) & (!sk[59]) & (g2454) & (g633)) + ((!g2144) & (sk[59]) & (!g2454) & (g633)) + ((!g2144) & (sk[59]) & (g2454) & (g633)) + ((g2144) & (!sk[59]) & (!g2454) & (g633)) + ((g2144) & (!sk[59]) & (g2454) & (!g633)) + ((g2144) & (!sk[59]) & (g2454) & (g633)) + ((g2144) & (sk[59]) & (g2454) & (!g633)) + ((g2144) & (sk[59]) & (g2454) & (g633)));
	assign g4344 = (((!sk[60]) & (!g2145) & (!g2454) & (g634)) + ((!sk[60]) & (!g2145) & (g2454) & (!g634)) + ((!sk[60]) & (!g2145) & (g2454) & (g634)) + ((!sk[60]) & (g2145) & (!g2454) & (g634)) + ((!sk[60]) & (g2145) & (g2454) & (!g634)) + ((!sk[60]) & (g2145) & (g2454) & (g634)) + ((sk[60]) & (!g2145) & (!g2454) & (g634)) + ((sk[60]) & (!g2145) & (g2454) & (g634)) + ((sk[60]) & (g2145) & (g2454) & (!g634)) + ((sk[60]) & (g2145) & (g2454) & (g634)));
	assign g635 = (((!g631) & (!g632) & (!g633) & (g634) & (g147) & (g148)) + ((!g631) & (!g632) & (g633) & (!g634) & (!g147) & (g148)) + ((!g631) & (!g632) & (g633) & (g634) & (!g147) & (g148)) + ((!g631) & (!g632) & (g633) & (g634) & (g147) & (g148)) + ((!g631) & (g632) & (!g633) & (!g634) & (g147) & (!g148)) + ((!g631) & (g632) & (!g633) & (g634) & (g147) & (!g148)) + ((!g631) & (g632) & (!g633) & (g634) & (g147) & (g148)) + ((!g631) & (g632) & (g633) & (!g634) & (!g147) & (g148)) + ((!g631) & (g632) & (g633) & (!g634) & (g147) & (!g148)) + ((!g631) & (g632) & (g633) & (g634) & (!g147) & (g148)) + ((!g631) & (g632) & (g633) & (g634) & (g147) & (!g148)) + ((!g631) & (g632) & (g633) & (g634) & (g147) & (g148)) + ((g631) & (!g632) & (!g633) & (!g634) & (!g147) & (!g148)) + ((g631) & (!g632) & (!g633) & (g634) & (!g147) & (!g148)) + ((g631) & (!g632) & (!g633) & (g634) & (g147) & (g148)) + ((g631) & (!g632) & (g633) & (!g634) & (!g147) & (!g148)) + ((g631) & (!g632) & (g633) & (!g634) & (!g147) & (g148)) + ((g631) & (!g632) & (g633) & (g634) & (!g147) & (!g148)) + ((g631) & (!g632) & (g633) & (g634) & (!g147) & (g148)) + ((g631) & (!g632) & (g633) & (g634) & (g147) & (g148)) + ((g631) & (g632) & (!g633) & (!g634) & (!g147) & (!g148)) + ((g631) & (g632) & (!g633) & (!g634) & (g147) & (!g148)) + ((g631) & (g632) & (!g633) & (g634) & (!g147) & (!g148)) + ((g631) & (g632) & (!g633) & (g634) & (g147) & (!g148)) + ((g631) & (g632) & (!g633) & (g634) & (g147) & (g148)) + ((g631) & (g632) & (g633) & (!g634) & (!g147) & (!g148)) + ((g631) & (g632) & (g633) & (!g634) & (!g147) & (g148)) + ((g631) & (g632) & (g633) & (!g634) & (g147) & (!g148)) + ((g631) & (g632) & (g633) & (g634) & (!g147) & (!g148)) + ((g631) & (g632) & (g633) & (g634) & (!g147) & (g148)) + ((g631) & (g632) & (g633) & (g634) & (g147) & (!g148)) + ((g631) & (g632) & (g633) & (g634) & (g147) & (g148)));
	assign g4345 = (((!g2146) & (!sk[62]) & (!g2454) & (g636)) + ((!g2146) & (!sk[62]) & (g2454) & (!g636)) + ((!g2146) & (!sk[62]) & (g2454) & (g636)) + ((!g2146) & (sk[62]) & (!g2454) & (g636)) + ((!g2146) & (sk[62]) & (g2454) & (g636)) + ((g2146) & (!sk[62]) & (!g2454) & (g636)) + ((g2146) & (!sk[62]) & (g2454) & (!g636)) + ((g2146) & (!sk[62]) & (g2454) & (g636)) + ((g2146) & (sk[62]) & (g2454) & (!g636)) + ((g2146) & (sk[62]) & (g2454) & (g636)));
	assign g4346 = (((!g2148) & (!sk[63]) & (!g2454) & (g637)) + ((!g2148) & (!sk[63]) & (g2454) & (!g637)) + ((!g2148) & (!sk[63]) & (g2454) & (g637)) + ((!g2148) & (sk[63]) & (!g2454) & (g637)) + ((!g2148) & (sk[63]) & (g2454) & (g637)) + ((g2148) & (!sk[63]) & (!g2454) & (g637)) + ((g2148) & (!sk[63]) & (g2454) & (!g637)) + ((g2148) & (!sk[63]) & (g2454) & (g637)) + ((g2148) & (sk[63]) & (g2454) & (!g637)) + ((g2148) & (sk[63]) & (g2454) & (g637)));
	assign g4347 = (((!sk[64]) & (!g2150) & (!g2454) & (g638)) + ((!sk[64]) & (!g2150) & (g2454) & (!g638)) + ((!sk[64]) & (!g2150) & (g2454) & (g638)) + ((!sk[64]) & (g2150) & (!g2454) & (g638)) + ((!sk[64]) & (g2150) & (g2454) & (!g638)) + ((!sk[64]) & (g2150) & (g2454) & (g638)) + ((sk[64]) & (!g2150) & (!g2454) & (g638)) + ((sk[64]) & (!g2150) & (g2454) & (g638)) + ((sk[64]) & (g2150) & (g2454) & (!g638)) + ((sk[64]) & (g2150) & (g2454) & (g638)));
	assign g4348 = (((!sk[65]) & (!g2151) & (!g2454) & (g639)) + ((!sk[65]) & (!g2151) & (g2454) & (!g639)) + ((!sk[65]) & (!g2151) & (g2454) & (g639)) + ((!sk[65]) & (g2151) & (!g2454) & (g639)) + ((!sk[65]) & (g2151) & (g2454) & (!g639)) + ((!sk[65]) & (g2151) & (g2454) & (g639)) + ((sk[65]) & (!g2151) & (!g2454) & (g639)) + ((sk[65]) & (!g2151) & (g2454) & (g639)) + ((sk[65]) & (g2151) & (g2454) & (!g639)) + ((sk[65]) & (g2151) & (g2454) & (g639)));
	assign g640 = (((!g636) & (!g637) & (!g638) & (g639) & (g147) & (g148)) + ((!g636) & (!g637) & (g638) & (!g639) & (!g147) & (g148)) + ((!g636) & (!g637) & (g638) & (g639) & (!g147) & (g148)) + ((!g636) & (!g637) & (g638) & (g639) & (g147) & (g148)) + ((!g636) & (g637) & (!g638) & (!g639) & (g147) & (!g148)) + ((!g636) & (g637) & (!g638) & (g639) & (g147) & (!g148)) + ((!g636) & (g637) & (!g638) & (g639) & (g147) & (g148)) + ((!g636) & (g637) & (g638) & (!g639) & (!g147) & (g148)) + ((!g636) & (g637) & (g638) & (!g639) & (g147) & (!g148)) + ((!g636) & (g637) & (g638) & (g639) & (!g147) & (g148)) + ((!g636) & (g637) & (g638) & (g639) & (g147) & (!g148)) + ((!g636) & (g637) & (g638) & (g639) & (g147) & (g148)) + ((g636) & (!g637) & (!g638) & (!g639) & (!g147) & (!g148)) + ((g636) & (!g637) & (!g638) & (g639) & (!g147) & (!g148)) + ((g636) & (!g637) & (!g638) & (g639) & (g147) & (g148)) + ((g636) & (!g637) & (g638) & (!g639) & (!g147) & (!g148)) + ((g636) & (!g637) & (g638) & (!g639) & (!g147) & (g148)) + ((g636) & (!g637) & (g638) & (g639) & (!g147) & (!g148)) + ((g636) & (!g637) & (g638) & (g639) & (!g147) & (g148)) + ((g636) & (!g637) & (g638) & (g639) & (g147) & (g148)) + ((g636) & (g637) & (!g638) & (!g639) & (!g147) & (!g148)) + ((g636) & (g637) & (!g638) & (!g639) & (g147) & (!g148)) + ((g636) & (g637) & (!g638) & (g639) & (!g147) & (!g148)) + ((g636) & (g637) & (!g638) & (g639) & (g147) & (!g148)) + ((g636) & (g637) & (!g638) & (g639) & (g147) & (g148)) + ((g636) & (g637) & (g638) & (!g639) & (!g147) & (!g148)) + ((g636) & (g637) & (g638) & (!g639) & (!g147) & (g148)) + ((g636) & (g637) & (g638) & (!g639) & (g147) & (!g148)) + ((g636) & (g637) & (g638) & (g639) & (!g147) & (!g148)) + ((g636) & (g637) & (g638) & (g639) & (!g147) & (g148)) + ((g636) & (g637) & (g638) & (g639) & (g147) & (!g148)) + ((g636) & (g637) & (g638) & (g639) & (g147) & (g148)));
	assign g4349 = (((!sk[67]) & (!g2152) & (!g2454) & (g641)) + ((!sk[67]) & (!g2152) & (g2454) & (!g641)) + ((!sk[67]) & (!g2152) & (g2454) & (g641)) + ((!sk[67]) & (g2152) & (!g2454) & (g641)) + ((!sk[67]) & (g2152) & (g2454) & (!g641)) + ((!sk[67]) & (g2152) & (g2454) & (g641)) + ((sk[67]) & (!g2152) & (!g2454) & (g641)) + ((sk[67]) & (!g2152) & (g2454) & (g641)) + ((sk[67]) & (g2152) & (g2454) & (!g641)) + ((sk[67]) & (g2152) & (g2454) & (g641)));
	assign g4350 = (((!g2153) & (!sk[68]) & (!g2454) & (g642)) + ((!g2153) & (!sk[68]) & (g2454) & (!g642)) + ((!g2153) & (!sk[68]) & (g2454) & (g642)) + ((!g2153) & (sk[68]) & (!g2454) & (g642)) + ((!g2153) & (sk[68]) & (g2454) & (g642)) + ((g2153) & (!sk[68]) & (!g2454) & (g642)) + ((g2153) & (!sk[68]) & (g2454) & (!g642)) + ((g2153) & (!sk[68]) & (g2454) & (g642)) + ((g2153) & (sk[68]) & (g2454) & (!g642)) + ((g2153) & (sk[68]) & (g2454) & (g642)));
	assign g4351 = (((!g2155) & (!g2454) & (!sk[69]) & (g643)) + ((!g2155) & (!g2454) & (sk[69]) & (g643)) + ((!g2155) & (g2454) & (!sk[69]) & (!g643)) + ((!g2155) & (g2454) & (!sk[69]) & (g643)) + ((!g2155) & (g2454) & (sk[69]) & (g643)) + ((g2155) & (!g2454) & (!sk[69]) & (g643)) + ((g2155) & (g2454) & (!sk[69]) & (!g643)) + ((g2155) & (g2454) & (!sk[69]) & (g643)) + ((g2155) & (g2454) & (sk[69]) & (!g643)) + ((g2155) & (g2454) & (sk[69]) & (g643)));
	assign g4352 = (((!g2157) & (!sk[70]) & (!g2454) & (g644)) + ((!g2157) & (!sk[70]) & (g2454) & (!g644)) + ((!g2157) & (!sk[70]) & (g2454) & (g644)) + ((!g2157) & (sk[70]) & (!g2454) & (g644)) + ((!g2157) & (sk[70]) & (g2454) & (g644)) + ((g2157) & (!sk[70]) & (!g2454) & (g644)) + ((g2157) & (!sk[70]) & (g2454) & (!g644)) + ((g2157) & (!sk[70]) & (g2454) & (g644)) + ((g2157) & (sk[70]) & (g2454) & (!g644)) + ((g2157) & (sk[70]) & (g2454) & (g644)));
	assign g645 = (((!g641) & (!g642) & (!g643) & (g644) & (g147) & (g148)) + ((!g641) & (!g642) & (g643) & (!g644) & (!g147) & (g148)) + ((!g641) & (!g642) & (g643) & (g644) & (!g147) & (g148)) + ((!g641) & (!g642) & (g643) & (g644) & (g147) & (g148)) + ((!g641) & (g642) & (!g643) & (!g644) & (g147) & (!g148)) + ((!g641) & (g642) & (!g643) & (g644) & (g147) & (!g148)) + ((!g641) & (g642) & (!g643) & (g644) & (g147) & (g148)) + ((!g641) & (g642) & (g643) & (!g644) & (!g147) & (g148)) + ((!g641) & (g642) & (g643) & (!g644) & (g147) & (!g148)) + ((!g641) & (g642) & (g643) & (g644) & (!g147) & (g148)) + ((!g641) & (g642) & (g643) & (g644) & (g147) & (!g148)) + ((!g641) & (g642) & (g643) & (g644) & (g147) & (g148)) + ((g641) & (!g642) & (!g643) & (!g644) & (!g147) & (!g148)) + ((g641) & (!g642) & (!g643) & (g644) & (!g147) & (!g148)) + ((g641) & (!g642) & (!g643) & (g644) & (g147) & (g148)) + ((g641) & (!g642) & (g643) & (!g644) & (!g147) & (!g148)) + ((g641) & (!g642) & (g643) & (!g644) & (!g147) & (g148)) + ((g641) & (!g642) & (g643) & (g644) & (!g147) & (!g148)) + ((g641) & (!g642) & (g643) & (g644) & (!g147) & (g148)) + ((g641) & (!g642) & (g643) & (g644) & (g147) & (g148)) + ((g641) & (g642) & (!g643) & (!g644) & (!g147) & (!g148)) + ((g641) & (g642) & (!g643) & (!g644) & (g147) & (!g148)) + ((g641) & (g642) & (!g643) & (g644) & (!g147) & (!g148)) + ((g641) & (g642) & (!g643) & (g644) & (g147) & (!g148)) + ((g641) & (g642) & (!g643) & (g644) & (g147) & (g148)) + ((g641) & (g642) & (g643) & (!g644) & (!g147) & (!g148)) + ((g641) & (g642) & (g643) & (!g644) & (!g147) & (g148)) + ((g641) & (g642) & (g643) & (!g644) & (g147) & (!g148)) + ((g641) & (g642) & (g643) & (g644) & (!g147) & (!g148)) + ((g641) & (g642) & (g643) & (g644) & (!g147) & (g148)) + ((g641) & (g642) & (g643) & (g644) & (g147) & (!g148)) + ((g641) & (g642) & (g643) & (g644) & (g147) & (g148)));
	assign g4353 = (((!sk[72]) & (!g2158) & (!g2454) & (g646)) + ((!sk[72]) & (!g2158) & (g2454) & (!g646)) + ((!sk[72]) & (!g2158) & (g2454) & (g646)) + ((!sk[72]) & (g2158) & (!g2454) & (g646)) + ((!sk[72]) & (g2158) & (g2454) & (!g646)) + ((!sk[72]) & (g2158) & (g2454) & (g646)) + ((sk[72]) & (!g2158) & (!g2454) & (g646)) + ((sk[72]) & (!g2158) & (g2454) & (g646)) + ((sk[72]) & (g2158) & (g2454) & (!g646)) + ((sk[72]) & (g2158) & (g2454) & (g646)));
	assign g4354 = (((!sk[73]) & (!g2159) & (!g2454) & (g647)) + ((!sk[73]) & (!g2159) & (g2454) & (!g647)) + ((!sk[73]) & (!g2159) & (g2454) & (g647)) + ((!sk[73]) & (g2159) & (!g2454) & (g647)) + ((!sk[73]) & (g2159) & (g2454) & (!g647)) + ((!sk[73]) & (g2159) & (g2454) & (g647)) + ((sk[73]) & (!g2159) & (!g2454) & (g647)) + ((sk[73]) & (!g2159) & (g2454) & (g647)) + ((sk[73]) & (g2159) & (g2454) & (!g647)) + ((sk[73]) & (g2159) & (g2454) & (g647)));
	assign g4355 = (((!sk[74]) & (!g2160) & (!g2454) & (g648)) + ((!sk[74]) & (!g2160) & (g2454) & (!g648)) + ((!sk[74]) & (!g2160) & (g2454) & (g648)) + ((!sk[74]) & (g2160) & (!g2454) & (g648)) + ((!sk[74]) & (g2160) & (g2454) & (!g648)) + ((!sk[74]) & (g2160) & (g2454) & (g648)) + ((sk[74]) & (!g2160) & (!g2454) & (g648)) + ((sk[74]) & (!g2160) & (g2454) & (g648)) + ((sk[74]) & (g2160) & (g2454) & (!g648)) + ((sk[74]) & (g2160) & (g2454) & (g648)));
	assign g4356 = (((!g2161) & (!sk[75]) & (!g2454) & (g649)) + ((!g2161) & (!sk[75]) & (g2454) & (!g649)) + ((!g2161) & (!sk[75]) & (g2454) & (g649)) + ((!g2161) & (sk[75]) & (!g2454) & (g649)) + ((!g2161) & (sk[75]) & (g2454) & (g649)) + ((g2161) & (!sk[75]) & (!g2454) & (g649)) + ((g2161) & (!sk[75]) & (g2454) & (!g649)) + ((g2161) & (!sk[75]) & (g2454) & (g649)) + ((g2161) & (sk[75]) & (g2454) & (!g649)) + ((g2161) & (sk[75]) & (g2454) & (g649)));
	assign g650 = (((!g646) & (!g647) & (!g648) & (g649) & (g147) & (g148)) + ((!g646) & (!g647) & (g648) & (!g649) & (!g147) & (g148)) + ((!g646) & (!g647) & (g648) & (g649) & (!g147) & (g148)) + ((!g646) & (!g647) & (g648) & (g649) & (g147) & (g148)) + ((!g646) & (g647) & (!g648) & (!g649) & (g147) & (!g148)) + ((!g646) & (g647) & (!g648) & (g649) & (g147) & (!g148)) + ((!g646) & (g647) & (!g648) & (g649) & (g147) & (g148)) + ((!g646) & (g647) & (g648) & (!g649) & (!g147) & (g148)) + ((!g646) & (g647) & (g648) & (!g649) & (g147) & (!g148)) + ((!g646) & (g647) & (g648) & (g649) & (!g147) & (g148)) + ((!g646) & (g647) & (g648) & (g649) & (g147) & (!g148)) + ((!g646) & (g647) & (g648) & (g649) & (g147) & (g148)) + ((g646) & (!g647) & (!g648) & (!g649) & (!g147) & (!g148)) + ((g646) & (!g647) & (!g648) & (g649) & (!g147) & (!g148)) + ((g646) & (!g647) & (!g648) & (g649) & (g147) & (g148)) + ((g646) & (!g647) & (g648) & (!g649) & (!g147) & (!g148)) + ((g646) & (!g647) & (g648) & (!g649) & (!g147) & (g148)) + ((g646) & (!g647) & (g648) & (g649) & (!g147) & (!g148)) + ((g646) & (!g647) & (g648) & (g649) & (!g147) & (g148)) + ((g646) & (!g647) & (g648) & (g649) & (g147) & (g148)) + ((g646) & (g647) & (!g648) & (!g649) & (!g147) & (!g148)) + ((g646) & (g647) & (!g648) & (!g649) & (g147) & (!g148)) + ((g646) & (g647) & (!g648) & (g649) & (!g147) & (!g148)) + ((g646) & (g647) & (!g648) & (g649) & (g147) & (!g148)) + ((g646) & (g647) & (!g648) & (g649) & (g147) & (g148)) + ((g646) & (g647) & (g648) & (!g649) & (!g147) & (!g148)) + ((g646) & (g647) & (g648) & (!g649) & (!g147) & (g148)) + ((g646) & (g647) & (g648) & (!g649) & (g147) & (!g148)) + ((g646) & (g647) & (g648) & (g649) & (!g147) & (!g148)) + ((g646) & (g647) & (g648) & (g649) & (!g147) & (g148)) + ((g646) & (g647) & (g648) & (g649) & (g147) & (!g148)) + ((g646) & (g647) & (g648) & (g649) & (g147) & (g148)));
	assign g651 = (((!g635) & (!g640) & (!g645) & (g650) & (g165) & (g166)) + ((!g635) & (!g640) & (g645) & (!g650) & (!g165) & (g166)) + ((!g635) & (!g640) & (g645) & (g650) & (!g165) & (g166)) + ((!g635) & (!g640) & (g645) & (g650) & (g165) & (g166)) + ((!g635) & (g640) & (!g645) & (!g650) & (g165) & (!g166)) + ((!g635) & (g640) & (!g645) & (g650) & (g165) & (!g166)) + ((!g635) & (g640) & (!g645) & (g650) & (g165) & (g166)) + ((!g635) & (g640) & (g645) & (!g650) & (!g165) & (g166)) + ((!g635) & (g640) & (g645) & (!g650) & (g165) & (!g166)) + ((!g635) & (g640) & (g645) & (g650) & (!g165) & (g166)) + ((!g635) & (g640) & (g645) & (g650) & (g165) & (!g166)) + ((!g635) & (g640) & (g645) & (g650) & (g165) & (g166)) + ((g635) & (!g640) & (!g645) & (!g650) & (!g165) & (!g166)) + ((g635) & (!g640) & (!g645) & (g650) & (!g165) & (!g166)) + ((g635) & (!g640) & (!g645) & (g650) & (g165) & (g166)) + ((g635) & (!g640) & (g645) & (!g650) & (!g165) & (!g166)) + ((g635) & (!g640) & (g645) & (!g650) & (!g165) & (g166)) + ((g635) & (!g640) & (g645) & (g650) & (!g165) & (!g166)) + ((g635) & (!g640) & (g645) & (g650) & (!g165) & (g166)) + ((g635) & (!g640) & (g645) & (g650) & (g165) & (g166)) + ((g635) & (g640) & (!g645) & (!g650) & (!g165) & (!g166)) + ((g635) & (g640) & (!g645) & (!g650) & (g165) & (!g166)) + ((g635) & (g640) & (!g645) & (g650) & (!g165) & (!g166)) + ((g635) & (g640) & (!g645) & (g650) & (g165) & (!g166)) + ((g635) & (g640) & (!g645) & (g650) & (g165) & (g166)) + ((g635) & (g640) & (g645) & (!g650) & (!g165) & (!g166)) + ((g635) & (g640) & (g645) & (!g650) & (!g165) & (g166)) + ((g635) & (g640) & (g645) & (!g650) & (g165) & (!g166)) + ((g635) & (g640) & (g645) & (g650) & (!g165) & (!g166)) + ((g635) & (g640) & (g645) & (g650) & (!g165) & (g166)) + ((g635) & (g640) & (g645) & (g650) & (g165) & (!g166)) + ((g635) & (g640) & (g645) & (g650) & (g165) & (g166)));
	assign g4357 = (((!g2173) & (!sk[78]) & (!g2454) & (g652)) + ((!g2173) & (!sk[78]) & (g2454) & (!g652)) + ((!g2173) & (!sk[78]) & (g2454) & (g652)) + ((!g2173) & (sk[78]) & (!g2454) & (g652)) + ((!g2173) & (sk[78]) & (g2454) & (g652)) + ((g2173) & (!sk[78]) & (!g2454) & (g652)) + ((g2173) & (!sk[78]) & (g2454) & (!g652)) + ((g2173) & (!sk[78]) & (g2454) & (g652)) + ((g2173) & (sk[78]) & (g2454) & (!g652)) + ((g2173) & (sk[78]) & (g2454) & (g652)));
	assign g4358 = (((!g2174) & (!sk[79]) & (!g2454) & (g653)) + ((!g2174) & (!sk[79]) & (g2454) & (!g653)) + ((!g2174) & (!sk[79]) & (g2454) & (g653)) + ((!g2174) & (sk[79]) & (!g2454) & (g653)) + ((!g2174) & (sk[79]) & (g2454) & (g653)) + ((g2174) & (!sk[79]) & (!g2454) & (g653)) + ((g2174) & (!sk[79]) & (g2454) & (!g653)) + ((g2174) & (!sk[79]) & (g2454) & (g653)) + ((g2174) & (sk[79]) & (g2454) & (!g653)) + ((g2174) & (sk[79]) & (g2454) & (g653)));
	assign g4359 = (((!g2175) & (!sk[80]) & (!g2454) & (g654)) + ((!g2175) & (!sk[80]) & (g2454) & (!g654)) + ((!g2175) & (!sk[80]) & (g2454) & (g654)) + ((!g2175) & (sk[80]) & (!g2454) & (g654)) + ((!g2175) & (sk[80]) & (g2454) & (g654)) + ((g2175) & (!sk[80]) & (!g2454) & (g654)) + ((g2175) & (!sk[80]) & (g2454) & (!g654)) + ((g2175) & (!sk[80]) & (g2454) & (g654)) + ((g2175) & (sk[80]) & (g2454) & (!g654)) + ((g2175) & (sk[80]) & (g2454) & (g654)));
	assign g4360 = (((!sk[81]) & (!g2176) & (!g2454) & (g655)) + ((!sk[81]) & (!g2176) & (g2454) & (!g655)) + ((!sk[81]) & (!g2176) & (g2454) & (g655)) + ((!sk[81]) & (g2176) & (!g2454) & (g655)) + ((!sk[81]) & (g2176) & (g2454) & (!g655)) + ((!sk[81]) & (g2176) & (g2454) & (g655)) + ((sk[81]) & (!g2176) & (!g2454) & (g655)) + ((sk[81]) & (!g2176) & (g2454) & (g655)) + ((sk[81]) & (g2176) & (g2454) & (!g655)) + ((sk[81]) & (g2176) & (g2454) & (g655)));
	assign g656 = (((!g652) & (!g653) & (!g654) & (g655) & (g165) & (g166)) + ((!g652) & (!g653) & (g654) & (!g655) & (!g165) & (g166)) + ((!g652) & (!g653) & (g654) & (g655) & (!g165) & (g166)) + ((!g652) & (!g653) & (g654) & (g655) & (g165) & (g166)) + ((!g652) & (g653) & (!g654) & (!g655) & (g165) & (!g166)) + ((!g652) & (g653) & (!g654) & (g655) & (g165) & (!g166)) + ((!g652) & (g653) & (!g654) & (g655) & (g165) & (g166)) + ((!g652) & (g653) & (g654) & (!g655) & (!g165) & (g166)) + ((!g652) & (g653) & (g654) & (!g655) & (g165) & (!g166)) + ((!g652) & (g653) & (g654) & (g655) & (!g165) & (g166)) + ((!g652) & (g653) & (g654) & (g655) & (g165) & (!g166)) + ((!g652) & (g653) & (g654) & (g655) & (g165) & (g166)) + ((g652) & (!g653) & (!g654) & (!g655) & (!g165) & (!g166)) + ((g652) & (!g653) & (!g654) & (g655) & (!g165) & (!g166)) + ((g652) & (!g653) & (!g654) & (g655) & (g165) & (g166)) + ((g652) & (!g653) & (g654) & (!g655) & (!g165) & (!g166)) + ((g652) & (!g653) & (g654) & (!g655) & (!g165) & (g166)) + ((g652) & (!g653) & (g654) & (g655) & (!g165) & (!g166)) + ((g652) & (!g653) & (g654) & (g655) & (!g165) & (g166)) + ((g652) & (!g653) & (g654) & (g655) & (g165) & (g166)) + ((g652) & (g653) & (!g654) & (!g655) & (!g165) & (!g166)) + ((g652) & (g653) & (!g654) & (!g655) & (g165) & (!g166)) + ((g652) & (g653) & (!g654) & (g655) & (!g165) & (!g166)) + ((g652) & (g653) & (!g654) & (g655) & (g165) & (!g166)) + ((g652) & (g653) & (!g654) & (g655) & (g165) & (g166)) + ((g652) & (g653) & (g654) & (!g655) & (!g165) & (!g166)) + ((g652) & (g653) & (g654) & (!g655) & (!g165) & (g166)) + ((g652) & (g653) & (g654) & (!g655) & (g165) & (!g166)) + ((g652) & (g653) & (g654) & (g655) & (!g165) & (!g166)) + ((g652) & (g653) & (g654) & (g655) & (!g165) & (g166)) + ((g652) & (g653) & (g654) & (g655) & (g165) & (!g166)) + ((g652) & (g653) & (g654) & (g655) & (g165) & (g166)));
	assign g4361 = (((!sk[83]) & (!g2177) & (!g2454) & (g657)) + ((!sk[83]) & (!g2177) & (g2454) & (!g657)) + ((!sk[83]) & (!g2177) & (g2454) & (g657)) + ((!sk[83]) & (g2177) & (!g2454) & (g657)) + ((!sk[83]) & (g2177) & (g2454) & (!g657)) + ((!sk[83]) & (g2177) & (g2454) & (g657)) + ((sk[83]) & (!g2177) & (!g2454) & (g657)) + ((sk[83]) & (!g2177) & (g2454) & (g657)) + ((sk[83]) & (g2177) & (g2454) & (!g657)) + ((sk[83]) & (g2177) & (g2454) & (g657)));
	assign g4362 = (((!g2178) & (!g2454) & (!sk[84]) & (g658)) + ((!g2178) & (!g2454) & (sk[84]) & (g658)) + ((!g2178) & (g2454) & (!sk[84]) & (!g658)) + ((!g2178) & (g2454) & (!sk[84]) & (g658)) + ((!g2178) & (g2454) & (sk[84]) & (g658)) + ((g2178) & (!g2454) & (!sk[84]) & (g658)) + ((g2178) & (g2454) & (!sk[84]) & (!g658)) + ((g2178) & (g2454) & (!sk[84]) & (g658)) + ((g2178) & (g2454) & (sk[84]) & (!g658)) + ((g2178) & (g2454) & (sk[84]) & (g658)));
	assign g4363 = (((!g2179) & (!g2454) & (!sk[85]) & (g659)) + ((!g2179) & (!g2454) & (sk[85]) & (g659)) + ((!g2179) & (g2454) & (!sk[85]) & (!g659)) + ((!g2179) & (g2454) & (!sk[85]) & (g659)) + ((!g2179) & (g2454) & (sk[85]) & (g659)) + ((g2179) & (!g2454) & (!sk[85]) & (g659)) + ((g2179) & (g2454) & (!sk[85]) & (!g659)) + ((g2179) & (g2454) & (!sk[85]) & (g659)) + ((g2179) & (g2454) & (sk[85]) & (!g659)) + ((g2179) & (g2454) & (sk[85]) & (g659)));
	assign g660 = (((!g165) & (!g166) & (!g657) & (g658) & (!sk[86]) & (!g659)) + ((!g165) & (!g166) & (!g657) & (g658) & (!sk[86]) & (g659)) + ((!g165) & (!g166) & (g657) & (!g658) & (!sk[86]) & (!g659)) + ((!g165) & (!g166) & (g657) & (!g658) & (!sk[86]) & (g659)) + ((!g165) & (!g166) & (g657) & (g658) & (!sk[86]) & (!g659)) + ((!g165) & (!g166) & (g657) & (g658) & (!sk[86]) & (g659)) + ((!g165) & (g166) & (!g657) & (!g658) & (!sk[86]) & (!g659)) + ((!g165) & (g166) & (!g657) & (!g658) & (!sk[86]) & (g659)) + ((!g165) & (g166) & (!g657) & (!g658) & (sk[86]) & (g659)) + ((!g165) & (g166) & (!g657) & (g658) & (!sk[86]) & (!g659)) + ((!g165) & (g166) & (!g657) & (g658) & (!sk[86]) & (g659)) + ((!g165) & (g166) & (!g657) & (g658) & (sk[86]) & (g659)) + ((!g165) & (g166) & (g657) & (!g658) & (!sk[86]) & (!g659)) + ((!g165) & (g166) & (g657) & (!g658) & (!sk[86]) & (g659)) + ((!g165) & (g166) & (g657) & (!g658) & (sk[86]) & (g659)) + ((!g165) & (g166) & (g657) & (g658) & (!sk[86]) & (!g659)) + ((!g165) & (g166) & (g657) & (g658) & (!sk[86]) & (g659)) + ((!g165) & (g166) & (g657) & (g658) & (sk[86]) & (g659)) + ((g165) & (!g166) & (!g657) & (g658) & (!sk[86]) & (!g659)) + ((g165) & (!g166) & (!g657) & (g658) & (!sk[86]) & (g659)) + ((g165) & (!g166) & (g657) & (!g658) & (!sk[86]) & (!g659)) + ((g165) & (!g166) & (g657) & (!g658) & (!sk[86]) & (g659)) + ((g165) & (!g166) & (g657) & (!g658) & (sk[86]) & (!g659)) + ((g165) & (!g166) & (g657) & (!g658) & (sk[86]) & (g659)) + ((g165) & (!g166) & (g657) & (g658) & (!sk[86]) & (!g659)) + ((g165) & (!g166) & (g657) & (g658) & (!sk[86]) & (g659)) + ((g165) & (!g166) & (g657) & (g658) & (sk[86]) & (!g659)) + ((g165) & (!g166) & (g657) & (g658) & (sk[86]) & (g659)) + ((g165) & (g166) & (!g657) & (!g658) & (!sk[86]) & (!g659)) + ((g165) & (g166) & (!g657) & (!g658) & (!sk[86]) & (g659)) + ((g165) & (g166) & (!g657) & (g658) & (!sk[86]) & (!g659)) + ((g165) & (g166) & (!g657) & (g658) & (!sk[86]) & (g659)) + ((g165) & (g166) & (!g657) & (g658) & (sk[86]) & (!g659)) + ((g165) & (g166) & (!g657) & (g658) & (sk[86]) & (g659)) + ((g165) & (g166) & (g657) & (!g658) & (!sk[86]) & (!g659)) + ((g165) & (g166) & (g657) & (!g658) & (!sk[86]) & (g659)) + ((g165) & (g166) & (g657) & (g658) & (!sk[86]) & (!g659)) + ((g165) & (g166) & (g657) & (g658) & (!sk[86]) & (g659)) + ((g165) & (g166) & (g657) & (g658) & (sk[86]) & (!g659)) + ((g165) & (g166) & (g657) & (g658) & (sk[86]) & (g659)));
	assign g4364 = (((!g2162) & (!sk[87]) & (!g2454) & (g661)) + ((!g2162) & (!sk[87]) & (g2454) & (!g661)) + ((!g2162) & (!sk[87]) & (g2454) & (g661)) + ((!g2162) & (sk[87]) & (!g2454) & (g661)) + ((!g2162) & (sk[87]) & (g2454) & (g661)) + ((g2162) & (!sk[87]) & (!g2454) & (g661)) + ((g2162) & (!sk[87]) & (g2454) & (!g661)) + ((g2162) & (!sk[87]) & (g2454) & (g661)) + ((g2162) & (sk[87]) & (g2454) & (!g661)) + ((g2162) & (sk[87]) & (g2454) & (g661)));
	assign g4365 = (((!sk[88]) & (!g2164) & (!g2454) & (g662)) + ((!sk[88]) & (!g2164) & (g2454) & (!g662)) + ((!sk[88]) & (!g2164) & (g2454) & (g662)) + ((!sk[88]) & (g2164) & (!g2454) & (g662)) + ((!sk[88]) & (g2164) & (g2454) & (!g662)) + ((!sk[88]) & (g2164) & (g2454) & (g662)) + ((sk[88]) & (!g2164) & (!g2454) & (g662)) + ((sk[88]) & (!g2164) & (g2454) & (g662)) + ((sk[88]) & (g2164) & (g2454) & (!g662)) + ((sk[88]) & (g2164) & (g2454) & (g662)));
	assign g4366 = (((!sk[89]) & (!g2166) & (!g2454) & (g663)) + ((!sk[89]) & (!g2166) & (g2454) & (!g663)) + ((!sk[89]) & (!g2166) & (g2454) & (g663)) + ((!sk[89]) & (g2166) & (!g2454) & (g663)) + ((!sk[89]) & (g2166) & (g2454) & (!g663)) + ((!sk[89]) & (g2166) & (g2454) & (g663)) + ((sk[89]) & (!g2166) & (!g2454) & (g663)) + ((sk[89]) & (!g2166) & (g2454) & (g663)) + ((sk[89]) & (g2166) & (g2454) & (!g663)) + ((sk[89]) & (g2166) & (g2454) & (g663)));
	assign g4367 = (((!g2168) & (!g2454) & (!sk[90]) & (g664)) + ((!g2168) & (!g2454) & (sk[90]) & (g664)) + ((!g2168) & (g2454) & (!sk[90]) & (!g664)) + ((!g2168) & (g2454) & (!sk[90]) & (g664)) + ((!g2168) & (g2454) & (sk[90]) & (g664)) + ((g2168) & (!g2454) & (!sk[90]) & (g664)) + ((g2168) & (g2454) & (!sk[90]) & (!g664)) + ((g2168) & (g2454) & (!sk[90]) & (g664)) + ((g2168) & (g2454) & (sk[90]) & (!g664)) + ((g2168) & (g2454) & (sk[90]) & (g664)));
	assign g665 = (((!g661) & (!g662) & (!g663) & (g664) & (g165) & (g166)) + ((!g661) & (!g662) & (g663) & (!g664) & (!g165) & (g166)) + ((!g661) & (!g662) & (g663) & (g664) & (!g165) & (g166)) + ((!g661) & (!g662) & (g663) & (g664) & (g165) & (g166)) + ((!g661) & (g662) & (!g663) & (!g664) & (g165) & (!g166)) + ((!g661) & (g662) & (!g663) & (g664) & (g165) & (!g166)) + ((!g661) & (g662) & (!g663) & (g664) & (g165) & (g166)) + ((!g661) & (g662) & (g663) & (!g664) & (!g165) & (g166)) + ((!g661) & (g662) & (g663) & (!g664) & (g165) & (!g166)) + ((!g661) & (g662) & (g663) & (g664) & (!g165) & (g166)) + ((!g661) & (g662) & (g663) & (g664) & (g165) & (!g166)) + ((!g661) & (g662) & (g663) & (g664) & (g165) & (g166)) + ((g661) & (!g662) & (!g663) & (!g664) & (!g165) & (!g166)) + ((g661) & (!g662) & (!g663) & (g664) & (!g165) & (!g166)) + ((g661) & (!g662) & (!g663) & (g664) & (g165) & (g166)) + ((g661) & (!g662) & (g663) & (!g664) & (!g165) & (!g166)) + ((g661) & (!g662) & (g663) & (!g664) & (!g165) & (g166)) + ((g661) & (!g662) & (g663) & (g664) & (!g165) & (!g166)) + ((g661) & (!g662) & (g663) & (g664) & (!g165) & (g166)) + ((g661) & (!g662) & (g663) & (g664) & (g165) & (g166)) + ((g661) & (g662) & (!g663) & (!g664) & (!g165) & (!g166)) + ((g661) & (g662) & (!g663) & (!g664) & (g165) & (!g166)) + ((g661) & (g662) & (!g663) & (g664) & (!g165) & (!g166)) + ((g661) & (g662) & (!g663) & (g664) & (g165) & (!g166)) + ((g661) & (g662) & (!g663) & (g664) & (g165) & (g166)) + ((g661) & (g662) & (g663) & (!g664) & (!g165) & (!g166)) + ((g661) & (g662) & (g663) & (!g664) & (!g165) & (g166)) + ((g661) & (g662) & (g663) & (!g664) & (g165) & (!g166)) + ((g661) & (g662) & (g663) & (g664) & (!g165) & (!g166)) + ((g661) & (g662) & (g663) & (g664) & (!g165) & (g166)) + ((g661) & (g662) & (g663) & (g664) & (g165) & (!g166)) + ((g661) & (g662) & (g663) & (g664) & (g165) & (g166)));
	assign g4368 = (((!sk[92]) & (!g2169) & (!g2454) & (g666)) + ((!sk[92]) & (!g2169) & (g2454) & (!g666)) + ((!sk[92]) & (!g2169) & (g2454) & (g666)) + ((!sk[92]) & (g2169) & (!g2454) & (g666)) + ((!sk[92]) & (g2169) & (g2454) & (!g666)) + ((!sk[92]) & (g2169) & (g2454) & (g666)) + ((sk[92]) & (!g2169) & (!g2454) & (g666)) + ((sk[92]) & (!g2169) & (g2454) & (g666)) + ((sk[92]) & (g2169) & (g2454) & (!g666)) + ((sk[92]) & (g2169) & (g2454) & (g666)));
	assign g4369 = (((!sk[93]) & (!g2170) & (!g2454) & (g667)) + ((!sk[93]) & (!g2170) & (g2454) & (!g667)) + ((!sk[93]) & (!g2170) & (g2454) & (g667)) + ((!sk[93]) & (g2170) & (!g2454) & (g667)) + ((!sk[93]) & (g2170) & (g2454) & (!g667)) + ((!sk[93]) & (g2170) & (g2454) & (g667)) + ((sk[93]) & (!g2170) & (!g2454) & (g667)) + ((sk[93]) & (!g2170) & (g2454) & (g667)) + ((sk[93]) & (g2170) & (g2454) & (!g667)) + ((sk[93]) & (g2170) & (g2454) & (g667)));
	assign g4370 = (((!g2171) & (!g2454) & (!sk[94]) & (g668)) + ((!g2171) & (!g2454) & (sk[94]) & (g668)) + ((!g2171) & (g2454) & (!sk[94]) & (!g668)) + ((!g2171) & (g2454) & (!sk[94]) & (g668)) + ((!g2171) & (g2454) & (sk[94]) & (g668)) + ((g2171) & (!g2454) & (!sk[94]) & (g668)) + ((g2171) & (g2454) & (!sk[94]) & (!g668)) + ((g2171) & (g2454) & (!sk[94]) & (g668)) + ((g2171) & (g2454) & (sk[94]) & (!g668)) + ((g2171) & (g2454) & (sk[94]) & (g668)));
	assign g4371 = (((!sk[95]) & (!g2172) & (!g2454) & (g669)) + ((!sk[95]) & (!g2172) & (g2454) & (!g669)) + ((!sk[95]) & (!g2172) & (g2454) & (g669)) + ((!sk[95]) & (g2172) & (!g2454) & (g669)) + ((!sk[95]) & (g2172) & (g2454) & (!g669)) + ((!sk[95]) & (g2172) & (g2454) & (g669)) + ((sk[95]) & (!g2172) & (!g2454) & (g669)) + ((sk[95]) & (!g2172) & (g2454) & (g669)) + ((sk[95]) & (g2172) & (g2454) & (!g669)) + ((sk[95]) & (g2172) & (g2454) & (g669)));
	assign g670 = (((!g666) & (!g667) & (!g668) & (g669) & (g165) & (g166)) + ((!g666) & (!g667) & (g668) & (!g669) & (!g165) & (g166)) + ((!g666) & (!g667) & (g668) & (g669) & (!g165) & (g166)) + ((!g666) & (!g667) & (g668) & (g669) & (g165) & (g166)) + ((!g666) & (g667) & (!g668) & (!g669) & (g165) & (!g166)) + ((!g666) & (g667) & (!g668) & (g669) & (g165) & (!g166)) + ((!g666) & (g667) & (!g668) & (g669) & (g165) & (g166)) + ((!g666) & (g667) & (g668) & (!g669) & (!g165) & (g166)) + ((!g666) & (g667) & (g668) & (!g669) & (g165) & (!g166)) + ((!g666) & (g667) & (g668) & (g669) & (!g165) & (g166)) + ((!g666) & (g667) & (g668) & (g669) & (g165) & (!g166)) + ((!g666) & (g667) & (g668) & (g669) & (g165) & (g166)) + ((g666) & (!g667) & (!g668) & (!g669) & (!g165) & (!g166)) + ((g666) & (!g667) & (!g668) & (g669) & (!g165) & (!g166)) + ((g666) & (!g667) & (!g668) & (g669) & (g165) & (g166)) + ((g666) & (!g667) & (g668) & (!g669) & (!g165) & (!g166)) + ((g666) & (!g667) & (g668) & (!g669) & (!g165) & (g166)) + ((g666) & (!g667) & (g668) & (g669) & (!g165) & (!g166)) + ((g666) & (!g667) & (g668) & (g669) & (!g165) & (g166)) + ((g666) & (!g667) & (g668) & (g669) & (g165) & (g166)) + ((g666) & (g667) & (!g668) & (!g669) & (!g165) & (!g166)) + ((g666) & (g667) & (!g668) & (!g669) & (g165) & (!g166)) + ((g666) & (g667) & (!g668) & (g669) & (!g165) & (!g166)) + ((g666) & (g667) & (!g668) & (g669) & (g165) & (!g166)) + ((g666) & (g667) & (!g668) & (g669) & (g165) & (g166)) + ((g666) & (g667) & (g668) & (!g669) & (!g165) & (!g166)) + ((g666) & (g667) & (g668) & (!g669) & (!g165) & (g166)) + ((g666) & (g667) & (g668) & (!g669) & (g165) & (!g166)) + ((g666) & (g667) & (g668) & (g669) & (!g165) & (!g166)) + ((g666) & (g667) & (g668) & (g669) & (!g165) & (g166)) + ((g666) & (g667) & (g668) & (g669) & (g165) & (!g166)) + ((g666) & (g667) & (g668) & (g669) & (g165) & (g166)));
	assign g671 = (((!g147) & (!g148) & (!g656) & (g660) & (!g665) & (!g670)) + ((!g147) & (!g148) & (!g656) & (g660) & (!g665) & (g670)) + ((!g147) & (!g148) & (!g656) & (g660) & (g665) & (!g670)) + ((!g147) & (!g148) & (!g656) & (g660) & (g665) & (g670)) + ((!g147) & (!g148) & (g656) & (g660) & (!g665) & (!g670)) + ((!g147) & (!g148) & (g656) & (g660) & (!g665) & (g670)) + ((!g147) & (!g148) & (g656) & (g660) & (g665) & (!g670)) + ((!g147) & (!g148) & (g656) & (g660) & (g665) & (g670)) + ((!g147) & (g148) & (!g656) & (!g660) & (!g665) & (g670)) + ((!g147) & (g148) & (!g656) & (!g660) & (g665) & (g670)) + ((!g147) & (g148) & (!g656) & (g660) & (!g665) & (g670)) + ((!g147) & (g148) & (!g656) & (g660) & (g665) & (g670)) + ((!g147) & (g148) & (g656) & (!g660) & (!g665) & (g670)) + ((!g147) & (g148) & (g656) & (!g660) & (g665) & (g670)) + ((!g147) & (g148) & (g656) & (g660) & (!g665) & (g670)) + ((!g147) & (g148) & (g656) & (g660) & (g665) & (g670)) + ((g147) & (!g148) & (g656) & (!g660) & (!g665) & (!g670)) + ((g147) & (!g148) & (g656) & (!g660) & (!g665) & (g670)) + ((g147) & (!g148) & (g656) & (!g660) & (g665) & (!g670)) + ((g147) & (!g148) & (g656) & (!g660) & (g665) & (g670)) + ((g147) & (!g148) & (g656) & (g660) & (!g665) & (!g670)) + ((g147) & (!g148) & (g656) & (g660) & (!g665) & (g670)) + ((g147) & (!g148) & (g656) & (g660) & (g665) & (!g670)) + ((g147) & (!g148) & (g656) & (g660) & (g665) & (g670)) + ((g147) & (g148) & (!g656) & (!g660) & (g665) & (!g670)) + ((g147) & (g148) & (!g656) & (!g660) & (g665) & (g670)) + ((g147) & (g148) & (!g656) & (g660) & (g665) & (!g670)) + ((g147) & (g148) & (!g656) & (g660) & (g665) & (g670)) + ((g147) & (g148) & (g656) & (!g660) & (g665) & (!g670)) + ((g147) & (g148) & (g656) & (!g660) & (g665) & (g670)) + ((g147) & (g148) & (g656) & (g660) & (g665) & (!g670)) + ((g147) & (g148) & (g656) & (g660) & (g665) & (g670)));
	assign g672 = (((!g142) & (!g651) & (!sk[98]) & (g671)) + ((!g142) & (!g651) & (sk[98]) & (g671)) + ((!g142) & (g651) & (!sk[98]) & (!g671)) + ((!g142) & (g651) & (!sk[98]) & (g671)) + ((!g142) & (g651) & (sk[98]) & (g671)) + ((g142) & (!g651) & (!sk[98]) & (g671)) + ((g142) & (g651) & (!sk[98]) & (!g671)) + ((g142) & (g651) & (!sk[98]) & (g671)) + ((g142) & (g651) & (sk[98]) & (!g671)) + ((g142) & (g651) & (sk[98]) & (g671)));
	assign g673 = (((!g586) & (sk[99]) & (g629)) + ((g586) & (!sk[99]) & (!g629)) + ((g586) & (!sk[99]) & (g629)) + ((g586) & (sk[99]) & (!g629)));
	assign g674 = (((!g91) & (!g92) & (g497) & (g539) & (g584) & (g673)) + ((!g91) & (g92) & (!g497) & (g539) & (g584) & (g673)) + ((!g91) & (g92) & (g497) & (!g539) & (g584) & (g673)) + ((!g91) & (g92) & (g497) & (g539) & (g584) & (g673)) + ((g91) & (!g92) & (!g497) & (!g539) & (g584) & (g673)) + ((g91) & (!g92) & (!g497) & (g539) & (g584) & (g673)) + ((g91) & (!g92) & (g497) & (!g539) & (g584) & (g673)) + ((g91) & (!g92) & (g497) & (g539) & (!g584) & (g673)) + ((g91) & (!g92) & (g497) & (g539) & (g584) & (g673)) + ((g91) & (g92) & (!g497) & (!g539) & (g584) & (g673)) + ((g91) & (g92) & (!g497) & (g539) & (!g584) & (g673)) + ((g91) & (g92) & (!g497) & (g539) & (g584) & (g673)) + ((g91) & (g92) & (g497) & (!g539) & (!g584) & (g673)) + ((g91) & (g92) & (g497) & (!g539) & (g584) & (g673)) + ((g91) & (g92) & (g497) & (g539) & (!g584) & (g673)) + ((g91) & (g92) & (g497) & (g539) & (g584) & (g673)));
	assign g675 = (((g586) & (!sk[101]) & (!g629)) + ((g586) & (!sk[101]) & (g629)) + ((g586) & (sk[101]) & (g629)));
	assign g676 = (((!sk[102]) & (g674) & (!g675)) + ((!sk[102]) & (g674) & (g675)) + ((sk[102]) & (!g674) & (!g675)));
	assign g4372 = (((!g2064) & (!sk[103]) & (!dmem_dat_ix11x) & (g677)) + ((!g2064) & (!sk[103]) & (dmem_dat_ix11x) & (!g677)) + ((!g2064) & (!sk[103]) & (dmem_dat_ix11x) & (g677)) + ((!g2064) & (sk[103]) & (!dmem_dat_ix11x) & (g677)) + ((!g2064) & (sk[103]) & (dmem_dat_ix11x) & (g677)) + ((g2064) & (!sk[103]) & (!dmem_dat_ix11x) & (g677)) + ((g2064) & (!sk[103]) & (dmem_dat_ix11x) & (!g677)) + ((g2064) & (!sk[103]) & (dmem_dat_ix11x) & (g677)) + ((g2064) & (sk[103]) & (dmem_dat_ix11x) & (!g677)) + ((g2064) & (sk[103]) & (dmem_dat_ix11x) & (g677)));
	assign g4373 = (((!g2064) & (!dmem_dat_ix21x) & (!sk[104]) & (g678)) + ((!g2064) & (!dmem_dat_ix21x) & (sk[104]) & (g678)) + ((!g2064) & (dmem_dat_ix21x) & (!sk[104]) & (!g678)) + ((!g2064) & (dmem_dat_ix21x) & (!sk[104]) & (g678)) + ((!g2064) & (dmem_dat_ix21x) & (sk[104]) & (g678)) + ((g2064) & (!dmem_dat_ix21x) & (!sk[104]) & (g678)) + ((g2064) & (dmem_dat_ix21x) & (!sk[104]) & (!g678)) + ((g2064) & (dmem_dat_ix21x) & (!sk[104]) & (g678)) + ((g2064) & (dmem_dat_ix21x) & (sk[104]) & (!g678)) + ((g2064) & (dmem_dat_ix21x) & (sk[104]) & (g678)));
	assign g679 = (((!sk[105]) & (g132) & (!g134)) + ((!sk[105]) & (g132) & (g134)) + ((sk[105]) & (!g132) & (!g134)));
	assign g680 = (((!g677) & (!sk[106]) & (!g678) & (g679)) + ((!g677) & (!sk[106]) & (g678) & (!g679)) + ((!g677) & (!sk[106]) & (g678) & (g679)) + ((!g677) & (sk[106]) & (!g678) & (!g679)) + ((!g677) & (sk[106]) & (!g678) & (g679)) + ((!g677) & (sk[106]) & (g678) & (g679)) + ((g677) & (!sk[106]) & (!g678) & (g679)) + ((g677) & (!sk[106]) & (g678) & (!g679)) + ((g677) & (!sk[106]) & (g678) & (g679)) + ((g677) & (sk[106]) & (!g678) & (!g679)));
	assign g681 = (((!g126) & (!sk[107]) & (!g630) & (!g672) & (g676) & (!g680)) + ((!g126) & (!sk[107]) & (!g630) & (!g672) & (g676) & (g680)) + ((!g126) & (!sk[107]) & (!g630) & (g672) & (!g676) & (!g680)) + ((!g126) & (!sk[107]) & (!g630) & (g672) & (!g676) & (g680)) + ((!g126) & (!sk[107]) & (!g630) & (g672) & (g676) & (!g680)) + ((!g126) & (!sk[107]) & (!g630) & (g672) & (g676) & (g680)) + ((!g126) & (!sk[107]) & (g630) & (!g672) & (!g676) & (!g680)) + ((!g126) & (!sk[107]) & (g630) & (!g672) & (!g676) & (g680)) + ((!g126) & (!sk[107]) & (g630) & (!g672) & (g676) & (!g680)) + ((!g126) & (!sk[107]) & (g630) & (!g672) & (g676) & (g680)) + ((!g126) & (!sk[107]) & (g630) & (g672) & (!g676) & (!g680)) + ((!g126) & (!sk[107]) & (g630) & (g672) & (!g676) & (g680)) + ((!g126) & (!sk[107]) & (g630) & (g672) & (g676) & (!g680)) + ((!g126) & (!sk[107]) & (g630) & (g672) & (g676) & (g680)) + ((!g126) & (sk[107]) & (g630) & (!g672) & (!g676) & (!g680)) + ((!g126) & (sk[107]) & (g630) & (!g672) & (!g676) & (g680)) + ((!g126) & (sk[107]) & (g630) & (!g672) & (g676) & (!g680)) + ((!g126) & (sk[107]) & (g630) & (!g672) & (g676) & (g680)) + ((!g126) & (sk[107]) & (g630) & (g672) & (!g676) & (!g680)) + ((!g126) & (sk[107]) & (g630) & (g672) & (!g676) & (g680)) + ((!g126) & (sk[107]) & (g630) & (g672) & (g676) & (!g680)) + ((!g126) & (sk[107]) & (g630) & (g672) & (g676) & (g680)) + ((g126) & (!sk[107]) & (!g630) & (!g672) & (g676) & (!g680)) + ((g126) & (!sk[107]) & (!g630) & (!g672) & (g676) & (g680)) + ((g126) & (!sk[107]) & (!g630) & (g672) & (!g676) & (!g680)) + ((g126) & (!sk[107]) & (!g630) & (g672) & (!g676) & (g680)) + ((g126) & (!sk[107]) & (!g630) & (g672) & (g676) & (!g680)) + ((g126) & (!sk[107]) & (!g630) & (g672) & (g676) & (g680)) + ((g126) & (!sk[107]) & (g630) & (!g672) & (!g676) & (!g680)) + ((g126) & (!sk[107]) & (g630) & (!g672) & (!g676) & (g680)) + ((g126) & (!sk[107]) & (g630) & (!g672) & (g676) & (!g680)) + ((g126) & (!sk[107]) & (g630) & (!g672) & (g676) & (g680)) + ((g126) & (!sk[107]) & (g630) & (g672) & (!g676) & (!g680)) + ((g126) & (!sk[107]) & (g630) & (g672) & (!g676) & (g680)) + ((g126) & (!sk[107]) & (g630) & (g672) & (g676) & (!g680)) + ((g126) & (!sk[107]) & (g630) & (g672) & (g676) & (g680)) + ((g126) & (sk[107]) & (!g630) & (!g672) & (!g676) & (g680)) + ((g126) & (sk[107]) & (!g630) & (!g672) & (g676) & (!g680)) + ((g126) & (sk[107]) & (!g630) & (g672) & (!g676) & (!g680)) + ((g126) & (sk[107]) & (!g630) & (g672) & (g676) & (g680)) + ((g126) & (sk[107]) & (g630) & (!g672) & (!g676) & (g680)) + ((g126) & (sk[107]) & (g630) & (!g672) & (g676) & (!g680)) + ((g126) & (sk[107]) & (g630) & (g672) & (!g676) & (!g680)) + ((g126) & (sk[107]) & (g630) & (g672) & (g676) & (g680)));
	assign g4374 = (((!g2140) & (!sk[108]) & (!g2473) & (g682)) + ((!g2140) & (!sk[108]) & (g2473) & (!g682)) + ((!g2140) & (!sk[108]) & (g2473) & (g682)) + ((!g2140) & (sk[108]) & (!g2473) & (g682)) + ((!g2140) & (sk[108]) & (g2473) & (g682)) + ((g2140) & (!sk[108]) & (!g2473) & (g682)) + ((g2140) & (!sk[108]) & (g2473) & (!g682)) + ((g2140) & (!sk[108]) & (g2473) & (g682)) + ((g2140) & (sk[108]) & (g2473) & (!g682)) + ((g2140) & (sk[108]) & (g2473) & (g682)));
	assign g4375 = (((!g2142) & (!g2473) & (!sk[109]) & (g683)) + ((!g2142) & (!g2473) & (sk[109]) & (g683)) + ((!g2142) & (g2473) & (!sk[109]) & (!g683)) + ((!g2142) & (g2473) & (!sk[109]) & (g683)) + ((!g2142) & (g2473) & (sk[109]) & (g683)) + ((g2142) & (!g2473) & (!sk[109]) & (g683)) + ((g2142) & (g2473) & (!sk[109]) & (!g683)) + ((g2142) & (g2473) & (!sk[109]) & (g683)) + ((g2142) & (g2473) & (sk[109]) & (!g683)) + ((g2142) & (g2473) & (sk[109]) & (g683)));
	assign g4376 = (((!g2144) & (!g2473) & (!sk[110]) & (g684)) + ((!g2144) & (!g2473) & (sk[110]) & (g684)) + ((!g2144) & (g2473) & (!sk[110]) & (!g684)) + ((!g2144) & (g2473) & (!sk[110]) & (g684)) + ((!g2144) & (g2473) & (sk[110]) & (g684)) + ((g2144) & (!g2473) & (!sk[110]) & (g684)) + ((g2144) & (g2473) & (!sk[110]) & (!g684)) + ((g2144) & (g2473) & (!sk[110]) & (g684)) + ((g2144) & (g2473) & (sk[110]) & (!g684)) + ((g2144) & (g2473) & (sk[110]) & (g684)));
	assign g4377 = (((!g2145) & (!g2473) & (!sk[111]) & (g685)) + ((!g2145) & (!g2473) & (sk[111]) & (g685)) + ((!g2145) & (g2473) & (!sk[111]) & (!g685)) + ((!g2145) & (g2473) & (!sk[111]) & (g685)) + ((!g2145) & (g2473) & (sk[111]) & (g685)) + ((g2145) & (!g2473) & (!sk[111]) & (g685)) + ((g2145) & (g2473) & (!sk[111]) & (!g685)) + ((g2145) & (g2473) & (!sk[111]) & (g685)) + ((g2145) & (g2473) & (sk[111]) & (!g685)) + ((g2145) & (g2473) & (sk[111]) & (g685)));
	assign g686 = (((!g682) & (!g683) & (!g684) & (g685) & (g147) & (g148)) + ((!g682) & (!g683) & (g684) & (!g685) & (!g147) & (g148)) + ((!g682) & (!g683) & (g684) & (g685) & (!g147) & (g148)) + ((!g682) & (!g683) & (g684) & (g685) & (g147) & (g148)) + ((!g682) & (g683) & (!g684) & (!g685) & (g147) & (!g148)) + ((!g682) & (g683) & (!g684) & (g685) & (g147) & (!g148)) + ((!g682) & (g683) & (!g684) & (g685) & (g147) & (g148)) + ((!g682) & (g683) & (g684) & (!g685) & (!g147) & (g148)) + ((!g682) & (g683) & (g684) & (!g685) & (g147) & (!g148)) + ((!g682) & (g683) & (g684) & (g685) & (!g147) & (g148)) + ((!g682) & (g683) & (g684) & (g685) & (g147) & (!g148)) + ((!g682) & (g683) & (g684) & (g685) & (g147) & (g148)) + ((g682) & (!g683) & (!g684) & (!g685) & (!g147) & (!g148)) + ((g682) & (!g683) & (!g684) & (g685) & (!g147) & (!g148)) + ((g682) & (!g683) & (!g684) & (g685) & (g147) & (g148)) + ((g682) & (!g683) & (g684) & (!g685) & (!g147) & (!g148)) + ((g682) & (!g683) & (g684) & (!g685) & (!g147) & (g148)) + ((g682) & (!g683) & (g684) & (g685) & (!g147) & (!g148)) + ((g682) & (!g683) & (g684) & (g685) & (!g147) & (g148)) + ((g682) & (!g683) & (g684) & (g685) & (g147) & (g148)) + ((g682) & (g683) & (!g684) & (!g685) & (!g147) & (!g148)) + ((g682) & (g683) & (!g684) & (!g685) & (g147) & (!g148)) + ((g682) & (g683) & (!g684) & (g685) & (!g147) & (!g148)) + ((g682) & (g683) & (!g684) & (g685) & (g147) & (!g148)) + ((g682) & (g683) & (!g684) & (g685) & (g147) & (g148)) + ((g682) & (g683) & (g684) & (!g685) & (!g147) & (!g148)) + ((g682) & (g683) & (g684) & (!g685) & (!g147) & (g148)) + ((g682) & (g683) & (g684) & (!g685) & (g147) & (!g148)) + ((g682) & (g683) & (g684) & (g685) & (!g147) & (!g148)) + ((g682) & (g683) & (g684) & (g685) & (!g147) & (g148)) + ((g682) & (g683) & (g684) & (g685) & (g147) & (!g148)) + ((g682) & (g683) & (g684) & (g685) & (g147) & (g148)));
	assign g4378 = (((!g2146) & (!sk[113]) & (!g2473) & (g687)) + ((!g2146) & (!sk[113]) & (g2473) & (!g687)) + ((!g2146) & (!sk[113]) & (g2473) & (g687)) + ((!g2146) & (sk[113]) & (!g2473) & (g687)) + ((!g2146) & (sk[113]) & (g2473) & (g687)) + ((g2146) & (!sk[113]) & (!g2473) & (g687)) + ((g2146) & (!sk[113]) & (g2473) & (!g687)) + ((g2146) & (!sk[113]) & (g2473) & (g687)) + ((g2146) & (sk[113]) & (g2473) & (!g687)) + ((g2146) & (sk[113]) & (g2473) & (g687)));
	assign g4379 = (((!sk[114]) & (!g2148) & (!g2473) & (g688)) + ((!sk[114]) & (!g2148) & (g2473) & (!g688)) + ((!sk[114]) & (!g2148) & (g2473) & (g688)) + ((!sk[114]) & (g2148) & (!g2473) & (g688)) + ((!sk[114]) & (g2148) & (g2473) & (!g688)) + ((!sk[114]) & (g2148) & (g2473) & (g688)) + ((sk[114]) & (!g2148) & (!g2473) & (g688)) + ((sk[114]) & (!g2148) & (g2473) & (g688)) + ((sk[114]) & (g2148) & (g2473) & (!g688)) + ((sk[114]) & (g2148) & (g2473) & (g688)));
	assign g4380 = (((!sk[115]) & (!g2150) & (!g2473) & (g689)) + ((!sk[115]) & (!g2150) & (g2473) & (!g689)) + ((!sk[115]) & (!g2150) & (g2473) & (g689)) + ((!sk[115]) & (g2150) & (!g2473) & (g689)) + ((!sk[115]) & (g2150) & (g2473) & (!g689)) + ((!sk[115]) & (g2150) & (g2473) & (g689)) + ((sk[115]) & (!g2150) & (!g2473) & (g689)) + ((sk[115]) & (!g2150) & (g2473) & (g689)) + ((sk[115]) & (g2150) & (g2473) & (!g689)) + ((sk[115]) & (g2150) & (g2473) & (g689)));
	assign g4381 = (((!g2151) & (!g2473) & (!sk[116]) & (g690)) + ((!g2151) & (!g2473) & (sk[116]) & (g690)) + ((!g2151) & (g2473) & (!sk[116]) & (!g690)) + ((!g2151) & (g2473) & (!sk[116]) & (g690)) + ((!g2151) & (g2473) & (sk[116]) & (g690)) + ((g2151) & (!g2473) & (!sk[116]) & (g690)) + ((g2151) & (g2473) & (!sk[116]) & (!g690)) + ((g2151) & (g2473) & (!sk[116]) & (g690)) + ((g2151) & (g2473) & (sk[116]) & (!g690)) + ((g2151) & (g2473) & (sk[116]) & (g690)));
	assign g691 = (((!g687) & (!g688) & (!g689) & (g690) & (g147) & (g148)) + ((!g687) & (!g688) & (g689) & (!g690) & (!g147) & (g148)) + ((!g687) & (!g688) & (g689) & (g690) & (!g147) & (g148)) + ((!g687) & (!g688) & (g689) & (g690) & (g147) & (g148)) + ((!g687) & (g688) & (!g689) & (!g690) & (g147) & (!g148)) + ((!g687) & (g688) & (!g689) & (g690) & (g147) & (!g148)) + ((!g687) & (g688) & (!g689) & (g690) & (g147) & (g148)) + ((!g687) & (g688) & (g689) & (!g690) & (!g147) & (g148)) + ((!g687) & (g688) & (g689) & (!g690) & (g147) & (!g148)) + ((!g687) & (g688) & (g689) & (g690) & (!g147) & (g148)) + ((!g687) & (g688) & (g689) & (g690) & (g147) & (!g148)) + ((!g687) & (g688) & (g689) & (g690) & (g147) & (g148)) + ((g687) & (!g688) & (!g689) & (!g690) & (!g147) & (!g148)) + ((g687) & (!g688) & (!g689) & (g690) & (!g147) & (!g148)) + ((g687) & (!g688) & (!g689) & (g690) & (g147) & (g148)) + ((g687) & (!g688) & (g689) & (!g690) & (!g147) & (!g148)) + ((g687) & (!g688) & (g689) & (!g690) & (!g147) & (g148)) + ((g687) & (!g688) & (g689) & (g690) & (!g147) & (!g148)) + ((g687) & (!g688) & (g689) & (g690) & (!g147) & (g148)) + ((g687) & (!g688) & (g689) & (g690) & (g147) & (g148)) + ((g687) & (g688) & (!g689) & (!g690) & (!g147) & (!g148)) + ((g687) & (g688) & (!g689) & (!g690) & (g147) & (!g148)) + ((g687) & (g688) & (!g689) & (g690) & (!g147) & (!g148)) + ((g687) & (g688) & (!g689) & (g690) & (g147) & (!g148)) + ((g687) & (g688) & (!g689) & (g690) & (g147) & (g148)) + ((g687) & (g688) & (g689) & (!g690) & (!g147) & (!g148)) + ((g687) & (g688) & (g689) & (!g690) & (!g147) & (g148)) + ((g687) & (g688) & (g689) & (!g690) & (g147) & (!g148)) + ((g687) & (g688) & (g689) & (g690) & (!g147) & (!g148)) + ((g687) & (g688) & (g689) & (g690) & (!g147) & (g148)) + ((g687) & (g688) & (g689) & (g690) & (g147) & (!g148)) + ((g687) & (g688) & (g689) & (g690) & (g147) & (g148)));
	assign g4382 = (((!g2152) & (!g2473) & (!sk[118]) & (g692)) + ((!g2152) & (!g2473) & (sk[118]) & (g692)) + ((!g2152) & (g2473) & (!sk[118]) & (!g692)) + ((!g2152) & (g2473) & (!sk[118]) & (g692)) + ((!g2152) & (g2473) & (sk[118]) & (g692)) + ((g2152) & (!g2473) & (!sk[118]) & (g692)) + ((g2152) & (g2473) & (!sk[118]) & (!g692)) + ((g2152) & (g2473) & (!sk[118]) & (g692)) + ((g2152) & (g2473) & (sk[118]) & (!g692)) + ((g2152) & (g2473) & (sk[118]) & (g692)));
	assign g4383 = (((!g2153) & (!g2473) & (!sk[119]) & (g693)) + ((!g2153) & (!g2473) & (sk[119]) & (g693)) + ((!g2153) & (g2473) & (!sk[119]) & (!g693)) + ((!g2153) & (g2473) & (!sk[119]) & (g693)) + ((!g2153) & (g2473) & (sk[119]) & (g693)) + ((g2153) & (!g2473) & (!sk[119]) & (g693)) + ((g2153) & (g2473) & (!sk[119]) & (!g693)) + ((g2153) & (g2473) & (!sk[119]) & (g693)) + ((g2153) & (g2473) & (sk[119]) & (!g693)) + ((g2153) & (g2473) & (sk[119]) & (g693)));
	assign g4384 = (((!sk[120]) & (!g2155) & (!g2473) & (g694)) + ((!sk[120]) & (!g2155) & (g2473) & (!g694)) + ((!sk[120]) & (!g2155) & (g2473) & (g694)) + ((!sk[120]) & (g2155) & (!g2473) & (g694)) + ((!sk[120]) & (g2155) & (g2473) & (!g694)) + ((!sk[120]) & (g2155) & (g2473) & (g694)) + ((sk[120]) & (!g2155) & (!g2473) & (g694)) + ((sk[120]) & (!g2155) & (g2473) & (g694)) + ((sk[120]) & (g2155) & (g2473) & (!g694)) + ((sk[120]) & (g2155) & (g2473) & (g694)));
	assign g4385 = (((!g2157) & (!g2473) & (!sk[121]) & (g695)) + ((!g2157) & (!g2473) & (sk[121]) & (g695)) + ((!g2157) & (g2473) & (!sk[121]) & (!g695)) + ((!g2157) & (g2473) & (!sk[121]) & (g695)) + ((!g2157) & (g2473) & (sk[121]) & (g695)) + ((g2157) & (!g2473) & (!sk[121]) & (g695)) + ((g2157) & (g2473) & (!sk[121]) & (!g695)) + ((g2157) & (g2473) & (!sk[121]) & (g695)) + ((g2157) & (g2473) & (sk[121]) & (!g695)) + ((g2157) & (g2473) & (sk[121]) & (g695)));
	assign g696 = (((!g692) & (!g693) & (!g694) & (g695) & (g147) & (g148)) + ((!g692) & (!g693) & (g694) & (!g695) & (!g147) & (g148)) + ((!g692) & (!g693) & (g694) & (g695) & (!g147) & (g148)) + ((!g692) & (!g693) & (g694) & (g695) & (g147) & (g148)) + ((!g692) & (g693) & (!g694) & (!g695) & (g147) & (!g148)) + ((!g692) & (g693) & (!g694) & (g695) & (g147) & (!g148)) + ((!g692) & (g693) & (!g694) & (g695) & (g147) & (g148)) + ((!g692) & (g693) & (g694) & (!g695) & (!g147) & (g148)) + ((!g692) & (g693) & (g694) & (!g695) & (g147) & (!g148)) + ((!g692) & (g693) & (g694) & (g695) & (!g147) & (g148)) + ((!g692) & (g693) & (g694) & (g695) & (g147) & (!g148)) + ((!g692) & (g693) & (g694) & (g695) & (g147) & (g148)) + ((g692) & (!g693) & (!g694) & (!g695) & (!g147) & (!g148)) + ((g692) & (!g693) & (!g694) & (g695) & (!g147) & (!g148)) + ((g692) & (!g693) & (!g694) & (g695) & (g147) & (g148)) + ((g692) & (!g693) & (g694) & (!g695) & (!g147) & (!g148)) + ((g692) & (!g693) & (g694) & (!g695) & (!g147) & (g148)) + ((g692) & (!g693) & (g694) & (g695) & (!g147) & (!g148)) + ((g692) & (!g693) & (g694) & (g695) & (!g147) & (g148)) + ((g692) & (!g693) & (g694) & (g695) & (g147) & (g148)) + ((g692) & (g693) & (!g694) & (!g695) & (!g147) & (!g148)) + ((g692) & (g693) & (!g694) & (!g695) & (g147) & (!g148)) + ((g692) & (g693) & (!g694) & (g695) & (!g147) & (!g148)) + ((g692) & (g693) & (!g694) & (g695) & (g147) & (!g148)) + ((g692) & (g693) & (!g694) & (g695) & (g147) & (g148)) + ((g692) & (g693) & (g694) & (!g695) & (!g147) & (!g148)) + ((g692) & (g693) & (g694) & (!g695) & (!g147) & (g148)) + ((g692) & (g693) & (g694) & (!g695) & (g147) & (!g148)) + ((g692) & (g693) & (g694) & (g695) & (!g147) & (!g148)) + ((g692) & (g693) & (g694) & (g695) & (!g147) & (g148)) + ((g692) & (g693) & (g694) & (g695) & (g147) & (!g148)) + ((g692) & (g693) & (g694) & (g695) & (g147) & (g148)));
	assign g4386 = (((!sk[123]) & (!g2158) & (!g2473) & (g697)) + ((!sk[123]) & (!g2158) & (g2473) & (!g697)) + ((!sk[123]) & (!g2158) & (g2473) & (g697)) + ((!sk[123]) & (g2158) & (!g2473) & (g697)) + ((!sk[123]) & (g2158) & (g2473) & (!g697)) + ((!sk[123]) & (g2158) & (g2473) & (g697)) + ((sk[123]) & (!g2158) & (!g2473) & (g697)) + ((sk[123]) & (!g2158) & (g2473) & (g697)) + ((sk[123]) & (g2158) & (g2473) & (!g697)) + ((sk[123]) & (g2158) & (g2473) & (g697)));
	assign g4387 = (((!sk[124]) & (!g2159) & (!g2473) & (g698)) + ((!sk[124]) & (!g2159) & (g2473) & (!g698)) + ((!sk[124]) & (!g2159) & (g2473) & (g698)) + ((!sk[124]) & (g2159) & (!g2473) & (g698)) + ((!sk[124]) & (g2159) & (g2473) & (!g698)) + ((!sk[124]) & (g2159) & (g2473) & (g698)) + ((sk[124]) & (!g2159) & (!g2473) & (g698)) + ((sk[124]) & (!g2159) & (g2473) & (g698)) + ((sk[124]) & (g2159) & (g2473) & (!g698)) + ((sk[124]) & (g2159) & (g2473) & (g698)));
	assign g4388 = (((!g2160) & (!g2473) & (!sk[125]) & (g699)) + ((!g2160) & (!g2473) & (sk[125]) & (g699)) + ((!g2160) & (g2473) & (!sk[125]) & (!g699)) + ((!g2160) & (g2473) & (!sk[125]) & (g699)) + ((!g2160) & (g2473) & (sk[125]) & (g699)) + ((g2160) & (!g2473) & (!sk[125]) & (g699)) + ((g2160) & (g2473) & (!sk[125]) & (!g699)) + ((g2160) & (g2473) & (!sk[125]) & (g699)) + ((g2160) & (g2473) & (sk[125]) & (!g699)) + ((g2160) & (g2473) & (sk[125]) & (g699)));
	assign g4389 = (((!g2161) & (!g2473) & (!sk[126]) & (g700)) + ((!g2161) & (!g2473) & (sk[126]) & (g700)) + ((!g2161) & (g2473) & (!sk[126]) & (!g700)) + ((!g2161) & (g2473) & (!sk[126]) & (g700)) + ((!g2161) & (g2473) & (sk[126]) & (g700)) + ((g2161) & (!g2473) & (!sk[126]) & (g700)) + ((g2161) & (g2473) & (!sk[126]) & (!g700)) + ((g2161) & (g2473) & (!sk[126]) & (g700)) + ((g2161) & (g2473) & (sk[126]) & (!g700)) + ((g2161) & (g2473) & (sk[126]) & (g700)));
	assign g701 = (((!g697) & (!g698) & (!g699) & (g700) & (g147) & (g148)) + ((!g697) & (!g698) & (g699) & (!g700) & (!g147) & (g148)) + ((!g697) & (!g698) & (g699) & (g700) & (!g147) & (g148)) + ((!g697) & (!g698) & (g699) & (g700) & (g147) & (g148)) + ((!g697) & (g698) & (!g699) & (!g700) & (g147) & (!g148)) + ((!g697) & (g698) & (!g699) & (g700) & (g147) & (!g148)) + ((!g697) & (g698) & (!g699) & (g700) & (g147) & (g148)) + ((!g697) & (g698) & (g699) & (!g700) & (!g147) & (g148)) + ((!g697) & (g698) & (g699) & (!g700) & (g147) & (!g148)) + ((!g697) & (g698) & (g699) & (g700) & (!g147) & (g148)) + ((!g697) & (g698) & (g699) & (g700) & (g147) & (!g148)) + ((!g697) & (g698) & (g699) & (g700) & (g147) & (g148)) + ((g697) & (!g698) & (!g699) & (!g700) & (!g147) & (!g148)) + ((g697) & (!g698) & (!g699) & (g700) & (!g147) & (!g148)) + ((g697) & (!g698) & (!g699) & (g700) & (g147) & (g148)) + ((g697) & (!g698) & (g699) & (!g700) & (!g147) & (!g148)) + ((g697) & (!g698) & (g699) & (!g700) & (!g147) & (g148)) + ((g697) & (!g698) & (g699) & (g700) & (!g147) & (!g148)) + ((g697) & (!g698) & (g699) & (g700) & (!g147) & (g148)) + ((g697) & (!g698) & (g699) & (g700) & (g147) & (g148)) + ((g697) & (g698) & (!g699) & (!g700) & (!g147) & (!g148)) + ((g697) & (g698) & (!g699) & (!g700) & (g147) & (!g148)) + ((g697) & (g698) & (!g699) & (g700) & (!g147) & (!g148)) + ((g697) & (g698) & (!g699) & (g700) & (g147) & (!g148)) + ((g697) & (g698) & (!g699) & (g700) & (g147) & (g148)) + ((g697) & (g698) & (g699) & (!g700) & (!g147) & (!g148)) + ((g697) & (g698) & (g699) & (!g700) & (!g147) & (g148)) + ((g697) & (g698) & (g699) & (!g700) & (g147) & (!g148)) + ((g697) & (g698) & (g699) & (g700) & (!g147) & (!g148)) + ((g697) & (g698) & (g699) & (g700) & (!g147) & (g148)) + ((g697) & (g698) & (g699) & (g700) & (g147) & (!g148)) + ((g697) & (g698) & (g699) & (g700) & (g147) & (g148)));
	assign g702 = (((!g686) & (!g691) & (!g696) & (g701) & (g165) & (g166)) + ((!g686) & (!g691) & (g696) & (!g701) & (!g165) & (g166)) + ((!g686) & (!g691) & (g696) & (g701) & (!g165) & (g166)) + ((!g686) & (!g691) & (g696) & (g701) & (g165) & (g166)) + ((!g686) & (g691) & (!g696) & (!g701) & (g165) & (!g166)) + ((!g686) & (g691) & (!g696) & (g701) & (g165) & (!g166)) + ((!g686) & (g691) & (!g696) & (g701) & (g165) & (g166)) + ((!g686) & (g691) & (g696) & (!g701) & (!g165) & (g166)) + ((!g686) & (g691) & (g696) & (!g701) & (g165) & (!g166)) + ((!g686) & (g691) & (g696) & (g701) & (!g165) & (g166)) + ((!g686) & (g691) & (g696) & (g701) & (g165) & (!g166)) + ((!g686) & (g691) & (g696) & (g701) & (g165) & (g166)) + ((g686) & (!g691) & (!g696) & (!g701) & (!g165) & (!g166)) + ((g686) & (!g691) & (!g696) & (g701) & (!g165) & (!g166)) + ((g686) & (!g691) & (!g696) & (g701) & (g165) & (g166)) + ((g686) & (!g691) & (g696) & (!g701) & (!g165) & (!g166)) + ((g686) & (!g691) & (g696) & (!g701) & (!g165) & (g166)) + ((g686) & (!g691) & (g696) & (g701) & (!g165) & (!g166)) + ((g686) & (!g691) & (g696) & (g701) & (!g165) & (g166)) + ((g686) & (!g691) & (g696) & (g701) & (g165) & (g166)) + ((g686) & (g691) & (!g696) & (!g701) & (!g165) & (!g166)) + ((g686) & (g691) & (!g696) & (!g701) & (g165) & (!g166)) + ((g686) & (g691) & (!g696) & (g701) & (!g165) & (!g166)) + ((g686) & (g691) & (!g696) & (g701) & (g165) & (!g166)) + ((g686) & (g691) & (!g696) & (g701) & (g165) & (g166)) + ((g686) & (g691) & (g696) & (!g701) & (!g165) & (!g166)) + ((g686) & (g691) & (g696) & (!g701) & (!g165) & (g166)) + ((g686) & (g691) & (g696) & (!g701) & (g165) & (!g166)) + ((g686) & (g691) & (g696) & (g701) & (!g165) & (!g166)) + ((g686) & (g691) & (g696) & (g701) & (!g165) & (g166)) + ((g686) & (g691) & (g696) & (g701) & (g165) & (!g166)) + ((g686) & (g691) & (g696) & (g701) & (g165) & (g166)));
	assign g4390 = (((!g2173) & (!g2473) & (!sk[1]) & (g703)) + ((!g2173) & (!g2473) & (sk[1]) & (g703)) + ((!g2173) & (g2473) & (!sk[1]) & (!g703)) + ((!g2173) & (g2473) & (!sk[1]) & (g703)) + ((!g2173) & (g2473) & (sk[1]) & (g703)) + ((g2173) & (!g2473) & (!sk[1]) & (g703)) + ((g2173) & (g2473) & (!sk[1]) & (!g703)) + ((g2173) & (g2473) & (!sk[1]) & (g703)) + ((g2173) & (g2473) & (sk[1]) & (!g703)) + ((g2173) & (g2473) & (sk[1]) & (g703)));
	assign g4391 = (((!g2174) & (!g2473) & (!sk[2]) & (g704)) + ((!g2174) & (!g2473) & (sk[2]) & (g704)) + ((!g2174) & (g2473) & (!sk[2]) & (!g704)) + ((!g2174) & (g2473) & (!sk[2]) & (g704)) + ((!g2174) & (g2473) & (sk[2]) & (g704)) + ((g2174) & (!g2473) & (!sk[2]) & (g704)) + ((g2174) & (g2473) & (!sk[2]) & (!g704)) + ((g2174) & (g2473) & (!sk[2]) & (g704)) + ((g2174) & (g2473) & (sk[2]) & (!g704)) + ((g2174) & (g2473) & (sk[2]) & (g704)));
	assign g4392 = (((!g2175) & (!sk[3]) & (!g2473) & (g705)) + ((!g2175) & (!sk[3]) & (g2473) & (!g705)) + ((!g2175) & (!sk[3]) & (g2473) & (g705)) + ((!g2175) & (sk[3]) & (!g2473) & (g705)) + ((!g2175) & (sk[3]) & (g2473) & (g705)) + ((g2175) & (!sk[3]) & (!g2473) & (g705)) + ((g2175) & (!sk[3]) & (g2473) & (!g705)) + ((g2175) & (!sk[3]) & (g2473) & (g705)) + ((g2175) & (sk[3]) & (g2473) & (!g705)) + ((g2175) & (sk[3]) & (g2473) & (g705)));
	assign g4393 = (((!sk[4]) & (!g2176) & (!g2473) & (g706)) + ((!sk[4]) & (!g2176) & (g2473) & (!g706)) + ((!sk[4]) & (!g2176) & (g2473) & (g706)) + ((!sk[4]) & (g2176) & (!g2473) & (g706)) + ((!sk[4]) & (g2176) & (g2473) & (!g706)) + ((!sk[4]) & (g2176) & (g2473) & (g706)) + ((sk[4]) & (!g2176) & (!g2473) & (g706)) + ((sk[4]) & (!g2176) & (g2473) & (g706)) + ((sk[4]) & (g2176) & (g2473) & (!g706)) + ((sk[4]) & (g2176) & (g2473) & (g706)));
	assign g707 = (((!g703) & (!g704) & (!g705) & (g706) & (g165) & (g166)) + ((!g703) & (!g704) & (g705) & (!g706) & (!g165) & (g166)) + ((!g703) & (!g704) & (g705) & (g706) & (!g165) & (g166)) + ((!g703) & (!g704) & (g705) & (g706) & (g165) & (g166)) + ((!g703) & (g704) & (!g705) & (!g706) & (g165) & (!g166)) + ((!g703) & (g704) & (!g705) & (g706) & (g165) & (!g166)) + ((!g703) & (g704) & (!g705) & (g706) & (g165) & (g166)) + ((!g703) & (g704) & (g705) & (!g706) & (!g165) & (g166)) + ((!g703) & (g704) & (g705) & (!g706) & (g165) & (!g166)) + ((!g703) & (g704) & (g705) & (g706) & (!g165) & (g166)) + ((!g703) & (g704) & (g705) & (g706) & (g165) & (!g166)) + ((!g703) & (g704) & (g705) & (g706) & (g165) & (g166)) + ((g703) & (!g704) & (!g705) & (!g706) & (!g165) & (!g166)) + ((g703) & (!g704) & (!g705) & (g706) & (!g165) & (!g166)) + ((g703) & (!g704) & (!g705) & (g706) & (g165) & (g166)) + ((g703) & (!g704) & (g705) & (!g706) & (!g165) & (!g166)) + ((g703) & (!g704) & (g705) & (!g706) & (!g165) & (g166)) + ((g703) & (!g704) & (g705) & (g706) & (!g165) & (!g166)) + ((g703) & (!g704) & (g705) & (g706) & (!g165) & (g166)) + ((g703) & (!g704) & (g705) & (g706) & (g165) & (g166)) + ((g703) & (g704) & (!g705) & (!g706) & (!g165) & (!g166)) + ((g703) & (g704) & (!g705) & (!g706) & (g165) & (!g166)) + ((g703) & (g704) & (!g705) & (g706) & (!g165) & (!g166)) + ((g703) & (g704) & (!g705) & (g706) & (g165) & (!g166)) + ((g703) & (g704) & (!g705) & (g706) & (g165) & (g166)) + ((g703) & (g704) & (g705) & (!g706) & (!g165) & (!g166)) + ((g703) & (g704) & (g705) & (!g706) & (!g165) & (g166)) + ((g703) & (g704) & (g705) & (!g706) & (g165) & (!g166)) + ((g703) & (g704) & (g705) & (g706) & (!g165) & (!g166)) + ((g703) & (g704) & (g705) & (g706) & (!g165) & (g166)) + ((g703) & (g704) & (g705) & (g706) & (g165) & (!g166)) + ((g703) & (g704) & (g705) & (g706) & (g165) & (g166)));
	assign g4394 = (((!sk[6]) & (!g2177) & (!g2473) & (g708)) + ((!sk[6]) & (!g2177) & (g2473) & (!g708)) + ((!sk[6]) & (!g2177) & (g2473) & (g708)) + ((!sk[6]) & (g2177) & (!g2473) & (g708)) + ((!sk[6]) & (g2177) & (g2473) & (!g708)) + ((!sk[6]) & (g2177) & (g2473) & (g708)) + ((sk[6]) & (!g2177) & (!g2473) & (g708)) + ((sk[6]) & (!g2177) & (g2473) & (g708)) + ((sk[6]) & (g2177) & (g2473) & (!g708)) + ((sk[6]) & (g2177) & (g2473) & (g708)));
	assign g4395 = (((!g2178) & (!g2473) & (!sk[7]) & (g709)) + ((!g2178) & (!g2473) & (sk[7]) & (g709)) + ((!g2178) & (g2473) & (!sk[7]) & (!g709)) + ((!g2178) & (g2473) & (!sk[7]) & (g709)) + ((!g2178) & (g2473) & (sk[7]) & (g709)) + ((g2178) & (!g2473) & (!sk[7]) & (g709)) + ((g2178) & (g2473) & (!sk[7]) & (!g709)) + ((g2178) & (g2473) & (!sk[7]) & (g709)) + ((g2178) & (g2473) & (sk[7]) & (!g709)) + ((g2178) & (g2473) & (sk[7]) & (g709)));
	assign g4396 = (((!sk[8]) & (!g2179) & (!g2473) & (g710)) + ((!sk[8]) & (!g2179) & (g2473) & (!g710)) + ((!sk[8]) & (!g2179) & (g2473) & (g710)) + ((!sk[8]) & (g2179) & (!g2473) & (g710)) + ((!sk[8]) & (g2179) & (g2473) & (!g710)) + ((!sk[8]) & (g2179) & (g2473) & (g710)) + ((sk[8]) & (!g2179) & (!g2473) & (g710)) + ((sk[8]) & (!g2179) & (g2473) & (g710)) + ((sk[8]) & (g2179) & (g2473) & (!g710)) + ((sk[8]) & (g2179) & (g2473) & (g710)));
	assign g711 = (((!g165) & (!g166) & (!sk[9]) & (!g708) & (g709) & (!g710)) + ((!g165) & (!g166) & (!sk[9]) & (!g708) & (g709) & (g710)) + ((!g165) & (!g166) & (!sk[9]) & (g708) & (!g709) & (!g710)) + ((!g165) & (!g166) & (!sk[9]) & (g708) & (!g709) & (g710)) + ((!g165) & (!g166) & (!sk[9]) & (g708) & (g709) & (!g710)) + ((!g165) & (!g166) & (!sk[9]) & (g708) & (g709) & (g710)) + ((!g165) & (g166) & (!sk[9]) & (!g708) & (!g709) & (!g710)) + ((!g165) & (g166) & (!sk[9]) & (!g708) & (!g709) & (g710)) + ((!g165) & (g166) & (!sk[9]) & (!g708) & (g709) & (!g710)) + ((!g165) & (g166) & (!sk[9]) & (!g708) & (g709) & (g710)) + ((!g165) & (g166) & (!sk[9]) & (g708) & (!g709) & (!g710)) + ((!g165) & (g166) & (!sk[9]) & (g708) & (!g709) & (g710)) + ((!g165) & (g166) & (!sk[9]) & (g708) & (g709) & (!g710)) + ((!g165) & (g166) & (!sk[9]) & (g708) & (g709) & (g710)) + ((!g165) & (g166) & (sk[9]) & (!g708) & (!g709) & (g710)) + ((!g165) & (g166) & (sk[9]) & (!g708) & (g709) & (g710)) + ((!g165) & (g166) & (sk[9]) & (g708) & (!g709) & (g710)) + ((!g165) & (g166) & (sk[9]) & (g708) & (g709) & (g710)) + ((g165) & (!g166) & (!sk[9]) & (!g708) & (g709) & (!g710)) + ((g165) & (!g166) & (!sk[9]) & (!g708) & (g709) & (g710)) + ((g165) & (!g166) & (!sk[9]) & (g708) & (!g709) & (!g710)) + ((g165) & (!g166) & (!sk[9]) & (g708) & (!g709) & (g710)) + ((g165) & (!g166) & (!sk[9]) & (g708) & (g709) & (!g710)) + ((g165) & (!g166) & (!sk[9]) & (g708) & (g709) & (g710)) + ((g165) & (!g166) & (sk[9]) & (g708) & (!g709) & (!g710)) + ((g165) & (!g166) & (sk[9]) & (g708) & (!g709) & (g710)) + ((g165) & (!g166) & (sk[9]) & (g708) & (g709) & (!g710)) + ((g165) & (!g166) & (sk[9]) & (g708) & (g709) & (g710)) + ((g165) & (g166) & (!sk[9]) & (!g708) & (!g709) & (!g710)) + ((g165) & (g166) & (!sk[9]) & (!g708) & (!g709) & (g710)) + ((g165) & (g166) & (!sk[9]) & (!g708) & (g709) & (!g710)) + ((g165) & (g166) & (!sk[9]) & (!g708) & (g709) & (g710)) + ((g165) & (g166) & (!sk[9]) & (g708) & (!g709) & (!g710)) + ((g165) & (g166) & (!sk[9]) & (g708) & (!g709) & (g710)) + ((g165) & (g166) & (!sk[9]) & (g708) & (g709) & (!g710)) + ((g165) & (g166) & (!sk[9]) & (g708) & (g709) & (g710)) + ((g165) & (g166) & (sk[9]) & (!g708) & (g709) & (!g710)) + ((g165) & (g166) & (sk[9]) & (!g708) & (g709) & (g710)) + ((g165) & (g166) & (sk[9]) & (g708) & (g709) & (!g710)) + ((g165) & (g166) & (sk[9]) & (g708) & (g709) & (g710)));
	assign g4397 = (((!g2162) & (!sk[10]) & (!g2473) & (g712)) + ((!g2162) & (!sk[10]) & (g2473) & (!g712)) + ((!g2162) & (!sk[10]) & (g2473) & (g712)) + ((!g2162) & (sk[10]) & (!g2473) & (g712)) + ((!g2162) & (sk[10]) & (g2473) & (g712)) + ((g2162) & (!sk[10]) & (!g2473) & (g712)) + ((g2162) & (!sk[10]) & (g2473) & (!g712)) + ((g2162) & (!sk[10]) & (g2473) & (g712)) + ((g2162) & (sk[10]) & (g2473) & (!g712)) + ((g2162) & (sk[10]) & (g2473) & (g712)));
	assign g4398 = (((!g2164) & (!sk[11]) & (!g2473) & (g713)) + ((!g2164) & (!sk[11]) & (g2473) & (!g713)) + ((!g2164) & (!sk[11]) & (g2473) & (g713)) + ((!g2164) & (sk[11]) & (!g2473) & (g713)) + ((!g2164) & (sk[11]) & (g2473) & (g713)) + ((g2164) & (!sk[11]) & (!g2473) & (g713)) + ((g2164) & (!sk[11]) & (g2473) & (!g713)) + ((g2164) & (!sk[11]) & (g2473) & (g713)) + ((g2164) & (sk[11]) & (g2473) & (!g713)) + ((g2164) & (sk[11]) & (g2473) & (g713)));
	assign g4399 = (((!g2166) & (!sk[12]) & (!g2473) & (g714)) + ((!g2166) & (!sk[12]) & (g2473) & (!g714)) + ((!g2166) & (!sk[12]) & (g2473) & (g714)) + ((!g2166) & (sk[12]) & (!g2473) & (g714)) + ((!g2166) & (sk[12]) & (g2473) & (g714)) + ((g2166) & (!sk[12]) & (!g2473) & (g714)) + ((g2166) & (!sk[12]) & (g2473) & (!g714)) + ((g2166) & (!sk[12]) & (g2473) & (g714)) + ((g2166) & (sk[12]) & (g2473) & (!g714)) + ((g2166) & (sk[12]) & (g2473) & (g714)));
	assign g4400 = (((!g2168) & (!sk[13]) & (!g2473) & (g715)) + ((!g2168) & (!sk[13]) & (g2473) & (!g715)) + ((!g2168) & (!sk[13]) & (g2473) & (g715)) + ((!g2168) & (sk[13]) & (!g2473) & (g715)) + ((!g2168) & (sk[13]) & (g2473) & (g715)) + ((g2168) & (!sk[13]) & (!g2473) & (g715)) + ((g2168) & (!sk[13]) & (g2473) & (!g715)) + ((g2168) & (!sk[13]) & (g2473) & (g715)) + ((g2168) & (sk[13]) & (g2473) & (!g715)) + ((g2168) & (sk[13]) & (g2473) & (g715)));
	assign g716 = (((!g712) & (!g713) & (!g714) & (g715) & (g165) & (g166)) + ((!g712) & (!g713) & (g714) & (!g715) & (!g165) & (g166)) + ((!g712) & (!g713) & (g714) & (g715) & (!g165) & (g166)) + ((!g712) & (!g713) & (g714) & (g715) & (g165) & (g166)) + ((!g712) & (g713) & (!g714) & (!g715) & (g165) & (!g166)) + ((!g712) & (g713) & (!g714) & (g715) & (g165) & (!g166)) + ((!g712) & (g713) & (!g714) & (g715) & (g165) & (g166)) + ((!g712) & (g713) & (g714) & (!g715) & (!g165) & (g166)) + ((!g712) & (g713) & (g714) & (!g715) & (g165) & (!g166)) + ((!g712) & (g713) & (g714) & (g715) & (!g165) & (g166)) + ((!g712) & (g713) & (g714) & (g715) & (g165) & (!g166)) + ((!g712) & (g713) & (g714) & (g715) & (g165) & (g166)) + ((g712) & (!g713) & (!g714) & (!g715) & (!g165) & (!g166)) + ((g712) & (!g713) & (!g714) & (g715) & (!g165) & (!g166)) + ((g712) & (!g713) & (!g714) & (g715) & (g165) & (g166)) + ((g712) & (!g713) & (g714) & (!g715) & (!g165) & (!g166)) + ((g712) & (!g713) & (g714) & (!g715) & (!g165) & (g166)) + ((g712) & (!g713) & (g714) & (g715) & (!g165) & (!g166)) + ((g712) & (!g713) & (g714) & (g715) & (!g165) & (g166)) + ((g712) & (!g713) & (g714) & (g715) & (g165) & (g166)) + ((g712) & (g713) & (!g714) & (!g715) & (!g165) & (!g166)) + ((g712) & (g713) & (!g714) & (!g715) & (g165) & (!g166)) + ((g712) & (g713) & (!g714) & (g715) & (!g165) & (!g166)) + ((g712) & (g713) & (!g714) & (g715) & (g165) & (!g166)) + ((g712) & (g713) & (!g714) & (g715) & (g165) & (g166)) + ((g712) & (g713) & (g714) & (!g715) & (!g165) & (!g166)) + ((g712) & (g713) & (g714) & (!g715) & (!g165) & (g166)) + ((g712) & (g713) & (g714) & (!g715) & (g165) & (!g166)) + ((g712) & (g713) & (g714) & (g715) & (!g165) & (!g166)) + ((g712) & (g713) & (g714) & (g715) & (!g165) & (g166)) + ((g712) & (g713) & (g714) & (g715) & (g165) & (!g166)) + ((g712) & (g713) & (g714) & (g715) & (g165) & (g166)));
	assign g4401 = (((!sk[15]) & (!g2169) & (!g2473) & (g717)) + ((!sk[15]) & (!g2169) & (g2473) & (!g717)) + ((!sk[15]) & (!g2169) & (g2473) & (g717)) + ((!sk[15]) & (g2169) & (!g2473) & (g717)) + ((!sk[15]) & (g2169) & (g2473) & (!g717)) + ((!sk[15]) & (g2169) & (g2473) & (g717)) + ((sk[15]) & (!g2169) & (!g2473) & (g717)) + ((sk[15]) & (!g2169) & (g2473) & (g717)) + ((sk[15]) & (g2169) & (g2473) & (!g717)) + ((sk[15]) & (g2169) & (g2473) & (g717)));
	assign g4402 = (((!sk[16]) & (!g2170) & (!g2473) & (g718)) + ((!sk[16]) & (!g2170) & (g2473) & (!g718)) + ((!sk[16]) & (!g2170) & (g2473) & (g718)) + ((!sk[16]) & (g2170) & (!g2473) & (g718)) + ((!sk[16]) & (g2170) & (g2473) & (!g718)) + ((!sk[16]) & (g2170) & (g2473) & (g718)) + ((sk[16]) & (!g2170) & (!g2473) & (g718)) + ((sk[16]) & (!g2170) & (g2473) & (g718)) + ((sk[16]) & (g2170) & (g2473) & (!g718)) + ((sk[16]) & (g2170) & (g2473) & (g718)));
	assign g4403 = (((!g2171) & (!g2473) & (!sk[17]) & (g719)) + ((!g2171) & (!g2473) & (sk[17]) & (g719)) + ((!g2171) & (g2473) & (!sk[17]) & (!g719)) + ((!g2171) & (g2473) & (!sk[17]) & (g719)) + ((!g2171) & (g2473) & (sk[17]) & (g719)) + ((g2171) & (!g2473) & (!sk[17]) & (g719)) + ((g2171) & (g2473) & (!sk[17]) & (!g719)) + ((g2171) & (g2473) & (!sk[17]) & (g719)) + ((g2171) & (g2473) & (sk[17]) & (!g719)) + ((g2171) & (g2473) & (sk[17]) & (g719)));
	assign g4404 = (((!g2172) & (!sk[18]) & (!g2473) & (g720)) + ((!g2172) & (!sk[18]) & (g2473) & (!g720)) + ((!g2172) & (!sk[18]) & (g2473) & (g720)) + ((!g2172) & (sk[18]) & (!g2473) & (g720)) + ((!g2172) & (sk[18]) & (g2473) & (g720)) + ((g2172) & (!sk[18]) & (!g2473) & (g720)) + ((g2172) & (!sk[18]) & (g2473) & (!g720)) + ((g2172) & (!sk[18]) & (g2473) & (g720)) + ((g2172) & (sk[18]) & (g2473) & (!g720)) + ((g2172) & (sk[18]) & (g2473) & (g720)));
	assign g721 = (((!g717) & (!g718) & (!g719) & (g720) & (g165) & (g166)) + ((!g717) & (!g718) & (g719) & (!g720) & (!g165) & (g166)) + ((!g717) & (!g718) & (g719) & (g720) & (!g165) & (g166)) + ((!g717) & (!g718) & (g719) & (g720) & (g165) & (g166)) + ((!g717) & (g718) & (!g719) & (!g720) & (g165) & (!g166)) + ((!g717) & (g718) & (!g719) & (g720) & (g165) & (!g166)) + ((!g717) & (g718) & (!g719) & (g720) & (g165) & (g166)) + ((!g717) & (g718) & (g719) & (!g720) & (!g165) & (g166)) + ((!g717) & (g718) & (g719) & (!g720) & (g165) & (!g166)) + ((!g717) & (g718) & (g719) & (g720) & (!g165) & (g166)) + ((!g717) & (g718) & (g719) & (g720) & (g165) & (!g166)) + ((!g717) & (g718) & (g719) & (g720) & (g165) & (g166)) + ((g717) & (!g718) & (!g719) & (!g720) & (!g165) & (!g166)) + ((g717) & (!g718) & (!g719) & (g720) & (!g165) & (!g166)) + ((g717) & (!g718) & (!g719) & (g720) & (g165) & (g166)) + ((g717) & (!g718) & (g719) & (!g720) & (!g165) & (!g166)) + ((g717) & (!g718) & (g719) & (!g720) & (!g165) & (g166)) + ((g717) & (!g718) & (g719) & (g720) & (!g165) & (!g166)) + ((g717) & (!g718) & (g719) & (g720) & (!g165) & (g166)) + ((g717) & (!g718) & (g719) & (g720) & (g165) & (g166)) + ((g717) & (g718) & (!g719) & (!g720) & (!g165) & (!g166)) + ((g717) & (g718) & (!g719) & (!g720) & (g165) & (!g166)) + ((g717) & (g718) & (!g719) & (g720) & (!g165) & (!g166)) + ((g717) & (g718) & (!g719) & (g720) & (g165) & (!g166)) + ((g717) & (g718) & (!g719) & (g720) & (g165) & (g166)) + ((g717) & (g718) & (g719) & (!g720) & (!g165) & (!g166)) + ((g717) & (g718) & (g719) & (!g720) & (!g165) & (g166)) + ((g717) & (g718) & (g719) & (!g720) & (g165) & (!g166)) + ((g717) & (g718) & (g719) & (g720) & (!g165) & (!g166)) + ((g717) & (g718) & (g719) & (g720) & (!g165) & (g166)) + ((g717) & (g718) & (g719) & (g720) & (g165) & (!g166)) + ((g717) & (g718) & (g719) & (g720) & (g165) & (g166)));
	assign g722 = (((!g147) & (!g148) & (!g707) & (g711) & (!g716) & (!g721)) + ((!g147) & (!g148) & (!g707) & (g711) & (!g716) & (g721)) + ((!g147) & (!g148) & (!g707) & (g711) & (g716) & (!g721)) + ((!g147) & (!g148) & (!g707) & (g711) & (g716) & (g721)) + ((!g147) & (!g148) & (g707) & (g711) & (!g716) & (!g721)) + ((!g147) & (!g148) & (g707) & (g711) & (!g716) & (g721)) + ((!g147) & (!g148) & (g707) & (g711) & (g716) & (!g721)) + ((!g147) & (!g148) & (g707) & (g711) & (g716) & (g721)) + ((!g147) & (g148) & (!g707) & (!g711) & (!g716) & (g721)) + ((!g147) & (g148) & (!g707) & (!g711) & (g716) & (g721)) + ((!g147) & (g148) & (!g707) & (g711) & (!g716) & (g721)) + ((!g147) & (g148) & (!g707) & (g711) & (g716) & (g721)) + ((!g147) & (g148) & (g707) & (!g711) & (!g716) & (g721)) + ((!g147) & (g148) & (g707) & (!g711) & (g716) & (g721)) + ((!g147) & (g148) & (g707) & (g711) & (!g716) & (g721)) + ((!g147) & (g148) & (g707) & (g711) & (g716) & (g721)) + ((g147) & (!g148) & (g707) & (!g711) & (!g716) & (!g721)) + ((g147) & (!g148) & (g707) & (!g711) & (!g716) & (g721)) + ((g147) & (!g148) & (g707) & (!g711) & (g716) & (!g721)) + ((g147) & (!g148) & (g707) & (!g711) & (g716) & (g721)) + ((g147) & (!g148) & (g707) & (g711) & (!g716) & (!g721)) + ((g147) & (!g148) & (g707) & (g711) & (!g716) & (g721)) + ((g147) & (!g148) & (g707) & (g711) & (g716) & (!g721)) + ((g147) & (!g148) & (g707) & (g711) & (g716) & (g721)) + ((g147) & (g148) & (!g707) & (!g711) & (g716) & (!g721)) + ((g147) & (g148) & (!g707) & (!g711) & (g716) & (g721)) + ((g147) & (g148) & (!g707) & (g711) & (g716) & (!g721)) + ((g147) & (g148) & (!g707) & (g711) & (g716) & (g721)) + ((g147) & (g148) & (g707) & (!g711) & (g716) & (!g721)) + ((g147) & (g148) & (g707) & (!g711) & (g716) & (g721)) + ((g147) & (g148) & (g707) & (g711) & (g716) & (!g721)) + ((g147) & (g148) & (g707) & (g711) & (g716) & (g721)));
	assign g723 = (((!g142) & (!g702) & (!sk[21]) & (g722)) + ((!g142) & (!g702) & (sk[21]) & (g722)) + ((!g142) & (g702) & (!sk[21]) & (!g722)) + ((!g142) & (g702) & (!sk[21]) & (g722)) + ((!g142) & (g702) & (sk[21]) & (g722)) + ((g142) & (!g702) & (!sk[21]) & (g722)) + ((g142) & (g702) & (!sk[21]) & (!g722)) + ((g142) & (g702) & (!sk[21]) & (g722)) + ((g142) & (g702) & (sk[21]) & (!g722)) + ((g142) & (g702) & (sk[21]) & (g722)));
	assign g4405 = (((!g2059) & (!g2479) & (!sk[22]) & (g724)) + ((!g2059) & (!g2479) & (sk[22]) & (g724)) + ((!g2059) & (g2479) & (!sk[22]) & (!g724)) + ((!g2059) & (g2479) & (!sk[22]) & (g724)) + ((!g2059) & (g2479) & (sk[22]) & (g724)) + ((g2059) & (!g2479) & (!sk[22]) & (g724)) + ((g2059) & (g2479) & (!sk[22]) & (!g724)) + ((g2059) & (g2479) & (!sk[22]) & (g724)) + ((g2059) & (g2479) & (sk[22]) & (!g724)) + ((g2059) & (g2479) & (sk[22]) & (g724)));
	assign g725 = (((!g672) & (!g676) & (!sk[23]) & (g680)) + ((!g672) & (!g676) & (sk[23]) & (!g680)) + ((!g672) & (g676) & (!sk[23]) & (!g680)) + ((!g672) & (g676) & (!sk[23]) & (g680)) + ((g672) & (!g676) & (!sk[23]) & (g680)) + ((g672) & (!g676) & (sk[23]) & (!g680)) + ((g672) & (!g676) & (sk[23]) & (g680)) + ((g672) & (g676) & (!sk[23]) & (!g680)) + ((g672) & (g676) & (!sk[23]) & (g680)) + ((g672) & (g676) & (sk[23]) & (!g680)));
	assign g4406 = (((!sk[24]) & (!g2064) & (!dmem_dat_ix12x) & (g726)) + ((!sk[24]) & (!g2064) & (dmem_dat_ix12x) & (!g726)) + ((!sk[24]) & (!g2064) & (dmem_dat_ix12x) & (g726)) + ((!sk[24]) & (g2064) & (!dmem_dat_ix12x) & (g726)) + ((!sk[24]) & (g2064) & (dmem_dat_ix12x) & (!g726)) + ((!sk[24]) & (g2064) & (dmem_dat_ix12x) & (g726)) + ((sk[24]) & (!g2064) & (!dmem_dat_ix12x) & (g726)) + ((sk[24]) & (!g2064) & (dmem_dat_ix12x) & (g726)) + ((sk[24]) & (g2064) & (dmem_dat_ix12x) & (!g726)) + ((sk[24]) & (g2064) & (dmem_dat_ix12x) & (g726)));
	assign g727 = (((!sk[25]) & (!g679) & (!g109) & (g726)) + ((!sk[25]) & (!g679) & (g109) & (!g726)) + ((!sk[25]) & (!g679) & (g109) & (g726)) + ((!sk[25]) & (g679) & (!g109) & (g726)) + ((!sk[25]) & (g679) & (g109) & (!g726)) + ((!sk[25]) & (g679) & (g109) & (g726)) + ((sk[25]) & (!g679) & (!g109) & (!g726)) + ((sk[25]) & (!g679) & (!g109) & (g726)) + ((sk[25]) & (g679) & (!g109) & (!g726)) + ((sk[25]) & (g679) & (g109) & (!g726)));
	assign g728 = (((!sk[26]) & (!g126) & (!g723) & (!g724) & (g725) & (!g727)) + ((!sk[26]) & (!g126) & (!g723) & (!g724) & (g725) & (g727)) + ((!sk[26]) & (!g126) & (!g723) & (g724) & (!g725) & (!g727)) + ((!sk[26]) & (!g126) & (!g723) & (g724) & (!g725) & (g727)) + ((!sk[26]) & (!g126) & (!g723) & (g724) & (g725) & (!g727)) + ((!sk[26]) & (!g126) & (!g723) & (g724) & (g725) & (g727)) + ((!sk[26]) & (!g126) & (g723) & (!g724) & (!g725) & (!g727)) + ((!sk[26]) & (!g126) & (g723) & (!g724) & (!g725) & (g727)) + ((!sk[26]) & (!g126) & (g723) & (!g724) & (g725) & (!g727)) + ((!sk[26]) & (!g126) & (g723) & (!g724) & (g725) & (g727)) + ((!sk[26]) & (!g126) & (g723) & (g724) & (!g725) & (!g727)) + ((!sk[26]) & (!g126) & (g723) & (g724) & (!g725) & (g727)) + ((!sk[26]) & (!g126) & (g723) & (g724) & (g725) & (!g727)) + ((!sk[26]) & (!g126) & (g723) & (g724) & (g725) & (g727)) + ((!sk[26]) & (g126) & (!g723) & (!g724) & (g725) & (!g727)) + ((!sk[26]) & (g126) & (!g723) & (!g724) & (g725) & (g727)) + ((!sk[26]) & (g126) & (!g723) & (g724) & (!g725) & (!g727)) + ((!sk[26]) & (g126) & (!g723) & (g724) & (!g725) & (g727)) + ((!sk[26]) & (g126) & (!g723) & (g724) & (g725) & (!g727)) + ((!sk[26]) & (g126) & (!g723) & (g724) & (g725) & (g727)) + ((!sk[26]) & (g126) & (g723) & (!g724) & (!g725) & (!g727)) + ((!sk[26]) & (g126) & (g723) & (!g724) & (!g725) & (g727)) + ((!sk[26]) & (g126) & (g723) & (!g724) & (g725) & (!g727)) + ((!sk[26]) & (g126) & (g723) & (!g724) & (g725) & (g727)) + ((!sk[26]) & (g126) & (g723) & (g724) & (!g725) & (!g727)) + ((!sk[26]) & (g126) & (g723) & (g724) & (!g725) & (g727)) + ((!sk[26]) & (g126) & (g723) & (g724) & (g725) & (!g727)) + ((!sk[26]) & (g126) & (g723) & (g724) & (g725) & (g727)) + ((sk[26]) & (!g126) & (!g723) & (g724) & (!g725) & (!g727)) + ((sk[26]) & (!g126) & (!g723) & (g724) & (!g725) & (g727)) + ((sk[26]) & (!g126) & (!g723) & (g724) & (g725) & (!g727)) + ((sk[26]) & (!g126) & (!g723) & (g724) & (g725) & (g727)) + ((sk[26]) & (!g126) & (g723) & (g724) & (!g725) & (!g727)) + ((sk[26]) & (!g126) & (g723) & (g724) & (!g725) & (g727)) + ((sk[26]) & (!g126) & (g723) & (g724) & (g725) & (!g727)) + ((sk[26]) & (!g126) & (g723) & (g724) & (g725) & (g727)) + ((sk[26]) & (g126) & (!g723) & (!g724) & (!g725) & (!g727)) + ((sk[26]) & (g126) & (!g723) & (!g724) & (g725) & (g727)) + ((sk[26]) & (g126) & (!g723) & (g724) & (!g725) & (!g727)) + ((sk[26]) & (g126) & (!g723) & (g724) & (g725) & (g727)) + ((sk[26]) & (g126) & (g723) & (!g724) & (!g725) & (g727)) + ((sk[26]) & (g126) & (g723) & (!g724) & (g725) & (!g727)) + ((sk[26]) & (g126) & (g723) & (g724) & (!g725) & (g727)) + ((sk[26]) & (g126) & (g723) & (g724) & (g725) & (!g727)));
	assign g4407 = (((!sk[27]) & (!g2140) & (!g2495) & (g729)) + ((!sk[27]) & (!g2140) & (g2495) & (!g729)) + ((!sk[27]) & (!g2140) & (g2495) & (g729)) + ((!sk[27]) & (g2140) & (!g2495) & (g729)) + ((!sk[27]) & (g2140) & (g2495) & (!g729)) + ((!sk[27]) & (g2140) & (g2495) & (g729)) + ((sk[27]) & (!g2140) & (!g2495) & (g729)) + ((sk[27]) & (!g2140) & (g2495) & (g729)) + ((sk[27]) & (g2140) & (g2495) & (!g729)) + ((sk[27]) & (g2140) & (g2495) & (g729)));
	assign g4408 = (((!sk[28]) & (!g2142) & (!g2495) & (g730)) + ((!sk[28]) & (!g2142) & (g2495) & (!g730)) + ((!sk[28]) & (!g2142) & (g2495) & (g730)) + ((!sk[28]) & (g2142) & (!g2495) & (g730)) + ((!sk[28]) & (g2142) & (g2495) & (!g730)) + ((!sk[28]) & (g2142) & (g2495) & (g730)) + ((sk[28]) & (!g2142) & (!g2495) & (g730)) + ((sk[28]) & (!g2142) & (g2495) & (g730)) + ((sk[28]) & (g2142) & (g2495) & (!g730)) + ((sk[28]) & (g2142) & (g2495) & (g730)));
	assign g4409 = (((!g2144) & (!g2495) & (!sk[29]) & (g731)) + ((!g2144) & (!g2495) & (sk[29]) & (g731)) + ((!g2144) & (g2495) & (!sk[29]) & (!g731)) + ((!g2144) & (g2495) & (!sk[29]) & (g731)) + ((!g2144) & (g2495) & (sk[29]) & (g731)) + ((g2144) & (!g2495) & (!sk[29]) & (g731)) + ((g2144) & (g2495) & (!sk[29]) & (!g731)) + ((g2144) & (g2495) & (!sk[29]) & (g731)) + ((g2144) & (g2495) & (sk[29]) & (!g731)) + ((g2144) & (g2495) & (sk[29]) & (g731)));
	assign g4410 = (((!g2145) & (!g2495) & (!sk[30]) & (g732)) + ((!g2145) & (!g2495) & (sk[30]) & (g732)) + ((!g2145) & (g2495) & (!sk[30]) & (!g732)) + ((!g2145) & (g2495) & (!sk[30]) & (g732)) + ((!g2145) & (g2495) & (sk[30]) & (g732)) + ((g2145) & (!g2495) & (!sk[30]) & (g732)) + ((g2145) & (g2495) & (!sk[30]) & (!g732)) + ((g2145) & (g2495) & (!sk[30]) & (g732)) + ((g2145) & (g2495) & (sk[30]) & (!g732)) + ((g2145) & (g2495) & (sk[30]) & (g732)));
	assign g733 = (((!g729) & (!g730) & (!g731) & (g732) & (g147) & (g148)) + ((!g729) & (!g730) & (g731) & (!g732) & (!g147) & (g148)) + ((!g729) & (!g730) & (g731) & (g732) & (!g147) & (g148)) + ((!g729) & (!g730) & (g731) & (g732) & (g147) & (g148)) + ((!g729) & (g730) & (!g731) & (!g732) & (g147) & (!g148)) + ((!g729) & (g730) & (!g731) & (g732) & (g147) & (!g148)) + ((!g729) & (g730) & (!g731) & (g732) & (g147) & (g148)) + ((!g729) & (g730) & (g731) & (!g732) & (!g147) & (g148)) + ((!g729) & (g730) & (g731) & (!g732) & (g147) & (!g148)) + ((!g729) & (g730) & (g731) & (g732) & (!g147) & (g148)) + ((!g729) & (g730) & (g731) & (g732) & (g147) & (!g148)) + ((!g729) & (g730) & (g731) & (g732) & (g147) & (g148)) + ((g729) & (!g730) & (!g731) & (!g732) & (!g147) & (!g148)) + ((g729) & (!g730) & (!g731) & (g732) & (!g147) & (!g148)) + ((g729) & (!g730) & (!g731) & (g732) & (g147) & (g148)) + ((g729) & (!g730) & (g731) & (!g732) & (!g147) & (!g148)) + ((g729) & (!g730) & (g731) & (!g732) & (!g147) & (g148)) + ((g729) & (!g730) & (g731) & (g732) & (!g147) & (!g148)) + ((g729) & (!g730) & (g731) & (g732) & (!g147) & (g148)) + ((g729) & (!g730) & (g731) & (g732) & (g147) & (g148)) + ((g729) & (g730) & (!g731) & (!g732) & (!g147) & (!g148)) + ((g729) & (g730) & (!g731) & (!g732) & (g147) & (!g148)) + ((g729) & (g730) & (!g731) & (g732) & (!g147) & (!g148)) + ((g729) & (g730) & (!g731) & (g732) & (g147) & (!g148)) + ((g729) & (g730) & (!g731) & (g732) & (g147) & (g148)) + ((g729) & (g730) & (g731) & (!g732) & (!g147) & (!g148)) + ((g729) & (g730) & (g731) & (!g732) & (!g147) & (g148)) + ((g729) & (g730) & (g731) & (!g732) & (g147) & (!g148)) + ((g729) & (g730) & (g731) & (g732) & (!g147) & (!g148)) + ((g729) & (g730) & (g731) & (g732) & (!g147) & (g148)) + ((g729) & (g730) & (g731) & (g732) & (g147) & (!g148)) + ((g729) & (g730) & (g731) & (g732) & (g147) & (g148)));
	assign g4411 = (((!g2146) & (!sk[32]) & (!g2495) & (g734)) + ((!g2146) & (!sk[32]) & (g2495) & (!g734)) + ((!g2146) & (!sk[32]) & (g2495) & (g734)) + ((!g2146) & (sk[32]) & (!g2495) & (g734)) + ((!g2146) & (sk[32]) & (g2495) & (g734)) + ((g2146) & (!sk[32]) & (!g2495) & (g734)) + ((g2146) & (!sk[32]) & (g2495) & (!g734)) + ((g2146) & (!sk[32]) & (g2495) & (g734)) + ((g2146) & (sk[32]) & (g2495) & (!g734)) + ((g2146) & (sk[32]) & (g2495) & (g734)));
	assign g4412 = (((!sk[33]) & (!g2148) & (!g2495) & (g735)) + ((!sk[33]) & (!g2148) & (g2495) & (!g735)) + ((!sk[33]) & (!g2148) & (g2495) & (g735)) + ((!sk[33]) & (g2148) & (!g2495) & (g735)) + ((!sk[33]) & (g2148) & (g2495) & (!g735)) + ((!sk[33]) & (g2148) & (g2495) & (g735)) + ((sk[33]) & (!g2148) & (!g2495) & (g735)) + ((sk[33]) & (!g2148) & (g2495) & (g735)) + ((sk[33]) & (g2148) & (g2495) & (!g735)) + ((sk[33]) & (g2148) & (g2495) & (g735)));
	assign g4413 = (((!g2150) & (!g2495) & (!sk[34]) & (g736)) + ((!g2150) & (!g2495) & (sk[34]) & (g736)) + ((!g2150) & (g2495) & (!sk[34]) & (!g736)) + ((!g2150) & (g2495) & (!sk[34]) & (g736)) + ((!g2150) & (g2495) & (sk[34]) & (g736)) + ((g2150) & (!g2495) & (!sk[34]) & (g736)) + ((g2150) & (g2495) & (!sk[34]) & (!g736)) + ((g2150) & (g2495) & (!sk[34]) & (g736)) + ((g2150) & (g2495) & (sk[34]) & (!g736)) + ((g2150) & (g2495) & (sk[34]) & (g736)));
	assign g4414 = (((!sk[35]) & (!g2151) & (!g2495) & (g737)) + ((!sk[35]) & (!g2151) & (g2495) & (!g737)) + ((!sk[35]) & (!g2151) & (g2495) & (g737)) + ((!sk[35]) & (g2151) & (!g2495) & (g737)) + ((!sk[35]) & (g2151) & (g2495) & (!g737)) + ((!sk[35]) & (g2151) & (g2495) & (g737)) + ((sk[35]) & (!g2151) & (!g2495) & (g737)) + ((sk[35]) & (!g2151) & (g2495) & (g737)) + ((sk[35]) & (g2151) & (g2495) & (!g737)) + ((sk[35]) & (g2151) & (g2495) & (g737)));
	assign g738 = (((!g734) & (!g735) & (!g736) & (g737) & (g147) & (g148)) + ((!g734) & (!g735) & (g736) & (!g737) & (!g147) & (g148)) + ((!g734) & (!g735) & (g736) & (g737) & (!g147) & (g148)) + ((!g734) & (!g735) & (g736) & (g737) & (g147) & (g148)) + ((!g734) & (g735) & (!g736) & (!g737) & (g147) & (!g148)) + ((!g734) & (g735) & (!g736) & (g737) & (g147) & (!g148)) + ((!g734) & (g735) & (!g736) & (g737) & (g147) & (g148)) + ((!g734) & (g735) & (g736) & (!g737) & (!g147) & (g148)) + ((!g734) & (g735) & (g736) & (!g737) & (g147) & (!g148)) + ((!g734) & (g735) & (g736) & (g737) & (!g147) & (g148)) + ((!g734) & (g735) & (g736) & (g737) & (g147) & (!g148)) + ((!g734) & (g735) & (g736) & (g737) & (g147) & (g148)) + ((g734) & (!g735) & (!g736) & (!g737) & (!g147) & (!g148)) + ((g734) & (!g735) & (!g736) & (g737) & (!g147) & (!g148)) + ((g734) & (!g735) & (!g736) & (g737) & (g147) & (g148)) + ((g734) & (!g735) & (g736) & (!g737) & (!g147) & (!g148)) + ((g734) & (!g735) & (g736) & (!g737) & (!g147) & (g148)) + ((g734) & (!g735) & (g736) & (g737) & (!g147) & (!g148)) + ((g734) & (!g735) & (g736) & (g737) & (!g147) & (g148)) + ((g734) & (!g735) & (g736) & (g737) & (g147) & (g148)) + ((g734) & (g735) & (!g736) & (!g737) & (!g147) & (!g148)) + ((g734) & (g735) & (!g736) & (!g737) & (g147) & (!g148)) + ((g734) & (g735) & (!g736) & (g737) & (!g147) & (!g148)) + ((g734) & (g735) & (!g736) & (g737) & (g147) & (!g148)) + ((g734) & (g735) & (!g736) & (g737) & (g147) & (g148)) + ((g734) & (g735) & (g736) & (!g737) & (!g147) & (!g148)) + ((g734) & (g735) & (g736) & (!g737) & (!g147) & (g148)) + ((g734) & (g735) & (g736) & (!g737) & (g147) & (!g148)) + ((g734) & (g735) & (g736) & (g737) & (!g147) & (!g148)) + ((g734) & (g735) & (g736) & (g737) & (!g147) & (g148)) + ((g734) & (g735) & (g736) & (g737) & (g147) & (!g148)) + ((g734) & (g735) & (g736) & (g737) & (g147) & (g148)));
	assign g4415 = (((!g2152) & (!sk[37]) & (!g2495) & (g739)) + ((!g2152) & (!sk[37]) & (g2495) & (!g739)) + ((!g2152) & (!sk[37]) & (g2495) & (g739)) + ((!g2152) & (sk[37]) & (!g2495) & (g739)) + ((!g2152) & (sk[37]) & (g2495) & (g739)) + ((g2152) & (!sk[37]) & (!g2495) & (g739)) + ((g2152) & (!sk[37]) & (g2495) & (!g739)) + ((g2152) & (!sk[37]) & (g2495) & (g739)) + ((g2152) & (sk[37]) & (g2495) & (!g739)) + ((g2152) & (sk[37]) & (g2495) & (g739)));
	assign g4416 = (((!g2153) & (!sk[38]) & (!g2495) & (g740)) + ((!g2153) & (!sk[38]) & (g2495) & (!g740)) + ((!g2153) & (!sk[38]) & (g2495) & (g740)) + ((!g2153) & (sk[38]) & (!g2495) & (g740)) + ((!g2153) & (sk[38]) & (g2495) & (g740)) + ((g2153) & (!sk[38]) & (!g2495) & (g740)) + ((g2153) & (!sk[38]) & (g2495) & (!g740)) + ((g2153) & (!sk[38]) & (g2495) & (g740)) + ((g2153) & (sk[38]) & (g2495) & (!g740)) + ((g2153) & (sk[38]) & (g2495) & (g740)));
	assign g4417 = (((!g2155) & (!g2495) & (!sk[39]) & (g741)) + ((!g2155) & (!g2495) & (sk[39]) & (g741)) + ((!g2155) & (g2495) & (!sk[39]) & (!g741)) + ((!g2155) & (g2495) & (!sk[39]) & (g741)) + ((!g2155) & (g2495) & (sk[39]) & (g741)) + ((g2155) & (!g2495) & (!sk[39]) & (g741)) + ((g2155) & (g2495) & (!sk[39]) & (!g741)) + ((g2155) & (g2495) & (!sk[39]) & (g741)) + ((g2155) & (g2495) & (sk[39]) & (!g741)) + ((g2155) & (g2495) & (sk[39]) & (g741)));
	assign g4418 = (((!g2157) & (!sk[40]) & (!g2495) & (g742)) + ((!g2157) & (!sk[40]) & (g2495) & (!g742)) + ((!g2157) & (!sk[40]) & (g2495) & (g742)) + ((!g2157) & (sk[40]) & (!g2495) & (g742)) + ((!g2157) & (sk[40]) & (g2495) & (g742)) + ((g2157) & (!sk[40]) & (!g2495) & (g742)) + ((g2157) & (!sk[40]) & (g2495) & (!g742)) + ((g2157) & (!sk[40]) & (g2495) & (g742)) + ((g2157) & (sk[40]) & (g2495) & (!g742)) + ((g2157) & (sk[40]) & (g2495) & (g742)));
	assign g743 = (((!g739) & (!g740) & (!g741) & (g742) & (g147) & (g148)) + ((!g739) & (!g740) & (g741) & (!g742) & (!g147) & (g148)) + ((!g739) & (!g740) & (g741) & (g742) & (!g147) & (g148)) + ((!g739) & (!g740) & (g741) & (g742) & (g147) & (g148)) + ((!g739) & (g740) & (!g741) & (!g742) & (g147) & (!g148)) + ((!g739) & (g740) & (!g741) & (g742) & (g147) & (!g148)) + ((!g739) & (g740) & (!g741) & (g742) & (g147) & (g148)) + ((!g739) & (g740) & (g741) & (!g742) & (!g147) & (g148)) + ((!g739) & (g740) & (g741) & (!g742) & (g147) & (!g148)) + ((!g739) & (g740) & (g741) & (g742) & (!g147) & (g148)) + ((!g739) & (g740) & (g741) & (g742) & (g147) & (!g148)) + ((!g739) & (g740) & (g741) & (g742) & (g147) & (g148)) + ((g739) & (!g740) & (!g741) & (!g742) & (!g147) & (!g148)) + ((g739) & (!g740) & (!g741) & (g742) & (!g147) & (!g148)) + ((g739) & (!g740) & (!g741) & (g742) & (g147) & (g148)) + ((g739) & (!g740) & (g741) & (!g742) & (!g147) & (!g148)) + ((g739) & (!g740) & (g741) & (!g742) & (!g147) & (g148)) + ((g739) & (!g740) & (g741) & (g742) & (!g147) & (!g148)) + ((g739) & (!g740) & (g741) & (g742) & (!g147) & (g148)) + ((g739) & (!g740) & (g741) & (g742) & (g147) & (g148)) + ((g739) & (g740) & (!g741) & (!g742) & (!g147) & (!g148)) + ((g739) & (g740) & (!g741) & (!g742) & (g147) & (!g148)) + ((g739) & (g740) & (!g741) & (g742) & (!g147) & (!g148)) + ((g739) & (g740) & (!g741) & (g742) & (g147) & (!g148)) + ((g739) & (g740) & (!g741) & (g742) & (g147) & (g148)) + ((g739) & (g740) & (g741) & (!g742) & (!g147) & (!g148)) + ((g739) & (g740) & (g741) & (!g742) & (!g147) & (g148)) + ((g739) & (g740) & (g741) & (!g742) & (g147) & (!g148)) + ((g739) & (g740) & (g741) & (g742) & (!g147) & (!g148)) + ((g739) & (g740) & (g741) & (g742) & (!g147) & (g148)) + ((g739) & (g740) & (g741) & (g742) & (g147) & (!g148)) + ((g739) & (g740) & (g741) & (g742) & (g147) & (g148)));
	assign g4419 = (((!g2158) & (!g2495) & (!sk[42]) & (g744)) + ((!g2158) & (!g2495) & (sk[42]) & (g744)) + ((!g2158) & (g2495) & (!sk[42]) & (!g744)) + ((!g2158) & (g2495) & (!sk[42]) & (g744)) + ((!g2158) & (g2495) & (sk[42]) & (g744)) + ((g2158) & (!g2495) & (!sk[42]) & (g744)) + ((g2158) & (g2495) & (!sk[42]) & (!g744)) + ((g2158) & (g2495) & (!sk[42]) & (g744)) + ((g2158) & (g2495) & (sk[42]) & (!g744)) + ((g2158) & (g2495) & (sk[42]) & (g744)));
	assign g4420 = (((!sk[43]) & (!g2159) & (!g2495) & (g745)) + ((!sk[43]) & (!g2159) & (g2495) & (!g745)) + ((!sk[43]) & (!g2159) & (g2495) & (g745)) + ((!sk[43]) & (g2159) & (!g2495) & (g745)) + ((!sk[43]) & (g2159) & (g2495) & (!g745)) + ((!sk[43]) & (g2159) & (g2495) & (g745)) + ((sk[43]) & (!g2159) & (!g2495) & (g745)) + ((sk[43]) & (!g2159) & (g2495) & (g745)) + ((sk[43]) & (g2159) & (g2495) & (!g745)) + ((sk[43]) & (g2159) & (g2495) & (g745)));
	assign g4421 = (((!g2160) & (!g2495) & (!sk[44]) & (g746)) + ((!g2160) & (!g2495) & (sk[44]) & (g746)) + ((!g2160) & (g2495) & (!sk[44]) & (!g746)) + ((!g2160) & (g2495) & (!sk[44]) & (g746)) + ((!g2160) & (g2495) & (sk[44]) & (g746)) + ((g2160) & (!g2495) & (!sk[44]) & (g746)) + ((g2160) & (g2495) & (!sk[44]) & (!g746)) + ((g2160) & (g2495) & (!sk[44]) & (g746)) + ((g2160) & (g2495) & (sk[44]) & (!g746)) + ((g2160) & (g2495) & (sk[44]) & (g746)));
	assign g4422 = (((!sk[45]) & (!g2161) & (!g2495) & (g747)) + ((!sk[45]) & (!g2161) & (g2495) & (!g747)) + ((!sk[45]) & (!g2161) & (g2495) & (g747)) + ((!sk[45]) & (g2161) & (!g2495) & (g747)) + ((!sk[45]) & (g2161) & (g2495) & (!g747)) + ((!sk[45]) & (g2161) & (g2495) & (g747)) + ((sk[45]) & (!g2161) & (!g2495) & (g747)) + ((sk[45]) & (!g2161) & (g2495) & (g747)) + ((sk[45]) & (g2161) & (g2495) & (!g747)) + ((sk[45]) & (g2161) & (g2495) & (g747)));
	assign g748 = (((!g744) & (!g745) & (!g746) & (g747) & (g147) & (g148)) + ((!g744) & (!g745) & (g746) & (!g747) & (!g147) & (g148)) + ((!g744) & (!g745) & (g746) & (g747) & (!g147) & (g148)) + ((!g744) & (!g745) & (g746) & (g747) & (g147) & (g148)) + ((!g744) & (g745) & (!g746) & (!g747) & (g147) & (!g148)) + ((!g744) & (g745) & (!g746) & (g747) & (g147) & (!g148)) + ((!g744) & (g745) & (!g746) & (g747) & (g147) & (g148)) + ((!g744) & (g745) & (g746) & (!g747) & (!g147) & (g148)) + ((!g744) & (g745) & (g746) & (!g747) & (g147) & (!g148)) + ((!g744) & (g745) & (g746) & (g747) & (!g147) & (g148)) + ((!g744) & (g745) & (g746) & (g747) & (g147) & (!g148)) + ((!g744) & (g745) & (g746) & (g747) & (g147) & (g148)) + ((g744) & (!g745) & (!g746) & (!g747) & (!g147) & (!g148)) + ((g744) & (!g745) & (!g746) & (g747) & (!g147) & (!g148)) + ((g744) & (!g745) & (!g746) & (g747) & (g147) & (g148)) + ((g744) & (!g745) & (g746) & (!g747) & (!g147) & (!g148)) + ((g744) & (!g745) & (g746) & (!g747) & (!g147) & (g148)) + ((g744) & (!g745) & (g746) & (g747) & (!g147) & (!g148)) + ((g744) & (!g745) & (g746) & (g747) & (!g147) & (g148)) + ((g744) & (!g745) & (g746) & (g747) & (g147) & (g148)) + ((g744) & (g745) & (!g746) & (!g747) & (!g147) & (!g148)) + ((g744) & (g745) & (!g746) & (!g747) & (g147) & (!g148)) + ((g744) & (g745) & (!g746) & (g747) & (!g147) & (!g148)) + ((g744) & (g745) & (!g746) & (g747) & (g147) & (!g148)) + ((g744) & (g745) & (!g746) & (g747) & (g147) & (g148)) + ((g744) & (g745) & (g746) & (!g747) & (!g147) & (!g148)) + ((g744) & (g745) & (g746) & (!g747) & (!g147) & (g148)) + ((g744) & (g745) & (g746) & (!g747) & (g147) & (!g148)) + ((g744) & (g745) & (g746) & (g747) & (!g147) & (!g148)) + ((g744) & (g745) & (g746) & (g747) & (!g147) & (g148)) + ((g744) & (g745) & (g746) & (g747) & (g147) & (!g148)) + ((g744) & (g745) & (g746) & (g747) & (g147) & (g148)));
	assign g749 = (((!g733) & (!g738) & (!g743) & (g748) & (g165) & (g166)) + ((!g733) & (!g738) & (g743) & (!g748) & (!g165) & (g166)) + ((!g733) & (!g738) & (g743) & (g748) & (!g165) & (g166)) + ((!g733) & (!g738) & (g743) & (g748) & (g165) & (g166)) + ((!g733) & (g738) & (!g743) & (!g748) & (g165) & (!g166)) + ((!g733) & (g738) & (!g743) & (g748) & (g165) & (!g166)) + ((!g733) & (g738) & (!g743) & (g748) & (g165) & (g166)) + ((!g733) & (g738) & (g743) & (!g748) & (!g165) & (g166)) + ((!g733) & (g738) & (g743) & (!g748) & (g165) & (!g166)) + ((!g733) & (g738) & (g743) & (g748) & (!g165) & (g166)) + ((!g733) & (g738) & (g743) & (g748) & (g165) & (!g166)) + ((!g733) & (g738) & (g743) & (g748) & (g165) & (g166)) + ((g733) & (!g738) & (!g743) & (!g748) & (!g165) & (!g166)) + ((g733) & (!g738) & (!g743) & (g748) & (!g165) & (!g166)) + ((g733) & (!g738) & (!g743) & (g748) & (g165) & (g166)) + ((g733) & (!g738) & (g743) & (!g748) & (!g165) & (!g166)) + ((g733) & (!g738) & (g743) & (!g748) & (!g165) & (g166)) + ((g733) & (!g738) & (g743) & (g748) & (!g165) & (!g166)) + ((g733) & (!g738) & (g743) & (g748) & (!g165) & (g166)) + ((g733) & (!g738) & (g743) & (g748) & (g165) & (g166)) + ((g733) & (g738) & (!g743) & (!g748) & (!g165) & (!g166)) + ((g733) & (g738) & (!g743) & (!g748) & (g165) & (!g166)) + ((g733) & (g738) & (!g743) & (g748) & (!g165) & (!g166)) + ((g733) & (g738) & (!g743) & (g748) & (g165) & (!g166)) + ((g733) & (g738) & (!g743) & (g748) & (g165) & (g166)) + ((g733) & (g738) & (g743) & (!g748) & (!g165) & (!g166)) + ((g733) & (g738) & (g743) & (!g748) & (!g165) & (g166)) + ((g733) & (g738) & (g743) & (!g748) & (g165) & (!g166)) + ((g733) & (g738) & (g743) & (g748) & (!g165) & (!g166)) + ((g733) & (g738) & (g743) & (g748) & (!g165) & (g166)) + ((g733) & (g738) & (g743) & (g748) & (g165) & (!g166)) + ((g733) & (g738) & (g743) & (g748) & (g165) & (g166)));
	assign g4423 = (((!g2173) & (!g2495) & (!sk[48]) & (g750)) + ((!g2173) & (!g2495) & (sk[48]) & (g750)) + ((!g2173) & (g2495) & (!sk[48]) & (!g750)) + ((!g2173) & (g2495) & (!sk[48]) & (g750)) + ((!g2173) & (g2495) & (sk[48]) & (g750)) + ((g2173) & (!g2495) & (!sk[48]) & (g750)) + ((g2173) & (g2495) & (!sk[48]) & (!g750)) + ((g2173) & (g2495) & (!sk[48]) & (g750)) + ((g2173) & (g2495) & (sk[48]) & (!g750)) + ((g2173) & (g2495) & (sk[48]) & (g750)));
	assign g4424 = (((!g2174) & (!sk[49]) & (!g2495) & (g751)) + ((!g2174) & (!sk[49]) & (g2495) & (!g751)) + ((!g2174) & (!sk[49]) & (g2495) & (g751)) + ((!g2174) & (sk[49]) & (!g2495) & (g751)) + ((!g2174) & (sk[49]) & (g2495) & (g751)) + ((g2174) & (!sk[49]) & (!g2495) & (g751)) + ((g2174) & (!sk[49]) & (g2495) & (!g751)) + ((g2174) & (!sk[49]) & (g2495) & (g751)) + ((g2174) & (sk[49]) & (g2495) & (!g751)) + ((g2174) & (sk[49]) & (g2495) & (g751)));
	assign g4425 = (((!g2175) & (!g2495) & (!sk[50]) & (g752)) + ((!g2175) & (!g2495) & (sk[50]) & (g752)) + ((!g2175) & (g2495) & (!sk[50]) & (!g752)) + ((!g2175) & (g2495) & (!sk[50]) & (g752)) + ((!g2175) & (g2495) & (sk[50]) & (g752)) + ((g2175) & (!g2495) & (!sk[50]) & (g752)) + ((g2175) & (g2495) & (!sk[50]) & (!g752)) + ((g2175) & (g2495) & (!sk[50]) & (g752)) + ((g2175) & (g2495) & (sk[50]) & (!g752)) + ((g2175) & (g2495) & (sk[50]) & (g752)));
	assign g4426 = (((!sk[51]) & (!g2176) & (!g2495) & (g753)) + ((!sk[51]) & (!g2176) & (g2495) & (!g753)) + ((!sk[51]) & (!g2176) & (g2495) & (g753)) + ((!sk[51]) & (g2176) & (!g2495) & (g753)) + ((!sk[51]) & (g2176) & (g2495) & (!g753)) + ((!sk[51]) & (g2176) & (g2495) & (g753)) + ((sk[51]) & (!g2176) & (!g2495) & (g753)) + ((sk[51]) & (!g2176) & (g2495) & (g753)) + ((sk[51]) & (g2176) & (g2495) & (!g753)) + ((sk[51]) & (g2176) & (g2495) & (g753)));
	assign g754 = (((!g750) & (!g751) & (!g752) & (g753) & (g165) & (g166)) + ((!g750) & (!g751) & (g752) & (!g753) & (!g165) & (g166)) + ((!g750) & (!g751) & (g752) & (g753) & (!g165) & (g166)) + ((!g750) & (!g751) & (g752) & (g753) & (g165) & (g166)) + ((!g750) & (g751) & (!g752) & (!g753) & (g165) & (!g166)) + ((!g750) & (g751) & (!g752) & (g753) & (g165) & (!g166)) + ((!g750) & (g751) & (!g752) & (g753) & (g165) & (g166)) + ((!g750) & (g751) & (g752) & (!g753) & (!g165) & (g166)) + ((!g750) & (g751) & (g752) & (!g753) & (g165) & (!g166)) + ((!g750) & (g751) & (g752) & (g753) & (!g165) & (g166)) + ((!g750) & (g751) & (g752) & (g753) & (g165) & (!g166)) + ((!g750) & (g751) & (g752) & (g753) & (g165) & (g166)) + ((g750) & (!g751) & (!g752) & (!g753) & (!g165) & (!g166)) + ((g750) & (!g751) & (!g752) & (g753) & (!g165) & (!g166)) + ((g750) & (!g751) & (!g752) & (g753) & (g165) & (g166)) + ((g750) & (!g751) & (g752) & (!g753) & (!g165) & (!g166)) + ((g750) & (!g751) & (g752) & (!g753) & (!g165) & (g166)) + ((g750) & (!g751) & (g752) & (g753) & (!g165) & (!g166)) + ((g750) & (!g751) & (g752) & (g753) & (!g165) & (g166)) + ((g750) & (!g751) & (g752) & (g753) & (g165) & (g166)) + ((g750) & (g751) & (!g752) & (!g753) & (!g165) & (!g166)) + ((g750) & (g751) & (!g752) & (!g753) & (g165) & (!g166)) + ((g750) & (g751) & (!g752) & (g753) & (!g165) & (!g166)) + ((g750) & (g751) & (!g752) & (g753) & (g165) & (!g166)) + ((g750) & (g751) & (!g752) & (g753) & (g165) & (g166)) + ((g750) & (g751) & (g752) & (!g753) & (!g165) & (!g166)) + ((g750) & (g751) & (g752) & (!g753) & (!g165) & (g166)) + ((g750) & (g751) & (g752) & (!g753) & (g165) & (!g166)) + ((g750) & (g751) & (g752) & (g753) & (!g165) & (!g166)) + ((g750) & (g751) & (g752) & (g753) & (!g165) & (g166)) + ((g750) & (g751) & (g752) & (g753) & (g165) & (!g166)) + ((g750) & (g751) & (g752) & (g753) & (g165) & (g166)));
	assign g4427 = (((!sk[53]) & (!g2177) & (!g2495) & (g755)) + ((!sk[53]) & (!g2177) & (g2495) & (!g755)) + ((!sk[53]) & (!g2177) & (g2495) & (g755)) + ((!sk[53]) & (g2177) & (!g2495) & (g755)) + ((!sk[53]) & (g2177) & (g2495) & (!g755)) + ((!sk[53]) & (g2177) & (g2495) & (g755)) + ((sk[53]) & (!g2177) & (!g2495) & (g755)) + ((sk[53]) & (!g2177) & (g2495) & (g755)) + ((sk[53]) & (g2177) & (g2495) & (!g755)) + ((sk[53]) & (g2177) & (g2495) & (g755)));
	assign g4428 = (((!g2178) & (!g2495) & (!sk[54]) & (g756)) + ((!g2178) & (!g2495) & (sk[54]) & (g756)) + ((!g2178) & (g2495) & (!sk[54]) & (!g756)) + ((!g2178) & (g2495) & (!sk[54]) & (g756)) + ((!g2178) & (g2495) & (sk[54]) & (g756)) + ((g2178) & (!g2495) & (!sk[54]) & (g756)) + ((g2178) & (g2495) & (!sk[54]) & (!g756)) + ((g2178) & (g2495) & (!sk[54]) & (g756)) + ((g2178) & (g2495) & (sk[54]) & (!g756)) + ((g2178) & (g2495) & (sk[54]) & (g756)));
	assign g4429 = (((!g2179) & (!sk[55]) & (!g2495) & (g757)) + ((!g2179) & (!sk[55]) & (g2495) & (!g757)) + ((!g2179) & (!sk[55]) & (g2495) & (g757)) + ((!g2179) & (sk[55]) & (!g2495) & (g757)) + ((!g2179) & (sk[55]) & (g2495) & (g757)) + ((g2179) & (!sk[55]) & (!g2495) & (g757)) + ((g2179) & (!sk[55]) & (g2495) & (!g757)) + ((g2179) & (!sk[55]) & (g2495) & (g757)) + ((g2179) & (sk[55]) & (g2495) & (!g757)) + ((g2179) & (sk[55]) & (g2495) & (g757)));
	assign g758 = (((!g165) & (!g166) & (!g755) & (g756) & (!sk[56]) & (!g757)) + ((!g165) & (!g166) & (!g755) & (g756) & (!sk[56]) & (g757)) + ((!g165) & (!g166) & (g755) & (!g756) & (!sk[56]) & (!g757)) + ((!g165) & (!g166) & (g755) & (!g756) & (!sk[56]) & (g757)) + ((!g165) & (!g166) & (g755) & (g756) & (!sk[56]) & (!g757)) + ((!g165) & (!g166) & (g755) & (g756) & (!sk[56]) & (g757)) + ((!g165) & (g166) & (!g755) & (!g756) & (!sk[56]) & (!g757)) + ((!g165) & (g166) & (!g755) & (!g756) & (!sk[56]) & (g757)) + ((!g165) & (g166) & (!g755) & (!g756) & (sk[56]) & (g757)) + ((!g165) & (g166) & (!g755) & (g756) & (!sk[56]) & (!g757)) + ((!g165) & (g166) & (!g755) & (g756) & (!sk[56]) & (g757)) + ((!g165) & (g166) & (!g755) & (g756) & (sk[56]) & (g757)) + ((!g165) & (g166) & (g755) & (!g756) & (!sk[56]) & (!g757)) + ((!g165) & (g166) & (g755) & (!g756) & (!sk[56]) & (g757)) + ((!g165) & (g166) & (g755) & (!g756) & (sk[56]) & (g757)) + ((!g165) & (g166) & (g755) & (g756) & (!sk[56]) & (!g757)) + ((!g165) & (g166) & (g755) & (g756) & (!sk[56]) & (g757)) + ((!g165) & (g166) & (g755) & (g756) & (sk[56]) & (g757)) + ((g165) & (!g166) & (!g755) & (g756) & (!sk[56]) & (!g757)) + ((g165) & (!g166) & (!g755) & (g756) & (!sk[56]) & (g757)) + ((g165) & (!g166) & (g755) & (!g756) & (!sk[56]) & (!g757)) + ((g165) & (!g166) & (g755) & (!g756) & (!sk[56]) & (g757)) + ((g165) & (!g166) & (g755) & (!g756) & (sk[56]) & (!g757)) + ((g165) & (!g166) & (g755) & (!g756) & (sk[56]) & (g757)) + ((g165) & (!g166) & (g755) & (g756) & (!sk[56]) & (!g757)) + ((g165) & (!g166) & (g755) & (g756) & (!sk[56]) & (g757)) + ((g165) & (!g166) & (g755) & (g756) & (sk[56]) & (!g757)) + ((g165) & (!g166) & (g755) & (g756) & (sk[56]) & (g757)) + ((g165) & (g166) & (!g755) & (!g756) & (!sk[56]) & (!g757)) + ((g165) & (g166) & (!g755) & (!g756) & (!sk[56]) & (g757)) + ((g165) & (g166) & (!g755) & (g756) & (!sk[56]) & (!g757)) + ((g165) & (g166) & (!g755) & (g756) & (!sk[56]) & (g757)) + ((g165) & (g166) & (!g755) & (g756) & (sk[56]) & (!g757)) + ((g165) & (g166) & (!g755) & (g756) & (sk[56]) & (g757)) + ((g165) & (g166) & (g755) & (!g756) & (!sk[56]) & (!g757)) + ((g165) & (g166) & (g755) & (!g756) & (!sk[56]) & (g757)) + ((g165) & (g166) & (g755) & (g756) & (!sk[56]) & (!g757)) + ((g165) & (g166) & (g755) & (g756) & (!sk[56]) & (g757)) + ((g165) & (g166) & (g755) & (g756) & (sk[56]) & (!g757)) + ((g165) & (g166) & (g755) & (g756) & (sk[56]) & (g757)));
	assign g4430 = (((!g2162) & (!g2495) & (!sk[57]) & (g759)) + ((!g2162) & (!g2495) & (sk[57]) & (g759)) + ((!g2162) & (g2495) & (!sk[57]) & (!g759)) + ((!g2162) & (g2495) & (!sk[57]) & (g759)) + ((!g2162) & (g2495) & (sk[57]) & (g759)) + ((g2162) & (!g2495) & (!sk[57]) & (g759)) + ((g2162) & (g2495) & (!sk[57]) & (!g759)) + ((g2162) & (g2495) & (!sk[57]) & (g759)) + ((g2162) & (g2495) & (sk[57]) & (!g759)) + ((g2162) & (g2495) & (sk[57]) & (g759)));
	assign g4431 = (((!g2164) & (!g2495) & (!sk[58]) & (g760)) + ((!g2164) & (!g2495) & (sk[58]) & (g760)) + ((!g2164) & (g2495) & (!sk[58]) & (!g760)) + ((!g2164) & (g2495) & (!sk[58]) & (g760)) + ((!g2164) & (g2495) & (sk[58]) & (g760)) + ((g2164) & (!g2495) & (!sk[58]) & (g760)) + ((g2164) & (g2495) & (!sk[58]) & (!g760)) + ((g2164) & (g2495) & (!sk[58]) & (g760)) + ((g2164) & (g2495) & (sk[58]) & (!g760)) + ((g2164) & (g2495) & (sk[58]) & (g760)));
	assign g4432 = (((!sk[59]) & (!g2166) & (!g2495) & (g761)) + ((!sk[59]) & (!g2166) & (g2495) & (!g761)) + ((!sk[59]) & (!g2166) & (g2495) & (g761)) + ((!sk[59]) & (g2166) & (!g2495) & (g761)) + ((!sk[59]) & (g2166) & (g2495) & (!g761)) + ((!sk[59]) & (g2166) & (g2495) & (g761)) + ((sk[59]) & (!g2166) & (!g2495) & (g761)) + ((sk[59]) & (!g2166) & (g2495) & (g761)) + ((sk[59]) & (g2166) & (g2495) & (!g761)) + ((sk[59]) & (g2166) & (g2495) & (g761)));
	assign g4433 = (((!g2168) & (!g2495) & (!sk[60]) & (g762)) + ((!g2168) & (!g2495) & (sk[60]) & (g762)) + ((!g2168) & (g2495) & (!sk[60]) & (!g762)) + ((!g2168) & (g2495) & (!sk[60]) & (g762)) + ((!g2168) & (g2495) & (sk[60]) & (g762)) + ((g2168) & (!g2495) & (!sk[60]) & (g762)) + ((g2168) & (g2495) & (!sk[60]) & (!g762)) + ((g2168) & (g2495) & (!sk[60]) & (g762)) + ((g2168) & (g2495) & (sk[60]) & (!g762)) + ((g2168) & (g2495) & (sk[60]) & (g762)));
	assign g763 = (((!g759) & (!g760) & (!g761) & (g762) & (g165) & (g166)) + ((!g759) & (!g760) & (g761) & (!g762) & (!g165) & (g166)) + ((!g759) & (!g760) & (g761) & (g762) & (!g165) & (g166)) + ((!g759) & (!g760) & (g761) & (g762) & (g165) & (g166)) + ((!g759) & (g760) & (!g761) & (!g762) & (g165) & (!g166)) + ((!g759) & (g760) & (!g761) & (g762) & (g165) & (!g166)) + ((!g759) & (g760) & (!g761) & (g762) & (g165) & (g166)) + ((!g759) & (g760) & (g761) & (!g762) & (!g165) & (g166)) + ((!g759) & (g760) & (g761) & (!g762) & (g165) & (!g166)) + ((!g759) & (g760) & (g761) & (g762) & (!g165) & (g166)) + ((!g759) & (g760) & (g761) & (g762) & (g165) & (!g166)) + ((!g759) & (g760) & (g761) & (g762) & (g165) & (g166)) + ((g759) & (!g760) & (!g761) & (!g762) & (!g165) & (!g166)) + ((g759) & (!g760) & (!g761) & (g762) & (!g165) & (!g166)) + ((g759) & (!g760) & (!g761) & (g762) & (g165) & (g166)) + ((g759) & (!g760) & (g761) & (!g762) & (!g165) & (!g166)) + ((g759) & (!g760) & (g761) & (!g762) & (!g165) & (g166)) + ((g759) & (!g760) & (g761) & (g762) & (!g165) & (!g166)) + ((g759) & (!g760) & (g761) & (g762) & (!g165) & (g166)) + ((g759) & (!g760) & (g761) & (g762) & (g165) & (g166)) + ((g759) & (g760) & (!g761) & (!g762) & (!g165) & (!g166)) + ((g759) & (g760) & (!g761) & (!g762) & (g165) & (!g166)) + ((g759) & (g760) & (!g761) & (g762) & (!g165) & (!g166)) + ((g759) & (g760) & (!g761) & (g762) & (g165) & (!g166)) + ((g759) & (g760) & (!g761) & (g762) & (g165) & (g166)) + ((g759) & (g760) & (g761) & (!g762) & (!g165) & (!g166)) + ((g759) & (g760) & (g761) & (!g762) & (!g165) & (g166)) + ((g759) & (g760) & (g761) & (!g762) & (g165) & (!g166)) + ((g759) & (g760) & (g761) & (g762) & (!g165) & (!g166)) + ((g759) & (g760) & (g761) & (g762) & (!g165) & (g166)) + ((g759) & (g760) & (g761) & (g762) & (g165) & (!g166)) + ((g759) & (g760) & (g761) & (g762) & (g165) & (g166)));
	assign g4434 = (((!sk[62]) & (!g2169) & (!g2495) & (g764)) + ((!sk[62]) & (!g2169) & (g2495) & (!g764)) + ((!sk[62]) & (!g2169) & (g2495) & (g764)) + ((!sk[62]) & (g2169) & (!g2495) & (g764)) + ((!sk[62]) & (g2169) & (g2495) & (!g764)) + ((!sk[62]) & (g2169) & (g2495) & (g764)) + ((sk[62]) & (!g2169) & (!g2495) & (g764)) + ((sk[62]) & (!g2169) & (g2495) & (g764)) + ((sk[62]) & (g2169) & (g2495) & (!g764)) + ((sk[62]) & (g2169) & (g2495) & (g764)));
	assign g4435 = (((!g2170) & (!sk[63]) & (!g2495) & (g765)) + ((!g2170) & (!sk[63]) & (g2495) & (!g765)) + ((!g2170) & (!sk[63]) & (g2495) & (g765)) + ((!g2170) & (sk[63]) & (!g2495) & (g765)) + ((!g2170) & (sk[63]) & (g2495) & (g765)) + ((g2170) & (!sk[63]) & (!g2495) & (g765)) + ((g2170) & (!sk[63]) & (g2495) & (!g765)) + ((g2170) & (!sk[63]) & (g2495) & (g765)) + ((g2170) & (sk[63]) & (g2495) & (!g765)) + ((g2170) & (sk[63]) & (g2495) & (g765)));
	assign g4436 = (((!sk[64]) & (!g2171) & (!g2495) & (g766)) + ((!sk[64]) & (!g2171) & (g2495) & (!g766)) + ((!sk[64]) & (!g2171) & (g2495) & (g766)) + ((!sk[64]) & (g2171) & (!g2495) & (g766)) + ((!sk[64]) & (g2171) & (g2495) & (!g766)) + ((!sk[64]) & (g2171) & (g2495) & (g766)) + ((sk[64]) & (!g2171) & (!g2495) & (g766)) + ((sk[64]) & (!g2171) & (g2495) & (g766)) + ((sk[64]) & (g2171) & (g2495) & (!g766)) + ((sk[64]) & (g2171) & (g2495) & (g766)));
	assign g4437 = (((!g2172) & (!g2495) & (!sk[65]) & (g767)) + ((!g2172) & (!g2495) & (sk[65]) & (g767)) + ((!g2172) & (g2495) & (!sk[65]) & (!g767)) + ((!g2172) & (g2495) & (!sk[65]) & (g767)) + ((!g2172) & (g2495) & (sk[65]) & (g767)) + ((g2172) & (!g2495) & (!sk[65]) & (g767)) + ((g2172) & (g2495) & (!sk[65]) & (!g767)) + ((g2172) & (g2495) & (!sk[65]) & (g767)) + ((g2172) & (g2495) & (sk[65]) & (!g767)) + ((g2172) & (g2495) & (sk[65]) & (g767)));
	assign g768 = (((!g764) & (!g765) & (!g766) & (g767) & (g165) & (g166)) + ((!g764) & (!g765) & (g766) & (!g767) & (!g165) & (g166)) + ((!g764) & (!g765) & (g766) & (g767) & (!g165) & (g166)) + ((!g764) & (!g765) & (g766) & (g767) & (g165) & (g166)) + ((!g764) & (g765) & (!g766) & (!g767) & (g165) & (!g166)) + ((!g764) & (g765) & (!g766) & (g767) & (g165) & (!g166)) + ((!g764) & (g765) & (!g766) & (g767) & (g165) & (g166)) + ((!g764) & (g765) & (g766) & (!g767) & (!g165) & (g166)) + ((!g764) & (g765) & (g766) & (!g767) & (g165) & (!g166)) + ((!g764) & (g765) & (g766) & (g767) & (!g165) & (g166)) + ((!g764) & (g765) & (g766) & (g767) & (g165) & (!g166)) + ((!g764) & (g765) & (g766) & (g767) & (g165) & (g166)) + ((g764) & (!g765) & (!g766) & (!g767) & (!g165) & (!g166)) + ((g764) & (!g765) & (!g766) & (g767) & (!g165) & (!g166)) + ((g764) & (!g765) & (!g766) & (g767) & (g165) & (g166)) + ((g764) & (!g765) & (g766) & (!g767) & (!g165) & (!g166)) + ((g764) & (!g765) & (g766) & (!g767) & (!g165) & (g166)) + ((g764) & (!g765) & (g766) & (g767) & (!g165) & (!g166)) + ((g764) & (!g765) & (g766) & (g767) & (!g165) & (g166)) + ((g764) & (!g765) & (g766) & (g767) & (g165) & (g166)) + ((g764) & (g765) & (!g766) & (!g767) & (!g165) & (!g166)) + ((g764) & (g765) & (!g766) & (!g767) & (g165) & (!g166)) + ((g764) & (g765) & (!g766) & (g767) & (!g165) & (!g166)) + ((g764) & (g765) & (!g766) & (g767) & (g165) & (!g166)) + ((g764) & (g765) & (!g766) & (g767) & (g165) & (g166)) + ((g764) & (g765) & (g766) & (!g767) & (!g165) & (!g166)) + ((g764) & (g765) & (g766) & (!g767) & (!g165) & (g166)) + ((g764) & (g765) & (g766) & (!g767) & (g165) & (!g166)) + ((g764) & (g765) & (g766) & (g767) & (!g165) & (!g166)) + ((g764) & (g765) & (g766) & (g767) & (!g165) & (g166)) + ((g764) & (g765) & (g766) & (g767) & (g165) & (!g166)) + ((g764) & (g765) & (g766) & (g767) & (g165) & (g166)));
	assign g769 = (((!g147) & (!g148) & (!g754) & (g758) & (!g763) & (!g768)) + ((!g147) & (!g148) & (!g754) & (g758) & (!g763) & (g768)) + ((!g147) & (!g148) & (!g754) & (g758) & (g763) & (!g768)) + ((!g147) & (!g148) & (!g754) & (g758) & (g763) & (g768)) + ((!g147) & (!g148) & (g754) & (g758) & (!g763) & (!g768)) + ((!g147) & (!g148) & (g754) & (g758) & (!g763) & (g768)) + ((!g147) & (!g148) & (g754) & (g758) & (g763) & (!g768)) + ((!g147) & (!g148) & (g754) & (g758) & (g763) & (g768)) + ((!g147) & (g148) & (!g754) & (!g758) & (!g763) & (g768)) + ((!g147) & (g148) & (!g754) & (!g758) & (g763) & (g768)) + ((!g147) & (g148) & (!g754) & (g758) & (!g763) & (g768)) + ((!g147) & (g148) & (!g754) & (g758) & (g763) & (g768)) + ((!g147) & (g148) & (g754) & (!g758) & (!g763) & (g768)) + ((!g147) & (g148) & (g754) & (!g758) & (g763) & (g768)) + ((!g147) & (g148) & (g754) & (g758) & (!g763) & (g768)) + ((!g147) & (g148) & (g754) & (g758) & (g763) & (g768)) + ((g147) & (!g148) & (g754) & (!g758) & (!g763) & (!g768)) + ((g147) & (!g148) & (g754) & (!g758) & (!g763) & (g768)) + ((g147) & (!g148) & (g754) & (!g758) & (g763) & (!g768)) + ((g147) & (!g148) & (g754) & (!g758) & (g763) & (g768)) + ((g147) & (!g148) & (g754) & (g758) & (!g763) & (!g768)) + ((g147) & (!g148) & (g754) & (g758) & (!g763) & (g768)) + ((g147) & (!g148) & (g754) & (g758) & (g763) & (!g768)) + ((g147) & (!g148) & (g754) & (g758) & (g763) & (g768)) + ((g147) & (g148) & (!g754) & (!g758) & (g763) & (!g768)) + ((g147) & (g148) & (!g754) & (!g758) & (g763) & (g768)) + ((g147) & (g148) & (!g754) & (g758) & (g763) & (!g768)) + ((g147) & (g148) & (!g754) & (g758) & (g763) & (g768)) + ((g147) & (g148) & (g754) & (!g758) & (g763) & (!g768)) + ((g147) & (g148) & (g754) & (!g758) & (g763) & (g768)) + ((g147) & (g148) & (g754) & (g758) & (g763) & (!g768)) + ((g147) & (g148) & (g754) & (g758) & (g763) & (g768)));
	assign g770 = (((!g142) & (!g749) & (!sk[68]) & (g769)) + ((!g142) & (!g749) & (sk[68]) & (g769)) + ((!g142) & (g749) & (!sk[68]) & (!g769)) + ((!g142) & (g749) & (!sk[68]) & (g769)) + ((!g142) & (g749) & (sk[68]) & (g769)) + ((g142) & (!g749) & (!sk[68]) & (g769)) + ((g142) & (g749) & (!sk[68]) & (!g769)) + ((g142) & (g749) & (!sk[68]) & (g769)) + ((g142) & (g749) & (sk[68]) & (!g769)) + ((g142) & (g749) & (sk[68]) & (g769)));
	assign g4438 = (((!g2059) & (!g2504) & (!sk[69]) & (g771)) + ((!g2059) & (!g2504) & (sk[69]) & (g771)) + ((!g2059) & (g2504) & (!sk[69]) & (!g771)) + ((!g2059) & (g2504) & (!sk[69]) & (g771)) + ((!g2059) & (g2504) & (sk[69]) & (g771)) + ((g2059) & (!g2504) & (!sk[69]) & (g771)) + ((g2059) & (g2504) & (!sk[69]) & (!g771)) + ((g2059) & (g2504) & (!sk[69]) & (g771)) + ((g2059) & (g2504) & (sk[69]) & (!g771)) + ((g2059) & (g2504) & (sk[69]) & (g771)));
	assign g772 = (((!g723) & (!g672) & (!g674) & (!g675) & (!g680) & (!g727)) + ((!g723) & (!g672) & (!g674) & (!g675) & (!g680) & (g727)) + ((!g723) & (!g672) & (!g674) & (!g675) & (g680) & (!g727)) + ((!g723) & (!g672) & (!g674) & (!g675) & (g680) & (g727)) + ((!g723) & (!g672) & (!g674) & (g675) & (!g680) & (g727)) + ((!g723) & (!g672) & (!g674) & (g675) & (g680) & (!g727)) + ((!g723) & (!g672) & (!g674) & (g675) & (g680) & (g727)) + ((!g723) & (!g672) & (g674) & (!g675) & (!g680) & (g727)) + ((!g723) & (!g672) & (g674) & (!g675) & (g680) & (!g727)) + ((!g723) & (!g672) & (g674) & (!g675) & (g680) & (g727)) + ((!g723) & (!g672) & (g674) & (g675) & (!g680) & (g727)) + ((!g723) & (!g672) & (g674) & (g675) & (g680) & (!g727)) + ((!g723) & (!g672) & (g674) & (g675) & (g680) & (g727)) + ((!g723) & (g672) & (!g674) & (!g675) & (!g680) & (g727)) + ((!g723) & (g672) & (!g674) & (!g675) & (g680) & (!g727)) + ((!g723) & (g672) & (!g674) & (!g675) & (g680) & (g727)) + ((!g723) & (g672) & (!g674) & (g675) & (!g680) & (g727)) + ((!g723) & (g672) & (!g674) & (g675) & (g680) & (g727)) + ((!g723) & (g672) & (g674) & (!g675) & (!g680) & (g727)) + ((!g723) & (g672) & (g674) & (!g675) & (g680) & (g727)) + ((!g723) & (g672) & (g674) & (g675) & (!g680) & (g727)) + ((!g723) & (g672) & (g674) & (g675) & (g680) & (g727)) + ((g723) & (!g672) & (!g674) & (!g675) & (!g680) & (g727)) + ((g723) & (!g672) & (!g674) & (!g675) & (g680) & (g727)) + ((g723) & (!g672) & (!g674) & (g675) & (g680) & (g727)) + ((g723) & (!g672) & (g674) & (!g675) & (g680) & (g727)) + ((g723) & (!g672) & (g674) & (g675) & (g680) & (g727)) + ((g723) & (g672) & (!g674) & (!g675) & (g680) & (g727)));
	assign g4439 = (((!g2064) & (!dmem_dat_ix13x) & (!sk[71]) & (g773)) + ((!g2064) & (!dmem_dat_ix13x) & (sk[71]) & (g773)) + ((!g2064) & (dmem_dat_ix13x) & (!sk[71]) & (!g773)) + ((!g2064) & (dmem_dat_ix13x) & (!sk[71]) & (g773)) + ((!g2064) & (dmem_dat_ix13x) & (sk[71]) & (g773)) + ((g2064) & (!dmem_dat_ix13x) & (!sk[71]) & (g773)) + ((g2064) & (dmem_dat_ix13x) & (!sk[71]) & (!g773)) + ((g2064) & (dmem_dat_ix13x) & (!sk[71]) & (g773)) + ((g2064) & (dmem_dat_ix13x) & (sk[71]) & (!g773)) + ((g2064) & (dmem_dat_ix13x) & (sk[71]) & (g773)));
	assign g774 = (((!sk[72]) & (!g679) & (!g108) & (g773)) + ((!sk[72]) & (!g679) & (g108) & (!g773)) + ((!sk[72]) & (!g679) & (g108) & (g773)) + ((!sk[72]) & (g679) & (!g108) & (g773)) + ((!sk[72]) & (g679) & (g108) & (!g773)) + ((!sk[72]) & (g679) & (g108) & (g773)) + ((sk[72]) & (!g679) & (!g108) & (!g773)) + ((sk[72]) & (!g679) & (!g108) & (g773)) + ((sk[72]) & (g679) & (!g108) & (!g773)) + ((sk[72]) & (g679) & (g108) & (!g773)));
	assign g775 = (((!g126) & (!sk[73]) & (!g770) & (!g771) & (g772) & (!g774)) + ((!g126) & (!sk[73]) & (!g770) & (!g771) & (g772) & (g774)) + ((!g126) & (!sk[73]) & (!g770) & (g771) & (!g772) & (!g774)) + ((!g126) & (!sk[73]) & (!g770) & (g771) & (!g772) & (g774)) + ((!g126) & (!sk[73]) & (!g770) & (g771) & (g772) & (!g774)) + ((!g126) & (!sk[73]) & (!g770) & (g771) & (g772) & (g774)) + ((!g126) & (!sk[73]) & (g770) & (!g771) & (!g772) & (!g774)) + ((!g126) & (!sk[73]) & (g770) & (!g771) & (!g772) & (g774)) + ((!g126) & (!sk[73]) & (g770) & (!g771) & (g772) & (!g774)) + ((!g126) & (!sk[73]) & (g770) & (!g771) & (g772) & (g774)) + ((!g126) & (!sk[73]) & (g770) & (g771) & (!g772) & (!g774)) + ((!g126) & (!sk[73]) & (g770) & (g771) & (!g772) & (g774)) + ((!g126) & (!sk[73]) & (g770) & (g771) & (g772) & (!g774)) + ((!g126) & (!sk[73]) & (g770) & (g771) & (g772) & (g774)) + ((!g126) & (sk[73]) & (!g770) & (g771) & (!g772) & (!g774)) + ((!g126) & (sk[73]) & (!g770) & (g771) & (!g772) & (g774)) + ((!g126) & (sk[73]) & (!g770) & (g771) & (g772) & (!g774)) + ((!g126) & (sk[73]) & (!g770) & (g771) & (g772) & (g774)) + ((!g126) & (sk[73]) & (g770) & (g771) & (!g772) & (!g774)) + ((!g126) & (sk[73]) & (g770) & (g771) & (!g772) & (g774)) + ((!g126) & (sk[73]) & (g770) & (g771) & (g772) & (!g774)) + ((!g126) & (sk[73]) & (g770) & (g771) & (g772) & (g774)) + ((g126) & (!sk[73]) & (!g770) & (!g771) & (g772) & (!g774)) + ((g126) & (!sk[73]) & (!g770) & (!g771) & (g772) & (g774)) + ((g126) & (!sk[73]) & (!g770) & (g771) & (!g772) & (!g774)) + ((g126) & (!sk[73]) & (!g770) & (g771) & (!g772) & (g774)) + ((g126) & (!sk[73]) & (!g770) & (g771) & (g772) & (!g774)) + ((g126) & (!sk[73]) & (!g770) & (g771) & (g772) & (g774)) + ((g126) & (!sk[73]) & (g770) & (!g771) & (!g772) & (!g774)) + ((g126) & (!sk[73]) & (g770) & (!g771) & (!g772) & (g774)) + ((g126) & (!sk[73]) & (g770) & (!g771) & (g772) & (!g774)) + ((g126) & (!sk[73]) & (g770) & (!g771) & (g772) & (g774)) + ((g126) & (!sk[73]) & (g770) & (g771) & (!g772) & (!g774)) + ((g126) & (!sk[73]) & (g770) & (g771) & (!g772) & (g774)) + ((g126) & (!sk[73]) & (g770) & (g771) & (g772) & (!g774)) + ((g126) & (!sk[73]) & (g770) & (g771) & (g772) & (g774)) + ((g126) & (sk[73]) & (!g770) & (!g771) & (!g772) & (g774)) + ((g126) & (sk[73]) & (!g770) & (!g771) & (g772) & (!g774)) + ((g126) & (sk[73]) & (!g770) & (g771) & (!g772) & (g774)) + ((g126) & (sk[73]) & (!g770) & (g771) & (g772) & (!g774)) + ((g126) & (sk[73]) & (g770) & (!g771) & (!g772) & (!g774)) + ((g126) & (sk[73]) & (g770) & (!g771) & (g772) & (g774)) + ((g126) & (sk[73]) & (g770) & (g771) & (!g772) & (!g774)) + ((g126) & (sk[73]) & (g770) & (g771) & (g772) & (g774)));
	assign g4440 = (((!g2140) & (!sk[74]) & (!g2520) & (g776)) + ((!g2140) & (!sk[74]) & (g2520) & (!g776)) + ((!g2140) & (!sk[74]) & (g2520) & (g776)) + ((!g2140) & (sk[74]) & (!g2520) & (g776)) + ((!g2140) & (sk[74]) & (g2520) & (g776)) + ((g2140) & (!sk[74]) & (!g2520) & (g776)) + ((g2140) & (!sk[74]) & (g2520) & (!g776)) + ((g2140) & (!sk[74]) & (g2520) & (g776)) + ((g2140) & (sk[74]) & (g2520) & (!g776)) + ((g2140) & (sk[74]) & (g2520) & (g776)));
	assign g4441 = (((!g2142) & (!sk[75]) & (!g2520) & (g777)) + ((!g2142) & (!sk[75]) & (g2520) & (!g777)) + ((!g2142) & (!sk[75]) & (g2520) & (g777)) + ((!g2142) & (sk[75]) & (!g2520) & (g777)) + ((!g2142) & (sk[75]) & (g2520) & (g777)) + ((g2142) & (!sk[75]) & (!g2520) & (g777)) + ((g2142) & (!sk[75]) & (g2520) & (!g777)) + ((g2142) & (!sk[75]) & (g2520) & (g777)) + ((g2142) & (sk[75]) & (g2520) & (!g777)) + ((g2142) & (sk[75]) & (g2520) & (g777)));
	assign g4442 = (((!g2144) & (!g2520) & (!sk[76]) & (g778)) + ((!g2144) & (!g2520) & (sk[76]) & (g778)) + ((!g2144) & (g2520) & (!sk[76]) & (!g778)) + ((!g2144) & (g2520) & (!sk[76]) & (g778)) + ((!g2144) & (g2520) & (sk[76]) & (g778)) + ((g2144) & (!g2520) & (!sk[76]) & (g778)) + ((g2144) & (g2520) & (!sk[76]) & (!g778)) + ((g2144) & (g2520) & (!sk[76]) & (g778)) + ((g2144) & (g2520) & (sk[76]) & (!g778)) + ((g2144) & (g2520) & (sk[76]) & (g778)));
	assign g4443 = (((!g2145) & (!g2520) & (!sk[77]) & (g779)) + ((!g2145) & (!g2520) & (sk[77]) & (g779)) + ((!g2145) & (g2520) & (!sk[77]) & (!g779)) + ((!g2145) & (g2520) & (!sk[77]) & (g779)) + ((!g2145) & (g2520) & (sk[77]) & (g779)) + ((g2145) & (!g2520) & (!sk[77]) & (g779)) + ((g2145) & (g2520) & (!sk[77]) & (!g779)) + ((g2145) & (g2520) & (!sk[77]) & (g779)) + ((g2145) & (g2520) & (sk[77]) & (!g779)) + ((g2145) & (g2520) & (sk[77]) & (g779)));
	assign g780 = (((!g776) & (!g777) & (!g778) & (g779) & (g147) & (g148)) + ((!g776) & (!g777) & (g778) & (!g779) & (!g147) & (g148)) + ((!g776) & (!g777) & (g778) & (g779) & (!g147) & (g148)) + ((!g776) & (!g777) & (g778) & (g779) & (g147) & (g148)) + ((!g776) & (g777) & (!g778) & (!g779) & (g147) & (!g148)) + ((!g776) & (g777) & (!g778) & (g779) & (g147) & (!g148)) + ((!g776) & (g777) & (!g778) & (g779) & (g147) & (g148)) + ((!g776) & (g777) & (g778) & (!g779) & (!g147) & (g148)) + ((!g776) & (g777) & (g778) & (!g779) & (g147) & (!g148)) + ((!g776) & (g777) & (g778) & (g779) & (!g147) & (g148)) + ((!g776) & (g777) & (g778) & (g779) & (g147) & (!g148)) + ((!g776) & (g777) & (g778) & (g779) & (g147) & (g148)) + ((g776) & (!g777) & (!g778) & (!g779) & (!g147) & (!g148)) + ((g776) & (!g777) & (!g778) & (g779) & (!g147) & (!g148)) + ((g776) & (!g777) & (!g778) & (g779) & (g147) & (g148)) + ((g776) & (!g777) & (g778) & (!g779) & (!g147) & (!g148)) + ((g776) & (!g777) & (g778) & (!g779) & (!g147) & (g148)) + ((g776) & (!g777) & (g778) & (g779) & (!g147) & (!g148)) + ((g776) & (!g777) & (g778) & (g779) & (!g147) & (g148)) + ((g776) & (!g777) & (g778) & (g779) & (g147) & (g148)) + ((g776) & (g777) & (!g778) & (!g779) & (!g147) & (!g148)) + ((g776) & (g777) & (!g778) & (!g779) & (g147) & (!g148)) + ((g776) & (g777) & (!g778) & (g779) & (!g147) & (!g148)) + ((g776) & (g777) & (!g778) & (g779) & (g147) & (!g148)) + ((g776) & (g777) & (!g778) & (g779) & (g147) & (g148)) + ((g776) & (g777) & (g778) & (!g779) & (!g147) & (!g148)) + ((g776) & (g777) & (g778) & (!g779) & (!g147) & (g148)) + ((g776) & (g777) & (g778) & (!g779) & (g147) & (!g148)) + ((g776) & (g777) & (g778) & (g779) & (!g147) & (!g148)) + ((g776) & (g777) & (g778) & (g779) & (!g147) & (g148)) + ((g776) & (g777) & (g778) & (g779) & (g147) & (!g148)) + ((g776) & (g777) & (g778) & (g779) & (g147) & (g148)));
	assign g4444 = (((!sk[79]) & (!g2146) & (!g2520) & (g781)) + ((!sk[79]) & (!g2146) & (g2520) & (!g781)) + ((!sk[79]) & (!g2146) & (g2520) & (g781)) + ((!sk[79]) & (g2146) & (!g2520) & (g781)) + ((!sk[79]) & (g2146) & (g2520) & (!g781)) + ((!sk[79]) & (g2146) & (g2520) & (g781)) + ((sk[79]) & (!g2146) & (!g2520) & (g781)) + ((sk[79]) & (!g2146) & (g2520) & (g781)) + ((sk[79]) & (g2146) & (g2520) & (!g781)) + ((sk[79]) & (g2146) & (g2520) & (g781)));
	assign g4445 = (((!g2148) & (!g2520) & (!sk[80]) & (g782)) + ((!g2148) & (!g2520) & (sk[80]) & (g782)) + ((!g2148) & (g2520) & (!sk[80]) & (!g782)) + ((!g2148) & (g2520) & (!sk[80]) & (g782)) + ((!g2148) & (g2520) & (sk[80]) & (g782)) + ((g2148) & (!g2520) & (!sk[80]) & (g782)) + ((g2148) & (g2520) & (!sk[80]) & (!g782)) + ((g2148) & (g2520) & (!sk[80]) & (g782)) + ((g2148) & (g2520) & (sk[80]) & (!g782)) + ((g2148) & (g2520) & (sk[80]) & (g782)));
	assign g4446 = (((!sk[81]) & (!g2150) & (!g2520) & (g783)) + ((!sk[81]) & (!g2150) & (g2520) & (!g783)) + ((!sk[81]) & (!g2150) & (g2520) & (g783)) + ((!sk[81]) & (g2150) & (!g2520) & (g783)) + ((!sk[81]) & (g2150) & (g2520) & (!g783)) + ((!sk[81]) & (g2150) & (g2520) & (g783)) + ((sk[81]) & (!g2150) & (!g2520) & (g783)) + ((sk[81]) & (!g2150) & (g2520) & (g783)) + ((sk[81]) & (g2150) & (g2520) & (!g783)) + ((sk[81]) & (g2150) & (g2520) & (g783)));
	assign g4447 = (((!g2151) & (!g2520) & (!sk[82]) & (g784)) + ((!g2151) & (!g2520) & (sk[82]) & (g784)) + ((!g2151) & (g2520) & (!sk[82]) & (!g784)) + ((!g2151) & (g2520) & (!sk[82]) & (g784)) + ((!g2151) & (g2520) & (sk[82]) & (g784)) + ((g2151) & (!g2520) & (!sk[82]) & (g784)) + ((g2151) & (g2520) & (!sk[82]) & (!g784)) + ((g2151) & (g2520) & (!sk[82]) & (g784)) + ((g2151) & (g2520) & (sk[82]) & (!g784)) + ((g2151) & (g2520) & (sk[82]) & (g784)));
	assign g785 = (((!g781) & (!g782) & (!g783) & (g784) & (g147) & (g148)) + ((!g781) & (!g782) & (g783) & (!g784) & (!g147) & (g148)) + ((!g781) & (!g782) & (g783) & (g784) & (!g147) & (g148)) + ((!g781) & (!g782) & (g783) & (g784) & (g147) & (g148)) + ((!g781) & (g782) & (!g783) & (!g784) & (g147) & (!g148)) + ((!g781) & (g782) & (!g783) & (g784) & (g147) & (!g148)) + ((!g781) & (g782) & (!g783) & (g784) & (g147) & (g148)) + ((!g781) & (g782) & (g783) & (!g784) & (!g147) & (g148)) + ((!g781) & (g782) & (g783) & (!g784) & (g147) & (!g148)) + ((!g781) & (g782) & (g783) & (g784) & (!g147) & (g148)) + ((!g781) & (g782) & (g783) & (g784) & (g147) & (!g148)) + ((!g781) & (g782) & (g783) & (g784) & (g147) & (g148)) + ((g781) & (!g782) & (!g783) & (!g784) & (!g147) & (!g148)) + ((g781) & (!g782) & (!g783) & (g784) & (!g147) & (!g148)) + ((g781) & (!g782) & (!g783) & (g784) & (g147) & (g148)) + ((g781) & (!g782) & (g783) & (!g784) & (!g147) & (!g148)) + ((g781) & (!g782) & (g783) & (!g784) & (!g147) & (g148)) + ((g781) & (!g782) & (g783) & (g784) & (!g147) & (!g148)) + ((g781) & (!g782) & (g783) & (g784) & (!g147) & (g148)) + ((g781) & (!g782) & (g783) & (g784) & (g147) & (g148)) + ((g781) & (g782) & (!g783) & (!g784) & (!g147) & (!g148)) + ((g781) & (g782) & (!g783) & (!g784) & (g147) & (!g148)) + ((g781) & (g782) & (!g783) & (g784) & (!g147) & (!g148)) + ((g781) & (g782) & (!g783) & (g784) & (g147) & (!g148)) + ((g781) & (g782) & (!g783) & (g784) & (g147) & (g148)) + ((g781) & (g782) & (g783) & (!g784) & (!g147) & (!g148)) + ((g781) & (g782) & (g783) & (!g784) & (!g147) & (g148)) + ((g781) & (g782) & (g783) & (!g784) & (g147) & (!g148)) + ((g781) & (g782) & (g783) & (g784) & (!g147) & (!g148)) + ((g781) & (g782) & (g783) & (g784) & (!g147) & (g148)) + ((g781) & (g782) & (g783) & (g784) & (g147) & (!g148)) + ((g781) & (g782) & (g783) & (g784) & (g147) & (g148)));
	assign g4448 = (((!g2152) & (!sk[84]) & (!g2520) & (g786)) + ((!g2152) & (!sk[84]) & (g2520) & (!g786)) + ((!g2152) & (!sk[84]) & (g2520) & (g786)) + ((!g2152) & (sk[84]) & (!g2520) & (g786)) + ((!g2152) & (sk[84]) & (g2520) & (g786)) + ((g2152) & (!sk[84]) & (!g2520) & (g786)) + ((g2152) & (!sk[84]) & (g2520) & (!g786)) + ((g2152) & (!sk[84]) & (g2520) & (g786)) + ((g2152) & (sk[84]) & (g2520) & (!g786)) + ((g2152) & (sk[84]) & (g2520) & (g786)));
	assign g4449 = (((!sk[85]) & (!g2153) & (!g2520) & (g787)) + ((!sk[85]) & (!g2153) & (g2520) & (!g787)) + ((!sk[85]) & (!g2153) & (g2520) & (g787)) + ((!sk[85]) & (g2153) & (!g2520) & (g787)) + ((!sk[85]) & (g2153) & (g2520) & (!g787)) + ((!sk[85]) & (g2153) & (g2520) & (g787)) + ((sk[85]) & (!g2153) & (!g2520) & (g787)) + ((sk[85]) & (!g2153) & (g2520) & (g787)) + ((sk[85]) & (g2153) & (g2520) & (!g787)) + ((sk[85]) & (g2153) & (g2520) & (g787)));
	assign g4450 = (((!g2155) & (!g2520) & (!sk[86]) & (g788)) + ((!g2155) & (!g2520) & (sk[86]) & (g788)) + ((!g2155) & (g2520) & (!sk[86]) & (!g788)) + ((!g2155) & (g2520) & (!sk[86]) & (g788)) + ((!g2155) & (g2520) & (sk[86]) & (g788)) + ((g2155) & (!g2520) & (!sk[86]) & (g788)) + ((g2155) & (g2520) & (!sk[86]) & (!g788)) + ((g2155) & (g2520) & (!sk[86]) & (g788)) + ((g2155) & (g2520) & (sk[86]) & (!g788)) + ((g2155) & (g2520) & (sk[86]) & (g788)));
	assign g4451 = (((!g2157) & (!sk[87]) & (!g2520) & (g789)) + ((!g2157) & (!sk[87]) & (g2520) & (!g789)) + ((!g2157) & (!sk[87]) & (g2520) & (g789)) + ((!g2157) & (sk[87]) & (!g2520) & (g789)) + ((!g2157) & (sk[87]) & (g2520) & (g789)) + ((g2157) & (!sk[87]) & (!g2520) & (g789)) + ((g2157) & (!sk[87]) & (g2520) & (!g789)) + ((g2157) & (!sk[87]) & (g2520) & (g789)) + ((g2157) & (sk[87]) & (g2520) & (!g789)) + ((g2157) & (sk[87]) & (g2520) & (g789)));
	assign g790 = (((!g786) & (!g787) & (!g788) & (g789) & (g147) & (g148)) + ((!g786) & (!g787) & (g788) & (!g789) & (!g147) & (g148)) + ((!g786) & (!g787) & (g788) & (g789) & (!g147) & (g148)) + ((!g786) & (!g787) & (g788) & (g789) & (g147) & (g148)) + ((!g786) & (g787) & (!g788) & (!g789) & (g147) & (!g148)) + ((!g786) & (g787) & (!g788) & (g789) & (g147) & (!g148)) + ((!g786) & (g787) & (!g788) & (g789) & (g147) & (g148)) + ((!g786) & (g787) & (g788) & (!g789) & (!g147) & (g148)) + ((!g786) & (g787) & (g788) & (!g789) & (g147) & (!g148)) + ((!g786) & (g787) & (g788) & (g789) & (!g147) & (g148)) + ((!g786) & (g787) & (g788) & (g789) & (g147) & (!g148)) + ((!g786) & (g787) & (g788) & (g789) & (g147) & (g148)) + ((g786) & (!g787) & (!g788) & (!g789) & (!g147) & (!g148)) + ((g786) & (!g787) & (!g788) & (g789) & (!g147) & (!g148)) + ((g786) & (!g787) & (!g788) & (g789) & (g147) & (g148)) + ((g786) & (!g787) & (g788) & (!g789) & (!g147) & (!g148)) + ((g786) & (!g787) & (g788) & (!g789) & (!g147) & (g148)) + ((g786) & (!g787) & (g788) & (g789) & (!g147) & (!g148)) + ((g786) & (!g787) & (g788) & (g789) & (!g147) & (g148)) + ((g786) & (!g787) & (g788) & (g789) & (g147) & (g148)) + ((g786) & (g787) & (!g788) & (!g789) & (!g147) & (!g148)) + ((g786) & (g787) & (!g788) & (!g789) & (g147) & (!g148)) + ((g786) & (g787) & (!g788) & (g789) & (!g147) & (!g148)) + ((g786) & (g787) & (!g788) & (g789) & (g147) & (!g148)) + ((g786) & (g787) & (!g788) & (g789) & (g147) & (g148)) + ((g786) & (g787) & (g788) & (!g789) & (!g147) & (!g148)) + ((g786) & (g787) & (g788) & (!g789) & (!g147) & (g148)) + ((g786) & (g787) & (g788) & (!g789) & (g147) & (!g148)) + ((g786) & (g787) & (g788) & (g789) & (!g147) & (!g148)) + ((g786) & (g787) & (g788) & (g789) & (!g147) & (g148)) + ((g786) & (g787) & (g788) & (g789) & (g147) & (!g148)) + ((g786) & (g787) & (g788) & (g789) & (g147) & (g148)));
	assign g4452 = (((!g2158) & (!sk[89]) & (!g2520) & (g791)) + ((!g2158) & (!sk[89]) & (g2520) & (!g791)) + ((!g2158) & (!sk[89]) & (g2520) & (g791)) + ((!g2158) & (sk[89]) & (!g2520) & (g791)) + ((!g2158) & (sk[89]) & (g2520) & (g791)) + ((g2158) & (!sk[89]) & (!g2520) & (g791)) + ((g2158) & (!sk[89]) & (g2520) & (!g791)) + ((g2158) & (!sk[89]) & (g2520) & (g791)) + ((g2158) & (sk[89]) & (g2520) & (!g791)) + ((g2158) & (sk[89]) & (g2520) & (g791)));
	assign g4453 = (((!sk[90]) & (!g2159) & (!g2520) & (g792)) + ((!sk[90]) & (!g2159) & (g2520) & (!g792)) + ((!sk[90]) & (!g2159) & (g2520) & (g792)) + ((!sk[90]) & (g2159) & (!g2520) & (g792)) + ((!sk[90]) & (g2159) & (g2520) & (!g792)) + ((!sk[90]) & (g2159) & (g2520) & (g792)) + ((sk[90]) & (!g2159) & (!g2520) & (g792)) + ((sk[90]) & (!g2159) & (g2520) & (g792)) + ((sk[90]) & (g2159) & (g2520) & (!g792)) + ((sk[90]) & (g2159) & (g2520) & (g792)));
	assign g4454 = (((!sk[91]) & (!g2160) & (!g2520) & (g793)) + ((!sk[91]) & (!g2160) & (g2520) & (!g793)) + ((!sk[91]) & (!g2160) & (g2520) & (g793)) + ((!sk[91]) & (g2160) & (!g2520) & (g793)) + ((!sk[91]) & (g2160) & (g2520) & (!g793)) + ((!sk[91]) & (g2160) & (g2520) & (g793)) + ((sk[91]) & (!g2160) & (!g2520) & (g793)) + ((sk[91]) & (!g2160) & (g2520) & (g793)) + ((sk[91]) & (g2160) & (g2520) & (!g793)) + ((sk[91]) & (g2160) & (g2520) & (g793)));
	assign g4455 = (((!sk[92]) & (!g2161) & (!g2520) & (g794)) + ((!sk[92]) & (!g2161) & (g2520) & (!g794)) + ((!sk[92]) & (!g2161) & (g2520) & (g794)) + ((!sk[92]) & (g2161) & (!g2520) & (g794)) + ((!sk[92]) & (g2161) & (g2520) & (!g794)) + ((!sk[92]) & (g2161) & (g2520) & (g794)) + ((sk[92]) & (!g2161) & (!g2520) & (g794)) + ((sk[92]) & (!g2161) & (g2520) & (g794)) + ((sk[92]) & (g2161) & (g2520) & (!g794)) + ((sk[92]) & (g2161) & (g2520) & (g794)));
	assign g795 = (((!g791) & (!g792) & (!g793) & (g794) & (g147) & (g148)) + ((!g791) & (!g792) & (g793) & (!g794) & (!g147) & (g148)) + ((!g791) & (!g792) & (g793) & (g794) & (!g147) & (g148)) + ((!g791) & (!g792) & (g793) & (g794) & (g147) & (g148)) + ((!g791) & (g792) & (!g793) & (!g794) & (g147) & (!g148)) + ((!g791) & (g792) & (!g793) & (g794) & (g147) & (!g148)) + ((!g791) & (g792) & (!g793) & (g794) & (g147) & (g148)) + ((!g791) & (g792) & (g793) & (!g794) & (!g147) & (g148)) + ((!g791) & (g792) & (g793) & (!g794) & (g147) & (!g148)) + ((!g791) & (g792) & (g793) & (g794) & (!g147) & (g148)) + ((!g791) & (g792) & (g793) & (g794) & (g147) & (!g148)) + ((!g791) & (g792) & (g793) & (g794) & (g147) & (g148)) + ((g791) & (!g792) & (!g793) & (!g794) & (!g147) & (!g148)) + ((g791) & (!g792) & (!g793) & (g794) & (!g147) & (!g148)) + ((g791) & (!g792) & (!g793) & (g794) & (g147) & (g148)) + ((g791) & (!g792) & (g793) & (!g794) & (!g147) & (!g148)) + ((g791) & (!g792) & (g793) & (!g794) & (!g147) & (g148)) + ((g791) & (!g792) & (g793) & (g794) & (!g147) & (!g148)) + ((g791) & (!g792) & (g793) & (g794) & (!g147) & (g148)) + ((g791) & (!g792) & (g793) & (g794) & (g147) & (g148)) + ((g791) & (g792) & (!g793) & (!g794) & (!g147) & (!g148)) + ((g791) & (g792) & (!g793) & (!g794) & (g147) & (!g148)) + ((g791) & (g792) & (!g793) & (g794) & (!g147) & (!g148)) + ((g791) & (g792) & (!g793) & (g794) & (g147) & (!g148)) + ((g791) & (g792) & (!g793) & (g794) & (g147) & (g148)) + ((g791) & (g792) & (g793) & (!g794) & (!g147) & (!g148)) + ((g791) & (g792) & (g793) & (!g794) & (!g147) & (g148)) + ((g791) & (g792) & (g793) & (!g794) & (g147) & (!g148)) + ((g791) & (g792) & (g793) & (g794) & (!g147) & (!g148)) + ((g791) & (g792) & (g793) & (g794) & (!g147) & (g148)) + ((g791) & (g792) & (g793) & (g794) & (g147) & (!g148)) + ((g791) & (g792) & (g793) & (g794) & (g147) & (g148)));
	assign g796 = (((!g780) & (!g785) & (!g790) & (g795) & (g165) & (g166)) + ((!g780) & (!g785) & (g790) & (!g795) & (!g165) & (g166)) + ((!g780) & (!g785) & (g790) & (g795) & (!g165) & (g166)) + ((!g780) & (!g785) & (g790) & (g795) & (g165) & (g166)) + ((!g780) & (g785) & (!g790) & (!g795) & (g165) & (!g166)) + ((!g780) & (g785) & (!g790) & (g795) & (g165) & (!g166)) + ((!g780) & (g785) & (!g790) & (g795) & (g165) & (g166)) + ((!g780) & (g785) & (g790) & (!g795) & (!g165) & (g166)) + ((!g780) & (g785) & (g790) & (!g795) & (g165) & (!g166)) + ((!g780) & (g785) & (g790) & (g795) & (!g165) & (g166)) + ((!g780) & (g785) & (g790) & (g795) & (g165) & (!g166)) + ((!g780) & (g785) & (g790) & (g795) & (g165) & (g166)) + ((g780) & (!g785) & (!g790) & (!g795) & (!g165) & (!g166)) + ((g780) & (!g785) & (!g790) & (g795) & (!g165) & (!g166)) + ((g780) & (!g785) & (!g790) & (g795) & (g165) & (g166)) + ((g780) & (!g785) & (g790) & (!g795) & (!g165) & (!g166)) + ((g780) & (!g785) & (g790) & (!g795) & (!g165) & (g166)) + ((g780) & (!g785) & (g790) & (g795) & (!g165) & (!g166)) + ((g780) & (!g785) & (g790) & (g795) & (!g165) & (g166)) + ((g780) & (!g785) & (g790) & (g795) & (g165) & (g166)) + ((g780) & (g785) & (!g790) & (!g795) & (!g165) & (!g166)) + ((g780) & (g785) & (!g790) & (!g795) & (g165) & (!g166)) + ((g780) & (g785) & (!g790) & (g795) & (!g165) & (!g166)) + ((g780) & (g785) & (!g790) & (g795) & (g165) & (!g166)) + ((g780) & (g785) & (!g790) & (g795) & (g165) & (g166)) + ((g780) & (g785) & (g790) & (!g795) & (!g165) & (!g166)) + ((g780) & (g785) & (g790) & (!g795) & (!g165) & (g166)) + ((g780) & (g785) & (g790) & (!g795) & (g165) & (!g166)) + ((g780) & (g785) & (g790) & (g795) & (!g165) & (!g166)) + ((g780) & (g785) & (g790) & (g795) & (!g165) & (g166)) + ((g780) & (g785) & (g790) & (g795) & (g165) & (!g166)) + ((g780) & (g785) & (g790) & (g795) & (g165) & (g166)));
	assign g4456 = (((!g2173) & (!g2520) & (!sk[95]) & (g797)) + ((!g2173) & (!g2520) & (sk[95]) & (g797)) + ((!g2173) & (g2520) & (!sk[95]) & (!g797)) + ((!g2173) & (g2520) & (!sk[95]) & (g797)) + ((!g2173) & (g2520) & (sk[95]) & (g797)) + ((g2173) & (!g2520) & (!sk[95]) & (g797)) + ((g2173) & (g2520) & (!sk[95]) & (!g797)) + ((g2173) & (g2520) & (!sk[95]) & (g797)) + ((g2173) & (g2520) & (sk[95]) & (!g797)) + ((g2173) & (g2520) & (sk[95]) & (g797)));
	assign g4457 = (((!g2174) & (!g2520) & (!sk[96]) & (g798)) + ((!g2174) & (!g2520) & (sk[96]) & (g798)) + ((!g2174) & (g2520) & (!sk[96]) & (!g798)) + ((!g2174) & (g2520) & (!sk[96]) & (g798)) + ((!g2174) & (g2520) & (sk[96]) & (g798)) + ((g2174) & (!g2520) & (!sk[96]) & (g798)) + ((g2174) & (g2520) & (!sk[96]) & (!g798)) + ((g2174) & (g2520) & (!sk[96]) & (g798)) + ((g2174) & (g2520) & (sk[96]) & (!g798)) + ((g2174) & (g2520) & (sk[96]) & (g798)));
	assign g4458 = (((!sk[97]) & (!g2175) & (!g2520) & (g799)) + ((!sk[97]) & (!g2175) & (g2520) & (!g799)) + ((!sk[97]) & (!g2175) & (g2520) & (g799)) + ((!sk[97]) & (g2175) & (!g2520) & (g799)) + ((!sk[97]) & (g2175) & (g2520) & (!g799)) + ((!sk[97]) & (g2175) & (g2520) & (g799)) + ((sk[97]) & (!g2175) & (!g2520) & (g799)) + ((sk[97]) & (!g2175) & (g2520) & (g799)) + ((sk[97]) & (g2175) & (g2520) & (!g799)) + ((sk[97]) & (g2175) & (g2520) & (g799)));
	assign g4459 = (((!g2176) & (!sk[98]) & (!g2520) & (g800)) + ((!g2176) & (!sk[98]) & (g2520) & (!g800)) + ((!g2176) & (!sk[98]) & (g2520) & (g800)) + ((!g2176) & (sk[98]) & (!g2520) & (g800)) + ((!g2176) & (sk[98]) & (g2520) & (g800)) + ((g2176) & (!sk[98]) & (!g2520) & (g800)) + ((g2176) & (!sk[98]) & (g2520) & (!g800)) + ((g2176) & (!sk[98]) & (g2520) & (g800)) + ((g2176) & (sk[98]) & (g2520) & (!g800)) + ((g2176) & (sk[98]) & (g2520) & (g800)));
	assign g801 = (((!g797) & (!g798) & (!g799) & (g800) & (g165) & (g166)) + ((!g797) & (!g798) & (g799) & (!g800) & (!g165) & (g166)) + ((!g797) & (!g798) & (g799) & (g800) & (!g165) & (g166)) + ((!g797) & (!g798) & (g799) & (g800) & (g165) & (g166)) + ((!g797) & (g798) & (!g799) & (!g800) & (g165) & (!g166)) + ((!g797) & (g798) & (!g799) & (g800) & (g165) & (!g166)) + ((!g797) & (g798) & (!g799) & (g800) & (g165) & (g166)) + ((!g797) & (g798) & (g799) & (!g800) & (!g165) & (g166)) + ((!g797) & (g798) & (g799) & (!g800) & (g165) & (!g166)) + ((!g797) & (g798) & (g799) & (g800) & (!g165) & (g166)) + ((!g797) & (g798) & (g799) & (g800) & (g165) & (!g166)) + ((!g797) & (g798) & (g799) & (g800) & (g165) & (g166)) + ((g797) & (!g798) & (!g799) & (!g800) & (!g165) & (!g166)) + ((g797) & (!g798) & (!g799) & (g800) & (!g165) & (!g166)) + ((g797) & (!g798) & (!g799) & (g800) & (g165) & (g166)) + ((g797) & (!g798) & (g799) & (!g800) & (!g165) & (!g166)) + ((g797) & (!g798) & (g799) & (!g800) & (!g165) & (g166)) + ((g797) & (!g798) & (g799) & (g800) & (!g165) & (!g166)) + ((g797) & (!g798) & (g799) & (g800) & (!g165) & (g166)) + ((g797) & (!g798) & (g799) & (g800) & (g165) & (g166)) + ((g797) & (g798) & (!g799) & (!g800) & (!g165) & (!g166)) + ((g797) & (g798) & (!g799) & (!g800) & (g165) & (!g166)) + ((g797) & (g798) & (!g799) & (g800) & (!g165) & (!g166)) + ((g797) & (g798) & (!g799) & (g800) & (g165) & (!g166)) + ((g797) & (g798) & (!g799) & (g800) & (g165) & (g166)) + ((g797) & (g798) & (g799) & (!g800) & (!g165) & (!g166)) + ((g797) & (g798) & (g799) & (!g800) & (!g165) & (g166)) + ((g797) & (g798) & (g799) & (!g800) & (g165) & (!g166)) + ((g797) & (g798) & (g799) & (g800) & (!g165) & (!g166)) + ((g797) & (g798) & (g799) & (g800) & (!g165) & (g166)) + ((g797) & (g798) & (g799) & (g800) & (g165) & (!g166)) + ((g797) & (g798) & (g799) & (g800) & (g165) & (g166)));
	assign g4460 = (((!sk[100]) & (!g2177) & (!g2520) & (g802)) + ((!sk[100]) & (!g2177) & (g2520) & (!g802)) + ((!sk[100]) & (!g2177) & (g2520) & (g802)) + ((!sk[100]) & (g2177) & (!g2520) & (g802)) + ((!sk[100]) & (g2177) & (g2520) & (!g802)) + ((!sk[100]) & (g2177) & (g2520) & (g802)) + ((sk[100]) & (!g2177) & (!g2520) & (g802)) + ((sk[100]) & (!g2177) & (g2520) & (g802)) + ((sk[100]) & (g2177) & (g2520) & (!g802)) + ((sk[100]) & (g2177) & (g2520) & (g802)));
	assign g4461 = (((!g2178) & (!g2520) & (!sk[101]) & (g803)) + ((!g2178) & (!g2520) & (sk[101]) & (g803)) + ((!g2178) & (g2520) & (!sk[101]) & (!g803)) + ((!g2178) & (g2520) & (!sk[101]) & (g803)) + ((!g2178) & (g2520) & (sk[101]) & (g803)) + ((g2178) & (!g2520) & (!sk[101]) & (g803)) + ((g2178) & (g2520) & (!sk[101]) & (!g803)) + ((g2178) & (g2520) & (!sk[101]) & (g803)) + ((g2178) & (g2520) & (sk[101]) & (!g803)) + ((g2178) & (g2520) & (sk[101]) & (g803)));
	assign g4462 = (((!g2179) & (!sk[102]) & (!g2520) & (g804)) + ((!g2179) & (!sk[102]) & (g2520) & (!g804)) + ((!g2179) & (!sk[102]) & (g2520) & (g804)) + ((!g2179) & (sk[102]) & (!g2520) & (g804)) + ((!g2179) & (sk[102]) & (g2520) & (g804)) + ((g2179) & (!sk[102]) & (!g2520) & (g804)) + ((g2179) & (!sk[102]) & (g2520) & (!g804)) + ((g2179) & (!sk[102]) & (g2520) & (g804)) + ((g2179) & (sk[102]) & (g2520) & (!g804)) + ((g2179) & (sk[102]) & (g2520) & (g804)));
	assign g805 = (((!sk[103]) & (!g165) & (!g166) & (!g802) & (g803) & (!g804)) + ((!sk[103]) & (!g165) & (!g166) & (!g802) & (g803) & (g804)) + ((!sk[103]) & (!g165) & (!g166) & (g802) & (!g803) & (!g804)) + ((!sk[103]) & (!g165) & (!g166) & (g802) & (!g803) & (g804)) + ((!sk[103]) & (!g165) & (!g166) & (g802) & (g803) & (!g804)) + ((!sk[103]) & (!g165) & (!g166) & (g802) & (g803) & (g804)) + ((!sk[103]) & (!g165) & (g166) & (!g802) & (!g803) & (!g804)) + ((!sk[103]) & (!g165) & (g166) & (!g802) & (!g803) & (g804)) + ((!sk[103]) & (!g165) & (g166) & (!g802) & (g803) & (!g804)) + ((!sk[103]) & (!g165) & (g166) & (!g802) & (g803) & (g804)) + ((!sk[103]) & (!g165) & (g166) & (g802) & (!g803) & (!g804)) + ((!sk[103]) & (!g165) & (g166) & (g802) & (!g803) & (g804)) + ((!sk[103]) & (!g165) & (g166) & (g802) & (g803) & (!g804)) + ((!sk[103]) & (!g165) & (g166) & (g802) & (g803) & (g804)) + ((!sk[103]) & (g165) & (!g166) & (!g802) & (g803) & (!g804)) + ((!sk[103]) & (g165) & (!g166) & (!g802) & (g803) & (g804)) + ((!sk[103]) & (g165) & (!g166) & (g802) & (!g803) & (!g804)) + ((!sk[103]) & (g165) & (!g166) & (g802) & (!g803) & (g804)) + ((!sk[103]) & (g165) & (!g166) & (g802) & (g803) & (!g804)) + ((!sk[103]) & (g165) & (!g166) & (g802) & (g803) & (g804)) + ((!sk[103]) & (g165) & (g166) & (!g802) & (!g803) & (!g804)) + ((!sk[103]) & (g165) & (g166) & (!g802) & (!g803) & (g804)) + ((!sk[103]) & (g165) & (g166) & (!g802) & (g803) & (!g804)) + ((!sk[103]) & (g165) & (g166) & (!g802) & (g803) & (g804)) + ((!sk[103]) & (g165) & (g166) & (g802) & (!g803) & (!g804)) + ((!sk[103]) & (g165) & (g166) & (g802) & (!g803) & (g804)) + ((!sk[103]) & (g165) & (g166) & (g802) & (g803) & (!g804)) + ((!sk[103]) & (g165) & (g166) & (g802) & (g803) & (g804)) + ((sk[103]) & (!g165) & (g166) & (!g802) & (!g803) & (g804)) + ((sk[103]) & (!g165) & (g166) & (!g802) & (g803) & (g804)) + ((sk[103]) & (!g165) & (g166) & (g802) & (!g803) & (g804)) + ((sk[103]) & (!g165) & (g166) & (g802) & (g803) & (g804)) + ((sk[103]) & (g165) & (!g166) & (g802) & (!g803) & (!g804)) + ((sk[103]) & (g165) & (!g166) & (g802) & (!g803) & (g804)) + ((sk[103]) & (g165) & (!g166) & (g802) & (g803) & (!g804)) + ((sk[103]) & (g165) & (!g166) & (g802) & (g803) & (g804)) + ((sk[103]) & (g165) & (g166) & (!g802) & (g803) & (!g804)) + ((sk[103]) & (g165) & (g166) & (!g802) & (g803) & (g804)) + ((sk[103]) & (g165) & (g166) & (g802) & (g803) & (!g804)) + ((sk[103]) & (g165) & (g166) & (g802) & (g803) & (g804)));
	assign g4463 = (((!g2162) & (!g2520) & (!sk[104]) & (g806)) + ((!g2162) & (!g2520) & (sk[104]) & (g806)) + ((!g2162) & (g2520) & (!sk[104]) & (!g806)) + ((!g2162) & (g2520) & (!sk[104]) & (g806)) + ((!g2162) & (g2520) & (sk[104]) & (g806)) + ((g2162) & (!g2520) & (!sk[104]) & (g806)) + ((g2162) & (g2520) & (!sk[104]) & (!g806)) + ((g2162) & (g2520) & (!sk[104]) & (g806)) + ((g2162) & (g2520) & (sk[104]) & (!g806)) + ((g2162) & (g2520) & (sk[104]) & (g806)));
	assign g4464 = (((!sk[105]) & (!g2164) & (!g2520) & (g807)) + ((!sk[105]) & (!g2164) & (g2520) & (!g807)) + ((!sk[105]) & (!g2164) & (g2520) & (g807)) + ((!sk[105]) & (g2164) & (!g2520) & (g807)) + ((!sk[105]) & (g2164) & (g2520) & (!g807)) + ((!sk[105]) & (g2164) & (g2520) & (g807)) + ((sk[105]) & (!g2164) & (!g2520) & (g807)) + ((sk[105]) & (!g2164) & (g2520) & (g807)) + ((sk[105]) & (g2164) & (g2520) & (!g807)) + ((sk[105]) & (g2164) & (g2520) & (g807)));
	assign g4465 = (((!sk[106]) & (!g2166) & (!g2520) & (g808)) + ((!sk[106]) & (!g2166) & (g2520) & (!g808)) + ((!sk[106]) & (!g2166) & (g2520) & (g808)) + ((!sk[106]) & (g2166) & (!g2520) & (g808)) + ((!sk[106]) & (g2166) & (g2520) & (!g808)) + ((!sk[106]) & (g2166) & (g2520) & (g808)) + ((sk[106]) & (!g2166) & (!g2520) & (g808)) + ((sk[106]) & (!g2166) & (g2520) & (g808)) + ((sk[106]) & (g2166) & (g2520) & (!g808)) + ((sk[106]) & (g2166) & (g2520) & (g808)));
	assign g4466 = (((!sk[107]) & (!g2168) & (!g2520) & (g809)) + ((!sk[107]) & (!g2168) & (g2520) & (!g809)) + ((!sk[107]) & (!g2168) & (g2520) & (g809)) + ((!sk[107]) & (g2168) & (!g2520) & (g809)) + ((!sk[107]) & (g2168) & (g2520) & (!g809)) + ((!sk[107]) & (g2168) & (g2520) & (g809)) + ((sk[107]) & (!g2168) & (!g2520) & (g809)) + ((sk[107]) & (!g2168) & (g2520) & (g809)) + ((sk[107]) & (g2168) & (g2520) & (!g809)) + ((sk[107]) & (g2168) & (g2520) & (g809)));
	assign g810 = (((!g806) & (!g807) & (!g808) & (g809) & (g165) & (g166)) + ((!g806) & (!g807) & (g808) & (!g809) & (!g165) & (g166)) + ((!g806) & (!g807) & (g808) & (g809) & (!g165) & (g166)) + ((!g806) & (!g807) & (g808) & (g809) & (g165) & (g166)) + ((!g806) & (g807) & (!g808) & (!g809) & (g165) & (!g166)) + ((!g806) & (g807) & (!g808) & (g809) & (g165) & (!g166)) + ((!g806) & (g807) & (!g808) & (g809) & (g165) & (g166)) + ((!g806) & (g807) & (g808) & (!g809) & (!g165) & (g166)) + ((!g806) & (g807) & (g808) & (!g809) & (g165) & (!g166)) + ((!g806) & (g807) & (g808) & (g809) & (!g165) & (g166)) + ((!g806) & (g807) & (g808) & (g809) & (g165) & (!g166)) + ((!g806) & (g807) & (g808) & (g809) & (g165) & (g166)) + ((g806) & (!g807) & (!g808) & (!g809) & (!g165) & (!g166)) + ((g806) & (!g807) & (!g808) & (g809) & (!g165) & (!g166)) + ((g806) & (!g807) & (!g808) & (g809) & (g165) & (g166)) + ((g806) & (!g807) & (g808) & (!g809) & (!g165) & (!g166)) + ((g806) & (!g807) & (g808) & (!g809) & (!g165) & (g166)) + ((g806) & (!g807) & (g808) & (g809) & (!g165) & (!g166)) + ((g806) & (!g807) & (g808) & (g809) & (!g165) & (g166)) + ((g806) & (!g807) & (g808) & (g809) & (g165) & (g166)) + ((g806) & (g807) & (!g808) & (!g809) & (!g165) & (!g166)) + ((g806) & (g807) & (!g808) & (!g809) & (g165) & (!g166)) + ((g806) & (g807) & (!g808) & (g809) & (!g165) & (!g166)) + ((g806) & (g807) & (!g808) & (g809) & (g165) & (!g166)) + ((g806) & (g807) & (!g808) & (g809) & (g165) & (g166)) + ((g806) & (g807) & (g808) & (!g809) & (!g165) & (!g166)) + ((g806) & (g807) & (g808) & (!g809) & (!g165) & (g166)) + ((g806) & (g807) & (g808) & (!g809) & (g165) & (!g166)) + ((g806) & (g807) & (g808) & (g809) & (!g165) & (!g166)) + ((g806) & (g807) & (g808) & (g809) & (!g165) & (g166)) + ((g806) & (g807) & (g808) & (g809) & (g165) & (!g166)) + ((g806) & (g807) & (g808) & (g809) & (g165) & (g166)));
	assign g4467 = (((!g2169) & (!g2520) & (!sk[109]) & (g811)) + ((!g2169) & (!g2520) & (sk[109]) & (g811)) + ((!g2169) & (g2520) & (!sk[109]) & (!g811)) + ((!g2169) & (g2520) & (!sk[109]) & (g811)) + ((!g2169) & (g2520) & (sk[109]) & (g811)) + ((g2169) & (!g2520) & (!sk[109]) & (g811)) + ((g2169) & (g2520) & (!sk[109]) & (!g811)) + ((g2169) & (g2520) & (!sk[109]) & (g811)) + ((g2169) & (g2520) & (sk[109]) & (!g811)) + ((g2169) & (g2520) & (sk[109]) & (g811)));
	assign g4468 = (((!g2170) & (!g2520) & (!sk[110]) & (g812)) + ((!g2170) & (!g2520) & (sk[110]) & (g812)) + ((!g2170) & (g2520) & (!sk[110]) & (!g812)) + ((!g2170) & (g2520) & (!sk[110]) & (g812)) + ((!g2170) & (g2520) & (sk[110]) & (g812)) + ((g2170) & (!g2520) & (!sk[110]) & (g812)) + ((g2170) & (g2520) & (!sk[110]) & (!g812)) + ((g2170) & (g2520) & (!sk[110]) & (g812)) + ((g2170) & (g2520) & (sk[110]) & (!g812)) + ((g2170) & (g2520) & (sk[110]) & (g812)));
	assign g4469 = (((!sk[111]) & (!g2171) & (!g2520) & (g813)) + ((!sk[111]) & (!g2171) & (g2520) & (!g813)) + ((!sk[111]) & (!g2171) & (g2520) & (g813)) + ((!sk[111]) & (g2171) & (!g2520) & (g813)) + ((!sk[111]) & (g2171) & (g2520) & (!g813)) + ((!sk[111]) & (g2171) & (g2520) & (g813)) + ((sk[111]) & (!g2171) & (!g2520) & (g813)) + ((sk[111]) & (!g2171) & (g2520) & (g813)) + ((sk[111]) & (g2171) & (g2520) & (!g813)) + ((sk[111]) & (g2171) & (g2520) & (g813)));
	assign g4470 = (((!sk[112]) & (!g2172) & (!g2520) & (g814)) + ((!sk[112]) & (!g2172) & (g2520) & (!g814)) + ((!sk[112]) & (!g2172) & (g2520) & (g814)) + ((!sk[112]) & (g2172) & (!g2520) & (g814)) + ((!sk[112]) & (g2172) & (g2520) & (!g814)) + ((!sk[112]) & (g2172) & (g2520) & (g814)) + ((sk[112]) & (!g2172) & (!g2520) & (g814)) + ((sk[112]) & (!g2172) & (g2520) & (g814)) + ((sk[112]) & (g2172) & (g2520) & (!g814)) + ((sk[112]) & (g2172) & (g2520) & (g814)));
	assign g815 = (((!g811) & (!g812) & (!g813) & (g814) & (g165) & (g166)) + ((!g811) & (!g812) & (g813) & (!g814) & (!g165) & (g166)) + ((!g811) & (!g812) & (g813) & (g814) & (!g165) & (g166)) + ((!g811) & (!g812) & (g813) & (g814) & (g165) & (g166)) + ((!g811) & (g812) & (!g813) & (!g814) & (g165) & (!g166)) + ((!g811) & (g812) & (!g813) & (g814) & (g165) & (!g166)) + ((!g811) & (g812) & (!g813) & (g814) & (g165) & (g166)) + ((!g811) & (g812) & (g813) & (!g814) & (!g165) & (g166)) + ((!g811) & (g812) & (g813) & (!g814) & (g165) & (!g166)) + ((!g811) & (g812) & (g813) & (g814) & (!g165) & (g166)) + ((!g811) & (g812) & (g813) & (g814) & (g165) & (!g166)) + ((!g811) & (g812) & (g813) & (g814) & (g165) & (g166)) + ((g811) & (!g812) & (!g813) & (!g814) & (!g165) & (!g166)) + ((g811) & (!g812) & (!g813) & (g814) & (!g165) & (!g166)) + ((g811) & (!g812) & (!g813) & (g814) & (g165) & (g166)) + ((g811) & (!g812) & (g813) & (!g814) & (!g165) & (!g166)) + ((g811) & (!g812) & (g813) & (!g814) & (!g165) & (g166)) + ((g811) & (!g812) & (g813) & (g814) & (!g165) & (!g166)) + ((g811) & (!g812) & (g813) & (g814) & (!g165) & (g166)) + ((g811) & (!g812) & (g813) & (g814) & (g165) & (g166)) + ((g811) & (g812) & (!g813) & (!g814) & (!g165) & (!g166)) + ((g811) & (g812) & (!g813) & (!g814) & (g165) & (!g166)) + ((g811) & (g812) & (!g813) & (g814) & (!g165) & (!g166)) + ((g811) & (g812) & (!g813) & (g814) & (g165) & (!g166)) + ((g811) & (g812) & (!g813) & (g814) & (g165) & (g166)) + ((g811) & (g812) & (g813) & (!g814) & (!g165) & (!g166)) + ((g811) & (g812) & (g813) & (!g814) & (!g165) & (g166)) + ((g811) & (g812) & (g813) & (!g814) & (g165) & (!g166)) + ((g811) & (g812) & (g813) & (g814) & (!g165) & (!g166)) + ((g811) & (g812) & (g813) & (g814) & (!g165) & (g166)) + ((g811) & (g812) & (g813) & (g814) & (g165) & (!g166)) + ((g811) & (g812) & (g813) & (g814) & (g165) & (g166)));
	assign g816 = (((!g147) & (!g148) & (!g801) & (g805) & (!g810) & (!g815)) + ((!g147) & (!g148) & (!g801) & (g805) & (!g810) & (g815)) + ((!g147) & (!g148) & (!g801) & (g805) & (g810) & (!g815)) + ((!g147) & (!g148) & (!g801) & (g805) & (g810) & (g815)) + ((!g147) & (!g148) & (g801) & (g805) & (!g810) & (!g815)) + ((!g147) & (!g148) & (g801) & (g805) & (!g810) & (g815)) + ((!g147) & (!g148) & (g801) & (g805) & (g810) & (!g815)) + ((!g147) & (!g148) & (g801) & (g805) & (g810) & (g815)) + ((!g147) & (g148) & (!g801) & (!g805) & (!g810) & (g815)) + ((!g147) & (g148) & (!g801) & (!g805) & (g810) & (g815)) + ((!g147) & (g148) & (!g801) & (g805) & (!g810) & (g815)) + ((!g147) & (g148) & (!g801) & (g805) & (g810) & (g815)) + ((!g147) & (g148) & (g801) & (!g805) & (!g810) & (g815)) + ((!g147) & (g148) & (g801) & (!g805) & (g810) & (g815)) + ((!g147) & (g148) & (g801) & (g805) & (!g810) & (g815)) + ((!g147) & (g148) & (g801) & (g805) & (g810) & (g815)) + ((g147) & (!g148) & (g801) & (!g805) & (!g810) & (!g815)) + ((g147) & (!g148) & (g801) & (!g805) & (!g810) & (g815)) + ((g147) & (!g148) & (g801) & (!g805) & (g810) & (!g815)) + ((g147) & (!g148) & (g801) & (!g805) & (g810) & (g815)) + ((g147) & (!g148) & (g801) & (g805) & (!g810) & (!g815)) + ((g147) & (!g148) & (g801) & (g805) & (!g810) & (g815)) + ((g147) & (!g148) & (g801) & (g805) & (g810) & (!g815)) + ((g147) & (!g148) & (g801) & (g805) & (g810) & (g815)) + ((g147) & (g148) & (!g801) & (!g805) & (g810) & (!g815)) + ((g147) & (g148) & (!g801) & (!g805) & (g810) & (g815)) + ((g147) & (g148) & (!g801) & (g805) & (g810) & (!g815)) + ((g147) & (g148) & (!g801) & (g805) & (g810) & (g815)) + ((g147) & (g148) & (g801) & (!g805) & (g810) & (!g815)) + ((g147) & (g148) & (g801) & (!g805) & (g810) & (g815)) + ((g147) & (g148) & (g801) & (g805) & (g810) & (!g815)) + ((g147) & (g148) & (g801) & (g805) & (g810) & (g815)));
	assign g817 = (((!g142) & (!sk[115]) & (!g796) & (g816)) + ((!g142) & (!sk[115]) & (g796) & (!g816)) + ((!g142) & (!sk[115]) & (g796) & (g816)) + ((!g142) & (sk[115]) & (!g796) & (g816)) + ((!g142) & (sk[115]) & (g796) & (g816)) + ((g142) & (!sk[115]) & (!g796) & (g816)) + ((g142) & (!sk[115]) & (g796) & (!g816)) + ((g142) & (!sk[115]) & (g796) & (g816)) + ((g142) & (sk[115]) & (g796) & (!g816)) + ((g142) & (sk[115]) & (g796) & (g816)));
	assign g4471 = (((!g2059) & (!g2526) & (!sk[116]) & (g818)) + ((!g2059) & (!g2526) & (sk[116]) & (g818)) + ((!g2059) & (g2526) & (!sk[116]) & (!g818)) + ((!g2059) & (g2526) & (!sk[116]) & (g818)) + ((!g2059) & (g2526) & (sk[116]) & (g818)) + ((g2059) & (!g2526) & (!sk[116]) & (g818)) + ((g2059) & (g2526) & (!sk[116]) & (!g818)) + ((g2059) & (g2526) & (!sk[116]) & (g818)) + ((g2059) & (g2526) & (sk[116]) & (!g818)) + ((g2059) & (g2526) & (sk[116]) & (g818)));
	assign g819 = (((!g770) & (!sk[117]) & (!g772) & (g774)) + ((!g770) & (!sk[117]) & (g772) & (!g774)) + ((!g770) & (!sk[117]) & (g772) & (g774)) + ((!g770) & (sk[117]) & (!g772) & (!g774)) + ((g770) & (!sk[117]) & (!g772) & (g774)) + ((g770) & (!sk[117]) & (g772) & (!g774)) + ((g770) & (!sk[117]) & (g772) & (g774)) + ((g770) & (sk[117]) & (!g772) & (!g774)) + ((g770) & (sk[117]) & (!g772) & (g774)) + ((g770) & (sk[117]) & (g772) & (!g774)));
	assign g4472 = (((!sk[118]) & (!g2064) & (!dmem_dat_ix14x) & (g820)) + ((!sk[118]) & (!g2064) & (dmem_dat_ix14x) & (!g820)) + ((!sk[118]) & (!g2064) & (dmem_dat_ix14x) & (g820)) + ((!sk[118]) & (g2064) & (!dmem_dat_ix14x) & (g820)) + ((!sk[118]) & (g2064) & (dmem_dat_ix14x) & (!g820)) + ((!sk[118]) & (g2064) & (dmem_dat_ix14x) & (g820)) + ((sk[118]) & (!g2064) & (!dmem_dat_ix14x) & (g820)) + ((sk[118]) & (!g2064) & (dmem_dat_ix14x) & (g820)) + ((sk[118]) & (g2064) & (dmem_dat_ix14x) & (!g820)) + ((sk[118]) & (g2064) & (dmem_dat_ix14x) & (g820)));
	assign g821 = (((!sk[119]) & (!g679) & (!g110) & (g820)) + ((!sk[119]) & (!g679) & (g110) & (!g820)) + ((!sk[119]) & (!g679) & (g110) & (g820)) + ((!sk[119]) & (g679) & (!g110) & (g820)) + ((!sk[119]) & (g679) & (g110) & (!g820)) + ((!sk[119]) & (g679) & (g110) & (g820)) + ((sk[119]) & (!g679) & (!g110) & (!g820)) + ((sk[119]) & (!g679) & (!g110) & (g820)) + ((sk[119]) & (g679) & (!g110) & (!g820)) + ((sk[119]) & (g679) & (g110) & (!g820)));
	assign g822 = (((!g126) & (!g817) & (!sk[120]) & (!g818) & (g819) & (!g821)) + ((!g126) & (!g817) & (!sk[120]) & (!g818) & (g819) & (g821)) + ((!g126) & (!g817) & (!sk[120]) & (g818) & (!g819) & (!g821)) + ((!g126) & (!g817) & (!sk[120]) & (g818) & (!g819) & (g821)) + ((!g126) & (!g817) & (!sk[120]) & (g818) & (g819) & (!g821)) + ((!g126) & (!g817) & (!sk[120]) & (g818) & (g819) & (g821)) + ((!g126) & (!g817) & (sk[120]) & (g818) & (!g819) & (!g821)) + ((!g126) & (!g817) & (sk[120]) & (g818) & (!g819) & (g821)) + ((!g126) & (!g817) & (sk[120]) & (g818) & (g819) & (!g821)) + ((!g126) & (!g817) & (sk[120]) & (g818) & (g819) & (g821)) + ((!g126) & (g817) & (!sk[120]) & (!g818) & (!g819) & (!g821)) + ((!g126) & (g817) & (!sk[120]) & (!g818) & (!g819) & (g821)) + ((!g126) & (g817) & (!sk[120]) & (!g818) & (g819) & (!g821)) + ((!g126) & (g817) & (!sk[120]) & (!g818) & (g819) & (g821)) + ((!g126) & (g817) & (!sk[120]) & (g818) & (!g819) & (!g821)) + ((!g126) & (g817) & (!sk[120]) & (g818) & (!g819) & (g821)) + ((!g126) & (g817) & (!sk[120]) & (g818) & (g819) & (!g821)) + ((!g126) & (g817) & (!sk[120]) & (g818) & (g819) & (g821)) + ((!g126) & (g817) & (sk[120]) & (g818) & (!g819) & (!g821)) + ((!g126) & (g817) & (sk[120]) & (g818) & (!g819) & (g821)) + ((!g126) & (g817) & (sk[120]) & (g818) & (g819) & (!g821)) + ((!g126) & (g817) & (sk[120]) & (g818) & (g819) & (g821)) + ((g126) & (!g817) & (!sk[120]) & (!g818) & (g819) & (!g821)) + ((g126) & (!g817) & (!sk[120]) & (!g818) & (g819) & (g821)) + ((g126) & (!g817) & (!sk[120]) & (g818) & (!g819) & (!g821)) + ((g126) & (!g817) & (!sk[120]) & (g818) & (!g819) & (g821)) + ((g126) & (!g817) & (!sk[120]) & (g818) & (g819) & (!g821)) + ((g126) & (!g817) & (!sk[120]) & (g818) & (g819) & (g821)) + ((g126) & (!g817) & (sk[120]) & (!g818) & (!g819) & (!g821)) + ((g126) & (!g817) & (sk[120]) & (!g818) & (g819) & (g821)) + ((g126) & (!g817) & (sk[120]) & (g818) & (!g819) & (!g821)) + ((g126) & (!g817) & (sk[120]) & (g818) & (g819) & (g821)) + ((g126) & (g817) & (!sk[120]) & (!g818) & (!g819) & (!g821)) + ((g126) & (g817) & (!sk[120]) & (!g818) & (!g819) & (g821)) + ((g126) & (g817) & (!sk[120]) & (!g818) & (g819) & (!g821)) + ((g126) & (g817) & (!sk[120]) & (!g818) & (g819) & (g821)) + ((g126) & (g817) & (!sk[120]) & (g818) & (!g819) & (!g821)) + ((g126) & (g817) & (!sk[120]) & (g818) & (!g819) & (g821)) + ((g126) & (g817) & (!sk[120]) & (g818) & (g819) & (!g821)) + ((g126) & (g817) & (!sk[120]) & (g818) & (g819) & (g821)) + ((g126) & (g817) & (sk[120]) & (!g818) & (!g819) & (g821)) + ((g126) & (g817) & (sk[120]) & (!g818) & (g819) & (!g821)) + ((g126) & (g817) & (sk[120]) & (g818) & (!g819) & (g821)) + ((g126) & (g817) & (sk[120]) & (g818) & (g819) & (!g821)));
	assign g4473 = (((!g2140) & (!g2542) & (!sk[121]) & (g823)) + ((!g2140) & (!g2542) & (sk[121]) & (g823)) + ((!g2140) & (g2542) & (!sk[121]) & (!g823)) + ((!g2140) & (g2542) & (!sk[121]) & (g823)) + ((!g2140) & (g2542) & (sk[121]) & (g823)) + ((g2140) & (!g2542) & (!sk[121]) & (g823)) + ((g2140) & (g2542) & (!sk[121]) & (!g823)) + ((g2140) & (g2542) & (!sk[121]) & (g823)) + ((g2140) & (g2542) & (sk[121]) & (!g823)) + ((g2140) & (g2542) & (sk[121]) & (g823)));
	assign g4474 = (((!sk[122]) & (!g2142) & (!g2542) & (g824)) + ((!sk[122]) & (!g2142) & (g2542) & (!g824)) + ((!sk[122]) & (!g2142) & (g2542) & (g824)) + ((!sk[122]) & (g2142) & (!g2542) & (g824)) + ((!sk[122]) & (g2142) & (g2542) & (!g824)) + ((!sk[122]) & (g2142) & (g2542) & (g824)) + ((sk[122]) & (!g2142) & (!g2542) & (g824)) + ((sk[122]) & (!g2142) & (g2542) & (g824)) + ((sk[122]) & (g2142) & (g2542) & (!g824)) + ((sk[122]) & (g2142) & (g2542) & (g824)));
	assign g4475 = (((!g2144) & (!sk[123]) & (!g2542) & (g825)) + ((!g2144) & (!sk[123]) & (g2542) & (!g825)) + ((!g2144) & (!sk[123]) & (g2542) & (g825)) + ((!g2144) & (sk[123]) & (!g2542) & (g825)) + ((!g2144) & (sk[123]) & (g2542) & (g825)) + ((g2144) & (!sk[123]) & (!g2542) & (g825)) + ((g2144) & (!sk[123]) & (g2542) & (!g825)) + ((g2144) & (!sk[123]) & (g2542) & (g825)) + ((g2144) & (sk[123]) & (g2542) & (!g825)) + ((g2144) & (sk[123]) & (g2542) & (g825)));
	assign g4476 = (((!sk[124]) & (!g2145) & (!g2542) & (g826)) + ((!sk[124]) & (!g2145) & (g2542) & (!g826)) + ((!sk[124]) & (!g2145) & (g2542) & (g826)) + ((!sk[124]) & (g2145) & (!g2542) & (g826)) + ((!sk[124]) & (g2145) & (g2542) & (!g826)) + ((!sk[124]) & (g2145) & (g2542) & (g826)) + ((sk[124]) & (!g2145) & (!g2542) & (g826)) + ((sk[124]) & (!g2145) & (g2542) & (g826)) + ((sk[124]) & (g2145) & (g2542) & (!g826)) + ((sk[124]) & (g2145) & (g2542) & (g826)));
	assign g827 = (((!g823) & (!g824) & (!g825) & (g826) & (g147) & (g148)) + ((!g823) & (!g824) & (g825) & (!g826) & (!g147) & (g148)) + ((!g823) & (!g824) & (g825) & (g826) & (!g147) & (g148)) + ((!g823) & (!g824) & (g825) & (g826) & (g147) & (g148)) + ((!g823) & (g824) & (!g825) & (!g826) & (g147) & (!g148)) + ((!g823) & (g824) & (!g825) & (g826) & (g147) & (!g148)) + ((!g823) & (g824) & (!g825) & (g826) & (g147) & (g148)) + ((!g823) & (g824) & (g825) & (!g826) & (!g147) & (g148)) + ((!g823) & (g824) & (g825) & (!g826) & (g147) & (!g148)) + ((!g823) & (g824) & (g825) & (g826) & (!g147) & (g148)) + ((!g823) & (g824) & (g825) & (g826) & (g147) & (!g148)) + ((!g823) & (g824) & (g825) & (g826) & (g147) & (g148)) + ((g823) & (!g824) & (!g825) & (!g826) & (!g147) & (!g148)) + ((g823) & (!g824) & (!g825) & (g826) & (!g147) & (!g148)) + ((g823) & (!g824) & (!g825) & (g826) & (g147) & (g148)) + ((g823) & (!g824) & (g825) & (!g826) & (!g147) & (!g148)) + ((g823) & (!g824) & (g825) & (!g826) & (!g147) & (g148)) + ((g823) & (!g824) & (g825) & (g826) & (!g147) & (!g148)) + ((g823) & (!g824) & (g825) & (g826) & (!g147) & (g148)) + ((g823) & (!g824) & (g825) & (g826) & (g147) & (g148)) + ((g823) & (g824) & (!g825) & (!g826) & (!g147) & (!g148)) + ((g823) & (g824) & (!g825) & (!g826) & (g147) & (!g148)) + ((g823) & (g824) & (!g825) & (g826) & (!g147) & (!g148)) + ((g823) & (g824) & (!g825) & (g826) & (g147) & (!g148)) + ((g823) & (g824) & (!g825) & (g826) & (g147) & (g148)) + ((g823) & (g824) & (g825) & (!g826) & (!g147) & (!g148)) + ((g823) & (g824) & (g825) & (!g826) & (!g147) & (g148)) + ((g823) & (g824) & (g825) & (!g826) & (g147) & (!g148)) + ((g823) & (g824) & (g825) & (g826) & (!g147) & (!g148)) + ((g823) & (g824) & (g825) & (g826) & (!g147) & (g148)) + ((g823) & (g824) & (g825) & (g826) & (g147) & (!g148)) + ((g823) & (g824) & (g825) & (g826) & (g147) & (g148)));
	assign g4477 = (((!sk[126]) & (!g2146) & (!g2542) & (g828)) + ((!sk[126]) & (!g2146) & (g2542) & (!g828)) + ((!sk[126]) & (!g2146) & (g2542) & (g828)) + ((!sk[126]) & (g2146) & (!g2542) & (g828)) + ((!sk[126]) & (g2146) & (g2542) & (!g828)) + ((!sk[126]) & (g2146) & (g2542) & (g828)) + ((sk[126]) & (!g2146) & (!g2542) & (g828)) + ((sk[126]) & (!g2146) & (g2542) & (g828)) + ((sk[126]) & (g2146) & (g2542) & (!g828)) + ((sk[126]) & (g2146) & (g2542) & (g828)));
	assign g4478 = (((!g2148) & (!sk[127]) & (!g2542) & (g829)) + ((!g2148) & (!sk[127]) & (g2542) & (!g829)) + ((!g2148) & (!sk[127]) & (g2542) & (g829)) + ((!g2148) & (sk[127]) & (!g2542) & (g829)) + ((!g2148) & (sk[127]) & (g2542) & (g829)) + ((g2148) & (!sk[127]) & (!g2542) & (g829)) + ((g2148) & (!sk[127]) & (g2542) & (!g829)) + ((g2148) & (!sk[127]) & (g2542) & (g829)) + ((g2148) & (sk[127]) & (g2542) & (!g829)) + ((g2148) & (sk[127]) & (g2542) & (g829)));
	assign g4479 = (((!g2150) & (!sk[0]) & (!g2542) & (g830)) + ((!g2150) & (!sk[0]) & (g2542) & (!g830)) + ((!g2150) & (!sk[0]) & (g2542) & (g830)) + ((!g2150) & (sk[0]) & (!g2542) & (g830)) + ((!g2150) & (sk[0]) & (g2542) & (g830)) + ((g2150) & (!sk[0]) & (!g2542) & (g830)) + ((g2150) & (!sk[0]) & (g2542) & (!g830)) + ((g2150) & (!sk[0]) & (g2542) & (g830)) + ((g2150) & (sk[0]) & (g2542) & (!g830)) + ((g2150) & (sk[0]) & (g2542) & (g830)));
	assign g4480 = (((!sk[1]) & (!g2151) & (!g2542) & (g831)) + ((!sk[1]) & (!g2151) & (g2542) & (!g831)) + ((!sk[1]) & (!g2151) & (g2542) & (g831)) + ((!sk[1]) & (g2151) & (!g2542) & (g831)) + ((!sk[1]) & (g2151) & (g2542) & (!g831)) + ((!sk[1]) & (g2151) & (g2542) & (g831)) + ((sk[1]) & (!g2151) & (!g2542) & (g831)) + ((sk[1]) & (!g2151) & (g2542) & (g831)) + ((sk[1]) & (g2151) & (g2542) & (!g831)) + ((sk[1]) & (g2151) & (g2542) & (g831)));
	assign g832 = (((!g828) & (!g829) & (!g830) & (g831) & (g147) & (g148)) + ((!g828) & (!g829) & (g830) & (!g831) & (!g147) & (g148)) + ((!g828) & (!g829) & (g830) & (g831) & (!g147) & (g148)) + ((!g828) & (!g829) & (g830) & (g831) & (g147) & (g148)) + ((!g828) & (g829) & (!g830) & (!g831) & (g147) & (!g148)) + ((!g828) & (g829) & (!g830) & (g831) & (g147) & (!g148)) + ((!g828) & (g829) & (!g830) & (g831) & (g147) & (g148)) + ((!g828) & (g829) & (g830) & (!g831) & (!g147) & (g148)) + ((!g828) & (g829) & (g830) & (!g831) & (g147) & (!g148)) + ((!g828) & (g829) & (g830) & (g831) & (!g147) & (g148)) + ((!g828) & (g829) & (g830) & (g831) & (g147) & (!g148)) + ((!g828) & (g829) & (g830) & (g831) & (g147) & (g148)) + ((g828) & (!g829) & (!g830) & (!g831) & (!g147) & (!g148)) + ((g828) & (!g829) & (!g830) & (g831) & (!g147) & (!g148)) + ((g828) & (!g829) & (!g830) & (g831) & (g147) & (g148)) + ((g828) & (!g829) & (g830) & (!g831) & (!g147) & (!g148)) + ((g828) & (!g829) & (g830) & (!g831) & (!g147) & (g148)) + ((g828) & (!g829) & (g830) & (g831) & (!g147) & (!g148)) + ((g828) & (!g829) & (g830) & (g831) & (!g147) & (g148)) + ((g828) & (!g829) & (g830) & (g831) & (g147) & (g148)) + ((g828) & (g829) & (!g830) & (!g831) & (!g147) & (!g148)) + ((g828) & (g829) & (!g830) & (!g831) & (g147) & (!g148)) + ((g828) & (g829) & (!g830) & (g831) & (!g147) & (!g148)) + ((g828) & (g829) & (!g830) & (g831) & (g147) & (!g148)) + ((g828) & (g829) & (!g830) & (g831) & (g147) & (g148)) + ((g828) & (g829) & (g830) & (!g831) & (!g147) & (!g148)) + ((g828) & (g829) & (g830) & (!g831) & (!g147) & (g148)) + ((g828) & (g829) & (g830) & (!g831) & (g147) & (!g148)) + ((g828) & (g829) & (g830) & (g831) & (!g147) & (!g148)) + ((g828) & (g829) & (g830) & (g831) & (!g147) & (g148)) + ((g828) & (g829) & (g830) & (g831) & (g147) & (!g148)) + ((g828) & (g829) & (g830) & (g831) & (g147) & (g148)));
	assign g4481 = (((!g2152) & (!sk[3]) & (!g2542) & (g833)) + ((!g2152) & (!sk[3]) & (g2542) & (!g833)) + ((!g2152) & (!sk[3]) & (g2542) & (g833)) + ((!g2152) & (sk[3]) & (!g2542) & (g833)) + ((!g2152) & (sk[3]) & (g2542) & (g833)) + ((g2152) & (!sk[3]) & (!g2542) & (g833)) + ((g2152) & (!sk[3]) & (g2542) & (!g833)) + ((g2152) & (!sk[3]) & (g2542) & (g833)) + ((g2152) & (sk[3]) & (g2542) & (!g833)) + ((g2152) & (sk[3]) & (g2542) & (g833)));
	assign g4482 = (((!sk[4]) & (!g2153) & (!g2542) & (g834)) + ((!sk[4]) & (!g2153) & (g2542) & (!g834)) + ((!sk[4]) & (!g2153) & (g2542) & (g834)) + ((!sk[4]) & (g2153) & (!g2542) & (g834)) + ((!sk[4]) & (g2153) & (g2542) & (!g834)) + ((!sk[4]) & (g2153) & (g2542) & (g834)) + ((sk[4]) & (!g2153) & (!g2542) & (g834)) + ((sk[4]) & (!g2153) & (g2542) & (g834)) + ((sk[4]) & (g2153) & (g2542) & (!g834)) + ((sk[4]) & (g2153) & (g2542) & (g834)));
	assign g4483 = (((!sk[5]) & (!g2155) & (!g2542) & (g835)) + ((!sk[5]) & (!g2155) & (g2542) & (!g835)) + ((!sk[5]) & (!g2155) & (g2542) & (g835)) + ((!sk[5]) & (g2155) & (!g2542) & (g835)) + ((!sk[5]) & (g2155) & (g2542) & (!g835)) + ((!sk[5]) & (g2155) & (g2542) & (g835)) + ((sk[5]) & (!g2155) & (!g2542) & (g835)) + ((sk[5]) & (!g2155) & (g2542) & (g835)) + ((sk[5]) & (g2155) & (g2542) & (!g835)) + ((sk[5]) & (g2155) & (g2542) & (g835)));
	assign g4484 = (((!g2157) & (!sk[6]) & (!g2542) & (g836)) + ((!g2157) & (!sk[6]) & (g2542) & (!g836)) + ((!g2157) & (!sk[6]) & (g2542) & (g836)) + ((!g2157) & (sk[6]) & (!g2542) & (g836)) + ((!g2157) & (sk[6]) & (g2542) & (g836)) + ((g2157) & (!sk[6]) & (!g2542) & (g836)) + ((g2157) & (!sk[6]) & (g2542) & (!g836)) + ((g2157) & (!sk[6]) & (g2542) & (g836)) + ((g2157) & (sk[6]) & (g2542) & (!g836)) + ((g2157) & (sk[6]) & (g2542) & (g836)));
	assign g837 = (((!g833) & (!g834) & (!g835) & (g836) & (g147) & (g148)) + ((!g833) & (!g834) & (g835) & (!g836) & (!g147) & (g148)) + ((!g833) & (!g834) & (g835) & (g836) & (!g147) & (g148)) + ((!g833) & (!g834) & (g835) & (g836) & (g147) & (g148)) + ((!g833) & (g834) & (!g835) & (!g836) & (g147) & (!g148)) + ((!g833) & (g834) & (!g835) & (g836) & (g147) & (!g148)) + ((!g833) & (g834) & (!g835) & (g836) & (g147) & (g148)) + ((!g833) & (g834) & (g835) & (!g836) & (!g147) & (g148)) + ((!g833) & (g834) & (g835) & (!g836) & (g147) & (!g148)) + ((!g833) & (g834) & (g835) & (g836) & (!g147) & (g148)) + ((!g833) & (g834) & (g835) & (g836) & (g147) & (!g148)) + ((!g833) & (g834) & (g835) & (g836) & (g147) & (g148)) + ((g833) & (!g834) & (!g835) & (!g836) & (!g147) & (!g148)) + ((g833) & (!g834) & (!g835) & (g836) & (!g147) & (!g148)) + ((g833) & (!g834) & (!g835) & (g836) & (g147) & (g148)) + ((g833) & (!g834) & (g835) & (!g836) & (!g147) & (!g148)) + ((g833) & (!g834) & (g835) & (!g836) & (!g147) & (g148)) + ((g833) & (!g834) & (g835) & (g836) & (!g147) & (!g148)) + ((g833) & (!g834) & (g835) & (g836) & (!g147) & (g148)) + ((g833) & (!g834) & (g835) & (g836) & (g147) & (g148)) + ((g833) & (g834) & (!g835) & (!g836) & (!g147) & (!g148)) + ((g833) & (g834) & (!g835) & (!g836) & (g147) & (!g148)) + ((g833) & (g834) & (!g835) & (g836) & (!g147) & (!g148)) + ((g833) & (g834) & (!g835) & (g836) & (g147) & (!g148)) + ((g833) & (g834) & (!g835) & (g836) & (g147) & (g148)) + ((g833) & (g834) & (g835) & (!g836) & (!g147) & (!g148)) + ((g833) & (g834) & (g835) & (!g836) & (!g147) & (g148)) + ((g833) & (g834) & (g835) & (!g836) & (g147) & (!g148)) + ((g833) & (g834) & (g835) & (g836) & (!g147) & (!g148)) + ((g833) & (g834) & (g835) & (g836) & (!g147) & (g148)) + ((g833) & (g834) & (g835) & (g836) & (g147) & (!g148)) + ((g833) & (g834) & (g835) & (g836) & (g147) & (g148)));
	assign g4485 = (((!g2158) & (!g2542) & (!sk[8]) & (g838)) + ((!g2158) & (!g2542) & (sk[8]) & (g838)) + ((!g2158) & (g2542) & (!sk[8]) & (!g838)) + ((!g2158) & (g2542) & (!sk[8]) & (g838)) + ((!g2158) & (g2542) & (sk[8]) & (g838)) + ((g2158) & (!g2542) & (!sk[8]) & (g838)) + ((g2158) & (g2542) & (!sk[8]) & (!g838)) + ((g2158) & (g2542) & (!sk[8]) & (g838)) + ((g2158) & (g2542) & (sk[8]) & (!g838)) + ((g2158) & (g2542) & (sk[8]) & (g838)));
	assign g4486 = (((!g2159) & (!g2542) & (!sk[9]) & (g839)) + ((!g2159) & (!g2542) & (sk[9]) & (g839)) + ((!g2159) & (g2542) & (!sk[9]) & (!g839)) + ((!g2159) & (g2542) & (!sk[9]) & (g839)) + ((!g2159) & (g2542) & (sk[9]) & (g839)) + ((g2159) & (!g2542) & (!sk[9]) & (g839)) + ((g2159) & (g2542) & (!sk[9]) & (!g839)) + ((g2159) & (g2542) & (!sk[9]) & (g839)) + ((g2159) & (g2542) & (sk[9]) & (!g839)) + ((g2159) & (g2542) & (sk[9]) & (g839)));
	assign g4487 = (((!g2160) & (!sk[10]) & (!g2542) & (g840)) + ((!g2160) & (!sk[10]) & (g2542) & (!g840)) + ((!g2160) & (!sk[10]) & (g2542) & (g840)) + ((!g2160) & (sk[10]) & (!g2542) & (g840)) + ((!g2160) & (sk[10]) & (g2542) & (g840)) + ((g2160) & (!sk[10]) & (!g2542) & (g840)) + ((g2160) & (!sk[10]) & (g2542) & (!g840)) + ((g2160) & (!sk[10]) & (g2542) & (g840)) + ((g2160) & (sk[10]) & (g2542) & (!g840)) + ((g2160) & (sk[10]) & (g2542) & (g840)));
	assign g4488 = (((!g2161) & (!g2542) & (!sk[11]) & (g841)) + ((!g2161) & (!g2542) & (sk[11]) & (g841)) + ((!g2161) & (g2542) & (!sk[11]) & (!g841)) + ((!g2161) & (g2542) & (!sk[11]) & (g841)) + ((!g2161) & (g2542) & (sk[11]) & (g841)) + ((g2161) & (!g2542) & (!sk[11]) & (g841)) + ((g2161) & (g2542) & (!sk[11]) & (!g841)) + ((g2161) & (g2542) & (!sk[11]) & (g841)) + ((g2161) & (g2542) & (sk[11]) & (!g841)) + ((g2161) & (g2542) & (sk[11]) & (g841)));
	assign g842 = (((!g838) & (!g839) & (!g840) & (g841) & (g147) & (g148)) + ((!g838) & (!g839) & (g840) & (!g841) & (!g147) & (g148)) + ((!g838) & (!g839) & (g840) & (g841) & (!g147) & (g148)) + ((!g838) & (!g839) & (g840) & (g841) & (g147) & (g148)) + ((!g838) & (g839) & (!g840) & (!g841) & (g147) & (!g148)) + ((!g838) & (g839) & (!g840) & (g841) & (g147) & (!g148)) + ((!g838) & (g839) & (!g840) & (g841) & (g147) & (g148)) + ((!g838) & (g839) & (g840) & (!g841) & (!g147) & (g148)) + ((!g838) & (g839) & (g840) & (!g841) & (g147) & (!g148)) + ((!g838) & (g839) & (g840) & (g841) & (!g147) & (g148)) + ((!g838) & (g839) & (g840) & (g841) & (g147) & (!g148)) + ((!g838) & (g839) & (g840) & (g841) & (g147) & (g148)) + ((g838) & (!g839) & (!g840) & (!g841) & (!g147) & (!g148)) + ((g838) & (!g839) & (!g840) & (g841) & (!g147) & (!g148)) + ((g838) & (!g839) & (!g840) & (g841) & (g147) & (g148)) + ((g838) & (!g839) & (g840) & (!g841) & (!g147) & (!g148)) + ((g838) & (!g839) & (g840) & (!g841) & (!g147) & (g148)) + ((g838) & (!g839) & (g840) & (g841) & (!g147) & (!g148)) + ((g838) & (!g839) & (g840) & (g841) & (!g147) & (g148)) + ((g838) & (!g839) & (g840) & (g841) & (g147) & (g148)) + ((g838) & (g839) & (!g840) & (!g841) & (!g147) & (!g148)) + ((g838) & (g839) & (!g840) & (!g841) & (g147) & (!g148)) + ((g838) & (g839) & (!g840) & (g841) & (!g147) & (!g148)) + ((g838) & (g839) & (!g840) & (g841) & (g147) & (!g148)) + ((g838) & (g839) & (!g840) & (g841) & (g147) & (g148)) + ((g838) & (g839) & (g840) & (!g841) & (!g147) & (!g148)) + ((g838) & (g839) & (g840) & (!g841) & (!g147) & (g148)) + ((g838) & (g839) & (g840) & (!g841) & (g147) & (!g148)) + ((g838) & (g839) & (g840) & (g841) & (!g147) & (!g148)) + ((g838) & (g839) & (g840) & (g841) & (!g147) & (g148)) + ((g838) & (g839) & (g840) & (g841) & (g147) & (!g148)) + ((g838) & (g839) & (g840) & (g841) & (g147) & (g148)));
	assign g843 = (((!g827) & (!g832) & (!g837) & (g842) & (g165) & (g166)) + ((!g827) & (!g832) & (g837) & (!g842) & (!g165) & (g166)) + ((!g827) & (!g832) & (g837) & (g842) & (!g165) & (g166)) + ((!g827) & (!g832) & (g837) & (g842) & (g165) & (g166)) + ((!g827) & (g832) & (!g837) & (!g842) & (g165) & (!g166)) + ((!g827) & (g832) & (!g837) & (g842) & (g165) & (!g166)) + ((!g827) & (g832) & (!g837) & (g842) & (g165) & (g166)) + ((!g827) & (g832) & (g837) & (!g842) & (!g165) & (g166)) + ((!g827) & (g832) & (g837) & (!g842) & (g165) & (!g166)) + ((!g827) & (g832) & (g837) & (g842) & (!g165) & (g166)) + ((!g827) & (g832) & (g837) & (g842) & (g165) & (!g166)) + ((!g827) & (g832) & (g837) & (g842) & (g165) & (g166)) + ((g827) & (!g832) & (!g837) & (!g842) & (!g165) & (!g166)) + ((g827) & (!g832) & (!g837) & (g842) & (!g165) & (!g166)) + ((g827) & (!g832) & (!g837) & (g842) & (g165) & (g166)) + ((g827) & (!g832) & (g837) & (!g842) & (!g165) & (!g166)) + ((g827) & (!g832) & (g837) & (!g842) & (!g165) & (g166)) + ((g827) & (!g832) & (g837) & (g842) & (!g165) & (!g166)) + ((g827) & (!g832) & (g837) & (g842) & (!g165) & (g166)) + ((g827) & (!g832) & (g837) & (g842) & (g165) & (g166)) + ((g827) & (g832) & (!g837) & (!g842) & (!g165) & (!g166)) + ((g827) & (g832) & (!g837) & (!g842) & (g165) & (!g166)) + ((g827) & (g832) & (!g837) & (g842) & (!g165) & (!g166)) + ((g827) & (g832) & (!g837) & (g842) & (g165) & (!g166)) + ((g827) & (g832) & (!g837) & (g842) & (g165) & (g166)) + ((g827) & (g832) & (g837) & (!g842) & (!g165) & (!g166)) + ((g827) & (g832) & (g837) & (!g842) & (!g165) & (g166)) + ((g827) & (g832) & (g837) & (!g842) & (g165) & (!g166)) + ((g827) & (g832) & (g837) & (g842) & (!g165) & (!g166)) + ((g827) & (g832) & (g837) & (g842) & (!g165) & (g166)) + ((g827) & (g832) & (g837) & (g842) & (g165) & (!g166)) + ((g827) & (g832) & (g837) & (g842) & (g165) & (g166)));
	assign g4489 = (((!sk[14]) & (!g2173) & (!g2542) & (g844)) + ((!sk[14]) & (!g2173) & (g2542) & (!g844)) + ((!sk[14]) & (!g2173) & (g2542) & (g844)) + ((!sk[14]) & (g2173) & (!g2542) & (g844)) + ((!sk[14]) & (g2173) & (g2542) & (!g844)) + ((!sk[14]) & (g2173) & (g2542) & (g844)) + ((sk[14]) & (!g2173) & (!g2542) & (g844)) + ((sk[14]) & (!g2173) & (g2542) & (g844)) + ((sk[14]) & (g2173) & (g2542) & (!g844)) + ((sk[14]) & (g2173) & (g2542) & (g844)));
	assign g4490 = (((!g2174) & (!sk[15]) & (!g2542) & (g845)) + ((!g2174) & (!sk[15]) & (g2542) & (!g845)) + ((!g2174) & (!sk[15]) & (g2542) & (g845)) + ((!g2174) & (sk[15]) & (!g2542) & (g845)) + ((!g2174) & (sk[15]) & (g2542) & (g845)) + ((g2174) & (!sk[15]) & (!g2542) & (g845)) + ((g2174) & (!sk[15]) & (g2542) & (!g845)) + ((g2174) & (!sk[15]) & (g2542) & (g845)) + ((g2174) & (sk[15]) & (g2542) & (!g845)) + ((g2174) & (sk[15]) & (g2542) & (g845)));
	assign g4491 = (((!g2175) & (!g2542) & (!sk[16]) & (g846)) + ((!g2175) & (!g2542) & (sk[16]) & (g846)) + ((!g2175) & (g2542) & (!sk[16]) & (!g846)) + ((!g2175) & (g2542) & (!sk[16]) & (g846)) + ((!g2175) & (g2542) & (sk[16]) & (g846)) + ((g2175) & (!g2542) & (!sk[16]) & (g846)) + ((g2175) & (g2542) & (!sk[16]) & (!g846)) + ((g2175) & (g2542) & (!sk[16]) & (g846)) + ((g2175) & (g2542) & (sk[16]) & (!g846)) + ((g2175) & (g2542) & (sk[16]) & (g846)));
	assign g4492 = (((!g2176) & (!sk[17]) & (!g2542) & (g847)) + ((!g2176) & (!sk[17]) & (g2542) & (!g847)) + ((!g2176) & (!sk[17]) & (g2542) & (g847)) + ((!g2176) & (sk[17]) & (!g2542) & (g847)) + ((!g2176) & (sk[17]) & (g2542) & (g847)) + ((g2176) & (!sk[17]) & (!g2542) & (g847)) + ((g2176) & (!sk[17]) & (g2542) & (!g847)) + ((g2176) & (!sk[17]) & (g2542) & (g847)) + ((g2176) & (sk[17]) & (g2542) & (!g847)) + ((g2176) & (sk[17]) & (g2542) & (g847)));
	assign g848 = (((!g844) & (!g845) & (!g846) & (g847) & (g165) & (g166)) + ((!g844) & (!g845) & (g846) & (!g847) & (!g165) & (g166)) + ((!g844) & (!g845) & (g846) & (g847) & (!g165) & (g166)) + ((!g844) & (!g845) & (g846) & (g847) & (g165) & (g166)) + ((!g844) & (g845) & (!g846) & (!g847) & (g165) & (!g166)) + ((!g844) & (g845) & (!g846) & (g847) & (g165) & (!g166)) + ((!g844) & (g845) & (!g846) & (g847) & (g165) & (g166)) + ((!g844) & (g845) & (g846) & (!g847) & (!g165) & (g166)) + ((!g844) & (g845) & (g846) & (!g847) & (g165) & (!g166)) + ((!g844) & (g845) & (g846) & (g847) & (!g165) & (g166)) + ((!g844) & (g845) & (g846) & (g847) & (g165) & (!g166)) + ((!g844) & (g845) & (g846) & (g847) & (g165) & (g166)) + ((g844) & (!g845) & (!g846) & (!g847) & (!g165) & (!g166)) + ((g844) & (!g845) & (!g846) & (g847) & (!g165) & (!g166)) + ((g844) & (!g845) & (!g846) & (g847) & (g165) & (g166)) + ((g844) & (!g845) & (g846) & (!g847) & (!g165) & (!g166)) + ((g844) & (!g845) & (g846) & (!g847) & (!g165) & (g166)) + ((g844) & (!g845) & (g846) & (g847) & (!g165) & (!g166)) + ((g844) & (!g845) & (g846) & (g847) & (!g165) & (g166)) + ((g844) & (!g845) & (g846) & (g847) & (g165) & (g166)) + ((g844) & (g845) & (!g846) & (!g847) & (!g165) & (!g166)) + ((g844) & (g845) & (!g846) & (!g847) & (g165) & (!g166)) + ((g844) & (g845) & (!g846) & (g847) & (!g165) & (!g166)) + ((g844) & (g845) & (!g846) & (g847) & (g165) & (!g166)) + ((g844) & (g845) & (!g846) & (g847) & (g165) & (g166)) + ((g844) & (g845) & (g846) & (!g847) & (!g165) & (!g166)) + ((g844) & (g845) & (g846) & (!g847) & (!g165) & (g166)) + ((g844) & (g845) & (g846) & (!g847) & (g165) & (!g166)) + ((g844) & (g845) & (g846) & (g847) & (!g165) & (!g166)) + ((g844) & (g845) & (g846) & (g847) & (!g165) & (g166)) + ((g844) & (g845) & (g846) & (g847) & (g165) & (!g166)) + ((g844) & (g845) & (g846) & (g847) & (g165) & (g166)));
	assign g4493 = (((!g2177) & (!g2542) & (!sk[19]) & (g849)) + ((!g2177) & (!g2542) & (sk[19]) & (g849)) + ((!g2177) & (g2542) & (!sk[19]) & (!g849)) + ((!g2177) & (g2542) & (!sk[19]) & (g849)) + ((!g2177) & (g2542) & (sk[19]) & (g849)) + ((g2177) & (!g2542) & (!sk[19]) & (g849)) + ((g2177) & (g2542) & (!sk[19]) & (!g849)) + ((g2177) & (g2542) & (!sk[19]) & (g849)) + ((g2177) & (g2542) & (sk[19]) & (!g849)) + ((g2177) & (g2542) & (sk[19]) & (g849)));
	assign g4494 = (((!sk[20]) & (!g2178) & (!g2542) & (g850)) + ((!sk[20]) & (!g2178) & (g2542) & (!g850)) + ((!sk[20]) & (!g2178) & (g2542) & (g850)) + ((!sk[20]) & (g2178) & (!g2542) & (g850)) + ((!sk[20]) & (g2178) & (g2542) & (!g850)) + ((!sk[20]) & (g2178) & (g2542) & (g850)) + ((sk[20]) & (!g2178) & (!g2542) & (g850)) + ((sk[20]) & (!g2178) & (g2542) & (g850)) + ((sk[20]) & (g2178) & (g2542) & (!g850)) + ((sk[20]) & (g2178) & (g2542) & (g850)));
	assign g4495 = (((!g2179) & (!sk[21]) & (!g2542) & (g851)) + ((!g2179) & (!sk[21]) & (g2542) & (!g851)) + ((!g2179) & (!sk[21]) & (g2542) & (g851)) + ((!g2179) & (sk[21]) & (!g2542) & (g851)) + ((!g2179) & (sk[21]) & (g2542) & (g851)) + ((g2179) & (!sk[21]) & (!g2542) & (g851)) + ((g2179) & (!sk[21]) & (g2542) & (!g851)) + ((g2179) & (!sk[21]) & (g2542) & (g851)) + ((g2179) & (sk[21]) & (g2542) & (!g851)) + ((g2179) & (sk[21]) & (g2542) & (g851)));
	assign g852 = (((!sk[22]) & (!g165) & (!g166) & (!g849) & (g850) & (!g851)) + ((!sk[22]) & (!g165) & (!g166) & (!g849) & (g850) & (g851)) + ((!sk[22]) & (!g165) & (!g166) & (g849) & (!g850) & (!g851)) + ((!sk[22]) & (!g165) & (!g166) & (g849) & (!g850) & (g851)) + ((!sk[22]) & (!g165) & (!g166) & (g849) & (g850) & (!g851)) + ((!sk[22]) & (!g165) & (!g166) & (g849) & (g850) & (g851)) + ((!sk[22]) & (!g165) & (g166) & (!g849) & (!g850) & (!g851)) + ((!sk[22]) & (!g165) & (g166) & (!g849) & (!g850) & (g851)) + ((!sk[22]) & (!g165) & (g166) & (!g849) & (g850) & (!g851)) + ((!sk[22]) & (!g165) & (g166) & (!g849) & (g850) & (g851)) + ((!sk[22]) & (!g165) & (g166) & (g849) & (!g850) & (!g851)) + ((!sk[22]) & (!g165) & (g166) & (g849) & (!g850) & (g851)) + ((!sk[22]) & (!g165) & (g166) & (g849) & (g850) & (!g851)) + ((!sk[22]) & (!g165) & (g166) & (g849) & (g850) & (g851)) + ((!sk[22]) & (g165) & (!g166) & (!g849) & (g850) & (!g851)) + ((!sk[22]) & (g165) & (!g166) & (!g849) & (g850) & (g851)) + ((!sk[22]) & (g165) & (!g166) & (g849) & (!g850) & (!g851)) + ((!sk[22]) & (g165) & (!g166) & (g849) & (!g850) & (g851)) + ((!sk[22]) & (g165) & (!g166) & (g849) & (g850) & (!g851)) + ((!sk[22]) & (g165) & (!g166) & (g849) & (g850) & (g851)) + ((!sk[22]) & (g165) & (g166) & (!g849) & (!g850) & (!g851)) + ((!sk[22]) & (g165) & (g166) & (!g849) & (!g850) & (g851)) + ((!sk[22]) & (g165) & (g166) & (!g849) & (g850) & (!g851)) + ((!sk[22]) & (g165) & (g166) & (!g849) & (g850) & (g851)) + ((!sk[22]) & (g165) & (g166) & (g849) & (!g850) & (!g851)) + ((!sk[22]) & (g165) & (g166) & (g849) & (!g850) & (g851)) + ((!sk[22]) & (g165) & (g166) & (g849) & (g850) & (!g851)) + ((!sk[22]) & (g165) & (g166) & (g849) & (g850) & (g851)) + ((sk[22]) & (!g165) & (g166) & (!g849) & (!g850) & (g851)) + ((sk[22]) & (!g165) & (g166) & (!g849) & (g850) & (g851)) + ((sk[22]) & (!g165) & (g166) & (g849) & (!g850) & (g851)) + ((sk[22]) & (!g165) & (g166) & (g849) & (g850) & (g851)) + ((sk[22]) & (g165) & (!g166) & (g849) & (!g850) & (!g851)) + ((sk[22]) & (g165) & (!g166) & (g849) & (!g850) & (g851)) + ((sk[22]) & (g165) & (!g166) & (g849) & (g850) & (!g851)) + ((sk[22]) & (g165) & (!g166) & (g849) & (g850) & (g851)) + ((sk[22]) & (g165) & (g166) & (!g849) & (g850) & (!g851)) + ((sk[22]) & (g165) & (g166) & (!g849) & (g850) & (g851)) + ((sk[22]) & (g165) & (g166) & (g849) & (g850) & (!g851)) + ((sk[22]) & (g165) & (g166) & (g849) & (g850) & (g851)));
	assign g4496 = (((!g2162) & (!g2542) & (!sk[23]) & (g853)) + ((!g2162) & (!g2542) & (sk[23]) & (g853)) + ((!g2162) & (g2542) & (!sk[23]) & (!g853)) + ((!g2162) & (g2542) & (!sk[23]) & (g853)) + ((!g2162) & (g2542) & (sk[23]) & (g853)) + ((g2162) & (!g2542) & (!sk[23]) & (g853)) + ((g2162) & (g2542) & (!sk[23]) & (!g853)) + ((g2162) & (g2542) & (!sk[23]) & (g853)) + ((g2162) & (g2542) & (sk[23]) & (!g853)) + ((g2162) & (g2542) & (sk[23]) & (g853)));
	assign g4497 = (((!g2164) & (!g2542) & (!sk[24]) & (g854)) + ((!g2164) & (!g2542) & (sk[24]) & (g854)) + ((!g2164) & (g2542) & (!sk[24]) & (!g854)) + ((!g2164) & (g2542) & (!sk[24]) & (g854)) + ((!g2164) & (g2542) & (sk[24]) & (g854)) + ((g2164) & (!g2542) & (!sk[24]) & (g854)) + ((g2164) & (g2542) & (!sk[24]) & (!g854)) + ((g2164) & (g2542) & (!sk[24]) & (g854)) + ((g2164) & (g2542) & (sk[24]) & (!g854)) + ((g2164) & (g2542) & (sk[24]) & (g854)));
	assign g4498 = (((!sk[25]) & (!g2166) & (!g2542) & (g855)) + ((!sk[25]) & (!g2166) & (g2542) & (!g855)) + ((!sk[25]) & (!g2166) & (g2542) & (g855)) + ((!sk[25]) & (g2166) & (!g2542) & (g855)) + ((!sk[25]) & (g2166) & (g2542) & (!g855)) + ((!sk[25]) & (g2166) & (g2542) & (g855)) + ((sk[25]) & (!g2166) & (!g2542) & (g855)) + ((sk[25]) & (!g2166) & (g2542) & (g855)) + ((sk[25]) & (g2166) & (g2542) & (!g855)) + ((sk[25]) & (g2166) & (g2542) & (g855)));
	assign g4499 = (((!g2168) & (!sk[26]) & (!g2542) & (g856)) + ((!g2168) & (!sk[26]) & (g2542) & (!g856)) + ((!g2168) & (!sk[26]) & (g2542) & (g856)) + ((!g2168) & (sk[26]) & (!g2542) & (g856)) + ((!g2168) & (sk[26]) & (g2542) & (g856)) + ((g2168) & (!sk[26]) & (!g2542) & (g856)) + ((g2168) & (!sk[26]) & (g2542) & (!g856)) + ((g2168) & (!sk[26]) & (g2542) & (g856)) + ((g2168) & (sk[26]) & (g2542) & (!g856)) + ((g2168) & (sk[26]) & (g2542) & (g856)));
	assign g857 = (((!g853) & (!g854) & (!g855) & (g856) & (g165) & (g166)) + ((!g853) & (!g854) & (g855) & (!g856) & (!g165) & (g166)) + ((!g853) & (!g854) & (g855) & (g856) & (!g165) & (g166)) + ((!g853) & (!g854) & (g855) & (g856) & (g165) & (g166)) + ((!g853) & (g854) & (!g855) & (!g856) & (g165) & (!g166)) + ((!g853) & (g854) & (!g855) & (g856) & (g165) & (!g166)) + ((!g853) & (g854) & (!g855) & (g856) & (g165) & (g166)) + ((!g853) & (g854) & (g855) & (!g856) & (!g165) & (g166)) + ((!g853) & (g854) & (g855) & (!g856) & (g165) & (!g166)) + ((!g853) & (g854) & (g855) & (g856) & (!g165) & (g166)) + ((!g853) & (g854) & (g855) & (g856) & (g165) & (!g166)) + ((!g853) & (g854) & (g855) & (g856) & (g165) & (g166)) + ((g853) & (!g854) & (!g855) & (!g856) & (!g165) & (!g166)) + ((g853) & (!g854) & (!g855) & (g856) & (!g165) & (!g166)) + ((g853) & (!g854) & (!g855) & (g856) & (g165) & (g166)) + ((g853) & (!g854) & (g855) & (!g856) & (!g165) & (!g166)) + ((g853) & (!g854) & (g855) & (!g856) & (!g165) & (g166)) + ((g853) & (!g854) & (g855) & (g856) & (!g165) & (!g166)) + ((g853) & (!g854) & (g855) & (g856) & (!g165) & (g166)) + ((g853) & (!g854) & (g855) & (g856) & (g165) & (g166)) + ((g853) & (g854) & (!g855) & (!g856) & (!g165) & (!g166)) + ((g853) & (g854) & (!g855) & (!g856) & (g165) & (!g166)) + ((g853) & (g854) & (!g855) & (g856) & (!g165) & (!g166)) + ((g853) & (g854) & (!g855) & (g856) & (g165) & (!g166)) + ((g853) & (g854) & (!g855) & (g856) & (g165) & (g166)) + ((g853) & (g854) & (g855) & (!g856) & (!g165) & (!g166)) + ((g853) & (g854) & (g855) & (!g856) & (!g165) & (g166)) + ((g853) & (g854) & (g855) & (!g856) & (g165) & (!g166)) + ((g853) & (g854) & (g855) & (g856) & (!g165) & (!g166)) + ((g853) & (g854) & (g855) & (g856) & (!g165) & (g166)) + ((g853) & (g854) & (g855) & (g856) & (g165) & (!g166)) + ((g853) & (g854) & (g855) & (g856) & (g165) & (g166)));
	assign g4500 = (((!sk[28]) & (!g2169) & (!g2542) & (g858)) + ((!sk[28]) & (!g2169) & (g2542) & (!g858)) + ((!sk[28]) & (!g2169) & (g2542) & (g858)) + ((!sk[28]) & (g2169) & (!g2542) & (g858)) + ((!sk[28]) & (g2169) & (g2542) & (!g858)) + ((!sk[28]) & (g2169) & (g2542) & (g858)) + ((sk[28]) & (!g2169) & (!g2542) & (g858)) + ((sk[28]) & (!g2169) & (g2542) & (g858)) + ((sk[28]) & (g2169) & (g2542) & (!g858)) + ((sk[28]) & (g2169) & (g2542) & (g858)));
	assign g4501 = (((!g2170) & (!sk[29]) & (!g2542) & (g859)) + ((!g2170) & (!sk[29]) & (g2542) & (!g859)) + ((!g2170) & (!sk[29]) & (g2542) & (g859)) + ((!g2170) & (sk[29]) & (!g2542) & (g859)) + ((!g2170) & (sk[29]) & (g2542) & (g859)) + ((g2170) & (!sk[29]) & (!g2542) & (g859)) + ((g2170) & (!sk[29]) & (g2542) & (!g859)) + ((g2170) & (!sk[29]) & (g2542) & (g859)) + ((g2170) & (sk[29]) & (g2542) & (!g859)) + ((g2170) & (sk[29]) & (g2542) & (g859)));
	assign g4502 = (((!g2171) & (!sk[30]) & (!g2542) & (g860)) + ((!g2171) & (!sk[30]) & (g2542) & (!g860)) + ((!g2171) & (!sk[30]) & (g2542) & (g860)) + ((!g2171) & (sk[30]) & (!g2542) & (g860)) + ((!g2171) & (sk[30]) & (g2542) & (g860)) + ((g2171) & (!sk[30]) & (!g2542) & (g860)) + ((g2171) & (!sk[30]) & (g2542) & (!g860)) + ((g2171) & (!sk[30]) & (g2542) & (g860)) + ((g2171) & (sk[30]) & (g2542) & (!g860)) + ((g2171) & (sk[30]) & (g2542) & (g860)));
	assign g4503 = (((!g2172) & (!g2542) & (!sk[31]) & (g861)) + ((!g2172) & (!g2542) & (sk[31]) & (g861)) + ((!g2172) & (g2542) & (!sk[31]) & (!g861)) + ((!g2172) & (g2542) & (!sk[31]) & (g861)) + ((!g2172) & (g2542) & (sk[31]) & (g861)) + ((g2172) & (!g2542) & (!sk[31]) & (g861)) + ((g2172) & (g2542) & (!sk[31]) & (!g861)) + ((g2172) & (g2542) & (!sk[31]) & (g861)) + ((g2172) & (g2542) & (sk[31]) & (!g861)) + ((g2172) & (g2542) & (sk[31]) & (g861)));
	assign g862 = (((!g858) & (!g859) & (!g860) & (g861) & (g165) & (g166)) + ((!g858) & (!g859) & (g860) & (!g861) & (!g165) & (g166)) + ((!g858) & (!g859) & (g860) & (g861) & (!g165) & (g166)) + ((!g858) & (!g859) & (g860) & (g861) & (g165) & (g166)) + ((!g858) & (g859) & (!g860) & (!g861) & (g165) & (!g166)) + ((!g858) & (g859) & (!g860) & (g861) & (g165) & (!g166)) + ((!g858) & (g859) & (!g860) & (g861) & (g165) & (g166)) + ((!g858) & (g859) & (g860) & (!g861) & (!g165) & (g166)) + ((!g858) & (g859) & (g860) & (!g861) & (g165) & (!g166)) + ((!g858) & (g859) & (g860) & (g861) & (!g165) & (g166)) + ((!g858) & (g859) & (g860) & (g861) & (g165) & (!g166)) + ((!g858) & (g859) & (g860) & (g861) & (g165) & (g166)) + ((g858) & (!g859) & (!g860) & (!g861) & (!g165) & (!g166)) + ((g858) & (!g859) & (!g860) & (g861) & (!g165) & (!g166)) + ((g858) & (!g859) & (!g860) & (g861) & (g165) & (g166)) + ((g858) & (!g859) & (g860) & (!g861) & (!g165) & (!g166)) + ((g858) & (!g859) & (g860) & (!g861) & (!g165) & (g166)) + ((g858) & (!g859) & (g860) & (g861) & (!g165) & (!g166)) + ((g858) & (!g859) & (g860) & (g861) & (!g165) & (g166)) + ((g858) & (!g859) & (g860) & (g861) & (g165) & (g166)) + ((g858) & (g859) & (!g860) & (!g861) & (!g165) & (!g166)) + ((g858) & (g859) & (!g860) & (!g861) & (g165) & (!g166)) + ((g858) & (g859) & (!g860) & (g861) & (!g165) & (!g166)) + ((g858) & (g859) & (!g860) & (g861) & (g165) & (!g166)) + ((g858) & (g859) & (!g860) & (g861) & (g165) & (g166)) + ((g858) & (g859) & (g860) & (!g861) & (!g165) & (!g166)) + ((g858) & (g859) & (g860) & (!g861) & (!g165) & (g166)) + ((g858) & (g859) & (g860) & (!g861) & (g165) & (!g166)) + ((g858) & (g859) & (g860) & (g861) & (!g165) & (!g166)) + ((g858) & (g859) & (g860) & (g861) & (!g165) & (g166)) + ((g858) & (g859) & (g860) & (g861) & (g165) & (!g166)) + ((g858) & (g859) & (g860) & (g861) & (g165) & (g166)));
	assign g863 = (((!g147) & (!g148) & (!g848) & (g852) & (!g857) & (!g862)) + ((!g147) & (!g148) & (!g848) & (g852) & (!g857) & (g862)) + ((!g147) & (!g148) & (!g848) & (g852) & (g857) & (!g862)) + ((!g147) & (!g148) & (!g848) & (g852) & (g857) & (g862)) + ((!g147) & (!g148) & (g848) & (g852) & (!g857) & (!g862)) + ((!g147) & (!g148) & (g848) & (g852) & (!g857) & (g862)) + ((!g147) & (!g148) & (g848) & (g852) & (g857) & (!g862)) + ((!g147) & (!g148) & (g848) & (g852) & (g857) & (g862)) + ((!g147) & (g148) & (!g848) & (!g852) & (!g857) & (g862)) + ((!g147) & (g148) & (!g848) & (!g852) & (g857) & (g862)) + ((!g147) & (g148) & (!g848) & (g852) & (!g857) & (g862)) + ((!g147) & (g148) & (!g848) & (g852) & (g857) & (g862)) + ((!g147) & (g148) & (g848) & (!g852) & (!g857) & (g862)) + ((!g147) & (g148) & (g848) & (!g852) & (g857) & (g862)) + ((!g147) & (g148) & (g848) & (g852) & (!g857) & (g862)) + ((!g147) & (g148) & (g848) & (g852) & (g857) & (g862)) + ((g147) & (!g148) & (g848) & (!g852) & (!g857) & (!g862)) + ((g147) & (!g148) & (g848) & (!g852) & (!g857) & (g862)) + ((g147) & (!g148) & (g848) & (!g852) & (g857) & (!g862)) + ((g147) & (!g148) & (g848) & (!g852) & (g857) & (g862)) + ((g147) & (!g148) & (g848) & (g852) & (!g857) & (!g862)) + ((g147) & (!g148) & (g848) & (g852) & (!g857) & (g862)) + ((g147) & (!g148) & (g848) & (g852) & (g857) & (!g862)) + ((g147) & (!g148) & (g848) & (g852) & (g857) & (g862)) + ((g147) & (g148) & (!g848) & (!g852) & (g857) & (!g862)) + ((g147) & (g148) & (!g848) & (!g852) & (g857) & (g862)) + ((g147) & (g148) & (!g848) & (g852) & (g857) & (!g862)) + ((g147) & (g148) & (!g848) & (g852) & (g857) & (g862)) + ((g147) & (g148) & (g848) & (!g852) & (g857) & (!g862)) + ((g147) & (g148) & (g848) & (!g852) & (g857) & (g862)) + ((g147) & (g148) & (g848) & (g852) & (g857) & (!g862)) + ((g147) & (g148) & (g848) & (g852) & (g857) & (g862)));
	assign g864 = (((!sk[34]) & (!g142) & (!g843) & (g863)) + ((!sk[34]) & (!g142) & (g843) & (!g863)) + ((!sk[34]) & (!g142) & (g843) & (g863)) + ((!sk[34]) & (g142) & (!g843) & (g863)) + ((!sk[34]) & (g142) & (g843) & (!g863)) + ((!sk[34]) & (g142) & (g843) & (g863)) + ((sk[34]) & (!g142) & (!g843) & (g863)) + ((sk[34]) & (!g142) & (g843) & (g863)) + ((sk[34]) & (g142) & (g843) & (!g863)) + ((sk[34]) & (g142) & (g843) & (g863)));
	assign g4504 = (((!g2059) & (!sk[35]) & (!g2548) & (g865)) + ((!g2059) & (!sk[35]) & (g2548) & (!g865)) + ((!g2059) & (!sk[35]) & (g2548) & (g865)) + ((!g2059) & (sk[35]) & (!g2548) & (g865)) + ((!g2059) & (sk[35]) & (g2548) & (g865)) + ((g2059) & (!sk[35]) & (!g2548) & (g865)) + ((g2059) & (!sk[35]) & (g2548) & (!g865)) + ((g2059) & (!sk[35]) & (g2548) & (g865)) + ((g2059) & (sk[35]) & (g2548) & (!g865)) + ((g2059) & (sk[35]) & (g2548) & (g865)));
	assign g866 = (((!g817) & (!g819) & (!sk[36]) & (g821)) + ((!g817) & (g819) & (!sk[36]) & (!g821)) + ((!g817) & (g819) & (!sk[36]) & (g821)) + ((!g817) & (g819) & (sk[36]) & (!g821)) + ((g817) & (!g819) & (!sk[36]) & (g821)) + ((g817) & (!g819) & (sk[36]) & (!g821)) + ((g817) & (g819) & (!sk[36]) & (!g821)) + ((g817) & (g819) & (!sk[36]) & (g821)) + ((g817) & (g819) & (sk[36]) & (!g821)) + ((g817) & (g819) & (sk[36]) & (g821)));
	assign g4505 = (((!sk[37]) & (!g2064) & (!dmem_dat_ix15x) & (g867)) + ((!sk[37]) & (!g2064) & (dmem_dat_ix15x) & (!g867)) + ((!sk[37]) & (!g2064) & (dmem_dat_ix15x) & (g867)) + ((!sk[37]) & (g2064) & (!dmem_dat_ix15x) & (g867)) + ((!sk[37]) & (g2064) & (dmem_dat_ix15x) & (!g867)) + ((!sk[37]) & (g2064) & (dmem_dat_ix15x) & (g867)) + ((sk[37]) & (!g2064) & (!dmem_dat_ix15x) & (g867)) + ((sk[37]) & (!g2064) & (dmem_dat_ix15x) & (g867)) + ((sk[37]) & (g2064) & (dmem_dat_ix15x) & (!g867)) + ((sk[37]) & (g2064) & (dmem_dat_ix15x) & (g867)));
	assign g868 = (((!sk[38]) & (!g679) & (!g107) & (g867)) + ((!sk[38]) & (!g679) & (g107) & (!g867)) + ((!sk[38]) & (!g679) & (g107) & (g867)) + ((!sk[38]) & (g679) & (!g107) & (g867)) + ((!sk[38]) & (g679) & (g107) & (!g867)) + ((!sk[38]) & (g679) & (g107) & (g867)) + ((sk[38]) & (!g679) & (!g107) & (!g867)) + ((sk[38]) & (!g679) & (!g107) & (g867)) + ((sk[38]) & (g679) & (!g107) & (!g867)) + ((sk[38]) & (g679) & (g107) & (!g867)));
	assign g869 = (((!sk[39]) & (!g126) & (!g864) & (!g865) & (g866) & (!g868)) + ((!sk[39]) & (!g126) & (!g864) & (!g865) & (g866) & (g868)) + ((!sk[39]) & (!g126) & (!g864) & (g865) & (!g866) & (!g868)) + ((!sk[39]) & (!g126) & (!g864) & (g865) & (!g866) & (g868)) + ((!sk[39]) & (!g126) & (!g864) & (g865) & (g866) & (!g868)) + ((!sk[39]) & (!g126) & (!g864) & (g865) & (g866) & (g868)) + ((!sk[39]) & (!g126) & (g864) & (!g865) & (!g866) & (!g868)) + ((!sk[39]) & (!g126) & (g864) & (!g865) & (!g866) & (g868)) + ((!sk[39]) & (!g126) & (g864) & (!g865) & (g866) & (!g868)) + ((!sk[39]) & (!g126) & (g864) & (!g865) & (g866) & (g868)) + ((!sk[39]) & (!g126) & (g864) & (g865) & (!g866) & (!g868)) + ((!sk[39]) & (!g126) & (g864) & (g865) & (!g866) & (g868)) + ((!sk[39]) & (!g126) & (g864) & (g865) & (g866) & (!g868)) + ((!sk[39]) & (!g126) & (g864) & (g865) & (g866) & (g868)) + ((!sk[39]) & (g126) & (!g864) & (!g865) & (g866) & (!g868)) + ((!sk[39]) & (g126) & (!g864) & (!g865) & (g866) & (g868)) + ((!sk[39]) & (g126) & (!g864) & (g865) & (!g866) & (!g868)) + ((!sk[39]) & (g126) & (!g864) & (g865) & (!g866) & (g868)) + ((!sk[39]) & (g126) & (!g864) & (g865) & (g866) & (!g868)) + ((!sk[39]) & (g126) & (!g864) & (g865) & (g866) & (g868)) + ((!sk[39]) & (g126) & (g864) & (!g865) & (!g866) & (!g868)) + ((!sk[39]) & (g126) & (g864) & (!g865) & (!g866) & (g868)) + ((!sk[39]) & (g126) & (g864) & (!g865) & (g866) & (!g868)) + ((!sk[39]) & (g126) & (g864) & (!g865) & (g866) & (g868)) + ((!sk[39]) & (g126) & (g864) & (g865) & (!g866) & (!g868)) + ((!sk[39]) & (g126) & (g864) & (g865) & (!g866) & (g868)) + ((!sk[39]) & (g126) & (g864) & (g865) & (g866) & (!g868)) + ((!sk[39]) & (g126) & (g864) & (g865) & (g866) & (g868)) + ((sk[39]) & (!g126) & (!g864) & (g865) & (!g866) & (!g868)) + ((sk[39]) & (!g126) & (!g864) & (g865) & (!g866) & (g868)) + ((sk[39]) & (!g126) & (!g864) & (g865) & (g866) & (!g868)) + ((sk[39]) & (!g126) & (!g864) & (g865) & (g866) & (g868)) + ((sk[39]) & (!g126) & (g864) & (g865) & (!g866) & (!g868)) + ((sk[39]) & (!g126) & (g864) & (g865) & (!g866) & (g868)) + ((sk[39]) & (!g126) & (g864) & (g865) & (g866) & (!g868)) + ((sk[39]) & (!g126) & (g864) & (g865) & (g866) & (g868)) + ((sk[39]) & (g126) & (!g864) & (!g865) & (!g866) & (!g868)) + ((sk[39]) & (g126) & (!g864) & (!g865) & (g866) & (g868)) + ((sk[39]) & (g126) & (!g864) & (g865) & (!g866) & (!g868)) + ((sk[39]) & (g126) & (!g864) & (g865) & (g866) & (g868)) + ((sk[39]) & (g126) & (g864) & (!g865) & (!g866) & (g868)) + ((sk[39]) & (g126) & (g864) & (!g865) & (g866) & (!g868)) + ((sk[39]) & (g126) & (g864) & (g865) & (!g866) & (g868)) + ((sk[39]) & (g126) & (g864) & (g865) & (g866) & (!g868)));
	assign g4506 = (((!g2140) & (!g3539) & (!sk[40]) & (g870)) + ((!g2140) & (!g3539) & (sk[40]) & (g870)) + ((!g2140) & (g3539) & (!sk[40]) & (!g870)) + ((!g2140) & (g3539) & (!sk[40]) & (g870)) + ((!g2140) & (g3539) & (sk[40]) & (g870)) + ((g2140) & (!g3539) & (!sk[40]) & (g870)) + ((g2140) & (g3539) & (!sk[40]) & (!g870)) + ((g2140) & (g3539) & (!sk[40]) & (g870)) + ((g2140) & (g3539) & (sk[40]) & (!g870)) + ((g2140) & (g3539) & (sk[40]) & (g870)));
	assign g4507 = (((!g2142) & (!g3539) & (!sk[41]) & (g871)) + ((!g2142) & (!g3539) & (sk[41]) & (g871)) + ((!g2142) & (g3539) & (!sk[41]) & (!g871)) + ((!g2142) & (g3539) & (!sk[41]) & (g871)) + ((!g2142) & (g3539) & (sk[41]) & (g871)) + ((g2142) & (!g3539) & (!sk[41]) & (g871)) + ((g2142) & (g3539) & (!sk[41]) & (!g871)) + ((g2142) & (g3539) & (!sk[41]) & (g871)) + ((g2142) & (g3539) & (sk[41]) & (!g871)) + ((g2142) & (g3539) & (sk[41]) & (g871)));
	assign g4508 = (((!g2144) & (!g3539) & (!sk[42]) & (g872)) + ((!g2144) & (!g3539) & (sk[42]) & (g872)) + ((!g2144) & (g3539) & (!sk[42]) & (!g872)) + ((!g2144) & (g3539) & (!sk[42]) & (g872)) + ((!g2144) & (g3539) & (sk[42]) & (g872)) + ((g2144) & (!g3539) & (!sk[42]) & (g872)) + ((g2144) & (g3539) & (!sk[42]) & (!g872)) + ((g2144) & (g3539) & (!sk[42]) & (g872)) + ((g2144) & (g3539) & (sk[42]) & (!g872)) + ((g2144) & (g3539) & (sk[42]) & (g872)));
	assign g4509 = (((!g2145) & (!g3539) & (!sk[43]) & (g873)) + ((!g2145) & (!g3539) & (sk[43]) & (g873)) + ((!g2145) & (g3539) & (!sk[43]) & (!g873)) + ((!g2145) & (g3539) & (!sk[43]) & (g873)) + ((!g2145) & (g3539) & (sk[43]) & (g873)) + ((g2145) & (!g3539) & (!sk[43]) & (g873)) + ((g2145) & (g3539) & (!sk[43]) & (!g873)) + ((g2145) & (g3539) & (!sk[43]) & (g873)) + ((g2145) & (g3539) & (sk[43]) & (!g873)) + ((g2145) & (g3539) & (sk[43]) & (g873)));
	assign g874 = (((!g870) & (!g871) & (!g872) & (g873) & (g147) & (g148)) + ((!g870) & (!g871) & (g872) & (!g873) & (!g147) & (g148)) + ((!g870) & (!g871) & (g872) & (g873) & (!g147) & (g148)) + ((!g870) & (!g871) & (g872) & (g873) & (g147) & (g148)) + ((!g870) & (g871) & (!g872) & (!g873) & (g147) & (!g148)) + ((!g870) & (g871) & (!g872) & (g873) & (g147) & (!g148)) + ((!g870) & (g871) & (!g872) & (g873) & (g147) & (g148)) + ((!g870) & (g871) & (g872) & (!g873) & (!g147) & (g148)) + ((!g870) & (g871) & (g872) & (!g873) & (g147) & (!g148)) + ((!g870) & (g871) & (g872) & (g873) & (!g147) & (g148)) + ((!g870) & (g871) & (g872) & (g873) & (g147) & (!g148)) + ((!g870) & (g871) & (g872) & (g873) & (g147) & (g148)) + ((g870) & (!g871) & (!g872) & (!g873) & (!g147) & (!g148)) + ((g870) & (!g871) & (!g872) & (g873) & (!g147) & (!g148)) + ((g870) & (!g871) & (!g872) & (g873) & (g147) & (g148)) + ((g870) & (!g871) & (g872) & (!g873) & (!g147) & (!g148)) + ((g870) & (!g871) & (g872) & (!g873) & (!g147) & (g148)) + ((g870) & (!g871) & (g872) & (g873) & (!g147) & (!g148)) + ((g870) & (!g871) & (g872) & (g873) & (!g147) & (g148)) + ((g870) & (!g871) & (g872) & (g873) & (g147) & (g148)) + ((g870) & (g871) & (!g872) & (!g873) & (!g147) & (!g148)) + ((g870) & (g871) & (!g872) & (!g873) & (g147) & (!g148)) + ((g870) & (g871) & (!g872) & (g873) & (!g147) & (!g148)) + ((g870) & (g871) & (!g872) & (g873) & (g147) & (!g148)) + ((g870) & (g871) & (!g872) & (g873) & (g147) & (g148)) + ((g870) & (g871) & (g872) & (!g873) & (!g147) & (!g148)) + ((g870) & (g871) & (g872) & (!g873) & (!g147) & (g148)) + ((g870) & (g871) & (g872) & (!g873) & (g147) & (!g148)) + ((g870) & (g871) & (g872) & (g873) & (!g147) & (!g148)) + ((g870) & (g871) & (g872) & (g873) & (!g147) & (g148)) + ((g870) & (g871) & (g872) & (g873) & (g147) & (!g148)) + ((g870) & (g871) & (g872) & (g873) & (g147) & (g148)));
	assign g4510 = (((!g2146) & (!sk[45]) & (!g3539) & (g875)) + ((!g2146) & (!sk[45]) & (g3539) & (!g875)) + ((!g2146) & (!sk[45]) & (g3539) & (g875)) + ((!g2146) & (sk[45]) & (!g3539) & (g875)) + ((!g2146) & (sk[45]) & (g3539) & (g875)) + ((g2146) & (!sk[45]) & (!g3539) & (g875)) + ((g2146) & (!sk[45]) & (g3539) & (!g875)) + ((g2146) & (!sk[45]) & (g3539) & (g875)) + ((g2146) & (sk[45]) & (g3539) & (!g875)) + ((g2146) & (sk[45]) & (g3539) & (g875)));
	assign g4511 = (((!g2148) & (!g3539) & (!sk[46]) & (g876)) + ((!g2148) & (!g3539) & (sk[46]) & (g876)) + ((!g2148) & (g3539) & (!sk[46]) & (!g876)) + ((!g2148) & (g3539) & (!sk[46]) & (g876)) + ((!g2148) & (g3539) & (sk[46]) & (g876)) + ((g2148) & (!g3539) & (!sk[46]) & (g876)) + ((g2148) & (g3539) & (!sk[46]) & (!g876)) + ((g2148) & (g3539) & (!sk[46]) & (g876)) + ((g2148) & (g3539) & (sk[46]) & (!g876)) + ((g2148) & (g3539) & (sk[46]) & (g876)));
	assign g4512 = (((!sk[47]) & (!g2150) & (!g3539) & (g877)) + ((!sk[47]) & (!g2150) & (g3539) & (!g877)) + ((!sk[47]) & (!g2150) & (g3539) & (g877)) + ((!sk[47]) & (g2150) & (!g3539) & (g877)) + ((!sk[47]) & (g2150) & (g3539) & (!g877)) + ((!sk[47]) & (g2150) & (g3539) & (g877)) + ((sk[47]) & (!g2150) & (!g3539) & (g877)) + ((sk[47]) & (!g2150) & (g3539) & (g877)) + ((sk[47]) & (g2150) & (g3539) & (!g877)) + ((sk[47]) & (g2150) & (g3539) & (g877)));
	assign g4513 = (((!sk[48]) & (!g2151) & (!g3539) & (g878)) + ((!sk[48]) & (!g2151) & (g3539) & (!g878)) + ((!sk[48]) & (!g2151) & (g3539) & (g878)) + ((!sk[48]) & (g2151) & (!g3539) & (g878)) + ((!sk[48]) & (g2151) & (g3539) & (!g878)) + ((!sk[48]) & (g2151) & (g3539) & (g878)) + ((sk[48]) & (!g2151) & (!g3539) & (g878)) + ((sk[48]) & (!g2151) & (g3539) & (g878)) + ((sk[48]) & (g2151) & (g3539) & (!g878)) + ((sk[48]) & (g2151) & (g3539) & (g878)));
	assign g879 = (((!g875) & (!g876) & (!g877) & (g878) & (g147) & (g148)) + ((!g875) & (!g876) & (g877) & (!g878) & (!g147) & (g148)) + ((!g875) & (!g876) & (g877) & (g878) & (!g147) & (g148)) + ((!g875) & (!g876) & (g877) & (g878) & (g147) & (g148)) + ((!g875) & (g876) & (!g877) & (!g878) & (g147) & (!g148)) + ((!g875) & (g876) & (!g877) & (g878) & (g147) & (!g148)) + ((!g875) & (g876) & (!g877) & (g878) & (g147) & (g148)) + ((!g875) & (g876) & (g877) & (!g878) & (!g147) & (g148)) + ((!g875) & (g876) & (g877) & (!g878) & (g147) & (!g148)) + ((!g875) & (g876) & (g877) & (g878) & (!g147) & (g148)) + ((!g875) & (g876) & (g877) & (g878) & (g147) & (!g148)) + ((!g875) & (g876) & (g877) & (g878) & (g147) & (g148)) + ((g875) & (!g876) & (!g877) & (!g878) & (!g147) & (!g148)) + ((g875) & (!g876) & (!g877) & (g878) & (!g147) & (!g148)) + ((g875) & (!g876) & (!g877) & (g878) & (g147) & (g148)) + ((g875) & (!g876) & (g877) & (!g878) & (!g147) & (!g148)) + ((g875) & (!g876) & (g877) & (!g878) & (!g147) & (g148)) + ((g875) & (!g876) & (g877) & (g878) & (!g147) & (!g148)) + ((g875) & (!g876) & (g877) & (g878) & (!g147) & (g148)) + ((g875) & (!g876) & (g877) & (g878) & (g147) & (g148)) + ((g875) & (g876) & (!g877) & (!g878) & (!g147) & (!g148)) + ((g875) & (g876) & (!g877) & (!g878) & (g147) & (!g148)) + ((g875) & (g876) & (!g877) & (g878) & (!g147) & (!g148)) + ((g875) & (g876) & (!g877) & (g878) & (g147) & (!g148)) + ((g875) & (g876) & (!g877) & (g878) & (g147) & (g148)) + ((g875) & (g876) & (g877) & (!g878) & (!g147) & (!g148)) + ((g875) & (g876) & (g877) & (!g878) & (!g147) & (g148)) + ((g875) & (g876) & (g877) & (!g878) & (g147) & (!g148)) + ((g875) & (g876) & (g877) & (g878) & (!g147) & (!g148)) + ((g875) & (g876) & (g877) & (g878) & (!g147) & (g148)) + ((g875) & (g876) & (g877) & (g878) & (g147) & (!g148)) + ((g875) & (g876) & (g877) & (g878) & (g147) & (g148)));
	assign g4514 = (((!g2152) & (!g3539) & (!sk[50]) & (g880)) + ((!g2152) & (!g3539) & (sk[50]) & (g880)) + ((!g2152) & (g3539) & (!sk[50]) & (!g880)) + ((!g2152) & (g3539) & (!sk[50]) & (g880)) + ((!g2152) & (g3539) & (sk[50]) & (g880)) + ((g2152) & (!g3539) & (!sk[50]) & (g880)) + ((g2152) & (g3539) & (!sk[50]) & (!g880)) + ((g2152) & (g3539) & (!sk[50]) & (g880)) + ((g2152) & (g3539) & (sk[50]) & (!g880)) + ((g2152) & (g3539) & (sk[50]) & (g880)));
	assign g4515 = (((!sk[51]) & (!g2153) & (!g3539) & (g881)) + ((!sk[51]) & (!g2153) & (g3539) & (!g881)) + ((!sk[51]) & (!g2153) & (g3539) & (g881)) + ((!sk[51]) & (g2153) & (!g3539) & (g881)) + ((!sk[51]) & (g2153) & (g3539) & (!g881)) + ((!sk[51]) & (g2153) & (g3539) & (g881)) + ((sk[51]) & (!g2153) & (!g3539) & (g881)) + ((sk[51]) & (!g2153) & (g3539) & (g881)) + ((sk[51]) & (g2153) & (g3539) & (!g881)) + ((sk[51]) & (g2153) & (g3539) & (g881)));
	assign g4516 = (((!g2155) & (!sk[52]) & (!g3539) & (g882)) + ((!g2155) & (!sk[52]) & (g3539) & (!g882)) + ((!g2155) & (!sk[52]) & (g3539) & (g882)) + ((!g2155) & (sk[52]) & (!g3539) & (g882)) + ((!g2155) & (sk[52]) & (g3539) & (g882)) + ((g2155) & (!sk[52]) & (!g3539) & (g882)) + ((g2155) & (!sk[52]) & (g3539) & (!g882)) + ((g2155) & (!sk[52]) & (g3539) & (g882)) + ((g2155) & (sk[52]) & (g3539) & (!g882)) + ((g2155) & (sk[52]) & (g3539) & (g882)));
	assign g4517 = (((!g2157) & (!g3539) & (!sk[53]) & (g883)) + ((!g2157) & (!g3539) & (sk[53]) & (g883)) + ((!g2157) & (g3539) & (!sk[53]) & (!g883)) + ((!g2157) & (g3539) & (!sk[53]) & (g883)) + ((!g2157) & (g3539) & (sk[53]) & (g883)) + ((g2157) & (!g3539) & (!sk[53]) & (g883)) + ((g2157) & (g3539) & (!sk[53]) & (!g883)) + ((g2157) & (g3539) & (!sk[53]) & (g883)) + ((g2157) & (g3539) & (sk[53]) & (!g883)) + ((g2157) & (g3539) & (sk[53]) & (g883)));
	assign g884 = (((!g880) & (!g881) & (!g882) & (g883) & (g147) & (g148)) + ((!g880) & (!g881) & (g882) & (!g883) & (!g147) & (g148)) + ((!g880) & (!g881) & (g882) & (g883) & (!g147) & (g148)) + ((!g880) & (!g881) & (g882) & (g883) & (g147) & (g148)) + ((!g880) & (g881) & (!g882) & (!g883) & (g147) & (!g148)) + ((!g880) & (g881) & (!g882) & (g883) & (g147) & (!g148)) + ((!g880) & (g881) & (!g882) & (g883) & (g147) & (g148)) + ((!g880) & (g881) & (g882) & (!g883) & (!g147) & (g148)) + ((!g880) & (g881) & (g882) & (!g883) & (g147) & (!g148)) + ((!g880) & (g881) & (g882) & (g883) & (!g147) & (g148)) + ((!g880) & (g881) & (g882) & (g883) & (g147) & (!g148)) + ((!g880) & (g881) & (g882) & (g883) & (g147) & (g148)) + ((g880) & (!g881) & (!g882) & (!g883) & (!g147) & (!g148)) + ((g880) & (!g881) & (!g882) & (g883) & (!g147) & (!g148)) + ((g880) & (!g881) & (!g882) & (g883) & (g147) & (g148)) + ((g880) & (!g881) & (g882) & (!g883) & (!g147) & (!g148)) + ((g880) & (!g881) & (g882) & (!g883) & (!g147) & (g148)) + ((g880) & (!g881) & (g882) & (g883) & (!g147) & (!g148)) + ((g880) & (!g881) & (g882) & (g883) & (!g147) & (g148)) + ((g880) & (!g881) & (g882) & (g883) & (g147) & (g148)) + ((g880) & (g881) & (!g882) & (!g883) & (!g147) & (!g148)) + ((g880) & (g881) & (!g882) & (!g883) & (g147) & (!g148)) + ((g880) & (g881) & (!g882) & (g883) & (!g147) & (!g148)) + ((g880) & (g881) & (!g882) & (g883) & (g147) & (!g148)) + ((g880) & (g881) & (!g882) & (g883) & (g147) & (g148)) + ((g880) & (g881) & (g882) & (!g883) & (!g147) & (!g148)) + ((g880) & (g881) & (g882) & (!g883) & (!g147) & (g148)) + ((g880) & (g881) & (g882) & (!g883) & (g147) & (!g148)) + ((g880) & (g881) & (g882) & (g883) & (!g147) & (!g148)) + ((g880) & (g881) & (g882) & (g883) & (!g147) & (g148)) + ((g880) & (g881) & (g882) & (g883) & (g147) & (!g148)) + ((g880) & (g881) & (g882) & (g883) & (g147) & (g148)));
	assign g4518 = (((!g2158) & (!sk[55]) & (!g3539) & (g885)) + ((!g2158) & (!sk[55]) & (g3539) & (!g885)) + ((!g2158) & (!sk[55]) & (g3539) & (g885)) + ((!g2158) & (sk[55]) & (!g3539) & (g885)) + ((!g2158) & (sk[55]) & (g3539) & (g885)) + ((g2158) & (!sk[55]) & (!g3539) & (g885)) + ((g2158) & (!sk[55]) & (g3539) & (!g885)) + ((g2158) & (!sk[55]) & (g3539) & (g885)) + ((g2158) & (sk[55]) & (g3539) & (!g885)) + ((g2158) & (sk[55]) & (g3539) & (g885)));
	assign g4519 = (((!g2159) & (!g3539) & (!sk[56]) & (g886)) + ((!g2159) & (!g3539) & (sk[56]) & (g886)) + ((!g2159) & (g3539) & (!sk[56]) & (!g886)) + ((!g2159) & (g3539) & (!sk[56]) & (g886)) + ((!g2159) & (g3539) & (sk[56]) & (g886)) + ((g2159) & (!g3539) & (!sk[56]) & (g886)) + ((g2159) & (g3539) & (!sk[56]) & (!g886)) + ((g2159) & (g3539) & (!sk[56]) & (g886)) + ((g2159) & (g3539) & (sk[56]) & (!g886)) + ((g2159) & (g3539) & (sk[56]) & (g886)));
	assign g4520 = (((!g2160) & (!sk[57]) & (!g3539) & (g887)) + ((!g2160) & (!sk[57]) & (g3539) & (!g887)) + ((!g2160) & (!sk[57]) & (g3539) & (g887)) + ((!g2160) & (sk[57]) & (!g3539) & (g887)) + ((!g2160) & (sk[57]) & (g3539) & (g887)) + ((g2160) & (!sk[57]) & (!g3539) & (g887)) + ((g2160) & (!sk[57]) & (g3539) & (!g887)) + ((g2160) & (!sk[57]) & (g3539) & (g887)) + ((g2160) & (sk[57]) & (g3539) & (!g887)) + ((g2160) & (sk[57]) & (g3539) & (g887)));
	assign g4521 = (((!g2161) & (!sk[58]) & (!g3539) & (g888)) + ((!g2161) & (!sk[58]) & (g3539) & (!g888)) + ((!g2161) & (!sk[58]) & (g3539) & (g888)) + ((!g2161) & (sk[58]) & (!g3539) & (g888)) + ((!g2161) & (sk[58]) & (g3539) & (g888)) + ((g2161) & (!sk[58]) & (!g3539) & (g888)) + ((g2161) & (!sk[58]) & (g3539) & (!g888)) + ((g2161) & (!sk[58]) & (g3539) & (g888)) + ((g2161) & (sk[58]) & (g3539) & (!g888)) + ((g2161) & (sk[58]) & (g3539) & (g888)));
	assign g889 = (((!g885) & (!g886) & (!g887) & (g888) & (g147) & (g148)) + ((!g885) & (!g886) & (g887) & (!g888) & (!g147) & (g148)) + ((!g885) & (!g886) & (g887) & (g888) & (!g147) & (g148)) + ((!g885) & (!g886) & (g887) & (g888) & (g147) & (g148)) + ((!g885) & (g886) & (!g887) & (!g888) & (g147) & (!g148)) + ((!g885) & (g886) & (!g887) & (g888) & (g147) & (!g148)) + ((!g885) & (g886) & (!g887) & (g888) & (g147) & (g148)) + ((!g885) & (g886) & (g887) & (!g888) & (!g147) & (g148)) + ((!g885) & (g886) & (g887) & (!g888) & (g147) & (!g148)) + ((!g885) & (g886) & (g887) & (g888) & (!g147) & (g148)) + ((!g885) & (g886) & (g887) & (g888) & (g147) & (!g148)) + ((!g885) & (g886) & (g887) & (g888) & (g147) & (g148)) + ((g885) & (!g886) & (!g887) & (!g888) & (!g147) & (!g148)) + ((g885) & (!g886) & (!g887) & (g888) & (!g147) & (!g148)) + ((g885) & (!g886) & (!g887) & (g888) & (g147) & (g148)) + ((g885) & (!g886) & (g887) & (!g888) & (!g147) & (!g148)) + ((g885) & (!g886) & (g887) & (!g888) & (!g147) & (g148)) + ((g885) & (!g886) & (g887) & (g888) & (!g147) & (!g148)) + ((g885) & (!g886) & (g887) & (g888) & (!g147) & (g148)) + ((g885) & (!g886) & (g887) & (g888) & (g147) & (g148)) + ((g885) & (g886) & (!g887) & (!g888) & (!g147) & (!g148)) + ((g885) & (g886) & (!g887) & (!g888) & (g147) & (!g148)) + ((g885) & (g886) & (!g887) & (g888) & (!g147) & (!g148)) + ((g885) & (g886) & (!g887) & (g888) & (g147) & (!g148)) + ((g885) & (g886) & (!g887) & (g888) & (g147) & (g148)) + ((g885) & (g886) & (g887) & (!g888) & (!g147) & (!g148)) + ((g885) & (g886) & (g887) & (!g888) & (!g147) & (g148)) + ((g885) & (g886) & (g887) & (!g888) & (g147) & (!g148)) + ((g885) & (g886) & (g887) & (g888) & (!g147) & (!g148)) + ((g885) & (g886) & (g887) & (g888) & (!g147) & (g148)) + ((g885) & (g886) & (g887) & (g888) & (g147) & (!g148)) + ((g885) & (g886) & (g887) & (g888) & (g147) & (g148)));
	assign g890 = (((!g874) & (!g879) & (!g884) & (g889) & (g165) & (g166)) + ((!g874) & (!g879) & (g884) & (!g889) & (!g165) & (g166)) + ((!g874) & (!g879) & (g884) & (g889) & (!g165) & (g166)) + ((!g874) & (!g879) & (g884) & (g889) & (g165) & (g166)) + ((!g874) & (g879) & (!g884) & (!g889) & (g165) & (!g166)) + ((!g874) & (g879) & (!g884) & (g889) & (g165) & (!g166)) + ((!g874) & (g879) & (!g884) & (g889) & (g165) & (g166)) + ((!g874) & (g879) & (g884) & (!g889) & (!g165) & (g166)) + ((!g874) & (g879) & (g884) & (!g889) & (g165) & (!g166)) + ((!g874) & (g879) & (g884) & (g889) & (!g165) & (g166)) + ((!g874) & (g879) & (g884) & (g889) & (g165) & (!g166)) + ((!g874) & (g879) & (g884) & (g889) & (g165) & (g166)) + ((g874) & (!g879) & (!g884) & (!g889) & (!g165) & (!g166)) + ((g874) & (!g879) & (!g884) & (g889) & (!g165) & (!g166)) + ((g874) & (!g879) & (!g884) & (g889) & (g165) & (g166)) + ((g874) & (!g879) & (g884) & (!g889) & (!g165) & (!g166)) + ((g874) & (!g879) & (g884) & (!g889) & (!g165) & (g166)) + ((g874) & (!g879) & (g884) & (g889) & (!g165) & (!g166)) + ((g874) & (!g879) & (g884) & (g889) & (!g165) & (g166)) + ((g874) & (!g879) & (g884) & (g889) & (g165) & (g166)) + ((g874) & (g879) & (!g884) & (!g889) & (!g165) & (!g166)) + ((g874) & (g879) & (!g884) & (!g889) & (g165) & (!g166)) + ((g874) & (g879) & (!g884) & (g889) & (!g165) & (!g166)) + ((g874) & (g879) & (!g884) & (g889) & (g165) & (!g166)) + ((g874) & (g879) & (!g884) & (g889) & (g165) & (g166)) + ((g874) & (g879) & (g884) & (!g889) & (!g165) & (!g166)) + ((g874) & (g879) & (g884) & (!g889) & (!g165) & (g166)) + ((g874) & (g879) & (g884) & (!g889) & (g165) & (!g166)) + ((g874) & (g879) & (g884) & (g889) & (!g165) & (!g166)) + ((g874) & (g879) & (g884) & (g889) & (!g165) & (g166)) + ((g874) & (g879) & (g884) & (g889) & (g165) & (!g166)) + ((g874) & (g879) & (g884) & (g889) & (g165) & (g166)));
	assign g4522 = (((!g2173) & (!sk[61]) & (!g3539) & (g891)) + ((!g2173) & (!sk[61]) & (g3539) & (!g891)) + ((!g2173) & (!sk[61]) & (g3539) & (g891)) + ((!g2173) & (sk[61]) & (!g3539) & (g891)) + ((!g2173) & (sk[61]) & (g3539) & (g891)) + ((g2173) & (!sk[61]) & (!g3539) & (g891)) + ((g2173) & (!sk[61]) & (g3539) & (!g891)) + ((g2173) & (!sk[61]) & (g3539) & (g891)) + ((g2173) & (sk[61]) & (g3539) & (!g891)) + ((g2173) & (sk[61]) & (g3539) & (g891)));
	assign g4523 = (((!g2174) & (!g3539) & (!sk[62]) & (g892)) + ((!g2174) & (!g3539) & (sk[62]) & (g892)) + ((!g2174) & (g3539) & (!sk[62]) & (!g892)) + ((!g2174) & (g3539) & (!sk[62]) & (g892)) + ((!g2174) & (g3539) & (sk[62]) & (g892)) + ((g2174) & (!g3539) & (!sk[62]) & (g892)) + ((g2174) & (g3539) & (!sk[62]) & (!g892)) + ((g2174) & (g3539) & (!sk[62]) & (g892)) + ((g2174) & (g3539) & (sk[62]) & (!g892)) + ((g2174) & (g3539) & (sk[62]) & (g892)));
	assign g4524 = (((!g2175) & (!sk[63]) & (!g3539) & (g893)) + ((!g2175) & (!sk[63]) & (g3539) & (!g893)) + ((!g2175) & (!sk[63]) & (g3539) & (g893)) + ((!g2175) & (sk[63]) & (!g3539) & (g893)) + ((!g2175) & (sk[63]) & (g3539) & (g893)) + ((g2175) & (!sk[63]) & (!g3539) & (g893)) + ((g2175) & (!sk[63]) & (g3539) & (!g893)) + ((g2175) & (!sk[63]) & (g3539) & (g893)) + ((g2175) & (sk[63]) & (g3539) & (!g893)) + ((g2175) & (sk[63]) & (g3539) & (g893)));
	assign g4525 = (((!g2176) & (!sk[64]) & (!g3539) & (g894)) + ((!g2176) & (!sk[64]) & (g3539) & (!g894)) + ((!g2176) & (!sk[64]) & (g3539) & (g894)) + ((!g2176) & (sk[64]) & (!g3539) & (g894)) + ((!g2176) & (sk[64]) & (g3539) & (g894)) + ((g2176) & (!sk[64]) & (!g3539) & (g894)) + ((g2176) & (!sk[64]) & (g3539) & (!g894)) + ((g2176) & (!sk[64]) & (g3539) & (g894)) + ((g2176) & (sk[64]) & (g3539) & (!g894)) + ((g2176) & (sk[64]) & (g3539) & (g894)));
	assign g895 = (((!g891) & (!g892) & (!g893) & (g894) & (g165) & (g166)) + ((!g891) & (!g892) & (g893) & (!g894) & (!g165) & (g166)) + ((!g891) & (!g892) & (g893) & (g894) & (!g165) & (g166)) + ((!g891) & (!g892) & (g893) & (g894) & (g165) & (g166)) + ((!g891) & (g892) & (!g893) & (!g894) & (g165) & (!g166)) + ((!g891) & (g892) & (!g893) & (g894) & (g165) & (!g166)) + ((!g891) & (g892) & (!g893) & (g894) & (g165) & (g166)) + ((!g891) & (g892) & (g893) & (!g894) & (!g165) & (g166)) + ((!g891) & (g892) & (g893) & (!g894) & (g165) & (!g166)) + ((!g891) & (g892) & (g893) & (g894) & (!g165) & (g166)) + ((!g891) & (g892) & (g893) & (g894) & (g165) & (!g166)) + ((!g891) & (g892) & (g893) & (g894) & (g165) & (g166)) + ((g891) & (!g892) & (!g893) & (!g894) & (!g165) & (!g166)) + ((g891) & (!g892) & (!g893) & (g894) & (!g165) & (!g166)) + ((g891) & (!g892) & (!g893) & (g894) & (g165) & (g166)) + ((g891) & (!g892) & (g893) & (!g894) & (!g165) & (!g166)) + ((g891) & (!g892) & (g893) & (!g894) & (!g165) & (g166)) + ((g891) & (!g892) & (g893) & (g894) & (!g165) & (!g166)) + ((g891) & (!g892) & (g893) & (g894) & (!g165) & (g166)) + ((g891) & (!g892) & (g893) & (g894) & (g165) & (g166)) + ((g891) & (g892) & (!g893) & (!g894) & (!g165) & (!g166)) + ((g891) & (g892) & (!g893) & (!g894) & (g165) & (!g166)) + ((g891) & (g892) & (!g893) & (g894) & (!g165) & (!g166)) + ((g891) & (g892) & (!g893) & (g894) & (g165) & (!g166)) + ((g891) & (g892) & (!g893) & (g894) & (g165) & (g166)) + ((g891) & (g892) & (g893) & (!g894) & (!g165) & (!g166)) + ((g891) & (g892) & (g893) & (!g894) & (!g165) & (g166)) + ((g891) & (g892) & (g893) & (!g894) & (g165) & (!g166)) + ((g891) & (g892) & (g893) & (g894) & (!g165) & (!g166)) + ((g891) & (g892) & (g893) & (g894) & (!g165) & (g166)) + ((g891) & (g892) & (g893) & (g894) & (g165) & (!g166)) + ((g891) & (g892) & (g893) & (g894) & (g165) & (g166)));
	assign g4526 = (((!sk[66]) & (!g2177) & (!g3539) & (g896)) + ((!sk[66]) & (!g2177) & (g3539) & (!g896)) + ((!sk[66]) & (!g2177) & (g3539) & (g896)) + ((!sk[66]) & (g2177) & (!g3539) & (g896)) + ((!sk[66]) & (g2177) & (g3539) & (!g896)) + ((!sk[66]) & (g2177) & (g3539) & (g896)) + ((sk[66]) & (!g2177) & (!g3539) & (g896)) + ((sk[66]) & (!g2177) & (g3539) & (g896)) + ((sk[66]) & (g2177) & (g3539) & (!g896)) + ((sk[66]) & (g2177) & (g3539) & (g896)));
	assign g4527 = (((!sk[67]) & (!g2178) & (!g3539) & (g897)) + ((!sk[67]) & (!g2178) & (g3539) & (!g897)) + ((!sk[67]) & (!g2178) & (g3539) & (g897)) + ((!sk[67]) & (g2178) & (!g3539) & (g897)) + ((!sk[67]) & (g2178) & (g3539) & (!g897)) + ((!sk[67]) & (g2178) & (g3539) & (g897)) + ((sk[67]) & (!g2178) & (!g3539) & (g897)) + ((sk[67]) & (!g2178) & (g3539) & (g897)) + ((sk[67]) & (g2178) & (g3539) & (!g897)) + ((sk[67]) & (g2178) & (g3539) & (g897)));
	assign g4528 = (((!sk[68]) & (!g2179) & (!g3539) & (g898)) + ((!sk[68]) & (!g2179) & (g3539) & (!g898)) + ((!sk[68]) & (!g2179) & (g3539) & (g898)) + ((!sk[68]) & (g2179) & (!g3539) & (g898)) + ((!sk[68]) & (g2179) & (g3539) & (!g898)) + ((!sk[68]) & (g2179) & (g3539) & (g898)) + ((sk[68]) & (!g2179) & (!g3539) & (g898)) + ((sk[68]) & (!g2179) & (g3539) & (g898)) + ((sk[68]) & (g2179) & (g3539) & (!g898)) + ((sk[68]) & (g2179) & (g3539) & (g898)));
	assign g899 = (((!g165) & (!g166) & (!g896) & (g897) & (!sk[69]) & (!g898)) + ((!g165) & (!g166) & (!g896) & (g897) & (!sk[69]) & (g898)) + ((!g165) & (!g166) & (g896) & (!g897) & (!sk[69]) & (!g898)) + ((!g165) & (!g166) & (g896) & (!g897) & (!sk[69]) & (g898)) + ((!g165) & (!g166) & (g896) & (g897) & (!sk[69]) & (!g898)) + ((!g165) & (!g166) & (g896) & (g897) & (!sk[69]) & (g898)) + ((!g165) & (g166) & (!g896) & (!g897) & (!sk[69]) & (!g898)) + ((!g165) & (g166) & (!g896) & (!g897) & (!sk[69]) & (g898)) + ((!g165) & (g166) & (!g896) & (!g897) & (sk[69]) & (g898)) + ((!g165) & (g166) & (!g896) & (g897) & (!sk[69]) & (!g898)) + ((!g165) & (g166) & (!g896) & (g897) & (!sk[69]) & (g898)) + ((!g165) & (g166) & (!g896) & (g897) & (sk[69]) & (g898)) + ((!g165) & (g166) & (g896) & (!g897) & (!sk[69]) & (!g898)) + ((!g165) & (g166) & (g896) & (!g897) & (!sk[69]) & (g898)) + ((!g165) & (g166) & (g896) & (!g897) & (sk[69]) & (g898)) + ((!g165) & (g166) & (g896) & (g897) & (!sk[69]) & (!g898)) + ((!g165) & (g166) & (g896) & (g897) & (!sk[69]) & (g898)) + ((!g165) & (g166) & (g896) & (g897) & (sk[69]) & (g898)) + ((g165) & (!g166) & (!g896) & (g897) & (!sk[69]) & (!g898)) + ((g165) & (!g166) & (!g896) & (g897) & (!sk[69]) & (g898)) + ((g165) & (!g166) & (g896) & (!g897) & (!sk[69]) & (!g898)) + ((g165) & (!g166) & (g896) & (!g897) & (!sk[69]) & (g898)) + ((g165) & (!g166) & (g896) & (!g897) & (sk[69]) & (!g898)) + ((g165) & (!g166) & (g896) & (!g897) & (sk[69]) & (g898)) + ((g165) & (!g166) & (g896) & (g897) & (!sk[69]) & (!g898)) + ((g165) & (!g166) & (g896) & (g897) & (!sk[69]) & (g898)) + ((g165) & (!g166) & (g896) & (g897) & (sk[69]) & (!g898)) + ((g165) & (!g166) & (g896) & (g897) & (sk[69]) & (g898)) + ((g165) & (g166) & (!g896) & (!g897) & (!sk[69]) & (!g898)) + ((g165) & (g166) & (!g896) & (!g897) & (!sk[69]) & (g898)) + ((g165) & (g166) & (!g896) & (g897) & (!sk[69]) & (!g898)) + ((g165) & (g166) & (!g896) & (g897) & (!sk[69]) & (g898)) + ((g165) & (g166) & (!g896) & (g897) & (sk[69]) & (!g898)) + ((g165) & (g166) & (!g896) & (g897) & (sk[69]) & (g898)) + ((g165) & (g166) & (g896) & (!g897) & (!sk[69]) & (!g898)) + ((g165) & (g166) & (g896) & (!g897) & (!sk[69]) & (g898)) + ((g165) & (g166) & (g896) & (g897) & (!sk[69]) & (!g898)) + ((g165) & (g166) & (g896) & (g897) & (!sk[69]) & (g898)) + ((g165) & (g166) & (g896) & (g897) & (sk[69]) & (!g898)) + ((g165) & (g166) & (g896) & (g897) & (sk[69]) & (g898)));
	assign g4529 = (((!sk[70]) & (!g2162) & (!g3539) & (g900)) + ((!sk[70]) & (!g2162) & (g3539) & (!g900)) + ((!sk[70]) & (!g2162) & (g3539) & (g900)) + ((!sk[70]) & (g2162) & (!g3539) & (g900)) + ((!sk[70]) & (g2162) & (g3539) & (!g900)) + ((!sk[70]) & (g2162) & (g3539) & (g900)) + ((sk[70]) & (!g2162) & (!g3539) & (g900)) + ((sk[70]) & (!g2162) & (g3539) & (g900)) + ((sk[70]) & (g2162) & (g3539) & (!g900)) + ((sk[70]) & (g2162) & (g3539) & (g900)));
	assign g4530 = (((!sk[71]) & (!g2164) & (!g3539) & (g901)) + ((!sk[71]) & (!g2164) & (g3539) & (!g901)) + ((!sk[71]) & (!g2164) & (g3539) & (g901)) + ((!sk[71]) & (g2164) & (!g3539) & (g901)) + ((!sk[71]) & (g2164) & (g3539) & (!g901)) + ((!sk[71]) & (g2164) & (g3539) & (g901)) + ((sk[71]) & (!g2164) & (!g3539) & (g901)) + ((sk[71]) & (!g2164) & (g3539) & (g901)) + ((sk[71]) & (g2164) & (g3539) & (!g901)) + ((sk[71]) & (g2164) & (g3539) & (g901)));
	assign g4531 = (((!g2166) & (!g3539) & (!sk[72]) & (g902)) + ((!g2166) & (!g3539) & (sk[72]) & (g902)) + ((!g2166) & (g3539) & (!sk[72]) & (!g902)) + ((!g2166) & (g3539) & (!sk[72]) & (g902)) + ((!g2166) & (g3539) & (sk[72]) & (g902)) + ((g2166) & (!g3539) & (!sk[72]) & (g902)) + ((g2166) & (g3539) & (!sk[72]) & (!g902)) + ((g2166) & (g3539) & (!sk[72]) & (g902)) + ((g2166) & (g3539) & (sk[72]) & (!g902)) + ((g2166) & (g3539) & (sk[72]) & (g902)));
	assign g4532 = (((!sk[73]) & (!g2168) & (!g3539) & (g903)) + ((!sk[73]) & (!g2168) & (g3539) & (!g903)) + ((!sk[73]) & (!g2168) & (g3539) & (g903)) + ((!sk[73]) & (g2168) & (!g3539) & (g903)) + ((!sk[73]) & (g2168) & (g3539) & (!g903)) + ((!sk[73]) & (g2168) & (g3539) & (g903)) + ((sk[73]) & (!g2168) & (!g3539) & (g903)) + ((sk[73]) & (!g2168) & (g3539) & (g903)) + ((sk[73]) & (g2168) & (g3539) & (!g903)) + ((sk[73]) & (g2168) & (g3539) & (g903)));
	assign g904 = (((!g900) & (!g901) & (!g902) & (g903) & (g165) & (g166)) + ((!g900) & (!g901) & (g902) & (!g903) & (!g165) & (g166)) + ((!g900) & (!g901) & (g902) & (g903) & (!g165) & (g166)) + ((!g900) & (!g901) & (g902) & (g903) & (g165) & (g166)) + ((!g900) & (g901) & (!g902) & (!g903) & (g165) & (!g166)) + ((!g900) & (g901) & (!g902) & (g903) & (g165) & (!g166)) + ((!g900) & (g901) & (!g902) & (g903) & (g165) & (g166)) + ((!g900) & (g901) & (g902) & (!g903) & (!g165) & (g166)) + ((!g900) & (g901) & (g902) & (!g903) & (g165) & (!g166)) + ((!g900) & (g901) & (g902) & (g903) & (!g165) & (g166)) + ((!g900) & (g901) & (g902) & (g903) & (g165) & (!g166)) + ((!g900) & (g901) & (g902) & (g903) & (g165) & (g166)) + ((g900) & (!g901) & (!g902) & (!g903) & (!g165) & (!g166)) + ((g900) & (!g901) & (!g902) & (g903) & (!g165) & (!g166)) + ((g900) & (!g901) & (!g902) & (g903) & (g165) & (g166)) + ((g900) & (!g901) & (g902) & (!g903) & (!g165) & (!g166)) + ((g900) & (!g901) & (g902) & (!g903) & (!g165) & (g166)) + ((g900) & (!g901) & (g902) & (g903) & (!g165) & (!g166)) + ((g900) & (!g901) & (g902) & (g903) & (!g165) & (g166)) + ((g900) & (!g901) & (g902) & (g903) & (g165) & (g166)) + ((g900) & (g901) & (!g902) & (!g903) & (!g165) & (!g166)) + ((g900) & (g901) & (!g902) & (!g903) & (g165) & (!g166)) + ((g900) & (g901) & (!g902) & (g903) & (!g165) & (!g166)) + ((g900) & (g901) & (!g902) & (g903) & (g165) & (!g166)) + ((g900) & (g901) & (!g902) & (g903) & (g165) & (g166)) + ((g900) & (g901) & (g902) & (!g903) & (!g165) & (!g166)) + ((g900) & (g901) & (g902) & (!g903) & (!g165) & (g166)) + ((g900) & (g901) & (g902) & (!g903) & (g165) & (!g166)) + ((g900) & (g901) & (g902) & (g903) & (!g165) & (!g166)) + ((g900) & (g901) & (g902) & (g903) & (!g165) & (g166)) + ((g900) & (g901) & (g902) & (g903) & (g165) & (!g166)) + ((g900) & (g901) & (g902) & (g903) & (g165) & (g166)));
	assign g4533 = (((!g2169) & (!sk[75]) & (!g3539) & (g905)) + ((!g2169) & (!sk[75]) & (g3539) & (!g905)) + ((!g2169) & (!sk[75]) & (g3539) & (g905)) + ((!g2169) & (sk[75]) & (!g3539) & (g905)) + ((!g2169) & (sk[75]) & (g3539) & (g905)) + ((g2169) & (!sk[75]) & (!g3539) & (g905)) + ((g2169) & (!sk[75]) & (g3539) & (!g905)) + ((g2169) & (!sk[75]) & (g3539) & (g905)) + ((g2169) & (sk[75]) & (g3539) & (!g905)) + ((g2169) & (sk[75]) & (g3539) & (g905)));
	assign g4534 = (((!g2170) & (!sk[76]) & (!g3539) & (g906)) + ((!g2170) & (!sk[76]) & (g3539) & (!g906)) + ((!g2170) & (!sk[76]) & (g3539) & (g906)) + ((!g2170) & (sk[76]) & (!g3539) & (g906)) + ((!g2170) & (sk[76]) & (g3539) & (g906)) + ((g2170) & (!sk[76]) & (!g3539) & (g906)) + ((g2170) & (!sk[76]) & (g3539) & (!g906)) + ((g2170) & (!sk[76]) & (g3539) & (g906)) + ((g2170) & (sk[76]) & (g3539) & (!g906)) + ((g2170) & (sk[76]) & (g3539) & (g906)));
	assign g4535 = (((!sk[77]) & (!g2171) & (!g3539) & (g907)) + ((!sk[77]) & (!g2171) & (g3539) & (!g907)) + ((!sk[77]) & (!g2171) & (g3539) & (g907)) + ((!sk[77]) & (g2171) & (!g3539) & (g907)) + ((!sk[77]) & (g2171) & (g3539) & (!g907)) + ((!sk[77]) & (g2171) & (g3539) & (g907)) + ((sk[77]) & (!g2171) & (!g3539) & (g907)) + ((sk[77]) & (!g2171) & (g3539) & (g907)) + ((sk[77]) & (g2171) & (g3539) & (!g907)) + ((sk[77]) & (g2171) & (g3539) & (g907)));
	assign g4536 = (((!g2172) & (!sk[78]) & (!g3539) & (g908)) + ((!g2172) & (!sk[78]) & (g3539) & (!g908)) + ((!g2172) & (!sk[78]) & (g3539) & (g908)) + ((!g2172) & (sk[78]) & (!g3539) & (g908)) + ((!g2172) & (sk[78]) & (g3539) & (g908)) + ((g2172) & (!sk[78]) & (!g3539) & (g908)) + ((g2172) & (!sk[78]) & (g3539) & (!g908)) + ((g2172) & (!sk[78]) & (g3539) & (g908)) + ((g2172) & (sk[78]) & (g3539) & (!g908)) + ((g2172) & (sk[78]) & (g3539) & (g908)));
	assign g909 = (((!g905) & (!g906) & (!g907) & (g908) & (g165) & (g166)) + ((!g905) & (!g906) & (g907) & (!g908) & (!g165) & (g166)) + ((!g905) & (!g906) & (g907) & (g908) & (!g165) & (g166)) + ((!g905) & (!g906) & (g907) & (g908) & (g165) & (g166)) + ((!g905) & (g906) & (!g907) & (!g908) & (g165) & (!g166)) + ((!g905) & (g906) & (!g907) & (g908) & (g165) & (!g166)) + ((!g905) & (g906) & (!g907) & (g908) & (g165) & (g166)) + ((!g905) & (g906) & (g907) & (!g908) & (!g165) & (g166)) + ((!g905) & (g906) & (g907) & (!g908) & (g165) & (!g166)) + ((!g905) & (g906) & (g907) & (g908) & (!g165) & (g166)) + ((!g905) & (g906) & (g907) & (g908) & (g165) & (!g166)) + ((!g905) & (g906) & (g907) & (g908) & (g165) & (g166)) + ((g905) & (!g906) & (!g907) & (!g908) & (!g165) & (!g166)) + ((g905) & (!g906) & (!g907) & (g908) & (!g165) & (!g166)) + ((g905) & (!g906) & (!g907) & (g908) & (g165) & (g166)) + ((g905) & (!g906) & (g907) & (!g908) & (!g165) & (!g166)) + ((g905) & (!g906) & (g907) & (!g908) & (!g165) & (g166)) + ((g905) & (!g906) & (g907) & (g908) & (!g165) & (!g166)) + ((g905) & (!g906) & (g907) & (g908) & (!g165) & (g166)) + ((g905) & (!g906) & (g907) & (g908) & (g165) & (g166)) + ((g905) & (g906) & (!g907) & (!g908) & (!g165) & (!g166)) + ((g905) & (g906) & (!g907) & (!g908) & (g165) & (!g166)) + ((g905) & (g906) & (!g907) & (g908) & (!g165) & (!g166)) + ((g905) & (g906) & (!g907) & (g908) & (g165) & (!g166)) + ((g905) & (g906) & (!g907) & (g908) & (g165) & (g166)) + ((g905) & (g906) & (g907) & (!g908) & (!g165) & (!g166)) + ((g905) & (g906) & (g907) & (!g908) & (!g165) & (g166)) + ((g905) & (g906) & (g907) & (!g908) & (g165) & (!g166)) + ((g905) & (g906) & (g907) & (g908) & (!g165) & (!g166)) + ((g905) & (g906) & (g907) & (g908) & (!g165) & (g166)) + ((g905) & (g906) & (g907) & (g908) & (g165) & (!g166)) + ((g905) & (g906) & (g907) & (g908) & (g165) & (g166)));
	assign g910 = (((!g147) & (!g148) & (!g895) & (g899) & (!g904) & (!g909)) + ((!g147) & (!g148) & (!g895) & (g899) & (!g904) & (g909)) + ((!g147) & (!g148) & (!g895) & (g899) & (g904) & (!g909)) + ((!g147) & (!g148) & (!g895) & (g899) & (g904) & (g909)) + ((!g147) & (!g148) & (g895) & (g899) & (!g904) & (!g909)) + ((!g147) & (!g148) & (g895) & (g899) & (!g904) & (g909)) + ((!g147) & (!g148) & (g895) & (g899) & (g904) & (!g909)) + ((!g147) & (!g148) & (g895) & (g899) & (g904) & (g909)) + ((!g147) & (g148) & (!g895) & (!g899) & (!g904) & (g909)) + ((!g147) & (g148) & (!g895) & (!g899) & (g904) & (g909)) + ((!g147) & (g148) & (!g895) & (g899) & (!g904) & (g909)) + ((!g147) & (g148) & (!g895) & (g899) & (g904) & (g909)) + ((!g147) & (g148) & (g895) & (!g899) & (!g904) & (g909)) + ((!g147) & (g148) & (g895) & (!g899) & (g904) & (g909)) + ((!g147) & (g148) & (g895) & (g899) & (!g904) & (g909)) + ((!g147) & (g148) & (g895) & (g899) & (g904) & (g909)) + ((g147) & (!g148) & (g895) & (!g899) & (!g904) & (!g909)) + ((g147) & (!g148) & (g895) & (!g899) & (!g904) & (g909)) + ((g147) & (!g148) & (g895) & (!g899) & (g904) & (!g909)) + ((g147) & (!g148) & (g895) & (!g899) & (g904) & (g909)) + ((g147) & (!g148) & (g895) & (g899) & (!g904) & (!g909)) + ((g147) & (!g148) & (g895) & (g899) & (!g904) & (g909)) + ((g147) & (!g148) & (g895) & (g899) & (g904) & (!g909)) + ((g147) & (!g148) & (g895) & (g899) & (g904) & (g909)) + ((g147) & (g148) & (!g895) & (!g899) & (g904) & (!g909)) + ((g147) & (g148) & (!g895) & (!g899) & (g904) & (g909)) + ((g147) & (g148) & (!g895) & (g899) & (g904) & (!g909)) + ((g147) & (g148) & (!g895) & (g899) & (g904) & (g909)) + ((g147) & (g148) & (g895) & (!g899) & (g904) & (!g909)) + ((g147) & (g148) & (g895) & (!g899) & (g904) & (g909)) + ((g147) & (g148) & (g895) & (g899) & (g904) & (!g909)) + ((g147) & (g148) & (g895) & (g899) & (g904) & (g909)));
	assign g911 = (((!g142) & (!sk[81]) & (!g890) & (g910)) + ((!g142) & (!sk[81]) & (g890) & (!g910)) + ((!g142) & (!sk[81]) & (g890) & (g910)) + ((!g142) & (sk[81]) & (!g890) & (g910)) + ((!g142) & (sk[81]) & (g890) & (g910)) + ((g142) & (!sk[81]) & (!g890) & (g910)) + ((g142) & (!sk[81]) & (g890) & (!g910)) + ((g142) & (!sk[81]) & (g890) & (g910)) + ((g142) & (sk[81]) & (g890) & (!g910)) + ((g142) & (sk[81]) & (g890) & (g910)));
	assign g4537 = (((!sk[82]) & (!g2059) & (!g2569) & (g912)) + ((!sk[82]) & (!g2059) & (g2569) & (!g912)) + ((!sk[82]) & (!g2059) & (g2569) & (g912)) + ((!sk[82]) & (g2059) & (!g2569) & (g912)) + ((!sk[82]) & (g2059) & (g2569) & (!g912)) + ((!sk[82]) & (g2059) & (g2569) & (g912)) + ((sk[82]) & (!g2059) & (!g2569) & (g912)) + ((sk[82]) & (!g2059) & (g2569) & (g912)) + ((sk[82]) & (g2059) & (g2569) & (!g912)) + ((sk[82]) & (g2059) & (g2569) & (g912)));
	assign g913 = (((!g672) & (!g674) & (!g675) & (!g680) & (!g3134) & (g3135)) + ((!g672) & (!g674) & (!g675) & (g680) & (!g3134) & (g3135)) + ((!g672) & (!g674) & (g675) & (!g680) & (!g3134) & (g3135)) + ((!g672) & (!g674) & (g675) & (!g680) & (g3134) & (g3135)) + ((!g672) & (!g674) & (g675) & (g680) & (!g3134) & (g3135)) + ((!g672) & (g674) & (!g675) & (!g680) & (!g3134) & (g3135)) + ((!g672) & (g674) & (!g675) & (!g680) & (g3134) & (g3135)) + ((!g672) & (g674) & (!g675) & (g680) & (!g3134) & (g3135)) + ((!g672) & (g674) & (g675) & (!g680) & (!g3134) & (g3135)) + ((!g672) & (g674) & (g675) & (!g680) & (g3134) & (g3135)) + ((!g672) & (g674) & (g675) & (g680) & (!g3134) & (g3135)) + ((g672) & (!g674) & (!g675) & (!g680) & (!g3134) & (g3135)) + ((g672) & (!g674) & (!g675) & (!g680) & (g3134) & (g3135)) + ((g672) & (!g674) & (!g675) & (g680) & (!g3134) & (g3135)) + ((g672) & (!g674) & (g675) & (!g680) & (!g3134) & (g3135)) + ((g672) & (!g674) & (g675) & (!g680) & (g3134) & (g3135)) + ((g672) & (!g674) & (g675) & (g680) & (!g3134) & (g3135)) + ((g672) & (!g674) & (g675) & (g680) & (g3134) & (g3135)) + ((g672) & (g674) & (!g675) & (!g680) & (!g3134) & (g3135)) + ((g672) & (g674) & (!g675) & (!g680) & (g3134) & (g3135)) + ((g672) & (g674) & (!g675) & (g680) & (!g3134) & (g3135)) + ((g672) & (g674) & (!g675) & (g680) & (g3134) & (g3135)) + ((g672) & (g674) & (g675) & (!g680) & (!g3134) & (g3135)) + ((g672) & (g674) & (g675) & (!g680) & (g3134) & (g3135)) + ((g672) & (g674) & (g675) & (g680) & (!g3134) & (g3135)) + ((g672) & (g674) & (g675) & (g680) & (g3134) & (g3135)));
	assign g914 = (((g864) & (!sk[84]) & (!g868)) + ((g864) & (!sk[84]) & (g868)) + ((g864) & (sk[84]) & (!g868)));
	assign g915 = (((!g913) & (sk[85]) & (!g914)) + ((g913) & (!sk[85]) & (!g914)) + ((g913) & (!sk[85]) & (g914)));
	assign g916 = (((!g867) & (!g107) & (!sk[86]) & (g679)) + ((!g867) & (!g107) & (sk[86]) & (!g679)) + ((!g867) & (!g107) & (sk[86]) & (g679)) + ((!g867) & (g107) & (!sk[86]) & (!g679)) + ((!g867) & (g107) & (!sk[86]) & (g679)) + ((!g867) & (g107) & (sk[86]) & (g679)) + ((g867) & (!g107) & (!sk[86]) & (g679)) + ((g867) & (!g107) & (sk[86]) & (!g679)) + ((g867) & (g107) & (!sk[86]) & (!g679)) + ((g867) & (g107) & (!sk[86]) & (g679)));
	assign g917 = (((!g126) & (!sk[87]) & (!g911) & (!g912) & (g915) & (!g916)) + ((!g126) & (!sk[87]) & (!g911) & (!g912) & (g915) & (g916)) + ((!g126) & (!sk[87]) & (!g911) & (g912) & (!g915) & (!g916)) + ((!g126) & (!sk[87]) & (!g911) & (g912) & (!g915) & (g916)) + ((!g126) & (!sk[87]) & (!g911) & (g912) & (g915) & (!g916)) + ((!g126) & (!sk[87]) & (!g911) & (g912) & (g915) & (g916)) + ((!g126) & (!sk[87]) & (g911) & (!g912) & (!g915) & (!g916)) + ((!g126) & (!sk[87]) & (g911) & (!g912) & (!g915) & (g916)) + ((!g126) & (!sk[87]) & (g911) & (!g912) & (g915) & (!g916)) + ((!g126) & (!sk[87]) & (g911) & (!g912) & (g915) & (g916)) + ((!g126) & (!sk[87]) & (g911) & (g912) & (!g915) & (!g916)) + ((!g126) & (!sk[87]) & (g911) & (g912) & (!g915) & (g916)) + ((!g126) & (!sk[87]) & (g911) & (g912) & (g915) & (!g916)) + ((!g126) & (!sk[87]) & (g911) & (g912) & (g915) & (g916)) + ((!g126) & (sk[87]) & (!g911) & (g912) & (!g915) & (!g916)) + ((!g126) & (sk[87]) & (!g911) & (g912) & (!g915) & (g916)) + ((!g126) & (sk[87]) & (!g911) & (g912) & (g915) & (!g916)) + ((!g126) & (sk[87]) & (!g911) & (g912) & (g915) & (g916)) + ((!g126) & (sk[87]) & (g911) & (g912) & (!g915) & (!g916)) + ((!g126) & (sk[87]) & (g911) & (g912) & (!g915) & (g916)) + ((!g126) & (sk[87]) & (g911) & (g912) & (g915) & (!g916)) + ((!g126) & (sk[87]) & (g911) & (g912) & (g915) & (g916)) + ((g126) & (!sk[87]) & (!g911) & (!g912) & (g915) & (!g916)) + ((g126) & (!sk[87]) & (!g911) & (!g912) & (g915) & (g916)) + ((g126) & (!sk[87]) & (!g911) & (g912) & (!g915) & (!g916)) + ((g126) & (!sk[87]) & (!g911) & (g912) & (!g915) & (g916)) + ((g126) & (!sk[87]) & (!g911) & (g912) & (g915) & (!g916)) + ((g126) & (!sk[87]) & (!g911) & (g912) & (g915) & (g916)) + ((g126) & (!sk[87]) & (g911) & (!g912) & (!g915) & (!g916)) + ((g126) & (!sk[87]) & (g911) & (!g912) & (!g915) & (g916)) + ((g126) & (!sk[87]) & (g911) & (!g912) & (g915) & (!g916)) + ((g126) & (!sk[87]) & (g911) & (!g912) & (g915) & (g916)) + ((g126) & (!sk[87]) & (g911) & (g912) & (!g915) & (!g916)) + ((g126) & (!sk[87]) & (g911) & (g912) & (!g915) & (g916)) + ((g126) & (!sk[87]) & (g911) & (g912) & (g915) & (!g916)) + ((g126) & (!sk[87]) & (g911) & (g912) & (g915) & (g916)) + ((g126) & (sk[87]) & (!g911) & (!g912) & (!g915) & (g916)) + ((g126) & (sk[87]) & (!g911) & (!g912) & (g915) & (!g916)) + ((g126) & (sk[87]) & (!g911) & (g912) & (!g915) & (g916)) + ((g126) & (sk[87]) & (!g911) & (g912) & (g915) & (!g916)) + ((g126) & (sk[87]) & (g911) & (!g912) & (!g915) & (!g916)) + ((g126) & (sk[87]) & (g911) & (!g912) & (g915) & (g916)) + ((g126) & (sk[87]) & (g911) & (g912) & (!g915) & (!g916)) + ((g126) & (sk[87]) & (g911) & (g912) & (g915) & (g916)));
	assign g4538 = (((!g2140) & (!sk[88]) & (!g3515) & (g918)) + ((!g2140) & (!sk[88]) & (g3515) & (!g918)) + ((!g2140) & (!sk[88]) & (g3515) & (g918)) + ((!g2140) & (sk[88]) & (!g3515) & (g918)) + ((!g2140) & (sk[88]) & (g3515) & (g918)) + ((g2140) & (!sk[88]) & (!g3515) & (g918)) + ((g2140) & (!sk[88]) & (g3515) & (!g918)) + ((g2140) & (!sk[88]) & (g3515) & (g918)) + ((g2140) & (sk[88]) & (g3515) & (!g918)) + ((g2140) & (sk[88]) & (g3515) & (g918)));
	assign g4539 = (((!g2142) & (!sk[89]) & (!g3515) & (g919)) + ((!g2142) & (!sk[89]) & (g3515) & (!g919)) + ((!g2142) & (!sk[89]) & (g3515) & (g919)) + ((!g2142) & (sk[89]) & (!g3515) & (g919)) + ((!g2142) & (sk[89]) & (g3515) & (g919)) + ((g2142) & (!sk[89]) & (!g3515) & (g919)) + ((g2142) & (!sk[89]) & (g3515) & (!g919)) + ((g2142) & (!sk[89]) & (g3515) & (g919)) + ((g2142) & (sk[89]) & (g3515) & (!g919)) + ((g2142) & (sk[89]) & (g3515) & (g919)));
	assign g4540 = (((!g2144) & (!g3515) & (!sk[90]) & (g920)) + ((!g2144) & (!g3515) & (sk[90]) & (g920)) + ((!g2144) & (g3515) & (!sk[90]) & (!g920)) + ((!g2144) & (g3515) & (!sk[90]) & (g920)) + ((!g2144) & (g3515) & (sk[90]) & (g920)) + ((g2144) & (!g3515) & (!sk[90]) & (g920)) + ((g2144) & (g3515) & (!sk[90]) & (!g920)) + ((g2144) & (g3515) & (!sk[90]) & (g920)) + ((g2144) & (g3515) & (sk[90]) & (!g920)) + ((g2144) & (g3515) & (sk[90]) & (g920)));
	assign g4541 = (((!g2145) & (!sk[91]) & (!g3515) & (g921)) + ((!g2145) & (!sk[91]) & (g3515) & (!g921)) + ((!g2145) & (!sk[91]) & (g3515) & (g921)) + ((!g2145) & (sk[91]) & (!g3515) & (g921)) + ((!g2145) & (sk[91]) & (g3515) & (g921)) + ((g2145) & (!sk[91]) & (!g3515) & (g921)) + ((g2145) & (!sk[91]) & (g3515) & (!g921)) + ((g2145) & (!sk[91]) & (g3515) & (g921)) + ((g2145) & (sk[91]) & (g3515) & (!g921)) + ((g2145) & (sk[91]) & (g3515) & (g921)));
	assign g922 = (((!g918) & (!g919) & (!g920) & (g921) & (g147) & (g148)) + ((!g918) & (!g919) & (g920) & (!g921) & (!g147) & (g148)) + ((!g918) & (!g919) & (g920) & (g921) & (!g147) & (g148)) + ((!g918) & (!g919) & (g920) & (g921) & (g147) & (g148)) + ((!g918) & (g919) & (!g920) & (!g921) & (g147) & (!g148)) + ((!g918) & (g919) & (!g920) & (g921) & (g147) & (!g148)) + ((!g918) & (g919) & (!g920) & (g921) & (g147) & (g148)) + ((!g918) & (g919) & (g920) & (!g921) & (!g147) & (g148)) + ((!g918) & (g919) & (g920) & (!g921) & (g147) & (!g148)) + ((!g918) & (g919) & (g920) & (g921) & (!g147) & (g148)) + ((!g918) & (g919) & (g920) & (g921) & (g147) & (!g148)) + ((!g918) & (g919) & (g920) & (g921) & (g147) & (g148)) + ((g918) & (!g919) & (!g920) & (!g921) & (!g147) & (!g148)) + ((g918) & (!g919) & (!g920) & (g921) & (!g147) & (!g148)) + ((g918) & (!g919) & (!g920) & (g921) & (g147) & (g148)) + ((g918) & (!g919) & (g920) & (!g921) & (!g147) & (!g148)) + ((g918) & (!g919) & (g920) & (!g921) & (!g147) & (g148)) + ((g918) & (!g919) & (g920) & (g921) & (!g147) & (!g148)) + ((g918) & (!g919) & (g920) & (g921) & (!g147) & (g148)) + ((g918) & (!g919) & (g920) & (g921) & (g147) & (g148)) + ((g918) & (g919) & (!g920) & (!g921) & (!g147) & (!g148)) + ((g918) & (g919) & (!g920) & (!g921) & (g147) & (!g148)) + ((g918) & (g919) & (!g920) & (g921) & (!g147) & (!g148)) + ((g918) & (g919) & (!g920) & (g921) & (g147) & (!g148)) + ((g918) & (g919) & (!g920) & (g921) & (g147) & (g148)) + ((g918) & (g919) & (g920) & (!g921) & (!g147) & (!g148)) + ((g918) & (g919) & (g920) & (!g921) & (!g147) & (g148)) + ((g918) & (g919) & (g920) & (!g921) & (g147) & (!g148)) + ((g918) & (g919) & (g920) & (g921) & (!g147) & (!g148)) + ((g918) & (g919) & (g920) & (g921) & (!g147) & (g148)) + ((g918) & (g919) & (g920) & (g921) & (g147) & (!g148)) + ((g918) & (g919) & (g920) & (g921) & (g147) & (g148)));
	assign g4542 = (((!sk[93]) & (!g2146) & (!g3515) & (g923)) + ((!sk[93]) & (!g2146) & (g3515) & (!g923)) + ((!sk[93]) & (!g2146) & (g3515) & (g923)) + ((!sk[93]) & (g2146) & (!g3515) & (g923)) + ((!sk[93]) & (g2146) & (g3515) & (!g923)) + ((!sk[93]) & (g2146) & (g3515) & (g923)) + ((sk[93]) & (!g2146) & (!g3515) & (g923)) + ((sk[93]) & (!g2146) & (g3515) & (g923)) + ((sk[93]) & (g2146) & (g3515) & (!g923)) + ((sk[93]) & (g2146) & (g3515) & (g923)));
	assign g4543 = (((!sk[94]) & (!g2148) & (!g3515) & (g924)) + ((!sk[94]) & (!g2148) & (g3515) & (!g924)) + ((!sk[94]) & (!g2148) & (g3515) & (g924)) + ((!sk[94]) & (g2148) & (!g3515) & (g924)) + ((!sk[94]) & (g2148) & (g3515) & (!g924)) + ((!sk[94]) & (g2148) & (g3515) & (g924)) + ((sk[94]) & (!g2148) & (!g3515) & (g924)) + ((sk[94]) & (!g2148) & (g3515) & (g924)) + ((sk[94]) & (g2148) & (g3515) & (!g924)) + ((sk[94]) & (g2148) & (g3515) & (g924)));
	assign g4544 = (((!g2150) & (!g3515) & (!sk[95]) & (g925)) + ((!g2150) & (!g3515) & (sk[95]) & (g925)) + ((!g2150) & (g3515) & (!sk[95]) & (!g925)) + ((!g2150) & (g3515) & (!sk[95]) & (g925)) + ((!g2150) & (g3515) & (sk[95]) & (g925)) + ((g2150) & (!g3515) & (!sk[95]) & (g925)) + ((g2150) & (g3515) & (!sk[95]) & (!g925)) + ((g2150) & (g3515) & (!sk[95]) & (g925)) + ((g2150) & (g3515) & (sk[95]) & (!g925)) + ((g2150) & (g3515) & (sk[95]) & (g925)));
	assign g4545 = (((!sk[96]) & (!g2151) & (!g3515) & (g926)) + ((!sk[96]) & (!g2151) & (g3515) & (!g926)) + ((!sk[96]) & (!g2151) & (g3515) & (g926)) + ((!sk[96]) & (g2151) & (!g3515) & (g926)) + ((!sk[96]) & (g2151) & (g3515) & (!g926)) + ((!sk[96]) & (g2151) & (g3515) & (g926)) + ((sk[96]) & (!g2151) & (!g3515) & (g926)) + ((sk[96]) & (!g2151) & (g3515) & (g926)) + ((sk[96]) & (g2151) & (g3515) & (!g926)) + ((sk[96]) & (g2151) & (g3515) & (g926)));
	assign g927 = (((!g923) & (!g924) & (!g925) & (g926) & (g147) & (g148)) + ((!g923) & (!g924) & (g925) & (!g926) & (!g147) & (g148)) + ((!g923) & (!g924) & (g925) & (g926) & (!g147) & (g148)) + ((!g923) & (!g924) & (g925) & (g926) & (g147) & (g148)) + ((!g923) & (g924) & (!g925) & (!g926) & (g147) & (!g148)) + ((!g923) & (g924) & (!g925) & (g926) & (g147) & (!g148)) + ((!g923) & (g924) & (!g925) & (g926) & (g147) & (g148)) + ((!g923) & (g924) & (g925) & (!g926) & (!g147) & (g148)) + ((!g923) & (g924) & (g925) & (!g926) & (g147) & (!g148)) + ((!g923) & (g924) & (g925) & (g926) & (!g147) & (g148)) + ((!g923) & (g924) & (g925) & (g926) & (g147) & (!g148)) + ((!g923) & (g924) & (g925) & (g926) & (g147) & (g148)) + ((g923) & (!g924) & (!g925) & (!g926) & (!g147) & (!g148)) + ((g923) & (!g924) & (!g925) & (g926) & (!g147) & (!g148)) + ((g923) & (!g924) & (!g925) & (g926) & (g147) & (g148)) + ((g923) & (!g924) & (g925) & (!g926) & (!g147) & (!g148)) + ((g923) & (!g924) & (g925) & (!g926) & (!g147) & (g148)) + ((g923) & (!g924) & (g925) & (g926) & (!g147) & (!g148)) + ((g923) & (!g924) & (g925) & (g926) & (!g147) & (g148)) + ((g923) & (!g924) & (g925) & (g926) & (g147) & (g148)) + ((g923) & (g924) & (!g925) & (!g926) & (!g147) & (!g148)) + ((g923) & (g924) & (!g925) & (!g926) & (g147) & (!g148)) + ((g923) & (g924) & (!g925) & (g926) & (!g147) & (!g148)) + ((g923) & (g924) & (!g925) & (g926) & (g147) & (!g148)) + ((g923) & (g924) & (!g925) & (g926) & (g147) & (g148)) + ((g923) & (g924) & (g925) & (!g926) & (!g147) & (!g148)) + ((g923) & (g924) & (g925) & (!g926) & (!g147) & (g148)) + ((g923) & (g924) & (g925) & (!g926) & (g147) & (!g148)) + ((g923) & (g924) & (g925) & (g926) & (!g147) & (!g148)) + ((g923) & (g924) & (g925) & (g926) & (!g147) & (g148)) + ((g923) & (g924) & (g925) & (g926) & (g147) & (!g148)) + ((g923) & (g924) & (g925) & (g926) & (g147) & (g148)));
	assign g4546 = (((!g2152) & (!g3515) & (!sk[98]) & (g928)) + ((!g2152) & (!g3515) & (sk[98]) & (g928)) + ((!g2152) & (g3515) & (!sk[98]) & (!g928)) + ((!g2152) & (g3515) & (!sk[98]) & (g928)) + ((!g2152) & (g3515) & (sk[98]) & (g928)) + ((g2152) & (!g3515) & (!sk[98]) & (g928)) + ((g2152) & (g3515) & (!sk[98]) & (!g928)) + ((g2152) & (g3515) & (!sk[98]) & (g928)) + ((g2152) & (g3515) & (sk[98]) & (!g928)) + ((g2152) & (g3515) & (sk[98]) & (g928)));
	assign g4547 = (((!g2153) & (!sk[99]) & (!g3515) & (g929)) + ((!g2153) & (!sk[99]) & (g3515) & (!g929)) + ((!g2153) & (!sk[99]) & (g3515) & (g929)) + ((!g2153) & (sk[99]) & (!g3515) & (g929)) + ((!g2153) & (sk[99]) & (g3515) & (g929)) + ((g2153) & (!sk[99]) & (!g3515) & (g929)) + ((g2153) & (!sk[99]) & (g3515) & (!g929)) + ((g2153) & (!sk[99]) & (g3515) & (g929)) + ((g2153) & (sk[99]) & (g3515) & (!g929)) + ((g2153) & (sk[99]) & (g3515) & (g929)));
	assign g4548 = (((!g2155) & (!sk[100]) & (!g3515) & (g930)) + ((!g2155) & (!sk[100]) & (g3515) & (!g930)) + ((!g2155) & (!sk[100]) & (g3515) & (g930)) + ((!g2155) & (sk[100]) & (!g3515) & (g930)) + ((!g2155) & (sk[100]) & (g3515) & (g930)) + ((g2155) & (!sk[100]) & (!g3515) & (g930)) + ((g2155) & (!sk[100]) & (g3515) & (!g930)) + ((g2155) & (!sk[100]) & (g3515) & (g930)) + ((g2155) & (sk[100]) & (g3515) & (!g930)) + ((g2155) & (sk[100]) & (g3515) & (g930)));
	assign g4549 = (((!g2157) & (!sk[101]) & (!g3515) & (g931)) + ((!g2157) & (!sk[101]) & (g3515) & (!g931)) + ((!g2157) & (!sk[101]) & (g3515) & (g931)) + ((!g2157) & (sk[101]) & (!g3515) & (g931)) + ((!g2157) & (sk[101]) & (g3515) & (g931)) + ((g2157) & (!sk[101]) & (!g3515) & (g931)) + ((g2157) & (!sk[101]) & (g3515) & (!g931)) + ((g2157) & (!sk[101]) & (g3515) & (g931)) + ((g2157) & (sk[101]) & (g3515) & (!g931)) + ((g2157) & (sk[101]) & (g3515) & (g931)));
	assign g932 = (((!g928) & (!g929) & (!g930) & (g931) & (g147) & (g148)) + ((!g928) & (!g929) & (g930) & (!g931) & (!g147) & (g148)) + ((!g928) & (!g929) & (g930) & (g931) & (!g147) & (g148)) + ((!g928) & (!g929) & (g930) & (g931) & (g147) & (g148)) + ((!g928) & (g929) & (!g930) & (!g931) & (g147) & (!g148)) + ((!g928) & (g929) & (!g930) & (g931) & (g147) & (!g148)) + ((!g928) & (g929) & (!g930) & (g931) & (g147) & (g148)) + ((!g928) & (g929) & (g930) & (!g931) & (!g147) & (g148)) + ((!g928) & (g929) & (g930) & (!g931) & (g147) & (!g148)) + ((!g928) & (g929) & (g930) & (g931) & (!g147) & (g148)) + ((!g928) & (g929) & (g930) & (g931) & (g147) & (!g148)) + ((!g928) & (g929) & (g930) & (g931) & (g147) & (g148)) + ((g928) & (!g929) & (!g930) & (!g931) & (!g147) & (!g148)) + ((g928) & (!g929) & (!g930) & (g931) & (!g147) & (!g148)) + ((g928) & (!g929) & (!g930) & (g931) & (g147) & (g148)) + ((g928) & (!g929) & (g930) & (!g931) & (!g147) & (!g148)) + ((g928) & (!g929) & (g930) & (!g931) & (!g147) & (g148)) + ((g928) & (!g929) & (g930) & (g931) & (!g147) & (!g148)) + ((g928) & (!g929) & (g930) & (g931) & (!g147) & (g148)) + ((g928) & (!g929) & (g930) & (g931) & (g147) & (g148)) + ((g928) & (g929) & (!g930) & (!g931) & (!g147) & (!g148)) + ((g928) & (g929) & (!g930) & (!g931) & (g147) & (!g148)) + ((g928) & (g929) & (!g930) & (g931) & (!g147) & (!g148)) + ((g928) & (g929) & (!g930) & (g931) & (g147) & (!g148)) + ((g928) & (g929) & (!g930) & (g931) & (g147) & (g148)) + ((g928) & (g929) & (g930) & (!g931) & (!g147) & (!g148)) + ((g928) & (g929) & (g930) & (!g931) & (!g147) & (g148)) + ((g928) & (g929) & (g930) & (!g931) & (g147) & (!g148)) + ((g928) & (g929) & (g930) & (g931) & (!g147) & (!g148)) + ((g928) & (g929) & (g930) & (g931) & (!g147) & (g148)) + ((g928) & (g929) & (g930) & (g931) & (g147) & (!g148)) + ((g928) & (g929) & (g930) & (g931) & (g147) & (g148)));
	assign g4550 = (((!g2158) & (!g3515) & (!sk[103]) & (g933)) + ((!g2158) & (!g3515) & (sk[103]) & (g933)) + ((!g2158) & (g3515) & (!sk[103]) & (!g933)) + ((!g2158) & (g3515) & (!sk[103]) & (g933)) + ((!g2158) & (g3515) & (sk[103]) & (g933)) + ((g2158) & (!g3515) & (!sk[103]) & (g933)) + ((g2158) & (g3515) & (!sk[103]) & (!g933)) + ((g2158) & (g3515) & (!sk[103]) & (g933)) + ((g2158) & (g3515) & (sk[103]) & (!g933)) + ((g2158) & (g3515) & (sk[103]) & (g933)));
	assign g4551 = (((!sk[104]) & (!g2159) & (!g3515) & (g934)) + ((!sk[104]) & (!g2159) & (g3515) & (!g934)) + ((!sk[104]) & (!g2159) & (g3515) & (g934)) + ((!sk[104]) & (g2159) & (!g3515) & (g934)) + ((!sk[104]) & (g2159) & (g3515) & (!g934)) + ((!sk[104]) & (g2159) & (g3515) & (g934)) + ((sk[104]) & (!g2159) & (!g3515) & (g934)) + ((sk[104]) & (!g2159) & (g3515) & (g934)) + ((sk[104]) & (g2159) & (g3515) & (!g934)) + ((sk[104]) & (g2159) & (g3515) & (g934)));
	assign g4552 = (((!g2160) & (!g3515) & (!sk[105]) & (g935)) + ((!g2160) & (!g3515) & (sk[105]) & (g935)) + ((!g2160) & (g3515) & (!sk[105]) & (!g935)) + ((!g2160) & (g3515) & (!sk[105]) & (g935)) + ((!g2160) & (g3515) & (sk[105]) & (g935)) + ((g2160) & (!g3515) & (!sk[105]) & (g935)) + ((g2160) & (g3515) & (!sk[105]) & (!g935)) + ((g2160) & (g3515) & (!sk[105]) & (g935)) + ((g2160) & (g3515) & (sk[105]) & (!g935)) + ((g2160) & (g3515) & (sk[105]) & (g935)));
	assign g4553 = (((!g2161) & (!g3515) & (!sk[106]) & (g936)) + ((!g2161) & (!g3515) & (sk[106]) & (g936)) + ((!g2161) & (g3515) & (!sk[106]) & (!g936)) + ((!g2161) & (g3515) & (!sk[106]) & (g936)) + ((!g2161) & (g3515) & (sk[106]) & (g936)) + ((g2161) & (!g3515) & (!sk[106]) & (g936)) + ((g2161) & (g3515) & (!sk[106]) & (!g936)) + ((g2161) & (g3515) & (!sk[106]) & (g936)) + ((g2161) & (g3515) & (sk[106]) & (!g936)) + ((g2161) & (g3515) & (sk[106]) & (g936)));
	assign g937 = (((!g933) & (!g934) & (!g935) & (g936) & (g147) & (g148)) + ((!g933) & (!g934) & (g935) & (!g936) & (!g147) & (g148)) + ((!g933) & (!g934) & (g935) & (g936) & (!g147) & (g148)) + ((!g933) & (!g934) & (g935) & (g936) & (g147) & (g148)) + ((!g933) & (g934) & (!g935) & (!g936) & (g147) & (!g148)) + ((!g933) & (g934) & (!g935) & (g936) & (g147) & (!g148)) + ((!g933) & (g934) & (!g935) & (g936) & (g147) & (g148)) + ((!g933) & (g934) & (g935) & (!g936) & (!g147) & (g148)) + ((!g933) & (g934) & (g935) & (!g936) & (g147) & (!g148)) + ((!g933) & (g934) & (g935) & (g936) & (!g147) & (g148)) + ((!g933) & (g934) & (g935) & (g936) & (g147) & (!g148)) + ((!g933) & (g934) & (g935) & (g936) & (g147) & (g148)) + ((g933) & (!g934) & (!g935) & (!g936) & (!g147) & (!g148)) + ((g933) & (!g934) & (!g935) & (g936) & (!g147) & (!g148)) + ((g933) & (!g934) & (!g935) & (g936) & (g147) & (g148)) + ((g933) & (!g934) & (g935) & (!g936) & (!g147) & (!g148)) + ((g933) & (!g934) & (g935) & (!g936) & (!g147) & (g148)) + ((g933) & (!g934) & (g935) & (g936) & (!g147) & (!g148)) + ((g933) & (!g934) & (g935) & (g936) & (!g147) & (g148)) + ((g933) & (!g934) & (g935) & (g936) & (g147) & (g148)) + ((g933) & (g934) & (!g935) & (!g936) & (!g147) & (!g148)) + ((g933) & (g934) & (!g935) & (!g936) & (g147) & (!g148)) + ((g933) & (g934) & (!g935) & (g936) & (!g147) & (!g148)) + ((g933) & (g934) & (!g935) & (g936) & (g147) & (!g148)) + ((g933) & (g934) & (!g935) & (g936) & (g147) & (g148)) + ((g933) & (g934) & (g935) & (!g936) & (!g147) & (!g148)) + ((g933) & (g934) & (g935) & (!g936) & (!g147) & (g148)) + ((g933) & (g934) & (g935) & (!g936) & (g147) & (!g148)) + ((g933) & (g934) & (g935) & (g936) & (!g147) & (!g148)) + ((g933) & (g934) & (g935) & (g936) & (!g147) & (g148)) + ((g933) & (g934) & (g935) & (g936) & (g147) & (!g148)) + ((g933) & (g934) & (g935) & (g936) & (g147) & (g148)));
	assign g938 = (((!g922) & (!g927) & (!g932) & (g937) & (g165) & (g166)) + ((!g922) & (!g927) & (g932) & (!g937) & (!g165) & (g166)) + ((!g922) & (!g927) & (g932) & (g937) & (!g165) & (g166)) + ((!g922) & (!g927) & (g932) & (g937) & (g165) & (g166)) + ((!g922) & (g927) & (!g932) & (!g937) & (g165) & (!g166)) + ((!g922) & (g927) & (!g932) & (g937) & (g165) & (!g166)) + ((!g922) & (g927) & (!g932) & (g937) & (g165) & (g166)) + ((!g922) & (g927) & (g932) & (!g937) & (!g165) & (g166)) + ((!g922) & (g927) & (g932) & (!g937) & (g165) & (!g166)) + ((!g922) & (g927) & (g932) & (g937) & (!g165) & (g166)) + ((!g922) & (g927) & (g932) & (g937) & (g165) & (!g166)) + ((!g922) & (g927) & (g932) & (g937) & (g165) & (g166)) + ((g922) & (!g927) & (!g932) & (!g937) & (!g165) & (!g166)) + ((g922) & (!g927) & (!g932) & (g937) & (!g165) & (!g166)) + ((g922) & (!g927) & (!g932) & (g937) & (g165) & (g166)) + ((g922) & (!g927) & (g932) & (!g937) & (!g165) & (!g166)) + ((g922) & (!g927) & (g932) & (!g937) & (!g165) & (g166)) + ((g922) & (!g927) & (g932) & (g937) & (!g165) & (!g166)) + ((g922) & (!g927) & (g932) & (g937) & (!g165) & (g166)) + ((g922) & (!g927) & (g932) & (g937) & (g165) & (g166)) + ((g922) & (g927) & (!g932) & (!g937) & (!g165) & (!g166)) + ((g922) & (g927) & (!g932) & (!g937) & (g165) & (!g166)) + ((g922) & (g927) & (!g932) & (g937) & (!g165) & (!g166)) + ((g922) & (g927) & (!g932) & (g937) & (g165) & (!g166)) + ((g922) & (g927) & (!g932) & (g937) & (g165) & (g166)) + ((g922) & (g927) & (g932) & (!g937) & (!g165) & (!g166)) + ((g922) & (g927) & (g932) & (!g937) & (!g165) & (g166)) + ((g922) & (g927) & (g932) & (!g937) & (g165) & (!g166)) + ((g922) & (g927) & (g932) & (g937) & (!g165) & (!g166)) + ((g922) & (g927) & (g932) & (g937) & (!g165) & (g166)) + ((g922) & (g927) & (g932) & (g937) & (g165) & (!g166)) + ((g922) & (g927) & (g932) & (g937) & (g165) & (g166)));
	assign g4554 = (((!g2173) & (!g3515) & (!sk[109]) & (g939)) + ((!g2173) & (!g3515) & (sk[109]) & (g939)) + ((!g2173) & (g3515) & (!sk[109]) & (!g939)) + ((!g2173) & (g3515) & (!sk[109]) & (g939)) + ((!g2173) & (g3515) & (sk[109]) & (g939)) + ((g2173) & (!g3515) & (!sk[109]) & (g939)) + ((g2173) & (g3515) & (!sk[109]) & (!g939)) + ((g2173) & (g3515) & (!sk[109]) & (g939)) + ((g2173) & (g3515) & (sk[109]) & (!g939)) + ((g2173) & (g3515) & (sk[109]) & (g939)));
	assign g4555 = (((!g2174) & (!sk[110]) & (!g3515) & (g940)) + ((!g2174) & (!sk[110]) & (g3515) & (!g940)) + ((!g2174) & (!sk[110]) & (g3515) & (g940)) + ((!g2174) & (sk[110]) & (!g3515) & (g940)) + ((!g2174) & (sk[110]) & (g3515) & (g940)) + ((g2174) & (!sk[110]) & (!g3515) & (g940)) + ((g2174) & (!sk[110]) & (g3515) & (!g940)) + ((g2174) & (!sk[110]) & (g3515) & (g940)) + ((g2174) & (sk[110]) & (g3515) & (!g940)) + ((g2174) & (sk[110]) & (g3515) & (g940)));
	assign g4556 = (((!g2175) & (!g3515) & (!sk[111]) & (g941)) + ((!g2175) & (!g3515) & (sk[111]) & (g941)) + ((!g2175) & (g3515) & (!sk[111]) & (!g941)) + ((!g2175) & (g3515) & (!sk[111]) & (g941)) + ((!g2175) & (g3515) & (sk[111]) & (g941)) + ((g2175) & (!g3515) & (!sk[111]) & (g941)) + ((g2175) & (g3515) & (!sk[111]) & (!g941)) + ((g2175) & (g3515) & (!sk[111]) & (g941)) + ((g2175) & (g3515) & (sk[111]) & (!g941)) + ((g2175) & (g3515) & (sk[111]) & (g941)));
	assign g4557 = (((!g2176) & (!g3515) & (!sk[112]) & (g942)) + ((!g2176) & (!g3515) & (sk[112]) & (g942)) + ((!g2176) & (g3515) & (!sk[112]) & (!g942)) + ((!g2176) & (g3515) & (!sk[112]) & (g942)) + ((!g2176) & (g3515) & (sk[112]) & (g942)) + ((g2176) & (!g3515) & (!sk[112]) & (g942)) + ((g2176) & (g3515) & (!sk[112]) & (!g942)) + ((g2176) & (g3515) & (!sk[112]) & (g942)) + ((g2176) & (g3515) & (sk[112]) & (!g942)) + ((g2176) & (g3515) & (sk[112]) & (g942)));
	assign g943 = (((!g939) & (!g940) & (!g941) & (g942) & (g165) & (g166)) + ((!g939) & (!g940) & (g941) & (!g942) & (!g165) & (g166)) + ((!g939) & (!g940) & (g941) & (g942) & (!g165) & (g166)) + ((!g939) & (!g940) & (g941) & (g942) & (g165) & (g166)) + ((!g939) & (g940) & (!g941) & (!g942) & (g165) & (!g166)) + ((!g939) & (g940) & (!g941) & (g942) & (g165) & (!g166)) + ((!g939) & (g940) & (!g941) & (g942) & (g165) & (g166)) + ((!g939) & (g940) & (g941) & (!g942) & (!g165) & (g166)) + ((!g939) & (g940) & (g941) & (!g942) & (g165) & (!g166)) + ((!g939) & (g940) & (g941) & (g942) & (!g165) & (g166)) + ((!g939) & (g940) & (g941) & (g942) & (g165) & (!g166)) + ((!g939) & (g940) & (g941) & (g942) & (g165) & (g166)) + ((g939) & (!g940) & (!g941) & (!g942) & (!g165) & (!g166)) + ((g939) & (!g940) & (!g941) & (g942) & (!g165) & (!g166)) + ((g939) & (!g940) & (!g941) & (g942) & (g165) & (g166)) + ((g939) & (!g940) & (g941) & (!g942) & (!g165) & (!g166)) + ((g939) & (!g940) & (g941) & (!g942) & (!g165) & (g166)) + ((g939) & (!g940) & (g941) & (g942) & (!g165) & (!g166)) + ((g939) & (!g940) & (g941) & (g942) & (!g165) & (g166)) + ((g939) & (!g940) & (g941) & (g942) & (g165) & (g166)) + ((g939) & (g940) & (!g941) & (!g942) & (!g165) & (!g166)) + ((g939) & (g940) & (!g941) & (!g942) & (g165) & (!g166)) + ((g939) & (g940) & (!g941) & (g942) & (!g165) & (!g166)) + ((g939) & (g940) & (!g941) & (g942) & (g165) & (!g166)) + ((g939) & (g940) & (!g941) & (g942) & (g165) & (g166)) + ((g939) & (g940) & (g941) & (!g942) & (!g165) & (!g166)) + ((g939) & (g940) & (g941) & (!g942) & (!g165) & (g166)) + ((g939) & (g940) & (g941) & (!g942) & (g165) & (!g166)) + ((g939) & (g940) & (g941) & (g942) & (!g165) & (!g166)) + ((g939) & (g940) & (g941) & (g942) & (!g165) & (g166)) + ((g939) & (g940) & (g941) & (g942) & (g165) & (!g166)) + ((g939) & (g940) & (g941) & (g942) & (g165) & (g166)));
	assign g4558 = (((!g2177) & (!sk[114]) & (!g3515) & (g944)) + ((!g2177) & (!sk[114]) & (g3515) & (!g944)) + ((!g2177) & (!sk[114]) & (g3515) & (g944)) + ((!g2177) & (sk[114]) & (!g3515) & (g944)) + ((!g2177) & (sk[114]) & (g3515) & (g944)) + ((g2177) & (!sk[114]) & (!g3515) & (g944)) + ((g2177) & (!sk[114]) & (g3515) & (!g944)) + ((g2177) & (!sk[114]) & (g3515) & (g944)) + ((g2177) & (sk[114]) & (g3515) & (!g944)) + ((g2177) & (sk[114]) & (g3515) & (g944)));
	assign g4559 = (((!g2178) & (!sk[115]) & (!g3515) & (g945)) + ((!g2178) & (!sk[115]) & (g3515) & (!g945)) + ((!g2178) & (!sk[115]) & (g3515) & (g945)) + ((!g2178) & (sk[115]) & (!g3515) & (g945)) + ((!g2178) & (sk[115]) & (g3515) & (g945)) + ((g2178) & (!sk[115]) & (!g3515) & (g945)) + ((g2178) & (!sk[115]) & (g3515) & (!g945)) + ((g2178) & (!sk[115]) & (g3515) & (g945)) + ((g2178) & (sk[115]) & (g3515) & (!g945)) + ((g2178) & (sk[115]) & (g3515) & (g945)));
	assign g4560 = (((!sk[116]) & (!g2179) & (!g3515) & (g946)) + ((!sk[116]) & (!g2179) & (g3515) & (!g946)) + ((!sk[116]) & (!g2179) & (g3515) & (g946)) + ((!sk[116]) & (g2179) & (!g3515) & (g946)) + ((!sk[116]) & (g2179) & (g3515) & (!g946)) + ((!sk[116]) & (g2179) & (g3515) & (g946)) + ((sk[116]) & (!g2179) & (!g3515) & (g946)) + ((sk[116]) & (!g2179) & (g3515) & (g946)) + ((sk[116]) & (g2179) & (g3515) & (!g946)) + ((sk[116]) & (g2179) & (g3515) & (g946)));
	assign g947 = (((!g165) & (!g166) & (!g944) & (g945) & (!sk[117]) & (!g946)) + ((!g165) & (!g166) & (!g944) & (g945) & (!sk[117]) & (g946)) + ((!g165) & (!g166) & (g944) & (!g945) & (!sk[117]) & (!g946)) + ((!g165) & (!g166) & (g944) & (!g945) & (!sk[117]) & (g946)) + ((!g165) & (!g166) & (g944) & (g945) & (!sk[117]) & (!g946)) + ((!g165) & (!g166) & (g944) & (g945) & (!sk[117]) & (g946)) + ((!g165) & (g166) & (!g944) & (!g945) & (!sk[117]) & (!g946)) + ((!g165) & (g166) & (!g944) & (!g945) & (!sk[117]) & (g946)) + ((!g165) & (g166) & (!g944) & (!g945) & (sk[117]) & (g946)) + ((!g165) & (g166) & (!g944) & (g945) & (!sk[117]) & (!g946)) + ((!g165) & (g166) & (!g944) & (g945) & (!sk[117]) & (g946)) + ((!g165) & (g166) & (!g944) & (g945) & (sk[117]) & (g946)) + ((!g165) & (g166) & (g944) & (!g945) & (!sk[117]) & (!g946)) + ((!g165) & (g166) & (g944) & (!g945) & (!sk[117]) & (g946)) + ((!g165) & (g166) & (g944) & (!g945) & (sk[117]) & (g946)) + ((!g165) & (g166) & (g944) & (g945) & (!sk[117]) & (!g946)) + ((!g165) & (g166) & (g944) & (g945) & (!sk[117]) & (g946)) + ((!g165) & (g166) & (g944) & (g945) & (sk[117]) & (g946)) + ((g165) & (!g166) & (!g944) & (g945) & (!sk[117]) & (!g946)) + ((g165) & (!g166) & (!g944) & (g945) & (!sk[117]) & (g946)) + ((g165) & (!g166) & (g944) & (!g945) & (!sk[117]) & (!g946)) + ((g165) & (!g166) & (g944) & (!g945) & (!sk[117]) & (g946)) + ((g165) & (!g166) & (g944) & (!g945) & (sk[117]) & (!g946)) + ((g165) & (!g166) & (g944) & (!g945) & (sk[117]) & (g946)) + ((g165) & (!g166) & (g944) & (g945) & (!sk[117]) & (!g946)) + ((g165) & (!g166) & (g944) & (g945) & (!sk[117]) & (g946)) + ((g165) & (!g166) & (g944) & (g945) & (sk[117]) & (!g946)) + ((g165) & (!g166) & (g944) & (g945) & (sk[117]) & (g946)) + ((g165) & (g166) & (!g944) & (!g945) & (!sk[117]) & (!g946)) + ((g165) & (g166) & (!g944) & (!g945) & (!sk[117]) & (g946)) + ((g165) & (g166) & (!g944) & (g945) & (!sk[117]) & (!g946)) + ((g165) & (g166) & (!g944) & (g945) & (!sk[117]) & (g946)) + ((g165) & (g166) & (!g944) & (g945) & (sk[117]) & (!g946)) + ((g165) & (g166) & (!g944) & (g945) & (sk[117]) & (g946)) + ((g165) & (g166) & (g944) & (!g945) & (!sk[117]) & (!g946)) + ((g165) & (g166) & (g944) & (!g945) & (!sk[117]) & (g946)) + ((g165) & (g166) & (g944) & (g945) & (!sk[117]) & (!g946)) + ((g165) & (g166) & (g944) & (g945) & (!sk[117]) & (g946)) + ((g165) & (g166) & (g944) & (g945) & (sk[117]) & (!g946)) + ((g165) & (g166) & (g944) & (g945) & (sk[117]) & (g946)));
	assign g4561 = (((!g2162) & (!g3515) & (!sk[118]) & (g948)) + ((!g2162) & (!g3515) & (sk[118]) & (g948)) + ((!g2162) & (g3515) & (!sk[118]) & (!g948)) + ((!g2162) & (g3515) & (!sk[118]) & (g948)) + ((!g2162) & (g3515) & (sk[118]) & (g948)) + ((g2162) & (!g3515) & (!sk[118]) & (g948)) + ((g2162) & (g3515) & (!sk[118]) & (!g948)) + ((g2162) & (g3515) & (!sk[118]) & (g948)) + ((g2162) & (g3515) & (sk[118]) & (!g948)) + ((g2162) & (g3515) & (sk[118]) & (g948)));
	assign g4562 = (((!sk[119]) & (!g2164) & (!g3515) & (g949)) + ((!sk[119]) & (!g2164) & (g3515) & (!g949)) + ((!sk[119]) & (!g2164) & (g3515) & (g949)) + ((!sk[119]) & (g2164) & (!g3515) & (g949)) + ((!sk[119]) & (g2164) & (g3515) & (!g949)) + ((!sk[119]) & (g2164) & (g3515) & (g949)) + ((sk[119]) & (!g2164) & (!g3515) & (g949)) + ((sk[119]) & (!g2164) & (g3515) & (g949)) + ((sk[119]) & (g2164) & (g3515) & (!g949)) + ((sk[119]) & (g2164) & (g3515) & (g949)));
	assign g4563 = (((!sk[120]) & (!g2166) & (!g3515) & (g950)) + ((!sk[120]) & (!g2166) & (g3515) & (!g950)) + ((!sk[120]) & (!g2166) & (g3515) & (g950)) + ((!sk[120]) & (g2166) & (!g3515) & (g950)) + ((!sk[120]) & (g2166) & (g3515) & (!g950)) + ((!sk[120]) & (g2166) & (g3515) & (g950)) + ((sk[120]) & (!g2166) & (!g3515) & (g950)) + ((sk[120]) & (!g2166) & (g3515) & (g950)) + ((sk[120]) & (g2166) & (g3515) & (!g950)) + ((sk[120]) & (g2166) & (g3515) & (g950)));
	assign g4564 = (((!sk[121]) & (!g2168) & (!g3515) & (g951)) + ((!sk[121]) & (!g2168) & (g3515) & (!g951)) + ((!sk[121]) & (!g2168) & (g3515) & (g951)) + ((!sk[121]) & (g2168) & (!g3515) & (g951)) + ((!sk[121]) & (g2168) & (g3515) & (!g951)) + ((!sk[121]) & (g2168) & (g3515) & (g951)) + ((sk[121]) & (!g2168) & (!g3515) & (g951)) + ((sk[121]) & (!g2168) & (g3515) & (g951)) + ((sk[121]) & (g2168) & (g3515) & (!g951)) + ((sk[121]) & (g2168) & (g3515) & (g951)));
	assign g952 = (((!g948) & (!g949) & (!g950) & (g951) & (g165) & (g166)) + ((!g948) & (!g949) & (g950) & (!g951) & (!g165) & (g166)) + ((!g948) & (!g949) & (g950) & (g951) & (!g165) & (g166)) + ((!g948) & (!g949) & (g950) & (g951) & (g165) & (g166)) + ((!g948) & (g949) & (!g950) & (!g951) & (g165) & (!g166)) + ((!g948) & (g949) & (!g950) & (g951) & (g165) & (!g166)) + ((!g948) & (g949) & (!g950) & (g951) & (g165) & (g166)) + ((!g948) & (g949) & (g950) & (!g951) & (!g165) & (g166)) + ((!g948) & (g949) & (g950) & (!g951) & (g165) & (!g166)) + ((!g948) & (g949) & (g950) & (g951) & (!g165) & (g166)) + ((!g948) & (g949) & (g950) & (g951) & (g165) & (!g166)) + ((!g948) & (g949) & (g950) & (g951) & (g165) & (g166)) + ((g948) & (!g949) & (!g950) & (!g951) & (!g165) & (!g166)) + ((g948) & (!g949) & (!g950) & (g951) & (!g165) & (!g166)) + ((g948) & (!g949) & (!g950) & (g951) & (g165) & (g166)) + ((g948) & (!g949) & (g950) & (!g951) & (!g165) & (!g166)) + ((g948) & (!g949) & (g950) & (!g951) & (!g165) & (g166)) + ((g948) & (!g949) & (g950) & (g951) & (!g165) & (!g166)) + ((g948) & (!g949) & (g950) & (g951) & (!g165) & (g166)) + ((g948) & (!g949) & (g950) & (g951) & (g165) & (g166)) + ((g948) & (g949) & (!g950) & (!g951) & (!g165) & (!g166)) + ((g948) & (g949) & (!g950) & (!g951) & (g165) & (!g166)) + ((g948) & (g949) & (!g950) & (g951) & (!g165) & (!g166)) + ((g948) & (g949) & (!g950) & (g951) & (g165) & (!g166)) + ((g948) & (g949) & (!g950) & (g951) & (g165) & (g166)) + ((g948) & (g949) & (g950) & (!g951) & (!g165) & (!g166)) + ((g948) & (g949) & (g950) & (!g951) & (!g165) & (g166)) + ((g948) & (g949) & (g950) & (!g951) & (g165) & (!g166)) + ((g948) & (g949) & (g950) & (g951) & (!g165) & (!g166)) + ((g948) & (g949) & (g950) & (g951) & (!g165) & (g166)) + ((g948) & (g949) & (g950) & (g951) & (g165) & (!g166)) + ((g948) & (g949) & (g950) & (g951) & (g165) & (g166)));
	assign g4565 = (((!sk[123]) & (!g2169) & (!g3515) & (g953)) + ((!sk[123]) & (!g2169) & (g3515) & (!g953)) + ((!sk[123]) & (!g2169) & (g3515) & (g953)) + ((!sk[123]) & (g2169) & (!g3515) & (g953)) + ((!sk[123]) & (g2169) & (g3515) & (!g953)) + ((!sk[123]) & (g2169) & (g3515) & (g953)) + ((sk[123]) & (!g2169) & (!g3515) & (g953)) + ((sk[123]) & (!g2169) & (g3515) & (g953)) + ((sk[123]) & (g2169) & (g3515) & (!g953)) + ((sk[123]) & (g2169) & (g3515) & (g953)));
	assign g4566 = (((!g2170) & (!sk[124]) & (!g3515) & (g954)) + ((!g2170) & (!sk[124]) & (g3515) & (!g954)) + ((!g2170) & (!sk[124]) & (g3515) & (g954)) + ((!g2170) & (sk[124]) & (!g3515) & (g954)) + ((!g2170) & (sk[124]) & (g3515) & (g954)) + ((g2170) & (!sk[124]) & (!g3515) & (g954)) + ((g2170) & (!sk[124]) & (g3515) & (!g954)) + ((g2170) & (!sk[124]) & (g3515) & (g954)) + ((g2170) & (sk[124]) & (g3515) & (!g954)) + ((g2170) & (sk[124]) & (g3515) & (g954)));
	assign g4567 = (((!sk[125]) & (!g2171) & (!g3515) & (g955)) + ((!sk[125]) & (!g2171) & (g3515) & (!g955)) + ((!sk[125]) & (!g2171) & (g3515) & (g955)) + ((!sk[125]) & (g2171) & (!g3515) & (g955)) + ((!sk[125]) & (g2171) & (g3515) & (!g955)) + ((!sk[125]) & (g2171) & (g3515) & (g955)) + ((sk[125]) & (!g2171) & (!g3515) & (g955)) + ((sk[125]) & (!g2171) & (g3515) & (g955)) + ((sk[125]) & (g2171) & (g3515) & (!g955)) + ((sk[125]) & (g2171) & (g3515) & (g955)));
	assign g4568 = (((!g2172) & (!sk[126]) & (!g3515) & (g956)) + ((!g2172) & (!sk[126]) & (g3515) & (!g956)) + ((!g2172) & (!sk[126]) & (g3515) & (g956)) + ((!g2172) & (sk[126]) & (!g3515) & (g956)) + ((!g2172) & (sk[126]) & (g3515) & (g956)) + ((g2172) & (!sk[126]) & (!g3515) & (g956)) + ((g2172) & (!sk[126]) & (g3515) & (!g956)) + ((g2172) & (!sk[126]) & (g3515) & (g956)) + ((g2172) & (sk[126]) & (g3515) & (!g956)) + ((g2172) & (sk[126]) & (g3515) & (g956)));
	assign g957 = (((!g953) & (!g954) & (!g955) & (g956) & (g165) & (g166)) + ((!g953) & (!g954) & (g955) & (!g956) & (!g165) & (g166)) + ((!g953) & (!g954) & (g955) & (g956) & (!g165) & (g166)) + ((!g953) & (!g954) & (g955) & (g956) & (g165) & (g166)) + ((!g953) & (g954) & (!g955) & (!g956) & (g165) & (!g166)) + ((!g953) & (g954) & (!g955) & (g956) & (g165) & (!g166)) + ((!g953) & (g954) & (!g955) & (g956) & (g165) & (g166)) + ((!g953) & (g954) & (g955) & (!g956) & (!g165) & (g166)) + ((!g953) & (g954) & (g955) & (!g956) & (g165) & (!g166)) + ((!g953) & (g954) & (g955) & (g956) & (!g165) & (g166)) + ((!g953) & (g954) & (g955) & (g956) & (g165) & (!g166)) + ((!g953) & (g954) & (g955) & (g956) & (g165) & (g166)) + ((g953) & (!g954) & (!g955) & (!g956) & (!g165) & (!g166)) + ((g953) & (!g954) & (!g955) & (g956) & (!g165) & (!g166)) + ((g953) & (!g954) & (!g955) & (g956) & (g165) & (g166)) + ((g953) & (!g954) & (g955) & (!g956) & (!g165) & (!g166)) + ((g953) & (!g954) & (g955) & (!g956) & (!g165) & (g166)) + ((g953) & (!g954) & (g955) & (g956) & (!g165) & (!g166)) + ((g953) & (!g954) & (g955) & (g956) & (!g165) & (g166)) + ((g953) & (!g954) & (g955) & (g956) & (g165) & (g166)) + ((g953) & (g954) & (!g955) & (!g956) & (!g165) & (!g166)) + ((g953) & (g954) & (!g955) & (!g956) & (g165) & (!g166)) + ((g953) & (g954) & (!g955) & (g956) & (!g165) & (!g166)) + ((g953) & (g954) & (!g955) & (g956) & (g165) & (!g166)) + ((g953) & (g954) & (!g955) & (g956) & (g165) & (g166)) + ((g953) & (g954) & (g955) & (!g956) & (!g165) & (!g166)) + ((g953) & (g954) & (g955) & (!g956) & (!g165) & (g166)) + ((g953) & (g954) & (g955) & (!g956) & (g165) & (!g166)) + ((g953) & (g954) & (g955) & (g956) & (!g165) & (!g166)) + ((g953) & (g954) & (g955) & (g956) & (!g165) & (g166)) + ((g953) & (g954) & (g955) & (g956) & (g165) & (!g166)) + ((g953) & (g954) & (g955) & (g956) & (g165) & (g166)));
	assign g958 = (((!g147) & (!g148) & (!g943) & (g947) & (!g952) & (!g957)) + ((!g147) & (!g148) & (!g943) & (g947) & (!g952) & (g957)) + ((!g147) & (!g148) & (!g943) & (g947) & (g952) & (!g957)) + ((!g147) & (!g148) & (!g943) & (g947) & (g952) & (g957)) + ((!g147) & (!g148) & (g943) & (g947) & (!g952) & (!g957)) + ((!g147) & (!g148) & (g943) & (g947) & (!g952) & (g957)) + ((!g147) & (!g148) & (g943) & (g947) & (g952) & (!g957)) + ((!g147) & (!g148) & (g943) & (g947) & (g952) & (g957)) + ((!g147) & (g148) & (!g943) & (!g947) & (!g952) & (g957)) + ((!g147) & (g148) & (!g943) & (!g947) & (g952) & (g957)) + ((!g147) & (g148) & (!g943) & (g947) & (!g952) & (g957)) + ((!g147) & (g148) & (!g943) & (g947) & (g952) & (g957)) + ((!g147) & (g148) & (g943) & (!g947) & (!g952) & (g957)) + ((!g147) & (g148) & (g943) & (!g947) & (g952) & (g957)) + ((!g147) & (g148) & (g943) & (g947) & (!g952) & (g957)) + ((!g147) & (g148) & (g943) & (g947) & (g952) & (g957)) + ((g147) & (!g148) & (g943) & (!g947) & (!g952) & (!g957)) + ((g147) & (!g148) & (g943) & (!g947) & (!g952) & (g957)) + ((g147) & (!g148) & (g943) & (!g947) & (g952) & (!g957)) + ((g147) & (!g148) & (g943) & (!g947) & (g952) & (g957)) + ((g147) & (!g148) & (g943) & (g947) & (!g952) & (!g957)) + ((g147) & (!g148) & (g943) & (g947) & (!g952) & (g957)) + ((g147) & (!g148) & (g943) & (g947) & (g952) & (!g957)) + ((g147) & (!g148) & (g943) & (g947) & (g952) & (g957)) + ((g147) & (g148) & (!g943) & (!g947) & (g952) & (!g957)) + ((g147) & (g148) & (!g943) & (!g947) & (g952) & (g957)) + ((g147) & (g148) & (!g943) & (g947) & (g952) & (!g957)) + ((g147) & (g148) & (!g943) & (g947) & (g952) & (g957)) + ((g147) & (g148) & (g943) & (!g947) & (g952) & (!g957)) + ((g147) & (g148) & (g943) & (!g947) & (g952) & (g957)) + ((g147) & (g148) & (g943) & (g947) & (g952) & (!g957)) + ((g147) & (g148) & (g943) & (g947) & (g952) & (g957)));
	assign g959 = (((!g142) & (!sk[1]) & (!g938) & (g958)) + ((!g142) & (!sk[1]) & (g938) & (!g958)) + ((!g142) & (!sk[1]) & (g938) & (g958)) + ((!g142) & (sk[1]) & (!g938) & (g958)) + ((!g142) & (sk[1]) & (g938) & (g958)) + ((g142) & (!sk[1]) & (!g938) & (g958)) + ((g142) & (!sk[1]) & (g938) & (!g958)) + ((g142) & (!sk[1]) & (g938) & (g958)) + ((g142) & (sk[1]) & (g938) & (!g958)) + ((g142) & (sk[1]) & (g938) & (g958)));
	assign g4569 = (((!sk[2]) & (!g2059) & (!g2589) & (g960)) + ((!sk[2]) & (!g2059) & (g2589) & (!g960)) + ((!sk[2]) & (!g2059) & (g2589) & (g960)) + ((!sk[2]) & (g2059) & (!g2589) & (g960)) + ((!sk[2]) & (g2059) & (g2589) & (!g960)) + ((!sk[2]) & (g2059) & (g2589) & (g960)) + ((sk[2]) & (!g2059) & (!g2589) & (g960)) + ((sk[2]) & (!g2059) & (g2589) & (g960)) + ((sk[2]) & (g2059) & (g2589) & (!g960)) + ((sk[2]) & (g2059) & (g2589) & (g960)));
	assign g961 = (((!sk[3]) & (!g911) & (!g915) & (g916)) + ((!sk[3]) & (!g911) & (g915) & (!g916)) + ((!sk[3]) & (!g911) & (g915) & (g916)) + ((!sk[3]) & (g911) & (!g915) & (g916)) + ((!sk[3]) & (g911) & (g915) & (!g916)) + ((!sk[3]) & (g911) & (g915) & (g916)) + ((sk[3]) & (!g911) & (!g915) & (!g916)) + ((sk[3]) & (g911) & (!g915) & (!g916)) + ((sk[3]) & (g911) & (!g915) & (g916)) + ((sk[3]) & (g911) & (g915) & (!g916)));
	assign g962 = (((!g126) & (!g959) & (!g960) & (g961) & (!sk[4]) & (!g916)) + ((!g126) & (!g959) & (!g960) & (g961) & (!sk[4]) & (g916)) + ((!g126) & (!g959) & (g960) & (!g961) & (!sk[4]) & (!g916)) + ((!g126) & (!g959) & (g960) & (!g961) & (!sk[4]) & (g916)) + ((!g126) & (!g959) & (g960) & (!g961) & (sk[4]) & (!g916)) + ((!g126) & (!g959) & (g960) & (!g961) & (sk[4]) & (g916)) + ((!g126) & (!g959) & (g960) & (g961) & (!sk[4]) & (!g916)) + ((!g126) & (!g959) & (g960) & (g961) & (!sk[4]) & (g916)) + ((!g126) & (!g959) & (g960) & (g961) & (sk[4]) & (!g916)) + ((!g126) & (!g959) & (g960) & (g961) & (sk[4]) & (g916)) + ((!g126) & (g959) & (!g960) & (!g961) & (!sk[4]) & (!g916)) + ((!g126) & (g959) & (!g960) & (!g961) & (!sk[4]) & (g916)) + ((!g126) & (g959) & (!g960) & (g961) & (!sk[4]) & (!g916)) + ((!g126) & (g959) & (!g960) & (g961) & (!sk[4]) & (g916)) + ((!g126) & (g959) & (g960) & (!g961) & (!sk[4]) & (!g916)) + ((!g126) & (g959) & (g960) & (!g961) & (!sk[4]) & (g916)) + ((!g126) & (g959) & (g960) & (!g961) & (sk[4]) & (!g916)) + ((!g126) & (g959) & (g960) & (!g961) & (sk[4]) & (g916)) + ((!g126) & (g959) & (g960) & (g961) & (!sk[4]) & (!g916)) + ((!g126) & (g959) & (g960) & (g961) & (!sk[4]) & (g916)) + ((!g126) & (g959) & (g960) & (g961) & (sk[4]) & (!g916)) + ((!g126) & (g959) & (g960) & (g961) & (sk[4]) & (g916)) + ((g126) & (!g959) & (!g960) & (!g961) & (sk[4]) & (!g916)) + ((g126) & (!g959) & (!g960) & (g961) & (!sk[4]) & (!g916)) + ((g126) & (!g959) & (!g960) & (g961) & (!sk[4]) & (g916)) + ((g126) & (!g959) & (!g960) & (g961) & (sk[4]) & (g916)) + ((g126) & (!g959) & (g960) & (!g961) & (!sk[4]) & (!g916)) + ((g126) & (!g959) & (g960) & (!g961) & (!sk[4]) & (g916)) + ((g126) & (!g959) & (g960) & (!g961) & (sk[4]) & (!g916)) + ((g126) & (!g959) & (g960) & (g961) & (!sk[4]) & (!g916)) + ((g126) & (!g959) & (g960) & (g961) & (!sk[4]) & (g916)) + ((g126) & (!g959) & (g960) & (g961) & (sk[4]) & (g916)) + ((g126) & (g959) & (!g960) & (!g961) & (!sk[4]) & (!g916)) + ((g126) & (g959) & (!g960) & (!g961) & (!sk[4]) & (g916)) + ((g126) & (g959) & (!g960) & (!g961) & (sk[4]) & (g916)) + ((g126) & (g959) & (!g960) & (g961) & (!sk[4]) & (!g916)) + ((g126) & (g959) & (!g960) & (g961) & (!sk[4]) & (g916)) + ((g126) & (g959) & (!g960) & (g961) & (sk[4]) & (!g916)) + ((g126) & (g959) & (g960) & (!g961) & (!sk[4]) & (!g916)) + ((g126) & (g959) & (g960) & (!g961) & (!sk[4]) & (g916)) + ((g126) & (g959) & (g960) & (!g961) & (sk[4]) & (g916)) + ((g126) & (g959) & (g960) & (g961) & (!sk[4]) & (!g916)) + ((g126) & (g959) & (g960) & (g961) & (!sk[4]) & (g916)) + ((g126) & (g959) & (g960) & (g961) & (sk[4]) & (!g916)));
	assign g4570 = (((!g2140) & (!sk[5]) & (!g3491) & (g963)) + ((!g2140) & (!sk[5]) & (g3491) & (!g963)) + ((!g2140) & (!sk[5]) & (g3491) & (g963)) + ((!g2140) & (sk[5]) & (!g3491) & (g963)) + ((!g2140) & (sk[5]) & (g3491) & (g963)) + ((g2140) & (!sk[5]) & (!g3491) & (g963)) + ((g2140) & (!sk[5]) & (g3491) & (!g963)) + ((g2140) & (!sk[5]) & (g3491) & (g963)) + ((g2140) & (sk[5]) & (g3491) & (!g963)) + ((g2140) & (sk[5]) & (g3491) & (g963)));
	assign g4571 = (((!g2142) & (!sk[6]) & (!g3491) & (g964)) + ((!g2142) & (!sk[6]) & (g3491) & (!g964)) + ((!g2142) & (!sk[6]) & (g3491) & (g964)) + ((!g2142) & (sk[6]) & (!g3491) & (g964)) + ((!g2142) & (sk[6]) & (g3491) & (g964)) + ((g2142) & (!sk[6]) & (!g3491) & (g964)) + ((g2142) & (!sk[6]) & (g3491) & (!g964)) + ((g2142) & (!sk[6]) & (g3491) & (g964)) + ((g2142) & (sk[6]) & (g3491) & (!g964)) + ((g2142) & (sk[6]) & (g3491) & (g964)));
	assign g4572 = (((!sk[7]) & (!g2144) & (!g3491) & (g965)) + ((!sk[7]) & (!g2144) & (g3491) & (!g965)) + ((!sk[7]) & (!g2144) & (g3491) & (g965)) + ((!sk[7]) & (g2144) & (!g3491) & (g965)) + ((!sk[7]) & (g2144) & (g3491) & (!g965)) + ((!sk[7]) & (g2144) & (g3491) & (g965)) + ((sk[7]) & (!g2144) & (!g3491) & (g965)) + ((sk[7]) & (!g2144) & (g3491) & (g965)) + ((sk[7]) & (g2144) & (g3491) & (!g965)) + ((sk[7]) & (g2144) & (g3491) & (g965)));
	assign g4573 = (((!sk[8]) & (!g2145) & (!g3491) & (g966)) + ((!sk[8]) & (!g2145) & (g3491) & (!g966)) + ((!sk[8]) & (!g2145) & (g3491) & (g966)) + ((!sk[8]) & (g2145) & (!g3491) & (g966)) + ((!sk[8]) & (g2145) & (g3491) & (!g966)) + ((!sk[8]) & (g2145) & (g3491) & (g966)) + ((sk[8]) & (!g2145) & (!g3491) & (g966)) + ((sk[8]) & (!g2145) & (g3491) & (g966)) + ((sk[8]) & (g2145) & (g3491) & (!g966)) + ((sk[8]) & (g2145) & (g3491) & (g966)));
	assign g967 = (((!g963) & (!g964) & (!g965) & (g966) & (g147) & (g148)) + ((!g963) & (!g964) & (g965) & (!g966) & (!g147) & (g148)) + ((!g963) & (!g964) & (g965) & (g966) & (!g147) & (g148)) + ((!g963) & (!g964) & (g965) & (g966) & (g147) & (g148)) + ((!g963) & (g964) & (!g965) & (!g966) & (g147) & (!g148)) + ((!g963) & (g964) & (!g965) & (g966) & (g147) & (!g148)) + ((!g963) & (g964) & (!g965) & (g966) & (g147) & (g148)) + ((!g963) & (g964) & (g965) & (!g966) & (!g147) & (g148)) + ((!g963) & (g964) & (g965) & (!g966) & (g147) & (!g148)) + ((!g963) & (g964) & (g965) & (g966) & (!g147) & (g148)) + ((!g963) & (g964) & (g965) & (g966) & (g147) & (!g148)) + ((!g963) & (g964) & (g965) & (g966) & (g147) & (g148)) + ((g963) & (!g964) & (!g965) & (!g966) & (!g147) & (!g148)) + ((g963) & (!g964) & (!g965) & (g966) & (!g147) & (!g148)) + ((g963) & (!g964) & (!g965) & (g966) & (g147) & (g148)) + ((g963) & (!g964) & (g965) & (!g966) & (!g147) & (!g148)) + ((g963) & (!g964) & (g965) & (!g966) & (!g147) & (g148)) + ((g963) & (!g964) & (g965) & (g966) & (!g147) & (!g148)) + ((g963) & (!g964) & (g965) & (g966) & (!g147) & (g148)) + ((g963) & (!g964) & (g965) & (g966) & (g147) & (g148)) + ((g963) & (g964) & (!g965) & (!g966) & (!g147) & (!g148)) + ((g963) & (g964) & (!g965) & (!g966) & (g147) & (!g148)) + ((g963) & (g964) & (!g965) & (g966) & (!g147) & (!g148)) + ((g963) & (g964) & (!g965) & (g966) & (g147) & (!g148)) + ((g963) & (g964) & (!g965) & (g966) & (g147) & (g148)) + ((g963) & (g964) & (g965) & (!g966) & (!g147) & (!g148)) + ((g963) & (g964) & (g965) & (!g966) & (!g147) & (g148)) + ((g963) & (g964) & (g965) & (!g966) & (g147) & (!g148)) + ((g963) & (g964) & (g965) & (g966) & (!g147) & (!g148)) + ((g963) & (g964) & (g965) & (g966) & (!g147) & (g148)) + ((g963) & (g964) & (g965) & (g966) & (g147) & (!g148)) + ((g963) & (g964) & (g965) & (g966) & (g147) & (g148)));
	assign g4574 = (((!sk[10]) & (!g2146) & (!g3491) & (g968)) + ((!sk[10]) & (!g2146) & (g3491) & (!g968)) + ((!sk[10]) & (!g2146) & (g3491) & (g968)) + ((!sk[10]) & (g2146) & (!g3491) & (g968)) + ((!sk[10]) & (g2146) & (g3491) & (!g968)) + ((!sk[10]) & (g2146) & (g3491) & (g968)) + ((sk[10]) & (!g2146) & (!g3491) & (g968)) + ((sk[10]) & (!g2146) & (g3491) & (g968)) + ((sk[10]) & (g2146) & (g3491) & (!g968)) + ((sk[10]) & (g2146) & (g3491) & (g968)));
	assign g4575 = (((!g2148) & (!g3491) & (!sk[11]) & (g969)) + ((!g2148) & (!g3491) & (sk[11]) & (g969)) + ((!g2148) & (g3491) & (!sk[11]) & (!g969)) + ((!g2148) & (g3491) & (!sk[11]) & (g969)) + ((!g2148) & (g3491) & (sk[11]) & (g969)) + ((g2148) & (!g3491) & (!sk[11]) & (g969)) + ((g2148) & (g3491) & (!sk[11]) & (!g969)) + ((g2148) & (g3491) & (!sk[11]) & (g969)) + ((g2148) & (g3491) & (sk[11]) & (!g969)) + ((g2148) & (g3491) & (sk[11]) & (g969)));
	assign g4576 = (((!sk[12]) & (!g2150) & (!g3491) & (g970)) + ((!sk[12]) & (!g2150) & (g3491) & (!g970)) + ((!sk[12]) & (!g2150) & (g3491) & (g970)) + ((!sk[12]) & (g2150) & (!g3491) & (g970)) + ((!sk[12]) & (g2150) & (g3491) & (!g970)) + ((!sk[12]) & (g2150) & (g3491) & (g970)) + ((sk[12]) & (!g2150) & (!g3491) & (g970)) + ((sk[12]) & (!g2150) & (g3491) & (g970)) + ((sk[12]) & (g2150) & (g3491) & (!g970)) + ((sk[12]) & (g2150) & (g3491) & (g970)));
	assign g4577 = (((!sk[13]) & (!g2151) & (!g3491) & (g971)) + ((!sk[13]) & (!g2151) & (g3491) & (!g971)) + ((!sk[13]) & (!g2151) & (g3491) & (g971)) + ((!sk[13]) & (g2151) & (!g3491) & (g971)) + ((!sk[13]) & (g2151) & (g3491) & (!g971)) + ((!sk[13]) & (g2151) & (g3491) & (g971)) + ((sk[13]) & (!g2151) & (!g3491) & (g971)) + ((sk[13]) & (!g2151) & (g3491) & (g971)) + ((sk[13]) & (g2151) & (g3491) & (!g971)) + ((sk[13]) & (g2151) & (g3491) & (g971)));
	assign g972 = (((!g968) & (!g969) & (!g970) & (g971) & (g147) & (g148)) + ((!g968) & (!g969) & (g970) & (!g971) & (!g147) & (g148)) + ((!g968) & (!g969) & (g970) & (g971) & (!g147) & (g148)) + ((!g968) & (!g969) & (g970) & (g971) & (g147) & (g148)) + ((!g968) & (g969) & (!g970) & (!g971) & (g147) & (!g148)) + ((!g968) & (g969) & (!g970) & (g971) & (g147) & (!g148)) + ((!g968) & (g969) & (!g970) & (g971) & (g147) & (g148)) + ((!g968) & (g969) & (g970) & (!g971) & (!g147) & (g148)) + ((!g968) & (g969) & (g970) & (!g971) & (g147) & (!g148)) + ((!g968) & (g969) & (g970) & (g971) & (!g147) & (g148)) + ((!g968) & (g969) & (g970) & (g971) & (g147) & (!g148)) + ((!g968) & (g969) & (g970) & (g971) & (g147) & (g148)) + ((g968) & (!g969) & (!g970) & (!g971) & (!g147) & (!g148)) + ((g968) & (!g969) & (!g970) & (g971) & (!g147) & (!g148)) + ((g968) & (!g969) & (!g970) & (g971) & (g147) & (g148)) + ((g968) & (!g969) & (g970) & (!g971) & (!g147) & (!g148)) + ((g968) & (!g969) & (g970) & (!g971) & (!g147) & (g148)) + ((g968) & (!g969) & (g970) & (g971) & (!g147) & (!g148)) + ((g968) & (!g969) & (g970) & (g971) & (!g147) & (g148)) + ((g968) & (!g969) & (g970) & (g971) & (g147) & (g148)) + ((g968) & (g969) & (!g970) & (!g971) & (!g147) & (!g148)) + ((g968) & (g969) & (!g970) & (!g971) & (g147) & (!g148)) + ((g968) & (g969) & (!g970) & (g971) & (!g147) & (!g148)) + ((g968) & (g969) & (!g970) & (g971) & (g147) & (!g148)) + ((g968) & (g969) & (!g970) & (g971) & (g147) & (g148)) + ((g968) & (g969) & (g970) & (!g971) & (!g147) & (!g148)) + ((g968) & (g969) & (g970) & (!g971) & (!g147) & (g148)) + ((g968) & (g969) & (g970) & (!g971) & (g147) & (!g148)) + ((g968) & (g969) & (g970) & (g971) & (!g147) & (!g148)) + ((g968) & (g969) & (g970) & (g971) & (!g147) & (g148)) + ((g968) & (g969) & (g970) & (g971) & (g147) & (!g148)) + ((g968) & (g969) & (g970) & (g971) & (g147) & (g148)));
	assign g4578 = (((!g2152) & (!sk[15]) & (!g3491) & (g973)) + ((!g2152) & (!sk[15]) & (g3491) & (!g973)) + ((!g2152) & (!sk[15]) & (g3491) & (g973)) + ((!g2152) & (sk[15]) & (!g3491) & (g973)) + ((!g2152) & (sk[15]) & (g3491) & (g973)) + ((g2152) & (!sk[15]) & (!g3491) & (g973)) + ((g2152) & (!sk[15]) & (g3491) & (!g973)) + ((g2152) & (!sk[15]) & (g3491) & (g973)) + ((g2152) & (sk[15]) & (g3491) & (!g973)) + ((g2152) & (sk[15]) & (g3491) & (g973)));
	assign g4579 = (((!g2153) & (!g3491) & (!sk[16]) & (g974)) + ((!g2153) & (!g3491) & (sk[16]) & (g974)) + ((!g2153) & (g3491) & (!sk[16]) & (!g974)) + ((!g2153) & (g3491) & (!sk[16]) & (g974)) + ((!g2153) & (g3491) & (sk[16]) & (g974)) + ((g2153) & (!g3491) & (!sk[16]) & (g974)) + ((g2153) & (g3491) & (!sk[16]) & (!g974)) + ((g2153) & (g3491) & (!sk[16]) & (g974)) + ((g2153) & (g3491) & (sk[16]) & (!g974)) + ((g2153) & (g3491) & (sk[16]) & (g974)));
	assign g4580 = (((!g2155) & (!sk[17]) & (!g3491) & (g975)) + ((!g2155) & (!sk[17]) & (g3491) & (!g975)) + ((!g2155) & (!sk[17]) & (g3491) & (g975)) + ((!g2155) & (sk[17]) & (!g3491) & (g975)) + ((!g2155) & (sk[17]) & (g3491) & (g975)) + ((g2155) & (!sk[17]) & (!g3491) & (g975)) + ((g2155) & (!sk[17]) & (g3491) & (!g975)) + ((g2155) & (!sk[17]) & (g3491) & (g975)) + ((g2155) & (sk[17]) & (g3491) & (!g975)) + ((g2155) & (sk[17]) & (g3491) & (g975)));
	assign g4581 = (((!sk[18]) & (!g2157) & (!g3491) & (g976)) + ((!sk[18]) & (!g2157) & (g3491) & (!g976)) + ((!sk[18]) & (!g2157) & (g3491) & (g976)) + ((!sk[18]) & (g2157) & (!g3491) & (g976)) + ((!sk[18]) & (g2157) & (g3491) & (!g976)) + ((!sk[18]) & (g2157) & (g3491) & (g976)) + ((sk[18]) & (!g2157) & (!g3491) & (g976)) + ((sk[18]) & (!g2157) & (g3491) & (g976)) + ((sk[18]) & (g2157) & (g3491) & (!g976)) + ((sk[18]) & (g2157) & (g3491) & (g976)));
	assign g977 = (((!g973) & (!g974) & (!g975) & (g976) & (g147) & (g148)) + ((!g973) & (!g974) & (g975) & (!g976) & (!g147) & (g148)) + ((!g973) & (!g974) & (g975) & (g976) & (!g147) & (g148)) + ((!g973) & (!g974) & (g975) & (g976) & (g147) & (g148)) + ((!g973) & (g974) & (!g975) & (!g976) & (g147) & (!g148)) + ((!g973) & (g974) & (!g975) & (g976) & (g147) & (!g148)) + ((!g973) & (g974) & (!g975) & (g976) & (g147) & (g148)) + ((!g973) & (g974) & (g975) & (!g976) & (!g147) & (g148)) + ((!g973) & (g974) & (g975) & (!g976) & (g147) & (!g148)) + ((!g973) & (g974) & (g975) & (g976) & (!g147) & (g148)) + ((!g973) & (g974) & (g975) & (g976) & (g147) & (!g148)) + ((!g973) & (g974) & (g975) & (g976) & (g147) & (g148)) + ((g973) & (!g974) & (!g975) & (!g976) & (!g147) & (!g148)) + ((g973) & (!g974) & (!g975) & (g976) & (!g147) & (!g148)) + ((g973) & (!g974) & (!g975) & (g976) & (g147) & (g148)) + ((g973) & (!g974) & (g975) & (!g976) & (!g147) & (!g148)) + ((g973) & (!g974) & (g975) & (!g976) & (!g147) & (g148)) + ((g973) & (!g974) & (g975) & (g976) & (!g147) & (!g148)) + ((g973) & (!g974) & (g975) & (g976) & (!g147) & (g148)) + ((g973) & (!g974) & (g975) & (g976) & (g147) & (g148)) + ((g973) & (g974) & (!g975) & (!g976) & (!g147) & (!g148)) + ((g973) & (g974) & (!g975) & (!g976) & (g147) & (!g148)) + ((g973) & (g974) & (!g975) & (g976) & (!g147) & (!g148)) + ((g973) & (g974) & (!g975) & (g976) & (g147) & (!g148)) + ((g973) & (g974) & (!g975) & (g976) & (g147) & (g148)) + ((g973) & (g974) & (g975) & (!g976) & (!g147) & (!g148)) + ((g973) & (g974) & (g975) & (!g976) & (!g147) & (g148)) + ((g973) & (g974) & (g975) & (!g976) & (g147) & (!g148)) + ((g973) & (g974) & (g975) & (g976) & (!g147) & (!g148)) + ((g973) & (g974) & (g975) & (g976) & (!g147) & (g148)) + ((g973) & (g974) & (g975) & (g976) & (g147) & (!g148)) + ((g973) & (g974) & (g975) & (g976) & (g147) & (g148)));
	assign g4582 = (((!g2158) & (!g3491) & (!sk[20]) & (g978)) + ((!g2158) & (!g3491) & (sk[20]) & (g978)) + ((!g2158) & (g3491) & (!sk[20]) & (!g978)) + ((!g2158) & (g3491) & (!sk[20]) & (g978)) + ((!g2158) & (g3491) & (sk[20]) & (g978)) + ((g2158) & (!g3491) & (!sk[20]) & (g978)) + ((g2158) & (g3491) & (!sk[20]) & (!g978)) + ((g2158) & (g3491) & (!sk[20]) & (g978)) + ((g2158) & (g3491) & (sk[20]) & (!g978)) + ((g2158) & (g3491) & (sk[20]) & (g978)));
	assign g4583 = (((!g2159) & (!g3491) & (!sk[21]) & (g979)) + ((!g2159) & (!g3491) & (sk[21]) & (g979)) + ((!g2159) & (g3491) & (!sk[21]) & (!g979)) + ((!g2159) & (g3491) & (!sk[21]) & (g979)) + ((!g2159) & (g3491) & (sk[21]) & (g979)) + ((g2159) & (!g3491) & (!sk[21]) & (g979)) + ((g2159) & (g3491) & (!sk[21]) & (!g979)) + ((g2159) & (g3491) & (!sk[21]) & (g979)) + ((g2159) & (g3491) & (sk[21]) & (!g979)) + ((g2159) & (g3491) & (sk[21]) & (g979)));
	assign g4584 = (((!sk[22]) & (!g2160) & (!g3491) & (g980)) + ((!sk[22]) & (!g2160) & (g3491) & (!g980)) + ((!sk[22]) & (!g2160) & (g3491) & (g980)) + ((!sk[22]) & (g2160) & (!g3491) & (g980)) + ((!sk[22]) & (g2160) & (g3491) & (!g980)) + ((!sk[22]) & (g2160) & (g3491) & (g980)) + ((sk[22]) & (!g2160) & (!g3491) & (g980)) + ((sk[22]) & (!g2160) & (g3491) & (g980)) + ((sk[22]) & (g2160) & (g3491) & (!g980)) + ((sk[22]) & (g2160) & (g3491) & (g980)));
	assign g4585 = (((!sk[23]) & (!g2161) & (!g3491) & (g981)) + ((!sk[23]) & (!g2161) & (g3491) & (!g981)) + ((!sk[23]) & (!g2161) & (g3491) & (g981)) + ((!sk[23]) & (g2161) & (!g3491) & (g981)) + ((!sk[23]) & (g2161) & (g3491) & (!g981)) + ((!sk[23]) & (g2161) & (g3491) & (g981)) + ((sk[23]) & (!g2161) & (!g3491) & (g981)) + ((sk[23]) & (!g2161) & (g3491) & (g981)) + ((sk[23]) & (g2161) & (g3491) & (!g981)) + ((sk[23]) & (g2161) & (g3491) & (g981)));
	assign g982 = (((!g978) & (!g979) & (!g980) & (g981) & (g147) & (g148)) + ((!g978) & (!g979) & (g980) & (!g981) & (!g147) & (g148)) + ((!g978) & (!g979) & (g980) & (g981) & (!g147) & (g148)) + ((!g978) & (!g979) & (g980) & (g981) & (g147) & (g148)) + ((!g978) & (g979) & (!g980) & (!g981) & (g147) & (!g148)) + ((!g978) & (g979) & (!g980) & (g981) & (g147) & (!g148)) + ((!g978) & (g979) & (!g980) & (g981) & (g147) & (g148)) + ((!g978) & (g979) & (g980) & (!g981) & (!g147) & (g148)) + ((!g978) & (g979) & (g980) & (!g981) & (g147) & (!g148)) + ((!g978) & (g979) & (g980) & (g981) & (!g147) & (g148)) + ((!g978) & (g979) & (g980) & (g981) & (g147) & (!g148)) + ((!g978) & (g979) & (g980) & (g981) & (g147) & (g148)) + ((g978) & (!g979) & (!g980) & (!g981) & (!g147) & (!g148)) + ((g978) & (!g979) & (!g980) & (g981) & (!g147) & (!g148)) + ((g978) & (!g979) & (!g980) & (g981) & (g147) & (g148)) + ((g978) & (!g979) & (g980) & (!g981) & (!g147) & (!g148)) + ((g978) & (!g979) & (g980) & (!g981) & (!g147) & (g148)) + ((g978) & (!g979) & (g980) & (g981) & (!g147) & (!g148)) + ((g978) & (!g979) & (g980) & (g981) & (!g147) & (g148)) + ((g978) & (!g979) & (g980) & (g981) & (g147) & (g148)) + ((g978) & (g979) & (!g980) & (!g981) & (!g147) & (!g148)) + ((g978) & (g979) & (!g980) & (!g981) & (g147) & (!g148)) + ((g978) & (g979) & (!g980) & (g981) & (!g147) & (!g148)) + ((g978) & (g979) & (!g980) & (g981) & (g147) & (!g148)) + ((g978) & (g979) & (!g980) & (g981) & (g147) & (g148)) + ((g978) & (g979) & (g980) & (!g981) & (!g147) & (!g148)) + ((g978) & (g979) & (g980) & (!g981) & (!g147) & (g148)) + ((g978) & (g979) & (g980) & (!g981) & (g147) & (!g148)) + ((g978) & (g979) & (g980) & (g981) & (!g147) & (!g148)) + ((g978) & (g979) & (g980) & (g981) & (!g147) & (g148)) + ((g978) & (g979) & (g980) & (g981) & (g147) & (!g148)) + ((g978) & (g979) & (g980) & (g981) & (g147) & (g148)));
	assign g983 = (((!g967) & (!g972) & (!g977) & (g982) & (g165) & (g166)) + ((!g967) & (!g972) & (g977) & (!g982) & (!g165) & (g166)) + ((!g967) & (!g972) & (g977) & (g982) & (!g165) & (g166)) + ((!g967) & (!g972) & (g977) & (g982) & (g165) & (g166)) + ((!g967) & (g972) & (!g977) & (!g982) & (g165) & (!g166)) + ((!g967) & (g972) & (!g977) & (g982) & (g165) & (!g166)) + ((!g967) & (g972) & (!g977) & (g982) & (g165) & (g166)) + ((!g967) & (g972) & (g977) & (!g982) & (!g165) & (g166)) + ((!g967) & (g972) & (g977) & (!g982) & (g165) & (!g166)) + ((!g967) & (g972) & (g977) & (g982) & (!g165) & (g166)) + ((!g967) & (g972) & (g977) & (g982) & (g165) & (!g166)) + ((!g967) & (g972) & (g977) & (g982) & (g165) & (g166)) + ((g967) & (!g972) & (!g977) & (!g982) & (!g165) & (!g166)) + ((g967) & (!g972) & (!g977) & (g982) & (!g165) & (!g166)) + ((g967) & (!g972) & (!g977) & (g982) & (g165) & (g166)) + ((g967) & (!g972) & (g977) & (!g982) & (!g165) & (!g166)) + ((g967) & (!g972) & (g977) & (!g982) & (!g165) & (g166)) + ((g967) & (!g972) & (g977) & (g982) & (!g165) & (!g166)) + ((g967) & (!g972) & (g977) & (g982) & (!g165) & (g166)) + ((g967) & (!g972) & (g977) & (g982) & (g165) & (g166)) + ((g967) & (g972) & (!g977) & (!g982) & (!g165) & (!g166)) + ((g967) & (g972) & (!g977) & (!g982) & (g165) & (!g166)) + ((g967) & (g972) & (!g977) & (g982) & (!g165) & (!g166)) + ((g967) & (g972) & (!g977) & (g982) & (g165) & (!g166)) + ((g967) & (g972) & (!g977) & (g982) & (g165) & (g166)) + ((g967) & (g972) & (g977) & (!g982) & (!g165) & (!g166)) + ((g967) & (g972) & (g977) & (!g982) & (!g165) & (g166)) + ((g967) & (g972) & (g977) & (!g982) & (g165) & (!g166)) + ((g967) & (g972) & (g977) & (g982) & (!g165) & (!g166)) + ((g967) & (g972) & (g977) & (g982) & (!g165) & (g166)) + ((g967) & (g972) & (g977) & (g982) & (g165) & (!g166)) + ((g967) & (g972) & (g977) & (g982) & (g165) & (g166)));
	assign g4586 = (((!sk[26]) & (!g2173) & (!g3491) & (g984)) + ((!sk[26]) & (!g2173) & (g3491) & (!g984)) + ((!sk[26]) & (!g2173) & (g3491) & (g984)) + ((!sk[26]) & (g2173) & (!g3491) & (g984)) + ((!sk[26]) & (g2173) & (g3491) & (!g984)) + ((!sk[26]) & (g2173) & (g3491) & (g984)) + ((sk[26]) & (!g2173) & (!g3491) & (g984)) + ((sk[26]) & (!g2173) & (g3491) & (g984)) + ((sk[26]) & (g2173) & (g3491) & (!g984)) + ((sk[26]) & (g2173) & (g3491) & (g984)));
	assign g4587 = (((!g2174) & (!g3491) & (!sk[27]) & (g985)) + ((!g2174) & (!g3491) & (sk[27]) & (g985)) + ((!g2174) & (g3491) & (!sk[27]) & (!g985)) + ((!g2174) & (g3491) & (!sk[27]) & (g985)) + ((!g2174) & (g3491) & (sk[27]) & (g985)) + ((g2174) & (!g3491) & (!sk[27]) & (g985)) + ((g2174) & (g3491) & (!sk[27]) & (!g985)) + ((g2174) & (g3491) & (!sk[27]) & (g985)) + ((g2174) & (g3491) & (sk[27]) & (!g985)) + ((g2174) & (g3491) & (sk[27]) & (g985)));
	assign g4588 = (((!g2175) & (!g3491) & (!sk[28]) & (g986)) + ((!g2175) & (!g3491) & (sk[28]) & (g986)) + ((!g2175) & (g3491) & (!sk[28]) & (!g986)) + ((!g2175) & (g3491) & (!sk[28]) & (g986)) + ((!g2175) & (g3491) & (sk[28]) & (g986)) + ((g2175) & (!g3491) & (!sk[28]) & (g986)) + ((g2175) & (g3491) & (!sk[28]) & (!g986)) + ((g2175) & (g3491) & (!sk[28]) & (g986)) + ((g2175) & (g3491) & (sk[28]) & (!g986)) + ((g2175) & (g3491) & (sk[28]) & (g986)));
	assign g4589 = (((!sk[29]) & (!g2176) & (!g3491) & (g987)) + ((!sk[29]) & (!g2176) & (g3491) & (!g987)) + ((!sk[29]) & (!g2176) & (g3491) & (g987)) + ((!sk[29]) & (g2176) & (!g3491) & (g987)) + ((!sk[29]) & (g2176) & (g3491) & (!g987)) + ((!sk[29]) & (g2176) & (g3491) & (g987)) + ((sk[29]) & (!g2176) & (!g3491) & (g987)) + ((sk[29]) & (!g2176) & (g3491) & (g987)) + ((sk[29]) & (g2176) & (g3491) & (!g987)) + ((sk[29]) & (g2176) & (g3491) & (g987)));
	assign g988 = (((!g984) & (!g985) & (!g986) & (g987) & (g165) & (g166)) + ((!g984) & (!g985) & (g986) & (!g987) & (!g165) & (g166)) + ((!g984) & (!g985) & (g986) & (g987) & (!g165) & (g166)) + ((!g984) & (!g985) & (g986) & (g987) & (g165) & (g166)) + ((!g984) & (g985) & (!g986) & (!g987) & (g165) & (!g166)) + ((!g984) & (g985) & (!g986) & (g987) & (g165) & (!g166)) + ((!g984) & (g985) & (!g986) & (g987) & (g165) & (g166)) + ((!g984) & (g985) & (g986) & (!g987) & (!g165) & (g166)) + ((!g984) & (g985) & (g986) & (!g987) & (g165) & (!g166)) + ((!g984) & (g985) & (g986) & (g987) & (!g165) & (g166)) + ((!g984) & (g985) & (g986) & (g987) & (g165) & (!g166)) + ((!g984) & (g985) & (g986) & (g987) & (g165) & (g166)) + ((g984) & (!g985) & (!g986) & (!g987) & (!g165) & (!g166)) + ((g984) & (!g985) & (!g986) & (g987) & (!g165) & (!g166)) + ((g984) & (!g985) & (!g986) & (g987) & (g165) & (g166)) + ((g984) & (!g985) & (g986) & (!g987) & (!g165) & (!g166)) + ((g984) & (!g985) & (g986) & (!g987) & (!g165) & (g166)) + ((g984) & (!g985) & (g986) & (g987) & (!g165) & (!g166)) + ((g984) & (!g985) & (g986) & (g987) & (!g165) & (g166)) + ((g984) & (!g985) & (g986) & (g987) & (g165) & (g166)) + ((g984) & (g985) & (!g986) & (!g987) & (!g165) & (!g166)) + ((g984) & (g985) & (!g986) & (!g987) & (g165) & (!g166)) + ((g984) & (g985) & (!g986) & (g987) & (!g165) & (!g166)) + ((g984) & (g985) & (!g986) & (g987) & (g165) & (!g166)) + ((g984) & (g985) & (!g986) & (g987) & (g165) & (g166)) + ((g984) & (g985) & (g986) & (!g987) & (!g165) & (!g166)) + ((g984) & (g985) & (g986) & (!g987) & (!g165) & (g166)) + ((g984) & (g985) & (g986) & (!g987) & (g165) & (!g166)) + ((g984) & (g985) & (g986) & (g987) & (!g165) & (!g166)) + ((g984) & (g985) & (g986) & (g987) & (!g165) & (g166)) + ((g984) & (g985) & (g986) & (g987) & (g165) & (!g166)) + ((g984) & (g985) & (g986) & (g987) & (g165) & (g166)));
	assign g4590 = (((!g2177) & (!sk[31]) & (!g3491) & (g989)) + ((!g2177) & (!sk[31]) & (g3491) & (!g989)) + ((!g2177) & (!sk[31]) & (g3491) & (g989)) + ((!g2177) & (sk[31]) & (!g3491) & (g989)) + ((!g2177) & (sk[31]) & (g3491) & (g989)) + ((g2177) & (!sk[31]) & (!g3491) & (g989)) + ((g2177) & (!sk[31]) & (g3491) & (!g989)) + ((g2177) & (!sk[31]) & (g3491) & (g989)) + ((g2177) & (sk[31]) & (g3491) & (!g989)) + ((g2177) & (sk[31]) & (g3491) & (g989)));
	assign g4591 = (((!sk[32]) & (!g2178) & (!g3491) & (g990)) + ((!sk[32]) & (!g2178) & (g3491) & (!g990)) + ((!sk[32]) & (!g2178) & (g3491) & (g990)) + ((!sk[32]) & (g2178) & (!g3491) & (g990)) + ((!sk[32]) & (g2178) & (g3491) & (!g990)) + ((!sk[32]) & (g2178) & (g3491) & (g990)) + ((sk[32]) & (!g2178) & (!g3491) & (g990)) + ((sk[32]) & (!g2178) & (g3491) & (g990)) + ((sk[32]) & (g2178) & (g3491) & (!g990)) + ((sk[32]) & (g2178) & (g3491) & (g990)));
	assign g4592 = (((!g2179) & (!g3491) & (!sk[33]) & (g991)) + ((!g2179) & (!g3491) & (sk[33]) & (g991)) + ((!g2179) & (g3491) & (!sk[33]) & (!g991)) + ((!g2179) & (g3491) & (!sk[33]) & (g991)) + ((!g2179) & (g3491) & (sk[33]) & (g991)) + ((g2179) & (!g3491) & (!sk[33]) & (g991)) + ((g2179) & (g3491) & (!sk[33]) & (!g991)) + ((g2179) & (g3491) & (!sk[33]) & (g991)) + ((g2179) & (g3491) & (sk[33]) & (!g991)) + ((g2179) & (g3491) & (sk[33]) & (g991)));
	assign g992 = (((!g165) & (!g166) & (!g989) & (g990) & (!sk[34]) & (!g991)) + ((!g165) & (!g166) & (!g989) & (g990) & (!sk[34]) & (g991)) + ((!g165) & (!g166) & (g989) & (!g990) & (!sk[34]) & (!g991)) + ((!g165) & (!g166) & (g989) & (!g990) & (!sk[34]) & (g991)) + ((!g165) & (!g166) & (g989) & (g990) & (!sk[34]) & (!g991)) + ((!g165) & (!g166) & (g989) & (g990) & (!sk[34]) & (g991)) + ((!g165) & (g166) & (!g989) & (!g990) & (!sk[34]) & (!g991)) + ((!g165) & (g166) & (!g989) & (!g990) & (!sk[34]) & (g991)) + ((!g165) & (g166) & (!g989) & (!g990) & (sk[34]) & (g991)) + ((!g165) & (g166) & (!g989) & (g990) & (!sk[34]) & (!g991)) + ((!g165) & (g166) & (!g989) & (g990) & (!sk[34]) & (g991)) + ((!g165) & (g166) & (!g989) & (g990) & (sk[34]) & (g991)) + ((!g165) & (g166) & (g989) & (!g990) & (!sk[34]) & (!g991)) + ((!g165) & (g166) & (g989) & (!g990) & (!sk[34]) & (g991)) + ((!g165) & (g166) & (g989) & (!g990) & (sk[34]) & (g991)) + ((!g165) & (g166) & (g989) & (g990) & (!sk[34]) & (!g991)) + ((!g165) & (g166) & (g989) & (g990) & (!sk[34]) & (g991)) + ((!g165) & (g166) & (g989) & (g990) & (sk[34]) & (g991)) + ((g165) & (!g166) & (!g989) & (g990) & (!sk[34]) & (!g991)) + ((g165) & (!g166) & (!g989) & (g990) & (!sk[34]) & (g991)) + ((g165) & (!g166) & (g989) & (!g990) & (!sk[34]) & (!g991)) + ((g165) & (!g166) & (g989) & (!g990) & (!sk[34]) & (g991)) + ((g165) & (!g166) & (g989) & (!g990) & (sk[34]) & (!g991)) + ((g165) & (!g166) & (g989) & (!g990) & (sk[34]) & (g991)) + ((g165) & (!g166) & (g989) & (g990) & (!sk[34]) & (!g991)) + ((g165) & (!g166) & (g989) & (g990) & (!sk[34]) & (g991)) + ((g165) & (!g166) & (g989) & (g990) & (sk[34]) & (!g991)) + ((g165) & (!g166) & (g989) & (g990) & (sk[34]) & (g991)) + ((g165) & (g166) & (!g989) & (!g990) & (!sk[34]) & (!g991)) + ((g165) & (g166) & (!g989) & (!g990) & (!sk[34]) & (g991)) + ((g165) & (g166) & (!g989) & (g990) & (!sk[34]) & (!g991)) + ((g165) & (g166) & (!g989) & (g990) & (!sk[34]) & (g991)) + ((g165) & (g166) & (!g989) & (g990) & (sk[34]) & (!g991)) + ((g165) & (g166) & (!g989) & (g990) & (sk[34]) & (g991)) + ((g165) & (g166) & (g989) & (!g990) & (!sk[34]) & (!g991)) + ((g165) & (g166) & (g989) & (!g990) & (!sk[34]) & (g991)) + ((g165) & (g166) & (g989) & (g990) & (!sk[34]) & (!g991)) + ((g165) & (g166) & (g989) & (g990) & (!sk[34]) & (g991)) + ((g165) & (g166) & (g989) & (g990) & (sk[34]) & (!g991)) + ((g165) & (g166) & (g989) & (g990) & (sk[34]) & (g991)));
	assign g4593 = (((!sk[35]) & (!g2162) & (!g3491) & (g993)) + ((!sk[35]) & (!g2162) & (g3491) & (!g993)) + ((!sk[35]) & (!g2162) & (g3491) & (g993)) + ((!sk[35]) & (g2162) & (!g3491) & (g993)) + ((!sk[35]) & (g2162) & (g3491) & (!g993)) + ((!sk[35]) & (g2162) & (g3491) & (g993)) + ((sk[35]) & (!g2162) & (!g3491) & (g993)) + ((sk[35]) & (!g2162) & (g3491) & (g993)) + ((sk[35]) & (g2162) & (g3491) & (!g993)) + ((sk[35]) & (g2162) & (g3491) & (g993)));
	assign g4594 = (((!g2164) & (!sk[36]) & (!g3491) & (g994)) + ((!g2164) & (!sk[36]) & (g3491) & (!g994)) + ((!g2164) & (!sk[36]) & (g3491) & (g994)) + ((!g2164) & (sk[36]) & (!g3491) & (g994)) + ((!g2164) & (sk[36]) & (g3491) & (g994)) + ((g2164) & (!sk[36]) & (!g3491) & (g994)) + ((g2164) & (!sk[36]) & (g3491) & (!g994)) + ((g2164) & (!sk[36]) & (g3491) & (g994)) + ((g2164) & (sk[36]) & (g3491) & (!g994)) + ((g2164) & (sk[36]) & (g3491) & (g994)));
	assign g4595 = (((!sk[37]) & (!g2166) & (!g3491) & (g995)) + ((!sk[37]) & (!g2166) & (g3491) & (!g995)) + ((!sk[37]) & (!g2166) & (g3491) & (g995)) + ((!sk[37]) & (g2166) & (!g3491) & (g995)) + ((!sk[37]) & (g2166) & (g3491) & (!g995)) + ((!sk[37]) & (g2166) & (g3491) & (g995)) + ((sk[37]) & (!g2166) & (!g3491) & (g995)) + ((sk[37]) & (!g2166) & (g3491) & (g995)) + ((sk[37]) & (g2166) & (g3491) & (!g995)) + ((sk[37]) & (g2166) & (g3491) & (g995)));
	assign g4596 = (((!g2168) & (!sk[38]) & (!g3491) & (g996)) + ((!g2168) & (!sk[38]) & (g3491) & (!g996)) + ((!g2168) & (!sk[38]) & (g3491) & (g996)) + ((!g2168) & (sk[38]) & (!g3491) & (g996)) + ((!g2168) & (sk[38]) & (g3491) & (g996)) + ((g2168) & (!sk[38]) & (!g3491) & (g996)) + ((g2168) & (!sk[38]) & (g3491) & (!g996)) + ((g2168) & (!sk[38]) & (g3491) & (g996)) + ((g2168) & (sk[38]) & (g3491) & (!g996)) + ((g2168) & (sk[38]) & (g3491) & (g996)));
	assign g997 = (((!g993) & (!g994) & (!g995) & (g996) & (g165) & (g166)) + ((!g993) & (!g994) & (g995) & (!g996) & (!g165) & (g166)) + ((!g993) & (!g994) & (g995) & (g996) & (!g165) & (g166)) + ((!g993) & (!g994) & (g995) & (g996) & (g165) & (g166)) + ((!g993) & (g994) & (!g995) & (!g996) & (g165) & (!g166)) + ((!g993) & (g994) & (!g995) & (g996) & (g165) & (!g166)) + ((!g993) & (g994) & (!g995) & (g996) & (g165) & (g166)) + ((!g993) & (g994) & (g995) & (!g996) & (!g165) & (g166)) + ((!g993) & (g994) & (g995) & (!g996) & (g165) & (!g166)) + ((!g993) & (g994) & (g995) & (g996) & (!g165) & (g166)) + ((!g993) & (g994) & (g995) & (g996) & (g165) & (!g166)) + ((!g993) & (g994) & (g995) & (g996) & (g165) & (g166)) + ((g993) & (!g994) & (!g995) & (!g996) & (!g165) & (!g166)) + ((g993) & (!g994) & (!g995) & (g996) & (!g165) & (!g166)) + ((g993) & (!g994) & (!g995) & (g996) & (g165) & (g166)) + ((g993) & (!g994) & (g995) & (!g996) & (!g165) & (!g166)) + ((g993) & (!g994) & (g995) & (!g996) & (!g165) & (g166)) + ((g993) & (!g994) & (g995) & (g996) & (!g165) & (!g166)) + ((g993) & (!g994) & (g995) & (g996) & (!g165) & (g166)) + ((g993) & (!g994) & (g995) & (g996) & (g165) & (g166)) + ((g993) & (g994) & (!g995) & (!g996) & (!g165) & (!g166)) + ((g993) & (g994) & (!g995) & (!g996) & (g165) & (!g166)) + ((g993) & (g994) & (!g995) & (g996) & (!g165) & (!g166)) + ((g993) & (g994) & (!g995) & (g996) & (g165) & (!g166)) + ((g993) & (g994) & (!g995) & (g996) & (g165) & (g166)) + ((g993) & (g994) & (g995) & (!g996) & (!g165) & (!g166)) + ((g993) & (g994) & (g995) & (!g996) & (!g165) & (g166)) + ((g993) & (g994) & (g995) & (!g996) & (g165) & (!g166)) + ((g993) & (g994) & (g995) & (g996) & (!g165) & (!g166)) + ((g993) & (g994) & (g995) & (g996) & (!g165) & (g166)) + ((g993) & (g994) & (g995) & (g996) & (g165) & (!g166)) + ((g993) & (g994) & (g995) & (g996) & (g165) & (g166)));
	assign g4597 = (((!g2169) & (!sk[40]) & (!g3491) & (g998)) + ((!g2169) & (!sk[40]) & (g3491) & (!g998)) + ((!g2169) & (!sk[40]) & (g3491) & (g998)) + ((!g2169) & (sk[40]) & (!g3491) & (g998)) + ((!g2169) & (sk[40]) & (g3491) & (g998)) + ((g2169) & (!sk[40]) & (!g3491) & (g998)) + ((g2169) & (!sk[40]) & (g3491) & (!g998)) + ((g2169) & (!sk[40]) & (g3491) & (g998)) + ((g2169) & (sk[40]) & (g3491) & (!g998)) + ((g2169) & (sk[40]) & (g3491) & (g998)));
	assign g4598 = (((!g2170) & (!g3491) & (!sk[41]) & (g999)) + ((!g2170) & (!g3491) & (sk[41]) & (g999)) + ((!g2170) & (g3491) & (!sk[41]) & (!g999)) + ((!g2170) & (g3491) & (!sk[41]) & (g999)) + ((!g2170) & (g3491) & (sk[41]) & (g999)) + ((g2170) & (!g3491) & (!sk[41]) & (g999)) + ((g2170) & (g3491) & (!sk[41]) & (!g999)) + ((g2170) & (g3491) & (!sk[41]) & (g999)) + ((g2170) & (g3491) & (sk[41]) & (!g999)) + ((g2170) & (g3491) & (sk[41]) & (g999)));
	assign g4599 = (((!sk[42]) & (!g2171) & (!g3491) & (g1000)) + ((!sk[42]) & (!g2171) & (g3491) & (!g1000)) + ((!sk[42]) & (!g2171) & (g3491) & (g1000)) + ((!sk[42]) & (g2171) & (!g3491) & (g1000)) + ((!sk[42]) & (g2171) & (g3491) & (!g1000)) + ((!sk[42]) & (g2171) & (g3491) & (g1000)) + ((sk[42]) & (!g2171) & (!g3491) & (g1000)) + ((sk[42]) & (!g2171) & (g3491) & (g1000)) + ((sk[42]) & (g2171) & (g3491) & (!g1000)) + ((sk[42]) & (g2171) & (g3491) & (g1000)));
	assign g4600 = (((!g2172) & (!g3491) & (!sk[43]) & (g1001)) + ((!g2172) & (!g3491) & (sk[43]) & (g1001)) + ((!g2172) & (g3491) & (!sk[43]) & (!g1001)) + ((!g2172) & (g3491) & (!sk[43]) & (g1001)) + ((!g2172) & (g3491) & (sk[43]) & (g1001)) + ((g2172) & (!g3491) & (!sk[43]) & (g1001)) + ((g2172) & (g3491) & (!sk[43]) & (!g1001)) + ((g2172) & (g3491) & (!sk[43]) & (g1001)) + ((g2172) & (g3491) & (sk[43]) & (!g1001)) + ((g2172) & (g3491) & (sk[43]) & (g1001)));
	assign g1002 = (((!g998) & (!g999) & (!g1000) & (g1001) & (g165) & (g166)) + ((!g998) & (!g999) & (g1000) & (!g1001) & (!g165) & (g166)) + ((!g998) & (!g999) & (g1000) & (g1001) & (!g165) & (g166)) + ((!g998) & (!g999) & (g1000) & (g1001) & (g165) & (g166)) + ((!g998) & (g999) & (!g1000) & (!g1001) & (g165) & (!g166)) + ((!g998) & (g999) & (!g1000) & (g1001) & (g165) & (!g166)) + ((!g998) & (g999) & (!g1000) & (g1001) & (g165) & (g166)) + ((!g998) & (g999) & (g1000) & (!g1001) & (!g165) & (g166)) + ((!g998) & (g999) & (g1000) & (!g1001) & (g165) & (!g166)) + ((!g998) & (g999) & (g1000) & (g1001) & (!g165) & (g166)) + ((!g998) & (g999) & (g1000) & (g1001) & (g165) & (!g166)) + ((!g998) & (g999) & (g1000) & (g1001) & (g165) & (g166)) + ((g998) & (!g999) & (!g1000) & (!g1001) & (!g165) & (!g166)) + ((g998) & (!g999) & (!g1000) & (g1001) & (!g165) & (!g166)) + ((g998) & (!g999) & (!g1000) & (g1001) & (g165) & (g166)) + ((g998) & (!g999) & (g1000) & (!g1001) & (!g165) & (!g166)) + ((g998) & (!g999) & (g1000) & (!g1001) & (!g165) & (g166)) + ((g998) & (!g999) & (g1000) & (g1001) & (!g165) & (!g166)) + ((g998) & (!g999) & (g1000) & (g1001) & (!g165) & (g166)) + ((g998) & (!g999) & (g1000) & (g1001) & (g165) & (g166)) + ((g998) & (g999) & (!g1000) & (!g1001) & (!g165) & (!g166)) + ((g998) & (g999) & (!g1000) & (!g1001) & (g165) & (!g166)) + ((g998) & (g999) & (!g1000) & (g1001) & (!g165) & (!g166)) + ((g998) & (g999) & (!g1000) & (g1001) & (g165) & (!g166)) + ((g998) & (g999) & (!g1000) & (g1001) & (g165) & (g166)) + ((g998) & (g999) & (g1000) & (!g1001) & (!g165) & (!g166)) + ((g998) & (g999) & (g1000) & (!g1001) & (!g165) & (g166)) + ((g998) & (g999) & (g1000) & (!g1001) & (g165) & (!g166)) + ((g998) & (g999) & (g1000) & (g1001) & (!g165) & (!g166)) + ((g998) & (g999) & (g1000) & (g1001) & (!g165) & (g166)) + ((g998) & (g999) & (g1000) & (g1001) & (g165) & (!g166)) + ((g998) & (g999) & (g1000) & (g1001) & (g165) & (g166)));
	assign g1003 = (((!g147) & (!g148) & (!g988) & (g992) & (!g997) & (!g1002)) + ((!g147) & (!g148) & (!g988) & (g992) & (!g997) & (g1002)) + ((!g147) & (!g148) & (!g988) & (g992) & (g997) & (!g1002)) + ((!g147) & (!g148) & (!g988) & (g992) & (g997) & (g1002)) + ((!g147) & (!g148) & (g988) & (g992) & (!g997) & (!g1002)) + ((!g147) & (!g148) & (g988) & (g992) & (!g997) & (g1002)) + ((!g147) & (!g148) & (g988) & (g992) & (g997) & (!g1002)) + ((!g147) & (!g148) & (g988) & (g992) & (g997) & (g1002)) + ((!g147) & (g148) & (!g988) & (!g992) & (!g997) & (g1002)) + ((!g147) & (g148) & (!g988) & (!g992) & (g997) & (g1002)) + ((!g147) & (g148) & (!g988) & (g992) & (!g997) & (g1002)) + ((!g147) & (g148) & (!g988) & (g992) & (g997) & (g1002)) + ((!g147) & (g148) & (g988) & (!g992) & (!g997) & (g1002)) + ((!g147) & (g148) & (g988) & (!g992) & (g997) & (g1002)) + ((!g147) & (g148) & (g988) & (g992) & (!g997) & (g1002)) + ((!g147) & (g148) & (g988) & (g992) & (g997) & (g1002)) + ((g147) & (!g148) & (g988) & (!g992) & (!g997) & (!g1002)) + ((g147) & (!g148) & (g988) & (!g992) & (!g997) & (g1002)) + ((g147) & (!g148) & (g988) & (!g992) & (g997) & (!g1002)) + ((g147) & (!g148) & (g988) & (!g992) & (g997) & (g1002)) + ((g147) & (!g148) & (g988) & (g992) & (!g997) & (!g1002)) + ((g147) & (!g148) & (g988) & (g992) & (!g997) & (g1002)) + ((g147) & (!g148) & (g988) & (g992) & (g997) & (!g1002)) + ((g147) & (!g148) & (g988) & (g992) & (g997) & (g1002)) + ((g147) & (g148) & (!g988) & (!g992) & (g997) & (!g1002)) + ((g147) & (g148) & (!g988) & (!g992) & (g997) & (g1002)) + ((g147) & (g148) & (!g988) & (g992) & (g997) & (!g1002)) + ((g147) & (g148) & (!g988) & (g992) & (g997) & (g1002)) + ((g147) & (g148) & (g988) & (!g992) & (g997) & (!g1002)) + ((g147) & (g148) & (g988) & (!g992) & (g997) & (g1002)) + ((g147) & (g148) & (g988) & (g992) & (g997) & (!g1002)) + ((g147) & (g148) & (g988) & (g992) & (g997) & (g1002)));
	assign g1004 = (((!g142) & (!g983) & (!sk[46]) & (g1003)) + ((!g142) & (!g983) & (sk[46]) & (g1003)) + ((!g142) & (g983) & (!sk[46]) & (!g1003)) + ((!g142) & (g983) & (!sk[46]) & (g1003)) + ((!g142) & (g983) & (sk[46]) & (g1003)) + ((g142) & (!g983) & (!sk[46]) & (g1003)) + ((g142) & (g983) & (!sk[46]) & (!g1003)) + ((g142) & (g983) & (!sk[46]) & (g1003)) + ((g142) & (g983) & (sk[46]) & (!g1003)) + ((g142) & (g983) & (sk[46]) & (g1003)));
	assign g4601 = (((!g2059) & (!g2607) & (!sk[47]) & (g1005)) + ((!g2059) & (!g2607) & (sk[47]) & (g1005)) + ((!g2059) & (g2607) & (!sk[47]) & (!g1005)) + ((!g2059) & (g2607) & (!sk[47]) & (g1005)) + ((!g2059) & (g2607) & (sk[47]) & (g1005)) + ((g2059) & (!g2607) & (!sk[47]) & (g1005)) + ((g2059) & (g2607) & (!sk[47]) & (!g1005)) + ((g2059) & (g2607) & (!sk[47]) & (g1005)) + ((g2059) & (g2607) & (sk[47]) & (!g1005)) + ((g2059) & (g2607) & (sk[47]) & (g1005)));
	assign g1006 = (((!g911) & (!sk[48]) & (!g959) & (!g913) & (g914) & (!g916)) + ((!g911) & (!sk[48]) & (!g959) & (!g913) & (g914) & (g916)) + ((!g911) & (!sk[48]) & (!g959) & (g913) & (!g914) & (!g916)) + ((!g911) & (!sk[48]) & (!g959) & (g913) & (!g914) & (g916)) + ((!g911) & (!sk[48]) & (!g959) & (g913) & (g914) & (!g916)) + ((!g911) & (!sk[48]) & (!g959) & (g913) & (g914) & (g916)) + ((!g911) & (!sk[48]) & (g959) & (!g913) & (!g914) & (!g916)) + ((!g911) & (!sk[48]) & (g959) & (!g913) & (!g914) & (g916)) + ((!g911) & (!sk[48]) & (g959) & (!g913) & (g914) & (!g916)) + ((!g911) & (!sk[48]) & (g959) & (!g913) & (g914) & (g916)) + ((!g911) & (!sk[48]) & (g959) & (g913) & (!g914) & (!g916)) + ((!g911) & (!sk[48]) & (g959) & (g913) & (!g914) & (g916)) + ((!g911) & (!sk[48]) & (g959) & (g913) & (g914) & (!g916)) + ((!g911) & (!sk[48]) & (g959) & (g913) & (g914) & (g916)) + ((!g911) & (sk[48]) & (!g959) & (!g913) & (g914) & (!g916)) + ((!g911) & (sk[48]) & (!g959) & (g913) & (!g914) & (!g916)) + ((!g911) & (sk[48]) & (!g959) & (g913) & (g914) & (!g916)) + ((!g911) & (sk[48]) & (g959) & (!g913) & (!g914) & (!g916)) + ((!g911) & (sk[48]) & (g959) & (!g913) & (g914) & (!g916)) + ((!g911) & (sk[48]) & (g959) & (g913) & (!g914) & (!g916)) + ((!g911) & (sk[48]) & (g959) & (g913) & (g914) & (!g916)) + ((g911) & (!sk[48]) & (!g959) & (!g913) & (g914) & (!g916)) + ((g911) & (!sk[48]) & (!g959) & (!g913) & (g914) & (g916)) + ((g911) & (!sk[48]) & (!g959) & (g913) & (!g914) & (!g916)) + ((g911) & (!sk[48]) & (!g959) & (g913) & (!g914) & (g916)) + ((g911) & (!sk[48]) & (!g959) & (g913) & (g914) & (!g916)) + ((g911) & (!sk[48]) & (!g959) & (g913) & (g914) & (g916)) + ((g911) & (!sk[48]) & (g959) & (!g913) & (!g914) & (!g916)) + ((g911) & (!sk[48]) & (g959) & (!g913) & (!g914) & (g916)) + ((g911) & (!sk[48]) & (g959) & (!g913) & (g914) & (!g916)) + ((g911) & (!sk[48]) & (g959) & (!g913) & (g914) & (g916)) + ((g911) & (!sk[48]) & (g959) & (g913) & (!g914) & (!g916)) + ((g911) & (!sk[48]) & (g959) & (g913) & (!g914) & (g916)) + ((g911) & (!sk[48]) & (g959) & (g913) & (g914) & (!g916)) + ((g911) & (!sk[48]) & (g959) & (g913) & (g914) & (g916)) + ((g911) & (sk[48]) & (!g959) & (!g913) & (!g914) & (!g916)) + ((g911) & (sk[48]) & (!g959) & (!g913) & (g914) & (!g916)) + ((g911) & (sk[48]) & (!g959) & (g913) & (!g914) & (!g916)) + ((g911) & (sk[48]) & (!g959) & (g913) & (g914) & (!g916)) + ((g911) & (sk[48]) & (g959) & (!g913) & (!g914) & (!g916)) + ((g911) & (sk[48]) & (g959) & (!g913) & (g914) & (!g916)) + ((g911) & (sk[48]) & (g959) & (!g913) & (g914) & (g916)) + ((g911) & (sk[48]) & (g959) & (g913) & (!g914) & (!g916)) + ((g911) & (sk[48]) & (g959) & (g913) & (!g914) & (g916)) + ((g911) & (sk[48]) & (g959) & (g913) & (g914) & (!g916)) + ((g911) & (sk[48]) & (g959) & (g913) & (g914) & (g916)));
	assign g1007 = (((!g126) & (!sk[49]) & (!g1004) & (!g1005) & (g1006) & (!g916)) + ((!g126) & (!sk[49]) & (!g1004) & (!g1005) & (g1006) & (g916)) + ((!g126) & (!sk[49]) & (!g1004) & (g1005) & (!g1006) & (!g916)) + ((!g126) & (!sk[49]) & (!g1004) & (g1005) & (!g1006) & (g916)) + ((!g126) & (!sk[49]) & (!g1004) & (g1005) & (g1006) & (!g916)) + ((!g126) & (!sk[49]) & (!g1004) & (g1005) & (g1006) & (g916)) + ((!g126) & (!sk[49]) & (g1004) & (!g1005) & (!g1006) & (!g916)) + ((!g126) & (!sk[49]) & (g1004) & (!g1005) & (!g1006) & (g916)) + ((!g126) & (!sk[49]) & (g1004) & (!g1005) & (g1006) & (!g916)) + ((!g126) & (!sk[49]) & (g1004) & (!g1005) & (g1006) & (g916)) + ((!g126) & (!sk[49]) & (g1004) & (g1005) & (!g1006) & (!g916)) + ((!g126) & (!sk[49]) & (g1004) & (g1005) & (!g1006) & (g916)) + ((!g126) & (!sk[49]) & (g1004) & (g1005) & (g1006) & (!g916)) + ((!g126) & (!sk[49]) & (g1004) & (g1005) & (g1006) & (g916)) + ((!g126) & (sk[49]) & (!g1004) & (g1005) & (!g1006) & (!g916)) + ((!g126) & (sk[49]) & (!g1004) & (g1005) & (!g1006) & (g916)) + ((!g126) & (sk[49]) & (!g1004) & (g1005) & (g1006) & (!g916)) + ((!g126) & (sk[49]) & (!g1004) & (g1005) & (g1006) & (g916)) + ((!g126) & (sk[49]) & (g1004) & (g1005) & (!g1006) & (!g916)) + ((!g126) & (sk[49]) & (g1004) & (g1005) & (!g1006) & (g916)) + ((!g126) & (sk[49]) & (g1004) & (g1005) & (g1006) & (!g916)) + ((!g126) & (sk[49]) & (g1004) & (g1005) & (g1006) & (g916)) + ((g126) & (!sk[49]) & (!g1004) & (!g1005) & (g1006) & (!g916)) + ((g126) & (!sk[49]) & (!g1004) & (!g1005) & (g1006) & (g916)) + ((g126) & (!sk[49]) & (!g1004) & (g1005) & (!g1006) & (!g916)) + ((g126) & (!sk[49]) & (!g1004) & (g1005) & (!g1006) & (g916)) + ((g126) & (!sk[49]) & (!g1004) & (g1005) & (g1006) & (!g916)) + ((g126) & (!sk[49]) & (!g1004) & (g1005) & (g1006) & (g916)) + ((g126) & (!sk[49]) & (g1004) & (!g1005) & (!g1006) & (!g916)) + ((g126) & (!sk[49]) & (g1004) & (!g1005) & (!g1006) & (g916)) + ((g126) & (!sk[49]) & (g1004) & (!g1005) & (g1006) & (!g916)) + ((g126) & (!sk[49]) & (g1004) & (!g1005) & (g1006) & (g916)) + ((g126) & (!sk[49]) & (g1004) & (g1005) & (!g1006) & (!g916)) + ((g126) & (!sk[49]) & (g1004) & (g1005) & (!g1006) & (g916)) + ((g126) & (!sk[49]) & (g1004) & (g1005) & (g1006) & (!g916)) + ((g126) & (!sk[49]) & (g1004) & (g1005) & (g1006) & (g916)) + ((g126) & (sk[49]) & (!g1004) & (!g1005) & (!g1006) & (!g916)) + ((g126) & (sk[49]) & (!g1004) & (!g1005) & (g1006) & (g916)) + ((g126) & (sk[49]) & (!g1004) & (g1005) & (!g1006) & (!g916)) + ((g126) & (sk[49]) & (!g1004) & (g1005) & (g1006) & (g916)) + ((g126) & (sk[49]) & (g1004) & (!g1005) & (!g1006) & (g916)) + ((g126) & (sk[49]) & (g1004) & (!g1005) & (g1006) & (!g916)) + ((g126) & (sk[49]) & (g1004) & (g1005) & (!g1006) & (g916)) + ((g126) & (sk[49]) & (g1004) & (g1005) & (g1006) & (!g916)));
	assign g4602 = (((!g2140) & (!sk[50]) & (!g3468) & (g1008)) + ((!g2140) & (!sk[50]) & (g3468) & (!g1008)) + ((!g2140) & (!sk[50]) & (g3468) & (g1008)) + ((!g2140) & (sk[50]) & (!g3468) & (g1008)) + ((!g2140) & (sk[50]) & (g3468) & (g1008)) + ((g2140) & (!sk[50]) & (!g3468) & (g1008)) + ((g2140) & (!sk[50]) & (g3468) & (!g1008)) + ((g2140) & (!sk[50]) & (g3468) & (g1008)) + ((g2140) & (sk[50]) & (g3468) & (!g1008)) + ((g2140) & (sk[50]) & (g3468) & (g1008)));
	assign g4603 = (((!g2142) & (!sk[51]) & (!g3468) & (g1009)) + ((!g2142) & (!sk[51]) & (g3468) & (!g1009)) + ((!g2142) & (!sk[51]) & (g3468) & (g1009)) + ((!g2142) & (sk[51]) & (!g3468) & (g1009)) + ((!g2142) & (sk[51]) & (g3468) & (g1009)) + ((g2142) & (!sk[51]) & (!g3468) & (g1009)) + ((g2142) & (!sk[51]) & (g3468) & (!g1009)) + ((g2142) & (!sk[51]) & (g3468) & (g1009)) + ((g2142) & (sk[51]) & (g3468) & (!g1009)) + ((g2142) & (sk[51]) & (g3468) & (g1009)));
	assign g4604 = (((!g2144) & (!g3468) & (!sk[52]) & (g1010)) + ((!g2144) & (!g3468) & (sk[52]) & (g1010)) + ((!g2144) & (g3468) & (!sk[52]) & (!g1010)) + ((!g2144) & (g3468) & (!sk[52]) & (g1010)) + ((!g2144) & (g3468) & (sk[52]) & (g1010)) + ((g2144) & (!g3468) & (!sk[52]) & (g1010)) + ((g2144) & (g3468) & (!sk[52]) & (!g1010)) + ((g2144) & (g3468) & (!sk[52]) & (g1010)) + ((g2144) & (g3468) & (sk[52]) & (!g1010)) + ((g2144) & (g3468) & (sk[52]) & (g1010)));
	assign g4605 = (((!g2145) & (!sk[53]) & (!g3468) & (g1011)) + ((!g2145) & (!sk[53]) & (g3468) & (!g1011)) + ((!g2145) & (!sk[53]) & (g3468) & (g1011)) + ((!g2145) & (sk[53]) & (!g3468) & (g1011)) + ((!g2145) & (sk[53]) & (g3468) & (g1011)) + ((g2145) & (!sk[53]) & (!g3468) & (g1011)) + ((g2145) & (!sk[53]) & (g3468) & (!g1011)) + ((g2145) & (!sk[53]) & (g3468) & (g1011)) + ((g2145) & (sk[53]) & (g3468) & (!g1011)) + ((g2145) & (sk[53]) & (g3468) & (g1011)));
	assign g1012 = (((!g1008) & (!g1009) & (!g1010) & (g1011) & (g147) & (g148)) + ((!g1008) & (!g1009) & (g1010) & (!g1011) & (!g147) & (g148)) + ((!g1008) & (!g1009) & (g1010) & (g1011) & (!g147) & (g148)) + ((!g1008) & (!g1009) & (g1010) & (g1011) & (g147) & (g148)) + ((!g1008) & (g1009) & (!g1010) & (!g1011) & (g147) & (!g148)) + ((!g1008) & (g1009) & (!g1010) & (g1011) & (g147) & (!g148)) + ((!g1008) & (g1009) & (!g1010) & (g1011) & (g147) & (g148)) + ((!g1008) & (g1009) & (g1010) & (!g1011) & (!g147) & (g148)) + ((!g1008) & (g1009) & (g1010) & (!g1011) & (g147) & (!g148)) + ((!g1008) & (g1009) & (g1010) & (g1011) & (!g147) & (g148)) + ((!g1008) & (g1009) & (g1010) & (g1011) & (g147) & (!g148)) + ((!g1008) & (g1009) & (g1010) & (g1011) & (g147) & (g148)) + ((g1008) & (!g1009) & (!g1010) & (!g1011) & (!g147) & (!g148)) + ((g1008) & (!g1009) & (!g1010) & (g1011) & (!g147) & (!g148)) + ((g1008) & (!g1009) & (!g1010) & (g1011) & (g147) & (g148)) + ((g1008) & (!g1009) & (g1010) & (!g1011) & (!g147) & (!g148)) + ((g1008) & (!g1009) & (g1010) & (!g1011) & (!g147) & (g148)) + ((g1008) & (!g1009) & (g1010) & (g1011) & (!g147) & (!g148)) + ((g1008) & (!g1009) & (g1010) & (g1011) & (!g147) & (g148)) + ((g1008) & (!g1009) & (g1010) & (g1011) & (g147) & (g148)) + ((g1008) & (g1009) & (!g1010) & (!g1011) & (!g147) & (!g148)) + ((g1008) & (g1009) & (!g1010) & (!g1011) & (g147) & (!g148)) + ((g1008) & (g1009) & (!g1010) & (g1011) & (!g147) & (!g148)) + ((g1008) & (g1009) & (!g1010) & (g1011) & (g147) & (!g148)) + ((g1008) & (g1009) & (!g1010) & (g1011) & (g147) & (g148)) + ((g1008) & (g1009) & (g1010) & (!g1011) & (!g147) & (!g148)) + ((g1008) & (g1009) & (g1010) & (!g1011) & (!g147) & (g148)) + ((g1008) & (g1009) & (g1010) & (!g1011) & (g147) & (!g148)) + ((g1008) & (g1009) & (g1010) & (g1011) & (!g147) & (!g148)) + ((g1008) & (g1009) & (g1010) & (g1011) & (!g147) & (g148)) + ((g1008) & (g1009) & (g1010) & (g1011) & (g147) & (!g148)) + ((g1008) & (g1009) & (g1010) & (g1011) & (g147) & (g148)));
	assign g4606 = (((!g2146) & (!sk[55]) & (!g3468) & (g1013)) + ((!g2146) & (!sk[55]) & (g3468) & (!g1013)) + ((!g2146) & (!sk[55]) & (g3468) & (g1013)) + ((!g2146) & (sk[55]) & (!g3468) & (g1013)) + ((!g2146) & (sk[55]) & (g3468) & (g1013)) + ((g2146) & (!sk[55]) & (!g3468) & (g1013)) + ((g2146) & (!sk[55]) & (g3468) & (!g1013)) + ((g2146) & (!sk[55]) & (g3468) & (g1013)) + ((g2146) & (sk[55]) & (g3468) & (!g1013)) + ((g2146) & (sk[55]) & (g3468) & (g1013)));
	assign g4607 = (((!sk[56]) & (!g2148) & (!g3468) & (g1014)) + ((!sk[56]) & (!g2148) & (g3468) & (!g1014)) + ((!sk[56]) & (!g2148) & (g3468) & (g1014)) + ((!sk[56]) & (g2148) & (!g3468) & (g1014)) + ((!sk[56]) & (g2148) & (g3468) & (!g1014)) + ((!sk[56]) & (g2148) & (g3468) & (g1014)) + ((sk[56]) & (!g2148) & (!g3468) & (g1014)) + ((sk[56]) & (!g2148) & (g3468) & (g1014)) + ((sk[56]) & (g2148) & (g3468) & (!g1014)) + ((sk[56]) & (g2148) & (g3468) & (g1014)));
	assign g4608 = (((!sk[57]) & (!g2150) & (!g3468) & (g1015)) + ((!sk[57]) & (!g2150) & (g3468) & (!g1015)) + ((!sk[57]) & (!g2150) & (g3468) & (g1015)) + ((!sk[57]) & (g2150) & (!g3468) & (g1015)) + ((!sk[57]) & (g2150) & (g3468) & (!g1015)) + ((!sk[57]) & (g2150) & (g3468) & (g1015)) + ((sk[57]) & (!g2150) & (!g3468) & (g1015)) + ((sk[57]) & (!g2150) & (g3468) & (g1015)) + ((sk[57]) & (g2150) & (g3468) & (!g1015)) + ((sk[57]) & (g2150) & (g3468) & (g1015)));
	assign g4609 = (((!g2151) & (!g3468) & (!sk[58]) & (g1016)) + ((!g2151) & (!g3468) & (sk[58]) & (g1016)) + ((!g2151) & (g3468) & (!sk[58]) & (!g1016)) + ((!g2151) & (g3468) & (!sk[58]) & (g1016)) + ((!g2151) & (g3468) & (sk[58]) & (g1016)) + ((g2151) & (!g3468) & (!sk[58]) & (g1016)) + ((g2151) & (g3468) & (!sk[58]) & (!g1016)) + ((g2151) & (g3468) & (!sk[58]) & (g1016)) + ((g2151) & (g3468) & (sk[58]) & (!g1016)) + ((g2151) & (g3468) & (sk[58]) & (g1016)));
	assign g1017 = (((!g1013) & (!g1014) & (!g1015) & (g1016) & (g147) & (g148)) + ((!g1013) & (!g1014) & (g1015) & (!g1016) & (!g147) & (g148)) + ((!g1013) & (!g1014) & (g1015) & (g1016) & (!g147) & (g148)) + ((!g1013) & (!g1014) & (g1015) & (g1016) & (g147) & (g148)) + ((!g1013) & (g1014) & (!g1015) & (!g1016) & (g147) & (!g148)) + ((!g1013) & (g1014) & (!g1015) & (g1016) & (g147) & (!g148)) + ((!g1013) & (g1014) & (!g1015) & (g1016) & (g147) & (g148)) + ((!g1013) & (g1014) & (g1015) & (!g1016) & (!g147) & (g148)) + ((!g1013) & (g1014) & (g1015) & (!g1016) & (g147) & (!g148)) + ((!g1013) & (g1014) & (g1015) & (g1016) & (!g147) & (g148)) + ((!g1013) & (g1014) & (g1015) & (g1016) & (g147) & (!g148)) + ((!g1013) & (g1014) & (g1015) & (g1016) & (g147) & (g148)) + ((g1013) & (!g1014) & (!g1015) & (!g1016) & (!g147) & (!g148)) + ((g1013) & (!g1014) & (!g1015) & (g1016) & (!g147) & (!g148)) + ((g1013) & (!g1014) & (!g1015) & (g1016) & (g147) & (g148)) + ((g1013) & (!g1014) & (g1015) & (!g1016) & (!g147) & (!g148)) + ((g1013) & (!g1014) & (g1015) & (!g1016) & (!g147) & (g148)) + ((g1013) & (!g1014) & (g1015) & (g1016) & (!g147) & (!g148)) + ((g1013) & (!g1014) & (g1015) & (g1016) & (!g147) & (g148)) + ((g1013) & (!g1014) & (g1015) & (g1016) & (g147) & (g148)) + ((g1013) & (g1014) & (!g1015) & (!g1016) & (!g147) & (!g148)) + ((g1013) & (g1014) & (!g1015) & (!g1016) & (g147) & (!g148)) + ((g1013) & (g1014) & (!g1015) & (g1016) & (!g147) & (!g148)) + ((g1013) & (g1014) & (!g1015) & (g1016) & (g147) & (!g148)) + ((g1013) & (g1014) & (!g1015) & (g1016) & (g147) & (g148)) + ((g1013) & (g1014) & (g1015) & (!g1016) & (!g147) & (!g148)) + ((g1013) & (g1014) & (g1015) & (!g1016) & (!g147) & (g148)) + ((g1013) & (g1014) & (g1015) & (!g1016) & (g147) & (!g148)) + ((g1013) & (g1014) & (g1015) & (g1016) & (!g147) & (!g148)) + ((g1013) & (g1014) & (g1015) & (g1016) & (!g147) & (g148)) + ((g1013) & (g1014) & (g1015) & (g1016) & (g147) & (!g148)) + ((g1013) & (g1014) & (g1015) & (g1016) & (g147) & (g148)));
	assign g4610 = (((!g2152) & (!sk[60]) & (!g3468) & (g1018)) + ((!g2152) & (!sk[60]) & (g3468) & (!g1018)) + ((!g2152) & (!sk[60]) & (g3468) & (g1018)) + ((!g2152) & (sk[60]) & (!g3468) & (g1018)) + ((!g2152) & (sk[60]) & (g3468) & (g1018)) + ((g2152) & (!sk[60]) & (!g3468) & (g1018)) + ((g2152) & (!sk[60]) & (g3468) & (!g1018)) + ((g2152) & (!sk[60]) & (g3468) & (g1018)) + ((g2152) & (sk[60]) & (g3468) & (!g1018)) + ((g2152) & (sk[60]) & (g3468) & (g1018)));
	assign g4611 = (((!sk[61]) & (!g2153) & (!g3468) & (g1019)) + ((!sk[61]) & (!g2153) & (g3468) & (!g1019)) + ((!sk[61]) & (!g2153) & (g3468) & (g1019)) + ((!sk[61]) & (g2153) & (!g3468) & (g1019)) + ((!sk[61]) & (g2153) & (g3468) & (!g1019)) + ((!sk[61]) & (g2153) & (g3468) & (g1019)) + ((sk[61]) & (!g2153) & (!g3468) & (g1019)) + ((sk[61]) & (!g2153) & (g3468) & (g1019)) + ((sk[61]) & (g2153) & (g3468) & (!g1019)) + ((sk[61]) & (g2153) & (g3468) & (g1019)));
	assign g4612 = (((!g2155) & (!sk[62]) & (!g3468) & (g1020)) + ((!g2155) & (!sk[62]) & (g3468) & (!g1020)) + ((!g2155) & (!sk[62]) & (g3468) & (g1020)) + ((!g2155) & (sk[62]) & (!g3468) & (g1020)) + ((!g2155) & (sk[62]) & (g3468) & (g1020)) + ((g2155) & (!sk[62]) & (!g3468) & (g1020)) + ((g2155) & (!sk[62]) & (g3468) & (!g1020)) + ((g2155) & (!sk[62]) & (g3468) & (g1020)) + ((g2155) & (sk[62]) & (g3468) & (!g1020)) + ((g2155) & (sk[62]) & (g3468) & (g1020)));
	assign g4613 = (((!sk[63]) & (!g2157) & (!g3468) & (g1021)) + ((!sk[63]) & (!g2157) & (g3468) & (!g1021)) + ((!sk[63]) & (!g2157) & (g3468) & (g1021)) + ((!sk[63]) & (g2157) & (!g3468) & (g1021)) + ((!sk[63]) & (g2157) & (g3468) & (!g1021)) + ((!sk[63]) & (g2157) & (g3468) & (g1021)) + ((sk[63]) & (!g2157) & (!g3468) & (g1021)) + ((sk[63]) & (!g2157) & (g3468) & (g1021)) + ((sk[63]) & (g2157) & (g3468) & (!g1021)) + ((sk[63]) & (g2157) & (g3468) & (g1021)));
	assign g1022 = (((!g1018) & (!g1019) & (!g1020) & (g1021) & (g147) & (g148)) + ((!g1018) & (!g1019) & (g1020) & (!g1021) & (!g147) & (g148)) + ((!g1018) & (!g1019) & (g1020) & (g1021) & (!g147) & (g148)) + ((!g1018) & (!g1019) & (g1020) & (g1021) & (g147) & (g148)) + ((!g1018) & (g1019) & (!g1020) & (!g1021) & (g147) & (!g148)) + ((!g1018) & (g1019) & (!g1020) & (g1021) & (g147) & (!g148)) + ((!g1018) & (g1019) & (!g1020) & (g1021) & (g147) & (g148)) + ((!g1018) & (g1019) & (g1020) & (!g1021) & (!g147) & (g148)) + ((!g1018) & (g1019) & (g1020) & (!g1021) & (g147) & (!g148)) + ((!g1018) & (g1019) & (g1020) & (g1021) & (!g147) & (g148)) + ((!g1018) & (g1019) & (g1020) & (g1021) & (g147) & (!g148)) + ((!g1018) & (g1019) & (g1020) & (g1021) & (g147) & (g148)) + ((g1018) & (!g1019) & (!g1020) & (!g1021) & (!g147) & (!g148)) + ((g1018) & (!g1019) & (!g1020) & (g1021) & (!g147) & (!g148)) + ((g1018) & (!g1019) & (!g1020) & (g1021) & (g147) & (g148)) + ((g1018) & (!g1019) & (g1020) & (!g1021) & (!g147) & (!g148)) + ((g1018) & (!g1019) & (g1020) & (!g1021) & (!g147) & (g148)) + ((g1018) & (!g1019) & (g1020) & (g1021) & (!g147) & (!g148)) + ((g1018) & (!g1019) & (g1020) & (g1021) & (!g147) & (g148)) + ((g1018) & (!g1019) & (g1020) & (g1021) & (g147) & (g148)) + ((g1018) & (g1019) & (!g1020) & (!g1021) & (!g147) & (!g148)) + ((g1018) & (g1019) & (!g1020) & (!g1021) & (g147) & (!g148)) + ((g1018) & (g1019) & (!g1020) & (g1021) & (!g147) & (!g148)) + ((g1018) & (g1019) & (!g1020) & (g1021) & (g147) & (!g148)) + ((g1018) & (g1019) & (!g1020) & (g1021) & (g147) & (g148)) + ((g1018) & (g1019) & (g1020) & (!g1021) & (!g147) & (!g148)) + ((g1018) & (g1019) & (g1020) & (!g1021) & (!g147) & (g148)) + ((g1018) & (g1019) & (g1020) & (!g1021) & (g147) & (!g148)) + ((g1018) & (g1019) & (g1020) & (g1021) & (!g147) & (!g148)) + ((g1018) & (g1019) & (g1020) & (g1021) & (!g147) & (g148)) + ((g1018) & (g1019) & (g1020) & (g1021) & (g147) & (!g148)) + ((g1018) & (g1019) & (g1020) & (g1021) & (g147) & (g148)));
	assign g4614 = (((!sk[65]) & (!g2158) & (!g3468) & (g1023)) + ((!sk[65]) & (!g2158) & (g3468) & (!g1023)) + ((!sk[65]) & (!g2158) & (g3468) & (g1023)) + ((!sk[65]) & (g2158) & (!g3468) & (g1023)) + ((!sk[65]) & (g2158) & (g3468) & (!g1023)) + ((!sk[65]) & (g2158) & (g3468) & (g1023)) + ((sk[65]) & (!g2158) & (!g3468) & (g1023)) + ((sk[65]) & (!g2158) & (g3468) & (g1023)) + ((sk[65]) & (g2158) & (g3468) & (!g1023)) + ((sk[65]) & (g2158) & (g3468) & (g1023)));
	assign g4615 = (((!sk[66]) & (!g2159) & (!g3468) & (g1024)) + ((!sk[66]) & (!g2159) & (g3468) & (!g1024)) + ((!sk[66]) & (!g2159) & (g3468) & (g1024)) + ((!sk[66]) & (g2159) & (!g3468) & (g1024)) + ((!sk[66]) & (g2159) & (g3468) & (!g1024)) + ((!sk[66]) & (g2159) & (g3468) & (g1024)) + ((sk[66]) & (!g2159) & (!g3468) & (g1024)) + ((sk[66]) & (!g2159) & (g3468) & (g1024)) + ((sk[66]) & (g2159) & (g3468) & (!g1024)) + ((sk[66]) & (g2159) & (g3468) & (g1024)));
	assign g4616 = (((!sk[67]) & (!g2160) & (!g3468) & (g1025)) + ((!sk[67]) & (!g2160) & (g3468) & (!g1025)) + ((!sk[67]) & (!g2160) & (g3468) & (g1025)) + ((!sk[67]) & (g2160) & (!g3468) & (g1025)) + ((!sk[67]) & (g2160) & (g3468) & (!g1025)) + ((!sk[67]) & (g2160) & (g3468) & (g1025)) + ((sk[67]) & (!g2160) & (!g3468) & (g1025)) + ((sk[67]) & (!g2160) & (g3468) & (g1025)) + ((sk[67]) & (g2160) & (g3468) & (!g1025)) + ((sk[67]) & (g2160) & (g3468) & (g1025)));
	assign g4617 = (((!g2161) & (!g3468) & (!sk[68]) & (g1026)) + ((!g2161) & (!g3468) & (sk[68]) & (g1026)) + ((!g2161) & (g3468) & (!sk[68]) & (!g1026)) + ((!g2161) & (g3468) & (!sk[68]) & (g1026)) + ((!g2161) & (g3468) & (sk[68]) & (g1026)) + ((g2161) & (!g3468) & (!sk[68]) & (g1026)) + ((g2161) & (g3468) & (!sk[68]) & (!g1026)) + ((g2161) & (g3468) & (!sk[68]) & (g1026)) + ((g2161) & (g3468) & (sk[68]) & (!g1026)) + ((g2161) & (g3468) & (sk[68]) & (g1026)));
	assign g1027 = (((!g1023) & (!g1024) & (!g1025) & (g1026) & (g147) & (g148)) + ((!g1023) & (!g1024) & (g1025) & (!g1026) & (!g147) & (g148)) + ((!g1023) & (!g1024) & (g1025) & (g1026) & (!g147) & (g148)) + ((!g1023) & (!g1024) & (g1025) & (g1026) & (g147) & (g148)) + ((!g1023) & (g1024) & (!g1025) & (!g1026) & (g147) & (!g148)) + ((!g1023) & (g1024) & (!g1025) & (g1026) & (g147) & (!g148)) + ((!g1023) & (g1024) & (!g1025) & (g1026) & (g147) & (g148)) + ((!g1023) & (g1024) & (g1025) & (!g1026) & (!g147) & (g148)) + ((!g1023) & (g1024) & (g1025) & (!g1026) & (g147) & (!g148)) + ((!g1023) & (g1024) & (g1025) & (g1026) & (!g147) & (g148)) + ((!g1023) & (g1024) & (g1025) & (g1026) & (g147) & (!g148)) + ((!g1023) & (g1024) & (g1025) & (g1026) & (g147) & (g148)) + ((g1023) & (!g1024) & (!g1025) & (!g1026) & (!g147) & (!g148)) + ((g1023) & (!g1024) & (!g1025) & (g1026) & (!g147) & (!g148)) + ((g1023) & (!g1024) & (!g1025) & (g1026) & (g147) & (g148)) + ((g1023) & (!g1024) & (g1025) & (!g1026) & (!g147) & (!g148)) + ((g1023) & (!g1024) & (g1025) & (!g1026) & (!g147) & (g148)) + ((g1023) & (!g1024) & (g1025) & (g1026) & (!g147) & (!g148)) + ((g1023) & (!g1024) & (g1025) & (g1026) & (!g147) & (g148)) + ((g1023) & (!g1024) & (g1025) & (g1026) & (g147) & (g148)) + ((g1023) & (g1024) & (!g1025) & (!g1026) & (!g147) & (!g148)) + ((g1023) & (g1024) & (!g1025) & (!g1026) & (g147) & (!g148)) + ((g1023) & (g1024) & (!g1025) & (g1026) & (!g147) & (!g148)) + ((g1023) & (g1024) & (!g1025) & (g1026) & (g147) & (!g148)) + ((g1023) & (g1024) & (!g1025) & (g1026) & (g147) & (g148)) + ((g1023) & (g1024) & (g1025) & (!g1026) & (!g147) & (!g148)) + ((g1023) & (g1024) & (g1025) & (!g1026) & (!g147) & (g148)) + ((g1023) & (g1024) & (g1025) & (!g1026) & (g147) & (!g148)) + ((g1023) & (g1024) & (g1025) & (g1026) & (!g147) & (!g148)) + ((g1023) & (g1024) & (g1025) & (g1026) & (!g147) & (g148)) + ((g1023) & (g1024) & (g1025) & (g1026) & (g147) & (!g148)) + ((g1023) & (g1024) & (g1025) & (g1026) & (g147) & (g148)));
	assign g1028 = (((!g1012) & (!g1017) & (!g1022) & (g1027) & (g165) & (g166)) + ((!g1012) & (!g1017) & (g1022) & (!g1027) & (!g165) & (g166)) + ((!g1012) & (!g1017) & (g1022) & (g1027) & (!g165) & (g166)) + ((!g1012) & (!g1017) & (g1022) & (g1027) & (g165) & (g166)) + ((!g1012) & (g1017) & (!g1022) & (!g1027) & (g165) & (!g166)) + ((!g1012) & (g1017) & (!g1022) & (g1027) & (g165) & (!g166)) + ((!g1012) & (g1017) & (!g1022) & (g1027) & (g165) & (g166)) + ((!g1012) & (g1017) & (g1022) & (!g1027) & (!g165) & (g166)) + ((!g1012) & (g1017) & (g1022) & (!g1027) & (g165) & (!g166)) + ((!g1012) & (g1017) & (g1022) & (g1027) & (!g165) & (g166)) + ((!g1012) & (g1017) & (g1022) & (g1027) & (g165) & (!g166)) + ((!g1012) & (g1017) & (g1022) & (g1027) & (g165) & (g166)) + ((g1012) & (!g1017) & (!g1022) & (!g1027) & (!g165) & (!g166)) + ((g1012) & (!g1017) & (!g1022) & (g1027) & (!g165) & (!g166)) + ((g1012) & (!g1017) & (!g1022) & (g1027) & (g165) & (g166)) + ((g1012) & (!g1017) & (g1022) & (!g1027) & (!g165) & (!g166)) + ((g1012) & (!g1017) & (g1022) & (!g1027) & (!g165) & (g166)) + ((g1012) & (!g1017) & (g1022) & (g1027) & (!g165) & (!g166)) + ((g1012) & (!g1017) & (g1022) & (g1027) & (!g165) & (g166)) + ((g1012) & (!g1017) & (g1022) & (g1027) & (g165) & (g166)) + ((g1012) & (g1017) & (!g1022) & (!g1027) & (!g165) & (!g166)) + ((g1012) & (g1017) & (!g1022) & (!g1027) & (g165) & (!g166)) + ((g1012) & (g1017) & (!g1022) & (g1027) & (!g165) & (!g166)) + ((g1012) & (g1017) & (!g1022) & (g1027) & (g165) & (!g166)) + ((g1012) & (g1017) & (!g1022) & (g1027) & (g165) & (g166)) + ((g1012) & (g1017) & (g1022) & (!g1027) & (!g165) & (!g166)) + ((g1012) & (g1017) & (g1022) & (!g1027) & (!g165) & (g166)) + ((g1012) & (g1017) & (g1022) & (!g1027) & (g165) & (!g166)) + ((g1012) & (g1017) & (g1022) & (g1027) & (!g165) & (!g166)) + ((g1012) & (g1017) & (g1022) & (g1027) & (!g165) & (g166)) + ((g1012) & (g1017) & (g1022) & (g1027) & (g165) & (!g166)) + ((g1012) & (g1017) & (g1022) & (g1027) & (g165) & (g166)));
	assign g4618 = (((!g2173) & (!sk[71]) & (!g3468) & (g1029)) + ((!g2173) & (!sk[71]) & (g3468) & (!g1029)) + ((!g2173) & (!sk[71]) & (g3468) & (g1029)) + ((!g2173) & (sk[71]) & (!g3468) & (g1029)) + ((!g2173) & (sk[71]) & (g3468) & (g1029)) + ((g2173) & (!sk[71]) & (!g3468) & (g1029)) + ((g2173) & (!sk[71]) & (g3468) & (!g1029)) + ((g2173) & (!sk[71]) & (g3468) & (g1029)) + ((g2173) & (sk[71]) & (g3468) & (!g1029)) + ((g2173) & (sk[71]) & (g3468) & (g1029)));
	assign g4619 = (((!g2174) & (!g3468) & (!sk[72]) & (g1030)) + ((!g2174) & (!g3468) & (sk[72]) & (g1030)) + ((!g2174) & (g3468) & (!sk[72]) & (!g1030)) + ((!g2174) & (g3468) & (!sk[72]) & (g1030)) + ((!g2174) & (g3468) & (sk[72]) & (g1030)) + ((g2174) & (!g3468) & (!sk[72]) & (g1030)) + ((g2174) & (g3468) & (!sk[72]) & (!g1030)) + ((g2174) & (g3468) & (!sk[72]) & (g1030)) + ((g2174) & (g3468) & (sk[72]) & (!g1030)) + ((g2174) & (g3468) & (sk[72]) & (g1030)));
	assign g4620 = (((!g2175) & (!sk[73]) & (!g3468) & (g1031)) + ((!g2175) & (!sk[73]) & (g3468) & (!g1031)) + ((!g2175) & (!sk[73]) & (g3468) & (g1031)) + ((!g2175) & (sk[73]) & (!g3468) & (g1031)) + ((!g2175) & (sk[73]) & (g3468) & (g1031)) + ((g2175) & (!sk[73]) & (!g3468) & (g1031)) + ((g2175) & (!sk[73]) & (g3468) & (!g1031)) + ((g2175) & (!sk[73]) & (g3468) & (g1031)) + ((g2175) & (sk[73]) & (g3468) & (!g1031)) + ((g2175) & (sk[73]) & (g3468) & (g1031)));
	assign g4621 = (((!g2176) & (!sk[74]) & (!g3468) & (g1032)) + ((!g2176) & (!sk[74]) & (g3468) & (!g1032)) + ((!g2176) & (!sk[74]) & (g3468) & (g1032)) + ((!g2176) & (sk[74]) & (!g3468) & (g1032)) + ((!g2176) & (sk[74]) & (g3468) & (g1032)) + ((g2176) & (!sk[74]) & (!g3468) & (g1032)) + ((g2176) & (!sk[74]) & (g3468) & (!g1032)) + ((g2176) & (!sk[74]) & (g3468) & (g1032)) + ((g2176) & (sk[74]) & (g3468) & (!g1032)) + ((g2176) & (sk[74]) & (g3468) & (g1032)));
	assign g1033 = (((!g1029) & (!g1030) & (!g1031) & (g1032) & (g165) & (g166)) + ((!g1029) & (!g1030) & (g1031) & (!g1032) & (!g165) & (g166)) + ((!g1029) & (!g1030) & (g1031) & (g1032) & (!g165) & (g166)) + ((!g1029) & (!g1030) & (g1031) & (g1032) & (g165) & (g166)) + ((!g1029) & (g1030) & (!g1031) & (!g1032) & (g165) & (!g166)) + ((!g1029) & (g1030) & (!g1031) & (g1032) & (g165) & (!g166)) + ((!g1029) & (g1030) & (!g1031) & (g1032) & (g165) & (g166)) + ((!g1029) & (g1030) & (g1031) & (!g1032) & (!g165) & (g166)) + ((!g1029) & (g1030) & (g1031) & (!g1032) & (g165) & (!g166)) + ((!g1029) & (g1030) & (g1031) & (g1032) & (!g165) & (g166)) + ((!g1029) & (g1030) & (g1031) & (g1032) & (g165) & (!g166)) + ((!g1029) & (g1030) & (g1031) & (g1032) & (g165) & (g166)) + ((g1029) & (!g1030) & (!g1031) & (!g1032) & (!g165) & (!g166)) + ((g1029) & (!g1030) & (!g1031) & (g1032) & (!g165) & (!g166)) + ((g1029) & (!g1030) & (!g1031) & (g1032) & (g165) & (g166)) + ((g1029) & (!g1030) & (g1031) & (!g1032) & (!g165) & (!g166)) + ((g1029) & (!g1030) & (g1031) & (!g1032) & (!g165) & (g166)) + ((g1029) & (!g1030) & (g1031) & (g1032) & (!g165) & (!g166)) + ((g1029) & (!g1030) & (g1031) & (g1032) & (!g165) & (g166)) + ((g1029) & (!g1030) & (g1031) & (g1032) & (g165) & (g166)) + ((g1029) & (g1030) & (!g1031) & (!g1032) & (!g165) & (!g166)) + ((g1029) & (g1030) & (!g1031) & (!g1032) & (g165) & (!g166)) + ((g1029) & (g1030) & (!g1031) & (g1032) & (!g165) & (!g166)) + ((g1029) & (g1030) & (!g1031) & (g1032) & (g165) & (!g166)) + ((g1029) & (g1030) & (!g1031) & (g1032) & (g165) & (g166)) + ((g1029) & (g1030) & (g1031) & (!g1032) & (!g165) & (!g166)) + ((g1029) & (g1030) & (g1031) & (!g1032) & (!g165) & (g166)) + ((g1029) & (g1030) & (g1031) & (!g1032) & (g165) & (!g166)) + ((g1029) & (g1030) & (g1031) & (g1032) & (!g165) & (!g166)) + ((g1029) & (g1030) & (g1031) & (g1032) & (!g165) & (g166)) + ((g1029) & (g1030) & (g1031) & (g1032) & (g165) & (!g166)) + ((g1029) & (g1030) & (g1031) & (g1032) & (g165) & (g166)));
	assign g4622 = (((!g2177) & (!g3468) & (!sk[76]) & (g1034)) + ((!g2177) & (!g3468) & (sk[76]) & (g1034)) + ((!g2177) & (g3468) & (!sk[76]) & (!g1034)) + ((!g2177) & (g3468) & (!sk[76]) & (g1034)) + ((!g2177) & (g3468) & (sk[76]) & (g1034)) + ((g2177) & (!g3468) & (!sk[76]) & (g1034)) + ((g2177) & (g3468) & (!sk[76]) & (!g1034)) + ((g2177) & (g3468) & (!sk[76]) & (g1034)) + ((g2177) & (g3468) & (sk[76]) & (!g1034)) + ((g2177) & (g3468) & (sk[76]) & (g1034)));
	assign g4623 = (((!sk[77]) & (!g2178) & (!g3468) & (g1035)) + ((!sk[77]) & (!g2178) & (g3468) & (!g1035)) + ((!sk[77]) & (!g2178) & (g3468) & (g1035)) + ((!sk[77]) & (g2178) & (!g3468) & (g1035)) + ((!sk[77]) & (g2178) & (g3468) & (!g1035)) + ((!sk[77]) & (g2178) & (g3468) & (g1035)) + ((sk[77]) & (!g2178) & (!g3468) & (g1035)) + ((sk[77]) & (!g2178) & (g3468) & (g1035)) + ((sk[77]) & (g2178) & (g3468) & (!g1035)) + ((sk[77]) & (g2178) & (g3468) & (g1035)));
	assign g4624 = (((!sk[78]) & (!g2179) & (!g3468) & (g1036)) + ((!sk[78]) & (!g2179) & (g3468) & (!g1036)) + ((!sk[78]) & (!g2179) & (g3468) & (g1036)) + ((!sk[78]) & (g2179) & (!g3468) & (g1036)) + ((!sk[78]) & (g2179) & (g3468) & (!g1036)) + ((!sk[78]) & (g2179) & (g3468) & (g1036)) + ((sk[78]) & (!g2179) & (!g3468) & (g1036)) + ((sk[78]) & (!g2179) & (g3468) & (g1036)) + ((sk[78]) & (g2179) & (g3468) & (!g1036)) + ((sk[78]) & (g2179) & (g3468) & (g1036)));
	assign g1037 = (((!g165) & (!g166) & (!sk[79]) & (!g1034) & (g1035) & (!g1036)) + ((!g165) & (!g166) & (!sk[79]) & (!g1034) & (g1035) & (g1036)) + ((!g165) & (!g166) & (!sk[79]) & (g1034) & (!g1035) & (!g1036)) + ((!g165) & (!g166) & (!sk[79]) & (g1034) & (!g1035) & (g1036)) + ((!g165) & (!g166) & (!sk[79]) & (g1034) & (g1035) & (!g1036)) + ((!g165) & (!g166) & (!sk[79]) & (g1034) & (g1035) & (g1036)) + ((!g165) & (g166) & (!sk[79]) & (!g1034) & (!g1035) & (!g1036)) + ((!g165) & (g166) & (!sk[79]) & (!g1034) & (!g1035) & (g1036)) + ((!g165) & (g166) & (!sk[79]) & (!g1034) & (g1035) & (!g1036)) + ((!g165) & (g166) & (!sk[79]) & (!g1034) & (g1035) & (g1036)) + ((!g165) & (g166) & (!sk[79]) & (g1034) & (!g1035) & (!g1036)) + ((!g165) & (g166) & (!sk[79]) & (g1034) & (!g1035) & (g1036)) + ((!g165) & (g166) & (!sk[79]) & (g1034) & (g1035) & (!g1036)) + ((!g165) & (g166) & (!sk[79]) & (g1034) & (g1035) & (g1036)) + ((!g165) & (g166) & (sk[79]) & (!g1034) & (!g1035) & (g1036)) + ((!g165) & (g166) & (sk[79]) & (!g1034) & (g1035) & (g1036)) + ((!g165) & (g166) & (sk[79]) & (g1034) & (!g1035) & (g1036)) + ((!g165) & (g166) & (sk[79]) & (g1034) & (g1035) & (g1036)) + ((g165) & (!g166) & (!sk[79]) & (!g1034) & (g1035) & (!g1036)) + ((g165) & (!g166) & (!sk[79]) & (!g1034) & (g1035) & (g1036)) + ((g165) & (!g166) & (!sk[79]) & (g1034) & (!g1035) & (!g1036)) + ((g165) & (!g166) & (!sk[79]) & (g1034) & (!g1035) & (g1036)) + ((g165) & (!g166) & (!sk[79]) & (g1034) & (g1035) & (!g1036)) + ((g165) & (!g166) & (!sk[79]) & (g1034) & (g1035) & (g1036)) + ((g165) & (!g166) & (sk[79]) & (g1034) & (!g1035) & (!g1036)) + ((g165) & (!g166) & (sk[79]) & (g1034) & (!g1035) & (g1036)) + ((g165) & (!g166) & (sk[79]) & (g1034) & (g1035) & (!g1036)) + ((g165) & (!g166) & (sk[79]) & (g1034) & (g1035) & (g1036)) + ((g165) & (g166) & (!sk[79]) & (!g1034) & (!g1035) & (!g1036)) + ((g165) & (g166) & (!sk[79]) & (!g1034) & (!g1035) & (g1036)) + ((g165) & (g166) & (!sk[79]) & (!g1034) & (g1035) & (!g1036)) + ((g165) & (g166) & (!sk[79]) & (!g1034) & (g1035) & (g1036)) + ((g165) & (g166) & (!sk[79]) & (g1034) & (!g1035) & (!g1036)) + ((g165) & (g166) & (!sk[79]) & (g1034) & (!g1035) & (g1036)) + ((g165) & (g166) & (!sk[79]) & (g1034) & (g1035) & (!g1036)) + ((g165) & (g166) & (!sk[79]) & (g1034) & (g1035) & (g1036)) + ((g165) & (g166) & (sk[79]) & (!g1034) & (g1035) & (!g1036)) + ((g165) & (g166) & (sk[79]) & (!g1034) & (g1035) & (g1036)) + ((g165) & (g166) & (sk[79]) & (g1034) & (g1035) & (!g1036)) + ((g165) & (g166) & (sk[79]) & (g1034) & (g1035) & (g1036)));
	assign g4625 = (((!g2162) & (!g3468) & (!sk[80]) & (g1038)) + ((!g2162) & (!g3468) & (sk[80]) & (g1038)) + ((!g2162) & (g3468) & (!sk[80]) & (!g1038)) + ((!g2162) & (g3468) & (!sk[80]) & (g1038)) + ((!g2162) & (g3468) & (sk[80]) & (g1038)) + ((g2162) & (!g3468) & (!sk[80]) & (g1038)) + ((g2162) & (g3468) & (!sk[80]) & (!g1038)) + ((g2162) & (g3468) & (!sk[80]) & (g1038)) + ((g2162) & (g3468) & (sk[80]) & (!g1038)) + ((g2162) & (g3468) & (sk[80]) & (g1038)));
	assign g4626 = (((!g2164) & (!sk[81]) & (!g3468) & (g1039)) + ((!g2164) & (!sk[81]) & (g3468) & (!g1039)) + ((!g2164) & (!sk[81]) & (g3468) & (g1039)) + ((!g2164) & (sk[81]) & (!g3468) & (g1039)) + ((!g2164) & (sk[81]) & (g3468) & (g1039)) + ((g2164) & (!sk[81]) & (!g3468) & (g1039)) + ((g2164) & (!sk[81]) & (g3468) & (!g1039)) + ((g2164) & (!sk[81]) & (g3468) & (g1039)) + ((g2164) & (sk[81]) & (g3468) & (!g1039)) + ((g2164) & (sk[81]) & (g3468) & (g1039)));
	assign g4627 = (((!g2166) & (!g3468) & (!sk[82]) & (g1040)) + ((!g2166) & (!g3468) & (sk[82]) & (g1040)) + ((!g2166) & (g3468) & (!sk[82]) & (!g1040)) + ((!g2166) & (g3468) & (!sk[82]) & (g1040)) + ((!g2166) & (g3468) & (sk[82]) & (g1040)) + ((g2166) & (!g3468) & (!sk[82]) & (g1040)) + ((g2166) & (g3468) & (!sk[82]) & (!g1040)) + ((g2166) & (g3468) & (!sk[82]) & (g1040)) + ((g2166) & (g3468) & (sk[82]) & (!g1040)) + ((g2166) & (g3468) & (sk[82]) & (g1040)));
	assign g4628 = (((!g2168) & (!g3468) & (!sk[83]) & (g1041)) + ((!g2168) & (!g3468) & (sk[83]) & (g1041)) + ((!g2168) & (g3468) & (!sk[83]) & (!g1041)) + ((!g2168) & (g3468) & (!sk[83]) & (g1041)) + ((!g2168) & (g3468) & (sk[83]) & (g1041)) + ((g2168) & (!g3468) & (!sk[83]) & (g1041)) + ((g2168) & (g3468) & (!sk[83]) & (!g1041)) + ((g2168) & (g3468) & (!sk[83]) & (g1041)) + ((g2168) & (g3468) & (sk[83]) & (!g1041)) + ((g2168) & (g3468) & (sk[83]) & (g1041)));
	assign g1042 = (((!g1038) & (!g1039) & (!g1040) & (g1041) & (g165) & (g166)) + ((!g1038) & (!g1039) & (g1040) & (!g1041) & (!g165) & (g166)) + ((!g1038) & (!g1039) & (g1040) & (g1041) & (!g165) & (g166)) + ((!g1038) & (!g1039) & (g1040) & (g1041) & (g165) & (g166)) + ((!g1038) & (g1039) & (!g1040) & (!g1041) & (g165) & (!g166)) + ((!g1038) & (g1039) & (!g1040) & (g1041) & (g165) & (!g166)) + ((!g1038) & (g1039) & (!g1040) & (g1041) & (g165) & (g166)) + ((!g1038) & (g1039) & (g1040) & (!g1041) & (!g165) & (g166)) + ((!g1038) & (g1039) & (g1040) & (!g1041) & (g165) & (!g166)) + ((!g1038) & (g1039) & (g1040) & (g1041) & (!g165) & (g166)) + ((!g1038) & (g1039) & (g1040) & (g1041) & (g165) & (!g166)) + ((!g1038) & (g1039) & (g1040) & (g1041) & (g165) & (g166)) + ((g1038) & (!g1039) & (!g1040) & (!g1041) & (!g165) & (!g166)) + ((g1038) & (!g1039) & (!g1040) & (g1041) & (!g165) & (!g166)) + ((g1038) & (!g1039) & (!g1040) & (g1041) & (g165) & (g166)) + ((g1038) & (!g1039) & (g1040) & (!g1041) & (!g165) & (!g166)) + ((g1038) & (!g1039) & (g1040) & (!g1041) & (!g165) & (g166)) + ((g1038) & (!g1039) & (g1040) & (g1041) & (!g165) & (!g166)) + ((g1038) & (!g1039) & (g1040) & (g1041) & (!g165) & (g166)) + ((g1038) & (!g1039) & (g1040) & (g1041) & (g165) & (g166)) + ((g1038) & (g1039) & (!g1040) & (!g1041) & (!g165) & (!g166)) + ((g1038) & (g1039) & (!g1040) & (!g1041) & (g165) & (!g166)) + ((g1038) & (g1039) & (!g1040) & (g1041) & (!g165) & (!g166)) + ((g1038) & (g1039) & (!g1040) & (g1041) & (g165) & (!g166)) + ((g1038) & (g1039) & (!g1040) & (g1041) & (g165) & (g166)) + ((g1038) & (g1039) & (g1040) & (!g1041) & (!g165) & (!g166)) + ((g1038) & (g1039) & (g1040) & (!g1041) & (!g165) & (g166)) + ((g1038) & (g1039) & (g1040) & (!g1041) & (g165) & (!g166)) + ((g1038) & (g1039) & (g1040) & (g1041) & (!g165) & (!g166)) + ((g1038) & (g1039) & (g1040) & (g1041) & (!g165) & (g166)) + ((g1038) & (g1039) & (g1040) & (g1041) & (g165) & (!g166)) + ((g1038) & (g1039) & (g1040) & (g1041) & (g165) & (g166)));
	assign g4629 = (((!g2169) & (!g3468) & (!sk[85]) & (g1043)) + ((!g2169) & (!g3468) & (sk[85]) & (g1043)) + ((!g2169) & (g3468) & (!sk[85]) & (!g1043)) + ((!g2169) & (g3468) & (!sk[85]) & (g1043)) + ((!g2169) & (g3468) & (sk[85]) & (g1043)) + ((g2169) & (!g3468) & (!sk[85]) & (g1043)) + ((g2169) & (g3468) & (!sk[85]) & (!g1043)) + ((g2169) & (g3468) & (!sk[85]) & (g1043)) + ((g2169) & (g3468) & (sk[85]) & (!g1043)) + ((g2169) & (g3468) & (sk[85]) & (g1043)));
	assign g4630 = (((!g2170) & (!g3468) & (!sk[86]) & (g1044)) + ((!g2170) & (!g3468) & (sk[86]) & (g1044)) + ((!g2170) & (g3468) & (!sk[86]) & (!g1044)) + ((!g2170) & (g3468) & (!sk[86]) & (g1044)) + ((!g2170) & (g3468) & (sk[86]) & (g1044)) + ((g2170) & (!g3468) & (!sk[86]) & (g1044)) + ((g2170) & (g3468) & (!sk[86]) & (!g1044)) + ((g2170) & (g3468) & (!sk[86]) & (g1044)) + ((g2170) & (g3468) & (sk[86]) & (!g1044)) + ((g2170) & (g3468) & (sk[86]) & (g1044)));
	assign g4631 = (((!sk[87]) & (!g2171) & (!g3468) & (g1045)) + ((!sk[87]) & (!g2171) & (g3468) & (!g1045)) + ((!sk[87]) & (!g2171) & (g3468) & (g1045)) + ((!sk[87]) & (g2171) & (!g3468) & (g1045)) + ((!sk[87]) & (g2171) & (g3468) & (!g1045)) + ((!sk[87]) & (g2171) & (g3468) & (g1045)) + ((sk[87]) & (!g2171) & (!g3468) & (g1045)) + ((sk[87]) & (!g2171) & (g3468) & (g1045)) + ((sk[87]) & (g2171) & (g3468) & (!g1045)) + ((sk[87]) & (g2171) & (g3468) & (g1045)));
	assign g4632 = (((!g2172) & (!g3468) & (!sk[88]) & (g1046)) + ((!g2172) & (!g3468) & (sk[88]) & (g1046)) + ((!g2172) & (g3468) & (!sk[88]) & (!g1046)) + ((!g2172) & (g3468) & (!sk[88]) & (g1046)) + ((!g2172) & (g3468) & (sk[88]) & (g1046)) + ((g2172) & (!g3468) & (!sk[88]) & (g1046)) + ((g2172) & (g3468) & (!sk[88]) & (!g1046)) + ((g2172) & (g3468) & (!sk[88]) & (g1046)) + ((g2172) & (g3468) & (sk[88]) & (!g1046)) + ((g2172) & (g3468) & (sk[88]) & (g1046)));
	assign g1047 = (((!g1043) & (!g1044) & (!g1045) & (g1046) & (g165) & (g166)) + ((!g1043) & (!g1044) & (g1045) & (!g1046) & (!g165) & (g166)) + ((!g1043) & (!g1044) & (g1045) & (g1046) & (!g165) & (g166)) + ((!g1043) & (!g1044) & (g1045) & (g1046) & (g165) & (g166)) + ((!g1043) & (g1044) & (!g1045) & (!g1046) & (g165) & (!g166)) + ((!g1043) & (g1044) & (!g1045) & (g1046) & (g165) & (!g166)) + ((!g1043) & (g1044) & (!g1045) & (g1046) & (g165) & (g166)) + ((!g1043) & (g1044) & (g1045) & (!g1046) & (!g165) & (g166)) + ((!g1043) & (g1044) & (g1045) & (!g1046) & (g165) & (!g166)) + ((!g1043) & (g1044) & (g1045) & (g1046) & (!g165) & (g166)) + ((!g1043) & (g1044) & (g1045) & (g1046) & (g165) & (!g166)) + ((!g1043) & (g1044) & (g1045) & (g1046) & (g165) & (g166)) + ((g1043) & (!g1044) & (!g1045) & (!g1046) & (!g165) & (!g166)) + ((g1043) & (!g1044) & (!g1045) & (g1046) & (!g165) & (!g166)) + ((g1043) & (!g1044) & (!g1045) & (g1046) & (g165) & (g166)) + ((g1043) & (!g1044) & (g1045) & (!g1046) & (!g165) & (!g166)) + ((g1043) & (!g1044) & (g1045) & (!g1046) & (!g165) & (g166)) + ((g1043) & (!g1044) & (g1045) & (g1046) & (!g165) & (!g166)) + ((g1043) & (!g1044) & (g1045) & (g1046) & (!g165) & (g166)) + ((g1043) & (!g1044) & (g1045) & (g1046) & (g165) & (g166)) + ((g1043) & (g1044) & (!g1045) & (!g1046) & (!g165) & (!g166)) + ((g1043) & (g1044) & (!g1045) & (!g1046) & (g165) & (!g166)) + ((g1043) & (g1044) & (!g1045) & (g1046) & (!g165) & (!g166)) + ((g1043) & (g1044) & (!g1045) & (g1046) & (g165) & (!g166)) + ((g1043) & (g1044) & (!g1045) & (g1046) & (g165) & (g166)) + ((g1043) & (g1044) & (g1045) & (!g1046) & (!g165) & (!g166)) + ((g1043) & (g1044) & (g1045) & (!g1046) & (!g165) & (g166)) + ((g1043) & (g1044) & (g1045) & (!g1046) & (g165) & (!g166)) + ((g1043) & (g1044) & (g1045) & (g1046) & (!g165) & (!g166)) + ((g1043) & (g1044) & (g1045) & (g1046) & (!g165) & (g166)) + ((g1043) & (g1044) & (g1045) & (g1046) & (g165) & (!g166)) + ((g1043) & (g1044) & (g1045) & (g1046) & (g165) & (g166)));
	assign g1048 = (((!g147) & (!g148) & (!g1033) & (g1037) & (!g1042) & (!g1047)) + ((!g147) & (!g148) & (!g1033) & (g1037) & (!g1042) & (g1047)) + ((!g147) & (!g148) & (!g1033) & (g1037) & (g1042) & (!g1047)) + ((!g147) & (!g148) & (!g1033) & (g1037) & (g1042) & (g1047)) + ((!g147) & (!g148) & (g1033) & (g1037) & (!g1042) & (!g1047)) + ((!g147) & (!g148) & (g1033) & (g1037) & (!g1042) & (g1047)) + ((!g147) & (!g148) & (g1033) & (g1037) & (g1042) & (!g1047)) + ((!g147) & (!g148) & (g1033) & (g1037) & (g1042) & (g1047)) + ((!g147) & (g148) & (!g1033) & (!g1037) & (!g1042) & (g1047)) + ((!g147) & (g148) & (!g1033) & (!g1037) & (g1042) & (g1047)) + ((!g147) & (g148) & (!g1033) & (g1037) & (!g1042) & (g1047)) + ((!g147) & (g148) & (!g1033) & (g1037) & (g1042) & (g1047)) + ((!g147) & (g148) & (g1033) & (!g1037) & (!g1042) & (g1047)) + ((!g147) & (g148) & (g1033) & (!g1037) & (g1042) & (g1047)) + ((!g147) & (g148) & (g1033) & (g1037) & (!g1042) & (g1047)) + ((!g147) & (g148) & (g1033) & (g1037) & (g1042) & (g1047)) + ((g147) & (!g148) & (g1033) & (!g1037) & (!g1042) & (!g1047)) + ((g147) & (!g148) & (g1033) & (!g1037) & (!g1042) & (g1047)) + ((g147) & (!g148) & (g1033) & (!g1037) & (g1042) & (!g1047)) + ((g147) & (!g148) & (g1033) & (!g1037) & (g1042) & (g1047)) + ((g147) & (!g148) & (g1033) & (g1037) & (!g1042) & (!g1047)) + ((g147) & (!g148) & (g1033) & (g1037) & (!g1042) & (g1047)) + ((g147) & (!g148) & (g1033) & (g1037) & (g1042) & (!g1047)) + ((g147) & (!g148) & (g1033) & (g1037) & (g1042) & (g1047)) + ((g147) & (g148) & (!g1033) & (!g1037) & (g1042) & (!g1047)) + ((g147) & (g148) & (!g1033) & (!g1037) & (g1042) & (g1047)) + ((g147) & (g148) & (!g1033) & (g1037) & (g1042) & (!g1047)) + ((g147) & (g148) & (!g1033) & (g1037) & (g1042) & (g1047)) + ((g147) & (g148) & (g1033) & (!g1037) & (g1042) & (!g1047)) + ((g147) & (g148) & (g1033) & (!g1037) & (g1042) & (g1047)) + ((g147) & (g148) & (g1033) & (g1037) & (g1042) & (!g1047)) + ((g147) & (g148) & (g1033) & (g1037) & (g1042) & (g1047)));
	assign g1049 = (((!g142) & (!sk[91]) & (!g1028) & (g1048)) + ((!g142) & (!sk[91]) & (g1028) & (!g1048)) + ((!g142) & (!sk[91]) & (g1028) & (g1048)) + ((!g142) & (sk[91]) & (!g1028) & (g1048)) + ((!g142) & (sk[91]) & (g1028) & (g1048)) + ((g142) & (!sk[91]) & (!g1028) & (g1048)) + ((g142) & (!sk[91]) & (g1028) & (!g1048)) + ((g142) & (!sk[91]) & (g1028) & (g1048)) + ((g142) & (sk[91]) & (g1028) & (!g1048)) + ((g142) & (sk[91]) & (g1028) & (g1048)));
	assign g4633 = (((!g2059) & (!g2624) & (!sk[92]) & (g1050)) + ((!g2059) & (!g2624) & (sk[92]) & (g1050)) + ((!g2059) & (g2624) & (!sk[92]) & (!g1050)) + ((!g2059) & (g2624) & (!sk[92]) & (g1050)) + ((!g2059) & (g2624) & (sk[92]) & (g1050)) + ((g2059) & (!g2624) & (!sk[92]) & (g1050)) + ((g2059) & (g2624) & (!sk[92]) & (!g1050)) + ((g2059) & (g2624) & (!sk[92]) & (g1050)) + ((g2059) & (g2624) & (sk[92]) & (!g1050)) + ((g2059) & (g2624) & (sk[92]) & (g1050)));
	assign g1051 = (((!g1004) & (!g1006) & (!sk[93]) & (g916)) + ((!g1004) & (g1006) & (!sk[93]) & (!g916)) + ((!g1004) & (g1006) & (!sk[93]) & (g916)) + ((!g1004) & (g1006) & (sk[93]) & (!g916)) + ((g1004) & (!g1006) & (!sk[93]) & (g916)) + ((g1004) & (!g1006) & (sk[93]) & (!g916)) + ((g1004) & (g1006) & (!sk[93]) & (!g916)) + ((g1004) & (g1006) & (!sk[93]) & (g916)) + ((g1004) & (g1006) & (sk[93]) & (!g916)) + ((g1004) & (g1006) & (sk[93]) & (g916)));
	assign g1052 = (((!g126) & (!g1049) & (!g1050) & (!sk[94]) & (g1051) & (!g916)) + ((!g126) & (!g1049) & (!g1050) & (!sk[94]) & (g1051) & (g916)) + ((!g126) & (!g1049) & (g1050) & (!sk[94]) & (!g1051) & (!g916)) + ((!g126) & (!g1049) & (g1050) & (!sk[94]) & (!g1051) & (g916)) + ((!g126) & (!g1049) & (g1050) & (!sk[94]) & (g1051) & (!g916)) + ((!g126) & (!g1049) & (g1050) & (!sk[94]) & (g1051) & (g916)) + ((!g126) & (!g1049) & (g1050) & (sk[94]) & (!g1051) & (!g916)) + ((!g126) & (!g1049) & (g1050) & (sk[94]) & (!g1051) & (g916)) + ((!g126) & (!g1049) & (g1050) & (sk[94]) & (g1051) & (!g916)) + ((!g126) & (!g1049) & (g1050) & (sk[94]) & (g1051) & (g916)) + ((!g126) & (g1049) & (!g1050) & (!sk[94]) & (!g1051) & (!g916)) + ((!g126) & (g1049) & (!g1050) & (!sk[94]) & (!g1051) & (g916)) + ((!g126) & (g1049) & (!g1050) & (!sk[94]) & (g1051) & (!g916)) + ((!g126) & (g1049) & (!g1050) & (!sk[94]) & (g1051) & (g916)) + ((!g126) & (g1049) & (g1050) & (!sk[94]) & (!g1051) & (!g916)) + ((!g126) & (g1049) & (g1050) & (!sk[94]) & (!g1051) & (g916)) + ((!g126) & (g1049) & (g1050) & (!sk[94]) & (g1051) & (!g916)) + ((!g126) & (g1049) & (g1050) & (!sk[94]) & (g1051) & (g916)) + ((!g126) & (g1049) & (g1050) & (sk[94]) & (!g1051) & (!g916)) + ((!g126) & (g1049) & (g1050) & (sk[94]) & (!g1051) & (g916)) + ((!g126) & (g1049) & (g1050) & (sk[94]) & (g1051) & (!g916)) + ((!g126) & (g1049) & (g1050) & (sk[94]) & (g1051) & (g916)) + ((g126) & (!g1049) & (!g1050) & (!sk[94]) & (g1051) & (!g916)) + ((g126) & (!g1049) & (!g1050) & (!sk[94]) & (g1051) & (g916)) + ((g126) & (!g1049) & (!g1050) & (sk[94]) & (!g1051) & (!g916)) + ((g126) & (!g1049) & (!g1050) & (sk[94]) & (g1051) & (g916)) + ((g126) & (!g1049) & (g1050) & (!sk[94]) & (!g1051) & (!g916)) + ((g126) & (!g1049) & (g1050) & (!sk[94]) & (!g1051) & (g916)) + ((g126) & (!g1049) & (g1050) & (!sk[94]) & (g1051) & (!g916)) + ((g126) & (!g1049) & (g1050) & (!sk[94]) & (g1051) & (g916)) + ((g126) & (!g1049) & (g1050) & (sk[94]) & (!g1051) & (!g916)) + ((g126) & (!g1049) & (g1050) & (sk[94]) & (g1051) & (g916)) + ((g126) & (g1049) & (!g1050) & (!sk[94]) & (!g1051) & (!g916)) + ((g126) & (g1049) & (!g1050) & (!sk[94]) & (!g1051) & (g916)) + ((g126) & (g1049) & (!g1050) & (!sk[94]) & (g1051) & (!g916)) + ((g126) & (g1049) & (!g1050) & (!sk[94]) & (g1051) & (g916)) + ((g126) & (g1049) & (!g1050) & (sk[94]) & (!g1051) & (g916)) + ((g126) & (g1049) & (!g1050) & (sk[94]) & (g1051) & (!g916)) + ((g126) & (g1049) & (g1050) & (!sk[94]) & (!g1051) & (!g916)) + ((g126) & (g1049) & (g1050) & (!sk[94]) & (!g1051) & (g916)) + ((g126) & (g1049) & (g1050) & (!sk[94]) & (g1051) & (!g916)) + ((g126) & (g1049) & (g1050) & (!sk[94]) & (g1051) & (g916)) + ((g126) & (g1049) & (g1050) & (sk[94]) & (!g1051) & (g916)) + ((g126) & (g1049) & (g1050) & (sk[94]) & (g1051) & (!g916)));
	assign g4634 = (((!sk[95]) & (!g2140) & (!g3444) & (g1053)) + ((!sk[95]) & (!g2140) & (g3444) & (!g1053)) + ((!sk[95]) & (!g2140) & (g3444) & (g1053)) + ((!sk[95]) & (g2140) & (!g3444) & (g1053)) + ((!sk[95]) & (g2140) & (g3444) & (!g1053)) + ((!sk[95]) & (g2140) & (g3444) & (g1053)) + ((sk[95]) & (!g2140) & (!g3444) & (g1053)) + ((sk[95]) & (!g2140) & (g3444) & (g1053)) + ((sk[95]) & (g2140) & (g3444) & (!g1053)) + ((sk[95]) & (g2140) & (g3444) & (g1053)));
	assign g4635 = (((!sk[96]) & (!g2142) & (!g3444) & (g1054)) + ((!sk[96]) & (!g2142) & (g3444) & (!g1054)) + ((!sk[96]) & (!g2142) & (g3444) & (g1054)) + ((!sk[96]) & (g2142) & (!g3444) & (g1054)) + ((!sk[96]) & (g2142) & (g3444) & (!g1054)) + ((!sk[96]) & (g2142) & (g3444) & (g1054)) + ((sk[96]) & (!g2142) & (!g3444) & (g1054)) + ((sk[96]) & (!g2142) & (g3444) & (g1054)) + ((sk[96]) & (g2142) & (g3444) & (!g1054)) + ((sk[96]) & (g2142) & (g3444) & (g1054)));
	assign g4636 = (((!g2144) & (!sk[97]) & (!g3444) & (g1055)) + ((!g2144) & (!sk[97]) & (g3444) & (!g1055)) + ((!g2144) & (!sk[97]) & (g3444) & (g1055)) + ((!g2144) & (sk[97]) & (!g3444) & (g1055)) + ((!g2144) & (sk[97]) & (g3444) & (g1055)) + ((g2144) & (!sk[97]) & (!g3444) & (g1055)) + ((g2144) & (!sk[97]) & (g3444) & (!g1055)) + ((g2144) & (!sk[97]) & (g3444) & (g1055)) + ((g2144) & (sk[97]) & (g3444) & (!g1055)) + ((g2144) & (sk[97]) & (g3444) & (g1055)));
	assign g4637 = (((!sk[98]) & (!g2145) & (!g3444) & (g1056)) + ((!sk[98]) & (!g2145) & (g3444) & (!g1056)) + ((!sk[98]) & (!g2145) & (g3444) & (g1056)) + ((!sk[98]) & (g2145) & (!g3444) & (g1056)) + ((!sk[98]) & (g2145) & (g3444) & (!g1056)) + ((!sk[98]) & (g2145) & (g3444) & (g1056)) + ((sk[98]) & (!g2145) & (!g3444) & (g1056)) + ((sk[98]) & (!g2145) & (g3444) & (g1056)) + ((sk[98]) & (g2145) & (g3444) & (!g1056)) + ((sk[98]) & (g2145) & (g3444) & (g1056)));
	assign g1057 = (((!g1053) & (!g1054) & (!g1055) & (g1056) & (g147) & (g148)) + ((!g1053) & (!g1054) & (g1055) & (!g1056) & (!g147) & (g148)) + ((!g1053) & (!g1054) & (g1055) & (g1056) & (!g147) & (g148)) + ((!g1053) & (!g1054) & (g1055) & (g1056) & (g147) & (g148)) + ((!g1053) & (g1054) & (!g1055) & (!g1056) & (g147) & (!g148)) + ((!g1053) & (g1054) & (!g1055) & (g1056) & (g147) & (!g148)) + ((!g1053) & (g1054) & (!g1055) & (g1056) & (g147) & (g148)) + ((!g1053) & (g1054) & (g1055) & (!g1056) & (!g147) & (g148)) + ((!g1053) & (g1054) & (g1055) & (!g1056) & (g147) & (!g148)) + ((!g1053) & (g1054) & (g1055) & (g1056) & (!g147) & (g148)) + ((!g1053) & (g1054) & (g1055) & (g1056) & (g147) & (!g148)) + ((!g1053) & (g1054) & (g1055) & (g1056) & (g147) & (g148)) + ((g1053) & (!g1054) & (!g1055) & (!g1056) & (!g147) & (!g148)) + ((g1053) & (!g1054) & (!g1055) & (g1056) & (!g147) & (!g148)) + ((g1053) & (!g1054) & (!g1055) & (g1056) & (g147) & (g148)) + ((g1053) & (!g1054) & (g1055) & (!g1056) & (!g147) & (!g148)) + ((g1053) & (!g1054) & (g1055) & (!g1056) & (!g147) & (g148)) + ((g1053) & (!g1054) & (g1055) & (g1056) & (!g147) & (!g148)) + ((g1053) & (!g1054) & (g1055) & (g1056) & (!g147) & (g148)) + ((g1053) & (!g1054) & (g1055) & (g1056) & (g147) & (g148)) + ((g1053) & (g1054) & (!g1055) & (!g1056) & (!g147) & (!g148)) + ((g1053) & (g1054) & (!g1055) & (!g1056) & (g147) & (!g148)) + ((g1053) & (g1054) & (!g1055) & (g1056) & (!g147) & (!g148)) + ((g1053) & (g1054) & (!g1055) & (g1056) & (g147) & (!g148)) + ((g1053) & (g1054) & (!g1055) & (g1056) & (g147) & (g148)) + ((g1053) & (g1054) & (g1055) & (!g1056) & (!g147) & (!g148)) + ((g1053) & (g1054) & (g1055) & (!g1056) & (!g147) & (g148)) + ((g1053) & (g1054) & (g1055) & (!g1056) & (g147) & (!g148)) + ((g1053) & (g1054) & (g1055) & (g1056) & (!g147) & (!g148)) + ((g1053) & (g1054) & (g1055) & (g1056) & (!g147) & (g148)) + ((g1053) & (g1054) & (g1055) & (g1056) & (g147) & (!g148)) + ((g1053) & (g1054) & (g1055) & (g1056) & (g147) & (g148)));
	assign g4638 = (((!g2146) & (!g3444) & (!sk[100]) & (g1058)) + ((!g2146) & (!g3444) & (sk[100]) & (g1058)) + ((!g2146) & (g3444) & (!sk[100]) & (!g1058)) + ((!g2146) & (g3444) & (!sk[100]) & (g1058)) + ((!g2146) & (g3444) & (sk[100]) & (g1058)) + ((g2146) & (!g3444) & (!sk[100]) & (g1058)) + ((g2146) & (g3444) & (!sk[100]) & (!g1058)) + ((g2146) & (g3444) & (!sk[100]) & (g1058)) + ((g2146) & (g3444) & (sk[100]) & (!g1058)) + ((g2146) & (g3444) & (sk[100]) & (g1058)));
	assign g4639 = (((!g2148) & (!g3444) & (!sk[101]) & (g1059)) + ((!g2148) & (!g3444) & (sk[101]) & (g1059)) + ((!g2148) & (g3444) & (!sk[101]) & (!g1059)) + ((!g2148) & (g3444) & (!sk[101]) & (g1059)) + ((!g2148) & (g3444) & (sk[101]) & (g1059)) + ((g2148) & (!g3444) & (!sk[101]) & (g1059)) + ((g2148) & (g3444) & (!sk[101]) & (!g1059)) + ((g2148) & (g3444) & (!sk[101]) & (g1059)) + ((g2148) & (g3444) & (sk[101]) & (!g1059)) + ((g2148) & (g3444) & (sk[101]) & (g1059)));
	assign g4640 = (((!g2150) & (!sk[102]) & (!g3444) & (g1060)) + ((!g2150) & (!sk[102]) & (g3444) & (!g1060)) + ((!g2150) & (!sk[102]) & (g3444) & (g1060)) + ((!g2150) & (sk[102]) & (!g3444) & (g1060)) + ((!g2150) & (sk[102]) & (g3444) & (g1060)) + ((g2150) & (!sk[102]) & (!g3444) & (g1060)) + ((g2150) & (!sk[102]) & (g3444) & (!g1060)) + ((g2150) & (!sk[102]) & (g3444) & (g1060)) + ((g2150) & (sk[102]) & (g3444) & (!g1060)) + ((g2150) & (sk[102]) & (g3444) & (g1060)));
	assign g4641 = (((!sk[103]) & (!g2151) & (!g3444) & (g1061)) + ((!sk[103]) & (!g2151) & (g3444) & (!g1061)) + ((!sk[103]) & (!g2151) & (g3444) & (g1061)) + ((!sk[103]) & (g2151) & (!g3444) & (g1061)) + ((!sk[103]) & (g2151) & (g3444) & (!g1061)) + ((!sk[103]) & (g2151) & (g3444) & (g1061)) + ((sk[103]) & (!g2151) & (!g3444) & (g1061)) + ((sk[103]) & (!g2151) & (g3444) & (g1061)) + ((sk[103]) & (g2151) & (g3444) & (!g1061)) + ((sk[103]) & (g2151) & (g3444) & (g1061)));
	assign g1062 = (((!g1058) & (!g1059) & (!g1060) & (g1061) & (g147) & (g148)) + ((!g1058) & (!g1059) & (g1060) & (!g1061) & (!g147) & (g148)) + ((!g1058) & (!g1059) & (g1060) & (g1061) & (!g147) & (g148)) + ((!g1058) & (!g1059) & (g1060) & (g1061) & (g147) & (g148)) + ((!g1058) & (g1059) & (!g1060) & (!g1061) & (g147) & (!g148)) + ((!g1058) & (g1059) & (!g1060) & (g1061) & (g147) & (!g148)) + ((!g1058) & (g1059) & (!g1060) & (g1061) & (g147) & (g148)) + ((!g1058) & (g1059) & (g1060) & (!g1061) & (!g147) & (g148)) + ((!g1058) & (g1059) & (g1060) & (!g1061) & (g147) & (!g148)) + ((!g1058) & (g1059) & (g1060) & (g1061) & (!g147) & (g148)) + ((!g1058) & (g1059) & (g1060) & (g1061) & (g147) & (!g148)) + ((!g1058) & (g1059) & (g1060) & (g1061) & (g147) & (g148)) + ((g1058) & (!g1059) & (!g1060) & (!g1061) & (!g147) & (!g148)) + ((g1058) & (!g1059) & (!g1060) & (g1061) & (!g147) & (!g148)) + ((g1058) & (!g1059) & (!g1060) & (g1061) & (g147) & (g148)) + ((g1058) & (!g1059) & (g1060) & (!g1061) & (!g147) & (!g148)) + ((g1058) & (!g1059) & (g1060) & (!g1061) & (!g147) & (g148)) + ((g1058) & (!g1059) & (g1060) & (g1061) & (!g147) & (!g148)) + ((g1058) & (!g1059) & (g1060) & (g1061) & (!g147) & (g148)) + ((g1058) & (!g1059) & (g1060) & (g1061) & (g147) & (g148)) + ((g1058) & (g1059) & (!g1060) & (!g1061) & (!g147) & (!g148)) + ((g1058) & (g1059) & (!g1060) & (!g1061) & (g147) & (!g148)) + ((g1058) & (g1059) & (!g1060) & (g1061) & (!g147) & (!g148)) + ((g1058) & (g1059) & (!g1060) & (g1061) & (g147) & (!g148)) + ((g1058) & (g1059) & (!g1060) & (g1061) & (g147) & (g148)) + ((g1058) & (g1059) & (g1060) & (!g1061) & (!g147) & (!g148)) + ((g1058) & (g1059) & (g1060) & (!g1061) & (!g147) & (g148)) + ((g1058) & (g1059) & (g1060) & (!g1061) & (g147) & (!g148)) + ((g1058) & (g1059) & (g1060) & (g1061) & (!g147) & (!g148)) + ((g1058) & (g1059) & (g1060) & (g1061) & (!g147) & (g148)) + ((g1058) & (g1059) & (g1060) & (g1061) & (g147) & (!g148)) + ((g1058) & (g1059) & (g1060) & (g1061) & (g147) & (g148)));
	assign g4642 = (((!sk[105]) & (!g2152) & (!g3444) & (g1063)) + ((!sk[105]) & (!g2152) & (g3444) & (!g1063)) + ((!sk[105]) & (!g2152) & (g3444) & (g1063)) + ((!sk[105]) & (g2152) & (!g3444) & (g1063)) + ((!sk[105]) & (g2152) & (g3444) & (!g1063)) + ((!sk[105]) & (g2152) & (g3444) & (g1063)) + ((sk[105]) & (!g2152) & (!g3444) & (g1063)) + ((sk[105]) & (!g2152) & (g3444) & (g1063)) + ((sk[105]) & (g2152) & (g3444) & (!g1063)) + ((sk[105]) & (g2152) & (g3444) & (g1063)));
	assign g4643 = (((!sk[106]) & (!g2153) & (!g3444) & (g1064)) + ((!sk[106]) & (!g2153) & (g3444) & (!g1064)) + ((!sk[106]) & (!g2153) & (g3444) & (g1064)) + ((!sk[106]) & (g2153) & (!g3444) & (g1064)) + ((!sk[106]) & (g2153) & (g3444) & (!g1064)) + ((!sk[106]) & (g2153) & (g3444) & (g1064)) + ((sk[106]) & (!g2153) & (!g3444) & (g1064)) + ((sk[106]) & (!g2153) & (g3444) & (g1064)) + ((sk[106]) & (g2153) & (g3444) & (!g1064)) + ((sk[106]) & (g2153) & (g3444) & (g1064)));
	assign g4644 = (((!sk[107]) & (!g2155) & (!g3444) & (g1065)) + ((!sk[107]) & (!g2155) & (g3444) & (!g1065)) + ((!sk[107]) & (!g2155) & (g3444) & (g1065)) + ((!sk[107]) & (g2155) & (!g3444) & (g1065)) + ((!sk[107]) & (g2155) & (g3444) & (!g1065)) + ((!sk[107]) & (g2155) & (g3444) & (g1065)) + ((sk[107]) & (!g2155) & (!g3444) & (g1065)) + ((sk[107]) & (!g2155) & (g3444) & (g1065)) + ((sk[107]) & (g2155) & (g3444) & (!g1065)) + ((sk[107]) & (g2155) & (g3444) & (g1065)));
	assign g4645 = (((!g2157) & (!sk[108]) & (!g3444) & (g1066)) + ((!g2157) & (!sk[108]) & (g3444) & (!g1066)) + ((!g2157) & (!sk[108]) & (g3444) & (g1066)) + ((!g2157) & (sk[108]) & (!g3444) & (g1066)) + ((!g2157) & (sk[108]) & (g3444) & (g1066)) + ((g2157) & (!sk[108]) & (!g3444) & (g1066)) + ((g2157) & (!sk[108]) & (g3444) & (!g1066)) + ((g2157) & (!sk[108]) & (g3444) & (g1066)) + ((g2157) & (sk[108]) & (g3444) & (!g1066)) + ((g2157) & (sk[108]) & (g3444) & (g1066)));
	assign g1067 = (((!g1063) & (!g1064) & (!g1065) & (g1066) & (g147) & (g148)) + ((!g1063) & (!g1064) & (g1065) & (!g1066) & (!g147) & (g148)) + ((!g1063) & (!g1064) & (g1065) & (g1066) & (!g147) & (g148)) + ((!g1063) & (!g1064) & (g1065) & (g1066) & (g147) & (g148)) + ((!g1063) & (g1064) & (!g1065) & (!g1066) & (g147) & (!g148)) + ((!g1063) & (g1064) & (!g1065) & (g1066) & (g147) & (!g148)) + ((!g1063) & (g1064) & (!g1065) & (g1066) & (g147) & (g148)) + ((!g1063) & (g1064) & (g1065) & (!g1066) & (!g147) & (g148)) + ((!g1063) & (g1064) & (g1065) & (!g1066) & (g147) & (!g148)) + ((!g1063) & (g1064) & (g1065) & (g1066) & (!g147) & (g148)) + ((!g1063) & (g1064) & (g1065) & (g1066) & (g147) & (!g148)) + ((!g1063) & (g1064) & (g1065) & (g1066) & (g147) & (g148)) + ((g1063) & (!g1064) & (!g1065) & (!g1066) & (!g147) & (!g148)) + ((g1063) & (!g1064) & (!g1065) & (g1066) & (!g147) & (!g148)) + ((g1063) & (!g1064) & (!g1065) & (g1066) & (g147) & (g148)) + ((g1063) & (!g1064) & (g1065) & (!g1066) & (!g147) & (!g148)) + ((g1063) & (!g1064) & (g1065) & (!g1066) & (!g147) & (g148)) + ((g1063) & (!g1064) & (g1065) & (g1066) & (!g147) & (!g148)) + ((g1063) & (!g1064) & (g1065) & (g1066) & (!g147) & (g148)) + ((g1063) & (!g1064) & (g1065) & (g1066) & (g147) & (g148)) + ((g1063) & (g1064) & (!g1065) & (!g1066) & (!g147) & (!g148)) + ((g1063) & (g1064) & (!g1065) & (!g1066) & (g147) & (!g148)) + ((g1063) & (g1064) & (!g1065) & (g1066) & (!g147) & (!g148)) + ((g1063) & (g1064) & (!g1065) & (g1066) & (g147) & (!g148)) + ((g1063) & (g1064) & (!g1065) & (g1066) & (g147) & (g148)) + ((g1063) & (g1064) & (g1065) & (!g1066) & (!g147) & (!g148)) + ((g1063) & (g1064) & (g1065) & (!g1066) & (!g147) & (g148)) + ((g1063) & (g1064) & (g1065) & (!g1066) & (g147) & (!g148)) + ((g1063) & (g1064) & (g1065) & (g1066) & (!g147) & (!g148)) + ((g1063) & (g1064) & (g1065) & (g1066) & (!g147) & (g148)) + ((g1063) & (g1064) & (g1065) & (g1066) & (g147) & (!g148)) + ((g1063) & (g1064) & (g1065) & (g1066) & (g147) & (g148)));
	assign g4646 = (((!g2158) & (!g3444) & (!sk[110]) & (g1068)) + ((!g2158) & (!g3444) & (sk[110]) & (g1068)) + ((!g2158) & (g3444) & (!sk[110]) & (!g1068)) + ((!g2158) & (g3444) & (!sk[110]) & (g1068)) + ((!g2158) & (g3444) & (sk[110]) & (g1068)) + ((g2158) & (!g3444) & (!sk[110]) & (g1068)) + ((g2158) & (g3444) & (!sk[110]) & (!g1068)) + ((g2158) & (g3444) & (!sk[110]) & (g1068)) + ((g2158) & (g3444) & (sk[110]) & (!g1068)) + ((g2158) & (g3444) & (sk[110]) & (g1068)));
	assign g4647 = (((!g2159) & (!sk[111]) & (!g3444) & (g1069)) + ((!g2159) & (!sk[111]) & (g3444) & (!g1069)) + ((!g2159) & (!sk[111]) & (g3444) & (g1069)) + ((!g2159) & (sk[111]) & (!g3444) & (g1069)) + ((!g2159) & (sk[111]) & (g3444) & (g1069)) + ((g2159) & (!sk[111]) & (!g3444) & (g1069)) + ((g2159) & (!sk[111]) & (g3444) & (!g1069)) + ((g2159) & (!sk[111]) & (g3444) & (g1069)) + ((g2159) & (sk[111]) & (g3444) & (!g1069)) + ((g2159) & (sk[111]) & (g3444) & (g1069)));
	assign g4648 = (((!sk[112]) & (!g2160) & (!g3444) & (g1070)) + ((!sk[112]) & (!g2160) & (g3444) & (!g1070)) + ((!sk[112]) & (!g2160) & (g3444) & (g1070)) + ((!sk[112]) & (g2160) & (!g3444) & (g1070)) + ((!sk[112]) & (g2160) & (g3444) & (!g1070)) + ((!sk[112]) & (g2160) & (g3444) & (g1070)) + ((sk[112]) & (!g2160) & (!g3444) & (g1070)) + ((sk[112]) & (!g2160) & (g3444) & (g1070)) + ((sk[112]) & (g2160) & (g3444) & (!g1070)) + ((sk[112]) & (g2160) & (g3444) & (g1070)));
	assign g4649 = (((!g2161) & (!g3444) & (!sk[113]) & (g1071)) + ((!g2161) & (!g3444) & (sk[113]) & (g1071)) + ((!g2161) & (g3444) & (!sk[113]) & (!g1071)) + ((!g2161) & (g3444) & (!sk[113]) & (g1071)) + ((!g2161) & (g3444) & (sk[113]) & (g1071)) + ((g2161) & (!g3444) & (!sk[113]) & (g1071)) + ((g2161) & (g3444) & (!sk[113]) & (!g1071)) + ((g2161) & (g3444) & (!sk[113]) & (g1071)) + ((g2161) & (g3444) & (sk[113]) & (!g1071)) + ((g2161) & (g3444) & (sk[113]) & (g1071)));
	assign g1072 = (((!g1068) & (!g1069) & (!g1070) & (g1071) & (g147) & (g148)) + ((!g1068) & (!g1069) & (g1070) & (!g1071) & (!g147) & (g148)) + ((!g1068) & (!g1069) & (g1070) & (g1071) & (!g147) & (g148)) + ((!g1068) & (!g1069) & (g1070) & (g1071) & (g147) & (g148)) + ((!g1068) & (g1069) & (!g1070) & (!g1071) & (g147) & (!g148)) + ((!g1068) & (g1069) & (!g1070) & (g1071) & (g147) & (!g148)) + ((!g1068) & (g1069) & (!g1070) & (g1071) & (g147) & (g148)) + ((!g1068) & (g1069) & (g1070) & (!g1071) & (!g147) & (g148)) + ((!g1068) & (g1069) & (g1070) & (!g1071) & (g147) & (!g148)) + ((!g1068) & (g1069) & (g1070) & (g1071) & (!g147) & (g148)) + ((!g1068) & (g1069) & (g1070) & (g1071) & (g147) & (!g148)) + ((!g1068) & (g1069) & (g1070) & (g1071) & (g147) & (g148)) + ((g1068) & (!g1069) & (!g1070) & (!g1071) & (!g147) & (!g148)) + ((g1068) & (!g1069) & (!g1070) & (g1071) & (!g147) & (!g148)) + ((g1068) & (!g1069) & (!g1070) & (g1071) & (g147) & (g148)) + ((g1068) & (!g1069) & (g1070) & (!g1071) & (!g147) & (!g148)) + ((g1068) & (!g1069) & (g1070) & (!g1071) & (!g147) & (g148)) + ((g1068) & (!g1069) & (g1070) & (g1071) & (!g147) & (!g148)) + ((g1068) & (!g1069) & (g1070) & (g1071) & (!g147) & (g148)) + ((g1068) & (!g1069) & (g1070) & (g1071) & (g147) & (g148)) + ((g1068) & (g1069) & (!g1070) & (!g1071) & (!g147) & (!g148)) + ((g1068) & (g1069) & (!g1070) & (!g1071) & (g147) & (!g148)) + ((g1068) & (g1069) & (!g1070) & (g1071) & (!g147) & (!g148)) + ((g1068) & (g1069) & (!g1070) & (g1071) & (g147) & (!g148)) + ((g1068) & (g1069) & (!g1070) & (g1071) & (g147) & (g148)) + ((g1068) & (g1069) & (g1070) & (!g1071) & (!g147) & (!g148)) + ((g1068) & (g1069) & (g1070) & (!g1071) & (!g147) & (g148)) + ((g1068) & (g1069) & (g1070) & (!g1071) & (g147) & (!g148)) + ((g1068) & (g1069) & (g1070) & (g1071) & (!g147) & (!g148)) + ((g1068) & (g1069) & (g1070) & (g1071) & (!g147) & (g148)) + ((g1068) & (g1069) & (g1070) & (g1071) & (g147) & (!g148)) + ((g1068) & (g1069) & (g1070) & (g1071) & (g147) & (g148)));
	assign g1073 = (((!g1057) & (!g1062) & (!g1067) & (g1072) & (g165) & (g166)) + ((!g1057) & (!g1062) & (g1067) & (!g1072) & (!g165) & (g166)) + ((!g1057) & (!g1062) & (g1067) & (g1072) & (!g165) & (g166)) + ((!g1057) & (!g1062) & (g1067) & (g1072) & (g165) & (g166)) + ((!g1057) & (g1062) & (!g1067) & (!g1072) & (g165) & (!g166)) + ((!g1057) & (g1062) & (!g1067) & (g1072) & (g165) & (!g166)) + ((!g1057) & (g1062) & (!g1067) & (g1072) & (g165) & (g166)) + ((!g1057) & (g1062) & (g1067) & (!g1072) & (!g165) & (g166)) + ((!g1057) & (g1062) & (g1067) & (!g1072) & (g165) & (!g166)) + ((!g1057) & (g1062) & (g1067) & (g1072) & (!g165) & (g166)) + ((!g1057) & (g1062) & (g1067) & (g1072) & (g165) & (!g166)) + ((!g1057) & (g1062) & (g1067) & (g1072) & (g165) & (g166)) + ((g1057) & (!g1062) & (!g1067) & (!g1072) & (!g165) & (!g166)) + ((g1057) & (!g1062) & (!g1067) & (g1072) & (!g165) & (!g166)) + ((g1057) & (!g1062) & (!g1067) & (g1072) & (g165) & (g166)) + ((g1057) & (!g1062) & (g1067) & (!g1072) & (!g165) & (!g166)) + ((g1057) & (!g1062) & (g1067) & (!g1072) & (!g165) & (g166)) + ((g1057) & (!g1062) & (g1067) & (g1072) & (!g165) & (!g166)) + ((g1057) & (!g1062) & (g1067) & (g1072) & (!g165) & (g166)) + ((g1057) & (!g1062) & (g1067) & (g1072) & (g165) & (g166)) + ((g1057) & (g1062) & (!g1067) & (!g1072) & (!g165) & (!g166)) + ((g1057) & (g1062) & (!g1067) & (!g1072) & (g165) & (!g166)) + ((g1057) & (g1062) & (!g1067) & (g1072) & (!g165) & (!g166)) + ((g1057) & (g1062) & (!g1067) & (g1072) & (g165) & (!g166)) + ((g1057) & (g1062) & (!g1067) & (g1072) & (g165) & (g166)) + ((g1057) & (g1062) & (g1067) & (!g1072) & (!g165) & (!g166)) + ((g1057) & (g1062) & (g1067) & (!g1072) & (!g165) & (g166)) + ((g1057) & (g1062) & (g1067) & (!g1072) & (g165) & (!g166)) + ((g1057) & (g1062) & (g1067) & (g1072) & (!g165) & (!g166)) + ((g1057) & (g1062) & (g1067) & (g1072) & (!g165) & (g166)) + ((g1057) & (g1062) & (g1067) & (g1072) & (g165) & (!g166)) + ((g1057) & (g1062) & (g1067) & (g1072) & (g165) & (g166)));
	assign g4650 = (((!g2173) & (!sk[116]) & (!g3444) & (g1074)) + ((!g2173) & (!sk[116]) & (g3444) & (!g1074)) + ((!g2173) & (!sk[116]) & (g3444) & (g1074)) + ((!g2173) & (sk[116]) & (!g3444) & (g1074)) + ((!g2173) & (sk[116]) & (g3444) & (g1074)) + ((g2173) & (!sk[116]) & (!g3444) & (g1074)) + ((g2173) & (!sk[116]) & (g3444) & (!g1074)) + ((g2173) & (!sk[116]) & (g3444) & (g1074)) + ((g2173) & (sk[116]) & (g3444) & (!g1074)) + ((g2173) & (sk[116]) & (g3444) & (g1074)));
	assign g4651 = (((!g2174) & (!g3444) & (!sk[117]) & (g1075)) + ((!g2174) & (!g3444) & (sk[117]) & (g1075)) + ((!g2174) & (g3444) & (!sk[117]) & (!g1075)) + ((!g2174) & (g3444) & (!sk[117]) & (g1075)) + ((!g2174) & (g3444) & (sk[117]) & (g1075)) + ((g2174) & (!g3444) & (!sk[117]) & (g1075)) + ((g2174) & (g3444) & (!sk[117]) & (!g1075)) + ((g2174) & (g3444) & (!sk[117]) & (g1075)) + ((g2174) & (g3444) & (sk[117]) & (!g1075)) + ((g2174) & (g3444) & (sk[117]) & (g1075)));
	assign g4652 = (((!g2175) & (!sk[118]) & (!g3444) & (g1076)) + ((!g2175) & (!sk[118]) & (g3444) & (!g1076)) + ((!g2175) & (!sk[118]) & (g3444) & (g1076)) + ((!g2175) & (sk[118]) & (!g3444) & (g1076)) + ((!g2175) & (sk[118]) & (g3444) & (g1076)) + ((g2175) & (!sk[118]) & (!g3444) & (g1076)) + ((g2175) & (!sk[118]) & (g3444) & (!g1076)) + ((g2175) & (!sk[118]) & (g3444) & (g1076)) + ((g2175) & (sk[118]) & (g3444) & (!g1076)) + ((g2175) & (sk[118]) & (g3444) & (g1076)));
	assign g4653 = (((!sk[119]) & (!g2176) & (!g3444) & (g1077)) + ((!sk[119]) & (!g2176) & (g3444) & (!g1077)) + ((!sk[119]) & (!g2176) & (g3444) & (g1077)) + ((!sk[119]) & (g2176) & (!g3444) & (g1077)) + ((!sk[119]) & (g2176) & (g3444) & (!g1077)) + ((!sk[119]) & (g2176) & (g3444) & (g1077)) + ((sk[119]) & (!g2176) & (!g3444) & (g1077)) + ((sk[119]) & (!g2176) & (g3444) & (g1077)) + ((sk[119]) & (g2176) & (g3444) & (!g1077)) + ((sk[119]) & (g2176) & (g3444) & (g1077)));
	assign g1078 = (((!g1074) & (!g1075) & (!g1076) & (g1077) & (g165) & (g166)) + ((!g1074) & (!g1075) & (g1076) & (!g1077) & (!g165) & (g166)) + ((!g1074) & (!g1075) & (g1076) & (g1077) & (!g165) & (g166)) + ((!g1074) & (!g1075) & (g1076) & (g1077) & (g165) & (g166)) + ((!g1074) & (g1075) & (!g1076) & (!g1077) & (g165) & (!g166)) + ((!g1074) & (g1075) & (!g1076) & (g1077) & (g165) & (!g166)) + ((!g1074) & (g1075) & (!g1076) & (g1077) & (g165) & (g166)) + ((!g1074) & (g1075) & (g1076) & (!g1077) & (!g165) & (g166)) + ((!g1074) & (g1075) & (g1076) & (!g1077) & (g165) & (!g166)) + ((!g1074) & (g1075) & (g1076) & (g1077) & (!g165) & (g166)) + ((!g1074) & (g1075) & (g1076) & (g1077) & (g165) & (!g166)) + ((!g1074) & (g1075) & (g1076) & (g1077) & (g165) & (g166)) + ((g1074) & (!g1075) & (!g1076) & (!g1077) & (!g165) & (!g166)) + ((g1074) & (!g1075) & (!g1076) & (g1077) & (!g165) & (!g166)) + ((g1074) & (!g1075) & (!g1076) & (g1077) & (g165) & (g166)) + ((g1074) & (!g1075) & (g1076) & (!g1077) & (!g165) & (!g166)) + ((g1074) & (!g1075) & (g1076) & (!g1077) & (!g165) & (g166)) + ((g1074) & (!g1075) & (g1076) & (g1077) & (!g165) & (!g166)) + ((g1074) & (!g1075) & (g1076) & (g1077) & (!g165) & (g166)) + ((g1074) & (!g1075) & (g1076) & (g1077) & (g165) & (g166)) + ((g1074) & (g1075) & (!g1076) & (!g1077) & (!g165) & (!g166)) + ((g1074) & (g1075) & (!g1076) & (!g1077) & (g165) & (!g166)) + ((g1074) & (g1075) & (!g1076) & (g1077) & (!g165) & (!g166)) + ((g1074) & (g1075) & (!g1076) & (g1077) & (g165) & (!g166)) + ((g1074) & (g1075) & (!g1076) & (g1077) & (g165) & (g166)) + ((g1074) & (g1075) & (g1076) & (!g1077) & (!g165) & (!g166)) + ((g1074) & (g1075) & (g1076) & (!g1077) & (!g165) & (g166)) + ((g1074) & (g1075) & (g1076) & (!g1077) & (g165) & (!g166)) + ((g1074) & (g1075) & (g1076) & (g1077) & (!g165) & (!g166)) + ((g1074) & (g1075) & (g1076) & (g1077) & (!g165) & (g166)) + ((g1074) & (g1075) & (g1076) & (g1077) & (g165) & (!g166)) + ((g1074) & (g1075) & (g1076) & (g1077) & (g165) & (g166)));
	assign g4654 = (((!g2177) & (!sk[121]) & (!g3444) & (g1079)) + ((!g2177) & (!sk[121]) & (g3444) & (!g1079)) + ((!g2177) & (!sk[121]) & (g3444) & (g1079)) + ((!g2177) & (sk[121]) & (!g3444) & (g1079)) + ((!g2177) & (sk[121]) & (g3444) & (g1079)) + ((g2177) & (!sk[121]) & (!g3444) & (g1079)) + ((g2177) & (!sk[121]) & (g3444) & (!g1079)) + ((g2177) & (!sk[121]) & (g3444) & (g1079)) + ((g2177) & (sk[121]) & (g3444) & (!g1079)) + ((g2177) & (sk[121]) & (g3444) & (g1079)));
	assign g4655 = (((!g2178) & (!sk[122]) & (!g3444) & (g1080)) + ((!g2178) & (!sk[122]) & (g3444) & (!g1080)) + ((!g2178) & (!sk[122]) & (g3444) & (g1080)) + ((!g2178) & (sk[122]) & (!g3444) & (g1080)) + ((!g2178) & (sk[122]) & (g3444) & (g1080)) + ((g2178) & (!sk[122]) & (!g3444) & (g1080)) + ((g2178) & (!sk[122]) & (g3444) & (!g1080)) + ((g2178) & (!sk[122]) & (g3444) & (g1080)) + ((g2178) & (sk[122]) & (g3444) & (!g1080)) + ((g2178) & (sk[122]) & (g3444) & (g1080)));
	assign g4656 = (((!g2179) & (!g3444) & (!sk[123]) & (g1081)) + ((!g2179) & (!g3444) & (sk[123]) & (g1081)) + ((!g2179) & (g3444) & (!sk[123]) & (!g1081)) + ((!g2179) & (g3444) & (!sk[123]) & (g1081)) + ((!g2179) & (g3444) & (sk[123]) & (g1081)) + ((g2179) & (!g3444) & (!sk[123]) & (g1081)) + ((g2179) & (g3444) & (!sk[123]) & (!g1081)) + ((g2179) & (g3444) & (!sk[123]) & (g1081)) + ((g2179) & (g3444) & (sk[123]) & (!g1081)) + ((g2179) & (g3444) & (sk[123]) & (g1081)));
	assign g1082 = (((!sk[124]) & (!g165) & (!g166) & (!g1079) & (g1080) & (!g1081)) + ((!sk[124]) & (!g165) & (!g166) & (!g1079) & (g1080) & (g1081)) + ((!sk[124]) & (!g165) & (!g166) & (g1079) & (!g1080) & (!g1081)) + ((!sk[124]) & (!g165) & (!g166) & (g1079) & (!g1080) & (g1081)) + ((!sk[124]) & (!g165) & (!g166) & (g1079) & (g1080) & (!g1081)) + ((!sk[124]) & (!g165) & (!g166) & (g1079) & (g1080) & (g1081)) + ((!sk[124]) & (!g165) & (g166) & (!g1079) & (!g1080) & (!g1081)) + ((!sk[124]) & (!g165) & (g166) & (!g1079) & (!g1080) & (g1081)) + ((!sk[124]) & (!g165) & (g166) & (!g1079) & (g1080) & (!g1081)) + ((!sk[124]) & (!g165) & (g166) & (!g1079) & (g1080) & (g1081)) + ((!sk[124]) & (!g165) & (g166) & (g1079) & (!g1080) & (!g1081)) + ((!sk[124]) & (!g165) & (g166) & (g1079) & (!g1080) & (g1081)) + ((!sk[124]) & (!g165) & (g166) & (g1079) & (g1080) & (!g1081)) + ((!sk[124]) & (!g165) & (g166) & (g1079) & (g1080) & (g1081)) + ((!sk[124]) & (g165) & (!g166) & (!g1079) & (g1080) & (!g1081)) + ((!sk[124]) & (g165) & (!g166) & (!g1079) & (g1080) & (g1081)) + ((!sk[124]) & (g165) & (!g166) & (g1079) & (!g1080) & (!g1081)) + ((!sk[124]) & (g165) & (!g166) & (g1079) & (!g1080) & (g1081)) + ((!sk[124]) & (g165) & (!g166) & (g1079) & (g1080) & (!g1081)) + ((!sk[124]) & (g165) & (!g166) & (g1079) & (g1080) & (g1081)) + ((!sk[124]) & (g165) & (g166) & (!g1079) & (!g1080) & (!g1081)) + ((!sk[124]) & (g165) & (g166) & (!g1079) & (!g1080) & (g1081)) + ((!sk[124]) & (g165) & (g166) & (!g1079) & (g1080) & (!g1081)) + ((!sk[124]) & (g165) & (g166) & (!g1079) & (g1080) & (g1081)) + ((!sk[124]) & (g165) & (g166) & (g1079) & (!g1080) & (!g1081)) + ((!sk[124]) & (g165) & (g166) & (g1079) & (!g1080) & (g1081)) + ((!sk[124]) & (g165) & (g166) & (g1079) & (g1080) & (!g1081)) + ((!sk[124]) & (g165) & (g166) & (g1079) & (g1080) & (g1081)) + ((sk[124]) & (!g165) & (g166) & (!g1079) & (!g1080) & (g1081)) + ((sk[124]) & (!g165) & (g166) & (!g1079) & (g1080) & (g1081)) + ((sk[124]) & (!g165) & (g166) & (g1079) & (!g1080) & (g1081)) + ((sk[124]) & (!g165) & (g166) & (g1079) & (g1080) & (g1081)) + ((sk[124]) & (g165) & (!g166) & (g1079) & (!g1080) & (!g1081)) + ((sk[124]) & (g165) & (!g166) & (g1079) & (!g1080) & (g1081)) + ((sk[124]) & (g165) & (!g166) & (g1079) & (g1080) & (!g1081)) + ((sk[124]) & (g165) & (!g166) & (g1079) & (g1080) & (g1081)) + ((sk[124]) & (g165) & (g166) & (!g1079) & (g1080) & (!g1081)) + ((sk[124]) & (g165) & (g166) & (!g1079) & (g1080) & (g1081)) + ((sk[124]) & (g165) & (g166) & (g1079) & (g1080) & (!g1081)) + ((sk[124]) & (g165) & (g166) & (g1079) & (g1080) & (g1081)));
	assign g4657 = (((!g2162) & (!sk[125]) & (!g3444) & (g1083)) + ((!g2162) & (!sk[125]) & (g3444) & (!g1083)) + ((!g2162) & (!sk[125]) & (g3444) & (g1083)) + ((!g2162) & (sk[125]) & (!g3444) & (g1083)) + ((!g2162) & (sk[125]) & (g3444) & (g1083)) + ((g2162) & (!sk[125]) & (!g3444) & (g1083)) + ((g2162) & (!sk[125]) & (g3444) & (!g1083)) + ((g2162) & (!sk[125]) & (g3444) & (g1083)) + ((g2162) & (sk[125]) & (g3444) & (!g1083)) + ((g2162) & (sk[125]) & (g3444) & (g1083)));
	assign g4658 = (((!g2164) & (!sk[126]) & (!g3444) & (g1084)) + ((!g2164) & (!sk[126]) & (g3444) & (!g1084)) + ((!g2164) & (!sk[126]) & (g3444) & (g1084)) + ((!g2164) & (sk[126]) & (!g3444) & (g1084)) + ((!g2164) & (sk[126]) & (g3444) & (g1084)) + ((g2164) & (!sk[126]) & (!g3444) & (g1084)) + ((g2164) & (!sk[126]) & (g3444) & (!g1084)) + ((g2164) & (!sk[126]) & (g3444) & (g1084)) + ((g2164) & (sk[126]) & (g3444) & (!g1084)) + ((g2164) & (sk[126]) & (g3444) & (g1084)));
	assign g4659 = (((!sk[127]) & (!g2166) & (!g3444) & (g1085)) + ((!sk[127]) & (!g2166) & (g3444) & (!g1085)) + ((!sk[127]) & (!g2166) & (g3444) & (g1085)) + ((!sk[127]) & (g2166) & (!g3444) & (g1085)) + ((!sk[127]) & (g2166) & (g3444) & (!g1085)) + ((!sk[127]) & (g2166) & (g3444) & (g1085)) + ((sk[127]) & (!g2166) & (!g3444) & (g1085)) + ((sk[127]) & (!g2166) & (g3444) & (g1085)) + ((sk[127]) & (g2166) & (g3444) & (!g1085)) + ((sk[127]) & (g2166) & (g3444) & (g1085)));
	assign g4660 = (((!g2168) & (!sk[0]) & (!g3444) & (g1086)) + ((!g2168) & (!sk[0]) & (g3444) & (!g1086)) + ((!g2168) & (!sk[0]) & (g3444) & (g1086)) + ((!g2168) & (sk[0]) & (!g3444) & (g1086)) + ((!g2168) & (sk[0]) & (g3444) & (g1086)) + ((g2168) & (!sk[0]) & (!g3444) & (g1086)) + ((g2168) & (!sk[0]) & (g3444) & (!g1086)) + ((g2168) & (!sk[0]) & (g3444) & (g1086)) + ((g2168) & (sk[0]) & (g3444) & (!g1086)) + ((g2168) & (sk[0]) & (g3444) & (g1086)));
	assign g1087 = (((!g1083) & (!g1084) & (!g1085) & (g1086) & (g165) & (g166)) + ((!g1083) & (!g1084) & (g1085) & (!g1086) & (!g165) & (g166)) + ((!g1083) & (!g1084) & (g1085) & (g1086) & (!g165) & (g166)) + ((!g1083) & (!g1084) & (g1085) & (g1086) & (g165) & (g166)) + ((!g1083) & (g1084) & (!g1085) & (!g1086) & (g165) & (!g166)) + ((!g1083) & (g1084) & (!g1085) & (g1086) & (g165) & (!g166)) + ((!g1083) & (g1084) & (!g1085) & (g1086) & (g165) & (g166)) + ((!g1083) & (g1084) & (g1085) & (!g1086) & (!g165) & (g166)) + ((!g1083) & (g1084) & (g1085) & (!g1086) & (g165) & (!g166)) + ((!g1083) & (g1084) & (g1085) & (g1086) & (!g165) & (g166)) + ((!g1083) & (g1084) & (g1085) & (g1086) & (g165) & (!g166)) + ((!g1083) & (g1084) & (g1085) & (g1086) & (g165) & (g166)) + ((g1083) & (!g1084) & (!g1085) & (!g1086) & (!g165) & (!g166)) + ((g1083) & (!g1084) & (!g1085) & (g1086) & (!g165) & (!g166)) + ((g1083) & (!g1084) & (!g1085) & (g1086) & (g165) & (g166)) + ((g1083) & (!g1084) & (g1085) & (!g1086) & (!g165) & (!g166)) + ((g1083) & (!g1084) & (g1085) & (!g1086) & (!g165) & (g166)) + ((g1083) & (!g1084) & (g1085) & (g1086) & (!g165) & (!g166)) + ((g1083) & (!g1084) & (g1085) & (g1086) & (!g165) & (g166)) + ((g1083) & (!g1084) & (g1085) & (g1086) & (g165) & (g166)) + ((g1083) & (g1084) & (!g1085) & (!g1086) & (!g165) & (!g166)) + ((g1083) & (g1084) & (!g1085) & (!g1086) & (g165) & (!g166)) + ((g1083) & (g1084) & (!g1085) & (g1086) & (!g165) & (!g166)) + ((g1083) & (g1084) & (!g1085) & (g1086) & (g165) & (!g166)) + ((g1083) & (g1084) & (!g1085) & (g1086) & (g165) & (g166)) + ((g1083) & (g1084) & (g1085) & (!g1086) & (!g165) & (!g166)) + ((g1083) & (g1084) & (g1085) & (!g1086) & (!g165) & (g166)) + ((g1083) & (g1084) & (g1085) & (!g1086) & (g165) & (!g166)) + ((g1083) & (g1084) & (g1085) & (g1086) & (!g165) & (!g166)) + ((g1083) & (g1084) & (g1085) & (g1086) & (!g165) & (g166)) + ((g1083) & (g1084) & (g1085) & (g1086) & (g165) & (!g166)) + ((g1083) & (g1084) & (g1085) & (g1086) & (g165) & (g166)));
	assign g4661 = (((!sk[2]) & (!g2169) & (!g3444) & (g1088)) + ((!sk[2]) & (!g2169) & (g3444) & (!g1088)) + ((!sk[2]) & (!g2169) & (g3444) & (g1088)) + ((!sk[2]) & (g2169) & (!g3444) & (g1088)) + ((!sk[2]) & (g2169) & (g3444) & (!g1088)) + ((!sk[2]) & (g2169) & (g3444) & (g1088)) + ((sk[2]) & (!g2169) & (!g3444) & (g1088)) + ((sk[2]) & (!g2169) & (g3444) & (g1088)) + ((sk[2]) & (g2169) & (g3444) & (!g1088)) + ((sk[2]) & (g2169) & (g3444) & (g1088)));
	assign g4662 = (((!g2170) & (!sk[3]) & (!g3444) & (g1089)) + ((!g2170) & (!sk[3]) & (g3444) & (!g1089)) + ((!g2170) & (!sk[3]) & (g3444) & (g1089)) + ((!g2170) & (sk[3]) & (!g3444) & (g1089)) + ((!g2170) & (sk[3]) & (g3444) & (g1089)) + ((g2170) & (!sk[3]) & (!g3444) & (g1089)) + ((g2170) & (!sk[3]) & (g3444) & (!g1089)) + ((g2170) & (!sk[3]) & (g3444) & (g1089)) + ((g2170) & (sk[3]) & (g3444) & (!g1089)) + ((g2170) & (sk[3]) & (g3444) & (g1089)));
	assign g4663 = (((!g2171) & (!sk[4]) & (!g3444) & (g1090)) + ((!g2171) & (!sk[4]) & (g3444) & (!g1090)) + ((!g2171) & (!sk[4]) & (g3444) & (g1090)) + ((!g2171) & (sk[4]) & (!g3444) & (g1090)) + ((!g2171) & (sk[4]) & (g3444) & (g1090)) + ((g2171) & (!sk[4]) & (!g3444) & (g1090)) + ((g2171) & (!sk[4]) & (g3444) & (!g1090)) + ((g2171) & (!sk[4]) & (g3444) & (g1090)) + ((g2171) & (sk[4]) & (g3444) & (!g1090)) + ((g2171) & (sk[4]) & (g3444) & (g1090)));
	assign g4664 = (((!g2172) & (!sk[5]) & (!g3444) & (g1091)) + ((!g2172) & (!sk[5]) & (g3444) & (!g1091)) + ((!g2172) & (!sk[5]) & (g3444) & (g1091)) + ((!g2172) & (sk[5]) & (!g3444) & (g1091)) + ((!g2172) & (sk[5]) & (g3444) & (g1091)) + ((g2172) & (!sk[5]) & (!g3444) & (g1091)) + ((g2172) & (!sk[5]) & (g3444) & (!g1091)) + ((g2172) & (!sk[5]) & (g3444) & (g1091)) + ((g2172) & (sk[5]) & (g3444) & (!g1091)) + ((g2172) & (sk[5]) & (g3444) & (g1091)));
	assign g1092 = (((!g1088) & (!g1089) & (!g1090) & (g1091) & (g165) & (g166)) + ((!g1088) & (!g1089) & (g1090) & (!g1091) & (!g165) & (g166)) + ((!g1088) & (!g1089) & (g1090) & (g1091) & (!g165) & (g166)) + ((!g1088) & (!g1089) & (g1090) & (g1091) & (g165) & (g166)) + ((!g1088) & (g1089) & (!g1090) & (!g1091) & (g165) & (!g166)) + ((!g1088) & (g1089) & (!g1090) & (g1091) & (g165) & (!g166)) + ((!g1088) & (g1089) & (!g1090) & (g1091) & (g165) & (g166)) + ((!g1088) & (g1089) & (g1090) & (!g1091) & (!g165) & (g166)) + ((!g1088) & (g1089) & (g1090) & (!g1091) & (g165) & (!g166)) + ((!g1088) & (g1089) & (g1090) & (g1091) & (!g165) & (g166)) + ((!g1088) & (g1089) & (g1090) & (g1091) & (g165) & (!g166)) + ((!g1088) & (g1089) & (g1090) & (g1091) & (g165) & (g166)) + ((g1088) & (!g1089) & (!g1090) & (!g1091) & (!g165) & (!g166)) + ((g1088) & (!g1089) & (!g1090) & (g1091) & (!g165) & (!g166)) + ((g1088) & (!g1089) & (!g1090) & (g1091) & (g165) & (g166)) + ((g1088) & (!g1089) & (g1090) & (!g1091) & (!g165) & (!g166)) + ((g1088) & (!g1089) & (g1090) & (!g1091) & (!g165) & (g166)) + ((g1088) & (!g1089) & (g1090) & (g1091) & (!g165) & (!g166)) + ((g1088) & (!g1089) & (g1090) & (g1091) & (!g165) & (g166)) + ((g1088) & (!g1089) & (g1090) & (g1091) & (g165) & (g166)) + ((g1088) & (g1089) & (!g1090) & (!g1091) & (!g165) & (!g166)) + ((g1088) & (g1089) & (!g1090) & (!g1091) & (g165) & (!g166)) + ((g1088) & (g1089) & (!g1090) & (g1091) & (!g165) & (!g166)) + ((g1088) & (g1089) & (!g1090) & (g1091) & (g165) & (!g166)) + ((g1088) & (g1089) & (!g1090) & (g1091) & (g165) & (g166)) + ((g1088) & (g1089) & (g1090) & (!g1091) & (!g165) & (!g166)) + ((g1088) & (g1089) & (g1090) & (!g1091) & (!g165) & (g166)) + ((g1088) & (g1089) & (g1090) & (!g1091) & (g165) & (!g166)) + ((g1088) & (g1089) & (g1090) & (g1091) & (!g165) & (!g166)) + ((g1088) & (g1089) & (g1090) & (g1091) & (!g165) & (g166)) + ((g1088) & (g1089) & (g1090) & (g1091) & (g165) & (!g166)) + ((g1088) & (g1089) & (g1090) & (g1091) & (g165) & (g166)));
	assign g1093 = (((!g147) & (!g148) & (!g1078) & (g1082) & (!g1087) & (!g1092)) + ((!g147) & (!g148) & (!g1078) & (g1082) & (!g1087) & (g1092)) + ((!g147) & (!g148) & (!g1078) & (g1082) & (g1087) & (!g1092)) + ((!g147) & (!g148) & (!g1078) & (g1082) & (g1087) & (g1092)) + ((!g147) & (!g148) & (g1078) & (g1082) & (!g1087) & (!g1092)) + ((!g147) & (!g148) & (g1078) & (g1082) & (!g1087) & (g1092)) + ((!g147) & (!g148) & (g1078) & (g1082) & (g1087) & (!g1092)) + ((!g147) & (!g148) & (g1078) & (g1082) & (g1087) & (g1092)) + ((!g147) & (g148) & (!g1078) & (!g1082) & (!g1087) & (g1092)) + ((!g147) & (g148) & (!g1078) & (!g1082) & (g1087) & (g1092)) + ((!g147) & (g148) & (!g1078) & (g1082) & (!g1087) & (g1092)) + ((!g147) & (g148) & (!g1078) & (g1082) & (g1087) & (g1092)) + ((!g147) & (g148) & (g1078) & (!g1082) & (!g1087) & (g1092)) + ((!g147) & (g148) & (g1078) & (!g1082) & (g1087) & (g1092)) + ((!g147) & (g148) & (g1078) & (g1082) & (!g1087) & (g1092)) + ((!g147) & (g148) & (g1078) & (g1082) & (g1087) & (g1092)) + ((g147) & (!g148) & (g1078) & (!g1082) & (!g1087) & (!g1092)) + ((g147) & (!g148) & (g1078) & (!g1082) & (!g1087) & (g1092)) + ((g147) & (!g148) & (g1078) & (!g1082) & (g1087) & (!g1092)) + ((g147) & (!g148) & (g1078) & (!g1082) & (g1087) & (g1092)) + ((g147) & (!g148) & (g1078) & (g1082) & (!g1087) & (!g1092)) + ((g147) & (!g148) & (g1078) & (g1082) & (!g1087) & (g1092)) + ((g147) & (!g148) & (g1078) & (g1082) & (g1087) & (!g1092)) + ((g147) & (!g148) & (g1078) & (g1082) & (g1087) & (g1092)) + ((g147) & (g148) & (!g1078) & (!g1082) & (g1087) & (!g1092)) + ((g147) & (g148) & (!g1078) & (!g1082) & (g1087) & (g1092)) + ((g147) & (g148) & (!g1078) & (g1082) & (g1087) & (!g1092)) + ((g147) & (g148) & (!g1078) & (g1082) & (g1087) & (g1092)) + ((g147) & (g148) & (g1078) & (!g1082) & (g1087) & (!g1092)) + ((g147) & (g148) & (g1078) & (!g1082) & (g1087) & (g1092)) + ((g147) & (g148) & (g1078) & (g1082) & (g1087) & (!g1092)) + ((g147) & (g148) & (g1078) & (g1082) & (g1087) & (g1092)));
	assign g1094 = (((!sk[8]) & (!g142) & (!g1073) & (g1093)) + ((!sk[8]) & (!g142) & (g1073) & (!g1093)) + ((!sk[8]) & (!g142) & (g1073) & (g1093)) + ((!sk[8]) & (g142) & (!g1073) & (g1093)) + ((!sk[8]) & (g142) & (g1073) & (!g1093)) + ((!sk[8]) & (g142) & (g1073) & (g1093)) + ((sk[8]) & (!g142) & (!g1073) & (g1093)) + ((sk[8]) & (!g142) & (g1073) & (g1093)) + ((sk[8]) & (g142) & (g1073) & (!g1093)) + ((sk[8]) & (g142) & (g1073) & (g1093)));
	assign g4665 = (((!g2059) & (!g2641) & (!sk[9]) & (g1095)) + ((!g2059) & (!g2641) & (sk[9]) & (g1095)) + ((!g2059) & (g2641) & (!sk[9]) & (!g1095)) + ((!g2059) & (g2641) & (!sk[9]) & (g1095)) + ((!g2059) & (g2641) & (sk[9]) & (g1095)) + ((g2059) & (!g2641) & (!sk[9]) & (g1095)) + ((g2059) & (g2641) & (!sk[9]) & (!g1095)) + ((g2059) & (g2641) & (!sk[9]) & (g1095)) + ((g2059) & (g2641) & (sk[9]) & (!g1095)) + ((g2059) & (g2641) & (sk[9]) & (g1095)));
	assign g1096 = (((!g1049) & (!sk[10]) & (!g1051) & (g916)) + ((!g1049) & (!sk[10]) & (g1051) & (!g916)) + ((!g1049) & (!sk[10]) & (g1051) & (g916)) + ((!g1049) & (sk[10]) & (g1051) & (!g916)) + ((g1049) & (!sk[10]) & (!g1051) & (g916)) + ((g1049) & (!sk[10]) & (g1051) & (!g916)) + ((g1049) & (!sk[10]) & (g1051) & (g916)) + ((g1049) & (sk[10]) & (!g1051) & (!g916)) + ((g1049) & (sk[10]) & (g1051) & (!g916)) + ((g1049) & (sk[10]) & (g1051) & (g916)));
	assign g1097 = (((!g126) & (!sk[11]) & (!g1094) & (!g1095) & (g1096) & (!g916)) + ((!g126) & (!sk[11]) & (!g1094) & (!g1095) & (g1096) & (g916)) + ((!g126) & (!sk[11]) & (!g1094) & (g1095) & (!g1096) & (!g916)) + ((!g126) & (!sk[11]) & (!g1094) & (g1095) & (!g1096) & (g916)) + ((!g126) & (!sk[11]) & (!g1094) & (g1095) & (g1096) & (!g916)) + ((!g126) & (!sk[11]) & (!g1094) & (g1095) & (g1096) & (g916)) + ((!g126) & (!sk[11]) & (g1094) & (!g1095) & (!g1096) & (!g916)) + ((!g126) & (!sk[11]) & (g1094) & (!g1095) & (!g1096) & (g916)) + ((!g126) & (!sk[11]) & (g1094) & (!g1095) & (g1096) & (!g916)) + ((!g126) & (!sk[11]) & (g1094) & (!g1095) & (g1096) & (g916)) + ((!g126) & (!sk[11]) & (g1094) & (g1095) & (!g1096) & (!g916)) + ((!g126) & (!sk[11]) & (g1094) & (g1095) & (!g1096) & (g916)) + ((!g126) & (!sk[11]) & (g1094) & (g1095) & (g1096) & (!g916)) + ((!g126) & (!sk[11]) & (g1094) & (g1095) & (g1096) & (g916)) + ((!g126) & (sk[11]) & (!g1094) & (g1095) & (!g1096) & (!g916)) + ((!g126) & (sk[11]) & (!g1094) & (g1095) & (!g1096) & (g916)) + ((!g126) & (sk[11]) & (!g1094) & (g1095) & (g1096) & (!g916)) + ((!g126) & (sk[11]) & (!g1094) & (g1095) & (g1096) & (g916)) + ((!g126) & (sk[11]) & (g1094) & (g1095) & (!g1096) & (!g916)) + ((!g126) & (sk[11]) & (g1094) & (g1095) & (!g1096) & (g916)) + ((!g126) & (sk[11]) & (g1094) & (g1095) & (g1096) & (!g916)) + ((!g126) & (sk[11]) & (g1094) & (g1095) & (g1096) & (g916)) + ((g126) & (!sk[11]) & (!g1094) & (!g1095) & (g1096) & (!g916)) + ((g126) & (!sk[11]) & (!g1094) & (!g1095) & (g1096) & (g916)) + ((g126) & (!sk[11]) & (!g1094) & (g1095) & (!g1096) & (!g916)) + ((g126) & (!sk[11]) & (!g1094) & (g1095) & (!g1096) & (g916)) + ((g126) & (!sk[11]) & (!g1094) & (g1095) & (g1096) & (!g916)) + ((g126) & (!sk[11]) & (!g1094) & (g1095) & (g1096) & (g916)) + ((g126) & (!sk[11]) & (g1094) & (!g1095) & (!g1096) & (!g916)) + ((g126) & (!sk[11]) & (g1094) & (!g1095) & (!g1096) & (g916)) + ((g126) & (!sk[11]) & (g1094) & (!g1095) & (g1096) & (!g916)) + ((g126) & (!sk[11]) & (g1094) & (!g1095) & (g1096) & (g916)) + ((g126) & (!sk[11]) & (g1094) & (g1095) & (!g1096) & (!g916)) + ((g126) & (!sk[11]) & (g1094) & (g1095) & (!g1096) & (g916)) + ((g126) & (!sk[11]) & (g1094) & (g1095) & (g1096) & (!g916)) + ((g126) & (!sk[11]) & (g1094) & (g1095) & (g1096) & (g916)) + ((g126) & (sk[11]) & (!g1094) & (!g1095) & (!g1096) & (!g916)) + ((g126) & (sk[11]) & (!g1094) & (!g1095) & (g1096) & (g916)) + ((g126) & (sk[11]) & (!g1094) & (g1095) & (!g1096) & (!g916)) + ((g126) & (sk[11]) & (!g1094) & (g1095) & (g1096) & (g916)) + ((g126) & (sk[11]) & (g1094) & (!g1095) & (!g1096) & (g916)) + ((g126) & (sk[11]) & (g1094) & (!g1095) & (g1096) & (!g916)) + ((g126) & (sk[11]) & (g1094) & (g1095) & (!g1096) & (g916)) + ((g126) & (sk[11]) & (g1094) & (g1095) & (g1096) & (!g916)));
	assign g4666 = (((!sk[12]) & (!g2140) & (!g3420) & (g1098)) + ((!sk[12]) & (!g2140) & (g3420) & (!g1098)) + ((!sk[12]) & (!g2140) & (g3420) & (g1098)) + ((!sk[12]) & (g2140) & (!g3420) & (g1098)) + ((!sk[12]) & (g2140) & (g3420) & (!g1098)) + ((!sk[12]) & (g2140) & (g3420) & (g1098)) + ((sk[12]) & (!g2140) & (!g3420) & (g1098)) + ((sk[12]) & (!g2140) & (g3420) & (g1098)) + ((sk[12]) & (g2140) & (g3420) & (!g1098)) + ((sk[12]) & (g2140) & (g3420) & (g1098)));
	assign g4667 = (((!sk[13]) & (!g2142) & (!g3420) & (g1099)) + ((!sk[13]) & (!g2142) & (g3420) & (!g1099)) + ((!sk[13]) & (!g2142) & (g3420) & (g1099)) + ((!sk[13]) & (g2142) & (!g3420) & (g1099)) + ((!sk[13]) & (g2142) & (g3420) & (!g1099)) + ((!sk[13]) & (g2142) & (g3420) & (g1099)) + ((sk[13]) & (!g2142) & (!g3420) & (g1099)) + ((sk[13]) & (!g2142) & (g3420) & (g1099)) + ((sk[13]) & (g2142) & (g3420) & (!g1099)) + ((sk[13]) & (g2142) & (g3420) & (g1099)));
	assign g4668 = (((!g2144) & (!sk[14]) & (!g3420) & (g1100)) + ((!g2144) & (!sk[14]) & (g3420) & (!g1100)) + ((!g2144) & (!sk[14]) & (g3420) & (g1100)) + ((!g2144) & (sk[14]) & (!g3420) & (g1100)) + ((!g2144) & (sk[14]) & (g3420) & (g1100)) + ((g2144) & (!sk[14]) & (!g3420) & (g1100)) + ((g2144) & (!sk[14]) & (g3420) & (!g1100)) + ((g2144) & (!sk[14]) & (g3420) & (g1100)) + ((g2144) & (sk[14]) & (g3420) & (!g1100)) + ((g2144) & (sk[14]) & (g3420) & (g1100)));
	assign g4669 = (((!g2145) & (!g3420) & (!sk[15]) & (g1101)) + ((!g2145) & (!g3420) & (sk[15]) & (g1101)) + ((!g2145) & (g3420) & (!sk[15]) & (!g1101)) + ((!g2145) & (g3420) & (!sk[15]) & (g1101)) + ((!g2145) & (g3420) & (sk[15]) & (g1101)) + ((g2145) & (!g3420) & (!sk[15]) & (g1101)) + ((g2145) & (g3420) & (!sk[15]) & (!g1101)) + ((g2145) & (g3420) & (!sk[15]) & (g1101)) + ((g2145) & (g3420) & (sk[15]) & (!g1101)) + ((g2145) & (g3420) & (sk[15]) & (g1101)));
	assign g1102 = (((!g1098) & (!g1099) & (!g1100) & (g1101) & (g147) & (g148)) + ((!g1098) & (!g1099) & (g1100) & (!g1101) & (!g147) & (g148)) + ((!g1098) & (!g1099) & (g1100) & (g1101) & (!g147) & (g148)) + ((!g1098) & (!g1099) & (g1100) & (g1101) & (g147) & (g148)) + ((!g1098) & (g1099) & (!g1100) & (!g1101) & (g147) & (!g148)) + ((!g1098) & (g1099) & (!g1100) & (g1101) & (g147) & (!g148)) + ((!g1098) & (g1099) & (!g1100) & (g1101) & (g147) & (g148)) + ((!g1098) & (g1099) & (g1100) & (!g1101) & (!g147) & (g148)) + ((!g1098) & (g1099) & (g1100) & (!g1101) & (g147) & (!g148)) + ((!g1098) & (g1099) & (g1100) & (g1101) & (!g147) & (g148)) + ((!g1098) & (g1099) & (g1100) & (g1101) & (g147) & (!g148)) + ((!g1098) & (g1099) & (g1100) & (g1101) & (g147) & (g148)) + ((g1098) & (!g1099) & (!g1100) & (!g1101) & (!g147) & (!g148)) + ((g1098) & (!g1099) & (!g1100) & (g1101) & (!g147) & (!g148)) + ((g1098) & (!g1099) & (!g1100) & (g1101) & (g147) & (g148)) + ((g1098) & (!g1099) & (g1100) & (!g1101) & (!g147) & (!g148)) + ((g1098) & (!g1099) & (g1100) & (!g1101) & (!g147) & (g148)) + ((g1098) & (!g1099) & (g1100) & (g1101) & (!g147) & (!g148)) + ((g1098) & (!g1099) & (g1100) & (g1101) & (!g147) & (g148)) + ((g1098) & (!g1099) & (g1100) & (g1101) & (g147) & (g148)) + ((g1098) & (g1099) & (!g1100) & (!g1101) & (!g147) & (!g148)) + ((g1098) & (g1099) & (!g1100) & (!g1101) & (g147) & (!g148)) + ((g1098) & (g1099) & (!g1100) & (g1101) & (!g147) & (!g148)) + ((g1098) & (g1099) & (!g1100) & (g1101) & (g147) & (!g148)) + ((g1098) & (g1099) & (!g1100) & (g1101) & (g147) & (g148)) + ((g1098) & (g1099) & (g1100) & (!g1101) & (!g147) & (!g148)) + ((g1098) & (g1099) & (g1100) & (!g1101) & (!g147) & (g148)) + ((g1098) & (g1099) & (g1100) & (!g1101) & (g147) & (!g148)) + ((g1098) & (g1099) & (g1100) & (g1101) & (!g147) & (!g148)) + ((g1098) & (g1099) & (g1100) & (g1101) & (!g147) & (g148)) + ((g1098) & (g1099) & (g1100) & (g1101) & (g147) & (!g148)) + ((g1098) & (g1099) & (g1100) & (g1101) & (g147) & (g148)));
	assign g4670 = (((!g2146) & (!sk[17]) & (!g3420) & (g1103)) + ((!g2146) & (!sk[17]) & (g3420) & (!g1103)) + ((!g2146) & (!sk[17]) & (g3420) & (g1103)) + ((!g2146) & (sk[17]) & (!g3420) & (g1103)) + ((!g2146) & (sk[17]) & (g3420) & (g1103)) + ((g2146) & (!sk[17]) & (!g3420) & (g1103)) + ((g2146) & (!sk[17]) & (g3420) & (!g1103)) + ((g2146) & (!sk[17]) & (g3420) & (g1103)) + ((g2146) & (sk[17]) & (g3420) & (!g1103)) + ((g2146) & (sk[17]) & (g3420) & (g1103)));
	assign g4671 = (((!g2148) & (!g3420) & (!sk[18]) & (g1104)) + ((!g2148) & (!g3420) & (sk[18]) & (g1104)) + ((!g2148) & (g3420) & (!sk[18]) & (!g1104)) + ((!g2148) & (g3420) & (!sk[18]) & (g1104)) + ((!g2148) & (g3420) & (sk[18]) & (g1104)) + ((g2148) & (!g3420) & (!sk[18]) & (g1104)) + ((g2148) & (g3420) & (!sk[18]) & (!g1104)) + ((g2148) & (g3420) & (!sk[18]) & (g1104)) + ((g2148) & (g3420) & (sk[18]) & (!g1104)) + ((g2148) & (g3420) & (sk[18]) & (g1104)));
	assign g4672 = (((!sk[19]) & (!g2150) & (!g3420) & (g1105)) + ((!sk[19]) & (!g2150) & (g3420) & (!g1105)) + ((!sk[19]) & (!g2150) & (g3420) & (g1105)) + ((!sk[19]) & (g2150) & (!g3420) & (g1105)) + ((!sk[19]) & (g2150) & (g3420) & (!g1105)) + ((!sk[19]) & (g2150) & (g3420) & (g1105)) + ((sk[19]) & (!g2150) & (!g3420) & (g1105)) + ((sk[19]) & (!g2150) & (g3420) & (g1105)) + ((sk[19]) & (g2150) & (g3420) & (!g1105)) + ((sk[19]) & (g2150) & (g3420) & (g1105)));
	assign g4673 = (((!g2151) & (!g3420) & (!sk[20]) & (g1106)) + ((!g2151) & (!g3420) & (sk[20]) & (g1106)) + ((!g2151) & (g3420) & (!sk[20]) & (!g1106)) + ((!g2151) & (g3420) & (!sk[20]) & (g1106)) + ((!g2151) & (g3420) & (sk[20]) & (g1106)) + ((g2151) & (!g3420) & (!sk[20]) & (g1106)) + ((g2151) & (g3420) & (!sk[20]) & (!g1106)) + ((g2151) & (g3420) & (!sk[20]) & (g1106)) + ((g2151) & (g3420) & (sk[20]) & (!g1106)) + ((g2151) & (g3420) & (sk[20]) & (g1106)));
	assign g1107 = (((!g1103) & (!g1104) & (!g1105) & (g1106) & (g147) & (g148)) + ((!g1103) & (!g1104) & (g1105) & (!g1106) & (!g147) & (g148)) + ((!g1103) & (!g1104) & (g1105) & (g1106) & (!g147) & (g148)) + ((!g1103) & (!g1104) & (g1105) & (g1106) & (g147) & (g148)) + ((!g1103) & (g1104) & (!g1105) & (!g1106) & (g147) & (!g148)) + ((!g1103) & (g1104) & (!g1105) & (g1106) & (g147) & (!g148)) + ((!g1103) & (g1104) & (!g1105) & (g1106) & (g147) & (g148)) + ((!g1103) & (g1104) & (g1105) & (!g1106) & (!g147) & (g148)) + ((!g1103) & (g1104) & (g1105) & (!g1106) & (g147) & (!g148)) + ((!g1103) & (g1104) & (g1105) & (g1106) & (!g147) & (g148)) + ((!g1103) & (g1104) & (g1105) & (g1106) & (g147) & (!g148)) + ((!g1103) & (g1104) & (g1105) & (g1106) & (g147) & (g148)) + ((g1103) & (!g1104) & (!g1105) & (!g1106) & (!g147) & (!g148)) + ((g1103) & (!g1104) & (!g1105) & (g1106) & (!g147) & (!g148)) + ((g1103) & (!g1104) & (!g1105) & (g1106) & (g147) & (g148)) + ((g1103) & (!g1104) & (g1105) & (!g1106) & (!g147) & (!g148)) + ((g1103) & (!g1104) & (g1105) & (!g1106) & (!g147) & (g148)) + ((g1103) & (!g1104) & (g1105) & (g1106) & (!g147) & (!g148)) + ((g1103) & (!g1104) & (g1105) & (g1106) & (!g147) & (g148)) + ((g1103) & (!g1104) & (g1105) & (g1106) & (g147) & (g148)) + ((g1103) & (g1104) & (!g1105) & (!g1106) & (!g147) & (!g148)) + ((g1103) & (g1104) & (!g1105) & (!g1106) & (g147) & (!g148)) + ((g1103) & (g1104) & (!g1105) & (g1106) & (!g147) & (!g148)) + ((g1103) & (g1104) & (!g1105) & (g1106) & (g147) & (!g148)) + ((g1103) & (g1104) & (!g1105) & (g1106) & (g147) & (g148)) + ((g1103) & (g1104) & (g1105) & (!g1106) & (!g147) & (!g148)) + ((g1103) & (g1104) & (g1105) & (!g1106) & (!g147) & (g148)) + ((g1103) & (g1104) & (g1105) & (!g1106) & (g147) & (!g148)) + ((g1103) & (g1104) & (g1105) & (g1106) & (!g147) & (!g148)) + ((g1103) & (g1104) & (g1105) & (g1106) & (!g147) & (g148)) + ((g1103) & (g1104) & (g1105) & (g1106) & (g147) & (!g148)) + ((g1103) & (g1104) & (g1105) & (g1106) & (g147) & (g148)));
	assign g4674 = (((!sk[22]) & (!g2152) & (!g3420) & (g1108)) + ((!sk[22]) & (!g2152) & (g3420) & (!g1108)) + ((!sk[22]) & (!g2152) & (g3420) & (g1108)) + ((!sk[22]) & (g2152) & (!g3420) & (g1108)) + ((!sk[22]) & (g2152) & (g3420) & (!g1108)) + ((!sk[22]) & (g2152) & (g3420) & (g1108)) + ((sk[22]) & (!g2152) & (!g3420) & (g1108)) + ((sk[22]) & (!g2152) & (g3420) & (g1108)) + ((sk[22]) & (g2152) & (g3420) & (!g1108)) + ((sk[22]) & (g2152) & (g3420) & (g1108)));
	assign g4675 = (((!g2153) & (!sk[23]) & (!g3420) & (g1109)) + ((!g2153) & (!sk[23]) & (g3420) & (!g1109)) + ((!g2153) & (!sk[23]) & (g3420) & (g1109)) + ((!g2153) & (sk[23]) & (!g3420) & (g1109)) + ((!g2153) & (sk[23]) & (g3420) & (g1109)) + ((g2153) & (!sk[23]) & (!g3420) & (g1109)) + ((g2153) & (!sk[23]) & (g3420) & (!g1109)) + ((g2153) & (!sk[23]) & (g3420) & (g1109)) + ((g2153) & (sk[23]) & (g3420) & (!g1109)) + ((g2153) & (sk[23]) & (g3420) & (g1109)));
	assign g4676 = (((!g2155) & (!g3420) & (!sk[24]) & (g1110)) + ((!g2155) & (!g3420) & (sk[24]) & (g1110)) + ((!g2155) & (g3420) & (!sk[24]) & (!g1110)) + ((!g2155) & (g3420) & (!sk[24]) & (g1110)) + ((!g2155) & (g3420) & (sk[24]) & (g1110)) + ((g2155) & (!g3420) & (!sk[24]) & (g1110)) + ((g2155) & (g3420) & (!sk[24]) & (!g1110)) + ((g2155) & (g3420) & (!sk[24]) & (g1110)) + ((g2155) & (g3420) & (sk[24]) & (!g1110)) + ((g2155) & (g3420) & (sk[24]) & (g1110)));
	assign g4677 = (((!g2157) & (!sk[25]) & (!g3420) & (g1111)) + ((!g2157) & (!sk[25]) & (g3420) & (!g1111)) + ((!g2157) & (!sk[25]) & (g3420) & (g1111)) + ((!g2157) & (sk[25]) & (!g3420) & (g1111)) + ((!g2157) & (sk[25]) & (g3420) & (g1111)) + ((g2157) & (!sk[25]) & (!g3420) & (g1111)) + ((g2157) & (!sk[25]) & (g3420) & (!g1111)) + ((g2157) & (!sk[25]) & (g3420) & (g1111)) + ((g2157) & (sk[25]) & (g3420) & (!g1111)) + ((g2157) & (sk[25]) & (g3420) & (g1111)));
	assign g1112 = (((!g1108) & (!g1109) & (!g1110) & (g1111) & (g147) & (g148)) + ((!g1108) & (!g1109) & (g1110) & (!g1111) & (!g147) & (g148)) + ((!g1108) & (!g1109) & (g1110) & (g1111) & (!g147) & (g148)) + ((!g1108) & (!g1109) & (g1110) & (g1111) & (g147) & (g148)) + ((!g1108) & (g1109) & (!g1110) & (!g1111) & (g147) & (!g148)) + ((!g1108) & (g1109) & (!g1110) & (g1111) & (g147) & (!g148)) + ((!g1108) & (g1109) & (!g1110) & (g1111) & (g147) & (g148)) + ((!g1108) & (g1109) & (g1110) & (!g1111) & (!g147) & (g148)) + ((!g1108) & (g1109) & (g1110) & (!g1111) & (g147) & (!g148)) + ((!g1108) & (g1109) & (g1110) & (g1111) & (!g147) & (g148)) + ((!g1108) & (g1109) & (g1110) & (g1111) & (g147) & (!g148)) + ((!g1108) & (g1109) & (g1110) & (g1111) & (g147) & (g148)) + ((g1108) & (!g1109) & (!g1110) & (!g1111) & (!g147) & (!g148)) + ((g1108) & (!g1109) & (!g1110) & (g1111) & (!g147) & (!g148)) + ((g1108) & (!g1109) & (!g1110) & (g1111) & (g147) & (g148)) + ((g1108) & (!g1109) & (g1110) & (!g1111) & (!g147) & (!g148)) + ((g1108) & (!g1109) & (g1110) & (!g1111) & (!g147) & (g148)) + ((g1108) & (!g1109) & (g1110) & (g1111) & (!g147) & (!g148)) + ((g1108) & (!g1109) & (g1110) & (g1111) & (!g147) & (g148)) + ((g1108) & (!g1109) & (g1110) & (g1111) & (g147) & (g148)) + ((g1108) & (g1109) & (!g1110) & (!g1111) & (!g147) & (!g148)) + ((g1108) & (g1109) & (!g1110) & (!g1111) & (g147) & (!g148)) + ((g1108) & (g1109) & (!g1110) & (g1111) & (!g147) & (!g148)) + ((g1108) & (g1109) & (!g1110) & (g1111) & (g147) & (!g148)) + ((g1108) & (g1109) & (!g1110) & (g1111) & (g147) & (g148)) + ((g1108) & (g1109) & (g1110) & (!g1111) & (!g147) & (!g148)) + ((g1108) & (g1109) & (g1110) & (!g1111) & (!g147) & (g148)) + ((g1108) & (g1109) & (g1110) & (!g1111) & (g147) & (!g148)) + ((g1108) & (g1109) & (g1110) & (g1111) & (!g147) & (!g148)) + ((g1108) & (g1109) & (g1110) & (g1111) & (!g147) & (g148)) + ((g1108) & (g1109) & (g1110) & (g1111) & (g147) & (!g148)) + ((g1108) & (g1109) & (g1110) & (g1111) & (g147) & (g148)));
	assign g4678 = (((!g2158) & (!g3420) & (!sk[27]) & (g1113)) + ((!g2158) & (!g3420) & (sk[27]) & (g1113)) + ((!g2158) & (g3420) & (!sk[27]) & (!g1113)) + ((!g2158) & (g3420) & (!sk[27]) & (g1113)) + ((!g2158) & (g3420) & (sk[27]) & (g1113)) + ((g2158) & (!g3420) & (!sk[27]) & (g1113)) + ((g2158) & (g3420) & (!sk[27]) & (!g1113)) + ((g2158) & (g3420) & (!sk[27]) & (g1113)) + ((g2158) & (g3420) & (sk[27]) & (!g1113)) + ((g2158) & (g3420) & (sk[27]) & (g1113)));
	assign g4679 = (((!sk[28]) & (!g2159) & (!g3420) & (g1114)) + ((!sk[28]) & (!g2159) & (g3420) & (!g1114)) + ((!sk[28]) & (!g2159) & (g3420) & (g1114)) + ((!sk[28]) & (g2159) & (!g3420) & (g1114)) + ((!sk[28]) & (g2159) & (g3420) & (!g1114)) + ((!sk[28]) & (g2159) & (g3420) & (g1114)) + ((sk[28]) & (!g2159) & (!g3420) & (g1114)) + ((sk[28]) & (!g2159) & (g3420) & (g1114)) + ((sk[28]) & (g2159) & (g3420) & (!g1114)) + ((sk[28]) & (g2159) & (g3420) & (g1114)));
	assign g4680 = (((!g2160) & (!sk[29]) & (!g3420) & (g1115)) + ((!g2160) & (!sk[29]) & (g3420) & (!g1115)) + ((!g2160) & (!sk[29]) & (g3420) & (g1115)) + ((!g2160) & (sk[29]) & (!g3420) & (g1115)) + ((!g2160) & (sk[29]) & (g3420) & (g1115)) + ((g2160) & (!sk[29]) & (!g3420) & (g1115)) + ((g2160) & (!sk[29]) & (g3420) & (!g1115)) + ((g2160) & (!sk[29]) & (g3420) & (g1115)) + ((g2160) & (sk[29]) & (g3420) & (!g1115)) + ((g2160) & (sk[29]) & (g3420) & (g1115)));
	assign g4681 = (((!g2161) & (!sk[30]) & (!g3420) & (g1116)) + ((!g2161) & (!sk[30]) & (g3420) & (!g1116)) + ((!g2161) & (!sk[30]) & (g3420) & (g1116)) + ((!g2161) & (sk[30]) & (!g3420) & (g1116)) + ((!g2161) & (sk[30]) & (g3420) & (g1116)) + ((g2161) & (!sk[30]) & (!g3420) & (g1116)) + ((g2161) & (!sk[30]) & (g3420) & (!g1116)) + ((g2161) & (!sk[30]) & (g3420) & (g1116)) + ((g2161) & (sk[30]) & (g3420) & (!g1116)) + ((g2161) & (sk[30]) & (g3420) & (g1116)));
	assign g1117 = (((!g1113) & (!g1114) & (!g1115) & (g1116) & (g147) & (g148)) + ((!g1113) & (!g1114) & (g1115) & (!g1116) & (!g147) & (g148)) + ((!g1113) & (!g1114) & (g1115) & (g1116) & (!g147) & (g148)) + ((!g1113) & (!g1114) & (g1115) & (g1116) & (g147) & (g148)) + ((!g1113) & (g1114) & (!g1115) & (!g1116) & (g147) & (!g148)) + ((!g1113) & (g1114) & (!g1115) & (g1116) & (g147) & (!g148)) + ((!g1113) & (g1114) & (!g1115) & (g1116) & (g147) & (g148)) + ((!g1113) & (g1114) & (g1115) & (!g1116) & (!g147) & (g148)) + ((!g1113) & (g1114) & (g1115) & (!g1116) & (g147) & (!g148)) + ((!g1113) & (g1114) & (g1115) & (g1116) & (!g147) & (g148)) + ((!g1113) & (g1114) & (g1115) & (g1116) & (g147) & (!g148)) + ((!g1113) & (g1114) & (g1115) & (g1116) & (g147) & (g148)) + ((g1113) & (!g1114) & (!g1115) & (!g1116) & (!g147) & (!g148)) + ((g1113) & (!g1114) & (!g1115) & (g1116) & (!g147) & (!g148)) + ((g1113) & (!g1114) & (!g1115) & (g1116) & (g147) & (g148)) + ((g1113) & (!g1114) & (g1115) & (!g1116) & (!g147) & (!g148)) + ((g1113) & (!g1114) & (g1115) & (!g1116) & (!g147) & (g148)) + ((g1113) & (!g1114) & (g1115) & (g1116) & (!g147) & (!g148)) + ((g1113) & (!g1114) & (g1115) & (g1116) & (!g147) & (g148)) + ((g1113) & (!g1114) & (g1115) & (g1116) & (g147) & (g148)) + ((g1113) & (g1114) & (!g1115) & (!g1116) & (!g147) & (!g148)) + ((g1113) & (g1114) & (!g1115) & (!g1116) & (g147) & (!g148)) + ((g1113) & (g1114) & (!g1115) & (g1116) & (!g147) & (!g148)) + ((g1113) & (g1114) & (!g1115) & (g1116) & (g147) & (!g148)) + ((g1113) & (g1114) & (!g1115) & (g1116) & (g147) & (g148)) + ((g1113) & (g1114) & (g1115) & (!g1116) & (!g147) & (!g148)) + ((g1113) & (g1114) & (g1115) & (!g1116) & (!g147) & (g148)) + ((g1113) & (g1114) & (g1115) & (!g1116) & (g147) & (!g148)) + ((g1113) & (g1114) & (g1115) & (g1116) & (!g147) & (!g148)) + ((g1113) & (g1114) & (g1115) & (g1116) & (!g147) & (g148)) + ((g1113) & (g1114) & (g1115) & (g1116) & (g147) & (!g148)) + ((g1113) & (g1114) & (g1115) & (g1116) & (g147) & (g148)));
	assign g1118 = (((!g1102) & (!g1107) & (!g1112) & (g1117) & (g165) & (g166)) + ((!g1102) & (!g1107) & (g1112) & (!g1117) & (!g165) & (g166)) + ((!g1102) & (!g1107) & (g1112) & (g1117) & (!g165) & (g166)) + ((!g1102) & (!g1107) & (g1112) & (g1117) & (g165) & (g166)) + ((!g1102) & (g1107) & (!g1112) & (!g1117) & (g165) & (!g166)) + ((!g1102) & (g1107) & (!g1112) & (g1117) & (g165) & (!g166)) + ((!g1102) & (g1107) & (!g1112) & (g1117) & (g165) & (g166)) + ((!g1102) & (g1107) & (g1112) & (!g1117) & (!g165) & (g166)) + ((!g1102) & (g1107) & (g1112) & (!g1117) & (g165) & (!g166)) + ((!g1102) & (g1107) & (g1112) & (g1117) & (!g165) & (g166)) + ((!g1102) & (g1107) & (g1112) & (g1117) & (g165) & (!g166)) + ((!g1102) & (g1107) & (g1112) & (g1117) & (g165) & (g166)) + ((g1102) & (!g1107) & (!g1112) & (!g1117) & (!g165) & (!g166)) + ((g1102) & (!g1107) & (!g1112) & (g1117) & (!g165) & (!g166)) + ((g1102) & (!g1107) & (!g1112) & (g1117) & (g165) & (g166)) + ((g1102) & (!g1107) & (g1112) & (!g1117) & (!g165) & (!g166)) + ((g1102) & (!g1107) & (g1112) & (!g1117) & (!g165) & (g166)) + ((g1102) & (!g1107) & (g1112) & (g1117) & (!g165) & (!g166)) + ((g1102) & (!g1107) & (g1112) & (g1117) & (!g165) & (g166)) + ((g1102) & (!g1107) & (g1112) & (g1117) & (g165) & (g166)) + ((g1102) & (g1107) & (!g1112) & (!g1117) & (!g165) & (!g166)) + ((g1102) & (g1107) & (!g1112) & (!g1117) & (g165) & (!g166)) + ((g1102) & (g1107) & (!g1112) & (g1117) & (!g165) & (!g166)) + ((g1102) & (g1107) & (!g1112) & (g1117) & (g165) & (!g166)) + ((g1102) & (g1107) & (!g1112) & (g1117) & (g165) & (g166)) + ((g1102) & (g1107) & (g1112) & (!g1117) & (!g165) & (!g166)) + ((g1102) & (g1107) & (g1112) & (!g1117) & (!g165) & (g166)) + ((g1102) & (g1107) & (g1112) & (!g1117) & (g165) & (!g166)) + ((g1102) & (g1107) & (g1112) & (g1117) & (!g165) & (!g166)) + ((g1102) & (g1107) & (g1112) & (g1117) & (!g165) & (g166)) + ((g1102) & (g1107) & (g1112) & (g1117) & (g165) & (!g166)) + ((g1102) & (g1107) & (g1112) & (g1117) & (g165) & (g166)));
	assign g4682 = (((!sk[33]) & (!g2173) & (!g3420) & (g1119)) + ((!sk[33]) & (!g2173) & (g3420) & (!g1119)) + ((!sk[33]) & (!g2173) & (g3420) & (g1119)) + ((!sk[33]) & (g2173) & (!g3420) & (g1119)) + ((!sk[33]) & (g2173) & (g3420) & (!g1119)) + ((!sk[33]) & (g2173) & (g3420) & (g1119)) + ((sk[33]) & (!g2173) & (!g3420) & (g1119)) + ((sk[33]) & (!g2173) & (g3420) & (g1119)) + ((sk[33]) & (g2173) & (g3420) & (!g1119)) + ((sk[33]) & (g2173) & (g3420) & (g1119)));
	assign g4683 = (((!g2174) & (!sk[34]) & (!g3420) & (g1120)) + ((!g2174) & (!sk[34]) & (g3420) & (!g1120)) + ((!g2174) & (!sk[34]) & (g3420) & (g1120)) + ((!g2174) & (sk[34]) & (!g3420) & (g1120)) + ((!g2174) & (sk[34]) & (g3420) & (g1120)) + ((g2174) & (!sk[34]) & (!g3420) & (g1120)) + ((g2174) & (!sk[34]) & (g3420) & (!g1120)) + ((g2174) & (!sk[34]) & (g3420) & (g1120)) + ((g2174) & (sk[34]) & (g3420) & (!g1120)) + ((g2174) & (sk[34]) & (g3420) & (g1120)));
	assign g4684 = (((!sk[35]) & (!g2175) & (!g3420) & (g1121)) + ((!sk[35]) & (!g2175) & (g3420) & (!g1121)) + ((!sk[35]) & (!g2175) & (g3420) & (g1121)) + ((!sk[35]) & (g2175) & (!g3420) & (g1121)) + ((!sk[35]) & (g2175) & (g3420) & (!g1121)) + ((!sk[35]) & (g2175) & (g3420) & (g1121)) + ((sk[35]) & (!g2175) & (!g3420) & (g1121)) + ((sk[35]) & (!g2175) & (g3420) & (g1121)) + ((sk[35]) & (g2175) & (g3420) & (!g1121)) + ((sk[35]) & (g2175) & (g3420) & (g1121)));
	assign g4685 = (((!g2176) & (!sk[36]) & (!g3420) & (g1122)) + ((!g2176) & (!sk[36]) & (g3420) & (!g1122)) + ((!g2176) & (!sk[36]) & (g3420) & (g1122)) + ((!g2176) & (sk[36]) & (!g3420) & (g1122)) + ((!g2176) & (sk[36]) & (g3420) & (g1122)) + ((g2176) & (!sk[36]) & (!g3420) & (g1122)) + ((g2176) & (!sk[36]) & (g3420) & (!g1122)) + ((g2176) & (!sk[36]) & (g3420) & (g1122)) + ((g2176) & (sk[36]) & (g3420) & (!g1122)) + ((g2176) & (sk[36]) & (g3420) & (g1122)));
	assign g1123 = (((!g1119) & (!g1120) & (!g1121) & (g1122) & (g165) & (g166)) + ((!g1119) & (!g1120) & (g1121) & (!g1122) & (!g165) & (g166)) + ((!g1119) & (!g1120) & (g1121) & (g1122) & (!g165) & (g166)) + ((!g1119) & (!g1120) & (g1121) & (g1122) & (g165) & (g166)) + ((!g1119) & (g1120) & (!g1121) & (!g1122) & (g165) & (!g166)) + ((!g1119) & (g1120) & (!g1121) & (g1122) & (g165) & (!g166)) + ((!g1119) & (g1120) & (!g1121) & (g1122) & (g165) & (g166)) + ((!g1119) & (g1120) & (g1121) & (!g1122) & (!g165) & (g166)) + ((!g1119) & (g1120) & (g1121) & (!g1122) & (g165) & (!g166)) + ((!g1119) & (g1120) & (g1121) & (g1122) & (!g165) & (g166)) + ((!g1119) & (g1120) & (g1121) & (g1122) & (g165) & (!g166)) + ((!g1119) & (g1120) & (g1121) & (g1122) & (g165) & (g166)) + ((g1119) & (!g1120) & (!g1121) & (!g1122) & (!g165) & (!g166)) + ((g1119) & (!g1120) & (!g1121) & (g1122) & (!g165) & (!g166)) + ((g1119) & (!g1120) & (!g1121) & (g1122) & (g165) & (g166)) + ((g1119) & (!g1120) & (g1121) & (!g1122) & (!g165) & (!g166)) + ((g1119) & (!g1120) & (g1121) & (!g1122) & (!g165) & (g166)) + ((g1119) & (!g1120) & (g1121) & (g1122) & (!g165) & (!g166)) + ((g1119) & (!g1120) & (g1121) & (g1122) & (!g165) & (g166)) + ((g1119) & (!g1120) & (g1121) & (g1122) & (g165) & (g166)) + ((g1119) & (g1120) & (!g1121) & (!g1122) & (!g165) & (!g166)) + ((g1119) & (g1120) & (!g1121) & (!g1122) & (g165) & (!g166)) + ((g1119) & (g1120) & (!g1121) & (g1122) & (!g165) & (!g166)) + ((g1119) & (g1120) & (!g1121) & (g1122) & (g165) & (!g166)) + ((g1119) & (g1120) & (!g1121) & (g1122) & (g165) & (g166)) + ((g1119) & (g1120) & (g1121) & (!g1122) & (!g165) & (!g166)) + ((g1119) & (g1120) & (g1121) & (!g1122) & (!g165) & (g166)) + ((g1119) & (g1120) & (g1121) & (!g1122) & (g165) & (!g166)) + ((g1119) & (g1120) & (g1121) & (g1122) & (!g165) & (!g166)) + ((g1119) & (g1120) & (g1121) & (g1122) & (!g165) & (g166)) + ((g1119) & (g1120) & (g1121) & (g1122) & (g165) & (!g166)) + ((g1119) & (g1120) & (g1121) & (g1122) & (g165) & (g166)));
	assign g4686 = (((!g2177) & (!sk[38]) & (!g3420) & (g1124)) + ((!g2177) & (!sk[38]) & (g3420) & (!g1124)) + ((!g2177) & (!sk[38]) & (g3420) & (g1124)) + ((!g2177) & (sk[38]) & (!g3420) & (g1124)) + ((!g2177) & (sk[38]) & (g3420) & (g1124)) + ((g2177) & (!sk[38]) & (!g3420) & (g1124)) + ((g2177) & (!sk[38]) & (g3420) & (!g1124)) + ((g2177) & (!sk[38]) & (g3420) & (g1124)) + ((g2177) & (sk[38]) & (g3420) & (!g1124)) + ((g2177) & (sk[38]) & (g3420) & (g1124)));
	assign g4687 = (((!g2178) & (!sk[39]) & (!g3420) & (g1125)) + ((!g2178) & (!sk[39]) & (g3420) & (!g1125)) + ((!g2178) & (!sk[39]) & (g3420) & (g1125)) + ((!g2178) & (sk[39]) & (!g3420) & (g1125)) + ((!g2178) & (sk[39]) & (g3420) & (g1125)) + ((g2178) & (!sk[39]) & (!g3420) & (g1125)) + ((g2178) & (!sk[39]) & (g3420) & (!g1125)) + ((g2178) & (!sk[39]) & (g3420) & (g1125)) + ((g2178) & (sk[39]) & (g3420) & (!g1125)) + ((g2178) & (sk[39]) & (g3420) & (g1125)));
	assign g4688 = (((!g2179) & (!g3420) & (!sk[40]) & (g1126)) + ((!g2179) & (!g3420) & (sk[40]) & (g1126)) + ((!g2179) & (g3420) & (!sk[40]) & (!g1126)) + ((!g2179) & (g3420) & (!sk[40]) & (g1126)) + ((!g2179) & (g3420) & (sk[40]) & (g1126)) + ((g2179) & (!g3420) & (!sk[40]) & (g1126)) + ((g2179) & (g3420) & (!sk[40]) & (!g1126)) + ((g2179) & (g3420) & (!sk[40]) & (g1126)) + ((g2179) & (g3420) & (sk[40]) & (!g1126)) + ((g2179) & (g3420) & (sk[40]) & (g1126)));
	assign g1127 = (((!g165) & (!sk[41]) & (!g166) & (!g1124) & (g1125) & (!g1126)) + ((!g165) & (!sk[41]) & (!g166) & (!g1124) & (g1125) & (g1126)) + ((!g165) & (!sk[41]) & (!g166) & (g1124) & (!g1125) & (!g1126)) + ((!g165) & (!sk[41]) & (!g166) & (g1124) & (!g1125) & (g1126)) + ((!g165) & (!sk[41]) & (!g166) & (g1124) & (g1125) & (!g1126)) + ((!g165) & (!sk[41]) & (!g166) & (g1124) & (g1125) & (g1126)) + ((!g165) & (!sk[41]) & (g166) & (!g1124) & (!g1125) & (!g1126)) + ((!g165) & (!sk[41]) & (g166) & (!g1124) & (!g1125) & (g1126)) + ((!g165) & (!sk[41]) & (g166) & (!g1124) & (g1125) & (!g1126)) + ((!g165) & (!sk[41]) & (g166) & (!g1124) & (g1125) & (g1126)) + ((!g165) & (!sk[41]) & (g166) & (g1124) & (!g1125) & (!g1126)) + ((!g165) & (!sk[41]) & (g166) & (g1124) & (!g1125) & (g1126)) + ((!g165) & (!sk[41]) & (g166) & (g1124) & (g1125) & (!g1126)) + ((!g165) & (!sk[41]) & (g166) & (g1124) & (g1125) & (g1126)) + ((!g165) & (sk[41]) & (g166) & (!g1124) & (!g1125) & (g1126)) + ((!g165) & (sk[41]) & (g166) & (!g1124) & (g1125) & (g1126)) + ((!g165) & (sk[41]) & (g166) & (g1124) & (!g1125) & (g1126)) + ((!g165) & (sk[41]) & (g166) & (g1124) & (g1125) & (g1126)) + ((g165) & (!sk[41]) & (!g166) & (!g1124) & (g1125) & (!g1126)) + ((g165) & (!sk[41]) & (!g166) & (!g1124) & (g1125) & (g1126)) + ((g165) & (!sk[41]) & (!g166) & (g1124) & (!g1125) & (!g1126)) + ((g165) & (!sk[41]) & (!g166) & (g1124) & (!g1125) & (g1126)) + ((g165) & (!sk[41]) & (!g166) & (g1124) & (g1125) & (!g1126)) + ((g165) & (!sk[41]) & (!g166) & (g1124) & (g1125) & (g1126)) + ((g165) & (!sk[41]) & (g166) & (!g1124) & (!g1125) & (!g1126)) + ((g165) & (!sk[41]) & (g166) & (!g1124) & (!g1125) & (g1126)) + ((g165) & (!sk[41]) & (g166) & (!g1124) & (g1125) & (!g1126)) + ((g165) & (!sk[41]) & (g166) & (!g1124) & (g1125) & (g1126)) + ((g165) & (!sk[41]) & (g166) & (g1124) & (!g1125) & (!g1126)) + ((g165) & (!sk[41]) & (g166) & (g1124) & (!g1125) & (g1126)) + ((g165) & (!sk[41]) & (g166) & (g1124) & (g1125) & (!g1126)) + ((g165) & (!sk[41]) & (g166) & (g1124) & (g1125) & (g1126)) + ((g165) & (sk[41]) & (!g166) & (g1124) & (!g1125) & (!g1126)) + ((g165) & (sk[41]) & (!g166) & (g1124) & (!g1125) & (g1126)) + ((g165) & (sk[41]) & (!g166) & (g1124) & (g1125) & (!g1126)) + ((g165) & (sk[41]) & (!g166) & (g1124) & (g1125) & (g1126)) + ((g165) & (sk[41]) & (g166) & (!g1124) & (g1125) & (!g1126)) + ((g165) & (sk[41]) & (g166) & (!g1124) & (g1125) & (g1126)) + ((g165) & (sk[41]) & (g166) & (g1124) & (g1125) & (!g1126)) + ((g165) & (sk[41]) & (g166) & (g1124) & (g1125) & (g1126)));
	assign g4689 = (((!g2162) & (!g3420) & (!sk[42]) & (g1128)) + ((!g2162) & (!g3420) & (sk[42]) & (g1128)) + ((!g2162) & (g3420) & (!sk[42]) & (!g1128)) + ((!g2162) & (g3420) & (!sk[42]) & (g1128)) + ((!g2162) & (g3420) & (sk[42]) & (g1128)) + ((g2162) & (!g3420) & (!sk[42]) & (g1128)) + ((g2162) & (g3420) & (!sk[42]) & (!g1128)) + ((g2162) & (g3420) & (!sk[42]) & (g1128)) + ((g2162) & (g3420) & (sk[42]) & (!g1128)) + ((g2162) & (g3420) & (sk[42]) & (g1128)));
	assign g4690 = (((!g2164) & (!g3420) & (!sk[43]) & (g1129)) + ((!g2164) & (!g3420) & (sk[43]) & (g1129)) + ((!g2164) & (g3420) & (!sk[43]) & (!g1129)) + ((!g2164) & (g3420) & (!sk[43]) & (g1129)) + ((!g2164) & (g3420) & (sk[43]) & (g1129)) + ((g2164) & (!g3420) & (!sk[43]) & (g1129)) + ((g2164) & (g3420) & (!sk[43]) & (!g1129)) + ((g2164) & (g3420) & (!sk[43]) & (g1129)) + ((g2164) & (g3420) & (sk[43]) & (!g1129)) + ((g2164) & (g3420) & (sk[43]) & (g1129)));
	assign g4691 = (((!sk[44]) & (!g2166) & (!g3420) & (g1130)) + ((!sk[44]) & (!g2166) & (g3420) & (!g1130)) + ((!sk[44]) & (!g2166) & (g3420) & (g1130)) + ((!sk[44]) & (g2166) & (!g3420) & (g1130)) + ((!sk[44]) & (g2166) & (g3420) & (!g1130)) + ((!sk[44]) & (g2166) & (g3420) & (g1130)) + ((sk[44]) & (!g2166) & (!g3420) & (g1130)) + ((sk[44]) & (!g2166) & (g3420) & (g1130)) + ((sk[44]) & (g2166) & (g3420) & (!g1130)) + ((sk[44]) & (g2166) & (g3420) & (g1130)));
	assign g4692 = (((!g2168) & (!g3420) & (!sk[45]) & (g1131)) + ((!g2168) & (!g3420) & (sk[45]) & (g1131)) + ((!g2168) & (g3420) & (!sk[45]) & (!g1131)) + ((!g2168) & (g3420) & (!sk[45]) & (g1131)) + ((!g2168) & (g3420) & (sk[45]) & (g1131)) + ((g2168) & (!g3420) & (!sk[45]) & (g1131)) + ((g2168) & (g3420) & (!sk[45]) & (!g1131)) + ((g2168) & (g3420) & (!sk[45]) & (g1131)) + ((g2168) & (g3420) & (sk[45]) & (!g1131)) + ((g2168) & (g3420) & (sk[45]) & (g1131)));
	assign g1132 = (((!g1128) & (!g1129) & (!g1130) & (g1131) & (g165) & (g166)) + ((!g1128) & (!g1129) & (g1130) & (!g1131) & (!g165) & (g166)) + ((!g1128) & (!g1129) & (g1130) & (g1131) & (!g165) & (g166)) + ((!g1128) & (!g1129) & (g1130) & (g1131) & (g165) & (g166)) + ((!g1128) & (g1129) & (!g1130) & (!g1131) & (g165) & (!g166)) + ((!g1128) & (g1129) & (!g1130) & (g1131) & (g165) & (!g166)) + ((!g1128) & (g1129) & (!g1130) & (g1131) & (g165) & (g166)) + ((!g1128) & (g1129) & (g1130) & (!g1131) & (!g165) & (g166)) + ((!g1128) & (g1129) & (g1130) & (!g1131) & (g165) & (!g166)) + ((!g1128) & (g1129) & (g1130) & (g1131) & (!g165) & (g166)) + ((!g1128) & (g1129) & (g1130) & (g1131) & (g165) & (!g166)) + ((!g1128) & (g1129) & (g1130) & (g1131) & (g165) & (g166)) + ((g1128) & (!g1129) & (!g1130) & (!g1131) & (!g165) & (!g166)) + ((g1128) & (!g1129) & (!g1130) & (g1131) & (!g165) & (!g166)) + ((g1128) & (!g1129) & (!g1130) & (g1131) & (g165) & (g166)) + ((g1128) & (!g1129) & (g1130) & (!g1131) & (!g165) & (!g166)) + ((g1128) & (!g1129) & (g1130) & (!g1131) & (!g165) & (g166)) + ((g1128) & (!g1129) & (g1130) & (g1131) & (!g165) & (!g166)) + ((g1128) & (!g1129) & (g1130) & (g1131) & (!g165) & (g166)) + ((g1128) & (!g1129) & (g1130) & (g1131) & (g165) & (g166)) + ((g1128) & (g1129) & (!g1130) & (!g1131) & (!g165) & (!g166)) + ((g1128) & (g1129) & (!g1130) & (!g1131) & (g165) & (!g166)) + ((g1128) & (g1129) & (!g1130) & (g1131) & (!g165) & (!g166)) + ((g1128) & (g1129) & (!g1130) & (g1131) & (g165) & (!g166)) + ((g1128) & (g1129) & (!g1130) & (g1131) & (g165) & (g166)) + ((g1128) & (g1129) & (g1130) & (!g1131) & (!g165) & (!g166)) + ((g1128) & (g1129) & (g1130) & (!g1131) & (!g165) & (g166)) + ((g1128) & (g1129) & (g1130) & (!g1131) & (g165) & (!g166)) + ((g1128) & (g1129) & (g1130) & (g1131) & (!g165) & (!g166)) + ((g1128) & (g1129) & (g1130) & (g1131) & (!g165) & (g166)) + ((g1128) & (g1129) & (g1130) & (g1131) & (g165) & (!g166)) + ((g1128) & (g1129) & (g1130) & (g1131) & (g165) & (g166)));
	assign g4693 = (((!g2169) & (!sk[47]) & (!g3420) & (g1133)) + ((!g2169) & (!sk[47]) & (g3420) & (!g1133)) + ((!g2169) & (!sk[47]) & (g3420) & (g1133)) + ((!g2169) & (sk[47]) & (!g3420) & (g1133)) + ((!g2169) & (sk[47]) & (g3420) & (g1133)) + ((g2169) & (!sk[47]) & (!g3420) & (g1133)) + ((g2169) & (!sk[47]) & (g3420) & (!g1133)) + ((g2169) & (!sk[47]) & (g3420) & (g1133)) + ((g2169) & (sk[47]) & (g3420) & (!g1133)) + ((g2169) & (sk[47]) & (g3420) & (g1133)));
	assign g4694 = (((!g2170) & (!g3420) & (!sk[48]) & (g1134)) + ((!g2170) & (!g3420) & (sk[48]) & (g1134)) + ((!g2170) & (g3420) & (!sk[48]) & (!g1134)) + ((!g2170) & (g3420) & (!sk[48]) & (g1134)) + ((!g2170) & (g3420) & (sk[48]) & (g1134)) + ((g2170) & (!g3420) & (!sk[48]) & (g1134)) + ((g2170) & (g3420) & (!sk[48]) & (!g1134)) + ((g2170) & (g3420) & (!sk[48]) & (g1134)) + ((g2170) & (g3420) & (sk[48]) & (!g1134)) + ((g2170) & (g3420) & (sk[48]) & (g1134)));
	assign g4695 = (((!sk[49]) & (!g2171) & (!g3420) & (g1135)) + ((!sk[49]) & (!g2171) & (g3420) & (!g1135)) + ((!sk[49]) & (!g2171) & (g3420) & (g1135)) + ((!sk[49]) & (g2171) & (!g3420) & (g1135)) + ((!sk[49]) & (g2171) & (g3420) & (!g1135)) + ((!sk[49]) & (g2171) & (g3420) & (g1135)) + ((sk[49]) & (!g2171) & (!g3420) & (g1135)) + ((sk[49]) & (!g2171) & (g3420) & (g1135)) + ((sk[49]) & (g2171) & (g3420) & (!g1135)) + ((sk[49]) & (g2171) & (g3420) & (g1135)));
	assign g4696 = (((!sk[50]) & (!g2172) & (!g3420) & (g1136)) + ((!sk[50]) & (!g2172) & (g3420) & (!g1136)) + ((!sk[50]) & (!g2172) & (g3420) & (g1136)) + ((!sk[50]) & (g2172) & (!g3420) & (g1136)) + ((!sk[50]) & (g2172) & (g3420) & (!g1136)) + ((!sk[50]) & (g2172) & (g3420) & (g1136)) + ((sk[50]) & (!g2172) & (!g3420) & (g1136)) + ((sk[50]) & (!g2172) & (g3420) & (g1136)) + ((sk[50]) & (g2172) & (g3420) & (!g1136)) + ((sk[50]) & (g2172) & (g3420) & (g1136)));
	assign g1137 = (((!g1133) & (!g1134) & (!g1135) & (g1136) & (g165) & (g166)) + ((!g1133) & (!g1134) & (g1135) & (!g1136) & (!g165) & (g166)) + ((!g1133) & (!g1134) & (g1135) & (g1136) & (!g165) & (g166)) + ((!g1133) & (!g1134) & (g1135) & (g1136) & (g165) & (g166)) + ((!g1133) & (g1134) & (!g1135) & (!g1136) & (g165) & (!g166)) + ((!g1133) & (g1134) & (!g1135) & (g1136) & (g165) & (!g166)) + ((!g1133) & (g1134) & (!g1135) & (g1136) & (g165) & (g166)) + ((!g1133) & (g1134) & (g1135) & (!g1136) & (!g165) & (g166)) + ((!g1133) & (g1134) & (g1135) & (!g1136) & (g165) & (!g166)) + ((!g1133) & (g1134) & (g1135) & (g1136) & (!g165) & (g166)) + ((!g1133) & (g1134) & (g1135) & (g1136) & (g165) & (!g166)) + ((!g1133) & (g1134) & (g1135) & (g1136) & (g165) & (g166)) + ((g1133) & (!g1134) & (!g1135) & (!g1136) & (!g165) & (!g166)) + ((g1133) & (!g1134) & (!g1135) & (g1136) & (!g165) & (!g166)) + ((g1133) & (!g1134) & (!g1135) & (g1136) & (g165) & (g166)) + ((g1133) & (!g1134) & (g1135) & (!g1136) & (!g165) & (!g166)) + ((g1133) & (!g1134) & (g1135) & (!g1136) & (!g165) & (g166)) + ((g1133) & (!g1134) & (g1135) & (g1136) & (!g165) & (!g166)) + ((g1133) & (!g1134) & (g1135) & (g1136) & (!g165) & (g166)) + ((g1133) & (!g1134) & (g1135) & (g1136) & (g165) & (g166)) + ((g1133) & (g1134) & (!g1135) & (!g1136) & (!g165) & (!g166)) + ((g1133) & (g1134) & (!g1135) & (!g1136) & (g165) & (!g166)) + ((g1133) & (g1134) & (!g1135) & (g1136) & (!g165) & (!g166)) + ((g1133) & (g1134) & (!g1135) & (g1136) & (g165) & (!g166)) + ((g1133) & (g1134) & (!g1135) & (g1136) & (g165) & (g166)) + ((g1133) & (g1134) & (g1135) & (!g1136) & (!g165) & (!g166)) + ((g1133) & (g1134) & (g1135) & (!g1136) & (!g165) & (g166)) + ((g1133) & (g1134) & (g1135) & (!g1136) & (g165) & (!g166)) + ((g1133) & (g1134) & (g1135) & (g1136) & (!g165) & (!g166)) + ((g1133) & (g1134) & (g1135) & (g1136) & (!g165) & (g166)) + ((g1133) & (g1134) & (g1135) & (g1136) & (g165) & (!g166)) + ((g1133) & (g1134) & (g1135) & (g1136) & (g165) & (g166)));
	assign g1138 = (((!g147) & (!g148) & (!g1123) & (g1127) & (!g1132) & (!g1137)) + ((!g147) & (!g148) & (!g1123) & (g1127) & (!g1132) & (g1137)) + ((!g147) & (!g148) & (!g1123) & (g1127) & (g1132) & (!g1137)) + ((!g147) & (!g148) & (!g1123) & (g1127) & (g1132) & (g1137)) + ((!g147) & (!g148) & (g1123) & (g1127) & (!g1132) & (!g1137)) + ((!g147) & (!g148) & (g1123) & (g1127) & (!g1132) & (g1137)) + ((!g147) & (!g148) & (g1123) & (g1127) & (g1132) & (!g1137)) + ((!g147) & (!g148) & (g1123) & (g1127) & (g1132) & (g1137)) + ((!g147) & (g148) & (!g1123) & (!g1127) & (!g1132) & (g1137)) + ((!g147) & (g148) & (!g1123) & (!g1127) & (g1132) & (g1137)) + ((!g147) & (g148) & (!g1123) & (g1127) & (!g1132) & (g1137)) + ((!g147) & (g148) & (!g1123) & (g1127) & (g1132) & (g1137)) + ((!g147) & (g148) & (g1123) & (!g1127) & (!g1132) & (g1137)) + ((!g147) & (g148) & (g1123) & (!g1127) & (g1132) & (g1137)) + ((!g147) & (g148) & (g1123) & (g1127) & (!g1132) & (g1137)) + ((!g147) & (g148) & (g1123) & (g1127) & (g1132) & (g1137)) + ((g147) & (!g148) & (g1123) & (!g1127) & (!g1132) & (!g1137)) + ((g147) & (!g148) & (g1123) & (!g1127) & (!g1132) & (g1137)) + ((g147) & (!g148) & (g1123) & (!g1127) & (g1132) & (!g1137)) + ((g147) & (!g148) & (g1123) & (!g1127) & (g1132) & (g1137)) + ((g147) & (!g148) & (g1123) & (g1127) & (!g1132) & (!g1137)) + ((g147) & (!g148) & (g1123) & (g1127) & (!g1132) & (g1137)) + ((g147) & (!g148) & (g1123) & (g1127) & (g1132) & (!g1137)) + ((g147) & (!g148) & (g1123) & (g1127) & (g1132) & (g1137)) + ((g147) & (g148) & (!g1123) & (!g1127) & (g1132) & (!g1137)) + ((g147) & (g148) & (!g1123) & (!g1127) & (g1132) & (g1137)) + ((g147) & (g148) & (!g1123) & (g1127) & (g1132) & (!g1137)) + ((g147) & (g148) & (!g1123) & (g1127) & (g1132) & (g1137)) + ((g147) & (g148) & (g1123) & (!g1127) & (g1132) & (!g1137)) + ((g147) & (g148) & (g1123) & (!g1127) & (g1132) & (g1137)) + ((g147) & (g148) & (g1123) & (g1127) & (g1132) & (!g1137)) + ((g147) & (g148) & (g1123) & (g1127) & (g1132) & (g1137)));
	assign g1139 = (((!g142) & (!g1118) & (!sk[53]) & (g1138)) + ((!g142) & (!g1118) & (sk[53]) & (g1138)) + ((!g142) & (g1118) & (!sk[53]) & (!g1138)) + ((!g142) & (g1118) & (!sk[53]) & (g1138)) + ((!g142) & (g1118) & (sk[53]) & (g1138)) + ((g142) & (!g1118) & (!sk[53]) & (g1138)) + ((g142) & (g1118) & (!sk[53]) & (!g1138)) + ((g142) & (g1118) & (!sk[53]) & (g1138)) + ((g142) & (g1118) & (sk[53]) & (!g1138)) + ((g142) & (g1118) & (sk[53]) & (g1138)));
	assign g4697 = (((!g2059) & (!g2659) & (!sk[54]) & (g1140)) + ((!g2059) & (!g2659) & (sk[54]) & (g1140)) + ((!g2059) & (g2659) & (!sk[54]) & (!g1140)) + ((!g2059) & (g2659) & (!sk[54]) & (g1140)) + ((!g2059) & (g2659) & (sk[54]) & (g1140)) + ((g2059) & (!g2659) & (!sk[54]) & (g1140)) + ((g2059) & (g2659) & (!sk[54]) & (!g1140)) + ((g2059) & (g2659) & (!sk[54]) & (g1140)) + ((g2059) & (g2659) & (sk[54]) & (!g1140)) + ((g2059) & (g2659) & (sk[54]) & (g1140)));
	assign g1141 = (((g1094) & (!sk[55]) & (!g916)) + ((g1094) & (!sk[55]) & (g916)) + ((g1094) & (sk[55]) & (!g916)));
	assign g1142 = (((!g126) & (!g1139) & (g1140) & (!g3836) & (!g1141) & (!g916)) + ((!g126) & (!g1139) & (g1140) & (!g3836) & (!g1141) & (g916)) + ((!g126) & (!g1139) & (g1140) & (!g3836) & (g1141) & (!g916)) + ((!g126) & (!g1139) & (g1140) & (!g3836) & (g1141) & (g916)) + ((!g126) & (!g1139) & (g1140) & (g3836) & (!g1141) & (!g916)) + ((!g126) & (!g1139) & (g1140) & (g3836) & (!g1141) & (g916)) + ((!g126) & (!g1139) & (g1140) & (g3836) & (g1141) & (!g916)) + ((!g126) & (!g1139) & (g1140) & (g3836) & (g1141) & (g916)) + ((!g126) & (g1139) & (g1140) & (!g3836) & (!g1141) & (!g916)) + ((!g126) & (g1139) & (g1140) & (!g3836) & (!g1141) & (g916)) + ((!g126) & (g1139) & (g1140) & (!g3836) & (g1141) & (!g916)) + ((!g126) & (g1139) & (g1140) & (!g3836) & (g1141) & (g916)) + ((!g126) & (g1139) & (g1140) & (g3836) & (!g1141) & (!g916)) + ((!g126) & (g1139) & (g1140) & (g3836) & (!g1141) & (g916)) + ((!g126) & (g1139) & (g1140) & (g3836) & (g1141) & (!g916)) + ((!g126) & (g1139) & (g1140) & (g3836) & (g1141) & (g916)) + ((g126) & (!g1139) & (!g1140) & (!g3836) & (!g1141) & (!g916)) + ((g126) & (!g1139) & (!g1140) & (!g3836) & (g1141) & (g916)) + ((g126) & (!g1139) & (!g1140) & (g3836) & (!g1141) & (g916)) + ((g126) & (!g1139) & (!g1140) & (g3836) & (g1141) & (g916)) + ((g126) & (!g1139) & (g1140) & (!g3836) & (!g1141) & (!g916)) + ((g126) & (!g1139) & (g1140) & (!g3836) & (g1141) & (g916)) + ((g126) & (!g1139) & (g1140) & (g3836) & (!g1141) & (g916)) + ((g126) & (!g1139) & (g1140) & (g3836) & (g1141) & (g916)) + ((g126) & (g1139) & (!g1140) & (!g3836) & (!g1141) & (g916)) + ((g126) & (g1139) & (!g1140) & (!g3836) & (g1141) & (!g916)) + ((g126) & (g1139) & (!g1140) & (g3836) & (!g1141) & (!g916)) + ((g126) & (g1139) & (!g1140) & (g3836) & (g1141) & (!g916)) + ((g126) & (g1139) & (g1140) & (!g3836) & (!g1141) & (g916)) + ((g126) & (g1139) & (g1140) & (!g3836) & (g1141) & (!g916)) + ((g126) & (g1139) & (g1140) & (g3836) & (!g1141) & (!g916)) + ((g126) & (g1139) & (g1140) & (g3836) & (g1141) & (!g916)));
	assign g4698 = (((!sk[57]) & (!g2140) & (!g3397) & (g1143)) + ((!sk[57]) & (!g2140) & (g3397) & (!g1143)) + ((!sk[57]) & (!g2140) & (g3397) & (g1143)) + ((!sk[57]) & (g2140) & (!g3397) & (g1143)) + ((!sk[57]) & (g2140) & (g3397) & (!g1143)) + ((!sk[57]) & (g2140) & (g3397) & (g1143)) + ((sk[57]) & (!g2140) & (!g3397) & (g1143)) + ((sk[57]) & (!g2140) & (g3397) & (g1143)) + ((sk[57]) & (g2140) & (g3397) & (!g1143)) + ((sk[57]) & (g2140) & (g3397) & (g1143)));
	assign g4699 = (((!g2142) & (!sk[58]) & (!g3397) & (g1144)) + ((!g2142) & (!sk[58]) & (g3397) & (!g1144)) + ((!g2142) & (!sk[58]) & (g3397) & (g1144)) + ((!g2142) & (sk[58]) & (!g3397) & (g1144)) + ((!g2142) & (sk[58]) & (g3397) & (g1144)) + ((g2142) & (!sk[58]) & (!g3397) & (g1144)) + ((g2142) & (!sk[58]) & (g3397) & (!g1144)) + ((g2142) & (!sk[58]) & (g3397) & (g1144)) + ((g2142) & (sk[58]) & (g3397) & (!g1144)) + ((g2142) & (sk[58]) & (g3397) & (g1144)));
	assign g4700 = (((!g2144) & (!g3397) & (!sk[59]) & (g1145)) + ((!g2144) & (!g3397) & (sk[59]) & (g1145)) + ((!g2144) & (g3397) & (!sk[59]) & (!g1145)) + ((!g2144) & (g3397) & (!sk[59]) & (g1145)) + ((!g2144) & (g3397) & (sk[59]) & (g1145)) + ((g2144) & (!g3397) & (!sk[59]) & (g1145)) + ((g2144) & (g3397) & (!sk[59]) & (!g1145)) + ((g2144) & (g3397) & (!sk[59]) & (g1145)) + ((g2144) & (g3397) & (sk[59]) & (!g1145)) + ((g2144) & (g3397) & (sk[59]) & (g1145)));
	assign g4701 = (((!g2145) & (!g3397) & (!sk[60]) & (g1146)) + ((!g2145) & (!g3397) & (sk[60]) & (g1146)) + ((!g2145) & (g3397) & (!sk[60]) & (!g1146)) + ((!g2145) & (g3397) & (!sk[60]) & (g1146)) + ((!g2145) & (g3397) & (sk[60]) & (g1146)) + ((g2145) & (!g3397) & (!sk[60]) & (g1146)) + ((g2145) & (g3397) & (!sk[60]) & (!g1146)) + ((g2145) & (g3397) & (!sk[60]) & (g1146)) + ((g2145) & (g3397) & (sk[60]) & (!g1146)) + ((g2145) & (g3397) & (sk[60]) & (g1146)));
	assign g1147 = (((!g1143) & (!g1144) & (!g1145) & (g1146) & (g147) & (g148)) + ((!g1143) & (!g1144) & (g1145) & (!g1146) & (!g147) & (g148)) + ((!g1143) & (!g1144) & (g1145) & (g1146) & (!g147) & (g148)) + ((!g1143) & (!g1144) & (g1145) & (g1146) & (g147) & (g148)) + ((!g1143) & (g1144) & (!g1145) & (!g1146) & (g147) & (!g148)) + ((!g1143) & (g1144) & (!g1145) & (g1146) & (g147) & (!g148)) + ((!g1143) & (g1144) & (!g1145) & (g1146) & (g147) & (g148)) + ((!g1143) & (g1144) & (g1145) & (!g1146) & (!g147) & (g148)) + ((!g1143) & (g1144) & (g1145) & (!g1146) & (g147) & (!g148)) + ((!g1143) & (g1144) & (g1145) & (g1146) & (!g147) & (g148)) + ((!g1143) & (g1144) & (g1145) & (g1146) & (g147) & (!g148)) + ((!g1143) & (g1144) & (g1145) & (g1146) & (g147) & (g148)) + ((g1143) & (!g1144) & (!g1145) & (!g1146) & (!g147) & (!g148)) + ((g1143) & (!g1144) & (!g1145) & (g1146) & (!g147) & (!g148)) + ((g1143) & (!g1144) & (!g1145) & (g1146) & (g147) & (g148)) + ((g1143) & (!g1144) & (g1145) & (!g1146) & (!g147) & (!g148)) + ((g1143) & (!g1144) & (g1145) & (!g1146) & (!g147) & (g148)) + ((g1143) & (!g1144) & (g1145) & (g1146) & (!g147) & (!g148)) + ((g1143) & (!g1144) & (g1145) & (g1146) & (!g147) & (g148)) + ((g1143) & (!g1144) & (g1145) & (g1146) & (g147) & (g148)) + ((g1143) & (g1144) & (!g1145) & (!g1146) & (!g147) & (!g148)) + ((g1143) & (g1144) & (!g1145) & (!g1146) & (g147) & (!g148)) + ((g1143) & (g1144) & (!g1145) & (g1146) & (!g147) & (!g148)) + ((g1143) & (g1144) & (!g1145) & (g1146) & (g147) & (!g148)) + ((g1143) & (g1144) & (!g1145) & (g1146) & (g147) & (g148)) + ((g1143) & (g1144) & (g1145) & (!g1146) & (!g147) & (!g148)) + ((g1143) & (g1144) & (g1145) & (!g1146) & (!g147) & (g148)) + ((g1143) & (g1144) & (g1145) & (!g1146) & (g147) & (!g148)) + ((g1143) & (g1144) & (g1145) & (g1146) & (!g147) & (!g148)) + ((g1143) & (g1144) & (g1145) & (g1146) & (!g147) & (g148)) + ((g1143) & (g1144) & (g1145) & (g1146) & (g147) & (!g148)) + ((g1143) & (g1144) & (g1145) & (g1146) & (g147) & (g148)));
	assign g4702 = (((!g2146) & (!sk[62]) & (!g3397) & (g1148)) + ((!g2146) & (!sk[62]) & (g3397) & (!g1148)) + ((!g2146) & (!sk[62]) & (g3397) & (g1148)) + ((!g2146) & (sk[62]) & (!g3397) & (g1148)) + ((!g2146) & (sk[62]) & (g3397) & (g1148)) + ((g2146) & (!sk[62]) & (!g3397) & (g1148)) + ((g2146) & (!sk[62]) & (g3397) & (!g1148)) + ((g2146) & (!sk[62]) & (g3397) & (g1148)) + ((g2146) & (sk[62]) & (g3397) & (!g1148)) + ((g2146) & (sk[62]) & (g3397) & (g1148)));
	assign g4703 = (((!sk[63]) & (!g2148) & (!g3397) & (g1149)) + ((!sk[63]) & (!g2148) & (g3397) & (!g1149)) + ((!sk[63]) & (!g2148) & (g3397) & (g1149)) + ((!sk[63]) & (g2148) & (!g3397) & (g1149)) + ((!sk[63]) & (g2148) & (g3397) & (!g1149)) + ((!sk[63]) & (g2148) & (g3397) & (g1149)) + ((sk[63]) & (!g2148) & (!g3397) & (g1149)) + ((sk[63]) & (!g2148) & (g3397) & (g1149)) + ((sk[63]) & (g2148) & (g3397) & (!g1149)) + ((sk[63]) & (g2148) & (g3397) & (g1149)));
	assign g4704 = (((!sk[64]) & (!g2150) & (!g3397) & (g1150)) + ((!sk[64]) & (!g2150) & (g3397) & (!g1150)) + ((!sk[64]) & (!g2150) & (g3397) & (g1150)) + ((!sk[64]) & (g2150) & (!g3397) & (g1150)) + ((!sk[64]) & (g2150) & (g3397) & (!g1150)) + ((!sk[64]) & (g2150) & (g3397) & (g1150)) + ((sk[64]) & (!g2150) & (!g3397) & (g1150)) + ((sk[64]) & (!g2150) & (g3397) & (g1150)) + ((sk[64]) & (g2150) & (g3397) & (!g1150)) + ((sk[64]) & (g2150) & (g3397) & (g1150)));
	assign g4705 = (((!g2151) & (!g3397) & (!sk[65]) & (g1151)) + ((!g2151) & (!g3397) & (sk[65]) & (g1151)) + ((!g2151) & (g3397) & (!sk[65]) & (!g1151)) + ((!g2151) & (g3397) & (!sk[65]) & (g1151)) + ((!g2151) & (g3397) & (sk[65]) & (g1151)) + ((g2151) & (!g3397) & (!sk[65]) & (g1151)) + ((g2151) & (g3397) & (!sk[65]) & (!g1151)) + ((g2151) & (g3397) & (!sk[65]) & (g1151)) + ((g2151) & (g3397) & (sk[65]) & (!g1151)) + ((g2151) & (g3397) & (sk[65]) & (g1151)));
	assign g1152 = (((!g1148) & (!g1149) & (!g1150) & (g1151) & (g147) & (g148)) + ((!g1148) & (!g1149) & (g1150) & (!g1151) & (!g147) & (g148)) + ((!g1148) & (!g1149) & (g1150) & (g1151) & (!g147) & (g148)) + ((!g1148) & (!g1149) & (g1150) & (g1151) & (g147) & (g148)) + ((!g1148) & (g1149) & (!g1150) & (!g1151) & (g147) & (!g148)) + ((!g1148) & (g1149) & (!g1150) & (g1151) & (g147) & (!g148)) + ((!g1148) & (g1149) & (!g1150) & (g1151) & (g147) & (g148)) + ((!g1148) & (g1149) & (g1150) & (!g1151) & (!g147) & (g148)) + ((!g1148) & (g1149) & (g1150) & (!g1151) & (g147) & (!g148)) + ((!g1148) & (g1149) & (g1150) & (g1151) & (!g147) & (g148)) + ((!g1148) & (g1149) & (g1150) & (g1151) & (g147) & (!g148)) + ((!g1148) & (g1149) & (g1150) & (g1151) & (g147) & (g148)) + ((g1148) & (!g1149) & (!g1150) & (!g1151) & (!g147) & (!g148)) + ((g1148) & (!g1149) & (!g1150) & (g1151) & (!g147) & (!g148)) + ((g1148) & (!g1149) & (!g1150) & (g1151) & (g147) & (g148)) + ((g1148) & (!g1149) & (g1150) & (!g1151) & (!g147) & (!g148)) + ((g1148) & (!g1149) & (g1150) & (!g1151) & (!g147) & (g148)) + ((g1148) & (!g1149) & (g1150) & (g1151) & (!g147) & (!g148)) + ((g1148) & (!g1149) & (g1150) & (g1151) & (!g147) & (g148)) + ((g1148) & (!g1149) & (g1150) & (g1151) & (g147) & (g148)) + ((g1148) & (g1149) & (!g1150) & (!g1151) & (!g147) & (!g148)) + ((g1148) & (g1149) & (!g1150) & (!g1151) & (g147) & (!g148)) + ((g1148) & (g1149) & (!g1150) & (g1151) & (!g147) & (!g148)) + ((g1148) & (g1149) & (!g1150) & (g1151) & (g147) & (!g148)) + ((g1148) & (g1149) & (!g1150) & (g1151) & (g147) & (g148)) + ((g1148) & (g1149) & (g1150) & (!g1151) & (!g147) & (!g148)) + ((g1148) & (g1149) & (g1150) & (!g1151) & (!g147) & (g148)) + ((g1148) & (g1149) & (g1150) & (!g1151) & (g147) & (!g148)) + ((g1148) & (g1149) & (g1150) & (g1151) & (!g147) & (!g148)) + ((g1148) & (g1149) & (g1150) & (g1151) & (!g147) & (g148)) + ((g1148) & (g1149) & (g1150) & (g1151) & (g147) & (!g148)) + ((g1148) & (g1149) & (g1150) & (g1151) & (g147) & (g148)));
	assign g4706 = (((!sk[67]) & (!g2152) & (!g3397) & (g1153)) + ((!sk[67]) & (!g2152) & (g3397) & (!g1153)) + ((!sk[67]) & (!g2152) & (g3397) & (g1153)) + ((!sk[67]) & (g2152) & (!g3397) & (g1153)) + ((!sk[67]) & (g2152) & (g3397) & (!g1153)) + ((!sk[67]) & (g2152) & (g3397) & (g1153)) + ((sk[67]) & (!g2152) & (!g3397) & (g1153)) + ((sk[67]) & (!g2152) & (g3397) & (g1153)) + ((sk[67]) & (g2152) & (g3397) & (!g1153)) + ((sk[67]) & (g2152) & (g3397) & (g1153)));
	assign g4707 = (((!g2153) & (!sk[68]) & (!g3397) & (g1154)) + ((!g2153) & (!sk[68]) & (g3397) & (!g1154)) + ((!g2153) & (!sk[68]) & (g3397) & (g1154)) + ((!g2153) & (sk[68]) & (!g3397) & (g1154)) + ((!g2153) & (sk[68]) & (g3397) & (g1154)) + ((g2153) & (!sk[68]) & (!g3397) & (g1154)) + ((g2153) & (!sk[68]) & (g3397) & (!g1154)) + ((g2153) & (!sk[68]) & (g3397) & (g1154)) + ((g2153) & (sk[68]) & (g3397) & (!g1154)) + ((g2153) & (sk[68]) & (g3397) & (g1154)));
	assign g4708 = (((!g2155) & (!sk[69]) & (!g3397) & (g1155)) + ((!g2155) & (!sk[69]) & (g3397) & (!g1155)) + ((!g2155) & (!sk[69]) & (g3397) & (g1155)) + ((!g2155) & (sk[69]) & (!g3397) & (g1155)) + ((!g2155) & (sk[69]) & (g3397) & (g1155)) + ((g2155) & (!sk[69]) & (!g3397) & (g1155)) + ((g2155) & (!sk[69]) & (g3397) & (!g1155)) + ((g2155) & (!sk[69]) & (g3397) & (g1155)) + ((g2155) & (sk[69]) & (g3397) & (!g1155)) + ((g2155) & (sk[69]) & (g3397) & (g1155)));
	assign g4709 = (((!g2157) & (!g3397) & (!sk[70]) & (g1156)) + ((!g2157) & (!g3397) & (sk[70]) & (g1156)) + ((!g2157) & (g3397) & (!sk[70]) & (!g1156)) + ((!g2157) & (g3397) & (!sk[70]) & (g1156)) + ((!g2157) & (g3397) & (sk[70]) & (g1156)) + ((g2157) & (!g3397) & (!sk[70]) & (g1156)) + ((g2157) & (g3397) & (!sk[70]) & (!g1156)) + ((g2157) & (g3397) & (!sk[70]) & (g1156)) + ((g2157) & (g3397) & (sk[70]) & (!g1156)) + ((g2157) & (g3397) & (sk[70]) & (g1156)));
	assign g1157 = (((!g1153) & (!g1154) & (!g1155) & (g1156) & (g147) & (g148)) + ((!g1153) & (!g1154) & (g1155) & (!g1156) & (!g147) & (g148)) + ((!g1153) & (!g1154) & (g1155) & (g1156) & (!g147) & (g148)) + ((!g1153) & (!g1154) & (g1155) & (g1156) & (g147) & (g148)) + ((!g1153) & (g1154) & (!g1155) & (!g1156) & (g147) & (!g148)) + ((!g1153) & (g1154) & (!g1155) & (g1156) & (g147) & (!g148)) + ((!g1153) & (g1154) & (!g1155) & (g1156) & (g147) & (g148)) + ((!g1153) & (g1154) & (g1155) & (!g1156) & (!g147) & (g148)) + ((!g1153) & (g1154) & (g1155) & (!g1156) & (g147) & (!g148)) + ((!g1153) & (g1154) & (g1155) & (g1156) & (!g147) & (g148)) + ((!g1153) & (g1154) & (g1155) & (g1156) & (g147) & (!g148)) + ((!g1153) & (g1154) & (g1155) & (g1156) & (g147) & (g148)) + ((g1153) & (!g1154) & (!g1155) & (!g1156) & (!g147) & (!g148)) + ((g1153) & (!g1154) & (!g1155) & (g1156) & (!g147) & (!g148)) + ((g1153) & (!g1154) & (!g1155) & (g1156) & (g147) & (g148)) + ((g1153) & (!g1154) & (g1155) & (!g1156) & (!g147) & (!g148)) + ((g1153) & (!g1154) & (g1155) & (!g1156) & (!g147) & (g148)) + ((g1153) & (!g1154) & (g1155) & (g1156) & (!g147) & (!g148)) + ((g1153) & (!g1154) & (g1155) & (g1156) & (!g147) & (g148)) + ((g1153) & (!g1154) & (g1155) & (g1156) & (g147) & (g148)) + ((g1153) & (g1154) & (!g1155) & (!g1156) & (!g147) & (!g148)) + ((g1153) & (g1154) & (!g1155) & (!g1156) & (g147) & (!g148)) + ((g1153) & (g1154) & (!g1155) & (g1156) & (!g147) & (!g148)) + ((g1153) & (g1154) & (!g1155) & (g1156) & (g147) & (!g148)) + ((g1153) & (g1154) & (!g1155) & (g1156) & (g147) & (g148)) + ((g1153) & (g1154) & (g1155) & (!g1156) & (!g147) & (!g148)) + ((g1153) & (g1154) & (g1155) & (!g1156) & (!g147) & (g148)) + ((g1153) & (g1154) & (g1155) & (!g1156) & (g147) & (!g148)) + ((g1153) & (g1154) & (g1155) & (g1156) & (!g147) & (!g148)) + ((g1153) & (g1154) & (g1155) & (g1156) & (!g147) & (g148)) + ((g1153) & (g1154) & (g1155) & (g1156) & (g147) & (!g148)) + ((g1153) & (g1154) & (g1155) & (g1156) & (g147) & (g148)));
	assign g4710 = (((!g2158) & (!g3397) & (!sk[72]) & (g1158)) + ((!g2158) & (!g3397) & (sk[72]) & (g1158)) + ((!g2158) & (g3397) & (!sk[72]) & (!g1158)) + ((!g2158) & (g3397) & (!sk[72]) & (g1158)) + ((!g2158) & (g3397) & (sk[72]) & (g1158)) + ((g2158) & (!g3397) & (!sk[72]) & (g1158)) + ((g2158) & (g3397) & (!sk[72]) & (!g1158)) + ((g2158) & (g3397) & (!sk[72]) & (g1158)) + ((g2158) & (g3397) & (sk[72]) & (!g1158)) + ((g2158) & (g3397) & (sk[72]) & (g1158)));
	assign g4711 = (((!g2159) & (!g3397) & (!sk[73]) & (g1159)) + ((!g2159) & (!g3397) & (sk[73]) & (g1159)) + ((!g2159) & (g3397) & (!sk[73]) & (!g1159)) + ((!g2159) & (g3397) & (!sk[73]) & (g1159)) + ((!g2159) & (g3397) & (sk[73]) & (g1159)) + ((g2159) & (!g3397) & (!sk[73]) & (g1159)) + ((g2159) & (g3397) & (!sk[73]) & (!g1159)) + ((g2159) & (g3397) & (!sk[73]) & (g1159)) + ((g2159) & (g3397) & (sk[73]) & (!g1159)) + ((g2159) & (g3397) & (sk[73]) & (g1159)));
	assign g4712 = (((!g2160) & (!g3397) & (!sk[74]) & (g1160)) + ((!g2160) & (!g3397) & (sk[74]) & (g1160)) + ((!g2160) & (g3397) & (!sk[74]) & (!g1160)) + ((!g2160) & (g3397) & (!sk[74]) & (g1160)) + ((!g2160) & (g3397) & (sk[74]) & (g1160)) + ((g2160) & (!g3397) & (!sk[74]) & (g1160)) + ((g2160) & (g3397) & (!sk[74]) & (!g1160)) + ((g2160) & (g3397) & (!sk[74]) & (g1160)) + ((g2160) & (g3397) & (sk[74]) & (!g1160)) + ((g2160) & (g3397) & (sk[74]) & (g1160)));
	assign g4713 = (((!sk[75]) & (!g2161) & (!g3397) & (g1161)) + ((!sk[75]) & (!g2161) & (g3397) & (!g1161)) + ((!sk[75]) & (!g2161) & (g3397) & (g1161)) + ((!sk[75]) & (g2161) & (!g3397) & (g1161)) + ((!sk[75]) & (g2161) & (g3397) & (!g1161)) + ((!sk[75]) & (g2161) & (g3397) & (g1161)) + ((sk[75]) & (!g2161) & (!g3397) & (g1161)) + ((sk[75]) & (!g2161) & (g3397) & (g1161)) + ((sk[75]) & (g2161) & (g3397) & (!g1161)) + ((sk[75]) & (g2161) & (g3397) & (g1161)));
	assign g1162 = (((!g1158) & (!g1159) & (!g1160) & (g1161) & (g147) & (g148)) + ((!g1158) & (!g1159) & (g1160) & (!g1161) & (!g147) & (g148)) + ((!g1158) & (!g1159) & (g1160) & (g1161) & (!g147) & (g148)) + ((!g1158) & (!g1159) & (g1160) & (g1161) & (g147) & (g148)) + ((!g1158) & (g1159) & (!g1160) & (!g1161) & (g147) & (!g148)) + ((!g1158) & (g1159) & (!g1160) & (g1161) & (g147) & (!g148)) + ((!g1158) & (g1159) & (!g1160) & (g1161) & (g147) & (g148)) + ((!g1158) & (g1159) & (g1160) & (!g1161) & (!g147) & (g148)) + ((!g1158) & (g1159) & (g1160) & (!g1161) & (g147) & (!g148)) + ((!g1158) & (g1159) & (g1160) & (g1161) & (!g147) & (g148)) + ((!g1158) & (g1159) & (g1160) & (g1161) & (g147) & (!g148)) + ((!g1158) & (g1159) & (g1160) & (g1161) & (g147) & (g148)) + ((g1158) & (!g1159) & (!g1160) & (!g1161) & (!g147) & (!g148)) + ((g1158) & (!g1159) & (!g1160) & (g1161) & (!g147) & (!g148)) + ((g1158) & (!g1159) & (!g1160) & (g1161) & (g147) & (g148)) + ((g1158) & (!g1159) & (g1160) & (!g1161) & (!g147) & (!g148)) + ((g1158) & (!g1159) & (g1160) & (!g1161) & (!g147) & (g148)) + ((g1158) & (!g1159) & (g1160) & (g1161) & (!g147) & (!g148)) + ((g1158) & (!g1159) & (g1160) & (g1161) & (!g147) & (g148)) + ((g1158) & (!g1159) & (g1160) & (g1161) & (g147) & (g148)) + ((g1158) & (g1159) & (!g1160) & (!g1161) & (!g147) & (!g148)) + ((g1158) & (g1159) & (!g1160) & (!g1161) & (g147) & (!g148)) + ((g1158) & (g1159) & (!g1160) & (g1161) & (!g147) & (!g148)) + ((g1158) & (g1159) & (!g1160) & (g1161) & (g147) & (!g148)) + ((g1158) & (g1159) & (!g1160) & (g1161) & (g147) & (g148)) + ((g1158) & (g1159) & (g1160) & (!g1161) & (!g147) & (!g148)) + ((g1158) & (g1159) & (g1160) & (!g1161) & (!g147) & (g148)) + ((g1158) & (g1159) & (g1160) & (!g1161) & (g147) & (!g148)) + ((g1158) & (g1159) & (g1160) & (g1161) & (!g147) & (!g148)) + ((g1158) & (g1159) & (g1160) & (g1161) & (!g147) & (g148)) + ((g1158) & (g1159) & (g1160) & (g1161) & (g147) & (!g148)) + ((g1158) & (g1159) & (g1160) & (g1161) & (g147) & (g148)));
	assign g1163 = (((!g1147) & (!g1152) & (!g1157) & (g1162) & (g165) & (g166)) + ((!g1147) & (!g1152) & (g1157) & (!g1162) & (!g165) & (g166)) + ((!g1147) & (!g1152) & (g1157) & (g1162) & (!g165) & (g166)) + ((!g1147) & (!g1152) & (g1157) & (g1162) & (g165) & (g166)) + ((!g1147) & (g1152) & (!g1157) & (!g1162) & (g165) & (!g166)) + ((!g1147) & (g1152) & (!g1157) & (g1162) & (g165) & (!g166)) + ((!g1147) & (g1152) & (!g1157) & (g1162) & (g165) & (g166)) + ((!g1147) & (g1152) & (g1157) & (!g1162) & (!g165) & (g166)) + ((!g1147) & (g1152) & (g1157) & (!g1162) & (g165) & (!g166)) + ((!g1147) & (g1152) & (g1157) & (g1162) & (!g165) & (g166)) + ((!g1147) & (g1152) & (g1157) & (g1162) & (g165) & (!g166)) + ((!g1147) & (g1152) & (g1157) & (g1162) & (g165) & (g166)) + ((g1147) & (!g1152) & (!g1157) & (!g1162) & (!g165) & (!g166)) + ((g1147) & (!g1152) & (!g1157) & (g1162) & (!g165) & (!g166)) + ((g1147) & (!g1152) & (!g1157) & (g1162) & (g165) & (g166)) + ((g1147) & (!g1152) & (g1157) & (!g1162) & (!g165) & (!g166)) + ((g1147) & (!g1152) & (g1157) & (!g1162) & (!g165) & (g166)) + ((g1147) & (!g1152) & (g1157) & (g1162) & (!g165) & (!g166)) + ((g1147) & (!g1152) & (g1157) & (g1162) & (!g165) & (g166)) + ((g1147) & (!g1152) & (g1157) & (g1162) & (g165) & (g166)) + ((g1147) & (g1152) & (!g1157) & (!g1162) & (!g165) & (!g166)) + ((g1147) & (g1152) & (!g1157) & (!g1162) & (g165) & (!g166)) + ((g1147) & (g1152) & (!g1157) & (g1162) & (!g165) & (!g166)) + ((g1147) & (g1152) & (!g1157) & (g1162) & (g165) & (!g166)) + ((g1147) & (g1152) & (!g1157) & (g1162) & (g165) & (g166)) + ((g1147) & (g1152) & (g1157) & (!g1162) & (!g165) & (!g166)) + ((g1147) & (g1152) & (g1157) & (!g1162) & (!g165) & (g166)) + ((g1147) & (g1152) & (g1157) & (!g1162) & (g165) & (!g166)) + ((g1147) & (g1152) & (g1157) & (g1162) & (!g165) & (!g166)) + ((g1147) & (g1152) & (g1157) & (g1162) & (!g165) & (g166)) + ((g1147) & (g1152) & (g1157) & (g1162) & (g165) & (!g166)) + ((g1147) & (g1152) & (g1157) & (g1162) & (g165) & (g166)));
	assign g4714 = (((!g2173) & (!g3397) & (!sk[78]) & (g1164)) + ((!g2173) & (!g3397) & (sk[78]) & (g1164)) + ((!g2173) & (g3397) & (!sk[78]) & (!g1164)) + ((!g2173) & (g3397) & (!sk[78]) & (g1164)) + ((!g2173) & (g3397) & (sk[78]) & (g1164)) + ((g2173) & (!g3397) & (!sk[78]) & (g1164)) + ((g2173) & (g3397) & (!sk[78]) & (!g1164)) + ((g2173) & (g3397) & (!sk[78]) & (g1164)) + ((g2173) & (g3397) & (sk[78]) & (!g1164)) + ((g2173) & (g3397) & (sk[78]) & (g1164)));
	assign g4715 = (((!g2174) & (!g3397) & (!sk[79]) & (g1165)) + ((!g2174) & (!g3397) & (sk[79]) & (g1165)) + ((!g2174) & (g3397) & (!sk[79]) & (!g1165)) + ((!g2174) & (g3397) & (!sk[79]) & (g1165)) + ((!g2174) & (g3397) & (sk[79]) & (g1165)) + ((g2174) & (!g3397) & (!sk[79]) & (g1165)) + ((g2174) & (g3397) & (!sk[79]) & (!g1165)) + ((g2174) & (g3397) & (!sk[79]) & (g1165)) + ((g2174) & (g3397) & (sk[79]) & (!g1165)) + ((g2174) & (g3397) & (sk[79]) & (g1165)));
	assign g4716 = (((!g2175) & (!g3397) & (!sk[80]) & (g1166)) + ((!g2175) & (!g3397) & (sk[80]) & (g1166)) + ((!g2175) & (g3397) & (!sk[80]) & (!g1166)) + ((!g2175) & (g3397) & (!sk[80]) & (g1166)) + ((!g2175) & (g3397) & (sk[80]) & (g1166)) + ((g2175) & (!g3397) & (!sk[80]) & (g1166)) + ((g2175) & (g3397) & (!sk[80]) & (!g1166)) + ((g2175) & (g3397) & (!sk[80]) & (g1166)) + ((g2175) & (g3397) & (sk[80]) & (!g1166)) + ((g2175) & (g3397) & (sk[80]) & (g1166)));
	assign g4717 = (((!g2176) & (!g3397) & (!sk[81]) & (g1167)) + ((!g2176) & (!g3397) & (sk[81]) & (g1167)) + ((!g2176) & (g3397) & (!sk[81]) & (!g1167)) + ((!g2176) & (g3397) & (!sk[81]) & (g1167)) + ((!g2176) & (g3397) & (sk[81]) & (g1167)) + ((g2176) & (!g3397) & (!sk[81]) & (g1167)) + ((g2176) & (g3397) & (!sk[81]) & (!g1167)) + ((g2176) & (g3397) & (!sk[81]) & (g1167)) + ((g2176) & (g3397) & (sk[81]) & (!g1167)) + ((g2176) & (g3397) & (sk[81]) & (g1167)));
	assign g1168 = (((!g1164) & (!g1165) & (!g1166) & (g1167) & (g165) & (g166)) + ((!g1164) & (!g1165) & (g1166) & (!g1167) & (!g165) & (g166)) + ((!g1164) & (!g1165) & (g1166) & (g1167) & (!g165) & (g166)) + ((!g1164) & (!g1165) & (g1166) & (g1167) & (g165) & (g166)) + ((!g1164) & (g1165) & (!g1166) & (!g1167) & (g165) & (!g166)) + ((!g1164) & (g1165) & (!g1166) & (g1167) & (g165) & (!g166)) + ((!g1164) & (g1165) & (!g1166) & (g1167) & (g165) & (g166)) + ((!g1164) & (g1165) & (g1166) & (!g1167) & (!g165) & (g166)) + ((!g1164) & (g1165) & (g1166) & (!g1167) & (g165) & (!g166)) + ((!g1164) & (g1165) & (g1166) & (g1167) & (!g165) & (g166)) + ((!g1164) & (g1165) & (g1166) & (g1167) & (g165) & (!g166)) + ((!g1164) & (g1165) & (g1166) & (g1167) & (g165) & (g166)) + ((g1164) & (!g1165) & (!g1166) & (!g1167) & (!g165) & (!g166)) + ((g1164) & (!g1165) & (!g1166) & (g1167) & (!g165) & (!g166)) + ((g1164) & (!g1165) & (!g1166) & (g1167) & (g165) & (g166)) + ((g1164) & (!g1165) & (g1166) & (!g1167) & (!g165) & (!g166)) + ((g1164) & (!g1165) & (g1166) & (!g1167) & (!g165) & (g166)) + ((g1164) & (!g1165) & (g1166) & (g1167) & (!g165) & (!g166)) + ((g1164) & (!g1165) & (g1166) & (g1167) & (!g165) & (g166)) + ((g1164) & (!g1165) & (g1166) & (g1167) & (g165) & (g166)) + ((g1164) & (g1165) & (!g1166) & (!g1167) & (!g165) & (!g166)) + ((g1164) & (g1165) & (!g1166) & (!g1167) & (g165) & (!g166)) + ((g1164) & (g1165) & (!g1166) & (g1167) & (!g165) & (!g166)) + ((g1164) & (g1165) & (!g1166) & (g1167) & (g165) & (!g166)) + ((g1164) & (g1165) & (!g1166) & (g1167) & (g165) & (g166)) + ((g1164) & (g1165) & (g1166) & (!g1167) & (!g165) & (!g166)) + ((g1164) & (g1165) & (g1166) & (!g1167) & (!g165) & (g166)) + ((g1164) & (g1165) & (g1166) & (!g1167) & (g165) & (!g166)) + ((g1164) & (g1165) & (g1166) & (g1167) & (!g165) & (!g166)) + ((g1164) & (g1165) & (g1166) & (g1167) & (!g165) & (g166)) + ((g1164) & (g1165) & (g1166) & (g1167) & (g165) & (!g166)) + ((g1164) & (g1165) & (g1166) & (g1167) & (g165) & (g166)));
	assign g4718 = (((!g2177) & (!g3397) & (!sk[83]) & (g1169)) + ((!g2177) & (!g3397) & (sk[83]) & (g1169)) + ((!g2177) & (g3397) & (!sk[83]) & (!g1169)) + ((!g2177) & (g3397) & (!sk[83]) & (g1169)) + ((!g2177) & (g3397) & (sk[83]) & (g1169)) + ((g2177) & (!g3397) & (!sk[83]) & (g1169)) + ((g2177) & (g3397) & (!sk[83]) & (!g1169)) + ((g2177) & (g3397) & (!sk[83]) & (g1169)) + ((g2177) & (g3397) & (sk[83]) & (!g1169)) + ((g2177) & (g3397) & (sk[83]) & (g1169)));
	assign g4719 = (((!g2178) & (!sk[84]) & (!g3397) & (g1170)) + ((!g2178) & (!sk[84]) & (g3397) & (!g1170)) + ((!g2178) & (!sk[84]) & (g3397) & (g1170)) + ((!g2178) & (sk[84]) & (!g3397) & (g1170)) + ((!g2178) & (sk[84]) & (g3397) & (g1170)) + ((g2178) & (!sk[84]) & (!g3397) & (g1170)) + ((g2178) & (!sk[84]) & (g3397) & (!g1170)) + ((g2178) & (!sk[84]) & (g3397) & (g1170)) + ((g2178) & (sk[84]) & (g3397) & (!g1170)) + ((g2178) & (sk[84]) & (g3397) & (g1170)));
	assign g4720 = (((!sk[85]) & (!g2179) & (!g3397) & (g1171)) + ((!sk[85]) & (!g2179) & (g3397) & (!g1171)) + ((!sk[85]) & (!g2179) & (g3397) & (g1171)) + ((!sk[85]) & (g2179) & (!g3397) & (g1171)) + ((!sk[85]) & (g2179) & (g3397) & (!g1171)) + ((!sk[85]) & (g2179) & (g3397) & (g1171)) + ((sk[85]) & (!g2179) & (!g3397) & (g1171)) + ((sk[85]) & (!g2179) & (g3397) & (g1171)) + ((sk[85]) & (g2179) & (g3397) & (!g1171)) + ((sk[85]) & (g2179) & (g3397) & (g1171)));
	assign g1172 = (((!g165) & (!g166) & (!g1169) & (g1170) & (!sk[86]) & (!g1171)) + ((!g165) & (!g166) & (!g1169) & (g1170) & (!sk[86]) & (g1171)) + ((!g165) & (!g166) & (g1169) & (!g1170) & (!sk[86]) & (!g1171)) + ((!g165) & (!g166) & (g1169) & (!g1170) & (!sk[86]) & (g1171)) + ((!g165) & (!g166) & (g1169) & (g1170) & (!sk[86]) & (!g1171)) + ((!g165) & (!g166) & (g1169) & (g1170) & (!sk[86]) & (g1171)) + ((!g165) & (g166) & (!g1169) & (!g1170) & (!sk[86]) & (!g1171)) + ((!g165) & (g166) & (!g1169) & (!g1170) & (!sk[86]) & (g1171)) + ((!g165) & (g166) & (!g1169) & (!g1170) & (sk[86]) & (g1171)) + ((!g165) & (g166) & (!g1169) & (g1170) & (!sk[86]) & (!g1171)) + ((!g165) & (g166) & (!g1169) & (g1170) & (!sk[86]) & (g1171)) + ((!g165) & (g166) & (!g1169) & (g1170) & (sk[86]) & (g1171)) + ((!g165) & (g166) & (g1169) & (!g1170) & (!sk[86]) & (!g1171)) + ((!g165) & (g166) & (g1169) & (!g1170) & (!sk[86]) & (g1171)) + ((!g165) & (g166) & (g1169) & (!g1170) & (sk[86]) & (g1171)) + ((!g165) & (g166) & (g1169) & (g1170) & (!sk[86]) & (!g1171)) + ((!g165) & (g166) & (g1169) & (g1170) & (!sk[86]) & (g1171)) + ((!g165) & (g166) & (g1169) & (g1170) & (sk[86]) & (g1171)) + ((g165) & (!g166) & (!g1169) & (g1170) & (!sk[86]) & (!g1171)) + ((g165) & (!g166) & (!g1169) & (g1170) & (!sk[86]) & (g1171)) + ((g165) & (!g166) & (g1169) & (!g1170) & (!sk[86]) & (!g1171)) + ((g165) & (!g166) & (g1169) & (!g1170) & (!sk[86]) & (g1171)) + ((g165) & (!g166) & (g1169) & (!g1170) & (sk[86]) & (!g1171)) + ((g165) & (!g166) & (g1169) & (!g1170) & (sk[86]) & (g1171)) + ((g165) & (!g166) & (g1169) & (g1170) & (!sk[86]) & (!g1171)) + ((g165) & (!g166) & (g1169) & (g1170) & (!sk[86]) & (g1171)) + ((g165) & (!g166) & (g1169) & (g1170) & (sk[86]) & (!g1171)) + ((g165) & (!g166) & (g1169) & (g1170) & (sk[86]) & (g1171)) + ((g165) & (g166) & (!g1169) & (!g1170) & (!sk[86]) & (!g1171)) + ((g165) & (g166) & (!g1169) & (!g1170) & (!sk[86]) & (g1171)) + ((g165) & (g166) & (!g1169) & (g1170) & (!sk[86]) & (!g1171)) + ((g165) & (g166) & (!g1169) & (g1170) & (!sk[86]) & (g1171)) + ((g165) & (g166) & (!g1169) & (g1170) & (sk[86]) & (!g1171)) + ((g165) & (g166) & (!g1169) & (g1170) & (sk[86]) & (g1171)) + ((g165) & (g166) & (g1169) & (!g1170) & (!sk[86]) & (!g1171)) + ((g165) & (g166) & (g1169) & (!g1170) & (!sk[86]) & (g1171)) + ((g165) & (g166) & (g1169) & (g1170) & (!sk[86]) & (!g1171)) + ((g165) & (g166) & (g1169) & (g1170) & (!sk[86]) & (g1171)) + ((g165) & (g166) & (g1169) & (g1170) & (sk[86]) & (!g1171)) + ((g165) & (g166) & (g1169) & (g1170) & (sk[86]) & (g1171)));
	assign g4721 = (((!g2162) & (!g3397) & (!sk[87]) & (g1173)) + ((!g2162) & (!g3397) & (sk[87]) & (g1173)) + ((!g2162) & (g3397) & (!sk[87]) & (!g1173)) + ((!g2162) & (g3397) & (!sk[87]) & (g1173)) + ((!g2162) & (g3397) & (sk[87]) & (g1173)) + ((g2162) & (!g3397) & (!sk[87]) & (g1173)) + ((g2162) & (g3397) & (!sk[87]) & (!g1173)) + ((g2162) & (g3397) & (!sk[87]) & (g1173)) + ((g2162) & (g3397) & (sk[87]) & (!g1173)) + ((g2162) & (g3397) & (sk[87]) & (g1173)));
	assign g4722 = (((!g2164) & (!g3397) & (!sk[88]) & (g1174)) + ((!g2164) & (!g3397) & (sk[88]) & (g1174)) + ((!g2164) & (g3397) & (!sk[88]) & (!g1174)) + ((!g2164) & (g3397) & (!sk[88]) & (g1174)) + ((!g2164) & (g3397) & (sk[88]) & (g1174)) + ((g2164) & (!g3397) & (!sk[88]) & (g1174)) + ((g2164) & (g3397) & (!sk[88]) & (!g1174)) + ((g2164) & (g3397) & (!sk[88]) & (g1174)) + ((g2164) & (g3397) & (sk[88]) & (!g1174)) + ((g2164) & (g3397) & (sk[88]) & (g1174)));
	assign g4723 = (((!g2166) & (!sk[89]) & (!g3397) & (g1175)) + ((!g2166) & (!sk[89]) & (g3397) & (!g1175)) + ((!g2166) & (!sk[89]) & (g3397) & (g1175)) + ((!g2166) & (sk[89]) & (!g3397) & (g1175)) + ((!g2166) & (sk[89]) & (g3397) & (g1175)) + ((g2166) & (!sk[89]) & (!g3397) & (g1175)) + ((g2166) & (!sk[89]) & (g3397) & (!g1175)) + ((g2166) & (!sk[89]) & (g3397) & (g1175)) + ((g2166) & (sk[89]) & (g3397) & (!g1175)) + ((g2166) & (sk[89]) & (g3397) & (g1175)));
	assign g4724 = (((!sk[90]) & (!g2168) & (!g3397) & (g1176)) + ((!sk[90]) & (!g2168) & (g3397) & (!g1176)) + ((!sk[90]) & (!g2168) & (g3397) & (g1176)) + ((!sk[90]) & (g2168) & (!g3397) & (g1176)) + ((!sk[90]) & (g2168) & (g3397) & (!g1176)) + ((!sk[90]) & (g2168) & (g3397) & (g1176)) + ((sk[90]) & (!g2168) & (!g3397) & (g1176)) + ((sk[90]) & (!g2168) & (g3397) & (g1176)) + ((sk[90]) & (g2168) & (g3397) & (!g1176)) + ((sk[90]) & (g2168) & (g3397) & (g1176)));
	assign g1177 = (((!g1173) & (!g1174) & (!g1175) & (g1176) & (g165) & (g166)) + ((!g1173) & (!g1174) & (g1175) & (!g1176) & (!g165) & (g166)) + ((!g1173) & (!g1174) & (g1175) & (g1176) & (!g165) & (g166)) + ((!g1173) & (!g1174) & (g1175) & (g1176) & (g165) & (g166)) + ((!g1173) & (g1174) & (!g1175) & (!g1176) & (g165) & (!g166)) + ((!g1173) & (g1174) & (!g1175) & (g1176) & (g165) & (!g166)) + ((!g1173) & (g1174) & (!g1175) & (g1176) & (g165) & (g166)) + ((!g1173) & (g1174) & (g1175) & (!g1176) & (!g165) & (g166)) + ((!g1173) & (g1174) & (g1175) & (!g1176) & (g165) & (!g166)) + ((!g1173) & (g1174) & (g1175) & (g1176) & (!g165) & (g166)) + ((!g1173) & (g1174) & (g1175) & (g1176) & (g165) & (!g166)) + ((!g1173) & (g1174) & (g1175) & (g1176) & (g165) & (g166)) + ((g1173) & (!g1174) & (!g1175) & (!g1176) & (!g165) & (!g166)) + ((g1173) & (!g1174) & (!g1175) & (g1176) & (!g165) & (!g166)) + ((g1173) & (!g1174) & (!g1175) & (g1176) & (g165) & (g166)) + ((g1173) & (!g1174) & (g1175) & (!g1176) & (!g165) & (!g166)) + ((g1173) & (!g1174) & (g1175) & (!g1176) & (!g165) & (g166)) + ((g1173) & (!g1174) & (g1175) & (g1176) & (!g165) & (!g166)) + ((g1173) & (!g1174) & (g1175) & (g1176) & (!g165) & (g166)) + ((g1173) & (!g1174) & (g1175) & (g1176) & (g165) & (g166)) + ((g1173) & (g1174) & (!g1175) & (!g1176) & (!g165) & (!g166)) + ((g1173) & (g1174) & (!g1175) & (!g1176) & (g165) & (!g166)) + ((g1173) & (g1174) & (!g1175) & (g1176) & (!g165) & (!g166)) + ((g1173) & (g1174) & (!g1175) & (g1176) & (g165) & (!g166)) + ((g1173) & (g1174) & (!g1175) & (g1176) & (g165) & (g166)) + ((g1173) & (g1174) & (g1175) & (!g1176) & (!g165) & (!g166)) + ((g1173) & (g1174) & (g1175) & (!g1176) & (!g165) & (g166)) + ((g1173) & (g1174) & (g1175) & (!g1176) & (g165) & (!g166)) + ((g1173) & (g1174) & (g1175) & (g1176) & (!g165) & (!g166)) + ((g1173) & (g1174) & (g1175) & (g1176) & (!g165) & (g166)) + ((g1173) & (g1174) & (g1175) & (g1176) & (g165) & (!g166)) + ((g1173) & (g1174) & (g1175) & (g1176) & (g165) & (g166)));
	assign g4725 = (((!sk[92]) & (!g2169) & (!g3397) & (g1178)) + ((!sk[92]) & (!g2169) & (g3397) & (!g1178)) + ((!sk[92]) & (!g2169) & (g3397) & (g1178)) + ((!sk[92]) & (g2169) & (!g3397) & (g1178)) + ((!sk[92]) & (g2169) & (g3397) & (!g1178)) + ((!sk[92]) & (g2169) & (g3397) & (g1178)) + ((sk[92]) & (!g2169) & (!g3397) & (g1178)) + ((sk[92]) & (!g2169) & (g3397) & (g1178)) + ((sk[92]) & (g2169) & (g3397) & (!g1178)) + ((sk[92]) & (g2169) & (g3397) & (g1178)));
	assign g4726 = (((!sk[93]) & (!g2170) & (!g3397) & (g1179)) + ((!sk[93]) & (!g2170) & (g3397) & (!g1179)) + ((!sk[93]) & (!g2170) & (g3397) & (g1179)) + ((!sk[93]) & (g2170) & (!g3397) & (g1179)) + ((!sk[93]) & (g2170) & (g3397) & (!g1179)) + ((!sk[93]) & (g2170) & (g3397) & (g1179)) + ((sk[93]) & (!g2170) & (!g3397) & (g1179)) + ((sk[93]) & (!g2170) & (g3397) & (g1179)) + ((sk[93]) & (g2170) & (g3397) & (!g1179)) + ((sk[93]) & (g2170) & (g3397) & (g1179)));
	assign g4727 = (((!g2171) & (!g3397) & (!sk[94]) & (g1180)) + ((!g2171) & (!g3397) & (sk[94]) & (g1180)) + ((!g2171) & (g3397) & (!sk[94]) & (!g1180)) + ((!g2171) & (g3397) & (!sk[94]) & (g1180)) + ((!g2171) & (g3397) & (sk[94]) & (g1180)) + ((g2171) & (!g3397) & (!sk[94]) & (g1180)) + ((g2171) & (g3397) & (!sk[94]) & (!g1180)) + ((g2171) & (g3397) & (!sk[94]) & (g1180)) + ((g2171) & (g3397) & (sk[94]) & (!g1180)) + ((g2171) & (g3397) & (sk[94]) & (g1180)));
	assign g4728 = (((!g2172) & (!g3397) & (!sk[95]) & (g1181)) + ((!g2172) & (!g3397) & (sk[95]) & (g1181)) + ((!g2172) & (g3397) & (!sk[95]) & (!g1181)) + ((!g2172) & (g3397) & (!sk[95]) & (g1181)) + ((!g2172) & (g3397) & (sk[95]) & (g1181)) + ((g2172) & (!g3397) & (!sk[95]) & (g1181)) + ((g2172) & (g3397) & (!sk[95]) & (!g1181)) + ((g2172) & (g3397) & (!sk[95]) & (g1181)) + ((g2172) & (g3397) & (sk[95]) & (!g1181)) + ((g2172) & (g3397) & (sk[95]) & (g1181)));
	assign g1182 = (((!g1178) & (!g1179) & (!g1180) & (g1181) & (g165) & (g166)) + ((!g1178) & (!g1179) & (g1180) & (!g1181) & (!g165) & (g166)) + ((!g1178) & (!g1179) & (g1180) & (g1181) & (!g165) & (g166)) + ((!g1178) & (!g1179) & (g1180) & (g1181) & (g165) & (g166)) + ((!g1178) & (g1179) & (!g1180) & (!g1181) & (g165) & (!g166)) + ((!g1178) & (g1179) & (!g1180) & (g1181) & (g165) & (!g166)) + ((!g1178) & (g1179) & (!g1180) & (g1181) & (g165) & (g166)) + ((!g1178) & (g1179) & (g1180) & (!g1181) & (!g165) & (g166)) + ((!g1178) & (g1179) & (g1180) & (!g1181) & (g165) & (!g166)) + ((!g1178) & (g1179) & (g1180) & (g1181) & (!g165) & (g166)) + ((!g1178) & (g1179) & (g1180) & (g1181) & (g165) & (!g166)) + ((!g1178) & (g1179) & (g1180) & (g1181) & (g165) & (g166)) + ((g1178) & (!g1179) & (!g1180) & (!g1181) & (!g165) & (!g166)) + ((g1178) & (!g1179) & (!g1180) & (g1181) & (!g165) & (!g166)) + ((g1178) & (!g1179) & (!g1180) & (g1181) & (g165) & (g166)) + ((g1178) & (!g1179) & (g1180) & (!g1181) & (!g165) & (!g166)) + ((g1178) & (!g1179) & (g1180) & (!g1181) & (!g165) & (g166)) + ((g1178) & (!g1179) & (g1180) & (g1181) & (!g165) & (!g166)) + ((g1178) & (!g1179) & (g1180) & (g1181) & (!g165) & (g166)) + ((g1178) & (!g1179) & (g1180) & (g1181) & (g165) & (g166)) + ((g1178) & (g1179) & (!g1180) & (!g1181) & (!g165) & (!g166)) + ((g1178) & (g1179) & (!g1180) & (!g1181) & (g165) & (!g166)) + ((g1178) & (g1179) & (!g1180) & (g1181) & (!g165) & (!g166)) + ((g1178) & (g1179) & (!g1180) & (g1181) & (g165) & (!g166)) + ((g1178) & (g1179) & (!g1180) & (g1181) & (g165) & (g166)) + ((g1178) & (g1179) & (g1180) & (!g1181) & (!g165) & (!g166)) + ((g1178) & (g1179) & (g1180) & (!g1181) & (!g165) & (g166)) + ((g1178) & (g1179) & (g1180) & (!g1181) & (g165) & (!g166)) + ((g1178) & (g1179) & (g1180) & (g1181) & (!g165) & (!g166)) + ((g1178) & (g1179) & (g1180) & (g1181) & (!g165) & (g166)) + ((g1178) & (g1179) & (g1180) & (g1181) & (g165) & (!g166)) + ((g1178) & (g1179) & (g1180) & (g1181) & (g165) & (g166)));
	assign g1183 = (((!g147) & (!g148) & (!g1168) & (g1172) & (!g1177) & (!g1182)) + ((!g147) & (!g148) & (!g1168) & (g1172) & (!g1177) & (g1182)) + ((!g147) & (!g148) & (!g1168) & (g1172) & (g1177) & (!g1182)) + ((!g147) & (!g148) & (!g1168) & (g1172) & (g1177) & (g1182)) + ((!g147) & (!g148) & (g1168) & (g1172) & (!g1177) & (!g1182)) + ((!g147) & (!g148) & (g1168) & (g1172) & (!g1177) & (g1182)) + ((!g147) & (!g148) & (g1168) & (g1172) & (g1177) & (!g1182)) + ((!g147) & (!g148) & (g1168) & (g1172) & (g1177) & (g1182)) + ((!g147) & (g148) & (!g1168) & (!g1172) & (!g1177) & (g1182)) + ((!g147) & (g148) & (!g1168) & (!g1172) & (g1177) & (g1182)) + ((!g147) & (g148) & (!g1168) & (g1172) & (!g1177) & (g1182)) + ((!g147) & (g148) & (!g1168) & (g1172) & (g1177) & (g1182)) + ((!g147) & (g148) & (g1168) & (!g1172) & (!g1177) & (g1182)) + ((!g147) & (g148) & (g1168) & (!g1172) & (g1177) & (g1182)) + ((!g147) & (g148) & (g1168) & (g1172) & (!g1177) & (g1182)) + ((!g147) & (g148) & (g1168) & (g1172) & (g1177) & (g1182)) + ((g147) & (!g148) & (g1168) & (!g1172) & (!g1177) & (!g1182)) + ((g147) & (!g148) & (g1168) & (!g1172) & (!g1177) & (g1182)) + ((g147) & (!g148) & (g1168) & (!g1172) & (g1177) & (!g1182)) + ((g147) & (!g148) & (g1168) & (!g1172) & (g1177) & (g1182)) + ((g147) & (!g148) & (g1168) & (g1172) & (!g1177) & (!g1182)) + ((g147) & (!g148) & (g1168) & (g1172) & (!g1177) & (g1182)) + ((g147) & (!g148) & (g1168) & (g1172) & (g1177) & (!g1182)) + ((g147) & (!g148) & (g1168) & (g1172) & (g1177) & (g1182)) + ((g147) & (g148) & (!g1168) & (!g1172) & (g1177) & (!g1182)) + ((g147) & (g148) & (!g1168) & (!g1172) & (g1177) & (g1182)) + ((g147) & (g148) & (!g1168) & (g1172) & (g1177) & (!g1182)) + ((g147) & (g148) & (!g1168) & (g1172) & (g1177) & (g1182)) + ((g147) & (g148) & (g1168) & (!g1172) & (g1177) & (!g1182)) + ((g147) & (g148) & (g1168) & (!g1172) & (g1177) & (g1182)) + ((g147) & (g148) & (g1168) & (g1172) & (g1177) & (!g1182)) + ((g147) & (g148) & (g1168) & (g1172) & (g1177) & (g1182)));
	assign g1184 = (((!g142) & (!g1163) & (!sk[98]) & (g1183)) + ((!g142) & (!g1163) & (sk[98]) & (g1183)) + ((!g142) & (g1163) & (!sk[98]) & (!g1183)) + ((!g142) & (g1163) & (!sk[98]) & (g1183)) + ((!g142) & (g1163) & (sk[98]) & (g1183)) + ((g142) & (!g1163) & (!sk[98]) & (g1183)) + ((g142) & (g1163) & (!sk[98]) & (!g1183)) + ((g142) & (g1163) & (!sk[98]) & (g1183)) + ((g142) & (g1163) & (sk[98]) & (!g1183)) + ((g142) & (g1163) & (sk[98]) & (g1183)));
	assign g4729 = (((!g2059) & (!sk[99]) & (!g2679) & (g1185)) + ((!g2059) & (!sk[99]) & (g2679) & (!g1185)) + ((!g2059) & (!sk[99]) & (g2679) & (g1185)) + ((!g2059) & (sk[99]) & (!g2679) & (g1185)) + ((!g2059) & (sk[99]) & (g2679) & (g1185)) + ((g2059) & (!sk[99]) & (!g2679) & (g1185)) + ((g2059) & (!sk[99]) & (g2679) & (!g1185)) + ((g2059) & (!sk[99]) & (g2679) & (g1185)) + ((g2059) & (sk[99]) & (g2679) & (!g1185)) + ((g2059) & (sk[99]) & (g2679) & (g1185)));
	assign g1186 = (((!g1139) & (!sk[100]) & (!g3836) & (!g1141) & (g916)) + ((!g1139) & (!sk[100]) & (!g3836) & (g1141) & (!g916)) + ((!g1139) & (!sk[100]) & (!g3836) & (g1141) & (g916)) + ((!g1139) & (!sk[100]) & (g3836) & (!g1141) & (!g916)) + ((!g1139) & (!sk[100]) & (g3836) & (!g1141) & (g916)) + ((!g1139) & (!sk[100]) & (g3836) & (g1141) & (!g916)) + ((!g1139) & (!sk[100]) & (g3836) & (g1141) & (g916)) + ((!g1139) & (sk[100]) & (!g3836) & (!g1141) & (!g916)) + ((!g1139) & (sk[100]) & (!g3836) & (!g1141) & (g916)) + ((!g1139) & (sk[100]) & (!g3836) & (g1141) & (g916)) + ((!g1139) & (sk[100]) & (g3836) & (!g1141) & (g916)) + ((!g1139) & (sk[100]) & (g3836) & (g1141) & (g916)) + ((g1139) & (!sk[100]) & (!g3836) & (!g1141) & (g916)) + ((g1139) & (!sk[100]) & (!g3836) & (g1141) & (!g916)) + ((g1139) & (!sk[100]) & (!g3836) & (g1141) & (g916)) + ((g1139) & (!sk[100]) & (g3836) & (!g1141) & (!g916)) + ((g1139) & (!sk[100]) & (g3836) & (!g1141) & (g916)) + ((g1139) & (!sk[100]) & (g3836) & (g1141) & (!g916)) + ((g1139) & (!sk[100]) & (g3836) & (g1141) & (g916)) + ((g1139) & (sk[100]) & (!g3836) & (!g1141) & (g916)));
	assign g1187 = (((!g126) & (!sk[101]) & (!g1184) & (!g1185) & (g1186) & (!g916)) + ((!g126) & (!sk[101]) & (!g1184) & (!g1185) & (g1186) & (g916)) + ((!g126) & (!sk[101]) & (!g1184) & (g1185) & (!g1186) & (!g916)) + ((!g126) & (!sk[101]) & (!g1184) & (g1185) & (!g1186) & (g916)) + ((!g126) & (!sk[101]) & (!g1184) & (g1185) & (g1186) & (!g916)) + ((!g126) & (!sk[101]) & (!g1184) & (g1185) & (g1186) & (g916)) + ((!g126) & (!sk[101]) & (g1184) & (!g1185) & (!g1186) & (!g916)) + ((!g126) & (!sk[101]) & (g1184) & (!g1185) & (!g1186) & (g916)) + ((!g126) & (!sk[101]) & (g1184) & (!g1185) & (g1186) & (!g916)) + ((!g126) & (!sk[101]) & (g1184) & (!g1185) & (g1186) & (g916)) + ((!g126) & (!sk[101]) & (g1184) & (g1185) & (!g1186) & (!g916)) + ((!g126) & (!sk[101]) & (g1184) & (g1185) & (!g1186) & (g916)) + ((!g126) & (!sk[101]) & (g1184) & (g1185) & (g1186) & (!g916)) + ((!g126) & (!sk[101]) & (g1184) & (g1185) & (g1186) & (g916)) + ((!g126) & (sk[101]) & (!g1184) & (g1185) & (!g1186) & (!g916)) + ((!g126) & (sk[101]) & (!g1184) & (g1185) & (!g1186) & (g916)) + ((!g126) & (sk[101]) & (!g1184) & (g1185) & (g1186) & (!g916)) + ((!g126) & (sk[101]) & (!g1184) & (g1185) & (g1186) & (g916)) + ((!g126) & (sk[101]) & (g1184) & (g1185) & (!g1186) & (!g916)) + ((!g126) & (sk[101]) & (g1184) & (g1185) & (!g1186) & (g916)) + ((!g126) & (sk[101]) & (g1184) & (g1185) & (g1186) & (!g916)) + ((!g126) & (sk[101]) & (g1184) & (g1185) & (g1186) & (g916)) + ((g126) & (!sk[101]) & (!g1184) & (!g1185) & (g1186) & (!g916)) + ((g126) & (!sk[101]) & (!g1184) & (!g1185) & (g1186) & (g916)) + ((g126) & (!sk[101]) & (!g1184) & (g1185) & (!g1186) & (!g916)) + ((g126) & (!sk[101]) & (!g1184) & (g1185) & (!g1186) & (g916)) + ((g126) & (!sk[101]) & (!g1184) & (g1185) & (g1186) & (!g916)) + ((g126) & (!sk[101]) & (!g1184) & (g1185) & (g1186) & (g916)) + ((g126) & (!sk[101]) & (g1184) & (!g1185) & (!g1186) & (!g916)) + ((g126) & (!sk[101]) & (g1184) & (!g1185) & (!g1186) & (g916)) + ((g126) & (!sk[101]) & (g1184) & (!g1185) & (g1186) & (!g916)) + ((g126) & (!sk[101]) & (g1184) & (!g1185) & (g1186) & (g916)) + ((g126) & (!sk[101]) & (g1184) & (g1185) & (!g1186) & (!g916)) + ((g126) & (!sk[101]) & (g1184) & (g1185) & (!g1186) & (g916)) + ((g126) & (!sk[101]) & (g1184) & (g1185) & (g1186) & (!g916)) + ((g126) & (!sk[101]) & (g1184) & (g1185) & (g1186) & (g916)) + ((g126) & (sk[101]) & (!g1184) & (!g1185) & (!g1186) & (g916)) + ((g126) & (sk[101]) & (!g1184) & (!g1185) & (g1186) & (!g916)) + ((g126) & (sk[101]) & (!g1184) & (g1185) & (!g1186) & (g916)) + ((g126) & (sk[101]) & (!g1184) & (g1185) & (g1186) & (!g916)) + ((g126) & (sk[101]) & (g1184) & (!g1185) & (!g1186) & (!g916)) + ((g126) & (sk[101]) & (g1184) & (!g1185) & (g1186) & (g916)) + ((g126) & (sk[101]) & (g1184) & (g1185) & (!g1186) & (!g916)) + ((g126) & (sk[101]) & (g1184) & (g1185) & (g1186) & (g916)));
	assign g4730 = (((!g2140) & (!sk[102]) & (!g3373) & (g1188)) + ((!g2140) & (!sk[102]) & (g3373) & (!g1188)) + ((!g2140) & (!sk[102]) & (g3373) & (g1188)) + ((!g2140) & (sk[102]) & (!g3373) & (g1188)) + ((!g2140) & (sk[102]) & (g3373) & (g1188)) + ((g2140) & (!sk[102]) & (!g3373) & (g1188)) + ((g2140) & (!sk[102]) & (g3373) & (!g1188)) + ((g2140) & (!sk[102]) & (g3373) & (g1188)) + ((g2140) & (sk[102]) & (g3373) & (!g1188)) + ((g2140) & (sk[102]) & (g3373) & (g1188)));
	assign g4731 = (((!g2142) & (!g3373) & (!sk[103]) & (g1189)) + ((!g2142) & (!g3373) & (sk[103]) & (g1189)) + ((!g2142) & (g3373) & (!sk[103]) & (!g1189)) + ((!g2142) & (g3373) & (!sk[103]) & (g1189)) + ((!g2142) & (g3373) & (sk[103]) & (g1189)) + ((g2142) & (!g3373) & (!sk[103]) & (g1189)) + ((g2142) & (g3373) & (!sk[103]) & (!g1189)) + ((g2142) & (g3373) & (!sk[103]) & (g1189)) + ((g2142) & (g3373) & (sk[103]) & (!g1189)) + ((g2142) & (g3373) & (sk[103]) & (g1189)));
	assign g4732 = (((!g2144) & (!sk[104]) & (!g3373) & (g1190)) + ((!g2144) & (!sk[104]) & (g3373) & (!g1190)) + ((!g2144) & (!sk[104]) & (g3373) & (g1190)) + ((!g2144) & (sk[104]) & (!g3373) & (g1190)) + ((!g2144) & (sk[104]) & (g3373) & (g1190)) + ((g2144) & (!sk[104]) & (!g3373) & (g1190)) + ((g2144) & (!sk[104]) & (g3373) & (!g1190)) + ((g2144) & (!sk[104]) & (g3373) & (g1190)) + ((g2144) & (sk[104]) & (g3373) & (!g1190)) + ((g2144) & (sk[104]) & (g3373) & (g1190)));
	assign g4733 = (((!g2145) & (!sk[105]) & (!g3373) & (g1191)) + ((!g2145) & (!sk[105]) & (g3373) & (!g1191)) + ((!g2145) & (!sk[105]) & (g3373) & (g1191)) + ((!g2145) & (sk[105]) & (!g3373) & (g1191)) + ((!g2145) & (sk[105]) & (g3373) & (g1191)) + ((g2145) & (!sk[105]) & (!g3373) & (g1191)) + ((g2145) & (!sk[105]) & (g3373) & (!g1191)) + ((g2145) & (!sk[105]) & (g3373) & (g1191)) + ((g2145) & (sk[105]) & (g3373) & (!g1191)) + ((g2145) & (sk[105]) & (g3373) & (g1191)));
	assign g1192 = (((!g1188) & (!g1189) & (!g1190) & (g1191) & (g147) & (g148)) + ((!g1188) & (!g1189) & (g1190) & (!g1191) & (!g147) & (g148)) + ((!g1188) & (!g1189) & (g1190) & (g1191) & (!g147) & (g148)) + ((!g1188) & (!g1189) & (g1190) & (g1191) & (g147) & (g148)) + ((!g1188) & (g1189) & (!g1190) & (!g1191) & (g147) & (!g148)) + ((!g1188) & (g1189) & (!g1190) & (g1191) & (g147) & (!g148)) + ((!g1188) & (g1189) & (!g1190) & (g1191) & (g147) & (g148)) + ((!g1188) & (g1189) & (g1190) & (!g1191) & (!g147) & (g148)) + ((!g1188) & (g1189) & (g1190) & (!g1191) & (g147) & (!g148)) + ((!g1188) & (g1189) & (g1190) & (g1191) & (!g147) & (g148)) + ((!g1188) & (g1189) & (g1190) & (g1191) & (g147) & (!g148)) + ((!g1188) & (g1189) & (g1190) & (g1191) & (g147) & (g148)) + ((g1188) & (!g1189) & (!g1190) & (!g1191) & (!g147) & (!g148)) + ((g1188) & (!g1189) & (!g1190) & (g1191) & (!g147) & (!g148)) + ((g1188) & (!g1189) & (!g1190) & (g1191) & (g147) & (g148)) + ((g1188) & (!g1189) & (g1190) & (!g1191) & (!g147) & (!g148)) + ((g1188) & (!g1189) & (g1190) & (!g1191) & (!g147) & (g148)) + ((g1188) & (!g1189) & (g1190) & (g1191) & (!g147) & (!g148)) + ((g1188) & (!g1189) & (g1190) & (g1191) & (!g147) & (g148)) + ((g1188) & (!g1189) & (g1190) & (g1191) & (g147) & (g148)) + ((g1188) & (g1189) & (!g1190) & (!g1191) & (!g147) & (!g148)) + ((g1188) & (g1189) & (!g1190) & (!g1191) & (g147) & (!g148)) + ((g1188) & (g1189) & (!g1190) & (g1191) & (!g147) & (!g148)) + ((g1188) & (g1189) & (!g1190) & (g1191) & (g147) & (!g148)) + ((g1188) & (g1189) & (!g1190) & (g1191) & (g147) & (g148)) + ((g1188) & (g1189) & (g1190) & (!g1191) & (!g147) & (!g148)) + ((g1188) & (g1189) & (g1190) & (!g1191) & (!g147) & (g148)) + ((g1188) & (g1189) & (g1190) & (!g1191) & (g147) & (!g148)) + ((g1188) & (g1189) & (g1190) & (g1191) & (!g147) & (!g148)) + ((g1188) & (g1189) & (g1190) & (g1191) & (!g147) & (g148)) + ((g1188) & (g1189) & (g1190) & (g1191) & (g147) & (!g148)) + ((g1188) & (g1189) & (g1190) & (g1191) & (g147) & (g148)));
	assign g4734 = (((!sk[107]) & (!g2146) & (!g3373) & (g1193)) + ((!sk[107]) & (!g2146) & (g3373) & (!g1193)) + ((!sk[107]) & (!g2146) & (g3373) & (g1193)) + ((!sk[107]) & (g2146) & (!g3373) & (g1193)) + ((!sk[107]) & (g2146) & (g3373) & (!g1193)) + ((!sk[107]) & (g2146) & (g3373) & (g1193)) + ((sk[107]) & (!g2146) & (!g3373) & (g1193)) + ((sk[107]) & (!g2146) & (g3373) & (g1193)) + ((sk[107]) & (g2146) & (g3373) & (!g1193)) + ((sk[107]) & (g2146) & (g3373) & (g1193)));
	assign g4735 = (((!g2148) & (!g3373) & (!sk[108]) & (g1194)) + ((!g2148) & (!g3373) & (sk[108]) & (g1194)) + ((!g2148) & (g3373) & (!sk[108]) & (!g1194)) + ((!g2148) & (g3373) & (!sk[108]) & (g1194)) + ((!g2148) & (g3373) & (sk[108]) & (g1194)) + ((g2148) & (!g3373) & (!sk[108]) & (g1194)) + ((g2148) & (g3373) & (!sk[108]) & (!g1194)) + ((g2148) & (g3373) & (!sk[108]) & (g1194)) + ((g2148) & (g3373) & (sk[108]) & (!g1194)) + ((g2148) & (g3373) & (sk[108]) & (g1194)));
	assign g4736 = (((!g2150) & (!g3373) & (!sk[109]) & (g1195)) + ((!g2150) & (!g3373) & (sk[109]) & (g1195)) + ((!g2150) & (g3373) & (!sk[109]) & (!g1195)) + ((!g2150) & (g3373) & (!sk[109]) & (g1195)) + ((!g2150) & (g3373) & (sk[109]) & (g1195)) + ((g2150) & (!g3373) & (!sk[109]) & (g1195)) + ((g2150) & (g3373) & (!sk[109]) & (!g1195)) + ((g2150) & (g3373) & (!sk[109]) & (g1195)) + ((g2150) & (g3373) & (sk[109]) & (!g1195)) + ((g2150) & (g3373) & (sk[109]) & (g1195)));
	assign g4737 = (((!g2151) & (!sk[110]) & (!g3373) & (g1196)) + ((!g2151) & (!sk[110]) & (g3373) & (!g1196)) + ((!g2151) & (!sk[110]) & (g3373) & (g1196)) + ((!g2151) & (sk[110]) & (!g3373) & (g1196)) + ((!g2151) & (sk[110]) & (g3373) & (g1196)) + ((g2151) & (!sk[110]) & (!g3373) & (g1196)) + ((g2151) & (!sk[110]) & (g3373) & (!g1196)) + ((g2151) & (!sk[110]) & (g3373) & (g1196)) + ((g2151) & (sk[110]) & (g3373) & (!g1196)) + ((g2151) & (sk[110]) & (g3373) & (g1196)));
	assign g1197 = (((!g1193) & (!g1194) & (!g1195) & (g1196) & (g147) & (g148)) + ((!g1193) & (!g1194) & (g1195) & (!g1196) & (!g147) & (g148)) + ((!g1193) & (!g1194) & (g1195) & (g1196) & (!g147) & (g148)) + ((!g1193) & (!g1194) & (g1195) & (g1196) & (g147) & (g148)) + ((!g1193) & (g1194) & (!g1195) & (!g1196) & (g147) & (!g148)) + ((!g1193) & (g1194) & (!g1195) & (g1196) & (g147) & (!g148)) + ((!g1193) & (g1194) & (!g1195) & (g1196) & (g147) & (g148)) + ((!g1193) & (g1194) & (g1195) & (!g1196) & (!g147) & (g148)) + ((!g1193) & (g1194) & (g1195) & (!g1196) & (g147) & (!g148)) + ((!g1193) & (g1194) & (g1195) & (g1196) & (!g147) & (g148)) + ((!g1193) & (g1194) & (g1195) & (g1196) & (g147) & (!g148)) + ((!g1193) & (g1194) & (g1195) & (g1196) & (g147) & (g148)) + ((g1193) & (!g1194) & (!g1195) & (!g1196) & (!g147) & (!g148)) + ((g1193) & (!g1194) & (!g1195) & (g1196) & (!g147) & (!g148)) + ((g1193) & (!g1194) & (!g1195) & (g1196) & (g147) & (g148)) + ((g1193) & (!g1194) & (g1195) & (!g1196) & (!g147) & (!g148)) + ((g1193) & (!g1194) & (g1195) & (!g1196) & (!g147) & (g148)) + ((g1193) & (!g1194) & (g1195) & (g1196) & (!g147) & (!g148)) + ((g1193) & (!g1194) & (g1195) & (g1196) & (!g147) & (g148)) + ((g1193) & (!g1194) & (g1195) & (g1196) & (g147) & (g148)) + ((g1193) & (g1194) & (!g1195) & (!g1196) & (!g147) & (!g148)) + ((g1193) & (g1194) & (!g1195) & (!g1196) & (g147) & (!g148)) + ((g1193) & (g1194) & (!g1195) & (g1196) & (!g147) & (!g148)) + ((g1193) & (g1194) & (!g1195) & (g1196) & (g147) & (!g148)) + ((g1193) & (g1194) & (!g1195) & (g1196) & (g147) & (g148)) + ((g1193) & (g1194) & (g1195) & (!g1196) & (!g147) & (!g148)) + ((g1193) & (g1194) & (g1195) & (!g1196) & (!g147) & (g148)) + ((g1193) & (g1194) & (g1195) & (!g1196) & (g147) & (!g148)) + ((g1193) & (g1194) & (g1195) & (g1196) & (!g147) & (!g148)) + ((g1193) & (g1194) & (g1195) & (g1196) & (!g147) & (g148)) + ((g1193) & (g1194) & (g1195) & (g1196) & (g147) & (!g148)) + ((g1193) & (g1194) & (g1195) & (g1196) & (g147) & (g148)));
	assign g4738 = (((!sk[112]) & (!g2152) & (!g3373) & (g1198)) + ((!sk[112]) & (!g2152) & (g3373) & (!g1198)) + ((!sk[112]) & (!g2152) & (g3373) & (g1198)) + ((!sk[112]) & (g2152) & (!g3373) & (g1198)) + ((!sk[112]) & (g2152) & (g3373) & (!g1198)) + ((!sk[112]) & (g2152) & (g3373) & (g1198)) + ((sk[112]) & (!g2152) & (!g3373) & (g1198)) + ((sk[112]) & (!g2152) & (g3373) & (g1198)) + ((sk[112]) & (g2152) & (g3373) & (!g1198)) + ((sk[112]) & (g2152) & (g3373) & (g1198)));
	assign g4739 = (((!sk[113]) & (!g2153) & (!g3373) & (g1199)) + ((!sk[113]) & (!g2153) & (g3373) & (!g1199)) + ((!sk[113]) & (!g2153) & (g3373) & (g1199)) + ((!sk[113]) & (g2153) & (!g3373) & (g1199)) + ((!sk[113]) & (g2153) & (g3373) & (!g1199)) + ((!sk[113]) & (g2153) & (g3373) & (g1199)) + ((sk[113]) & (!g2153) & (!g3373) & (g1199)) + ((sk[113]) & (!g2153) & (g3373) & (g1199)) + ((sk[113]) & (g2153) & (g3373) & (!g1199)) + ((sk[113]) & (g2153) & (g3373) & (g1199)));
	assign g4740 = (((!sk[114]) & (!g2155) & (!g3373) & (g1200)) + ((!sk[114]) & (!g2155) & (g3373) & (!g1200)) + ((!sk[114]) & (!g2155) & (g3373) & (g1200)) + ((!sk[114]) & (g2155) & (!g3373) & (g1200)) + ((!sk[114]) & (g2155) & (g3373) & (!g1200)) + ((!sk[114]) & (g2155) & (g3373) & (g1200)) + ((sk[114]) & (!g2155) & (!g3373) & (g1200)) + ((sk[114]) & (!g2155) & (g3373) & (g1200)) + ((sk[114]) & (g2155) & (g3373) & (!g1200)) + ((sk[114]) & (g2155) & (g3373) & (g1200)));
	assign g4741 = (((!g2157) & (!g3373) & (!sk[115]) & (g1201)) + ((!g2157) & (!g3373) & (sk[115]) & (g1201)) + ((!g2157) & (g3373) & (!sk[115]) & (!g1201)) + ((!g2157) & (g3373) & (!sk[115]) & (g1201)) + ((!g2157) & (g3373) & (sk[115]) & (g1201)) + ((g2157) & (!g3373) & (!sk[115]) & (g1201)) + ((g2157) & (g3373) & (!sk[115]) & (!g1201)) + ((g2157) & (g3373) & (!sk[115]) & (g1201)) + ((g2157) & (g3373) & (sk[115]) & (!g1201)) + ((g2157) & (g3373) & (sk[115]) & (g1201)));
	assign g1202 = (((!g1198) & (!g1199) & (!g1200) & (g1201) & (g147) & (g148)) + ((!g1198) & (!g1199) & (g1200) & (!g1201) & (!g147) & (g148)) + ((!g1198) & (!g1199) & (g1200) & (g1201) & (!g147) & (g148)) + ((!g1198) & (!g1199) & (g1200) & (g1201) & (g147) & (g148)) + ((!g1198) & (g1199) & (!g1200) & (!g1201) & (g147) & (!g148)) + ((!g1198) & (g1199) & (!g1200) & (g1201) & (g147) & (!g148)) + ((!g1198) & (g1199) & (!g1200) & (g1201) & (g147) & (g148)) + ((!g1198) & (g1199) & (g1200) & (!g1201) & (!g147) & (g148)) + ((!g1198) & (g1199) & (g1200) & (!g1201) & (g147) & (!g148)) + ((!g1198) & (g1199) & (g1200) & (g1201) & (!g147) & (g148)) + ((!g1198) & (g1199) & (g1200) & (g1201) & (g147) & (!g148)) + ((!g1198) & (g1199) & (g1200) & (g1201) & (g147) & (g148)) + ((g1198) & (!g1199) & (!g1200) & (!g1201) & (!g147) & (!g148)) + ((g1198) & (!g1199) & (!g1200) & (g1201) & (!g147) & (!g148)) + ((g1198) & (!g1199) & (!g1200) & (g1201) & (g147) & (g148)) + ((g1198) & (!g1199) & (g1200) & (!g1201) & (!g147) & (!g148)) + ((g1198) & (!g1199) & (g1200) & (!g1201) & (!g147) & (g148)) + ((g1198) & (!g1199) & (g1200) & (g1201) & (!g147) & (!g148)) + ((g1198) & (!g1199) & (g1200) & (g1201) & (!g147) & (g148)) + ((g1198) & (!g1199) & (g1200) & (g1201) & (g147) & (g148)) + ((g1198) & (g1199) & (!g1200) & (!g1201) & (!g147) & (!g148)) + ((g1198) & (g1199) & (!g1200) & (!g1201) & (g147) & (!g148)) + ((g1198) & (g1199) & (!g1200) & (g1201) & (!g147) & (!g148)) + ((g1198) & (g1199) & (!g1200) & (g1201) & (g147) & (!g148)) + ((g1198) & (g1199) & (!g1200) & (g1201) & (g147) & (g148)) + ((g1198) & (g1199) & (g1200) & (!g1201) & (!g147) & (!g148)) + ((g1198) & (g1199) & (g1200) & (!g1201) & (!g147) & (g148)) + ((g1198) & (g1199) & (g1200) & (!g1201) & (g147) & (!g148)) + ((g1198) & (g1199) & (g1200) & (g1201) & (!g147) & (!g148)) + ((g1198) & (g1199) & (g1200) & (g1201) & (!g147) & (g148)) + ((g1198) & (g1199) & (g1200) & (g1201) & (g147) & (!g148)) + ((g1198) & (g1199) & (g1200) & (g1201) & (g147) & (g148)));
	assign g4742 = (((!g2158) & (!sk[117]) & (!g3373) & (g1203)) + ((!g2158) & (!sk[117]) & (g3373) & (!g1203)) + ((!g2158) & (!sk[117]) & (g3373) & (g1203)) + ((!g2158) & (sk[117]) & (!g3373) & (g1203)) + ((!g2158) & (sk[117]) & (g3373) & (g1203)) + ((g2158) & (!sk[117]) & (!g3373) & (g1203)) + ((g2158) & (!sk[117]) & (g3373) & (!g1203)) + ((g2158) & (!sk[117]) & (g3373) & (g1203)) + ((g2158) & (sk[117]) & (g3373) & (!g1203)) + ((g2158) & (sk[117]) & (g3373) & (g1203)));
	assign g4743 = (((!g2159) & (!g3373) & (!sk[118]) & (g1204)) + ((!g2159) & (!g3373) & (sk[118]) & (g1204)) + ((!g2159) & (g3373) & (!sk[118]) & (!g1204)) + ((!g2159) & (g3373) & (!sk[118]) & (g1204)) + ((!g2159) & (g3373) & (sk[118]) & (g1204)) + ((g2159) & (!g3373) & (!sk[118]) & (g1204)) + ((g2159) & (g3373) & (!sk[118]) & (!g1204)) + ((g2159) & (g3373) & (!sk[118]) & (g1204)) + ((g2159) & (g3373) & (sk[118]) & (!g1204)) + ((g2159) & (g3373) & (sk[118]) & (g1204)));
	assign g4744 = (((!g2160) & (!sk[119]) & (!g3373) & (g1205)) + ((!g2160) & (!sk[119]) & (g3373) & (!g1205)) + ((!g2160) & (!sk[119]) & (g3373) & (g1205)) + ((!g2160) & (sk[119]) & (!g3373) & (g1205)) + ((!g2160) & (sk[119]) & (g3373) & (g1205)) + ((g2160) & (!sk[119]) & (!g3373) & (g1205)) + ((g2160) & (!sk[119]) & (g3373) & (!g1205)) + ((g2160) & (!sk[119]) & (g3373) & (g1205)) + ((g2160) & (sk[119]) & (g3373) & (!g1205)) + ((g2160) & (sk[119]) & (g3373) & (g1205)));
	assign g4745 = (((!sk[120]) & (!g2161) & (!g3373) & (g1206)) + ((!sk[120]) & (!g2161) & (g3373) & (!g1206)) + ((!sk[120]) & (!g2161) & (g3373) & (g1206)) + ((!sk[120]) & (g2161) & (!g3373) & (g1206)) + ((!sk[120]) & (g2161) & (g3373) & (!g1206)) + ((!sk[120]) & (g2161) & (g3373) & (g1206)) + ((sk[120]) & (!g2161) & (!g3373) & (g1206)) + ((sk[120]) & (!g2161) & (g3373) & (g1206)) + ((sk[120]) & (g2161) & (g3373) & (!g1206)) + ((sk[120]) & (g2161) & (g3373) & (g1206)));
	assign g1207 = (((!g1203) & (!g1204) & (!g1205) & (g1206) & (g147) & (g148)) + ((!g1203) & (!g1204) & (g1205) & (!g1206) & (!g147) & (g148)) + ((!g1203) & (!g1204) & (g1205) & (g1206) & (!g147) & (g148)) + ((!g1203) & (!g1204) & (g1205) & (g1206) & (g147) & (g148)) + ((!g1203) & (g1204) & (!g1205) & (!g1206) & (g147) & (!g148)) + ((!g1203) & (g1204) & (!g1205) & (g1206) & (g147) & (!g148)) + ((!g1203) & (g1204) & (!g1205) & (g1206) & (g147) & (g148)) + ((!g1203) & (g1204) & (g1205) & (!g1206) & (!g147) & (g148)) + ((!g1203) & (g1204) & (g1205) & (!g1206) & (g147) & (!g148)) + ((!g1203) & (g1204) & (g1205) & (g1206) & (!g147) & (g148)) + ((!g1203) & (g1204) & (g1205) & (g1206) & (g147) & (!g148)) + ((!g1203) & (g1204) & (g1205) & (g1206) & (g147) & (g148)) + ((g1203) & (!g1204) & (!g1205) & (!g1206) & (!g147) & (!g148)) + ((g1203) & (!g1204) & (!g1205) & (g1206) & (!g147) & (!g148)) + ((g1203) & (!g1204) & (!g1205) & (g1206) & (g147) & (g148)) + ((g1203) & (!g1204) & (g1205) & (!g1206) & (!g147) & (!g148)) + ((g1203) & (!g1204) & (g1205) & (!g1206) & (!g147) & (g148)) + ((g1203) & (!g1204) & (g1205) & (g1206) & (!g147) & (!g148)) + ((g1203) & (!g1204) & (g1205) & (g1206) & (!g147) & (g148)) + ((g1203) & (!g1204) & (g1205) & (g1206) & (g147) & (g148)) + ((g1203) & (g1204) & (!g1205) & (!g1206) & (!g147) & (!g148)) + ((g1203) & (g1204) & (!g1205) & (!g1206) & (g147) & (!g148)) + ((g1203) & (g1204) & (!g1205) & (g1206) & (!g147) & (!g148)) + ((g1203) & (g1204) & (!g1205) & (g1206) & (g147) & (!g148)) + ((g1203) & (g1204) & (!g1205) & (g1206) & (g147) & (g148)) + ((g1203) & (g1204) & (g1205) & (!g1206) & (!g147) & (!g148)) + ((g1203) & (g1204) & (g1205) & (!g1206) & (!g147) & (g148)) + ((g1203) & (g1204) & (g1205) & (!g1206) & (g147) & (!g148)) + ((g1203) & (g1204) & (g1205) & (g1206) & (!g147) & (!g148)) + ((g1203) & (g1204) & (g1205) & (g1206) & (!g147) & (g148)) + ((g1203) & (g1204) & (g1205) & (g1206) & (g147) & (!g148)) + ((g1203) & (g1204) & (g1205) & (g1206) & (g147) & (g148)));
	assign g1208 = (((!g1192) & (!g1197) & (!g1202) & (g1207) & (g165) & (g166)) + ((!g1192) & (!g1197) & (g1202) & (!g1207) & (!g165) & (g166)) + ((!g1192) & (!g1197) & (g1202) & (g1207) & (!g165) & (g166)) + ((!g1192) & (!g1197) & (g1202) & (g1207) & (g165) & (g166)) + ((!g1192) & (g1197) & (!g1202) & (!g1207) & (g165) & (!g166)) + ((!g1192) & (g1197) & (!g1202) & (g1207) & (g165) & (!g166)) + ((!g1192) & (g1197) & (!g1202) & (g1207) & (g165) & (g166)) + ((!g1192) & (g1197) & (g1202) & (!g1207) & (!g165) & (g166)) + ((!g1192) & (g1197) & (g1202) & (!g1207) & (g165) & (!g166)) + ((!g1192) & (g1197) & (g1202) & (g1207) & (!g165) & (g166)) + ((!g1192) & (g1197) & (g1202) & (g1207) & (g165) & (!g166)) + ((!g1192) & (g1197) & (g1202) & (g1207) & (g165) & (g166)) + ((g1192) & (!g1197) & (!g1202) & (!g1207) & (!g165) & (!g166)) + ((g1192) & (!g1197) & (!g1202) & (g1207) & (!g165) & (!g166)) + ((g1192) & (!g1197) & (!g1202) & (g1207) & (g165) & (g166)) + ((g1192) & (!g1197) & (g1202) & (!g1207) & (!g165) & (!g166)) + ((g1192) & (!g1197) & (g1202) & (!g1207) & (!g165) & (g166)) + ((g1192) & (!g1197) & (g1202) & (g1207) & (!g165) & (!g166)) + ((g1192) & (!g1197) & (g1202) & (g1207) & (!g165) & (g166)) + ((g1192) & (!g1197) & (g1202) & (g1207) & (g165) & (g166)) + ((g1192) & (g1197) & (!g1202) & (!g1207) & (!g165) & (!g166)) + ((g1192) & (g1197) & (!g1202) & (!g1207) & (g165) & (!g166)) + ((g1192) & (g1197) & (!g1202) & (g1207) & (!g165) & (!g166)) + ((g1192) & (g1197) & (!g1202) & (g1207) & (g165) & (!g166)) + ((g1192) & (g1197) & (!g1202) & (g1207) & (g165) & (g166)) + ((g1192) & (g1197) & (g1202) & (!g1207) & (!g165) & (!g166)) + ((g1192) & (g1197) & (g1202) & (!g1207) & (!g165) & (g166)) + ((g1192) & (g1197) & (g1202) & (!g1207) & (g165) & (!g166)) + ((g1192) & (g1197) & (g1202) & (g1207) & (!g165) & (!g166)) + ((g1192) & (g1197) & (g1202) & (g1207) & (!g165) & (g166)) + ((g1192) & (g1197) & (g1202) & (g1207) & (g165) & (!g166)) + ((g1192) & (g1197) & (g1202) & (g1207) & (g165) & (g166)));
	assign g4746 = (((!g2173) & (!g3373) & (!sk[123]) & (g1209)) + ((!g2173) & (!g3373) & (sk[123]) & (g1209)) + ((!g2173) & (g3373) & (!sk[123]) & (!g1209)) + ((!g2173) & (g3373) & (!sk[123]) & (g1209)) + ((!g2173) & (g3373) & (sk[123]) & (g1209)) + ((g2173) & (!g3373) & (!sk[123]) & (g1209)) + ((g2173) & (g3373) & (!sk[123]) & (!g1209)) + ((g2173) & (g3373) & (!sk[123]) & (g1209)) + ((g2173) & (g3373) & (sk[123]) & (!g1209)) + ((g2173) & (g3373) & (sk[123]) & (g1209)));
	assign g4747 = (((!sk[124]) & (!g2174) & (!g3373) & (g1210)) + ((!sk[124]) & (!g2174) & (g3373) & (!g1210)) + ((!sk[124]) & (!g2174) & (g3373) & (g1210)) + ((!sk[124]) & (g2174) & (!g3373) & (g1210)) + ((!sk[124]) & (g2174) & (g3373) & (!g1210)) + ((!sk[124]) & (g2174) & (g3373) & (g1210)) + ((sk[124]) & (!g2174) & (!g3373) & (g1210)) + ((sk[124]) & (!g2174) & (g3373) & (g1210)) + ((sk[124]) & (g2174) & (g3373) & (!g1210)) + ((sk[124]) & (g2174) & (g3373) & (g1210)));
	assign g4748 = (((!g2175) & (!g3373) & (!sk[125]) & (g1211)) + ((!g2175) & (!g3373) & (sk[125]) & (g1211)) + ((!g2175) & (g3373) & (!sk[125]) & (!g1211)) + ((!g2175) & (g3373) & (!sk[125]) & (g1211)) + ((!g2175) & (g3373) & (sk[125]) & (g1211)) + ((g2175) & (!g3373) & (!sk[125]) & (g1211)) + ((g2175) & (g3373) & (!sk[125]) & (!g1211)) + ((g2175) & (g3373) & (!sk[125]) & (g1211)) + ((g2175) & (g3373) & (sk[125]) & (!g1211)) + ((g2175) & (g3373) & (sk[125]) & (g1211)));
	assign g4749 = (((!g2176) & (!g3373) & (!sk[126]) & (g1212)) + ((!g2176) & (!g3373) & (sk[126]) & (g1212)) + ((!g2176) & (g3373) & (!sk[126]) & (!g1212)) + ((!g2176) & (g3373) & (!sk[126]) & (g1212)) + ((!g2176) & (g3373) & (sk[126]) & (g1212)) + ((g2176) & (!g3373) & (!sk[126]) & (g1212)) + ((g2176) & (g3373) & (!sk[126]) & (!g1212)) + ((g2176) & (g3373) & (!sk[126]) & (g1212)) + ((g2176) & (g3373) & (sk[126]) & (!g1212)) + ((g2176) & (g3373) & (sk[126]) & (g1212)));
	assign g1213 = (((!g1209) & (!g1210) & (!g1211) & (g1212) & (g165) & (g166)) + ((!g1209) & (!g1210) & (g1211) & (!g1212) & (!g165) & (g166)) + ((!g1209) & (!g1210) & (g1211) & (g1212) & (!g165) & (g166)) + ((!g1209) & (!g1210) & (g1211) & (g1212) & (g165) & (g166)) + ((!g1209) & (g1210) & (!g1211) & (!g1212) & (g165) & (!g166)) + ((!g1209) & (g1210) & (!g1211) & (g1212) & (g165) & (!g166)) + ((!g1209) & (g1210) & (!g1211) & (g1212) & (g165) & (g166)) + ((!g1209) & (g1210) & (g1211) & (!g1212) & (!g165) & (g166)) + ((!g1209) & (g1210) & (g1211) & (!g1212) & (g165) & (!g166)) + ((!g1209) & (g1210) & (g1211) & (g1212) & (!g165) & (g166)) + ((!g1209) & (g1210) & (g1211) & (g1212) & (g165) & (!g166)) + ((!g1209) & (g1210) & (g1211) & (g1212) & (g165) & (g166)) + ((g1209) & (!g1210) & (!g1211) & (!g1212) & (!g165) & (!g166)) + ((g1209) & (!g1210) & (!g1211) & (g1212) & (!g165) & (!g166)) + ((g1209) & (!g1210) & (!g1211) & (g1212) & (g165) & (g166)) + ((g1209) & (!g1210) & (g1211) & (!g1212) & (!g165) & (!g166)) + ((g1209) & (!g1210) & (g1211) & (!g1212) & (!g165) & (g166)) + ((g1209) & (!g1210) & (g1211) & (g1212) & (!g165) & (!g166)) + ((g1209) & (!g1210) & (g1211) & (g1212) & (!g165) & (g166)) + ((g1209) & (!g1210) & (g1211) & (g1212) & (g165) & (g166)) + ((g1209) & (g1210) & (!g1211) & (!g1212) & (!g165) & (!g166)) + ((g1209) & (g1210) & (!g1211) & (!g1212) & (g165) & (!g166)) + ((g1209) & (g1210) & (!g1211) & (g1212) & (!g165) & (!g166)) + ((g1209) & (g1210) & (!g1211) & (g1212) & (g165) & (!g166)) + ((g1209) & (g1210) & (!g1211) & (g1212) & (g165) & (g166)) + ((g1209) & (g1210) & (g1211) & (!g1212) & (!g165) & (!g166)) + ((g1209) & (g1210) & (g1211) & (!g1212) & (!g165) & (g166)) + ((g1209) & (g1210) & (g1211) & (!g1212) & (g165) & (!g166)) + ((g1209) & (g1210) & (g1211) & (g1212) & (!g165) & (!g166)) + ((g1209) & (g1210) & (g1211) & (g1212) & (!g165) & (g166)) + ((g1209) & (g1210) & (g1211) & (g1212) & (g165) & (!g166)) + ((g1209) & (g1210) & (g1211) & (g1212) & (g165) & (g166)));
	assign g4750 = (((!sk[0]) & (!g2177) & (!g3373) & (g1214)) + ((!sk[0]) & (!g2177) & (g3373) & (!g1214)) + ((!sk[0]) & (!g2177) & (g3373) & (g1214)) + ((!sk[0]) & (g2177) & (!g3373) & (g1214)) + ((!sk[0]) & (g2177) & (g3373) & (!g1214)) + ((!sk[0]) & (g2177) & (g3373) & (g1214)) + ((sk[0]) & (!g2177) & (!g3373) & (g1214)) + ((sk[0]) & (!g2177) & (g3373) & (g1214)) + ((sk[0]) & (g2177) & (g3373) & (!g1214)) + ((sk[0]) & (g2177) & (g3373) & (g1214)));
	assign g4751 = (((!g2178) & (!g3373) & (!sk[1]) & (g1215)) + ((!g2178) & (!g3373) & (sk[1]) & (g1215)) + ((!g2178) & (g3373) & (!sk[1]) & (!g1215)) + ((!g2178) & (g3373) & (!sk[1]) & (g1215)) + ((!g2178) & (g3373) & (sk[1]) & (g1215)) + ((g2178) & (!g3373) & (!sk[1]) & (g1215)) + ((g2178) & (g3373) & (!sk[1]) & (!g1215)) + ((g2178) & (g3373) & (!sk[1]) & (g1215)) + ((g2178) & (g3373) & (sk[1]) & (!g1215)) + ((g2178) & (g3373) & (sk[1]) & (g1215)));
	assign g4752 = (((!g2179) & (!g3373) & (!sk[2]) & (g1216)) + ((!g2179) & (!g3373) & (sk[2]) & (g1216)) + ((!g2179) & (g3373) & (!sk[2]) & (!g1216)) + ((!g2179) & (g3373) & (!sk[2]) & (g1216)) + ((!g2179) & (g3373) & (sk[2]) & (g1216)) + ((g2179) & (!g3373) & (!sk[2]) & (g1216)) + ((g2179) & (g3373) & (!sk[2]) & (!g1216)) + ((g2179) & (g3373) & (!sk[2]) & (g1216)) + ((g2179) & (g3373) & (sk[2]) & (!g1216)) + ((g2179) & (g3373) & (sk[2]) & (g1216)));
	assign g1217 = (((!g165) & (!g166) & (!g1214) & (!sk[3]) & (g1215) & (!g1216)) + ((!g165) & (!g166) & (!g1214) & (!sk[3]) & (g1215) & (g1216)) + ((!g165) & (!g166) & (g1214) & (!sk[3]) & (!g1215) & (!g1216)) + ((!g165) & (!g166) & (g1214) & (!sk[3]) & (!g1215) & (g1216)) + ((!g165) & (!g166) & (g1214) & (!sk[3]) & (g1215) & (!g1216)) + ((!g165) & (!g166) & (g1214) & (!sk[3]) & (g1215) & (g1216)) + ((!g165) & (g166) & (!g1214) & (!sk[3]) & (!g1215) & (!g1216)) + ((!g165) & (g166) & (!g1214) & (!sk[3]) & (!g1215) & (g1216)) + ((!g165) & (g166) & (!g1214) & (!sk[3]) & (g1215) & (!g1216)) + ((!g165) & (g166) & (!g1214) & (!sk[3]) & (g1215) & (g1216)) + ((!g165) & (g166) & (!g1214) & (sk[3]) & (!g1215) & (g1216)) + ((!g165) & (g166) & (!g1214) & (sk[3]) & (g1215) & (g1216)) + ((!g165) & (g166) & (g1214) & (!sk[3]) & (!g1215) & (!g1216)) + ((!g165) & (g166) & (g1214) & (!sk[3]) & (!g1215) & (g1216)) + ((!g165) & (g166) & (g1214) & (!sk[3]) & (g1215) & (!g1216)) + ((!g165) & (g166) & (g1214) & (!sk[3]) & (g1215) & (g1216)) + ((!g165) & (g166) & (g1214) & (sk[3]) & (!g1215) & (g1216)) + ((!g165) & (g166) & (g1214) & (sk[3]) & (g1215) & (g1216)) + ((g165) & (!g166) & (!g1214) & (!sk[3]) & (g1215) & (!g1216)) + ((g165) & (!g166) & (!g1214) & (!sk[3]) & (g1215) & (g1216)) + ((g165) & (!g166) & (g1214) & (!sk[3]) & (!g1215) & (!g1216)) + ((g165) & (!g166) & (g1214) & (!sk[3]) & (!g1215) & (g1216)) + ((g165) & (!g166) & (g1214) & (!sk[3]) & (g1215) & (!g1216)) + ((g165) & (!g166) & (g1214) & (!sk[3]) & (g1215) & (g1216)) + ((g165) & (!g166) & (g1214) & (sk[3]) & (!g1215) & (!g1216)) + ((g165) & (!g166) & (g1214) & (sk[3]) & (!g1215) & (g1216)) + ((g165) & (!g166) & (g1214) & (sk[3]) & (g1215) & (!g1216)) + ((g165) & (!g166) & (g1214) & (sk[3]) & (g1215) & (g1216)) + ((g165) & (g166) & (!g1214) & (!sk[3]) & (!g1215) & (!g1216)) + ((g165) & (g166) & (!g1214) & (!sk[3]) & (!g1215) & (g1216)) + ((g165) & (g166) & (!g1214) & (!sk[3]) & (g1215) & (!g1216)) + ((g165) & (g166) & (!g1214) & (!sk[3]) & (g1215) & (g1216)) + ((g165) & (g166) & (!g1214) & (sk[3]) & (g1215) & (!g1216)) + ((g165) & (g166) & (!g1214) & (sk[3]) & (g1215) & (g1216)) + ((g165) & (g166) & (g1214) & (!sk[3]) & (!g1215) & (!g1216)) + ((g165) & (g166) & (g1214) & (!sk[3]) & (!g1215) & (g1216)) + ((g165) & (g166) & (g1214) & (!sk[3]) & (g1215) & (!g1216)) + ((g165) & (g166) & (g1214) & (!sk[3]) & (g1215) & (g1216)) + ((g165) & (g166) & (g1214) & (sk[3]) & (g1215) & (!g1216)) + ((g165) & (g166) & (g1214) & (sk[3]) & (g1215) & (g1216)));
	assign g4753 = (((!g2162) & (!g3373) & (!sk[4]) & (g1218)) + ((!g2162) & (!g3373) & (sk[4]) & (g1218)) + ((!g2162) & (g3373) & (!sk[4]) & (!g1218)) + ((!g2162) & (g3373) & (!sk[4]) & (g1218)) + ((!g2162) & (g3373) & (sk[4]) & (g1218)) + ((g2162) & (!g3373) & (!sk[4]) & (g1218)) + ((g2162) & (g3373) & (!sk[4]) & (!g1218)) + ((g2162) & (g3373) & (!sk[4]) & (g1218)) + ((g2162) & (g3373) & (sk[4]) & (!g1218)) + ((g2162) & (g3373) & (sk[4]) & (g1218)));
	assign g4754 = (((!g2164) & (!g3373) & (!sk[5]) & (g1219)) + ((!g2164) & (!g3373) & (sk[5]) & (g1219)) + ((!g2164) & (g3373) & (!sk[5]) & (!g1219)) + ((!g2164) & (g3373) & (!sk[5]) & (g1219)) + ((!g2164) & (g3373) & (sk[5]) & (g1219)) + ((g2164) & (!g3373) & (!sk[5]) & (g1219)) + ((g2164) & (g3373) & (!sk[5]) & (!g1219)) + ((g2164) & (g3373) & (!sk[5]) & (g1219)) + ((g2164) & (g3373) & (sk[5]) & (!g1219)) + ((g2164) & (g3373) & (sk[5]) & (g1219)));
	assign g4755 = (((!g2166) & (!sk[6]) & (!g3373) & (g1220)) + ((!g2166) & (!sk[6]) & (g3373) & (!g1220)) + ((!g2166) & (!sk[6]) & (g3373) & (g1220)) + ((!g2166) & (sk[6]) & (!g3373) & (g1220)) + ((!g2166) & (sk[6]) & (g3373) & (g1220)) + ((g2166) & (!sk[6]) & (!g3373) & (g1220)) + ((g2166) & (!sk[6]) & (g3373) & (!g1220)) + ((g2166) & (!sk[6]) & (g3373) & (g1220)) + ((g2166) & (sk[6]) & (g3373) & (!g1220)) + ((g2166) & (sk[6]) & (g3373) & (g1220)));
	assign g4756 = (((!g2168) & (!g3373) & (!sk[7]) & (g1221)) + ((!g2168) & (!g3373) & (sk[7]) & (g1221)) + ((!g2168) & (g3373) & (!sk[7]) & (!g1221)) + ((!g2168) & (g3373) & (!sk[7]) & (g1221)) + ((!g2168) & (g3373) & (sk[7]) & (g1221)) + ((g2168) & (!g3373) & (!sk[7]) & (g1221)) + ((g2168) & (g3373) & (!sk[7]) & (!g1221)) + ((g2168) & (g3373) & (!sk[7]) & (g1221)) + ((g2168) & (g3373) & (sk[7]) & (!g1221)) + ((g2168) & (g3373) & (sk[7]) & (g1221)));
	assign g1222 = (((!g1218) & (!g1219) & (!g1220) & (g1221) & (g165) & (g166)) + ((!g1218) & (!g1219) & (g1220) & (!g1221) & (!g165) & (g166)) + ((!g1218) & (!g1219) & (g1220) & (g1221) & (!g165) & (g166)) + ((!g1218) & (!g1219) & (g1220) & (g1221) & (g165) & (g166)) + ((!g1218) & (g1219) & (!g1220) & (!g1221) & (g165) & (!g166)) + ((!g1218) & (g1219) & (!g1220) & (g1221) & (g165) & (!g166)) + ((!g1218) & (g1219) & (!g1220) & (g1221) & (g165) & (g166)) + ((!g1218) & (g1219) & (g1220) & (!g1221) & (!g165) & (g166)) + ((!g1218) & (g1219) & (g1220) & (!g1221) & (g165) & (!g166)) + ((!g1218) & (g1219) & (g1220) & (g1221) & (!g165) & (g166)) + ((!g1218) & (g1219) & (g1220) & (g1221) & (g165) & (!g166)) + ((!g1218) & (g1219) & (g1220) & (g1221) & (g165) & (g166)) + ((g1218) & (!g1219) & (!g1220) & (!g1221) & (!g165) & (!g166)) + ((g1218) & (!g1219) & (!g1220) & (g1221) & (!g165) & (!g166)) + ((g1218) & (!g1219) & (!g1220) & (g1221) & (g165) & (g166)) + ((g1218) & (!g1219) & (g1220) & (!g1221) & (!g165) & (!g166)) + ((g1218) & (!g1219) & (g1220) & (!g1221) & (!g165) & (g166)) + ((g1218) & (!g1219) & (g1220) & (g1221) & (!g165) & (!g166)) + ((g1218) & (!g1219) & (g1220) & (g1221) & (!g165) & (g166)) + ((g1218) & (!g1219) & (g1220) & (g1221) & (g165) & (g166)) + ((g1218) & (g1219) & (!g1220) & (!g1221) & (!g165) & (!g166)) + ((g1218) & (g1219) & (!g1220) & (!g1221) & (g165) & (!g166)) + ((g1218) & (g1219) & (!g1220) & (g1221) & (!g165) & (!g166)) + ((g1218) & (g1219) & (!g1220) & (g1221) & (g165) & (!g166)) + ((g1218) & (g1219) & (!g1220) & (g1221) & (g165) & (g166)) + ((g1218) & (g1219) & (g1220) & (!g1221) & (!g165) & (!g166)) + ((g1218) & (g1219) & (g1220) & (!g1221) & (!g165) & (g166)) + ((g1218) & (g1219) & (g1220) & (!g1221) & (g165) & (!g166)) + ((g1218) & (g1219) & (g1220) & (g1221) & (!g165) & (!g166)) + ((g1218) & (g1219) & (g1220) & (g1221) & (!g165) & (g166)) + ((g1218) & (g1219) & (g1220) & (g1221) & (g165) & (!g166)) + ((g1218) & (g1219) & (g1220) & (g1221) & (g165) & (g166)));
	assign g4757 = (((!g2169) & (!sk[9]) & (!g3373) & (g1223)) + ((!g2169) & (!sk[9]) & (g3373) & (!g1223)) + ((!g2169) & (!sk[9]) & (g3373) & (g1223)) + ((!g2169) & (sk[9]) & (!g3373) & (g1223)) + ((!g2169) & (sk[9]) & (g3373) & (g1223)) + ((g2169) & (!sk[9]) & (!g3373) & (g1223)) + ((g2169) & (!sk[9]) & (g3373) & (!g1223)) + ((g2169) & (!sk[9]) & (g3373) & (g1223)) + ((g2169) & (sk[9]) & (g3373) & (!g1223)) + ((g2169) & (sk[9]) & (g3373) & (g1223)));
	assign g4758 = (((!g2170) & (!g3373) & (!sk[10]) & (g1224)) + ((!g2170) & (!g3373) & (sk[10]) & (g1224)) + ((!g2170) & (g3373) & (!sk[10]) & (!g1224)) + ((!g2170) & (g3373) & (!sk[10]) & (g1224)) + ((!g2170) & (g3373) & (sk[10]) & (g1224)) + ((g2170) & (!g3373) & (!sk[10]) & (g1224)) + ((g2170) & (g3373) & (!sk[10]) & (!g1224)) + ((g2170) & (g3373) & (!sk[10]) & (g1224)) + ((g2170) & (g3373) & (sk[10]) & (!g1224)) + ((g2170) & (g3373) & (sk[10]) & (g1224)));
	assign g4759 = (((!sk[11]) & (!g2171) & (!g3373) & (g1225)) + ((!sk[11]) & (!g2171) & (g3373) & (!g1225)) + ((!sk[11]) & (!g2171) & (g3373) & (g1225)) + ((!sk[11]) & (g2171) & (!g3373) & (g1225)) + ((!sk[11]) & (g2171) & (g3373) & (!g1225)) + ((!sk[11]) & (g2171) & (g3373) & (g1225)) + ((sk[11]) & (!g2171) & (!g3373) & (g1225)) + ((sk[11]) & (!g2171) & (g3373) & (g1225)) + ((sk[11]) & (g2171) & (g3373) & (!g1225)) + ((sk[11]) & (g2171) & (g3373) & (g1225)));
	assign g4760 = (((!g2172) & (!sk[12]) & (!g3373) & (g1226)) + ((!g2172) & (!sk[12]) & (g3373) & (!g1226)) + ((!g2172) & (!sk[12]) & (g3373) & (g1226)) + ((!g2172) & (sk[12]) & (!g3373) & (g1226)) + ((!g2172) & (sk[12]) & (g3373) & (g1226)) + ((g2172) & (!sk[12]) & (!g3373) & (g1226)) + ((g2172) & (!sk[12]) & (g3373) & (!g1226)) + ((g2172) & (!sk[12]) & (g3373) & (g1226)) + ((g2172) & (sk[12]) & (g3373) & (!g1226)) + ((g2172) & (sk[12]) & (g3373) & (g1226)));
	assign g1227 = (((!g1223) & (!g1224) & (!g1225) & (g1226) & (g165) & (g166)) + ((!g1223) & (!g1224) & (g1225) & (!g1226) & (!g165) & (g166)) + ((!g1223) & (!g1224) & (g1225) & (g1226) & (!g165) & (g166)) + ((!g1223) & (!g1224) & (g1225) & (g1226) & (g165) & (g166)) + ((!g1223) & (g1224) & (!g1225) & (!g1226) & (g165) & (!g166)) + ((!g1223) & (g1224) & (!g1225) & (g1226) & (g165) & (!g166)) + ((!g1223) & (g1224) & (!g1225) & (g1226) & (g165) & (g166)) + ((!g1223) & (g1224) & (g1225) & (!g1226) & (!g165) & (g166)) + ((!g1223) & (g1224) & (g1225) & (!g1226) & (g165) & (!g166)) + ((!g1223) & (g1224) & (g1225) & (g1226) & (!g165) & (g166)) + ((!g1223) & (g1224) & (g1225) & (g1226) & (g165) & (!g166)) + ((!g1223) & (g1224) & (g1225) & (g1226) & (g165) & (g166)) + ((g1223) & (!g1224) & (!g1225) & (!g1226) & (!g165) & (!g166)) + ((g1223) & (!g1224) & (!g1225) & (g1226) & (!g165) & (!g166)) + ((g1223) & (!g1224) & (!g1225) & (g1226) & (g165) & (g166)) + ((g1223) & (!g1224) & (g1225) & (!g1226) & (!g165) & (!g166)) + ((g1223) & (!g1224) & (g1225) & (!g1226) & (!g165) & (g166)) + ((g1223) & (!g1224) & (g1225) & (g1226) & (!g165) & (!g166)) + ((g1223) & (!g1224) & (g1225) & (g1226) & (!g165) & (g166)) + ((g1223) & (!g1224) & (g1225) & (g1226) & (g165) & (g166)) + ((g1223) & (g1224) & (!g1225) & (!g1226) & (!g165) & (!g166)) + ((g1223) & (g1224) & (!g1225) & (!g1226) & (g165) & (!g166)) + ((g1223) & (g1224) & (!g1225) & (g1226) & (!g165) & (!g166)) + ((g1223) & (g1224) & (!g1225) & (g1226) & (g165) & (!g166)) + ((g1223) & (g1224) & (!g1225) & (g1226) & (g165) & (g166)) + ((g1223) & (g1224) & (g1225) & (!g1226) & (!g165) & (!g166)) + ((g1223) & (g1224) & (g1225) & (!g1226) & (!g165) & (g166)) + ((g1223) & (g1224) & (g1225) & (!g1226) & (g165) & (!g166)) + ((g1223) & (g1224) & (g1225) & (g1226) & (!g165) & (!g166)) + ((g1223) & (g1224) & (g1225) & (g1226) & (!g165) & (g166)) + ((g1223) & (g1224) & (g1225) & (g1226) & (g165) & (!g166)) + ((g1223) & (g1224) & (g1225) & (g1226) & (g165) & (g166)));
	assign g1228 = (((!g147) & (!g148) & (!g1213) & (g1217) & (!g1222) & (!g1227)) + ((!g147) & (!g148) & (!g1213) & (g1217) & (!g1222) & (g1227)) + ((!g147) & (!g148) & (!g1213) & (g1217) & (g1222) & (!g1227)) + ((!g147) & (!g148) & (!g1213) & (g1217) & (g1222) & (g1227)) + ((!g147) & (!g148) & (g1213) & (g1217) & (!g1222) & (!g1227)) + ((!g147) & (!g148) & (g1213) & (g1217) & (!g1222) & (g1227)) + ((!g147) & (!g148) & (g1213) & (g1217) & (g1222) & (!g1227)) + ((!g147) & (!g148) & (g1213) & (g1217) & (g1222) & (g1227)) + ((!g147) & (g148) & (!g1213) & (!g1217) & (!g1222) & (g1227)) + ((!g147) & (g148) & (!g1213) & (!g1217) & (g1222) & (g1227)) + ((!g147) & (g148) & (!g1213) & (g1217) & (!g1222) & (g1227)) + ((!g147) & (g148) & (!g1213) & (g1217) & (g1222) & (g1227)) + ((!g147) & (g148) & (g1213) & (!g1217) & (!g1222) & (g1227)) + ((!g147) & (g148) & (g1213) & (!g1217) & (g1222) & (g1227)) + ((!g147) & (g148) & (g1213) & (g1217) & (!g1222) & (g1227)) + ((!g147) & (g148) & (g1213) & (g1217) & (g1222) & (g1227)) + ((g147) & (!g148) & (g1213) & (!g1217) & (!g1222) & (!g1227)) + ((g147) & (!g148) & (g1213) & (!g1217) & (!g1222) & (g1227)) + ((g147) & (!g148) & (g1213) & (!g1217) & (g1222) & (!g1227)) + ((g147) & (!g148) & (g1213) & (!g1217) & (g1222) & (g1227)) + ((g147) & (!g148) & (g1213) & (g1217) & (!g1222) & (!g1227)) + ((g147) & (!g148) & (g1213) & (g1217) & (!g1222) & (g1227)) + ((g147) & (!g148) & (g1213) & (g1217) & (g1222) & (!g1227)) + ((g147) & (!g148) & (g1213) & (g1217) & (g1222) & (g1227)) + ((g147) & (g148) & (!g1213) & (!g1217) & (g1222) & (!g1227)) + ((g147) & (g148) & (!g1213) & (!g1217) & (g1222) & (g1227)) + ((g147) & (g148) & (!g1213) & (g1217) & (g1222) & (!g1227)) + ((g147) & (g148) & (!g1213) & (g1217) & (g1222) & (g1227)) + ((g147) & (g148) & (g1213) & (!g1217) & (g1222) & (!g1227)) + ((g147) & (g148) & (g1213) & (!g1217) & (g1222) & (g1227)) + ((g147) & (g148) & (g1213) & (g1217) & (g1222) & (!g1227)) + ((g147) & (g148) & (g1213) & (g1217) & (g1222) & (g1227)));
	assign g1229 = (((!g142) & (!sk[15]) & (!g1208) & (g1228)) + ((!g142) & (!sk[15]) & (g1208) & (!g1228)) + ((!g142) & (!sk[15]) & (g1208) & (g1228)) + ((!g142) & (sk[15]) & (!g1208) & (g1228)) + ((!g142) & (sk[15]) & (g1208) & (g1228)) + ((g142) & (!sk[15]) & (!g1208) & (g1228)) + ((g142) & (!sk[15]) & (g1208) & (!g1228)) + ((g142) & (!sk[15]) & (g1208) & (g1228)) + ((g142) & (sk[15]) & (g1208) & (!g1228)) + ((g142) & (sk[15]) & (g1208) & (g1228)));
	assign g4761 = (((!g2059) & (!sk[16]) & (!g2698) & (g1230)) + ((!g2059) & (!sk[16]) & (g2698) & (!g1230)) + ((!g2059) & (!sk[16]) & (g2698) & (g1230)) + ((!g2059) & (sk[16]) & (!g2698) & (g1230)) + ((!g2059) & (sk[16]) & (g2698) & (g1230)) + ((g2059) & (!sk[16]) & (!g2698) & (g1230)) + ((g2059) & (!sk[16]) & (g2698) & (!g1230)) + ((g2059) & (!sk[16]) & (g2698) & (g1230)) + ((g2059) & (sk[16]) & (g2698) & (!g1230)) + ((g2059) & (sk[16]) & (g2698) & (g1230)));
	assign g1231 = (((!g1139) & (!g1184) & (!g3836) & (!sk[17]) & (g1141) & (!g916)) + ((!g1139) & (!g1184) & (!g3836) & (!sk[17]) & (g1141) & (g916)) + ((!g1139) & (!g1184) & (!g3836) & (sk[17]) & (g1141) & (!g916)) + ((!g1139) & (!g1184) & (g3836) & (!sk[17]) & (!g1141) & (!g916)) + ((!g1139) & (!g1184) & (g3836) & (!sk[17]) & (!g1141) & (g916)) + ((!g1139) & (!g1184) & (g3836) & (!sk[17]) & (g1141) & (!g916)) + ((!g1139) & (!g1184) & (g3836) & (!sk[17]) & (g1141) & (g916)) + ((!g1139) & (!g1184) & (g3836) & (sk[17]) & (!g1141) & (!g916)) + ((!g1139) & (!g1184) & (g3836) & (sk[17]) & (g1141) & (!g916)) + ((!g1139) & (g1184) & (!g3836) & (!sk[17]) & (!g1141) & (!g916)) + ((!g1139) & (g1184) & (!g3836) & (!sk[17]) & (!g1141) & (g916)) + ((!g1139) & (g1184) & (!g3836) & (!sk[17]) & (g1141) & (!g916)) + ((!g1139) & (g1184) & (!g3836) & (!sk[17]) & (g1141) & (g916)) + ((!g1139) & (g1184) & (!g3836) & (sk[17]) & (!g1141) & (!g916)) + ((!g1139) & (g1184) & (!g3836) & (sk[17]) & (g1141) & (!g916)) + ((!g1139) & (g1184) & (g3836) & (!sk[17]) & (!g1141) & (!g916)) + ((!g1139) & (g1184) & (g3836) & (!sk[17]) & (!g1141) & (g916)) + ((!g1139) & (g1184) & (g3836) & (!sk[17]) & (g1141) & (!g916)) + ((!g1139) & (g1184) & (g3836) & (!sk[17]) & (g1141) & (g916)) + ((!g1139) & (g1184) & (g3836) & (sk[17]) & (!g1141) & (!g916)) + ((!g1139) & (g1184) & (g3836) & (sk[17]) & (g1141) & (!g916)) + ((g1139) & (!g1184) & (!g3836) & (!sk[17]) & (g1141) & (!g916)) + ((g1139) & (!g1184) & (!g3836) & (!sk[17]) & (g1141) & (g916)) + ((g1139) & (!g1184) & (!g3836) & (sk[17]) & (!g1141) & (!g916)) + ((g1139) & (!g1184) & (!g3836) & (sk[17]) & (g1141) & (!g916)) + ((g1139) & (!g1184) & (g3836) & (!sk[17]) & (!g1141) & (!g916)) + ((g1139) & (!g1184) & (g3836) & (!sk[17]) & (!g1141) & (g916)) + ((g1139) & (!g1184) & (g3836) & (!sk[17]) & (g1141) & (!g916)) + ((g1139) & (!g1184) & (g3836) & (!sk[17]) & (g1141) & (g916)) + ((g1139) & (!g1184) & (g3836) & (sk[17]) & (!g1141) & (!g916)) + ((g1139) & (!g1184) & (g3836) & (sk[17]) & (g1141) & (!g916)) + ((g1139) & (g1184) & (!g3836) & (!sk[17]) & (!g1141) & (!g916)) + ((g1139) & (g1184) & (!g3836) & (!sk[17]) & (!g1141) & (g916)) + ((g1139) & (g1184) & (!g3836) & (!sk[17]) & (g1141) & (!g916)) + ((g1139) & (g1184) & (!g3836) & (!sk[17]) & (g1141) & (g916)) + ((g1139) & (g1184) & (!g3836) & (sk[17]) & (!g1141) & (!g916)) + ((g1139) & (g1184) & (!g3836) & (sk[17]) & (g1141) & (!g916)) + ((g1139) & (g1184) & (!g3836) & (sk[17]) & (g1141) & (g916)) + ((g1139) & (g1184) & (g3836) & (!sk[17]) & (!g1141) & (!g916)) + ((g1139) & (g1184) & (g3836) & (!sk[17]) & (!g1141) & (g916)) + ((g1139) & (g1184) & (g3836) & (!sk[17]) & (g1141) & (!g916)) + ((g1139) & (g1184) & (g3836) & (!sk[17]) & (g1141) & (g916)) + ((g1139) & (g1184) & (g3836) & (sk[17]) & (!g1141) & (!g916)) + ((g1139) & (g1184) & (g3836) & (sk[17]) & (!g1141) & (g916)) + ((g1139) & (g1184) & (g3836) & (sk[17]) & (g1141) & (!g916)) + ((g1139) & (g1184) & (g3836) & (sk[17]) & (g1141) & (g916)));
	assign g1232 = (((!g126) & (!g1229) & (!g1230) & (g1231) & (!sk[18]) & (!g916)) + ((!g126) & (!g1229) & (!g1230) & (g1231) & (!sk[18]) & (g916)) + ((!g126) & (!g1229) & (g1230) & (!g1231) & (!sk[18]) & (!g916)) + ((!g126) & (!g1229) & (g1230) & (!g1231) & (!sk[18]) & (g916)) + ((!g126) & (!g1229) & (g1230) & (!g1231) & (sk[18]) & (!g916)) + ((!g126) & (!g1229) & (g1230) & (!g1231) & (sk[18]) & (g916)) + ((!g126) & (!g1229) & (g1230) & (g1231) & (!sk[18]) & (!g916)) + ((!g126) & (!g1229) & (g1230) & (g1231) & (!sk[18]) & (g916)) + ((!g126) & (!g1229) & (g1230) & (g1231) & (sk[18]) & (!g916)) + ((!g126) & (!g1229) & (g1230) & (g1231) & (sk[18]) & (g916)) + ((!g126) & (g1229) & (!g1230) & (!g1231) & (!sk[18]) & (!g916)) + ((!g126) & (g1229) & (!g1230) & (!g1231) & (!sk[18]) & (g916)) + ((!g126) & (g1229) & (!g1230) & (g1231) & (!sk[18]) & (!g916)) + ((!g126) & (g1229) & (!g1230) & (g1231) & (!sk[18]) & (g916)) + ((!g126) & (g1229) & (g1230) & (!g1231) & (!sk[18]) & (!g916)) + ((!g126) & (g1229) & (g1230) & (!g1231) & (!sk[18]) & (g916)) + ((!g126) & (g1229) & (g1230) & (!g1231) & (sk[18]) & (!g916)) + ((!g126) & (g1229) & (g1230) & (!g1231) & (sk[18]) & (g916)) + ((!g126) & (g1229) & (g1230) & (g1231) & (!sk[18]) & (!g916)) + ((!g126) & (g1229) & (g1230) & (g1231) & (!sk[18]) & (g916)) + ((!g126) & (g1229) & (g1230) & (g1231) & (sk[18]) & (!g916)) + ((!g126) & (g1229) & (g1230) & (g1231) & (sk[18]) & (g916)) + ((g126) & (!g1229) & (!g1230) & (!g1231) & (sk[18]) & (!g916)) + ((g126) & (!g1229) & (!g1230) & (g1231) & (!sk[18]) & (!g916)) + ((g126) & (!g1229) & (!g1230) & (g1231) & (!sk[18]) & (g916)) + ((g126) & (!g1229) & (!g1230) & (g1231) & (sk[18]) & (g916)) + ((g126) & (!g1229) & (g1230) & (!g1231) & (!sk[18]) & (!g916)) + ((g126) & (!g1229) & (g1230) & (!g1231) & (!sk[18]) & (g916)) + ((g126) & (!g1229) & (g1230) & (!g1231) & (sk[18]) & (!g916)) + ((g126) & (!g1229) & (g1230) & (g1231) & (!sk[18]) & (!g916)) + ((g126) & (!g1229) & (g1230) & (g1231) & (!sk[18]) & (g916)) + ((g126) & (!g1229) & (g1230) & (g1231) & (sk[18]) & (g916)) + ((g126) & (g1229) & (!g1230) & (!g1231) & (!sk[18]) & (!g916)) + ((g126) & (g1229) & (!g1230) & (!g1231) & (!sk[18]) & (g916)) + ((g126) & (g1229) & (!g1230) & (!g1231) & (sk[18]) & (g916)) + ((g126) & (g1229) & (!g1230) & (g1231) & (!sk[18]) & (!g916)) + ((g126) & (g1229) & (!g1230) & (g1231) & (!sk[18]) & (g916)) + ((g126) & (g1229) & (!g1230) & (g1231) & (sk[18]) & (!g916)) + ((g126) & (g1229) & (g1230) & (!g1231) & (!sk[18]) & (!g916)) + ((g126) & (g1229) & (g1230) & (!g1231) & (!sk[18]) & (g916)) + ((g126) & (g1229) & (g1230) & (!g1231) & (sk[18]) & (g916)) + ((g126) & (g1229) & (g1230) & (g1231) & (!sk[18]) & (!g916)) + ((g126) & (g1229) & (g1230) & (g1231) & (!sk[18]) & (g916)) + ((g126) & (g1229) & (g1230) & (g1231) & (sk[18]) & (!g916)));
	assign g4762 = (((!sk[19]) & (!g2140) & (!g3349) & (g1233)) + ((!sk[19]) & (!g2140) & (g3349) & (!g1233)) + ((!sk[19]) & (!g2140) & (g3349) & (g1233)) + ((!sk[19]) & (g2140) & (!g3349) & (g1233)) + ((!sk[19]) & (g2140) & (g3349) & (!g1233)) + ((!sk[19]) & (g2140) & (g3349) & (g1233)) + ((sk[19]) & (!g2140) & (!g3349) & (g1233)) + ((sk[19]) & (!g2140) & (g3349) & (g1233)) + ((sk[19]) & (g2140) & (g3349) & (!g1233)) + ((sk[19]) & (g2140) & (g3349) & (g1233)));
	assign g4763 = (((!g2142) & (!sk[20]) & (!g3349) & (g1234)) + ((!g2142) & (!sk[20]) & (g3349) & (!g1234)) + ((!g2142) & (!sk[20]) & (g3349) & (g1234)) + ((!g2142) & (sk[20]) & (!g3349) & (g1234)) + ((!g2142) & (sk[20]) & (g3349) & (g1234)) + ((g2142) & (!sk[20]) & (!g3349) & (g1234)) + ((g2142) & (!sk[20]) & (g3349) & (!g1234)) + ((g2142) & (!sk[20]) & (g3349) & (g1234)) + ((g2142) & (sk[20]) & (g3349) & (!g1234)) + ((g2142) & (sk[20]) & (g3349) & (g1234)));
	assign g4764 = (((!g2144) & (!sk[21]) & (!g3349) & (g1235)) + ((!g2144) & (!sk[21]) & (g3349) & (!g1235)) + ((!g2144) & (!sk[21]) & (g3349) & (g1235)) + ((!g2144) & (sk[21]) & (!g3349) & (g1235)) + ((!g2144) & (sk[21]) & (g3349) & (g1235)) + ((g2144) & (!sk[21]) & (!g3349) & (g1235)) + ((g2144) & (!sk[21]) & (g3349) & (!g1235)) + ((g2144) & (!sk[21]) & (g3349) & (g1235)) + ((g2144) & (sk[21]) & (g3349) & (!g1235)) + ((g2144) & (sk[21]) & (g3349) & (g1235)));
	assign g4765 = (((!g2145) & (!g3349) & (!sk[22]) & (g1236)) + ((!g2145) & (!g3349) & (sk[22]) & (g1236)) + ((!g2145) & (g3349) & (!sk[22]) & (!g1236)) + ((!g2145) & (g3349) & (!sk[22]) & (g1236)) + ((!g2145) & (g3349) & (sk[22]) & (g1236)) + ((g2145) & (!g3349) & (!sk[22]) & (g1236)) + ((g2145) & (g3349) & (!sk[22]) & (!g1236)) + ((g2145) & (g3349) & (!sk[22]) & (g1236)) + ((g2145) & (g3349) & (sk[22]) & (!g1236)) + ((g2145) & (g3349) & (sk[22]) & (g1236)));
	assign g1237 = (((!g1233) & (!g1234) & (!g1235) & (g1236) & (g147) & (g148)) + ((!g1233) & (!g1234) & (g1235) & (!g1236) & (!g147) & (g148)) + ((!g1233) & (!g1234) & (g1235) & (g1236) & (!g147) & (g148)) + ((!g1233) & (!g1234) & (g1235) & (g1236) & (g147) & (g148)) + ((!g1233) & (g1234) & (!g1235) & (!g1236) & (g147) & (!g148)) + ((!g1233) & (g1234) & (!g1235) & (g1236) & (g147) & (!g148)) + ((!g1233) & (g1234) & (!g1235) & (g1236) & (g147) & (g148)) + ((!g1233) & (g1234) & (g1235) & (!g1236) & (!g147) & (g148)) + ((!g1233) & (g1234) & (g1235) & (!g1236) & (g147) & (!g148)) + ((!g1233) & (g1234) & (g1235) & (g1236) & (!g147) & (g148)) + ((!g1233) & (g1234) & (g1235) & (g1236) & (g147) & (!g148)) + ((!g1233) & (g1234) & (g1235) & (g1236) & (g147) & (g148)) + ((g1233) & (!g1234) & (!g1235) & (!g1236) & (!g147) & (!g148)) + ((g1233) & (!g1234) & (!g1235) & (g1236) & (!g147) & (!g148)) + ((g1233) & (!g1234) & (!g1235) & (g1236) & (g147) & (g148)) + ((g1233) & (!g1234) & (g1235) & (!g1236) & (!g147) & (!g148)) + ((g1233) & (!g1234) & (g1235) & (!g1236) & (!g147) & (g148)) + ((g1233) & (!g1234) & (g1235) & (g1236) & (!g147) & (!g148)) + ((g1233) & (!g1234) & (g1235) & (g1236) & (!g147) & (g148)) + ((g1233) & (!g1234) & (g1235) & (g1236) & (g147) & (g148)) + ((g1233) & (g1234) & (!g1235) & (!g1236) & (!g147) & (!g148)) + ((g1233) & (g1234) & (!g1235) & (!g1236) & (g147) & (!g148)) + ((g1233) & (g1234) & (!g1235) & (g1236) & (!g147) & (!g148)) + ((g1233) & (g1234) & (!g1235) & (g1236) & (g147) & (!g148)) + ((g1233) & (g1234) & (!g1235) & (g1236) & (g147) & (g148)) + ((g1233) & (g1234) & (g1235) & (!g1236) & (!g147) & (!g148)) + ((g1233) & (g1234) & (g1235) & (!g1236) & (!g147) & (g148)) + ((g1233) & (g1234) & (g1235) & (!g1236) & (g147) & (!g148)) + ((g1233) & (g1234) & (g1235) & (g1236) & (!g147) & (!g148)) + ((g1233) & (g1234) & (g1235) & (g1236) & (!g147) & (g148)) + ((g1233) & (g1234) & (g1235) & (g1236) & (g147) & (!g148)) + ((g1233) & (g1234) & (g1235) & (g1236) & (g147) & (g148)));
	assign g4766 = (((!g2146) & (!sk[24]) & (!g3349) & (g1238)) + ((!g2146) & (!sk[24]) & (g3349) & (!g1238)) + ((!g2146) & (!sk[24]) & (g3349) & (g1238)) + ((!g2146) & (sk[24]) & (!g3349) & (g1238)) + ((!g2146) & (sk[24]) & (g3349) & (g1238)) + ((g2146) & (!sk[24]) & (!g3349) & (g1238)) + ((g2146) & (!sk[24]) & (g3349) & (!g1238)) + ((g2146) & (!sk[24]) & (g3349) & (g1238)) + ((g2146) & (sk[24]) & (g3349) & (!g1238)) + ((g2146) & (sk[24]) & (g3349) & (g1238)));
	assign g4767 = (((!g2148) & (!g3349) & (!sk[25]) & (g1239)) + ((!g2148) & (!g3349) & (sk[25]) & (g1239)) + ((!g2148) & (g3349) & (!sk[25]) & (!g1239)) + ((!g2148) & (g3349) & (!sk[25]) & (g1239)) + ((!g2148) & (g3349) & (sk[25]) & (g1239)) + ((g2148) & (!g3349) & (!sk[25]) & (g1239)) + ((g2148) & (g3349) & (!sk[25]) & (!g1239)) + ((g2148) & (g3349) & (!sk[25]) & (g1239)) + ((g2148) & (g3349) & (sk[25]) & (!g1239)) + ((g2148) & (g3349) & (sk[25]) & (g1239)));
	assign g4768 = (((!g2150) & (!g3349) & (!sk[26]) & (g1240)) + ((!g2150) & (!g3349) & (sk[26]) & (g1240)) + ((!g2150) & (g3349) & (!sk[26]) & (!g1240)) + ((!g2150) & (g3349) & (!sk[26]) & (g1240)) + ((!g2150) & (g3349) & (sk[26]) & (g1240)) + ((g2150) & (!g3349) & (!sk[26]) & (g1240)) + ((g2150) & (g3349) & (!sk[26]) & (!g1240)) + ((g2150) & (g3349) & (!sk[26]) & (g1240)) + ((g2150) & (g3349) & (sk[26]) & (!g1240)) + ((g2150) & (g3349) & (sk[26]) & (g1240)));
	assign g4769 = (((!g2151) & (!sk[27]) & (!g3349) & (g1241)) + ((!g2151) & (!sk[27]) & (g3349) & (!g1241)) + ((!g2151) & (!sk[27]) & (g3349) & (g1241)) + ((!g2151) & (sk[27]) & (!g3349) & (g1241)) + ((!g2151) & (sk[27]) & (g3349) & (g1241)) + ((g2151) & (!sk[27]) & (!g3349) & (g1241)) + ((g2151) & (!sk[27]) & (g3349) & (!g1241)) + ((g2151) & (!sk[27]) & (g3349) & (g1241)) + ((g2151) & (sk[27]) & (g3349) & (!g1241)) + ((g2151) & (sk[27]) & (g3349) & (g1241)));
	assign g1242 = (((!g1238) & (!g1239) & (!g1240) & (g1241) & (g147) & (g148)) + ((!g1238) & (!g1239) & (g1240) & (!g1241) & (!g147) & (g148)) + ((!g1238) & (!g1239) & (g1240) & (g1241) & (!g147) & (g148)) + ((!g1238) & (!g1239) & (g1240) & (g1241) & (g147) & (g148)) + ((!g1238) & (g1239) & (!g1240) & (!g1241) & (g147) & (!g148)) + ((!g1238) & (g1239) & (!g1240) & (g1241) & (g147) & (!g148)) + ((!g1238) & (g1239) & (!g1240) & (g1241) & (g147) & (g148)) + ((!g1238) & (g1239) & (g1240) & (!g1241) & (!g147) & (g148)) + ((!g1238) & (g1239) & (g1240) & (!g1241) & (g147) & (!g148)) + ((!g1238) & (g1239) & (g1240) & (g1241) & (!g147) & (g148)) + ((!g1238) & (g1239) & (g1240) & (g1241) & (g147) & (!g148)) + ((!g1238) & (g1239) & (g1240) & (g1241) & (g147) & (g148)) + ((g1238) & (!g1239) & (!g1240) & (!g1241) & (!g147) & (!g148)) + ((g1238) & (!g1239) & (!g1240) & (g1241) & (!g147) & (!g148)) + ((g1238) & (!g1239) & (!g1240) & (g1241) & (g147) & (g148)) + ((g1238) & (!g1239) & (g1240) & (!g1241) & (!g147) & (!g148)) + ((g1238) & (!g1239) & (g1240) & (!g1241) & (!g147) & (g148)) + ((g1238) & (!g1239) & (g1240) & (g1241) & (!g147) & (!g148)) + ((g1238) & (!g1239) & (g1240) & (g1241) & (!g147) & (g148)) + ((g1238) & (!g1239) & (g1240) & (g1241) & (g147) & (g148)) + ((g1238) & (g1239) & (!g1240) & (!g1241) & (!g147) & (!g148)) + ((g1238) & (g1239) & (!g1240) & (!g1241) & (g147) & (!g148)) + ((g1238) & (g1239) & (!g1240) & (g1241) & (!g147) & (!g148)) + ((g1238) & (g1239) & (!g1240) & (g1241) & (g147) & (!g148)) + ((g1238) & (g1239) & (!g1240) & (g1241) & (g147) & (g148)) + ((g1238) & (g1239) & (g1240) & (!g1241) & (!g147) & (!g148)) + ((g1238) & (g1239) & (g1240) & (!g1241) & (!g147) & (g148)) + ((g1238) & (g1239) & (g1240) & (!g1241) & (g147) & (!g148)) + ((g1238) & (g1239) & (g1240) & (g1241) & (!g147) & (!g148)) + ((g1238) & (g1239) & (g1240) & (g1241) & (!g147) & (g148)) + ((g1238) & (g1239) & (g1240) & (g1241) & (g147) & (!g148)) + ((g1238) & (g1239) & (g1240) & (g1241) & (g147) & (g148)));
	assign g4770 = (((!g2152) & (!g3349) & (!sk[29]) & (g1243)) + ((!g2152) & (!g3349) & (sk[29]) & (g1243)) + ((!g2152) & (g3349) & (!sk[29]) & (!g1243)) + ((!g2152) & (g3349) & (!sk[29]) & (g1243)) + ((!g2152) & (g3349) & (sk[29]) & (g1243)) + ((g2152) & (!g3349) & (!sk[29]) & (g1243)) + ((g2152) & (g3349) & (!sk[29]) & (!g1243)) + ((g2152) & (g3349) & (!sk[29]) & (g1243)) + ((g2152) & (g3349) & (sk[29]) & (!g1243)) + ((g2152) & (g3349) & (sk[29]) & (g1243)));
	assign g4771 = (((!g2153) & (!sk[30]) & (!g3349) & (g1244)) + ((!g2153) & (!sk[30]) & (g3349) & (!g1244)) + ((!g2153) & (!sk[30]) & (g3349) & (g1244)) + ((!g2153) & (sk[30]) & (!g3349) & (g1244)) + ((!g2153) & (sk[30]) & (g3349) & (g1244)) + ((g2153) & (!sk[30]) & (!g3349) & (g1244)) + ((g2153) & (!sk[30]) & (g3349) & (!g1244)) + ((g2153) & (!sk[30]) & (g3349) & (g1244)) + ((g2153) & (sk[30]) & (g3349) & (!g1244)) + ((g2153) & (sk[30]) & (g3349) & (g1244)));
	assign g4772 = (((!g2155) & (!g3349) & (!sk[31]) & (g1245)) + ((!g2155) & (!g3349) & (sk[31]) & (g1245)) + ((!g2155) & (g3349) & (!sk[31]) & (!g1245)) + ((!g2155) & (g3349) & (!sk[31]) & (g1245)) + ((!g2155) & (g3349) & (sk[31]) & (g1245)) + ((g2155) & (!g3349) & (!sk[31]) & (g1245)) + ((g2155) & (g3349) & (!sk[31]) & (!g1245)) + ((g2155) & (g3349) & (!sk[31]) & (g1245)) + ((g2155) & (g3349) & (sk[31]) & (!g1245)) + ((g2155) & (g3349) & (sk[31]) & (g1245)));
	assign g4773 = (((!g2157) & (!sk[32]) & (!g3349) & (g1246)) + ((!g2157) & (!sk[32]) & (g3349) & (!g1246)) + ((!g2157) & (!sk[32]) & (g3349) & (g1246)) + ((!g2157) & (sk[32]) & (!g3349) & (g1246)) + ((!g2157) & (sk[32]) & (g3349) & (g1246)) + ((g2157) & (!sk[32]) & (!g3349) & (g1246)) + ((g2157) & (!sk[32]) & (g3349) & (!g1246)) + ((g2157) & (!sk[32]) & (g3349) & (g1246)) + ((g2157) & (sk[32]) & (g3349) & (!g1246)) + ((g2157) & (sk[32]) & (g3349) & (g1246)));
	assign g1247 = (((!g1243) & (!g1244) & (!g1245) & (g1246) & (g147) & (g148)) + ((!g1243) & (!g1244) & (g1245) & (!g1246) & (!g147) & (g148)) + ((!g1243) & (!g1244) & (g1245) & (g1246) & (!g147) & (g148)) + ((!g1243) & (!g1244) & (g1245) & (g1246) & (g147) & (g148)) + ((!g1243) & (g1244) & (!g1245) & (!g1246) & (g147) & (!g148)) + ((!g1243) & (g1244) & (!g1245) & (g1246) & (g147) & (!g148)) + ((!g1243) & (g1244) & (!g1245) & (g1246) & (g147) & (g148)) + ((!g1243) & (g1244) & (g1245) & (!g1246) & (!g147) & (g148)) + ((!g1243) & (g1244) & (g1245) & (!g1246) & (g147) & (!g148)) + ((!g1243) & (g1244) & (g1245) & (g1246) & (!g147) & (g148)) + ((!g1243) & (g1244) & (g1245) & (g1246) & (g147) & (!g148)) + ((!g1243) & (g1244) & (g1245) & (g1246) & (g147) & (g148)) + ((g1243) & (!g1244) & (!g1245) & (!g1246) & (!g147) & (!g148)) + ((g1243) & (!g1244) & (!g1245) & (g1246) & (!g147) & (!g148)) + ((g1243) & (!g1244) & (!g1245) & (g1246) & (g147) & (g148)) + ((g1243) & (!g1244) & (g1245) & (!g1246) & (!g147) & (!g148)) + ((g1243) & (!g1244) & (g1245) & (!g1246) & (!g147) & (g148)) + ((g1243) & (!g1244) & (g1245) & (g1246) & (!g147) & (!g148)) + ((g1243) & (!g1244) & (g1245) & (g1246) & (!g147) & (g148)) + ((g1243) & (!g1244) & (g1245) & (g1246) & (g147) & (g148)) + ((g1243) & (g1244) & (!g1245) & (!g1246) & (!g147) & (!g148)) + ((g1243) & (g1244) & (!g1245) & (!g1246) & (g147) & (!g148)) + ((g1243) & (g1244) & (!g1245) & (g1246) & (!g147) & (!g148)) + ((g1243) & (g1244) & (!g1245) & (g1246) & (g147) & (!g148)) + ((g1243) & (g1244) & (!g1245) & (g1246) & (g147) & (g148)) + ((g1243) & (g1244) & (g1245) & (!g1246) & (!g147) & (!g148)) + ((g1243) & (g1244) & (g1245) & (!g1246) & (!g147) & (g148)) + ((g1243) & (g1244) & (g1245) & (!g1246) & (g147) & (!g148)) + ((g1243) & (g1244) & (g1245) & (g1246) & (!g147) & (!g148)) + ((g1243) & (g1244) & (g1245) & (g1246) & (!g147) & (g148)) + ((g1243) & (g1244) & (g1245) & (g1246) & (g147) & (!g148)) + ((g1243) & (g1244) & (g1245) & (g1246) & (g147) & (g148)));
	assign g4774 = (((!g2158) & (!g3349) & (!sk[34]) & (g1248)) + ((!g2158) & (!g3349) & (sk[34]) & (g1248)) + ((!g2158) & (g3349) & (!sk[34]) & (!g1248)) + ((!g2158) & (g3349) & (!sk[34]) & (g1248)) + ((!g2158) & (g3349) & (sk[34]) & (g1248)) + ((g2158) & (!g3349) & (!sk[34]) & (g1248)) + ((g2158) & (g3349) & (!sk[34]) & (!g1248)) + ((g2158) & (g3349) & (!sk[34]) & (g1248)) + ((g2158) & (g3349) & (sk[34]) & (!g1248)) + ((g2158) & (g3349) & (sk[34]) & (g1248)));
	assign g4775 = (((!g2159) & (!sk[35]) & (!g3349) & (g1249)) + ((!g2159) & (!sk[35]) & (g3349) & (!g1249)) + ((!g2159) & (!sk[35]) & (g3349) & (g1249)) + ((!g2159) & (sk[35]) & (!g3349) & (g1249)) + ((!g2159) & (sk[35]) & (g3349) & (g1249)) + ((g2159) & (!sk[35]) & (!g3349) & (g1249)) + ((g2159) & (!sk[35]) & (g3349) & (!g1249)) + ((g2159) & (!sk[35]) & (g3349) & (g1249)) + ((g2159) & (sk[35]) & (g3349) & (!g1249)) + ((g2159) & (sk[35]) & (g3349) & (g1249)));
	assign g4776 = (((!g2160) & (!g3349) & (!sk[36]) & (g1250)) + ((!g2160) & (!g3349) & (sk[36]) & (g1250)) + ((!g2160) & (g3349) & (!sk[36]) & (!g1250)) + ((!g2160) & (g3349) & (!sk[36]) & (g1250)) + ((!g2160) & (g3349) & (sk[36]) & (g1250)) + ((g2160) & (!g3349) & (!sk[36]) & (g1250)) + ((g2160) & (g3349) & (!sk[36]) & (!g1250)) + ((g2160) & (g3349) & (!sk[36]) & (g1250)) + ((g2160) & (g3349) & (sk[36]) & (!g1250)) + ((g2160) & (g3349) & (sk[36]) & (g1250)));
	assign g4777 = (((!g2161) & (!sk[37]) & (!g3349) & (g1251)) + ((!g2161) & (!sk[37]) & (g3349) & (!g1251)) + ((!g2161) & (!sk[37]) & (g3349) & (g1251)) + ((!g2161) & (sk[37]) & (!g3349) & (g1251)) + ((!g2161) & (sk[37]) & (g3349) & (g1251)) + ((g2161) & (!sk[37]) & (!g3349) & (g1251)) + ((g2161) & (!sk[37]) & (g3349) & (!g1251)) + ((g2161) & (!sk[37]) & (g3349) & (g1251)) + ((g2161) & (sk[37]) & (g3349) & (!g1251)) + ((g2161) & (sk[37]) & (g3349) & (g1251)));
	assign g1252 = (((!g1248) & (!g1249) & (!g1250) & (g1251) & (g147) & (g148)) + ((!g1248) & (!g1249) & (g1250) & (!g1251) & (!g147) & (g148)) + ((!g1248) & (!g1249) & (g1250) & (g1251) & (!g147) & (g148)) + ((!g1248) & (!g1249) & (g1250) & (g1251) & (g147) & (g148)) + ((!g1248) & (g1249) & (!g1250) & (!g1251) & (g147) & (!g148)) + ((!g1248) & (g1249) & (!g1250) & (g1251) & (g147) & (!g148)) + ((!g1248) & (g1249) & (!g1250) & (g1251) & (g147) & (g148)) + ((!g1248) & (g1249) & (g1250) & (!g1251) & (!g147) & (g148)) + ((!g1248) & (g1249) & (g1250) & (!g1251) & (g147) & (!g148)) + ((!g1248) & (g1249) & (g1250) & (g1251) & (!g147) & (g148)) + ((!g1248) & (g1249) & (g1250) & (g1251) & (g147) & (!g148)) + ((!g1248) & (g1249) & (g1250) & (g1251) & (g147) & (g148)) + ((g1248) & (!g1249) & (!g1250) & (!g1251) & (!g147) & (!g148)) + ((g1248) & (!g1249) & (!g1250) & (g1251) & (!g147) & (!g148)) + ((g1248) & (!g1249) & (!g1250) & (g1251) & (g147) & (g148)) + ((g1248) & (!g1249) & (g1250) & (!g1251) & (!g147) & (!g148)) + ((g1248) & (!g1249) & (g1250) & (!g1251) & (!g147) & (g148)) + ((g1248) & (!g1249) & (g1250) & (g1251) & (!g147) & (!g148)) + ((g1248) & (!g1249) & (g1250) & (g1251) & (!g147) & (g148)) + ((g1248) & (!g1249) & (g1250) & (g1251) & (g147) & (g148)) + ((g1248) & (g1249) & (!g1250) & (!g1251) & (!g147) & (!g148)) + ((g1248) & (g1249) & (!g1250) & (!g1251) & (g147) & (!g148)) + ((g1248) & (g1249) & (!g1250) & (g1251) & (!g147) & (!g148)) + ((g1248) & (g1249) & (!g1250) & (g1251) & (g147) & (!g148)) + ((g1248) & (g1249) & (!g1250) & (g1251) & (g147) & (g148)) + ((g1248) & (g1249) & (g1250) & (!g1251) & (!g147) & (!g148)) + ((g1248) & (g1249) & (g1250) & (!g1251) & (!g147) & (g148)) + ((g1248) & (g1249) & (g1250) & (!g1251) & (g147) & (!g148)) + ((g1248) & (g1249) & (g1250) & (g1251) & (!g147) & (!g148)) + ((g1248) & (g1249) & (g1250) & (g1251) & (!g147) & (g148)) + ((g1248) & (g1249) & (g1250) & (g1251) & (g147) & (!g148)) + ((g1248) & (g1249) & (g1250) & (g1251) & (g147) & (g148)));
	assign g1253 = (((!g1237) & (!g1242) & (!g1247) & (g1252) & (g165) & (g166)) + ((!g1237) & (!g1242) & (g1247) & (!g1252) & (!g165) & (g166)) + ((!g1237) & (!g1242) & (g1247) & (g1252) & (!g165) & (g166)) + ((!g1237) & (!g1242) & (g1247) & (g1252) & (g165) & (g166)) + ((!g1237) & (g1242) & (!g1247) & (!g1252) & (g165) & (!g166)) + ((!g1237) & (g1242) & (!g1247) & (g1252) & (g165) & (!g166)) + ((!g1237) & (g1242) & (!g1247) & (g1252) & (g165) & (g166)) + ((!g1237) & (g1242) & (g1247) & (!g1252) & (!g165) & (g166)) + ((!g1237) & (g1242) & (g1247) & (!g1252) & (g165) & (!g166)) + ((!g1237) & (g1242) & (g1247) & (g1252) & (!g165) & (g166)) + ((!g1237) & (g1242) & (g1247) & (g1252) & (g165) & (!g166)) + ((!g1237) & (g1242) & (g1247) & (g1252) & (g165) & (g166)) + ((g1237) & (!g1242) & (!g1247) & (!g1252) & (!g165) & (!g166)) + ((g1237) & (!g1242) & (!g1247) & (g1252) & (!g165) & (!g166)) + ((g1237) & (!g1242) & (!g1247) & (g1252) & (g165) & (g166)) + ((g1237) & (!g1242) & (g1247) & (!g1252) & (!g165) & (!g166)) + ((g1237) & (!g1242) & (g1247) & (!g1252) & (!g165) & (g166)) + ((g1237) & (!g1242) & (g1247) & (g1252) & (!g165) & (!g166)) + ((g1237) & (!g1242) & (g1247) & (g1252) & (!g165) & (g166)) + ((g1237) & (!g1242) & (g1247) & (g1252) & (g165) & (g166)) + ((g1237) & (g1242) & (!g1247) & (!g1252) & (!g165) & (!g166)) + ((g1237) & (g1242) & (!g1247) & (!g1252) & (g165) & (!g166)) + ((g1237) & (g1242) & (!g1247) & (g1252) & (!g165) & (!g166)) + ((g1237) & (g1242) & (!g1247) & (g1252) & (g165) & (!g166)) + ((g1237) & (g1242) & (!g1247) & (g1252) & (g165) & (g166)) + ((g1237) & (g1242) & (g1247) & (!g1252) & (!g165) & (!g166)) + ((g1237) & (g1242) & (g1247) & (!g1252) & (!g165) & (g166)) + ((g1237) & (g1242) & (g1247) & (!g1252) & (g165) & (!g166)) + ((g1237) & (g1242) & (g1247) & (g1252) & (!g165) & (!g166)) + ((g1237) & (g1242) & (g1247) & (g1252) & (!g165) & (g166)) + ((g1237) & (g1242) & (g1247) & (g1252) & (g165) & (!g166)) + ((g1237) & (g1242) & (g1247) & (g1252) & (g165) & (g166)));
	assign g4778 = (((!g2173) & (!sk[40]) & (!g3349) & (g1254)) + ((!g2173) & (!sk[40]) & (g3349) & (!g1254)) + ((!g2173) & (!sk[40]) & (g3349) & (g1254)) + ((!g2173) & (sk[40]) & (!g3349) & (g1254)) + ((!g2173) & (sk[40]) & (g3349) & (g1254)) + ((g2173) & (!sk[40]) & (!g3349) & (g1254)) + ((g2173) & (!sk[40]) & (g3349) & (!g1254)) + ((g2173) & (!sk[40]) & (g3349) & (g1254)) + ((g2173) & (sk[40]) & (g3349) & (!g1254)) + ((g2173) & (sk[40]) & (g3349) & (g1254)));
	assign g4779 = (((!g2174) & (!sk[41]) & (!g3349) & (g1255)) + ((!g2174) & (!sk[41]) & (g3349) & (!g1255)) + ((!g2174) & (!sk[41]) & (g3349) & (g1255)) + ((!g2174) & (sk[41]) & (!g3349) & (g1255)) + ((!g2174) & (sk[41]) & (g3349) & (g1255)) + ((g2174) & (!sk[41]) & (!g3349) & (g1255)) + ((g2174) & (!sk[41]) & (g3349) & (!g1255)) + ((g2174) & (!sk[41]) & (g3349) & (g1255)) + ((g2174) & (sk[41]) & (g3349) & (!g1255)) + ((g2174) & (sk[41]) & (g3349) & (g1255)));
	assign g4780 = (((!sk[42]) & (!g2175) & (!g3349) & (g1256)) + ((!sk[42]) & (!g2175) & (g3349) & (!g1256)) + ((!sk[42]) & (!g2175) & (g3349) & (g1256)) + ((!sk[42]) & (g2175) & (!g3349) & (g1256)) + ((!sk[42]) & (g2175) & (g3349) & (!g1256)) + ((!sk[42]) & (g2175) & (g3349) & (g1256)) + ((sk[42]) & (!g2175) & (!g3349) & (g1256)) + ((sk[42]) & (!g2175) & (g3349) & (g1256)) + ((sk[42]) & (g2175) & (g3349) & (!g1256)) + ((sk[42]) & (g2175) & (g3349) & (g1256)));
	assign g4781 = (((!g2176) & (!g3349) & (!sk[43]) & (g1257)) + ((!g2176) & (!g3349) & (sk[43]) & (g1257)) + ((!g2176) & (g3349) & (!sk[43]) & (!g1257)) + ((!g2176) & (g3349) & (!sk[43]) & (g1257)) + ((!g2176) & (g3349) & (sk[43]) & (g1257)) + ((g2176) & (!g3349) & (!sk[43]) & (g1257)) + ((g2176) & (g3349) & (!sk[43]) & (!g1257)) + ((g2176) & (g3349) & (!sk[43]) & (g1257)) + ((g2176) & (g3349) & (sk[43]) & (!g1257)) + ((g2176) & (g3349) & (sk[43]) & (g1257)));
	assign g1258 = (((!g1254) & (!g1255) & (!g1256) & (g1257) & (g165) & (g166)) + ((!g1254) & (!g1255) & (g1256) & (!g1257) & (!g165) & (g166)) + ((!g1254) & (!g1255) & (g1256) & (g1257) & (!g165) & (g166)) + ((!g1254) & (!g1255) & (g1256) & (g1257) & (g165) & (g166)) + ((!g1254) & (g1255) & (!g1256) & (!g1257) & (g165) & (!g166)) + ((!g1254) & (g1255) & (!g1256) & (g1257) & (g165) & (!g166)) + ((!g1254) & (g1255) & (!g1256) & (g1257) & (g165) & (g166)) + ((!g1254) & (g1255) & (g1256) & (!g1257) & (!g165) & (g166)) + ((!g1254) & (g1255) & (g1256) & (!g1257) & (g165) & (!g166)) + ((!g1254) & (g1255) & (g1256) & (g1257) & (!g165) & (g166)) + ((!g1254) & (g1255) & (g1256) & (g1257) & (g165) & (!g166)) + ((!g1254) & (g1255) & (g1256) & (g1257) & (g165) & (g166)) + ((g1254) & (!g1255) & (!g1256) & (!g1257) & (!g165) & (!g166)) + ((g1254) & (!g1255) & (!g1256) & (g1257) & (!g165) & (!g166)) + ((g1254) & (!g1255) & (!g1256) & (g1257) & (g165) & (g166)) + ((g1254) & (!g1255) & (g1256) & (!g1257) & (!g165) & (!g166)) + ((g1254) & (!g1255) & (g1256) & (!g1257) & (!g165) & (g166)) + ((g1254) & (!g1255) & (g1256) & (g1257) & (!g165) & (!g166)) + ((g1254) & (!g1255) & (g1256) & (g1257) & (!g165) & (g166)) + ((g1254) & (!g1255) & (g1256) & (g1257) & (g165) & (g166)) + ((g1254) & (g1255) & (!g1256) & (!g1257) & (!g165) & (!g166)) + ((g1254) & (g1255) & (!g1256) & (!g1257) & (g165) & (!g166)) + ((g1254) & (g1255) & (!g1256) & (g1257) & (!g165) & (!g166)) + ((g1254) & (g1255) & (!g1256) & (g1257) & (g165) & (!g166)) + ((g1254) & (g1255) & (!g1256) & (g1257) & (g165) & (g166)) + ((g1254) & (g1255) & (g1256) & (!g1257) & (!g165) & (!g166)) + ((g1254) & (g1255) & (g1256) & (!g1257) & (!g165) & (g166)) + ((g1254) & (g1255) & (g1256) & (!g1257) & (g165) & (!g166)) + ((g1254) & (g1255) & (g1256) & (g1257) & (!g165) & (!g166)) + ((g1254) & (g1255) & (g1256) & (g1257) & (!g165) & (g166)) + ((g1254) & (g1255) & (g1256) & (g1257) & (g165) & (!g166)) + ((g1254) & (g1255) & (g1256) & (g1257) & (g165) & (g166)));
	assign g4782 = (((!g2177) & (!g3349) & (!sk[45]) & (g1259)) + ((!g2177) & (!g3349) & (sk[45]) & (g1259)) + ((!g2177) & (g3349) & (!sk[45]) & (!g1259)) + ((!g2177) & (g3349) & (!sk[45]) & (g1259)) + ((!g2177) & (g3349) & (sk[45]) & (g1259)) + ((g2177) & (!g3349) & (!sk[45]) & (g1259)) + ((g2177) & (g3349) & (!sk[45]) & (!g1259)) + ((g2177) & (g3349) & (!sk[45]) & (g1259)) + ((g2177) & (g3349) & (sk[45]) & (!g1259)) + ((g2177) & (g3349) & (sk[45]) & (g1259)));
	assign g4783 = (((!g2178) & (!g3349) & (!sk[46]) & (g1260)) + ((!g2178) & (!g3349) & (sk[46]) & (g1260)) + ((!g2178) & (g3349) & (!sk[46]) & (!g1260)) + ((!g2178) & (g3349) & (!sk[46]) & (g1260)) + ((!g2178) & (g3349) & (sk[46]) & (g1260)) + ((g2178) & (!g3349) & (!sk[46]) & (g1260)) + ((g2178) & (g3349) & (!sk[46]) & (!g1260)) + ((g2178) & (g3349) & (!sk[46]) & (g1260)) + ((g2178) & (g3349) & (sk[46]) & (!g1260)) + ((g2178) & (g3349) & (sk[46]) & (g1260)));
	assign g4784 = (((!g2179) & (!sk[47]) & (!g3349) & (g1261)) + ((!g2179) & (!sk[47]) & (g3349) & (!g1261)) + ((!g2179) & (!sk[47]) & (g3349) & (g1261)) + ((!g2179) & (sk[47]) & (!g3349) & (g1261)) + ((!g2179) & (sk[47]) & (g3349) & (g1261)) + ((g2179) & (!sk[47]) & (!g3349) & (g1261)) + ((g2179) & (!sk[47]) & (g3349) & (!g1261)) + ((g2179) & (!sk[47]) & (g3349) & (g1261)) + ((g2179) & (sk[47]) & (g3349) & (!g1261)) + ((g2179) & (sk[47]) & (g3349) & (g1261)));
	assign g1262 = (((!g165) & (!g166) & (!sk[48]) & (!g1259) & (g1260) & (!g1261)) + ((!g165) & (!g166) & (!sk[48]) & (!g1259) & (g1260) & (g1261)) + ((!g165) & (!g166) & (!sk[48]) & (g1259) & (!g1260) & (!g1261)) + ((!g165) & (!g166) & (!sk[48]) & (g1259) & (!g1260) & (g1261)) + ((!g165) & (!g166) & (!sk[48]) & (g1259) & (g1260) & (!g1261)) + ((!g165) & (!g166) & (!sk[48]) & (g1259) & (g1260) & (g1261)) + ((!g165) & (g166) & (!sk[48]) & (!g1259) & (!g1260) & (!g1261)) + ((!g165) & (g166) & (!sk[48]) & (!g1259) & (!g1260) & (g1261)) + ((!g165) & (g166) & (!sk[48]) & (!g1259) & (g1260) & (!g1261)) + ((!g165) & (g166) & (!sk[48]) & (!g1259) & (g1260) & (g1261)) + ((!g165) & (g166) & (!sk[48]) & (g1259) & (!g1260) & (!g1261)) + ((!g165) & (g166) & (!sk[48]) & (g1259) & (!g1260) & (g1261)) + ((!g165) & (g166) & (!sk[48]) & (g1259) & (g1260) & (!g1261)) + ((!g165) & (g166) & (!sk[48]) & (g1259) & (g1260) & (g1261)) + ((!g165) & (g166) & (sk[48]) & (!g1259) & (!g1260) & (g1261)) + ((!g165) & (g166) & (sk[48]) & (!g1259) & (g1260) & (g1261)) + ((!g165) & (g166) & (sk[48]) & (g1259) & (!g1260) & (g1261)) + ((!g165) & (g166) & (sk[48]) & (g1259) & (g1260) & (g1261)) + ((g165) & (!g166) & (!sk[48]) & (!g1259) & (g1260) & (!g1261)) + ((g165) & (!g166) & (!sk[48]) & (!g1259) & (g1260) & (g1261)) + ((g165) & (!g166) & (!sk[48]) & (g1259) & (!g1260) & (!g1261)) + ((g165) & (!g166) & (!sk[48]) & (g1259) & (!g1260) & (g1261)) + ((g165) & (!g166) & (!sk[48]) & (g1259) & (g1260) & (!g1261)) + ((g165) & (!g166) & (!sk[48]) & (g1259) & (g1260) & (g1261)) + ((g165) & (!g166) & (sk[48]) & (g1259) & (!g1260) & (!g1261)) + ((g165) & (!g166) & (sk[48]) & (g1259) & (!g1260) & (g1261)) + ((g165) & (!g166) & (sk[48]) & (g1259) & (g1260) & (!g1261)) + ((g165) & (!g166) & (sk[48]) & (g1259) & (g1260) & (g1261)) + ((g165) & (g166) & (!sk[48]) & (!g1259) & (!g1260) & (!g1261)) + ((g165) & (g166) & (!sk[48]) & (!g1259) & (!g1260) & (g1261)) + ((g165) & (g166) & (!sk[48]) & (!g1259) & (g1260) & (!g1261)) + ((g165) & (g166) & (!sk[48]) & (!g1259) & (g1260) & (g1261)) + ((g165) & (g166) & (!sk[48]) & (g1259) & (!g1260) & (!g1261)) + ((g165) & (g166) & (!sk[48]) & (g1259) & (!g1260) & (g1261)) + ((g165) & (g166) & (!sk[48]) & (g1259) & (g1260) & (!g1261)) + ((g165) & (g166) & (!sk[48]) & (g1259) & (g1260) & (g1261)) + ((g165) & (g166) & (sk[48]) & (!g1259) & (g1260) & (!g1261)) + ((g165) & (g166) & (sk[48]) & (!g1259) & (g1260) & (g1261)) + ((g165) & (g166) & (sk[48]) & (g1259) & (g1260) & (!g1261)) + ((g165) & (g166) & (sk[48]) & (g1259) & (g1260) & (g1261)));
	assign g4785 = (((!sk[49]) & (!g2162) & (!g3349) & (g1263)) + ((!sk[49]) & (!g2162) & (g3349) & (!g1263)) + ((!sk[49]) & (!g2162) & (g3349) & (g1263)) + ((!sk[49]) & (g2162) & (!g3349) & (g1263)) + ((!sk[49]) & (g2162) & (g3349) & (!g1263)) + ((!sk[49]) & (g2162) & (g3349) & (g1263)) + ((sk[49]) & (!g2162) & (!g3349) & (g1263)) + ((sk[49]) & (!g2162) & (g3349) & (g1263)) + ((sk[49]) & (g2162) & (g3349) & (!g1263)) + ((sk[49]) & (g2162) & (g3349) & (g1263)));
	assign g4786 = (((!sk[50]) & (!g2164) & (!g3349) & (g1264)) + ((!sk[50]) & (!g2164) & (g3349) & (!g1264)) + ((!sk[50]) & (!g2164) & (g3349) & (g1264)) + ((!sk[50]) & (g2164) & (!g3349) & (g1264)) + ((!sk[50]) & (g2164) & (g3349) & (!g1264)) + ((!sk[50]) & (g2164) & (g3349) & (g1264)) + ((sk[50]) & (!g2164) & (!g3349) & (g1264)) + ((sk[50]) & (!g2164) & (g3349) & (g1264)) + ((sk[50]) & (g2164) & (g3349) & (!g1264)) + ((sk[50]) & (g2164) & (g3349) & (g1264)));
	assign g4787 = (((!sk[51]) & (!g2166) & (!g3349) & (g1265)) + ((!sk[51]) & (!g2166) & (g3349) & (!g1265)) + ((!sk[51]) & (!g2166) & (g3349) & (g1265)) + ((!sk[51]) & (g2166) & (!g3349) & (g1265)) + ((!sk[51]) & (g2166) & (g3349) & (!g1265)) + ((!sk[51]) & (g2166) & (g3349) & (g1265)) + ((sk[51]) & (!g2166) & (!g3349) & (g1265)) + ((sk[51]) & (!g2166) & (g3349) & (g1265)) + ((sk[51]) & (g2166) & (g3349) & (!g1265)) + ((sk[51]) & (g2166) & (g3349) & (g1265)));
	assign g4788 = (((!g2168) & (!sk[52]) & (!g3349) & (g1266)) + ((!g2168) & (!sk[52]) & (g3349) & (!g1266)) + ((!g2168) & (!sk[52]) & (g3349) & (g1266)) + ((!g2168) & (sk[52]) & (!g3349) & (g1266)) + ((!g2168) & (sk[52]) & (g3349) & (g1266)) + ((g2168) & (!sk[52]) & (!g3349) & (g1266)) + ((g2168) & (!sk[52]) & (g3349) & (!g1266)) + ((g2168) & (!sk[52]) & (g3349) & (g1266)) + ((g2168) & (sk[52]) & (g3349) & (!g1266)) + ((g2168) & (sk[52]) & (g3349) & (g1266)));
	assign g1267 = (((!g1263) & (!g1264) & (!g1265) & (g1266) & (g165) & (g166)) + ((!g1263) & (!g1264) & (g1265) & (!g1266) & (!g165) & (g166)) + ((!g1263) & (!g1264) & (g1265) & (g1266) & (!g165) & (g166)) + ((!g1263) & (!g1264) & (g1265) & (g1266) & (g165) & (g166)) + ((!g1263) & (g1264) & (!g1265) & (!g1266) & (g165) & (!g166)) + ((!g1263) & (g1264) & (!g1265) & (g1266) & (g165) & (!g166)) + ((!g1263) & (g1264) & (!g1265) & (g1266) & (g165) & (g166)) + ((!g1263) & (g1264) & (g1265) & (!g1266) & (!g165) & (g166)) + ((!g1263) & (g1264) & (g1265) & (!g1266) & (g165) & (!g166)) + ((!g1263) & (g1264) & (g1265) & (g1266) & (!g165) & (g166)) + ((!g1263) & (g1264) & (g1265) & (g1266) & (g165) & (!g166)) + ((!g1263) & (g1264) & (g1265) & (g1266) & (g165) & (g166)) + ((g1263) & (!g1264) & (!g1265) & (!g1266) & (!g165) & (!g166)) + ((g1263) & (!g1264) & (!g1265) & (g1266) & (!g165) & (!g166)) + ((g1263) & (!g1264) & (!g1265) & (g1266) & (g165) & (g166)) + ((g1263) & (!g1264) & (g1265) & (!g1266) & (!g165) & (!g166)) + ((g1263) & (!g1264) & (g1265) & (!g1266) & (!g165) & (g166)) + ((g1263) & (!g1264) & (g1265) & (g1266) & (!g165) & (!g166)) + ((g1263) & (!g1264) & (g1265) & (g1266) & (!g165) & (g166)) + ((g1263) & (!g1264) & (g1265) & (g1266) & (g165) & (g166)) + ((g1263) & (g1264) & (!g1265) & (!g1266) & (!g165) & (!g166)) + ((g1263) & (g1264) & (!g1265) & (!g1266) & (g165) & (!g166)) + ((g1263) & (g1264) & (!g1265) & (g1266) & (!g165) & (!g166)) + ((g1263) & (g1264) & (!g1265) & (g1266) & (g165) & (!g166)) + ((g1263) & (g1264) & (!g1265) & (g1266) & (g165) & (g166)) + ((g1263) & (g1264) & (g1265) & (!g1266) & (!g165) & (!g166)) + ((g1263) & (g1264) & (g1265) & (!g1266) & (!g165) & (g166)) + ((g1263) & (g1264) & (g1265) & (!g1266) & (g165) & (!g166)) + ((g1263) & (g1264) & (g1265) & (g1266) & (!g165) & (!g166)) + ((g1263) & (g1264) & (g1265) & (g1266) & (!g165) & (g166)) + ((g1263) & (g1264) & (g1265) & (g1266) & (g165) & (!g166)) + ((g1263) & (g1264) & (g1265) & (g1266) & (g165) & (g166)));
	assign g4789 = (((!sk[54]) & (!g2169) & (!g3349) & (g1268)) + ((!sk[54]) & (!g2169) & (g3349) & (!g1268)) + ((!sk[54]) & (!g2169) & (g3349) & (g1268)) + ((!sk[54]) & (g2169) & (!g3349) & (g1268)) + ((!sk[54]) & (g2169) & (g3349) & (!g1268)) + ((!sk[54]) & (g2169) & (g3349) & (g1268)) + ((sk[54]) & (!g2169) & (!g3349) & (g1268)) + ((sk[54]) & (!g2169) & (g3349) & (g1268)) + ((sk[54]) & (g2169) & (g3349) & (!g1268)) + ((sk[54]) & (g2169) & (g3349) & (g1268)));
	assign g4790 = (((!g2170) & (!sk[55]) & (!g3349) & (g1269)) + ((!g2170) & (!sk[55]) & (g3349) & (!g1269)) + ((!g2170) & (!sk[55]) & (g3349) & (g1269)) + ((!g2170) & (sk[55]) & (!g3349) & (g1269)) + ((!g2170) & (sk[55]) & (g3349) & (g1269)) + ((g2170) & (!sk[55]) & (!g3349) & (g1269)) + ((g2170) & (!sk[55]) & (g3349) & (!g1269)) + ((g2170) & (!sk[55]) & (g3349) & (g1269)) + ((g2170) & (sk[55]) & (g3349) & (!g1269)) + ((g2170) & (sk[55]) & (g3349) & (g1269)));
	assign g4791 = (((!sk[56]) & (!g2171) & (!g3349) & (g1270)) + ((!sk[56]) & (!g2171) & (g3349) & (!g1270)) + ((!sk[56]) & (!g2171) & (g3349) & (g1270)) + ((!sk[56]) & (g2171) & (!g3349) & (g1270)) + ((!sk[56]) & (g2171) & (g3349) & (!g1270)) + ((!sk[56]) & (g2171) & (g3349) & (g1270)) + ((sk[56]) & (!g2171) & (!g3349) & (g1270)) + ((sk[56]) & (!g2171) & (g3349) & (g1270)) + ((sk[56]) & (g2171) & (g3349) & (!g1270)) + ((sk[56]) & (g2171) & (g3349) & (g1270)));
	assign g4792 = (((!g2172) & (!g3349) & (!sk[57]) & (g1271)) + ((!g2172) & (!g3349) & (sk[57]) & (g1271)) + ((!g2172) & (g3349) & (!sk[57]) & (!g1271)) + ((!g2172) & (g3349) & (!sk[57]) & (g1271)) + ((!g2172) & (g3349) & (sk[57]) & (g1271)) + ((g2172) & (!g3349) & (!sk[57]) & (g1271)) + ((g2172) & (g3349) & (!sk[57]) & (!g1271)) + ((g2172) & (g3349) & (!sk[57]) & (g1271)) + ((g2172) & (g3349) & (sk[57]) & (!g1271)) + ((g2172) & (g3349) & (sk[57]) & (g1271)));
	assign g1272 = (((!g1268) & (!g1269) & (!g1270) & (g1271) & (g165) & (g166)) + ((!g1268) & (!g1269) & (g1270) & (!g1271) & (!g165) & (g166)) + ((!g1268) & (!g1269) & (g1270) & (g1271) & (!g165) & (g166)) + ((!g1268) & (!g1269) & (g1270) & (g1271) & (g165) & (g166)) + ((!g1268) & (g1269) & (!g1270) & (!g1271) & (g165) & (!g166)) + ((!g1268) & (g1269) & (!g1270) & (g1271) & (g165) & (!g166)) + ((!g1268) & (g1269) & (!g1270) & (g1271) & (g165) & (g166)) + ((!g1268) & (g1269) & (g1270) & (!g1271) & (!g165) & (g166)) + ((!g1268) & (g1269) & (g1270) & (!g1271) & (g165) & (!g166)) + ((!g1268) & (g1269) & (g1270) & (g1271) & (!g165) & (g166)) + ((!g1268) & (g1269) & (g1270) & (g1271) & (g165) & (!g166)) + ((!g1268) & (g1269) & (g1270) & (g1271) & (g165) & (g166)) + ((g1268) & (!g1269) & (!g1270) & (!g1271) & (!g165) & (!g166)) + ((g1268) & (!g1269) & (!g1270) & (g1271) & (!g165) & (!g166)) + ((g1268) & (!g1269) & (!g1270) & (g1271) & (g165) & (g166)) + ((g1268) & (!g1269) & (g1270) & (!g1271) & (!g165) & (!g166)) + ((g1268) & (!g1269) & (g1270) & (!g1271) & (!g165) & (g166)) + ((g1268) & (!g1269) & (g1270) & (g1271) & (!g165) & (!g166)) + ((g1268) & (!g1269) & (g1270) & (g1271) & (!g165) & (g166)) + ((g1268) & (!g1269) & (g1270) & (g1271) & (g165) & (g166)) + ((g1268) & (g1269) & (!g1270) & (!g1271) & (!g165) & (!g166)) + ((g1268) & (g1269) & (!g1270) & (!g1271) & (g165) & (!g166)) + ((g1268) & (g1269) & (!g1270) & (g1271) & (!g165) & (!g166)) + ((g1268) & (g1269) & (!g1270) & (g1271) & (g165) & (!g166)) + ((g1268) & (g1269) & (!g1270) & (g1271) & (g165) & (g166)) + ((g1268) & (g1269) & (g1270) & (!g1271) & (!g165) & (!g166)) + ((g1268) & (g1269) & (g1270) & (!g1271) & (!g165) & (g166)) + ((g1268) & (g1269) & (g1270) & (!g1271) & (g165) & (!g166)) + ((g1268) & (g1269) & (g1270) & (g1271) & (!g165) & (!g166)) + ((g1268) & (g1269) & (g1270) & (g1271) & (!g165) & (g166)) + ((g1268) & (g1269) & (g1270) & (g1271) & (g165) & (!g166)) + ((g1268) & (g1269) & (g1270) & (g1271) & (g165) & (g166)));
	assign g1273 = (((!g147) & (!g148) & (!g1258) & (g1262) & (!g1267) & (!g1272)) + ((!g147) & (!g148) & (!g1258) & (g1262) & (!g1267) & (g1272)) + ((!g147) & (!g148) & (!g1258) & (g1262) & (g1267) & (!g1272)) + ((!g147) & (!g148) & (!g1258) & (g1262) & (g1267) & (g1272)) + ((!g147) & (!g148) & (g1258) & (g1262) & (!g1267) & (!g1272)) + ((!g147) & (!g148) & (g1258) & (g1262) & (!g1267) & (g1272)) + ((!g147) & (!g148) & (g1258) & (g1262) & (g1267) & (!g1272)) + ((!g147) & (!g148) & (g1258) & (g1262) & (g1267) & (g1272)) + ((!g147) & (g148) & (!g1258) & (!g1262) & (!g1267) & (g1272)) + ((!g147) & (g148) & (!g1258) & (!g1262) & (g1267) & (g1272)) + ((!g147) & (g148) & (!g1258) & (g1262) & (!g1267) & (g1272)) + ((!g147) & (g148) & (!g1258) & (g1262) & (g1267) & (g1272)) + ((!g147) & (g148) & (g1258) & (!g1262) & (!g1267) & (g1272)) + ((!g147) & (g148) & (g1258) & (!g1262) & (g1267) & (g1272)) + ((!g147) & (g148) & (g1258) & (g1262) & (!g1267) & (g1272)) + ((!g147) & (g148) & (g1258) & (g1262) & (g1267) & (g1272)) + ((g147) & (!g148) & (g1258) & (!g1262) & (!g1267) & (!g1272)) + ((g147) & (!g148) & (g1258) & (!g1262) & (!g1267) & (g1272)) + ((g147) & (!g148) & (g1258) & (!g1262) & (g1267) & (!g1272)) + ((g147) & (!g148) & (g1258) & (!g1262) & (g1267) & (g1272)) + ((g147) & (!g148) & (g1258) & (g1262) & (!g1267) & (!g1272)) + ((g147) & (!g148) & (g1258) & (g1262) & (!g1267) & (g1272)) + ((g147) & (!g148) & (g1258) & (g1262) & (g1267) & (!g1272)) + ((g147) & (!g148) & (g1258) & (g1262) & (g1267) & (g1272)) + ((g147) & (g148) & (!g1258) & (!g1262) & (g1267) & (!g1272)) + ((g147) & (g148) & (!g1258) & (!g1262) & (g1267) & (g1272)) + ((g147) & (g148) & (!g1258) & (g1262) & (g1267) & (!g1272)) + ((g147) & (g148) & (!g1258) & (g1262) & (g1267) & (g1272)) + ((g147) & (g148) & (g1258) & (!g1262) & (g1267) & (!g1272)) + ((g147) & (g148) & (g1258) & (!g1262) & (g1267) & (g1272)) + ((g147) & (g148) & (g1258) & (g1262) & (g1267) & (!g1272)) + ((g147) & (g148) & (g1258) & (g1262) & (g1267) & (g1272)));
	assign g1274 = (((!sk[60]) & (!g142) & (!g1253) & (g1273)) + ((!sk[60]) & (!g142) & (g1253) & (!g1273)) + ((!sk[60]) & (!g142) & (g1253) & (g1273)) + ((!sk[60]) & (g142) & (!g1253) & (g1273)) + ((!sk[60]) & (g142) & (g1253) & (!g1273)) + ((!sk[60]) & (g142) & (g1253) & (g1273)) + ((sk[60]) & (!g142) & (!g1253) & (g1273)) + ((sk[60]) & (!g142) & (g1253) & (g1273)) + ((sk[60]) & (g142) & (g1253) & (!g1273)) + ((sk[60]) & (g142) & (g1253) & (g1273)));
	assign g4793 = (((!g2059) & (!sk[61]) & (!g2714) & (g1275)) + ((!g2059) & (!sk[61]) & (g2714) & (!g1275)) + ((!g2059) & (!sk[61]) & (g2714) & (g1275)) + ((!g2059) & (sk[61]) & (!g2714) & (g1275)) + ((!g2059) & (sk[61]) & (g2714) & (g1275)) + ((g2059) & (!sk[61]) & (!g2714) & (g1275)) + ((g2059) & (!sk[61]) & (g2714) & (!g1275)) + ((g2059) & (!sk[61]) & (g2714) & (g1275)) + ((g2059) & (sk[61]) & (g2714) & (!g1275)) + ((g2059) & (sk[61]) & (g2714) & (g1275)));
	assign g1276 = (((!sk[62]) & (!g1229) & (!g1231) & (g916)) + ((!sk[62]) & (!g1229) & (g1231) & (!g916)) + ((!sk[62]) & (!g1229) & (g1231) & (g916)) + ((!sk[62]) & (g1229) & (!g1231) & (g916)) + ((!sk[62]) & (g1229) & (g1231) & (!g916)) + ((!sk[62]) & (g1229) & (g1231) & (g916)) + ((sk[62]) & (!g1229) & (g1231) & (!g916)) + ((sk[62]) & (g1229) & (!g1231) & (!g916)) + ((sk[62]) & (g1229) & (g1231) & (!g916)) + ((sk[62]) & (g1229) & (g1231) & (g916)));
	assign g1277 = (((!sk[63]) & (!g126) & (!g1274) & (!g1275) & (g1276) & (!g916)) + ((!sk[63]) & (!g126) & (!g1274) & (!g1275) & (g1276) & (g916)) + ((!sk[63]) & (!g126) & (!g1274) & (g1275) & (!g1276) & (!g916)) + ((!sk[63]) & (!g126) & (!g1274) & (g1275) & (!g1276) & (g916)) + ((!sk[63]) & (!g126) & (!g1274) & (g1275) & (g1276) & (!g916)) + ((!sk[63]) & (!g126) & (!g1274) & (g1275) & (g1276) & (g916)) + ((!sk[63]) & (!g126) & (g1274) & (!g1275) & (!g1276) & (!g916)) + ((!sk[63]) & (!g126) & (g1274) & (!g1275) & (!g1276) & (g916)) + ((!sk[63]) & (!g126) & (g1274) & (!g1275) & (g1276) & (!g916)) + ((!sk[63]) & (!g126) & (g1274) & (!g1275) & (g1276) & (g916)) + ((!sk[63]) & (!g126) & (g1274) & (g1275) & (!g1276) & (!g916)) + ((!sk[63]) & (!g126) & (g1274) & (g1275) & (!g1276) & (g916)) + ((!sk[63]) & (!g126) & (g1274) & (g1275) & (g1276) & (!g916)) + ((!sk[63]) & (!g126) & (g1274) & (g1275) & (g1276) & (g916)) + ((!sk[63]) & (g126) & (!g1274) & (!g1275) & (g1276) & (!g916)) + ((!sk[63]) & (g126) & (!g1274) & (!g1275) & (g1276) & (g916)) + ((!sk[63]) & (g126) & (!g1274) & (g1275) & (!g1276) & (!g916)) + ((!sk[63]) & (g126) & (!g1274) & (g1275) & (!g1276) & (g916)) + ((!sk[63]) & (g126) & (!g1274) & (g1275) & (g1276) & (!g916)) + ((!sk[63]) & (g126) & (!g1274) & (g1275) & (g1276) & (g916)) + ((!sk[63]) & (g126) & (g1274) & (!g1275) & (!g1276) & (!g916)) + ((!sk[63]) & (g126) & (g1274) & (!g1275) & (!g1276) & (g916)) + ((!sk[63]) & (g126) & (g1274) & (!g1275) & (g1276) & (!g916)) + ((!sk[63]) & (g126) & (g1274) & (!g1275) & (g1276) & (g916)) + ((!sk[63]) & (g126) & (g1274) & (g1275) & (!g1276) & (!g916)) + ((!sk[63]) & (g126) & (g1274) & (g1275) & (!g1276) & (g916)) + ((!sk[63]) & (g126) & (g1274) & (g1275) & (g1276) & (!g916)) + ((!sk[63]) & (g126) & (g1274) & (g1275) & (g1276) & (g916)) + ((sk[63]) & (!g126) & (!g1274) & (g1275) & (!g1276) & (!g916)) + ((sk[63]) & (!g126) & (!g1274) & (g1275) & (!g1276) & (g916)) + ((sk[63]) & (!g126) & (!g1274) & (g1275) & (g1276) & (!g916)) + ((sk[63]) & (!g126) & (!g1274) & (g1275) & (g1276) & (g916)) + ((sk[63]) & (!g126) & (g1274) & (g1275) & (!g1276) & (!g916)) + ((sk[63]) & (!g126) & (g1274) & (g1275) & (!g1276) & (g916)) + ((sk[63]) & (!g126) & (g1274) & (g1275) & (g1276) & (!g916)) + ((sk[63]) & (!g126) & (g1274) & (g1275) & (g1276) & (g916)) + ((sk[63]) & (g126) & (!g1274) & (!g1275) & (!g1276) & (!g916)) + ((sk[63]) & (g126) & (!g1274) & (!g1275) & (g1276) & (g916)) + ((sk[63]) & (g126) & (!g1274) & (g1275) & (!g1276) & (!g916)) + ((sk[63]) & (g126) & (!g1274) & (g1275) & (g1276) & (g916)) + ((sk[63]) & (g126) & (g1274) & (!g1275) & (!g1276) & (g916)) + ((sk[63]) & (g126) & (g1274) & (!g1275) & (g1276) & (!g916)) + ((sk[63]) & (g126) & (g1274) & (g1275) & (!g1276) & (g916)) + ((sk[63]) & (g126) & (g1274) & (g1275) & (g1276) & (!g916)));
	assign g4794 = (((!g2140) & (!g3325) & (!sk[64]) & (g1278)) + ((!g2140) & (!g3325) & (sk[64]) & (g1278)) + ((!g2140) & (g3325) & (!sk[64]) & (!g1278)) + ((!g2140) & (g3325) & (!sk[64]) & (g1278)) + ((!g2140) & (g3325) & (sk[64]) & (g1278)) + ((g2140) & (!g3325) & (!sk[64]) & (g1278)) + ((g2140) & (g3325) & (!sk[64]) & (!g1278)) + ((g2140) & (g3325) & (!sk[64]) & (g1278)) + ((g2140) & (g3325) & (sk[64]) & (!g1278)) + ((g2140) & (g3325) & (sk[64]) & (g1278)));
	assign g4795 = (((!sk[65]) & (!g2142) & (!g3325) & (g1279)) + ((!sk[65]) & (!g2142) & (g3325) & (!g1279)) + ((!sk[65]) & (!g2142) & (g3325) & (g1279)) + ((!sk[65]) & (g2142) & (!g3325) & (g1279)) + ((!sk[65]) & (g2142) & (g3325) & (!g1279)) + ((!sk[65]) & (g2142) & (g3325) & (g1279)) + ((sk[65]) & (!g2142) & (!g3325) & (g1279)) + ((sk[65]) & (!g2142) & (g3325) & (g1279)) + ((sk[65]) & (g2142) & (g3325) & (!g1279)) + ((sk[65]) & (g2142) & (g3325) & (g1279)));
	assign g4796 = (((!sk[66]) & (!g2144) & (!g3325) & (g1280)) + ((!sk[66]) & (!g2144) & (g3325) & (!g1280)) + ((!sk[66]) & (!g2144) & (g3325) & (g1280)) + ((!sk[66]) & (g2144) & (!g3325) & (g1280)) + ((!sk[66]) & (g2144) & (g3325) & (!g1280)) + ((!sk[66]) & (g2144) & (g3325) & (g1280)) + ((sk[66]) & (!g2144) & (!g3325) & (g1280)) + ((sk[66]) & (!g2144) & (g3325) & (g1280)) + ((sk[66]) & (g2144) & (g3325) & (!g1280)) + ((sk[66]) & (g2144) & (g3325) & (g1280)));
	assign g4797 = (((!g2145) & (!sk[67]) & (!g3325) & (g1281)) + ((!g2145) & (!sk[67]) & (g3325) & (!g1281)) + ((!g2145) & (!sk[67]) & (g3325) & (g1281)) + ((!g2145) & (sk[67]) & (!g3325) & (g1281)) + ((!g2145) & (sk[67]) & (g3325) & (g1281)) + ((g2145) & (!sk[67]) & (!g3325) & (g1281)) + ((g2145) & (!sk[67]) & (g3325) & (!g1281)) + ((g2145) & (!sk[67]) & (g3325) & (g1281)) + ((g2145) & (sk[67]) & (g3325) & (!g1281)) + ((g2145) & (sk[67]) & (g3325) & (g1281)));
	assign g1282 = (((!g1278) & (!g1279) & (!g1280) & (g1281) & (g147) & (g148)) + ((!g1278) & (!g1279) & (g1280) & (!g1281) & (!g147) & (g148)) + ((!g1278) & (!g1279) & (g1280) & (g1281) & (!g147) & (g148)) + ((!g1278) & (!g1279) & (g1280) & (g1281) & (g147) & (g148)) + ((!g1278) & (g1279) & (!g1280) & (!g1281) & (g147) & (!g148)) + ((!g1278) & (g1279) & (!g1280) & (g1281) & (g147) & (!g148)) + ((!g1278) & (g1279) & (!g1280) & (g1281) & (g147) & (g148)) + ((!g1278) & (g1279) & (g1280) & (!g1281) & (!g147) & (g148)) + ((!g1278) & (g1279) & (g1280) & (!g1281) & (g147) & (!g148)) + ((!g1278) & (g1279) & (g1280) & (g1281) & (!g147) & (g148)) + ((!g1278) & (g1279) & (g1280) & (g1281) & (g147) & (!g148)) + ((!g1278) & (g1279) & (g1280) & (g1281) & (g147) & (g148)) + ((g1278) & (!g1279) & (!g1280) & (!g1281) & (!g147) & (!g148)) + ((g1278) & (!g1279) & (!g1280) & (g1281) & (!g147) & (!g148)) + ((g1278) & (!g1279) & (!g1280) & (g1281) & (g147) & (g148)) + ((g1278) & (!g1279) & (g1280) & (!g1281) & (!g147) & (!g148)) + ((g1278) & (!g1279) & (g1280) & (!g1281) & (!g147) & (g148)) + ((g1278) & (!g1279) & (g1280) & (g1281) & (!g147) & (!g148)) + ((g1278) & (!g1279) & (g1280) & (g1281) & (!g147) & (g148)) + ((g1278) & (!g1279) & (g1280) & (g1281) & (g147) & (g148)) + ((g1278) & (g1279) & (!g1280) & (!g1281) & (!g147) & (!g148)) + ((g1278) & (g1279) & (!g1280) & (!g1281) & (g147) & (!g148)) + ((g1278) & (g1279) & (!g1280) & (g1281) & (!g147) & (!g148)) + ((g1278) & (g1279) & (!g1280) & (g1281) & (g147) & (!g148)) + ((g1278) & (g1279) & (!g1280) & (g1281) & (g147) & (g148)) + ((g1278) & (g1279) & (g1280) & (!g1281) & (!g147) & (!g148)) + ((g1278) & (g1279) & (g1280) & (!g1281) & (!g147) & (g148)) + ((g1278) & (g1279) & (g1280) & (!g1281) & (g147) & (!g148)) + ((g1278) & (g1279) & (g1280) & (g1281) & (!g147) & (!g148)) + ((g1278) & (g1279) & (g1280) & (g1281) & (!g147) & (g148)) + ((g1278) & (g1279) & (g1280) & (g1281) & (g147) & (!g148)) + ((g1278) & (g1279) & (g1280) & (g1281) & (g147) & (g148)));
	assign g4798 = (((!sk[69]) & (!g2146) & (!g3325) & (g1283)) + ((!sk[69]) & (!g2146) & (g3325) & (!g1283)) + ((!sk[69]) & (!g2146) & (g3325) & (g1283)) + ((!sk[69]) & (g2146) & (!g3325) & (g1283)) + ((!sk[69]) & (g2146) & (g3325) & (!g1283)) + ((!sk[69]) & (g2146) & (g3325) & (g1283)) + ((sk[69]) & (!g2146) & (!g3325) & (g1283)) + ((sk[69]) & (!g2146) & (g3325) & (g1283)) + ((sk[69]) & (g2146) & (g3325) & (!g1283)) + ((sk[69]) & (g2146) & (g3325) & (g1283)));
	assign g4799 = (((!sk[70]) & (!g2148) & (!g3325) & (g1284)) + ((!sk[70]) & (!g2148) & (g3325) & (!g1284)) + ((!sk[70]) & (!g2148) & (g3325) & (g1284)) + ((!sk[70]) & (g2148) & (!g3325) & (g1284)) + ((!sk[70]) & (g2148) & (g3325) & (!g1284)) + ((!sk[70]) & (g2148) & (g3325) & (g1284)) + ((sk[70]) & (!g2148) & (!g3325) & (g1284)) + ((sk[70]) & (!g2148) & (g3325) & (g1284)) + ((sk[70]) & (g2148) & (g3325) & (!g1284)) + ((sk[70]) & (g2148) & (g3325) & (g1284)));
	assign g4800 = (((!g2150) & (!g3325) & (!sk[71]) & (g1285)) + ((!g2150) & (!g3325) & (sk[71]) & (g1285)) + ((!g2150) & (g3325) & (!sk[71]) & (!g1285)) + ((!g2150) & (g3325) & (!sk[71]) & (g1285)) + ((!g2150) & (g3325) & (sk[71]) & (g1285)) + ((g2150) & (!g3325) & (!sk[71]) & (g1285)) + ((g2150) & (g3325) & (!sk[71]) & (!g1285)) + ((g2150) & (g3325) & (!sk[71]) & (g1285)) + ((g2150) & (g3325) & (sk[71]) & (!g1285)) + ((g2150) & (g3325) & (sk[71]) & (g1285)));
	assign g4801 = (((!sk[72]) & (!g2151) & (!g3325) & (g1286)) + ((!sk[72]) & (!g2151) & (g3325) & (!g1286)) + ((!sk[72]) & (!g2151) & (g3325) & (g1286)) + ((!sk[72]) & (g2151) & (!g3325) & (g1286)) + ((!sk[72]) & (g2151) & (g3325) & (!g1286)) + ((!sk[72]) & (g2151) & (g3325) & (g1286)) + ((sk[72]) & (!g2151) & (!g3325) & (g1286)) + ((sk[72]) & (!g2151) & (g3325) & (g1286)) + ((sk[72]) & (g2151) & (g3325) & (!g1286)) + ((sk[72]) & (g2151) & (g3325) & (g1286)));
	assign g1287 = (((!g1283) & (!g1284) & (!g1285) & (g1286) & (g147) & (g148)) + ((!g1283) & (!g1284) & (g1285) & (!g1286) & (!g147) & (g148)) + ((!g1283) & (!g1284) & (g1285) & (g1286) & (!g147) & (g148)) + ((!g1283) & (!g1284) & (g1285) & (g1286) & (g147) & (g148)) + ((!g1283) & (g1284) & (!g1285) & (!g1286) & (g147) & (!g148)) + ((!g1283) & (g1284) & (!g1285) & (g1286) & (g147) & (!g148)) + ((!g1283) & (g1284) & (!g1285) & (g1286) & (g147) & (g148)) + ((!g1283) & (g1284) & (g1285) & (!g1286) & (!g147) & (g148)) + ((!g1283) & (g1284) & (g1285) & (!g1286) & (g147) & (!g148)) + ((!g1283) & (g1284) & (g1285) & (g1286) & (!g147) & (g148)) + ((!g1283) & (g1284) & (g1285) & (g1286) & (g147) & (!g148)) + ((!g1283) & (g1284) & (g1285) & (g1286) & (g147) & (g148)) + ((g1283) & (!g1284) & (!g1285) & (!g1286) & (!g147) & (!g148)) + ((g1283) & (!g1284) & (!g1285) & (g1286) & (!g147) & (!g148)) + ((g1283) & (!g1284) & (!g1285) & (g1286) & (g147) & (g148)) + ((g1283) & (!g1284) & (g1285) & (!g1286) & (!g147) & (!g148)) + ((g1283) & (!g1284) & (g1285) & (!g1286) & (!g147) & (g148)) + ((g1283) & (!g1284) & (g1285) & (g1286) & (!g147) & (!g148)) + ((g1283) & (!g1284) & (g1285) & (g1286) & (!g147) & (g148)) + ((g1283) & (!g1284) & (g1285) & (g1286) & (g147) & (g148)) + ((g1283) & (g1284) & (!g1285) & (!g1286) & (!g147) & (!g148)) + ((g1283) & (g1284) & (!g1285) & (!g1286) & (g147) & (!g148)) + ((g1283) & (g1284) & (!g1285) & (g1286) & (!g147) & (!g148)) + ((g1283) & (g1284) & (!g1285) & (g1286) & (g147) & (!g148)) + ((g1283) & (g1284) & (!g1285) & (g1286) & (g147) & (g148)) + ((g1283) & (g1284) & (g1285) & (!g1286) & (!g147) & (!g148)) + ((g1283) & (g1284) & (g1285) & (!g1286) & (!g147) & (g148)) + ((g1283) & (g1284) & (g1285) & (!g1286) & (g147) & (!g148)) + ((g1283) & (g1284) & (g1285) & (g1286) & (!g147) & (!g148)) + ((g1283) & (g1284) & (g1285) & (g1286) & (!g147) & (g148)) + ((g1283) & (g1284) & (g1285) & (g1286) & (g147) & (!g148)) + ((g1283) & (g1284) & (g1285) & (g1286) & (g147) & (g148)));
	assign g4802 = (((!g2152) & (!g3325) & (!sk[74]) & (g1288)) + ((!g2152) & (!g3325) & (sk[74]) & (g1288)) + ((!g2152) & (g3325) & (!sk[74]) & (!g1288)) + ((!g2152) & (g3325) & (!sk[74]) & (g1288)) + ((!g2152) & (g3325) & (sk[74]) & (g1288)) + ((g2152) & (!g3325) & (!sk[74]) & (g1288)) + ((g2152) & (g3325) & (!sk[74]) & (!g1288)) + ((g2152) & (g3325) & (!sk[74]) & (g1288)) + ((g2152) & (g3325) & (sk[74]) & (!g1288)) + ((g2152) & (g3325) & (sk[74]) & (g1288)));
	assign g4803 = (((!sk[75]) & (!g2153) & (!g3325) & (g1289)) + ((!sk[75]) & (!g2153) & (g3325) & (!g1289)) + ((!sk[75]) & (!g2153) & (g3325) & (g1289)) + ((!sk[75]) & (g2153) & (!g3325) & (g1289)) + ((!sk[75]) & (g2153) & (g3325) & (!g1289)) + ((!sk[75]) & (g2153) & (g3325) & (g1289)) + ((sk[75]) & (!g2153) & (!g3325) & (g1289)) + ((sk[75]) & (!g2153) & (g3325) & (g1289)) + ((sk[75]) & (g2153) & (g3325) & (!g1289)) + ((sk[75]) & (g2153) & (g3325) & (g1289)));
	assign g4804 = (((!sk[76]) & (!g2155) & (!g3325) & (g1290)) + ((!sk[76]) & (!g2155) & (g3325) & (!g1290)) + ((!sk[76]) & (!g2155) & (g3325) & (g1290)) + ((!sk[76]) & (g2155) & (!g3325) & (g1290)) + ((!sk[76]) & (g2155) & (g3325) & (!g1290)) + ((!sk[76]) & (g2155) & (g3325) & (g1290)) + ((sk[76]) & (!g2155) & (!g3325) & (g1290)) + ((sk[76]) & (!g2155) & (g3325) & (g1290)) + ((sk[76]) & (g2155) & (g3325) & (!g1290)) + ((sk[76]) & (g2155) & (g3325) & (g1290)));
	assign g4805 = (((!g2157) & (!g3325) & (!sk[77]) & (g1291)) + ((!g2157) & (!g3325) & (sk[77]) & (g1291)) + ((!g2157) & (g3325) & (!sk[77]) & (!g1291)) + ((!g2157) & (g3325) & (!sk[77]) & (g1291)) + ((!g2157) & (g3325) & (sk[77]) & (g1291)) + ((g2157) & (!g3325) & (!sk[77]) & (g1291)) + ((g2157) & (g3325) & (!sk[77]) & (!g1291)) + ((g2157) & (g3325) & (!sk[77]) & (g1291)) + ((g2157) & (g3325) & (sk[77]) & (!g1291)) + ((g2157) & (g3325) & (sk[77]) & (g1291)));
	assign g1292 = (((!g1288) & (!g1289) & (!g1290) & (g1291) & (g147) & (g148)) + ((!g1288) & (!g1289) & (g1290) & (!g1291) & (!g147) & (g148)) + ((!g1288) & (!g1289) & (g1290) & (g1291) & (!g147) & (g148)) + ((!g1288) & (!g1289) & (g1290) & (g1291) & (g147) & (g148)) + ((!g1288) & (g1289) & (!g1290) & (!g1291) & (g147) & (!g148)) + ((!g1288) & (g1289) & (!g1290) & (g1291) & (g147) & (!g148)) + ((!g1288) & (g1289) & (!g1290) & (g1291) & (g147) & (g148)) + ((!g1288) & (g1289) & (g1290) & (!g1291) & (!g147) & (g148)) + ((!g1288) & (g1289) & (g1290) & (!g1291) & (g147) & (!g148)) + ((!g1288) & (g1289) & (g1290) & (g1291) & (!g147) & (g148)) + ((!g1288) & (g1289) & (g1290) & (g1291) & (g147) & (!g148)) + ((!g1288) & (g1289) & (g1290) & (g1291) & (g147) & (g148)) + ((g1288) & (!g1289) & (!g1290) & (!g1291) & (!g147) & (!g148)) + ((g1288) & (!g1289) & (!g1290) & (g1291) & (!g147) & (!g148)) + ((g1288) & (!g1289) & (!g1290) & (g1291) & (g147) & (g148)) + ((g1288) & (!g1289) & (g1290) & (!g1291) & (!g147) & (!g148)) + ((g1288) & (!g1289) & (g1290) & (!g1291) & (!g147) & (g148)) + ((g1288) & (!g1289) & (g1290) & (g1291) & (!g147) & (!g148)) + ((g1288) & (!g1289) & (g1290) & (g1291) & (!g147) & (g148)) + ((g1288) & (!g1289) & (g1290) & (g1291) & (g147) & (g148)) + ((g1288) & (g1289) & (!g1290) & (!g1291) & (!g147) & (!g148)) + ((g1288) & (g1289) & (!g1290) & (!g1291) & (g147) & (!g148)) + ((g1288) & (g1289) & (!g1290) & (g1291) & (!g147) & (!g148)) + ((g1288) & (g1289) & (!g1290) & (g1291) & (g147) & (!g148)) + ((g1288) & (g1289) & (!g1290) & (g1291) & (g147) & (g148)) + ((g1288) & (g1289) & (g1290) & (!g1291) & (!g147) & (!g148)) + ((g1288) & (g1289) & (g1290) & (!g1291) & (!g147) & (g148)) + ((g1288) & (g1289) & (g1290) & (!g1291) & (g147) & (!g148)) + ((g1288) & (g1289) & (g1290) & (g1291) & (!g147) & (!g148)) + ((g1288) & (g1289) & (g1290) & (g1291) & (!g147) & (g148)) + ((g1288) & (g1289) & (g1290) & (g1291) & (g147) & (!g148)) + ((g1288) & (g1289) & (g1290) & (g1291) & (g147) & (g148)));
	assign g4806 = (((!g2158) & (!g3325) & (!sk[79]) & (g1293)) + ((!g2158) & (!g3325) & (sk[79]) & (g1293)) + ((!g2158) & (g3325) & (!sk[79]) & (!g1293)) + ((!g2158) & (g3325) & (!sk[79]) & (g1293)) + ((!g2158) & (g3325) & (sk[79]) & (g1293)) + ((g2158) & (!g3325) & (!sk[79]) & (g1293)) + ((g2158) & (g3325) & (!sk[79]) & (!g1293)) + ((g2158) & (g3325) & (!sk[79]) & (g1293)) + ((g2158) & (g3325) & (sk[79]) & (!g1293)) + ((g2158) & (g3325) & (sk[79]) & (g1293)));
	assign g4807 = (((!g2159) & (!sk[80]) & (!g3325) & (g1294)) + ((!g2159) & (!sk[80]) & (g3325) & (!g1294)) + ((!g2159) & (!sk[80]) & (g3325) & (g1294)) + ((!g2159) & (sk[80]) & (!g3325) & (g1294)) + ((!g2159) & (sk[80]) & (g3325) & (g1294)) + ((g2159) & (!sk[80]) & (!g3325) & (g1294)) + ((g2159) & (!sk[80]) & (g3325) & (!g1294)) + ((g2159) & (!sk[80]) & (g3325) & (g1294)) + ((g2159) & (sk[80]) & (g3325) & (!g1294)) + ((g2159) & (sk[80]) & (g3325) & (g1294)));
	assign g4808 = (((!sk[81]) & (!g2160) & (!g3325) & (g1295)) + ((!sk[81]) & (!g2160) & (g3325) & (!g1295)) + ((!sk[81]) & (!g2160) & (g3325) & (g1295)) + ((!sk[81]) & (g2160) & (!g3325) & (g1295)) + ((!sk[81]) & (g2160) & (g3325) & (!g1295)) + ((!sk[81]) & (g2160) & (g3325) & (g1295)) + ((sk[81]) & (!g2160) & (!g3325) & (g1295)) + ((sk[81]) & (!g2160) & (g3325) & (g1295)) + ((sk[81]) & (g2160) & (g3325) & (!g1295)) + ((sk[81]) & (g2160) & (g3325) & (g1295)));
	assign g4809 = (((!sk[82]) & (!g2161) & (!g3325) & (g1296)) + ((!sk[82]) & (!g2161) & (g3325) & (!g1296)) + ((!sk[82]) & (!g2161) & (g3325) & (g1296)) + ((!sk[82]) & (g2161) & (!g3325) & (g1296)) + ((!sk[82]) & (g2161) & (g3325) & (!g1296)) + ((!sk[82]) & (g2161) & (g3325) & (g1296)) + ((sk[82]) & (!g2161) & (!g3325) & (g1296)) + ((sk[82]) & (!g2161) & (g3325) & (g1296)) + ((sk[82]) & (g2161) & (g3325) & (!g1296)) + ((sk[82]) & (g2161) & (g3325) & (g1296)));
	assign g1297 = (((!g1293) & (!g1294) & (!g1295) & (g1296) & (g147) & (g148)) + ((!g1293) & (!g1294) & (g1295) & (!g1296) & (!g147) & (g148)) + ((!g1293) & (!g1294) & (g1295) & (g1296) & (!g147) & (g148)) + ((!g1293) & (!g1294) & (g1295) & (g1296) & (g147) & (g148)) + ((!g1293) & (g1294) & (!g1295) & (!g1296) & (g147) & (!g148)) + ((!g1293) & (g1294) & (!g1295) & (g1296) & (g147) & (!g148)) + ((!g1293) & (g1294) & (!g1295) & (g1296) & (g147) & (g148)) + ((!g1293) & (g1294) & (g1295) & (!g1296) & (!g147) & (g148)) + ((!g1293) & (g1294) & (g1295) & (!g1296) & (g147) & (!g148)) + ((!g1293) & (g1294) & (g1295) & (g1296) & (!g147) & (g148)) + ((!g1293) & (g1294) & (g1295) & (g1296) & (g147) & (!g148)) + ((!g1293) & (g1294) & (g1295) & (g1296) & (g147) & (g148)) + ((g1293) & (!g1294) & (!g1295) & (!g1296) & (!g147) & (!g148)) + ((g1293) & (!g1294) & (!g1295) & (g1296) & (!g147) & (!g148)) + ((g1293) & (!g1294) & (!g1295) & (g1296) & (g147) & (g148)) + ((g1293) & (!g1294) & (g1295) & (!g1296) & (!g147) & (!g148)) + ((g1293) & (!g1294) & (g1295) & (!g1296) & (!g147) & (g148)) + ((g1293) & (!g1294) & (g1295) & (g1296) & (!g147) & (!g148)) + ((g1293) & (!g1294) & (g1295) & (g1296) & (!g147) & (g148)) + ((g1293) & (!g1294) & (g1295) & (g1296) & (g147) & (g148)) + ((g1293) & (g1294) & (!g1295) & (!g1296) & (!g147) & (!g148)) + ((g1293) & (g1294) & (!g1295) & (!g1296) & (g147) & (!g148)) + ((g1293) & (g1294) & (!g1295) & (g1296) & (!g147) & (!g148)) + ((g1293) & (g1294) & (!g1295) & (g1296) & (g147) & (!g148)) + ((g1293) & (g1294) & (!g1295) & (g1296) & (g147) & (g148)) + ((g1293) & (g1294) & (g1295) & (!g1296) & (!g147) & (!g148)) + ((g1293) & (g1294) & (g1295) & (!g1296) & (!g147) & (g148)) + ((g1293) & (g1294) & (g1295) & (!g1296) & (g147) & (!g148)) + ((g1293) & (g1294) & (g1295) & (g1296) & (!g147) & (!g148)) + ((g1293) & (g1294) & (g1295) & (g1296) & (!g147) & (g148)) + ((g1293) & (g1294) & (g1295) & (g1296) & (g147) & (!g148)) + ((g1293) & (g1294) & (g1295) & (g1296) & (g147) & (g148)));
	assign g1298 = (((!g1282) & (!g1287) & (!g1292) & (g1297) & (g165) & (g166)) + ((!g1282) & (!g1287) & (g1292) & (!g1297) & (!g165) & (g166)) + ((!g1282) & (!g1287) & (g1292) & (g1297) & (!g165) & (g166)) + ((!g1282) & (!g1287) & (g1292) & (g1297) & (g165) & (g166)) + ((!g1282) & (g1287) & (!g1292) & (!g1297) & (g165) & (!g166)) + ((!g1282) & (g1287) & (!g1292) & (g1297) & (g165) & (!g166)) + ((!g1282) & (g1287) & (!g1292) & (g1297) & (g165) & (g166)) + ((!g1282) & (g1287) & (g1292) & (!g1297) & (!g165) & (g166)) + ((!g1282) & (g1287) & (g1292) & (!g1297) & (g165) & (!g166)) + ((!g1282) & (g1287) & (g1292) & (g1297) & (!g165) & (g166)) + ((!g1282) & (g1287) & (g1292) & (g1297) & (g165) & (!g166)) + ((!g1282) & (g1287) & (g1292) & (g1297) & (g165) & (g166)) + ((g1282) & (!g1287) & (!g1292) & (!g1297) & (!g165) & (!g166)) + ((g1282) & (!g1287) & (!g1292) & (g1297) & (!g165) & (!g166)) + ((g1282) & (!g1287) & (!g1292) & (g1297) & (g165) & (g166)) + ((g1282) & (!g1287) & (g1292) & (!g1297) & (!g165) & (!g166)) + ((g1282) & (!g1287) & (g1292) & (!g1297) & (!g165) & (g166)) + ((g1282) & (!g1287) & (g1292) & (g1297) & (!g165) & (!g166)) + ((g1282) & (!g1287) & (g1292) & (g1297) & (!g165) & (g166)) + ((g1282) & (!g1287) & (g1292) & (g1297) & (g165) & (g166)) + ((g1282) & (g1287) & (!g1292) & (!g1297) & (!g165) & (!g166)) + ((g1282) & (g1287) & (!g1292) & (!g1297) & (g165) & (!g166)) + ((g1282) & (g1287) & (!g1292) & (g1297) & (!g165) & (!g166)) + ((g1282) & (g1287) & (!g1292) & (g1297) & (g165) & (!g166)) + ((g1282) & (g1287) & (!g1292) & (g1297) & (g165) & (g166)) + ((g1282) & (g1287) & (g1292) & (!g1297) & (!g165) & (!g166)) + ((g1282) & (g1287) & (g1292) & (!g1297) & (!g165) & (g166)) + ((g1282) & (g1287) & (g1292) & (!g1297) & (g165) & (!g166)) + ((g1282) & (g1287) & (g1292) & (g1297) & (!g165) & (!g166)) + ((g1282) & (g1287) & (g1292) & (g1297) & (!g165) & (g166)) + ((g1282) & (g1287) & (g1292) & (g1297) & (g165) & (!g166)) + ((g1282) & (g1287) & (g1292) & (g1297) & (g165) & (g166)));
	assign g4810 = (((!g2173) & (!sk[85]) & (!g3325) & (g1299)) + ((!g2173) & (!sk[85]) & (g3325) & (!g1299)) + ((!g2173) & (!sk[85]) & (g3325) & (g1299)) + ((!g2173) & (sk[85]) & (!g3325) & (g1299)) + ((!g2173) & (sk[85]) & (g3325) & (g1299)) + ((g2173) & (!sk[85]) & (!g3325) & (g1299)) + ((g2173) & (!sk[85]) & (g3325) & (!g1299)) + ((g2173) & (!sk[85]) & (g3325) & (g1299)) + ((g2173) & (sk[85]) & (g3325) & (!g1299)) + ((g2173) & (sk[85]) & (g3325) & (g1299)));
	assign g4811 = (((!g2174) & (!g3325) & (!sk[86]) & (g1300)) + ((!g2174) & (!g3325) & (sk[86]) & (g1300)) + ((!g2174) & (g3325) & (!sk[86]) & (!g1300)) + ((!g2174) & (g3325) & (!sk[86]) & (g1300)) + ((!g2174) & (g3325) & (sk[86]) & (g1300)) + ((g2174) & (!g3325) & (!sk[86]) & (g1300)) + ((g2174) & (g3325) & (!sk[86]) & (!g1300)) + ((g2174) & (g3325) & (!sk[86]) & (g1300)) + ((g2174) & (g3325) & (sk[86]) & (!g1300)) + ((g2174) & (g3325) & (sk[86]) & (g1300)));
	assign g4812 = (((!g2175) & (!g3325) & (!sk[87]) & (g1301)) + ((!g2175) & (!g3325) & (sk[87]) & (g1301)) + ((!g2175) & (g3325) & (!sk[87]) & (!g1301)) + ((!g2175) & (g3325) & (!sk[87]) & (g1301)) + ((!g2175) & (g3325) & (sk[87]) & (g1301)) + ((g2175) & (!g3325) & (!sk[87]) & (g1301)) + ((g2175) & (g3325) & (!sk[87]) & (!g1301)) + ((g2175) & (g3325) & (!sk[87]) & (g1301)) + ((g2175) & (g3325) & (sk[87]) & (!g1301)) + ((g2175) & (g3325) & (sk[87]) & (g1301)));
	assign g4813 = (((!g2176) & (!sk[88]) & (!g3325) & (g1302)) + ((!g2176) & (!sk[88]) & (g3325) & (!g1302)) + ((!g2176) & (!sk[88]) & (g3325) & (g1302)) + ((!g2176) & (sk[88]) & (!g3325) & (g1302)) + ((!g2176) & (sk[88]) & (g3325) & (g1302)) + ((g2176) & (!sk[88]) & (!g3325) & (g1302)) + ((g2176) & (!sk[88]) & (g3325) & (!g1302)) + ((g2176) & (!sk[88]) & (g3325) & (g1302)) + ((g2176) & (sk[88]) & (g3325) & (!g1302)) + ((g2176) & (sk[88]) & (g3325) & (g1302)));
	assign g1303 = (((!g1299) & (!g1300) & (!g1301) & (g1302) & (g165) & (g166)) + ((!g1299) & (!g1300) & (g1301) & (!g1302) & (!g165) & (g166)) + ((!g1299) & (!g1300) & (g1301) & (g1302) & (!g165) & (g166)) + ((!g1299) & (!g1300) & (g1301) & (g1302) & (g165) & (g166)) + ((!g1299) & (g1300) & (!g1301) & (!g1302) & (g165) & (!g166)) + ((!g1299) & (g1300) & (!g1301) & (g1302) & (g165) & (!g166)) + ((!g1299) & (g1300) & (!g1301) & (g1302) & (g165) & (g166)) + ((!g1299) & (g1300) & (g1301) & (!g1302) & (!g165) & (g166)) + ((!g1299) & (g1300) & (g1301) & (!g1302) & (g165) & (!g166)) + ((!g1299) & (g1300) & (g1301) & (g1302) & (!g165) & (g166)) + ((!g1299) & (g1300) & (g1301) & (g1302) & (g165) & (!g166)) + ((!g1299) & (g1300) & (g1301) & (g1302) & (g165) & (g166)) + ((g1299) & (!g1300) & (!g1301) & (!g1302) & (!g165) & (!g166)) + ((g1299) & (!g1300) & (!g1301) & (g1302) & (!g165) & (!g166)) + ((g1299) & (!g1300) & (!g1301) & (g1302) & (g165) & (g166)) + ((g1299) & (!g1300) & (g1301) & (!g1302) & (!g165) & (!g166)) + ((g1299) & (!g1300) & (g1301) & (!g1302) & (!g165) & (g166)) + ((g1299) & (!g1300) & (g1301) & (g1302) & (!g165) & (!g166)) + ((g1299) & (!g1300) & (g1301) & (g1302) & (!g165) & (g166)) + ((g1299) & (!g1300) & (g1301) & (g1302) & (g165) & (g166)) + ((g1299) & (g1300) & (!g1301) & (!g1302) & (!g165) & (!g166)) + ((g1299) & (g1300) & (!g1301) & (!g1302) & (g165) & (!g166)) + ((g1299) & (g1300) & (!g1301) & (g1302) & (!g165) & (!g166)) + ((g1299) & (g1300) & (!g1301) & (g1302) & (g165) & (!g166)) + ((g1299) & (g1300) & (!g1301) & (g1302) & (g165) & (g166)) + ((g1299) & (g1300) & (g1301) & (!g1302) & (!g165) & (!g166)) + ((g1299) & (g1300) & (g1301) & (!g1302) & (!g165) & (g166)) + ((g1299) & (g1300) & (g1301) & (!g1302) & (g165) & (!g166)) + ((g1299) & (g1300) & (g1301) & (g1302) & (!g165) & (!g166)) + ((g1299) & (g1300) & (g1301) & (g1302) & (!g165) & (g166)) + ((g1299) & (g1300) & (g1301) & (g1302) & (g165) & (!g166)) + ((g1299) & (g1300) & (g1301) & (g1302) & (g165) & (g166)));
	assign g4814 = (((!g2177) & (!g3325) & (!sk[90]) & (g1304)) + ((!g2177) & (!g3325) & (sk[90]) & (g1304)) + ((!g2177) & (g3325) & (!sk[90]) & (!g1304)) + ((!g2177) & (g3325) & (!sk[90]) & (g1304)) + ((!g2177) & (g3325) & (sk[90]) & (g1304)) + ((g2177) & (!g3325) & (!sk[90]) & (g1304)) + ((g2177) & (g3325) & (!sk[90]) & (!g1304)) + ((g2177) & (g3325) & (!sk[90]) & (g1304)) + ((g2177) & (g3325) & (sk[90]) & (!g1304)) + ((g2177) & (g3325) & (sk[90]) & (g1304)));
	assign g4815 = (((!g2178) & (!g3325) & (!sk[91]) & (g1305)) + ((!g2178) & (!g3325) & (sk[91]) & (g1305)) + ((!g2178) & (g3325) & (!sk[91]) & (!g1305)) + ((!g2178) & (g3325) & (!sk[91]) & (g1305)) + ((!g2178) & (g3325) & (sk[91]) & (g1305)) + ((g2178) & (!g3325) & (!sk[91]) & (g1305)) + ((g2178) & (g3325) & (!sk[91]) & (!g1305)) + ((g2178) & (g3325) & (!sk[91]) & (g1305)) + ((g2178) & (g3325) & (sk[91]) & (!g1305)) + ((g2178) & (g3325) & (sk[91]) & (g1305)));
	assign g4816 = (((!g2179) & (!sk[92]) & (!g3325) & (g1306)) + ((!g2179) & (!sk[92]) & (g3325) & (!g1306)) + ((!g2179) & (!sk[92]) & (g3325) & (g1306)) + ((!g2179) & (sk[92]) & (!g3325) & (g1306)) + ((!g2179) & (sk[92]) & (g3325) & (g1306)) + ((g2179) & (!sk[92]) & (!g3325) & (g1306)) + ((g2179) & (!sk[92]) & (g3325) & (!g1306)) + ((g2179) & (!sk[92]) & (g3325) & (g1306)) + ((g2179) & (sk[92]) & (g3325) & (!g1306)) + ((g2179) & (sk[92]) & (g3325) & (g1306)));
	assign g1307 = (((!g165) & (!g166) & (!sk[93]) & (!g1304) & (g1305) & (!g1306)) + ((!g165) & (!g166) & (!sk[93]) & (!g1304) & (g1305) & (g1306)) + ((!g165) & (!g166) & (!sk[93]) & (g1304) & (!g1305) & (!g1306)) + ((!g165) & (!g166) & (!sk[93]) & (g1304) & (!g1305) & (g1306)) + ((!g165) & (!g166) & (!sk[93]) & (g1304) & (g1305) & (!g1306)) + ((!g165) & (!g166) & (!sk[93]) & (g1304) & (g1305) & (g1306)) + ((!g165) & (g166) & (!sk[93]) & (!g1304) & (!g1305) & (!g1306)) + ((!g165) & (g166) & (!sk[93]) & (!g1304) & (!g1305) & (g1306)) + ((!g165) & (g166) & (!sk[93]) & (!g1304) & (g1305) & (!g1306)) + ((!g165) & (g166) & (!sk[93]) & (!g1304) & (g1305) & (g1306)) + ((!g165) & (g166) & (!sk[93]) & (g1304) & (!g1305) & (!g1306)) + ((!g165) & (g166) & (!sk[93]) & (g1304) & (!g1305) & (g1306)) + ((!g165) & (g166) & (!sk[93]) & (g1304) & (g1305) & (!g1306)) + ((!g165) & (g166) & (!sk[93]) & (g1304) & (g1305) & (g1306)) + ((!g165) & (g166) & (sk[93]) & (!g1304) & (!g1305) & (g1306)) + ((!g165) & (g166) & (sk[93]) & (!g1304) & (g1305) & (g1306)) + ((!g165) & (g166) & (sk[93]) & (g1304) & (!g1305) & (g1306)) + ((!g165) & (g166) & (sk[93]) & (g1304) & (g1305) & (g1306)) + ((g165) & (!g166) & (!sk[93]) & (!g1304) & (g1305) & (!g1306)) + ((g165) & (!g166) & (!sk[93]) & (!g1304) & (g1305) & (g1306)) + ((g165) & (!g166) & (!sk[93]) & (g1304) & (!g1305) & (!g1306)) + ((g165) & (!g166) & (!sk[93]) & (g1304) & (!g1305) & (g1306)) + ((g165) & (!g166) & (!sk[93]) & (g1304) & (g1305) & (!g1306)) + ((g165) & (!g166) & (!sk[93]) & (g1304) & (g1305) & (g1306)) + ((g165) & (!g166) & (sk[93]) & (g1304) & (!g1305) & (!g1306)) + ((g165) & (!g166) & (sk[93]) & (g1304) & (!g1305) & (g1306)) + ((g165) & (!g166) & (sk[93]) & (g1304) & (g1305) & (!g1306)) + ((g165) & (!g166) & (sk[93]) & (g1304) & (g1305) & (g1306)) + ((g165) & (g166) & (!sk[93]) & (!g1304) & (!g1305) & (!g1306)) + ((g165) & (g166) & (!sk[93]) & (!g1304) & (!g1305) & (g1306)) + ((g165) & (g166) & (!sk[93]) & (!g1304) & (g1305) & (!g1306)) + ((g165) & (g166) & (!sk[93]) & (!g1304) & (g1305) & (g1306)) + ((g165) & (g166) & (!sk[93]) & (g1304) & (!g1305) & (!g1306)) + ((g165) & (g166) & (!sk[93]) & (g1304) & (!g1305) & (g1306)) + ((g165) & (g166) & (!sk[93]) & (g1304) & (g1305) & (!g1306)) + ((g165) & (g166) & (!sk[93]) & (g1304) & (g1305) & (g1306)) + ((g165) & (g166) & (sk[93]) & (!g1304) & (g1305) & (!g1306)) + ((g165) & (g166) & (sk[93]) & (!g1304) & (g1305) & (g1306)) + ((g165) & (g166) & (sk[93]) & (g1304) & (g1305) & (!g1306)) + ((g165) & (g166) & (sk[93]) & (g1304) & (g1305) & (g1306)));
	assign g4817 = (((!g2162) & (!sk[94]) & (!g3325) & (g1308)) + ((!g2162) & (!sk[94]) & (g3325) & (!g1308)) + ((!g2162) & (!sk[94]) & (g3325) & (g1308)) + ((!g2162) & (sk[94]) & (!g3325) & (g1308)) + ((!g2162) & (sk[94]) & (g3325) & (g1308)) + ((g2162) & (!sk[94]) & (!g3325) & (g1308)) + ((g2162) & (!sk[94]) & (g3325) & (!g1308)) + ((g2162) & (!sk[94]) & (g3325) & (g1308)) + ((g2162) & (sk[94]) & (g3325) & (!g1308)) + ((g2162) & (sk[94]) & (g3325) & (g1308)));
	assign g4818 = (((!sk[95]) & (!g2164) & (!g3325) & (g1309)) + ((!sk[95]) & (!g2164) & (g3325) & (!g1309)) + ((!sk[95]) & (!g2164) & (g3325) & (g1309)) + ((!sk[95]) & (g2164) & (!g3325) & (g1309)) + ((!sk[95]) & (g2164) & (g3325) & (!g1309)) + ((!sk[95]) & (g2164) & (g3325) & (g1309)) + ((sk[95]) & (!g2164) & (!g3325) & (g1309)) + ((sk[95]) & (!g2164) & (g3325) & (g1309)) + ((sk[95]) & (g2164) & (g3325) & (!g1309)) + ((sk[95]) & (g2164) & (g3325) & (g1309)));
	assign g4819 = (((!g2166) & (!sk[96]) & (!g3325) & (g1310)) + ((!g2166) & (!sk[96]) & (g3325) & (!g1310)) + ((!g2166) & (!sk[96]) & (g3325) & (g1310)) + ((!g2166) & (sk[96]) & (!g3325) & (g1310)) + ((!g2166) & (sk[96]) & (g3325) & (g1310)) + ((g2166) & (!sk[96]) & (!g3325) & (g1310)) + ((g2166) & (!sk[96]) & (g3325) & (!g1310)) + ((g2166) & (!sk[96]) & (g3325) & (g1310)) + ((g2166) & (sk[96]) & (g3325) & (!g1310)) + ((g2166) & (sk[96]) & (g3325) & (g1310)));
	assign g4820 = (((!sk[97]) & (!g2168) & (!g3325) & (g1311)) + ((!sk[97]) & (!g2168) & (g3325) & (!g1311)) + ((!sk[97]) & (!g2168) & (g3325) & (g1311)) + ((!sk[97]) & (g2168) & (!g3325) & (g1311)) + ((!sk[97]) & (g2168) & (g3325) & (!g1311)) + ((!sk[97]) & (g2168) & (g3325) & (g1311)) + ((sk[97]) & (!g2168) & (!g3325) & (g1311)) + ((sk[97]) & (!g2168) & (g3325) & (g1311)) + ((sk[97]) & (g2168) & (g3325) & (!g1311)) + ((sk[97]) & (g2168) & (g3325) & (g1311)));
	assign g1312 = (((!g1308) & (!g1309) & (!g1310) & (g1311) & (g165) & (g166)) + ((!g1308) & (!g1309) & (g1310) & (!g1311) & (!g165) & (g166)) + ((!g1308) & (!g1309) & (g1310) & (g1311) & (!g165) & (g166)) + ((!g1308) & (!g1309) & (g1310) & (g1311) & (g165) & (g166)) + ((!g1308) & (g1309) & (!g1310) & (!g1311) & (g165) & (!g166)) + ((!g1308) & (g1309) & (!g1310) & (g1311) & (g165) & (!g166)) + ((!g1308) & (g1309) & (!g1310) & (g1311) & (g165) & (g166)) + ((!g1308) & (g1309) & (g1310) & (!g1311) & (!g165) & (g166)) + ((!g1308) & (g1309) & (g1310) & (!g1311) & (g165) & (!g166)) + ((!g1308) & (g1309) & (g1310) & (g1311) & (!g165) & (g166)) + ((!g1308) & (g1309) & (g1310) & (g1311) & (g165) & (!g166)) + ((!g1308) & (g1309) & (g1310) & (g1311) & (g165) & (g166)) + ((g1308) & (!g1309) & (!g1310) & (!g1311) & (!g165) & (!g166)) + ((g1308) & (!g1309) & (!g1310) & (g1311) & (!g165) & (!g166)) + ((g1308) & (!g1309) & (!g1310) & (g1311) & (g165) & (g166)) + ((g1308) & (!g1309) & (g1310) & (!g1311) & (!g165) & (!g166)) + ((g1308) & (!g1309) & (g1310) & (!g1311) & (!g165) & (g166)) + ((g1308) & (!g1309) & (g1310) & (g1311) & (!g165) & (!g166)) + ((g1308) & (!g1309) & (g1310) & (g1311) & (!g165) & (g166)) + ((g1308) & (!g1309) & (g1310) & (g1311) & (g165) & (g166)) + ((g1308) & (g1309) & (!g1310) & (!g1311) & (!g165) & (!g166)) + ((g1308) & (g1309) & (!g1310) & (!g1311) & (g165) & (!g166)) + ((g1308) & (g1309) & (!g1310) & (g1311) & (!g165) & (!g166)) + ((g1308) & (g1309) & (!g1310) & (g1311) & (g165) & (!g166)) + ((g1308) & (g1309) & (!g1310) & (g1311) & (g165) & (g166)) + ((g1308) & (g1309) & (g1310) & (!g1311) & (!g165) & (!g166)) + ((g1308) & (g1309) & (g1310) & (!g1311) & (!g165) & (g166)) + ((g1308) & (g1309) & (g1310) & (!g1311) & (g165) & (!g166)) + ((g1308) & (g1309) & (g1310) & (g1311) & (!g165) & (!g166)) + ((g1308) & (g1309) & (g1310) & (g1311) & (!g165) & (g166)) + ((g1308) & (g1309) & (g1310) & (g1311) & (g165) & (!g166)) + ((g1308) & (g1309) & (g1310) & (g1311) & (g165) & (g166)));
	assign g4821 = (((!g2169) & (!sk[99]) & (!g3325) & (g1313)) + ((!g2169) & (!sk[99]) & (g3325) & (!g1313)) + ((!g2169) & (!sk[99]) & (g3325) & (g1313)) + ((!g2169) & (sk[99]) & (!g3325) & (g1313)) + ((!g2169) & (sk[99]) & (g3325) & (g1313)) + ((g2169) & (!sk[99]) & (!g3325) & (g1313)) + ((g2169) & (!sk[99]) & (g3325) & (!g1313)) + ((g2169) & (!sk[99]) & (g3325) & (g1313)) + ((g2169) & (sk[99]) & (g3325) & (!g1313)) + ((g2169) & (sk[99]) & (g3325) & (g1313)));
	assign g4822 = (((!sk[100]) & (!g2170) & (!g3325) & (g1314)) + ((!sk[100]) & (!g2170) & (g3325) & (!g1314)) + ((!sk[100]) & (!g2170) & (g3325) & (g1314)) + ((!sk[100]) & (g2170) & (!g3325) & (g1314)) + ((!sk[100]) & (g2170) & (g3325) & (!g1314)) + ((!sk[100]) & (g2170) & (g3325) & (g1314)) + ((sk[100]) & (!g2170) & (!g3325) & (g1314)) + ((sk[100]) & (!g2170) & (g3325) & (g1314)) + ((sk[100]) & (g2170) & (g3325) & (!g1314)) + ((sk[100]) & (g2170) & (g3325) & (g1314)));
	assign g4823 = (((!g2171) & (!sk[101]) & (!g3325) & (g1315)) + ((!g2171) & (!sk[101]) & (g3325) & (!g1315)) + ((!g2171) & (!sk[101]) & (g3325) & (g1315)) + ((!g2171) & (sk[101]) & (!g3325) & (g1315)) + ((!g2171) & (sk[101]) & (g3325) & (g1315)) + ((g2171) & (!sk[101]) & (!g3325) & (g1315)) + ((g2171) & (!sk[101]) & (g3325) & (!g1315)) + ((g2171) & (!sk[101]) & (g3325) & (g1315)) + ((g2171) & (sk[101]) & (g3325) & (!g1315)) + ((g2171) & (sk[101]) & (g3325) & (g1315)));
	assign g4824 = (((!sk[102]) & (!g2172) & (!g3325) & (g1316)) + ((!sk[102]) & (!g2172) & (g3325) & (!g1316)) + ((!sk[102]) & (!g2172) & (g3325) & (g1316)) + ((!sk[102]) & (g2172) & (!g3325) & (g1316)) + ((!sk[102]) & (g2172) & (g3325) & (!g1316)) + ((!sk[102]) & (g2172) & (g3325) & (g1316)) + ((sk[102]) & (!g2172) & (!g3325) & (g1316)) + ((sk[102]) & (!g2172) & (g3325) & (g1316)) + ((sk[102]) & (g2172) & (g3325) & (!g1316)) + ((sk[102]) & (g2172) & (g3325) & (g1316)));
	assign g1317 = (((!g1313) & (!g1314) & (!g1315) & (g1316) & (g165) & (g166)) + ((!g1313) & (!g1314) & (g1315) & (!g1316) & (!g165) & (g166)) + ((!g1313) & (!g1314) & (g1315) & (g1316) & (!g165) & (g166)) + ((!g1313) & (!g1314) & (g1315) & (g1316) & (g165) & (g166)) + ((!g1313) & (g1314) & (!g1315) & (!g1316) & (g165) & (!g166)) + ((!g1313) & (g1314) & (!g1315) & (g1316) & (g165) & (!g166)) + ((!g1313) & (g1314) & (!g1315) & (g1316) & (g165) & (g166)) + ((!g1313) & (g1314) & (g1315) & (!g1316) & (!g165) & (g166)) + ((!g1313) & (g1314) & (g1315) & (!g1316) & (g165) & (!g166)) + ((!g1313) & (g1314) & (g1315) & (g1316) & (!g165) & (g166)) + ((!g1313) & (g1314) & (g1315) & (g1316) & (g165) & (!g166)) + ((!g1313) & (g1314) & (g1315) & (g1316) & (g165) & (g166)) + ((g1313) & (!g1314) & (!g1315) & (!g1316) & (!g165) & (!g166)) + ((g1313) & (!g1314) & (!g1315) & (g1316) & (!g165) & (!g166)) + ((g1313) & (!g1314) & (!g1315) & (g1316) & (g165) & (g166)) + ((g1313) & (!g1314) & (g1315) & (!g1316) & (!g165) & (!g166)) + ((g1313) & (!g1314) & (g1315) & (!g1316) & (!g165) & (g166)) + ((g1313) & (!g1314) & (g1315) & (g1316) & (!g165) & (!g166)) + ((g1313) & (!g1314) & (g1315) & (g1316) & (!g165) & (g166)) + ((g1313) & (!g1314) & (g1315) & (g1316) & (g165) & (g166)) + ((g1313) & (g1314) & (!g1315) & (!g1316) & (!g165) & (!g166)) + ((g1313) & (g1314) & (!g1315) & (!g1316) & (g165) & (!g166)) + ((g1313) & (g1314) & (!g1315) & (g1316) & (!g165) & (!g166)) + ((g1313) & (g1314) & (!g1315) & (g1316) & (g165) & (!g166)) + ((g1313) & (g1314) & (!g1315) & (g1316) & (g165) & (g166)) + ((g1313) & (g1314) & (g1315) & (!g1316) & (!g165) & (!g166)) + ((g1313) & (g1314) & (g1315) & (!g1316) & (!g165) & (g166)) + ((g1313) & (g1314) & (g1315) & (!g1316) & (g165) & (!g166)) + ((g1313) & (g1314) & (g1315) & (g1316) & (!g165) & (!g166)) + ((g1313) & (g1314) & (g1315) & (g1316) & (!g165) & (g166)) + ((g1313) & (g1314) & (g1315) & (g1316) & (g165) & (!g166)) + ((g1313) & (g1314) & (g1315) & (g1316) & (g165) & (g166)));
	assign g1318 = (((!g147) & (!g148) & (!g1303) & (g1307) & (!g1312) & (!g1317)) + ((!g147) & (!g148) & (!g1303) & (g1307) & (!g1312) & (g1317)) + ((!g147) & (!g148) & (!g1303) & (g1307) & (g1312) & (!g1317)) + ((!g147) & (!g148) & (!g1303) & (g1307) & (g1312) & (g1317)) + ((!g147) & (!g148) & (g1303) & (g1307) & (!g1312) & (!g1317)) + ((!g147) & (!g148) & (g1303) & (g1307) & (!g1312) & (g1317)) + ((!g147) & (!g148) & (g1303) & (g1307) & (g1312) & (!g1317)) + ((!g147) & (!g148) & (g1303) & (g1307) & (g1312) & (g1317)) + ((!g147) & (g148) & (!g1303) & (!g1307) & (!g1312) & (g1317)) + ((!g147) & (g148) & (!g1303) & (!g1307) & (g1312) & (g1317)) + ((!g147) & (g148) & (!g1303) & (g1307) & (!g1312) & (g1317)) + ((!g147) & (g148) & (!g1303) & (g1307) & (g1312) & (g1317)) + ((!g147) & (g148) & (g1303) & (!g1307) & (!g1312) & (g1317)) + ((!g147) & (g148) & (g1303) & (!g1307) & (g1312) & (g1317)) + ((!g147) & (g148) & (g1303) & (g1307) & (!g1312) & (g1317)) + ((!g147) & (g148) & (g1303) & (g1307) & (g1312) & (g1317)) + ((g147) & (!g148) & (g1303) & (!g1307) & (!g1312) & (!g1317)) + ((g147) & (!g148) & (g1303) & (!g1307) & (!g1312) & (g1317)) + ((g147) & (!g148) & (g1303) & (!g1307) & (g1312) & (!g1317)) + ((g147) & (!g148) & (g1303) & (!g1307) & (g1312) & (g1317)) + ((g147) & (!g148) & (g1303) & (g1307) & (!g1312) & (!g1317)) + ((g147) & (!g148) & (g1303) & (g1307) & (!g1312) & (g1317)) + ((g147) & (!g148) & (g1303) & (g1307) & (g1312) & (!g1317)) + ((g147) & (!g148) & (g1303) & (g1307) & (g1312) & (g1317)) + ((g147) & (g148) & (!g1303) & (!g1307) & (g1312) & (!g1317)) + ((g147) & (g148) & (!g1303) & (!g1307) & (g1312) & (g1317)) + ((g147) & (g148) & (!g1303) & (g1307) & (g1312) & (!g1317)) + ((g147) & (g148) & (!g1303) & (g1307) & (g1312) & (g1317)) + ((g147) & (g148) & (g1303) & (!g1307) & (g1312) & (!g1317)) + ((g147) & (g148) & (g1303) & (!g1307) & (g1312) & (g1317)) + ((g147) & (g148) & (g1303) & (g1307) & (g1312) & (!g1317)) + ((g147) & (g148) & (g1303) & (g1307) & (g1312) & (g1317)));
	assign g1319 = (((!g142) & (!sk[105]) & (!g1298) & (g1318)) + ((!g142) & (!sk[105]) & (g1298) & (!g1318)) + ((!g142) & (!sk[105]) & (g1298) & (g1318)) + ((!g142) & (sk[105]) & (!g1298) & (g1318)) + ((!g142) & (sk[105]) & (g1298) & (g1318)) + ((g142) & (!sk[105]) & (!g1298) & (g1318)) + ((g142) & (!sk[105]) & (g1298) & (!g1318)) + ((g142) & (!sk[105]) & (g1298) & (g1318)) + ((g142) & (sk[105]) & (g1298) & (!g1318)) + ((g142) & (sk[105]) & (g1298) & (g1318)));
	assign g4825 = (((!g2059) & (!g2733) & (!sk[106]) & (g1320)) + ((!g2059) & (!g2733) & (sk[106]) & (g1320)) + ((!g2059) & (g2733) & (!sk[106]) & (!g1320)) + ((!g2059) & (g2733) & (!sk[106]) & (g1320)) + ((!g2059) & (g2733) & (sk[106]) & (g1320)) + ((g2059) & (!g2733) & (!sk[106]) & (g1320)) + ((g2059) & (g2733) & (!sk[106]) & (!g1320)) + ((g2059) & (g2733) & (!sk[106]) & (g1320)) + ((g2059) & (g2733) & (sk[106]) & (!g1320)) + ((g2059) & (g2733) & (sk[106]) & (g1320)));
	assign g1321 = (((!g1274) & (!g1276) & (!sk[107]) & (g916)) + ((!g1274) & (g1276) & (!sk[107]) & (!g916)) + ((!g1274) & (g1276) & (!sk[107]) & (g916)) + ((!g1274) & (g1276) & (sk[107]) & (!g916)) + ((g1274) & (!g1276) & (!sk[107]) & (g916)) + ((g1274) & (!g1276) & (sk[107]) & (!g916)) + ((g1274) & (g1276) & (!sk[107]) & (!g916)) + ((g1274) & (g1276) & (!sk[107]) & (g916)) + ((g1274) & (g1276) & (sk[107]) & (!g916)) + ((g1274) & (g1276) & (sk[107]) & (g916)));
	assign g1322 = (((!g126) & (!g1319) & (!sk[108]) & (!g1320) & (g1321) & (!g916)) + ((!g126) & (!g1319) & (!sk[108]) & (!g1320) & (g1321) & (g916)) + ((!g126) & (!g1319) & (!sk[108]) & (g1320) & (!g1321) & (!g916)) + ((!g126) & (!g1319) & (!sk[108]) & (g1320) & (!g1321) & (g916)) + ((!g126) & (!g1319) & (!sk[108]) & (g1320) & (g1321) & (!g916)) + ((!g126) & (!g1319) & (!sk[108]) & (g1320) & (g1321) & (g916)) + ((!g126) & (!g1319) & (sk[108]) & (g1320) & (!g1321) & (!g916)) + ((!g126) & (!g1319) & (sk[108]) & (g1320) & (!g1321) & (g916)) + ((!g126) & (!g1319) & (sk[108]) & (g1320) & (g1321) & (!g916)) + ((!g126) & (!g1319) & (sk[108]) & (g1320) & (g1321) & (g916)) + ((!g126) & (g1319) & (!sk[108]) & (!g1320) & (!g1321) & (!g916)) + ((!g126) & (g1319) & (!sk[108]) & (!g1320) & (!g1321) & (g916)) + ((!g126) & (g1319) & (!sk[108]) & (!g1320) & (g1321) & (!g916)) + ((!g126) & (g1319) & (!sk[108]) & (!g1320) & (g1321) & (g916)) + ((!g126) & (g1319) & (!sk[108]) & (g1320) & (!g1321) & (!g916)) + ((!g126) & (g1319) & (!sk[108]) & (g1320) & (!g1321) & (g916)) + ((!g126) & (g1319) & (!sk[108]) & (g1320) & (g1321) & (!g916)) + ((!g126) & (g1319) & (!sk[108]) & (g1320) & (g1321) & (g916)) + ((!g126) & (g1319) & (sk[108]) & (g1320) & (!g1321) & (!g916)) + ((!g126) & (g1319) & (sk[108]) & (g1320) & (!g1321) & (g916)) + ((!g126) & (g1319) & (sk[108]) & (g1320) & (g1321) & (!g916)) + ((!g126) & (g1319) & (sk[108]) & (g1320) & (g1321) & (g916)) + ((g126) & (!g1319) & (!sk[108]) & (!g1320) & (g1321) & (!g916)) + ((g126) & (!g1319) & (!sk[108]) & (!g1320) & (g1321) & (g916)) + ((g126) & (!g1319) & (!sk[108]) & (g1320) & (!g1321) & (!g916)) + ((g126) & (!g1319) & (!sk[108]) & (g1320) & (!g1321) & (g916)) + ((g126) & (!g1319) & (!sk[108]) & (g1320) & (g1321) & (!g916)) + ((g126) & (!g1319) & (!sk[108]) & (g1320) & (g1321) & (g916)) + ((g126) & (!g1319) & (sk[108]) & (!g1320) & (!g1321) & (!g916)) + ((g126) & (!g1319) & (sk[108]) & (!g1320) & (g1321) & (g916)) + ((g126) & (!g1319) & (sk[108]) & (g1320) & (!g1321) & (!g916)) + ((g126) & (!g1319) & (sk[108]) & (g1320) & (g1321) & (g916)) + ((g126) & (g1319) & (!sk[108]) & (!g1320) & (!g1321) & (!g916)) + ((g126) & (g1319) & (!sk[108]) & (!g1320) & (!g1321) & (g916)) + ((g126) & (g1319) & (!sk[108]) & (!g1320) & (g1321) & (!g916)) + ((g126) & (g1319) & (!sk[108]) & (!g1320) & (g1321) & (g916)) + ((g126) & (g1319) & (!sk[108]) & (g1320) & (!g1321) & (!g916)) + ((g126) & (g1319) & (!sk[108]) & (g1320) & (!g1321) & (g916)) + ((g126) & (g1319) & (!sk[108]) & (g1320) & (g1321) & (!g916)) + ((g126) & (g1319) & (!sk[108]) & (g1320) & (g1321) & (g916)) + ((g126) & (g1319) & (sk[108]) & (!g1320) & (!g1321) & (g916)) + ((g126) & (g1319) & (sk[108]) & (!g1320) & (g1321) & (!g916)) + ((g126) & (g1319) & (sk[108]) & (g1320) & (!g1321) & (g916)) + ((g126) & (g1319) & (sk[108]) & (g1320) & (g1321) & (!g916)));
	assign g4826 = (((!sk[109]) & (!g2140) & (!g3302) & (g1323)) + ((!sk[109]) & (!g2140) & (g3302) & (!g1323)) + ((!sk[109]) & (!g2140) & (g3302) & (g1323)) + ((!sk[109]) & (g2140) & (!g3302) & (g1323)) + ((!sk[109]) & (g2140) & (g3302) & (!g1323)) + ((!sk[109]) & (g2140) & (g3302) & (g1323)) + ((sk[109]) & (!g2140) & (!g3302) & (g1323)) + ((sk[109]) & (!g2140) & (g3302) & (g1323)) + ((sk[109]) & (g2140) & (g3302) & (!g1323)) + ((sk[109]) & (g2140) & (g3302) & (g1323)));
	assign g4827 = (((!g2142) & (!g3302) & (!sk[110]) & (g1324)) + ((!g2142) & (!g3302) & (sk[110]) & (g1324)) + ((!g2142) & (g3302) & (!sk[110]) & (!g1324)) + ((!g2142) & (g3302) & (!sk[110]) & (g1324)) + ((!g2142) & (g3302) & (sk[110]) & (g1324)) + ((g2142) & (!g3302) & (!sk[110]) & (g1324)) + ((g2142) & (g3302) & (!sk[110]) & (!g1324)) + ((g2142) & (g3302) & (!sk[110]) & (g1324)) + ((g2142) & (g3302) & (sk[110]) & (!g1324)) + ((g2142) & (g3302) & (sk[110]) & (g1324)));
	assign g4828 = (((!g2144) & (!sk[111]) & (!g3302) & (g1325)) + ((!g2144) & (!sk[111]) & (g3302) & (!g1325)) + ((!g2144) & (!sk[111]) & (g3302) & (g1325)) + ((!g2144) & (sk[111]) & (!g3302) & (g1325)) + ((!g2144) & (sk[111]) & (g3302) & (g1325)) + ((g2144) & (!sk[111]) & (!g3302) & (g1325)) + ((g2144) & (!sk[111]) & (g3302) & (!g1325)) + ((g2144) & (!sk[111]) & (g3302) & (g1325)) + ((g2144) & (sk[111]) & (g3302) & (!g1325)) + ((g2144) & (sk[111]) & (g3302) & (g1325)));
	assign g4829 = (((!g2145) & (!sk[112]) & (!g3302) & (g1326)) + ((!g2145) & (!sk[112]) & (g3302) & (!g1326)) + ((!g2145) & (!sk[112]) & (g3302) & (g1326)) + ((!g2145) & (sk[112]) & (!g3302) & (g1326)) + ((!g2145) & (sk[112]) & (g3302) & (g1326)) + ((g2145) & (!sk[112]) & (!g3302) & (g1326)) + ((g2145) & (!sk[112]) & (g3302) & (!g1326)) + ((g2145) & (!sk[112]) & (g3302) & (g1326)) + ((g2145) & (sk[112]) & (g3302) & (!g1326)) + ((g2145) & (sk[112]) & (g3302) & (g1326)));
	assign g1327 = (((!g1323) & (!g1324) & (!g1325) & (g1326) & (g147) & (g148)) + ((!g1323) & (!g1324) & (g1325) & (!g1326) & (!g147) & (g148)) + ((!g1323) & (!g1324) & (g1325) & (g1326) & (!g147) & (g148)) + ((!g1323) & (!g1324) & (g1325) & (g1326) & (g147) & (g148)) + ((!g1323) & (g1324) & (!g1325) & (!g1326) & (g147) & (!g148)) + ((!g1323) & (g1324) & (!g1325) & (g1326) & (g147) & (!g148)) + ((!g1323) & (g1324) & (!g1325) & (g1326) & (g147) & (g148)) + ((!g1323) & (g1324) & (g1325) & (!g1326) & (!g147) & (g148)) + ((!g1323) & (g1324) & (g1325) & (!g1326) & (g147) & (!g148)) + ((!g1323) & (g1324) & (g1325) & (g1326) & (!g147) & (g148)) + ((!g1323) & (g1324) & (g1325) & (g1326) & (g147) & (!g148)) + ((!g1323) & (g1324) & (g1325) & (g1326) & (g147) & (g148)) + ((g1323) & (!g1324) & (!g1325) & (!g1326) & (!g147) & (!g148)) + ((g1323) & (!g1324) & (!g1325) & (g1326) & (!g147) & (!g148)) + ((g1323) & (!g1324) & (!g1325) & (g1326) & (g147) & (g148)) + ((g1323) & (!g1324) & (g1325) & (!g1326) & (!g147) & (!g148)) + ((g1323) & (!g1324) & (g1325) & (!g1326) & (!g147) & (g148)) + ((g1323) & (!g1324) & (g1325) & (g1326) & (!g147) & (!g148)) + ((g1323) & (!g1324) & (g1325) & (g1326) & (!g147) & (g148)) + ((g1323) & (!g1324) & (g1325) & (g1326) & (g147) & (g148)) + ((g1323) & (g1324) & (!g1325) & (!g1326) & (!g147) & (!g148)) + ((g1323) & (g1324) & (!g1325) & (!g1326) & (g147) & (!g148)) + ((g1323) & (g1324) & (!g1325) & (g1326) & (!g147) & (!g148)) + ((g1323) & (g1324) & (!g1325) & (g1326) & (g147) & (!g148)) + ((g1323) & (g1324) & (!g1325) & (g1326) & (g147) & (g148)) + ((g1323) & (g1324) & (g1325) & (!g1326) & (!g147) & (!g148)) + ((g1323) & (g1324) & (g1325) & (!g1326) & (!g147) & (g148)) + ((g1323) & (g1324) & (g1325) & (!g1326) & (g147) & (!g148)) + ((g1323) & (g1324) & (g1325) & (g1326) & (!g147) & (!g148)) + ((g1323) & (g1324) & (g1325) & (g1326) & (!g147) & (g148)) + ((g1323) & (g1324) & (g1325) & (g1326) & (g147) & (!g148)) + ((g1323) & (g1324) & (g1325) & (g1326) & (g147) & (g148)));
	assign g4830 = (((!sk[114]) & (!g2146) & (!g3302) & (g1328)) + ((!sk[114]) & (!g2146) & (g3302) & (!g1328)) + ((!sk[114]) & (!g2146) & (g3302) & (g1328)) + ((!sk[114]) & (g2146) & (!g3302) & (g1328)) + ((!sk[114]) & (g2146) & (g3302) & (!g1328)) + ((!sk[114]) & (g2146) & (g3302) & (g1328)) + ((sk[114]) & (!g2146) & (!g3302) & (g1328)) + ((sk[114]) & (!g2146) & (g3302) & (g1328)) + ((sk[114]) & (g2146) & (g3302) & (!g1328)) + ((sk[114]) & (g2146) & (g3302) & (g1328)));
	assign g4831 = (((!g2148) & (!sk[115]) & (!g3302) & (g1329)) + ((!g2148) & (!sk[115]) & (g3302) & (!g1329)) + ((!g2148) & (!sk[115]) & (g3302) & (g1329)) + ((!g2148) & (sk[115]) & (!g3302) & (g1329)) + ((!g2148) & (sk[115]) & (g3302) & (g1329)) + ((g2148) & (!sk[115]) & (!g3302) & (g1329)) + ((g2148) & (!sk[115]) & (g3302) & (!g1329)) + ((g2148) & (!sk[115]) & (g3302) & (g1329)) + ((g2148) & (sk[115]) & (g3302) & (!g1329)) + ((g2148) & (sk[115]) & (g3302) & (g1329)));
	assign g4832 = (((!g2150) & (!sk[116]) & (!g3302) & (g1330)) + ((!g2150) & (!sk[116]) & (g3302) & (!g1330)) + ((!g2150) & (!sk[116]) & (g3302) & (g1330)) + ((!g2150) & (sk[116]) & (!g3302) & (g1330)) + ((!g2150) & (sk[116]) & (g3302) & (g1330)) + ((g2150) & (!sk[116]) & (!g3302) & (g1330)) + ((g2150) & (!sk[116]) & (g3302) & (!g1330)) + ((g2150) & (!sk[116]) & (g3302) & (g1330)) + ((g2150) & (sk[116]) & (g3302) & (!g1330)) + ((g2150) & (sk[116]) & (g3302) & (g1330)));
	assign g4833 = (((!sk[117]) & (!g2151) & (!g3302) & (g1331)) + ((!sk[117]) & (!g2151) & (g3302) & (!g1331)) + ((!sk[117]) & (!g2151) & (g3302) & (g1331)) + ((!sk[117]) & (g2151) & (!g3302) & (g1331)) + ((!sk[117]) & (g2151) & (g3302) & (!g1331)) + ((!sk[117]) & (g2151) & (g3302) & (g1331)) + ((sk[117]) & (!g2151) & (!g3302) & (g1331)) + ((sk[117]) & (!g2151) & (g3302) & (g1331)) + ((sk[117]) & (g2151) & (g3302) & (!g1331)) + ((sk[117]) & (g2151) & (g3302) & (g1331)));
	assign g1332 = (((!g1328) & (!g1329) & (!g1330) & (g1331) & (g147) & (g148)) + ((!g1328) & (!g1329) & (g1330) & (!g1331) & (!g147) & (g148)) + ((!g1328) & (!g1329) & (g1330) & (g1331) & (!g147) & (g148)) + ((!g1328) & (!g1329) & (g1330) & (g1331) & (g147) & (g148)) + ((!g1328) & (g1329) & (!g1330) & (!g1331) & (g147) & (!g148)) + ((!g1328) & (g1329) & (!g1330) & (g1331) & (g147) & (!g148)) + ((!g1328) & (g1329) & (!g1330) & (g1331) & (g147) & (g148)) + ((!g1328) & (g1329) & (g1330) & (!g1331) & (!g147) & (g148)) + ((!g1328) & (g1329) & (g1330) & (!g1331) & (g147) & (!g148)) + ((!g1328) & (g1329) & (g1330) & (g1331) & (!g147) & (g148)) + ((!g1328) & (g1329) & (g1330) & (g1331) & (g147) & (!g148)) + ((!g1328) & (g1329) & (g1330) & (g1331) & (g147) & (g148)) + ((g1328) & (!g1329) & (!g1330) & (!g1331) & (!g147) & (!g148)) + ((g1328) & (!g1329) & (!g1330) & (g1331) & (!g147) & (!g148)) + ((g1328) & (!g1329) & (!g1330) & (g1331) & (g147) & (g148)) + ((g1328) & (!g1329) & (g1330) & (!g1331) & (!g147) & (!g148)) + ((g1328) & (!g1329) & (g1330) & (!g1331) & (!g147) & (g148)) + ((g1328) & (!g1329) & (g1330) & (g1331) & (!g147) & (!g148)) + ((g1328) & (!g1329) & (g1330) & (g1331) & (!g147) & (g148)) + ((g1328) & (!g1329) & (g1330) & (g1331) & (g147) & (g148)) + ((g1328) & (g1329) & (!g1330) & (!g1331) & (!g147) & (!g148)) + ((g1328) & (g1329) & (!g1330) & (!g1331) & (g147) & (!g148)) + ((g1328) & (g1329) & (!g1330) & (g1331) & (!g147) & (!g148)) + ((g1328) & (g1329) & (!g1330) & (g1331) & (g147) & (!g148)) + ((g1328) & (g1329) & (!g1330) & (g1331) & (g147) & (g148)) + ((g1328) & (g1329) & (g1330) & (!g1331) & (!g147) & (!g148)) + ((g1328) & (g1329) & (g1330) & (!g1331) & (!g147) & (g148)) + ((g1328) & (g1329) & (g1330) & (!g1331) & (g147) & (!g148)) + ((g1328) & (g1329) & (g1330) & (g1331) & (!g147) & (!g148)) + ((g1328) & (g1329) & (g1330) & (g1331) & (!g147) & (g148)) + ((g1328) & (g1329) & (g1330) & (g1331) & (g147) & (!g148)) + ((g1328) & (g1329) & (g1330) & (g1331) & (g147) & (g148)));
	assign g4834 = (((!g2152) & (!g3302) & (!sk[119]) & (g1333)) + ((!g2152) & (!g3302) & (sk[119]) & (g1333)) + ((!g2152) & (g3302) & (!sk[119]) & (!g1333)) + ((!g2152) & (g3302) & (!sk[119]) & (g1333)) + ((!g2152) & (g3302) & (sk[119]) & (g1333)) + ((g2152) & (!g3302) & (!sk[119]) & (g1333)) + ((g2152) & (g3302) & (!sk[119]) & (!g1333)) + ((g2152) & (g3302) & (!sk[119]) & (g1333)) + ((g2152) & (g3302) & (sk[119]) & (!g1333)) + ((g2152) & (g3302) & (sk[119]) & (g1333)));
	assign g4835 = (((!sk[120]) & (!g2153) & (!g3302) & (g1334)) + ((!sk[120]) & (!g2153) & (g3302) & (!g1334)) + ((!sk[120]) & (!g2153) & (g3302) & (g1334)) + ((!sk[120]) & (g2153) & (!g3302) & (g1334)) + ((!sk[120]) & (g2153) & (g3302) & (!g1334)) + ((!sk[120]) & (g2153) & (g3302) & (g1334)) + ((sk[120]) & (!g2153) & (!g3302) & (g1334)) + ((sk[120]) & (!g2153) & (g3302) & (g1334)) + ((sk[120]) & (g2153) & (g3302) & (!g1334)) + ((sk[120]) & (g2153) & (g3302) & (g1334)));
	assign g4836 = (((!g2155) & (!sk[121]) & (!g3302) & (g1335)) + ((!g2155) & (!sk[121]) & (g3302) & (!g1335)) + ((!g2155) & (!sk[121]) & (g3302) & (g1335)) + ((!g2155) & (sk[121]) & (!g3302) & (g1335)) + ((!g2155) & (sk[121]) & (g3302) & (g1335)) + ((g2155) & (!sk[121]) & (!g3302) & (g1335)) + ((g2155) & (!sk[121]) & (g3302) & (!g1335)) + ((g2155) & (!sk[121]) & (g3302) & (g1335)) + ((g2155) & (sk[121]) & (g3302) & (!g1335)) + ((g2155) & (sk[121]) & (g3302) & (g1335)));
	assign g4837 = (((!g2157) & (!sk[122]) & (!g3302) & (g1336)) + ((!g2157) & (!sk[122]) & (g3302) & (!g1336)) + ((!g2157) & (!sk[122]) & (g3302) & (g1336)) + ((!g2157) & (sk[122]) & (!g3302) & (g1336)) + ((!g2157) & (sk[122]) & (g3302) & (g1336)) + ((g2157) & (!sk[122]) & (!g3302) & (g1336)) + ((g2157) & (!sk[122]) & (g3302) & (!g1336)) + ((g2157) & (!sk[122]) & (g3302) & (g1336)) + ((g2157) & (sk[122]) & (g3302) & (!g1336)) + ((g2157) & (sk[122]) & (g3302) & (g1336)));
	assign g1337 = (((!g1333) & (!g1334) & (!g1335) & (g1336) & (g147) & (g148)) + ((!g1333) & (!g1334) & (g1335) & (!g1336) & (!g147) & (g148)) + ((!g1333) & (!g1334) & (g1335) & (g1336) & (!g147) & (g148)) + ((!g1333) & (!g1334) & (g1335) & (g1336) & (g147) & (g148)) + ((!g1333) & (g1334) & (!g1335) & (!g1336) & (g147) & (!g148)) + ((!g1333) & (g1334) & (!g1335) & (g1336) & (g147) & (!g148)) + ((!g1333) & (g1334) & (!g1335) & (g1336) & (g147) & (g148)) + ((!g1333) & (g1334) & (g1335) & (!g1336) & (!g147) & (g148)) + ((!g1333) & (g1334) & (g1335) & (!g1336) & (g147) & (!g148)) + ((!g1333) & (g1334) & (g1335) & (g1336) & (!g147) & (g148)) + ((!g1333) & (g1334) & (g1335) & (g1336) & (g147) & (!g148)) + ((!g1333) & (g1334) & (g1335) & (g1336) & (g147) & (g148)) + ((g1333) & (!g1334) & (!g1335) & (!g1336) & (!g147) & (!g148)) + ((g1333) & (!g1334) & (!g1335) & (g1336) & (!g147) & (!g148)) + ((g1333) & (!g1334) & (!g1335) & (g1336) & (g147) & (g148)) + ((g1333) & (!g1334) & (g1335) & (!g1336) & (!g147) & (!g148)) + ((g1333) & (!g1334) & (g1335) & (!g1336) & (!g147) & (g148)) + ((g1333) & (!g1334) & (g1335) & (g1336) & (!g147) & (!g148)) + ((g1333) & (!g1334) & (g1335) & (g1336) & (!g147) & (g148)) + ((g1333) & (!g1334) & (g1335) & (g1336) & (g147) & (g148)) + ((g1333) & (g1334) & (!g1335) & (!g1336) & (!g147) & (!g148)) + ((g1333) & (g1334) & (!g1335) & (!g1336) & (g147) & (!g148)) + ((g1333) & (g1334) & (!g1335) & (g1336) & (!g147) & (!g148)) + ((g1333) & (g1334) & (!g1335) & (g1336) & (g147) & (!g148)) + ((g1333) & (g1334) & (!g1335) & (g1336) & (g147) & (g148)) + ((g1333) & (g1334) & (g1335) & (!g1336) & (!g147) & (!g148)) + ((g1333) & (g1334) & (g1335) & (!g1336) & (!g147) & (g148)) + ((g1333) & (g1334) & (g1335) & (!g1336) & (g147) & (!g148)) + ((g1333) & (g1334) & (g1335) & (g1336) & (!g147) & (!g148)) + ((g1333) & (g1334) & (g1335) & (g1336) & (!g147) & (g148)) + ((g1333) & (g1334) & (g1335) & (g1336) & (g147) & (!g148)) + ((g1333) & (g1334) & (g1335) & (g1336) & (g147) & (g148)));
	assign g4838 = (((!g2158) & (!sk[124]) & (!g3302) & (g1338)) + ((!g2158) & (!sk[124]) & (g3302) & (!g1338)) + ((!g2158) & (!sk[124]) & (g3302) & (g1338)) + ((!g2158) & (sk[124]) & (!g3302) & (g1338)) + ((!g2158) & (sk[124]) & (g3302) & (g1338)) + ((g2158) & (!sk[124]) & (!g3302) & (g1338)) + ((g2158) & (!sk[124]) & (g3302) & (!g1338)) + ((g2158) & (!sk[124]) & (g3302) & (g1338)) + ((g2158) & (sk[124]) & (g3302) & (!g1338)) + ((g2158) & (sk[124]) & (g3302) & (g1338)));
	assign g4839 = (((!sk[125]) & (!g2159) & (!g3302) & (g1339)) + ((!sk[125]) & (!g2159) & (g3302) & (!g1339)) + ((!sk[125]) & (!g2159) & (g3302) & (g1339)) + ((!sk[125]) & (g2159) & (!g3302) & (g1339)) + ((!sk[125]) & (g2159) & (g3302) & (!g1339)) + ((!sk[125]) & (g2159) & (g3302) & (g1339)) + ((sk[125]) & (!g2159) & (!g3302) & (g1339)) + ((sk[125]) & (!g2159) & (g3302) & (g1339)) + ((sk[125]) & (g2159) & (g3302) & (!g1339)) + ((sk[125]) & (g2159) & (g3302) & (g1339)));
	assign g4840 = (((!g2160) & (!sk[126]) & (!g3302) & (g1340)) + ((!g2160) & (!sk[126]) & (g3302) & (!g1340)) + ((!g2160) & (!sk[126]) & (g3302) & (g1340)) + ((!g2160) & (sk[126]) & (!g3302) & (g1340)) + ((!g2160) & (sk[126]) & (g3302) & (g1340)) + ((g2160) & (!sk[126]) & (!g3302) & (g1340)) + ((g2160) & (!sk[126]) & (g3302) & (!g1340)) + ((g2160) & (!sk[126]) & (g3302) & (g1340)) + ((g2160) & (sk[126]) & (g3302) & (!g1340)) + ((g2160) & (sk[126]) & (g3302) & (g1340)));
	assign g4841 = (((!sk[127]) & (!g2161) & (!g3302) & (g1341)) + ((!sk[127]) & (!g2161) & (g3302) & (!g1341)) + ((!sk[127]) & (!g2161) & (g3302) & (g1341)) + ((!sk[127]) & (g2161) & (!g3302) & (g1341)) + ((!sk[127]) & (g2161) & (g3302) & (!g1341)) + ((!sk[127]) & (g2161) & (g3302) & (g1341)) + ((sk[127]) & (!g2161) & (!g3302) & (g1341)) + ((sk[127]) & (!g2161) & (g3302) & (g1341)) + ((sk[127]) & (g2161) & (g3302) & (!g1341)) + ((sk[127]) & (g2161) & (g3302) & (g1341)));
	assign g1342 = (((!g1338) & (!g1339) & (!g1340) & (g1341) & (g147) & (g148)) + ((!g1338) & (!g1339) & (g1340) & (!g1341) & (!g147) & (g148)) + ((!g1338) & (!g1339) & (g1340) & (g1341) & (!g147) & (g148)) + ((!g1338) & (!g1339) & (g1340) & (g1341) & (g147) & (g148)) + ((!g1338) & (g1339) & (!g1340) & (!g1341) & (g147) & (!g148)) + ((!g1338) & (g1339) & (!g1340) & (g1341) & (g147) & (!g148)) + ((!g1338) & (g1339) & (!g1340) & (g1341) & (g147) & (g148)) + ((!g1338) & (g1339) & (g1340) & (!g1341) & (!g147) & (g148)) + ((!g1338) & (g1339) & (g1340) & (!g1341) & (g147) & (!g148)) + ((!g1338) & (g1339) & (g1340) & (g1341) & (!g147) & (g148)) + ((!g1338) & (g1339) & (g1340) & (g1341) & (g147) & (!g148)) + ((!g1338) & (g1339) & (g1340) & (g1341) & (g147) & (g148)) + ((g1338) & (!g1339) & (!g1340) & (!g1341) & (!g147) & (!g148)) + ((g1338) & (!g1339) & (!g1340) & (g1341) & (!g147) & (!g148)) + ((g1338) & (!g1339) & (!g1340) & (g1341) & (g147) & (g148)) + ((g1338) & (!g1339) & (g1340) & (!g1341) & (!g147) & (!g148)) + ((g1338) & (!g1339) & (g1340) & (!g1341) & (!g147) & (g148)) + ((g1338) & (!g1339) & (g1340) & (g1341) & (!g147) & (!g148)) + ((g1338) & (!g1339) & (g1340) & (g1341) & (!g147) & (g148)) + ((g1338) & (!g1339) & (g1340) & (g1341) & (g147) & (g148)) + ((g1338) & (g1339) & (!g1340) & (!g1341) & (!g147) & (!g148)) + ((g1338) & (g1339) & (!g1340) & (!g1341) & (g147) & (!g148)) + ((g1338) & (g1339) & (!g1340) & (g1341) & (!g147) & (!g148)) + ((g1338) & (g1339) & (!g1340) & (g1341) & (g147) & (!g148)) + ((g1338) & (g1339) & (!g1340) & (g1341) & (g147) & (g148)) + ((g1338) & (g1339) & (g1340) & (!g1341) & (!g147) & (!g148)) + ((g1338) & (g1339) & (g1340) & (!g1341) & (!g147) & (g148)) + ((g1338) & (g1339) & (g1340) & (!g1341) & (g147) & (!g148)) + ((g1338) & (g1339) & (g1340) & (g1341) & (!g147) & (!g148)) + ((g1338) & (g1339) & (g1340) & (g1341) & (!g147) & (g148)) + ((g1338) & (g1339) & (g1340) & (g1341) & (g147) & (!g148)) + ((g1338) & (g1339) & (g1340) & (g1341) & (g147) & (g148)));
	assign g1343 = (((!g1327) & (!g1332) & (!g1337) & (g1342) & (g165) & (g166)) + ((!g1327) & (!g1332) & (g1337) & (!g1342) & (!g165) & (g166)) + ((!g1327) & (!g1332) & (g1337) & (g1342) & (!g165) & (g166)) + ((!g1327) & (!g1332) & (g1337) & (g1342) & (g165) & (g166)) + ((!g1327) & (g1332) & (!g1337) & (!g1342) & (g165) & (!g166)) + ((!g1327) & (g1332) & (!g1337) & (g1342) & (g165) & (!g166)) + ((!g1327) & (g1332) & (!g1337) & (g1342) & (g165) & (g166)) + ((!g1327) & (g1332) & (g1337) & (!g1342) & (!g165) & (g166)) + ((!g1327) & (g1332) & (g1337) & (!g1342) & (g165) & (!g166)) + ((!g1327) & (g1332) & (g1337) & (g1342) & (!g165) & (g166)) + ((!g1327) & (g1332) & (g1337) & (g1342) & (g165) & (!g166)) + ((!g1327) & (g1332) & (g1337) & (g1342) & (g165) & (g166)) + ((g1327) & (!g1332) & (!g1337) & (!g1342) & (!g165) & (!g166)) + ((g1327) & (!g1332) & (!g1337) & (g1342) & (!g165) & (!g166)) + ((g1327) & (!g1332) & (!g1337) & (g1342) & (g165) & (g166)) + ((g1327) & (!g1332) & (g1337) & (!g1342) & (!g165) & (!g166)) + ((g1327) & (!g1332) & (g1337) & (!g1342) & (!g165) & (g166)) + ((g1327) & (!g1332) & (g1337) & (g1342) & (!g165) & (!g166)) + ((g1327) & (!g1332) & (g1337) & (g1342) & (!g165) & (g166)) + ((g1327) & (!g1332) & (g1337) & (g1342) & (g165) & (g166)) + ((g1327) & (g1332) & (!g1337) & (!g1342) & (!g165) & (!g166)) + ((g1327) & (g1332) & (!g1337) & (!g1342) & (g165) & (!g166)) + ((g1327) & (g1332) & (!g1337) & (g1342) & (!g165) & (!g166)) + ((g1327) & (g1332) & (!g1337) & (g1342) & (g165) & (!g166)) + ((g1327) & (g1332) & (!g1337) & (g1342) & (g165) & (g166)) + ((g1327) & (g1332) & (g1337) & (!g1342) & (!g165) & (!g166)) + ((g1327) & (g1332) & (g1337) & (!g1342) & (!g165) & (g166)) + ((g1327) & (g1332) & (g1337) & (!g1342) & (g165) & (!g166)) + ((g1327) & (g1332) & (g1337) & (g1342) & (!g165) & (!g166)) + ((g1327) & (g1332) & (g1337) & (g1342) & (!g165) & (g166)) + ((g1327) & (g1332) & (g1337) & (g1342) & (g165) & (!g166)) + ((g1327) & (g1332) & (g1337) & (g1342) & (g165) & (g166)));
	assign g4842 = (((!g2173) & (!g3302) & (!sk[2]) & (g1344)) + ((!g2173) & (!g3302) & (sk[2]) & (g1344)) + ((!g2173) & (g3302) & (!sk[2]) & (!g1344)) + ((!g2173) & (g3302) & (!sk[2]) & (g1344)) + ((!g2173) & (g3302) & (sk[2]) & (g1344)) + ((g2173) & (!g3302) & (!sk[2]) & (g1344)) + ((g2173) & (g3302) & (!sk[2]) & (!g1344)) + ((g2173) & (g3302) & (!sk[2]) & (g1344)) + ((g2173) & (g3302) & (sk[2]) & (!g1344)) + ((g2173) & (g3302) & (sk[2]) & (g1344)));
	assign g4843 = (((!g2174) & (!sk[3]) & (!g3302) & (g1345)) + ((!g2174) & (!sk[3]) & (g3302) & (!g1345)) + ((!g2174) & (!sk[3]) & (g3302) & (g1345)) + ((!g2174) & (sk[3]) & (!g3302) & (g1345)) + ((!g2174) & (sk[3]) & (g3302) & (g1345)) + ((g2174) & (!sk[3]) & (!g3302) & (g1345)) + ((g2174) & (!sk[3]) & (g3302) & (!g1345)) + ((g2174) & (!sk[3]) & (g3302) & (g1345)) + ((g2174) & (sk[3]) & (g3302) & (!g1345)) + ((g2174) & (sk[3]) & (g3302) & (g1345)));
	assign g4844 = (((!sk[4]) & (!g2175) & (!g3302) & (g1346)) + ((!sk[4]) & (!g2175) & (g3302) & (!g1346)) + ((!sk[4]) & (!g2175) & (g3302) & (g1346)) + ((!sk[4]) & (g2175) & (!g3302) & (g1346)) + ((!sk[4]) & (g2175) & (g3302) & (!g1346)) + ((!sk[4]) & (g2175) & (g3302) & (g1346)) + ((sk[4]) & (!g2175) & (!g3302) & (g1346)) + ((sk[4]) & (!g2175) & (g3302) & (g1346)) + ((sk[4]) & (g2175) & (g3302) & (!g1346)) + ((sk[4]) & (g2175) & (g3302) & (g1346)));
	assign g4845 = (((!g2176) & (!g3302) & (!sk[5]) & (g1347)) + ((!g2176) & (!g3302) & (sk[5]) & (g1347)) + ((!g2176) & (g3302) & (!sk[5]) & (!g1347)) + ((!g2176) & (g3302) & (!sk[5]) & (g1347)) + ((!g2176) & (g3302) & (sk[5]) & (g1347)) + ((g2176) & (!g3302) & (!sk[5]) & (g1347)) + ((g2176) & (g3302) & (!sk[5]) & (!g1347)) + ((g2176) & (g3302) & (!sk[5]) & (g1347)) + ((g2176) & (g3302) & (sk[5]) & (!g1347)) + ((g2176) & (g3302) & (sk[5]) & (g1347)));
	assign g1348 = (((!g1344) & (!g1345) & (!g1346) & (g1347) & (g165) & (g166)) + ((!g1344) & (!g1345) & (g1346) & (!g1347) & (!g165) & (g166)) + ((!g1344) & (!g1345) & (g1346) & (g1347) & (!g165) & (g166)) + ((!g1344) & (!g1345) & (g1346) & (g1347) & (g165) & (g166)) + ((!g1344) & (g1345) & (!g1346) & (!g1347) & (g165) & (!g166)) + ((!g1344) & (g1345) & (!g1346) & (g1347) & (g165) & (!g166)) + ((!g1344) & (g1345) & (!g1346) & (g1347) & (g165) & (g166)) + ((!g1344) & (g1345) & (g1346) & (!g1347) & (!g165) & (g166)) + ((!g1344) & (g1345) & (g1346) & (!g1347) & (g165) & (!g166)) + ((!g1344) & (g1345) & (g1346) & (g1347) & (!g165) & (g166)) + ((!g1344) & (g1345) & (g1346) & (g1347) & (g165) & (!g166)) + ((!g1344) & (g1345) & (g1346) & (g1347) & (g165) & (g166)) + ((g1344) & (!g1345) & (!g1346) & (!g1347) & (!g165) & (!g166)) + ((g1344) & (!g1345) & (!g1346) & (g1347) & (!g165) & (!g166)) + ((g1344) & (!g1345) & (!g1346) & (g1347) & (g165) & (g166)) + ((g1344) & (!g1345) & (g1346) & (!g1347) & (!g165) & (!g166)) + ((g1344) & (!g1345) & (g1346) & (!g1347) & (!g165) & (g166)) + ((g1344) & (!g1345) & (g1346) & (g1347) & (!g165) & (!g166)) + ((g1344) & (!g1345) & (g1346) & (g1347) & (!g165) & (g166)) + ((g1344) & (!g1345) & (g1346) & (g1347) & (g165) & (g166)) + ((g1344) & (g1345) & (!g1346) & (!g1347) & (!g165) & (!g166)) + ((g1344) & (g1345) & (!g1346) & (!g1347) & (g165) & (!g166)) + ((g1344) & (g1345) & (!g1346) & (g1347) & (!g165) & (!g166)) + ((g1344) & (g1345) & (!g1346) & (g1347) & (g165) & (!g166)) + ((g1344) & (g1345) & (!g1346) & (g1347) & (g165) & (g166)) + ((g1344) & (g1345) & (g1346) & (!g1347) & (!g165) & (!g166)) + ((g1344) & (g1345) & (g1346) & (!g1347) & (!g165) & (g166)) + ((g1344) & (g1345) & (g1346) & (!g1347) & (g165) & (!g166)) + ((g1344) & (g1345) & (g1346) & (g1347) & (!g165) & (!g166)) + ((g1344) & (g1345) & (g1346) & (g1347) & (!g165) & (g166)) + ((g1344) & (g1345) & (g1346) & (g1347) & (g165) & (!g166)) + ((g1344) & (g1345) & (g1346) & (g1347) & (g165) & (g166)));
	assign g4846 = (((!g2177) & (!sk[7]) & (!g3302) & (g1349)) + ((!g2177) & (!sk[7]) & (g3302) & (!g1349)) + ((!g2177) & (!sk[7]) & (g3302) & (g1349)) + ((!g2177) & (sk[7]) & (!g3302) & (g1349)) + ((!g2177) & (sk[7]) & (g3302) & (g1349)) + ((g2177) & (!sk[7]) & (!g3302) & (g1349)) + ((g2177) & (!sk[7]) & (g3302) & (!g1349)) + ((g2177) & (!sk[7]) & (g3302) & (g1349)) + ((g2177) & (sk[7]) & (g3302) & (!g1349)) + ((g2177) & (sk[7]) & (g3302) & (g1349)));
	assign g4847 = (((!g2178) & (!g3302) & (!sk[8]) & (g1350)) + ((!g2178) & (!g3302) & (sk[8]) & (g1350)) + ((!g2178) & (g3302) & (!sk[8]) & (!g1350)) + ((!g2178) & (g3302) & (!sk[8]) & (g1350)) + ((!g2178) & (g3302) & (sk[8]) & (g1350)) + ((g2178) & (!g3302) & (!sk[8]) & (g1350)) + ((g2178) & (g3302) & (!sk[8]) & (!g1350)) + ((g2178) & (g3302) & (!sk[8]) & (g1350)) + ((g2178) & (g3302) & (sk[8]) & (!g1350)) + ((g2178) & (g3302) & (sk[8]) & (g1350)));
	assign g4848 = (((!g2179) & (!g3302) & (!sk[9]) & (g1351)) + ((!g2179) & (!g3302) & (sk[9]) & (g1351)) + ((!g2179) & (g3302) & (!sk[9]) & (!g1351)) + ((!g2179) & (g3302) & (!sk[9]) & (g1351)) + ((!g2179) & (g3302) & (sk[9]) & (g1351)) + ((g2179) & (!g3302) & (!sk[9]) & (g1351)) + ((g2179) & (g3302) & (!sk[9]) & (!g1351)) + ((g2179) & (g3302) & (!sk[9]) & (g1351)) + ((g2179) & (g3302) & (sk[9]) & (!g1351)) + ((g2179) & (g3302) & (sk[9]) & (g1351)));
	assign g1352 = (((!g165) & (!g166) & (!g1349) & (g1350) & (!sk[10]) & (!g1351)) + ((!g165) & (!g166) & (!g1349) & (g1350) & (!sk[10]) & (g1351)) + ((!g165) & (!g166) & (g1349) & (!g1350) & (!sk[10]) & (!g1351)) + ((!g165) & (!g166) & (g1349) & (!g1350) & (!sk[10]) & (g1351)) + ((!g165) & (!g166) & (g1349) & (g1350) & (!sk[10]) & (!g1351)) + ((!g165) & (!g166) & (g1349) & (g1350) & (!sk[10]) & (g1351)) + ((!g165) & (g166) & (!g1349) & (!g1350) & (!sk[10]) & (!g1351)) + ((!g165) & (g166) & (!g1349) & (!g1350) & (!sk[10]) & (g1351)) + ((!g165) & (g166) & (!g1349) & (!g1350) & (sk[10]) & (g1351)) + ((!g165) & (g166) & (!g1349) & (g1350) & (!sk[10]) & (!g1351)) + ((!g165) & (g166) & (!g1349) & (g1350) & (!sk[10]) & (g1351)) + ((!g165) & (g166) & (!g1349) & (g1350) & (sk[10]) & (g1351)) + ((!g165) & (g166) & (g1349) & (!g1350) & (!sk[10]) & (!g1351)) + ((!g165) & (g166) & (g1349) & (!g1350) & (!sk[10]) & (g1351)) + ((!g165) & (g166) & (g1349) & (!g1350) & (sk[10]) & (g1351)) + ((!g165) & (g166) & (g1349) & (g1350) & (!sk[10]) & (!g1351)) + ((!g165) & (g166) & (g1349) & (g1350) & (!sk[10]) & (g1351)) + ((!g165) & (g166) & (g1349) & (g1350) & (sk[10]) & (g1351)) + ((g165) & (!g166) & (!g1349) & (g1350) & (!sk[10]) & (!g1351)) + ((g165) & (!g166) & (!g1349) & (g1350) & (!sk[10]) & (g1351)) + ((g165) & (!g166) & (g1349) & (!g1350) & (!sk[10]) & (!g1351)) + ((g165) & (!g166) & (g1349) & (!g1350) & (!sk[10]) & (g1351)) + ((g165) & (!g166) & (g1349) & (!g1350) & (sk[10]) & (!g1351)) + ((g165) & (!g166) & (g1349) & (!g1350) & (sk[10]) & (g1351)) + ((g165) & (!g166) & (g1349) & (g1350) & (!sk[10]) & (!g1351)) + ((g165) & (!g166) & (g1349) & (g1350) & (!sk[10]) & (g1351)) + ((g165) & (!g166) & (g1349) & (g1350) & (sk[10]) & (!g1351)) + ((g165) & (!g166) & (g1349) & (g1350) & (sk[10]) & (g1351)) + ((g165) & (g166) & (!g1349) & (!g1350) & (!sk[10]) & (!g1351)) + ((g165) & (g166) & (!g1349) & (!g1350) & (!sk[10]) & (g1351)) + ((g165) & (g166) & (!g1349) & (g1350) & (!sk[10]) & (!g1351)) + ((g165) & (g166) & (!g1349) & (g1350) & (!sk[10]) & (g1351)) + ((g165) & (g166) & (!g1349) & (g1350) & (sk[10]) & (!g1351)) + ((g165) & (g166) & (!g1349) & (g1350) & (sk[10]) & (g1351)) + ((g165) & (g166) & (g1349) & (!g1350) & (!sk[10]) & (!g1351)) + ((g165) & (g166) & (g1349) & (!g1350) & (!sk[10]) & (g1351)) + ((g165) & (g166) & (g1349) & (g1350) & (!sk[10]) & (!g1351)) + ((g165) & (g166) & (g1349) & (g1350) & (!sk[10]) & (g1351)) + ((g165) & (g166) & (g1349) & (g1350) & (sk[10]) & (!g1351)) + ((g165) & (g166) & (g1349) & (g1350) & (sk[10]) & (g1351)));
	assign g4849 = (((!g2162) & (!sk[11]) & (!g3302) & (g1353)) + ((!g2162) & (!sk[11]) & (g3302) & (!g1353)) + ((!g2162) & (!sk[11]) & (g3302) & (g1353)) + ((!g2162) & (sk[11]) & (!g3302) & (g1353)) + ((!g2162) & (sk[11]) & (g3302) & (g1353)) + ((g2162) & (!sk[11]) & (!g3302) & (g1353)) + ((g2162) & (!sk[11]) & (g3302) & (!g1353)) + ((g2162) & (!sk[11]) & (g3302) & (g1353)) + ((g2162) & (sk[11]) & (g3302) & (!g1353)) + ((g2162) & (sk[11]) & (g3302) & (g1353)));
	assign g4850 = (((!g2164) & (!sk[12]) & (!g3302) & (g1354)) + ((!g2164) & (!sk[12]) & (g3302) & (!g1354)) + ((!g2164) & (!sk[12]) & (g3302) & (g1354)) + ((!g2164) & (sk[12]) & (!g3302) & (g1354)) + ((!g2164) & (sk[12]) & (g3302) & (g1354)) + ((g2164) & (!sk[12]) & (!g3302) & (g1354)) + ((g2164) & (!sk[12]) & (g3302) & (!g1354)) + ((g2164) & (!sk[12]) & (g3302) & (g1354)) + ((g2164) & (sk[12]) & (g3302) & (!g1354)) + ((g2164) & (sk[12]) & (g3302) & (g1354)));
	assign g4851 = (((!g2166) & (!g3302) & (!sk[13]) & (g1355)) + ((!g2166) & (!g3302) & (sk[13]) & (g1355)) + ((!g2166) & (g3302) & (!sk[13]) & (!g1355)) + ((!g2166) & (g3302) & (!sk[13]) & (g1355)) + ((!g2166) & (g3302) & (sk[13]) & (g1355)) + ((g2166) & (!g3302) & (!sk[13]) & (g1355)) + ((g2166) & (g3302) & (!sk[13]) & (!g1355)) + ((g2166) & (g3302) & (!sk[13]) & (g1355)) + ((g2166) & (g3302) & (sk[13]) & (!g1355)) + ((g2166) & (g3302) & (sk[13]) & (g1355)));
	assign g4852 = (((!g2168) & (!g3302) & (!sk[14]) & (g1356)) + ((!g2168) & (!g3302) & (sk[14]) & (g1356)) + ((!g2168) & (g3302) & (!sk[14]) & (!g1356)) + ((!g2168) & (g3302) & (!sk[14]) & (g1356)) + ((!g2168) & (g3302) & (sk[14]) & (g1356)) + ((g2168) & (!g3302) & (!sk[14]) & (g1356)) + ((g2168) & (g3302) & (!sk[14]) & (!g1356)) + ((g2168) & (g3302) & (!sk[14]) & (g1356)) + ((g2168) & (g3302) & (sk[14]) & (!g1356)) + ((g2168) & (g3302) & (sk[14]) & (g1356)));
	assign g1357 = (((!g1353) & (!g1354) & (!g1355) & (g1356) & (g165) & (g166)) + ((!g1353) & (!g1354) & (g1355) & (!g1356) & (!g165) & (g166)) + ((!g1353) & (!g1354) & (g1355) & (g1356) & (!g165) & (g166)) + ((!g1353) & (!g1354) & (g1355) & (g1356) & (g165) & (g166)) + ((!g1353) & (g1354) & (!g1355) & (!g1356) & (g165) & (!g166)) + ((!g1353) & (g1354) & (!g1355) & (g1356) & (g165) & (!g166)) + ((!g1353) & (g1354) & (!g1355) & (g1356) & (g165) & (g166)) + ((!g1353) & (g1354) & (g1355) & (!g1356) & (!g165) & (g166)) + ((!g1353) & (g1354) & (g1355) & (!g1356) & (g165) & (!g166)) + ((!g1353) & (g1354) & (g1355) & (g1356) & (!g165) & (g166)) + ((!g1353) & (g1354) & (g1355) & (g1356) & (g165) & (!g166)) + ((!g1353) & (g1354) & (g1355) & (g1356) & (g165) & (g166)) + ((g1353) & (!g1354) & (!g1355) & (!g1356) & (!g165) & (!g166)) + ((g1353) & (!g1354) & (!g1355) & (g1356) & (!g165) & (!g166)) + ((g1353) & (!g1354) & (!g1355) & (g1356) & (g165) & (g166)) + ((g1353) & (!g1354) & (g1355) & (!g1356) & (!g165) & (!g166)) + ((g1353) & (!g1354) & (g1355) & (!g1356) & (!g165) & (g166)) + ((g1353) & (!g1354) & (g1355) & (g1356) & (!g165) & (!g166)) + ((g1353) & (!g1354) & (g1355) & (g1356) & (!g165) & (g166)) + ((g1353) & (!g1354) & (g1355) & (g1356) & (g165) & (g166)) + ((g1353) & (g1354) & (!g1355) & (!g1356) & (!g165) & (!g166)) + ((g1353) & (g1354) & (!g1355) & (!g1356) & (g165) & (!g166)) + ((g1353) & (g1354) & (!g1355) & (g1356) & (!g165) & (!g166)) + ((g1353) & (g1354) & (!g1355) & (g1356) & (g165) & (!g166)) + ((g1353) & (g1354) & (!g1355) & (g1356) & (g165) & (g166)) + ((g1353) & (g1354) & (g1355) & (!g1356) & (!g165) & (!g166)) + ((g1353) & (g1354) & (g1355) & (!g1356) & (!g165) & (g166)) + ((g1353) & (g1354) & (g1355) & (!g1356) & (g165) & (!g166)) + ((g1353) & (g1354) & (g1355) & (g1356) & (!g165) & (!g166)) + ((g1353) & (g1354) & (g1355) & (g1356) & (!g165) & (g166)) + ((g1353) & (g1354) & (g1355) & (g1356) & (g165) & (!g166)) + ((g1353) & (g1354) & (g1355) & (g1356) & (g165) & (g166)));
	assign g4853 = (((!g2169) & (!sk[16]) & (!g3302) & (g1358)) + ((!g2169) & (!sk[16]) & (g3302) & (!g1358)) + ((!g2169) & (!sk[16]) & (g3302) & (g1358)) + ((!g2169) & (sk[16]) & (!g3302) & (g1358)) + ((!g2169) & (sk[16]) & (g3302) & (g1358)) + ((g2169) & (!sk[16]) & (!g3302) & (g1358)) + ((g2169) & (!sk[16]) & (g3302) & (!g1358)) + ((g2169) & (!sk[16]) & (g3302) & (g1358)) + ((g2169) & (sk[16]) & (g3302) & (!g1358)) + ((g2169) & (sk[16]) & (g3302) & (g1358)));
	assign g4854 = (((!g2170) & (!g3302) & (!sk[17]) & (g1359)) + ((!g2170) & (!g3302) & (sk[17]) & (g1359)) + ((!g2170) & (g3302) & (!sk[17]) & (!g1359)) + ((!g2170) & (g3302) & (!sk[17]) & (g1359)) + ((!g2170) & (g3302) & (sk[17]) & (g1359)) + ((g2170) & (!g3302) & (!sk[17]) & (g1359)) + ((g2170) & (g3302) & (!sk[17]) & (!g1359)) + ((g2170) & (g3302) & (!sk[17]) & (g1359)) + ((g2170) & (g3302) & (sk[17]) & (!g1359)) + ((g2170) & (g3302) & (sk[17]) & (g1359)));
	assign g4855 = (((!g2171) & (!sk[18]) & (!g3302) & (g1360)) + ((!g2171) & (!sk[18]) & (g3302) & (!g1360)) + ((!g2171) & (!sk[18]) & (g3302) & (g1360)) + ((!g2171) & (sk[18]) & (!g3302) & (g1360)) + ((!g2171) & (sk[18]) & (g3302) & (g1360)) + ((g2171) & (!sk[18]) & (!g3302) & (g1360)) + ((g2171) & (!sk[18]) & (g3302) & (!g1360)) + ((g2171) & (!sk[18]) & (g3302) & (g1360)) + ((g2171) & (sk[18]) & (g3302) & (!g1360)) + ((g2171) & (sk[18]) & (g3302) & (g1360)));
	assign g4856 = (((!sk[19]) & (!g2172) & (!g3302) & (g1361)) + ((!sk[19]) & (!g2172) & (g3302) & (!g1361)) + ((!sk[19]) & (!g2172) & (g3302) & (g1361)) + ((!sk[19]) & (g2172) & (!g3302) & (g1361)) + ((!sk[19]) & (g2172) & (g3302) & (!g1361)) + ((!sk[19]) & (g2172) & (g3302) & (g1361)) + ((sk[19]) & (!g2172) & (!g3302) & (g1361)) + ((sk[19]) & (!g2172) & (g3302) & (g1361)) + ((sk[19]) & (g2172) & (g3302) & (!g1361)) + ((sk[19]) & (g2172) & (g3302) & (g1361)));
	assign g1362 = (((!g1358) & (!g1359) & (!g1360) & (g1361) & (g165) & (g166)) + ((!g1358) & (!g1359) & (g1360) & (!g1361) & (!g165) & (g166)) + ((!g1358) & (!g1359) & (g1360) & (g1361) & (!g165) & (g166)) + ((!g1358) & (!g1359) & (g1360) & (g1361) & (g165) & (g166)) + ((!g1358) & (g1359) & (!g1360) & (!g1361) & (g165) & (!g166)) + ((!g1358) & (g1359) & (!g1360) & (g1361) & (g165) & (!g166)) + ((!g1358) & (g1359) & (!g1360) & (g1361) & (g165) & (g166)) + ((!g1358) & (g1359) & (g1360) & (!g1361) & (!g165) & (g166)) + ((!g1358) & (g1359) & (g1360) & (!g1361) & (g165) & (!g166)) + ((!g1358) & (g1359) & (g1360) & (g1361) & (!g165) & (g166)) + ((!g1358) & (g1359) & (g1360) & (g1361) & (g165) & (!g166)) + ((!g1358) & (g1359) & (g1360) & (g1361) & (g165) & (g166)) + ((g1358) & (!g1359) & (!g1360) & (!g1361) & (!g165) & (!g166)) + ((g1358) & (!g1359) & (!g1360) & (g1361) & (!g165) & (!g166)) + ((g1358) & (!g1359) & (!g1360) & (g1361) & (g165) & (g166)) + ((g1358) & (!g1359) & (g1360) & (!g1361) & (!g165) & (!g166)) + ((g1358) & (!g1359) & (g1360) & (!g1361) & (!g165) & (g166)) + ((g1358) & (!g1359) & (g1360) & (g1361) & (!g165) & (!g166)) + ((g1358) & (!g1359) & (g1360) & (g1361) & (!g165) & (g166)) + ((g1358) & (!g1359) & (g1360) & (g1361) & (g165) & (g166)) + ((g1358) & (g1359) & (!g1360) & (!g1361) & (!g165) & (!g166)) + ((g1358) & (g1359) & (!g1360) & (!g1361) & (g165) & (!g166)) + ((g1358) & (g1359) & (!g1360) & (g1361) & (!g165) & (!g166)) + ((g1358) & (g1359) & (!g1360) & (g1361) & (g165) & (!g166)) + ((g1358) & (g1359) & (!g1360) & (g1361) & (g165) & (g166)) + ((g1358) & (g1359) & (g1360) & (!g1361) & (!g165) & (!g166)) + ((g1358) & (g1359) & (g1360) & (!g1361) & (!g165) & (g166)) + ((g1358) & (g1359) & (g1360) & (!g1361) & (g165) & (!g166)) + ((g1358) & (g1359) & (g1360) & (g1361) & (!g165) & (!g166)) + ((g1358) & (g1359) & (g1360) & (g1361) & (!g165) & (g166)) + ((g1358) & (g1359) & (g1360) & (g1361) & (g165) & (!g166)) + ((g1358) & (g1359) & (g1360) & (g1361) & (g165) & (g166)));
	assign g1363 = (((!g147) & (!g148) & (!g1348) & (g1352) & (!g1357) & (!g1362)) + ((!g147) & (!g148) & (!g1348) & (g1352) & (!g1357) & (g1362)) + ((!g147) & (!g148) & (!g1348) & (g1352) & (g1357) & (!g1362)) + ((!g147) & (!g148) & (!g1348) & (g1352) & (g1357) & (g1362)) + ((!g147) & (!g148) & (g1348) & (g1352) & (!g1357) & (!g1362)) + ((!g147) & (!g148) & (g1348) & (g1352) & (!g1357) & (g1362)) + ((!g147) & (!g148) & (g1348) & (g1352) & (g1357) & (!g1362)) + ((!g147) & (!g148) & (g1348) & (g1352) & (g1357) & (g1362)) + ((!g147) & (g148) & (!g1348) & (!g1352) & (!g1357) & (g1362)) + ((!g147) & (g148) & (!g1348) & (!g1352) & (g1357) & (g1362)) + ((!g147) & (g148) & (!g1348) & (g1352) & (!g1357) & (g1362)) + ((!g147) & (g148) & (!g1348) & (g1352) & (g1357) & (g1362)) + ((!g147) & (g148) & (g1348) & (!g1352) & (!g1357) & (g1362)) + ((!g147) & (g148) & (g1348) & (!g1352) & (g1357) & (g1362)) + ((!g147) & (g148) & (g1348) & (g1352) & (!g1357) & (g1362)) + ((!g147) & (g148) & (g1348) & (g1352) & (g1357) & (g1362)) + ((g147) & (!g148) & (g1348) & (!g1352) & (!g1357) & (!g1362)) + ((g147) & (!g148) & (g1348) & (!g1352) & (!g1357) & (g1362)) + ((g147) & (!g148) & (g1348) & (!g1352) & (g1357) & (!g1362)) + ((g147) & (!g148) & (g1348) & (!g1352) & (g1357) & (g1362)) + ((g147) & (!g148) & (g1348) & (g1352) & (!g1357) & (!g1362)) + ((g147) & (!g148) & (g1348) & (g1352) & (!g1357) & (g1362)) + ((g147) & (!g148) & (g1348) & (g1352) & (g1357) & (!g1362)) + ((g147) & (!g148) & (g1348) & (g1352) & (g1357) & (g1362)) + ((g147) & (g148) & (!g1348) & (!g1352) & (g1357) & (!g1362)) + ((g147) & (g148) & (!g1348) & (!g1352) & (g1357) & (g1362)) + ((g147) & (g148) & (!g1348) & (g1352) & (g1357) & (!g1362)) + ((g147) & (g148) & (!g1348) & (g1352) & (g1357) & (g1362)) + ((g147) & (g148) & (g1348) & (!g1352) & (g1357) & (!g1362)) + ((g147) & (g148) & (g1348) & (!g1352) & (g1357) & (g1362)) + ((g147) & (g148) & (g1348) & (g1352) & (g1357) & (!g1362)) + ((g147) & (g148) & (g1348) & (g1352) & (g1357) & (g1362)));
	assign g1364 = (((!g142) & (!sk[22]) & (!g1343) & (g1363)) + ((!g142) & (!sk[22]) & (g1343) & (!g1363)) + ((!g142) & (!sk[22]) & (g1343) & (g1363)) + ((!g142) & (sk[22]) & (!g1343) & (g1363)) + ((!g142) & (sk[22]) & (g1343) & (g1363)) + ((g142) & (!sk[22]) & (!g1343) & (g1363)) + ((g142) & (!sk[22]) & (g1343) & (!g1363)) + ((g142) & (!sk[22]) & (g1343) & (g1363)) + ((g142) & (sk[22]) & (g1343) & (!g1363)) + ((g142) & (sk[22]) & (g1343) & (g1363)));
	assign g4857 = (((!g2059) & (!sk[23]) & (!g2750) & (g1365)) + ((!g2059) & (!sk[23]) & (g2750) & (!g1365)) + ((!g2059) & (!sk[23]) & (g2750) & (g1365)) + ((!g2059) & (sk[23]) & (!g2750) & (g1365)) + ((!g2059) & (sk[23]) & (g2750) & (g1365)) + ((g2059) & (!sk[23]) & (!g2750) & (g1365)) + ((g2059) & (!sk[23]) & (g2750) & (!g1365)) + ((g2059) & (!sk[23]) & (g2750) & (g1365)) + ((g2059) & (sk[23]) & (g2750) & (!g1365)) + ((g2059) & (sk[23]) & (g2750) & (g1365)));
	assign g1366 = (((g1319) & (!sk[24]) & (!g916)) + ((g1319) & (!sk[24]) & (g916)) + ((g1319) & (sk[24]) & (!g916)));
	assign g1367 = (((!g126) & (!g1364) & (g1365) & (!g3823) & (!g1366) & (!g916)) + ((!g126) & (!g1364) & (g1365) & (!g3823) & (!g1366) & (g916)) + ((!g126) & (!g1364) & (g1365) & (!g3823) & (g1366) & (!g916)) + ((!g126) & (!g1364) & (g1365) & (!g3823) & (g1366) & (g916)) + ((!g126) & (!g1364) & (g1365) & (g3823) & (!g1366) & (!g916)) + ((!g126) & (!g1364) & (g1365) & (g3823) & (!g1366) & (g916)) + ((!g126) & (!g1364) & (g1365) & (g3823) & (g1366) & (!g916)) + ((!g126) & (!g1364) & (g1365) & (g3823) & (g1366) & (g916)) + ((!g126) & (g1364) & (g1365) & (!g3823) & (!g1366) & (!g916)) + ((!g126) & (g1364) & (g1365) & (!g3823) & (!g1366) & (g916)) + ((!g126) & (g1364) & (g1365) & (!g3823) & (g1366) & (!g916)) + ((!g126) & (g1364) & (g1365) & (!g3823) & (g1366) & (g916)) + ((!g126) & (g1364) & (g1365) & (g3823) & (!g1366) & (!g916)) + ((!g126) & (g1364) & (g1365) & (g3823) & (!g1366) & (g916)) + ((!g126) & (g1364) & (g1365) & (g3823) & (g1366) & (!g916)) + ((!g126) & (g1364) & (g1365) & (g3823) & (g1366) & (g916)) + ((g126) & (!g1364) & (!g1365) & (!g3823) & (!g1366) & (!g916)) + ((g126) & (!g1364) & (!g1365) & (!g3823) & (g1366) & (g916)) + ((g126) & (!g1364) & (!g1365) & (g3823) & (!g1366) & (g916)) + ((g126) & (!g1364) & (!g1365) & (g3823) & (g1366) & (g916)) + ((g126) & (!g1364) & (g1365) & (!g3823) & (!g1366) & (!g916)) + ((g126) & (!g1364) & (g1365) & (!g3823) & (g1366) & (g916)) + ((g126) & (!g1364) & (g1365) & (g3823) & (!g1366) & (g916)) + ((g126) & (!g1364) & (g1365) & (g3823) & (g1366) & (g916)) + ((g126) & (g1364) & (!g1365) & (!g3823) & (!g1366) & (g916)) + ((g126) & (g1364) & (!g1365) & (!g3823) & (g1366) & (!g916)) + ((g126) & (g1364) & (!g1365) & (g3823) & (!g1366) & (!g916)) + ((g126) & (g1364) & (!g1365) & (g3823) & (g1366) & (!g916)) + ((g126) & (g1364) & (g1365) & (!g3823) & (!g1366) & (g916)) + ((g126) & (g1364) & (g1365) & (!g3823) & (g1366) & (!g916)) + ((g126) & (g1364) & (g1365) & (g3823) & (!g1366) & (!g916)) + ((g126) & (g1364) & (g1365) & (g3823) & (g1366) & (!g916)));
	assign g4858 = (((!g2140) & (!sk[26]) & (!g3278) & (g1368)) + ((!g2140) & (!sk[26]) & (g3278) & (!g1368)) + ((!g2140) & (!sk[26]) & (g3278) & (g1368)) + ((!g2140) & (sk[26]) & (!g3278) & (g1368)) + ((!g2140) & (sk[26]) & (g3278) & (g1368)) + ((g2140) & (!sk[26]) & (!g3278) & (g1368)) + ((g2140) & (!sk[26]) & (g3278) & (!g1368)) + ((g2140) & (!sk[26]) & (g3278) & (g1368)) + ((g2140) & (sk[26]) & (g3278) & (!g1368)) + ((g2140) & (sk[26]) & (g3278) & (g1368)));
	assign g4859 = (((!g2142) & (!sk[27]) & (!g3278) & (g1369)) + ((!g2142) & (!sk[27]) & (g3278) & (!g1369)) + ((!g2142) & (!sk[27]) & (g3278) & (g1369)) + ((!g2142) & (sk[27]) & (!g3278) & (g1369)) + ((!g2142) & (sk[27]) & (g3278) & (g1369)) + ((g2142) & (!sk[27]) & (!g3278) & (g1369)) + ((g2142) & (!sk[27]) & (g3278) & (!g1369)) + ((g2142) & (!sk[27]) & (g3278) & (g1369)) + ((g2142) & (sk[27]) & (g3278) & (!g1369)) + ((g2142) & (sk[27]) & (g3278) & (g1369)));
	assign g4860 = (((!sk[28]) & (!g2144) & (!g3278) & (g1370)) + ((!sk[28]) & (!g2144) & (g3278) & (!g1370)) + ((!sk[28]) & (!g2144) & (g3278) & (g1370)) + ((!sk[28]) & (g2144) & (!g3278) & (g1370)) + ((!sk[28]) & (g2144) & (g3278) & (!g1370)) + ((!sk[28]) & (g2144) & (g3278) & (g1370)) + ((sk[28]) & (!g2144) & (!g3278) & (g1370)) + ((sk[28]) & (!g2144) & (g3278) & (g1370)) + ((sk[28]) & (g2144) & (g3278) & (!g1370)) + ((sk[28]) & (g2144) & (g3278) & (g1370)));
	assign g4861 = (((!sk[29]) & (!g2145) & (!g3278) & (g1371)) + ((!sk[29]) & (!g2145) & (g3278) & (!g1371)) + ((!sk[29]) & (!g2145) & (g3278) & (g1371)) + ((!sk[29]) & (g2145) & (!g3278) & (g1371)) + ((!sk[29]) & (g2145) & (g3278) & (!g1371)) + ((!sk[29]) & (g2145) & (g3278) & (g1371)) + ((sk[29]) & (!g2145) & (!g3278) & (g1371)) + ((sk[29]) & (!g2145) & (g3278) & (g1371)) + ((sk[29]) & (g2145) & (g3278) & (!g1371)) + ((sk[29]) & (g2145) & (g3278) & (g1371)));
	assign g1372 = (((!g1368) & (!g1369) & (!g1370) & (g1371) & (g147) & (g148)) + ((!g1368) & (!g1369) & (g1370) & (!g1371) & (!g147) & (g148)) + ((!g1368) & (!g1369) & (g1370) & (g1371) & (!g147) & (g148)) + ((!g1368) & (!g1369) & (g1370) & (g1371) & (g147) & (g148)) + ((!g1368) & (g1369) & (!g1370) & (!g1371) & (g147) & (!g148)) + ((!g1368) & (g1369) & (!g1370) & (g1371) & (g147) & (!g148)) + ((!g1368) & (g1369) & (!g1370) & (g1371) & (g147) & (g148)) + ((!g1368) & (g1369) & (g1370) & (!g1371) & (!g147) & (g148)) + ((!g1368) & (g1369) & (g1370) & (!g1371) & (g147) & (!g148)) + ((!g1368) & (g1369) & (g1370) & (g1371) & (!g147) & (g148)) + ((!g1368) & (g1369) & (g1370) & (g1371) & (g147) & (!g148)) + ((!g1368) & (g1369) & (g1370) & (g1371) & (g147) & (g148)) + ((g1368) & (!g1369) & (!g1370) & (!g1371) & (!g147) & (!g148)) + ((g1368) & (!g1369) & (!g1370) & (g1371) & (!g147) & (!g148)) + ((g1368) & (!g1369) & (!g1370) & (g1371) & (g147) & (g148)) + ((g1368) & (!g1369) & (g1370) & (!g1371) & (!g147) & (!g148)) + ((g1368) & (!g1369) & (g1370) & (!g1371) & (!g147) & (g148)) + ((g1368) & (!g1369) & (g1370) & (g1371) & (!g147) & (!g148)) + ((g1368) & (!g1369) & (g1370) & (g1371) & (!g147) & (g148)) + ((g1368) & (!g1369) & (g1370) & (g1371) & (g147) & (g148)) + ((g1368) & (g1369) & (!g1370) & (!g1371) & (!g147) & (!g148)) + ((g1368) & (g1369) & (!g1370) & (!g1371) & (g147) & (!g148)) + ((g1368) & (g1369) & (!g1370) & (g1371) & (!g147) & (!g148)) + ((g1368) & (g1369) & (!g1370) & (g1371) & (g147) & (!g148)) + ((g1368) & (g1369) & (!g1370) & (g1371) & (g147) & (g148)) + ((g1368) & (g1369) & (g1370) & (!g1371) & (!g147) & (!g148)) + ((g1368) & (g1369) & (g1370) & (!g1371) & (!g147) & (g148)) + ((g1368) & (g1369) & (g1370) & (!g1371) & (g147) & (!g148)) + ((g1368) & (g1369) & (g1370) & (g1371) & (!g147) & (!g148)) + ((g1368) & (g1369) & (g1370) & (g1371) & (!g147) & (g148)) + ((g1368) & (g1369) & (g1370) & (g1371) & (g147) & (!g148)) + ((g1368) & (g1369) & (g1370) & (g1371) & (g147) & (g148)));
	assign g4862 = (((!g2146) & (!sk[31]) & (!g3278) & (g1373)) + ((!g2146) & (!sk[31]) & (g3278) & (!g1373)) + ((!g2146) & (!sk[31]) & (g3278) & (g1373)) + ((!g2146) & (sk[31]) & (!g3278) & (g1373)) + ((!g2146) & (sk[31]) & (g3278) & (g1373)) + ((g2146) & (!sk[31]) & (!g3278) & (g1373)) + ((g2146) & (!sk[31]) & (g3278) & (!g1373)) + ((g2146) & (!sk[31]) & (g3278) & (g1373)) + ((g2146) & (sk[31]) & (g3278) & (!g1373)) + ((g2146) & (sk[31]) & (g3278) & (g1373)));
	assign g4863 = (((!g2148) & (!sk[32]) & (!g3278) & (g1374)) + ((!g2148) & (!sk[32]) & (g3278) & (!g1374)) + ((!g2148) & (!sk[32]) & (g3278) & (g1374)) + ((!g2148) & (sk[32]) & (!g3278) & (g1374)) + ((!g2148) & (sk[32]) & (g3278) & (g1374)) + ((g2148) & (!sk[32]) & (!g3278) & (g1374)) + ((g2148) & (!sk[32]) & (g3278) & (!g1374)) + ((g2148) & (!sk[32]) & (g3278) & (g1374)) + ((g2148) & (sk[32]) & (g3278) & (!g1374)) + ((g2148) & (sk[32]) & (g3278) & (g1374)));
	assign g4864 = (((!g2150) & (!sk[33]) & (!g3278) & (g1375)) + ((!g2150) & (!sk[33]) & (g3278) & (!g1375)) + ((!g2150) & (!sk[33]) & (g3278) & (g1375)) + ((!g2150) & (sk[33]) & (!g3278) & (g1375)) + ((!g2150) & (sk[33]) & (g3278) & (g1375)) + ((g2150) & (!sk[33]) & (!g3278) & (g1375)) + ((g2150) & (!sk[33]) & (g3278) & (!g1375)) + ((g2150) & (!sk[33]) & (g3278) & (g1375)) + ((g2150) & (sk[33]) & (g3278) & (!g1375)) + ((g2150) & (sk[33]) & (g3278) & (g1375)));
	assign g4865 = (((!g2151) & (!sk[34]) & (!g3278) & (g1376)) + ((!g2151) & (!sk[34]) & (g3278) & (!g1376)) + ((!g2151) & (!sk[34]) & (g3278) & (g1376)) + ((!g2151) & (sk[34]) & (!g3278) & (g1376)) + ((!g2151) & (sk[34]) & (g3278) & (g1376)) + ((g2151) & (!sk[34]) & (!g3278) & (g1376)) + ((g2151) & (!sk[34]) & (g3278) & (!g1376)) + ((g2151) & (!sk[34]) & (g3278) & (g1376)) + ((g2151) & (sk[34]) & (g3278) & (!g1376)) + ((g2151) & (sk[34]) & (g3278) & (g1376)));
	assign g1377 = (((!g1373) & (!g1374) & (!g1375) & (g1376) & (g147) & (g148)) + ((!g1373) & (!g1374) & (g1375) & (!g1376) & (!g147) & (g148)) + ((!g1373) & (!g1374) & (g1375) & (g1376) & (!g147) & (g148)) + ((!g1373) & (!g1374) & (g1375) & (g1376) & (g147) & (g148)) + ((!g1373) & (g1374) & (!g1375) & (!g1376) & (g147) & (!g148)) + ((!g1373) & (g1374) & (!g1375) & (g1376) & (g147) & (!g148)) + ((!g1373) & (g1374) & (!g1375) & (g1376) & (g147) & (g148)) + ((!g1373) & (g1374) & (g1375) & (!g1376) & (!g147) & (g148)) + ((!g1373) & (g1374) & (g1375) & (!g1376) & (g147) & (!g148)) + ((!g1373) & (g1374) & (g1375) & (g1376) & (!g147) & (g148)) + ((!g1373) & (g1374) & (g1375) & (g1376) & (g147) & (!g148)) + ((!g1373) & (g1374) & (g1375) & (g1376) & (g147) & (g148)) + ((g1373) & (!g1374) & (!g1375) & (!g1376) & (!g147) & (!g148)) + ((g1373) & (!g1374) & (!g1375) & (g1376) & (!g147) & (!g148)) + ((g1373) & (!g1374) & (!g1375) & (g1376) & (g147) & (g148)) + ((g1373) & (!g1374) & (g1375) & (!g1376) & (!g147) & (!g148)) + ((g1373) & (!g1374) & (g1375) & (!g1376) & (!g147) & (g148)) + ((g1373) & (!g1374) & (g1375) & (g1376) & (!g147) & (!g148)) + ((g1373) & (!g1374) & (g1375) & (g1376) & (!g147) & (g148)) + ((g1373) & (!g1374) & (g1375) & (g1376) & (g147) & (g148)) + ((g1373) & (g1374) & (!g1375) & (!g1376) & (!g147) & (!g148)) + ((g1373) & (g1374) & (!g1375) & (!g1376) & (g147) & (!g148)) + ((g1373) & (g1374) & (!g1375) & (g1376) & (!g147) & (!g148)) + ((g1373) & (g1374) & (!g1375) & (g1376) & (g147) & (!g148)) + ((g1373) & (g1374) & (!g1375) & (g1376) & (g147) & (g148)) + ((g1373) & (g1374) & (g1375) & (!g1376) & (!g147) & (!g148)) + ((g1373) & (g1374) & (g1375) & (!g1376) & (!g147) & (g148)) + ((g1373) & (g1374) & (g1375) & (!g1376) & (g147) & (!g148)) + ((g1373) & (g1374) & (g1375) & (g1376) & (!g147) & (!g148)) + ((g1373) & (g1374) & (g1375) & (g1376) & (!g147) & (g148)) + ((g1373) & (g1374) & (g1375) & (g1376) & (g147) & (!g148)) + ((g1373) & (g1374) & (g1375) & (g1376) & (g147) & (g148)));
	assign g4866 = (((!g2152) & (!sk[36]) & (!g3278) & (g1378)) + ((!g2152) & (!sk[36]) & (g3278) & (!g1378)) + ((!g2152) & (!sk[36]) & (g3278) & (g1378)) + ((!g2152) & (sk[36]) & (!g3278) & (g1378)) + ((!g2152) & (sk[36]) & (g3278) & (g1378)) + ((g2152) & (!sk[36]) & (!g3278) & (g1378)) + ((g2152) & (!sk[36]) & (g3278) & (!g1378)) + ((g2152) & (!sk[36]) & (g3278) & (g1378)) + ((g2152) & (sk[36]) & (g3278) & (!g1378)) + ((g2152) & (sk[36]) & (g3278) & (g1378)));
	assign g4867 = (((!g2153) & (!g3278) & (!sk[37]) & (g1379)) + ((!g2153) & (!g3278) & (sk[37]) & (g1379)) + ((!g2153) & (g3278) & (!sk[37]) & (!g1379)) + ((!g2153) & (g3278) & (!sk[37]) & (g1379)) + ((!g2153) & (g3278) & (sk[37]) & (g1379)) + ((g2153) & (!g3278) & (!sk[37]) & (g1379)) + ((g2153) & (g3278) & (!sk[37]) & (!g1379)) + ((g2153) & (g3278) & (!sk[37]) & (g1379)) + ((g2153) & (g3278) & (sk[37]) & (!g1379)) + ((g2153) & (g3278) & (sk[37]) & (g1379)));
	assign g4868 = (((!sk[38]) & (!g2155) & (!g3278) & (g1380)) + ((!sk[38]) & (!g2155) & (g3278) & (!g1380)) + ((!sk[38]) & (!g2155) & (g3278) & (g1380)) + ((!sk[38]) & (g2155) & (!g3278) & (g1380)) + ((!sk[38]) & (g2155) & (g3278) & (!g1380)) + ((!sk[38]) & (g2155) & (g3278) & (g1380)) + ((sk[38]) & (!g2155) & (!g3278) & (g1380)) + ((sk[38]) & (!g2155) & (g3278) & (g1380)) + ((sk[38]) & (g2155) & (g3278) & (!g1380)) + ((sk[38]) & (g2155) & (g3278) & (g1380)));
	assign g4869 = (((!g2157) & (!g3278) & (!sk[39]) & (g1381)) + ((!g2157) & (!g3278) & (sk[39]) & (g1381)) + ((!g2157) & (g3278) & (!sk[39]) & (!g1381)) + ((!g2157) & (g3278) & (!sk[39]) & (g1381)) + ((!g2157) & (g3278) & (sk[39]) & (g1381)) + ((g2157) & (!g3278) & (!sk[39]) & (g1381)) + ((g2157) & (g3278) & (!sk[39]) & (!g1381)) + ((g2157) & (g3278) & (!sk[39]) & (g1381)) + ((g2157) & (g3278) & (sk[39]) & (!g1381)) + ((g2157) & (g3278) & (sk[39]) & (g1381)));
	assign g1382 = (((!g1378) & (!g1379) & (!g1380) & (g1381) & (g147) & (g148)) + ((!g1378) & (!g1379) & (g1380) & (!g1381) & (!g147) & (g148)) + ((!g1378) & (!g1379) & (g1380) & (g1381) & (!g147) & (g148)) + ((!g1378) & (!g1379) & (g1380) & (g1381) & (g147) & (g148)) + ((!g1378) & (g1379) & (!g1380) & (!g1381) & (g147) & (!g148)) + ((!g1378) & (g1379) & (!g1380) & (g1381) & (g147) & (!g148)) + ((!g1378) & (g1379) & (!g1380) & (g1381) & (g147) & (g148)) + ((!g1378) & (g1379) & (g1380) & (!g1381) & (!g147) & (g148)) + ((!g1378) & (g1379) & (g1380) & (!g1381) & (g147) & (!g148)) + ((!g1378) & (g1379) & (g1380) & (g1381) & (!g147) & (g148)) + ((!g1378) & (g1379) & (g1380) & (g1381) & (g147) & (!g148)) + ((!g1378) & (g1379) & (g1380) & (g1381) & (g147) & (g148)) + ((g1378) & (!g1379) & (!g1380) & (!g1381) & (!g147) & (!g148)) + ((g1378) & (!g1379) & (!g1380) & (g1381) & (!g147) & (!g148)) + ((g1378) & (!g1379) & (!g1380) & (g1381) & (g147) & (g148)) + ((g1378) & (!g1379) & (g1380) & (!g1381) & (!g147) & (!g148)) + ((g1378) & (!g1379) & (g1380) & (!g1381) & (!g147) & (g148)) + ((g1378) & (!g1379) & (g1380) & (g1381) & (!g147) & (!g148)) + ((g1378) & (!g1379) & (g1380) & (g1381) & (!g147) & (g148)) + ((g1378) & (!g1379) & (g1380) & (g1381) & (g147) & (g148)) + ((g1378) & (g1379) & (!g1380) & (!g1381) & (!g147) & (!g148)) + ((g1378) & (g1379) & (!g1380) & (!g1381) & (g147) & (!g148)) + ((g1378) & (g1379) & (!g1380) & (g1381) & (!g147) & (!g148)) + ((g1378) & (g1379) & (!g1380) & (g1381) & (g147) & (!g148)) + ((g1378) & (g1379) & (!g1380) & (g1381) & (g147) & (g148)) + ((g1378) & (g1379) & (g1380) & (!g1381) & (!g147) & (!g148)) + ((g1378) & (g1379) & (g1380) & (!g1381) & (!g147) & (g148)) + ((g1378) & (g1379) & (g1380) & (!g1381) & (g147) & (!g148)) + ((g1378) & (g1379) & (g1380) & (g1381) & (!g147) & (!g148)) + ((g1378) & (g1379) & (g1380) & (g1381) & (!g147) & (g148)) + ((g1378) & (g1379) & (g1380) & (g1381) & (g147) & (!g148)) + ((g1378) & (g1379) & (g1380) & (g1381) & (g147) & (g148)));
	assign g4870 = (((!sk[41]) & (!g2158) & (!g3278) & (g1383)) + ((!sk[41]) & (!g2158) & (g3278) & (!g1383)) + ((!sk[41]) & (!g2158) & (g3278) & (g1383)) + ((!sk[41]) & (g2158) & (!g3278) & (g1383)) + ((!sk[41]) & (g2158) & (g3278) & (!g1383)) + ((!sk[41]) & (g2158) & (g3278) & (g1383)) + ((sk[41]) & (!g2158) & (!g3278) & (g1383)) + ((sk[41]) & (!g2158) & (g3278) & (g1383)) + ((sk[41]) & (g2158) & (g3278) & (!g1383)) + ((sk[41]) & (g2158) & (g3278) & (g1383)));
	assign g4871 = (((!g2159) & (!sk[42]) & (!g3278) & (g1384)) + ((!g2159) & (!sk[42]) & (g3278) & (!g1384)) + ((!g2159) & (!sk[42]) & (g3278) & (g1384)) + ((!g2159) & (sk[42]) & (!g3278) & (g1384)) + ((!g2159) & (sk[42]) & (g3278) & (g1384)) + ((g2159) & (!sk[42]) & (!g3278) & (g1384)) + ((g2159) & (!sk[42]) & (g3278) & (!g1384)) + ((g2159) & (!sk[42]) & (g3278) & (g1384)) + ((g2159) & (sk[42]) & (g3278) & (!g1384)) + ((g2159) & (sk[42]) & (g3278) & (g1384)));
	assign g4872 = (((!g2160) & (!sk[43]) & (!g3278) & (g1385)) + ((!g2160) & (!sk[43]) & (g3278) & (!g1385)) + ((!g2160) & (!sk[43]) & (g3278) & (g1385)) + ((!g2160) & (sk[43]) & (!g3278) & (g1385)) + ((!g2160) & (sk[43]) & (g3278) & (g1385)) + ((g2160) & (!sk[43]) & (!g3278) & (g1385)) + ((g2160) & (!sk[43]) & (g3278) & (!g1385)) + ((g2160) & (!sk[43]) & (g3278) & (g1385)) + ((g2160) & (sk[43]) & (g3278) & (!g1385)) + ((g2160) & (sk[43]) & (g3278) & (g1385)));
	assign g4873 = (((!g2161) & (!sk[44]) & (!g3278) & (g1386)) + ((!g2161) & (!sk[44]) & (g3278) & (!g1386)) + ((!g2161) & (!sk[44]) & (g3278) & (g1386)) + ((!g2161) & (sk[44]) & (!g3278) & (g1386)) + ((!g2161) & (sk[44]) & (g3278) & (g1386)) + ((g2161) & (!sk[44]) & (!g3278) & (g1386)) + ((g2161) & (!sk[44]) & (g3278) & (!g1386)) + ((g2161) & (!sk[44]) & (g3278) & (g1386)) + ((g2161) & (sk[44]) & (g3278) & (!g1386)) + ((g2161) & (sk[44]) & (g3278) & (g1386)));
	assign g1387 = (((!g1383) & (!g1384) & (!g1385) & (g1386) & (g147) & (g148)) + ((!g1383) & (!g1384) & (g1385) & (!g1386) & (!g147) & (g148)) + ((!g1383) & (!g1384) & (g1385) & (g1386) & (!g147) & (g148)) + ((!g1383) & (!g1384) & (g1385) & (g1386) & (g147) & (g148)) + ((!g1383) & (g1384) & (!g1385) & (!g1386) & (g147) & (!g148)) + ((!g1383) & (g1384) & (!g1385) & (g1386) & (g147) & (!g148)) + ((!g1383) & (g1384) & (!g1385) & (g1386) & (g147) & (g148)) + ((!g1383) & (g1384) & (g1385) & (!g1386) & (!g147) & (g148)) + ((!g1383) & (g1384) & (g1385) & (!g1386) & (g147) & (!g148)) + ((!g1383) & (g1384) & (g1385) & (g1386) & (!g147) & (g148)) + ((!g1383) & (g1384) & (g1385) & (g1386) & (g147) & (!g148)) + ((!g1383) & (g1384) & (g1385) & (g1386) & (g147) & (g148)) + ((g1383) & (!g1384) & (!g1385) & (!g1386) & (!g147) & (!g148)) + ((g1383) & (!g1384) & (!g1385) & (g1386) & (!g147) & (!g148)) + ((g1383) & (!g1384) & (!g1385) & (g1386) & (g147) & (g148)) + ((g1383) & (!g1384) & (g1385) & (!g1386) & (!g147) & (!g148)) + ((g1383) & (!g1384) & (g1385) & (!g1386) & (!g147) & (g148)) + ((g1383) & (!g1384) & (g1385) & (g1386) & (!g147) & (!g148)) + ((g1383) & (!g1384) & (g1385) & (g1386) & (!g147) & (g148)) + ((g1383) & (!g1384) & (g1385) & (g1386) & (g147) & (g148)) + ((g1383) & (g1384) & (!g1385) & (!g1386) & (!g147) & (!g148)) + ((g1383) & (g1384) & (!g1385) & (!g1386) & (g147) & (!g148)) + ((g1383) & (g1384) & (!g1385) & (g1386) & (!g147) & (!g148)) + ((g1383) & (g1384) & (!g1385) & (g1386) & (g147) & (!g148)) + ((g1383) & (g1384) & (!g1385) & (g1386) & (g147) & (g148)) + ((g1383) & (g1384) & (g1385) & (!g1386) & (!g147) & (!g148)) + ((g1383) & (g1384) & (g1385) & (!g1386) & (!g147) & (g148)) + ((g1383) & (g1384) & (g1385) & (!g1386) & (g147) & (!g148)) + ((g1383) & (g1384) & (g1385) & (g1386) & (!g147) & (!g148)) + ((g1383) & (g1384) & (g1385) & (g1386) & (!g147) & (g148)) + ((g1383) & (g1384) & (g1385) & (g1386) & (g147) & (!g148)) + ((g1383) & (g1384) & (g1385) & (g1386) & (g147) & (g148)));
	assign g1388 = (((!g1372) & (!g1377) & (!g1382) & (g1387) & (g165) & (g166)) + ((!g1372) & (!g1377) & (g1382) & (!g1387) & (!g165) & (g166)) + ((!g1372) & (!g1377) & (g1382) & (g1387) & (!g165) & (g166)) + ((!g1372) & (!g1377) & (g1382) & (g1387) & (g165) & (g166)) + ((!g1372) & (g1377) & (!g1382) & (!g1387) & (g165) & (!g166)) + ((!g1372) & (g1377) & (!g1382) & (g1387) & (g165) & (!g166)) + ((!g1372) & (g1377) & (!g1382) & (g1387) & (g165) & (g166)) + ((!g1372) & (g1377) & (g1382) & (!g1387) & (!g165) & (g166)) + ((!g1372) & (g1377) & (g1382) & (!g1387) & (g165) & (!g166)) + ((!g1372) & (g1377) & (g1382) & (g1387) & (!g165) & (g166)) + ((!g1372) & (g1377) & (g1382) & (g1387) & (g165) & (!g166)) + ((!g1372) & (g1377) & (g1382) & (g1387) & (g165) & (g166)) + ((g1372) & (!g1377) & (!g1382) & (!g1387) & (!g165) & (!g166)) + ((g1372) & (!g1377) & (!g1382) & (g1387) & (!g165) & (!g166)) + ((g1372) & (!g1377) & (!g1382) & (g1387) & (g165) & (g166)) + ((g1372) & (!g1377) & (g1382) & (!g1387) & (!g165) & (!g166)) + ((g1372) & (!g1377) & (g1382) & (!g1387) & (!g165) & (g166)) + ((g1372) & (!g1377) & (g1382) & (g1387) & (!g165) & (!g166)) + ((g1372) & (!g1377) & (g1382) & (g1387) & (!g165) & (g166)) + ((g1372) & (!g1377) & (g1382) & (g1387) & (g165) & (g166)) + ((g1372) & (g1377) & (!g1382) & (!g1387) & (!g165) & (!g166)) + ((g1372) & (g1377) & (!g1382) & (!g1387) & (g165) & (!g166)) + ((g1372) & (g1377) & (!g1382) & (g1387) & (!g165) & (!g166)) + ((g1372) & (g1377) & (!g1382) & (g1387) & (g165) & (!g166)) + ((g1372) & (g1377) & (!g1382) & (g1387) & (g165) & (g166)) + ((g1372) & (g1377) & (g1382) & (!g1387) & (!g165) & (!g166)) + ((g1372) & (g1377) & (g1382) & (!g1387) & (!g165) & (g166)) + ((g1372) & (g1377) & (g1382) & (!g1387) & (g165) & (!g166)) + ((g1372) & (g1377) & (g1382) & (g1387) & (!g165) & (!g166)) + ((g1372) & (g1377) & (g1382) & (g1387) & (!g165) & (g166)) + ((g1372) & (g1377) & (g1382) & (g1387) & (g165) & (!g166)) + ((g1372) & (g1377) & (g1382) & (g1387) & (g165) & (g166)));
	assign g4874 = (((!g2173) & (!g3278) & (!sk[47]) & (g1389)) + ((!g2173) & (!g3278) & (sk[47]) & (g1389)) + ((!g2173) & (g3278) & (!sk[47]) & (!g1389)) + ((!g2173) & (g3278) & (!sk[47]) & (g1389)) + ((!g2173) & (g3278) & (sk[47]) & (g1389)) + ((g2173) & (!g3278) & (!sk[47]) & (g1389)) + ((g2173) & (g3278) & (!sk[47]) & (!g1389)) + ((g2173) & (g3278) & (!sk[47]) & (g1389)) + ((g2173) & (g3278) & (sk[47]) & (!g1389)) + ((g2173) & (g3278) & (sk[47]) & (g1389)));
	assign g4875 = (((!g2174) & (!sk[48]) & (!g3278) & (g1390)) + ((!g2174) & (!sk[48]) & (g3278) & (!g1390)) + ((!g2174) & (!sk[48]) & (g3278) & (g1390)) + ((!g2174) & (sk[48]) & (!g3278) & (g1390)) + ((!g2174) & (sk[48]) & (g3278) & (g1390)) + ((g2174) & (!sk[48]) & (!g3278) & (g1390)) + ((g2174) & (!sk[48]) & (g3278) & (!g1390)) + ((g2174) & (!sk[48]) & (g3278) & (g1390)) + ((g2174) & (sk[48]) & (g3278) & (!g1390)) + ((g2174) & (sk[48]) & (g3278) & (g1390)));
	assign g4876 = (((!sk[49]) & (!g2175) & (!g3278) & (g1391)) + ((!sk[49]) & (!g2175) & (g3278) & (!g1391)) + ((!sk[49]) & (!g2175) & (g3278) & (g1391)) + ((!sk[49]) & (g2175) & (!g3278) & (g1391)) + ((!sk[49]) & (g2175) & (g3278) & (!g1391)) + ((!sk[49]) & (g2175) & (g3278) & (g1391)) + ((sk[49]) & (!g2175) & (!g3278) & (g1391)) + ((sk[49]) & (!g2175) & (g3278) & (g1391)) + ((sk[49]) & (g2175) & (g3278) & (!g1391)) + ((sk[49]) & (g2175) & (g3278) & (g1391)));
	assign g4877 = (((!sk[50]) & (!g2176) & (!g3278) & (g1392)) + ((!sk[50]) & (!g2176) & (g3278) & (!g1392)) + ((!sk[50]) & (!g2176) & (g3278) & (g1392)) + ((!sk[50]) & (g2176) & (!g3278) & (g1392)) + ((!sk[50]) & (g2176) & (g3278) & (!g1392)) + ((!sk[50]) & (g2176) & (g3278) & (g1392)) + ((sk[50]) & (!g2176) & (!g3278) & (g1392)) + ((sk[50]) & (!g2176) & (g3278) & (g1392)) + ((sk[50]) & (g2176) & (g3278) & (!g1392)) + ((sk[50]) & (g2176) & (g3278) & (g1392)));
	assign g1393 = (((!g1389) & (!g1390) & (!g1391) & (g1392) & (g165) & (g166)) + ((!g1389) & (!g1390) & (g1391) & (!g1392) & (!g165) & (g166)) + ((!g1389) & (!g1390) & (g1391) & (g1392) & (!g165) & (g166)) + ((!g1389) & (!g1390) & (g1391) & (g1392) & (g165) & (g166)) + ((!g1389) & (g1390) & (!g1391) & (!g1392) & (g165) & (!g166)) + ((!g1389) & (g1390) & (!g1391) & (g1392) & (g165) & (!g166)) + ((!g1389) & (g1390) & (!g1391) & (g1392) & (g165) & (g166)) + ((!g1389) & (g1390) & (g1391) & (!g1392) & (!g165) & (g166)) + ((!g1389) & (g1390) & (g1391) & (!g1392) & (g165) & (!g166)) + ((!g1389) & (g1390) & (g1391) & (g1392) & (!g165) & (g166)) + ((!g1389) & (g1390) & (g1391) & (g1392) & (g165) & (!g166)) + ((!g1389) & (g1390) & (g1391) & (g1392) & (g165) & (g166)) + ((g1389) & (!g1390) & (!g1391) & (!g1392) & (!g165) & (!g166)) + ((g1389) & (!g1390) & (!g1391) & (g1392) & (!g165) & (!g166)) + ((g1389) & (!g1390) & (!g1391) & (g1392) & (g165) & (g166)) + ((g1389) & (!g1390) & (g1391) & (!g1392) & (!g165) & (!g166)) + ((g1389) & (!g1390) & (g1391) & (!g1392) & (!g165) & (g166)) + ((g1389) & (!g1390) & (g1391) & (g1392) & (!g165) & (!g166)) + ((g1389) & (!g1390) & (g1391) & (g1392) & (!g165) & (g166)) + ((g1389) & (!g1390) & (g1391) & (g1392) & (g165) & (g166)) + ((g1389) & (g1390) & (!g1391) & (!g1392) & (!g165) & (!g166)) + ((g1389) & (g1390) & (!g1391) & (!g1392) & (g165) & (!g166)) + ((g1389) & (g1390) & (!g1391) & (g1392) & (!g165) & (!g166)) + ((g1389) & (g1390) & (!g1391) & (g1392) & (g165) & (!g166)) + ((g1389) & (g1390) & (!g1391) & (g1392) & (g165) & (g166)) + ((g1389) & (g1390) & (g1391) & (!g1392) & (!g165) & (!g166)) + ((g1389) & (g1390) & (g1391) & (!g1392) & (!g165) & (g166)) + ((g1389) & (g1390) & (g1391) & (!g1392) & (g165) & (!g166)) + ((g1389) & (g1390) & (g1391) & (g1392) & (!g165) & (!g166)) + ((g1389) & (g1390) & (g1391) & (g1392) & (!g165) & (g166)) + ((g1389) & (g1390) & (g1391) & (g1392) & (g165) & (!g166)) + ((g1389) & (g1390) & (g1391) & (g1392) & (g165) & (g166)));
	assign g4878 = (((!g2177) & (!sk[52]) & (!g3278) & (g1394)) + ((!g2177) & (!sk[52]) & (g3278) & (!g1394)) + ((!g2177) & (!sk[52]) & (g3278) & (g1394)) + ((!g2177) & (sk[52]) & (!g3278) & (g1394)) + ((!g2177) & (sk[52]) & (g3278) & (g1394)) + ((g2177) & (!sk[52]) & (!g3278) & (g1394)) + ((g2177) & (!sk[52]) & (g3278) & (!g1394)) + ((g2177) & (!sk[52]) & (g3278) & (g1394)) + ((g2177) & (sk[52]) & (g3278) & (!g1394)) + ((g2177) & (sk[52]) & (g3278) & (g1394)));
	assign g4879 = (((!sk[53]) & (!g2178) & (!g3278) & (g1395)) + ((!sk[53]) & (!g2178) & (g3278) & (!g1395)) + ((!sk[53]) & (!g2178) & (g3278) & (g1395)) + ((!sk[53]) & (g2178) & (!g3278) & (g1395)) + ((!sk[53]) & (g2178) & (g3278) & (!g1395)) + ((!sk[53]) & (g2178) & (g3278) & (g1395)) + ((sk[53]) & (!g2178) & (!g3278) & (g1395)) + ((sk[53]) & (!g2178) & (g3278) & (g1395)) + ((sk[53]) & (g2178) & (g3278) & (!g1395)) + ((sk[53]) & (g2178) & (g3278) & (g1395)));
	assign g4880 = (((!g2179) & (!g3278) & (!sk[54]) & (g1396)) + ((!g2179) & (!g3278) & (sk[54]) & (g1396)) + ((!g2179) & (g3278) & (!sk[54]) & (!g1396)) + ((!g2179) & (g3278) & (!sk[54]) & (g1396)) + ((!g2179) & (g3278) & (sk[54]) & (g1396)) + ((g2179) & (!g3278) & (!sk[54]) & (g1396)) + ((g2179) & (g3278) & (!sk[54]) & (!g1396)) + ((g2179) & (g3278) & (!sk[54]) & (g1396)) + ((g2179) & (g3278) & (sk[54]) & (!g1396)) + ((g2179) & (g3278) & (sk[54]) & (g1396)));
	assign g1397 = (((!g165) & (!g166) & (!g1394) & (g1395) & (!sk[55]) & (!g1396)) + ((!g165) & (!g166) & (!g1394) & (g1395) & (!sk[55]) & (g1396)) + ((!g165) & (!g166) & (g1394) & (!g1395) & (!sk[55]) & (!g1396)) + ((!g165) & (!g166) & (g1394) & (!g1395) & (!sk[55]) & (g1396)) + ((!g165) & (!g166) & (g1394) & (g1395) & (!sk[55]) & (!g1396)) + ((!g165) & (!g166) & (g1394) & (g1395) & (!sk[55]) & (g1396)) + ((!g165) & (g166) & (!g1394) & (!g1395) & (!sk[55]) & (!g1396)) + ((!g165) & (g166) & (!g1394) & (!g1395) & (!sk[55]) & (g1396)) + ((!g165) & (g166) & (!g1394) & (!g1395) & (sk[55]) & (g1396)) + ((!g165) & (g166) & (!g1394) & (g1395) & (!sk[55]) & (!g1396)) + ((!g165) & (g166) & (!g1394) & (g1395) & (!sk[55]) & (g1396)) + ((!g165) & (g166) & (!g1394) & (g1395) & (sk[55]) & (g1396)) + ((!g165) & (g166) & (g1394) & (!g1395) & (!sk[55]) & (!g1396)) + ((!g165) & (g166) & (g1394) & (!g1395) & (!sk[55]) & (g1396)) + ((!g165) & (g166) & (g1394) & (!g1395) & (sk[55]) & (g1396)) + ((!g165) & (g166) & (g1394) & (g1395) & (!sk[55]) & (!g1396)) + ((!g165) & (g166) & (g1394) & (g1395) & (!sk[55]) & (g1396)) + ((!g165) & (g166) & (g1394) & (g1395) & (sk[55]) & (g1396)) + ((g165) & (!g166) & (!g1394) & (g1395) & (!sk[55]) & (!g1396)) + ((g165) & (!g166) & (!g1394) & (g1395) & (!sk[55]) & (g1396)) + ((g165) & (!g166) & (g1394) & (!g1395) & (!sk[55]) & (!g1396)) + ((g165) & (!g166) & (g1394) & (!g1395) & (!sk[55]) & (g1396)) + ((g165) & (!g166) & (g1394) & (!g1395) & (sk[55]) & (!g1396)) + ((g165) & (!g166) & (g1394) & (!g1395) & (sk[55]) & (g1396)) + ((g165) & (!g166) & (g1394) & (g1395) & (!sk[55]) & (!g1396)) + ((g165) & (!g166) & (g1394) & (g1395) & (!sk[55]) & (g1396)) + ((g165) & (!g166) & (g1394) & (g1395) & (sk[55]) & (!g1396)) + ((g165) & (!g166) & (g1394) & (g1395) & (sk[55]) & (g1396)) + ((g165) & (g166) & (!g1394) & (!g1395) & (!sk[55]) & (!g1396)) + ((g165) & (g166) & (!g1394) & (!g1395) & (!sk[55]) & (g1396)) + ((g165) & (g166) & (!g1394) & (g1395) & (!sk[55]) & (!g1396)) + ((g165) & (g166) & (!g1394) & (g1395) & (!sk[55]) & (g1396)) + ((g165) & (g166) & (!g1394) & (g1395) & (sk[55]) & (!g1396)) + ((g165) & (g166) & (!g1394) & (g1395) & (sk[55]) & (g1396)) + ((g165) & (g166) & (g1394) & (!g1395) & (!sk[55]) & (!g1396)) + ((g165) & (g166) & (g1394) & (!g1395) & (!sk[55]) & (g1396)) + ((g165) & (g166) & (g1394) & (g1395) & (!sk[55]) & (!g1396)) + ((g165) & (g166) & (g1394) & (g1395) & (!sk[55]) & (g1396)) + ((g165) & (g166) & (g1394) & (g1395) & (sk[55]) & (!g1396)) + ((g165) & (g166) & (g1394) & (g1395) & (sk[55]) & (g1396)));
	assign g4881 = (((!g2162) & (!g3278) & (!sk[56]) & (g1398)) + ((!g2162) & (!g3278) & (sk[56]) & (g1398)) + ((!g2162) & (g3278) & (!sk[56]) & (!g1398)) + ((!g2162) & (g3278) & (!sk[56]) & (g1398)) + ((!g2162) & (g3278) & (sk[56]) & (g1398)) + ((g2162) & (!g3278) & (!sk[56]) & (g1398)) + ((g2162) & (g3278) & (!sk[56]) & (!g1398)) + ((g2162) & (g3278) & (!sk[56]) & (g1398)) + ((g2162) & (g3278) & (sk[56]) & (!g1398)) + ((g2162) & (g3278) & (sk[56]) & (g1398)));
	assign g4882 = (((!g2164) & (!sk[57]) & (!g3278) & (g1399)) + ((!g2164) & (!sk[57]) & (g3278) & (!g1399)) + ((!g2164) & (!sk[57]) & (g3278) & (g1399)) + ((!g2164) & (sk[57]) & (!g3278) & (g1399)) + ((!g2164) & (sk[57]) & (g3278) & (g1399)) + ((g2164) & (!sk[57]) & (!g3278) & (g1399)) + ((g2164) & (!sk[57]) & (g3278) & (!g1399)) + ((g2164) & (!sk[57]) & (g3278) & (g1399)) + ((g2164) & (sk[57]) & (g3278) & (!g1399)) + ((g2164) & (sk[57]) & (g3278) & (g1399)));
	assign g4883 = (((!g2166) & (!sk[58]) & (!g3278) & (g1400)) + ((!g2166) & (!sk[58]) & (g3278) & (!g1400)) + ((!g2166) & (!sk[58]) & (g3278) & (g1400)) + ((!g2166) & (sk[58]) & (!g3278) & (g1400)) + ((!g2166) & (sk[58]) & (g3278) & (g1400)) + ((g2166) & (!sk[58]) & (!g3278) & (g1400)) + ((g2166) & (!sk[58]) & (g3278) & (!g1400)) + ((g2166) & (!sk[58]) & (g3278) & (g1400)) + ((g2166) & (sk[58]) & (g3278) & (!g1400)) + ((g2166) & (sk[58]) & (g3278) & (g1400)));
	assign g4884 = (((!g2168) & (!g3278) & (!sk[59]) & (g1401)) + ((!g2168) & (!g3278) & (sk[59]) & (g1401)) + ((!g2168) & (g3278) & (!sk[59]) & (!g1401)) + ((!g2168) & (g3278) & (!sk[59]) & (g1401)) + ((!g2168) & (g3278) & (sk[59]) & (g1401)) + ((g2168) & (!g3278) & (!sk[59]) & (g1401)) + ((g2168) & (g3278) & (!sk[59]) & (!g1401)) + ((g2168) & (g3278) & (!sk[59]) & (g1401)) + ((g2168) & (g3278) & (sk[59]) & (!g1401)) + ((g2168) & (g3278) & (sk[59]) & (g1401)));
	assign g1402 = (((!g1398) & (!g1399) & (!g1400) & (g1401) & (g165) & (g166)) + ((!g1398) & (!g1399) & (g1400) & (!g1401) & (!g165) & (g166)) + ((!g1398) & (!g1399) & (g1400) & (g1401) & (!g165) & (g166)) + ((!g1398) & (!g1399) & (g1400) & (g1401) & (g165) & (g166)) + ((!g1398) & (g1399) & (!g1400) & (!g1401) & (g165) & (!g166)) + ((!g1398) & (g1399) & (!g1400) & (g1401) & (g165) & (!g166)) + ((!g1398) & (g1399) & (!g1400) & (g1401) & (g165) & (g166)) + ((!g1398) & (g1399) & (g1400) & (!g1401) & (!g165) & (g166)) + ((!g1398) & (g1399) & (g1400) & (!g1401) & (g165) & (!g166)) + ((!g1398) & (g1399) & (g1400) & (g1401) & (!g165) & (g166)) + ((!g1398) & (g1399) & (g1400) & (g1401) & (g165) & (!g166)) + ((!g1398) & (g1399) & (g1400) & (g1401) & (g165) & (g166)) + ((g1398) & (!g1399) & (!g1400) & (!g1401) & (!g165) & (!g166)) + ((g1398) & (!g1399) & (!g1400) & (g1401) & (!g165) & (!g166)) + ((g1398) & (!g1399) & (!g1400) & (g1401) & (g165) & (g166)) + ((g1398) & (!g1399) & (g1400) & (!g1401) & (!g165) & (!g166)) + ((g1398) & (!g1399) & (g1400) & (!g1401) & (!g165) & (g166)) + ((g1398) & (!g1399) & (g1400) & (g1401) & (!g165) & (!g166)) + ((g1398) & (!g1399) & (g1400) & (g1401) & (!g165) & (g166)) + ((g1398) & (!g1399) & (g1400) & (g1401) & (g165) & (g166)) + ((g1398) & (g1399) & (!g1400) & (!g1401) & (!g165) & (!g166)) + ((g1398) & (g1399) & (!g1400) & (!g1401) & (g165) & (!g166)) + ((g1398) & (g1399) & (!g1400) & (g1401) & (!g165) & (!g166)) + ((g1398) & (g1399) & (!g1400) & (g1401) & (g165) & (!g166)) + ((g1398) & (g1399) & (!g1400) & (g1401) & (g165) & (g166)) + ((g1398) & (g1399) & (g1400) & (!g1401) & (!g165) & (!g166)) + ((g1398) & (g1399) & (g1400) & (!g1401) & (!g165) & (g166)) + ((g1398) & (g1399) & (g1400) & (!g1401) & (g165) & (!g166)) + ((g1398) & (g1399) & (g1400) & (g1401) & (!g165) & (!g166)) + ((g1398) & (g1399) & (g1400) & (g1401) & (!g165) & (g166)) + ((g1398) & (g1399) & (g1400) & (g1401) & (g165) & (!g166)) + ((g1398) & (g1399) & (g1400) & (g1401) & (g165) & (g166)));
	assign g4885 = (((!sk[61]) & (!g2169) & (!g3278) & (g1403)) + ((!sk[61]) & (!g2169) & (g3278) & (!g1403)) + ((!sk[61]) & (!g2169) & (g3278) & (g1403)) + ((!sk[61]) & (g2169) & (!g3278) & (g1403)) + ((!sk[61]) & (g2169) & (g3278) & (!g1403)) + ((!sk[61]) & (g2169) & (g3278) & (g1403)) + ((sk[61]) & (!g2169) & (!g3278) & (g1403)) + ((sk[61]) & (!g2169) & (g3278) & (g1403)) + ((sk[61]) & (g2169) & (g3278) & (!g1403)) + ((sk[61]) & (g2169) & (g3278) & (g1403)));
	assign g4886 = (((!g2170) & (!sk[62]) & (!g3278) & (g1404)) + ((!g2170) & (!sk[62]) & (g3278) & (!g1404)) + ((!g2170) & (!sk[62]) & (g3278) & (g1404)) + ((!g2170) & (sk[62]) & (!g3278) & (g1404)) + ((!g2170) & (sk[62]) & (g3278) & (g1404)) + ((g2170) & (!sk[62]) & (!g3278) & (g1404)) + ((g2170) & (!sk[62]) & (g3278) & (!g1404)) + ((g2170) & (!sk[62]) & (g3278) & (g1404)) + ((g2170) & (sk[62]) & (g3278) & (!g1404)) + ((g2170) & (sk[62]) & (g3278) & (g1404)));
	assign g4887 = (((!sk[63]) & (!g2171) & (!g3278) & (g1405)) + ((!sk[63]) & (!g2171) & (g3278) & (!g1405)) + ((!sk[63]) & (!g2171) & (g3278) & (g1405)) + ((!sk[63]) & (g2171) & (!g3278) & (g1405)) + ((!sk[63]) & (g2171) & (g3278) & (!g1405)) + ((!sk[63]) & (g2171) & (g3278) & (g1405)) + ((sk[63]) & (!g2171) & (!g3278) & (g1405)) + ((sk[63]) & (!g2171) & (g3278) & (g1405)) + ((sk[63]) & (g2171) & (g3278) & (!g1405)) + ((sk[63]) & (g2171) & (g3278) & (g1405)));
	assign g4888 = (((!sk[64]) & (!g2172) & (!g3278) & (g1406)) + ((!sk[64]) & (!g2172) & (g3278) & (!g1406)) + ((!sk[64]) & (!g2172) & (g3278) & (g1406)) + ((!sk[64]) & (g2172) & (!g3278) & (g1406)) + ((!sk[64]) & (g2172) & (g3278) & (!g1406)) + ((!sk[64]) & (g2172) & (g3278) & (g1406)) + ((sk[64]) & (!g2172) & (!g3278) & (g1406)) + ((sk[64]) & (!g2172) & (g3278) & (g1406)) + ((sk[64]) & (g2172) & (g3278) & (!g1406)) + ((sk[64]) & (g2172) & (g3278) & (g1406)));
	assign g1407 = (((!g1403) & (!g1404) & (!g1405) & (g1406) & (g165) & (g166)) + ((!g1403) & (!g1404) & (g1405) & (!g1406) & (!g165) & (g166)) + ((!g1403) & (!g1404) & (g1405) & (g1406) & (!g165) & (g166)) + ((!g1403) & (!g1404) & (g1405) & (g1406) & (g165) & (g166)) + ((!g1403) & (g1404) & (!g1405) & (!g1406) & (g165) & (!g166)) + ((!g1403) & (g1404) & (!g1405) & (g1406) & (g165) & (!g166)) + ((!g1403) & (g1404) & (!g1405) & (g1406) & (g165) & (g166)) + ((!g1403) & (g1404) & (g1405) & (!g1406) & (!g165) & (g166)) + ((!g1403) & (g1404) & (g1405) & (!g1406) & (g165) & (!g166)) + ((!g1403) & (g1404) & (g1405) & (g1406) & (!g165) & (g166)) + ((!g1403) & (g1404) & (g1405) & (g1406) & (g165) & (!g166)) + ((!g1403) & (g1404) & (g1405) & (g1406) & (g165) & (g166)) + ((g1403) & (!g1404) & (!g1405) & (!g1406) & (!g165) & (!g166)) + ((g1403) & (!g1404) & (!g1405) & (g1406) & (!g165) & (!g166)) + ((g1403) & (!g1404) & (!g1405) & (g1406) & (g165) & (g166)) + ((g1403) & (!g1404) & (g1405) & (!g1406) & (!g165) & (!g166)) + ((g1403) & (!g1404) & (g1405) & (!g1406) & (!g165) & (g166)) + ((g1403) & (!g1404) & (g1405) & (g1406) & (!g165) & (!g166)) + ((g1403) & (!g1404) & (g1405) & (g1406) & (!g165) & (g166)) + ((g1403) & (!g1404) & (g1405) & (g1406) & (g165) & (g166)) + ((g1403) & (g1404) & (!g1405) & (!g1406) & (!g165) & (!g166)) + ((g1403) & (g1404) & (!g1405) & (!g1406) & (g165) & (!g166)) + ((g1403) & (g1404) & (!g1405) & (g1406) & (!g165) & (!g166)) + ((g1403) & (g1404) & (!g1405) & (g1406) & (g165) & (!g166)) + ((g1403) & (g1404) & (!g1405) & (g1406) & (g165) & (g166)) + ((g1403) & (g1404) & (g1405) & (!g1406) & (!g165) & (!g166)) + ((g1403) & (g1404) & (g1405) & (!g1406) & (!g165) & (g166)) + ((g1403) & (g1404) & (g1405) & (!g1406) & (g165) & (!g166)) + ((g1403) & (g1404) & (g1405) & (g1406) & (!g165) & (!g166)) + ((g1403) & (g1404) & (g1405) & (g1406) & (!g165) & (g166)) + ((g1403) & (g1404) & (g1405) & (g1406) & (g165) & (!g166)) + ((g1403) & (g1404) & (g1405) & (g1406) & (g165) & (g166)));
	assign g1408 = (((!g147) & (!g148) & (!g1393) & (g1397) & (!g1402) & (!g1407)) + ((!g147) & (!g148) & (!g1393) & (g1397) & (!g1402) & (g1407)) + ((!g147) & (!g148) & (!g1393) & (g1397) & (g1402) & (!g1407)) + ((!g147) & (!g148) & (!g1393) & (g1397) & (g1402) & (g1407)) + ((!g147) & (!g148) & (g1393) & (g1397) & (!g1402) & (!g1407)) + ((!g147) & (!g148) & (g1393) & (g1397) & (!g1402) & (g1407)) + ((!g147) & (!g148) & (g1393) & (g1397) & (g1402) & (!g1407)) + ((!g147) & (!g148) & (g1393) & (g1397) & (g1402) & (g1407)) + ((!g147) & (g148) & (!g1393) & (!g1397) & (!g1402) & (g1407)) + ((!g147) & (g148) & (!g1393) & (!g1397) & (g1402) & (g1407)) + ((!g147) & (g148) & (!g1393) & (g1397) & (!g1402) & (g1407)) + ((!g147) & (g148) & (!g1393) & (g1397) & (g1402) & (g1407)) + ((!g147) & (g148) & (g1393) & (!g1397) & (!g1402) & (g1407)) + ((!g147) & (g148) & (g1393) & (!g1397) & (g1402) & (g1407)) + ((!g147) & (g148) & (g1393) & (g1397) & (!g1402) & (g1407)) + ((!g147) & (g148) & (g1393) & (g1397) & (g1402) & (g1407)) + ((g147) & (!g148) & (g1393) & (!g1397) & (!g1402) & (!g1407)) + ((g147) & (!g148) & (g1393) & (!g1397) & (!g1402) & (g1407)) + ((g147) & (!g148) & (g1393) & (!g1397) & (g1402) & (!g1407)) + ((g147) & (!g148) & (g1393) & (!g1397) & (g1402) & (g1407)) + ((g147) & (!g148) & (g1393) & (g1397) & (!g1402) & (!g1407)) + ((g147) & (!g148) & (g1393) & (g1397) & (!g1402) & (g1407)) + ((g147) & (!g148) & (g1393) & (g1397) & (g1402) & (!g1407)) + ((g147) & (!g148) & (g1393) & (g1397) & (g1402) & (g1407)) + ((g147) & (g148) & (!g1393) & (!g1397) & (g1402) & (!g1407)) + ((g147) & (g148) & (!g1393) & (!g1397) & (g1402) & (g1407)) + ((g147) & (g148) & (!g1393) & (g1397) & (g1402) & (!g1407)) + ((g147) & (g148) & (!g1393) & (g1397) & (g1402) & (g1407)) + ((g147) & (g148) & (g1393) & (!g1397) & (g1402) & (!g1407)) + ((g147) & (g148) & (g1393) & (!g1397) & (g1402) & (g1407)) + ((g147) & (g148) & (g1393) & (g1397) & (g1402) & (!g1407)) + ((g147) & (g148) & (g1393) & (g1397) & (g1402) & (g1407)));
	assign g1409 = (((!g142) & (!g1388) & (!sk[67]) & (g1408)) + ((!g142) & (!g1388) & (sk[67]) & (g1408)) + ((!g142) & (g1388) & (!sk[67]) & (!g1408)) + ((!g142) & (g1388) & (!sk[67]) & (g1408)) + ((!g142) & (g1388) & (sk[67]) & (g1408)) + ((g142) & (!g1388) & (!sk[67]) & (g1408)) + ((g142) & (g1388) & (!sk[67]) & (!g1408)) + ((g142) & (g1388) & (!sk[67]) & (g1408)) + ((g142) & (g1388) & (sk[67]) & (!g1408)) + ((g142) & (g1388) & (sk[67]) & (g1408)));
	assign g4889 = (((!g2059) & (!sk[68]) & (!g2769) & (g1410)) + ((!g2059) & (!sk[68]) & (g2769) & (!g1410)) + ((!g2059) & (!sk[68]) & (g2769) & (g1410)) + ((!g2059) & (sk[68]) & (!g2769) & (g1410)) + ((!g2059) & (sk[68]) & (g2769) & (g1410)) + ((g2059) & (!sk[68]) & (!g2769) & (g1410)) + ((g2059) & (!sk[68]) & (g2769) & (!g1410)) + ((g2059) & (!sk[68]) & (g2769) & (g1410)) + ((g2059) & (sk[68]) & (g2769) & (!g1410)) + ((g2059) & (sk[68]) & (g2769) & (g1410)));
	assign g1411 = (((!sk[69]) & (!g1364) & (!g3823) & (!g1366) & (g916)) + ((!sk[69]) & (!g1364) & (!g3823) & (g1366) & (!g916)) + ((!sk[69]) & (!g1364) & (!g3823) & (g1366) & (g916)) + ((!sk[69]) & (!g1364) & (g3823) & (!g1366) & (!g916)) + ((!sk[69]) & (!g1364) & (g3823) & (!g1366) & (g916)) + ((!sk[69]) & (!g1364) & (g3823) & (g1366) & (!g916)) + ((!sk[69]) & (!g1364) & (g3823) & (g1366) & (g916)) + ((!sk[69]) & (g1364) & (!g3823) & (!g1366) & (g916)) + ((!sk[69]) & (g1364) & (!g3823) & (g1366) & (!g916)) + ((!sk[69]) & (g1364) & (!g3823) & (g1366) & (g916)) + ((!sk[69]) & (g1364) & (g3823) & (!g1366) & (!g916)) + ((!sk[69]) & (g1364) & (g3823) & (!g1366) & (g916)) + ((!sk[69]) & (g1364) & (g3823) & (g1366) & (!g916)) + ((!sk[69]) & (g1364) & (g3823) & (g1366) & (g916)) + ((sk[69]) & (!g1364) & (!g3823) & (!g1366) & (!g916)) + ((sk[69]) & (!g1364) & (!g3823) & (!g1366) & (g916)) + ((sk[69]) & (!g1364) & (!g3823) & (g1366) & (g916)) + ((sk[69]) & (!g1364) & (g3823) & (!g1366) & (g916)) + ((sk[69]) & (!g1364) & (g3823) & (g1366) & (g916)) + ((sk[69]) & (g1364) & (!g3823) & (!g1366) & (g916)));
	assign g1412 = (((!g126) & (!g1409) & (!g1410) & (!sk[70]) & (g1411) & (!g916)) + ((!g126) & (!g1409) & (!g1410) & (!sk[70]) & (g1411) & (g916)) + ((!g126) & (!g1409) & (g1410) & (!sk[70]) & (!g1411) & (!g916)) + ((!g126) & (!g1409) & (g1410) & (!sk[70]) & (!g1411) & (g916)) + ((!g126) & (!g1409) & (g1410) & (!sk[70]) & (g1411) & (!g916)) + ((!g126) & (!g1409) & (g1410) & (!sk[70]) & (g1411) & (g916)) + ((!g126) & (!g1409) & (g1410) & (sk[70]) & (!g1411) & (!g916)) + ((!g126) & (!g1409) & (g1410) & (sk[70]) & (!g1411) & (g916)) + ((!g126) & (!g1409) & (g1410) & (sk[70]) & (g1411) & (!g916)) + ((!g126) & (!g1409) & (g1410) & (sk[70]) & (g1411) & (g916)) + ((!g126) & (g1409) & (!g1410) & (!sk[70]) & (!g1411) & (!g916)) + ((!g126) & (g1409) & (!g1410) & (!sk[70]) & (!g1411) & (g916)) + ((!g126) & (g1409) & (!g1410) & (!sk[70]) & (g1411) & (!g916)) + ((!g126) & (g1409) & (!g1410) & (!sk[70]) & (g1411) & (g916)) + ((!g126) & (g1409) & (g1410) & (!sk[70]) & (!g1411) & (!g916)) + ((!g126) & (g1409) & (g1410) & (!sk[70]) & (!g1411) & (g916)) + ((!g126) & (g1409) & (g1410) & (!sk[70]) & (g1411) & (!g916)) + ((!g126) & (g1409) & (g1410) & (!sk[70]) & (g1411) & (g916)) + ((!g126) & (g1409) & (g1410) & (sk[70]) & (!g1411) & (!g916)) + ((!g126) & (g1409) & (g1410) & (sk[70]) & (!g1411) & (g916)) + ((!g126) & (g1409) & (g1410) & (sk[70]) & (g1411) & (!g916)) + ((!g126) & (g1409) & (g1410) & (sk[70]) & (g1411) & (g916)) + ((g126) & (!g1409) & (!g1410) & (!sk[70]) & (g1411) & (!g916)) + ((g126) & (!g1409) & (!g1410) & (!sk[70]) & (g1411) & (g916)) + ((g126) & (!g1409) & (!g1410) & (sk[70]) & (!g1411) & (g916)) + ((g126) & (!g1409) & (!g1410) & (sk[70]) & (g1411) & (!g916)) + ((g126) & (!g1409) & (g1410) & (!sk[70]) & (!g1411) & (!g916)) + ((g126) & (!g1409) & (g1410) & (!sk[70]) & (!g1411) & (g916)) + ((g126) & (!g1409) & (g1410) & (!sk[70]) & (g1411) & (!g916)) + ((g126) & (!g1409) & (g1410) & (!sk[70]) & (g1411) & (g916)) + ((g126) & (!g1409) & (g1410) & (sk[70]) & (!g1411) & (g916)) + ((g126) & (!g1409) & (g1410) & (sk[70]) & (g1411) & (!g916)) + ((g126) & (g1409) & (!g1410) & (!sk[70]) & (!g1411) & (!g916)) + ((g126) & (g1409) & (!g1410) & (!sk[70]) & (!g1411) & (g916)) + ((g126) & (g1409) & (!g1410) & (!sk[70]) & (g1411) & (!g916)) + ((g126) & (g1409) & (!g1410) & (!sk[70]) & (g1411) & (g916)) + ((g126) & (g1409) & (!g1410) & (sk[70]) & (!g1411) & (!g916)) + ((g126) & (g1409) & (!g1410) & (sk[70]) & (g1411) & (g916)) + ((g126) & (g1409) & (g1410) & (!sk[70]) & (!g1411) & (!g916)) + ((g126) & (g1409) & (g1410) & (!sk[70]) & (!g1411) & (g916)) + ((g126) & (g1409) & (g1410) & (!sk[70]) & (g1411) & (!g916)) + ((g126) & (g1409) & (g1410) & (!sk[70]) & (g1411) & (g916)) + ((g126) & (g1409) & (g1410) & (sk[70]) & (!g1411) & (!g916)) + ((g126) & (g1409) & (g1410) & (sk[70]) & (g1411) & (g916)));
	assign g4890 = (((!g2140) & (!sk[71]) & (!g2787) & (g1413)) + ((!g2140) & (!sk[71]) & (g2787) & (!g1413)) + ((!g2140) & (!sk[71]) & (g2787) & (g1413)) + ((!g2140) & (sk[71]) & (!g2787) & (g1413)) + ((!g2140) & (sk[71]) & (g2787) & (g1413)) + ((g2140) & (!sk[71]) & (!g2787) & (g1413)) + ((g2140) & (!sk[71]) & (g2787) & (!g1413)) + ((g2140) & (!sk[71]) & (g2787) & (g1413)) + ((g2140) & (sk[71]) & (g2787) & (!g1413)) + ((g2140) & (sk[71]) & (g2787) & (g1413)));
	assign g4891 = (((!sk[72]) & (!g2142) & (!g2787) & (g1414)) + ((!sk[72]) & (!g2142) & (g2787) & (!g1414)) + ((!sk[72]) & (!g2142) & (g2787) & (g1414)) + ((!sk[72]) & (g2142) & (!g2787) & (g1414)) + ((!sk[72]) & (g2142) & (g2787) & (!g1414)) + ((!sk[72]) & (g2142) & (g2787) & (g1414)) + ((sk[72]) & (!g2142) & (!g2787) & (g1414)) + ((sk[72]) & (!g2142) & (g2787) & (g1414)) + ((sk[72]) & (g2142) & (g2787) & (!g1414)) + ((sk[72]) & (g2142) & (g2787) & (g1414)));
	assign g4892 = (((!g2144) & (!g2787) & (!sk[73]) & (g1415)) + ((!g2144) & (!g2787) & (sk[73]) & (g1415)) + ((!g2144) & (g2787) & (!sk[73]) & (!g1415)) + ((!g2144) & (g2787) & (!sk[73]) & (g1415)) + ((!g2144) & (g2787) & (sk[73]) & (g1415)) + ((g2144) & (!g2787) & (!sk[73]) & (g1415)) + ((g2144) & (g2787) & (!sk[73]) & (!g1415)) + ((g2144) & (g2787) & (!sk[73]) & (g1415)) + ((g2144) & (g2787) & (sk[73]) & (!g1415)) + ((g2144) & (g2787) & (sk[73]) & (g1415)));
	assign g4893 = (((!sk[74]) & (!g2145) & (!g2787) & (g1416)) + ((!sk[74]) & (!g2145) & (g2787) & (!g1416)) + ((!sk[74]) & (!g2145) & (g2787) & (g1416)) + ((!sk[74]) & (g2145) & (!g2787) & (g1416)) + ((!sk[74]) & (g2145) & (g2787) & (!g1416)) + ((!sk[74]) & (g2145) & (g2787) & (g1416)) + ((sk[74]) & (!g2145) & (!g2787) & (g1416)) + ((sk[74]) & (!g2145) & (g2787) & (g1416)) + ((sk[74]) & (g2145) & (g2787) & (!g1416)) + ((sk[74]) & (g2145) & (g2787) & (g1416)));
	assign g1417 = (((!g1413) & (!g1414) & (!g1415) & (g1416) & (g147) & (g148)) + ((!g1413) & (!g1414) & (g1415) & (!g1416) & (!g147) & (g148)) + ((!g1413) & (!g1414) & (g1415) & (g1416) & (!g147) & (g148)) + ((!g1413) & (!g1414) & (g1415) & (g1416) & (g147) & (g148)) + ((!g1413) & (g1414) & (!g1415) & (!g1416) & (g147) & (!g148)) + ((!g1413) & (g1414) & (!g1415) & (g1416) & (g147) & (!g148)) + ((!g1413) & (g1414) & (!g1415) & (g1416) & (g147) & (g148)) + ((!g1413) & (g1414) & (g1415) & (!g1416) & (!g147) & (g148)) + ((!g1413) & (g1414) & (g1415) & (!g1416) & (g147) & (!g148)) + ((!g1413) & (g1414) & (g1415) & (g1416) & (!g147) & (g148)) + ((!g1413) & (g1414) & (g1415) & (g1416) & (g147) & (!g148)) + ((!g1413) & (g1414) & (g1415) & (g1416) & (g147) & (g148)) + ((g1413) & (!g1414) & (!g1415) & (!g1416) & (!g147) & (!g148)) + ((g1413) & (!g1414) & (!g1415) & (g1416) & (!g147) & (!g148)) + ((g1413) & (!g1414) & (!g1415) & (g1416) & (g147) & (g148)) + ((g1413) & (!g1414) & (g1415) & (!g1416) & (!g147) & (!g148)) + ((g1413) & (!g1414) & (g1415) & (!g1416) & (!g147) & (g148)) + ((g1413) & (!g1414) & (g1415) & (g1416) & (!g147) & (!g148)) + ((g1413) & (!g1414) & (g1415) & (g1416) & (!g147) & (g148)) + ((g1413) & (!g1414) & (g1415) & (g1416) & (g147) & (g148)) + ((g1413) & (g1414) & (!g1415) & (!g1416) & (!g147) & (!g148)) + ((g1413) & (g1414) & (!g1415) & (!g1416) & (g147) & (!g148)) + ((g1413) & (g1414) & (!g1415) & (g1416) & (!g147) & (!g148)) + ((g1413) & (g1414) & (!g1415) & (g1416) & (g147) & (!g148)) + ((g1413) & (g1414) & (!g1415) & (g1416) & (g147) & (g148)) + ((g1413) & (g1414) & (g1415) & (!g1416) & (!g147) & (!g148)) + ((g1413) & (g1414) & (g1415) & (!g1416) & (!g147) & (g148)) + ((g1413) & (g1414) & (g1415) & (!g1416) & (g147) & (!g148)) + ((g1413) & (g1414) & (g1415) & (g1416) & (!g147) & (!g148)) + ((g1413) & (g1414) & (g1415) & (g1416) & (!g147) & (g148)) + ((g1413) & (g1414) & (g1415) & (g1416) & (g147) & (!g148)) + ((g1413) & (g1414) & (g1415) & (g1416) & (g147) & (g148)));
	assign g4894 = (((!sk[76]) & (!g2146) & (!g2787) & (g1418)) + ((!sk[76]) & (!g2146) & (g2787) & (!g1418)) + ((!sk[76]) & (!g2146) & (g2787) & (g1418)) + ((!sk[76]) & (g2146) & (!g2787) & (g1418)) + ((!sk[76]) & (g2146) & (g2787) & (!g1418)) + ((!sk[76]) & (g2146) & (g2787) & (g1418)) + ((sk[76]) & (!g2146) & (!g2787) & (g1418)) + ((sk[76]) & (!g2146) & (g2787) & (g1418)) + ((sk[76]) & (g2146) & (g2787) & (!g1418)) + ((sk[76]) & (g2146) & (g2787) & (g1418)));
	assign g4895 = (((!g2148) & (!sk[77]) & (!g2787) & (g1419)) + ((!g2148) & (!sk[77]) & (g2787) & (!g1419)) + ((!g2148) & (!sk[77]) & (g2787) & (g1419)) + ((!g2148) & (sk[77]) & (!g2787) & (g1419)) + ((!g2148) & (sk[77]) & (g2787) & (g1419)) + ((g2148) & (!sk[77]) & (!g2787) & (g1419)) + ((g2148) & (!sk[77]) & (g2787) & (!g1419)) + ((g2148) & (!sk[77]) & (g2787) & (g1419)) + ((g2148) & (sk[77]) & (g2787) & (!g1419)) + ((g2148) & (sk[77]) & (g2787) & (g1419)));
	assign g4896 = (((!sk[78]) & (!g2150) & (!g2787) & (g1420)) + ((!sk[78]) & (!g2150) & (g2787) & (!g1420)) + ((!sk[78]) & (!g2150) & (g2787) & (g1420)) + ((!sk[78]) & (g2150) & (!g2787) & (g1420)) + ((!sk[78]) & (g2150) & (g2787) & (!g1420)) + ((!sk[78]) & (g2150) & (g2787) & (g1420)) + ((sk[78]) & (!g2150) & (!g2787) & (g1420)) + ((sk[78]) & (!g2150) & (g2787) & (g1420)) + ((sk[78]) & (g2150) & (g2787) & (!g1420)) + ((sk[78]) & (g2150) & (g2787) & (g1420)));
	assign g4897 = (((!sk[79]) & (!g2151) & (!g2787) & (g1421)) + ((!sk[79]) & (!g2151) & (g2787) & (!g1421)) + ((!sk[79]) & (!g2151) & (g2787) & (g1421)) + ((!sk[79]) & (g2151) & (!g2787) & (g1421)) + ((!sk[79]) & (g2151) & (g2787) & (!g1421)) + ((!sk[79]) & (g2151) & (g2787) & (g1421)) + ((sk[79]) & (!g2151) & (!g2787) & (g1421)) + ((sk[79]) & (!g2151) & (g2787) & (g1421)) + ((sk[79]) & (g2151) & (g2787) & (!g1421)) + ((sk[79]) & (g2151) & (g2787) & (g1421)));
	assign g1422 = (((!g1418) & (!g1419) & (!g1420) & (g1421) & (g147) & (g148)) + ((!g1418) & (!g1419) & (g1420) & (!g1421) & (!g147) & (g148)) + ((!g1418) & (!g1419) & (g1420) & (g1421) & (!g147) & (g148)) + ((!g1418) & (!g1419) & (g1420) & (g1421) & (g147) & (g148)) + ((!g1418) & (g1419) & (!g1420) & (!g1421) & (g147) & (!g148)) + ((!g1418) & (g1419) & (!g1420) & (g1421) & (g147) & (!g148)) + ((!g1418) & (g1419) & (!g1420) & (g1421) & (g147) & (g148)) + ((!g1418) & (g1419) & (g1420) & (!g1421) & (!g147) & (g148)) + ((!g1418) & (g1419) & (g1420) & (!g1421) & (g147) & (!g148)) + ((!g1418) & (g1419) & (g1420) & (g1421) & (!g147) & (g148)) + ((!g1418) & (g1419) & (g1420) & (g1421) & (g147) & (!g148)) + ((!g1418) & (g1419) & (g1420) & (g1421) & (g147) & (g148)) + ((g1418) & (!g1419) & (!g1420) & (!g1421) & (!g147) & (!g148)) + ((g1418) & (!g1419) & (!g1420) & (g1421) & (!g147) & (!g148)) + ((g1418) & (!g1419) & (!g1420) & (g1421) & (g147) & (g148)) + ((g1418) & (!g1419) & (g1420) & (!g1421) & (!g147) & (!g148)) + ((g1418) & (!g1419) & (g1420) & (!g1421) & (!g147) & (g148)) + ((g1418) & (!g1419) & (g1420) & (g1421) & (!g147) & (!g148)) + ((g1418) & (!g1419) & (g1420) & (g1421) & (!g147) & (g148)) + ((g1418) & (!g1419) & (g1420) & (g1421) & (g147) & (g148)) + ((g1418) & (g1419) & (!g1420) & (!g1421) & (!g147) & (!g148)) + ((g1418) & (g1419) & (!g1420) & (!g1421) & (g147) & (!g148)) + ((g1418) & (g1419) & (!g1420) & (g1421) & (!g147) & (!g148)) + ((g1418) & (g1419) & (!g1420) & (g1421) & (g147) & (!g148)) + ((g1418) & (g1419) & (!g1420) & (g1421) & (g147) & (g148)) + ((g1418) & (g1419) & (g1420) & (!g1421) & (!g147) & (!g148)) + ((g1418) & (g1419) & (g1420) & (!g1421) & (!g147) & (g148)) + ((g1418) & (g1419) & (g1420) & (!g1421) & (g147) & (!g148)) + ((g1418) & (g1419) & (g1420) & (g1421) & (!g147) & (!g148)) + ((g1418) & (g1419) & (g1420) & (g1421) & (!g147) & (g148)) + ((g1418) & (g1419) & (g1420) & (g1421) & (g147) & (!g148)) + ((g1418) & (g1419) & (g1420) & (g1421) & (g147) & (g148)));
	assign g4898 = (((!g2152) & (!sk[81]) & (!g2787) & (g1423)) + ((!g2152) & (!sk[81]) & (g2787) & (!g1423)) + ((!g2152) & (!sk[81]) & (g2787) & (g1423)) + ((!g2152) & (sk[81]) & (!g2787) & (g1423)) + ((!g2152) & (sk[81]) & (g2787) & (g1423)) + ((g2152) & (!sk[81]) & (!g2787) & (g1423)) + ((g2152) & (!sk[81]) & (g2787) & (!g1423)) + ((g2152) & (!sk[81]) & (g2787) & (g1423)) + ((g2152) & (sk[81]) & (g2787) & (!g1423)) + ((g2152) & (sk[81]) & (g2787) & (g1423)));
	assign g4899 = (((!g2153) & (!g2787) & (!sk[82]) & (g1424)) + ((!g2153) & (!g2787) & (sk[82]) & (g1424)) + ((!g2153) & (g2787) & (!sk[82]) & (!g1424)) + ((!g2153) & (g2787) & (!sk[82]) & (g1424)) + ((!g2153) & (g2787) & (sk[82]) & (g1424)) + ((g2153) & (!g2787) & (!sk[82]) & (g1424)) + ((g2153) & (g2787) & (!sk[82]) & (!g1424)) + ((g2153) & (g2787) & (!sk[82]) & (g1424)) + ((g2153) & (g2787) & (sk[82]) & (!g1424)) + ((g2153) & (g2787) & (sk[82]) & (g1424)));
	assign g4900 = (((!g2155) & (!sk[83]) & (!g2787) & (g1425)) + ((!g2155) & (!sk[83]) & (g2787) & (!g1425)) + ((!g2155) & (!sk[83]) & (g2787) & (g1425)) + ((!g2155) & (sk[83]) & (!g2787) & (g1425)) + ((!g2155) & (sk[83]) & (g2787) & (g1425)) + ((g2155) & (!sk[83]) & (!g2787) & (g1425)) + ((g2155) & (!sk[83]) & (g2787) & (!g1425)) + ((g2155) & (!sk[83]) & (g2787) & (g1425)) + ((g2155) & (sk[83]) & (g2787) & (!g1425)) + ((g2155) & (sk[83]) & (g2787) & (g1425)));
	assign g4901 = (((!g2157) & (!sk[84]) & (!g2787) & (g1426)) + ((!g2157) & (!sk[84]) & (g2787) & (!g1426)) + ((!g2157) & (!sk[84]) & (g2787) & (g1426)) + ((!g2157) & (sk[84]) & (!g2787) & (g1426)) + ((!g2157) & (sk[84]) & (g2787) & (g1426)) + ((g2157) & (!sk[84]) & (!g2787) & (g1426)) + ((g2157) & (!sk[84]) & (g2787) & (!g1426)) + ((g2157) & (!sk[84]) & (g2787) & (g1426)) + ((g2157) & (sk[84]) & (g2787) & (!g1426)) + ((g2157) & (sk[84]) & (g2787) & (g1426)));
	assign g1427 = (((!g1423) & (!g1424) & (!g1425) & (g1426) & (g147) & (g148)) + ((!g1423) & (!g1424) & (g1425) & (!g1426) & (!g147) & (g148)) + ((!g1423) & (!g1424) & (g1425) & (g1426) & (!g147) & (g148)) + ((!g1423) & (!g1424) & (g1425) & (g1426) & (g147) & (g148)) + ((!g1423) & (g1424) & (!g1425) & (!g1426) & (g147) & (!g148)) + ((!g1423) & (g1424) & (!g1425) & (g1426) & (g147) & (!g148)) + ((!g1423) & (g1424) & (!g1425) & (g1426) & (g147) & (g148)) + ((!g1423) & (g1424) & (g1425) & (!g1426) & (!g147) & (g148)) + ((!g1423) & (g1424) & (g1425) & (!g1426) & (g147) & (!g148)) + ((!g1423) & (g1424) & (g1425) & (g1426) & (!g147) & (g148)) + ((!g1423) & (g1424) & (g1425) & (g1426) & (g147) & (!g148)) + ((!g1423) & (g1424) & (g1425) & (g1426) & (g147) & (g148)) + ((g1423) & (!g1424) & (!g1425) & (!g1426) & (!g147) & (!g148)) + ((g1423) & (!g1424) & (!g1425) & (g1426) & (!g147) & (!g148)) + ((g1423) & (!g1424) & (!g1425) & (g1426) & (g147) & (g148)) + ((g1423) & (!g1424) & (g1425) & (!g1426) & (!g147) & (!g148)) + ((g1423) & (!g1424) & (g1425) & (!g1426) & (!g147) & (g148)) + ((g1423) & (!g1424) & (g1425) & (g1426) & (!g147) & (!g148)) + ((g1423) & (!g1424) & (g1425) & (g1426) & (!g147) & (g148)) + ((g1423) & (!g1424) & (g1425) & (g1426) & (g147) & (g148)) + ((g1423) & (g1424) & (!g1425) & (!g1426) & (!g147) & (!g148)) + ((g1423) & (g1424) & (!g1425) & (!g1426) & (g147) & (!g148)) + ((g1423) & (g1424) & (!g1425) & (g1426) & (!g147) & (!g148)) + ((g1423) & (g1424) & (!g1425) & (g1426) & (g147) & (!g148)) + ((g1423) & (g1424) & (!g1425) & (g1426) & (g147) & (g148)) + ((g1423) & (g1424) & (g1425) & (!g1426) & (!g147) & (!g148)) + ((g1423) & (g1424) & (g1425) & (!g1426) & (!g147) & (g148)) + ((g1423) & (g1424) & (g1425) & (!g1426) & (g147) & (!g148)) + ((g1423) & (g1424) & (g1425) & (g1426) & (!g147) & (!g148)) + ((g1423) & (g1424) & (g1425) & (g1426) & (!g147) & (g148)) + ((g1423) & (g1424) & (g1425) & (g1426) & (g147) & (!g148)) + ((g1423) & (g1424) & (g1425) & (g1426) & (g147) & (g148)));
	assign g4902 = (((!sk[86]) & (!g2158) & (!g2787) & (g1428)) + ((!sk[86]) & (!g2158) & (g2787) & (!g1428)) + ((!sk[86]) & (!g2158) & (g2787) & (g1428)) + ((!sk[86]) & (g2158) & (!g2787) & (g1428)) + ((!sk[86]) & (g2158) & (g2787) & (!g1428)) + ((!sk[86]) & (g2158) & (g2787) & (g1428)) + ((sk[86]) & (!g2158) & (!g2787) & (g1428)) + ((sk[86]) & (!g2158) & (g2787) & (g1428)) + ((sk[86]) & (g2158) & (g2787) & (!g1428)) + ((sk[86]) & (g2158) & (g2787) & (g1428)));
	assign g4903 = (((!g2159) & (!sk[87]) & (!g2787) & (g1429)) + ((!g2159) & (!sk[87]) & (g2787) & (!g1429)) + ((!g2159) & (!sk[87]) & (g2787) & (g1429)) + ((!g2159) & (sk[87]) & (!g2787) & (g1429)) + ((!g2159) & (sk[87]) & (g2787) & (g1429)) + ((g2159) & (!sk[87]) & (!g2787) & (g1429)) + ((g2159) & (!sk[87]) & (g2787) & (!g1429)) + ((g2159) & (!sk[87]) & (g2787) & (g1429)) + ((g2159) & (sk[87]) & (g2787) & (!g1429)) + ((g2159) & (sk[87]) & (g2787) & (g1429)));
	assign g4904 = (((!g2160) & (!sk[88]) & (!g2787) & (g1430)) + ((!g2160) & (!sk[88]) & (g2787) & (!g1430)) + ((!g2160) & (!sk[88]) & (g2787) & (g1430)) + ((!g2160) & (sk[88]) & (!g2787) & (g1430)) + ((!g2160) & (sk[88]) & (g2787) & (g1430)) + ((g2160) & (!sk[88]) & (!g2787) & (g1430)) + ((g2160) & (!sk[88]) & (g2787) & (!g1430)) + ((g2160) & (!sk[88]) & (g2787) & (g1430)) + ((g2160) & (sk[88]) & (g2787) & (!g1430)) + ((g2160) & (sk[88]) & (g2787) & (g1430)));
	assign g4905 = (((!g2161) & (!g2787) & (!sk[89]) & (g1431)) + ((!g2161) & (!g2787) & (sk[89]) & (g1431)) + ((!g2161) & (g2787) & (!sk[89]) & (!g1431)) + ((!g2161) & (g2787) & (!sk[89]) & (g1431)) + ((!g2161) & (g2787) & (sk[89]) & (g1431)) + ((g2161) & (!g2787) & (!sk[89]) & (g1431)) + ((g2161) & (g2787) & (!sk[89]) & (!g1431)) + ((g2161) & (g2787) & (!sk[89]) & (g1431)) + ((g2161) & (g2787) & (sk[89]) & (!g1431)) + ((g2161) & (g2787) & (sk[89]) & (g1431)));
	assign g1432 = (((!g1428) & (!g1429) & (!g1430) & (g1431) & (g147) & (g148)) + ((!g1428) & (!g1429) & (g1430) & (!g1431) & (!g147) & (g148)) + ((!g1428) & (!g1429) & (g1430) & (g1431) & (!g147) & (g148)) + ((!g1428) & (!g1429) & (g1430) & (g1431) & (g147) & (g148)) + ((!g1428) & (g1429) & (!g1430) & (!g1431) & (g147) & (!g148)) + ((!g1428) & (g1429) & (!g1430) & (g1431) & (g147) & (!g148)) + ((!g1428) & (g1429) & (!g1430) & (g1431) & (g147) & (g148)) + ((!g1428) & (g1429) & (g1430) & (!g1431) & (!g147) & (g148)) + ((!g1428) & (g1429) & (g1430) & (!g1431) & (g147) & (!g148)) + ((!g1428) & (g1429) & (g1430) & (g1431) & (!g147) & (g148)) + ((!g1428) & (g1429) & (g1430) & (g1431) & (g147) & (!g148)) + ((!g1428) & (g1429) & (g1430) & (g1431) & (g147) & (g148)) + ((g1428) & (!g1429) & (!g1430) & (!g1431) & (!g147) & (!g148)) + ((g1428) & (!g1429) & (!g1430) & (g1431) & (!g147) & (!g148)) + ((g1428) & (!g1429) & (!g1430) & (g1431) & (g147) & (g148)) + ((g1428) & (!g1429) & (g1430) & (!g1431) & (!g147) & (!g148)) + ((g1428) & (!g1429) & (g1430) & (!g1431) & (!g147) & (g148)) + ((g1428) & (!g1429) & (g1430) & (g1431) & (!g147) & (!g148)) + ((g1428) & (!g1429) & (g1430) & (g1431) & (!g147) & (g148)) + ((g1428) & (!g1429) & (g1430) & (g1431) & (g147) & (g148)) + ((g1428) & (g1429) & (!g1430) & (!g1431) & (!g147) & (!g148)) + ((g1428) & (g1429) & (!g1430) & (!g1431) & (g147) & (!g148)) + ((g1428) & (g1429) & (!g1430) & (g1431) & (!g147) & (!g148)) + ((g1428) & (g1429) & (!g1430) & (g1431) & (g147) & (!g148)) + ((g1428) & (g1429) & (!g1430) & (g1431) & (g147) & (g148)) + ((g1428) & (g1429) & (g1430) & (!g1431) & (!g147) & (!g148)) + ((g1428) & (g1429) & (g1430) & (!g1431) & (!g147) & (g148)) + ((g1428) & (g1429) & (g1430) & (!g1431) & (g147) & (!g148)) + ((g1428) & (g1429) & (g1430) & (g1431) & (!g147) & (!g148)) + ((g1428) & (g1429) & (g1430) & (g1431) & (!g147) & (g148)) + ((g1428) & (g1429) & (g1430) & (g1431) & (g147) & (!g148)) + ((g1428) & (g1429) & (g1430) & (g1431) & (g147) & (g148)));
	assign g1433 = (((!g1417) & (!g1422) & (!g1427) & (g1432) & (g165) & (g166)) + ((!g1417) & (!g1422) & (g1427) & (!g1432) & (!g165) & (g166)) + ((!g1417) & (!g1422) & (g1427) & (g1432) & (!g165) & (g166)) + ((!g1417) & (!g1422) & (g1427) & (g1432) & (g165) & (g166)) + ((!g1417) & (g1422) & (!g1427) & (!g1432) & (g165) & (!g166)) + ((!g1417) & (g1422) & (!g1427) & (g1432) & (g165) & (!g166)) + ((!g1417) & (g1422) & (!g1427) & (g1432) & (g165) & (g166)) + ((!g1417) & (g1422) & (g1427) & (!g1432) & (!g165) & (g166)) + ((!g1417) & (g1422) & (g1427) & (!g1432) & (g165) & (!g166)) + ((!g1417) & (g1422) & (g1427) & (g1432) & (!g165) & (g166)) + ((!g1417) & (g1422) & (g1427) & (g1432) & (g165) & (!g166)) + ((!g1417) & (g1422) & (g1427) & (g1432) & (g165) & (g166)) + ((g1417) & (!g1422) & (!g1427) & (!g1432) & (!g165) & (!g166)) + ((g1417) & (!g1422) & (!g1427) & (g1432) & (!g165) & (!g166)) + ((g1417) & (!g1422) & (!g1427) & (g1432) & (g165) & (g166)) + ((g1417) & (!g1422) & (g1427) & (!g1432) & (!g165) & (!g166)) + ((g1417) & (!g1422) & (g1427) & (!g1432) & (!g165) & (g166)) + ((g1417) & (!g1422) & (g1427) & (g1432) & (!g165) & (!g166)) + ((g1417) & (!g1422) & (g1427) & (g1432) & (!g165) & (g166)) + ((g1417) & (!g1422) & (g1427) & (g1432) & (g165) & (g166)) + ((g1417) & (g1422) & (!g1427) & (!g1432) & (!g165) & (!g166)) + ((g1417) & (g1422) & (!g1427) & (!g1432) & (g165) & (!g166)) + ((g1417) & (g1422) & (!g1427) & (g1432) & (!g165) & (!g166)) + ((g1417) & (g1422) & (!g1427) & (g1432) & (g165) & (!g166)) + ((g1417) & (g1422) & (!g1427) & (g1432) & (g165) & (g166)) + ((g1417) & (g1422) & (g1427) & (!g1432) & (!g165) & (!g166)) + ((g1417) & (g1422) & (g1427) & (!g1432) & (!g165) & (g166)) + ((g1417) & (g1422) & (g1427) & (!g1432) & (g165) & (!g166)) + ((g1417) & (g1422) & (g1427) & (g1432) & (!g165) & (!g166)) + ((g1417) & (g1422) & (g1427) & (g1432) & (!g165) & (g166)) + ((g1417) & (g1422) & (g1427) & (g1432) & (g165) & (!g166)) + ((g1417) & (g1422) & (g1427) & (g1432) & (g165) & (g166)));
	assign g4906 = (((!g2173) & (!sk[92]) & (!g2787) & (g1434)) + ((!g2173) & (!sk[92]) & (g2787) & (!g1434)) + ((!g2173) & (!sk[92]) & (g2787) & (g1434)) + ((!g2173) & (sk[92]) & (!g2787) & (g1434)) + ((!g2173) & (sk[92]) & (g2787) & (g1434)) + ((g2173) & (!sk[92]) & (!g2787) & (g1434)) + ((g2173) & (!sk[92]) & (g2787) & (!g1434)) + ((g2173) & (!sk[92]) & (g2787) & (g1434)) + ((g2173) & (sk[92]) & (g2787) & (!g1434)) + ((g2173) & (sk[92]) & (g2787) & (g1434)));
	assign g4907 = (((!g2174) & (!sk[93]) & (!g2787) & (g1435)) + ((!g2174) & (!sk[93]) & (g2787) & (!g1435)) + ((!g2174) & (!sk[93]) & (g2787) & (g1435)) + ((!g2174) & (sk[93]) & (!g2787) & (g1435)) + ((!g2174) & (sk[93]) & (g2787) & (g1435)) + ((g2174) & (!sk[93]) & (!g2787) & (g1435)) + ((g2174) & (!sk[93]) & (g2787) & (!g1435)) + ((g2174) & (!sk[93]) & (g2787) & (g1435)) + ((g2174) & (sk[93]) & (g2787) & (!g1435)) + ((g2174) & (sk[93]) & (g2787) & (g1435)));
	assign g4908 = (((!g2175) & (!sk[94]) & (!g2787) & (g1436)) + ((!g2175) & (!sk[94]) & (g2787) & (!g1436)) + ((!g2175) & (!sk[94]) & (g2787) & (g1436)) + ((!g2175) & (sk[94]) & (!g2787) & (g1436)) + ((!g2175) & (sk[94]) & (g2787) & (g1436)) + ((g2175) & (!sk[94]) & (!g2787) & (g1436)) + ((g2175) & (!sk[94]) & (g2787) & (!g1436)) + ((g2175) & (!sk[94]) & (g2787) & (g1436)) + ((g2175) & (sk[94]) & (g2787) & (!g1436)) + ((g2175) & (sk[94]) & (g2787) & (g1436)));
	assign g4909 = (((!sk[95]) & (!g2176) & (!g2787) & (g1437)) + ((!sk[95]) & (!g2176) & (g2787) & (!g1437)) + ((!sk[95]) & (!g2176) & (g2787) & (g1437)) + ((!sk[95]) & (g2176) & (!g2787) & (g1437)) + ((!sk[95]) & (g2176) & (g2787) & (!g1437)) + ((!sk[95]) & (g2176) & (g2787) & (g1437)) + ((sk[95]) & (!g2176) & (!g2787) & (g1437)) + ((sk[95]) & (!g2176) & (g2787) & (g1437)) + ((sk[95]) & (g2176) & (g2787) & (!g1437)) + ((sk[95]) & (g2176) & (g2787) & (g1437)));
	assign g1438 = (((!g1434) & (!g1435) & (!g1436) & (g1437) & (g165) & (g166)) + ((!g1434) & (!g1435) & (g1436) & (!g1437) & (!g165) & (g166)) + ((!g1434) & (!g1435) & (g1436) & (g1437) & (!g165) & (g166)) + ((!g1434) & (!g1435) & (g1436) & (g1437) & (g165) & (g166)) + ((!g1434) & (g1435) & (!g1436) & (!g1437) & (g165) & (!g166)) + ((!g1434) & (g1435) & (!g1436) & (g1437) & (g165) & (!g166)) + ((!g1434) & (g1435) & (!g1436) & (g1437) & (g165) & (g166)) + ((!g1434) & (g1435) & (g1436) & (!g1437) & (!g165) & (g166)) + ((!g1434) & (g1435) & (g1436) & (!g1437) & (g165) & (!g166)) + ((!g1434) & (g1435) & (g1436) & (g1437) & (!g165) & (g166)) + ((!g1434) & (g1435) & (g1436) & (g1437) & (g165) & (!g166)) + ((!g1434) & (g1435) & (g1436) & (g1437) & (g165) & (g166)) + ((g1434) & (!g1435) & (!g1436) & (!g1437) & (!g165) & (!g166)) + ((g1434) & (!g1435) & (!g1436) & (g1437) & (!g165) & (!g166)) + ((g1434) & (!g1435) & (!g1436) & (g1437) & (g165) & (g166)) + ((g1434) & (!g1435) & (g1436) & (!g1437) & (!g165) & (!g166)) + ((g1434) & (!g1435) & (g1436) & (!g1437) & (!g165) & (g166)) + ((g1434) & (!g1435) & (g1436) & (g1437) & (!g165) & (!g166)) + ((g1434) & (!g1435) & (g1436) & (g1437) & (!g165) & (g166)) + ((g1434) & (!g1435) & (g1436) & (g1437) & (g165) & (g166)) + ((g1434) & (g1435) & (!g1436) & (!g1437) & (!g165) & (!g166)) + ((g1434) & (g1435) & (!g1436) & (!g1437) & (g165) & (!g166)) + ((g1434) & (g1435) & (!g1436) & (g1437) & (!g165) & (!g166)) + ((g1434) & (g1435) & (!g1436) & (g1437) & (g165) & (!g166)) + ((g1434) & (g1435) & (!g1436) & (g1437) & (g165) & (g166)) + ((g1434) & (g1435) & (g1436) & (!g1437) & (!g165) & (!g166)) + ((g1434) & (g1435) & (g1436) & (!g1437) & (!g165) & (g166)) + ((g1434) & (g1435) & (g1436) & (!g1437) & (g165) & (!g166)) + ((g1434) & (g1435) & (g1436) & (g1437) & (!g165) & (!g166)) + ((g1434) & (g1435) & (g1436) & (g1437) & (!g165) & (g166)) + ((g1434) & (g1435) & (g1436) & (g1437) & (g165) & (!g166)) + ((g1434) & (g1435) & (g1436) & (g1437) & (g165) & (g166)));
	assign g4910 = (((!g2177) & (!g2787) & (!sk[97]) & (g1439)) + ((!g2177) & (!g2787) & (sk[97]) & (g1439)) + ((!g2177) & (g2787) & (!sk[97]) & (!g1439)) + ((!g2177) & (g2787) & (!sk[97]) & (g1439)) + ((!g2177) & (g2787) & (sk[97]) & (g1439)) + ((g2177) & (!g2787) & (!sk[97]) & (g1439)) + ((g2177) & (g2787) & (!sk[97]) & (!g1439)) + ((g2177) & (g2787) & (!sk[97]) & (g1439)) + ((g2177) & (g2787) & (sk[97]) & (!g1439)) + ((g2177) & (g2787) & (sk[97]) & (g1439)));
	assign g4911 = (((!g2178) & (!sk[98]) & (!g2787) & (g1440)) + ((!g2178) & (!sk[98]) & (g2787) & (!g1440)) + ((!g2178) & (!sk[98]) & (g2787) & (g1440)) + ((!g2178) & (sk[98]) & (!g2787) & (g1440)) + ((!g2178) & (sk[98]) & (g2787) & (g1440)) + ((g2178) & (!sk[98]) & (!g2787) & (g1440)) + ((g2178) & (!sk[98]) & (g2787) & (!g1440)) + ((g2178) & (!sk[98]) & (g2787) & (g1440)) + ((g2178) & (sk[98]) & (g2787) & (!g1440)) + ((g2178) & (sk[98]) & (g2787) & (g1440)));
	assign g4912 = (((!g2179) & (!sk[99]) & (!g2787) & (g1441)) + ((!g2179) & (!sk[99]) & (g2787) & (!g1441)) + ((!g2179) & (!sk[99]) & (g2787) & (g1441)) + ((!g2179) & (sk[99]) & (!g2787) & (g1441)) + ((!g2179) & (sk[99]) & (g2787) & (g1441)) + ((g2179) & (!sk[99]) & (!g2787) & (g1441)) + ((g2179) & (!sk[99]) & (g2787) & (!g1441)) + ((g2179) & (!sk[99]) & (g2787) & (g1441)) + ((g2179) & (sk[99]) & (g2787) & (!g1441)) + ((g2179) & (sk[99]) & (g2787) & (g1441)));
	assign g1442 = (((!g165) & (!g166) & (!g1439) & (g1440) & (!sk[100]) & (!g1441)) + ((!g165) & (!g166) & (!g1439) & (g1440) & (!sk[100]) & (g1441)) + ((!g165) & (!g166) & (g1439) & (!g1440) & (!sk[100]) & (!g1441)) + ((!g165) & (!g166) & (g1439) & (!g1440) & (!sk[100]) & (g1441)) + ((!g165) & (!g166) & (g1439) & (g1440) & (!sk[100]) & (!g1441)) + ((!g165) & (!g166) & (g1439) & (g1440) & (!sk[100]) & (g1441)) + ((!g165) & (g166) & (!g1439) & (!g1440) & (!sk[100]) & (!g1441)) + ((!g165) & (g166) & (!g1439) & (!g1440) & (!sk[100]) & (g1441)) + ((!g165) & (g166) & (!g1439) & (!g1440) & (sk[100]) & (g1441)) + ((!g165) & (g166) & (!g1439) & (g1440) & (!sk[100]) & (!g1441)) + ((!g165) & (g166) & (!g1439) & (g1440) & (!sk[100]) & (g1441)) + ((!g165) & (g166) & (!g1439) & (g1440) & (sk[100]) & (g1441)) + ((!g165) & (g166) & (g1439) & (!g1440) & (!sk[100]) & (!g1441)) + ((!g165) & (g166) & (g1439) & (!g1440) & (!sk[100]) & (g1441)) + ((!g165) & (g166) & (g1439) & (!g1440) & (sk[100]) & (g1441)) + ((!g165) & (g166) & (g1439) & (g1440) & (!sk[100]) & (!g1441)) + ((!g165) & (g166) & (g1439) & (g1440) & (!sk[100]) & (g1441)) + ((!g165) & (g166) & (g1439) & (g1440) & (sk[100]) & (g1441)) + ((g165) & (!g166) & (!g1439) & (g1440) & (!sk[100]) & (!g1441)) + ((g165) & (!g166) & (!g1439) & (g1440) & (!sk[100]) & (g1441)) + ((g165) & (!g166) & (g1439) & (!g1440) & (!sk[100]) & (!g1441)) + ((g165) & (!g166) & (g1439) & (!g1440) & (!sk[100]) & (g1441)) + ((g165) & (!g166) & (g1439) & (!g1440) & (sk[100]) & (!g1441)) + ((g165) & (!g166) & (g1439) & (!g1440) & (sk[100]) & (g1441)) + ((g165) & (!g166) & (g1439) & (g1440) & (!sk[100]) & (!g1441)) + ((g165) & (!g166) & (g1439) & (g1440) & (!sk[100]) & (g1441)) + ((g165) & (!g166) & (g1439) & (g1440) & (sk[100]) & (!g1441)) + ((g165) & (!g166) & (g1439) & (g1440) & (sk[100]) & (g1441)) + ((g165) & (g166) & (!g1439) & (!g1440) & (!sk[100]) & (!g1441)) + ((g165) & (g166) & (!g1439) & (!g1440) & (!sk[100]) & (g1441)) + ((g165) & (g166) & (!g1439) & (g1440) & (!sk[100]) & (!g1441)) + ((g165) & (g166) & (!g1439) & (g1440) & (!sk[100]) & (g1441)) + ((g165) & (g166) & (!g1439) & (g1440) & (sk[100]) & (!g1441)) + ((g165) & (g166) & (!g1439) & (g1440) & (sk[100]) & (g1441)) + ((g165) & (g166) & (g1439) & (!g1440) & (!sk[100]) & (!g1441)) + ((g165) & (g166) & (g1439) & (!g1440) & (!sk[100]) & (g1441)) + ((g165) & (g166) & (g1439) & (g1440) & (!sk[100]) & (!g1441)) + ((g165) & (g166) & (g1439) & (g1440) & (!sk[100]) & (g1441)) + ((g165) & (g166) & (g1439) & (g1440) & (sk[100]) & (!g1441)) + ((g165) & (g166) & (g1439) & (g1440) & (sk[100]) & (g1441)));
	assign g4913 = (((!g2162) & (!g2787) & (!sk[101]) & (g1443)) + ((!g2162) & (!g2787) & (sk[101]) & (g1443)) + ((!g2162) & (g2787) & (!sk[101]) & (!g1443)) + ((!g2162) & (g2787) & (!sk[101]) & (g1443)) + ((!g2162) & (g2787) & (sk[101]) & (g1443)) + ((g2162) & (!g2787) & (!sk[101]) & (g1443)) + ((g2162) & (g2787) & (!sk[101]) & (!g1443)) + ((g2162) & (g2787) & (!sk[101]) & (g1443)) + ((g2162) & (g2787) & (sk[101]) & (!g1443)) + ((g2162) & (g2787) & (sk[101]) & (g1443)));
	assign g4914 = (((!g2164) & (!g2787) & (!sk[102]) & (g1444)) + ((!g2164) & (!g2787) & (sk[102]) & (g1444)) + ((!g2164) & (g2787) & (!sk[102]) & (!g1444)) + ((!g2164) & (g2787) & (!sk[102]) & (g1444)) + ((!g2164) & (g2787) & (sk[102]) & (g1444)) + ((g2164) & (!g2787) & (!sk[102]) & (g1444)) + ((g2164) & (g2787) & (!sk[102]) & (!g1444)) + ((g2164) & (g2787) & (!sk[102]) & (g1444)) + ((g2164) & (g2787) & (sk[102]) & (!g1444)) + ((g2164) & (g2787) & (sk[102]) & (g1444)));
	assign g4915 = (((!g2166) & (!sk[103]) & (!g2787) & (g1445)) + ((!g2166) & (!sk[103]) & (g2787) & (!g1445)) + ((!g2166) & (!sk[103]) & (g2787) & (g1445)) + ((!g2166) & (sk[103]) & (!g2787) & (g1445)) + ((!g2166) & (sk[103]) & (g2787) & (g1445)) + ((g2166) & (!sk[103]) & (!g2787) & (g1445)) + ((g2166) & (!sk[103]) & (g2787) & (!g1445)) + ((g2166) & (!sk[103]) & (g2787) & (g1445)) + ((g2166) & (sk[103]) & (g2787) & (!g1445)) + ((g2166) & (sk[103]) & (g2787) & (g1445)));
	assign g4916 = (((!g2168) & (!g2787) & (!sk[104]) & (g1446)) + ((!g2168) & (!g2787) & (sk[104]) & (g1446)) + ((!g2168) & (g2787) & (!sk[104]) & (!g1446)) + ((!g2168) & (g2787) & (!sk[104]) & (g1446)) + ((!g2168) & (g2787) & (sk[104]) & (g1446)) + ((g2168) & (!g2787) & (!sk[104]) & (g1446)) + ((g2168) & (g2787) & (!sk[104]) & (!g1446)) + ((g2168) & (g2787) & (!sk[104]) & (g1446)) + ((g2168) & (g2787) & (sk[104]) & (!g1446)) + ((g2168) & (g2787) & (sk[104]) & (g1446)));
	assign g1447 = (((!g1443) & (!g1444) & (!g1445) & (g1446) & (g165) & (g166)) + ((!g1443) & (!g1444) & (g1445) & (!g1446) & (!g165) & (g166)) + ((!g1443) & (!g1444) & (g1445) & (g1446) & (!g165) & (g166)) + ((!g1443) & (!g1444) & (g1445) & (g1446) & (g165) & (g166)) + ((!g1443) & (g1444) & (!g1445) & (!g1446) & (g165) & (!g166)) + ((!g1443) & (g1444) & (!g1445) & (g1446) & (g165) & (!g166)) + ((!g1443) & (g1444) & (!g1445) & (g1446) & (g165) & (g166)) + ((!g1443) & (g1444) & (g1445) & (!g1446) & (!g165) & (g166)) + ((!g1443) & (g1444) & (g1445) & (!g1446) & (g165) & (!g166)) + ((!g1443) & (g1444) & (g1445) & (g1446) & (!g165) & (g166)) + ((!g1443) & (g1444) & (g1445) & (g1446) & (g165) & (!g166)) + ((!g1443) & (g1444) & (g1445) & (g1446) & (g165) & (g166)) + ((g1443) & (!g1444) & (!g1445) & (!g1446) & (!g165) & (!g166)) + ((g1443) & (!g1444) & (!g1445) & (g1446) & (!g165) & (!g166)) + ((g1443) & (!g1444) & (!g1445) & (g1446) & (g165) & (g166)) + ((g1443) & (!g1444) & (g1445) & (!g1446) & (!g165) & (!g166)) + ((g1443) & (!g1444) & (g1445) & (!g1446) & (!g165) & (g166)) + ((g1443) & (!g1444) & (g1445) & (g1446) & (!g165) & (!g166)) + ((g1443) & (!g1444) & (g1445) & (g1446) & (!g165) & (g166)) + ((g1443) & (!g1444) & (g1445) & (g1446) & (g165) & (g166)) + ((g1443) & (g1444) & (!g1445) & (!g1446) & (!g165) & (!g166)) + ((g1443) & (g1444) & (!g1445) & (!g1446) & (g165) & (!g166)) + ((g1443) & (g1444) & (!g1445) & (g1446) & (!g165) & (!g166)) + ((g1443) & (g1444) & (!g1445) & (g1446) & (g165) & (!g166)) + ((g1443) & (g1444) & (!g1445) & (g1446) & (g165) & (g166)) + ((g1443) & (g1444) & (g1445) & (!g1446) & (!g165) & (!g166)) + ((g1443) & (g1444) & (g1445) & (!g1446) & (!g165) & (g166)) + ((g1443) & (g1444) & (g1445) & (!g1446) & (g165) & (!g166)) + ((g1443) & (g1444) & (g1445) & (g1446) & (!g165) & (!g166)) + ((g1443) & (g1444) & (g1445) & (g1446) & (!g165) & (g166)) + ((g1443) & (g1444) & (g1445) & (g1446) & (g165) & (!g166)) + ((g1443) & (g1444) & (g1445) & (g1446) & (g165) & (g166)));
	assign g4917 = (((!g2169) & (!sk[106]) & (!g2787) & (g1448)) + ((!g2169) & (!sk[106]) & (g2787) & (!g1448)) + ((!g2169) & (!sk[106]) & (g2787) & (g1448)) + ((!g2169) & (sk[106]) & (!g2787) & (g1448)) + ((!g2169) & (sk[106]) & (g2787) & (g1448)) + ((g2169) & (!sk[106]) & (!g2787) & (g1448)) + ((g2169) & (!sk[106]) & (g2787) & (!g1448)) + ((g2169) & (!sk[106]) & (g2787) & (g1448)) + ((g2169) & (sk[106]) & (g2787) & (!g1448)) + ((g2169) & (sk[106]) & (g2787) & (g1448)));
	assign g4918 = (((!g2170) & (!g2787) & (!sk[107]) & (g1449)) + ((!g2170) & (!g2787) & (sk[107]) & (g1449)) + ((!g2170) & (g2787) & (!sk[107]) & (!g1449)) + ((!g2170) & (g2787) & (!sk[107]) & (g1449)) + ((!g2170) & (g2787) & (sk[107]) & (g1449)) + ((g2170) & (!g2787) & (!sk[107]) & (g1449)) + ((g2170) & (g2787) & (!sk[107]) & (!g1449)) + ((g2170) & (g2787) & (!sk[107]) & (g1449)) + ((g2170) & (g2787) & (sk[107]) & (!g1449)) + ((g2170) & (g2787) & (sk[107]) & (g1449)));
	assign g4919 = (((!g2171) & (!g2787) & (!sk[108]) & (g1450)) + ((!g2171) & (!g2787) & (sk[108]) & (g1450)) + ((!g2171) & (g2787) & (!sk[108]) & (!g1450)) + ((!g2171) & (g2787) & (!sk[108]) & (g1450)) + ((!g2171) & (g2787) & (sk[108]) & (g1450)) + ((g2171) & (!g2787) & (!sk[108]) & (g1450)) + ((g2171) & (g2787) & (!sk[108]) & (!g1450)) + ((g2171) & (g2787) & (!sk[108]) & (g1450)) + ((g2171) & (g2787) & (sk[108]) & (!g1450)) + ((g2171) & (g2787) & (sk[108]) & (g1450)));
	assign g4920 = (((!g2172) & (!g2787) & (!sk[109]) & (g1451)) + ((!g2172) & (!g2787) & (sk[109]) & (g1451)) + ((!g2172) & (g2787) & (!sk[109]) & (!g1451)) + ((!g2172) & (g2787) & (!sk[109]) & (g1451)) + ((!g2172) & (g2787) & (sk[109]) & (g1451)) + ((g2172) & (!g2787) & (!sk[109]) & (g1451)) + ((g2172) & (g2787) & (!sk[109]) & (!g1451)) + ((g2172) & (g2787) & (!sk[109]) & (g1451)) + ((g2172) & (g2787) & (sk[109]) & (!g1451)) + ((g2172) & (g2787) & (sk[109]) & (g1451)));
	assign g1452 = (((!g1448) & (!g1449) & (!g1450) & (g1451) & (g165) & (g166)) + ((!g1448) & (!g1449) & (g1450) & (!g1451) & (!g165) & (g166)) + ((!g1448) & (!g1449) & (g1450) & (g1451) & (!g165) & (g166)) + ((!g1448) & (!g1449) & (g1450) & (g1451) & (g165) & (g166)) + ((!g1448) & (g1449) & (!g1450) & (!g1451) & (g165) & (!g166)) + ((!g1448) & (g1449) & (!g1450) & (g1451) & (g165) & (!g166)) + ((!g1448) & (g1449) & (!g1450) & (g1451) & (g165) & (g166)) + ((!g1448) & (g1449) & (g1450) & (!g1451) & (!g165) & (g166)) + ((!g1448) & (g1449) & (g1450) & (!g1451) & (g165) & (!g166)) + ((!g1448) & (g1449) & (g1450) & (g1451) & (!g165) & (g166)) + ((!g1448) & (g1449) & (g1450) & (g1451) & (g165) & (!g166)) + ((!g1448) & (g1449) & (g1450) & (g1451) & (g165) & (g166)) + ((g1448) & (!g1449) & (!g1450) & (!g1451) & (!g165) & (!g166)) + ((g1448) & (!g1449) & (!g1450) & (g1451) & (!g165) & (!g166)) + ((g1448) & (!g1449) & (!g1450) & (g1451) & (g165) & (g166)) + ((g1448) & (!g1449) & (g1450) & (!g1451) & (!g165) & (!g166)) + ((g1448) & (!g1449) & (g1450) & (!g1451) & (!g165) & (g166)) + ((g1448) & (!g1449) & (g1450) & (g1451) & (!g165) & (!g166)) + ((g1448) & (!g1449) & (g1450) & (g1451) & (!g165) & (g166)) + ((g1448) & (!g1449) & (g1450) & (g1451) & (g165) & (g166)) + ((g1448) & (g1449) & (!g1450) & (!g1451) & (!g165) & (!g166)) + ((g1448) & (g1449) & (!g1450) & (!g1451) & (g165) & (!g166)) + ((g1448) & (g1449) & (!g1450) & (g1451) & (!g165) & (!g166)) + ((g1448) & (g1449) & (!g1450) & (g1451) & (g165) & (!g166)) + ((g1448) & (g1449) & (!g1450) & (g1451) & (g165) & (g166)) + ((g1448) & (g1449) & (g1450) & (!g1451) & (!g165) & (!g166)) + ((g1448) & (g1449) & (g1450) & (!g1451) & (!g165) & (g166)) + ((g1448) & (g1449) & (g1450) & (!g1451) & (g165) & (!g166)) + ((g1448) & (g1449) & (g1450) & (g1451) & (!g165) & (!g166)) + ((g1448) & (g1449) & (g1450) & (g1451) & (!g165) & (g166)) + ((g1448) & (g1449) & (g1450) & (g1451) & (g165) & (!g166)) + ((g1448) & (g1449) & (g1450) & (g1451) & (g165) & (g166)));
	assign g1453 = (((!g147) & (!g148) & (!g1438) & (g1442) & (!g1447) & (!g1452)) + ((!g147) & (!g148) & (!g1438) & (g1442) & (!g1447) & (g1452)) + ((!g147) & (!g148) & (!g1438) & (g1442) & (g1447) & (!g1452)) + ((!g147) & (!g148) & (!g1438) & (g1442) & (g1447) & (g1452)) + ((!g147) & (!g148) & (g1438) & (g1442) & (!g1447) & (!g1452)) + ((!g147) & (!g148) & (g1438) & (g1442) & (!g1447) & (g1452)) + ((!g147) & (!g148) & (g1438) & (g1442) & (g1447) & (!g1452)) + ((!g147) & (!g148) & (g1438) & (g1442) & (g1447) & (g1452)) + ((!g147) & (g148) & (!g1438) & (!g1442) & (!g1447) & (g1452)) + ((!g147) & (g148) & (!g1438) & (!g1442) & (g1447) & (g1452)) + ((!g147) & (g148) & (!g1438) & (g1442) & (!g1447) & (g1452)) + ((!g147) & (g148) & (!g1438) & (g1442) & (g1447) & (g1452)) + ((!g147) & (g148) & (g1438) & (!g1442) & (!g1447) & (g1452)) + ((!g147) & (g148) & (g1438) & (!g1442) & (g1447) & (g1452)) + ((!g147) & (g148) & (g1438) & (g1442) & (!g1447) & (g1452)) + ((!g147) & (g148) & (g1438) & (g1442) & (g1447) & (g1452)) + ((g147) & (!g148) & (g1438) & (!g1442) & (!g1447) & (!g1452)) + ((g147) & (!g148) & (g1438) & (!g1442) & (!g1447) & (g1452)) + ((g147) & (!g148) & (g1438) & (!g1442) & (g1447) & (!g1452)) + ((g147) & (!g148) & (g1438) & (!g1442) & (g1447) & (g1452)) + ((g147) & (!g148) & (g1438) & (g1442) & (!g1447) & (!g1452)) + ((g147) & (!g148) & (g1438) & (g1442) & (!g1447) & (g1452)) + ((g147) & (!g148) & (g1438) & (g1442) & (g1447) & (!g1452)) + ((g147) & (!g148) & (g1438) & (g1442) & (g1447) & (g1452)) + ((g147) & (g148) & (!g1438) & (!g1442) & (g1447) & (!g1452)) + ((g147) & (g148) & (!g1438) & (!g1442) & (g1447) & (g1452)) + ((g147) & (g148) & (!g1438) & (g1442) & (g1447) & (!g1452)) + ((g147) & (g148) & (!g1438) & (g1442) & (g1447) & (g1452)) + ((g147) & (g148) & (g1438) & (!g1442) & (g1447) & (!g1452)) + ((g147) & (g148) & (g1438) & (!g1442) & (g1447) & (g1452)) + ((g147) & (g148) & (g1438) & (g1442) & (g1447) & (!g1452)) + ((g147) & (g148) & (g1438) & (g1442) & (g1447) & (g1452)));
	assign g1454 = (((!g142) & (!sk[112]) & (!g1433) & (g1453)) + ((!g142) & (!sk[112]) & (g1433) & (!g1453)) + ((!g142) & (!sk[112]) & (g1433) & (g1453)) + ((!g142) & (sk[112]) & (!g1433) & (g1453)) + ((!g142) & (sk[112]) & (g1433) & (g1453)) + ((g142) & (!sk[112]) & (!g1433) & (g1453)) + ((g142) & (!sk[112]) & (g1433) & (!g1453)) + ((g142) & (!sk[112]) & (g1433) & (g1453)) + ((g142) & (sk[112]) & (g1433) & (!g1453)) + ((g142) & (sk[112]) & (g1433) & (g1453)));
	assign g4921 = (((!g2059) & (!g2793) & (!sk[113]) & (g1455)) + ((!g2059) & (!g2793) & (sk[113]) & (g1455)) + ((!g2059) & (g2793) & (!sk[113]) & (!g1455)) + ((!g2059) & (g2793) & (!sk[113]) & (g1455)) + ((!g2059) & (g2793) & (sk[113]) & (g1455)) + ((g2059) & (!g2793) & (!sk[113]) & (g1455)) + ((g2059) & (g2793) & (!sk[113]) & (!g1455)) + ((g2059) & (g2793) & (!sk[113]) & (g1455)) + ((g2059) & (g2793) & (sk[113]) & (!g1455)) + ((g2059) & (g2793) & (sk[113]) & (g1455)));
	assign g1456 = (((!sk[114]) & (!g1364) & (!g1409) & (!g3823) & (g1366) & (!g916)) + ((!sk[114]) & (!g1364) & (!g1409) & (!g3823) & (g1366) & (g916)) + ((!sk[114]) & (!g1364) & (!g1409) & (g3823) & (!g1366) & (!g916)) + ((!sk[114]) & (!g1364) & (!g1409) & (g3823) & (!g1366) & (g916)) + ((!sk[114]) & (!g1364) & (!g1409) & (g3823) & (g1366) & (!g916)) + ((!sk[114]) & (!g1364) & (!g1409) & (g3823) & (g1366) & (g916)) + ((!sk[114]) & (!g1364) & (g1409) & (!g3823) & (!g1366) & (!g916)) + ((!sk[114]) & (!g1364) & (g1409) & (!g3823) & (!g1366) & (g916)) + ((!sk[114]) & (!g1364) & (g1409) & (!g3823) & (g1366) & (!g916)) + ((!sk[114]) & (!g1364) & (g1409) & (!g3823) & (g1366) & (g916)) + ((!sk[114]) & (!g1364) & (g1409) & (g3823) & (!g1366) & (!g916)) + ((!sk[114]) & (!g1364) & (g1409) & (g3823) & (!g1366) & (g916)) + ((!sk[114]) & (!g1364) & (g1409) & (g3823) & (g1366) & (!g916)) + ((!sk[114]) & (!g1364) & (g1409) & (g3823) & (g1366) & (g916)) + ((!sk[114]) & (g1364) & (!g1409) & (!g3823) & (g1366) & (!g916)) + ((!sk[114]) & (g1364) & (!g1409) & (!g3823) & (g1366) & (g916)) + ((!sk[114]) & (g1364) & (!g1409) & (g3823) & (!g1366) & (!g916)) + ((!sk[114]) & (g1364) & (!g1409) & (g3823) & (!g1366) & (g916)) + ((!sk[114]) & (g1364) & (!g1409) & (g3823) & (g1366) & (!g916)) + ((!sk[114]) & (g1364) & (!g1409) & (g3823) & (g1366) & (g916)) + ((!sk[114]) & (g1364) & (g1409) & (!g3823) & (!g1366) & (!g916)) + ((!sk[114]) & (g1364) & (g1409) & (!g3823) & (!g1366) & (g916)) + ((!sk[114]) & (g1364) & (g1409) & (!g3823) & (g1366) & (!g916)) + ((!sk[114]) & (g1364) & (g1409) & (!g3823) & (g1366) & (g916)) + ((!sk[114]) & (g1364) & (g1409) & (g3823) & (!g1366) & (!g916)) + ((!sk[114]) & (g1364) & (g1409) & (g3823) & (!g1366) & (g916)) + ((!sk[114]) & (g1364) & (g1409) & (g3823) & (g1366) & (!g916)) + ((!sk[114]) & (g1364) & (g1409) & (g3823) & (g1366) & (g916)) + ((sk[114]) & (!g1364) & (!g1409) & (!g3823) & (!g1366) & (!g916)) + ((sk[114]) & (!g1364) & (!g1409) & (!g3823) & (!g1366) & (g916)) + ((sk[114]) & (!g1364) & (!g1409) & (!g3823) & (g1366) & (g916)) + ((sk[114]) & (!g1364) & (!g1409) & (g3823) & (!g1366) & (g916)) + ((sk[114]) & (!g1364) & (!g1409) & (g3823) & (g1366) & (g916)) + ((sk[114]) & (!g1364) & (g1409) & (!g3823) & (!g1366) & (g916)) + ((sk[114]) & (!g1364) & (g1409) & (!g3823) & (g1366) & (g916)) + ((sk[114]) & (!g1364) & (g1409) & (g3823) & (!g1366) & (g916)) + ((sk[114]) & (!g1364) & (g1409) & (g3823) & (g1366) & (g916)) + ((sk[114]) & (g1364) & (!g1409) & (!g3823) & (!g1366) & (g916)) + ((sk[114]) & (g1364) & (!g1409) & (!g3823) & (g1366) & (g916)) + ((sk[114]) & (g1364) & (!g1409) & (g3823) & (!g1366) & (g916)) + ((sk[114]) & (g1364) & (!g1409) & (g3823) & (g1366) & (g916)) + ((sk[114]) & (g1364) & (g1409) & (!g3823) & (!g1366) & (g916)));
	assign g1457 = (((!g126) & (!g1454) & (!sk[115]) & (!g1455) & (g1456) & (!g916)) + ((!g126) & (!g1454) & (!sk[115]) & (!g1455) & (g1456) & (g916)) + ((!g126) & (!g1454) & (!sk[115]) & (g1455) & (!g1456) & (!g916)) + ((!g126) & (!g1454) & (!sk[115]) & (g1455) & (!g1456) & (g916)) + ((!g126) & (!g1454) & (!sk[115]) & (g1455) & (g1456) & (!g916)) + ((!g126) & (!g1454) & (!sk[115]) & (g1455) & (g1456) & (g916)) + ((!g126) & (!g1454) & (sk[115]) & (g1455) & (!g1456) & (!g916)) + ((!g126) & (!g1454) & (sk[115]) & (g1455) & (!g1456) & (g916)) + ((!g126) & (!g1454) & (sk[115]) & (g1455) & (g1456) & (!g916)) + ((!g126) & (!g1454) & (sk[115]) & (g1455) & (g1456) & (g916)) + ((!g126) & (g1454) & (!sk[115]) & (!g1455) & (!g1456) & (!g916)) + ((!g126) & (g1454) & (!sk[115]) & (!g1455) & (!g1456) & (g916)) + ((!g126) & (g1454) & (!sk[115]) & (!g1455) & (g1456) & (!g916)) + ((!g126) & (g1454) & (!sk[115]) & (!g1455) & (g1456) & (g916)) + ((!g126) & (g1454) & (!sk[115]) & (g1455) & (!g1456) & (!g916)) + ((!g126) & (g1454) & (!sk[115]) & (g1455) & (!g1456) & (g916)) + ((!g126) & (g1454) & (!sk[115]) & (g1455) & (g1456) & (!g916)) + ((!g126) & (g1454) & (!sk[115]) & (g1455) & (g1456) & (g916)) + ((!g126) & (g1454) & (sk[115]) & (g1455) & (!g1456) & (!g916)) + ((!g126) & (g1454) & (sk[115]) & (g1455) & (!g1456) & (g916)) + ((!g126) & (g1454) & (sk[115]) & (g1455) & (g1456) & (!g916)) + ((!g126) & (g1454) & (sk[115]) & (g1455) & (g1456) & (g916)) + ((g126) & (!g1454) & (!sk[115]) & (!g1455) & (g1456) & (!g916)) + ((g126) & (!g1454) & (!sk[115]) & (!g1455) & (g1456) & (g916)) + ((g126) & (!g1454) & (!sk[115]) & (g1455) & (!g1456) & (!g916)) + ((g126) & (!g1454) & (!sk[115]) & (g1455) & (!g1456) & (g916)) + ((g126) & (!g1454) & (!sk[115]) & (g1455) & (g1456) & (!g916)) + ((g126) & (!g1454) & (!sk[115]) & (g1455) & (g1456) & (g916)) + ((g126) & (!g1454) & (sk[115]) & (!g1455) & (!g1456) & (g916)) + ((g126) & (!g1454) & (sk[115]) & (!g1455) & (g1456) & (!g916)) + ((g126) & (!g1454) & (sk[115]) & (g1455) & (!g1456) & (g916)) + ((g126) & (!g1454) & (sk[115]) & (g1455) & (g1456) & (!g916)) + ((g126) & (g1454) & (!sk[115]) & (!g1455) & (!g1456) & (!g916)) + ((g126) & (g1454) & (!sk[115]) & (!g1455) & (!g1456) & (g916)) + ((g126) & (g1454) & (!sk[115]) & (!g1455) & (g1456) & (!g916)) + ((g126) & (g1454) & (!sk[115]) & (!g1455) & (g1456) & (g916)) + ((g126) & (g1454) & (!sk[115]) & (g1455) & (!g1456) & (!g916)) + ((g126) & (g1454) & (!sk[115]) & (g1455) & (!g1456) & (g916)) + ((g126) & (g1454) & (!sk[115]) & (g1455) & (g1456) & (!g916)) + ((g126) & (g1454) & (!sk[115]) & (g1455) & (g1456) & (g916)) + ((g126) & (g1454) & (sk[115]) & (!g1455) & (!g1456) & (!g916)) + ((g126) & (g1454) & (sk[115]) & (!g1455) & (g1456) & (g916)) + ((g126) & (g1454) & (sk[115]) & (g1455) & (!g1456) & (!g916)) + ((g126) & (g1454) & (sk[115]) & (g1455) & (g1456) & (g916)));
	assign g4922 = (((!g2140) & (!g2805) & (!sk[116]) & (g1458)) + ((!g2140) & (!g2805) & (sk[116]) & (g1458)) + ((!g2140) & (g2805) & (!sk[116]) & (!g1458)) + ((!g2140) & (g2805) & (!sk[116]) & (g1458)) + ((!g2140) & (g2805) & (sk[116]) & (g1458)) + ((g2140) & (!g2805) & (!sk[116]) & (g1458)) + ((g2140) & (g2805) & (!sk[116]) & (!g1458)) + ((g2140) & (g2805) & (!sk[116]) & (g1458)) + ((g2140) & (g2805) & (sk[116]) & (!g1458)) + ((g2140) & (g2805) & (sk[116]) & (g1458)));
	assign g4923 = (((!g2142) & (!g2805) & (!sk[117]) & (g1459)) + ((!g2142) & (!g2805) & (sk[117]) & (g1459)) + ((!g2142) & (g2805) & (!sk[117]) & (!g1459)) + ((!g2142) & (g2805) & (!sk[117]) & (g1459)) + ((!g2142) & (g2805) & (sk[117]) & (g1459)) + ((g2142) & (!g2805) & (!sk[117]) & (g1459)) + ((g2142) & (g2805) & (!sk[117]) & (!g1459)) + ((g2142) & (g2805) & (!sk[117]) & (g1459)) + ((g2142) & (g2805) & (sk[117]) & (!g1459)) + ((g2142) & (g2805) & (sk[117]) & (g1459)));
	assign g4924 = (((!g2144) & (!g2805) & (!sk[118]) & (g1460)) + ((!g2144) & (!g2805) & (sk[118]) & (g1460)) + ((!g2144) & (g2805) & (!sk[118]) & (!g1460)) + ((!g2144) & (g2805) & (!sk[118]) & (g1460)) + ((!g2144) & (g2805) & (sk[118]) & (g1460)) + ((g2144) & (!g2805) & (!sk[118]) & (g1460)) + ((g2144) & (g2805) & (!sk[118]) & (!g1460)) + ((g2144) & (g2805) & (!sk[118]) & (g1460)) + ((g2144) & (g2805) & (sk[118]) & (!g1460)) + ((g2144) & (g2805) & (sk[118]) & (g1460)));
	assign g4925 = (((!g2145) & (!g2805) & (!sk[119]) & (g1461)) + ((!g2145) & (!g2805) & (sk[119]) & (g1461)) + ((!g2145) & (g2805) & (!sk[119]) & (!g1461)) + ((!g2145) & (g2805) & (!sk[119]) & (g1461)) + ((!g2145) & (g2805) & (sk[119]) & (g1461)) + ((g2145) & (!g2805) & (!sk[119]) & (g1461)) + ((g2145) & (g2805) & (!sk[119]) & (!g1461)) + ((g2145) & (g2805) & (!sk[119]) & (g1461)) + ((g2145) & (g2805) & (sk[119]) & (!g1461)) + ((g2145) & (g2805) & (sk[119]) & (g1461)));
	assign g1462 = (((!g1458) & (!g1459) & (!g1460) & (g1461) & (g147) & (g148)) + ((!g1458) & (!g1459) & (g1460) & (!g1461) & (!g147) & (g148)) + ((!g1458) & (!g1459) & (g1460) & (g1461) & (!g147) & (g148)) + ((!g1458) & (!g1459) & (g1460) & (g1461) & (g147) & (g148)) + ((!g1458) & (g1459) & (!g1460) & (!g1461) & (g147) & (!g148)) + ((!g1458) & (g1459) & (!g1460) & (g1461) & (g147) & (!g148)) + ((!g1458) & (g1459) & (!g1460) & (g1461) & (g147) & (g148)) + ((!g1458) & (g1459) & (g1460) & (!g1461) & (!g147) & (g148)) + ((!g1458) & (g1459) & (g1460) & (!g1461) & (g147) & (!g148)) + ((!g1458) & (g1459) & (g1460) & (g1461) & (!g147) & (g148)) + ((!g1458) & (g1459) & (g1460) & (g1461) & (g147) & (!g148)) + ((!g1458) & (g1459) & (g1460) & (g1461) & (g147) & (g148)) + ((g1458) & (!g1459) & (!g1460) & (!g1461) & (!g147) & (!g148)) + ((g1458) & (!g1459) & (!g1460) & (g1461) & (!g147) & (!g148)) + ((g1458) & (!g1459) & (!g1460) & (g1461) & (g147) & (g148)) + ((g1458) & (!g1459) & (g1460) & (!g1461) & (!g147) & (!g148)) + ((g1458) & (!g1459) & (g1460) & (!g1461) & (!g147) & (g148)) + ((g1458) & (!g1459) & (g1460) & (g1461) & (!g147) & (!g148)) + ((g1458) & (!g1459) & (g1460) & (g1461) & (!g147) & (g148)) + ((g1458) & (!g1459) & (g1460) & (g1461) & (g147) & (g148)) + ((g1458) & (g1459) & (!g1460) & (!g1461) & (!g147) & (!g148)) + ((g1458) & (g1459) & (!g1460) & (!g1461) & (g147) & (!g148)) + ((g1458) & (g1459) & (!g1460) & (g1461) & (!g147) & (!g148)) + ((g1458) & (g1459) & (!g1460) & (g1461) & (g147) & (!g148)) + ((g1458) & (g1459) & (!g1460) & (g1461) & (g147) & (g148)) + ((g1458) & (g1459) & (g1460) & (!g1461) & (!g147) & (!g148)) + ((g1458) & (g1459) & (g1460) & (!g1461) & (!g147) & (g148)) + ((g1458) & (g1459) & (g1460) & (!g1461) & (g147) & (!g148)) + ((g1458) & (g1459) & (g1460) & (g1461) & (!g147) & (!g148)) + ((g1458) & (g1459) & (g1460) & (g1461) & (!g147) & (g148)) + ((g1458) & (g1459) & (g1460) & (g1461) & (g147) & (!g148)) + ((g1458) & (g1459) & (g1460) & (g1461) & (g147) & (g148)));
	assign g4926 = (((!sk[121]) & (!g2146) & (!g2805) & (g1463)) + ((!sk[121]) & (!g2146) & (g2805) & (!g1463)) + ((!sk[121]) & (!g2146) & (g2805) & (g1463)) + ((!sk[121]) & (g2146) & (!g2805) & (g1463)) + ((!sk[121]) & (g2146) & (g2805) & (!g1463)) + ((!sk[121]) & (g2146) & (g2805) & (g1463)) + ((sk[121]) & (!g2146) & (!g2805) & (g1463)) + ((sk[121]) & (!g2146) & (g2805) & (g1463)) + ((sk[121]) & (g2146) & (g2805) & (!g1463)) + ((sk[121]) & (g2146) & (g2805) & (g1463)));
	assign g4927 = (((!g2148) & (!sk[122]) & (!g2805) & (g1464)) + ((!g2148) & (!sk[122]) & (g2805) & (!g1464)) + ((!g2148) & (!sk[122]) & (g2805) & (g1464)) + ((!g2148) & (sk[122]) & (!g2805) & (g1464)) + ((!g2148) & (sk[122]) & (g2805) & (g1464)) + ((g2148) & (!sk[122]) & (!g2805) & (g1464)) + ((g2148) & (!sk[122]) & (g2805) & (!g1464)) + ((g2148) & (!sk[122]) & (g2805) & (g1464)) + ((g2148) & (sk[122]) & (g2805) & (!g1464)) + ((g2148) & (sk[122]) & (g2805) & (g1464)));
	assign g4928 = (((!g2150) & (!sk[123]) & (!g2805) & (g1465)) + ((!g2150) & (!sk[123]) & (g2805) & (!g1465)) + ((!g2150) & (!sk[123]) & (g2805) & (g1465)) + ((!g2150) & (sk[123]) & (!g2805) & (g1465)) + ((!g2150) & (sk[123]) & (g2805) & (g1465)) + ((g2150) & (!sk[123]) & (!g2805) & (g1465)) + ((g2150) & (!sk[123]) & (g2805) & (!g1465)) + ((g2150) & (!sk[123]) & (g2805) & (g1465)) + ((g2150) & (sk[123]) & (g2805) & (!g1465)) + ((g2150) & (sk[123]) & (g2805) & (g1465)));
	assign g4929 = (((!g2151) & (!g2805) & (!sk[124]) & (g1466)) + ((!g2151) & (!g2805) & (sk[124]) & (g1466)) + ((!g2151) & (g2805) & (!sk[124]) & (!g1466)) + ((!g2151) & (g2805) & (!sk[124]) & (g1466)) + ((!g2151) & (g2805) & (sk[124]) & (g1466)) + ((g2151) & (!g2805) & (!sk[124]) & (g1466)) + ((g2151) & (g2805) & (!sk[124]) & (!g1466)) + ((g2151) & (g2805) & (!sk[124]) & (g1466)) + ((g2151) & (g2805) & (sk[124]) & (!g1466)) + ((g2151) & (g2805) & (sk[124]) & (g1466)));
	assign g1467 = (((!g1463) & (!g1464) & (!g1465) & (g1466) & (g147) & (g148)) + ((!g1463) & (!g1464) & (g1465) & (!g1466) & (!g147) & (g148)) + ((!g1463) & (!g1464) & (g1465) & (g1466) & (!g147) & (g148)) + ((!g1463) & (!g1464) & (g1465) & (g1466) & (g147) & (g148)) + ((!g1463) & (g1464) & (!g1465) & (!g1466) & (g147) & (!g148)) + ((!g1463) & (g1464) & (!g1465) & (g1466) & (g147) & (!g148)) + ((!g1463) & (g1464) & (!g1465) & (g1466) & (g147) & (g148)) + ((!g1463) & (g1464) & (g1465) & (!g1466) & (!g147) & (g148)) + ((!g1463) & (g1464) & (g1465) & (!g1466) & (g147) & (!g148)) + ((!g1463) & (g1464) & (g1465) & (g1466) & (!g147) & (g148)) + ((!g1463) & (g1464) & (g1465) & (g1466) & (g147) & (!g148)) + ((!g1463) & (g1464) & (g1465) & (g1466) & (g147) & (g148)) + ((g1463) & (!g1464) & (!g1465) & (!g1466) & (!g147) & (!g148)) + ((g1463) & (!g1464) & (!g1465) & (g1466) & (!g147) & (!g148)) + ((g1463) & (!g1464) & (!g1465) & (g1466) & (g147) & (g148)) + ((g1463) & (!g1464) & (g1465) & (!g1466) & (!g147) & (!g148)) + ((g1463) & (!g1464) & (g1465) & (!g1466) & (!g147) & (g148)) + ((g1463) & (!g1464) & (g1465) & (g1466) & (!g147) & (!g148)) + ((g1463) & (!g1464) & (g1465) & (g1466) & (!g147) & (g148)) + ((g1463) & (!g1464) & (g1465) & (g1466) & (g147) & (g148)) + ((g1463) & (g1464) & (!g1465) & (!g1466) & (!g147) & (!g148)) + ((g1463) & (g1464) & (!g1465) & (!g1466) & (g147) & (!g148)) + ((g1463) & (g1464) & (!g1465) & (g1466) & (!g147) & (!g148)) + ((g1463) & (g1464) & (!g1465) & (g1466) & (g147) & (!g148)) + ((g1463) & (g1464) & (!g1465) & (g1466) & (g147) & (g148)) + ((g1463) & (g1464) & (g1465) & (!g1466) & (!g147) & (!g148)) + ((g1463) & (g1464) & (g1465) & (!g1466) & (!g147) & (g148)) + ((g1463) & (g1464) & (g1465) & (!g1466) & (g147) & (!g148)) + ((g1463) & (g1464) & (g1465) & (g1466) & (!g147) & (!g148)) + ((g1463) & (g1464) & (g1465) & (g1466) & (!g147) & (g148)) + ((g1463) & (g1464) & (g1465) & (g1466) & (g147) & (!g148)) + ((g1463) & (g1464) & (g1465) & (g1466) & (g147) & (g148)));
	assign g4930 = (((!sk[126]) & (!g2152) & (!g2805) & (g1468)) + ((!sk[126]) & (!g2152) & (g2805) & (!g1468)) + ((!sk[126]) & (!g2152) & (g2805) & (g1468)) + ((!sk[126]) & (g2152) & (!g2805) & (g1468)) + ((!sk[126]) & (g2152) & (g2805) & (!g1468)) + ((!sk[126]) & (g2152) & (g2805) & (g1468)) + ((sk[126]) & (!g2152) & (!g2805) & (g1468)) + ((sk[126]) & (!g2152) & (g2805) & (g1468)) + ((sk[126]) & (g2152) & (g2805) & (!g1468)) + ((sk[126]) & (g2152) & (g2805) & (g1468)));
	assign g4931 = (((!sk[127]) & (!g2153) & (!g2805) & (g1469)) + ((!sk[127]) & (!g2153) & (g2805) & (!g1469)) + ((!sk[127]) & (!g2153) & (g2805) & (g1469)) + ((!sk[127]) & (g2153) & (!g2805) & (g1469)) + ((!sk[127]) & (g2153) & (g2805) & (!g1469)) + ((!sk[127]) & (g2153) & (g2805) & (g1469)) + ((sk[127]) & (!g2153) & (!g2805) & (g1469)) + ((sk[127]) & (!g2153) & (g2805) & (g1469)) + ((sk[127]) & (g2153) & (g2805) & (!g1469)) + ((sk[127]) & (g2153) & (g2805) & (g1469)));
	assign g4932 = (((!g2155) & (!sk[0]) & (!g2805) & (g1470)) + ((!g2155) & (!sk[0]) & (g2805) & (!g1470)) + ((!g2155) & (!sk[0]) & (g2805) & (g1470)) + ((!g2155) & (sk[0]) & (!g2805) & (g1470)) + ((!g2155) & (sk[0]) & (g2805) & (g1470)) + ((g2155) & (!sk[0]) & (!g2805) & (g1470)) + ((g2155) & (!sk[0]) & (g2805) & (!g1470)) + ((g2155) & (!sk[0]) & (g2805) & (g1470)) + ((g2155) & (sk[0]) & (g2805) & (!g1470)) + ((g2155) & (sk[0]) & (g2805) & (g1470)));
	assign g4933 = (((!g2157) & (!sk[1]) & (!g2805) & (g1471)) + ((!g2157) & (!sk[1]) & (g2805) & (!g1471)) + ((!g2157) & (!sk[1]) & (g2805) & (g1471)) + ((!g2157) & (sk[1]) & (!g2805) & (g1471)) + ((!g2157) & (sk[1]) & (g2805) & (g1471)) + ((g2157) & (!sk[1]) & (!g2805) & (g1471)) + ((g2157) & (!sk[1]) & (g2805) & (!g1471)) + ((g2157) & (!sk[1]) & (g2805) & (g1471)) + ((g2157) & (sk[1]) & (g2805) & (!g1471)) + ((g2157) & (sk[1]) & (g2805) & (g1471)));
	assign g1472 = (((!g1468) & (!g1469) & (!g1470) & (g1471) & (g147) & (g148)) + ((!g1468) & (!g1469) & (g1470) & (!g1471) & (!g147) & (g148)) + ((!g1468) & (!g1469) & (g1470) & (g1471) & (!g147) & (g148)) + ((!g1468) & (!g1469) & (g1470) & (g1471) & (g147) & (g148)) + ((!g1468) & (g1469) & (!g1470) & (!g1471) & (g147) & (!g148)) + ((!g1468) & (g1469) & (!g1470) & (g1471) & (g147) & (!g148)) + ((!g1468) & (g1469) & (!g1470) & (g1471) & (g147) & (g148)) + ((!g1468) & (g1469) & (g1470) & (!g1471) & (!g147) & (g148)) + ((!g1468) & (g1469) & (g1470) & (!g1471) & (g147) & (!g148)) + ((!g1468) & (g1469) & (g1470) & (g1471) & (!g147) & (g148)) + ((!g1468) & (g1469) & (g1470) & (g1471) & (g147) & (!g148)) + ((!g1468) & (g1469) & (g1470) & (g1471) & (g147) & (g148)) + ((g1468) & (!g1469) & (!g1470) & (!g1471) & (!g147) & (!g148)) + ((g1468) & (!g1469) & (!g1470) & (g1471) & (!g147) & (!g148)) + ((g1468) & (!g1469) & (!g1470) & (g1471) & (g147) & (g148)) + ((g1468) & (!g1469) & (g1470) & (!g1471) & (!g147) & (!g148)) + ((g1468) & (!g1469) & (g1470) & (!g1471) & (!g147) & (g148)) + ((g1468) & (!g1469) & (g1470) & (g1471) & (!g147) & (!g148)) + ((g1468) & (!g1469) & (g1470) & (g1471) & (!g147) & (g148)) + ((g1468) & (!g1469) & (g1470) & (g1471) & (g147) & (g148)) + ((g1468) & (g1469) & (!g1470) & (!g1471) & (!g147) & (!g148)) + ((g1468) & (g1469) & (!g1470) & (!g1471) & (g147) & (!g148)) + ((g1468) & (g1469) & (!g1470) & (g1471) & (!g147) & (!g148)) + ((g1468) & (g1469) & (!g1470) & (g1471) & (g147) & (!g148)) + ((g1468) & (g1469) & (!g1470) & (g1471) & (g147) & (g148)) + ((g1468) & (g1469) & (g1470) & (!g1471) & (!g147) & (!g148)) + ((g1468) & (g1469) & (g1470) & (!g1471) & (!g147) & (g148)) + ((g1468) & (g1469) & (g1470) & (!g1471) & (g147) & (!g148)) + ((g1468) & (g1469) & (g1470) & (g1471) & (!g147) & (!g148)) + ((g1468) & (g1469) & (g1470) & (g1471) & (!g147) & (g148)) + ((g1468) & (g1469) & (g1470) & (g1471) & (g147) & (!g148)) + ((g1468) & (g1469) & (g1470) & (g1471) & (g147) & (g148)));
	assign g4934 = (((!sk[3]) & (!g2158) & (!g2805) & (g1473)) + ((!sk[3]) & (!g2158) & (g2805) & (!g1473)) + ((!sk[3]) & (!g2158) & (g2805) & (g1473)) + ((!sk[3]) & (g2158) & (!g2805) & (g1473)) + ((!sk[3]) & (g2158) & (g2805) & (!g1473)) + ((!sk[3]) & (g2158) & (g2805) & (g1473)) + ((sk[3]) & (!g2158) & (!g2805) & (g1473)) + ((sk[3]) & (!g2158) & (g2805) & (g1473)) + ((sk[3]) & (g2158) & (g2805) & (!g1473)) + ((sk[3]) & (g2158) & (g2805) & (g1473)));
	assign g4935 = (((!g2159) & (!sk[4]) & (!g2805) & (g1474)) + ((!g2159) & (!sk[4]) & (g2805) & (!g1474)) + ((!g2159) & (!sk[4]) & (g2805) & (g1474)) + ((!g2159) & (sk[4]) & (!g2805) & (g1474)) + ((!g2159) & (sk[4]) & (g2805) & (g1474)) + ((g2159) & (!sk[4]) & (!g2805) & (g1474)) + ((g2159) & (!sk[4]) & (g2805) & (!g1474)) + ((g2159) & (!sk[4]) & (g2805) & (g1474)) + ((g2159) & (sk[4]) & (g2805) & (!g1474)) + ((g2159) & (sk[4]) & (g2805) & (g1474)));
	assign g4936 = (((!g2160) & (!sk[5]) & (!g2805) & (g1475)) + ((!g2160) & (!sk[5]) & (g2805) & (!g1475)) + ((!g2160) & (!sk[5]) & (g2805) & (g1475)) + ((!g2160) & (sk[5]) & (!g2805) & (g1475)) + ((!g2160) & (sk[5]) & (g2805) & (g1475)) + ((g2160) & (!sk[5]) & (!g2805) & (g1475)) + ((g2160) & (!sk[5]) & (g2805) & (!g1475)) + ((g2160) & (!sk[5]) & (g2805) & (g1475)) + ((g2160) & (sk[5]) & (g2805) & (!g1475)) + ((g2160) & (sk[5]) & (g2805) & (g1475)));
	assign g4937 = (((!g2161) & (!sk[6]) & (!g2805) & (g1476)) + ((!g2161) & (!sk[6]) & (g2805) & (!g1476)) + ((!g2161) & (!sk[6]) & (g2805) & (g1476)) + ((!g2161) & (sk[6]) & (!g2805) & (g1476)) + ((!g2161) & (sk[6]) & (g2805) & (g1476)) + ((g2161) & (!sk[6]) & (!g2805) & (g1476)) + ((g2161) & (!sk[6]) & (g2805) & (!g1476)) + ((g2161) & (!sk[6]) & (g2805) & (g1476)) + ((g2161) & (sk[6]) & (g2805) & (!g1476)) + ((g2161) & (sk[6]) & (g2805) & (g1476)));
	assign g1477 = (((!g1473) & (!g1474) & (!g1475) & (g1476) & (g147) & (g148)) + ((!g1473) & (!g1474) & (g1475) & (!g1476) & (!g147) & (g148)) + ((!g1473) & (!g1474) & (g1475) & (g1476) & (!g147) & (g148)) + ((!g1473) & (!g1474) & (g1475) & (g1476) & (g147) & (g148)) + ((!g1473) & (g1474) & (!g1475) & (!g1476) & (g147) & (!g148)) + ((!g1473) & (g1474) & (!g1475) & (g1476) & (g147) & (!g148)) + ((!g1473) & (g1474) & (!g1475) & (g1476) & (g147) & (g148)) + ((!g1473) & (g1474) & (g1475) & (!g1476) & (!g147) & (g148)) + ((!g1473) & (g1474) & (g1475) & (!g1476) & (g147) & (!g148)) + ((!g1473) & (g1474) & (g1475) & (g1476) & (!g147) & (g148)) + ((!g1473) & (g1474) & (g1475) & (g1476) & (g147) & (!g148)) + ((!g1473) & (g1474) & (g1475) & (g1476) & (g147) & (g148)) + ((g1473) & (!g1474) & (!g1475) & (!g1476) & (!g147) & (!g148)) + ((g1473) & (!g1474) & (!g1475) & (g1476) & (!g147) & (!g148)) + ((g1473) & (!g1474) & (!g1475) & (g1476) & (g147) & (g148)) + ((g1473) & (!g1474) & (g1475) & (!g1476) & (!g147) & (!g148)) + ((g1473) & (!g1474) & (g1475) & (!g1476) & (!g147) & (g148)) + ((g1473) & (!g1474) & (g1475) & (g1476) & (!g147) & (!g148)) + ((g1473) & (!g1474) & (g1475) & (g1476) & (!g147) & (g148)) + ((g1473) & (!g1474) & (g1475) & (g1476) & (g147) & (g148)) + ((g1473) & (g1474) & (!g1475) & (!g1476) & (!g147) & (!g148)) + ((g1473) & (g1474) & (!g1475) & (!g1476) & (g147) & (!g148)) + ((g1473) & (g1474) & (!g1475) & (g1476) & (!g147) & (!g148)) + ((g1473) & (g1474) & (!g1475) & (g1476) & (g147) & (!g148)) + ((g1473) & (g1474) & (!g1475) & (g1476) & (g147) & (g148)) + ((g1473) & (g1474) & (g1475) & (!g1476) & (!g147) & (!g148)) + ((g1473) & (g1474) & (g1475) & (!g1476) & (!g147) & (g148)) + ((g1473) & (g1474) & (g1475) & (!g1476) & (g147) & (!g148)) + ((g1473) & (g1474) & (g1475) & (g1476) & (!g147) & (!g148)) + ((g1473) & (g1474) & (g1475) & (g1476) & (!g147) & (g148)) + ((g1473) & (g1474) & (g1475) & (g1476) & (g147) & (!g148)) + ((g1473) & (g1474) & (g1475) & (g1476) & (g147) & (g148)));
	assign g1478 = (((!g1462) & (!g1467) & (!g1472) & (g1477) & (g165) & (g166)) + ((!g1462) & (!g1467) & (g1472) & (!g1477) & (!g165) & (g166)) + ((!g1462) & (!g1467) & (g1472) & (g1477) & (!g165) & (g166)) + ((!g1462) & (!g1467) & (g1472) & (g1477) & (g165) & (g166)) + ((!g1462) & (g1467) & (!g1472) & (!g1477) & (g165) & (!g166)) + ((!g1462) & (g1467) & (!g1472) & (g1477) & (g165) & (!g166)) + ((!g1462) & (g1467) & (!g1472) & (g1477) & (g165) & (g166)) + ((!g1462) & (g1467) & (g1472) & (!g1477) & (!g165) & (g166)) + ((!g1462) & (g1467) & (g1472) & (!g1477) & (g165) & (!g166)) + ((!g1462) & (g1467) & (g1472) & (g1477) & (!g165) & (g166)) + ((!g1462) & (g1467) & (g1472) & (g1477) & (g165) & (!g166)) + ((!g1462) & (g1467) & (g1472) & (g1477) & (g165) & (g166)) + ((g1462) & (!g1467) & (!g1472) & (!g1477) & (!g165) & (!g166)) + ((g1462) & (!g1467) & (!g1472) & (g1477) & (!g165) & (!g166)) + ((g1462) & (!g1467) & (!g1472) & (g1477) & (g165) & (g166)) + ((g1462) & (!g1467) & (g1472) & (!g1477) & (!g165) & (!g166)) + ((g1462) & (!g1467) & (g1472) & (!g1477) & (!g165) & (g166)) + ((g1462) & (!g1467) & (g1472) & (g1477) & (!g165) & (!g166)) + ((g1462) & (!g1467) & (g1472) & (g1477) & (!g165) & (g166)) + ((g1462) & (!g1467) & (g1472) & (g1477) & (g165) & (g166)) + ((g1462) & (g1467) & (!g1472) & (!g1477) & (!g165) & (!g166)) + ((g1462) & (g1467) & (!g1472) & (!g1477) & (g165) & (!g166)) + ((g1462) & (g1467) & (!g1472) & (g1477) & (!g165) & (!g166)) + ((g1462) & (g1467) & (!g1472) & (g1477) & (g165) & (!g166)) + ((g1462) & (g1467) & (!g1472) & (g1477) & (g165) & (g166)) + ((g1462) & (g1467) & (g1472) & (!g1477) & (!g165) & (!g166)) + ((g1462) & (g1467) & (g1472) & (!g1477) & (!g165) & (g166)) + ((g1462) & (g1467) & (g1472) & (!g1477) & (g165) & (!g166)) + ((g1462) & (g1467) & (g1472) & (g1477) & (!g165) & (!g166)) + ((g1462) & (g1467) & (g1472) & (g1477) & (!g165) & (g166)) + ((g1462) & (g1467) & (g1472) & (g1477) & (g165) & (!g166)) + ((g1462) & (g1467) & (g1472) & (g1477) & (g165) & (g166)));
	assign g4938 = (((!g2173) & (!g2805) & (!sk[9]) & (g1479)) + ((!g2173) & (!g2805) & (sk[9]) & (g1479)) + ((!g2173) & (g2805) & (!sk[9]) & (!g1479)) + ((!g2173) & (g2805) & (!sk[9]) & (g1479)) + ((!g2173) & (g2805) & (sk[9]) & (g1479)) + ((g2173) & (!g2805) & (!sk[9]) & (g1479)) + ((g2173) & (g2805) & (!sk[9]) & (!g1479)) + ((g2173) & (g2805) & (!sk[9]) & (g1479)) + ((g2173) & (g2805) & (sk[9]) & (!g1479)) + ((g2173) & (g2805) & (sk[9]) & (g1479)));
	assign g4939 = (((!g2174) & (!g2805) & (!sk[10]) & (g1480)) + ((!g2174) & (!g2805) & (sk[10]) & (g1480)) + ((!g2174) & (g2805) & (!sk[10]) & (!g1480)) + ((!g2174) & (g2805) & (!sk[10]) & (g1480)) + ((!g2174) & (g2805) & (sk[10]) & (g1480)) + ((g2174) & (!g2805) & (!sk[10]) & (g1480)) + ((g2174) & (g2805) & (!sk[10]) & (!g1480)) + ((g2174) & (g2805) & (!sk[10]) & (g1480)) + ((g2174) & (g2805) & (sk[10]) & (!g1480)) + ((g2174) & (g2805) & (sk[10]) & (g1480)));
	assign g4940 = (((!g2175) & (!g2805) & (!sk[11]) & (g1481)) + ((!g2175) & (!g2805) & (sk[11]) & (g1481)) + ((!g2175) & (g2805) & (!sk[11]) & (!g1481)) + ((!g2175) & (g2805) & (!sk[11]) & (g1481)) + ((!g2175) & (g2805) & (sk[11]) & (g1481)) + ((g2175) & (!g2805) & (!sk[11]) & (g1481)) + ((g2175) & (g2805) & (!sk[11]) & (!g1481)) + ((g2175) & (g2805) & (!sk[11]) & (g1481)) + ((g2175) & (g2805) & (sk[11]) & (!g1481)) + ((g2175) & (g2805) & (sk[11]) & (g1481)));
	assign g4941 = (((!sk[12]) & (!g2176) & (!g2805) & (g1482)) + ((!sk[12]) & (!g2176) & (g2805) & (!g1482)) + ((!sk[12]) & (!g2176) & (g2805) & (g1482)) + ((!sk[12]) & (g2176) & (!g2805) & (g1482)) + ((!sk[12]) & (g2176) & (g2805) & (!g1482)) + ((!sk[12]) & (g2176) & (g2805) & (g1482)) + ((sk[12]) & (!g2176) & (!g2805) & (g1482)) + ((sk[12]) & (!g2176) & (g2805) & (g1482)) + ((sk[12]) & (g2176) & (g2805) & (!g1482)) + ((sk[12]) & (g2176) & (g2805) & (g1482)));
	assign g1483 = (((!g1479) & (!g1480) & (!g1481) & (g1482) & (g165) & (g166)) + ((!g1479) & (!g1480) & (g1481) & (!g1482) & (!g165) & (g166)) + ((!g1479) & (!g1480) & (g1481) & (g1482) & (!g165) & (g166)) + ((!g1479) & (!g1480) & (g1481) & (g1482) & (g165) & (g166)) + ((!g1479) & (g1480) & (!g1481) & (!g1482) & (g165) & (!g166)) + ((!g1479) & (g1480) & (!g1481) & (g1482) & (g165) & (!g166)) + ((!g1479) & (g1480) & (!g1481) & (g1482) & (g165) & (g166)) + ((!g1479) & (g1480) & (g1481) & (!g1482) & (!g165) & (g166)) + ((!g1479) & (g1480) & (g1481) & (!g1482) & (g165) & (!g166)) + ((!g1479) & (g1480) & (g1481) & (g1482) & (!g165) & (g166)) + ((!g1479) & (g1480) & (g1481) & (g1482) & (g165) & (!g166)) + ((!g1479) & (g1480) & (g1481) & (g1482) & (g165) & (g166)) + ((g1479) & (!g1480) & (!g1481) & (!g1482) & (!g165) & (!g166)) + ((g1479) & (!g1480) & (!g1481) & (g1482) & (!g165) & (!g166)) + ((g1479) & (!g1480) & (!g1481) & (g1482) & (g165) & (g166)) + ((g1479) & (!g1480) & (g1481) & (!g1482) & (!g165) & (!g166)) + ((g1479) & (!g1480) & (g1481) & (!g1482) & (!g165) & (g166)) + ((g1479) & (!g1480) & (g1481) & (g1482) & (!g165) & (!g166)) + ((g1479) & (!g1480) & (g1481) & (g1482) & (!g165) & (g166)) + ((g1479) & (!g1480) & (g1481) & (g1482) & (g165) & (g166)) + ((g1479) & (g1480) & (!g1481) & (!g1482) & (!g165) & (!g166)) + ((g1479) & (g1480) & (!g1481) & (!g1482) & (g165) & (!g166)) + ((g1479) & (g1480) & (!g1481) & (g1482) & (!g165) & (!g166)) + ((g1479) & (g1480) & (!g1481) & (g1482) & (g165) & (!g166)) + ((g1479) & (g1480) & (!g1481) & (g1482) & (g165) & (g166)) + ((g1479) & (g1480) & (g1481) & (!g1482) & (!g165) & (!g166)) + ((g1479) & (g1480) & (g1481) & (!g1482) & (!g165) & (g166)) + ((g1479) & (g1480) & (g1481) & (!g1482) & (g165) & (!g166)) + ((g1479) & (g1480) & (g1481) & (g1482) & (!g165) & (!g166)) + ((g1479) & (g1480) & (g1481) & (g1482) & (!g165) & (g166)) + ((g1479) & (g1480) & (g1481) & (g1482) & (g165) & (!g166)) + ((g1479) & (g1480) & (g1481) & (g1482) & (g165) & (g166)));
	assign g4942 = (((!g2177) & (!g2805) & (!sk[14]) & (g1484)) + ((!g2177) & (!g2805) & (sk[14]) & (g1484)) + ((!g2177) & (g2805) & (!sk[14]) & (!g1484)) + ((!g2177) & (g2805) & (!sk[14]) & (g1484)) + ((!g2177) & (g2805) & (sk[14]) & (g1484)) + ((g2177) & (!g2805) & (!sk[14]) & (g1484)) + ((g2177) & (g2805) & (!sk[14]) & (!g1484)) + ((g2177) & (g2805) & (!sk[14]) & (g1484)) + ((g2177) & (g2805) & (sk[14]) & (!g1484)) + ((g2177) & (g2805) & (sk[14]) & (g1484)));
	assign g4943 = (((!g2178) & (!g2805) & (!sk[15]) & (g1485)) + ((!g2178) & (!g2805) & (sk[15]) & (g1485)) + ((!g2178) & (g2805) & (!sk[15]) & (!g1485)) + ((!g2178) & (g2805) & (!sk[15]) & (g1485)) + ((!g2178) & (g2805) & (sk[15]) & (g1485)) + ((g2178) & (!g2805) & (!sk[15]) & (g1485)) + ((g2178) & (g2805) & (!sk[15]) & (!g1485)) + ((g2178) & (g2805) & (!sk[15]) & (g1485)) + ((g2178) & (g2805) & (sk[15]) & (!g1485)) + ((g2178) & (g2805) & (sk[15]) & (g1485)));
	assign g4944 = (((!g2179) & (!sk[16]) & (!g2805) & (g1486)) + ((!g2179) & (!sk[16]) & (g2805) & (!g1486)) + ((!g2179) & (!sk[16]) & (g2805) & (g1486)) + ((!g2179) & (sk[16]) & (!g2805) & (g1486)) + ((!g2179) & (sk[16]) & (g2805) & (g1486)) + ((g2179) & (!sk[16]) & (!g2805) & (g1486)) + ((g2179) & (!sk[16]) & (g2805) & (!g1486)) + ((g2179) & (!sk[16]) & (g2805) & (g1486)) + ((g2179) & (sk[16]) & (g2805) & (!g1486)) + ((g2179) & (sk[16]) & (g2805) & (g1486)));
	assign g1487 = (((!g165) & (!sk[17]) & (!g166) & (!g1484) & (g1485) & (!g1486)) + ((!g165) & (!sk[17]) & (!g166) & (!g1484) & (g1485) & (g1486)) + ((!g165) & (!sk[17]) & (!g166) & (g1484) & (!g1485) & (!g1486)) + ((!g165) & (!sk[17]) & (!g166) & (g1484) & (!g1485) & (g1486)) + ((!g165) & (!sk[17]) & (!g166) & (g1484) & (g1485) & (!g1486)) + ((!g165) & (!sk[17]) & (!g166) & (g1484) & (g1485) & (g1486)) + ((!g165) & (!sk[17]) & (g166) & (!g1484) & (!g1485) & (!g1486)) + ((!g165) & (!sk[17]) & (g166) & (!g1484) & (!g1485) & (g1486)) + ((!g165) & (!sk[17]) & (g166) & (!g1484) & (g1485) & (!g1486)) + ((!g165) & (!sk[17]) & (g166) & (!g1484) & (g1485) & (g1486)) + ((!g165) & (!sk[17]) & (g166) & (g1484) & (!g1485) & (!g1486)) + ((!g165) & (!sk[17]) & (g166) & (g1484) & (!g1485) & (g1486)) + ((!g165) & (!sk[17]) & (g166) & (g1484) & (g1485) & (!g1486)) + ((!g165) & (!sk[17]) & (g166) & (g1484) & (g1485) & (g1486)) + ((!g165) & (sk[17]) & (g166) & (!g1484) & (!g1485) & (g1486)) + ((!g165) & (sk[17]) & (g166) & (!g1484) & (g1485) & (g1486)) + ((!g165) & (sk[17]) & (g166) & (g1484) & (!g1485) & (g1486)) + ((!g165) & (sk[17]) & (g166) & (g1484) & (g1485) & (g1486)) + ((g165) & (!sk[17]) & (!g166) & (!g1484) & (g1485) & (!g1486)) + ((g165) & (!sk[17]) & (!g166) & (!g1484) & (g1485) & (g1486)) + ((g165) & (!sk[17]) & (!g166) & (g1484) & (!g1485) & (!g1486)) + ((g165) & (!sk[17]) & (!g166) & (g1484) & (!g1485) & (g1486)) + ((g165) & (!sk[17]) & (!g166) & (g1484) & (g1485) & (!g1486)) + ((g165) & (!sk[17]) & (!g166) & (g1484) & (g1485) & (g1486)) + ((g165) & (!sk[17]) & (g166) & (!g1484) & (!g1485) & (!g1486)) + ((g165) & (!sk[17]) & (g166) & (!g1484) & (!g1485) & (g1486)) + ((g165) & (!sk[17]) & (g166) & (!g1484) & (g1485) & (!g1486)) + ((g165) & (!sk[17]) & (g166) & (!g1484) & (g1485) & (g1486)) + ((g165) & (!sk[17]) & (g166) & (g1484) & (!g1485) & (!g1486)) + ((g165) & (!sk[17]) & (g166) & (g1484) & (!g1485) & (g1486)) + ((g165) & (!sk[17]) & (g166) & (g1484) & (g1485) & (!g1486)) + ((g165) & (!sk[17]) & (g166) & (g1484) & (g1485) & (g1486)) + ((g165) & (sk[17]) & (!g166) & (g1484) & (!g1485) & (!g1486)) + ((g165) & (sk[17]) & (!g166) & (g1484) & (!g1485) & (g1486)) + ((g165) & (sk[17]) & (!g166) & (g1484) & (g1485) & (!g1486)) + ((g165) & (sk[17]) & (!g166) & (g1484) & (g1485) & (g1486)) + ((g165) & (sk[17]) & (g166) & (!g1484) & (g1485) & (!g1486)) + ((g165) & (sk[17]) & (g166) & (!g1484) & (g1485) & (g1486)) + ((g165) & (sk[17]) & (g166) & (g1484) & (g1485) & (!g1486)) + ((g165) & (sk[17]) & (g166) & (g1484) & (g1485) & (g1486)));
	assign g4945 = (((!sk[18]) & (!g2162) & (!g2805) & (g1488)) + ((!sk[18]) & (!g2162) & (g2805) & (!g1488)) + ((!sk[18]) & (!g2162) & (g2805) & (g1488)) + ((!sk[18]) & (g2162) & (!g2805) & (g1488)) + ((!sk[18]) & (g2162) & (g2805) & (!g1488)) + ((!sk[18]) & (g2162) & (g2805) & (g1488)) + ((sk[18]) & (!g2162) & (!g2805) & (g1488)) + ((sk[18]) & (!g2162) & (g2805) & (g1488)) + ((sk[18]) & (g2162) & (g2805) & (!g1488)) + ((sk[18]) & (g2162) & (g2805) & (g1488)));
	assign g4946 = (((!sk[19]) & (!g2164) & (!g2805) & (g1489)) + ((!sk[19]) & (!g2164) & (g2805) & (!g1489)) + ((!sk[19]) & (!g2164) & (g2805) & (g1489)) + ((!sk[19]) & (g2164) & (!g2805) & (g1489)) + ((!sk[19]) & (g2164) & (g2805) & (!g1489)) + ((!sk[19]) & (g2164) & (g2805) & (g1489)) + ((sk[19]) & (!g2164) & (!g2805) & (g1489)) + ((sk[19]) & (!g2164) & (g2805) & (g1489)) + ((sk[19]) & (g2164) & (g2805) & (!g1489)) + ((sk[19]) & (g2164) & (g2805) & (g1489)));
	assign g4947 = (((!g2166) & (!g2805) & (!sk[20]) & (g1490)) + ((!g2166) & (!g2805) & (sk[20]) & (g1490)) + ((!g2166) & (g2805) & (!sk[20]) & (!g1490)) + ((!g2166) & (g2805) & (!sk[20]) & (g1490)) + ((!g2166) & (g2805) & (sk[20]) & (g1490)) + ((g2166) & (!g2805) & (!sk[20]) & (g1490)) + ((g2166) & (g2805) & (!sk[20]) & (!g1490)) + ((g2166) & (g2805) & (!sk[20]) & (g1490)) + ((g2166) & (g2805) & (sk[20]) & (!g1490)) + ((g2166) & (g2805) & (sk[20]) & (g1490)));
	assign g4948 = (((!g2168) & (!sk[21]) & (!g2805) & (g1491)) + ((!g2168) & (!sk[21]) & (g2805) & (!g1491)) + ((!g2168) & (!sk[21]) & (g2805) & (g1491)) + ((!g2168) & (sk[21]) & (!g2805) & (g1491)) + ((!g2168) & (sk[21]) & (g2805) & (g1491)) + ((g2168) & (!sk[21]) & (!g2805) & (g1491)) + ((g2168) & (!sk[21]) & (g2805) & (!g1491)) + ((g2168) & (!sk[21]) & (g2805) & (g1491)) + ((g2168) & (sk[21]) & (g2805) & (!g1491)) + ((g2168) & (sk[21]) & (g2805) & (g1491)));
	assign g1492 = (((!g1488) & (!g1489) & (!g1490) & (g1491) & (g165) & (g166)) + ((!g1488) & (!g1489) & (g1490) & (!g1491) & (!g165) & (g166)) + ((!g1488) & (!g1489) & (g1490) & (g1491) & (!g165) & (g166)) + ((!g1488) & (!g1489) & (g1490) & (g1491) & (g165) & (g166)) + ((!g1488) & (g1489) & (!g1490) & (!g1491) & (g165) & (!g166)) + ((!g1488) & (g1489) & (!g1490) & (g1491) & (g165) & (!g166)) + ((!g1488) & (g1489) & (!g1490) & (g1491) & (g165) & (g166)) + ((!g1488) & (g1489) & (g1490) & (!g1491) & (!g165) & (g166)) + ((!g1488) & (g1489) & (g1490) & (!g1491) & (g165) & (!g166)) + ((!g1488) & (g1489) & (g1490) & (g1491) & (!g165) & (g166)) + ((!g1488) & (g1489) & (g1490) & (g1491) & (g165) & (!g166)) + ((!g1488) & (g1489) & (g1490) & (g1491) & (g165) & (g166)) + ((g1488) & (!g1489) & (!g1490) & (!g1491) & (!g165) & (!g166)) + ((g1488) & (!g1489) & (!g1490) & (g1491) & (!g165) & (!g166)) + ((g1488) & (!g1489) & (!g1490) & (g1491) & (g165) & (g166)) + ((g1488) & (!g1489) & (g1490) & (!g1491) & (!g165) & (!g166)) + ((g1488) & (!g1489) & (g1490) & (!g1491) & (!g165) & (g166)) + ((g1488) & (!g1489) & (g1490) & (g1491) & (!g165) & (!g166)) + ((g1488) & (!g1489) & (g1490) & (g1491) & (!g165) & (g166)) + ((g1488) & (!g1489) & (g1490) & (g1491) & (g165) & (g166)) + ((g1488) & (g1489) & (!g1490) & (!g1491) & (!g165) & (!g166)) + ((g1488) & (g1489) & (!g1490) & (!g1491) & (g165) & (!g166)) + ((g1488) & (g1489) & (!g1490) & (g1491) & (!g165) & (!g166)) + ((g1488) & (g1489) & (!g1490) & (g1491) & (g165) & (!g166)) + ((g1488) & (g1489) & (!g1490) & (g1491) & (g165) & (g166)) + ((g1488) & (g1489) & (g1490) & (!g1491) & (!g165) & (!g166)) + ((g1488) & (g1489) & (g1490) & (!g1491) & (!g165) & (g166)) + ((g1488) & (g1489) & (g1490) & (!g1491) & (g165) & (!g166)) + ((g1488) & (g1489) & (g1490) & (g1491) & (!g165) & (!g166)) + ((g1488) & (g1489) & (g1490) & (g1491) & (!g165) & (g166)) + ((g1488) & (g1489) & (g1490) & (g1491) & (g165) & (!g166)) + ((g1488) & (g1489) & (g1490) & (g1491) & (g165) & (g166)));
	assign g4949 = (((!g2169) & (!g2805) & (!sk[23]) & (g1493)) + ((!g2169) & (!g2805) & (sk[23]) & (g1493)) + ((!g2169) & (g2805) & (!sk[23]) & (!g1493)) + ((!g2169) & (g2805) & (!sk[23]) & (g1493)) + ((!g2169) & (g2805) & (sk[23]) & (g1493)) + ((g2169) & (!g2805) & (!sk[23]) & (g1493)) + ((g2169) & (g2805) & (!sk[23]) & (!g1493)) + ((g2169) & (g2805) & (!sk[23]) & (g1493)) + ((g2169) & (g2805) & (sk[23]) & (!g1493)) + ((g2169) & (g2805) & (sk[23]) & (g1493)));
	assign g4950 = (((!g2170) & (!g2805) & (!sk[24]) & (g1494)) + ((!g2170) & (!g2805) & (sk[24]) & (g1494)) + ((!g2170) & (g2805) & (!sk[24]) & (!g1494)) + ((!g2170) & (g2805) & (!sk[24]) & (g1494)) + ((!g2170) & (g2805) & (sk[24]) & (g1494)) + ((g2170) & (!g2805) & (!sk[24]) & (g1494)) + ((g2170) & (g2805) & (!sk[24]) & (!g1494)) + ((g2170) & (g2805) & (!sk[24]) & (g1494)) + ((g2170) & (g2805) & (sk[24]) & (!g1494)) + ((g2170) & (g2805) & (sk[24]) & (g1494)));
	assign g4951 = (((!g2171) & (!g2805) & (!sk[25]) & (g1495)) + ((!g2171) & (!g2805) & (sk[25]) & (g1495)) + ((!g2171) & (g2805) & (!sk[25]) & (!g1495)) + ((!g2171) & (g2805) & (!sk[25]) & (g1495)) + ((!g2171) & (g2805) & (sk[25]) & (g1495)) + ((g2171) & (!g2805) & (!sk[25]) & (g1495)) + ((g2171) & (g2805) & (!sk[25]) & (!g1495)) + ((g2171) & (g2805) & (!sk[25]) & (g1495)) + ((g2171) & (g2805) & (sk[25]) & (!g1495)) + ((g2171) & (g2805) & (sk[25]) & (g1495)));
	assign g4952 = (((!sk[26]) & (!g2172) & (!g2805) & (g1496)) + ((!sk[26]) & (!g2172) & (g2805) & (!g1496)) + ((!sk[26]) & (!g2172) & (g2805) & (g1496)) + ((!sk[26]) & (g2172) & (!g2805) & (g1496)) + ((!sk[26]) & (g2172) & (g2805) & (!g1496)) + ((!sk[26]) & (g2172) & (g2805) & (g1496)) + ((sk[26]) & (!g2172) & (!g2805) & (g1496)) + ((sk[26]) & (!g2172) & (g2805) & (g1496)) + ((sk[26]) & (g2172) & (g2805) & (!g1496)) + ((sk[26]) & (g2172) & (g2805) & (g1496)));
	assign g1497 = (((!g1493) & (!g1494) & (!g1495) & (g1496) & (g165) & (g166)) + ((!g1493) & (!g1494) & (g1495) & (!g1496) & (!g165) & (g166)) + ((!g1493) & (!g1494) & (g1495) & (g1496) & (!g165) & (g166)) + ((!g1493) & (!g1494) & (g1495) & (g1496) & (g165) & (g166)) + ((!g1493) & (g1494) & (!g1495) & (!g1496) & (g165) & (!g166)) + ((!g1493) & (g1494) & (!g1495) & (g1496) & (g165) & (!g166)) + ((!g1493) & (g1494) & (!g1495) & (g1496) & (g165) & (g166)) + ((!g1493) & (g1494) & (g1495) & (!g1496) & (!g165) & (g166)) + ((!g1493) & (g1494) & (g1495) & (!g1496) & (g165) & (!g166)) + ((!g1493) & (g1494) & (g1495) & (g1496) & (!g165) & (g166)) + ((!g1493) & (g1494) & (g1495) & (g1496) & (g165) & (!g166)) + ((!g1493) & (g1494) & (g1495) & (g1496) & (g165) & (g166)) + ((g1493) & (!g1494) & (!g1495) & (!g1496) & (!g165) & (!g166)) + ((g1493) & (!g1494) & (!g1495) & (g1496) & (!g165) & (!g166)) + ((g1493) & (!g1494) & (!g1495) & (g1496) & (g165) & (g166)) + ((g1493) & (!g1494) & (g1495) & (!g1496) & (!g165) & (!g166)) + ((g1493) & (!g1494) & (g1495) & (!g1496) & (!g165) & (g166)) + ((g1493) & (!g1494) & (g1495) & (g1496) & (!g165) & (!g166)) + ((g1493) & (!g1494) & (g1495) & (g1496) & (!g165) & (g166)) + ((g1493) & (!g1494) & (g1495) & (g1496) & (g165) & (g166)) + ((g1493) & (g1494) & (!g1495) & (!g1496) & (!g165) & (!g166)) + ((g1493) & (g1494) & (!g1495) & (!g1496) & (g165) & (!g166)) + ((g1493) & (g1494) & (!g1495) & (g1496) & (!g165) & (!g166)) + ((g1493) & (g1494) & (!g1495) & (g1496) & (g165) & (!g166)) + ((g1493) & (g1494) & (!g1495) & (g1496) & (g165) & (g166)) + ((g1493) & (g1494) & (g1495) & (!g1496) & (!g165) & (!g166)) + ((g1493) & (g1494) & (g1495) & (!g1496) & (!g165) & (g166)) + ((g1493) & (g1494) & (g1495) & (!g1496) & (g165) & (!g166)) + ((g1493) & (g1494) & (g1495) & (g1496) & (!g165) & (!g166)) + ((g1493) & (g1494) & (g1495) & (g1496) & (!g165) & (g166)) + ((g1493) & (g1494) & (g1495) & (g1496) & (g165) & (!g166)) + ((g1493) & (g1494) & (g1495) & (g1496) & (g165) & (g166)));
	assign g1498 = (((!g147) & (!g148) & (!g1483) & (g1487) & (!g1492) & (!g1497)) + ((!g147) & (!g148) & (!g1483) & (g1487) & (!g1492) & (g1497)) + ((!g147) & (!g148) & (!g1483) & (g1487) & (g1492) & (!g1497)) + ((!g147) & (!g148) & (!g1483) & (g1487) & (g1492) & (g1497)) + ((!g147) & (!g148) & (g1483) & (g1487) & (!g1492) & (!g1497)) + ((!g147) & (!g148) & (g1483) & (g1487) & (!g1492) & (g1497)) + ((!g147) & (!g148) & (g1483) & (g1487) & (g1492) & (!g1497)) + ((!g147) & (!g148) & (g1483) & (g1487) & (g1492) & (g1497)) + ((!g147) & (g148) & (!g1483) & (!g1487) & (!g1492) & (g1497)) + ((!g147) & (g148) & (!g1483) & (!g1487) & (g1492) & (g1497)) + ((!g147) & (g148) & (!g1483) & (g1487) & (!g1492) & (g1497)) + ((!g147) & (g148) & (!g1483) & (g1487) & (g1492) & (g1497)) + ((!g147) & (g148) & (g1483) & (!g1487) & (!g1492) & (g1497)) + ((!g147) & (g148) & (g1483) & (!g1487) & (g1492) & (g1497)) + ((!g147) & (g148) & (g1483) & (g1487) & (!g1492) & (g1497)) + ((!g147) & (g148) & (g1483) & (g1487) & (g1492) & (g1497)) + ((g147) & (!g148) & (g1483) & (!g1487) & (!g1492) & (!g1497)) + ((g147) & (!g148) & (g1483) & (!g1487) & (!g1492) & (g1497)) + ((g147) & (!g148) & (g1483) & (!g1487) & (g1492) & (!g1497)) + ((g147) & (!g148) & (g1483) & (!g1487) & (g1492) & (g1497)) + ((g147) & (!g148) & (g1483) & (g1487) & (!g1492) & (!g1497)) + ((g147) & (!g148) & (g1483) & (g1487) & (!g1492) & (g1497)) + ((g147) & (!g148) & (g1483) & (g1487) & (g1492) & (!g1497)) + ((g147) & (!g148) & (g1483) & (g1487) & (g1492) & (g1497)) + ((g147) & (g148) & (!g1483) & (!g1487) & (g1492) & (!g1497)) + ((g147) & (g148) & (!g1483) & (!g1487) & (g1492) & (g1497)) + ((g147) & (g148) & (!g1483) & (g1487) & (g1492) & (!g1497)) + ((g147) & (g148) & (!g1483) & (g1487) & (g1492) & (g1497)) + ((g147) & (g148) & (g1483) & (!g1487) & (g1492) & (!g1497)) + ((g147) & (g148) & (g1483) & (!g1487) & (g1492) & (g1497)) + ((g147) & (g148) & (g1483) & (g1487) & (g1492) & (!g1497)) + ((g147) & (g148) & (g1483) & (g1487) & (g1492) & (g1497)));
	assign g1499 = (((!g142) & (!sk[29]) & (!g1478) & (g1498)) + ((!g142) & (!sk[29]) & (g1478) & (!g1498)) + ((!g142) & (!sk[29]) & (g1478) & (g1498)) + ((!g142) & (sk[29]) & (!g1478) & (g1498)) + ((!g142) & (sk[29]) & (g1478) & (g1498)) + ((g142) & (!sk[29]) & (!g1478) & (g1498)) + ((g142) & (!sk[29]) & (g1478) & (!g1498)) + ((g142) & (!sk[29]) & (g1478) & (g1498)) + ((g142) & (sk[29]) & (g1478) & (!g1498)) + ((g142) & (sk[29]) & (g1478) & (g1498)));
	assign g4953 = (((!g2059) & (!g2810) & (!sk[30]) & (g1500)) + ((!g2059) & (!g2810) & (sk[30]) & (g1500)) + ((!g2059) & (g2810) & (!sk[30]) & (!g1500)) + ((!g2059) & (g2810) & (!sk[30]) & (g1500)) + ((!g2059) & (g2810) & (sk[30]) & (g1500)) + ((g2059) & (!g2810) & (!sk[30]) & (g1500)) + ((g2059) & (g2810) & (!sk[30]) & (!g1500)) + ((g2059) & (g2810) & (!sk[30]) & (g1500)) + ((g2059) & (g2810) & (sk[30]) & (!g1500)) + ((g2059) & (g2810) & (sk[30]) & (g1500)));
	assign g1501 = (((!g126) & (!g1499) & (!g916) & (!g1456) & (sk[31]) & (g3118)) + ((!g126) & (!g1499) & (!g916) & (g1456) & (!sk[31]) & (!g3118)) + ((!g126) & (!g1499) & (!g916) & (g1456) & (!sk[31]) & (g3118)) + ((!g126) & (!g1499) & (!g916) & (g1456) & (sk[31]) & (g3118)) + ((!g126) & (!g1499) & (g916) & (!g1456) & (!sk[31]) & (!g3118)) + ((!g126) & (!g1499) & (g916) & (!g1456) & (!sk[31]) & (g3118)) + ((!g126) & (!g1499) & (g916) & (!g1456) & (sk[31]) & (g3118)) + ((!g126) & (!g1499) & (g916) & (g1456) & (!sk[31]) & (!g3118)) + ((!g126) & (!g1499) & (g916) & (g1456) & (!sk[31]) & (g3118)) + ((!g126) & (!g1499) & (g916) & (g1456) & (sk[31]) & (g3118)) + ((!g126) & (g1499) & (!g916) & (!g1456) & (!sk[31]) & (!g3118)) + ((!g126) & (g1499) & (!g916) & (!g1456) & (!sk[31]) & (g3118)) + ((!g126) & (g1499) & (!g916) & (!g1456) & (sk[31]) & (g3118)) + ((!g126) & (g1499) & (!g916) & (g1456) & (!sk[31]) & (!g3118)) + ((!g126) & (g1499) & (!g916) & (g1456) & (!sk[31]) & (g3118)) + ((!g126) & (g1499) & (!g916) & (g1456) & (sk[31]) & (g3118)) + ((!g126) & (g1499) & (g916) & (!g1456) & (!sk[31]) & (!g3118)) + ((!g126) & (g1499) & (g916) & (!g1456) & (!sk[31]) & (g3118)) + ((!g126) & (g1499) & (g916) & (!g1456) & (sk[31]) & (g3118)) + ((!g126) & (g1499) & (g916) & (g1456) & (!sk[31]) & (!g3118)) + ((!g126) & (g1499) & (g916) & (g1456) & (!sk[31]) & (g3118)) + ((!g126) & (g1499) & (g916) & (g1456) & (sk[31]) & (g3118)) + ((g126) & (!g1499) & (!g916) & (g1456) & (!sk[31]) & (!g3118)) + ((g126) & (!g1499) & (!g916) & (g1456) & (!sk[31]) & (g3118)) + ((g126) & (!g1499) & (!g916) & (g1456) & (sk[31]) & (g3118)) + ((g126) & (!g1499) & (g916) & (!g1456) & (!sk[31]) & (!g3118)) + ((g126) & (!g1499) & (g916) & (!g1456) & (!sk[31]) & (g3118)) + ((g126) & (!g1499) & (g916) & (!g1456) & (sk[31]) & (!g3118)) + ((g126) & (!g1499) & (g916) & (g1456) & (!sk[31]) & (!g3118)) + ((g126) & (!g1499) & (g916) & (g1456) & (!sk[31]) & (g3118)) + ((g126) & (g1499) & (!g916) & (!g1456) & (!sk[31]) & (!g3118)) + ((g126) & (g1499) & (!g916) & (!g1456) & (!sk[31]) & (g3118)) + ((g126) & (g1499) & (!g916) & (!g1456) & (sk[31]) & (!g3118)) + ((g126) & (g1499) & (!g916) & (!g1456) & (sk[31]) & (g3118)) + ((g126) & (g1499) & (!g916) & (g1456) & (!sk[31]) & (!g3118)) + ((g126) & (g1499) & (!g916) & (g1456) & (!sk[31]) & (g3118)) + ((g126) & (g1499) & (!g916) & (g1456) & (sk[31]) & (!g3118)) + ((g126) & (g1499) & (g916) & (!g1456) & (!sk[31]) & (!g3118)) + ((g126) & (g1499) & (g916) & (!g1456) & (!sk[31]) & (g3118)) + ((g126) & (g1499) & (g916) & (!g1456) & (sk[31]) & (g3118)) + ((g126) & (g1499) & (g916) & (g1456) & (!sk[31]) & (!g3118)) + ((g126) & (g1499) & (g916) & (g1456) & (!sk[31]) & (g3118)) + ((g126) & (g1499) & (g916) & (g1456) & (sk[31]) & (!g3118)) + ((g126) & (g1499) & (g916) & (g1456) & (sk[31]) & (g3118)));
	assign g4954 = (((!g2140) & (!sk[32]) & (!g2821) & (g1502)) + ((!g2140) & (!sk[32]) & (g2821) & (!g1502)) + ((!g2140) & (!sk[32]) & (g2821) & (g1502)) + ((!g2140) & (sk[32]) & (!g2821) & (g1502)) + ((!g2140) & (sk[32]) & (g2821) & (g1502)) + ((g2140) & (!sk[32]) & (!g2821) & (g1502)) + ((g2140) & (!sk[32]) & (g2821) & (!g1502)) + ((g2140) & (!sk[32]) & (g2821) & (g1502)) + ((g2140) & (sk[32]) & (g2821) & (!g1502)) + ((g2140) & (sk[32]) & (g2821) & (g1502)));
	assign g4955 = (((!g2142) & (!sk[33]) & (!g2821) & (g1503)) + ((!g2142) & (!sk[33]) & (g2821) & (!g1503)) + ((!g2142) & (!sk[33]) & (g2821) & (g1503)) + ((!g2142) & (sk[33]) & (!g2821) & (g1503)) + ((!g2142) & (sk[33]) & (g2821) & (g1503)) + ((g2142) & (!sk[33]) & (!g2821) & (g1503)) + ((g2142) & (!sk[33]) & (g2821) & (!g1503)) + ((g2142) & (!sk[33]) & (g2821) & (g1503)) + ((g2142) & (sk[33]) & (g2821) & (!g1503)) + ((g2142) & (sk[33]) & (g2821) & (g1503)));
	assign g4956 = (((!g2144) & (!sk[34]) & (!g2821) & (g1504)) + ((!g2144) & (!sk[34]) & (g2821) & (!g1504)) + ((!g2144) & (!sk[34]) & (g2821) & (g1504)) + ((!g2144) & (sk[34]) & (!g2821) & (g1504)) + ((!g2144) & (sk[34]) & (g2821) & (g1504)) + ((g2144) & (!sk[34]) & (!g2821) & (g1504)) + ((g2144) & (!sk[34]) & (g2821) & (!g1504)) + ((g2144) & (!sk[34]) & (g2821) & (g1504)) + ((g2144) & (sk[34]) & (g2821) & (!g1504)) + ((g2144) & (sk[34]) & (g2821) & (g1504)));
	assign g4957 = (((!sk[35]) & (!g2145) & (!g2821) & (g1505)) + ((!sk[35]) & (!g2145) & (g2821) & (!g1505)) + ((!sk[35]) & (!g2145) & (g2821) & (g1505)) + ((!sk[35]) & (g2145) & (!g2821) & (g1505)) + ((!sk[35]) & (g2145) & (g2821) & (!g1505)) + ((!sk[35]) & (g2145) & (g2821) & (g1505)) + ((sk[35]) & (!g2145) & (!g2821) & (g1505)) + ((sk[35]) & (!g2145) & (g2821) & (g1505)) + ((sk[35]) & (g2145) & (g2821) & (!g1505)) + ((sk[35]) & (g2145) & (g2821) & (g1505)));
	assign g1506 = (((!g1502) & (!g1503) & (!g1504) & (g1505) & (g147) & (g148)) + ((!g1502) & (!g1503) & (g1504) & (!g1505) & (!g147) & (g148)) + ((!g1502) & (!g1503) & (g1504) & (g1505) & (!g147) & (g148)) + ((!g1502) & (!g1503) & (g1504) & (g1505) & (g147) & (g148)) + ((!g1502) & (g1503) & (!g1504) & (!g1505) & (g147) & (!g148)) + ((!g1502) & (g1503) & (!g1504) & (g1505) & (g147) & (!g148)) + ((!g1502) & (g1503) & (!g1504) & (g1505) & (g147) & (g148)) + ((!g1502) & (g1503) & (g1504) & (!g1505) & (!g147) & (g148)) + ((!g1502) & (g1503) & (g1504) & (!g1505) & (g147) & (!g148)) + ((!g1502) & (g1503) & (g1504) & (g1505) & (!g147) & (g148)) + ((!g1502) & (g1503) & (g1504) & (g1505) & (g147) & (!g148)) + ((!g1502) & (g1503) & (g1504) & (g1505) & (g147) & (g148)) + ((g1502) & (!g1503) & (!g1504) & (!g1505) & (!g147) & (!g148)) + ((g1502) & (!g1503) & (!g1504) & (g1505) & (!g147) & (!g148)) + ((g1502) & (!g1503) & (!g1504) & (g1505) & (g147) & (g148)) + ((g1502) & (!g1503) & (g1504) & (!g1505) & (!g147) & (!g148)) + ((g1502) & (!g1503) & (g1504) & (!g1505) & (!g147) & (g148)) + ((g1502) & (!g1503) & (g1504) & (g1505) & (!g147) & (!g148)) + ((g1502) & (!g1503) & (g1504) & (g1505) & (!g147) & (g148)) + ((g1502) & (!g1503) & (g1504) & (g1505) & (g147) & (g148)) + ((g1502) & (g1503) & (!g1504) & (!g1505) & (!g147) & (!g148)) + ((g1502) & (g1503) & (!g1504) & (!g1505) & (g147) & (!g148)) + ((g1502) & (g1503) & (!g1504) & (g1505) & (!g147) & (!g148)) + ((g1502) & (g1503) & (!g1504) & (g1505) & (g147) & (!g148)) + ((g1502) & (g1503) & (!g1504) & (g1505) & (g147) & (g148)) + ((g1502) & (g1503) & (g1504) & (!g1505) & (!g147) & (!g148)) + ((g1502) & (g1503) & (g1504) & (!g1505) & (!g147) & (g148)) + ((g1502) & (g1503) & (g1504) & (!g1505) & (g147) & (!g148)) + ((g1502) & (g1503) & (g1504) & (g1505) & (!g147) & (!g148)) + ((g1502) & (g1503) & (g1504) & (g1505) & (!g147) & (g148)) + ((g1502) & (g1503) & (g1504) & (g1505) & (g147) & (!g148)) + ((g1502) & (g1503) & (g1504) & (g1505) & (g147) & (g148)));
	assign g4958 = (((!sk[37]) & (!g2146) & (!g2821) & (g1507)) + ((!sk[37]) & (!g2146) & (g2821) & (!g1507)) + ((!sk[37]) & (!g2146) & (g2821) & (g1507)) + ((!sk[37]) & (g2146) & (!g2821) & (g1507)) + ((!sk[37]) & (g2146) & (g2821) & (!g1507)) + ((!sk[37]) & (g2146) & (g2821) & (g1507)) + ((sk[37]) & (!g2146) & (!g2821) & (g1507)) + ((sk[37]) & (!g2146) & (g2821) & (g1507)) + ((sk[37]) & (g2146) & (g2821) & (!g1507)) + ((sk[37]) & (g2146) & (g2821) & (g1507)));
	assign g4959 = (((!g2148) & (!g2821) & (!sk[38]) & (g1508)) + ((!g2148) & (!g2821) & (sk[38]) & (g1508)) + ((!g2148) & (g2821) & (!sk[38]) & (!g1508)) + ((!g2148) & (g2821) & (!sk[38]) & (g1508)) + ((!g2148) & (g2821) & (sk[38]) & (g1508)) + ((g2148) & (!g2821) & (!sk[38]) & (g1508)) + ((g2148) & (g2821) & (!sk[38]) & (!g1508)) + ((g2148) & (g2821) & (!sk[38]) & (g1508)) + ((g2148) & (g2821) & (sk[38]) & (!g1508)) + ((g2148) & (g2821) & (sk[38]) & (g1508)));
	assign g4960 = (((!g2150) & (!g2821) & (!sk[39]) & (g1509)) + ((!g2150) & (!g2821) & (sk[39]) & (g1509)) + ((!g2150) & (g2821) & (!sk[39]) & (!g1509)) + ((!g2150) & (g2821) & (!sk[39]) & (g1509)) + ((!g2150) & (g2821) & (sk[39]) & (g1509)) + ((g2150) & (!g2821) & (!sk[39]) & (g1509)) + ((g2150) & (g2821) & (!sk[39]) & (!g1509)) + ((g2150) & (g2821) & (!sk[39]) & (g1509)) + ((g2150) & (g2821) & (sk[39]) & (!g1509)) + ((g2150) & (g2821) & (sk[39]) & (g1509)));
	assign g4961 = (((!g2151) & (!g2821) & (!sk[40]) & (g1510)) + ((!g2151) & (!g2821) & (sk[40]) & (g1510)) + ((!g2151) & (g2821) & (!sk[40]) & (!g1510)) + ((!g2151) & (g2821) & (!sk[40]) & (g1510)) + ((!g2151) & (g2821) & (sk[40]) & (g1510)) + ((g2151) & (!g2821) & (!sk[40]) & (g1510)) + ((g2151) & (g2821) & (!sk[40]) & (!g1510)) + ((g2151) & (g2821) & (!sk[40]) & (g1510)) + ((g2151) & (g2821) & (sk[40]) & (!g1510)) + ((g2151) & (g2821) & (sk[40]) & (g1510)));
	assign g1511 = (((!g1507) & (!g1508) & (!g1509) & (g1510) & (g147) & (g148)) + ((!g1507) & (!g1508) & (g1509) & (!g1510) & (!g147) & (g148)) + ((!g1507) & (!g1508) & (g1509) & (g1510) & (!g147) & (g148)) + ((!g1507) & (!g1508) & (g1509) & (g1510) & (g147) & (g148)) + ((!g1507) & (g1508) & (!g1509) & (!g1510) & (g147) & (!g148)) + ((!g1507) & (g1508) & (!g1509) & (g1510) & (g147) & (!g148)) + ((!g1507) & (g1508) & (!g1509) & (g1510) & (g147) & (g148)) + ((!g1507) & (g1508) & (g1509) & (!g1510) & (!g147) & (g148)) + ((!g1507) & (g1508) & (g1509) & (!g1510) & (g147) & (!g148)) + ((!g1507) & (g1508) & (g1509) & (g1510) & (!g147) & (g148)) + ((!g1507) & (g1508) & (g1509) & (g1510) & (g147) & (!g148)) + ((!g1507) & (g1508) & (g1509) & (g1510) & (g147) & (g148)) + ((g1507) & (!g1508) & (!g1509) & (!g1510) & (!g147) & (!g148)) + ((g1507) & (!g1508) & (!g1509) & (g1510) & (!g147) & (!g148)) + ((g1507) & (!g1508) & (!g1509) & (g1510) & (g147) & (g148)) + ((g1507) & (!g1508) & (g1509) & (!g1510) & (!g147) & (!g148)) + ((g1507) & (!g1508) & (g1509) & (!g1510) & (!g147) & (g148)) + ((g1507) & (!g1508) & (g1509) & (g1510) & (!g147) & (!g148)) + ((g1507) & (!g1508) & (g1509) & (g1510) & (!g147) & (g148)) + ((g1507) & (!g1508) & (g1509) & (g1510) & (g147) & (g148)) + ((g1507) & (g1508) & (!g1509) & (!g1510) & (!g147) & (!g148)) + ((g1507) & (g1508) & (!g1509) & (!g1510) & (g147) & (!g148)) + ((g1507) & (g1508) & (!g1509) & (g1510) & (!g147) & (!g148)) + ((g1507) & (g1508) & (!g1509) & (g1510) & (g147) & (!g148)) + ((g1507) & (g1508) & (!g1509) & (g1510) & (g147) & (g148)) + ((g1507) & (g1508) & (g1509) & (!g1510) & (!g147) & (!g148)) + ((g1507) & (g1508) & (g1509) & (!g1510) & (!g147) & (g148)) + ((g1507) & (g1508) & (g1509) & (!g1510) & (g147) & (!g148)) + ((g1507) & (g1508) & (g1509) & (g1510) & (!g147) & (!g148)) + ((g1507) & (g1508) & (g1509) & (g1510) & (!g147) & (g148)) + ((g1507) & (g1508) & (g1509) & (g1510) & (g147) & (!g148)) + ((g1507) & (g1508) & (g1509) & (g1510) & (g147) & (g148)));
	assign g4962 = (((!g2152) & (!sk[42]) & (!g2821) & (g1512)) + ((!g2152) & (!sk[42]) & (g2821) & (!g1512)) + ((!g2152) & (!sk[42]) & (g2821) & (g1512)) + ((!g2152) & (sk[42]) & (!g2821) & (g1512)) + ((!g2152) & (sk[42]) & (g2821) & (g1512)) + ((g2152) & (!sk[42]) & (!g2821) & (g1512)) + ((g2152) & (!sk[42]) & (g2821) & (!g1512)) + ((g2152) & (!sk[42]) & (g2821) & (g1512)) + ((g2152) & (sk[42]) & (g2821) & (!g1512)) + ((g2152) & (sk[42]) & (g2821) & (g1512)));
	assign g4963 = (((!sk[43]) & (!g2153) & (!g2821) & (g1513)) + ((!sk[43]) & (!g2153) & (g2821) & (!g1513)) + ((!sk[43]) & (!g2153) & (g2821) & (g1513)) + ((!sk[43]) & (g2153) & (!g2821) & (g1513)) + ((!sk[43]) & (g2153) & (g2821) & (!g1513)) + ((!sk[43]) & (g2153) & (g2821) & (g1513)) + ((sk[43]) & (!g2153) & (!g2821) & (g1513)) + ((sk[43]) & (!g2153) & (g2821) & (g1513)) + ((sk[43]) & (g2153) & (g2821) & (!g1513)) + ((sk[43]) & (g2153) & (g2821) & (g1513)));
	assign g4964 = (((!g2155) & (!g2821) & (!sk[44]) & (g1514)) + ((!g2155) & (!g2821) & (sk[44]) & (g1514)) + ((!g2155) & (g2821) & (!sk[44]) & (!g1514)) + ((!g2155) & (g2821) & (!sk[44]) & (g1514)) + ((!g2155) & (g2821) & (sk[44]) & (g1514)) + ((g2155) & (!g2821) & (!sk[44]) & (g1514)) + ((g2155) & (g2821) & (!sk[44]) & (!g1514)) + ((g2155) & (g2821) & (!sk[44]) & (g1514)) + ((g2155) & (g2821) & (sk[44]) & (!g1514)) + ((g2155) & (g2821) & (sk[44]) & (g1514)));
	assign g4965 = (((!g2157) & (!g2821) & (!sk[45]) & (g1515)) + ((!g2157) & (!g2821) & (sk[45]) & (g1515)) + ((!g2157) & (g2821) & (!sk[45]) & (!g1515)) + ((!g2157) & (g2821) & (!sk[45]) & (g1515)) + ((!g2157) & (g2821) & (sk[45]) & (g1515)) + ((g2157) & (!g2821) & (!sk[45]) & (g1515)) + ((g2157) & (g2821) & (!sk[45]) & (!g1515)) + ((g2157) & (g2821) & (!sk[45]) & (g1515)) + ((g2157) & (g2821) & (sk[45]) & (!g1515)) + ((g2157) & (g2821) & (sk[45]) & (g1515)));
	assign g1516 = (((!g1512) & (!g1513) & (!g1514) & (g1515) & (g147) & (g148)) + ((!g1512) & (!g1513) & (g1514) & (!g1515) & (!g147) & (g148)) + ((!g1512) & (!g1513) & (g1514) & (g1515) & (!g147) & (g148)) + ((!g1512) & (!g1513) & (g1514) & (g1515) & (g147) & (g148)) + ((!g1512) & (g1513) & (!g1514) & (!g1515) & (g147) & (!g148)) + ((!g1512) & (g1513) & (!g1514) & (g1515) & (g147) & (!g148)) + ((!g1512) & (g1513) & (!g1514) & (g1515) & (g147) & (g148)) + ((!g1512) & (g1513) & (g1514) & (!g1515) & (!g147) & (g148)) + ((!g1512) & (g1513) & (g1514) & (!g1515) & (g147) & (!g148)) + ((!g1512) & (g1513) & (g1514) & (g1515) & (!g147) & (g148)) + ((!g1512) & (g1513) & (g1514) & (g1515) & (g147) & (!g148)) + ((!g1512) & (g1513) & (g1514) & (g1515) & (g147) & (g148)) + ((g1512) & (!g1513) & (!g1514) & (!g1515) & (!g147) & (!g148)) + ((g1512) & (!g1513) & (!g1514) & (g1515) & (!g147) & (!g148)) + ((g1512) & (!g1513) & (!g1514) & (g1515) & (g147) & (g148)) + ((g1512) & (!g1513) & (g1514) & (!g1515) & (!g147) & (!g148)) + ((g1512) & (!g1513) & (g1514) & (!g1515) & (!g147) & (g148)) + ((g1512) & (!g1513) & (g1514) & (g1515) & (!g147) & (!g148)) + ((g1512) & (!g1513) & (g1514) & (g1515) & (!g147) & (g148)) + ((g1512) & (!g1513) & (g1514) & (g1515) & (g147) & (g148)) + ((g1512) & (g1513) & (!g1514) & (!g1515) & (!g147) & (!g148)) + ((g1512) & (g1513) & (!g1514) & (!g1515) & (g147) & (!g148)) + ((g1512) & (g1513) & (!g1514) & (g1515) & (!g147) & (!g148)) + ((g1512) & (g1513) & (!g1514) & (g1515) & (g147) & (!g148)) + ((g1512) & (g1513) & (!g1514) & (g1515) & (g147) & (g148)) + ((g1512) & (g1513) & (g1514) & (!g1515) & (!g147) & (!g148)) + ((g1512) & (g1513) & (g1514) & (!g1515) & (!g147) & (g148)) + ((g1512) & (g1513) & (g1514) & (!g1515) & (g147) & (!g148)) + ((g1512) & (g1513) & (g1514) & (g1515) & (!g147) & (!g148)) + ((g1512) & (g1513) & (g1514) & (g1515) & (!g147) & (g148)) + ((g1512) & (g1513) & (g1514) & (g1515) & (g147) & (!g148)) + ((g1512) & (g1513) & (g1514) & (g1515) & (g147) & (g148)));
	assign g4966 = (((!g2158) & (!g2821) & (!sk[47]) & (g1517)) + ((!g2158) & (!g2821) & (sk[47]) & (g1517)) + ((!g2158) & (g2821) & (!sk[47]) & (!g1517)) + ((!g2158) & (g2821) & (!sk[47]) & (g1517)) + ((!g2158) & (g2821) & (sk[47]) & (g1517)) + ((g2158) & (!g2821) & (!sk[47]) & (g1517)) + ((g2158) & (g2821) & (!sk[47]) & (!g1517)) + ((g2158) & (g2821) & (!sk[47]) & (g1517)) + ((g2158) & (g2821) & (sk[47]) & (!g1517)) + ((g2158) & (g2821) & (sk[47]) & (g1517)));
	assign g4967 = (((!g2159) & (!sk[48]) & (!g2821) & (g1518)) + ((!g2159) & (!sk[48]) & (g2821) & (!g1518)) + ((!g2159) & (!sk[48]) & (g2821) & (g1518)) + ((!g2159) & (sk[48]) & (!g2821) & (g1518)) + ((!g2159) & (sk[48]) & (g2821) & (g1518)) + ((g2159) & (!sk[48]) & (!g2821) & (g1518)) + ((g2159) & (!sk[48]) & (g2821) & (!g1518)) + ((g2159) & (!sk[48]) & (g2821) & (g1518)) + ((g2159) & (sk[48]) & (g2821) & (!g1518)) + ((g2159) & (sk[48]) & (g2821) & (g1518)));
	assign g4968 = (((!g2160) & (!sk[49]) & (!g2821) & (g1519)) + ((!g2160) & (!sk[49]) & (g2821) & (!g1519)) + ((!g2160) & (!sk[49]) & (g2821) & (g1519)) + ((!g2160) & (sk[49]) & (!g2821) & (g1519)) + ((!g2160) & (sk[49]) & (g2821) & (g1519)) + ((g2160) & (!sk[49]) & (!g2821) & (g1519)) + ((g2160) & (!sk[49]) & (g2821) & (!g1519)) + ((g2160) & (!sk[49]) & (g2821) & (g1519)) + ((g2160) & (sk[49]) & (g2821) & (!g1519)) + ((g2160) & (sk[49]) & (g2821) & (g1519)));
	assign g4969 = (((!g2161) & (!g2821) & (!sk[50]) & (g1520)) + ((!g2161) & (!g2821) & (sk[50]) & (g1520)) + ((!g2161) & (g2821) & (!sk[50]) & (!g1520)) + ((!g2161) & (g2821) & (!sk[50]) & (g1520)) + ((!g2161) & (g2821) & (sk[50]) & (g1520)) + ((g2161) & (!g2821) & (!sk[50]) & (g1520)) + ((g2161) & (g2821) & (!sk[50]) & (!g1520)) + ((g2161) & (g2821) & (!sk[50]) & (g1520)) + ((g2161) & (g2821) & (sk[50]) & (!g1520)) + ((g2161) & (g2821) & (sk[50]) & (g1520)));
	assign g1521 = (((!g1517) & (!g1518) & (!g1519) & (g1520) & (g147) & (g148)) + ((!g1517) & (!g1518) & (g1519) & (!g1520) & (!g147) & (g148)) + ((!g1517) & (!g1518) & (g1519) & (g1520) & (!g147) & (g148)) + ((!g1517) & (!g1518) & (g1519) & (g1520) & (g147) & (g148)) + ((!g1517) & (g1518) & (!g1519) & (!g1520) & (g147) & (!g148)) + ((!g1517) & (g1518) & (!g1519) & (g1520) & (g147) & (!g148)) + ((!g1517) & (g1518) & (!g1519) & (g1520) & (g147) & (g148)) + ((!g1517) & (g1518) & (g1519) & (!g1520) & (!g147) & (g148)) + ((!g1517) & (g1518) & (g1519) & (!g1520) & (g147) & (!g148)) + ((!g1517) & (g1518) & (g1519) & (g1520) & (!g147) & (g148)) + ((!g1517) & (g1518) & (g1519) & (g1520) & (g147) & (!g148)) + ((!g1517) & (g1518) & (g1519) & (g1520) & (g147) & (g148)) + ((g1517) & (!g1518) & (!g1519) & (!g1520) & (!g147) & (!g148)) + ((g1517) & (!g1518) & (!g1519) & (g1520) & (!g147) & (!g148)) + ((g1517) & (!g1518) & (!g1519) & (g1520) & (g147) & (g148)) + ((g1517) & (!g1518) & (g1519) & (!g1520) & (!g147) & (!g148)) + ((g1517) & (!g1518) & (g1519) & (!g1520) & (!g147) & (g148)) + ((g1517) & (!g1518) & (g1519) & (g1520) & (!g147) & (!g148)) + ((g1517) & (!g1518) & (g1519) & (g1520) & (!g147) & (g148)) + ((g1517) & (!g1518) & (g1519) & (g1520) & (g147) & (g148)) + ((g1517) & (g1518) & (!g1519) & (!g1520) & (!g147) & (!g148)) + ((g1517) & (g1518) & (!g1519) & (!g1520) & (g147) & (!g148)) + ((g1517) & (g1518) & (!g1519) & (g1520) & (!g147) & (!g148)) + ((g1517) & (g1518) & (!g1519) & (g1520) & (g147) & (!g148)) + ((g1517) & (g1518) & (!g1519) & (g1520) & (g147) & (g148)) + ((g1517) & (g1518) & (g1519) & (!g1520) & (!g147) & (!g148)) + ((g1517) & (g1518) & (g1519) & (!g1520) & (!g147) & (g148)) + ((g1517) & (g1518) & (g1519) & (!g1520) & (g147) & (!g148)) + ((g1517) & (g1518) & (g1519) & (g1520) & (!g147) & (!g148)) + ((g1517) & (g1518) & (g1519) & (g1520) & (!g147) & (g148)) + ((g1517) & (g1518) & (g1519) & (g1520) & (g147) & (!g148)) + ((g1517) & (g1518) & (g1519) & (g1520) & (g147) & (g148)));
	assign g1522 = (((!g1506) & (!g1511) & (!g1516) & (g1521) & (g165) & (g166)) + ((!g1506) & (!g1511) & (g1516) & (!g1521) & (!g165) & (g166)) + ((!g1506) & (!g1511) & (g1516) & (g1521) & (!g165) & (g166)) + ((!g1506) & (!g1511) & (g1516) & (g1521) & (g165) & (g166)) + ((!g1506) & (g1511) & (!g1516) & (!g1521) & (g165) & (!g166)) + ((!g1506) & (g1511) & (!g1516) & (g1521) & (g165) & (!g166)) + ((!g1506) & (g1511) & (!g1516) & (g1521) & (g165) & (g166)) + ((!g1506) & (g1511) & (g1516) & (!g1521) & (!g165) & (g166)) + ((!g1506) & (g1511) & (g1516) & (!g1521) & (g165) & (!g166)) + ((!g1506) & (g1511) & (g1516) & (g1521) & (!g165) & (g166)) + ((!g1506) & (g1511) & (g1516) & (g1521) & (g165) & (!g166)) + ((!g1506) & (g1511) & (g1516) & (g1521) & (g165) & (g166)) + ((g1506) & (!g1511) & (!g1516) & (!g1521) & (!g165) & (!g166)) + ((g1506) & (!g1511) & (!g1516) & (g1521) & (!g165) & (!g166)) + ((g1506) & (!g1511) & (!g1516) & (g1521) & (g165) & (g166)) + ((g1506) & (!g1511) & (g1516) & (!g1521) & (!g165) & (!g166)) + ((g1506) & (!g1511) & (g1516) & (!g1521) & (!g165) & (g166)) + ((g1506) & (!g1511) & (g1516) & (g1521) & (!g165) & (!g166)) + ((g1506) & (!g1511) & (g1516) & (g1521) & (!g165) & (g166)) + ((g1506) & (!g1511) & (g1516) & (g1521) & (g165) & (g166)) + ((g1506) & (g1511) & (!g1516) & (!g1521) & (!g165) & (!g166)) + ((g1506) & (g1511) & (!g1516) & (!g1521) & (g165) & (!g166)) + ((g1506) & (g1511) & (!g1516) & (g1521) & (!g165) & (!g166)) + ((g1506) & (g1511) & (!g1516) & (g1521) & (g165) & (!g166)) + ((g1506) & (g1511) & (!g1516) & (g1521) & (g165) & (g166)) + ((g1506) & (g1511) & (g1516) & (!g1521) & (!g165) & (!g166)) + ((g1506) & (g1511) & (g1516) & (!g1521) & (!g165) & (g166)) + ((g1506) & (g1511) & (g1516) & (!g1521) & (g165) & (!g166)) + ((g1506) & (g1511) & (g1516) & (g1521) & (!g165) & (!g166)) + ((g1506) & (g1511) & (g1516) & (g1521) & (!g165) & (g166)) + ((g1506) & (g1511) & (g1516) & (g1521) & (g165) & (!g166)) + ((g1506) & (g1511) & (g1516) & (g1521) & (g165) & (g166)));
	assign g4970 = (((!g2173) & (!sk[53]) & (!g2821) & (g1523)) + ((!g2173) & (!sk[53]) & (g2821) & (!g1523)) + ((!g2173) & (!sk[53]) & (g2821) & (g1523)) + ((!g2173) & (sk[53]) & (!g2821) & (g1523)) + ((!g2173) & (sk[53]) & (g2821) & (g1523)) + ((g2173) & (!sk[53]) & (!g2821) & (g1523)) + ((g2173) & (!sk[53]) & (g2821) & (!g1523)) + ((g2173) & (!sk[53]) & (g2821) & (g1523)) + ((g2173) & (sk[53]) & (g2821) & (!g1523)) + ((g2173) & (sk[53]) & (g2821) & (g1523)));
	assign g4971 = (((!g2174) & (!g2821) & (!sk[54]) & (g1524)) + ((!g2174) & (!g2821) & (sk[54]) & (g1524)) + ((!g2174) & (g2821) & (!sk[54]) & (!g1524)) + ((!g2174) & (g2821) & (!sk[54]) & (g1524)) + ((!g2174) & (g2821) & (sk[54]) & (g1524)) + ((g2174) & (!g2821) & (!sk[54]) & (g1524)) + ((g2174) & (g2821) & (!sk[54]) & (!g1524)) + ((g2174) & (g2821) & (!sk[54]) & (g1524)) + ((g2174) & (g2821) & (sk[54]) & (!g1524)) + ((g2174) & (g2821) & (sk[54]) & (g1524)));
	assign g4972 = (((!sk[55]) & (!g2175) & (!g2821) & (g1525)) + ((!sk[55]) & (!g2175) & (g2821) & (!g1525)) + ((!sk[55]) & (!g2175) & (g2821) & (g1525)) + ((!sk[55]) & (g2175) & (!g2821) & (g1525)) + ((!sk[55]) & (g2175) & (g2821) & (!g1525)) + ((!sk[55]) & (g2175) & (g2821) & (g1525)) + ((sk[55]) & (!g2175) & (!g2821) & (g1525)) + ((sk[55]) & (!g2175) & (g2821) & (g1525)) + ((sk[55]) & (g2175) & (g2821) & (!g1525)) + ((sk[55]) & (g2175) & (g2821) & (g1525)));
	assign g4973 = (((!g2176) & (!g2821) & (!sk[56]) & (g1526)) + ((!g2176) & (!g2821) & (sk[56]) & (g1526)) + ((!g2176) & (g2821) & (!sk[56]) & (!g1526)) + ((!g2176) & (g2821) & (!sk[56]) & (g1526)) + ((!g2176) & (g2821) & (sk[56]) & (g1526)) + ((g2176) & (!g2821) & (!sk[56]) & (g1526)) + ((g2176) & (g2821) & (!sk[56]) & (!g1526)) + ((g2176) & (g2821) & (!sk[56]) & (g1526)) + ((g2176) & (g2821) & (sk[56]) & (!g1526)) + ((g2176) & (g2821) & (sk[56]) & (g1526)));
	assign g1527 = (((!g1523) & (!g1524) & (!g1525) & (g1526) & (g165) & (g166)) + ((!g1523) & (!g1524) & (g1525) & (!g1526) & (!g165) & (g166)) + ((!g1523) & (!g1524) & (g1525) & (g1526) & (!g165) & (g166)) + ((!g1523) & (!g1524) & (g1525) & (g1526) & (g165) & (g166)) + ((!g1523) & (g1524) & (!g1525) & (!g1526) & (g165) & (!g166)) + ((!g1523) & (g1524) & (!g1525) & (g1526) & (g165) & (!g166)) + ((!g1523) & (g1524) & (!g1525) & (g1526) & (g165) & (g166)) + ((!g1523) & (g1524) & (g1525) & (!g1526) & (!g165) & (g166)) + ((!g1523) & (g1524) & (g1525) & (!g1526) & (g165) & (!g166)) + ((!g1523) & (g1524) & (g1525) & (g1526) & (!g165) & (g166)) + ((!g1523) & (g1524) & (g1525) & (g1526) & (g165) & (!g166)) + ((!g1523) & (g1524) & (g1525) & (g1526) & (g165) & (g166)) + ((g1523) & (!g1524) & (!g1525) & (!g1526) & (!g165) & (!g166)) + ((g1523) & (!g1524) & (!g1525) & (g1526) & (!g165) & (!g166)) + ((g1523) & (!g1524) & (!g1525) & (g1526) & (g165) & (g166)) + ((g1523) & (!g1524) & (g1525) & (!g1526) & (!g165) & (!g166)) + ((g1523) & (!g1524) & (g1525) & (!g1526) & (!g165) & (g166)) + ((g1523) & (!g1524) & (g1525) & (g1526) & (!g165) & (!g166)) + ((g1523) & (!g1524) & (g1525) & (g1526) & (!g165) & (g166)) + ((g1523) & (!g1524) & (g1525) & (g1526) & (g165) & (g166)) + ((g1523) & (g1524) & (!g1525) & (!g1526) & (!g165) & (!g166)) + ((g1523) & (g1524) & (!g1525) & (!g1526) & (g165) & (!g166)) + ((g1523) & (g1524) & (!g1525) & (g1526) & (!g165) & (!g166)) + ((g1523) & (g1524) & (!g1525) & (g1526) & (g165) & (!g166)) + ((g1523) & (g1524) & (!g1525) & (g1526) & (g165) & (g166)) + ((g1523) & (g1524) & (g1525) & (!g1526) & (!g165) & (!g166)) + ((g1523) & (g1524) & (g1525) & (!g1526) & (!g165) & (g166)) + ((g1523) & (g1524) & (g1525) & (!g1526) & (g165) & (!g166)) + ((g1523) & (g1524) & (g1525) & (g1526) & (!g165) & (!g166)) + ((g1523) & (g1524) & (g1525) & (g1526) & (!g165) & (g166)) + ((g1523) & (g1524) & (g1525) & (g1526) & (g165) & (!g166)) + ((g1523) & (g1524) & (g1525) & (g1526) & (g165) & (g166)));
	assign g4974 = (((!sk[58]) & (!g2177) & (!g2821) & (g1528)) + ((!sk[58]) & (!g2177) & (g2821) & (!g1528)) + ((!sk[58]) & (!g2177) & (g2821) & (g1528)) + ((!sk[58]) & (g2177) & (!g2821) & (g1528)) + ((!sk[58]) & (g2177) & (g2821) & (!g1528)) + ((!sk[58]) & (g2177) & (g2821) & (g1528)) + ((sk[58]) & (!g2177) & (!g2821) & (g1528)) + ((sk[58]) & (!g2177) & (g2821) & (g1528)) + ((sk[58]) & (g2177) & (g2821) & (!g1528)) + ((sk[58]) & (g2177) & (g2821) & (g1528)));
	assign g4975 = (((!sk[59]) & (!g2178) & (!g2821) & (g1529)) + ((!sk[59]) & (!g2178) & (g2821) & (!g1529)) + ((!sk[59]) & (!g2178) & (g2821) & (g1529)) + ((!sk[59]) & (g2178) & (!g2821) & (g1529)) + ((!sk[59]) & (g2178) & (g2821) & (!g1529)) + ((!sk[59]) & (g2178) & (g2821) & (g1529)) + ((sk[59]) & (!g2178) & (!g2821) & (g1529)) + ((sk[59]) & (!g2178) & (g2821) & (g1529)) + ((sk[59]) & (g2178) & (g2821) & (!g1529)) + ((sk[59]) & (g2178) & (g2821) & (g1529)));
	assign g4976 = (((!g2179) & (!sk[60]) & (!g2821) & (g1530)) + ((!g2179) & (!sk[60]) & (g2821) & (!g1530)) + ((!g2179) & (!sk[60]) & (g2821) & (g1530)) + ((!g2179) & (sk[60]) & (!g2821) & (g1530)) + ((!g2179) & (sk[60]) & (g2821) & (g1530)) + ((g2179) & (!sk[60]) & (!g2821) & (g1530)) + ((g2179) & (!sk[60]) & (g2821) & (!g1530)) + ((g2179) & (!sk[60]) & (g2821) & (g1530)) + ((g2179) & (sk[60]) & (g2821) & (!g1530)) + ((g2179) & (sk[60]) & (g2821) & (g1530)));
	assign g1531 = (((!g165) & (!g166) & (!g1528) & (g1529) & (!sk[61]) & (!g1530)) + ((!g165) & (!g166) & (!g1528) & (g1529) & (!sk[61]) & (g1530)) + ((!g165) & (!g166) & (g1528) & (!g1529) & (!sk[61]) & (!g1530)) + ((!g165) & (!g166) & (g1528) & (!g1529) & (!sk[61]) & (g1530)) + ((!g165) & (!g166) & (g1528) & (g1529) & (!sk[61]) & (!g1530)) + ((!g165) & (!g166) & (g1528) & (g1529) & (!sk[61]) & (g1530)) + ((!g165) & (g166) & (!g1528) & (!g1529) & (!sk[61]) & (!g1530)) + ((!g165) & (g166) & (!g1528) & (!g1529) & (!sk[61]) & (g1530)) + ((!g165) & (g166) & (!g1528) & (!g1529) & (sk[61]) & (g1530)) + ((!g165) & (g166) & (!g1528) & (g1529) & (!sk[61]) & (!g1530)) + ((!g165) & (g166) & (!g1528) & (g1529) & (!sk[61]) & (g1530)) + ((!g165) & (g166) & (!g1528) & (g1529) & (sk[61]) & (g1530)) + ((!g165) & (g166) & (g1528) & (!g1529) & (!sk[61]) & (!g1530)) + ((!g165) & (g166) & (g1528) & (!g1529) & (!sk[61]) & (g1530)) + ((!g165) & (g166) & (g1528) & (!g1529) & (sk[61]) & (g1530)) + ((!g165) & (g166) & (g1528) & (g1529) & (!sk[61]) & (!g1530)) + ((!g165) & (g166) & (g1528) & (g1529) & (!sk[61]) & (g1530)) + ((!g165) & (g166) & (g1528) & (g1529) & (sk[61]) & (g1530)) + ((g165) & (!g166) & (!g1528) & (g1529) & (!sk[61]) & (!g1530)) + ((g165) & (!g166) & (!g1528) & (g1529) & (!sk[61]) & (g1530)) + ((g165) & (!g166) & (g1528) & (!g1529) & (!sk[61]) & (!g1530)) + ((g165) & (!g166) & (g1528) & (!g1529) & (!sk[61]) & (g1530)) + ((g165) & (!g166) & (g1528) & (!g1529) & (sk[61]) & (!g1530)) + ((g165) & (!g166) & (g1528) & (!g1529) & (sk[61]) & (g1530)) + ((g165) & (!g166) & (g1528) & (g1529) & (!sk[61]) & (!g1530)) + ((g165) & (!g166) & (g1528) & (g1529) & (!sk[61]) & (g1530)) + ((g165) & (!g166) & (g1528) & (g1529) & (sk[61]) & (!g1530)) + ((g165) & (!g166) & (g1528) & (g1529) & (sk[61]) & (g1530)) + ((g165) & (g166) & (!g1528) & (!g1529) & (!sk[61]) & (!g1530)) + ((g165) & (g166) & (!g1528) & (!g1529) & (!sk[61]) & (g1530)) + ((g165) & (g166) & (!g1528) & (g1529) & (!sk[61]) & (!g1530)) + ((g165) & (g166) & (!g1528) & (g1529) & (!sk[61]) & (g1530)) + ((g165) & (g166) & (!g1528) & (g1529) & (sk[61]) & (!g1530)) + ((g165) & (g166) & (!g1528) & (g1529) & (sk[61]) & (g1530)) + ((g165) & (g166) & (g1528) & (!g1529) & (!sk[61]) & (!g1530)) + ((g165) & (g166) & (g1528) & (!g1529) & (!sk[61]) & (g1530)) + ((g165) & (g166) & (g1528) & (g1529) & (!sk[61]) & (!g1530)) + ((g165) & (g166) & (g1528) & (g1529) & (!sk[61]) & (g1530)) + ((g165) & (g166) & (g1528) & (g1529) & (sk[61]) & (!g1530)) + ((g165) & (g166) & (g1528) & (g1529) & (sk[61]) & (g1530)));
	assign g4977 = (((!g2162) & (!g2821) & (!sk[62]) & (g1532)) + ((!g2162) & (!g2821) & (sk[62]) & (g1532)) + ((!g2162) & (g2821) & (!sk[62]) & (!g1532)) + ((!g2162) & (g2821) & (!sk[62]) & (g1532)) + ((!g2162) & (g2821) & (sk[62]) & (g1532)) + ((g2162) & (!g2821) & (!sk[62]) & (g1532)) + ((g2162) & (g2821) & (!sk[62]) & (!g1532)) + ((g2162) & (g2821) & (!sk[62]) & (g1532)) + ((g2162) & (g2821) & (sk[62]) & (!g1532)) + ((g2162) & (g2821) & (sk[62]) & (g1532)));
	assign g4978 = (((!g2164) & (!g2821) & (!sk[63]) & (g1533)) + ((!g2164) & (!g2821) & (sk[63]) & (g1533)) + ((!g2164) & (g2821) & (!sk[63]) & (!g1533)) + ((!g2164) & (g2821) & (!sk[63]) & (g1533)) + ((!g2164) & (g2821) & (sk[63]) & (g1533)) + ((g2164) & (!g2821) & (!sk[63]) & (g1533)) + ((g2164) & (g2821) & (!sk[63]) & (!g1533)) + ((g2164) & (g2821) & (!sk[63]) & (g1533)) + ((g2164) & (g2821) & (sk[63]) & (!g1533)) + ((g2164) & (g2821) & (sk[63]) & (g1533)));
	assign g4979 = (((!g2166) & (!g2821) & (!sk[64]) & (g1534)) + ((!g2166) & (!g2821) & (sk[64]) & (g1534)) + ((!g2166) & (g2821) & (!sk[64]) & (!g1534)) + ((!g2166) & (g2821) & (!sk[64]) & (g1534)) + ((!g2166) & (g2821) & (sk[64]) & (g1534)) + ((g2166) & (!g2821) & (!sk[64]) & (g1534)) + ((g2166) & (g2821) & (!sk[64]) & (!g1534)) + ((g2166) & (g2821) & (!sk[64]) & (g1534)) + ((g2166) & (g2821) & (sk[64]) & (!g1534)) + ((g2166) & (g2821) & (sk[64]) & (g1534)));
	assign g4980 = (((!sk[65]) & (!g2168) & (!g2821) & (g1535)) + ((!sk[65]) & (!g2168) & (g2821) & (!g1535)) + ((!sk[65]) & (!g2168) & (g2821) & (g1535)) + ((!sk[65]) & (g2168) & (!g2821) & (g1535)) + ((!sk[65]) & (g2168) & (g2821) & (!g1535)) + ((!sk[65]) & (g2168) & (g2821) & (g1535)) + ((sk[65]) & (!g2168) & (!g2821) & (g1535)) + ((sk[65]) & (!g2168) & (g2821) & (g1535)) + ((sk[65]) & (g2168) & (g2821) & (!g1535)) + ((sk[65]) & (g2168) & (g2821) & (g1535)));
	assign g1536 = (((!g1532) & (!g1533) & (!g1534) & (g1535) & (g165) & (g166)) + ((!g1532) & (!g1533) & (g1534) & (!g1535) & (!g165) & (g166)) + ((!g1532) & (!g1533) & (g1534) & (g1535) & (!g165) & (g166)) + ((!g1532) & (!g1533) & (g1534) & (g1535) & (g165) & (g166)) + ((!g1532) & (g1533) & (!g1534) & (!g1535) & (g165) & (!g166)) + ((!g1532) & (g1533) & (!g1534) & (g1535) & (g165) & (!g166)) + ((!g1532) & (g1533) & (!g1534) & (g1535) & (g165) & (g166)) + ((!g1532) & (g1533) & (g1534) & (!g1535) & (!g165) & (g166)) + ((!g1532) & (g1533) & (g1534) & (!g1535) & (g165) & (!g166)) + ((!g1532) & (g1533) & (g1534) & (g1535) & (!g165) & (g166)) + ((!g1532) & (g1533) & (g1534) & (g1535) & (g165) & (!g166)) + ((!g1532) & (g1533) & (g1534) & (g1535) & (g165) & (g166)) + ((g1532) & (!g1533) & (!g1534) & (!g1535) & (!g165) & (!g166)) + ((g1532) & (!g1533) & (!g1534) & (g1535) & (!g165) & (!g166)) + ((g1532) & (!g1533) & (!g1534) & (g1535) & (g165) & (g166)) + ((g1532) & (!g1533) & (g1534) & (!g1535) & (!g165) & (!g166)) + ((g1532) & (!g1533) & (g1534) & (!g1535) & (!g165) & (g166)) + ((g1532) & (!g1533) & (g1534) & (g1535) & (!g165) & (!g166)) + ((g1532) & (!g1533) & (g1534) & (g1535) & (!g165) & (g166)) + ((g1532) & (!g1533) & (g1534) & (g1535) & (g165) & (g166)) + ((g1532) & (g1533) & (!g1534) & (!g1535) & (!g165) & (!g166)) + ((g1532) & (g1533) & (!g1534) & (!g1535) & (g165) & (!g166)) + ((g1532) & (g1533) & (!g1534) & (g1535) & (!g165) & (!g166)) + ((g1532) & (g1533) & (!g1534) & (g1535) & (g165) & (!g166)) + ((g1532) & (g1533) & (!g1534) & (g1535) & (g165) & (g166)) + ((g1532) & (g1533) & (g1534) & (!g1535) & (!g165) & (!g166)) + ((g1532) & (g1533) & (g1534) & (!g1535) & (!g165) & (g166)) + ((g1532) & (g1533) & (g1534) & (!g1535) & (g165) & (!g166)) + ((g1532) & (g1533) & (g1534) & (g1535) & (!g165) & (!g166)) + ((g1532) & (g1533) & (g1534) & (g1535) & (!g165) & (g166)) + ((g1532) & (g1533) & (g1534) & (g1535) & (g165) & (!g166)) + ((g1532) & (g1533) & (g1534) & (g1535) & (g165) & (g166)));
	assign g4981 = (((!sk[67]) & (!g2169) & (!g2821) & (g1537)) + ((!sk[67]) & (!g2169) & (g2821) & (!g1537)) + ((!sk[67]) & (!g2169) & (g2821) & (g1537)) + ((!sk[67]) & (g2169) & (!g2821) & (g1537)) + ((!sk[67]) & (g2169) & (g2821) & (!g1537)) + ((!sk[67]) & (g2169) & (g2821) & (g1537)) + ((sk[67]) & (!g2169) & (!g2821) & (g1537)) + ((sk[67]) & (!g2169) & (g2821) & (g1537)) + ((sk[67]) & (g2169) & (g2821) & (!g1537)) + ((sk[67]) & (g2169) & (g2821) & (g1537)));
	assign g4982 = (((!g2170) & (!sk[68]) & (!g2821) & (g1538)) + ((!g2170) & (!sk[68]) & (g2821) & (!g1538)) + ((!g2170) & (!sk[68]) & (g2821) & (g1538)) + ((!g2170) & (sk[68]) & (!g2821) & (g1538)) + ((!g2170) & (sk[68]) & (g2821) & (g1538)) + ((g2170) & (!sk[68]) & (!g2821) & (g1538)) + ((g2170) & (!sk[68]) & (g2821) & (!g1538)) + ((g2170) & (!sk[68]) & (g2821) & (g1538)) + ((g2170) & (sk[68]) & (g2821) & (!g1538)) + ((g2170) & (sk[68]) & (g2821) & (g1538)));
	assign g4983 = (((!sk[69]) & (!g2171) & (!g2821) & (g1539)) + ((!sk[69]) & (!g2171) & (g2821) & (!g1539)) + ((!sk[69]) & (!g2171) & (g2821) & (g1539)) + ((!sk[69]) & (g2171) & (!g2821) & (g1539)) + ((!sk[69]) & (g2171) & (g2821) & (!g1539)) + ((!sk[69]) & (g2171) & (g2821) & (g1539)) + ((sk[69]) & (!g2171) & (!g2821) & (g1539)) + ((sk[69]) & (!g2171) & (g2821) & (g1539)) + ((sk[69]) & (g2171) & (g2821) & (!g1539)) + ((sk[69]) & (g2171) & (g2821) & (g1539)));
	assign g4984 = (((!sk[70]) & (!g2172) & (!g2821) & (g1540)) + ((!sk[70]) & (!g2172) & (g2821) & (!g1540)) + ((!sk[70]) & (!g2172) & (g2821) & (g1540)) + ((!sk[70]) & (g2172) & (!g2821) & (g1540)) + ((!sk[70]) & (g2172) & (g2821) & (!g1540)) + ((!sk[70]) & (g2172) & (g2821) & (g1540)) + ((sk[70]) & (!g2172) & (!g2821) & (g1540)) + ((sk[70]) & (!g2172) & (g2821) & (g1540)) + ((sk[70]) & (g2172) & (g2821) & (!g1540)) + ((sk[70]) & (g2172) & (g2821) & (g1540)));
	assign g1541 = (((!g1537) & (!g1538) & (!g1539) & (g1540) & (g165) & (g166)) + ((!g1537) & (!g1538) & (g1539) & (!g1540) & (!g165) & (g166)) + ((!g1537) & (!g1538) & (g1539) & (g1540) & (!g165) & (g166)) + ((!g1537) & (!g1538) & (g1539) & (g1540) & (g165) & (g166)) + ((!g1537) & (g1538) & (!g1539) & (!g1540) & (g165) & (!g166)) + ((!g1537) & (g1538) & (!g1539) & (g1540) & (g165) & (!g166)) + ((!g1537) & (g1538) & (!g1539) & (g1540) & (g165) & (g166)) + ((!g1537) & (g1538) & (g1539) & (!g1540) & (!g165) & (g166)) + ((!g1537) & (g1538) & (g1539) & (!g1540) & (g165) & (!g166)) + ((!g1537) & (g1538) & (g1539) & (g1540) & (!g165) & (g166)) + ((!g1537) & (g1538) & (g1539) & (g1540) & (g165) & (!g166)) + ((!g1537) & (g1538) & (g1539) & (g1540) & (g165) & (g166)) + ((g1537) & (!g1538) & (!g1539) & (!g1540) & (!g165) & (!g166)) + ((g1537) & (!g1538) & (!g1539) & (g1540) & (!g165) & (!g166)) + ((g1537) & (!g1538) & (!g1539) & (g1540) & (g165) & (g166)) + ((g1537) & (!g1538) & (g1539) & (!g1540) & (!g165) & (!g166)) + ((g1537) & (!g1538) & (g1539) & (!g1540) & (!g165) & (g166)) + ((g1537) & (!g1538) & (g1539) & (g1540) & (!g165) & (!g166)) + ((g1537) & (!g1538) & (g1539) & (g1540) & (!g165) & (g166)) + ((g1537) & (!g1538) & (g1539) & (g1540) & (g165) & (g166)) + ((g1537) & (g1538) & (!g1539) & (!g1540) & (!g165) & (!g166)) + ((g1537) & (g1538) & (!g1539) & (!g1540) & (g165) & (!g166)) + ((g1537) & (g1538) & (!g1539) & (g1540) & (!g165) & (!g166)) + ((g1537) & (g1538) & (!g1539) & (g1540) & (g165) & (!g166)) + ((g1537) & (g1538) & (!g1539) & (g1540) & (g165) & (g166)) + ((g1537) & (g1538) & (g1539) & (!g1540) & (!g165) & (!g166)) + ((g1537) & (g1538) & (g1539) & (!g1540) & (!g165) & (g166)) + ((g1537) & (g1538) & (g1539) & (!g1540) & (g165) & (!g166)) + ((g1537) & (g1538) & (g1539) & (g1540) & (!g165) & (!g166)) + ((g1537) & (g1538) & (g1539) & (g1540) & (!g165) & (g166)) + ((g1537) & (g1538) & (g1539) & (g1540) & (g165) & (!g166)) + ((g1537) & (g1538) & (g1539) & (g1540) & (g165) & (g166)));
	assign g1542 = (((!g147) & (!g148) & (!g1527) & (g1531) & (!g1536) & (!g1541)) + ((!g147) & (!g148) & (!g1527) & (g1531) & (!g1536) & (g1541)) + ((!g147) & (!g148) & (!g1527) & (g1531) & (g1536) & (!g1541)) + ((!g147) & (!g148) & (!g1527) & (g1531) & (g1536) & (g1541)) + ((!g147) & (!g148) & (g1527) & (g1531) & (!g1536) & (!g1541)) + ((!g147) & (!g148) & (g1527) & (g1531) & (!g1536) & (g1541)) + ((!g147) & (!g148) & (g1527) & (g1531) & (g1536) & (!g1541)) + ((!g147) & (!g148) & (g1527) & (g1531) & (g1536) & (g1541)) + ((!g147) & (g148) & (!g1527) & (!g1531) & (!g1536) & (g1541)) + ((!g147) & (g148) & (!g1527) & (!g1531) & (g1536) & (g1541)) + ((!g147) & (g148) & (!g1527) & (g1531) & (!g1536) & (g1541)) + ((!g147) & (g148) & (!g1527) & (g1531) & (g1536) & (g1541)) + ((!g147) & (g148) & (g1527) & (!g1531) & (!g1536) & (g1541)) + ((!g147) & (g148) & (g1527) & (!g1531) & (g1536) & (g1541)) + ((!g147) & (g148) & (g1527) & (g1531) & (!g1536) & (g1541)) + ((!g147) & (g148) & (g1527) & (g1531) & (g1536) & (g1541)) + ((g147) & (!g148) & (g1527) & (!g1531) & (!g1536) & (!g1541)) + ((g147) & (!g148) & (g1527) & (!g1531) & (!g1536) & (g1541)) + ((g147) & (!g148) & (g1527) & (!g1531) & (g1536) & (!g1541)) + ((g147) & (!g148) & (g1527) & (!g1531) & (g1536) & (g1541)) + ((g147) & (!g148) & (g1527) & (g1531) & (!g1536) & (!g1541)) + ((g147) & (!g148) & (g1527) & (g1531) & (!g1536) & (g1541)) + ((g147) & (!g148) & (g1527) & (g1531) & (g1536) & (!g1541)) + ((g147) & (!g148) & (g1527) & (g1531) & (g1536) & (g1541)) + ((g147) & (g148) & (!g1527) & (!g1531) & (g1536) & (!g1541)) + ((g147) & (g148) & (!g1527) & (!g1531) & (g1536) & (g1541)) + ((g147) & (g148) & (!g1527) & (g1531) & (g1536) & (!g1541)) + ((g147) & (g148) & (!g1527) & (g1531) & (g1536) & (g1541)) + ((g147) & (g148) & (g1527) & (!g1531) & (g1536) & (!g1541)) + ((g147) & (g148) & (g1527) & (!g1531) & (g1536) & (g1541)) + ((g147) & (g148) & (g1527) & (g1531) & (g1536) & (!g1541)) + ((g147) & (g148) & (g1527) & (g1531) & (g1536) & (g1541)));
	assign g1543 = (((!sk[73]) & (!g142) & (!g1522) & (g1542)) + ((!sk[73]) & (!g142) & (g1522) & (!g1542)) + ((!sk[73]) & (!g142) & (g1522) & (g1542)) + ((!sk[73]) & (g142) & (!g1522) & (g1542)) + ((!sk[73]) & (g142) & (g1522) & (!g1542)) + ((!sk[73]) & (g142) & (g1522) & (g1542)) + ((sk[73]) & (!g142) & (!g1522) & (g1542)) + ((sk[73]) & (!g142) & (g1522) & (g1542)) + ((sk[73]) & (g142) & (g1522) & (!g1542)) + ((sk[73]) & (g142) & (g1522) & (g1542)));
	assign g4985 = (((!g2059) & (!g2825) & (!sk[74]) & (g1544)) + ((!g2059) & (!g2825) & (sk[74]) & (g1544)) + ((!g2059) & (g2825) & (!sk[74]) & (!g1544)) + ((!g2059) & (g2825) & (!sk[74]) & (g1544)) + ((!g2059) & (g2825) & (sk[74]) & (g1544)) + ((g2059) & (!g2825) & (!sk[74]) & (g1544)) + ((g2059) & (g2825) & (!sk[74]) & (!g1544)) + ((g2059) & (g2825) & (!sk[74]) & (g1544)) + ((g2059) & (g2825) & (sk[74]) & (!g1544)) + ((g2059) & (g2825) & (sk[74]) & (g1544)));
	assign g1545 = (((!sk[75]) & (!g1454) & (!g1499) & (!g1456) & (g916)) + ((!sk[75]) & (!g1454) & (!g1499) & (g1456) & (!g916)) + ((!sk[75]) & (!g1454) & (!g1499) & (g1456) & (g916)) + ((!sk[75]) & (!g1454) & (g1499) & (!g1456) & (!g916)) + ((!sk[75]) & (!g1454) & (g1499) & (!g1456) & (g916)) + ((!sk[75]) & (!g1454) & (g1499) & (g1456) & (!g916)) + ((!sk[75]) & (!g1454) & (g1499) & (g1456) & (g916)) + ((!sk[75]) & (g1454) & (!g1499) & (!g1456) & (g916)) + ((!sk[75]) & (g1454) & (!g1499) & (g1456) & (!g916)) + ((!sk[75]) & (g1454) & (!g1499) & (g1456) & (g916)) + ((!sk[75]) & (g1454) & (g1499) & (!g1456) & (!g916)) + ((!sk[75]) & (g1454) & (g1499) & (!g1456) & (g916)) + ((!sk[75]) & (g1454) & (g1499) & (g1456) & (!g916)) + ((!sk[75]) & (g1454) & (g1499) & (g1456) & (g916)) + ((sk[75]) & (!g1454) & (!g1499) & (!g1456) & (!g916)) + ((sk[75]) & (!g1454) & (g1499) & (!g1456) & (!g916)) + ((sk[75]) & (!g1454) & (g1499) & (g1456) & (!g916)) + ((sk[75]) & (g1454) & (!g1499) & (!g1456) & (!g916)) + ((sk[75]) & (g1454) & (!g1499) & (g1456) & (!g916)) + ((sk[75]) & (g1454) & (g1499) & (!g1456) & (!g916)) + ((sk[75]) & (g1454) & (g1499) & (!g1456) & (g916)) + ((sk[75]) & (g1454) & (g1499) & (g1456) & (!g916)));
	assign g1546 = (((!g126) & (!g1543) & (!g1544) & (!sk[76]) & (g1545) & (!g916)) + ((!g126) & (!g1543) & (!g1544) & (!sk[76]) & (g1545) & (g916)) + ((!g126) & (!g1543) & (g1544) & (!sk[76]) & (!g1545) & (!g916)) + ((!g126) & (!g1543) & (g1544) & (!sk[76]) & (!g1545) & (g916)) + ((!g126) & (!g1543) & (g1544) & (!sk[76]) & (g1545) & (!g916)) + ((!g126) & (!g1543) & (g1544) & (!sk[76]) & (g1545) & (g916)) + ((!g126) & (!g1543) & (g1544) & (sk[76]) & (!g1545) & (!g916)) + ((!g126) & (!g1543) & (g1544) & (sk[76]) & (!g1545) & (g916)) + ((!g126) & (!g1543) & (g1544) & (sk[76]) & (g1545) & (!g916)) + ((!g126) & (!g1543) & (g1544) & (sk[76]) & (g1545) & (g916)) + ((!g126) & (g1543) & (!g1544) & (!sk[76]) & (!g1545) & (!g916)) + ((!g126) & (g1543) & (!g1544) & (!sk[76]) & (!g1545) & (g916)) + ((!g126) & (g1543) & (!g1544) & (!sk[76]) & (g1545) & (!g916)) + ((!g126) & (g1543) & (!g1544) & (!sk[76]) & (g1545) & (g916)) + ((!g126) & (g1543) & (g1544) & (!sk[76]) & (!g1545) & (!g916)) + ((!g126) & (g1543) & (g1544) & (!sk[76]) & (!g1545) & (g916)) + ((!g126) & (g1543) & (g1544) & (!sk[76]) & (g1545) & (!g916)) + ((!g126) & (g1543) & (g1544) & (!sk[76]) & (g1545) & (g916)) + ((!g126) & (g1543) & (g1544) & (sk[76]) & (!g1545) & (!g916)) + ((!g126) & (g1543) & (g1544) & (sk[76]) & (!g1545) & (g916)) + ((!g126) & (g1543) & (g1544) & (sk[76]) & (g1545) & (!g916)) + ((!g126) & (g1543) & (g1544) & (sk[76]) & (g1545) & (g916)) + ((g126) & (!g1543) & (!g1544) & (!sk[76]) & (g1545) & (!g916)) + ((g126) & (!g1543) & (!g1544) & (!sk[76]) & (g1545) & (g916)) + ((g126) & (!g1543) & (!g1544) & (sk[76]) & (!g1545) & (!g916)) + ((g126) & (!g1543) & (!g1544) & (sk[76]) & (g1545) & (g916)) + ((g126) & (!g1543) & (g1544) & (!sk[76]) & (!g1545) & (!g916)) + ((g126) & (!g1543) & (g1544) & (!sk[76]) & (!g1545) & (g916)) + ((g126) & (!g1543) & (g1544) & (!sk[76]) & (g1545) & (!g916)) + ((g126) & (!g1543) & (g1544) & (!sk[76]) & (g1545) & (g916)) + ((g126) & (!g1543) & (g1544) & (sk[76]) & (!g1545) & (!g916)) + ((g126) & (!g1543) & (g1544) & (sk[76]) & (g1545) & (g916)) + ((g126) & (g1543) & (!g1544) & (!sk[76]) & (!g1545) & (!g916)) + ((g126) & (g1543) & (!g1544) & (!sk[76]) & (!g1545) & (g916)) + ((g126) & (g1543) & (!g1544) & (!sk[76]) & (g1545) & (!g916)) + ((g126) & (g1543) & (!g1544) & (!sk[76]) & (g1545) & (g916)) + ((g126) & (g1543) & (!g1544) & (sk[76]) & (!g1545) & (g916)) + ((g126) & (g1543) & (!g1544) & (sk[76]) & (g1545) & (!g916)) + ((g126) & (g1543) & (g1544) & (!sk[76]) & (!g1545) & (!g916)) + ((g126) & (g1543) & (g1544) & (!sk[76]) & (!g1545) & (g916)) + ((g126) & (g1543) & (g1544) & (!sk[76]) & (g1545) & (!g916)) + ((g126) & (g1543) & (g1544) & (!sk[76]) & (g1545) & (g916)) + ((g126) & (g1543) & (g1544) & (sk[76]) & (!g1545) & (g916)) + ((g126) & (g1543) & (g1544) & (sk[76]) & (g1545) & (!g916)));
	assign g4986 = (((!g2059) & (!sk[77]) & (!g2830) & (g1547)) + ((!g2059) & (!sk[77]) & (g2830) & (!g1547)) + ((!g2059) & (!sk[77]) & (g2830) & (g1547)) + ((!g2059) & (sk[77]) & (!g2830) & (g1547)) + ((!g2059) & (sk[77]) & (g2830) & (g1547)) + ((g2059) & (!sk[77]) & (!g2830) & (g1547)) + ((g2059) & (!sk[77]) & (g2830) & (!g1547)) + ((g2059) & (!sk[77]) & (g2830) & (g1547)) + ((g2059) & (sk[77]) & (g2830) & (!g1547)) + ((g2059) & (sk[77]) & (g2830) & (g1547)));
	assign g4987 = (((!g2140) & (!g2841) & (!sk[78]) & (g1548)) + ((!g2140) & (!g2841) & (sk[78]) & (g1548)) + ((!g2140) & (g2841) & (!sk[78]) & (!g1548)) + ((!g2140) & (g2841) & (!sk[78]) & (g1548)) + ((!g2140) & (g2841) & (sk[78]) & (g1548)) + ((g2140) & (!g2841) & (!sk[78]) & (g1548)) + ((g2140) & (g2841) & (!sk[78]) & (!g1548)) + ((g2140) & (g2841) & (!sk[78]) & (g1548)) + ((g2140) & (g2841) & (sk[78]) & (!g1548)) + ((g2140) & (g2841) & (sk[78]) & (g1548)));
	assign g4988 = (((!g2142) & (!g2841) & (!sk[79]) & (g1549)) + ((!g2142) & (!g2841) & (sk[79]) & (g1549)) + ((!g2142) & (g2841) & (!sk[79]) & (!g1549)) + ((!g2142) & (g2841) & (!sk[79]) & (g1549)) + ((!g2142) & (g2841) & (sk[79]) & (g1549)) + ((g2142) & (!g2841) & (!sk[79]) & (g1549)) + ((g2142) & (g2841) & (!sk[79]) & (!g1549)) + ((g2142) & (g2841) & (!sk[79]) & (g1549)) + ((g2142) & (g2841) & (sk[79]) & (!g1549)) + ((g2142) & (g2841) & (sk[79]) & (g1549)));
	assign g4989 = (((!sk[80]) & (!g2144) & (!g2841) & (g1550)) + ((!sk[80]) & (!g2144) & (g2841) & (!g1550)) + ((!sk[80]) & (!g2144) & (g2841) & (g1550)) + ((!sk[80]) & (g2144) & (!g2841) & (g1550)) + ((!sk[80]) & (g2144) & (g2841) & (!g1550)) + ((!sk[80]) & (g2144) & (g2841) & (g1550)) + ((sk[80]) & (!g2144) & (!g2841) & (g1550)) + ((sk[80]) & (!g2144) & (g2841) & (g1550)) + ((sk[80]) & (g2144) & (g2841) & (!g1550)) + ((sk[80]) & (g2144) & (g2841) & (g1550)));
	assign g4990 = (((!sk[81]) & (!g2145) & (!g2841) & (g1551)) + ((!sk[81]) & (!g2145) & (g2841) & (!g1551)) + ((!sk[81]) & (!g2145) & (g2841) & (g1551)) + ((!sk[81]) & (g2145) & (!g2841) & (g1551)) + ((!sk[81]) & (g2145) & (g2841) & (!g1551)) + ((!sk[81]) & (g2145) & (g2841) & (g1551)) + ((sk[81]) & (!g2145) & (!g2841) & (g1551)) + ((sk[81]) & (!g2145) & (g2841) & (g1551)) + ((sk[81]) & (g2145) & (g2841) & (!g1551)) + ((sk[81]) & (g2145) & (g2841) & (g1551)));
	assign g1552 = (((!g1548) & (!g1549) & (!g1550) & (g1551) & (g147) & (g148)) + ((!g1548) & (!g1549) & (g1550) & (!g1551) & (!g147) & (g148)) + ((!g1548) & (!g1549) & (g1550) & (g1551) & (!g147) & (g148)) + ((!g1548) & (!g1549) & (g1550) & (g1551) & (g147) & (g148)) + ((!g1548) & (g1549) & (!g1550) & (!g1551) & (g147) & (!g148)) + ((!g1548) & (g1549) & (!g1550) & (g1551) & (g147) & (!g148)) + ((!g1548) & (g1549) & (!g1550) & (g1551) & (g147) & (g148)) + ((!g1548) & (g1549) & (g1550) & (!g1551) & (!g147) & (g148)) + ((!g1548) & (g1549) & (g1550) & (!g1551) & (g147) & (!g148)) + ((!g1548) & (g1549) & (g1550) & (g1551) & (!g147) & (g148)) + ((!g1548) & (g1549) & (g1550) & (g1551) & (g147) & (!g148)) + ((!g1548) & (g1549) & (g1550) & (g1551) & (g147) & (g148)) + ((g1548) & (!g1549) & (!g1550) & (!g1551) & (!g147) & (!g148)) + ((g1548) & (!g1549) & (!g1550) & (g1551) & (!g147) & (!g148)) + ((g1548) & (!g1549) & (!g1550) & (g1551) & (g147) & (g148)) + ((g1548) & (!g1549) & (g1550) & (!g1551) & (!g147) & (!g148)) + ((g1548) & (!g1549) & (g1550) & (!g1551) & (!g147) & (g148)) + ((g1548) & (!g1549) & (g1550) & (g1551) & (!g147) & (!g148)) + ((g1548) & (!g1549) & (g1550) & (g1551) & (!g147) & (g148)) + ((g1548) & (!g1549) & (g1550) & (g1551) & (g147) & (g148)) + ((g1548) & (g1549) & (!g1550) & (!g1551) & (!g147) & (!g148)) + ((g1548) & (g1549) & (!g1550) & (!g1551) & (g147) & (!g148)) + ((g1548) & (g1549) & (!g1550) & (g1551) & (!g147) & (!g148)) + ((g1548) & (g1549) & (!g1550) & (g1551) & (g147) & (!g148)) + ((g1548) & (g1549) & (!g1550) & (g1551) & (g147) & (g148)) + ((g1548) & (g1549) & (g1550) & (!g1551) & (!g147) & (!g148)) + ((g1548) & (g1549) & (g1550) & (!g1551) & (!g147) & (g148)) + ((g1548) & (g1549) & (g1550) & (!g1551) & (g147) & (!g148)) + ((g1548) & (g1549) & (g1550) & (g1551) & (!g147) & (!g148)) + ((g1548) & (g1549) & (g1550) & (g1551) & (!g147) & (g148)) + ((g1548) & (g1549) & (g1550) & (g1551) & (g147) & (!g148)) + ((g1548) & (g1549) & (g1550) & (g1551) & (g147) & (g148)));
	assign g4991 = (((!g2146) & (!g2841) & (!sk[83]) & (g1553)) + ((!g2146) & (!g2841) & (sk[83]) & (g1553)) + ((!g2146) & (g2841) & (!sk[83]) & (!g1553)) + ((!g2146) & (g2841) & (!sk[83]) & (g1553)) + ((!g2146) & (g2841) & (sk[83]) & (g1553)) + ((g2146) & (!g2841) & (!sk[83]) & (g1553)) + ((g2146) & (g2841) & (!sk[83]) & (!g1553)) + ((g2146) & (g2841) & (!sk[83]) & (g1553)) + ((g2146) & (g2841) & (sk[83]) & (!g1553)) + ((g2146) & (g2841) & (sk[83]) & (g1553)));
	assign g4992 = (((!g2148) & (!g2841) & (!sk[84]) & (g1554)) + ((!g2148) & (!g2841) & (sk[84]) & (g1554)) + ((!g2148) & (g2841) & (!sk[84]) & (!g1554)) + ((!g2148) & (g2841) & (!sk[84]) & (g1554)) + ((!g2148) & (g2841) & (sk[84]) & (g1554)) + ((g2148) & (!g2841) & (!sk[84]) & (g1554)) + ((g2148) & (g2841) & (!sk[84]) & (!g1554)) + ((g2148) & (g2841) & (!sk[84]) & (g1554)) + ((g2148) & (g2841) & (sk[84]) & (!g1554)) + ((g2148) & (g2841) & (sk[84]) & (g1554)));
	assign g4993 = (((!sk[85]) & (!g2150) & (!g2841) & (g1555)) + ((!sk[85]) & (!g2150) & (g2841) & (!g1555)) + ((!sk[85]) & (!g2150) & (g2841) & (g1555)) + ((!sk[85]) & (g2150) & (!g2841) & (g1555)) + ((!sk[85]) & (g2150) & (g2841) & (!g1555)) + ((!sk[85]) & (g2150) & (g2841) & (g1555)) + ((sk[85]) & (!g2150) & (!g2841) & (g1555)) + ((sk[85]) & (!g2150) & (g2841) & (g1555)) + ((sk[85]) & (g2150) & (g2841) & (!g1555)) + ((sk[85]) & (g2150) & (g2841) & (g1555)));
	assign g4994 = (((!sk[86]) & (!g2151) & (!g2841) & (g1556)) + ((!sk[86]) & (!g2151) & (g2841) & (!g1556)) + ((!sk[86]) & (!g2151) & (g2841) & (g1556)) + ((!sk[86]) & (g2151) & (!g2841) & (g1556)) + ((!sk[86]) & (g2151) & (g2841) & (!g1556)) + ((!sk[86]) & (g2151) & (g2841) & (g1556)) + ((sk[86]) & (!g2151) & (!g2841) & (g1556)) + ((sk[86]) & (!g2151) & (g2841) & (g1556)) + ((sk[86]) & (g2151) & (g2841) & (!g1556)) + ((sk[86]) & (g2151) & (g2841) & (g1556)));
	assign g1557 = (((!g1553) & (!g1554) & (!g1555) & (g1556) & (g147) & (g148)) + ((!g1553) & (!g1554) & (g1555) & (!g1556) & (!g147) & (g148)) + ((!g1553) & (!g1554) & (g1555) & (g1556) & (!g147) & (g148)) + ((!g1553) & (!g1554) & (g1555) & (g1556) & (g147) & (g148)) + ((!g1553) & (g1554) & (!g1555) & (!g1556) & (g147) & (!g148)) + ((!g1553) & (g1554) & (!g1555) & (g1556) & (g147) & (!g148)) + ((!g1553) & (g1554) & (!g1555) & (g1556) & (g147) & (g148)) + ((!g1553) & (g1554) & (g1555) & (!g1556) & (!g147) & (g148)) + ((!g1553) & (g1554) & (g1555) & (!g1556) & (g147) & (!g148)) + ((!g1553) & (g1554) & (g1555) & (g1556) & (!g147) & (g148)) + ((!g1553) & (g1554) & (g1555) & (g1556) & (g147) & (!g148)) + ((!g1553) & (g1554) & (g1555) & (g1556) & (g147) & (g148)) + ((g1553) & (!g1554) & (!g1555) & (!g1556) & (!g147) & (!g148)) + ((g1553) & (!g1554) & (!g1555) & (g1556) & (!g147) & (!g148)) + ((g1553) & (!g1554) & (!g1555) & (g1556) & (g147) & (g148)) + ((g1553) & (!g1554) & (g1555) & (!g1556) & (!g147) & (!g148)) + ((g1553) & (!g1554) & (g1555) & (!g1556) & (!g147) & (g148)) + ((g1553) & (!g1554) & (g1555) & (g1556) & (!g147) & (!g148)) + ((g1553) & (!g1554) & (g1555) & (g1556) & (!g147) & (g148)) + ((g1553) & (!g1554) & (g1555) & (g1556) & (g147) & (g148)) + ((g1553) & (g1554) & (!g1555) & (!g1556) & (!g147) & (!g148)) + ((g1553) & (g1554) & (!g1555) & (!g1556) & (g147) & (!g148)) + ((g1553) & (g1554) & (!g1555) & (g1556) & (!g147) & (!g148)) + ((g1553) & (g1554) & (!g1555) & (g1556) & (g147) & (!g148)) + ((g1553) & (g1554) & (!g1555) & (g1556) & (g147) & (g148)) + ((g1553) & (g1554) & (g1555) & (!g1556) & (!g147) & (!g148)) + ((g1553) & (g1554) & (g1555) & (!g1556) & (!g147) & (g148)) + ((g1553) & (g1554) & (g1555) & (!g1556) & (g147) & (!g148)) + ((g1553) & (g1554) & (g1555) & (g1556) & (!g147) & (!g148)) + ((g1553) & (g1554) & (g1555) & (g1556) & (!g147) & (g148)) + ((g1553) & (g1554) & (g1555) & (g1556) & (g147) & (!g148)) + ((g1553) & (g1554) & (g1555) & (g1556) & (g147) & (g148)));
	assign g4995 = (((!g2152) & (!sk[88]) & (!g2841) & (g1558)) + ((!g2152) & (!sk[88]) & (g2841) & (!g1558)) + ((!g2152) & (!sk[88]) & (g2841) & (g1558)) + ((!g2152) & (sk[88]) & (!g2841) & (g1558)) + ((!g2152) & (sk[88]) & (g2841) & (g1558)) + ((g2152) & (!sk[88]) & (!g2841) & (g1558)) + ((g2152) & (!sk[88]) & (g2841) & (!g1558)) + ((g2152) & (!sk[88]) & (g2841) & (g1558)) + ((g2152) & (sk[88]) & (g2841) & (!g1558)) + ((g2152) & (sk[88]) & (g2841) & (g1558)));
	assign g4996 = (((!g2153) & (!g2841) & (!sk[89]) & (g1559)) + ((!g2153) & (!g2841) & (sk[89]) & (g1559)) + ((!g2153) & (g2841) & (!sk[89]) & (!g1559)) + ((!g2153) & (g2841) & (!sk[89]) & (g1559)) + ((!g2153) & (g2841) & (sk[89]) & (g1559)) + ((g2153) & (!g2841) & (!sk[89]) & (g1559)) + ((g2153) & (g2841) & (!sk[89]) & (!g1559)) + ((g2153) & (g2841) & (!sk[89]) & (g1559)) + ((g2153) & (g2841) & (sk[89]) & (!g1559)) + ((g2153) & (g2841) & (sk[89]) & (g1559)));
	assign g4997 = (((!sk[90]) & (!g2155) & (!g2841) & (g1560)) + ((!sk[90]) & (!g2155) & (g2841) & (!g1560)) + ((!sk[90]) & (!g2155) & (g2841) & (g1560)) + ((!sk[90]) & (g2155) & (!g2841) & (g1560)) + ((!sk[90]) & (g2155) & (g2841) & (!g1560)) + ((!sk[90]) & (g2155) & (g2841) & (g1560)) + ((sk[90]) & (!g2155) & (!g2841) & (g1560)) + ((sk[90]) & (!g2155) & (g2841) & (g1560)) + ((sk[90]) & (g2155) & (g2841) & (!g1560)) + ((sk[90]) & (g2155) & (g2841) & (g1560)));
	assign g4998 = (((!g2157) & (!sk[91]) & (!g2841) & (g1561)) + ((!g2157) & (!sk[91]) & (g2841) & (!g1561)) + ((!g2157) & (!sk[91]) & (g2841) & (g1561)) + ((!g2157) & (sk[91]) & (!g2841) & (g1561)) + ((!g2157) & (sk[91]) & (g2841) & (g1561)) + ((g2157) & (!sk[91]) & (!g2841) & (g1561)) + ((g2157) & (!sk[91]) & (g2841) & (!g1561)) + ((g2157) & (!sk[91]) & (g2841) & (g1561)) + ((g2157) & (sk[91]) & (g2841) & (!g1561)) + ((g2157) & (sk[91]) & (g2841) & (g1561)));
	assign g1562 = (((!g1558) & (!g1559) & (!g1560) & (g1561) & (g147) & (g148)) + ((!g1558) & (!g1559) & (g1560) & (!g1561) & (!g147) & (g148)) + ((!g1558) & (!g1559) & (g1560) & (g1561) & (!g147) & (g148)) + ((!g1558) & (!g1559) & (g1560) & (g1561) & (g147) & (g148)) + ((!g1558) & (g1559) & (!g1560) & (!g1561) & (g147) & (!g148)) + ((!g1558) & (g1559) & (!g1560) & (g1561) & (g147) & (!g148)) + ((!g1558) & (g1559) & (!g1560) & (g1561) & (g147) & (g148)) + ((!g1558) & (g1559) & (g1560) & (!g1561) & (!g147) & (g148)) + ((!g1558) & (g1559) & (g1560) & (!g1561) & (g147) & (!g148)) + ((!g1558) & (g1559) & (g1560) & (g1561) & (!g147) & (g148)) + ((!g1558) & (g1559) & (g1560) & (g1561) & (g147) & (!g148)) + ((!g1558) & (g1559) & (g1560) & (g1561) & (g147) & (g148)) + ((g1558) & (!g1559) & (!g1560) & (!g1561) & (!g147) & (!g148)) + ((g1558) & (!g1559) & (!g1560) & (g1561) & (!g147) & (!g148)) + ((g1558) & (!g1559) & (!g1560) & (g1561) & (g147) & (g148)) + ((g1558) & (!g1559) & (g1560) & (!g1561) & (!g147) & (!g148)) + ((g1558) & (!g1559) & (g1560) & (!g1561) & (!g147) & (g148)) + ((g1558) & (!g1559) & (g1560) & (g1561) & (!g147) & (!g148)) + ((g1558) & (!g1559) & (g1560) & (g1561) & (!g147) & (g148)) + ((g1558) & (!g1559) & (g1560) & (g1561) & (g147) & (g148)) + ((g1558) & (g1559) & (!g1560) & (!g1561) & (!g147) & (!g148)) + ((g1558) & (g1559) & (!g1560) & (!g1561) & (g147) & (!g148)) + ((g1558) & (g1559) & (!g1560) & (g1561) & (!g147) & (!g148)) + ((g1558) & (g1559) & (!g1560) & (g1561) & (g147) & (!g148)) + ((g1558) & (g1559) & (!g1560) & (g1561) & (g147) & (g148)) + ((g1558) & (g1559) & (g1560) & (!g1561) & (!g147) & (!g148)) + ((g1558) & (g1559) & (g1560) & (!g1561) & (!g147) & (g148)) + ((g1558) & (g1559) & (g1560) & (!g1561) & (g147) & (!g148)) + ((g1558) & (g1559) & (g1560) & (g1561) & (!g147) & (!g148)) + ((g1558) & (g1559) & (g1560) & (g1561) & (!g147) & (g148)) + ((g1558) & (g1559) & (g1560) & (g1561) & (g147) & (!g148)) + ((g1558) & (g1559) & (g1560) & (g1561) & (g147) & (g148)));
	assign g4999 = (((!sk[93]) & (!g2158) & (!g2841) & (g1563)) + ((!sk[93]) & (!g2158) & (g2841) & (!g1563)) + ((!sk[93]) & (!g2158) & (g2841) & (g1563)) + ((!sk[93]) & (g2158) & (!g2841) & (g1563)) + ((!sk[93]) & (g2158) & (g2841) & (!g1563)) + ((!sk[93]) & (g2158) & (g2841) & (g1563)) + ((sk[93]) & (!g2158) & (!g2841) & (g1563)) + ((sk[93]) & (!g2158) & (g2841) & (g1563)) + ((sk[93]) & (g2158) & (g2841) & (!g1563)) + ((sk[93]) & (g2158) & (g2841) & (g1563)));
	assign g5000 = (((!sk[94]) & (!g2159) & (!g2841) & (g1564)) + ((!sk[94]) & (!g2159) & (g2841) & (!g1564)) + ((!sk[94]) & (!g2159) & (g2841) & (g1564)) + ((!sk[94]) & (g2159) & (!g2841) & (g1564)) + ((!sk[94]) & (g2159) & (g2841) & (!g1564)) + ((!sk[94]) & (g2159) & (g2841) & (g1564)) + ((sk[94]) & (!g2159) & (!g2841) & (g1564)) + ((sk[94]) & (!g2159) & (g2841) & (g1564)) + ((sk[94]) & (g2159) & (g2841) & (!g1564)) + ((sk[94]) & (g2159) & (g2841) & (g1564)));
	assign g5001 = (((!g2160) & (!sk[95]) & (!g2841) & (g1565)) + ((!g2160) & (!sk[95]) & (g2841) & (!g1565)) + ((!g2160) & (!sk[95]) & (g2841) & (g1565)) + ((!g2160) & (sk[95]) & (!g2841) & (g1565)) + ((!g2160) & (sk[95]) & (g2841) & (g1565)) + ((g2160) & (!sk[95]) & (!g2841) & (g1565)) + ((g2160) & (!sk[95]) & (g2841) & (!g1565)) + ((g2160) & (!sk[95]) & (g2841) & (g1565)) + ((g2160) & (sk[95]) & (g2841) & (!g1565)) + ((g2160) & (sk[95]) & (g2841) & (g1565)));
	assign g5002 = (((!g2161) & (!sk[96]) & (!g2841) & (g1566)) + ((!g2161) & (!sk[96]) & (g2841) & (!g1566)) + ((!g2161) & (!sk[96]) & (g2841) & (g1566)) + ((!g2161) & (sk[96]) & (!g2841) & (g1566)) + ((!g2161) & (sk[96]) & (g2841) & (g1566)) + ((g2161) & (!sk[96]) & (!g2841) & (g1566)) + ((g2161) & (!sk[96]) & (g2841) & (!g1566)) + ((g2161) & (!sk[96]) & (g2841) & (g1566)) + ((g2161) & (sk[96]) & (g2841) & (!g1566)) + ((g2161) & (sk[96]) & (g2841) & (g1566)));
	assign g1567 = (((!g1563) & (!g1564) & (!g1565) & (g1566) & (g147) & (g148)) + ((!g1563) & (!g1564) & (g1565) & (!g1566) & (!g147) & (g148)) + ((!g1563) & (!g1564) & (g1565) & (g1566) & (!g147) & (g148)) + ((!g1563) & (!g1564) & (g1565) & (g1566) & (g147) & (g148)) + ((!g1563) & (g1564) & (!g1565) & (!g1566) & (g147) & (!g148)) + ((!g1563) & (g1564) & (!g1565) & (g1566) & (g147) & (!g148)) + ((!g1563) & (g1564) & (!g1565) & (g1566) & (g147) & (g148)) + ((!g1563) & (g1564) & (g1565) & (!g1566) & (!g147) & (g148)) + ((!g1563) & (g1564) & (g1565) & (!g1566) & (g147) & (!g148)) + ((!g1563) & (g1564) & (g1565) & (g1566) & (!g147) & (g148)) + ((!g1563) & (g1564) & (g1565) & (g1566) & (g147) & (!g148)) + ((!g1563) & (g1564) & (g1565) & (g1566) & (g147) & (g148)) + ((g1563) & (!g1564) & (!g1565) & (!g1566) & (!g147) & (!g148)) + ((g1563) & (!g1564) & (!g1565) & (g1566) & (!g147) & (!g148)) + ((g1563) & (!g1564) & (!g1565) & (g1566) & (g147) & (g148)) + ((g1563) & (!g1564) & (g1565) & (!g1566) & (!g147) & (!g148)) + ((g1563) & (!g1564) & (g1565) & (!g1566) & (!g147) & (g148)) + ((g1563) & (!g1564) & (g1565) & (g1566) & (!g147) & (!g148)) + ((g1563) & (!g1564) & (g1565) & (g1566) & (!g147) & (g148)) + ((g1563) & (!g1564) & (g1565) & (g1566) & (g147) & (g148)) + ((g1563) & (g1564) & (!g1565) & (!g1566) & (!g147) & (!g148)) + ((g1563) & (g1564) & (!g1565) & (!g1566) & (g147) & (!g148)) + ((g1563) & (g1564) & (!g1565) & (g1566) & (!g147) & (!g148)) + ((g1563) & (g1564) & (!g1565) & (g1566) & (g147) & (!g148)) + ((g1563) & (g1564) & (!g1565) & (g1566) & (g147) & (g148)) + ((g1563) & (g1564) & (g1565) & (!g1566) & (!g147) & (!g148)) + ((g1563) & (g1564) & (g1565) & (!g1566) & (!g147) & (g148)) + ((g1563) & (g1564) & (g1565) & (!g1566) & (g147) & (!g148)) + ((g1563) & (g1564) & (g1565) & (g1566) & (!g147) & (!g148)) + ((g1563) & (g1564) & (g1565) & (g1566) & (!g147) & (g148)) + ((g1563) & (g1564) & (g1565) & (g1566) & (g147) & (!g148)) + ((g1563) & (g1564) & (g1565) & (g1566) & (g147) & (g148)));
	assign g1568 = (((!g1552) & (!g1557) & (!g1562) & (g1567) & (g165) & (g166)) + ((!g1552) & (!g1557) & (g1562) & (!g1567) & (!g165) & (g166)) + ((!g1552) & (!g1557) & (g1562) & (g1567) & (!g165) & (g166)) + ((!g1552) & (!g1557) & (g1562) & (g1567) & (g165) & (g166)) + ((!g1552) & (g1557) & (!g1562) & (!g1567) & (g165) & (!g166)) + ((!g1552) & (g1557) & (!g1562) & (g1567) & (g165) & (!g166)) + ((!g1552) & (g1557) & (!g1562) & (g1567) & (g165) & (g166)) + ((!g1552) & (g1557) & (g1562) & (!g1567) & (!g165) & (g166)) + ((!g1552) & (g1557) & (g1562) & (!g1567) & (g165) & (!g166)) + ((!g1552) & (g1557) & (g1562) & (g1567) & (!g165) & (g166)) + ((!g1552) & (g1557) & (g1562) & (g1567) & (g165) & (!g166)) + ((!g1552) & (g1557) & (g1562) & (g1567) & (g165) & (g166)) + ((g1552) & (!g1557) & (!g1562) & (!g1567) & (!g165) & (!g166)) + ((g1552) & (!g1557) & (!g1562) & (g1567) & (!g165) & (!g166)) + ((g1552) & (!g1557) & (!g1562) & (g1567) & (g165) & (g166)) + ((g1552) & (!g1557) & (g1562) & (!g1567) & (!g165) & (!g166)) + ((g1552) & (!g1557) & (g1562) & (!g1567) & (!g165) & (g166)) + ((g1552) & (!g1557) & (g1562) & (g1567) & (!g165) & (!g166)) + ((g1552) & (!g1557) & (g1562) & (g1567) & (!g165) & (g166)) + ((g1552) & (!g1557) & (g1562) & (g1567) & (g165) & (g166)) + ((g1552) & (g1557) & (!g1562) & (!g1567) & (!g165) & (!g166)) + ((g1552) & (g1557) & (!g1562) & (!g1567) & (g165) & (!g166)) + ((g1552) & (g1557) & (!g1562) & (g1567) & (!g165) & (!g166)) + ((g1552) & (g1557) & (!g1562) & (g1567) & (g165) & (!g166)) + ((g1552) & (g1557) & (!g1562) & (g1567) & (g165) & (g166)) + ((g1552) & (g1557) & (g1562) & (!g1567) & (!g165) & (!g166)) + ((g1552) & (g1557) & (g1562) & (!g1567) & (!g165) & (g166)) + ((g1552) & (g1557) & (g1562) & (!g1567) & (g165) & (!g166)) + ((g1552) & (g1557) & (g1562) & (g1567) & (!g165) & (!g166)) + ((g1552) & (g1557) & (g1562) & (g1567) & (!g165) & (g166)) + ((g1552) & (g1557) & (g1562) & (g1567) & (g165) & (!g166)) + ((g1552) & (g1557) & (g1562) & (g1567) & (g165) & (g166)));
	assign g5003 = (((!g2173) & (!g2841) & (!sk[99]) & (g1569)) + ((!g2173) & (!g2841) & (sk[99]) & (g1569)) + ((!g2173) & (g2841) & (!sk[99]) & (!g1569)) + ((!g2173) & (g2841) & (!sk[99]) & (g1569)) + ((!g2173) & (g2841) & (sk[99]) & (g1569)) + ((g2173) & (!g2841) & (!sk[99]) & (g1569)) + ((g2173) & (g2841) & (!sk[99]) & (!g1569)) + ((g2173) & (g2841) & (!sk[99]) & (g1569)) + ((g2173) & (g2841) & (sk[99]) & (!g1569)) + ((g2173) & (g2841) & (sk[99]) & (g1569)));
	assign g5004 = (((!g2174) & (!g2841) & (!sk[100]) & (g1570)) + ((!g2174) & (!g2841) & (sk[100]) & (g1570)) + ((!g2174) & (g2841) & (!sk[100]) & (!g1570)) + ((!g2174) & (g2841) & (!sk[100]) & (g1570)) + ((!g2174) & (g2841) & (sk[100]) & (g1570)) + ((g2174) & (!g2841) & (!sk[100]) & (g1570)) + ((g2174) & (g2841) & (!sk[100]) & (!g1570)) + ((g2174) & (g2841) & (!sk[100]) & (g1570)) + ((g2174) & (g2841) & (sk[100]) & (!g1570)) + ((g2174) & (g2841) & (sk[100]) & (g1570)));
	assign g5005 = (((!sk[101]) & (!g2175) & (!g2841) & (g1571)) + ((!sk[101]) & (!g2175) & (g2841) & (!g1571)) + ((!sk[101]) & (!g2175) & (g2841) & (g1571)) + ((!sk[101]) & (g2175) & (!g2841) & (g1571)) + ((!sk[101]) & (g2175) & (g2841) & (!g1571)) + ((!sk[101]) & (g2175) & (g2841) & (g1571)) + ((sk[101]) & (!g2175) & (!g2841) & (g1571)) + ((sk[101]) & (!g2175) & (g2841) & (g1571)) + ((sk[101]) & (g2175) & (g2841) & (!g1571)) + ((sk[101]) & (g2175) & (g2841) & (g1571)));
	assign g5006 = (((!g2176) & (!g2841) & (!sk[102]) & (g1572)) + ((!g2176) & (!g2841) & (sk[102]) & (g1572)) + ((!g2176) & (g2841) & (!sk[102]) & (!g1572)) + ((!g2176) & (g2841) & (!sk[102]) & (g1572)) + ((!g2176) & (g2841) & (sk[102]) & (g1572)) + ((g2176) & (!g2841) & (!sk[102]) & (g1572)) + ((g2176) & (g2841) & (!sk[102]) & (!g1572)) + ((g2176) & (g2841) & (!sk[102]) & (g1572)) + ((g2176) & (g2841) & (sk[102]) & (!g1572)) + ((g2176) & (g2841) & (sk[102]) & (g1572)));
	assign g1573 = (((!g1569) & (!g1570) & (!g1571) & (g1572) & (g165) & (g166)) + ((!g1569) & (!g1570) & (g1571) & (!g1572) & (!g165) & (g166)) + ((!g1569) & (!g1570) & (g1571) & (g1572) & (!g165) & (g166)) + ((!g1569) & (!g1570) & (g1571) & (g1572) & (g165) & (g166)) + ((!g1569) & (g1570) & (!g1571) & (!g1572) & (g165) & (!g166)) + ((!g1569) & (g1570) & (!g1571) & (g1572) & (g165) & (!g166)) + ((!g1569) & (g1570) & (!g1571) & (g1572) & (g165) & (g166)) + ((!g1569) & (g1570) & (g1571) & (!g1572) & (!g165) & (g166)) + ((!g1569) & (g1570) & (g1571) & (!g1572) & (g165) & (!g166)) + ((!g1569) & (g1570) & (g1571) & (g1572) & (!g165) & (g166)) + ((!g1569) & (g1570) & (g1571) & (g1572) & (g165) & (!g166)) + ((!g1569) & (g1570) & (g1571) & (g1572) & (g165) & (g166)) + ((g1569) & (!g1570) & (!g1571) & (!g1572) & (!g165) & (!g166)) + ((g1569) & (!g1570) & (!g1571) & (g1572) & (!g165) & (!g166)) + ((g1569) & (!g1570) & (!g1571) & (g1572) & (g165) & (g166)) + ((g1569) & (!g1570) & (g1571) & (!g1572) & (!g165) & (!g166)) + ((g1569) & (!g1570) & (g1571) & (!g1572) & (!g165) & (g166)) + ((g1569) & (!g1570) & (g1571) & (g1572) & (!g165) & (!g166)) + ((g1569) & (!g1570) & (g1571) & (g1572) & (!g165) & (g166)) + ((g1569) & (!g1570) & (g1571) & (g1572) & (g165) & (g166)) + ((g1569) & (g1570) & (!g1571) & (!g1572) & (!g165) & (!g166)) + ((g1569) & (g1570) & (!g1571) & (!g1572) & (g165) & (!g166)) + ((g1569) & (g1570) & (!g1571) & (g1572) & (!g165) & (!g166)) + ((g1569) & (g1570) & (!g1571) & (g1572) & (g165) & (!g166)) + ((g1569) & (g1570) & (!g1571) & (g1572) & (g165) & (g166)) + ((g1569) & (g1570) & (g1571) & (!g1572) & (!g165) & (!g166)) + ((g1569) & (g1570) & (g1571) & (!g1572) & (!g165) & (g166)) + ((g1569) & (g1570) & (g1571) & (!g1572) & (g165) & (!g166)) + ((g1569) & (g1570) & (g1571) & (g1572) & (!g165) & (!g166)) + ((g1569) & (g1570) & (g1571) & (g1572) & (!g165) & (g166)) + ((g1569) & (g1570) & (g1571) & (g1572) & (g165) & (!g166)) + ((g1569) & (g1570) & (g1571) & (g1572) & (g165) & (g166)));
	assign g5007 = (((!g2177) & (!g2841) & (!sk[104]) & (g1574)) + ((!g2177) & (!g2841) & (sk[104]) & (g1574)) + ((!g2177) & (g2841) & (!sk[104]) & (!g1574)) + ((!g2177) & (g2841) & (!sk[104]) & (g1574)) + ((!g2177) & (g2841) & (sk[104]) & (g1574)) + ((g2177) & (!g2841) & (!sk[104]) & (g1574)) + ((g2177) & (g2841) & (!sk[104]) & (!g1574)) + ((g2177) & (g2841) & (!sk[104]) & (g1574)) + ((g2177) & (g2841) & (sk[104]) & (!g1574)) + ((g2177) & (g2841) & (sk[104]) & (g1574)));
	assign g5008 = (((!sk[105]) & (!g2178) & (!g2841) & (g1575)) + ((!sk[105]) & (!g2178) & (g2841) & (!g1575)) + ((!sk[105]) & (!g2178) & (g2841) & (g1575)) + ((!sk[105]) & (g2178) & (!g2841) & (g1575)) + ((!sk[105]) & (g2178) & (g2841) & (!g1575)) + ((!sk[105]) & (g2178) & (g2841) & (g1575)) + ((sk[105]) & (!g2178) & (!g2841) & (g1575)) + ((sk[105]) & (!g2178) & (g2841) & (g1575)) + ((sk[105]) & (g2178) & (g2841) & (!g1575)) + ((sk[105]) & (g2178) & (g2841) & (g1575)));
	assign g5009 = (((!sk[106]) & (!g2179) & (!g2841) & (g1576)) + ((!sk[106]) & (!g2179) & (g2841) & (!g1576)) + ((!sk[106]) & (!g2179) & (g2841) & (g1576)) + ((!sk[106]) & (g2179) & (!g2841) & (g1576)) + ((!sk[106]) & (g2179) & (g2841) & (!g1576)) + ((!sk[106]) & (g2179) & (g2841) & (g1576)) + ((sk[106]) & (!g2179) & (!g2841) & (g1576)) + ((sk[106]) & (!g2179) & (g2841) & (g1576)) + ((sk[106]) & (g2179) & (g2841) & (!g1576)) + ((sk[106]) & (g2179) & (g2841) & (g1576)));
	assign g1577 = (((!g165) & (!sk[107]) & (!g166) & (!g1574) & (g1575) & (!g1576)) + ((!g165) & (!sk[107]) & (!g166) & (!g1574) & (g1575) & (g1576)) + ((!g165) & (!sk[107]) & (!g166) & (g1574) & (!g1575) & (!g1576)) + ((!g165) & (!sk[107]) & (!g166) & (g1574) & (!g1575) & (g1576)) + ((!g165) & (!sk[107]) & (!g166) & (g1574) & (g1575) & (!g1576)) + ((!g165) & (!sk[107]) & (!g166) & (g1574) & (g1575) & (g1576)) + ((!g165) & (!sk[107]) & (g166) & (!g1574) & (!g1575) & (!g1576)) + ((!g165) & (!sk[107]) & (g166) & (!g1574) & (!g1575) & (g1576)) + ((!g165) & (!sk[107]) & (g166) & (!g1574) & (g1575) & (!g1576)) + ((!g165) & (!sk[107]) & (g166) & (!g1574) & (g1575) & (g1576)) + ((!g165) & (!sk[107]) & (g166) & (g1574) & (!g1575) & (!g1576)) + ((!g165) & (!sk[107]) & (g166) & (g1574) & (!g1575) & (g1576)) + ((!g165) & (!sk[107]) & (g166) & (g1574) & (g1575) & (!g1576)) + ((!g165) & (!sk[107]) & (g166) & (g1574) & (g1575) & (g1576)) + ((!g165) & (sk[107]) & (g166) & (!g1574) & (!g1575) & (g1576)) + ((!g165) & (sk[107]) & (g166) & (!g1574) & (g1575) & (g1576)) + ((!g165) & (sk[107]) & (g166) & (g1574) & (!g1575) & (g1576)) + ((!g165) & (sk[107]) & (g166) & (g1574) & (g1575) & (g1576)) + ((g165) & (!sk[107]) & (!g166) & (!g1574) & (g1575) & (!g1576)) + ((g165) & (!sk[107]) & (!g166) & (!g1574) & (g1575) & (g1576)) + ((g165) & (!sk[107]) & (!g166) & (g1574) & (!g1575) & (!g1576)) + ((g165) & (!sk[107]) & (!g166) & (g1574) & (!g1575) & (g1576)) + ((g165) & (!sk[107]) & (!g166) & (g1574) & (g1575) & (!g1576)) + ((g165) & (!sk[107]) & (!g166) & (g1574) & (g1575) & (g1576)) + ((g165) & (!sk[107]) & (g166) & (!g1574) & (!g1575) & (!g1576)) + ((g165) & (!sk[107]) & (g166) & (!g1574) & (!g1575) & (g1576)) + ((g165) & (!sk[107]) & (g166) & (!g1574) & (g1575) & (!g1576)) + ((g165) & (!sk[107]) & (g166) & (!g1574) & (g1575) & (g1576)) + ((g165) & (!sk[107]) & (g166) & (g1574) & (!g1575) & (!g1576)) + ((g165) & (!sk[107]) & (g166) & (g1574) & (!g1575) & (g1576)) + ((g165) & (!sk[107]) & (g166) & (g1574) & (g1575) & (!g1576)) + ((g165) & (!sk[107]) & (g166) & (g1574) & (g1575) & (g1576)) + ((g165) & (sk[107]) & (!g166) & (g1574) & (!g1575) & (!g1576)) + ((g165) & (sk[107]) & (!g166) & (g1574) & (!g1575) & (g1576)) + ((g165) & (sk[107]) & (!g166) & (g1574) & (g1575) & (!g1576)) + ((g165) & (sk[107]) & (!g166) & (g1574) & (g1575) & (g1576)) + ((g165) & (sk[107]) & (g166) & (!g1574) & (g1575) & (!g1576)) + ((g165) & (sk[107]) & (g166) & (!g1574) & (g1575) & (g1576)) + ((g165) & (sk[107]) & (g166) & (g1574) & (g1575) & (!g1576)) + ((g165) & (sk[107]) & (g166) & (g1574) & (g1575) & (g1576)));
	assign g5010 = (((!g2162) & (!sk[108]) & (!g2841) & (g1578)) + ((!g2162) & (!sk[108]) & (g2841) & (!g1578)) + ((!g2162) & (!sk[108]) & (g2841) & (g1578)) + ((!g2162) & (sk[108]) & (!g2841) & (g1578)) + ((!g2162) & (sk[108]) & (g2841) & (g1578)) + ((g2162) & (!sk[108]) & (!g2841) & (g1578)) + ((g2162) & (!sk[108]) & (g2841) & (!g1578)) + ((g2162) & (!sk[108]) & (g2841) & (g1578)) + ((g2162) & (sk[108]) & (g2841) & (!g1578)) + ((g2162) & (sk[108]) & (g2841) & (g1578)));
	assign g5011 = (((!g2164) & (!g2841) & (!sk[109]) & (g1579)) + ((!g2164) & (!g2841) & (sk[109]) & (g1579)) + ((!g2164) & (g2841) & (!sk[109]) & (!g1579)) + ((!g2164) & (g2841) & (!sk[109]) & (g1579)) + ((!g2164) & (g2841) & (sk[109]) & (g1579)) + ((g2164) & (!g2841) & (!sk[109]) & (g1579)) + ((g2164) & (g2841) & (!sk[109]) & (!g1579)) + ((g2164) & (g2841) & (!sk[109]) & (g1579)) + ((g2164) & (g2841) & (sk[109]) & (!g1579)) + ((g2164) & (g2841) & (sk[109]) & (g1579)));
	assign g5012 = (((!sk[110]) & (!g2166) & (!g2841) & (g1580)) + ((!sk[110]) & (!g2166) & (g2841) & (!g1580)) + ((!sk[110]) & (!g2166) & (g2841) & (g1580)) + ((!sk[110]) & (g2166) & (!g2841) & (g1580)) + ((!sk[110]) & (g2166) & (g2841) & (!g1580)) + ((!sk[110]) & (g2166) & (g2841) & (g1580)) + ((sk[110]) & (!g2166) & (!g2841) & (g1580)) + ((sk[110]) & (!g2166) & (g2841) & (g1580)) + ((sk[110]) & (g2166) & (g2841) & (!g1580)) + ((sk[110]) & (g2166) & (g2841) & (g1580)));
	assign g5013 = (((!g2168) & (!g2841) & (!sk[111]) & (g1581)) + ((!g2168) & (!g2841) & (sk[111]) & (g1581)) + ((!g2168) & (g2841) & (!sk[111]) & (!g1581)) + ((!g2168) & (g2841) & (!sk[111]) & (g1581)) + ((!g2168) & (g2841) & (sk[111]) & (g1581)) + ((g2168) & (!g2841) & (!sk[111]) & (g1581)) + ((g2168) & (g2841) & (!sk[111]) & (!g1581)) + ((g2168) & (g2841) & (!sk[111]) & (g1581)) + ((g2168) & (g2841) & (sk[111]) & (!g1581)) + ((g2168) & (g2841) & (sk[111]) & (g1581)));
	assign g1582 = (((!g1578) & (!g1579) & (!g1580) & (g1581) & (g165) & (g166)) + ((!g1578) & (!g1579) & (g1580) & (!g1581) & (!g165) & (g166)) + ((!g1578) & (!g1579) & (g1580) & (g1581) & (!g165) & (g166)) + ((!g1578) & (!g1579) & (g1580) & (g1581) & (g165) & (g166)) + ((!g1578) & (g1579) & (!g1580) & (!g1581) & (g165) & (!g166)) + ((!g1578) & (g1579) & (!g1580) & (g1581) & (g165) & (!g166)) + ((!g1578) & (g1579) & (!g1580) & (g1581) & (g165) & (g166)) + ((!g1578) & (g1579) & (g1580) & (!g1581) & (!g165) & (g166)) + ((!g1578) & (g1579) & (g1580) & (!g1581) & (g165) & (!g166)) + ((!g1578) & (g1579) & (g1580) & (g1581) & (!g165) & (g166)) + ((!g1578) & (g1579) & (g1580) & (g1581) & (g165) & (!g166)) + ((!g1578) & (g1579) & (g1580) & (g1581) & (g165) & (g166)) + ((g1578) & (!g1579) & (!g1580) & (!g1581) & (!g165) & (!g166)) + ((g1578) & (!g1579) & (!g1580) & (g1581) & (!g165) & (!g166)) + ((g1578) & (!g1579) & (!g1580) & (g1581) & (g165) & (g166)) + ((g1578) & (!g1579) & (g1580) & (!g1581) & (!g165) & (!g166)) + ((g1578) & (!g1579) & (g1580) & (!g1581) & (!g165) & (g166)) + ((g1578) & (!g1579) & (g1580) & (g1581) & (!g165) & (!g166)) + ((g1578) & (!g1579) & (g1580) & (g1581) & (!g165) & (g166)) + ((g1578) & (!g1579) & (g1580) & (g1581) & (g165) & (g166)) + ((g1578) & (g1579) & (!g1580) & (!g1581) & (!g165) & (!g166)) + ((g1578) & (g1579) & (!g1580) & (!g1581) & (g165) & (!g166)) + ((g1578) & (g1579) & (!g1580) & (g1581) & (!g165) & (!g166)) + ((g1578) & (g1579) & (!g1580) & (g1581) & (g165) & (!g166)) + ((g1578) & (g1579) & (!g1580) & (g1581) & (g165) & (g166)) + ((g1578) & (g1579) & (g1580) & (!g1581) & (!g165) & (!g166)) + ((g1578) & (g1579) & (g1580) & (!g1581) & (!g165) & (g166)) + ((g1578) & (g1579) & (g1580) & (!g1581) & (g165) & (!g166)) + ((g1578) & (g1579) & (g1580) & (g1581) & (!g165) & (!g166)) + ((g1578) & (g1579) & (g1580) & (g1581) & (!g165) & (g166)) + ((g1578) & (g1579) & (g1580) & (g1581) & (g165) & (!g166)) + ((g1578) & (g1579) & (g1580) & (g1581) & (g165) & (g166)));
	assign g5014 = (((!g2169) & (!g2841) & (!sk[113]) & (g1583)) + ((!g2169) & (!g2841) & (sk[113]) & (g1583)) + ((!g2169) & (g2841) & (!sk[113]) & (!g1583)) + ((!g2169) & (g2841) & (!sk[113]) & (g1583)) + ((!g2169) & (g2841) & (sk[113]) & (g1583)) + ((g2169) & (!g2841) & (!sk[113]) & (g1583)) + ((g2169) & (g2841) & (!sk[113]) & (!g1583)) + ((g2169) & (g2841) & (!sk[113]) & (g1583)) + ((g2169) & (g2841) & (sk[113]) & (!g1583)) + ((g2169) & (g2841) & (sk[113]) & (g1583)));
	assign g5015 = (((!g2170) & (!sk[114]) & (!g2841) & (g1584)) + ((!g2170) & (!sk[114]) & (g2841) & (!g1584)) + ((!g2170) & (!sk[114]) & (g2841) & (g1584)) + ((!g2170) & (sk[114]) & (!g2841) & (g1584)) + ((!g2170) & (sk[114]) & (g2841) & (g1584)) + ((g2170) & (!sk[114]) & (!g2841) & (g1584)) + ((g2170) & (!sk[114]) & (g2841) & (!g1584)) + ((g2170) & (!sk[114]) & (g2841) & (g1584)) + ((g2170) & (sk[114]) & (g2841) & (!g1584)) + ((g2170) & (sk[114]) & (g2841) & (g1584)));
	assign g5016 = (((!sk[115]) & (!g2171) & (!g2841) & (g1585)) + ((!sk[115]) & (!g2171) & (g2841) & (!g1585)) + ((!sk[115]) & (!g2171) & (g2841) & (g1585)) + ((!sk[115]) & (g2171) & (!g2841) & (g1585)) + ((!sk[115]) & (g2171) & (g2841) & (!g1585)) + ((!sk[115]) & (g2171) & (g2841) & (g1585)) + ((sk[115]) & (!g2171) & (!g2841) & (g1585)) + ((sk[115]) & (!g2171) & (g2841) & (g1585)) + ((sk[115]) & (g2171) & (g2841) & (!g1585)) + ((sk[115]) & (g2171) & (g2841) & (g1585)));
	assign g5017 = (((!sk[116]) & (!g2172) & (!g2841) & (g1586)) + ((!sk[116]) & (!g2172) & (g2841) & (!g1586)) + ((!sk[116]) & (!g2172) & (g2841) & (g1586)) + ((!sk[116]) & (g2172) & (!g2841) & (g1586)) + ((!sk[116]) & (g2172) & (g2841) & (!g1586)) + ((!sk[116]) & (g2172) & (g2841) & (g1586)) + ((sk[116]) & (!g2172) & (!g2841) & (g1586)) + ((sk[116]) & (!g2172) & (g2841) & (g1586)) + ((sk[116]) & (g2172) & (g2841) & (!g1586)) + ((sk[116]) & (g2172) & (g2841) & (g1586)));
	assign g1587 = (((!g1583) & (!g1584) & (!g1585) & (g1586) & (g165) & (g166)) + ((!g1583) & (!g1584) & (g1585) & (!g1586) & (!g165) & (g166)) + ((!g1583) & (!g1584) & (g1585) & (g1586) & (!g165) & (g166)) + ((!g1583) & (!g1584) & (g1585) & (g1586) & (g165) & (g166)) + ((!g1583) & (g1584) & (!g1585) & (!g1586) & (g165) & (!g166)) + ((!g1583) & (g1584) & (!g1585) & (g1586) & (g165) & (!g166)) + ((!g1583) & (g1584) & (!g1585) & (g1586) & (g165) & (g166)) + ((!g1583) & (g1584) & (g1585) & (!g1586) & (!g165) & (g166)) + ((!g1583) & (g1584) & (g1585) & (!g1586) & (g165) & (!g166)) + ((!g1583) & (g1584) & (g1585) & (g1586) & (!g165) & (g166)) + ((!g1583) & (g1584) & (g1585) & (g1586) & (g165) & (!g166)) + ((!g1583) & (g1584) & (g1585) & (g1586) & (g165) & (g166)) + ((g1583) & (!g1584) & (!g1585) & (!g1586) & (!g165) & (!g166)) + ((g1583) & (!g1584) & (!g1585) & (g1586) & (!g165) & (!g166)) + ((g1583) & (!g1584) & (!g1585) & (g1586) & (g165) & (g166)) + ((g1583) & (!g1584) & (g1585) & (!g1586) & (!g165) & (!g166)) + ((g1583) & (!g1584) & (g1585) & (!g1586) & (!g165) & (g166)) + ((g1583) & (!g1584) & (g1585) & (g1586) & (!g165) & (!g166)) + ((g1583) & (!g1584) & (g1585) & (g1586) & (!g165) & (g166)) + ((g1583) & (!g1584) & (g1585) & (g1586) & (g165) & (g166)) + ((g1583) & (g1584) & (!g1585) & (!g1586) & (!g165) & (!g166)) + ((g1583) & (g1584) & (!g1585) & (!g1586) & (g165) & (!g166)) + ((g1583) & (g1584) & (!g1585) & (g1586) & (!g165) & (!g166)) + ((g1583) & (g1584) & (!g1585) & (g1586) & (g165) & (!g166)) + ((g1583) & (g1584) & (!g1585) & (g1586) & (g165) & (g166)) + ((g1583) & (g1584) & (g1585) & (!g1586) & (!g165) & (!g166)) + ((g1583) & (g1584) & (g1585) & (!g1586) & (!g165) & (g166)) + ((g1583) & (g1584) & (g1585) & (!g1586) & (g165) & (!g166)) + ((g1583) & (g1584) & (g1585) & (g1586) & (!g165) & (!g166)) + ((g1583) & (g1584) & (g1585) & (g1586) & (!g165) & (g166)) + ((g1583) & (g1584) & (g1585) & (g1586) & (g165) & (!g166)) + ((g1583) & (g1584) & (g1585) & (g1586) & (g165) & (g166)));
	assign g1588 = (((!g147) & (!g148) & (!g1573) & (g1577) & (!g1582) & (!g1587)) + ((!g147) & (!g148) & (!g1573) & (g1577) & (!g1582) & (g1587)) + ((!g147) & (!g148) & (!g1573) & (g1577) & (g1582) & (!g1587)) + ((!g147) & (!g148) & (!g1573) & (g1577) & (g1582) & (g1587)) + ((!g147) & (!g148) & (g1573) & (g1577) & (!g1582) & (!g1587)) + ((!g147) & (!g148) & (g1573) & (g1577) & (!g1582) & (g1587)) + ((!g147) & (!g148) & (g1573) & (g1577) & (g1582) & (!g1587)) + ((!g147) & (!g148) & (g1573) & (g1577) & (g1582) & (g1587)) + ((!g147) & (g148) & (!g1573) & (!g1577) & (!g1582) & (g1587)) + ((!g147) & (g148) & (!g1573) & (!g1577) & (g1582) & (g1587)) + ((!g147) & (g148) & (!g1573) & (g1577) & (!g1582) & (g1587)) + ((!g147) & (g148) & (!g1573) & (g1577) & (g1582) & (g1587)) + ((!g147) & (g148) & (g1573) & (!g1577) & (!g1582) & (g1587)) + ((!g147) & (g148) & (g1573) & (!g1577) & (g1582) & (g1587)) + ((!g147) & (g148) & (g1573) & (g1577) & (!g1582) & (g1587)) + ((!g147) & (g148) & (g1573) & (g1577) & (g1582) & (g1587)) + ((g147) & (!g148) & (g1573) & (!g1577) & (!g1582) & (!g1587)) + ((g147) & (!g148) & (g1573) & (!g1577) & (!g1582) & (g1587)) + ((g147) & (!g148) & (g1573) & (!g1577) & (g1582) & (!g1587)) + ((g147) & (!g148) & (g1573) & (!g1577) & (g1582) & (g1587)) + ((g147) & (!g148) & (g1573) & (g1577) & (!g1582) & (!g1587)) + ((g147) & (!g148) & (g1573) & (g1577) & (!g1582) & (g1587)) + ((g147) & (!g148) & (g1573) & (g1577) & (g1582) & (!g1587)) + ((g147) & (!g148) & (g1573) & (g1577) & (g1582) & (g1587)) + ((g147) & (g148) & (!g1573) & (!g1577) & (g1582) & (!g1587)) + ((g147) & (g148) & (!g1573) & (!g1577) & (g1582) & (g1587)) + ((g147) & (g148) & (!g1573) & (g1577) & (g1582) & (!g1587)) + ((g147) & (g148) & (!g1573) & (g1577) & (g1582) & (g1587)) + ((g147) & (g148) & (g1573) & (!g1577) & (g1582) & (!g1587)) + ((g147) & (g148) & (g1573) & (!g1577) & (g1582) & (g1587)) + ((g147) & (g148) & (g1573) & (g1577) & (g1582) & (!g1587)) + ((g147) & (g148) & (g1573) & (g1577) & (g1582) & (g1587)));
	assign g1589 = (((!g142) & (!sk[119]) & (!g1568) & (g1588)) + ((!g142) & (!sk[119]) & (g1568) & (!g1588)) + ((!g142) & (!sk[119]) & (g1568) & (g1588)) + ((!g142) & (sk[119]) & (!g1568) & (g1588)) + ((!g142) & (sk[119]) & (g1568) & (g1588)) + ((g142) & (!sk[119]) & (!g1568) & (g1588)) + ((g142) & (!sk[119]) & (g1568) & (!g1588)) + ((g142) & (!sk[119]) & (g1568) & (g1588)) + ((g142) & (sk[119]) & (g1568) & (!g1588)) + ((g142) & (sk[119]) & (g1568) & (g1588)));
	assign g1590 = (((!g867) & (!sk[120]) & (!g107) & (!g679) & (g1589)) + ((!g867) & (!sk[120]) & (!g107) & (g679) & (!g1589)) + ((!g867) & (!sk[120]) & (!g107) & (g679) & (g1589)) + ((!g867) & (!sk[120]) & (g107) & (!g679) & (!g1589)) + ((!g867) & (!sk[120]) & (g107) & (!g679) & (g1589)) + ((!g867) & (!sk[120]) & (g107) & (g679) & (!g1589)) + ((!g867) & (!sk[120]) & (g107) & (g679) & (g1589)) + ((!g867) & (sk[120]) & (!g107) & (!g679) & (g1589)) + ((!g867) & (sk[120]) & (!g107) & (g679) & (g1589)) + ((!g867) & (sk[120]) & (g107) & (!g679) & (!g1589)) + ((!g867) & (sk[120]) & (g107) & (g679) & (g1589)) + ((g867) & (!sk[120]) & (!g107) & (!g679) & (g1589)) + ((g867) & (!sk[120]) & (!g107) & (g679) & (!g1589)) + ((g867) & (!sk[120]) & (!g107) & (g679) & (g1589)) + ((g867) & (!sk[120]) & (g107) & (!g679) & (!g1589)) + ((g867) & (!sk[120]) & (g107) & (!g679) & (g1589)) + ((g867) & (!sk[120]) & (g107) & (g679) & (!g1589)) + ((g867) & (!sk[120]) & (g107) & (g679) & (g1589)) + ((g867) & (sk[120]) & (!g107) & (!g679) & (g1589)) + ((g867) & (sk[120]) & (!g107) & (g679) & (!g1589)) + ((g867) & (sk[120]) & (g107) & (!g679) & (!g1589)) + ((g867) & (sk[120]) & (g107) & (g679) & (!g1589)));
	assign g1591 = (((!g126) & (!g1543) & (g1547) & (!g1545) & (!g916) & (!g1590)) + ((!g126) & (!g1543) & (g1547) & (!g1545) & (!g916) & (g1590)) + ((!g126) & (!g1543) & (g1547) & (!g1545) & (g916) & (!g1590)) + ((!g126) & (!g1543) & (g1547) & (!g1545) & (g916) & (g1590)) + ((!g126) & (!g1543) & (g1547) & (g1545) & (!g916) & (!g1590)) + ((!g126) & (!g1543) & (g1547) & (g1545) & (!g916) & (g1590)) + ((!g126) & (!g1543) & (g1547) & (g1545) & (g916) & (!g1590)) + ((!g126) & (!g1543) & (g1547) & (g1545) & (g916) & (g1590)) + ((!g126) & (g1543) & (g1547) & (!g1545) & (!g916) & (!g1590)) + ((!g126) & (g1543) & (g1547) & (!g1545) & (!g916) & (g1590)) + ((!g126) & (g1543) & (g1547) & (!g1545) & (g916) & (!g1590)) + ((!g126) & (g1543) & (g1547) & (!g1545) & (g916) & (g1590)) + ((!g126) & (g1543) & (g1547) & (g1545) & (!g916) & (!g1590)) + ((!g126) & (g1543) & (g1547) & (g1545) & (!g916) & (g1590)) + ((!g126) & (g1543) & (g1547) & (g1545) & (g916) & (!g1590)) + ((!g126) & (g1543) & (g1547) & (g1545) & (g916) & (g1590)) + ((g126) & (!g1543) & (!g1547) & (!g1545) & (!g916) & (g1590)) + ((g126) & (!g1543) & (!g1547) & (!g1545) & (g916) & (g1590)) + ((g126) & (!g1543) & (!g1547) & (g1545) & (!g916) & (!g1590)) + ((g126) & (!g1543) & (!g1547) & (g1545) & (g916) & (g1590)) + ((g126) & (!g1543) & (g1547) & (!g1545) & (!g916) & (g1590)) + ((g126) & (!g1543) & (g1547) & (!g1545) & (g916) & (g1590)) + ((g126) & (!g1543) & (g1547) & (g1545) & (!g916) & (!g1590)) + ((g126) & (!g1543) & (g1547) & (g1545) & (g916) & (g1590)) + ((g126) & (g1543) & (!g1547) & (!g1545) & (!g916) & (!g1590)) + ((g126) & (g1543) & (!g1547) & (!g1545) & (g916) & (g1590)) + ((g126) & (g1543) & (!g1547) & (g1545) & (!g916) & (!g1590)) + ((g126) & (g1543) & (!g1547) & (g1545) & (g916) & (!g1590)) + ((g126) & (g1543) & (g1547) & (!g1545) & (!g916) & (!g1590)) + ((g126) & (g1543) & (g1547) & (!g1545) & (g916) & (g1590)) + ((g126) & (g1543) & (g1547) & (g1545) & (!g916) & (!g1590)) + ((g126) & (g1543) & (g1547) & (g1545) & (g916) & (!g1590)));
	assign g1592 = (((!g79) & (!g80) & (!sk[122]) & (!g81) & (g131)) + ((!g79) & (!g80) & (!sk[122]) & (g81) & (!g131)) + ((!g79) & (!g80) & (!sk[122]) & (g81) & (g131)) + ((!g79) & (g80) & (!sk[122]) & (!g81) & (!g131)) + ((!g79) & (g80) & (!sk[122]) & (!g81) & (g131)) + ((!g79) & (g80) & (!sk[122]) & (g81) & (!g131)) + ((!g79) & (g80) & (!sk[122]) & (g81) & (g131)) + ((g79) & (!g80) & (!sk[122]) & (!g81) & (g131)) + ((g79) & (!g80) & (!sk[122]) & (g81) & (!g131)) + ((g79) & (!g80) & (!sk[122]) & (g81) & (g131)) + ((g79) & (g80) & (!sk[122]) & (!g81) & (!g131)) + ((g79) & (g80) & (!sk[122]) & (!g81) & (g131)) + ((g79) & (g80) & (!sk[122]) & (g81) & (!g131)) + ((g79) & (g80) & (!sk[122]) & (g81) & (g131)) + ((g79) & (g80) & (sk[122]) & (g81) & (g131)));
	assign g1593 = (((!sk[123]) & (g89) & (!g188)) + ((!sk[123]) & (g89) & (g188)) + ((sk[123]) & (!g89) & (g188)) + ((sk[123]) & (g89) & (!g188)));
	assign g1594 = (((!g143) & (!g144) & (!g145) & (g146) & (g820) & (g773)) + ((!g143) & (!g144) & (g145) & (!g146) & (!g820) & (g773)) + ((!g143) & (!g144) & (g145) & (g146) & (!g820) & (g773)) + ((!g143) & (!g144) & (g145) & (g146) & (g820) & (g773)) + ((!g143) & (g144) & (!g145) & (!g146) & (g820) & (!g773)) + ((!g143) & (g144) & (!g145) & (g146) & (g820) & (!g773)) + ((!g143) & (g144) & (!g145) & (g146) & (g820) & (g773)) + ((!g143) & (g144) & (g145) & (!g146) & (!g820) & (g773)) + ((!g143) & (g144) & (g145) & (!g146) & (g820) & (!g773)) + ((!g143) & (g144) & (g145) & (g146) & (!g820) & (g773)) + ((!g143) & (g144) & (g145) & (g146) & (g820) & (!g773)) + ((!g143) & (g144) & (g145) & (g146) & (g820) & (g773)) + ((g143) & (!g144) & (!g145) & (!g146) & (!g820) & (!g773)) + ((g143) & (!g144) & (!g145) & (g146) & (!g820) & (!g773)) + ((g143) & (!g144) & (!g145) & (g146) & (g820) & (g773)) + ((g143) & (!g144) & (g145) & (!g146) & (!g820) & (!g773)) + ((g143) & (!g144) & (g145) & (!g146) & (!g820) & (g773)) + ((g143) & (!g144) & (g145) & (g146) & (!g820) & (!g773)) + ((g143) & (!g144) & (g145) & (g146) & (!g820) & (g773)) + ((g143) & (!g144) & (g145) & (g146) & (g820) & (g773)) + ((g143) & (g144) & (!g145) & (!g146) & (!g820) & (!g773)) + ((g143) & (g144) & (!g145) & (!g146) & (g820) & (!g773)) + ((g143) & (g144) & (!g145) & (g146) & (!g820) & (!g773)) + ((g143) & (g144) & (!g145) & (g146) & (g820) & (!g773)) + ((g143) & (g144) & (!g145) & (g146) & (g820) & (g773)) + ((g143) & (g144) & (g145) & (!g146) & (!g820) & (!g773)) + ((g143) & (g144) & (g145) & (!g146) & (!g820) & (g773)) + ((g143) & (g144) & (g145) & (!g146) & (g820) & (!g773)) + ((g143) & (g144) & (g145) & (g146) & (!g820) & (!g773)) + ((g143) & (g144) & (g145) & (g146) & (!g820) & (g773)) + ((g143) & (g144) & (g145) & (g146) & (g820) & (!g773)) + ((g143) & (g144) & (g145) & (g146) & (g820) & (g773)));
	assign g1595 = (((!g150) & (!g151) & (!g152) & (g153) & (g820) & (g773)) + ((!g150) & (!g151) & (g152) & (!g153) & (!g820) & (g773)) + ((!g150) & (!g151) & (g152) & (g153) & (!g820) & (g773)) + ((!g150) & (!g151) & (g152) & (g153) & (g820) & (g773)) + ((!g150) & (g151) & (!g152) & (!g153) & (g820) & (!g773)) + ((!g150) & (g151) & (!g152) & (g153) & (g820) & (!g773)) + ((!g150) & (g151) & (!g152) & (g153) & (g820) & (g773)) + ((!g150) & (g151) & (g152) & (!g153) & (!g820) & (g773)) + ((!g150) & (g151) & (g152) & (!g153) & (g820) & (!g773)) + ((!g150) & (g151) & (g152) & (g153) & (!g820) & (g773)) + ((!g150) & (g151) & (g152) & (g153) & (g820) & (!g773)) + ((!g150) & (g151) & (g152) & (g153) & (g820) & (g773)) + ((g150) & (!g151) & (!g152) & (!g153) & (!g820) & (!g773)) + ((g150) & (!g151) & (!g152) & (g153) & (!g820) & (!g773)) + ((g150) & (!g151) & (!g152) & (g153) & (g820) & (g773)) + ((g150) & (!g151) & (g152) & (!g153) & (!g820) & (!g773)) + ((g150) & (!g151) & (g152) & (!g153) & (!g820) & (g773)) + ((g150) & (!g151) & (g152) & (g153) & (!g820) & (!g773)) + ((g150) & (!g151) & (g152) & (g153) & (!g820) & (g773)) + ((g150) & (!g151) & (g152) & (g153) & (g820) & (g773)) + ((g150) & (g151) & (!g152) & (!g153) & (!g820) & (!g773)) + ((g150) & (g151) & (!g152) & (!g153) & (g820) & (!g773)) + ((g150) & (g151) & (!g152) & (g153) & (!g820) & (!g773)) + ((g150) & (g151) & (!g152) & (g153) & (g820) & (!g773)) + ((g150) & (g151) & (!g152) & (g153) & (g820) & (g773)) + ((g150) & (g151) & (g152) & (!g153) & (!g820) & (!g773)) + ((g150) & (g151) & (g152) & (!g153) & (!g820) & (g773)) + ((g150) & (g151) & (g152) & (!g153) & (g820) & (!g773)) + ((g150) & (g151) & (g152) & (g153) & (!g820) & (!g773)) + ((g150) & (g151) & (g152) & (g153) & (!g820) & (g773)) + ((g150) & (g151) & (g152) & (g153) & (g820) & (!g773)) + ((g150) & (g151) & (g152) & (g153) & (g820) & (g773)));
	assign g1596 = (((!g155) & (!g156) & (!g157) & (g158) & (g820) & (g773)) + ((!g155) & (!g156) & (g157) & (!g158) & (!g820) & (g773)) + ((!g155) & (!g156) & (g157) & (g158) & (!g820) & (g773)) + ((!g155) & (!g156) & (g157) & (g158) & (g820) & (g773)) + ((!g155) & (g156) & (!g157) & (!g158) & (g820) & (!g773)) + ((!g155) & (g156) & (!g157) & (g158) & (g820) & (!g773)) + ((!g155) & (g156) & (!g157) & (g158) & (g820) & (g773)) + ((!g155) & (g156) & (g157) & (!g158) & (!g820) & (g773)) + ((!g155) & (g156) & (g157) & (!g158) & (g820) & (!g773)) + ((!g155) & (g156) & (g157) & (g158) & (!g820) & (g773)) + ((!g155) & (g156) & (g157) & (g158) & (g820) & (!g773)) + ((!g155) & (g156) & (g157) & (g158) & (g820) & (g773)) + ((g155) & (!g156) & (!g157) & (!g158) & (!g820) & (!g773)) + ((g155) & (!g156) & (!g157) & (g158) & (!g820) & (!g773)) + ((g155) & (!g156) & (!g157) & (g158) & (g820) & (g773)) + ((g155) & (!g156) & (g157) & (!g158) & (!g820) & (!g773)) + ((g155) & (!g156) & (g157) & (!g158) & (!g820) & (g773)) + ((g155) & (!g156) & (g157) & (g158) & (!g820) & (!g773)) + ((g155) & (!g156) & (g157) & (g158) & (!g820) & (g773)) + ((g155) & (!g156) & (g157) & (g158) & (g820) & (g773)) + ((g155) & (g156) & (!g157) & (!g158) & (!g820) & (!g773)) + ((g155) & (g156) & (!g157) & (!g158) & (g820) & (!g773)) + ((g155) & (g156) & (!g157) & (g158) & (!g820) & (!g773)) + ((g155) & (g156) & (!g157) & (g158) & (g820) & (!g773)) + ((g155) & (g156) & (!g157) & (g158) & (g820) & (g773)) + ((g155) & (g156) & (g157) & (!g158) & (!g820) & (!g773)) + ((g155) & (g156) & (g157) & (!g158) & (!g820) & (g773)) + ((g155) & (g156) & (g157) & (!g158) & (g820) & (!g773)) + ((g155) & (g156) & (g157) & (g158) & (!g820) & (!g773)) + ((g155) & (g156) & (g157) & (g158) & (!g820) & (g773)) + ((g155) & (g156) & (g157) & (g158) & (g820) & (!g773)) + ((g155) & (g156) & (g157) & (g158) & (g820) & (g773)));
	assign g1597 = (((!g160) & (!g161) & (!g162) & (g163) & (g820) & (g773)) + ((!g160) & (!g161) & (g162) & (!g163) & (!g820) & (g773)) + ((!g160) & (!g161) & (g162) & (g163) & (!g820) & (g773)) + ((!g160) & (!g161) & (g162) & (g163) & (g820) & (g773)) + ((!g160) & (g161) & (!g162) & (!g163) & (g820) & (!g773)) + ((!g160) & (g161) & (!g162) & (g163) & (g820) & (!g773)) + ((!g160) & (g161) & (!g162) & (g163) & (g820) & (g773)) + ((!g160) & (g161) & (g162) & (!g163) & (!g820) & (g773)) + ((!g160) & (g161) & (g162) & (!g163) & (g820) & (!g773)) + ((!g160) & (g161) & (g162) & (g163) & (!g820) & (g773)) + ((!g160) & (g161) & (g162) & (g163) & (g820) & (!g773)) + ((!g160) & (g161) & (g162) & (g163) & (g820) & (g773)) + ((g160) & (!g161) & (!g162) & (!g163) & (!g820) & (!g773)) + ((g160) & (!g161) & (!g162) & (g163) & (!g820) & (!g773)) + ((g160) & (!g161) & (!g162) & (g163) & (g820) & (g773)) + ((g160) & (!g161) & (g162) & (!g163) & (!g820) & (!g773)) + ((g160) & (!g161) & (g162) & (!g163) & (!g820) & (g773)) + ((g160) & (!g161) & (g162) & (g163) & (!g820) & (!g773)) + ((g160) & (!g161) & (g162) & (g163) & (!g820) & (g773)) + ((g160) & (!g161) & (g162) & (g163) & (g820) & (g773)) + ((g160) & (g161) & (!g162) & (!g163) & (!g820) & (!g773)) + ((g160) & (g161) & (!g162) & (!g163) & (g820) & (!g773)) + ((g160) & (g161) & (!g162) & (g163) & (!g820) & (!g773)) + ((g160) & (g161) & (!g162) & (g163) & (g820) & (!g773)) + ((g160) & (g161) & (!g162) & (g163) & (g820) & (g773)) + ((g160) & (g161) & (g162) & (!g163) & (!g820) & (!g773)) + ((g160) & (g161) & (g162) & (!g163) & (!g820) & (g773)) + ((g160) & (g161) & (g162) & (!g163) & (g820) & (!g773)) + ((g160) & (g161) & (g162) & (g163) & (!g820) & (!g773)) + ((g160) & (g161) & (g162) & (g163) & (!g820) & (g773)) + ((g160) & (g161) & (g162) & (g163) & (g820) & (!g773)) + ((g160) & (g161) & (g162) & (g163) & (g820) & (g773)));
	assign g1598 = (((!g1594) & (!g1595) & (!g1596) & (g1597) & (g677) & (g726)) + ((!g1594) & (!g1595) & (g1596) & (!g1597) & (!g677) & (g726)) + ((!g1594) & (!g1595) & (g1596) & (g1597) & (!g677) & (g726)) + ((!g1594) & (!g1595) & (g1596) & (g1597) & (g677) & (g726)) + ((!g1594) & (g1595) & (!g1596) & (!g1597) & (g677) & (!g726)) + ((!g1594) & (g1595) & (!g1596) & (g1597) & (g677) & (!g726)) + ((!g1594) & (g1595) & (!g1596) & (g1597) & (g677) & (g726)) + ((!g1594) & (g1595) & (g1596) & (!g1597) & (!g677) & (g726)) + ((!g1594) & (g1595) & (g1596) & (!g1597) & (g677) & (!g726)) + ((!g1594) & (g1595) & (g1596) & (g1597) & (!g677) & (g726)) + ((!g1594) & (g1595) & (g1596) & (g1597) & (g677) & (!g726)) + ((!g1594) & (g1595) & (g1596) & (g1597) & (g677) & (g726)) + ((g1594) & (!g1595) & (!g1596) & (!g1597) & (!g677) & (!g726)) + ((g1594) & (!g1595) & (!g1596) & (g1597) & (!g677) & (!g726)) + ((g1594) & (!g1595) & (!g1596) & (g1597) & (g677) & (g726)) + ((g1594) & (!g1595) & (g1596) & (!g1597) & (!g677) & (!g726)) + ((g1594) & (!g1595) & (g1596) & (!g1597) & (!g677) & (g726)) + ((g1594) & (!g1595) & (g1596) & (g1597) & (!g677) & (!g726)) + ((g1594) & (!g1595) & (g1596) & (g1597) & (!g677) & (g726)) + ((g1594) & (!g1595) & (g1596) & (g1597) & (g677) & (g726)) + ((g1594) & (g1595) & (!g1596) & (!g1597) & (!g677) & (!g726)) + ((g1594) & (g1595) & (!g1596) & (!g1597) & (g677) & (!g726)) + ((g1594) & (g1595) & (!g1596) & (g1597) & (!g677) & (!g726)) + ((g1594) & (g1595) & (!g1596) & (g1597) & (g677) & (!g726)) + ((g1594) & (g1595) & (!g1596) & (g1597) & (g677) & (g726)) + ((g1594) & (g1595) & (g1596) & (!g1597) & (!g677) & (!g726)) + ((g1594) & (g1595) & (g1596) & (!g1597) & (!g677) & (g726)) + ((g1594) & (g1595) & (g1596) & (!g1597) & (g677) & (!g726)) + ((g1594) & (g1595) & (g1596) & (g1597) & (!g677) & (!g726)) + ((g1594) & (g1595) & (g1596) & (g1597) & (!g677) & (g726)) + ((g1594) & (g1595) & (g1596) & (g1597) & (g677) & (!g726)) + ((g1594) & (g1595) & (g1596) & (g1597) & (g677) & (g726)));
	assign g1599 = (((!g178) & (!g179) & (!g180) & (g181) & (g677) & (g726)) + ((!g178) & (!g179) & (g180) & (!g181) & (!g677) & (g726)) + ((!g178) & (!g179) & (g180) & (g181) & (!g677) & (g726)) + ((!g178) & (!g179) & (g180) & (g181) & (g677) & (g726)) + ((!g178) & (g179) & (!g180) & (!g181) & (g677) & (!g726)) + ((!g178) & (g179) & (!g180) & (g181) & (g677) & (!g726)) + ((!g178) & (g179) & (!g180) & (g181) & (g677) & (g726)) + ((!g178) & (g179) & (g180) & (!g181) & (!g677) & (g726)) + ((!g178) & (g179) & (g180) & (!g181) & (g677) & (!g726)) + ((!g178) & (g179) & (g180) & (g181) & (!g677) & (g726)) + ((!g178) & (g179) & (g180) & (g181) & (g677) & (!g726)) + ((!g178) & (g179) & (g180) & (g181) & (g677) & (g726)) + ((g178) & (!g179) & (!g180) & (!g181) & (!g677) & (!g726)) + ((g178) & (!g179) & (!g180) & (g181) & (!g677) & (!g726)) + ((g178) & (!g179) & (!g180) & (g181) & (g677) & (g726)) + ((g178) & (!g179) & (g180) & (!g181) & (!g677) & (!g726)) + ((g178) & (!g179) & (g180) & (!g181) & (!g677) & (g726)) + ((g178) & (!g179) & (g180) & (g181) & (!g677) & (!g726)) + ((g178) & (!g179) & (g180) & (g181) & (!g677) & (g726)) + ((g178) & (!g179) & (g180) & (g181) & (g677) & (g726)) + ((g178) & (g179) & (!g180) & (!g181) & (!g677) & (!g726)) + ((g178) & (g179) & (!g180) & (!g181) & (g677) & (!g726)) + ((g178) & (g179) & (!g180) & (g181) & (!g677) & (!g726)) + ((g178) & (g179) & (!g180) & (g181) & (g677) & (!g726)) + ((g178) & (g179) & (!g180) & (g181) & (g677) & (g726)) + ((g178) & (g179) & (g180) & (!g181) & (!g677) & (!g726)) + ((g178) & (g179) & (g180) & (!g181) & (!g677) & (g726)) + ((g178) & (g179) & (g180) & (!g181) & (g677) & (!g726)) + ((g178) & (g179) & (g180) & (g181) & (!g677) & (!g726)) + ((g178) & (g179) & (g180) & (g181) & (!g677) & (g726)) + ((g178) & (g179) & (g180) & (g181) & (g677) & (!g726)) + ((g178) & (g179) & (g180) & (g181) & (g677) & (g726)));
	assign g1600 = (((!sk[2]) & (!g183) & (!g184) & (!g185) & (g677) & (!g726)) + ((!sk[2]) & (!g183) & (!g184) & (!g185) & (g677) & (g726)) + ((!sk[2]) & (!g183) & (!g184) & (g185) & (!g677) & (!g726)) + ((!sk[2]) & (!g183) & (!g184) & (g185) & (!g677) & (g726)) + ((!sk[2]) & (!g183) & (!g184) & (g185) & (g677) & (!g726)) + ((!sk[2]) & (!g183) & (!g184) & (g185) & (g677) & (g726)) + ((!sk[2]) & (!g183) & (g184) & (!g185) & (!g677) & (!g726)) + ((!sk[2]) & (!g183) & (g184) & (!g185) & (!g677) & (g726)) + ((!sk[2]) & (!g183) & (g184) & (!g185) & (g677) & (!g726)) + ((!sk[2]) & (!g183) & (g184) & (!g185) & (g677) & (g726)) + ((!sk[2]) & (!g183) & (g184) & (g185) & (!g677) & (!g726)) + ((!sk[2]) & (!g183) & (g184) & (g185) & (!g677) & (g726)) + ((!sk[2]) & (!g183) & (g184) & (g185) & (g677) & (!g726)) + ((!sk[2]) & (!g183) & (g184) & (g185) & (g677) & (g726)) + ((!sk[2]) & (g183) & (!g184) & (!g185) & (g677) & (!g726)) + ((!sk[2]) & (g183) & (!g184) & (!g185) & (g677) & (g726)) + ((!sk[2]) & (g183) & (!g184) & (g185) & (!g677) & (!g726)) + ((!sk[2]) & (g183) & (!g184) & (g185) & (!g677) & (g726)) + ((!sk[2]) & (g183) & (!g184) & (g185) & (g677) & (!g726)) + ((!sk[2]) & (g183) & (!g184) & (g185) & (g677) & (g726)) + ((!sk[2]) & (g183) & (g184) & (!g185) & (!g677) & (!g726)) + ((!sk[2]) & (g183) & (g184) & (!g185) & (!g677) & (g726)) + ((!sk[2]) & (g183) & (g184) & (!g185) & (g677) & (!g726)) + ((!sk[2]) & (g183) & (g184) & (!g185) & (g677) & (g726)) + ((!sk[2]) & (g183) & (g184) & (g185) & (!g677) & (!g726)) + ((!sk[2]) & (g183) & (g184) & (g185) & (!g677) & (g726)) + ((!sk[2]) & (g183) & (g184) & (g185) & (g677) & (!g726)) + ((!sk[2]) & (g183) & (g184) & (g185) & (g677) & (g726)) + ((sk[2]) & (!g183) & (!g184) & (g185) & (!g677) & (g726)) + ((sk[2]) & (!g183) & (g184) & (!g185) & (g677) & (g726)) + ((sk[2]) & (!g183) & (g184) & (g185) & (!g677) & (g726)) + ((sk[2]) & (!g183) & (g184) & (g185) & (g677) & (g726)) + ((sk[2]) & (g183) & (!g184) & (!g185) & (g677) & (!g726)) + ((sk[2]) & (g183) & (!g184) & (g185) & (!g677) & (g726)) + ((sk[2]) & (g183) & (!g184) & (g185) & (g677) & (!g726)) + ((sk[2]) & (g183) & (g184) & (!g185) & (g677) & (!g726)) + ((sk[2]) & (g183) & (g184) & (!g185) & (g677) & (g726)) + ((sk[2]) & (g183) & (g184) & (g185) & (!g677) & (g726)) + ((sk[2]) & (g183) & (g184) & (g185) & (g677) & (!g726)) + ((sk[2]) & (g183) & (g184) & (g185) & (g677) & (g726)));
	assign g1601 = (((!g168) & (!g169) & (!g170) & (g171) & (g677) & (g726)) + ((!g168) & (!g169) & (g170) & (!g171) & (!g677) & (g726)) + ((!g168) & (!g169) & (g170) & (g171) & (!g677) & (g726)) + ((!g168) & (!g169) & (g170) & (g171) & (g677) & (g726)) + ((!g168) & (g169) & (!g170) & (!g171) & (g677) & (!g726)) + ((!g168) & (g169) & (!g170) & (g171) & (g677) & (!g726)) + ((!g168) & (g169) & (!g170) & (g171) & (g677) & (g726)) + ((!g168) & (g169) & (g170) & (!g171) & (!g677) & (g726)) + ((!g168) & (g169) & (g170) & (!g171) & (g677) & (!g726)) + ((!g168) & (g169) & (g170) & (g171) & (!g677) & (g726)) + ((!g168) & (g169) & (g170) & (g171) & (g677) & (!g726)) + ((!g168) & (g169) & (g170) & (g171) & (g677) & (g726)) + ((g168) & (!g169) & (!g170) & (!g171) & (!g677) & (!g726)) + ((g168) & (!g169) & (!g170) & (g171) & (!g677) & (!g726)) + ((g168) & (!g169) & (!g170) & (g171) & (g677) & (g726)) + ((g168) & (!g169) & (g170) & (!g171) & (!g677) & (!g726)) + ((g168) & (!g169) & (g170) & (!g171) & (!g677) & (g726)) + ((g168) & (!g169) & (g170) & (g171) & (!g677) & (!g726)) + ((g168) & (!g169) & (g170) & (g171) & (!g677) & (g726)) + ((g168) & (!g169) & (g170) & (g171) & (g677) & (g726)) + ((g168) & (g169) & (!g170) & (!g171) & (!g677) & (!g726)) + ((g168) & (g169) & (!g170) & (!g171) & (g677) & (!g726)) + ((g168) & (g169) & (!g170) & (g171) & (!g677) & (!g726)) + ((g168) & (g169) & (!g170) & (g171) & (g677) & (!g726)) + ((g168) & (g169) & (!g170) & (g171) & (g677) & (g726)) + ((g168) & (g169) & (g170) & (!g171) & (!g677) & (!g726)) + ((g168) & (g169) & (g170) & (!g171) & (!g677) & (g726)) + ((g168) & (g169) & (g170) & (!g171) & (g677) & (!g726)) + ((g168) & (g169) & (g170) & (g171) & (!g677) & (!g726)) + ((g168) & (g169) & (g170) & (g171) & (!g677) & (g726)) + ((g168) & (g169) & (g170) & (g171) & (g677) & (!g726)) + ((g168) & (g169) & (g170) & (g171) & (g677) & (g726)));
	assign g1602 = (((!g173) & (!g174) & (!g175) & (g176) & (g677) & (g726)) + ((!g173) & (!g174) & (g175) & (!g176) & (!g677) & (g726)) + ((!g173) & (!g174) & (g175) & (g176) & (!g677) & (g726)) + ((!g173) & (!g174) & (g175) & (g176) & (g677) & (g726)) + ((!g173) & (g174) & (!g175) & (!g176) & (g677) & (!g726)) + ((!g173) & (g174) & (!g175) & (g176) & (g677) & (!g726)) + ((!g173) & (g174) & (!g175) & (g176) & (g677) & (g726)) + ((!g173) & (g174) & (g175) & (!g176) & (!g677) & (g726)) + ((!g173) & (g174) & (g175) & (!g176) & (g677) & (!g726)) + ((!g173) & (g174) & (g175) & (g176) & (!g677) & (g726)) + ((!g173) & (g174) & (g175) & (g176) & (g677) & (!g726)) + ((!g173) & (g174) & (g175) & (g176) & (g677) & (g726)) + ((g173) & (!g174) & (!g175) & (!g176) & (!g677) & (!g726)) + ((g173) & (!g174) & (!g175) & (g176) & (!g677) & (!g726)) + ((g173) & (!g174) & (!g175) & (g176) & (g677) & (g726)) + ((g173) & (!g174) & (g175) & (!g176) & (!g677) & (!g726)) + ((g173) & (!g174) & (g175) & (!g176) & (!g677) & (g726)) + ((g173) & (!g174) & (g175) & (g176) & (!g677) & (!g726)) + ((g173) & (!g174) & (g175) & (g176) & (!g677) & (g726)) + ((g173) & (!g174) & (g175) & (g176) & (g677) & (g726)) + ((g173) & (g174) & (!g175) & (!g176) & (!g677) & (!g726)) + ((g173) & (g174) & (!g175) & (!g176) & (g677) & (!g726)) + ((g173) & (g174) & (!g175) & (g176) & (!g677) & (!g726)) + ((g173) & (g174) & (!g175) & (g176) & (g677) & (!g726)) + ((g173) & (g174) & (!g175) & (g176) & (g677) & (g726)) + ((g173) & (g174) & (g175) & (!g176) & (!g677) & (!g726)) + ((g173) & (g174) & (g175) & (!g176) & (!g677) & (g726)) + ((g173) & (g174) & (g175) & (!g176) & (g677) & (!g726)) + ((g173) & (g174) & (g175) & (g176) & (!g677) & (!g726)) + ((g173) & (g174) & (g175) & (g176) & (!g677) & (g726)) + ((g173) & (g174) & (g175) & (g176) & (g677) & (!g726)) + ((g173) & (g174) & (g175) & (g176) & (g677) & (g726)));
	assign g1603 = (((!g820) & (!g773) & (!g1599) & (g1600) & (!g1601) & (!g1602)) + ((!g820) & (!g773) & (!g1599) & (g1600) & (!g1601) & (g1602)) + ((!g820) & (!g773) & (!g1599) & (g1600) & (g1601) & (!g1602)) + ((!g820) & (!g773) & (!g1599) & (g1600) & (g1601) & (g1602)) + ((!g820) & (!g773) & (g1599) & (g1600) & (!g1601) & (!g1602)) + ((!g820) & (!g773) & (g1599) & (g1600) & (!g1601) & (g1602)) + ((!g820) & (!g773) & (g1599) & (g1600) & (g1601) & (!g1602)) + ((!g820) & (!g773) & (g1599) & (g1600) & (g1601) & (g1602)) + ((!g820) & (g773) & (!g1599) & (!g1600) & (!g1601) & (g1602)) + ((!g820) & (g773) & (!g1599) & (!g1600) & (g1601) & (g1602)) + ((!g820) & (g773) & (!g1599) & (g1600) & (!g1601) & (g1602)) + ((!g820) & (g773) & (!g1599) & (g1600) & (g1601) & (g1602)) + ((!g820) & (g773) & (g1599) & (!g1600) & (!g1601) & (g1602)) + ((!g820) & (g773) & (g1599) & (!g1600) & (g1601) & (g1602)) + ((!g820) & (g773) & (g1599) & (g1600) & (!g1601) & (g1602)) + ((!g820) & (g773) & (g1599) & (g1600) & (g1601) & (g1602)) + ((g820) & (!g773) & (g1599) & (!g1600) & (!g1601) & (!g1602)) + ((g820) & (!g773) & (g1599) & (!g1600) & (!g1601) & (g1602)) + ((g820) & (!g773) & (g1599) & (!g1600) & (g1601) & (!g1602)) + ((g820) & (!g773) & (g1599) & (!g1600) & (g1601) & (g1602)) + ((g820) & (!g773) & (g1599) & (g1600) & (!g1601) & (!g1602)) + ((g820) & (!g773) & (g1599) & (g1600) & (!g1601) & (g1602)) + ((g820) & (!g773) & (g1599) & (g1600) & (g1601) & (!g1602)) + ((g820) & (!g773) & (g1599) & (g1600) & (g1601) & (g1602)) + ((g820) & (g773) & (!g1599) & (!g1600) & (g1601) & (!g1602)) + ((g820) & (g773) & (!g1599) & (!g1600) & (g1601) & (g1602)) + ((g820) & (g773) & (!g1599) & (g1600) & (g1601) & (!g1602)) + ((g820) & (g773) & (!g1599) & (g1600) & (g1601) & (g1602)) + ((g820) & (g773) & (g1599) & (!g1600) & (g1601) & (!g1602)) + ((g820) & (g773) & (g1599) & (!g1600) & (g1601) & (g1602)) + ((g820) & (g773) & (g1599) & (g1600) & (g1601) & (!g1602)) + ((g820) & (g773) & (g1599) & (g1600) & (g1601) & (g1602)));
	assign g1604 = (((!g867) & (!g1598) & (!sk[6]) & (g1603)) + ((!g867) & (!g1598) & (sk[6]) & (g1603)) + ((!g867) & (g1598) & (!sk[6]) & (!g1603)) + ((!g867) & (g1598) & (!sk[6]) & (g1603)) + ((!g867) & (g1598) & (sk[6]) & (g1603)) + ((g867) & (!g1598) & (!sk[6]) & (g1603)) + ((g867) & (g1598) & (!sk[6]) & (!g1603)) + ((g867) & (g1598) & (!sk[6]) & (g1603)) + ((g867) & (g1598) & (sk[6]) & (!g1603)) + ((g867) & (g1598) & (sk[6]) & (g1603)));
	assign g1605 = (((!sk[7]) & (!g88) & (!g89) & (!g188) & (g230)) + ((!sk[7]) & (!g88) & (!g89) & (g188) & (!g230)) + ((!sk[7]) & (!g88) & (!g89) & (g188) & (g230)) + ((!sk[7]) & (!g88) & (g89) & (!g188) & (!g230)) + ((!sk[7]) & (!g88) & (g89) & (!g188) & (g230)) + ((!sk[7]) & (!g88) & (g89) & (g188) & (!g230)) + ((!sk[7]) & (!g88) & (g89) & (g188) & (g230)) + ((!sk[7]) & (g88) & (!g89) & (!g188) & (g230)) + ((!sk[7]) & (g88) & (!g89) & (g188) & (!g230)) + ((!sk[7]) & (g88) & (!g89) & (g188) & (g230)) + ((!sk[7]) & (g88) & (g89) & (!g188) & (!g230)) + ((!sk[7]) & (g88) & (g89) & (!g188) & (g230)) + ((!sk[7]) & (g88) & (g89) & (g188) & (!g230)) + ((!sk[7]) & (g88) & (g89) & (g188) & (g230)) + ((sk[7]) & (!g88) & (!g89) & (!g188) & (g230)) + ((sk[7]) & (!g88) & (!g89) & (g188) & (g230)) + ((sk[7]) & (!g88) & (g89) & (!g188) & (g230)) + ((sk[7]) & (!g88) & (g89) & (g188) & (!g230)) + ((sk[7]) & (g88) & (!g89) & (!g188) & (!g230)) + ((sk[7]) & (g88) & (!g89) & (g188) & (!g230)) + ((sk[7]) & (g88) & (g89) & (!g188) & (!g230)) + ((sk[7]) & (g88) & (g89) & (g188) & (g230)));
	assign g1606 = (((!g79) & (!sk[8]) & (!g80) & (!g81) & (g133)) + ((!g79) & (!sk[8]) & (!g80) & (g81) & (!g133)) + ((!g79) & (!sk[8]) & (!g80) & (g81) & (g133)) + ((!g79) & (!sk[8]) & (g80) & (!g81) & (!g133)) + ((!g79) & (!sk[8]) & (g80) & (!g81) & (g133)) + ((!g79) & (!sk[8]) & (g80) & (g81) & (!g133)) + ((!g79) & (!sk[8]) & (g80) & (g81) & (g133)) + ((g79) & (!sk[8]) & (!g80) & (!g81) & (g133)) + ((g79) & (!sk[8]) & (!g80) & (g81) & (!g133)) + ((g79) & (!sk[8]) & (!g80) & (g81) & (g133)) + ((g79) & (!sk[8]) & (g80) & (!g81) & (!g133)) + ((g79) & (!sk[8]) & (g80) & (!g81) & (g133)) + ((g79) & (!sk[8]) & (g80) & (g81) & (!g133)) + ((g79) & (!sk[8]) & (g80) & (g81) & (g133)) + ((g79) & (sk[8]) & (g80) & (g81) & (g133)));
	assign g1607 = (((!g1606) & (!sk[9]) & (!g136) & (!g1593) & (g1605)) + ((!g1606) & (!sk[9]) & (!g136) & (g1593) & (!g1605)) + ((!g1606) & (!sk[9]) & (!g136) & (g1593) & (g1605)) + ((!g1606) & (!sk[9]) & (g136) & (!g1593) & (!g1605)) + ((!g1606) & (!sk[9]) & (g136) & (!g1593) & (g1605)) + ((!g1606) & (!sk[9]) & (g136) & (g1593) & (!g1605)) + ((!g1606) & (!sk[9]) & (g136) & (g1593) & (g1605)) + ((!g1606) & (sk[9]) & (!g136) & (!g1593) & (!g1605)) + ((!g1606) & (sk[9]) & (!g136) & (!g1593) & (g1605)) + ((!g1606) & (sk[9]) & (!g136) & (g1593) & (!g1605)) + ((!g1606) & (sk[9]) & (!g136) & (g1593) & (g1605)) + ((g1606) & (!sk[9]) & (!g136) & (!g1593) & (g1605)) + ((g1606) & (!sk[9]) & (!g136) & (g1593) & (!g1605)) + ((g1606) & (!sk[9]) & (!g136) & (g1593) & (g1605)) + ((g1606) & (!sk[9]) & (g136) & (!g1593) & (!g1605)) + ((g1606) & (!sk[9]) & (g136) & (!g1593) & (g1605)) + ((g1606) & (!sk[9]) & (g136) & (g1593) & (!g1605)) + ((g1606) & (!sk[9]) & (g136) & (g1593) & (g1605)) + ((g1606) & (sk[9]) & (!g136) & (g1593) & (g1605)));
	assign g1608 = (((!g1592) & (!g35) & (!g1593) & (g1604) & (!g1605) & (g1607)) + ((!g1592) & (!g35) & (!g1593) & (g1604) & (g1605) & (g1607)) + ((!g1592) & (!g35) & (g1593) & (g1604) & (!g1605) & (g1607)) + ((!g1592) & (!g35) & (g1593) & (g1604) & (g1605) & (g1607)) + ((!g1592) & (g35) & (!g1593) & (g1604) & (!g1605) & (g1607)) + ((!g1592) & (g35) & (!g1593) & (g1604) & (g1605) & (g1607)) + ((!g1592) & (g35) & (g1593) & (g1604) & (!g1605) & (g1607)) + ((!g1592) & (g35) & (g1593) & (g1604) & (g1605) & (g1607)) + ((g1592) & (!g35) & (!g1593) & (g1604) & (g1605) & (g1607)) + ((g1592) & (g35) & (!g1593) & (g1604) & (g1605) & (g1607)) + ((g1592) & (g35) & (g1593) & (!g1604) & (!g1605) & (g1607)) + ((g1592) & (g35) & (g1593) & (!g1604) & (g1605) & (g1607)) + ((g1592) & (g35) & (g1593) & (g1604) & (!g1605) & (g1607)) + ((g1592) & (g35) & (g1593) & (g1604) & (g1605) & (g1607)));
	assign g1609 = (((!g137) & (sk[11]) & (g126)) + ((g137) & (!sk[11]) & (!g126)) + ((g137) & (!sk[11]) & (g126)));
	assign g1610 = (((!g189) & (!g194) & (!g199) & (g204) & (g820) & (g773)) + ((!g189) & (!g194) & (g199) & (!g204) & (!g820) & (g773)) + ((!g189) & (!g194) & (g199) & (g204) & (!g820) & (g773)) + ((!g189) & (!g194) & (g199) & (g204) & (g820) & (g773)) + ((!g189) & (g194) & (!g199) & (!g204) & (g820) & (!g773)) + ((!g189) & (g194) & (!g199) & (g204) & (g820) & (!g773)) + ((!g189) & (g194) & (!g199) & (g204) & (g820) & (g773)) + ((!g189) & (g194) & (g199) & (!g204) & (!g820) & (g773)) + ((!g189) & (g194) & (g199) & (!g204) & (g820) & (!g773)) + ((!g189) & (g194) & (g199) & (g204) & (!g820) & (g773)) + ((!g189) & (g194) & (g199) & (g204) & (g820) & (!g773)) + ((!g189) & (g194) & (g199) & (g204) & (g820) & (g773)) + ((g189) & (!g194) & (!g199) & (!g204) & (!g820) & (!g773)) + ((g189) & (!g194) & (!g199) & (g204) & (!g820) & (!g773)) + ((g189) & (!g194) & (!g199) & (g204) & (g820) & (g773)) + ((g189) & (!g194) & (g199) & (!g204) & (!g820) & (!g773)) + ((g189) & (!g194) & (g199) & (!g204) & (!g820) & (g773)) + ((g189) & (!g194) & (g199) & (g204) & (!g820) & (!g773)) + ((g189) & (!g194) & (g199) & (g204) & (!g820) & (g773)) + ((g189) & (!g194) & (g199) & (g204) & (g820) & (g773)) + ((g189) & (g194) & (!g199) & (!g204) & (!g820) & (!g773)) + ((g189) & (g194) & (!g199) & (!g204) & (g820) & (!g773)) + ((g189) & (g194) & (!g199) & (g204) & (!g820) & (!g773)) + ((g189) & (g194) & (!g199) & (g204) & (g820) & (!g773)) + ((g189) & (g194) & (!g199) & (g204) & (g820) & (g773)) + ((g189) & (g194) & (g199) & (!g204) & (!g820) & (!g773)) + ((g189) & (g194) & (g199) & (!g204) & (!g820) & (g773)) + ((g189) & (g194) & (g199) & (!g204) & (g820) & (!g773)) + ((g189) & (g194) & (g199) & (g204) & (!g820) & (!g773)) + ((g189) & (g194) & (g199) & (g204) & (!g820) & (g773)) + ((g189) & (g194) & (g199) & (g204) & (g820) & (!g773)) + ((g189) & (g194) & (g199) & (g204) & (g820) & (g773)));
	assign g1611 = (((!g190) & (!g195) & (!g200) & (g205) & (g820) & (g773)) + ((!g190) & (!g195) & (g200) & (!g205) & (!g820) & (g773)) + ((!g190) & (!g195) & (g200) & (g205) & (!g820) & (g773)) + ((!g190) & (!g195) & (g200) & (g205) & (g820) & (g773)) + ((!g190) & (g195) & (!g200) & (!g205) & (g820) & (!g773)) + ((!g190) & (g195) & (!g200) & (g205) & (g820) & (!g773)) + ((!g190) & (g195) & (!g200) & (g205) & (g820) & (g773)) + ((!g190) & (g195) & (g200) & (!g205) & (!g820) & (g773)) + ((!g190) & (g195) & (g200) & (!g205) & (g820) & (!g773)) + ((!g190) & (g195) & (g200) & (g205) & (!g820) & (g773)) + ((!g190) & (g195) & (g200) & (g205) & (g820) & (!g773)) + ((!g190) & (g195) & (g200) & (g205) & (g820) & (g773)) + ((g190) & (!g195) & (!g200) & (!g205) & (!g820) & (!g773)) + ((g190) & (!g195) & (!g200) & (g205) & (!g820) & (!g773)) + ((g190) & (!g195) & (!g200) & (g205) & (g820) & (g773)) + ((g190) & (!g195) & (g200) & (!g205) & (!g820) & (!g773)) + ((g190) & (!g195) & (g200) & (!g205) & (!g820) & (g773)) + ((g190) & (!g195) & (g200) & (g205) & (!g820) & (!g773)) + ((g190) & (!g195) & (g200) & (g205) & (!g820) & (g773)) + ((g190) & (!g195) & (g200) & (g205) & (g820) & (g773)) + ((g190) & (g195) & (!g200) & (!g205) & (!g820) & (!g773)) + ((g190) & (g195) & (!g200) & (!g205) & (g820) & (!g773)) + ((g190) & (g195) & (!g200) & (g205) & (!g820) & (!g773)) + ((g190) & (g195) & (!g200) & (g205) & (g820) & (!g773)) + ((g190) & (g195) & (!g200) & (g205) & (g820) & (g773)) + ((g190) & (g195) & (g200) & (!g205) & (!g820) & (!g773)) + ((g190) & (g195) & (g200) & (!g205) & (!g820) & (g773)) + ((g190) & (g195) & (g200) & (!g205) & (g820) & (!g773)) + ((g190) & (g195) & (g200) & (g205) & (!g820) & (!g773)) + ((g190) & (g195) & (g200) & (g205) & (!g820) & (g773)) + ((g190) & (g195) & (g200) & (g205) & (g820) & (!g773)) + ((g190) & (g195) & (g200) & (g205) & (g820) & (g773)));
	assign g1612 = (((!g191) & (!g196) & (!g201) & (g206) & (g820) & (g773)) + ((!g191) & (!g196) & (g201) & (!g206) & (!g820) & (g773)) + ((!g191) & (!g196) & (g201) & (g206) & (!g820) & (g773)) + ((!g191) & (!g196) & (g201) & (g206) & (g820) & (g773)) + ((!g191) & (g196) & (!g201) & (!g206) & (g820) & (!g773)) + ((!g191) & (g196) & (!g201) & (g206) & (g820) & (!g773)) + ((!g191) & (g196) & (!g201) & (g206) & (g820) & (g773)) + ((!g191) & (g196) & (g201) & (!g206) & (!g820) & (g773)) + ((!g191) & (g196) & (g201) & (!g206) & (g820) & (!g773)) + ((!g191) & (g196) & (g201) & (g206) & (!g820) & (g773)) + ((!g191) & (g196) & (g201) & (g206) & (g820) & (!g773)) + ((!g191) & (g196) & (g201) & (g206) & (g820) & (g773)) + ((g191) & (!g196) & (!g201) & (!g206) & (!g820) & (!g773)) + ((g191) & (!g196) & (!g201) & (g206) & (!g820) & (!g773)) + ((g191) & (!g196) & (!g201) & (g206) & (g820) & (g773)) + ((g191) & (!g196) & (g201) & (!g206) & (!g820) & (!g773)) + ((g191) & (!g196) & (g201) & (!g206) & (!g820) & (g773)) + ((g191) & (!g196) & (g201) & (g206) & (!g820) & (!g773)) + ((g191) & (!g196) & (g201) & (g206) & (!g820) & (g773)) + ((g191) & (!g196) & (g201) & (g206) & (g820) & (g773)) + ((g191) & (g196) & (!g201) & (!g206) & (!g820) & (!g773)) + ((g191) & (g196) & (!g201) & (!g206) & (g820) & (!g773)) + ((g191) & (g196) & (!g201) & (g206) & (!g820) & (!g773)) + ((g191) & (g196) & (!g201) & (g206) & (g820) & (!g773)) + ((g191) & (g196) & (!g201) & (g206) & (g820) & (g773)) + ((g191) & (g196) & (g201) & (!g206) & (!g820) & (!g773)) + ((g191) & (g196) & (g201) & (!g206) & (!g820) & (g773)) + ((g191) & (g196) & (g201) & (!g206) & (g820) & (!g773)) + ((g191) & (g196) & (g201) & (g206) & (!g820) & (!g773)) + ((g191) & (g196) & (g201) & (g206) & (!g820) & (g773)) + ((g191) & (g196) & (g201) & (g206) & (g820) & (!g773)) + ((g191) & (g196) & (g201) & (g206) & (g820) & (g773)));
	assign g1613 = (((!g192) & (!g197) & (!g202) & (g207) & (g820) & (g773)) + ((!g192) & (!g197) & (g202) & (!g207) & (!g820) & (g773)) + ((!g192) & (!g197) & (g202) & (g207) & (!g820) & (g773)) + ((!g192) & (!g197) & (g202) & (g207) & (g820) & (g773)) + ((!g192) & (g197) & (!g202) & (!g207) & (g820) & (!g773)) + ((!g192) & (g197) & (!g202) & (g207) & (g820) & (!g773)) + ((!g192) & (g197) & (!g202) & (g207) & (g820) & (g773)) + ((!g192) & (g197) & (g202) & (!g207) & (!g820) & (g773)) + ((!g192) & (g197) & (g202) & (!g207) & (g820) & (!g773)) + ((!g192) & (g197) & (g202) & (g207) & (!g820) & (g773)) + ((!g192) & (g197) & (g202) & (g207) & (g820) & (!g773)) + ((!g192) & (g197) & (g202) & (g207) & (g820) & (g773)) + ((g192) & (!g197) & (!g202) & (!g207) & (!g820) & (!g773)) + ((g192) & (!g197) & (!g202) & (g207) & (!g820) & (!g773)) + ((g192) & (!g197) & (!g202) & (g207) & (g820) & (g773)) + ((g192) & (!g197) & (g202) & (!g207) & (!g820) & (!g773)) + ((g192) & (!g197) & (g202) & (!g207) & (!g820) & (g773)) + ((g192) & (!g197) & (g202) & (g207) & (!g820) & (!g773)) + ((g192) & (!g197) & (g202) & (g207) & (!g820) & (g773)) + ((g192) & (!g197) & (g202) & (g207) & (g820) & (g773)) + ((g192) & (g197) & (!g202) & (!g207) & (!g820) & (!g773)) + ((g192) & (g197) & (!g202) & (!g207) & (g820) & (!g773)) + ((g192) & (g197) & (!g202) & (g207) & (!g820) & (!g773)) + ((g192) & (g197) & (!g202) & (g207) & (g820) & (!g773)) + ((g192) & (g197) & (!g202) & (g207) & (g820) & (g773)) + ((g192) & (g197) & (g202) & (!g207) & (!g820) & (!g773)) + ((g192) & (g197) & (g202) & (!g207) & (!g820) & (g773)) + ((g192) & (g197) & (g202) & (!g207) & (g820) & (!g773)) + ((g192) & (g197) & (g202) & (g207) & (!g820) & (!g773)) + ((g192) & (g197) & (g202) & (g207) & (!g820) & (g773)) + ((g192) & (g197) & (g202) & (g207) & (g820) & (!g773)) + ((g192) & (g197) & (g202) & (g207) & (g820) & (g773)));
	assign g1614 = (((!g1610) & (!g1611) & (!g1612) & (g1613) & (g677) & (g726)) + ((!g1610) & (!g1611) & (g1612) & (!g1613) & (!g677) & (g726)) + ((!g1610) & (!g1611) & (g1612) & (g1613) & (!g677) & (g726)) + ((!g1610) & (!g1611) & (g1612) & (g1613) & (g677) & (g726)) + ((!g1610) & (g1611) & (!g1612) & (!g1613) & (g677) & (!g726)) + ((!g1610) & (g1611) & (!g1612) & (g1613) & (g677) & (!g726)) + ((!g1610) & (g1611) & (!g1612) & (g1613) & (g677) & (g726)) + ((!g1610) & (g1611) & (g1612) & (!g1613) & (!g677) & (g726)) + ((!g1610) & (g1611) & (g1612) & (!g1613) & (g677) & (!g726)) + ((!g1610) & (g1611) & (g1612) & (g1613) & (!g677) & (g726)) + ((!g1610) & (g1611) & (g1612) & (g1613) & (g677) & (!g726)) + ((!g1610) & (g1611) & (g1612) & (g1613) & (g677) & (g726)) + ((g1610) & (!g1611) & (!g1612) & (!g1613) & (!g677) & (!g726)) + ((g1610) & (!g1611) & (!g1612) & (g1613) & (!g677) & (!g726)) + ((g1610) & (!g1611) & (!g1612) & (g1613) & (g677) & (g726)) + ((g1610) & (!g1611) & (g1612) & (!g1613) & (!g677) & (!g726)) + ((g1610) & (!g1611) & (g1612) & (!g1613) & (!g677) & (g726)) + ((g1610) & (!g1611) & (g1612) & (g1613) & (!g677) & (!g726)) + ((g1610) & (!g1611) & (g1612) & (g1613) & (!g677) & (g726)) + ((g1610) & (!g1611) & (g1612) & (g1613) & (g677) & (g726)) + ((g1610) & (g1611) & (!g1612) & (!g1613) & (!g677) & (!g726)) + ((g1610) & (g1611) & (!g1612) & (!g1613) & (g677) & (!g726)) + ((g1610) & (g1611) & (!g1612) & (g1613) & (!g677) & (!g726)) + ((g1610) & (g1611) & (!g1612) & (g1613) & (g677) & (!g726)) + ((g1610) & (g1611) & (!g1612) & (g1613) & (g677) & (g726)) + ((g1610) & (g1611) & (g1612) & (!g1613) & (!g677) & (!g726)) + ((g1610) & (g1611) & (g1612) & (!g1613) & (!g677) & (g726)) + ((g1610) & (g1611) & (g1612) & (!g1613) & (g677) & (!g726)) + ((g1610) & (g1611) & (g1612) & (g1613) & (!g677) & (!g726)) + ((g1610) & (g1611) & (g1612) & (g1613) & (!g677) & (g726)) + ((g1610) & (g1611) & (g1612) & (g1613) & (g677) & (!g726)) + ((g1610) & (g1611) & (g1612) & (g1613) & (g677) & (g726)));
	assign g1615 = (((!g220) & (!g221) & (!g222) & (g223) & (g677) & (g726)) + ((!g220) & (!g221) & (g222) & (!g223) & (!g677) & (g726)) + ((!g220) & (!g221) & (g222) & (g223) & (!g677) & (g726)) + ((!g220) & (!g221) & (g222) & (g223) & (g677) & (g726)) + ((!g220) & (g221) & (!g222) & (!g223) & (g677) & (!g726)) + ((!g220) & (g221) & (!g222) & (g223) & (g677) & (!g726)) + ((!g220) & (g221) & (!g222) & (g223) & (g677) & (g726)) + ((!g220) & (g221) & (g222) & (!g223) & (!g677) & (g726)) + ((!g220) & (g221) & (g222) & (!g223) & (g677) & (!g726)) + ((!g220) & (g221) & (g222) & (g223) & (!g677) & (g726)) + ((!g220) & (g221) & (g222) & (g223) & (g677) & (!g726)) + ((!g220) & (g221) & (g222) & (g223) & (g677) & (g726)) + ((g220) & (!g221) & (!g222) & (!g223) & (!g677) & (!g726)) + ((g220) & (!g221) & (!g222) & (g223) & (!g677) & (!g726)) + ((g220) & (!g221) & (!g222) & (g223) & (g677) & (g726)) + ((g220) & (!g221) & (g222) & (!g223) & (!g677) & (!g726)) + ((g220) & (!g221) & (g222) & (!g223) & (!g677) & (g726)) + ((g220) & (!g221) & (g222) & (g223) & (!g677) & (!g726)) + ((g220) & (!g221) & (g222) & (g223) & (!g677) & (g726)) + ((g220) & (!g221) & (g222) & (g223) & (g677) & (g726)) + ((g220) & (g221) & (!g222) & (!g223) & (!g677) & (!g726)) + ((g220) & (g221) & (!g222) & (!g223) & (g677) & (!g726)) + ((g220) & (g221) & (!g222) & (g223) & (!g677) & (!g726)) + ((g220) & (g221) & (!g222) & (g223) & (g677) & (!g726)) + ((g220) & (g221) & (!g222) & (g223) & (g677) & (g726)) + ((g220) & (g221) & (g222) & (!g223) & (!g677) & (!g726)) + ((g220) & (g221) & (g222) & (!g223) & (!g677) & (g726)) + ((g220) & (g221) & (g222) & (!g223) & (g677) & (!g726)) + ((g220) & (g221) & (g222) & (g223) & (!g677) & (!g726)) + ((g220) & (g221) & (g222) & (g223) & (!g677) & (g726)) + ((g220) & (g221) & (g222) & (g223) & (g677) & (!g726)) + ((g220) & (g221) & (g222) & (g223) & (g677) & (g726)));
	assign g1616 = (((!g677) & (!g726) & (!sk[18]) & (!g225) & (g226) & (!g227)) + ((!g677) & (!g726) & (!sk[18]) & (!g225) & (g226) & (g227)) + ((!g677) & (!g726) & (!sk[18]) & (g225) & (!g226) & (!g227)) + ((!g677) & (!g726) & (!sk[18]) & (g225) & (!g226) & (g227)) + ((!g677) & (!g726) & (!sk[18]) & (g225) & (g226) & (!g227)) + ((!g677) & (!g726) & (!sk[18]) & (g225) & (g226) & (g227)) + ((!g677) & (g726) & (!sk[18]) & (!g225) & (!g226) & (!g227)) + ((!g677) & (g726) & (!sk[18]) & (!g225) & (!g226) & (g227)) + ((!g677) & (g726) & (!sk[18]) & (!g225) & (g226) & (!g227)) + ((!g677) & (g726) & (!sk[18]) & (!g225) & (g226) & (g227)) + ((!g677) & (g726) & (!sk[18]) & (g225) & (!g226) & (!g227)) + ((!g677) & (g726) & (!sk[18]) & (g225) & (!g226) & (g227)) + ((!g677) & (g726) & (!sk[18]) & (g225) & (g226) & (!g227)) + ((!g677) & (g726) & (!sk[18]) & (g225) & (g226) & (g227)) + ((!g677) & (g726) & (sk[18]) & (!g225) & (!g226) & (g227)) + ((!g677) & (g726) & (sk[18]) & (!g225) & (g226) & (g227)) + ((!g677) & (g726) & (sk[18]) & (g225) & (!g226) & (g227)) + ((!g677) & (g726) & (sk[18]) & (g225) & (g226) & (g227)) + ((g677) & (!g726) & (!sk[18]) & (!g225) & (g226) & (!g227)) + ((g677) & (!g726) & (!sk[18]) & (!g225) & (g226) & (g227)) + ((g677) & (!g726) & (!sk[18]) & (g225) & (!g226) & (!g227)) + ((g677) & (!g726) & (!sk[18]) & (g225) & (!g226) & (g227)) + ((g677) & (!g726) & (!sk[18]) & (g225) & (g226) & (!g227)) + ((g677) & (!g726) & (!sk[18]) & (g225) & (g226) & (g227)) + ((g677) & (!g726) & (sk[18]) & (g225) & (!g226) & (!g227)) + ((g677) & (!g726) & (sk[18]) & (g225) & (!g226) & (g227)) + ((g677) & (!g726) & (sk[18]) & (g225) & (g226) & (!g227)) + ((g677) & (!g726) & (sk[18]) & (g225) & (g226) & (g227)) + ((g677) & (g726) & (!sk[18]) & (!g225) & (!g226) & (!g227)) + ((g677) & (g726) & (!sk[18]) & (!g225) & (!g226) & (g227)) + ((g677) & (g726) & (!sk[18]) & (!g225) & (g226) & (!g227)) + ((g677) & (g726) & (!sk[18]) & (!g225) & (g226) & (g227)) + ((g677) & (g726) & (!sk[18]) & (g225) & (!g226) & (!g227)) + ((g677) & (g726) & (!sk[18]) & (g225) & (!g226) & (g227)) + ((g677) & (g726) & (!sk[18]) & (g225) & (g226) & (!g227)) + ((g677) & (g726) & (!sk[18]) & (g225) & (g226) & (g227)) + ((g677) & (g726) & (sk[18]) & (!g225) & (g226) & (!g227)) + ((g677) & (g726) & (sk[18]) & (!g225) & (g226) & (g227)) + ((g677) & (g726) & (sk[18]) & (g225) & (g226) & (!g227)) + ((g677) & (g726) & (sk[18]) & (g225) & (g226) & (g227)));
	assign g1617 = (((!g210) & (!g211) & (!g212) & (g213) & (g677) & (g726)) + ((!g210) & (!g211) & (g212) & (!g213) & (!g677) & (g726)) + ((!g210) & (!g211) & (g212) & (g213) & (!g677) & (g726)) + ((!g210) & (!g211) & (g212) & (g213) & (g677) & (g726)) + ((!g210) & (g211) & (!g212) & (!g213) & (g677) & (!g726)) + ((!g210) & (g211) & (!g212) & (g213) & (g677) & (!g726)) + ((!g210) & (g211) & (!g212) & (g213) & (g677) & (g726)) + ((!g210) & (g211) & (g212) & (!g213) & (!g677) & (g726)) + ((!g210) & (g211) & (g212) & (!g213) & (g677) & (!g726)) + ((!g210) & (g211) & (g212) & (g213) & (!g677) & (g726)) + ((!g210) & (g211) & (g212) & (g213) & (g677) & (!g726)) + ((!g210) & (g211) & (g212) & (g213) & (g677) & (g726)) + ((g210) & (!g211) & (!g212) & (!g213) & (!g677) & (!g726)) + ((g210) & (!g211) & (!g212) & (g213) & (!g677) & (!g726)) + ((g210) & (!g211) & (!g212) & (g213) & (g677) & (g726)) + ((g210) & (!g211) & (g212) & (!g213) & (!g677) & (!g726)) + ((g210) & (!g211) & (g212) & (!g213) & (!g677) & (g726)) + ((g210) & (!g211) & (g212) & (g213) & (!g677) & (!g726)) + ((g210) & (!g211) & (g212) & (g213) & (!g677) & (g726)) + ((g210) & (!g211) & (g212) & (g213) & (g677) & (g726)) + ((g210) & (g211) & (!g212) & (!g213) & (!g677) & (!g726)) + ((g210) & (g211) & (!g212) & (!g213) & (g677) & (!g726)) + ((g210) & (g211) & (!g212) & (g213) & (!g677) & (!g726)) + ((g210) & (g211) & (!g212) & (g213) & (g677) & (!g726)) + ((g210) & (g211) & (!g212) & (g213) & (g677) & (g726)) + ((g210) & (g211) & (g212) & (!g213) & (!g677) & (!g726)) + ((g210) & (g211) & (g212) & (!g213) & (!g677) & (g726)) + ((g210) & (g211) & (g212) & (!g213) & (g677) & (!g726)) + ((g210) & (g211) & (g212) & (g213) & (!g677) & (!g726)) + ((g210) & (g211) & (g212) & (g213) & (!g677) & (g726)) + ((g210) & (g211) & (g212) & (g213) & (g677) & (!g726)) + ((g210) & (g211) & (g212) & (g213) & (g677) & (g726)));
	assign g1618 = (((!g215) & (!g216) & (!g217) & (g218) & (g677) & (g726)) + ((!g215) & (!g216) & (g217) & (!g218) & (!g677) & (g726)) + ((!g215) & (!g216) & (g217) & (g218) & (!g677) & (g726)) + ((!g215) & (!g216) & (g217) & (g218) & (g677) & (g726)) + ((!g215) & (g216) & (!g217) & (!g218) & (g677) & (!g726)) + ((!g215) & (g216) & (!g217) & (g218) & (g677) & (!g726)) + ((!g215) & (g216) & (!g217) & (g218) & (g677) & (g726)) + ((!g215) & (g216) & (g217) & (!g218) & (!g677) & (g726)) + ((!g215) & (g216) & (g217) & (!g218) & (g677) & (!g726)) + ((!g215) & (g216) & (g217) & (g218) & (!g677) & (g726)) + ((!g215) & (g216) & (g217) & (g218) & (g677) & (!g726)) + ((!g215) & (g216) & (g217) & (g218) & (g677) & (g726)) + ((g215) & (!g216) & (!g217) & (!g218) & (!g677) & (!g726)) + ((g215) & (!g216) & (!g217) & (g218) & (!g677) & (!g726)) + ((g215) & (!g216) & (!g217) & (g218) & (g677) & (g726)) + ((g215) & (!g216) & (g217) & (!g218) & (!g677) & (!g726)) + ((g215) & (!g216) & (g217) & (!g218) & (!g677) & (g726)) + ((g215) & (!g216) & (g217) & (g218) & (!g677) & (!g726)) + ((g215) & (!g216) & (g217) & (g218) & (!g677) & (g726)) + ((g215) & (!g216) & (g217) & (g218) & (g677) & (g726)) + ((g215) & (g216) & (!g217) & (!g218) & (!g677) & (!g726)) + ((g215) & (g216) & (!g217) & (!g218) & (g677) & (!g726)) + ((g215) & (g216) & (!g217) & (g218) & (!g677) & (!g726)) + ((g215) & (g216) & (!g217) & (g218) & (g677) & (!g726)) + ((g215) & (g216) & (!g217) & (g218) & (g677) & (g726)) + ((g215) & (g216) & (g217) & (!g218) & (!g677) & (!g726)) + ((g215) & (g216) & (g217) & (!g218) & (!g677) & (g726)) + ((g215) & (g216) & (g217) & (!g218) & (g677) & (!g726)) + ((g215) & (g216) & (g217) & (g218) & (!g677) & (!g726)) + ((g215) & (g216) & (g217) & (g218) & (!g677) & (g726)) + ((g215) & (g216) & (g217) & (g218) & (g677) & (!g726)) + ((g215) & (g216) & (g217) & (g218) & (g677) & (g726)));
	assign g1619 = (((!g820) & (!g773) & (!g1615) & (g1616) & (!g1617) & (!g1618)) + ((!g820) & (!g773) & (!g1615) & (g1616) & (!g1617) & (g1618)) + ((!g820) & (!g773) & (!g1615) & (g1616) & (g1617) & (!g1618)) + ((!g820) & (!g773) & (!g1615) & (g1616) & (g1617) & (g1618)) + ((!g820) & (!g773) & (g1615) & (g1616) & (!g1617) & (!g1618)) + ((!g820) & (!g773) & (g1615) & (g1616) & (!g1617) & (g1618)) + ((!g820) & (!g773) & (g1615) & (g1616) & (g1617) & (!g1618)) + ((!g820) & (!g773) & (g1615) & (g1616) & (g1617) & (g1618)) + ((!g820) & (g773) & (!g1615) & (!g1616) & (!g1617) & (g1618)) + ((!g820) & (g773) & (!g1615) & (!g1616) & (g1617) & (g1618)) + ((!g820) & (g773) & (!g1615) & (g1616) & (!g1617) & (g1618)) + ((!g820) & (g773) & (!g1615) & (g1616) & (g1617) & (g1618)) + ((!g820) & (g773) & (g1615) & (!g1616) & (!g1617) & (g1618)) + ((!g820) & (g773) & (g1615) & (!g1616) & (g1617) & (g1618)) + ((!g820) & (g773) & (g1615) & (g1616) & (!g1617) & (g1618)) + ((!g820) & (g773) & (g1615) & (g1616) & (g1617) & (g1618)) + ((g820) & (!g773) & (g1615) & (!g1616) & (!g1617) & (!g1618)) + ((g820) & (!g773) & (g1615) & (!g1616) & (!g1617) & (g1618)) + ((g820) & (!g773) & (g1615) & (!g1616) & (g1617) & (!g1618)) + ((g820) & (!g773) & (g1615) & (!g1616) & (g1617) & (g1618)) + ((g820) & (!g773) & (g1615) & (g1616) & (!g1617) & (!g1618)) + ((g820) & (!g773) & (g1615) & (g1616) & (!g1617) & (g1618)) + ((g820) & (!g773) & (g1615) & (g1616) & (g1617) & (!g1618)) + ((g820) & (!g773) & (g1615) & (g1616) & (g1617) & (g1618)) + ((g820) & (g773) & (!g1615) & (!g1616) & (g1617) & (!g1618)) + ((g820) & (g773) & (!g1615) & (!g1616) & (g1617) & (g1618)) + ((g820) & (g773) & (!g1615) & (g1616) & (g1617) & (!g1618)) + ((g820) & (g773) & (!g1615) & (g1616) & (g1617) & (g1618)) + ((g820) & (g773) & (g1615) & (!g1616) & (g1617) & (!g1618)) + ((g820) & (g773) & (g1615) & (!g1616) & (g1617) & (g1618)) + ((g820) & (g773) & (g1615) & (g1616) & (g1617) & (!g1618)) + ((g820) & (g773) & (g1615) & (g1616) & (g1617) & (g1618)));
	assign g1620 = (((!sk[22]) & (!g867) & (!g1614) & (g1619)) + ((!sk[22]) & (!g867) & (g1614) & (!g1619)) + ((!sk[22]) & (!g867) & (g1614) & (g1619)) + ((!sk[22]) & (g867) & (!g1614) & (g1619)) + ((!sk[22]) & (g867) & (g1614) & (!g1619)) + ((!sk[22]) & (g867) & (g1614) & (g1619)) + ((sk[22]) & (!g867) & (!g1614) & (g1619)) + ((sk[22]) & (!g867) & (g1614) & (g1619)) + ((sk[22]) & (g867) & (g1614) & (!g1619)) + ((sk[22]) & (g867) & (g1614) & (g1619)));
	assign g1621 = (((!g1592) & (!g1593) & (!g1605) & (g1607) & (!g36) & (g1620)) + ((!g1592) & (!g1593) & (!g1605) & (g1607) & (g36) & (g1620)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (!g36) & (g1620)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (g36) & (g1620)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (!g36) & (g1620)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (g36) & (g1620)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (!g36) & (g1620)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (g36) & (g1620)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (!g36) & (g1620)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (g36) & (g1620)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g36) & (!g1620)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g36) & (g1620)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g36) & (!g1620)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g36) & (g1620)));
	assign g1622 = (((!g232) & (!g233) & (!g234) & (g235) & (g820) & (g773)) + ((!g232) & (!g233) & (g234) & (!g235) & (!g820) & (g773)) + ((!g232) & (!g233) & (g234) & (g235) & (!g820) & (g773)) + ((!g232) & (!g233) & (g234) & (g235) & (g820) & (g773)) + ((!g232) & (g233) & (!g234) & (!g235) & (g820) & (!g773)) + ((!g232) & (g233) & (!g234) & (g235) & (g820) & (!g773)) + ((!g232) & (g233) & (!g234) & (g235) & (g820) & (g773)) + ((!g232) & (g233) & (g234) & (!g235) & (!g820) & (g773)) + ((!g232) & (g233) & (g234) & (!g235) & (g820) & (!g773)) + ((!g232) & (g233) & (g234) & (g235) & (!g820) & (g773)) + ((!g232) & (g233) & (g234) & (g235) & (g820) & (!g773)) + ((!g232) & (g233) & (g234) & (g235) & (g820) & (g773)) + ((g232) & (!g233) & (!g234) & (!g235) & (!g820) & (!g773)) + ((g232) & (!g233) & (!g234) & (g235) & (!g820) & (!g773)) + ((g232) & (!g233) & (!g234) & (g235) & (g820) & (g773)) + ((g232) & (!g233) & (g234) & (!g235) & (!g820) & (!g773)) + ((g232) & (!g233) & (g234) & (!g235) & (!g820) & (g773)) + ((g232) & (!g233) & (g234) & (g235) & (!g820) & (!g773)) + ((g232) & (!g233) & (g234) & (g235) & (!g820) & (g773)) + ((g232) & (!g233) & (g234) & (g235) & (g820) & (g773)) + ((g232) & (g233) & (!g234) & (!g235) & (!g820) & (!g773)) + ((g232) & (g233) & (!g234) & (!g235) & (g820) & (!g773)) + ((g232) & (g233) & (!g234) & (g235) & (!g820) & (!g773)) + ((g232) & (g233) & (!g234) & (g235) & (g820) & (!g773)) + ((g232) & (g233) & (!g234) & (g235) & (g820) & (g773)) + ((g232) & (g233) & (g234) & (!g235) & (!g820) & (!g773)) + ((g232) & (g233) & (g234) & (!g235) & (!g820) & (g773)) + ((g232) & (g233) & (g234) & (!g235) & (g820) & (!g773)) + ((g232) & (g233) & (g234) & (g235) & (!g820) & (!g773)) + ((g232) & (g233) & (g234) & (g235) & (!g820) & (g773)) + ((g232) & (g233) & (g234) & (g235) & (g820) & (!g773)) + ((g232) & (g233) & (g234) & (g235) & (g820) & (g773)));
	assign g1623 = (((!g237) & (!g238) & (!g239) & (g240) & (g820) & (g773)) + ((!g237) & (!g238) & (g239) & (!g240) & (!g820) & (g773)) + ((!g237) & (!g238) & (g239) & (g240) & (!g820) & (g773)) + ((!g237) & (!g238) & (g239) & (g240) & (g820) & (g773)) + ((!g237) & (g238) & (!g239) & (!g240) & (g820) & (!g773)) + ((!g237) & (g238) & (!g239) & (g240) & (g820) & (!g773)) + ((!g237) & (g238) & (!g239) & (g240) & (g820) & (g773)) + ((!g237) & (g238) & (g239) & (!g240) & (!g820) & (g773)) + ((!g237) & (g238) & (g239) & (!g240) & (g820) & (!g773)) + ((!g237) & (g238) & (g239) & (g240) & (!g820) & (g773)) + ((!g237) & (g238) & (g239) & (g240) & (g820) & (!g773)) + ((!g237) & (g238) & (g239) & (g240) & (g820) & (g773)) + ((g237) & (!g238) & (!g239) & (!g240) & (!g820) & (!g773)) + ((g237) & (!g238) & (!g239) & (g240) & (!g820) & (!g773)) + ((g237) & (!g238) & (!g239) & (g240) & (g820) & (g773)) + ((g237) & (!g238) & (g239) & (!g240) & (!g820) & (!g773)) + ((g237) & (!g238) & (g239) & (!g240) & (!g820) & (g773)) + ((g237) & (!g238) & (g239) & (g240) & (!g820) & (!g773)) + ((g237) & (!g238) & (g239) & (g240) & (!g820) & (g773)) + ((g237) & (!g238) & (g239) & (g240) & (g820) & (g773)) + ((g237) & (g238) & (!g239) & (!g240) & (!g820) & (!g773)) + ((g237) & (g238) & (!g239) & (!g240) & (g820) & (!g773)) + ((g237) & (g238) & (!g239) & (g240) & (!g820) & (!g773)) + ((g237) & (g238) & (!g239) & (g240) & (g820) & (!g773)) + ((g237) & (g238) & (!g239) & (g240) & (g820) & (g773)) + ((g237) & (g238) & (g239) & (!g240) & (!g820) & (!g773)) + ((g237) & (g238) & (g239) & (!g240) & (!g820) & (g773)) + ((g237) & (g238) & (g239) & (!g240) & (g820) & (!g773)) + ((g237) & (g238) & (g239) & (g240) & (!g820) & (!g773)) + ((g237) & (g238) & (g239) & (g240) & (!g820) & (g773)) + ((g237) & (g238) & (g239) & (g240) & (g820) & (!g773)) + ((g237) & (g238) & (g239) & (g240) & (g820) & (g773)));
	assign g1624 = (((!g242) & (!g243) & (!g244) & (g245) & (g820) & (g773)) + ((!g242) & (!g243) & (g244) & (!g245) & (!g820) & (g773)) + ((!g242) & (!g243) & (g244) & (g245) & (!g820) & (g773)) + ((!g242) & (!g243) & (g244) & (g245) & (g820) & (g773)) + ((!g242) & (g243) & (!g244) & (!g245) & (g820) & (!g773)) + ((!g242) & (g243) & (!g244) & (g245) & (g820) & (!g773)) + ((!g242) & (g243) & (!g244) & (g245) & (g820) & (g773)) + ((!g242) & (g243) & (g244) & (!g245) & (!g820) & (g773)) + ((!g242) & (g243) & (g244) & (!g245) & (g820) & (!g773)) + ((!g242) & (g243) & (g244) & (g245) & (!g820) & (g773)) + ((!g242) & (g243) & (g244) & (g245) & (g820) & (!g773)) + ((!g242) & (g243) & (g244) & (g245) & (g820) & (g773)) + ((g242) & (!g243) & (!g244) & (!g245) & (!g820) & (!g773)) + ((g242) & (!g243) & (!g244) & (g245) & (!g820) & (!g773)) + ((g242) & (!g243) & (!g244) & (g245) & (g820) & (g773)) + ((g242) & (!g243) & (g244) & (!g245) & (!g820) & (!g773)) + ((g242) & (!g243) & (g244) & (!g245) & (!g820) & (g773)) + ((g242) & (!g243) & (g244) & (g245) & (!g820) & (!g773)) + ((g242) & (!g243) & (g244) & (g245) & (!g820) & (g773)) + ((g242) & (!g243) & (g244) & (g245) & (g820) & (g773)) + ((g242) & (g243) & (!g244) & (!g245) & (!g820) & (!g773)) + ((g242) & (g243) & (!g244) & (!g245) & (g820) & (!g773)) + ((g242) & (g243) & (!g244) & (g245) & (!g820) & (!g773)) + ((g242) & (g243) & (!g244) & (g245) & (g820) & (!g773)) + ((g242) & (g243) & (!g244) & (g245) & (g820) & (g773)) + ((g242) & (g243) & (g244) & (!g245) & (!g820) & (!g773)) + ((g242) & (g243) & (g244) & (!g245) & (!g820) & (g773)) + ((g242) & (g243) & (g244) & (!g245) & (g820) & (!g773)) + ((g242) & (g243) & (g244) & (g245) & (!g820) & (!g773)) + ((g242) & (g243) & (g244) & (g245) & (!g820) & (g773)) + ((g242) & (g243) & (g244) & (g245) & (g820) & (!g773)) + ((g242) & (g243) & (g244) & (g245) & (g820) & (g773)));
	assign g1625 = (((!g247) & (!g248) & (!g249) & (g250) & (g820) & (g773)) + ((!g247) & (!g248) & (g249) & (!g250) & (!g820) & (g773)) + ((!g247) & (!g248) & (g249) & (g250) & (!g820) & (g773)) + ((!g247) & (!g248) & (g249) & (g250) & (g820) & (g773)) + ((!g247) & (g248) & (!g249) & (!g250) & (g820) & (!g773)) + ((!g247) & (g248) & (!g249) & (g250) & (g820) & (!g773)) + ((!g247) & (g248) & (!g249) & (g250) & (g820) & (g773)) + ((!g247) & (g248) & (g249) & (!g250) & (!g820) & (g773)) + ((!g247) & (g248) & (g249) & (!g250) & (g820) & (!g773)) + ((!g247) & (g248) & (g249) & (g250) & (!g820) & (g773)) + ((!g247) & (g248) & (g249) & (g250) & (g820) & (!g773)) + ((!g247) & (g248) & (g249) & (g250) & (g820) & (g773)) + ((g247) & (!g248) & (!g249) & (!g250) & (!g820) & (!g773)) + ((g247) & (!g248) & (!g249) & (g250) & (!g820) & (!g773)) + ((g247) & (!g248) & (!g249) & (g250) & (g820) & (g773)) + ((g247) & (!g248) & (g249) & (!g250) & (!g820) & (!g773)) + ((g247) & (!g248) & (g249) & (!g250) & (!g820) & (g773)) + ((g247) & (!g248) & (g249) & (g250) & (!g820) & (!g773)) + ((g247) & (!g248) & (g249) & (g250) & (!g820) & (g773)) + ((g247) & (!g248) & (g249) & (g250) & (g820) & (g773)) + ((g247) & (g248) & (!g249) & (!g250) & (!g820) & (!g773)) + ((g247) & (g248) & (!g249) & (!g250) & (g820) & (!g773)) + ((g247) & (g248) & (!g249) & (g250) & (!g820) & (!g773)) + ((g247) & (g248) & (!g249) & (g250) & (g820) & (!g773)) + ((g247) & (g248) & (!g249) & (g250) & (g820) & (g773)) + ((g247) & (g248) & (g249) & (!g250) & (!g820) & (!g773)) + ((g247) & (g248) & (g249) & (!g250) & (!g820) & (g773)) + ((g247) & (g248) & (g249) & (!g250) & (g820) & (!g773)) + ((g247) & (g248) & (g249) & (g250) & (!g820) & (!g773)) + ((g247) & (g248) & (g249) & (g250) & (!g820) & (g773)) + ((g247) & (g248) & (g249) & (g250) & (g820) & (!g773)) + ((g247) & (g248) & (g249) & (g250) & (g820) & (g773)));
	assign g1626 = (((!g1622) & (!g1623) & (!g1624) & (g1625) & (g677) & (g726)) + ((!g1622) & (!g1623) & (g1624) & (!g1625) & (!g677) & (g726)) + ((!g1622) & (!g1623) & (g1624) & (g1625) & (!g677) & (g726)) + ((!g1622) & (!g1623) & (g1624) & (g1625) & (g677) & (g726)) + ((!g1622) & (g1623) & (!g1624) & (!g1625) & (g677) & (!g726)) + ((!g1622) & (g1623) & (!g1624) & (g1625) & (g677) & (!g726)) + ((!g1622) & (g1623) & (!g1624) & (g1625) & (g677) & (g726)) + ((!g1622) & (g1623) & (g1624) & (!g1625) & (!g677) & (g726)) + ((!g1622) & (g1623) & (g1624) & (!g1625) & (g677) & (!g726)) + ((!g1622) & (g1623) & (g1624) & (g1625) & (!g677) & (g726)) + ((!g1622) & (g1623) & (g1624) & (g1625) & (g677) & (!g726)) + ((!g1622) & (g1623) & (g1624) & (g1625) & (g677) & (g726)) + ((g1622) & (!g1623) & (!g1624) & (!g1625) & (!g677) & (!g726)) + ((g1622) & (!g1623) & (!g1624) & (g1625) & (!g677) & (!g726)) + ((g1622) & (!g1623) & (!g1624) & (g1625) & (g677) & (g726)) + ((g1622) & (!g1623) & (g1624) & (!g1625) & (!g677) & (!g726)) + ((g1622) & (!g1623) & (g1624) & (!g1625) & (!g677) & (g726)) + ((g1622) & (!g1623) & (g1624) & (g1625) & (!g677) & (!g726)) + ((g1622) & (!g1623) & (g1624) & (g1625) & (!g677) & (g726)) + ((g1622) & (!g1623) & (g1624) & (g1625) & (g677) & (g726)) + ((g1622) & (g1623) & (!g1624) & (!g1625) & (!g677) & (!g726)) + ((g1622) & (g1623) & (!g1624) & (!g1625) & (g677) & (!g726)) + ((g1622) & (g1623) & (!g1624) & (g1625) & (!g677) & (!g726)) + ((g1622) & (g1623) & (!g1624) & (g1625) & (g677) & (!g726)) + ((g1622) & (g1623) & (!g1624) & (g1625) & (g677) & (g726)) + ((g1622) & (g1623) & (g1624) & (!g1625) & (!g677) & (!g726)) + ((g1622) & (g1623) & (g1624) & (!g1625) & (!g677) & (g726)) + ((g1622) & (g1623) & (g1624) & (!g1625) & (g677) & (!g726)) + ((g1622) & (g1623) & (g1624) & (g1625) & (!g677) & (!g726)) + ((g1622) & (g1623) & (g1624) & (g1625) & (!g677) & (g726)) + ((g1622) & (g1623) & (g1624) & (g1625) & (g677) & (!g726)) + ((g1622) & (g1623) & (g1624) & (g1625) & (g677) & (g726)));
	assign g1627 = (((!g253) & (!g254) & (!g255) & (g256) & (g677) & (g726)) + ((!g253) & (!g254) & (g255) & (!g256) & (!g677) & (g726)) + ((!g253) & (!g254) & (g255) & (g256) & (!g677) & (g726)) + ((!g253) & (!g254) & (g255) & (g256) & (g677) & (g726)) + ((!g253) & (g254) & (!g255) & (!g256) & (g677) & (!g726)) + ((!g253) & (g254) & (!g255) & (g256) & (g677) & (!g726)) + ((!g253) & (g254) & (!g255) & (g256) & (g677) & (g726)) + ((!g253) & (g254) & (g255) & (!g256) & (!g677) & (g726)) + ((!g253) & (g254) & (g255) & (!g256) & (g677) & (!g726)) + ((!g253) & (g254) & (g255) & (g256) & (!g677) & (g726)) + ((!g253) & (g254) & (g255) & (g256) & (g677) & (!g726)) + ((!g253) & (g254) & (g255) & (g256) & (g677) & (g726)) + ((g253) & (!g254) & (!g255) & (!g256) & (!g677) & (!g726)) + ((g253) & (!g254) & (!g255) & (g256) & (!g677) & (!g726)) + ((g253) & (!g254) & (!g255) & (g256) & (g677) & (g726)) + ((g253) & (!g254) & (g255) & (!g256) & (!g677) & (!g726)) + ((g253) & (!g254) & (g255) & (!g256) & (!g677) & (g726)) + ((g253) & (!g254) & (g255) & (g256) & (!g677) & (!g726)) + ((g253) & (!g254) & (g255) & (g256) & (!g677) & (g726)) + ((g253) & (!g254) & (g255) & (g256) & (g677) & (g726)) + ((g253) & (g254) & (!g255) & (!g256) & (!g677) & (!g726)) + ((g253) & (g254) & (!g255) & (!g256) & (g677) & (!g726)) + ((g253) & (g254) & (!g255) & (g256) & (!g677) & (!g726)) + ((g253) & (g254) & (!g255) & (g256) & (g677) & (!g726)) + ((g253) & (g254) & (!g255) & (g256) & (g677) & (g726)) + ((g253) & (g254) & (g255) & (!g256) & (!g677) & (!g726)) + ((g253) & (g254) & (g255) & (!g256) & (!g677) & (g726)) + ((g253) & (g254) & (g255) & (!g256) & (g677) & (!g726)) + ((g253) & (g254) & (g255) & (g256) & (!g677) & (!g726)) + ((g253) & (g254) & (g255) & (g256) & (!g677) & (g726)) + ((g253) & (g254) & (g255) & (g256) & (g677) & (!g726)) + ((g253) & (g254) & (g255) & (g256) & (g677) & (g726)));
	assign g1628 = (((!g677) & (!sk[30]) & (!g726) & (!g258) & (g259) & (!g260)) + ((!g677) & (!sk[30]) & (!g726) & (!g258) & (g259) & (g260)) + ((!g677) & (!sk[30]) & (!g726) & (g258) & (!g259) & (!g260)) + ((!g677) & (!sk[30]) & (!g726) & (g258) & (!g259) & (g260)) + ((!g677) & (!sk[30]) & (!g726) & (g258) & (g259) & (!g260)) + ((!g677) & (!sk[30]) & (!g726) & (g258) & (g259) & (g260)) + ((!g677) & (!sk[30]) & (g726) & (!g258) & (!g259) & (!g260)) + ((!g677) & (!sk[30]) & (g726) & (!g258) & (!g259) & (g260)) + ((!g677) & (!sk[30]) & (g726) & (!g258) & (g259) & (!g260)) + ((!g677) & (!sk[30]) & (g726) & (!g258) & (g259) & (g260)) + ((!g677) & (!sk[30]) & (g726) & (g258) & (!g259) & (!g260)) + ((!g677) & (!sk[30]) & (g726) & (g258) & (!g259) & (g260)) + ((!g677) & (!sk[30]) & (g726) & (g258) & (g259) & (!g260)) + ((!g677) & (!sk[30]) & (g726) & (g258) & (g259) & (g260)) + ((!g677) & (sk[30]) & (g726) & (!g258) & (!g259) & (g260)) + ((!g677) & (sk[30]) & (g726) & (!g258) & (g259) & (g260)) + ((!g677) & (sk[30]) & (g726) & (g258) & (!g259) & (g260)) + ((!g677) & (sk[30]) & (g726) & (g258) & (g259) & (g260)) + ((g677) & (!sk[30]) & (!g726) & (!g258) & (g259) & (!g260)) + ((g677) & (!sk[30]) & (!g726) & (!g258) & (g259) & (g260)) + ((g677) & (!sk[30]) & (!g726) & (g258) & (!g259) & (!g260)) + ((g677) & (!sk[30]) & (!g726) & (g258) & (!g259) & (g260)) + ((g677) & (!sk[30]) & (!g726) & (g258) & (g259) & (!g260)) + ((g677) & (!sk[30]) & (!g726) & (g258) & (g259) & (g260)) + ((g677) & (!sk[30]) & (g726) & (!g258) & (!g259) & (!g260)) + ((g677) & (!sk[30]) & (g726) & (!g258) & (!g259) & (g260)) + ((g677) & (!sk[30]) & (g726) & (!g258) & (g259) & (!g260)) + ((g677) & (!sk[30]) & (g726) & (!g258) & (g259) & (g260)) + ((g677) & (!sk[30]) & (g726) & (g258) & (!g259) & (!g260)) + ((g677) & (!sk[30]) & (g726) & (g258) & (!g259) & (g260)) + ((g677) & (!sk[30]) & (g726) & (g258) & (g259) & (!g260)) + ((g677) & (!sk[30]) & (g726) & (g258) & (g259) & (g260)) + ((g677) & (sk[30]) & (!g726) & (g258) & (!g259) & (!g260)) + ((g677) & (sk[30]) & (!g726) & (g258) & (!g259) & (g260)) + ((g677) & (sk[30]) & (!g726) & (g258) & (g259) & (!g260)) + ((g677) & (sk[30]) & (!g726) & (g258) & (g259) & (g260)) + ((g677) & (sk[30]) & (g726) & (!g258) & (g259) & (!g260)) + ((g677) & (sk[30]) & (g726) & (!g258) & (g259) & (g260)) + ((g677) & (sk[30]) & (g726) & (g258) & (g259) & (!g260)) + ((g677) & (sk[30]) & (g726) & (g258) & (g259) & (g260)));
	assign g1629 = (((!g262) & (!g263) & (!g264) & (g265) & (g677) & (g726)) + ((!g262) & (!g263) & (g264) & (!g265) & (!g677) & (g726)) + ((!g262) & (!g263) & (g264) & (g265) & (!g677) & (g726)) + ((!g262) & (!g263) & (g264) & (g265) & (g677) & (g726)) + ((!g262) & (g263) & (!g264) & (!g265) & (g677) & (!g726)) + ((!g262) & (g263) & (!g264) & (g265) & (g677) & (!g726)) + ((!g262) & (g263) & (!g264) & (g265) & (g677) & (g726)) + ((!g262) & (g263) & (g264) & (!g265) & (!g677) & (g726)) + ((!g262) & (g263) & (g264) & (!g265) & (g677) & (!g726)) + ((!g262) & (g263) & (g264) & (g265) & (!g677) & (g726)) + ((!g262) & (g263) & (g264) & (g265) & (g677) & (!g726)) + ((!g262) & (g263) & (g264) & (g265) & (g677) & (g726)) + ((g262) & (!g263) & (!g264) & (!g265) & (!g677) & (!g726)) + ((g262) & (!g263) & (!g264) & (g265) & (!g677) & (!g726)) + ((g262) & (!g263) & (!g264) & (g265) & (g677) & (g726)) + ((g262) & (!g263) & (g264) & (!g265) & (!g677) & (!g726)) + ((g262) & (!g263) & (g264) & (!g265) & (!g677) & (g726)) + ((g262) & (!g263) & (g264) & (g265) & (!g677) & (!g726)) + ((g262) & (!g263) & (g264) & (g265) & (!g677) & (g726)) + ((g262) & (!g263) & (g264) & (g265) & (g677) & (g726)) + ((g262) & (g263) & (!g264) & (!g265) & (!g677) & (!g726)) + ((g262) & (g263) & (!g264) & (!g265) & (g677) & (!g726)) + ((g262) & (g263) & (!g264) & (g265) & (!g677) & (!g726)) + ((g262) & (g263) & (!g264) & (g265) & (g677) & (!g726)) + ((g262) & (g263) & (!g264) & (g265) & (g677) & (g726)) + ((g262) & (g263) & (g264) & (!g265) & (!g677) & (!g726)) + ((g262) & (g263) & (g264) & (!g265) & (!g677) & (g726)) + ((g262) & (g263) & (g264) & (!g265) & (g677) & (!g726)) + ((g262) & (g263) & (g264) & (g265) & (!g677) & (!g726)) + ((g262) & (g263) & (g264) & (g265) & (!g677) & (g726)) + ((g262) & (g263) & (g264) & (g265) & (g677) & (!g726)) + ((g262) & (g263) & (g264) & (g265) & (g677) & (g726)));
	assign g1630 = (((!g267) & (!g268) & (!g269) & (g270) & (g677) & (g726)) + ((!g267) & (!g268) & (g269) & (!g270) & (!g677) & (g726)) + ((!g267) & (!g268) & (g269) & (g270) & (!g677) & (g726)) + ((!g267) & (!g268) & (g269) & (g270) & (g677) & (g726)) + ((!g267) & (g268) & (!g269) & (!g270) & (g677) & (!g726)) + ((!g267) & (g268) & (!g269) & (g270) & (g677) & (!g726)) + ((!g267) & (g268) & (!g269) & (g270) & (g677) & (g726)) + ((!g267) & (g268) & (g269) & (!g270) & (!g677) & (g726)) + ((!g267) & (g268) & (g269) & (!g270) & (g677) & (!g726)) + ((!g267) & (g268) & (g269) & (g270) & (!g677) & (g726)) + ((!g267) & (g268) & (g269) & (g270) & (g677) & (!g726)) + ((!g267) & (g268) & (g269) & (g270) & (g677) & (g726)) + ((g267) & (!g268) & (!g269) & (!g270) & (!g677) & (!g726)) + ((g267) & (!g268) & (!g269) & (g270) & (!g677) & (!g726)) + ((g267) & (!g268) & (!g269) & (g270) & (g677) & (g726)) + ((g267) & (!g268) & (g269) & (!g270) & (!g677) & (!g726)) + ((g267) & (!g268) & (g269) & (!g270) & (!g677) & (g726)) + ((g267) & (!g268) & (g269) & (g270) & (!g677) & (!g726)) + ((g267) & (!g268) & (g269) & (g270) & (!g677) & (g726)) + ((g267) & (!g268) & (g269) & (g270) & (g677) & (g726)) + ((g267) & (g268) & (!g269) & (!g270) & (!g677) & (!g726)) + ((g267) & (g268) & (!g269) & (!g270) & (g677) & (!g726)) + ((g267) & (g268) & (!g269) & (g270) & (!g677) & (!g726)) + ((g267) & (g268) & (!g269) & (g270) & (g677) & (!g726)) + ((g267) & (g268) & (!g269) & (g270) & (g677) & (g726)) + ((g267) & (g268) & (g269) & (!g270) & (!g677) & (!g726)) + ((g267) & (g268) & (g269) & (!g270) & (!g677) & (g726)) + ((g267) & (g268) & (g269) & (!g270) & (g677) & (!g726)) + ((g267) & (g268) & (g269) & (g270) & (!g677) & (!g726)) + ((g267) & (g268) & (g269) & (g270) & (!g677) & (g726)) + ((g267) & (g268) & (g269) & (g270) & (g677) & (!g726)) + ((g267) & (g268) & (g269) & (g270) & (g677) & (g726)));
	assign g1631 = (((!g820) & (!g773) & (!g1627) & (g1628) & (!g1629) & (!g1630)) + ((!g820) & (!g773) & (!g1627) & (g1628) & (!g1629) & (g1630)) + ((!g820) & (!g773) & (!g1627) & (g1628) & (g1629) & (!g1630)) + ((!g820) & (!g773) & (!g1627) & (g1628) & (g1629) & (g1630)) + ((!g820) & (!g773) & (g1627) & (g1628) & (!g1629) & (!g1630)) + ((!g820) & (!g773) & (g1627) & (g1628) & (!g1629) & (g1630)) + ((!g820) & (!g773) & (g1627) & (g1628) & (g1629) & (!g1630)) + ((!g820) & (!g773) & (g1627) & (g1628) & (g1629) & (g1630)) + ((!g820) & (g773) & (!g1627) & (!g1628) & (!g1629) & (g1630)) + ((!g820) & (g773) & (!g1627) & (!g1628) & (g1629) & (g1630)) + ((!g820) & (g773) & (!g1627) & (g1628) & (!g1629) & (g1630)) + ((!g820) & (g773) & (!g1627) & (g1628) & (g1629) & (g1630)) + ((!g820) & (g773) & (g1627) & (!g1628) & (!g1629) & (g1630)) + ((!g820) & (g773) & (g1627) & (!g1628) & (g1629) & (g1630)) + ((!g820) & (g773) & (g1627) & (g1628) & (!g1629) & (g1630)) + ((!g820) & (g773) & (g1627) & (g1628) & (g1629) & (g1630)) + ((g820) & (!g773) & (g1627) & (!g1628) & (!g1629) & (!g1630)) + ((g820) & (!g773) & (g1627) & (!g1628) & (!g1629) & (g1630)) + ((g820) & (!g773) & (g1627) & (!g1628) & (g1629) & (!g1630)) + ((g820) & (!g773) & (g1627) & (!g1628) & (g1629) & (g1630)) + ((g820) & (!g773) & (g1627) & (g1628) & (!g1629) & (!g1630)) + ((g820) & (!g773) & (g1627) & (g1628) & (!g1629) & (g1630)) + ((g820) & (!g773) & (g1627) & (g1628) & (g1629) & (!g1630)) + ((g820) & (!g773) & (g1627) & (g1628) & (g1629) & (g1630)) + ((g820) & (g773) & (!g1627) & (!g1628) & (g1629) & (!g1630)) + ((g820) & (g773) & (!g1627) & (!g1628) & (g1629) & (g1630)) + ((g820) & (g773) & (!g1627) & (g1628) & (g1629) & (!g1630)) + ((g820) & (g773) & (!g1627) & (g1628) & (g1629) & (g1630)) + ((g820) & (g773) & (g1627) & (!g1628) & (g1629) & (!g1630)) + ((g820) & (g773) & (g1627) & (!g1628) & (g1629) & (g1630)) + ((g820) & (g773) & (g1627) & (g1628) & (g1629) & (!g1630)) + ((g820) & (g773) & (g1627) & (g1628) & (g1629) & (g1630)));
	assign g1632 = (((!g867) & (!sk[34]) & (!g1626) & (g1631)) + ((!g867) & (!sk[34]) & (g1626) & (!g1631)) + ((!g867) & (!sk[34]) & (g1626) & (g1631)) + ((!g867) & (sk[34]) & (!g1626) & (g1631)) + ((!g867) & (sk[34]) & (g1626) & (g1631)) + ((g867) & (!sk[34]) & (!g1626) & (g1631)) + ((g867) & (!sk[34]) & (g1626) & (!g1631)) + ((g867) & (!sk[34]) & (g1626) & (g1631)) + ((g867) & (sk[34]) & (g1626) & (!g1631)) + ((g867) & (sk[34]) & (g1626) & (g1631)));
	assign g1633 = (((!g1592) & (!g1593) & (!g1605) & (g1607) & (!g37) & (g1632)) + ((!g1592) & (!g1593) & (!g1605) & (g1607) & (g37) & (g1632)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (!g37) & (g1632)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (g37) & (g1632)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (!g37) & (g1632)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (g37) & (g1632)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (!g37) & (g1632)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (g37) & (g1632)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (!g37) & (g1632)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (g37) & (g1632)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g37) & (!g1632)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g37) & (g1632)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g37) & (!g1632)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g37) & (g1632)));
	assign g1634 = (((!g276) & (!g281) & (!g286) & (g291) & (g820) & (g773)) + ((!g276) & (!g281) & (g286) & (!g291) & (!g820) & (g773)) + ((!g276) & (!g281) & (g286) & (g291) & (!g820) & (g773)) + ((!g276) & (!g281) & (g286) & (g291) & (g820) & (g773)) + ((!g276) & (g281) & (!g286) & (!g291) & (g820) & (!g773)) + ((!g276) & (g281) & (!g286) & (g291) & (g820) & (!g773)) + ((!g276) & (g281) & (!g286) & (g291) & (g820) & (g773)) + ((!g276) & (g281) & (g286) & (!g291) & (!g820) & (g773)) + ((!g276) & (g281) & (g286) & (!g291) & (g820) & (!g773)) + ((!g276) & (g281) & (g286) & (g291) & (!g820) & (g773)) + ((!g276) & (g281) & (g286) & (g291) & (g820) & (!g773)) + ((!g276) & (g281) & (g286) & (g291) & (g820) & (g773)) + ((g276) & (!g281) & (!g286) & (!g291) & (!g820) & (!g773)) + ((g276) & (!g281) & (!g286) & (g291) & (!g820) & (!g773)) + ((g276) & (!g281) & (!g286) & (g291) & (g820) & (g773)) + ((g276) & (!g281) & (g286) & (!g291) & (!g820) & (!g773)) + ((g276) & (!g281) & (g286) & (!g291) & (!g820) & (g773)) + ((g276) & (!g281) & (g286) & (g291) & (!g820) & (!g773)) + ((g276) & (!g281) & (g286) & (g291) & (!g820) & (g773)) + ((g276) & (!g281) & (g286) & (g291) & (g820) & (g773)) + ((g276) & (g281) & (!g286) & (!g291) & (!g820) & (!g773)) + ((g276) & (g281) & (!g286) & (!g291) & (g820) & (!g773)) + ((g276) & (g281) & (!g286) & (g291) & (!g820) & (!g773)) + ((g276) & (g281) & (!g286) & (g291) & (g820) & (!g773)) + ((g276) & (g281) & (!g286) & (g291) & (g820) & (g773)) + ((g276) & (g281) & (g286) & (!g291) & (!g820) & (!g773)) + ((g276) & (g281) & (g286) & (!g291) & (!g820) & (g773)) + ((g276) & (g281) & (g286) & (!g291) & (g820) & (!g773)) + ((g276) & (g281) & (g286) & (g291) & (!g820) & (!g773)) + ((g276) & (g281) & (g286) & (g291) & (!g820) & (g773)) + ((g276) & (g281) & (g286) & (g291) & (g820) & (!g773)) + ((g276) & (g281) & (g286) & (g291) & (g820) & (g773)));
	assign g1635 = (((!g277) & (!g282) & (!g287) & (g292) & (g820) & (g773)) + ((!g277) & (!g282) & (g287) & (!g292) & (!g820) & (g773)) + ((!g277) & (!g282) & (g287) & (g292) & (!g820) & (g773)) + ((!g277) & (!g282) & (g287) & (g292) & (g820) & (g773)) + ((!g277) & (g282) & (!g287) & (!g292) & (g820) & (!g773)) + ((!g277) & (g282) & (!g287) & (g292) & (g820) & (!g773)) + ((!g277) & (g282) & (!g287) & (g292) & (g820) & (g773)) + ((!g277) & (g282) & (g287) & (!g292) & (!g820) & (g773)) + ((!g277) & (g282) & (g287) & (!g292) & (g820) & (!g773)) + ((!g277) & (g282) & (g287) & (g292) & (!g820) & (g773)) + ((!g277) & (g282) & (g287) & (g292) & (g820) & (!g773)) + ((!g277) & (g282) & (g287) & (g292) & (g820) & (g773)) + ((g277) & (!g282) & (!g287) & (!g292) & (!g820) & (!g773)) + ((g277) & (!g282) & (!g287) & (g292) & (!g820) & (!g773)) + ((g277) & (!g282) & (!g287) & (g292) & (g820) & (g773)) + ((g277) & (!g282) & (g287) & (!g292) & (!g820) & (!g773)) + ((g277) & (!g282) & (g287) & (!g292) & (!g820) & (g773)) + ((g277) & (!g282) & (g287) & (g292) & (!g820) & (!g773)) + ((g277) & (!g282) & (g287) & (g292) & (!g820) & (g773)) + ((g277) & (!g282) & (g287) & (g292) & (g820) & (g773)) + ((g277) & (g282) & (!g287) & (!g292) & (!g820) & (!g773)) + ((g277) & (g282) & (!g287) & (!g292) & (g820) & (!g773)) + ((g277) & (g282) & (!g287) & (g292) & (!g820) & (!g773)) + ((g277) & (g282) & (!g287) & (g292) & (g820) & (!g773)) + ((g277) & (g282) & (!g287) & (g292) & (g820) & (g773)) + ((g277) & (g282) & (g287) & (!g292) & (!g820) & (!g773)) + ((g277) & (g282) & (g287) & (!g292) & (!g820) & (g773)) + ((g277) & (g282) & (g287) & (!g292) & (g820) & (!g773)) + ((g277) & (g282) & (g287) & (g292) & (!g820) & (!g773)) + ((g277) & (g282) & (g287) & (g292) & (!g820) & (g773)) + ((g277) & (g282) & (g287) & (g292) & (g820) & (!g773)) + ((g277) & (g282) & (g287) & (g292) & (g820) & (g773)));
	assign g1636 = (((!g278) & (!g283) & (!g288) & (g293) & (g820) & (g773)) + ((!g278) & (!g283) & (g288) & (!g293) & (!g820) & (g773)) + ((!g278) & (!g283) & (g288) & (g293) & (!g820) & (g773)) + ((!g278) & (!g283) & (g288) & (g293) & (g820) & (g773)) + ((!g278) & (g283) & (!g288) & (!g293) & (g820) & (!g773)) + ((!g278) & (g283) & (!g288) & (g293) & (g820) & (!g773)) + ((!g278) & (g283) & (!g288) & (g293) & (g820) & (g773)) + ((!g278) & (g283) & (g288) & (!g293) & (!g820) & (g773)) + ((!g278) & (g283) & (g288) & (!g293) & (g820) & (!g773)) + ((!g278) & (g283) & (g288) & (g293) & (!g820) & (g773)) + ((!g278) & (g283) & (g288) & (g293) & (g820) & (!g773)) + ((!g278) & (g283) & (g288) & (g293) & (g820) & (g773)) + ((g278) & (!g283) & (!g288) & (!g293) & (!g820) & (!g773)) + ((g278) & (!g283) & (!g288) & (g293) & (!g820) & (!g773)) + ((g278) & (!g283) & (!g288) & (g293) & (g820) & (g773)) + ((g278) & (!g283) & (g288) & (!g293) & (!g820) & (!g773)) + ((g278) & (!g283) & (g288) & (!g293) & (!g820) & (g773)) + ((g278) & (!g283) & (g288) & (g293) & (!g820) & (!g773)) + ((g278) & (!g283) & (g288) & (g293) & (!g820) & (g773)) + ((g278) & (!g283) & (g288) & (g293) & (g820) & (g773)) + ((g278) & (g283) & (!g288) & (!g293) & (!g820) & (!g773)) + ((g278) & (g283) & (!g288) & (!g293) & (g820) & (!g773)) + ((g278) & (g283) & (!g288) & (g293) & (!g820) & (!g773)) + ((g278) & (g283) & (!g288) & (g293) & (g820) & (!g773)) + ((g278) & (g283) & (!g288) & (g293) & (g820) & (g773)) + ((g278) & (g283) & (g288) & (!g293) & (!g820) & (!g773)) + ((g278) & (g283) & (g288) & (!g293) & (!g820) & (g773)) + ((g278) & (g283) & (g288) & (!g293) & (g820) & (!g773)) + ((g278) & (g283) & (g288) & (g293) & (!g820) & (!g773)) + ((g278) & (g283) & (g288) & (g293) & (!g820) & (g773)) + ((g278) & (g283) & (g288) & (g293) & (g820) & (!g773)) + ((g278) & (g283) & (g288) & (g293) & (g820) & (g773)));
	assign g1637 = (((!g279) & (!g284) & (!g289) & (g294) & (g820) & (g773)) + ((!g279) & (!g284) & (g289) & (!g294) & (!g820) & (g773)) + ((!g279) & (!g284) & (g289) & (g294) & (!g820) & (g773)) + ((!g279) & (!g284) & (g289) & (g294) & (g820) & (g773)) + ((!g279) & (g284) & (!g289) & (!g294) & (g820) & (!g773)) + ((!g279) & (g284) & (!g289) & (g294) & (g820) & (!g773)) + ((!g279) & (g284) & (!g289) & (g294) & (g820) & (g773)) + ((!g279) & (g284) & (g289) & (!g294) & (!g820) & (g773)) + ((!g279) & (g284) & (g289) & (!g294) & (g820) & (!g773)) + ((!g279) & (g284) & (g289) & (g294) & (!g820) & (g773)) + ((!g279) & (g284) & (g289) & (g294) & (g820) & (!g773)) + ((!g279) & (g284) & (g289) & (g294) & (g820) & (g773)) + ((g279) & (!g284) & (!g289) & (!g294) & (!g820) & (!g773)) + ((g279) & (!g284) & (!g289) & (g294) & (!g820) & (!g773)) + ((g279) & (!g284) & (!g289) & (g294) & (g820) & (g773)) + ((g279) & (!g284) & (g289) & (!g294) & (!g820) & (!g773)) + ((g279) & (!g284) & (g289) & (!g294) & (!g820) & (g773)) + ((g279) & (!g284) & (g289) & (g294) & (!g820) & (!g773)) + ((g279) & (!g284) & (g289) & (g294) & (!g820) & (g773)) + ((g279) & (!g284) & (g289) & (g294) & (g820) & (g773)) + ((g279) & (g284) & (!g289) & (!g294) & (!g820) & (!g773)) + ((g279) & (g284) & (!g289) & (!g294) & (g820) & (!g773)) + ((g279) & (g284) & (!g289) & (g294) & (!g820) & (!g773)) + ((g279) & (g284) & (!g289) & (g294) & (g820) & (!g773)) + ((g279) & (g284) & (!g289) & (g294) & (g820) & (g773)) + ((g279) & (g284) & (g289) & (!g294) & (!g820) & (!g773)) + ((g279) & (g284) & (g289) & (!g294) & (!g820) & (g773)) + ((g279) & (g284) & (g289) & (!g294) & (g820) & (!g773)) + ((g279) & (g284) & (g289) & (g294) & (!g820) & (!g773)) + ((g279) & (g284) & (g289) & (g294) & (!g820) & (g773)) + ((g279) & (g284) & (g289) & (g294) & (g820) & (!g773)) + ((g279) & (g284) & (g289) & (g294) & (g820) & (g773)));
	assign g1638 = (((!g1634) & (!g1635) & (!g1636) & (g1637) & (g677) & (g726)) + ((!g1634) & (!g1635) & (g1636) & (!g1637) & (!g677) & (g726)) + ((!g1634) & (!g1635) & (g1636) & (g1637) & (!g677) & (g726)) + ((!g1634) & (!g1635) & (g1636) & (g1637) & (g677) & (g726)) + ((!g1634) & (g1635) & (!g1636) & (!g1637) & (g677) & (!g726)) + ((!g1634) & (g1635) & (!g1636) & (g1637) & (g677) & (!g726)) + ((!g1634) & (g1635) & (!g1636) & (g1637) & (g677) & (g726)) + ((!g1634) & (g1635) & (g1636) & (!g1637) & (!g677) & (g726)) + ((!g1634) & (g1635) & (g1636) & (!g1637) & (g677) & (!g726)) + ((!g1634) & (g1635) & (g1636) & (g1637) & (!g677) & (g726)) + ((!g1634) & (g1635) & (g1636) & (g1637) & (g677) & (!g726)) + ((!g1634) & (g1635) & (g1636) & (g1637) & (g677) & (g726)) + ((g1634) & (!g1635) & (!g1636) & (!g1637) & (!g677) & (!g726)) + ((g1634) & (!g1635) & (!g1636) & (g1637) & (!g677) & (!g726)) + ((g1634) & (!g1635) & (!g1636) & (g1637) & (g677) & (g726)) + ((g1634) & (!g1635) & (g1636) & (!g1637) & (!g677) & (!g726)) + ((g1634) & (!g1635) & (g1636) & (!g1637) & (!g677) & (g726)) + ((g1634) & (!g1635) & (g1636) & (g1637) & (!g677) & (!g726)) + ((g1634) & (!g1635) & (g1636) & (g1637) & (!g677) & (g726)) + ((g1634) & (!g1635) & (g1636) & (g1637) & (g677) & (g726)) + ((g1634) & (g1635) & (!g1636) & (!g1637) & (!g677) & (!g726)) + ((g1634) & (g1635) & (!g1636) & (!g1637) & (g677) & (!g726)) + ((g1634) & (g1635) & (!g1636) & (g1637) & (!g677) & (!g726)) + ((g1634) & (g1635) & (!g1636) & (g1637) & (g677) & (!g726)) + ((g1634) & (g1635) & (!g1636) & (g1637) & (g677) & (g726)) + ((g1634) & (g1635) & (g1636) & (!g1637) & (!g677) & (!g726)) + ((g1634) & (g1635) & (g1636) & (!g1637) & (!g677) & (g726)) + ((g1634) & (g1635) & (g1636) & (!g1637) & (g677) & (!g726)) + ((g1634) & (g1635) & (g1636) & (g1637) & (!g677) & (!g726)) + ((g1634) & (g1635) & (g1636) & (g1637) & (!g677) & (g726)) + ((g1634) & (g1635) & (g1636) & (g1637) & (g677) & (!g726)) + ((g1634) & (g1635) & (g1636) & (g1637) & (g677) & (g726)));
	assign g1639 = (((!g297) & (!g298) & (!g299) & (g300) & (g677) & (g726)) + ((!g297) & (!g298) & (g299) & (!g300) & (!g677) & (g726)) + ((!g297) & (!g298) & (g299) & (g300) & (!g677) & (g726)) + ((!g297) & (!g298) & (g299) & (g300) & (g677) & (g726)) + ((!g297) & (g298) & (!g299) & (!g300) & (g677) & (!g726)) + ((!g297) & (g298) & (!g299) & (g300) & (g677) & (!g726)) + ((!g297) & (g298) & (!g299) & (g300) & (g677) & (g726)) + ((!g297) & (g298) & (g299) & (!g300) & (!g677) & (g726)) + ((!g297) & (g298) & (g299) & (!g300) & (g677) & (!g726)) + ((!g297) & (g298) & (g299) & (g300) & (!g677) & (g726)) + ((!g297) & (g298) & (g299) & (g300) & (g677) & (!g726)) + ((!g297) & (g298) & (g299) & (g300) & (g677) & (g726)) + ((g297) & (!g298) & (!g299) & (!g300) & (!g677) & (!g726)) + ((g297) & (!g298) & (!g299) & (g300) & (!g677) & (!g726)) + ((g297) & (!g298) & (!g299) & (g300) & (g677) & (g726)) + ((g297) & (!g298) & (g299) & (!g300) & (!g677) & (!g726)) + ((g297) & (!g298) & (g299) & (!g300) & (!g677) & (g726)) + ((g297) & (!g298) & (g299) & (g300) & (!g677) & (!g726)) + ((g297) & (!g298) & (g299) & (g300) & (!g677) & (g726)) + ((g297) & (!g298) & (g299) & (g300) & (g677) & (g726)) + ((g297) & (g298) & (!g299) & (!g300) & (!g677) & (!g726)) + ((g297) & (g298) & (!g299) & (!g300) & (g677) & (!g726)) + ((g297) & (g298) & (!g299) & (g300) & (!g677) & (!g726)) + ((g297) & (g298) & (!g299) & (g300) & (g677) & (!g726)) + ((g297) & (g298) & (!g299) & (g300) & (g677) & (g726)) + ((g297) & (g298) & (g299) & (!g300) & (!g677) & (!g726)) + ((g297) & (g298) & (g299) & (!g300) & (!g677) & (g726)) + ((g297) & (g298) & (g299) & (!g300) & (g677) & (!g726)) + ((g297) & (g298) & (g299) & (g300) & (!g677) & (!g726)) + ((g297) & (g298) & (g299) & (g300) & (!g677) & (g726)) + ((g297) & (g298) & (g299) & (g300) & (g677) & (!g726)) + ((g297) & (g298) & (g299) & (g300) & (g677) & (g726)));
	assign g1640 = (((!g677) & (!g726) & (!g302) & (g303) & (!sk[42]) & (!g304)) + ((!g677) & (!g726) & (!g302) & (g303) & (!sk[42]) & (g304)) + ((!g677) & (!g726) & (g302) & (!g303) & (!sk[42]) & (!g304)) + ((!g677) & (!g726) & (g302) & (!g303) & (!sk[42]) & (g304)) + ((!g677) & (!g726) & (g302) & (g303) & (!sk[42]) & (!g304)) + ((!g677) & (!g726) & (g302) & (g303) & (!sk[42]) & (g304)) + ((!g677) & (g726) & (!g302) & (!g303) & (!sk[42]) & (!g304)) + ((!g677) & (g726) & (!g302) & (!g303) & (!sk[42]) & (g304)) + ((!g677) & (g726) & (!g302) & (!g303) & (sk[42]) & (g304)) + ((!g677) & (g726) & (!g302) & (g303) & (!sk[42]) & (!g304)) + ((!g677) & (g726) & (!g302) & (g303) & (!sk[42]) & (g304)) + ((!g677) & (g726) & (!g302) & (g303) & (sk[42]) & (g304)) + ((!g677) & (g726) & (g302) & (!g303) & (!sk[42]) & (!g304)) + ((!g677) & (g726) & (g302) & (!g303) & (!sk[42]) & (g304)) + ((!g677) & (g726) & (g302) & (!g303) & (sk[42]) & (g304)) + ((!g677) & (g726) & (g302) & (g303) & (!sk[42]) & (!g304)) + ((!g677) & (g726) & (g302) & (g303) & (!sk[42]) & (g304)) + ((!g677) & (g726) & (g302) & (g303) & (sk[42]) & (g304)) + ((g677) & (!g726) & (!g302) & (g303) & (!sk[42]) & (!g304)) + ((g677) & (!g726) & (!g302) & (g303) & (!sk[42]) & (g304)) + ((g677) & (!g726) & (g302) & (!g303) & (!sk[42]) & (!g304)) + ((g677) & (!g726) & (g302) & (!g303) & (!sk[42]) & (g304)) + ((g677) & (!g726) & (g302) & (!g303) & (sk[42]) & (!g304)) + ((g677) & (!g726) & (g302) & (!g303) & (sk[42]) & (g304)) + ((g677) & (!g726) & (g302) & (g303) & (!sk[42]) & (!g304)) + ((g677) & (!g726) & (g302) & (g303) & (!sk[42]) & (g304)) + ((g677) & (!g726) & (g302) & (g303) & (sk[42]) & (!g304)) + ((g677) & (!g726) & (g302) & (g303) & (sk[42]) & (g304)) + ((g677) & (g726) & (!g302) & (!g303) & (!sk[42]) & (!g304)) + ((g677) & (g726) & (!g302) & (!g303) & (!sk[42]) & (g304)) + ((g677) & (g726) & (!g302) & (g303) & (!sk[42]) & (!g304)) + ((g677) & (g726) & (!g302) & (g303) & (!sk[42]) & (g304)) + ((g677) & (g726) & (!g302) & (g303) & (sk[42]) & (!g304)) + ((g677) & (g726) & (!g302) & (g303) & (sk[42]) & (g304)) + ((g677) & (g726) & (g302) & (!g303) & (!sk[42]) & (!g304)) + ((g677) & (g726) & (g302) & (!g303) & (!sk[42]) & (g304)) + ((g677) & (g726) & (g302) & (g303) & (!sk[42]) & (!g304)) + ((g677) & (g726) & (g302) & (g303) & (!sk[42]) & (g304)) + ((g677) & (g726) & (g302) & (g303) & (sk[42]) & (!g304)) + ((g677) & (g726) & (g302) & (g303) & (sk[42]) & (g304)));
	assign g1641 = (((!g306) & (!g307) & (!g308) & (g309) & (g677) & (g726)) + ((!g306) & (!g307) & (g308) & (!g309) & (!g677) & (g726)) + ((!g306) & (!g307) & (g308) & (g309) & (!g677) & (g726)) + ((!g306) & (!g307) & (g308) & (g309) & (g677) & (g726)) + ((!g306) & (g307) & (!g308) & (!g309) & (g677) & (!g726)) + ((!g306) & (g307) & (!g308) & (g309) & (g677) & (!g726)) + ((!g306) & (g307) & (!g308) & (g309) & (g677) & (g726)) + ((!g306) & (g307) & (g308) & (!g309) & (!g677) & (g726)) + ((!g306) & (g307) & (g308) & (!g309) & (g677) & (!g726)) + ((!g306) & (g307) & (g308) & (g309) & (!g677) & (g726)) + ((!g306) & (g307) & (g308) & (g309) & (g677) & (!g726)) + ((!g306) & (g307) & (g308) & (g309) & (g677) & (g726)) + ((g306) & (!g307) & (!g308) & (!g309) & (!g677) & (!g726)) + ((g306) & (!g307) & (!g308) & (g309) & (!g677) & (!g726)) + ((g306) & (!g307) & (!g308) & (g309) & (g677) & (g726)) + ((g306) & (!g307) & (g308) & (!g309) & (!g677) & (!g726)) + ((g306) & (!g307) & (g308) & (!g309) & (!g677) & (g726)) + ((g306) & (!g307) & (g308) & (g309) & (!g677) & (!g726)) + ((g306) & (!g307) & (g308) & (g309) & (!g677) & (g726)) + ((g306) & (!g307) & (g308) & (g309) & (g677) & (g726)) + ((g306) & (g307) & (!g308) & (!g309) & (!g677) & (!g726)) + ((g306) & (g307) & (!g308) & (!g309) & (g677) & (!g726)) + ((g306) & (g307) & (!g308) & (g309) & (!g677) & (!g726)) + ((g306) & (g307) & (!g308) & (g309) & (g677) & (!g726)) + ((g306) & (g307) & (!g308) & (g309) & (g677) & (g726)) + ((g306) & (g307) & (g308) & (!g309) & (!g677) & (!g726)) + ((g306) & (g307) & (g308) & (!g309) & (!g677) & (g726)) + ((g306) & (g307) & (g308) & (!g309) & (g677) & (!g726)) + ((g306) & (g307) & (g308) & (g309) & (!g677) & (!g726)) + ((g306) & (g307) & (g308) & (g309) & (!g677) & (g726)) + ((g306) & (g307) & (g308) & (g309) & (g677) & (!g726)) + ((g306) & (g307) & (g308) & (g309) & (g677) & (g726)));
	assign g1642 = (((!g311) & (!g312) & (!g313) & (g314) & (g677) & (g726)) + ((!g311) & (!g312) & (g313) & (!g314) & (!g677) & (g726)) + ((!g311) & (!g312) & (g313) & (g314) & (!g677) & (g726)) + ((!g311) & (!g312) & (g313) & (g314) & (g677) & (g726)) + ((!g311) & (g312) & (!g313) & (!g314) & (g677) & (!g726)) + ((!g311) & (g312) & (!g313) & (g314) & (g677) & (!g726)) + ((!g311) & (g312) & (!g313) & (g314) & (g677) & (g726)) + ((!g311) & (g312) & (g313) & (!g314) & (!g677) & (g726)) + ((!g311) & (g312) & (g313) & (!g314) & (g677) & (!g726)) + ((!g311) & (g312) & (g313) & (g314) & (!g677) & (g726)) + ((!g311) & (g312) & (g313) & (g314) & (g677) & (!g726)) + ((!g311) & (g312) & (g313) & (g314) & (g677) & (g726)) + ((g311) & (!g312) & (!g313) & (!g314) & (!g677) & (!g726)) + ((g311) & (!g312) & (!g313) & (g314) & (!g677) & (!g726)) + ((g311) & (!g312) & (!g313) & (g314) & (g677) & (g726)) + ((g311) & (!g312) & (g313) & (!g314) & (!g677) & (!g726)) + ((g311) & (!g312) & (g313) & (!g314) & (!g677) & (g726)) + ((g311) & (!g312) & (g313) & (g314) & (!g677) & (!g726)) + ((g311) & (!g312) & (g313) & (g314) & (!g677) & (g726)) + ((g311) & (!g312) & (g313) & (g314) & (g677) & (g726)) + ((g311) & (g312) & (!g313) & (!g314) & (!g677) & (!g726)) + ((g311) & (g312) & (!g313) & (!g314) & (g677) & (!g726)) + ((g311) & (g312) & (!g313) & (g314) & (!g677) & (!g726)) + ((g311) & (g312) & (!g313) & (g314) & (g677) & (!g726)) + ((g311) & (g312) & (!g313) & (g314) & (g677) & (g726)) + ((g311) & (g312) & (g313) & (!g314) & (!g677) & (!g726)) + ((g311) & (g312) & (g313) & (!g314) & (!g677) & (g726)) + ((g311) & (g312) & (g313) & (!g314) & (g677) & (!g726)) + ((g311) & (g312) & (g313) & (g314) & (!g677) & (!g726)) + ((g311) & (g312) & (g313) & (g314) & (!g677) & (g726)) + ((g311) & (g312) & (g313) & (g314) & (g677) & (!g726)) + ((g311) & (g312) & (g313) & (g314) & (g677) & (g726)));
	assign g1643 = (((!g820) & (!g773) & (!g1639) & (g1640) & (!g1641) & (!g1642)) + ((!g820) & (!g773) & (!g1639) & (g1640) & (!g1641) & (g1642)) + ((!g820) & (!g773) & (!g1639) & (g1640) & (g1641) & (!g1642)) + ((!g820) & (!g773) & (!g1639) & (g1640) & (g1641) & (g1642)) + ((!g820) & (!g773) & (g1639) & (g1640) & (!g1641) & (!g1642)) + ((!g820) & (!g773) & (g1639) & (g1640) & (!g1641) & (g1642)) + ((!g820) & (!g773) & (g1639) & (g1640) & (g1641) & (!g1642)) + ((!g820) & (!g773) & (g1639) & (g1640) & (g1641) & (g1642)) + ((!g820) & (g773) & (!g1639) & (!g1640) & (!g1641) & (g1642)) + ((!g820) & (g773) & (!g1639) & (!g1640) & (g1641) & (g1642)) + ((!g820) & (g773) & (!g1639) & (g1640) & (!g1641) & (g1642)) + ((!g820) & (g773) & (!g1639) & (g1640) & (g1641) & (g1642)) + ((!g820) & (g773) & (g1639) & (!g1640) & (!g1641) & (g1642)) + ((!g820) & (g773) & (g1639) & (!g1640) & (g1641) & (g1642)) + ((!g820) & (g773) & (g1639) & (g1640) & (!g1641) & (g1642)) + ((!g820) & (g773) & (g1639) & (g1640) & (g1641) & (g1642)) + ((g820) & (!g773) & (g1639) & (!g1640) & (!g1641) & (!g1642)) + ((g820) & (!g773) & (g1639) & (!g1640) & (!g1641) & (g1642)) + ((g820) & (!g773) & (g1639) & (!g1640) & (g1641) & (!g1642)) + ((g820) & (!g773) & (g1639) & (!g1640) & (g1641) & (g1642)) + ((g820) & (!g773) & (g1639) & (g1640) & (!g1641) & (!g1642)) + ((g820) & (!g773) & (g1639) & (g1640) & (!g1641) & (g1642)) + ((g820) & (!g773) & (g1639) & (g1640) & (g1641) & (!g1642)) + ((g820) & (!g773) & (g1639) & (g1640) & (g1641) & (g1642)) + ((g820) & (g773) & (!g1639) & (!g1640) & (g1641) & (!g1642)) + ((g820) & (g773) & (!g1639) & (!g1640) & (g1641) & (g1642)) + ((g820) & (g773) & (!g1639) & (g1640) & (g1641) & (!g1642)) + ((g820) & (g773) & (!g1639) & (g1640) & (g1641) & (g1642)) + ((g820) & (g773) & (g1639) & (!g1640) & (g1641) & (!g1642)) + ((g820) & (g773) & (g1639) & (!g1640) & (g1641) & (g1642)) + ((g820) & (g773) & (g1639) & (g1640) & (g1641) & (!g1642)) + ((g820) & (g773) & (g1639) & (g1640) & (g1641) & (g1642)));
	assign g1644 = (((!sk[46]) & (!g867) & (!g1638) & (g1643)) + ((!sk[46]) & (!g867) & (g1638) & (!g1643)) + ((!sk[46]) & (!g867) & (g1638) & (g1643)) + ((!sk[46]) & (g867) & (!g1638) & (g1643)) + ((!sk[46]) & (g867) & (g1638) & (!g1643)) + ((!sk[46]) & (g867) & (g1638) & (g1643)) + ((sk[46]) & (!g867) & (!g1638) & (g1643)) + ((sk[46]) & (!g867) & (g1638) & (g1643)) + ((sk[46]) & (g867) & (g1638) & (!g1643)) + ((sk[46]) & (g867) & (g1638) & (g1643)));
	assign g1645 = (((!g1592) & (!g1593) & (!g1605) & (g1607) & (!g38) & (g1644)) + ((!g1592) & (!g1593) & (!g1605) & (g1607) & (g38) & (g1644)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (!g38) & (g1644)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (g38) & (g1644)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (!g38) & (g1644)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (g38) & (g1644)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (!g38) & (g1644)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (g38) & (g1644)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (!g38) & (g1644)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (g38) & (g1644)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g38) & (!g1644)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g38) & (g1644)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g38) & (!g1644)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g38) & (g1644)));
	assign g1646 = (((!g321) & (!g322) & (!g323) & (g324) & (g820) & (g773)) + ((!g321) & (!g322) & (g323) & (!g324) & (!g820) & (g773)) + ((!g321) & (!g322) & (g323) & (g324) & (!g820) & (g773)) + ((!g321) & (!g322) & (g323) & (g324) & (g820) & (g773)) + ((!g321) & (g322) & (!g323) & (!g324) & (g820) & (!g773)) + ((!g321) & (g322) & (!g323) & (g324) & (g820) & (!g773)) + ((!g321) & (g322) & (!g323) & (g324) & (g820) & (g773)) + ((!g321) & (g322) & (g323) & (!g324) & (!g820) & (g773)) + ((!g321) & (g322) & (g323) & (!g324) & (g820) & (!g773)) + ((!g321) & (g322) & (g323) & (g324) & (!g820) & (g773)) + ((!g321) & (g322) & (g323) & (g324) & (g820) & (!g773)) + ((!g321) & (g322) & (g323) & (g324) & (g820) & (g773)) + ((g321) & (!g322) & (!g323) & (!g324) & (!g820) & (!g773)) + ((g321) & (!g322) & (!g323) & (g324) & (!g820) & (!g773)) + ((g321) & (!g322) & (!g323) & (g324) & (g820) & (g773)) + ((g321) & (!g322) & (g323) & (!g324) & (!g820) & (!g773)) + ((g321) & (!g322) & (g323) & (!g324) & (!g820) & (g773)) + ((g321) & (!g322) & (g323) & (g324) & (!g820) & (!g773)) + ((g321) & (!g322) & (g323) & (g324) & (!g820) & (g773)) + ((g321) & (!g322) & (g323) & (g324) & (g820) & (g773)) + ((g321) & (g322) & (!g323) & (!g324) & (!g820) & (!g773)) + ((g321) & (g322) & (!g323) & (!g324) & (g820) & (!g773)) + ((g321) & (g322) & (!g323) & (g324) & (!g820) & (!g773)) + ((g321) & (g322) & (!g323) & (g324) & (g820) & (!g773)) + ((g321) & (g322) & (!g323) & (g324) & (g820) & (g773)) + ((g321) & (g322) & (g323) & (!g324) & (!g820) & (!g773)) + ((g321) & (g322) & (g323) & (!g324) & (!g820) & (g773)) + ((g321) & (g322) & (g323) & (!g324) & (g820) & (!g773)) + ((g321) & (g322) & (g323) & (g324) & (!g820) & (!g773)) + ((g321) & (g322) & (g323) & (g324) & (!g820) & (g773)) + ((g321) & (g322) & (g323) & (g324) & (g820) & (!g773)) + ((g321) & (g322) & (g323) & (g324) & (g820) & (g773)));
	assign g1647 = (((!g326) & (!g327) & (!g328) & (g329) & (g820) & (g773)) + ((!g326) & (!g327) & (g328) & (!g329) & (!g820) & (g773)) + ((!g326) & (!g327) & (g328) & (g329) & (!g820) & (g773)) + ((!g326) & (!g327) & (g328) & (g329) & (g820) & (g773)) + ((!g326) & (g327) & (!g328) & (!g329) & (g820) & (!g773)) + ((!g326) & (g327) & (!g328) & (g329) & (g820) & (!g773)) + ((!g326) & (g327) & (!g328) & (g329) & (g820) & (g773)) + ((!g326) & (g327) & (g328) & (!g329) & (!g820) & (g773)) + ((!g326) & (g327) & (g328) & (!g329) & (g820) & (!g773)) + ((!g326) & (g327) & (g328) & (g329) & (!g820) & (g773)) + ((!g326) & (g327) & (g328) & (g329) & (g820) & (!g773)) + ((!g326) & (g327) & (g328) & (g329) & (g820) & (g773)) + ((g326) & (!g327) & (!g328) & (!g329) & (!g820) & (!g773)) + ((g326) & (!g327) & (!g328) & (g329) & (!g820) & (!g773)) + ((g326) & (!g327) & (!g328) & (g329) & (g820) & (g773)) + ((g326) & (!g327) & (g328) & (!g329) & (!g820) & (!g773)) + ((g326) & (!g327) & (g328) & (!g329) & (!g820) & (g773)) + ((g326) & (!g327) & (g328) & (g329) & (!g820) & (!g773)) + ((g326) & (!g327) & (g328) & (g329) & (!g820) & (g773)) + ((g326) & (!g327) & (g328) & (g329) & (g820) & (g773)) + ((g326) & (g327) & (!g328) & (!g329) & (!g820) & (!g773)) + ((g326) & (g327) & (!g328) & (!g329) & (g820) & (!g773)) + ((g326) & (g327) & (!g328) & (g329) & (!g820) & (!g773)) + ((g326) & (g327) & (!g328) & (g329) & (g820) & (!g773)) + ((g326) & (g327) & (!g328) & (g329) & (g820) & (g773)) + ((g326) & (g327) & (g328) & (!g329) & (!g820) & (!g773)) + ((g326) & (g327) & (g328) & (!g329) & (!g820) & (g773)) + ((g326) & (g327) & (g328) & (!g329) & (g820) & (!g773)) + ((g326) & (g327) & (g328) & (g329) & (!g820) & (!g773)) + ((g326) & (g327) & (g328) & (g329) & (!g820) & (g773)) + ((g326) & (g327) & (g328) & (g329) & (g820) & (!g773)) + ((g326) & (g327) & (g328) & (g329) & (g820) & (g773)));
	assign g1648 = (((!g331) & (!g332) & (!g333) & (g334) & (g820) & (g773)) + ((!g331) & (!g332) & (g333) & (!g334) & (!g820) & (g773)) + ((!g331) & (!g332) & (g333) & (g334) & (!g820) & (g773)) + ((!g331) & (!g332) & (g333) & (g334) & (g820) & (g773)) + ((!g331) & (g332) & (!g333) & (!g334) & (g820) & (!g773)) + ((!g331) & (g332) & (!g333) & (g334) & (g820) & (!g773)) + ((!g331) & (g332) & (!g333) & (g334) & (g820) & (g773)) + ((!g331) & (g332) & (g333) & (!g334) & (!g820) & (g773)) + ((!g331) & (g332) & (g333) & (!g334) & (g820) & (!g773)) + ((!g331) & (g332) & (g333) & (g334) & (!g820) & (g773)) + ((!g331) & (g332) & (g333) & (g334) & (g820) & (!g773)) + ((!g331) & (g332) & (g333) & (g334) & (g820) & (g773)) + ((g331) & (!g332) & (!g333) & (!g334) & (!g820) & (!g773)) + ((g331) & (!g332) & (!g333) & (g334) & (!g820) & (!g773)) + ((g331) & (!g332) & (!g333) & (g334) & (g820) & (g773)) + ((g331) & (!g332) & (g333) & (!g334) & (!g820) & (!g773)) + ((g331) & (!g332) & (g333) & (!g334) & (!g820) & (g773)) + ((g331) & (!g332) & (g333) & (g334) & (!g820) & (!g773)) + ((g331) & (!g332) & (g333) & (g334) & (!g820) & (g773)) + ((g331) & (!g332) & (g333) & (g334) & (g820) & (g773)) + ((g331) & (g332) & (!g333) & (!g334) & (!g820) & (!g773)) + ((g331) & (g332) & (!g333) & (!g334) & (g820) & (!g773)) + ((g331) & (g332) & (!g333) & (g334) & (!g820) & (!g773)) + ((g331) & (g332) & (!g333) & (g334) & (g820) & (!g773)) + ((g331) & (g332) & (!g333) & (g334) & (g820) & (g773)) + ((g331) & (g332) & (g333) & (!g334) & (!g820) & (!g773)) + ((g331) & (g332) & (g333) & (!g334) & (!g820) & (g773)) + ((g331) & (g332) & (g333) & (!g334) & (g820) & (!g773)) + ((g331) & (g332) & (g333) & (g334) & (!g820) & (!g773)) + ((g331) & (g332) & (g333) & (g334) & (!g820) & (g773)) + ((g331) & (g332) & (g333) & (g334) & (g820) & (!g773)) + ((g331) & (g332) & (g333) & (g334) & (g820) & (g773)));
	assign g1649 = (((!g336) & (!g337) & (!g338) & (g339) & (g820) & (g773)) + ((!g336) & (!g337) & (g338) & (!g339) & (!g820) & (g773)) + ((!g336) & (!g337) & (g338) & (g339) & (!g820) & (g773)) + ((!g336) & (!g337) & (g338) & (g339) & (g820) & (g773)) + ((!g336) & (g337) & (!g338) & (!g339) & (g820) & (!g773)) + ((!g336) & (g337) & (!g338) & (g339) & (g820) & (!g773)) + ((!g336) & (g337) & (!g338) & (g339) & (g820) & (g773)) + ((!g336) & (g337) & (g338) & (!g339) & (!g820) & (g773)) + ((!g336) & (g337) & (g338) & (!g339) & (g820) & (!g773)) + ((!g336) & (g337) & (g338) & (g339) & (!g820) & (g773)) + ((!g336) & (g337) & (g338) & (g339) & (g820) & (!g773)) + ((!g336) & (g337) & (g338) & (g339) & (g820) & (g773)) + ((g336) & (!g337) & (!g338) & (!g339) & (!g820) & (!g773)) + ((g336) & (!g337) & (!g338) & (g339) & (!g820) & (!g773)) + ((g336) & (!g337) & (!g338) & (g339) & (g820) & (g773)) + ((g336) & (!g337) & (g338) & (!g339) & (!g820) & (!g773)) + ((g336) & (!g337) & (g338) & (!g339) & (!g820) & (g773)) + ((g336) & (!g337) & (g338) & (g339) & (!g820) & (!g773)) + ((g336) & (!g337) & (g338) & (g339) & (!g820) & (g773)) + ((g336) & (!g337) & (g338) & (g339) & (g820) & (g773)) + ((g336) & (g337) & (!g338) & (!g339) & (!g820) & (!g773)) + ((g336) & (g337) & (!g338) & (!g339) & (g820) & (!g773)) + ((g336) & (g337) & (!g338) & (g339) & (!g820) & (!g773)) + ((g336) & (g337) & (!g338) & (g339) & (g820) & (!g773)) + ((g336) & (g337) & (!g338) & (g339) & (g820) & (g773)) + ((g336) & (g337) & (g338) & (!g339) & (!g820) & (!g773)) + ((g336) & (g337) & (g338) & (!g339) & (!g820) & (g773)) + ((g336) & (g337) & (g338) & (!g339) & (g820) & (!g773)) + ((g336) & (g337) & (g338) & (g339) & (!g820) & (!g773)) + ((g336) & (g337) & (g338) & (g339) & (!g820) & (g773)) + ((g336) & (g337) & (g338) & (g339) & (g820) & (!g773)) + ((g336) & (g337) & (g338) & (g339) & (g820) & (g773)));
	assign g1650 = (((!g1646) & (!g1647) & (!g1648) & (g1649) & (g677) & (g726)) + ((!g1646) & (!g1647) & (g1648) & (!g1649) & (!g677) & (g726)) + ((!g1646) & (!g1647) & (g1648) & (g1649) & (!g677) & (g726)) + ((!g1646) & (!g1647) & (g1648) & (g1649) & (g677) & (g726)) + ((!g1646) & (g1647) & (!g1648) & (!g1649) & (g677) & (!g726)) + ((!g1646) & (g1647) & (!g1648) & (g1649) & (g677) & (!g726)) + ((!g1646) & (g1647) & (!g1648) & (g1649) & (g677) & (g726)) + ((!g1646) & (g1647) & (g1648) & (!g1649) & (!g677) & (g726)) + ((!g1646) & (g1647) & (g1648) & (!g1649) & (g677) & (!g726)) + ((!g1646) & (g1647) & (g1648) & (g1649) & (!g677) & (g726)) + ((!g1646) & (g1647) & (g1648) & (g1649) & (g677) & (!g726)) + ((!g1646) & (g1647) & (g1648) & (g1649) & (g677) & (g726)) + ((g1646) & (!g1647) & (!g1648) & (!g1649) & (!g677) & (!g726)) + ((g1646) & (!g1647) & (!g1648) & (g1649) & (!g677) & (!g726)) + ((g1646) & (!g1647) & (!g1648) & (g1649) & (g677) & (g726)) + ((g1646) & (!g1647) & (g1648) & (!g1649) & (!g677) & (!g726)) + ((g1646) & (!g1647) & (g1648) & (!g1649) & (!g677) & (g726)) + ((g1646) & (!g1647) & (g1648) & (g1649) & (!g677) & (!g726)) + ((g1646) & (!g1647) & (g1648) & (g1649) & (!g677) & (g726)) + ((g1646) & (!g1647) & (g1648) & (g1649) & (g677) & (g726)) + ((g1646) & (g1647) & (!g1648) & (!g1649) & (!g677) & (!g726)) + ((g1646) & (g1647) & (!g1648) & (!g1649) & (g677) & (!g726)) + ((g1646) & (g1647) & (!g1648) & (g1649) & (!g677) & (!g726)) + ((g1646) & (g1647) & (!g1648) & (g1649) & (g677) & (!g726)) + ((g1646) & (g1647) & (!g1648) & (g1649) & (g677) & (g726)) + ((g1646) & (g1647) & (g1648) & (!g1649) & (!g677) & (!g726)) + ((g1646) & (g1647) & (g1648) & (!g1649) & (!g677) & (g726)) + ((g1646) & (g1647) & (g1648) & (!g1649) & (g677) & (!g726)) + ((g1646) & (g1647) & (g1648) & (g1649) & (!g677) & (!g726)) + ((g1646) & (g1647) & (g1648) & (g1649) & (!g677) & (g726)) + ((g1646) & (g1647) & (g1648) & (g1649) & (g677) & (!g726)) + ((g1646) & (g1647) & (g1648) & (g1649) & (g677) & (g726)));
	assign g1651 = (((!g342) & (!g343) & (!g344) & (g345) & (g677) & (g726)) + ((!g342) & (!g343) & (g344) & (!g345) & (!g677) & (g726)) + ((!g342) & (!g343) & (g344) & (g345) & (!g677) & (g726)) + ((!g342) & (!g343) & (g344) & (g345) & (g677) & (g726)) + ((!g342) & (g343) & (!g344) & (!g345) & (g677) & (!g726)) + ((!g342) & (g343) & (!g344) & (g345) & (g677) & (!g726)) + ((!g342) & (g343) & (!g344) & (g345) & (g677) & (g726)) + ((!g342) & (g343) & (g344) & (!g345) & (!g677) & (g726)) + ((!g342) & (g343) & (g344) & (!g345) & (g677) & (!g726)) + ((!g342) & (g343) & (g344) & (g345) & (!g677) & (g726)) + ((!g342) & (g343) & (g344) & (g345) & (g677) & (!g726)) + ((!g342) & (g343) & (g344) & (g345) & (g677) & (g726)) + ((g342) & (!g343) & (!g344) & (!g345) & (!g677) & (!g726)) + ((g342) & (!g343) & (!g344) & (g345) & (!g677) & (!g726)) + ((g342) & (!g343) & (!g344) & (g345) & (g677) & (g726)) + ((g342) & (!g343) & (g344) & (!g345) & (!g677) & (!g726)) + ((g342) & (!g343) & (g344) & (!g345) & (!g677) & (g726)) + ((g342) & (!g343) & (g344) & (g345) & (!g677) & (!g726)) + ((g342) & (!g343) & (g344) & (g345) & (!g677) & (g726)) + ((g342) & (!g343) & (g344) & (g345) & (g677) & (g726)) + ((g342) & (g343) & (!g344) & (!g345) & (!g677) & (!g726)) + ((g342) & (g343) & (!g344) & (!g345) & (g677) & (!g726)) + ((g342) & (g343) & (!g344) & (g345) & (!g677) & (!g726)) + ((g342) & (g343) & (!g344) & (g345) & (g677) & (!g726)) + ((g342) & (g343) & (!g344) & (g345) & (g677) & (g726)) + ((g342) & (g343) & (g344) & (!g345) & (!g677) & (!g726)) + ((g342) & (g343) & (g344) & (!g345) & (!g677) & (g726)) + ((g342) & (g343) & (g344) & (!g345) & (g677) & (!g726)) + ((g342) & (g343) & (g344) & (g345) & (!g677) & (!g726)) + ((g342) & (g343) & (g344) & (g345) & (!g677) & (g726)) + ((g342) & (g343) & (g344) & (g345) & (g677) & (!g726)) + ((g342) & (g343) & (g344) & (g345) & (g677) & (g726)));
	assign g1652 = (((!g677) & (!g726) & (!g347) & (g348) & (!sk[54]) & (!g349)) + ((!g677) & (!g726) & (!g347) & (g348) & (!sk[54]) & (g349)) + ((!g677) & (!g726) & (g347) & (!g348) & (!sk[54]) & (!g349)) + ((!g677) & (!g726) & (g347) & (!g348) & (!sk[54]) & (g349)) + ((!g677) & (!g726) & (g347) & (g348) & (!sk[54]) & (!g349)) + ((!g677) & (!g726) & (g347) & (g348) & (!sk[54]) & (g349)) + ((!g677) & (g726) & (!g347) & (!g348) & (!sk[54]) & (!g349)) + ((!g677) & (g726) & (!g347) & (!g348) & (!sk[54]) & (g349)) + ((!g677) & (g726) & (!g347) & (!g348) & (sk[54]) & (g349)) + ((!g677) & (g726) & (!g347) & (g348) & (!sk[54]) & (!g349)) + ((!g677) & (g726) & (!g347) & (g348) & (!sk[54]) & (g349)) + ((!g677) & (g726) & (!g347) & (g348) & (sk[54]) & (g349)) + ((!g677) & (g726) & (g347) & (!g348) & (!sk[54]) & (!g349)) + ((!g677) & (g726) & (g347) & (!g348) & (!sk[54]) & (g349)) + ((!g677) & (g726) & (g347) & (!g348) & (sk[54]) & (g349)) + ((!g677) & (g726) & (g347) & (g348) & (!sk[54]) & (!g349)) + ((!g677) & (g726) & (g347) & (g348) & (!sk[54]) & (g349)) + ((!g677) & (g726) & (g347) & (g348) & (sk[54]) & (g349)) + ((g677) & (!g726) & (!g347) & (g348) & (!sk[54]) & (!g349)) + ((g677) & (!g726) & (!g347) & (g348) & (!sk[54]) & (g349)) + ((g677) & (!g726) & (g347) & (!g348) & (!sk[54]) & (!g349)) + ((g677) & (!g726) & (g347) & (!g348) & (!sk[54]) & (g349)) + ((g677) & (!g726) & (g347) & (!g348) & (sk[54]) & (!g349)) + ((g677) & (!g726) & (g347) & (!g348) & (sk[54]) & (g349)) + ((g677) & (!g726) & (g347) & (g348) & (!sk[54]) & (!g349)) + ((g677) & (!g726) & (g347) & (g348) & (!sk[54]) & (g349)) + ((g677) & (!g726) & (g347) & (g348) & (sk[54]) & (!g349)) + ((g677) & (!g726) & (g347) & (g348) & (sk[54]) & (g349)) + ((g677) & (g726) & (!g347) & (!g348) & (!sk[54]) & (!g349)) + ((g677) & (g726) & (!g347) & (!g348) & (!sk[54]) & (g349)) + ((g677) & (g726) & (!g347) & (g348) & (!sk[54]) & (!g349)) + ((g677) & (g726) & (!g347) & (g348) & (!sk[54]) & (g349)) + ((g677) & (g726) & (!g347) & (g348) & (sk[54]) & (!g349)) + ((g677) & (g726) & (!g347) & (g348) & (sk[54]) & (g349)) + ((g677) & (g726) & (g347) & (!g348) & (!sk[54]) & (!g349)) + ((g677) & (g726) & (g347) & (!g348) & (!sk[54]) & (g349)) + ((g677) & (g726) & (g347) & (g348) & (!sk[54]) & (!g349)) + ((g677) & (g726) & (g347) & (g348) & (!sk[54]) & (g349)) + ((g677) & (g726) & (g347) & (g348) & (sk[54]) & (!g349)) + ((g677) & (g726) & (g347) & (g348) & (sk[54]) & (g349)));
	assign g1653 = (((!g351) & (!g352) & (!g353) & (g354) & (g677) & (g726)) + ((!g351) & (!g352) & (g353) & (!g354) & (!g677) & (g726)) + ((!g351) & (!g352) & (g353) & (g354) & (!g677) & (g726)) + ((!g351) & (!g352) & (g353) & (g354) & (g677) & (g726)) + ((!g351) & (g352) & (!g353) & (!g354) & (g677) & (!g726)) + ((!g351) & (g352) & (!g353) & (g354) & (g677) & (!g726)) + ((!g351) & (g352) & (!g353) & (g354) & (g677) & (g726)) + ((!g351) & (g352) & (g353) & (!g354) & (!g677) & (g726)) + ((!g351) & (g352) & (g353) & (!g354) & (g677) & (!g726)) + ((!g351) & (g352) & (g353) & (g354) & (!g677) & (g726)) + ((!g351) & (g352) & (g353) & (g354) & (g677) & (!g726)) + ((!g351) & (g352) & (g353) & (g354) & (g677) & (g726)) + ((g351) & (!g352) & (!g353) & (!g354) & (!g677) & (!g726)) + ((g351) & (!g352) & (!g353) & (g354) & (!g677) & (!g726)) + ((g351) & (!g352) & (!g353) & (g354) & (g677) & (g726)) + ((g351) & (!g352) & (g353) & (!g354) & (!g677) & (!g726)) + ((g351) & (!g352) & (g353) & (!g354) & (!g677) & (g726)) + ((g351) & (!g352) & (g353) & (g354) & (!g677) & (!g726)) + ((g351) & (!g352) & (g353) & (g354) & (!g677) & (g726)) + ((g351) & (!g352) & (g353) & (g354) & (g677) & (g726)) + ((g351) & (g352) & (!g353) & (!g354) & (!g677) & (!g726)) + ((g351) & (g352) & (!g353) & (!g354) & (g677) & (!g726)) + ((g351) & (g352) & (!g353) & (g354) & (!g677) & (!g726)) + ((g351) & (g352) & (!g353) & (g354) & (g677) & (!g726)) + ((g351) & (g352) & (!g353) & (g354) & (g677) & (g726)) + ((g351) & (g352) & (g353) & (!g354) & (!g677) & (!g726)) + ((g351) & (g352) & (g353) & (!g354) & (!g677) & (g726)) + ((g351) & (g352) & (g353) & (!g354) & (g677) & (!g726)) + ((g351) & (g352) & (g353) & (g354) & (!g677) & (!g726)) + ((g351) & (g352) & (g353) & (g354) & (!g677) & (g726)) + ((g351) & (g352) & (g353) & (g354) & (g677) & (!g726)) + ((g351) & (g352) & (g353) & (g354) & (g677) & (g726)));
	assign g1654 = (((!g356) & (!g357) & (!g358) & (g359) & (g677) & (g726)) + ((!g356) & (!g357) & (g358) & (!g359) & (!g677) & (g726)) + ((!g356) & (!g357) & (g358) & (g359) & (!g677) & (g726)) + ((!g356) & (!g357) & (g358) & (g359) & (g677) & (g726)) + ((!g356) & (g357) & (!g358) & (!g359) & (g677) & (!g726)) + ((!g356) & (g357) & (!g358) & (g359) & (g677) & (!g726)) + ((!g356) & (g357) & (!g358) & (g359) & (g677) & (g726)) + ((!g356) & (g357) & (g358) & (!g359) & (!g677) & (g726)) + ((!g356) & (g357) & (g358) & (!g359) & (g677) & (!g726)) + ((!g356) & (g357) & (g358) & (g359) & (!g677) & (g726)) + ((!g356) & (g357) & (g358) & (g359) & (g677) & (!g726)) + ((!g356) & (g357) & (g358) & (g359) & (g677) & (g726)) + ((g356) & (!g357) & (!g358) & (!g359) & (!g677) & (!g726)) + ((g356) & (!g357) & (!g358) & (g359) & (!g677) & (!g726)) + ((g356) & (!g357) & (!g358) & (g359) & (g677) & (g726)) + ((g356) & (!g357) & (g358) & (!g359) & (!g677) & (!g726)) + ((g356) & (!g357) & (g358) & (!g359) & (!g677) & (g726)) + ((g356) & (!g357) & (g358) & (g359) & (!g677) & (!g726)) + ((g356) & (!g357) & (g358) & (g359) & (!g677) & (g726)) + ((g356) & (!g357) & (g358) & (g359) & (g677) & (g726)) + ((g356) & (g357) & (!g358) & (!g359) & (!g677) & (!g726)) + ((g356) & (g357) & (!g358) & (!g359) & (g677) & (!g726)) + ((g356) & (g357) & (!g358) & (g359) & (!g677) & (!g726)) + ((g356) & (g357) & (!g358) & (g359) & (g677) & (!g726)) + ((g356) & (g357) & (!g358) & (g359) & (g677) & (g726)) + ((g356) & (g357) & (g358) & (!g359) & (!g677) & (!g726)) + ((g356) & (g357) & (g358) & (!g359) & (!g677) & (g726)) + ((g356) & (g357) & (g358) & (!g359) & (g677) & (!g726)) + ((g356) & (g357) & (g358) & (g359) & (!g677) & (!g726)) + ((g356) & (g357) & (g358) & (g359) & (!g677) & (g726)) + ((g356) & (g357) & (g358) & (g359) & (g677) & (!g726)) + ((g356) & (g357) & (g358) & (g359) & (g677) & (g726)));
	assign g1655 = (((!g820) & (!g773) & (!g1651) & (g1652) & (!g1653) & (!g1654)) + ((!g820) & (!g773) & (!g1651) & (g1652) & (!g1653) & (g1654)) + ((!g820) & (!g773) & (!g1651) & (g1652) & (g1653) & (!g1654)) + ((!g820) & (!g773) & (!g1651) & (g1652) & (g1653) & (g1654)) + ((!g820) & (!g773) & (g1651) & (g1652) & (!g1653) & (!g1654)) + ((!g820) & (!g773) & (g1651) & (g1652) & (!g1653) & (g1654)) + ((!g820) & (!g773) & (g1651) & (g1652) & (g1653) & (!g1654)) + ((!g820) & (!g773) & (g1651) & (g1652) & (g1653) & (g1654)) + ((!g820) & (g773) & (!g1651) & (!g1652) & (!g1653) & (g1654)) + ((!g820) & (g773) & (!g1651) & (!g1652) & (g1653) & (g1654)) + ((!g820) & (g773) & (!g1651) & (g1652) & (!g1653) & (g1654)) + ((!g820) & (g773) & (!g1651) & (g1652) & (g1653) & (g1654)) + ((!g820) & (g773) & (g1651) & (!g1652) & (!g1653) & (g1654)) + ((!g820) & (g773) & (g1651) & (!g1652) & (g1653) & (g1654)) + ((!g820) & (g773) & (g1651) & (g1652) & (!g1653) & (g1654)) + ((!g820) & (g773) & (g1651) & (g1652) & (g1653) & (g1654)) + ((g820) & (!g773) & (g1651) & (!g1652) & (!g1653) & (!g1654)) + ((g820) & (!g773) & (g1651) & (!g1652) & (!g1653) & (g1654)) + ((g820) & (!g773) & (g1651) & (!g1652) & (g1653) & (!g1654)) + ((g820) & (!g773) & (g1651) & (!g1652) & (g1653) & (g1654)) + ((g820) & (!g773) & (g1651) & (g1652) & (!g1653) & (!g1654)) + ((g820) & (!g773) & (g1651) & (g1652) & (!g1653) & (g1654)) + ((g820) & (!g773) & (g1651) & (g1652) & (g1653) & (!g1654)) + ((g820) & (!g773) & (g1651) & (g1652) & (g1653) & (g1654)) + ((g820) & (g773) & (!g1651) & (!g1652) & (g1653) & (!g1654)) + ((g820) & (g773) & (!g1651) & (!g1652) & (g1653) & (g1654)) + ((g820) & (g773) & (!g1651) & (g1652) & (g1653) & (!g1654)) + ((g820) & (g773) & (!g1651) & (g1652) & (g1653) & (g1654)) + ((g820) & (g773) & (g1651) & (!g1652) & (g1653) & (!g1654)) + ((g820) & (g773) & (g1651) & (!g1652) & (g1653) & (g1654)) + ((g820) & (g773) & (g1651) & (g1652) & (g1653) & (!g1654)) + ((g820) & (g773) & (g1651) & (g1652) & (g1653) & (g1654)));
	assign g1656 = (((!g867) & (!g1650) & (!sk[58]) & (g1655)) + ((!g867) & (!g1650) & (sk[58]) & (g1655)) + ((!g867) & (g1650) & (!sk[58]) & (!g1655)) + ((!g867) & (g1650) & (!sk[58]) & (g1655)) + ((!g867) & (g1650) & (sk[58]) & (g1655)) + ((g867) & (!g1650) & (!sk[58]) & (g1655)) + ((g867) & (g1650) & (!sk[58]) & (!g1655)) + ((g867) & (g1650) & (!sk[58]) & (g1655)) + ((g867) & (g1650) & (sk[58]) & (!g1655)) + ((g867) & (g1650) & (sk[58]) & (g1655)));
	assign g1657 = (((!g1592) & (!g1593) & (!g1605) & (g1607) & (!g39) & (g1656)) + ((!g1592) & (!g1593) & (!g1605) & (g1607) & (g39) & (g1656)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (!g39) & (g1656)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (g39) & (g1656)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (!g39) & (g1656)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (g39) & (g1656)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (!g39) & (g1656)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (g39) & (g1656)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (!g39) & (g1656)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (g39) & (g1656)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g39) & (!g1656)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g39) & (g1656)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g39) & (!g1656)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g39) & (g1656)));
	assign g1658 = (((!g366) & (!g371) & (!g376) & (g381) & (g820) & (g773)) + ((!g366) & (!g371) & (g376) & (!g381) & (!g820) & (g773)) + ((!g366) & (!g371) & (g376) & (g381) & (!g820) & (g773)) + ((!g366) & (!g371) & (g376) & (g381) & (g820) & (g773)) + ((!g366) & (g371) & (!g376) & (!g381) & (g820) & (!g773)) + ((!g366) & (g371) & (!g376) & (g381) & (g820) & (!g773)) + ((!g366) & (g371) & (!g376) & (g381) & (g820) & (g773)) + ((!g366) & (g371) & (g376) & (!g381) & (!g820) & (g773)) + ((!g366) & (g371) & (g376) & (!g381) & (g820) & (!g773)) + ((!g366) & (g371) & (g376) & (g381) & (!g820) & (g773)) + ((!g366) & (g371) & (g376) & (g381) & (g820) & (!g773)) + ((!g366) & (g371) & (g376) & (g381) & (g820) & (g773)) + ((g366) & (!g371) & (!g376) & (!g381) & (!g820) & (!g773)) + ((g366) & (!g371) & (!g376) & (g381) & (!g820) & (!g773)) + ((g366) & (!g371) & (!g376) & (g381) & (g820) & (g773)) + ((g366) & (!g371) & (g376) & (!g381) & (!g820) & (!g773)) + ((g366) & (!g371) & (g376) & (!g381) & (!g820) & (g773)) + ((g366) & (!g371) & (g376) & (g381) & (!g820) & (!g773)) + ((g366) & (!g371) & (g376) & (g381) & (!g820) & (g773)) + ((g366) & (!g371) & (g376) & (g381) & (g820) & (g773)) + ((g366) & (g371) & (!g376) & (!g381) & (!g820) & (!g773)) + ((g366) & (g371) & (!g376) & (!g381) & (g820) & (!g773)) + ((g366) & (g371) & (!g376) & (g381) & (!g820) & (!g773)) + ((g366) & (g371) & (!g376) & (g381) & (g820) & (!g773)) + ((g366) & (g371) & (!g376) & (g381) & (g820) & (g773)) + ((g366) & (g371) & (g376) & (!g381) & (!g820) & (!g773)) + ((g366) & (g371) & (g376) & (!g381) & (!g820) & (g773)) + ((g366) & (g371) & (g376) & (!g381) & (g820) & (!g773)) + ((g366) & (g371) & (g376) & (g381) & (!g820) & (!g773)) + ((g366) & (g371) & (g376) & (g381) & (!g820) & (g773)) + ((g366) & (g371) & (g376) & (g381) & (g820) & (!g773)) + ((g366) & (g371) & (g376) & (g381) & (g820) & (g773)));
	assign g1659 = (((!g367) & (!g372) & (!g377) & (g382) & (g820) & (g773)) + ((!g367) & (!g372) & (g377) & (!g382) & (!g820) & (g773)) + ((!g367) & (!g372) & (g377) & (g382) & (!g820) & (g773)) + ((!g367) & (!g372) & (g377) & (g382) & (g820) & (g773)) + ((!g367) & (g372) & (!g377) & (!g382) & (g820) & (!g773)) + ((!g367) & (g372) & (!g377) & (g382) & (g820) & (!g773)) + ((!g367) & (g372) & (!g377) & (g382) & (g820) & (g773)) + ((!g367) & (g372) & (g377) & (!g382) & (!g820) & (g773)) + ((!g367) & (g372) & (g377) & (!g382) & (g820) & (!g773)) + ((!g367) & (g372) & (g377) & (g382) & (!g820) & (g773)) + ((!g367) & (g372) & (g377) & (g382) & (g820) & (!g773)) + ((!g367) & (g372) & (g377) & (g382) & (g820) & (g773)) + ((g367) & (!g372) & (!g377) & (!g382) & (!g820) & (!g773)) + ((g367) & (!g372) & (!g377) & (g382) & (!g820) & (!g773)) + ((g367) & (!g372) & (!g377) & (g382) & (g820) & (g773)) + ((g367) & (!g372) & (g377) & (!g382) & (!g820) & (!g773)) + ((g367) & (!g372) & (g377) & (!g382) & (!g820) & (g773)) + ((g367) & (!g372) & (g377) & (g382) & (!g820) & (!g773)) + ((g367) & (!g372) & (g377) & (g382) & (!g820) & (g773)) + ((g367) & (!g372) & (g377) & (g382) & (g820) & (g773)) + ((g367) & (g372) & (!g377) & (!g382) & (!g820) & (!g773)) + ((g367) & (g372) & (!g377) & (!g382) & (g820) & (!g773)) + ((g367) & (g372) & (!g377) & (g382) & (!g820) & (!g773)) + ((g367) & (g372) & (!g377) & (g382) & (g820) & (!g773)) + ((g367) & (g372) & (!g377) & (g382) & (g820) & (g773)) + ((g367) & (g372) & (g377) & (!g382) & (!g820) & (!g773)) + ((g367) & (g372) & (g377) & (!g382) & (!g820) & (g773)) + ((g367) & (g372) & (g377) & (!g382) & (g820) & (!g773)) + ((g367) & (g372) & (g377) & (g382) & (!g820) & (!g773)) + ((g367) & (g372) & (g377) & (g382) & (!g820) & (g773)) + ((g367) & (g372) & (g377) & (g382) & (g820) & (!g773)) + ((g367) & (g372) & (g377) & (g382) & (g820) & (g773)));
	assign g1660 = (((!g368) & (!g373) & (!g378) & (g383) & (g820) & (g773)) + ((!g368) & (!g373) & (g378) & (!g383) & (!g820) & (g773)) + ((!g368) & (!g373) & (g378) & (g383) & (!g820) & (g773)) + ((!g368) & (!g373) & (g378) & (g383) & (g820) & (g773)) + ((!g368) & (g373) & (!g378) & (!g383) & (g820) & (!g773)) + ((!g368) & (g373) & (!g378) & (g383) & (g820) & (!g773)) + ((!g368) & (g373) & (!g378) & (g383) & (g820) & (g773)) + ((!g368) & (g373) & (g378) & (!g383) & (!g820) & (g773)) + ((!g368) & (g373) & (g378) & (!g383) & (g820) & (!g773)) + ((!g368) & (g373) & (g378) & (g383) & (!g820) & (g773)) + ((!g368) & (g373) & (g378) & (g383) & (g820) & (!g773)) + ((!g368) & (g373) & (g378) & (g383) & (g820) & (g773)) + ((g368) & (!g373) & (!g378) & (!g383) & (!g820) & (!g773)) + ((g368) & (!g373) & (!g378) & (g383) & (!g820) & (!g773)) + ((g368) & (!g373) & (!g378) & (g383) & (g820) & (g773)) + ((g368) & (!g373) & (g378) & (!g383) & (!g820) & (!g773)) + ((g368) & (!g373) & (g378) & (!g383) & (!g820) & (g773)) + ((g368) & (!g373) & (g378) & (g383) & (!g820) & (!g773)) + ((g368) & (!g373) & (g378) & (g383) & (!g820) & (g773)) + ((g368) & (!g373) & (g378) & (g383) & (g820) & (g773)) + ((g368) & (g373) & (!g378) & (!g383) & (!g820) & (!g773)) + ((g368) & (g373) & (!g378) & (!g383) & (g820) & (!g773)) + ((g368) & (g373) & (!g378) & (g383) & (!g820) & (!g773)) + ((g368) & (g373) & (!g378) & (g383) & (g820) & (!g773)) + ((g368) & (g373) & (!g378) & (g383) & (g820) & (g773)) + ((g368) & (g373) & (g378) & (!g383) & (!g820) & (!g773)) + ((g368) & (g373) & (g378) & (!g383) & (!g820) & (g773)) + ((g368) & (g373) & (g378) & (!g383) & (g820) & (!g773)) + ((g368) & (g373) & (g378) & (g383) & (!g820) & (!g773)) + ((g368) & (g373) & (g378) & (g383) & (!g820) & (g773)) + ((g368) & (g373) & (g378) & (g383) & (g820) & (!g773)) + ((g368) & (g373) & (g378) & (g383) & (g820) & (g773)));
	assign g1661 = (((!g369) & (!g374) & (!g379) & (g384) & (g820) & (g773)) + ((!g369) & (!g374) & (g379) & (!g384) & (!g820) & (g773)) + ((!g369) & (!g374) & (g379) & (g384) & (!g820) & (g773)) + ((!g369) & (!g374) & (g379) & (g384) & (g820) & (g773)) + ((!g369) & (g374) & (!g379) & (!g384) & (g820) & (!g773)) + ((!g369) & (g374) & (!g379) & (g384) & (g820) & (!g773)) + ((!g369) & (g374) & (!g379) & (g384) & (g820) & (g773)) + ((!g369) & (g374) & (g379) & (!g384) & (!g820) & (g773)) + ((!g369) & (g374) & (g379) & (!g384) & (g820) & (!g773)) + ((!g369) & (g374) & (g379) & (g384) & (!g820) & (g773)) + ((!g369) & (g374) & (g379) & (g384) & (g820) & (!g773)) + ((!g369) & (g374) & (g379) & (g384) & (g820) & (g773)) + ((g369) & (!g374) & (!g379) & (!g384) & (!g820) & (!g773)) + ((g369) & (!g374) & (!g379) & (g384) & (!g820) & (!g773)) + ((g369) & (!g374) & (!g379) & (g384) & (g820) & (g773)) + ((g369) & (!g374) & (g379) & (!g384) & (!g820) & (!g773)) + ((g369) & (!g374) & (g379) & (!g384) & (!g820) & (g773)) + ((g369) & (!g374) & (g379) & (g384) & (!g820) & (!g773)) + ((g369) & (!g374) & (g379) & (g384) & (!g820) & (g773)) + ((g369) & (!g374) & (g379) & (g384) & (g820) & (g773)) + ((g369) & (g374) & (!g379) & (!g384) & (!g820) & (!g773)) + ((g369) & (g374) & (!g379) & (!g384) & (g820) & (!g773)) + ((g369) & (g374) & (!g379) & (g384) & (!g820) & (!g773)) + ((g369) & (g374) & (!g379) & (g384) & (g820) & (!g773)) + ((g369) & (g374) & (!g379) & (g384) & (g820) & (g773)) + ((g369) & (g374) & (g379) & (!g384) & (!g820) & (!g773)) + ((g369) & (g374) & (g379) & (!g384) & (!g820) & (g773)) + ((g369) & (g374) & (g379) & (!g384) & (g820) & (!g773)) + ((g369) & (g374) & (g379) & (g384) & (!g820) & (!g773)) + ((g369) & (g374) & (g379) & (g384) & (!g820) & (g773)) + ((g369) & (g374) & (g379) & (g384) & (g820) & (!g773)) + ((g369) & (g374) & (g379) & (g384) & (g820) & (g773)));
	assign g1662 = (((!g1658) & (!g1659) & (!g1660) & (g1661) & (g677) & (g726)) + ((!g1658) & (!g1659) & (g1660) & (!g1661) & (!g677) & (g726)) + ((!g1658) & (!g1659) & (g1660) & (g1661) & (!g677) & (g726)) + ((!g1658) & (!g1659) & (g1660) & (g1661) & (g677) & (g726)) + ((!g1658) & (g1659) & (!g1660) & (!g1661) & (g677) & (!g726)) + ((!g1658) & (g1659) & (!g1660) & (g1661) & (g677) & (!g726)) + ((!g1658) & (g1659) & (!g1660) & (g1661) & (g677) & (g726)) + ((!g1658) & (g1659) & (g1660) & (!g1661) & (!g677) & (g726)) + ((!g1658) & (g1659) & (g1660) & (!g1661) & (g677) & (!g726)) + ((!g1658) & (g1659) & (g1660) & (g1661) & (!g677) & (g726)) + ((!g1658) & (g1659) & (g1660) & (g1661) & (g677) & (!g726)) + ((!g1658) & (g1659) & (g1660) & (g1661) & (g677) & (g726)) + ((g1658) & (!g1659) & (!g1660) & (!g1661) & (!g677) & (!g726)) + ((g1658) & (!g1659) & (!g1660) & (g1661) & (!g677) & (!g726)) + ((g1658) & (!g1659) & (!g1660) & (g1661) & (g677) & (g726)) + ((g1658) & (!g1659) & (g1660) & (!g1661) & (!g677) & (!g726)) + ((g1658) & (!g1659) & (g1660) & (!g1661) & (!g677) & (g726)) + ((g1658) & (!g1659) & (g1660) & (g1661) & (!g677) & (!g726)) + ((g1658) & (!g1659) & (g1660) & (g1661) & (!g677) & (g726)) + ((g1658) & (!g1659) & (g1660) & (g1661) & (g677) & (g726)) + ((g1658) & (g1659) & (!g1660) & (!g1661) & (!g677) & (!g726)) + ((g1658) & (g1659) & (!g1660) & (!g1661) & (g677) & (!g726)) + ((g1658) & (g1659) & (!g1660) & (g1661) & (!g677) & (!g726)) + ((g1658) & (g1659) & (!g1660) & (g1661) & (g677) & (!g726)) + ((g1658) & (g1659) & (!g1660) & (g1661) & (g677) & (g726)) + ((g1658) & (g1659) & (g1660) & (!g1661) & (!g677) & (!g726)) + ((g1658) & (g1659) & (g1660) & (!g1661) & (!g677) & (g726)) + ((g1658) & (g1659) & (g1660) & (!g1661) & (g677) & (!g726)) + ((g1658) & (g1659) & (g1660) & (g1661) & (!g677) & (!g726)) + ((g1658) & (g1659) & (g1660) & (g1661) & (!g677) & (g726)) + ((g1658) & (g1659) & (g1660) & (g1661) & (g677) & (!g726)) + ((g1658) & (g1659) & (g1660) & (g1661) & (g677) & (g726)));
	assign g1663 = (((!g387) & (!g388) & (!g389) & (g390) & (g677) & (g726)) + ((!g387) & (!g388) & (g389) & (!g390) & (!g677) & (g726)) + ((!g387) & (!g388) & (g389) & (g390) & (!g677) & (g726)) + ((!g387) & (!g388) & (g389) & (g390) & (g677) & (g726)) + ((!g387) & (g388) & (!g389) & (!g390) & (g677) & (!g726)) + ((!g387) & (g388) & (!g389) & (g390) & (g677) & (!g726)) + ((!g387) & (g388) & (!g389) & (g390) & (g677) & (g726)) + ((!g387) & (g388) & (g389) & (!g390) & (!g677) & (g726)) + ((!g387) & (g388) & (g389) & (!g390) & (g677) & (!g726)) + ((!g387) & (g388) & (g389) & (g390) & (!g677) & (g726)) + ((!g387) & (g388) & (g389) & (g390) & (g677) & (!g726)) + ((!g387) & (g388) & (g389) & (g390) & (g677) & (g726)) + ((g387) & (!g388) & (!g389) & (!g390) & (!g677) & (!g726)) + ((g387) & (!g388) & (!g389) & (g390) & (!g677) & (!g726)) + ((g387) & (!g388) & (!g389) & (g390) & (g677) & (g726)) + ((g387) & (!g388) & (g389) & (!g390) & (!g677) & (!g726)) + ((g387) & (!g388) & (g389) & (!g390) & (!g677) & (g726)) + ((g387) & (!g388) & (g389) & (g390) & (!g677) & (!g726)) + ((g387) & (!g388) & (g389) & (g390) & (!g677) & (g726)) + ((g387) & (!g388) & (g389) & (g390) & (g677) & (g726)) + ((g387) & (g388) & (!g389) & (!g390) & (!g677) & (!g726)) + ((g387) & (g388) & (!g389) & (!g390) & (g677) & (!g726)) + ((g387) & (g388) & (!g389) & (g390) & (!g677) & (!g726)) + ((g387) & (g388) & (!g389) & (g390) & (g677) & (!g726)) + ((g387) & (g388) & (!g389) & (g390) & (g677) & (g726)) + ((g387) & (g388) & (g389) & (!g390) & (!g677) & (!g726)) + ((g387) & (g388) & (g389) & (!g390) & (!g677) & (g726)) + ((g387) & (g388) & (g389) & (!g390) & (g677) & (!g726)) + ((g387) & (g388) & (g389) & (g390) & (!g677) & (!g726)) + ((g387) & (g388) & (g389) & (g390) & (!g677) & (g726)) + ((g387) & (g388) & (g389) & (g390) & (g677) & (!g726)) + ((g387) & (g388) & (g389) & (g390) & (g677) & (g726)));
	assign g1664 = (((!g677) & (!sk[66]) & (!g726) & (!g392) & (g393) & (!g394)) + ((!g677) & (!sk[66]) & (!g726) & (!g392) & (g393) & (g394)) + ((!g677) & (!sk[66]) & (!g726) & (g392) & (!g393) & (!g394)) + ((!g677) & (!sk[66]) & (!g726) & (g392) & (!g393) & (g394)) + ((!g677) & (!sk[66]) & (!g726) & (g392) & (g393) & (!g394)) + ((!g677) & (!sk[66]) & (!g726) & (g392) & (g393) & (g394)) + ((!g677) & (!sk[66]) & (g726) & (!g392) & (!g393) & (!g394)) + ((!g677) & (!sk[66]) & (g726) & (!g392) & (!g393) & (g394)) + ((!g677) & (!sk[66]) & (g726) & (!g392) & (g393) & (!g394)) + ((!g677) & (!sk[66]) & (g726) & (!g392) & (g393) & (g394)) + ((!g677) & (!sk[66]) & (g726) & (g392) & (!g393) & (!g394)) + ((!g677) & (!sk[66]) & (g726) & (g392) & (!g393) & (g394)) + ((!g677) & (!sk[66]) & (g726) & (g392) & (g393) & (!g394)) + ((!g677) & (!sk[66]) & (g726) & (g392) & (g393) & (g394)) + ((!g677) & (sk[66]) & (g726) & (!g392) & (!g393) & (g394)) + ((!g677) & (sk[66]) & (g726) & (!g392) & (g393) & (g394)) + ((!g677) & (sk[66]) & (g726) & (g392) & (!g393) & (g394)) + ((!g677) & (sk[66]) & (g726) & (g392) & (g393) & (g394)) + ((g677) & (!sk[66]) & (!g726) & (!g392) & (g393) & (!g394)) + ((g677) & (!sk[66]) & (!g726) & (!g392) & (g393) & (g394)) + ((g677) & (!sk[66]) & (!g726) & (g392) & (!g393) & (!g394)) + ((g677) & (!sk[66]) & (!g726) & (g392) & (!g393) & (g394)) + ((g677) & (!sk[66]) & (!g726) & (g392) & (g393) & (!g394)) + ((g677) & (!sk[66]) & (!g726) & (g392) & (g393) & (g394)) + ((g677) & (!sk[66]) & (g726) & (!g392) & (!g393) & (!g394)) + ((g677) & (!sk[66]) & (g726) & (!g392) & (!g393) & (g394)) + ((g677) & (!sk[66]) & (g726) & (!g392) & (g393) & (!g394)) + ((g677) & (!sk[66]) & (g726) & (!g392) & (g393) & (g394)) + ((g677) & (!sk[66]) & (g726) & (g392) & (!g393) & (!g394)) + ((g677) & (!sk[66]) & (g726) & (g392) & (!g393) & (g394)) + ((g677) & (!sk[66]) & (g726) & (g392) & (g393) & (!g394)) + ((g677) & (!sk[66]) & (g726) & (g392) & (g393) & (g394)) + ((g677) & (sk[66]) & (!g726) & (g392) & (!g393) & (!g394)) + ((g677) & (sk[66]) & (!g726) & (g392) & (!g393) & (g394)) + ((g677) & (sk[66]) & (!g726) & (g392) & (g393) & (!g394)) + ((g677) & (sk[66]) & (!g726) & (g392) & (g393) & (g394)) + ((g677) & (sk[66]) & (g726) & (!g392) & (g393) & (!g394)) + ((g677) & (sk[66]) & (g726) & (!g392) & (g393) & (g394)) + ((g677) & (sk[66]) & (g726) & (g392) & (g393) & (!g394)) + ((g677) & (sk[66]) & (g726) & (g392) & (g393) & (g394)));
	assign g1665 = (((!g396) & (!g397) & (!g398) & (g399) & (g677) & (g726)) + ((!g396) & (!g397) & (g398) & (!g399) & (!g677) & (g726)) + ((!g396) & (!g397) & (g398) & (g399) & (!g677) & (g726)) + ((!g396) & (!g397) & (g398) & (g399) & (g677) & (g726)) + ((!g396) & (g397) & (!g398) & (!g399) & (g677) & (!g726)) + ((!g396) & (g397) & (!g398) & (g399) & (g677) & (!g726)) + ((!g396) & (g397) & (!g398) & (g399) & (g677) & (g726)) + ((!g396) & (g397) & (g398) & (!g399) & (!g677) & (g726)) + ((!g396) & (g397) & (g398) & (!g399) & (g677) & (!g726)) + ((!g396) & (g397) & (g398) & (g399) & (!g677) & (g726)) + ((!g396) & (g397) & (g398) & (g399) & (g677) & (!g726)) + ((!g396) & (g397) & (g398) & (g399) & (g677) & (g726)) + ((g396) & (!g397) & (!g398) & (!g399) & (!g677) & (!g726)) + ((g396) & (!g397) & (!g398) & (g399) & (!g677) & (!g726)) + ((g396) & (!g397) & (!g398) & (g399) & (g677) & (g726)) + ((g396) & (!g397) & (g398) & (!g399) & (!g677) & (!g726)) + ((g396) & (!g397) & (g398) & (!g399) & (!g677) & (g726)) + ((g396) & (!g397) & (g398) & (g399) & (!g677) & (!g726)) + ((g396) & (!g397) & (g398) & (g399) & (!g677) & (g726)) + ((g396) & (!g397) & (g398) & (g399) & (g677) & (g726)) + ((g396) & (g397) & (!g398) & (!g399) & (!g677) & (!g726)) + ((g396) & (g397) & (!g398) & (!g399) & (g677) & (!g726)) + ((g396) & (g397) & (!g398) & (g399) & (!g677) & (!g726)) + ((g396) & (g397) & (!g398) & (g399) & (g677) & (!g726)) + ((g396) & (g397) & (!g398) & (g399) & (g677) & (g726)) + ((g396) & (g397) & (g398) & (!g399) & (!g677) & (!g726)) + ((g396) & (g397) & (g398) & (!g399) & (!g677) & (g726)) + ((g396) & (g397) & (g398) & (!g399) & (g677) & (!g726)) + ((g396) & (g397) & (g398) & (g399) & (!g677) & (!g726)) + ((g396) & (g397) & (g398) & (g399) & (!g677) & (g726)) + ((g396) & (g397) & (g398) & (g399) & (g677) & (!g726)) + ((g396) & (g397) & (g398) & (g399) & (g677) & (g726)));
	assign g1666 = (((!g401) & (!g402) & (!g403) & (g404) & (g677) & (g726)) + ((!g401) & (!g402) & (g403) & (!g404) & (!g677) & (g726)) + ((!g401) & (!g402) & (g403) & (g404) & (!g677) & (g726)) + ((!g401) & (!g402) & (g403) & (g404) & (g677) & (g726)) + ((!g401) & (g402) & (!g403) & (!g404) & (g677) & (!g726)) + ((!g401) & (g402) & (!g403) & (g404) & (g677) & (!g726)) + ((!g401) & (g402) & (!g403) & (g404) & (g677) & (g726)) + ((!g401) & (g402) & (g403) & (!g404) & (!g677) & (g726)) + ((!g401) & (g402) & (g403) & (!g404) & (g677) & (!g726)) + ((!g401) & (g402) & (g403) & (g404) & (!g677) & (g726)) + ((!g401) & (g402) & (g403) & (g404) & (g677) & (!g726)) + ((!g401) & (g402) & (g403) & (g404) & (g677) & (g726)) + ((g401) & (!g402) & (!g403) & (!g404) & (!g677) & (!g726)) + ((g401) & (!g402) & (!g403) & (g404) & (!g677) & (!g726)) + ((g401) & (!g402) & (!g403) & (g404) & (g677) & (g726)) + ((g401) & (!g402) & (g403) & (!g404) & (!g677) & (!g726)) + ((g401) & (!g402) & (g403) & (!g404) & (!g677) & (g726)) + ((g401) & (!g402) & (g403) & (g404) & (!g677) & (!g726)) + ((g401) & (!g402) & (g403) & (g404) & (!g677) & (g726)) + ((g401) & (!g402) & (g403) & (g404) & (g677) & (g726)) + ((g401) & (g402) & (!g403) & (!g404) & (!g677) & (!g726)) + ((g401) & (g402) & (!g403) & (!g404) & (g677) & (!g726)) + ((g401) & (g402) & (!g403) & (g404) & (!g677) & (!g726)) + ((g401) & (g402) & (!g403) & (g404) & (g677) & (!g726)) + ((g401) & (g402) & (!g403) & (g404) & (g677) & (g726)) + ((g401) & (g402) & (g403) & (!g404) & (!g677) & (!g726)) + ((g401) & (g402) & (g403) & (!g404) & (!g677) & (g726)) + ((g401) & (g402) & (g403) & (!g404) & (g677) & (!g726)) + ((g401) & (g402) & (g403) & (g404) & (!g677) & (!g726)) + ((g401) & (g402) & (g403) & (g404) & (!g677) & (g726)) + ((g401) & (g402) & (g403) & (g404) & (g677) & (!g726)) + ((g401) & (g402) & (g403) & (g404) & (g677) & (g726)));
	assign g1667 = (((!g820) & (!g773) & (!g1663) & (g1664) & (!g1665) & (!g1666)) + ((!g820) & (!g773) & (!g1663) & (g1664) & (!g1665) & (g1666)) + ((!g820) & (!g773) & (!g1663) & (g1664) & (g1665) & (!g1666)) + ((!g820) & (!g773) & (!g1663) & (g1664) & (g1665) & (g1666)) + ((!g820) & (!g773) & (g1663) & (g1664) & (!g1665) & (!g1666)) + ((!g820) & (!g773) & (g1663) & (g1664) & (!g1665) & (g1666)) + ((!g820) & (!g773) & (g1663) & (g1664) & (g1665) & (!g1666)) + ((!g820) & (!g773) & (g1663) & (g1664) & (g1665) & (g1666)) + ((!g820) & (g773) & (!g1663) & (!g1664) & (!g1665) & (g1666)) + ((!g820) & (g773) & (!g1663) & (!g1664) & (g1665) & (g1666)) + ((!g820) & (g773) & (!g1663) & (g1664) & (!g1665) & (g1666)) + ((!g820) & (g773) & (!g1663) & (g1664) & (g1665) & (g1666)) + ((!g820) & (g773) & (g1663) & (!g1664) & (!g1665) & (g1666)) + ((!g820) & (g773) & (g1663) & (!g1664) & (g1665) & (g1666)) + ((!g820) & (g773) & (g1663) & (g1664) & (!g1665) & (g1666)) + ((!g820) & (g773) & (g1663) & (g1664) & (g1665) & (g1666)) + ((g820) & (!g773) & (g1663) & (!g1664) & (!g1665) & (!g1666)) + ((g820) & (!g773) & (g1663) & (!g1664) & (!g1665) & (g1666)) + ((g820) & (!g773) & (g1663) & (!g1664) & (g1665) & (!g1666)) + ((g820) & (!g773) & (g1663) & (!g1664) & (g1665) & (g1666)) + ((g820) & (!g773) & (g1663) & (g1664) & (!g1665) & (!g1666)) + ((g820) & (!g773) & (g1663) & (g1664) & (!g1665) & (g1666)) + ((g820) & (!g773) & (g1663) & (g1664) & (g1665) & (!g1666)) + ((g820) & (!g773) & (g1663) & (g1664) & (g1665) & (g1666)) + ((g820) & (g773) & (!g1663) & (!g1664) & (g1665) & (!g1666)) + ((g820) & (g773) & (!g1663) & (!g1664) & (g1665) & (g1666)) + ((g820) & (g773) & (!g1663) & (g1664) & (g1665) & (!g1666)) + ((g820) & (g773) & (!g1663) & (g1664) & (g1665) & (g1666)) + ((g820) & (g773) & (g1663) & (!g1664) & (g1665) & (!g1666)) + ((g820) & (g773) & (g1663) & (!g1664) & (g1665) & (g1666)) + ((g820) & (g773) & (g1663) & (g1664) & (g1665) & (!g1666)) + ((g820) & (g773) & (g1663) & (g1664) & (g1665) & (g1666)));
	assign g1668 = (((!g867) & (!g1662) & (!sk[70]) & (g1667)) + ((!g867) & (!g1662) & (sk[70]) & (g1667)) + ((!g867) & (g1662) & (!sk[70]) & (!g1667)) + ((!g867) & (g1662) & (!sk[70]) & (g1667)) + ((!g867) & (g1662) & (sk[70]) & (g1667)) + ((g867) & (!g1662) & (!sk[70]) & (g1667)) + ((g867) & (g1662) & (!sk[70]) & (!g1667)) + ((g867) & (g1662) & (!sk[70]) & (g1667)) + ((g867) & (g1662) & (sk[70]) & (!g1667)) + ((g867) & (g1662) & (sk[70]) & (g1667)));
	assign g1669 = (((!g1592) & (!g1593) & (!g1605) & (g1607) & (!g40) & (g1668)) + ((!g1592) & (!g1593) & (!g1605) & (g1607) & (g40) & (g1668)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (!g40) & (g1668)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (g40) & (g1668)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (!g40) & (g1668)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (g40) & (g1668)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (!g40) & (g1668)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (g40) & (g1668)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (!g40) & (g1668)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (g40) & (g1668)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g40) & (!g1668)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g40) & (g1668)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g40) & (!g1668)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g40) & (g1668)));
	assign g1670 = (((!g410) & (!g411) & (!g412) & (g413) & (g820) & (g773)) + ((!g410) & (!g411) & (g412) & (!g413) & (!g820) & (g773)) + ((!g410) & (!g411) & (g412) & (g413) & (!g820) & (g773)) + ((!g410) & (!g411) & (g412) & (g413) & (g820) & (g773)) + ((!g410) & (g411) & (!g412) & (!g413) & (g820) & (!g773)) + ((!g410) & (g411) & (!g412) & (g413) & (g820) & (!g773)) + ((!g410) & (g411) & (!g412) & (g413) & (g820) & (g773)) + ((!g410) & (g411) & (g412) & (!g413) & (!g820) & (g773)) + ((!g410) & (g411) & (g412) & (!g413) & (g820) & (!g773)) + ((!g410) & (g411) & (g412) & (g413) & (!g820) & (g773)) + ((!g410) & (g411) & (g412) & (g413) & (g820) & (!g773)) + ((!g410) & (g411) & (g412) & (g413) & (g820) & (g773)) + ((g410) & (!g411) & (!g412) & (!g413) & (!g820) & (!g773)) + ((g410) & (!g411) & (!g412) & (g413) & (!g820) & (!g773)) + ((g410) & (!g411) & (!g412) & (g413) & (g820) & (g773)) + ((g410) & (!g411) & (g412) & (!g413) & (!g820) & (!g773)) + ((g410) & (!g411) & (g412) & (!g413) & (!g820) & (g773)) + ((g410) & (!g411) & (g412) & (g413) & (!g820) & (!g773)) + ((g410) & (!g411) & (g412) & (g413) & (!g820) & (g773)) + ((g410) & (!g411) & (g412) & (g413) & (g820) & (g773)) + ((g410) & (g411) & (!g412) & (!g413) & (!g820) & (!g773)) + ((g410) & (g411) & (!g412) & (!g413) & (g820) & (!g773)) + ((g410) & (g411) & (!g412) & (g413) & (!g820) & (!g773)) + ((g410) & (g411) & (!g412) & (g413) & (g820) & (!g773)) + ((g410) & (g411) & (!g412) & (g413) & (g820) & (g773)) + ((g410) & (g411) & (g412) & (!g413) & (!g820) & (!g773)) + ((g410) & (g411) & (g412) & (!g413) & (!g820) & (g773)) + ((g410) & (g411) & (g412) & (!g413) & (g820) & (!g773)) + ((g410) & (g411) & (g412) & (g413) & (!g820) & (!g773)) + ((g410) & (g411) & (g412) & (g413) & (!g820) & (g773)) + ((g410) & (g411) & (g412) & (g413) & (g820) & (!g773)) + ((g410) & (g411) & (g412) & (g413) & (g820) & (g773)));
	assign g1671 = (((!g415) & (!g416) & (!g417) & (g418) & (g820) & (g773)) + ((!g415) & (!g416) & (g417) & (!g418) & (!g820) & (g773)) + ((!g415) & (!g416) & (g417) & (g418) & (!g820) & (g773)) + ((!g415) & (!g416) & (g417) & (g418) & (g820) & (g773)) + ((!g415) & (g416) & (!g417) & (!g418) & (g820) & (!g773)) + ((!g415) & (g416) & (!g417) & (g418) & (g820) & (!g773)) + ((!g415) & (g416) & (!g417) & (g418) & (g820) & (g773)) + ((!g415) & (g416) & (g417) & (!g418) & (!g820) & (g773)) + ((!g415) & (g416) & (g417) & (!g418) & (g820) & (!g773)) + ((!g415) & (g416) & (g417) & (g418) & (!g820) & (g773)) + ((!g415) & (g416) & (g417) & (g418) & (g820) & (!g773)) + ((!g415) & (g416) & (g417) & (g418) & (g820) & (g773)) + ((g415) & (!g416) & (!g417) & (!g418) & (!g820) & (!g773)) + ((g415) & (!g416) & (!g417) & (g418) & (!g820) & (!g773)) + ((g415) & (!g416) & (!g417) & (g418) & (g820) & (g773)) + ((g415) & (!g416) & (g417) & (!g418) & (!g820) & (!g773)) + ((g415) & (!g416) & (g417) & (!g418) & (!g820) & (g773)) + ((g415) & (!g416) & (g417) & (g418) & (!g820) & (!g773)) + ((g415) & (!g416) & (g417) & (g418) & (!g820) & (g773)) + ((g415) & (!g416) & (g417) & (g418) & (g820) & (g773)) + ((g415) & (g416) & (!g417) & (!g418) & (!g820) & (!g773)) + ((g415) & (g416) & (!g417) & (!g418) & (g820) & (!g773)) + ((g415) & (g416) & (!g417) & (g418) & (!g820) & (!g773)) + ((g415) & (g416) & (!g417) & (g418) & (g820) & (!g773)) + ((g415) & (g416) & (!g417) & (g418) & (g820) & (g773)) + ((g415) & (g416) & (g417) & (!g418) & (!g820) & (!g773)) + ((g415) & (g416) & (g417) & (!g418) & (!g820) & (g773)) + ((g415) & (g416) & (g417) & (!g418) & (g820) & (!g773)) + ((g415) & (g416) & (g417) & (g418) & (!g820) & (!g773)) + ((g415) & (g416) & (g417) & (g418) & (!g820) & (g773)) + ((g415) & (g416) & (g417) & (g418) & (g820) & (!g773)) + ((g415) & (g416) & (g417) & (g418) & (g820) & (g773)));
	assign g1672 = (((!g420) & (!g421) & (!g422) & (g423) & (g820) & (g773)) + ((!g420) & (!g421) & (g422) & (!g423) & (!g820) & (g773)) + ((!g420) & (!g421) & (g422) & (g423) & (!g820) & (g773)) + ((!g420) & (!g421) & (g422) & (g423) & (g820) & (g773)) + ((!g420) & (g421) & (!g422) & (!g423) & (g820) & (!g773)) + ((!g420) & (g421) & (!g422) & (g423) & (g820) & (!g773)) + ((!g420) & (g421) & (!g422) & (g423) & (g820) & (g773)) + ((!g420) & (g421) & (g422) & (!g423) & (!g820) & (g773)) + ((!g420) & (g421) & (g422) & (!g423) & (g820) & (!g773)) + ((!g420) & (g421) & (g422) & (g423) & (!g820) & (g773)) + ((!g420) & (g421) & (g422) & (g423) & (g820) & (!g773)) + ((!g420) & (g421) & (g422) & (g423) & (g820) & (g773)) + ((g420) & (!g421) & (!g422) & (!g423) & (!g820) & (!g773)) + ((g420) & (!g421) & (!g422) & (g423) & (!g820) & (!g773)) + ((g420) & (!g421) & (!g422) & (g423) & (g820) & (g773)) + ((g420) & (!g421) & (g422) & (!g423) & (!g820) & (!g773)) + ((g420) & (!g421) & (g422) & (!g423) & (!g820) & (g773)) + ((g420) & (!g421) & (g422) & (g423) & (!g820) & (!g773)) + ((g420) & (!g421) & (g422) & (g423) & (!g820) & (g773)) + ((g420) & (!g421) & (g422) & (g423) & (g820) & (g773)) + ((g420) & (g421) & (!g422) & (!g423) & (!g820) & (!g773)) + ((g420) & (g421) & (!g422) & (!g423) & (g820) & (!g773)) + ((g420) & (g421) & (!g422) & (g423) & (!g820) & (!g773)) + ((g420) & (g421) & (!g422) & (g423) & (g820) & (!g773)) + ((g420) & (g421) & (!g422) & (g423) & (g820) & (g773)) + ((g420) & (g421) & (g422) & (!g423) & (!g820) & (!g773)) + ((g420) & (g421) & (g422) & (!g423) & (!g820) & (g773)) + ((g420) & (g421) & (g422) & (!g423) & (g820) & (!g773)) + ((g420) & (g421) & (g422) & (g423) & (!g820) & (!g773)) + ((g420) & (g421) & (g422) & (g423) & (!g820) & (g773)) + ((g420) & (g421) & (g422) & (g423) & (g820) & (!g773)) + ((g420) & (g421) & (g422) & (g423) & (g820) & (g773)));
	assign g1673 = (((!g425) & (!g426) & (!g427) & (g428) & (g820) & (g773)) + ((!g425) & (!g426) & (g427) & (!g428) & (!g820) & (g773)) + ((!g425) & (!g426) & (g427) & (g428) & (!g820) & (g773)) + ((!g425) & (!g426) & (g427) & (g428) & (g820) & (g773)) + ((!g425) & (g426) & (!g427) & (!g428) & (g820) & (!g773)) + ((!g425) & (g426) & (!g427) & (g428) & (g820) & (!g773)) + ((!g425) & (g426) & (!g427) & (g428) & (g820) & (g773)) + ((!g425) & (g426) & (g427) & (!g428) & (!g820) & (g773)) + ((!g425) & (g426) & (g427) & (!g428) & (g820) & (!g773)) + ((!g425) & (g426) & (g427) & (g428) & (!g820) & (g773)) + ((!g425) & (g426) & (g427) & (g428) & (g820) & (!g773)) + ((!g425) & (g426) & (g427) & (g428) & (g820) & (g773)) + ((g425) & (!g426) & (!g427) & (!g428) & (!g820) & (!g773)) + ((g425) & (!g426) & (!g427) & (g428) & (!g820) & (!g773)) + ((g425) & (!g426) & (!g427) & (g428) & (g820) & (g773)) + ((g425) & (!g426) & (g427) & (!g428) & (!g820) & (!g773)) + ((g425) & (!g426) & (g427) & (!g428) & (!g820) & (g773)) + ((g425) & (!g426) & (g427) & (g428) & (!g820) & (!g773)) + ((g425) & (!g426) & (g427) & (g428) & (!g820) & (g773)) + ((g425) & (!g426) & (g427) & (g428) & (g820) & (g773)) + ((g425) & (g426) & (!g427) & (!g428) & (!g820) & (!g773)) + ((g425) & (g426) & (!g427) & (!g428) & (g820) & (!g773)) + ((g425) & (g426) & (!g427) & (g428) & (!g820) & (!g773)) + ((g425) & (g426) & (!g427) & (g428) & (g820) & (!g773)) + ((g425) & (g426) & (!g427) & (g428) & (g820) & (g773)) + ((g425) & (g426) & (g427) & (!g428) & (!g820) & (!g773)) + ((g425) & (g426) & (g427) & (!g428) & (!g820) & (g773)) + ((g425) & (g426) & (g427) & (!g428) & (g820) & (!g773)) + ((g425) & (g426) & (g427) & (g428) & (!g820) & (!g773)) + ((g425) & (g426) & (g427) & (g428) & (!g820) & (g773)) + ((g425) & (g426) & (g427) & (g428) & (g820) & (!g773)) + ((g425) & (g426) & (g427) & (g428) & (g820) & (g773)));
	assign g1674 = (((!g1670) & (!g1671) & (!g1672) & (g1673) & (g677) & (g726)) + ((!g1670) & (!g1671) & (g1672) & (!g1673) & (!g677) & (g726)) + ((!g1670) & (!g1671) & (g1672) & (g1673) & (!g677) & (g726)) + ((!g1670) & (!g1671) & (g1672) & (g1673) & (g677) & (g726)) + ((!g1670) & (g1671) & (!g1672) & (!g1673) & (g677) & (!g726)) + ((!g1670) & (g1671) & (!g1672) & (g1673) & (g677) & (!g726)) + ((!g1670) & (g1671) & (!g1672) & (g1673) & (g677) & (g726)) + ((!g1670) & (g1671) & (g1672) & (!g1673) & (!g677) & (g726)) + ((!g1670) & (g1671) & (g1672) & (!g1673) & (g677) & (!g726)) + ((!g1670) & (g1671) & (g1672) & (g1673) & (!g677) & (g726)) + ((!g1670) & (g1671) & (g1672) & (g1673) & (g677) & (!g726)) + ((!g1670) & (g1671) & (g1672) & (g1673) & (g677) & (g726)) + ((g1670) & (!g1671) & (!g1672) & (!g1673) & (!g677) & (!g726)) + ((g1670) & (!g1671) & (!g1672) & (g1673) & (!g677) & (!g726)) + ((g1670) & (!g1671) & (!g1672) & (g1673) & (g677) & (g726)) + ((g1670) & (!g1671) & (g1672) & (!g1673) & (!g677) & (!g726)) + ((g1670) & (!g1671) & (g1672) & (!g1673) & (!g677) & (g726)) + ((g1670) & (!g1671) & (g1672) & (g1673) & (!g677) & (!g726)) + ((g1670) & (!g1671) & (g1672) & (g1673) & (!g677) & (g726)) + ((g1670) & (!g1671) & (g1672) & (g1673) & (g677) & (g726)) + ((g1670) & (g1671) & (!g1672) & (!g1673) & (!g677) & (!g726)) + ((g1670) & (g1671) & (!g1672) & (!g1673) & (g677) & (!g726)) + ((g1670) & (g1671) & (!g1672) & (g1673) & (!g677) & (!g726)) + ((g1670) & (g1671) & (!g1672) & (g1673) & (g677) & (!g726)) + ((g1670) & (g1671) & (!g1672) & (g1673) & (g677) & (g726)) + ((g1670) & (g1671) & (g1672) & (!g1673) & (!g677) & (!g726)) + ((g1670) & (g1671) & (g1672) & (!g1673) & (!g677) & (g726)) + ((g1670) & (g1671) & (g1672) & (!g1673) & (g677) & (!g726)) + ((g1670) & (g1671) & (g1672) & (g1673) & (!g677) & (!g726)) + ((g1670) & (g1671) & (g1672) & (g1673) & (!g677) & (g726)) + ((g1670) & (g1671) & (g1672) & (g1673) & (g677) & (!g726)) + ((g1670) & (g1671) & (g1672) & (g1673) & (g677) & (g726)));
	assign g1675 = (((!g431) & (!g432) & (!g433) & (g434) & (g677) & (g726)) + ((!g431) & (!g432) & (g433) & (!g434) & (!g677) & (g726)) + ((!g431) & (!g432) & (g433) & (g434) & (!g677) & (g726)) + ((!g431) & (!g432) & (g433) & (g434) & (g677) & (g726)) + ((!g431) & (g432) & (!g433) & (!g434) & (g677) & (!g726)) + ((!g431) & (g432) & (!g433) & (g434) & (g677) & (!g726)) + ((!g431) & (g432) & (!g433) & (g434) & (g677) & (g726)) + ((!g431) & (g432) & (g433) & (!g434) & (!g677) & (g726)) + ((!g431) & (g432) & (g433) & (!g434) & (g677) & (!g726)) + ((!g431) & (g432) & (g433) & (g434) & (!g677) & (g726)) + ((!g431) & (g432) & (g433) & (g434) & (g677) & (!g726)) + ((!g431) & (g432) & (g433) & (g434) & (g677) & (g726)) + ((g431) & (!g432) & (!g433) & (!g434) & (!g677) & (!g726)) + ((g431) & (!g432) & (!g433) & (g434) & (!g677) & (!g726)) + ((g431) & (!g432) & (!g433) & (g434) & (g677) & (g726)) + ((g431) & (!g432) & (g433) & (!g434) & (!g677) & (!g726)) + ((g431) & (!g432) & (g433) & (!g434) & (!g677) & (g726)) + ((g431) & (!g432) & (g433) & (g434) & (!g677) & (!g726)) + ((g431) & (!g432) & (g433) & (g434) & (!g677) & (g726)) + ((g431) & (!g432) & (g433) & (g434) & (g677) & (g726)) + ((g431) & (g432) & (!g433) & (!g434) & (!g677) & (!g726)) + ((g431) & (g432) & (!g433) & (!g434) & (g677) & (!g726)) + ((g431) & (g432) & (!g433) & (g434) & (!g677) & (!g726)) + ((g431) & (g432) & (!g433) & (g434) & (g677) & (!g726)) + ((g431) & (g432) & (!g433) & (g434) & (g677) & (g726)) + ((g431) & (g432) & (g433) & (!g434) & (!g677) & (!g726)) + ((g431) & (g432) & (g433) & (!g434) & (!g677) & (g726)) + ((g431) & (g432) & (g433) & (!g434) & (g677) & (!g726)) + ((g431) & (g432) & (g433) & (g434) & (!g677) & (!g726)) + ((g431) & (g432) & (g433) & (g434) & (!g677) & (g726)) + ((g431) & (g432) & (g433) & (g434) & (g677) & (!g726)) + ((g431) & (g432) & (g433) & (g434) & (g677) & (g726)));
	assign g1676 = (((!g677) & (!g726) & (!g436) & (g437) & (!sk[78]) & (!g438)) + ((!g677) & (!g726) & (!g436) & (g437) & (!sk[78]) & (g438)) + ((!g677) & (!g726) & (g436) & (!g437) & (!sk[78]) & (!g438)) + ((!g677) & (!g726) & (g436) & (!g437) & (!sk[78]) & (g438)) + ((!g677) & (!g726) & (g436) & (g437) & (!sk[78]) & (!g438)) + ((!g677) & (!g726) & (g436) & (g437) & (!sk[78]) & (g438)) + ((!g677) & (g726) & (!g436) & (!g437) & (!sk[78]) & (!g438)) + ((!g677) & (g726) & (!g436) & (!g437) & (!sk[78]) & (g438)) + ((!g677) & (g726) & (!g436) & (!g437) & (sk[78]) & (g438)) + ((!g677) & (g726) & (!g436) & (g437) & (!sk[78]) & (!g438)) + ((!g677) & (g726) & (!g436) & (g437) & (!sk[78]) & (g438)) + ((!g677) & (g726) & (!g436) & (g437) & (sk[78]) & (g438)) + ((!g677) & (g726) & (g436) & (!g437) & (!sk[78]) & (!g438)) + ((!g677) & (g726) & (g436) & (!g437) & (!sk[78]) & (g438)) + ((!g677) & (g726) & (g436) & (!g437) & (sk[78]) & (g438)) + ((!g677) & (g726) & (g436) & (g437) & (!sk[78]) & (!g438)) + ((!g677) & (g726) & (g436) & (g437) & (!sk[78]) & (g438)) + ((!g677) & (g726) & (g436) & (g437) & (sk[78]) & (g438)) + ((g677) & (!g726) & (!g436) & (g437) & (!sk[78]) & (!g438)) + ((g677) & (!g726) & (!g436) & (g437) & (!sk[78]) & (g438)) + ((g677) & (!g726) & (g436) & (!g437) & (!sk[78]) & (!g438)) + ((g677) & (!g726) & (g436) & (!g437) & (!sk[78]) & (g438)) + ((g677) & (!g726) & (g436) & (!g437) & (sk[78]) & (!g438)) + ((g677) & (!g726) & (g436) & (!g437) & (sk[78]) & (g438)) + ((g677) & (!g726) & (g436) & (g437) & (!sk[78]) & (!g438)) + ((g677) & (!g726) & (g436) & (g437) & (!sk[78]) & (g438)) + ((g677) & (!g726) & (g436) & (g437) & (sk[78]) & (!g438)) + ((g677) & (!g726) & (g436) & (g437) & (sk[78]) & (g438)) + ((g677) & (g726) & (!g436) & (!g437) & (!sk[78]) & (!g438)) + ((g677) & (g726) & (!g436) & (!g437) & (!sk[78]) & (g438)) + ((g677) & (g726) & (!g436) & (g437) & (!sk[78]) & (!g438)) + ((g677) & (g726) & (!g436) & (g437) & (!sk[78]) & (g438)) + ((g677) & (g726) & (!g436) & (g437) & (sk[78]) & (!g438)) + ((g677) & (g726) & (!g436) & (g437) & (sk[78]) & (g438)) + ((g677) & (g726) & (g436) & (!g437) & (!sk[78]) & (!g438)) + ((g677) & (g726) & (g436) & (!g437) & (!sk[78]) & (g438)) + ((g677) & (g726) & (g436) & (g437) & (!sk[78]) & (!g438)) + ((g677) & (g726) & (g436) & (g437) & (!sk[78]) & (g438)) + ((g677) & (g726) & (g436) & (g437) & (sk[78]) & (!g438)) + ((g677) & (g726) & (g436) & (g437) & (sk[78]) & (g438)));
	assign g1677 = (((!g440) & (!g441) & (!g442) & (g443) & (g677) & (g726)) + ((!g440) & (!g441) & (g442) & (!g443) & (!g677) & (g726)) + ((!g440) & (!g441) & (g442) & (g443) & (!g677) & (g726)) + ((!g440) & (!g441) & (g442) & (g443) & (g677) & (g726)) + ((!g440) & (g441) & (!g442) & (!g443) & (g677) & (!g726)) + ((!g440) & (g441) & (!g442) & (g443) & (g677) & (!g726)) + ((!g440) & (g441) & (!g442) & (g443) & (g677) & (g726)) + ((!g440) & (g441) & (g442) & (!g443) & (!g677) & (g726)) + ((!g440) & (g441) & (g442) & (!g443) & (g677) & (!g726)) + ((!g440) & (g441) & (g442) & (g443) & (!g677) & (g726)) + ((!g440) & (g441) & (g442) & (g443) & (g677) & (!g726)) + ((!g440) & (g441) & (g442) & (g443) & (g677) & (g726)) + ((g440) & (!g441) & (!g442) & (!g443) & (!g677) & (!g726)) + ((g440) & (!g441) & (!g442) & (g443) & (!g677) & (!g726)) + ((g440) & (!g441) & (!g442) & (g443) & (g677) & (g726)) + ((g440) & (!g441) & (g442) & (!g443) & (!g677) & (!g726)) + ((g440) & (!g441) & (g442) & (!g443) & (!g677) & (g726)) + ((g440) & (!g441) & (g442) & (g443) & (!g677) & (!g726)) + ((g440) & (!g441) & (g442) & (g443) & (!g677) & (g726)) + ((g440) & (!g441) & (g442) & (g443) & (g677) & (g726)) + ((g440) & (g441) & (!g442) & (!g443) & (!g677) & (!g726)) + ((g440) & (g441) & (!g442) & (!g443) & (g677) & (!g726)) + ((g440) & (g441) & (!g442) & (g443) & (!g677) & (!g726)) + ((g440) & (g441) & (!g442) & (g443) & (g677) & (!g726)) + ((g440) & (g441) & (!g442) & (g443) & (g677) & (g726)) + ((g440) & (g441) & (g442) & (!g443) & (!g677) & (!g726)) + ((g440) & (g441) & (g442) & (!g443) & (!g677) & (g726)) + ((g440) & (g441) & (g442) & (!g443) & (g677) & (!g726)) + ((g440) & (g441) & (g442) & (g443) & (!g677) & (!g726)) + ((g440) & (g441) & (g442) & (g443) & (!g677) & (g726)) + ((g440) & (g441) & (g442) & (g443) & (g677) & (!g726)) + ((g440) & (g441) & (g442) & (g443) & (g677) & (g726)));
	assign g1678 = (((!g445) & (!g446) & (!g447) & (g448) & (g677) & (g726)) + ((!g445) & (!g446) & (g447) & (!g448) & (!g677) & (g726)) + ((!g445) & (!g446) & (g447) & (g448) & (!g677) & (g726)) + ((!g445) & (!g446) & (g447) & (g448) & (g677) & (g726)) + ((!g445) & (g446) & (!g447) & (!g448) & (g677) & (!g726)) + ((!g445) & (g446) & (!g447) & (g448) & (g677) & (!g726)) + ((!g445) & (g446) & (!g447) & (g448) & (g677) & (g726)) + ((!g445) & (g446) & (g447) & (!g448) & (!g677) & (g726)) + ((!g445) & (g446) & (g447) & (!g448) & (g677) & (!g726)) + ((!g445) & (g446) & (g447) & (g448) & (!g677) & (g726)) + ((!g445) & (g446) & (g447) & (g448) & (g677) & (!g726)) + ((!g445) & (g446) & (g447) & (g448) & (g677) & (g726)) + ((g445) & (!g446) & (!g447) & (!g448) & (!g677) & (!g726)) + ((g445) & (!g446) & (!g447) & (g448) & (!g677) & (!g726)) + ((g445) & (!g446) & (!g447) & (g448) & (g677) & (g726)) + ((g445) & (!g446) & (g447) & (!g448) & (!g677) & (!g726)) + ((g445) & (!g446) & (g447) & (!g448) & (!g677) & (g726)) + ((g445) & (!g446) & (g447) & (g448) & (!g677) & (!g726)) + ((g445) & (!g446) & (g447) & (g448) & (!g677) & (g726)) + ((g445) & (!g446) & (g447) & (g448) & (g677) & (g726)) + ((g445) & (g446) & (!g447) & (!g448) & (!g677) & (!g726)) + ((g445) & (g446) & (!g447) & (!g448) & (g677) & (!g726)) + ((g445) & (g446) & (!g447) & (g448) & (!g677) & (!g726)) + ((g445) & (g446) & (!g447) & (g448) & (g677) & (!g726)) + ((g445) & (g446) & (!g447) & (g448) & (g677) & (g726)) + ((g445) & (g446) & (g447) & (!g448) & (!g677) & (!g726)) + ((g445) & (g446) & (g447) & (!g448) & (!g677) & (g726)) + ((g445) & (g446) & (g447) & (!g448) & (g677) & (!g726)) + ((g445) & (g446) & (g447) & (g448) & (!g677) & (!g726)) + ((g445) & (g446) & (g447) & (g448) & (!g677) & (g726)) + ((g445) & (g446) & (g447) & (g448) & (g677) & (!g726)) + ((g445) & (g446) & (g447) & (g448) & (g677) & (g726)));
	assign g1679 = (((!g820) & (!g773) & (!g1675) & (g1676) & (!g1677) & (!g1678)) + ((!g820) & (!g773) & (!g1675) & (g1676) & (!g1677) & (g1678)) + ((!g820) & (!g773) & (!g1675) & (g1676) & (g1677) & (!g1678)) + ((!g820) & (!g773) & (!g1675) & (g1676) & (g1677) & (g1678)) + ((!g820) & (!g773) & (g1675) & (g1676) & (!g1677) & (!g1678)) + ((!g820) & (!g773) & (g1675) & (g1676) & (!g1677) & (g1678)) + ((!g820) & (!g773) & (g1675) & (g1676) & (g1677) & (!g1678)) + ((!g820) & (!g773) & (g1675) & (g1676) & (g1677) & (g1678)) + ((!g820) & (g773) & (!g1675) & (!g1676) & (!g1677) & (g1678)) + ((!g820) & (g773) & (!g1675) & (!g1676) & (g1677) & (g1678)) + ((!g820) & (g773) & (!g1675) & (g1676) & (!g1677) & (g1678)) + ((!g820) & (g773) & (!g1675) & (g1676) & (g1677) & (g1678)) + ((!g820) & (g773) & (g1675) & (!g1676) & (!g1677) & (g1678)) + ((!g820) & (g773) & (g1675) & (!g1676) & (g1677) & (g1678)) + ((!g820) & (g773) & (g1675) & (g1676) & (!g1677) & (g1678)) + ((!g820) & (g773) & (g1675) & (g1676) & (g1677) & (g1678)) + ((g820) & (!g773) & (g1675) & (!g1676) & (!g1677) & (!g1678)) + ((g820) & (!g773) & (g1675) & (!g1676) & (!g1677) & (g1678)) + ((g820) & (!g773) & (g1675) & (!g1676) & (g1677) & (!g1678)) + ((g820) & (!g773) & (g1675) & (!g1676) & (g1677) & (g1678)) + ((g820) & (!g773) & (g1675) & (g1676) & (!g1677) & (!g1678)) + ((g820) & (!g773) & (g1675) & (g1676) & (!g1677) & (g1678)) + ((g820) & (!g773) & (g1675) & (g1676) & (g1677) & (!g1678)) + ((g820) & (!g773) & (g1675) & (g1676) & (g1677) & (g1678)) + ((g820) & (g773) & (!g1675) & (!g1676) & (g1677) & (!g1678)) + ((g820) & (g773) & (!g1675) & (!g1676) & (g1677) & (g1678)) + ((g820) & (g773) & (!g1675) & (g1676) & (g1677) & (!g1678)) + ((g820) & (g773) & (!g1675) & (g1676) & (g1677) & (g1678)) + ((g820) & (g773) & (g1675) & (!g1676) & (g1677) & (!g1678)) + ((g820) & (g773) & (g1675) & (!g1676) & (g1677) & (g1678)) + ((g820) & (g773) & (g1675) & (g1676) & (g1677) & (!g1678)) + ((g820) & (g773) & (g1675) & (g1676) & (g1677) & (g1678)));
	assign g1680 = (((!g867) & (!g1674) & (!sk[82]) & (g1679)) + ((!g867) & (!g1674) & (sk[82]) & (g1679)) + ((!g867) & (g1674) & (!sk[82]) & (!g1679)) + ((!g867) & (g1674) & (!sk[82]) & (g1679)) + ((!g867) & (g1674) & (sk[82]) & (g1679)) + ((g867) & (!g1674) & (!sk[82]) & (g1679)) + ((g867) & (g1674) & (!sk[82]) & (!g1679)) + ((g867) & (g1674) & (!sk[82]) & (g1679)) + ((g867) & (g1674) & (sk[82]) & (!g1679)) + ((g867) & (g1674) & (sk[82]) & (g1679)));
	assign g1681 = (((!g1592) & (!g1593) & (!g1605) & (g1607) & (!g41) & (g1680)) + ((!g1592) & (!g1593) & (!g1605) & (g1607) & (g41) & (g1680)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (!g41) & (g1680)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (g41) & (g1680)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (!g41) & (g1680)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (g41) & (g1680)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (!g41) & (g1680)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (g41) & (g1680)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (!g41) & (g1680)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (g41) & (g1680)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g41) & (!g1680)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g41) & (g1680)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g41) & (!g1680)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g41) & (g1680)));
	assign g1682 = (((!g454) & (!g459) & (!g464) & (g469) & (g820) & (g773)) + ((!g454) & (!g459) & (g464) & (!g469) & (!g820) & (g773)) + ((!g454) & (!g459) & (g464) & (g469) & (!g820) & (g773)) + ((!g454) & (!g459) & (g464) & (g469) & (g820) & (g773)) + ((!g454) & (g459) & (!g464) & (!g469) & (g820) & (!g773)) + ((!g454) & (g459) & (!g464) & (g469) & (g820) & (!g773)) + ((!g454) & (g459) & (!g464) & (g469) & (g820) & (g773)) + ((!g454) & (g459) & (g464) & (!g469) & (!g820) & (g773)) + ((!g454) & (g459) & (g464) & (!g469) & (g820) & (!g773)) + ((!g454) & (g459) & (g464) & (g469) & (!g820) & (g773)) + ((!g454) & (g459) & (g464) & (g469) & (g820) & (!g773)) + ((!g454) & (g459) & (g464) & (g469) & (g820) & (g773)) + ((g454) & (!g459) & (!g464) & (!g469) & (!g820) & (!g773)) + ((g454) & (!g459) & (!g464) & (g469) & (!g820) & (!g773)) + ((g454) & (!g459) & (!g464) & (g469) & (g820) & (g773)) + ((g454) & (!g459) & (g464) & (!g469) & (!g820) & (!g773)) + ((g454) & (!g459) & (g464) & (!g469) & (!g820) & (g773)) + ((g454) & (!g459) & (g464) & (g469) & (!g820) & (!g773)) + ((g454) & (!g459) & (g464) & (g469) & (!g820) & (g773)) + ((g454) & (!g459) & (g464) & (g469) & (g820) & (g773)) + ((g454) & (g459) & (!g464) & (!g469) & (!g820) & (!g773)) + ((g454) & (g459) & (!g464) & (!g469) & (g820) & (!g773)) + ((g454) & (g459) & (!g464) & (g469) & (!g820) & (!g773)) + ((g454) & (g459) & (!g464) & (g469) & (g820) & (!g773)) + ((g454) & (g459) & (!g464) & (g469) & (g820) & (g773)) + ((g454) & (g459) & (g464) & (!g469) & (!g820) & (!g773)) + ((g454) & (g459) & (g464) & (!g469) & (!g820) & (g773)) + ((g454) & (g459) & (g464) & (!g469) & (g820) & (!g773)) + ((g454) & (g459) & (g464) & (g469) & (!g820) & (!g773)) + ((g454) & (g459) & (g464) & (g469) & (!g820) & (g773)) + ((g454) & (g459) & (g464) & (g469) & (g820) & (!g773)) + ((g454) & (g459) & (g464) & (g469) & (g820) & (g773)));
	assign g1683 = (((!g455) & (!g460) & (!g465) & (g470) & (g820) & (g773)) + ((!g455) & (!g460) & (g465) & (!g470) & (!g820) & (g773)) + ((!g455) & (!g460) & (g465) & (g470) & (!g820) & (g773)) + ((!g455) & (!g460) & (g465) & (g470) & (g820) & (g773)) + ((!g455) & (g460) & (!g465) & (!g470) & (g820) & (!g773)) + ((!g455) & (g460) & (!g465) & (g470) & (g820) & (!g773)) + ((!g455) & (g460) & (!g465) & (g470) & (g820) & (g773)) + ((!g455) & (g460) & (g465) & (!g470) & (!g820) & (g773)) + ((!g455) & (g460) & (g465) & (!g470) & (g820) & (!g773)) + ((!g455) & (g460) & (g465) & (g470) & (!g820) & (g773)) + ((!g455) & (g460) & (g465) & (g470) & (g820) & (!g773)) + ((!g455) & (g460) & (g465) & (g470) & (g820) & (g773)) + ((g455) & (!g460) & (!g465) & (!g470) & (!g820) & (!g773)) + ((g455) & (!g460) & (!g465) & (g470) & (!g820) & (!g773)) + ((g455) & (!g460) & (!g465) & (g470) & (g820) & (g773)) + ((g455) & (!g460) & (g465) & (!g470) & (!g820) & (!g773)) + ((g455) & (!g460) & (g465) & (!g470) & (!g820) & (g773)) + ((g455) & (!g460) & (g465) & (g470) & (!g820) & (!g773)) + ((g455) & (!g460) & (g465) & (g470) & (!g820) & (g773)) + ((g455) & (!g460) & (g465) & (g470) & (g820) & (g773)) + ((g455) & (g460) & (!g465) & (!g470) & (!g820) & (!g773)) + ((g455) & (g460) & (!g465) & (!g470) & (g820) & (!g773)) + ((g455) & (g460) & (!g465) & (g470) & (!g820) & (!g773)) + ((g455) & (g460) & (!g465) & (g470) & (g820) & (!g773)) + ((g455) & (g460) & (!g465) & (g470) & (g820) & (g773)) + ((g455) & (g460) & (g465) & (!g470) & (!g820) & (!g773)) + ((g455) & (g460) & (g465) & (!g470) & (!g820) & (g773)) + ((g455) & (g460) & (g465) & (!g470) & (g820) & (!g773)) + ((g455) & (g460) & (g465) & (g470) & (!g820) & (!g773)) + ((g455) & (g460) & (g465) & (g470) & (!g820) & (g773)) + ((g455) & (g460) & (g465) & (g470) & (g820) & (!g773)) + ((g455) & (g460) & (g465) & (g470) & (g820) & (g773)));
	assign g1684 = (((!g456) & (!g461) & (!g466) & (g471) & (g820) & (g773)) + ((!g456) & (!g461) & (g466) & (!g471) & (!g820) & (g773)) + ((!g456) & (!g461) & (g466) & (g471) & (!g820) & (g773)) + ((!g456) & (!g461) & (g466) & (g471) & (g820) & (g773)) + ((!g456) & (g461) & (!g466) & (!g471) & (g820) & (!g773)) + ((!g456) & (g461) & (!g466) & (g471) & (g820) & (!g773)) + ((!g456) & (g461) & (!g466) & (g471) & (g820) & (g773)) + ((!g456) & (g461) & (g466) & (!g471) & (!g820) & (g773)) + ((!g456) & (g461) & (g466) & (!g471) & (g820) & (!g773)) + ((!g456) & (g461) & (g466) & (g471) & (!g820) & (g773)) + ((!g456) & (g461) & (g466) & (g471) & (g820) & (!g773)) + ((!g456) & (g461) & (g466) & (g471) & (g820) & (g773)) + ((g456) & (!g461) & (!g466) & (!g471) & (!g820) & (!g773)) + ((g456) & (!g461) & (!g466) & (g471) & (!g820) & (!g773)) + ((g456) & (!g461) & (!g466) & (g471) & (g820) & (g773)) + ((g456) & (!g461) & (g466) & (!g471) & (!g820) & (!g773)) + ((g456) & (!g461) & (g466) & (!g471) & (!g820) & (g773)) + ((g456) & (!g461) & (g466) & (g471) & (!g820) & (!g773)) + ((g456) & (!g461) & (g466) & (g471) & (!g820) & (g773)) + ((g456) & (!g461) & (g466) & (g471) & (g820) & (g773)) + ((g456) & (g461) & (!g466) & (!g471) & (!g820) & (!g773)) + ((g456) & (g461) & (!g466) & (!g471) & (g820) & (!g773)) + ((g456) & (g461) & (!g466) & (g471) & (!g820) & (!g773)) + ((g456) & (g461) & (!g466) & (g471) & (g820) & (!g773)) + ((g456) & (g461) & (!g466) & (g471) & (g820) & (g773)) + ((g456) & (g461) & (g466) & (!g471) & (!g820) & (!g773)) + ((g456) & (g461) & (g466) & (!g471) & (!g820) & (g773)) + ((g456) & (g461) & (g466) & (!g471) & (g820) & (!g773)) + ((g456) & (g461) & (g466) & (g471) & (!g820) & (!g773)) + ((g456) & (g461) & (g466) & (g471) & (!g820) & (g773)) + ((g456) & (g461) & (g466) & (g471) & (g820) & (!g773)) + ((g456) & (g461) & (g466) & (g471) & (g820) & (g773)));
	assign g1685 = (((!g457) & (!g462) & (!g467) & (g472) & (g820) & (g773)) + ((!g457) & (!g462) & (g467) & (!g472) & (!g820) & (g773)) + ((!g457) & (!g462) & (g467) & (g472) & (!g820) & (g773)) + ((!g457) & (!g462) & (g467) & (g472) & (g820) & (g773)) + ((!g457) & (g462) & (!g467) & (!g472) & (g820) & (!g773)) + ((!g457) & (g462) & (!g467) & (g472) & (g820) & (!g773)) + ((!g457) & (g462) & (!g467) & (g472) & (g820) & (g773)) + ((!g457) & (g462) & (g467) & (!g472) & (!g820) & (g773)) + ((!g457) & (g462) & (g467) & (!g472) & (g820) & (!g773)) + ((!g457) & (g462) & (g467) & (g472) & (!g820) & (g773)) + ((!g457) & (g462) & (g467) & (g472) & (g820) & (!g773)) + ((!g457) & (g462) & (g467) & (g472) & (g820) & (g773)) + ((g457) & (!g462) & (!g467) & (!g472) & (!g820) & (!g773)) + ((g457) & (!g462) & (!g467) & (g472) & (!g820) & (!g773)) + ((g457) & (!g462) & (!g467) & (g472) & (g820) & (g773)) + ((g457) & (!g462) & (g467) & (!g472) & (!g820) & (!g773)) + ((g457) & (!g462) & (g467) & (!g472) & (!g820) & (g773)) + ((g457) & (!g462) & (g467) & (g472) & (!g820) & (!g773)) + ((g457) & (!g462) & (g467) & (g472) & (!g820) & (g773)) + ((g457) & (!g462) & (g467) & (g472) & (g820) & (g773)) + ((g457) & (g462) & (!g467) & (!g472) & (!g820) & (!g773)) + ((g457) & (g462) & (!g467) & (!g472) & (g820) & (!g773)) + ((g457) & (g462) & (!g467) & (g472) & (!g820) & (!g773)) + ((g457) & (g462) & (!g467) & (g472) & (g820) & (!g773)) + ((g457) & (g462) & (!g467) & (g472) & (g820) & (g773)) + ((g457) & (g462) & (g467) & (!g472) & (!g820) & (!g773)) + ((g457) & (g462) & (g467) & (!g472) & (!g820) & (g773)) + ((g457) & (g462) & (g467) & (!g472) & (g820) & (!g773)) + ((g457) & (g462) & (g467) & (g472) & (!g820) & (!g773)) + ((g457) & (g462) & (g467) & (g472) & (!g820) & (g773)) + ((g457) & (g462) & (g467) & (g472) & (g820) & (!g773)) + ((g457) & (g462) & (g467) & (g472) & (g820) & (g773)));
	assign g1686 = (((!g1682) & (!g1683) & (!g1684) & (g1685) & (g677) & (g726)) + ((!g1682) & (!g1683) & (g1684) & (!g1685) & (!g677) & (g726)) + ((!g1682) & (!g1683) & (g1684) & (g1685) & (!g677) & (g726)) + ((!g1682) & (!g1683) & (g1684) & (g1685) & (g677) & (g726)) + ((!g1682) & (g1683) & (!g1684) & (!g1685) & (g677) & (!g726)) + ((!g1682) & (g1683) & (!g1684) & (g1685) & (g677) & (!g726)) + ((!g1682) & (g1683) & (!g1684) & (g1685) & (g677) & (g726)) + ((!g1682) & (g1683) & (g1684) & (!g1685) & (!g677) & (g726)) + ((!g1682) & (g1683) & (g1684) & (!g1685) & (g677) & (!g726)) + ((!g1682) & (g1683) & (g1684) & (g1685) & (!g677) & (g726)) + ((!g1682) & (g1683) & (g1684) & (g1685) & (g677) & (!g726)) + ((!g1682) & (g1683) & (g1684) & (g1685) & (g677) & (g726)) + ((g1682) & (!g1683) & (!g1684) & (!g1685) & (!g677) & (!g726)) + ((g1682) & (!g1683) & (!g1684) & (g1685) & (!g677) & (!g726)) + ((g1682) & (!g1683) & (!g1684) & (g1685) & (g677) & (g726)) + ((g1682) & (!g1683) & (g1684) & (!g1685) & (!g677) & (!g726)) + ((g1682) & (!g1683) & (g1684) & (!g1685) & (!g677) & (g726)) + ((g1682) & (!g1683) & (g1684) & (g1685) & (!g677) & (!g726)) + ((g1682) & (!g1683) & (g1684) & (g1685) & (!g677) & (g726)) + ((g1682) & (!g1683) & (g1684) & (g1685) & (g677) & (g726)) + ((g1682) & (g1683) & (!g1684) & (!g1685) & (!g677) & (!g726)) + ((g1682) & (g1683) & (!g1684) & (!g1685) & (g677) & (!g726)) + ((g1682) & (g1683) & (!g1684) & (g1685) & (!g677) & (!g726)) + ((g1682) & (g1683) & (!g1684) & (g1685) & (g677) & (!g726)) + ((g1682) & (g1683) & (!g1684) & (g1685) & (g677) & (g726)) + ((g1682) & (g1683) & (g1684) & (!g1685) & (!g677) & (!g726)) + ((g1682) & (g1683) & (g1684) & (!g1685) & (!g677) & (g726)) + ((g1682) & (g1683) & (g1684) & (!g1685) & (g677) & (!g726)) + ((g1682) & (g1683) & (g1684) & (g1685) & (!g677) & (!g726)) + ((g1682) & (g1683) & (g1684) & (g1685) & (!g677) & (g726)) + ((g1682) & (g1683) & (g1684) & (g1685) & (g677) & (!g726)) + ((g1682) & (g1683) & (g1684) & (g1685) & (g677) & (g726)));
	assign g1687 = (((!g475) & (!g476) & (!g477) & (g478) & (g677) & (g726)) + ((!g475) & (!g476) & (g477) & (!g478) & (!g677) & (g726)) + ((!g475) & (!g476) & (g477) & (g478) & (!g677) & (g726)) + ((!g475) & (!g476) & (g477) & (g478) & (g677) & (g726)) + ((!g475) & (g476) & (!g477) & (!g478) & (g677) & (!g726)) + ((!g475) & (g476) & (!g477) & (g478) & (g677) & (!g726)) + ((!g475) & (g476) & (!g477) & (g478) & (g677) & (g726)) + ((!g475) & (g476) & (g477) & (!g478) & (!g677) & (g726)) + ((!g475) & (g476) & (g477) & (!g478) & (g677) & (!g726)) + ((!g475) & (g476) & (g477) & (g478) & (!g677) & (g726)) + ((!g475) & (g476) & (g477) & (g478) & (g677) & (!g726)) + ((!g475) & (g476) & (g477) & (g478) & (g677) & (g726)) + ((g475) & (!g476) & (!g477) & (!g478) & (!g677) & (!g726)) + ((g475) & (!g476) & (!g477) & (g478) & (!g677) & (!g726)) + ((g475) & (!g476) & (!g477) & (g478) & (g677) & (g726)) + ((g475) & (!g476) & (g477) & (!g478) & (!g677) & (!g726)) + ((g475) & (!g476) & (g477) & (!g478) & (!g677) & (g726)) + ((g475) & (!g476) & (g477) & (g478) & (!g677) & (!g726)) + ((g475) & (!g476) & (g477) & (g478) & (!g677) & (g726)) + ((g475) & (!g476) & (g477) & (g478) & (g677) & (g726)) + ((g475) & (g476) & (!g477) & (!g478) & (!g677) & (!g726)) + ((g475) & (g476) & (!g477) & (!g478) & (g677) & (!g726)) + ((g475) & (g476) & (!g477) & (g478) & (!g677) & (!g726)) + ((g475) & (g476) & (!g477) & (g478) & (g677) & (!g726)) + ((g475) & (g476) & (!g477) & (g478) & (g677) & (g726)) + ((g475) & (g476) & (g477) & (!g478) & (!g677) & (!g726)) + ((g475) & (g476) & (g477) & (!g478) & (!g677) & (g726)) + ((g475) & (g476) & (g477) & (!g478) & (g677) & (!g726)) + ((g475) & (g476) & (g477) & (g478) & (!g677) & (!g726)) + ((g475) & (g476) & (g477) & (g478) & (!g677) & (g726)) + ((g475) & (g476) & (g477) & (g478) & (g677) & (!g726)) + ((g475) & (g476) & (g477) & (g478) & (g677) & (g726)));
	assign g1688 = (((!g677) & (!g726) & (!g480) & (!sk[90]) & (g481) & (!g482)) + ((!g677) & (!g726) & (!g480) & (!sk[90]) & (g481) & (g482)) + ((!g677) & (!g726) & (g480) & (!sk[90]) & (!g481) & (!g482)) + ((!g677) & (!g726) & (g480) & (!sk[90]) & (!g481) & (g482)) + ((!g677) & (!g726) & (g480) & (!sk[90]) & (g481) & (!g482)) + ((!g677) & (!g726) & (g480) & (!sk[90]) & (g481) & (g482)) + ((!g677) & (g726) & (!g480) & (!sk[90]) & (!g481) & (!g482)) + ((!g677) & (g726) & (!g480) & (!sk[90]) & (!g481) & (g482)) + ((!g677) & (g726) & (!g480) & (!sk[90]) & (g481) & (!g482)) + ((!g677) & (g726) & (!g480) & (!sk[90]) & (g481) & (g482)) + ((!g677) & (g726) & (!g480) & (sk[90]) & (!g481) & (g482)) + ((!g677) & (g726) & (!g480) & (sk[90]) & (g481) & (g482)) + ((!g677) & (g726) & (g480) & (!sk[90]) & (!g481) & (!g482)) + ((!g677) & (g726) & (g480) & (!sk[90]) & (!g481) & (g482)) + ((!g677) & (g726) & (g480) & (!sk[90]) & (g481) & (!g482)) + ((!g677) & (g726) & (g480) & (!sk[90]) & (g481) & (g482)) + ((!g677) & (g726) & (g480) & (sk[90]) & (!g481) & (g482)) + ((!g677) & (g726) & (g480) & (sk[90]) & (g481) & (g482)) + ((g677) & (!g726) & (!g480) & (!sk[90]) & (g481) & (!g482)) + ((g677) & (!g726) & (!g480) & (!sk[90]) & (g481) & (g482)) + ((g677) & (!g726) & (g480) & (!sk[90]) & (!g481) & (!g482)) + ((g677) & (!g726) & (g480) & (!sk[90]) & (!g481) & (g482)) + ((g677) & (!g726) & (g480) & (!sk[90]) & (g481) & (!g482)) + ((g677) & (!g726) & (g480) & (!sk[90]) & (g481) & (g482)) + ((g677) & (!g726) & (g480) & (sk[90]) & (!g481) & (!g482)) + ((g677) & (!g726) & (g480) & (sk[90]) & (!g481) & (g482)) + ((g677) & (!g726) & (g480) & (sk[90]) & (g481) & (!g482)) + ((g677) & (!g726) & (g480) & (sk[90]) & (g481) & (g482)) + ((g677) & (g726) & (!g480) & (!sk[90]) & (!g481) & (!g482)) + ((g677) & (g726) & (!g480) & (!sk[90]) & (!g481) & (g482)) + ((g677) & (g726) & (!g480) & (!sk[90]) & (g481) & (!g482)) + ((g677) & (g726) & (!g480) & (!sk[90]) & (g481) & (g482)) + ((g677) & (g726) & (!g480) & (sk[90]) & (g481) & (!g482)) + ((g677) & (g726) & (!g480) & (sk[90]) & (g481) & (g482)) + ((g677) & (g726) & (g480) & (!sk[90]) & (!g481) & (!g482)) + ((g677) & (g726) & (g480) & (!sk[90]) & (!g481) & (g482)) + ((g677) & (g726) & (g480) & (!sk[90]) & (g481) & (!g482)) + ((g677) & (g726) & (g480) & (!sk[90]) & (g481) & (g482)) + ((g677) & (g726) & (g480) & (sk[90]) & (g481) & (!g482)) + ((g677) & (g726) & (g480) & (sk[90]) & (g481) & (g482)));
	assign g1689 = (((!g484) & (!g485) & (!g486) & (g487) & (g677) & (g726)) + ((!g484) & (!g485) & (g486) & (!g487) & (!g677) & (g726)) + ((!g484) & (!g485) & (g486) & (g487) & (!g677) & (g726)) + ((!g484) & (!g485) & (g486) & (g487) & (g677) & (g726)) + ((!g484) & (g485) & (!g486) & (!g487) & (g677) & (!g726)) + ((!g484) & (g485) & (!g486) & (g487) & (g677) & (!g726)) + ((!g484) & (g485) & (!g486) & (g487) & (g677) & (g726)) + ((!g484) & (g485) & (g486) & (!g487) & (!g677) & (g726)) + ((!g484) & (g485) & (g486) & (!g487) & (g677) & (!g726)) + ((!g484) & (g485) & (g486) & (g487) & (!g677) & (g726)) + ((!g484) & (g485) & (g486) & (g487) & (g677) & (!g726)) + ((!g484) & (g485) & (g486) & (g487) & (g677) & (g726)) + ((g484) & (!g485) & (!g486) & (!g487) & (!g677) & (!g726)) + ((g484) & (!g485) & (!g486) & (g487) & (!g677) & (!g726)) + ((g484) & (!g485) & (!g486) & (g487) & (g677) & (g726)) + ((g484) & (!g485) & (g486) & (!g487) & (!g677) & (!g726)) + ((g484) & (!g485) & (g486) & (!g487) & (!g677) & (g726)) + ((g484) & (!g485) & (g486) & (g487) & (!g677) & (!g726)) + ((g484) & (!g485) & (g486) & (g487) & (!g677) & (g726)) + ((g484) & (!g485) & (g486) & (g487) & (g677) & (g726)) + ((g484) & (g485) & (!g486) & (!g487) & (!g677) & (!g726)) + ((g484) & (g485) & (!g486) & (!g487) & (g677) & (!g726)) + ((g484) & (g485) & (!g486) & (g487) & (!g677) & (!g726)) + ((g484) & (g485) & (!g486) & (g487) & (g677) & (!g726)) + ((g484) & (g485) & (!g486) & (g487) & (g677) & (g726)) + ((g484) & (g485) & (g486) & (!g487) & (!g677) & (!g726)) + ((g484) & (g485) & (g486) & (!g487) & (!g677) & (g726)) + ((g484) & (g485) & (g486) & (!g487) & (g677) & (!g726)) + ((g484) & (g485) & (g486) & (g487) & (!g677) & (!g726)) + ((g484) & (g485) & (g486) & (g487) & (!g677) & (g726)) + ((g484) & (g485) & (g486) & (g487) & (g677) & (!g726)) + ((g484) & (g485) & (g486) & (g487) & (g677) & (g726)));
	assign g1690 = (((!g489) & (!g490) & (!g491) & (g492) & (g677) & (g726)) + ((!g489) & (!g490) & (g491) & (!g492) & (!g677) & (g726)) + ((!g489) & (!g490) & (g491) & (g492) & (!g677) & (g726)) + ((!g489) & (!g490) & (g491) & (g492) & (g677) & (g726)) + ((!g489) & (g490) & (!g491) & (!g492) & (g677) & (!g726)) + ((!g489) & (g490) & (!g491) & (g492) & (g677) & (!g726)) + ((!g489) & (g490) & (!g491) & (g492) & (g677) & (g726)) + ((!g489) & (g490) & (g491) & (!g492) & (!g677) & (g726)) + ((!g489) & (g490) & (g491) & (!g492) & (g677) & (!g726)) + ((!g489) & (g490) & (g491) & (g492) & (!g677) & (g726)) + ((!g489) & (g490) & (g491) & (g492) & (g677) & (!g726)) + ((!g489) & (g490) & (g491) & (g492) & (g677) & (g726)) + ((g489) & (!g490) & (!g491) & (!g492) & (!g677) & (!g726)) + ((g489) & (!g490) & (!g491) & (g492) & (!g677) & (!g726)) + ((g489) & (!g490) & (!g491) & (g492) & (g677) & (g726)) + ((g489) & (!g490) & (g491) & (!g492) & (!g677) & (!g726)) + ((g489) & (!g490) & (g491) & (!g492) & (!g677) & (g726)) + ((g489) & (!g490) & (g491) & (g492) & (!g677) & (!g726)) + ((g489) & (!g490) & (g491) & (g492) & (!g677) & (g726)) + ((g489) & (!g490) & (g491) & (g492) & (g677) & (g726)) + ((g489) & (g490) & (!g491) & (!g492) & (!g677) & (!g726)) + ((g489) & (g490) & (!g491) & (!g492) & (g677) & (!g726)) + ((g489) & (g490) & (!g491) & (g492) & (!g677) & (!g726)) + ((g489) & (g490) & (!g491) & (g492) & (g677) & (!g726)) + ((g489) & (g490) & (!g491) & (g492) & (g677) & (g726)) + ((g489) & (g490) & (g491) & (!g492) & (!g677) & (!g726)) + ((g489) & (g490) & (g491) & (!g492) & (!g677) & (g726)) + ((g489) & (g490) & (g491) & (!g492) & (g677) & (!g726)) + ((g489) & (g490) & (g491) & (g492) & (!g677) & (!g726)) + ((g489) & (g490) & (g491) & (g492) & (!g677) & (g726)) + ((g489) & (g490) & (g491) & (g492) & (g677) & (!g726)) + ((g489) & (g490) & (g491) & (g492) & (g677) & (g726)));
	assign g1691 = (((!g820) & (!g773) & (!g1687) & (g1688) & (!g1689) & (!g1690)) + ((!g820) & (!g773) & (!g1687) & (g1688) & (!g1689) & (g1690)) + ((!g820) & (!g773) & (!g1687) & (g1688) & (g1689) & (!g1690)) + ((!g820) & (!g773) & (!g1687) & (g1688) & (g1689) & (g1690)) + ((!g820) & (!g773) & (g1687) & (g1688) & (!g1689) & (!g1690)) + ((!g820) & (!g773) & (g1687) & (g1688) & (!g1689) & (g1690)) + ((!g820) & (!g773) & (g1687) & (g1688) & (g1689) & (!g1690)) + ((!g820) & (!g773) & (g1687) & (g1688) & (g1689) & (g1690)) + ((!g820) & (g773) & (!g1687) & (!g1688) & (!g1689) & (g1690)) + ((!g820) & (g773) & (!g1687) & (!g1688) & (g1689) & (g1690)) + ((!g820) & (g773) & (!g1687) & (g1688) & (!g1689) & (g1690)) + ((!g820) & (g773) & (!g1687) & (g1688) & (g1689) & (g1690)) + ((!g820) & (g773) & (g1687) & (!g1688) & (!g1689) & (g1690)) + ((!g820) & (g773) & (g1687) & (!g1688) & (g1689) & (g1690)) + ((!g820) & (g773) & (g1687) & (g1688) & (!g1689) & (g1690)) + ((!g820) & (g773) & (g1687) & (g1688) & (g1689) & (g1690)) + ((g820) & (!g773) & (g1687) & (!g1688) & (!g1689) & (!g1690)) + ((g820) & (!g773) & (g1687) & (!g1688) & (!g1689) & (g1690)) + ((g820) & (!g773) & (g1687) & (!g1688) & (g1689) & (!g1690)) + ((g820) & (!g773) & (g1687) & (!g1688) & (g1689) & (g1690)) + ((g820) & (!g773) & (g1687) & (g1688) & (!g1689) & (!g1690)) + ((g820) & (!g773) & (g1687) & (g1688) & (!g1689) & (g1690)) + ((g820) & (!g773) & (g1687) & (g1688) & (g1689) & (!g1690)) + ((g820) & (!g773) & (g1687) & (g1688) & (g1689) & (g1690)) + ((g820) & (g773) & (!g1687) & (!g1688) & (g1689) & (!g1690)) + ((g820) & (g773) & (!g1687) & (!g1688) & (g1689) & (g1690)) + ((g820) & (g773) & (!g1687) & (g1688) & (g1689) & (!g1690)) + ((g820) & (g773) & (!g1687) & (g1688) & (g1689) & (g1690)) + ((g820) & (g773) & (g1687) & (!g1688) & (g1689) & (!g1690)) + ((g820) & (g773) & (g1687) & (!g1688) & (g1689) & (g1690)) + ((g820) & (g773) & (g1687) & (g1688) & (g1689) & (!g1690)) + ((g820) & (g773) & (g1687) & (g1688) & (g1689) & (g1690)));
	assign g1692 = (((!g867) & (!g1686) & (!sk[94]) & (g1691)) + ((!g867) & (!g1686) & (sk[94]) & (g1691)) + ((!g867) & (g1686) & (!sk[94]) & (!g1691)) + ((!g867) & (g1686) & (!sk[94]) & (g1691)) + ((!g867) & (g1686) & (sk[94]) & (g1691)) + ((g867) & (!g1686) & (!sk[94]) & (g1691)) + ((g867) & (g1686) & (!sk[94]) & (!g1691)) + ((g867) & (g1686) & (!sk[94]) & (g1691)) + ((g867) & (g1686) & (sk[94]) & (!g1691)) + ((g867) & (g1686) & (sk[94]) & (g1691)));
	assign g1693 = (((!g1592) & (!g1593) & (!g1605) & (g1607) & (!g42) & (g1692)) + ((!g1592) & (!g1593) & (!g1605) & (g1607) & (g42) & (g1692)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (!g42) & (g1692)) + ((!g1592) & (!g1593) & (g1605) & (g1607) & (g42) & (g1692)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (!g42) & (g1692)) + ((!g1592) & (g1593) & (!g1605) & (g1607) & (g42) & (g1692)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (!g42) & (g1692)) + ((!g1592) & (g1593) & (g1605) & (g1607) & (g42) & (g1692)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (!g42) & (g1692)) + ((g1592) & (!g1593) & (g1605) & (g1607) & (g42) & (g1692)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g42) & (!g1692)) + ((g1592) & (g1593) & (!g1605) & (g1607) & (g42) & (g1692)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g42) & (!g1692)) + ((g1592) & (g1593) & (g1605) & (g1607) & (g42) & (g1692)));
	assign g1694 = (((!g1592) & (!sk[96]) & (!g1593) & (!g1604) & (g43)) + ((!g1592) & (!sk[96]) & (!g1593) & (g1604) & (!g43)) + ((!g1592) & (!sk[96]) & (!g1593) & (g1604) & (g43)) + ((!g1592) & (!sk[96]) & (g1593) & (!g1604) & (!g43)) + ((!g1592) & (!sk[96]) & (g1593) & (!g1604) & (g43)) + ((!g1592) & (!sk[96]) & (g1593) & (g1604) & (!g43)) + ((!g1592) & (!sk[96]) & (g1593) & (g1604) & (g43)) + ((!g1592) & (sk[96]) & (!g1593) & (g1604) & (!g43)) + ((!g1592) & (sk[96]) & (!g1593) & (g1604) & (g43)) + ((!g1592) & (sk[96]) & (g1593) & (g1604) & (!g43)) + ((!g1592) & (sk[96]) & (g1593) & (g1604) & (g43)) + ((g1592) & (!sk[96]) & (!g1593) & (!g1604) & (g43)) + ((g1592) & (!sk[96]) & (!g1593) & (g1604) & (!g43)) + ((g1592) & (!sk[96]) & (!g1593) & (g1604) & (g43)) + ((g1592) & (!sk[96]) & (g1593) & (!g1604) & (!g43)) + ((g1592) & (!sk[96]) & (g1593) & (!g1604) & (g43)) + ((g1592) & (!sk[96]) & (g1593) & (g1604) & (!g43)) + ((g1592) & (!sk[96]) & (g1593) & (g1604) & (g43)) + ((g1592) & (sk[96]) & (g1593) & (!g1604) & (g43)) + ((g1592) & (sk[96]) & (g1593) & (g1604) & (g43)));
	assign g1695 = (((!g498) & (!g499) & (!g500) & (g501) & (g820) & (g773)) + ((!g498) & (!g499) & (g500) & (!g501) & (!g820) & (g773)) + ((!g498) & (!g499) & (g500) & (g501) & (!g820) & (g773)) + ((!g498) & (!g499) & (g500) & (g501) & (g820) & (g773)) + ((!g498) & (g499) & (!g500) & (!g501) & (g820) & (!g773)) + ((!g498) & (g499) & (!g500) & (g501) & (g820) & (!g773)) + ((!g498) & (g499) & (!g500) & (g501) & (g820) & (g773)) + ((!g498) & (g499) & (g500) & (!g501) & (!g820) & (g773)) + ((!g498) & (g499) & (g500) & (!g501) & (g820) & (!g773)) + ((!g498) & (g499) & (g500) & (g501) & (!g820) & (g773)) + ((!g498) & (g499) & (g500) & (g501) & (g820) & (!g773)) + ((!g498) & (g499) & (g500) & (g501) & (g820) & (g773)) + ((g498) & (!g499) & (!g500) & (!g501) & (!g820) & (!g773)) + ((g498) & (!g499) & (!g500) & (g501) & (!g820) & (!g773)) + ((g498) & (!g499) & (!g500) & (g501) & (g820) & (g773)) + ((g498) & (!g499) & (g500) & (!g501) & (!g820) & (!g773)) + ((g498) & (!g499) & (g500) & (!g501) & (!g820) & (g773)) + ((g498) & (!g499) & (g500) & (g501) & (!g820) & (!g773)) + ((g498) & (!g499) & (g500) & (g501) & (!g820) & (g773)) + ((g498) & (!g499) & (g500) & (g501) & (g820) & (g773)) + ((g498) & (g499) & (!g500) & (!g501) & (!g820) & (!g773)) + ((g498) & (g499) & (!g500) & (!g501) & (g820) & (!g773)) + ((g498) & (g499) & (!g500) & (g501) & (!g820) & (!g773)) + ((g498) & (g499) & (!g500) & (g501) & (g820) & (!g773)) + ((g498) & (g499) & (!g500) & (g501) & (g820) & (g773)) + ((g498) & (g499) & (g500) & (!g501) & (!g820) & (!g773)) + ((g498) & (g499) & (g500) & (!g501) & (!g820) & (g773)) + ((g498) & (g499) & (g500) & (!g501) & (g820) & (!g773)) + ((g498) & (g499) & (g500) & (g501) & (!g820) & (!g773)) + ((g498) & (g499) & (g500) & (g501) & (!g820) & (g773)) + ((g498) & (g499) & (g500) & (g501) & (g820) & (!g773)) + ((g498) & (g499) & (g500) & (g501) & (g820) & (g773)));
	assign g1696 = (((!g503) & (!g504) & (!g505) & (g506) & (g820) & (g773)) + ((!g503) & (!g504) & (g505) & (!g506) & (!g820) & (g773)) + ((!g503) & (!g504) & (g505) & (g506) & (!g820) & (g773)) + ((!g503) & (!g504) & (g505) & (g506) & (g820) & (g773)) + ((!g503) & (g504) & (!g505) & (!g506) & (g820) & (!g773)) + ((!g503) & (g504) & (!g505) & (g506) & (g820) & (!g773)) + ((!g503) & (g504) & (!g505) & (g506) & (g820) & (g773)) + ((!g503) & (g504) & (g505) & (!g506) & (!g820) & (g773)) + ((!g503) & (g504) & (g505) & (!g506) & (g820) & (!g773)) + ((!g503) & (g504) & (g505) & (g506) & (!g820) & (g773)) + ((!g503) & (g504) & (g505) & (g506) & (g820) & (!g773)) + ((!g503) & (g504) & (g505) & (g506) & (g820) & (g773)) + ((g503) & (!g504) & (!g505) & (!g506) & (!g820) & (!g773)) + ((g503) & (!g504) & (!g505) & (g506) & (!g820) & (!g773)) + ((g503) & (!g504) & (!g505) & (g506) & (g820) & (g773)) + ((g503) & (!g504) & (g505) & (!g506) & (!g820) & (!g773)) + ((g503) & (!g504) & (g505) & (!g506) & (!g820) & (g773)) + ((g503) & (!g504) & (g505) & (g506) & (!g820) & (!g773)) + ((g503) & (!g504) & (g505) & (g506) & (!g820) & (g773)) + ((g503) & (!g504) & (g505) & (g506) & (g820) & (g773)) + ((g503) & (g504) & (!g505) & (!g506) & (!g820) & (!g773)) + ((g503) & (g504) & (!g505) & (!g506) & (g820) & (!g773)) + ((g503) & (g504) & (!g505) & (g506) & (!g820) & (!g773)) + ((g503) & (g504) & (!g505) & (g506) & (g820) & (!g773)) + ((g503) & (g504) & (!g505) & (g506) & (g820) & (g773)) + ((g503) & (g504) & (g505) & (!g506) & (!g820) & (!g773)) + ((g503) & (g504) & (g505) & (!g506) & (!g820) & (g773)) + ((g503) & (g504) & (g505) & (!g506) & (g820) & (!g773)) + ((g503) & (g504) & (g505) & (g506) & (!g820) & (!g773)) + ((g503) & (g504) & (g505) & (g506) & (!g820) & (g773)) + ((g503) & (g504) & (g505) & (g506) & (g820) & (!g773)) + ((g503) & (g504) & (g505) & (g506) & (g820) & (g773)));
	assign g1697 = (((!g508) & (!g509) & (!g510) & (g511) & (g820) & (g773)) + ((!g508) & (!g509) & (g510) & (!g511) & (!g820) & (g773)) + ((!g508) & (!g509) & (g510) & (g511) & (!g820) & (g773)) + ((!g508) & (!g509) & (g510) & (g511) & (g820) & (g773)) + ((!g508) & (g509) & (!g510) & (!g511) & (g820) & (!g773)) + ((!g508) & (g509) & (!g510) & (g511) & (g820) & (!g773)) + ((!g508) & (g509) & (!g510) & (g511) & (g820) & (g773)) + ((!g508) & (g509) & (g510) & (!g511) & (!g820) & (g773)) + ((!g508) & (g509) & (g510) & (!g511) & (g820) & (!g773)) + ((!g508) & (g509) & (g510) & (g511) & (!g820) & (g773)) + ((!g508) & (g509) & (g510) & (g511) & (g820) & (!g773)) + ((!g508) & (g509) & (g510) & (g511) & (g820) & (g773)) + ((g508) & (!g509) & (!g510) & (!g511) & (!g820) & (!g773)) + ((g508) & (!g509) & (!g510) & (g511) & (!g820) & (!g773)) + ((g508) & (!g509) & (!g510) & (g511) & (g820) & (g773)) + ((g508) & (!g509) & (g510) & (!g511) & (!g820) & (!g773)) + ((g508) & (!g509) & (g510) & (!g511) & (!g820) & (g773)) + ((g508) & (!g509) & (g510) & (g511) & (!g820) & (!g773)) + ((g508) & (!g509) & (g510) & (g511) & (!g820) & (g773)) + ((g508) & (!g509) & (g510) & (g511) & (g820) & (g773)) + ((g508) & (g509) & (!g510) & (!g511) & (!g820) & (!g773)) + ((g508) & (g509) & (!g510) & (!g511) & (g820) & (!g773)) + ((g508) & (g509) & (!g510) & (g511) & (!g820) & (!g773)) + ((g508) & (g509) & (!g510) & (g511) & (g820) & (!g773)) + ((g508) & (g509) & (!g510) & (g511) & (g820) & (g773)) + ((g508) & (g509) & (g510) & (!g511) & (!g820) & (!g773)) + ((g508) & (g509) & (g510) & (!g511) & (!g820) & (g773)) + ((g508) & (g509) & (g510) & (!g511) & (g820) & (!g773)) + ((g508) & (g509) & (g510) & (g511) & (!g820) & (!g773)) + ((g508) & (g509) & (g510) & (g511) & (!g820) & (g773)) + ((g508) & (g509) & (g510) & (g511) & (g820) & (!g773)) + ((g508) & (g509) & (g510) & (g511) & (g820) & (g773)));
	assign g1698 = (((!g513) & (!g514) & (!g515) & (g516) & (g820) & (g773)) + ((!g513) & (!g514) & (g515) & (!g516) & (!g820) & (g773)) + ((!g513) & (!g514) & (g515) & (g516) & (!g820) & (g773)) + ((!g513) & (!g514) & (g515) & (g516) & (g820) & (g773)) + ((!g513) & (g514) & (!g515) & (!g516) & (g820) & (!g773)) + ((!g513) & (g514) & (!g515) & (g516) & (g820) & (!g773)) + ((!g513) & (g514) & (!g515) & (g516) & (g820) & (g773)) + ((!g513) & (g514) & (g515) & (!g516) & (!g820) & (g773)) + ((!g513) & (g514) & (g515) & (!g516) & (g820) & (!g773)) + ((!g513) & (g514) & (g515) & (g516) & (!g820) & (g773)) + ((!g513) & (g514) & (g515) & (g516) & (g820) & (!g773)) + ((!g513) & (g514) & (g515) & (g516) & (g820) & (g773)) + ((g513) & (!g514) & (!g515) & (!g516) & (!g820) & (!g773)) + ((g513) & (!g514) & (!g515) & (g516) & (!g820) & (!g773)) + ((g513) & (!g514) & (!g515) & (g516) & (g820) & (g773)) + ((g513) & (!g514) & (g515) & (!g516) & (!g820) & (!g773)) + ((g513) & (!g514) & (g515) & (!g516) & (!g820) & (g773)) + ((g513) & (!g514) & (g515) & (g516) & (!g820) & (!g773)) + ((g513) & (!g514) & (g515) & (g516) & (!g820) & (g773)) + ((g513) & (!g514) & (g515) & (g516) & (g820) & (g773)) + ((g513) & (g514) & (!g515) & (!g516) & (!g820) & (!g773)) + ((g513) & (g514) & (!g515) & (!g516) & (g820) & (!g773)) + ((g513) & (g514) & (!g515) & (g516) & (!g820) & (!g773)) + ((g513) & (g514) & (!g515) & (g516) & (g820) & (!g773)) + ((g513) & (g514) & (!g515) & (g516) & (g820) & (g773)) + ((g513) & (g514) & (g515) & (!g516) & (!g820) & (!g773)) + ((g513) & (g514) & (g515) & (!g516) & (!g820) & (g773)) + ((g513) & (g514) & (g515) & (!g516) & (g820) & (!g773)) + ((g513) & (g514) & (g515) & (g516) & (!g820) & (!g773)) + ((g513) & (g514) & (g515) & (g516) & (!g820) & (g773)) + ((g513) & (g514) & (g515) & (g516) & (g820) & (!g773)) + ((g513) & (g514) & (g515) & (g516) & (g820) & (g773)));
	assign g1699 = (((!g1695) & (!g1696) & (!g1697) & (g1698) & (g677) & (g726)) + ((!g1695) & (!g1696) & (g1697) & (!g1698) & (!g677) & (g726)) + ((!g1695) & (!g1696) & (g1697) & (g1698) & (!g677) & (g726)) + ((!g1695) & (!g1696) & (g1697) & (g1698) & (g677) & (g726)) + ((!g1695) & (g1696) & (!g1697) & (!g1698) & (g677) & (!g726)) + ((!g1695) & (g1696) & (!g1697) & (g1698) & (g677) & (!g726)) + ((!g1695) & (g1696) & (!g1697) & (g1698) & (g677) & (g726)) + ((!g1695) & (g1696) & (g1697) & (!g1698) & (!g677) & (g726)) + ((!g1695) & (g1696) & (g1697) & (!g1698) & (g677) & (!g726)) + ((!g1695) & (g1696) & (g1697) & (g1698) & (!g677) & (g726)) + ((!g1695) & (g1696) & (g1697) & (g1698) & (g677) & (!g726)) + ((!g1695) & (g1696) & (g1697) & (g1698) & (g677) & (g726)) + ((g1695) & (!g1696) & (!g1697) & (!g1698) & (!g677) & (!g726)) + ((g1695) & (!g1696) & (!g1697) & (g1698) & (!g677) & (!g726)) + ((g1695) & (!g1696) & (!g1697) & (g1698) & (g677) & (g726)) + ((g1695) & (!g1696) & (g1697) & (!g1698) & (!g677) & (!g726)) + ((g1695) & (!g1696) & (g1697) & (!g1698) & (!g677) & (g726)) + ((g1695) & (!g1696) & (g1697) & (g1698) & (!g677) & (!g726)) + ((g1695) & (!g1696) & (g1697) & (g1698) & (!g677) & (g726)) + ((g1695) & (!g1696) & (g1697) & (g1698) & (g677) & (g726)) + ((g1695) & (g1696) & (!g1697) & (!g1698) & (!g677) & (!g726)) + ((g1695) & (g1696) & (!g1697) & (!g1698) & (g677) & (!g726)) + ((g1695) & (g1696) & (!g1697) & (g1698) & (!g677) & (!g726)) + ((g1695) & (g1696) & (!g1697) & (g1698) & (g677) & (!g726)) + ((g1695) & (g1696) & (!g1697) & (g1698) & (g677) & (g726)) + ((g1695) & (g1696) & (g1697) & (!g1698) & (!g677) & (!g726)) + ((g1695) & (g1696) & (g1697) & (!g1698) & (!g677) & (g726)) + ((g1695) & (g1696) & (g1697) & (!g1698) & (g677) & (!g726)) + ((g1695) & (g1696) & (g1697) & (g1698) & (!g677) & (!g726)) + ((g1695) & (g1696) & (g1697) & (g1698) & (!g677) & (g726)) + ((g1695) & (g1696) & (g1697) & (g1698) & (g677) & (!g726)) + ((g1695) & (g1696) & (g1697) & (g1698) & (g677) & (g726)));
	assign g1700 = (((!g519) & (!g520) & (!g521) & (g522) & (g677) & (g726)) + ((!g519) & (!g520) & (g521) & (!g522) & (!g677) & (g726)) + ((!g519) & (!g520) & (g521) & (g522) & (!g677) & (g726)) + ((!g519) & (!g520) & (g521) & (g522) & (g677) & (g726)) + ((!g519) & (g520) & (!g521) & (!g522) & (g677) & (!g726)) + ((!g519) & (g520) & (!g521) & (g522) & (g677) & (!g726)) + ((!g519) & (g520) & (!g521) & (g522) & (g677) & (g726)) + ((!g519) & (g520) & (g521) & (!g522) & (!g677) & (g726)) + ((!g519) & (g520) & (g521) & (!g522) & (g677) & (!g726)) + ((!g519) & (g520) & (g521) & (g522) & (!g677) & (g726)) + ((!g519) & (g520) & (g521) & (g522) & (g677) & (!g726)) + ((!g519) & (g520) & (g521) & (g522) & (g677) & (g726)) + ((g519) & (!g520) & (!g521) & (!g522) & (!g677) & (!g726)) + ((g519) & (!g520) & (!g521) & (g522) & (!g677) & (!g726)) + ((g519) & (!g520) & (!g521) & (g522) & (g677) & (g726)) + ((g519) & (!g520) & (g521) & (!g522) & (!g677) & (!g726)) + ((g519) & (!g520) & (g521) & (!g522) & (!g677) & (g726)) + ((g519) & (!g520) & (g521) & (g522) & (!g677) & (!g726)) + ((g519) & (!g520) & (g521) & (g522) & (!g677) & (g726)) + ((g519) & (!g520) & (g521) & (g522) & (g677) & (g726)) + ((g519) & (g520) & (!g521) & (!g522) & (!g677) & (!g726)) + ((g519) & (g520) & (!g521) & (!g522) & (g677) & (!g726)) + ((g519) & (g520) & (!g521) & (g522) & (!g677) & (!g726)) + ((g519) & (g520) & (!g521) & (g522) & (g677) & (!g726)) + ((g519) & (g520) & (!g521) & (g522) & (g677) & (g726)) + ((g519) & (g520) & (g521) & (!g522) & (!g677) & (!g726)) + ((g519) & (g520) & (g521) & (!g522) & (!g677) & (g726)) + ((g519) & (g520) & (g521) & (!g522) & (g677) & (!g726)) + ((g519) & (g520) & (g521) & (g522) & (!g677) & (!g726)) + ((g519) & (g520) & (g521) & (g522) & (!g677) & (g726)) + ((g519) & (g520) & (g521) & (g522) & (g677) & (!g726)) + ((g519) & (g520) & (g521) & (g522) & (g677) & (g726)));
	assign g1701 = (((!g677) & (!g726) & (!g524) & (!sk[103]) & (g525) & (!g526)) + ((!g677) & (!g726) & (!g524) & (!sk[103]) & (g525) & (g526)) + ((!g677) & (!g726) & (g524) & (!sk[103]) & (!g525) & (!g526)) + ((!g677) & (!g726) & (g524) & (!sk[103]) & (!g525) & (g526)) + ((!g677) & (!g726) & (g524) & (!sk[103]) & (g525) & (!g526)) + ((!g677) & (!g726) & (g524) & (!sk[103]) & (g525) & (g526)) + ((!g677) & (g726) & (!g524) & (!sk[103]) & (!g525) & (!g526)) + ((!g677) & (g726) & (!g524) & (!sk[103]) & (!g525) & (g526)) + ((!g677) & (g726) & (!g524) & (!sk[103]) & (g525) & (!g526)) + ((!g677) & (g726) & (!g524) & (!sk[103]) & (g525) & (g526)) + ((!g677) & (g726) & (!g524) & (sk[103]) & (!g525) & (g526)) + ((!g677) & (g726) & (!g524) & (sk[103]) & (g525) & (g526)) + ((!g677) & (g726) & (g524) & (!sk[103]) & (!g525) & (!g526)) + ((!g677) & (g726) & (g524) & (!sk[103]) & (!g525) & (g526)) + ((!g677) & (g726) & (g524) & (!sk[103]) & (g525) & (!g526)) + ((!g677) & (g726) & (g524) & (!sk[103]) & (g525) & (g526)) + ((!g677) & (g726) & (g524) & (sk[103]) & (!g525) & (g526)) + ((!g677) & (g726) & (g524) & (sk[103]) & (g525) & (g526)) + ((g677) & (!g726) & (!g524) & (!sk[103]) & (g525) & (!g526)) + ((g677) & (!g726) & (!g524) & (!sk[103]) & (g525) & (g526)) + ((g677) & (!g726) & (g524) & (!sk[103]) & (!g525) & (!g526)) + ((g677) & (!g726) & (g524) & (!sk[103]) & (!g525) & (g526)) + ((g677) & (!g726) & (g524) & (!sk[103]) & (g525) & (!g526)) + ((g677) & (!g726) & (g524) & (!sk[103]) & (g525) & (g526)) + ((g677) & (!g726) & (g524) & (sk[103]) & (!g525) & (!g526)) + ((g677) & (!g726) & (g524) & (sk[103]) & (!g525) & (g526)) + ((g677) & (!g726) & (g524) & (sk[103]) & (g525) & (!g526)) + ((g677) & (!g726) & (g524) & (sk[103]) & (g525) & (g526)) + ((g677) & (g726) & (!g524) & (!sk[103]) & (!g525) & (!g526)) + ((g677) & (g726) & (!g524) & (!sk[103]) & (!g525) & (g526)) + ((g677) & (g726) & (!g524) & (!sk[103]) & (g525) & (!g526)) + ((g677) & (g726) & (!g524) & (!sk[103]) & (g525) & (g526)) + ((g677) & (g726) & (!g524) & (sk[103]) & (g525) & (!g526)) + ((g677) & (g726) & (!g524) & (sk[103]) & (g525) & (g526)) + ((g677) & (g726) & (g524) & (!sk[103]) & (!g525) & (!g526)) + ((g677) & (g726) & (g524) & (!sk[103]) & (!g525) & (g526)) + ((g677) & (g726) & (g524) & (!sk[103]) & (g525) & (!g526)) + ((g677) & (g726) & (g524) & (!sk[103]) & (g525) & (g526)) + ((g677) & (g726) & (g524) & (sk[103]) & (g525) & (!g526)) + ((g677) & (g726) & (g524) & (sk[103]) & (g525) & (g526)));
	assign g1702 = (((!g528) & (!g529) & (!g530) & (g531) & (g677) & (g726)) + ((!g528) & (!g529) & (g530) & (!g531) & (!g677) & (g726)) + ((!g528) & (!g529) & (g530) & (g531) & (!g677) & (g726)) + ((!g528) & (!g529) & (g530) & (g531) & (g677) & (g726)) + ((!g528) & (g529) & (!g530) & (!g531) & (g677) & (!g726)) + ((!g528) & (g529) & (!g530) & (g531) & (g677) & (!g726)) + ((!g528) & (g529) & (!g530) & (g531) & (g677) & (g726)) + ((!g528) & (g529) & (g530) & (!g531) & (!g677) & (g726)) + ((!g528) & (g529) & (g530) & (!g531) & (g677) & (!g726)) + ((!g528) & (g529) & (g530) & (g531) & (!g677) & (g726)) + ((!g528) & (g529) & (g530) & (g531) & (g677) & (!g726)) + ((!g528) & (g529) & (g530) & (g531) & (g677) & (g726)) + ((g528) & (!g529) & (!g530) & (!g531) & (!g677) & (!g726)) + ((g528) & (!g529) & (!g530) & (g531) & (!g677) & (!g726)) + ((g528) & (!g529) & (!g530) & (g531) & (g677) & (g726)) + ((g528) & (!g529) & (g530) & (!g531) & (!g677) & (!g726)) + ((g528) & (!g529) & (g530) & (!g531) & (!g677) & (g726)) + ((g528) & (!g529) & (g530) & (g531) & (!g677) & (!g726)) + ((g528) & (!g529) & (g530) & (g531) & (!g677) & (g726)) + ((g528) & (!g529) & (g530) & (g531) & (g677) & (g726)) + ((g528) & (g529) & (!g530) & (!g531) & (!g677) & (!g726)) + ((g528) & (g529) & (!g530) & (!g531) & (g677) & (!g726)) + ((g528) & (g529) & (!g530) & (g531) & (!g677) & (!g726)) + ((g528) & (g529) & (!g530) & (g531) & (g677) & (!g726)) + ((g528) & (g529) & (!g530) & (g531) & (g677) & (g726)) + ((g528) & (g529) & (g530) & (!g531) & (!g677) & (!g726)) + ((g528) & (g529) & (g530) & (!g531) & (!g677) & (g726)) + ((g528) & (g529) & (g530) & (!g531) & (g677) & (!g726)) + ((g528) & (g529) & (g530) & (g531) & (!g677) & (!g726)) + ((g528) & (g529) & (g530) & (g531) & (!g677) & (g726)) + ((g528) & (g529) & (g530) & (g531) & (g677) & (!g726)) + ((g528) & (g529) & (g530) & (g531) & (g677) & (g726)));
	assign g1703 = (((!g533) & (!g534) & (!g535) & (g536) & (g677) & (g726)) + ((!g533) & (!g534) & (g535) & (!g536) & (!g677) & (g726)) + ((!g533) & (!g534) & (g535) & (g536) & (!g677) & (g726)) + ((!g533) & (!g534) & (g535) & (g536) & (g677) & (g726)) + ((!g533) & (g534) & (!g535) & (!g536) & (g677) & (!g726)) + ((!g533) & (g534) & (!g535) & (g536) & (g677) & (!g726)) + ((!g533) & (g534) & (!g535) & (g536) & (g677) & (g726)) + ((!g533) & (g534) & (g535) & (!g536) & (!g677) & (g726)) + ((!g533) & (g534) & (g535) & (!g536) & (g677) & (!g726)) + ((!g533) & (g534) & (g535) & (g536) & (!g677) & (g726)) + ((!g533) & (g534) & (g535) & (g536) & (g677) & (!g726)) + ((!g533) & (g534) & (g535) & (g536) & (g677) & (g726)) + ((g533) & (!g534) & (!g535) & (!g536) & (!g677) & (!g726)) + ((g533) & (!g534) & (!g535) & (g536) & (!g677) & (!g726)) + ((g533) & (!g534) & (!g535) & (g536) & (g677) & (g726)) + ((g533) & (!g534) & (g535) & (!g536) & (!g677) & (!g726)) + ((g533) & (!g534) & (g535) & (!g536) & (!g677) & (g726)) + ((g533) & (!g534) & (g535) & (g536) & (!g677) & (!g726)) + ((g533) & (!g534) & (g535) & (g536) & (!g677) & (g726)) + ((g533) & (!g534) & (g535) & (g536) & (g677) & (g726)) + ((g533) & (g534) & (!g535) & (!g536) & (!g677) & (!g726)) + ((g533) & (g534) & (!g535) & (!g536) & (g677) & (!g726)) + ((g533) & (g534) & (!g535) & (g536) & (!g677) & (!g726)) + ((g533) & (g534) & (!g535) & (g536) & (g677) & (!g726)) + ((g533) & (g534) & (!g535) & (g536) & (g677) & (g726)) + ((g533) & (g534) & (g535) & (!g536) & (!g677) & (!g726)) + ((g533) & (g534) & (g535) & (!g536) & (!g677) & (g726)) + ((g533) & (g534) & (g535) & (!g536) & (g677) & (!g726)) + ((g533) & (g534) & (g535) & (g536) & (!g677) & (!g726)) + ((g533) & (g534) & (g535) & (g536) & (!g677) & (g726)) + ((g533) & (g534) & (g535) & (g536) & (g677) & (!g726)) + ((g533) & (g534) & (g535) & (g536) & (g677) & (g726)));
	assign g1704 = (((!g820) & (!g773) & (!g1700) & (g1701) & (!g1702) & (!g1703)) + ((!g820) & (!g773) & (!g1700) & (g1701) & (!g1702) & (g1703)) + ((!g820) & (!g773) & (!g1700) & (g1701) & (g1702) & (!g1703)) + ((!g820) & (!g773) & (!g1700) & (g1701) & (g1702) & (g1703)) + ((!g820) & (!g773) & (g1700) & (g1701) & (!g1702) & (!g1703)) + ((!g820) & (!g773) & (g1700) & (g1701) & (!g1702) & (g1703)) + ((!g820) & (!g773) & (g1700) & (g1701) & (g1702) & (!g1703)) + ((!g820) & (!g773) & (g1700) & (g1701) & (g1702) & (g1703)) + ((!g820) & (g773) & (!g1700) & (!g1701) & (!g1702) & (g1703)) + ((!g820) & (g773) & (!g1700) & (!g1701) & (g1702) & (g1703)) + ((!g820) & (g773) & (!g1700) & (g1701) & (!g1702) & (g1703)) + ((!g820) & (g773) & (!g1700) & (g1701) & (g1702) & (g1703)) + ((!g820) & (g773) & (g1700) & (!g1701) & (!g1702) & (g1703)) + ((!g820) & (g773) & (g1700) & (!g1701) & (g1702) & (g1703)) + ((!g820) & (g773) & (g1700) & (g1701) & (!g1702) & (g1703)) + ((!g820) & (g773) & (g1700) & (g1701) & (g1702) & (g1703)) + ((g820) & (!g773) & (g1700) & (!g1701) & (!g1702) & (!g1703)) + ((g820) & (!g773) & (g1700) & (!g1701) & (!g1702) & (g1703)) + ((g820) & (!g773) & (g1700) & (!g1701) & (g1702) & (!g1703)) + ((g820) & (!g773) & (g1700) & (!g1701) & (g1702) & (g1703)) + ((g820) & (!g773) & (g1700) & (g1701) & (!g1702) & (!g1703)) + ((g820) & (!g773) & (g1700) & (g1701) & (!g1702) & (g1703)) + ((g820) & (!g773) & (g1700) & (g1701) & (g1702) & (!g1703)) + ((g820) & (!g773) & (g1700) & (g1701) & (g1702) & (g1703)) + ((g820) & (g773) & (!g1700) & (!g1701) & (g1702) & (!g1703)) + ((g820) & (g773) & (!g1700) & (!g1701) & (g1702) & (g1703)) + ((g820) & (g773) & (!g1700) & (g1701) & (g1702) & (!g1703)) + ((g820) & (g773) & (!g1700) & (g1701) & (g1702) & (g1703)) + ((g820) & (g773) & (g1700) & (!g1701) & (g1702) & (!g1703)) + ((g820) & (g773) & (g1700) & (!g1701) & (g1702) & (g1703)) + ((g820) & (g773) & (g1700) & (g1701) & (g1702) & (!g1703)) + ((g820) & (g773) & (g1700) & (g1701) & (g1702) & (g1703)));
	assign g1705 = (((!g867) & (!sk[107]) & (!g1699) & (g1704)) + ((!g867) & (!sk[107]) & (g1699) & (!g1704)) + ((!g867) & (!sk[107]) & (g1699) & (g1704)) + ((!g867) & (sk[107]) & (!g1699) & (g1704)) + ((!g867) & (sk[107]) & (g1699) & (g1704)) + ((g867) & (!sk[107]) & (!g1699) & (g1704)) + ((g867) & (!sk[107]) & (g1699) & (!g1704)) + ((g867) & (!sk[107]) & (g1699) & (g1704)) + ((g867) & (sk[107]) & (g1699) & (!g1704)) + ((g867) & (sk[107]) & (g1699) & (g1704)));
	assign g1706 = (((!sk[108]) & (!g132) & (!g1592) & (!g1593) & (g1605)) + ((!sk[108]) & (!g132) & (!g1592) & (g1593) & (!g1605)) + ((!sk[108]) & (!g132) & (!g1592) & (g1593) & (g1605)) + ((!sk[108]) & (!g132) & (g1592) & (!g1593) & (!g1605)) + ((!sk[108]) & (!g132) & (g1592) & (!g1593) & (g1605)) + ((!sk[108]) & (!g132) & (g1592) & (g1593) & (!g1605)) + ((!sk[108]) & (!g132) & (g1592) & (g1593) & (g1605)) + ((!sk[108]) & (g132) & (!g1592) & (!g1593) & (g1605)) + ((!sk[108]) & (g132) & (!g1592) & (g1593) & (!g1605)) + ((!sk[108]) & (g132) & (!g1592) & (g1593) & (g1605)) + ((!sk[108]) & (g132) & (g1592) & (!g1593) & (!g1605)) + ((!sk[108]) & (g132) & (g1592) & (!g1593) & (g1605)) + ((!sk[108]) & (g132) & (g1592) & (g1593) & (!g1605)) + ((!sk[108]) & (g132) & (g1592) & (g1593) & (g1605)) + ((sk[108]) & (!g132) & (!g1592) & (!g1593) & (!g1605)) + ((sk[108]) & (!g132) & (!g1592) & (!g1593) & (g1605)) + ((sk[108]) & (!g132) & (!g1592) & (g1593) & (!g1605)) + ((sk[108]) & (!g132) & (!g1592) & (g1593) & (g1605)) + ((sk[108]) & (!g132) & (g1592) & (!g1593) & (!g1605)) + ((sk[108]) & (!g132) & (g1592) & (g1593) & (!g1605)) + ((sk[108]) & (!g132) & (g1592) & (g1593) & (g1605)));
	assign g1707 = (((!g132) & (!g1592) & (g1606) & (!g136) & (!g1593) & (g1605)) + ((!g132) & (g1592) & (!g1606) & (!g136) & (!g1593) & (!g1605)) + ((!g132) & (g1592) & (!g1606) & (!g136) & (!g1593) & (g1605)) + ((!g132) & (g1592) & (!g1606) & (!g136) & (g1593) & (!g1605)) + ((!g132) & (g1592) & (!g1606) & (!g136) & (g1593) & (g1605)) + ((!g132) & (g1592) & (g1606) & (!g136) & (!g1593) & (g1605)) + ((g132) & (!g1592) & (!g1606) & (!g136) & (!g1593) & (!g1605)) + ((g132) & (!g1592) & (!g1606) & (!g136) & (!g1593) & (g1605)) + ((g132) & (!g1592) & (!g1606) & (!g136) & (g1593) & (!g1605)) + ((g132) & (!g1592) & (!g1606) & (!g136) & (g1593) & (g1605)) + ((g132) & (!g1592) & (g1606) & (!g136) & (!g1593) & (g1605)) + ((g132) & (g1592) & (!g1606) & (!g136) & (!g1593) & (!g1605)) + ((g132) & (g1592) & (!g1606) & (!g136) & (!g1593) & (g1605)) + ((g132) & (g1592) & (!g1606) & (!g136) & (g1593) & (!g1605)) + ((g132) & (g1592) & (!g1606) & (!g136) & (g1593) & (g1605)) + ((g132) & (g1592) & (g1606) & (!g136) & (!g1593) & (g1605)));
	assign g1708 = (((!g132) & (!g1694) & (!g1705) & (g1706) & (!sk[110]) & (!g1707)) + ((!g132) & (!g1694) & (!g1705) & (g1706) & (!sk[110]) & (g1707)) + ((!g132) & (!g1694) & (g1705) & (!g1706) & (!sk[110]) & (!g1707)) + ((!g132) & (!g1694) & (g1705) & (!g1706) & (!sk[110]) & (g1707)) + ((!g132) & (!g1694) & (g1705) & (!g1706) & (sk[110]) & (g1707)) + ((!g132) & (!g1694) & (g1705) & (g1706) & (!sk[110]) & (!g1707)) + ((!g132) & (!g1694) & (g1705) & (g1706) & (!sk[110]) & (g1707)) + ((!g132) & (g1694) & (!g1705) & (!g1706) & (!sk[110]) & (!g1707)) + ((!g132) & (g1694) & (!g1705) & (!g1706) & (!sk[110]) & (g1707)) + ((!g132) & (g1694) & (!g1705) & (!g1706) & (sk[110]) & (g1707)) + ((!g132) & (g1694) & (!g1705) & (g1706) & (!sk[110]) & (!g1707)) + ((!g132) & (g1694) & (!g1705) & (g1706) & (!sk[110]) & (g1707)) + ((!g132) & (g1694) & (!g1705) & (g1706) & (sk[110]) & (g1707)) + ((!g132) & (g1694) & (g1705) & (!g1706) & (!sk[110]) & (!g1707)) + ((!g132) & (g1694) & (g1705) & (!g1706) & (!sk[110]) & (g1707)) + ((!g132) & (g1694) & (g1705) & (!g1706) & (sk[110]) & (g1707)) + ((!g132) & (g1694) & (g1705) & (g1706) & (!sk[110]) & (!g1707)) + ((!g132) & (g1694) & (g1705) & (g1706) & (!sk[110]) & (g1707)) + ((!g132) & (g1694) & (g1705) & (g1706) & (sk[110]) & (g1707)) + ((g132) & (!g1694) & (!g1705) & (g1706) & (!sk[110]) & (!g1707)) + ((g132) & (!g1694) & (!g1705) & (g1706) & (!sk[110]) & (g1707)) + ((g132) & (!g1694) & (g1705) & (!g1706) & (!sk[110]) & (!g1707)) + ((g132) & (!g1694) & (g1705) & (!g1706) & (!sk[110]) & (g1707)) + ((g132) & (!g1694) & (g1705) & (!g1706) & (sk[110]) & (g1707)) + ((g132) & (!g1694) & (g1705) & (g1706) & (!sk[110]) & (!g1707)) + ((g132) & (!g1694) & (g1705) & (g1706) & (!sk[110]) & (g1707)) + ((g132) & (g1694) & (!g1705) & (!g1706) & (!sk[110]) & (!g1707)) + ((g132) & (g1694) & (!g1705) & (!g1706) & (!sk[110]) & (g1707)) + ((g132) & (g1694) & (!g1705) & (g1706) & (!sk[110]) & (!g1707)) + ((g132) & (g1694) & (!g1705) & (g1706) & (!sk[110]) & (g1707)) + ((g132) & (g1694) & (g1705) & (!g1706) & (!sk[110]) & (!g1707)) + ((g132) & (g1694) & (g1705) & (!g1706) & (!sk[110]) & (g1707)) + ((g132) & (g1694) & (g1705) & (!g1706) & (sk[110]) & (g1707)) + ((g132) & (g1694) & (g1705) & (g1706) & (!sk[110]) & (!g1707)) + ((g132) & (g1694) & (g1705) & (g1706) & (!sk[110]) & (g1707)));
	assign g1709 = (((!g1592) & (!sk[111]) & (!g1593) & (!g1620) & (g44)) + ((!g1592) & (!sk[111]) & (!g1593) & (g1620) & (!g44)) + ((!g1592) & (!sk[111]) & (!g1593) & (g1620) & (g44)) + ((!g1592) & (!sk[111]) & (g1593) & (!g1620) & (!g44)) + ((!g1592) & (!sk[111]) & (g1593) & (!g1620) & (g44)) + ((!g1592) & (!sk[111]) & (g1593) & (g1620) & (!g44)) + ((!g1592) & (!sk[111]) & (g1593) & (g1620) & (g44)) + ((!g1592) & (sk[111]) & (!g1593) & (g1620) & (!g44)) + ((!g1592) & (sk[111]) & (!g1593) & (g1620) & (g44)) + ((!g1592) & (sk[111]) & (g1593) & (g1620) & (!g44)) + ((!g1592) & (sk[111]) & (g1593) & (g1620) & (g44)) + ((g1592) & (!sk[111]) & (!g1593) & (!g1620) & (g44)) + ((g1592) & (!sk[111]) & (!g1593) & (g1620) & (!g44)) + ((g1592) & (!sk[111]) & (!g1593) & (g1620) & (g44)) + ((g1592) & (!sk[111]) & (g1593) & (!g1620) & (!g44)) + ((g1592) & (!sk[111]) & (g1593) & (!g1620) & (g44)) + ((g1592) & (!sk[111]) & (g1593) & (g1620) & (!g44)) + ((g1592) & (!sk[111]) & (g1593) & (g1620) & (g44)) + ((g1592) & (sk[111]) & (g1593) & (!g1620) & (g44)) + ((g1592) & (sk[111]) & (g1593) & (g1620) & (g44)));
	assign g1710 = (((!g543) & (!g548) & (!g553) & (g558) & (g820) & (g773)) + ((!g543) & (!g548) & (g553) & (!g558) & (!g820) & (g773)) + ((!g543) & (!g548) & (g553) & (g558) & (!g820) & (g773)) + ((!g543) & (!g548) & (g553) & (g558) & (g820) & (g773)) + ((!g543) & (g548) & (!g553) & (!g558) & (g820) & (!g773)) + ((!g543) & (g548) & (!g553) & (g558) & (g820) & (!g773)) + ((!g543) & (g548) & (!g553) & (g558) & (g820) & (g773)) + ((!g543) & (g548) & (g553) & (!g558) & (!g820) & (g773)) + ((!g543) & (g548) & (g553) & (!g558) & (g820) & (!g773)) + ((!g543) & (g548) & (g553) & (g558) & (!g820) & (g773)) + ((!g543) & (g548) & (g553) & (g558) & (g820) & (!g773)) + ((!g543) & (g548) & (g553) & (g558) & (g820) & (g773)) + ((g543) & (!g548) & (!g553) & (!g558) & (!g820) & (!g773)) + ((g543) & (!g548) & (!g553) & (g558) & (!g820) & (!g773)) + ((g543) & (!g548) & (!g553) & (g558) & (g820) & (g773)) + ((g543) & (!g548) & (g553) & (!g558) & (!g820) & (!g773)) + ((g543) & (!g548) & (g553) & (!g558) & (!g820) & (g773)) + ((g543) & (!g548) & (g553) & (g558) & (!g820) & (!g773)) + ((g543) & (!g548) & (g553) & (g558) & (!g820) & (g773)) + ((g543) & (!g548) & (g553) & (g558) & (g820) & (g773)) + ((g543) & (g548) & (!g553) & (!g558) & (!g820) & (!g773)) + ((g543) & (g548) & (!g553) & (!g558) & (g820) & (!g773)) + ((g543) & (g548) & (!g553) & (g558) & (!g820) & (!g773)) + ((g543) & (g548) & (!g553) & (g558) & (g820) & (!g773)) + ((g543) & (g548) & (!g553) & (g558) & (g820) & (g773)) + ((g543) & (g548) & (g553) & (!g558) & (!g820) & (!g773)) + ((g543) & (g548) & (g553) & (!g558) & (!g820) & (g773)) + ((g543) & (g548) & (g553) & (!g558) & (g820) & (!g773)) + ((g543) & (g548) & (g553) & (g558) & (!g820) & (!g773)) + ((g543) & (g548) & (g553) & (g558) & (!g820) & (g773)) + ((g543) & (g548) & (g553) & (g558) & (g820) & (!g773)) + ((g543) & (g548) & (g553) & (g558) & (g820) & (g773)));
	assign g1711 = (((!g544) & (!g549) & (!g554) & (g559) & (g820) & (g773)) + ((!g544) & (!g549) & (g554) & (!g559) & (!g820) & (g773)) + ((!g544) & (!g549) & (g554) & (g559) & (!g820) & (g773)) + ((!g544) & (!g549) & (g554) & (g559) & (g820) & (g773)) + ((!g544) & (g549) & (!g554) & (!g559) & (g820) & (!g773)) + ((!g544) & (g549) & (!g554) & (g559) & (g820) & (!g773)) + ((!g544) & (g549) & (!g554) & (g559) & (g820) & (g773)) + ((!g544) & (g549) & (g554) & (!g559) & (!g820) & (g773)) + ((!g544) & (g549) & (g554) & (!g559) & (g820) & (!g773)) + ((!g544) & (g549) & (g554) & (g559) & (!g820) & (g773)) + ((!g544) & (g549) & (g554) & (g559) & (g820) & (!g773)) + ((!g544) & (g549) & (g554) & (g559) & (g820) & (g773)) + ((g544) & (!g549) & (!g554) & (!g559) & (!g820) & (!g773)) + ((g544) & (!g549) & (!g554) & (g559) & (!g820) & (!g773)) + ((g544) & (!g549) & (!g554) & (g559) & (g820) & (g773)) + ((g544) & (!g549) & (g554) & (!g559) & (!g820) & (!g773)) + ((g544) & (!g549) & (g554) & (!g559) & (!g820) & (g773)) + ((g544) & (!g549) & (g554) & (g559) & (!g820) & (!g773)) + ((g544) & (!g549) & (g554) & (g559) & (!g820) & (g773)) + ((g544) & (!g549) & (g554) & (g559) & (g820) & (g773)) + ((g544) & (g549) & (!g554) & (!g559) & (!g820) & (!g773)) + ((g544) & (g549) & (!g554) & (!g559) & (g820) & (!g773)) + ((g544) & (g549) & (!g554) & (g559) & (!g820) & (!g773)) + ((g544) & (g549) & (!g554) & (g559) & (g820) & (!g773)) + ((g544) & (g549) & (!g554) & (g559) & (g820) & (g773)) + ((g544) & (g549) & (g554) & (!g559) & (!g820) & (!g773)) + ((g544) & (g549) & (g554) & (!g559) & (!g820) & (g773)) + ((g544) & (g549) & (g554) & (!g559) & (g820) & (!g773)) + ((g544) & (g549) & (g554) & (g559) & (!g820) & (!g773)) + ((g544) & (g549) & (g554) & (g559) & (!g820) & (g773)) + ((g544) & (g549) & (g554) & (g559) & (g820) & (!g773)) + ((g544) & (g549) & (g554) & (g559) & (g820) & (g773)));
	assign g1712 = (((!g545) & (!g550) & (!g555) & (g560) & (g820) & (g773)) + ((!g545) & (!g550) & (g555) & (!g560) & (!g820) & (g773)) + ((!g545) & (!g550) & (g555) & (g560) & (!g820) & (g773)) + ((!g545) & (!g550) & (g555) & (g560) & (g820) & (g773)) + ((!g545) & (g550) & (!g555) & (!g560) & (g820) & (!g773)) + ((!g545) & (g550) & (!g555) & (g560) & (g820) & (!g773)) + ((!g545) & (g550) & (!g555) & (g560) & (g820) & (g773)) + ((!g545) & (g550) & (g555) & (!g560) & (!g820) & (g773)) + ((!g545) & (g550) & (g555) & (!g560) & (g820) & (!g773)) + ((!g545) & (g550) & (g555) & (g560) & (!g820) & (g773)) + ((!g545) & (g550) & (g555) & (g560) & (g820) & (!g773)) + ((!g545) & (g550) & (g555) & (g560) & (g820) & (g773)) + ((g545) & (!g550) & (!g555) & (!g560) & (!g820) & (!g773)) + ((g545) & (!g550) & (!g555) & (g560) & (!g820) & (!g773)) + ((g545) & (!g550) & (!g555) & (g560) & (g820) & (g773)) + ((g545) & (!g550) & (g555) & (!g560) & (!g820) & (!g773)) + ((g545) & (!g550) & (g555) & (!g560) & (!g820) & (g773)) + ((g545) & (!g550) & (g555) & (g560) & (!g820) & (!g773)) + ((g545) & (!g550) & (g555) & (g560) & (!g820) & (g773)) + ((g545) & (!g550) & (g555) & (g560) & (g820) & (g773)) + ((g545) & (g550) & (!g555) & (!g560) & (!g820) & (!g773)) + ((g545) & (g550) & (!g555) & (!g560) & (g820) & (!g773)) + ((g545) & (g550) & (!g555) & (g560) & (!g820) & (!g773)) + ((g545) & (g550) & (!g555) & (g560) & (g820) & (!g773)) + ((g545) & (g550) & (!g555) & (g560) & (g820) & (g773)) + ((g545) & (g550) & (g555) & (!g560) & (!g820) & (!g773)) + ((g545) & (g550) & (g555) & (!g560) & (!g820) & (g773)) + ((g545) & (g550) & (g555) & (!g560) & (g820) & (!g773)) + ((g545) & (g550) & (g555) & (g560) & (!g820) & (!g773)) + ((g545) & (g550) & (g555) & (g560) & (!g820) & (g773)) + ((g545) & (g550) & (g555) & (g560) & (g820) & (!g773)) + ((g545) & (g550) & (g555) & (g560) & (g820) & (g773)));
	assign g1713 = (((!g546) & (!g551) & (!g556) & (g561) & (g820) & (g773)) + ((!g546) & (!g551) & (g556) & (!g561) & (!g820) & (g773)) + ((!g546) & (!g551) & (g556) & (g561) & (!g820) & (g773)) + ((!g546) & (!g551) & (g556) & (g561) & (g820) & (g773)) + ((!g546) & (g551) & (!g556) & (!g561) & (g820) & (!g773)) + ((!g546) & (g551) & (!g556) & (g561) & (g820) & (!g773)) + ((!g546) & (g551) & (!g556) & (g561) & (g820) & (g773)) + ((!g546) & (g551) & (g556) & (!g561) & (!g820) & (g773)) + ((!g546) & (g551) & (g556) & (!g561) & (g820) & (!g773)) + ((!g546) & (g551) & (g556) & (g561) & (!g820) & (g773)) + ((!g546) & (g551) & (g556) & (g561) & (g820) & (!g773)) + ((!g546) & (g551) & (g556) & (g561) & (g820) & (g773)) + ((g546) & (!g551) & (!g556) & (!g561) & (!g820) & (!g773)) + ((g546) & (!g551) & (!g556) & (g561) & (!g820) & (!g773)) + ((g546) & (!g551) & (!g556) & (g561) & (g820) & (g773)) + ((g546) & (!g551) & (g556) & (!g561) & (!g820) & (!g773)) + ((g546) & (!g551) & (g556) & (!g561) & (!g820) & (g773)) + ((g546) & (!g551) & (g556) & (g561) & (!g820) & (!g773)) + ((g546) & (!g551) & (g556) & (g561) & (!g820) & (g773)) + ((g546) & (!g551) & (g556) & (g561) & (g820) & (g773)) + ((g546) & (g551) & (!g556) & (!g561) & (!g820) & (!g773)) + ((g546) & (g551) & (!g556) & (!g561) & (g820) & (!g773)) + ((g546) & (g551) & (!g556) & (g561) & (!g820) & (!g773)) + ((g546) & (g551) & (!g556) & (g561) & (g820) & (!g773)) + ((g546) & (g551) & (!g556) & (g561) & (g820) & (g773)) + ((g546) & (g551) & (g556) & (!g561) & (!g820) & (!g773)) + ((g546) & (g551) & (g556) & (!g561) & (!g820) & (g773)) + ((g546) & (g551) & (g556) & (!g561) & (g820) & (!g773)) + ((g546) & (g551) & (g556) & (g561) & (!g820) & (!g773)) + ((g546) & (g551) & (g556) & (g561) & (!g820) & (g773)) + ((g546) & (g551) & (g556) & (g561) & (g820) & (!g773)) + ((g546) & (g551) & (g556) & (g561) & (g820) & (g773)));
	assign g1714 = (((!g1710) & (!g1711) & (!g1712) & (g1713) & (g677) & (g726)) + ((!g1710) & (!g1711) & (g1712) & (!g1713) & (!g677) & (g726)) + ((!g1710) & (!g1711) & (g1712) & (g1713) & (!g677) & (g726)) + ((!g1710) & (!g1711) & (g1712) & (g1713) & (g677) & (g726)) + ((!g1710) & (g1711) & (!g1712) & (!g1713) & (g677) & (!g726)) + ((!g1710) & (g1711) & (!g1712) & (g1713) & (g677) & (!g726)) + ((!g1710) & (g1711) & (!g1712) & (g1713) & (g677) & (g726)) + ((!g1710) & (g1711) & (g1712) & (!g1713) & (!g677) & (g726)) + ((!g1710) & (g1711) & (g1712) & (!g1713) & (g677) & (!g726)) + ((!g1710) & (g1711) & (g1712) & (g1713) & (!g677) & (g726)) + ((!g1710) & (g1711) & (g1712) & (g1713) & (g677) & (!g726)) + ((!g1710) & (g1711) & (g1712) & (g1713) & (g677) & (g726)) + ((g1710) & (!g1711) & (!g1712) & (!g1713) & (!g677) & (!g726)) + ((g1710) & (!g1711) & (!g1712) & (g1713) & (!g677) & (!g726)) + ((g1710) & (!g1711) & (!g1712) & (g1713) & (g677) & (g726)) + ((g1710) & (!g1711) & (g1712) & (!g1713) & (!g677) & (!g726)) + ((g1710) & (!g1711) & (g1712) & (!g1713) & (!g677) & (g726)) + ((g1710) & (!g1711) & (g1712) & (g1713) & (!g677) & (!g726)) + ((g1710) & (!g1711) & (g1712) & (g1713) & (!g677) & (g726)) + ((g1710) & (!g1711) & (g1712) & (g1713) & (g677) & (g726)) + ((g1710) & (g1711) & (!g1712) & (!g1713) & (!g677) & (!g726)) + ((g1710) & (g1711) & (!g1712) & (!g1713) & (g677) & (!g726)) + ((g1710) & (g1711) & (!g1712) & (g1713) & (!g677) & (!g726)) + ((g1710) & (g1711) & (!g1712) & (g1713) & (g677) & (!g726)) + ((g1710) & (g1711) & (!g1712) & (g1713) & (g677) & (g726)) + ((g1710) & (g1711) & (g1712) & (!g1713) & (!g677) & (!g726)) + ((g1710) & (g1711) & (g1712) & (!g1713) & (!g677) & (g726)) + ((g1710) & (g1711) & (g1712) & (!g1713) & (g677) & (!g726)) + ((g1710) & (g1711) & (g1712) & (g1713) & (!g677) & (!g726)) + ((g1710) & (g1711) & (g1712) & (g1713) & (!g677) & (g726)) + ((g1710) & (g1711) & (g1712) & (g1713) & (g677) & (!g726)) + ((g1710) & (g1711) & (g1712) & (g1713) & (g677) & (g726)));
	assign g1715 = (((!g564) & (!g565) & (!g566) & (g567) & (g677) & (g726)) + ((!g564) & (!g565) & (g566) & (!g567) & (!g677) & (g726)) + ((!g564) & (!g565) & (g566) & (g567) & (!g677) & (g726)) + ((!g564) & (!g565) & (g566) & (g567) & (g677) & (g726)) + ((!g564) & (g565) & (!g566) & (!g567) & (g677) & (!g726)) + ((!g564) & (g565) & (!g566) & (g567) & (g677) & (!g726)) + ((!g564) & (g565) & (!g566) & (g567) & (g677) & (g726)) + ((!g564) & (g565) & (g566) & (!g567) & (!g677) & (g726)) + ((!g564) & (g565) & (g566) & (!g567) & (g677) & (!g726)) + ((!g564) & (g565) & (g566) & (g567) & (!g677) & (g726)) + ((!g564) & (g565) & (g566) & (g567) & (g677) & (!g726)) + ((!g564) & (g565) & (g566) & (g567) & (g677) & (g726)) + ((g564) & (!g565) & (!g566) & (!g567) & (!g677) & (!g726)) + ((g564) & (!g565) & (!g566) & (g567) & (!g677) & (!g726)) + ((g564) & (!g565) & (!g566) & (g567) & (g677) & (g726)) + ((g564) & (!g565) & (g566) & (!g567) & (!g677) & (!g726)) + ((g564) & (!g565) & (g566) & (!g567) & (!g677) & (g726)) + ((g564) & (!g565) & (g566) & (g567) & (!g677) & (!g726)) + ((g564) & (!g565) & (g566) & (g567) & (!g677) & (g726)) + ((g564) & (!g565) & (g566) & (g567) & (g677) & (g726)) + ((g564) & (g565) & (!g566) & (!g567) & (!g677) & (!g726)) + ((g564) & (g565) & (!g566) & (!g567) & (g677) & (!g726)) + ((g564) & (g565) & (!g566) & (g567) & (!g677) & (!g726)) + ((g564) & (g565) & (!g566) & (g567) & (g677) & (!g726)) + ((g564) & (g565) & (!g566) & (g567) & (g677) & (g726)) + ((g564) & (g565) & (g566) & (!g567) & (!g677) & (!g726)) + ((g564) & (g565) & (g566) & (!g567) & (!g677) & (g726)) + ((g564) & (g565) & (g566) & (!g567) & (g677) & (!g726)) + ((g564) & (g565) & (g566) & (g567) & (!g677) & (!g726)) + ((g564) & (g565) & (g566) & (g567) & (!g677) & (g726)) + ((g564) & (g565) & (g566) & (g567) & (g677) & (!g726)) + ((g564) & (g565) & (g566) & (g567) & (g677) & (g726)));
	assign g1716 = (((!g677) & (!g726) & (!sk[118]) & (!g569) & (g570) & (!g571)) + ((!g677) & (!g726) & (!sk[118]) & (!g569) & (g570) & (g571)) + ((!g677) & (!g726) & (!sk[118]) & (g569) & (!g570) & (!g571)) + ((!g677) & (!g726) & (!sk[118]) & (g569) & (!g570) & (g571)) + ((!g677) & (!g726) & (!sk[118]) & (g569) & (g570) & (!g571)) + ((!g677) & (!g726) & (!sk[118]) & (g569) & (g570) & (g571)) + ((!g677) & (g726) & (!sk[118]) & (!g569) & (!g570) & (!g571)) + ((!g677) & (g726) & (!sk[118]) & (!g569) & (!g570) & (g571)) + ((!g677) & (g726) & (!sk[118]) & (!g569) & (g570) & (!g571)) + ((!g677) & (g726) & (!sk[118]) & (!g569) & (g570) & (g571)) + ((!g677) & (g726) & (!sk[118]) & (g569) & (!g570) & (!g571)) + ((!g677) & (g726) & (!sk[118]) & (g569) & (!g570) & (g571)) + ((!g677) & (g726) & (!sk[118]) & (g569) & (g570) & (!g571)) + ((!g677) & (g726) & (!sk[118]) & (g569) & (g570) & (g571)) + ((!g677) & (g726) & (sk[118]) & (!g569) & (!g570) & (g571)) + ((!g677) & (g726) & (sk[118]) & (!g569) & (g570) & (g571)) + ((!g677) & (g726) & (sk[118]) & (g569) & (!g570) & (g571)) + ((!g677) & (g726) & (sk[118]) & (g569) & (g570) & (g571)) + ((g677) & (!g726) & (!sk[118]) & (!g569) & (g570) & (!g571)) + ((g677) & (!g726) & (!sk[118]) & (!g569) & (g570) & (g571)) + ((g677) & (!g726) & (!sk[118]) & (g569) & (!g570) & (!g571)) + ((g677) & (!g726) & (!sk[118]) & (g569) & (!g570) & (g571)) + ((g677) & (!g726) & (!sk[118]) & (g569) & (g570) & (!g571)) + ((g677) & (!g726) & (!sk[118]) & (g569) & (g570) & (g571)) + ((g677) & (!g726) & (sk[118]) & (g569) & (!g570) & (!g571)) + ((g677) & (!g726) & (sk[118]) & (g569) & (!g570) & (g571)) + ((g677) & (!g726) & (sk[118]) & (g569) & (g570) & (!g571)) + ((g677) & (!g726) & (sk[118]) & (g569) & (g570) & (g571)) + ((g677) & (g726) & (!sk[118]) & (!g569) & (!g570) & (!g571)) + ((g677) & (g726) & (!sk[118]) & (!g569) & (!g570) & (g571)) + ((g677) & (g726) & (!sk[118]) & (!g569) & (g570) & (!g571)) + ((g677) & (g726) & (!sk[118]) & (!g569) & (g570) & (g571)) + ((g677) & (g726) & (!sk[118]) & (g569) & (!g570) & (!g571)) + ((g677) & (g726) & (!sk[118]) & (g569) & (!g570) & (g571)) + ((g677) & (g726) & (!sk[118]) & (g569) & (g570) & (!g571)) + ((g677) & (g726) & (!sk[118]) & (g569) & (g570) & (g571)) + ((g677) & (g726) & (sk[118]) & (!g569) & (g570) & (!g571)) + ((g677) & (g726) & (sk[118]) & (!g569) & (g570) & (g571)) + ((g677) & (g726) & (sk[118]) & (g569) & (g570) & (!g571)) + ((g677) & (g726) & (sk[118]) & (g569) & (g570) & (g571)));
	assign g1717 = (((!g573) & (!g574) & (!g575) & (g576) & (g677) & (g726)) + ((!g573) & (!g574) & (g575) & (!g576) & (!g677) & (g726)) + ((!g573) & (!g574) & (g575) & (g576) & (!g677) & (g726)) + ((!g573) & (!g574) & (g575) & (g576) & (g677) & (g726)) + ((!g573) & (g574) & (!g575) & (!g576) & (g677) & (!g726)) + ((!g573) & (g574) & (!g575) & (g576) & (g677) & (!g726)) + ((!g573) & (g574) & (!g575) & (g576) & (g677) & (g726)) + ((!g573) & (g574) & (g575) & (!g576) & (!g677) & (g726)) + ((!g573) & (g574) & (g575) & (!g576) & (g677) & (!g726)) + ((!g573) & (g574) & (g575) & (g576) & (!g677) & (g726)) + ((!g573) & (g574) & (g575) & (g576) & (g677) & (!g726)) + ((!g573) & (g574) & (g575) & (g576) & (g677) & (g726)) + ((g573) & (!g574) & (!g575) & (!g576) & (!g677) & (!g726)) + ((g573) & (!g574) & (!g575) & (g576) & (!g677) & (!g726)) + ((g573) & (!g574) & (!g575) & (g576) & (g677) & (g726)) + ((g573) & (!g574) & (g575) & (!g576) & (!g677) & (!g726)) + ((g573) & (!g574) & (g575) & (!g576) & (!g677) & (g726)) + ((g573) & (!g574) & (g575) & (g576) & (!g677) & (!g726)) + ((g573) & (!g574) & (g575) & (g576) & (!g677) & (g726)) + ((g573) & (!g574) & (g575) & (g576) & (g677) & (g726)) + ((g573) & (g574) & (!g575) & (!g576) & (!g677) & (!g726)) + ((g573) & (g574) & (!g575) & (!g576) & (g677) & (!g726)) + ((g573) & (g574) & (!g575) & (g576) & (!g677) & (!g726)) + ((g573) & (g574) & (!g575) & (g576) & (g677) & (!g726)) + ((g573) & (g574) & (!g575) & (g576) & (g677) & (g726)) + ((g573) & (g574) & (g575) & (!g576) & (!g677) & (!g726)) + ((g573) & (g574) & (g575) & (!g576) & (!g677) & (g726)) + ((g573) & (g574) & (g575) & (!g576) & (g677) & (!g726)) + ((g573) & (g574) & (g575) & (g576) & (!g677) & (!g726)) + ((g573) & (g574) & (g575) & (g576) & (!g677) & (g726)) + ((g573) & (g574) & (g575) & (g576) & (g677) & (!g726)) + ((g573) & (g574) & (g575) & (g576) & (g677) & (g726)));
	assign g1718 = (((!g578) & (!g579) & (!g580) & (g581) & (g677) & (g726)) + ((!g578) & (!g579) & (g580) & (!g581) & (!g677) & (g726)) + ((!g578) & (!g579) & (g580) & (g581) & (!g677) & (g726)) + ((!g578) & (!g579) & (g580) & (g581) & (g677) & (g726)) + ((!g578) & (g579) & (!g580) & (!g581) & (g677) & (!g726)) + ((!g578) & (g579) & (!g580) & (g581) & (g677) & (!g726)) + ((!g578) & (g579) & (!g580) & (g581) & (g677) & (g726)) + ((!g578) & (g579) & (g580) & (!g581) & (!g677) & (g726)) + ((!g578) & (g579) & (g580) & (!g581) & (g677) & (!g726)) + ((!g578) & (g579) & (g580) & (g581) & (!g677) & (g726)) + ((!g578) & (g579) & (g580) & (g581) & (g677) & (!g726)) + ((!g578) & (g579) & (g580) & (g581) & (g677) & (g726)) + ((g578) & (!g579) & (!g580) & (!g581) & (!g677) & (!g726)) + ((g578) & (!g579) & (!g580) & (g581) & (!g677) & (!g726)) + ((g578) & (!g579) & (!g580) & (g581) & (g677) & (g726)) + ((g578) & (!g579) & (g580) & (!g581) & (!g677) & (!g726)) + ((g578) & (!g579) & (g580) & (!g581) & (!g677) & (g726)) + ((g578) & (!g579) & (g580) & (g581) & (!g677) & (!g726)) + ((g578) & (!g579) & (g580) & (g581) & (!g677) & (g726)) + ((g578) & (!g579) & (g580) & (g581) & (g677) & (g726)) + ((g578) & (g579) & (!g580) & (!g581) & (!g677) & (!g726)) + ((g578) & (g579) & (!g580) & (!g581) & (g677) & (!g726)) + ((g578) & (g579) & (!g580) & (g581) & (!g677) & (!g726)) + ((g578) & (g579) & (!g580) & (g581) & (g677) & (!g726)) + ((g578) & (g579) & (!g580) & (g581) & (g677) & (g726)) + ((g578) & (g579) & (g580) & (!g581) & (!g677) & (!g726)) + ((g578) & (g579) & (g580) & (!g581) & (!g677) & (g726)) + ((g578) & (g579) & (g580) & (!g581) & (g677) & (!g726)) + ((g578) & (g579) & (g580) & (g581) & (!g677) & (!g726)) + ((g578) & (g579) & (g580) & (g581) & (!g677) & (g726)) + ((g578) & (g579) & (g580) & (g581) & (g677) & (!g726)) + ((g578) & (g579) & (g580) & (g581) & (g677) & (g726)));
	assign g1719 = (((!g820) & (!g773) & (!g1715) & (g1716) & (!g1717) & (!g1718)) + ((!g820) & (!g773) & (!g1715) & (g1716) & (!g1717) & (g1718)) + ((!g820) & (!g773) & (!g1715) & (g1716) & (g1717) & (!g1718)) + ((!g820) & (!g773) & (!g1715) & (g1716) & (g1717) & (g1718)) + ((!g820) & (!g773) & (g1715) & (g1716) & (!g1717) & (!g1718)) + ((!g820) & (!g773) & (g1715) & (g1716) & (!g1717) & (g1718)) + ((!g820) & (!g773) & (g1715) & (g1716) & (g1717) & (!g1718)) + ((!g820) & (!g773) & (g1715) & (g1716) & (g1717) & (g1718)) + ((!g820) & (g773) & (!g1715) & (!g1716) & (!g1717) & (g1718)) + ((!g820) & (g773) & (!g1715) & (!g1716) & (g1717) & (g1718)) + ((!g820) & (g773) & (!g1715) & (g1716) & (!g1717) & (g1718)) + ((!g820) & (g773) & (!g1715) & (g1716) & (g1717) & (g1718)) + ((!g820) & (g773) & (g1715) & (!g1716) & (!g1717) & (g1718)) + ((!g820) & (g773) & (g1715) & (!g1716) & (g1717) & (g1718)) + ((!g820) & (g773) & (g1715) & (g1716) & (!g1717) & (g1718)) + ((!g820) & (g773) & (g1715) & (g1716) & (g1717) & (g1718)) + ((g820) & (!g773) & (g1715) & (!g1716) & (!g1717) & (!g1718)) + ((g820) & (!g773) & (g1715) & (!g1716) & (!g1717) & (g1718)) + ((g820) & (!g773) & (g1715) & (!g1716) & (g1717) & (!g1718)) + ((g820) & (!g773) & (g1715) & (!g1716) & (g1717) & (g1718)) + ((g820) & (!g773) & (g1715) & (g1716) & (!g1717) & (!g1718)) + ((g820) & (!g773) & (g1715) & (g1716) & (!g1717) & (g1718)) + ((g820) & (!g773) & (g1715) & (g1716) & (g1717) & (!g1718)) + ((g820) & (!g773) & (g1715) & (g1716) & (g1717) & (g1718)) + ((g820) & (g773) & (!g1715) & (!g1716) & (g1717) & (!g1718)) + ((g820) & (g773) & (!g1715) & (!g1716) & (g1717) & (g1718)) + ((g820) & (g773) & (!g1715) & (g1716) & (g1717) & (!g1718)) + ((g820) & (g773) & (!g1715) & (g1716) & (g1717) & (g1718)) + ((g820) & (g773) & (g1715) & (!g1716) & (g1717) & (!g1718)) + ((g820) & (g773) & (g1715) & (!g1716) & (g1717) & (g1718)) + ((g820) & (g773) & (g1715) & (g1716) & (g1717) & (!g1718)) + ((g820) & (g773) & (g1715) & (g1716) & (g1717) & (g1718)));
	assign g1720 = (((!g867) & (!g1714) & (!sk[122]) & (g1719)) + ((!g867) & (!g1714) & (sk[122]) & (g1719)) + ((!g867) & (g1714) & (!sk[122]) & (!g1719)) + ((!g867) & (g1714) & (!sk[122]) & (g1719)) + ((!g867) & (g1714) & (sk[122]) & (g1719)) + ((g867) & (!g1714) & (!sk[122]) & (g1719)) + ((g867) & (g1714) & (!sk[122]) & (!g1719)) + ((g867) & (g1714) & (!sk[122]) & (g1719)) + ((g867) & (g1714) & (sk[122]) & (!g1719)) + ((g867) & (g1714) & (sk[122]) & (g1719)));
	assign g1721 = (((!g132) & (!g1706) & (!g1707) & (!sk[123]) & (g1709) & (!g1720)) + ((!g132) & (!g1706) & (!g1707) & (!sk[123]) & (g1709) & (g1720)) + ((!g132) & (!g1706) & (g1707) & (!sk[123]) & (!g1709) & (!g1720)) + ((!g132) & (!g1706) & (g1707) & (!sk[123]) & (!g1709) & (g1720)) + ((!g132) & (!g1706) & (g1707) & (!sk[123]) & (g1709) & (!g1720)) + ((!g132) & (!g1706) & (g1707) & (!sk[123]) & (g1709) & (g1720)) + ((!g132) & (!g1706) & (g1707) & (sk[123]) & (!g1709) & (g1720)) + ((!g132) & (!g1706) & (g1707) & (sk[123]) & (g1709) & (!g1720)) + ((!g132) & (!g1706) & (g1707) & (sk[123]) & (g1709) & (g1720)) + ((!g132) & (g1706) & (!g1707) & (!sk[123]) & (!g1709) & (!g1720)) + ((!g132) & (g1706) & (!g1707) & (!sk[123]) & (!g1709) & (g1720)) + ((!g132) & (g1706) & (!g1707) & (!sk[123]) & (g1709) & (!g1720)) + ((!g132) & (g1706) & (!g1707) & (!sk[123]) & (g1709) & (g1720)) + ((!g132) & (g1706) & (g1707) & (!sk[123]) & (!g1709) & (!g1720)) + ((!g132) & (g1706) & (g1707) & (!sk[123]) & (!g1709) & (g1720)) + ((!g132) & (g1706) & (g1707) & (!sk[123]) & (g1709) & (!g1720)) + ((!g132) & (g1706) & (g1707) & (!sk[123]) & (g1709) & (g1720)) + ((!g132) & (g1706) & (g1707) & (sk[123]) & (g1709) & (!g1720)) + ((!g132) & (g1706) & (g1707) & (sk[123]) & (g1709) & (g1720)) + ((g132) & (!g1706) & (!g1707) & (!sk[123]) & (g1709) & (!g1720)) + ((g132) & (!g1706) & (!g1707) & (!sk[123]) & (g1709) & (g1720)) + ((g132) & (!g1706) & (g1707) & (!sk[123]) & (!g1709) & (!g1720)) + ((g132) & (!g1706) & (g1707) & (!sk[123]) & (!g1709) & (g1720)) + ((g132) & (!g1706) & (g1707) & (!sk[123]) & (g1709) & (!g1720)) + ((g132) & (!g1706) & (g1707) & (!sk[123]) & (g1709) & (g1720)) + ((g132) & (!g1706) & (g1707) & (sk[123]) & (!g1709) & (g1720)) + ((g132) & (!g1706) & (g1707) & (sk[123]) & (g1709) & (g1720)) + ((g132) & (g1706) & (!g1707) & (!sk[123]) & (!g1709) & (!g1720)) + ((g132) & (g1706) & (!g1707) & (!sk[123]) & (!g1709) & (g1720)) + ((g132) & (g1706) & (!g1707) & (!sk[123]) & (g1709) & (!g1720)) + ((g132) & (g1706) & (!g1707) & (!sk[123]) & (g1709) & (g1720)) + ((g132) & (g1706) & (g1707) & (!sk[123]) & (!g1709) & (!g1720)) + ((g132) & (g1706) & (g1707) & (!sk[123]) & (!g1709) & (g1720)) + ((g132) & (g1706) & (g1707) & (!sk[123]) & (g1709) & (!g1720)) + ((g132) & (g1706) & (g1707) & (!sk[123]) & (g1709) & (g1720)));
	assign g1722 = (((!sk[124]) & (!g1592) & (!g1593) & (!g1632) & (g45)) + ((!sk[124]) & (!g1592) & (!g1593) & (g1632) & (!g45)) + ((!sk[124]) & (!g1592) & (!g1593) & (g1632) & (g45)) + ((!sk[124]) & (!g1592) & (g1593) & (!g1632) & (!g45)) + ((!sk[124]) & (!g1592) & (g1593) & (!g1632) & (g45)) + ((!sk[124]) & (!g1592) & (g1593) & (g1632) & (!g45)) + ((!sk[124]) & (!g1592) & (g1593) & (g1632) & (g45)) + ((!sk[124]) & (g1592) & (!g1593) & (!g1632) & (g45)) + ((!sk[124]) & (g1592) & (!g1593) & (g1632) & (!g45)) + ((!sk[124]) & (g1592) & (!g1593) & (g1632) & (g45)) + ((!sk[124]) & (g1592) & (g1593) & (!g1632) & (!g45)) + ((!sk[124]) & (g1592) & (g1593) & (!g1632) & (g45)) + ((!sk[124]) & (g1592) & (g1593) & (g1632) & (!g45)) + ((!sk[124]) & (g1592) & (g1593) & (g1632) & (g45)) + ((sk[124]) & (!g1592) & (!g1593) & (g1632) & (!g45)) + ((sk[124]) & (!g1592) & (!g1593) & (g1632) & (g45)) + ((sk[124]) & (!g1592) & (g1593) & (g1632) & (!g45)) + ((sk[124]) & (!g1592) & (g1593) & (g1632) & (g45)) + ((sk[124]) & (g1592) & (g1593) & (!g1632) & (g45)) + ((sk[124]) & (g1592) & (g1593) & (g1632) & (g45)));
	assign g1723 = (((!g588) & (!g589) & (!g590) & (g591) & (g820) & (g773)) + ((!g588) & (!g589) & (g590) & (!g591) & (!g820) & (g773)) + ((!g588) & (!g589) & (g590) & (g591) & (!g820) & (g773)) + ((!g588) & (!g589) & (g590) & (g591) & (g820) & (g773)) + ((!g588) & (g589) & (!g590) & (!g591) & (g820) & (!g773)) + ((!g588) & (g589) & (!g590) & (g591) & (g820) & (!g773)) + ((!g588) & (g589) & (!g590) & (g591) & (g820) & (g773)) + ((!g588) & (g589) & (g590) & (!g591) & (!g820) & (g773)) + ((!g588) & (g589) & (g590) & (!g591) & (g820) & (!g773)) + ((!g588) & (g589) & (g590) & (g591) & (!g820) & (g773)) + ((!g588) & (g589) & (g590) & (g591) & (g820) & (!g773)) + ((!g588) & (g589) & (g590) & (g591) & (g820) & (g773)) + ((g588) & (!g589) & (!g590) & (!g591) & (!g820) & (!g773)) + ((g588) & (!g589) & (!g590) & (g591) & (!g820) & (!g773)) + ((g588) & (!g589) & (!g590) & (g591) & (g820) & (g773)) + ((g588) & (!g589) & (g590) & (!g591) & (!g820) & (!g773)) + ((g588) & (!g589) & (g590) & (!g591) & (!g820) & (g773)) + ((g588) & (!g589) & (g590) & (g591) & (!g820) & (!g773)) + ((g588) & (!g589) & (g590) & (g591) & (!g820) & (g773)) + ((g588) & (!g589) & (g590) & (g591) & (g820) & (g773)) + ((g588) & (g589) & (!g590) & (!g591) & (!g820) & (!g773)) + ((g588) & (g589) & (!g590) & (!g591) & (g820) & (!g773)) + ((g588) & (g589) & (!g590) & (g591) & (!g820) & (!g773)) + ((g588) & (g589) & (!g590) & (g591) & (g820) & (!g773)) + ((g588) & (g589) & (!g590) & (g591) & (g820) & (g773)) + ((g588) & (g589) & (g590) & (!g591) & (!g820) & (!g773)) + ((g588) & (g589) & (g590) & (!g591) & (!g820) & (g773)) + ((g588) & (g589) & (g590) & (!g591) & (g820) & (!g773)) + ((g588) & (g589) & (g590) & (g591) & (!g820) & (!g773)) + ((g588) & (g589) & (g590) & (g591) & (!g820) & (g773)) + ((g588) & (g589) & (g590) & (g591) & (g820) & (!g773)) + ((g588) & (g589) & (g590) & (g591) & (g820) & (g773)));
	assign g1724 = (((!g593) & (!g594) & (!g595) & (g596) & (g820) & (g773)) + ((!g593) & (!g594) & (g595) & (!g596) & (!g820) & (g773)) + ((!g593) & (!g594) & (g595) & (g596) & (!g820) & (g773)) + ((!g593) & (!g594) & (g595) & (g596) & (g820) & (g773)) + ((!g593) & (g594) & (!g595) & (!g596) & (g820) & (!g773)) + ((!g593) & (g594) & (!g595) & (g596) & (g820) & (!g773)) + ((!g593) & (g594) & (!g595) & (g596) & (g820) & (g773)) + ((!g593) & (g594) & (g595) & (!g596) & (!g820) & (g773)) + ((!g593) & (g594) & (g595) & (!g596) & (g820) & (!g773)) + ((!g593) & (g594) & (g595) & (g596) & (!g820) & (g773)) + ((!g593) & (g594) & (g595) & (g596) & (g820) & (!g773)) + ((!g593) & (g594) & (g595) & (g596) & (g820) & (g773)) + ((g593) & (!g594) & (!g595) & (!g596) & (!g820) & (!g773)) + ((g593) & (!g594) & (!g595) & (g596) & (!g820) & (!g773)) + ((g593) & (!g594) & (!g595) & (g596) & (g820) & (g773)) + ((g593) & (!g594) & (g595) & (!g596) & (!g820) & (!g773)) + ((g593) & (!g594) & (g595) & (!g596) & (!g820) & (g773)) + ((g593) & (!g594) & (g595) & (g596) & (!g820) & (!g773)) + ((g593) & (!g594) & (g595) & (g596) & (!g820) & (g773)) + ((g593) & (!g594) & (g595) & (g596) & (g820) & (g773)) + ((g593) & (g594) & (!g595) & (!g596) & (!g820) & (!g773)) + ((g593) & (g594) & (!g595) & (!g596) & (g820) & (!g773)) + ((g593) & (g594) & (!g595) & (g596) & (!g820) & (!g773)) + ((g593) & (g594) & (!g595) & (g596) & (g820) & (!g773)) + ((g593) & (g594) & (!g595) & (g596) & (g820) & (g773)) + ((g593) & (g594) & (g595) & (!g596) & (!g820) & (!g773)) + ((g593) & (g594) & (g595) & (!g596) & (!g820) & (g773)) + ((g593) & (g594) & (g595) & (!g596) & (g820) & (!g773)) + ((g593) & (g594) & (g595) & (g596) & (!g820) & (!g773)) + ((g593) & (g594) & (g595) & (g596) & (!g820) & (g773)) + ((g593) & (g594) & (g595) & (g596) & (g820) & (!g773)) + ((g593) & (g594) & (g595) & (g596) & (g820) & (g773)));
	assign g1725 = (((!g598) & (!g599) & (!g600) & (g601) & (g820) & (g773)) + ((!g598) & (!g599) & (g600) & (!g601) & (!g820) & (g773)) + ((!g598) & (!g599) & (g600) & (g601) & (!g820) & (g773)) + ((!g598) & (!g599) & (g600) & (g601) & (g820) & (g773)) + ((!g598) & (g599) & (!g600) & (!g601) & (g820) & (!g773)) + ((!g598) & (g599) & (!g600) & (g601) & (g820) & (!g773)) + ((!g598) & (g599) & (!g600) & (g601) & (g820) & (g773)) + ((!g598) & (g599) & (g600) & (!g601) & (!g820) & (g773)) + ((!g598) & (g599) & (g600) & (!g601) & (g820) & (!g773)) + ((!g598) & (g599) & (g600) & (g601) & (!g820) & (g773)) + ((!g598) & (g599) & (g600) & (g601) & (g820) & (!g773)) + ((!g598) & (g599) & (g600) & (g601) & (g820) & (g773)) + ((g598) & (!g599) & (!g600) & (!g601) & (!g820) & (!g773)) + ((g598) & (!g599) & (!g600) & (g601) & (!g820) & (!g773)) + ((g598) & (!g599) & (!g600) & (g601) & (g820) & (g773)) + ((g598) & (!g599) & (g600) & (!g601) & (!g820) & (!g773)) + ((g598) & (!g599) & (g600) & (!g601) & (!g820) & (g773)) + ((g598) & (!g599) & (g600) & (g601) & (!g820) & (!g773)) + ((g598) & (!g599) & (g600) & (g601) & (!g820) & (g773)) + ((g598) & (!g599) & (g600) & (g601) & (g820) & (g773)) + ((g598) & (g599) & (!g600) & (!g601) & (!g820) & (!g773)) + ((g598) & (g599) & (!g600) & (!g601) & (g820) & (!g773)) + ((g598) & (g599) & (!g600) & (g601) & (!g820) & (!g773)) + ((g598) & (g599) & (!g600) & (g601) & (g820) & (!g773)) + ((g598) & (g599) & (!g600) & (g601) & (g820) & (g773)) + ((g598) & (g599) & (g600) & (!g601) & (!g820) & (!g773)) + ((g598) & (g599) & (g600) & (!g601) & (!g820) & (g773)) + ((g598) & (g599) & (g600) & (!g601) & (g820) & (!g773)) + ((g598) & (g599) & (g600) & (g601) & (!g820) & (!g773)) + ((g598) & (g599) & (g600) & (g601) & (!g820) & (g773)) + ((g598) & (g599) & (g600) & (g601) & (g820) & (!g773)) + ((g598) & (g599) & (g600) & (g601) & (g820) & (g773)));
	assign g1726 = (((!g603) & (!g604) & (!g605) & (g606) & (g820) & (g773)) + ((!g603) & (!g604) & (g605) & (!g606) & (!g820) & (g773)) + ((!g603) & (!g604) & (g605) & (g606) & (!g820) & (g773)) + ((!g603) & (!g604) & (g605) & (g606) & (g820) & (g773)) + ((!g603) & (g604) & (!g605) & (!g606) & (g820) & (!g773)) + ((!g603) & (g604) & (!g605) & (g606) & (g820) & (!g773)) + ((!g603) & (g604) & (!g605) & (g606) & (g820) & (g773)) + ((!g603) & (g604) & (g605) & (!g606) & (!g820) & (g773)) + ((!g603) & (g604) & (g605) & (!g606) & (g820) & (!g773)) + ((!g603) & (g604) & (g605) & (g606) & (!g820) & (g773)) + ((!g603) & (g604) & (g605) & (g606) & (g820) & (!g773)) + ((!g603) & (g604) & (g605) & (g606) & (g820) & (g773)) + ((g603) & (!g604) & (!g605) & (!g606) & (!g820) & (!g773)) + ((g603) & (!g604) & (!g605) & (g606) & (!g820) & (!g773)) + ((g603) & (!g604) & (!g605) & (g606) & (g820) & (g773)) + ((g603) & (!g604) & (g605) & (!g606) & (!g820) & (!g773)) + ((g603) & (!g604) & (g605) & (!g606) & (!g820) & (g773)) + ((g603) & (!g604) & (g605) & (g606) & (!g820) & (!g773)) + ((g603) & (!g604) & (g605) & (g606) & (!g820) & (g773)) + ((g603) & (!g604) & (g605) & (g606) & (g820) & (g773)) + ((g603) & (g604) & (!g605) & (!g606) & (!g820) & (!g773)) + ((g603) & (g604) & (!g605) & (!g606) & (g820) & (!g773)) + ((g603) & (g604) & (!g605) & (g606) & (!g820) & (!g773)) + ((g603) & (g604) & (!g605) & (g606) & (g820) & (!g773)) + ((g603) & (g604) & (!g605) & (g606) & (g820) & (g773)) + ((g603) & (g604) & (g605) & (!g606) & (!g820) & (!g773)) + ((g603) & (g604) & (g605) & (!g606) & (!g820) & (g773)) + ((g603) & (g604) & (g605) & (!g606) & (g820) & (!g773)) + ((g603) & (g604) & (g605) & (g606) & (!g820) & (!g773)) + ((g603) & (g604) & (g605) & (g606) & (!g820) & (g773)) + ((g603) & (g604) & (g605) & (g606) & (g820) & (!g773)) + ((g603) & (g604) & (g605) & (g606) & (g820) & (g773)));
	assign g1727 = (((!g1723) & (!g1724) & (!g1725) & (g1726) & (g677) & (g726)) + ((!g1723) & (!g1724) & (g1725) & (!g1726) & (!g677) & (g726)) + ((!g1723) & (!g1724) & (g1725) & (g1726) & (!g677) & (g726)) + ((!g1723) & (!g1724) & (g1725) & (g1726) & (g677) & (g726)) + ((!g1723) & (g1724) & (!g1725) & (!g1726) & (g677) & (!g726)) + ((!g1723) & (g1724) & (!g1725) & (g1726) & (g677) & (!g726)) + ((!g1723) & (g1724) & (!g1725) & (g1726) & (g677) & (g726)) + ((!g1723) & (g1724) & (g1725) & (!g1726) & (!g677) & (g726)) + ((!g1723) & (g1724) & (g1725) & (!g1726) & (g677) & (!g726)) + ((!g1723) & (g1724) & (g1725) & (g1726) & (!g677) & (g726)) + ((!g1723) & (g1724) & (g1725) & (g1726) & (g677) & (!g726)) + ((!g1723) & (g1724) & (g1725) & (g1726) & (g677) & (g726)) + ((g1723) & (!g1724) & (!g1725) & (!g1726) & (!g677) & (!g726)) + ((g1723) & (!g1724) & (!g1725) & (g1726) & (!g677) & (!g726)) + ((g1723) & (!g1724) & (!g1725) & (g1726) & (g677) & (g726)) + ((g1723) & (!g1724) & (g1725) & (!g1726) & (!g677) & (!g726)) + ((g1723) & (!g1724) & (g1725) & (!g1726) & (!g677) & (g726)) + ((g1723) & (!g1724) & (g1725) & (g1726) & (!g677) & (!g726)) + ((g1723) & (!g1724) & (g1725) & (g1726) & (!g677) & (g726)) + ((g1723) & (!g1724) & (g1725) & (g1726) & (g677) & (g726)) + ((g1723) & (g1724) & (!g1725) & (!g1726) & (!g677) & (!g726)) + ((g1723) & (g1724) & (!g1725) & (!g1726) & (g677) & (!g726)) + ((g1723) & (g1724) & (!g1725) & (g1726) & (!g677) & (!g726)) + ((g1723) & (g1724) & (!g1725) & (g1726) & (g677) & (!g726)) + ((g1723) & (g1724) & (!g1725) & (g1726) & (g677) & (g726)) + ((g1723) & (g1724) & (g1725) & (!g1726) & (!g677) & (!g726)) + ((g1723) & (g1724) & (g1725) & (!g1726) & (!g677) & (g726)) + ((g1723) & (g1724) & (g1725) & (!g1726) & (g677) & (!g726)) + ((g1723) & (g1724) & (g1725) & (g1726) & (!g677) & (!g726)) + ((g1723) & (g1724) & (g1725) & (g1726) & (!g677) & (g726)) + ((g1723) & (g1724) & (g1725) & (g1726) & (g677) & (!g726)) + ((g1723) & (g1724) & (g1725) & (g1726) & (g677) & (g726)));
	assign g1728 = (((!g609) & (!g610) & (!g611) & (g612) & (g677) & (g726)) + ((!g609) & (!g610) & (g611) & (!g612) & (!g677) & (g726)) + ((!g609) & (!g610) & (g611) & (g612) & (!g677) & (g726)) + ((!g609) & (!g610) & (g611) & (g612) & (g677) & (g726)) + ((!g609) & (g610) & (!g611) & (!g612) & (g677) & (!g726)) + ((!g609) & (g610) & (!g611) & (g612) & (g677) & (!g726)) + ((!g609) & (g610) & (!g611) & (g612) & (g677) & (g726)) + ((!g609) & (g610) & (g611) & (!g612) & (!g677) & (g726)) + ((!g609) & (g610) & (g611) & (!g612) & (g677) & (!g726)) + ((!g609) & (g610) & (g611) & (g612) & (!g677) & (g726)) + ((!g609) & (g610) & (g611) & (g612) & (g677) & (!g726)) + ((!g609) & (g610) & (g611) & (g612) & (g677) & (g726)) + ((g609) & (!g610) & (!g611) & (!g612) & (!g677) & (!g726)) + ((g609) & (!g610) & (!g611) & (g612) & (!g677) & (!g726)) + ((g609) & (!g610) & (!g611) & (g612) & (g677) & (g726)) + ((g609) & (!g610) & (g611) & (!g612) & (!g677) & (!g726)) + ((g609) & (!g610) & (g611) & (!g612) & (!g677) & (g726)) + ((g609) & (!g610) & (g611) & (g612) & (!g677) & (!g726)) + ((g609) & (!g610) & (g611) & (g612) & (!g677) & (g726)) + ((g609) & (!g610) & (g611) & (g612) & (g677) & (g726)) + ((g609) & (g610) & (!g611) & (!g612) & (!g677) & (!g726)) + ((g609) & (g610) & (!g611) & (!g612) & (g677) & (!g726)) + ((g609) & (g610) & (!g611) & (g612) & (!g677) & (!g726)) + ((g609) & (g610) & (!g611) & (g612) & (g677) & (!g726)) + ((g609) & (g610) & (!g611) & (g612) & (g677) & (g726)) + ((g609) & (g610) & (g611) & (!g612) & (!g677) & (!g726)) + ((g609) & (g610) & (g611) & (!g612) & (!g677) & (g726)) + ((g609) & (g610) & (g611) & (!g612) & (g677) & (!g726)) + ((g609) & (g610) & (g611) & (g612) & (!g677) & (!g726)) + ((g609) & (g610) & (g611) & (g612) & (!g677) & (g726)) + ((g609) & (g610) & (g611) & (g612) & (g677) & (!g726)) + ((g609) & (g610) & (g611) & (g612) & (g677) & (g726)));
	assign g1729 = (((!g677) & (!g726) & (!g614) & (g615) & (!sk[3]) & (!g616)) + ((!g677) & (!g726) & (!g614) & (g615) & (!sk[3]) & (g616)) + ((!g677) & (!g726) & (g614) & (!g615) & (!sk[3]) & (!g616)) + ((!g677) & (!g726) & (g614) & (!g615) & (!sk[3]) & (g616)) + ((!g677) & (!g726) & (g614) & (g615) & (!sk[3]) & (!g616)) + ((!g677) & (!g726) & (g614) & (g615) & (!sk[3]) & (g616)) + ((!g677) & (g726) & (!g614) & (!g615) & (!sk[3]) & (!g616)) + ((!g677) & (g726) & (!g614) & (!g615) & (!sk[3]) & (g616)) + ((!g677) & (g726) & (!g614) & (!g615) & (sk[3]) & (g616)) + ((!g677) & (g726) & (!g614) & (g615) & (!sk[3]) & (!g616)) + ((!g677) & (g726) & (!g614) & (g615) & (!sk[3]) & (g616)) + ((!g677) & (g726) & (!g614) & (g615) & (sk[3]) & (g616)) + ((!g677) & (g726) & (g614) & (!g615) & (!sk[3]) & (!g616)) + ((!g677) & (g726) & (g614) & (!g615) & (!sk[3]) & (g616)) + ((!g677) & (g726) & (g614) & (!g615) & (sk[3]) & (g616)) + ((!g677) & (g726) & (g614) & (g615) & (!sk[3]) & (!g616)) + ((!g677) & (g726) & (g614) & (g615) & (!sk[3]) & (g616)) + ((!g677) & (g726) & (g614) & (g615) & (sk[3]) & (g616)) + ((g677) & (!g726) & (!g614) & (g615) & (!sk[3]) & (!g616)) + ((g677) & (!g726) & (!g614) & (g615) & (!sk[3]) & (g616)) + ((g677) & (!g726) & (g614) & (!g615) & (!sk[3]) & (!g616)) + ((g677) & (!g726) & (g614) & (!g615) & (!sk[3]) & (g616)) + ((g677) & (!g726) & (g614) & (!g615) & (sk[3]) & (!g616)) + ((g677) & (!g726) & (g614) & (!g615) & (sk[3]) & (g616)) + ((g677) & (!g726) & (g614) & (g615) & (!sk[3]) & (!g616)) + ((g677) & (!g726) & (g614) & (g615) & (!sk[3]) & (g616)) + ((g677) & (!g726) & (g614) & (g615) & (sk[3]) & (!g616)) + ((g677) & (!g726) & (g614) & (g615) & (sk[3]) & (g616)) + ((g677) & (g726) & (!g614) & (!g615) & (!sk[3]) & (!g616)) + ((g677) & (g726) & (!g614) & (!g615) & (!sk[3]) & (g616)) + ((g677) & (g726) & (!g614) & (g615) & (!sk[3]) & (!g616)) + ((g677) & (g726) & (!g614) & (g615) & (!sk[3]) & (g616)) + ((g677) & (g726) & (!g614) & (g615) & (sk[3]) & (!g616)) + ((g677) & (g726) & (!g614) & (g615) & (sk[3]) & (g616)) + ((g677) & (g726) & (g614) & (!g615) & (!sk[3]) & (!g616)) + ((g677) & (g726) & (g614) & (!g615) & (!sk[3]) & (g616)) + ((g677) & (g726) & (g614) & (g615) & (!sk[3]) & (!g616)) + ((g677) & (g726) & (g614) & (g615) & (!sk[3]) & (g616)) + ((g677) & (g726) & (g614) & (g615) & (sk[3]) & (!g616)) + ((g677) & (g726) & (g614) & (g615) & (sk[3]) & (g616)));
	assign g1730 = (((!g618) & (!g619) & (!g620) & (g621) & (g677) & (g726)) + ((!g618) & (!g619) & (g620) & (!g621) & (!g677) & (g726)) + ((!g618) & (!g619) & (g620) & (g621) & (!g677) & (g726)) + ((!g618) & (!g619) & (g620) & (g621) & (g677) & (g726)) + ((!g618) & (g619) & (!g620) & (!g621) & (g677) & (!g726)) + ((!g618) & (g619) & (!g620) & (g621) & (g677) & (!g726)) + ((!g618) & (g619) & (!g620) & (g621) & (g677) & (g726)) + ((!g618) & (g619) & (g620) & (!g621) & (!g677) & (g726)) + ((!g618) & (g619) & (g620) & (!g621) & (g677) & (!g726)) + ((!g618) & (g619) & (g620) & (g621) & (!g677) & (g726)) + ((!g618) & (g619) & (g620) & (g621) & (g677) & (!g726)) + ((!g618) & (g619) & (g620) & (g621) & (g677) & (g726)) + ((g618) & (!g619) & (!g620) & (!g621) & (!g677) & (!g726)) + ((g618) & (!g619) & (!g620) & (g621) & (!g677) & (!g726)) + ((g618) & (!g619) & (!g620) & (g621) & (g677) & (g726)) + ((g618) & (!g619) & (g620) & (!g621) & (!g677) & (!g726)) + ((g618) & (!g619) & (g620) & (!g621) & (!g677) & (g726)) + ((g618) & (!g619) & (g620) & (g621) & (!g677) & (!g726)) + ((g618) & (!g619) & (g620) & (g621) & (!g677) & (g726)) + ((g618) & (!g619) & (g620) & (g621) & (g677) & (g726)) + ((g618) & (g619) & (!g620) & (!g621) & (!g677) & (!g726)) + ((g618) & (g619) & (!g620) & (!g621) & (g677) & (!g726)) + ((g618) & (g619) & (!g620) & (g621) & (!g677) & (!g726)) + ((g618) & (g619) & (!g620) & (g621) & (g677) & (!g726)) + ((g618) & (g619) & (!g620) & (g621) & (g677) & (g726)) + ((g618) & (g619) & (g620) & (!g621) & (!g677) & (!g726)) + ((g618) & (g619) & (g620) & (!g621) & (!g677) & (g726)) + ((g618) & (g619) & (g620) & (!g621) & (g677) & (!g726)) + ((g618) & (g619) & (g620) & (g621) & (!g677) & (!g726)) + ((g618) & (g619) & (g620) & (g621) & (!g677) & (g726)) + ((g618) & (g619) & (g620) & (g621) & (g677) & (!g726)) + ((g618) & (g619) & (g620) & (g621) & (g677) & (g726)));
	assign g1731 = (((!g623) & (!g624) & (!g625) & (g626) & (g677) & (g726)) + ((!g623) & (!g624) & (g625) & (!g626) & (!g677) & (g726)) + ((!g623) & (!g624) & (g625) & (g626) & (!g677) & (g726)) + ((!g623) & (!g624) & (g625) & (g626) & (g677) & (g726)) + ((!g623) & (g624) & (!g625) & (!g626) & (g677) & (!g726)) + ((!g623) & (g624) & (!g625) & (g626) & (g677) & (!g726)) + ((!g623) & (g624) & (!g625) & (g626) & (g677) & (g726)) + ((!g623) & (g624) & (g625) & (!g626) & (!g677) & (g726)) + ((!g623) & (g624) & (g625) & (!g626) & (g677) & (!g726)) + ((!g623) & (g624) & (g625) & (g626) & (!g677) & (g726)) + ((!g623) & (g624) & (g625) & (g626) & (g677) & (!g726)) + ((!g623) & (g624) & (g625) & (g626) & (g677) & (g726)) + ((g623) & (!g624) & (!g625) & (!g626) & (!g677) & (!g726)) + ((g623) & (!g624) & (!g625) & (g626) & (!g677) & (!g726)) + ((g623) & (!g624) & (!g625) & (g626) & (g677) & (g726)) + ((g623) & (!g624) & (g625) & (!g626) & (!g677) & (!g726)) + ((g623) & (!g624) & (g625) & (!g626) & (!g677) & (g726)) + ((g623) & (!g624) & (g625) & (g626) & (!g677) & (!g726)) + ((g623) & (!g624) & (g625) & (g626) & (!g677) & (g726)) + ((g623) & (!g624) & (g625) & (g626) & (g677) & (g726)) + ((g623) & (g624) & (!g625) & (!g626) & (!g677) & (!g726)) + ((g623) & (g624) & (!g625) & (!g626) & (g677) & (!g726)) + ((g623) & (g624) & (!g625) & (g626) & (!g677) & (!g726)) + ((g623) & (g624) & (!g625) & (g626) & (g677) & (!g726)) + ((g623) & (g624) & (!g625) & (g626) & (g677) & (g726)) + ((g623) & (g624) & (g625) & (!g626) & (!g677) & (!g726)) + ((g623) & (g624) & (g625) & (!g626) & (!g677) & (g726)) + ((g623) & (g624) & (g625) & (!g626) & (g677) & (!g726)) + ((g623) & (g624) & (g625) & (g626) & (!g677) & (!g726)) + ((g623) & (g624) & (g625) & (g626) & (!g677) & (g726)) + ((g623) & (g624) & (g625) & (g626) & (g677) & (!g726)) + ((g623) & (g624) & (g625) & (g626) & (g677) & (g726)));
	assign g1732 = (((!g820) & (!g773) & (!g1728) & (g1729) & (!g1730) & (!g1731)) + ((!g820) & (!g773) & (!g1728) & (g1729) & (!g1730) & (g1731)) + ((!g820) & (!g773) & (!g1728) & (g1729) & (g1730) & (!g1731)) + ((!g820) & (!g773) & (!g1728) & (g1729) & (g1730) & (g1731)) + ((!g820) & (!g773) & (g1728) & (g1729) & (!g1730) & (!g1731)) + ((!g820) & (!g773) & (g1728) & (g1729) & (!g1730) & (g1731)) + ((!g820) & (!g773) & (g1728) & (g1729) & (g1730) & (!g1731)) + ((!g820) & (!g773) & (g1728) & (g1729) & (g1730) & (g1731)) + ((!g820) & (g773) & (!g1728) & (!g1729) & (!g1730) & (g1731)) + ((!g820) & (g773) & (!g1728) & (!g1729) & (g1730) & (g1731)) + ((!g820) & (g773) & (!g1728) & (g1729) & (!g1730) & (g1731)) + ((!g820) & (g773) & (!g1728) & (g1729) & (g1730) & (g1731)) + ((!g820) & (g773) & (g1728) & (!g1729) & (!g1730) & (g1731)) + ((!g820) & (g773) & (g1728) & (!g1729) & (g1730) & (g1731)) + ((!g820) & (g773) & (g1728) & (g1729) & (!g1730) & (g1731)) + ((!g820) & (g773) & (g1728) & (g1729) & (g1730) & (g1731)) + ((g820) & (!g773) & (g1728) & (!g1729) & (!g1730) & (!g1731)) + ((g820) & (!g773) & (g1728) & (!g1729) & (!g1730) & (g1731)) + ((g820) & (!g773) & (g1728) & (!g1729) & (g1730) & (!g1731)) + ((g820) & (!g773) & (g1728) & (!g1729) & (g1730) & (g1731)) + ((g820) & (!g773) & (g1728) & (g1729) & (!g1730) & (!g1731)) + ((g820) & (!g773) & (g1728) & (g1729) & (!g1730) & (g1731)) + ((g820) & (!g773) & (g1728) & (g1729) & (g1730) & (!g1731)) + ((g820) & (!g773) & (g1728) & (g1729) & (g1730) & (g1731)) + ((g820) & (g773) & (!g1728) & (!g1729) & (g1730) & (!g1731)) + ((g820) & (g773) & (!g1728) & (!g1729) & (g1730) & (g1731)) + ((g820) & (g773) & (!g1728) & (g1729) & (g1730) & (!g1731)) + ((g820) & (g773) & (!g1728) & (g1729) & (g1730) & (g1731)) + ((g820) & (g773) & (g1728) & (!g1729) & (g1730) & (!g1731)) + ((g820) & (g773) & (g1728) & (!g1729) & (g1730) & (g1731)) + ((g820) & (g773) & (g1728) & (g1729) & (g1730) & (!g1731)) + ((g820) & (g773) & (g1728) & (g1729) & (g1730) & (g1731)));
	assign g1733 = (((!g867) & (!g1727) & (!sk[7]) & (g1732)) + ((!g867) & (!g1727) & (sk[7]) & (g1732)) + ((!g867) & (g1727) & (!sk[7]) & (!g1732)) + ((!g867) & (g1727) & (!sk[7]) & (g1732)) + ((!g867) & (g1727) & (sk[7]) & (g1732)) + ((g867) & (!g1727) & (!sk[7]) & (g1732)) + ((g867) & (g1727) & (!sk[7]) & (!g1732)) + ((g867) & (g1727) & (!sk[7]) & (g1732)) + ((g867) & (g1727) & (sk[7]) & (!g1732)) + ((g867) & (g1727) & (sk[7]) & (g1732)));
	assign g1734 = (((!g132) & (!g1706) & (!sk[8]) & (!g1707) & (g1722) & (!g1733)) + ((!g132) & (!g1706) & (!sk[8]) & (!g1707) & (g1722) & (g1733)) + ((!g132) & (!g1706) & (!sk[8]) & (g1707) & (!g1722) & (!g1733)) + ((!g132) & (!g1706) & (!sk[8]) & (g1707) & (!g1722) & (g1733)) + ((!g132) & (!g1706) & (!sk[8]) & (g1707) & (g1722) & (!g1733)) + ((!g132) & (!g1706) & (!sk[8]) & (g1707) & (g1722) & (g1733)) + ((!g132) & (!g1706) & (sk[8]) & (g1707) & (!g1722) & (g1733)) + ((!g132) & (!g1706) & (sk[8]) & (g1707) & (g1722) & (!g1733)) + ((!g132) & (!g1706) & (sk[8]) & (g1707) & (g1722) & (g1733)) + ((!g132) & (g1706) & (!sk[8]) & (!g1707) & (!g1722) & (!g1733)) + ((!g132) & (g1706) & (!sk[8]) & (!g1707) & (!g1722) & (g1733)) + ((!g132) & (g1706) & (!sk[8]) & (!g1707) & (g1722) & (!g1733)) + ((!g132) & (g1706) & (!sk[8]) & (!g1707) & (g1722) & (g1733)) + ((!g132) & (g1706) & (!sk[8]) & (g1707) & (!g1722) & (!g1733)) + ((!g132) & (g1706) & (!sk[8]) & (g1707) & (!g1722) & (g1733)) + ((!g132) & (g1706) & (!sk[8]) & (g1707) & (g1722) & (!g1733)) + ((!g132) & (g1706) & (!sk[8]) & (g1707) & (g1722) & (g1733)) + ((!g132) & (g1706) & (sk[8]) & (g1707) & (g1722) & (!g1733)) + ((!g132) & (g1706) & (sk[8]) & (g1707) & (g1722) & (g1733)) + ((g132) & (!g1706) & (!sk[8]) & (!g1707) & (g1722) & (!g1733)) + ((g132) & (!g1706) & (!sk[8]) & (!g1707) & (g1722) & (g1733)) + ((g132) & (!g1706) & (!sk[8]) & (g1707) & (!g1722) & (!g1733)) + ((g132) & (!g1706) & (!sk[8]) & (g1707) & (!g1722) & (g1733)) + ((g132) & (!g1706) & (!sk[8]) & (g1707) & (g1722) & (!g1733)) + ((g132) & (!g1706) & (!sk[8]) & (g1707) & (g1722) & (g1733)) + ((g132) & (!g1706) & (sk[8]) & (g1707) & (!g1722) & (g1733)) + ((g132) & (!g1706) & (sk[8]) & (g1707) & (g1722) & (g1733)) + ((g132) & (g1706) & (!sk[8]) & (!g1707) & (!g1722) & (!g1733)) + ((g132) & (g1706) & (!sk[8]) & (!g1707) & (!g1722) & (g1733)) + ((g132) & (g1706) & (!sk[8]) & (!g1707) & (g1722) & (!g1733)) + ((g132) & (g1706) & (!sk[8]) & (!g1707) & (g1722) & (g1733)) + ((g132) & (g1706) & (!sk[8]) & (g1707) & (!g1722) & (!g1733)) + ((g132) & (g1706) & (!sk[8]) & (g1707) & (!g1722) & (g1733)) + ((g132) & (g1706) & (!sk[8]) & (g1707) & (g1722) & (!g1733)) + ((g132) & (g1706) & (!sk[8]) & (g1707) & (g1722) & (g1733)));
	assign g1735 = (((!g1592) & (!sk[9]) & (!g1593) & (!g1644) & (g46)) + ((!g1592) & (!sk[9]) & (!g1593) & (g1644) & (!g46)) + ((!g1592) & (!sk[9]) & (!g1593) & (g1644) & (g46)) + ((!g1592) & (!sk[9]) & (g1593) & (!g1644) & (!g46)) + ((!g1592) & (!sk[9]) & (g1593) & (!g1644) & (g46)) + ((!g1592) & (!sk[9]) & (g1593) & (g1644) & (!g46)) + ((!g1592) & (!sk[9]) & (g1593) & (g1644) & (g46)) + ((!g1592) & (sk[9]) & (!g1593) & (g1644) & (!g46)) + ((!g1592) & (sk[9]) & (!g1593) & (g1644) & (g46)) + ((!g1592) & (sk[9]) & (g1593) & (g1644) & (!g46)) + ((!g1592) & (sk[9]) & (g1593) & (g1644) & (g46)) + ((g1592) & (!sk[9]) & (!g1593) & (!g1644) & (g46)) + ((g1592) & (!sk[9]) & (!g1593) & (g1644) & (!g46)) + ((g1592) & (!sk[9]) & (!g1593) & (g1644) & (g46)) + ((g1592) & (!sk[9]) & (g1593) & (!g1644) & (!g46)) + ((g1592) & (!sk[9]) & (g1593) & (!g1644) & (g46)) + ((g1592) & (!sk[9]) & (g1593) & (g1644) & (!g46)) + ((g1592) & (!sk[9]) & (g1593) & (g1644) & (g46)) + ((g1592) & (sk[9]) & (g1593) & (!g1644) & (g46)) + ((g1592) & (sk[9]) & (g1593) & (g1644) & (g46)));
	assign g1736 = (((!g631) & (!g632) & (!g633) & (g634) & (g820) & (g773)) + ((!g631) & (!g632) & (g633) & (!g634) & (!g820) & (g773)) + ((!g631) & (!g632) & (g633) & (g634) & (!g820) & (g773)) + ((!g631) & (!g632) & (g633) & (g634) & (g820) & (g773)) + ((!g631) & (g632) & (!g633) & (!g634) & (g820) & (!g773)) + ((!g631) & (g632) & (!g633) & (g634) & (g820) & (!g773)) + ((!g631) & (g632) & (!g633) & (g634) & (g820) & (g773)) + ((!g631) & (g632) & (g633) & (!g634) & (!g820) & (g773)) + ((!g631) & (g632) & (g633) & (!g634) & (g820) & (!g773)) + ((!g631) & (g632) & (g633) & (g634) & (!g820) & (g773)) + ((!g631) & (g632) & (g633) & (g634) & (g820) & (!g773)) + ((!g631) & (g632) & (g633) & (g634) & (g820) & (g773)) + ((g631) & (!g632) & (!g633) & (!g634) & (!g820) & (!g773)) + ((g631) & (!g632) & (!g633) & (g634) & (!g820) & (!g773)) + ((g631) & (!g632) & (!g633) & (g634) & (g820) & (g773)) + ((g631) & (!g632) & (g633) & (!g634) & (!g820) & (!g773)) + ((g631) & (!g632) & (g633) & (!g634) & (!g820) & (g773)) + ((g631) & (!g632) & (g633) & (g634) & (!g820) & (!g773)) + ((g631) & (!g632) & (g633) & (g634) & (!g820) & (g773)) + ((g631) & (!g632) & (g633) & (g634) & (g820) & (g773)) + ((g631) & (g632) & (!g633) & (!g634) & (!g820) & (!g773)) + ((g631) & (g632) & (!g633) & (!g634) & (g820) & (!g773)) + ((g631) & (g632) & (!g633) & (g634) & (!g820) & (!g773)) + ((g631) & (g632) & (!g633) & (g634) & (g820) & (!g773)) + ((g631) & (g632) & (!g633) & (g634) & (g820) & (g773)) + ((g631) & (g632) & (g633) & (!g634) & (!g820) & (!g773)) + ((g631) & (g632) & (g633) & (!g634) & (!g820) & (g773)) + ((g631) & (g632) & (g633) & (!g634) & (g820) & (!g773)) + ((g631) & (g632) & (g633) & (g634) & (!g820) & (!g773)) + ((g631) & (g632) & (g633) & (g634) & (!g820) & (g773)) + ((g631) & (g632) & (g633) & (g634) & (g820) & (!g773)) + ((g631) & (g632) & (g633) & (g634) & (g820) & (g773)));
	assign g1737 = (((!g636) & (!g637) & (!g638) & (g639) & (g820) & (g773)) + ((!g636) & (!g637) & (g638) & (!g639) & (!g820) & (g773)) + ((!g636) & (!g637) & (g638) & (g639) & (!g820) & (g773)) + ((!g636) & (!g637) & (g638) & (g639) & (g820) & (g773)) + ((!g636) & (g637) & (!g638) & (!g639) & (g820) & (!g773)) + ((!g636) & (g637) & (!g638) & (g639) & (g820) & (!g773)) + ((!g636) & (g637) & (!g638) & (g639) & (g820) & (g773)) + ((!g636) & (g637) & (g638) & (!g639) & (!g820) & (g773)) + ((!g636) & (g637) & (g638) & (!g639) & (g820) & (!g773)) + ((!g636) & (g637) & (g638) & (g639) & (!g820) & (g773)) + ((!g636) & (g637) & (g638) & (g639) & (g820) & (!g773)) + ((!g636) & (g637) & (g638) & (g639) & (g820) & (g773)) + ((g636) & (!g637) & (!g638) & (!g639) & (!g820) & (!g773)) + ((g636) & (!g637) & (!g638) & (g639) & (!g820) & (!g773)) + ((g636) & (!g637) & (!g638) & (g639) & (g820) & (g773)) + ((g636) & (!g637) & (g638) & (!g639) & (!g820) & (!g773)) + ((g636) & (!g637) & (g638) & (!g639) & (!g820) & (g773)) + ((g636) & (!g637) & (g638) & (g639) & (!g820) & (!g773)) + ((g636) & (!g637) & (g638) & (g639) & (!g820) & (g773)) + ((g636) & (!g637) & (g638) & (g639) & (g820) & (g773)) + ((g636) & (g637) & (!g638) & (!g639) & (!g820) & (!g773)) + ((g636) & (g637) & (!g638) & (!g639) & (g820) & (!g773)) + ((g636) & (g637) & (!g638) & (g639) & (!g820) & (!g773)) + ((g636) & (g637) & (!g638) & (g639) & (g820) & (!g773)) + ((g636) & (g637) & (!g638) & (g639) & (g820) & (g773)) + ((g636) & (g637) & (g638) & (!g639) & (!g820) & (!g773)) + ((g636) & (g637) & (g638) & (!g639) & (!g820) & (g773)) + ((g636) & (g637) & (g638) & (!g639) & (g820) & (!g773)) + ((g636) & (g637) & (g638) & (g639) & (!g820) & (!g773)) + ((g636) & (g637) & (g638) & (g639) & (!g820) & (g773)) + ((g636) & (g637) & (g638) & (g639) & (g820) & (!g773)) + ((g636) & (g637) & (g638) & (g639) & (g820) & (g773)));
	assign g1738 = (((!g641) & (!g642) & (!g643) & (g644) & (g820) & (g773)) + ((!g641) & (!g642) & (g643) & (!g644) & (!g820) & (g773)) + ((!g641) & (!g642) & (g643) & (g644) & (!g820) & (g773)) + ((!g641) & (!g642) & (g643) & (g644) & (g820) & (g773)) + ((!g641) & (g642) & (!g643) & (!g644) & (g820) & (!g773)) + ((!g641) & (g642) & (!g643) & (g644) & (g820) & (!g773)) + ((!g641) & (g642) & (!g643) & (g644) & (g820) & (g773)) + ((!g641) & (g642) & (g643) & (!g644) & (!g820) & (g773)) + ((!g641) & (g642) & (g643) & (!g644) & (g820) & (!g773)) + ((!g641) & (g642) & (g643) & (g644) & (!g820) & (g773)) + ((!g641) & (g642) & (g643) & (g644) & (g820) & (!g773)) + ((!g641) & (g642) & (g643) & (g644) & (g820) & (g773)) + ((g641) & (!g642) & (!g643) & (!g644) & (!g820) & (!g773)) + ((g641) & (!g642) & (!g643) & (g644) & (!g820) & (!g773)) + ((g641) & (!g642) & (!g643) & (g644) & (g820) & (g773)) + ((g641) & (!g642) & (g643) & (!g644) & (!g820) & (!g773)) + ((g641) & (!g642) & (g643) & (!g644) & (!g820) & (g773)) + ((g641) & (!g642) & (g643) & (g644) & (!g820) & (!g773)) + ((g641) & (!g642) & (g643) & (g644) & (!g820) & (g773)) + ((g641) & (!g642) & (g643) & (g644) & (g820) & (g773)) + ((g641) & (g642) & (!g643) & (!g644) & (!g820) & (!g773)) + ((g641) & (g642) & (!g643) & (!g644) & (g820) & (!g773)) + ((g641) & (g642) & (!g643) & (g644) & (!g820) & (!g773)) + ((g641) & (g642) & (!g643) & (g644) & (g820) & (!g773)) + ((g641) & (g642) & (!g643) & (g644) & (g820) & (g773)) + ((g641) & (g642) & (g643) & (!g644) & (!g820) & (!g773)) + ((g641) & (g642) & (g643) & (!g644) & (!g820) & (g773)) + ((g641) & (g642) & (g643) & (!g644) & (g820) & (!g773)) + ((g641) & (g642) & (g643) & (g644) & (!g820) & (!g773)) + ((g641) & (g642) & (g643) & (g644) & (!g820) & (g773)) + ((g641) & (g642) & (g643) & (g644) & (g820) & (!g773)) + ((g641) & (g642) & (g643) & (g644) & (g820) & (g773)));
	assign g1739 = (((!g646) & (!g647) & (!g648) & (g649) & (g820) & (g773)) + ((!g646) & (!g647) & (g648) & (!g649) & (!g820) & (g773)) + ((!g646) & (!g647) & (g648) & (g649) & (!g820) & (g773)) + ((!g646) & (!g647) & (g648) & (g649) & (g820) & (g773)) + ((!g646) & (g647) & (!g648) & (!g649) & (g820) & (!g773)) + ((!g646) & (g647) & (!g648) & (g649) & (g820) & (!g773)) + ((!g646) & (g647) & (!g648) & (g649) & (g820) & (g773)) + ((!g646) & (g647) & (g648) & (!g649) & (!g820) & (g773)) + ((!g646) & (g647) & (g648) & (!g649) & (g820) & (!g773)) + ((!g646) & (g647) & (g648) & (g649) & (!g820) & (g773)) + ((!g646) & (g647) & (g648) & (g649) & (g820) & (!g773)) + ((!g646) & (g647) & (g648) & (g649) & (g820) & (g773)) + ((g646) & (!g647) & (!g648) & (!g649) & (!g820) & (!g773)) + ((g646) & (!g647) & (!g648) & (g649) & (!g820) & (!g773)) + ((g646) & (!g647) & (!g648) & (g649) & (g820) & (g773)) + ((g646) & (!g647) & (g648) & (!g649) & (!g820) & (!g773)) + ((g646) & (!g647) & (g648) & (!g649) & (!g820) & (g773)) + ((g646) & (!g647) & (g648) & (g649) & (!g820) & (!g773)) + ((g646) & (!g647) & (g648) & (g649) & (!g820) & (g773)) + ((g646) & (!g647) & (g648) & (g649) & (g820) & (g773)) + ((g646) & (g647) & (!g648) & (!g649) & (!g820) & (!g773)) + ((g646) & (g647) & (!g648) & (!g649) & (g820) & (!g773)) + ((g646) & (g647) & (!g648) & (g649) & (!g820) & (!g773)) + ((g646) & (g647) & (!g648) & (g649) & (g820) & (!g773)) + ((g646) & (g647) & (!g648) & (g649) & (g820) & (g773)) + ((g646) & (g647) & (g648) & (!g649) & (!g820) & (!g773)) + ((g646) & (g647) & (g648) & (!g649) & (!g820) & (g773)) + ((g646) & (g647) & (g648) & (!g649) & (g820) & (!g773)) + ((g646) & (g647) & (g648) & (g649) & (!g820) & (!g773)) + ((g646) & (g647) & (g648) & (g649) & (!g820) & (g773)) + ((g646) & (g647) & (g648) & (g649) & (g820) & (!g773)) + ((g646) & (g647) & (g648) & (g649) & (g820) & (g773)));
	assign g1740 = (((!g1736) & (!g1737) & (!g1738) & (g1739) & (g677) & (g726)) + ((!g1736) & (!g1737) & (g1738) & (!g1739) & (!g677) & (g726)) + ((!g1736) & (!g1737) & (g1738) & (g1739) & (!g677) & (g726)) + ((!g1736) & (!g1737) & (g1738) & (g1739) & (g677) & (g726)) + ((!g1736) & (g1737) & (!g1738) & (!g1739) & (g677) & (!g726)) + ((!g1736) & (g1737) & (!g1738) & (g1739) & (g677) & (!g726)) + ((!g1736) & (g1737) & (!g1738) & (g1739) & (g677) & (g726)) + ((!g1736) & (g1737) & (g1738) & (!g1739) & (!g677) & (g726)) + ((!g1736) & (g1737) & (g1738) & (!g1739) & (g677) & (!g726)) + ((!g1736) & (g1737) & (g1738) & (g1739) & (!g677) & (g726)) + ((!g1736) & (g1737) & (g1738) & (g1739) & (g677) & (!g726)) + ((!g1736) & (g1737) & (g1738) & (g1739) & (g677) & (g726)) + ((g1736) & (!g1737) & (!g1738) & (!g1739) & (!g677) & (!g726)) + ((g1736) & (!g1737) & (!g1738) & (g1739) & (!g677) & (!g726)) + ((g1736) & (!g1737) & (!g1738) & (g1739) & (g677) & (g726)) + ((g1736) & (!g1737) & (g1738) & (!g1739) & (!g677) & (!g726)) + ((g1736) & (!g1737) & (g1738) & (!g1739) & (!g677) & (g726)) + ((g1736) & (!g1737) & (g1738) & (g1739) & (!g677) & (!g726)) + ((g1736) & (!g1737) & (g1738) & (g1739) & (!g677) & (g726)) + ((g1736) & (!g1737) & (g1738) & (g1739) & (g677) & (g726)) + ((g1736) & (g1737) & (!g1738) & (!g1739) & (!g677) & (!g726)) + ((g1736) & (g1737) & (!g1738) & (!g1739) & (g677) & (!g726)) + ((g1736) & (g1737) & (!g1738) & (g1739) & (!g677) & (!g726)) + ((g1736) & (g1737) & (!g1738) & (g1739) & (g677) & (!g726)) + ((g1736) & (g1737) & (!g1738) & (g1739) & (g677) & (g726)) + ((g1736) & (g1737) & (g1738) & (!g1739) & (!g677) & (!g726)) + ((g1736) & (g1737) & (g1738) & (!g1739) & (!g677) & (g726)) + ((g1736) & (g1737) & (g1738) & (!g1739) & (g677) & (!g726)) + ((g1736) & (g1737) & (g1738) & (g1739) & (!g677) & (!g726)) + ((g1736) & (g1737) & (g1738) & (g1739) & (!g677) & (g726)) + ((g1736) & (g1737) & (g1738) & (g1739) & (g677) & (!g726)) + ((g1736) & (g1737) & (g1738) & (g1739) & (g677) & (g726)));
	assign g1741 = (((!g652) & (!g653) & (!g654) & (g655) & (g677) & (g726)) + ((!g652) & (!g653) & (g654) & (!g655) & (!g677) & (g726)) + ((!g652) & (!g653) & (g654) & (g655) & (!g677) & (g726)) + ((!g652) & (!g653) & (g654) & (g655) & (g677) & (g726)) + ((!g652) & (g653) & (!g654) & (!g655) & (g677) & (!g726)) + ((!g652) & (g653) & (!g654) & (g655) & (g677) & (!g726)) + ((!g652) & (g653) & (!g654) & (g655) & (g677) & (g726)) + ((!g652) & (g653) & (g654) & (!g655) & (!g677) & (g726)) + ((!g652) & (g653) & (g654) & (!g655) & (g677) & (!g726)) + ((!g652) & (g653) & (g654) & (g655) & (!g677) & (g726)) + ((!g652) & (g653) & (g654) & (g655) & (g677) & (!g726)) + ((!g652) & (g653) & (g654) & (g655) & (g677) & (g726)) + ((g652) & (!g653) & (!g654) & (!g655) & (!g677) & (!g726)) + ((g652) & (!g653) & (!g654) & (g655) & (!g677) & (!g726)) + ((g652) & (!g653) & (!g654) & (g655) & (g677) & (g726)) + ((g652) & (!g653) & (g654) & (!g655) & (!g677) & (!g726)) + ((g652) & (!g653) & (g654) & (!g655) & (!g677) & (g726)) + ((g652) & (!g653) & (g654) & (g655) & (!g677) & (!g726)) + ((g652) & (!g653) & (g654) & (g655) & (!g677) & (g726)) + ((g652) & (!g653) & (g654) & (g655) & (g677) & (g726)) + ((g652) & (g653) & (!g654) & (!g655) & (!g677) & (!g726)) + ((g652) & (g653) & (!g654) & (!g655) & (g677) & (!g726)) + ((g652) & (g653) & (!g654) & (g655) & (!g677) & (!g726)) + ((g652) & (g653) & (!g654) & (g655) & (g677) & (!g726)) + ((g652) & (g653) & (!g654) & (g655) & (g677) & (g726)) + ((g652) & (g653) & (g654) & (!g655) & (!g677) & (!g726)) + ((g652) & (g653) & (g654) & (!g655) & (!g677) & (g726)) + ((g652) & (g653) & (g654) & (!g655) & (g677) & (!g726)) + ((g652) & (g653) & (g654) & (g655) & (!g677) & (!g726)) + ((g652) & (g653) & (g654) & (g655) & (!g677) & (g726)) + ((g652) & (g653) & (g654) & (g655) & (g677) & (!g726)) + ((g652) & (g653) & (g654) & (g655) & (g677) & (g726)));
	assign g1742 = (((!g677) & (!sk[16]) & (!g726) & (!g657) & (g658) & (!g659)) + ((!g677) & (!sk[16]) & (!g726) & (!g657) & (g658) & (g659)) + ((!g677) & (!sk[16]) & (!g726) & (g657) & (!g658) & (!g659)) + ((!g677) & (!sk[16]) & (!g726) & (g657) & (!g658) & (g659)) + ((!g677) & (!sk[16]) & (!g726) & (g657) & (g658) & (!g659)) + ((!g677) & (!sk[16]) & (!g726) & (g657) & (g658) & (g659)) + ((!g677) & (!sk[16]) & (g726) & (!g657) & (!g658) & (!g659)) + ((!g677) & (!sk[16]) & (g726) & (!g657) & (!g658) & (g659)) + ((!g677) & (!sk[16]) & (g726) & (!g657) & (g658) & (!g659)) + ((!g677) & (!sk[16]) & (g726) & (!g657) & (g658) & (g659)) + ((!g677) & (!sk[16]) & (g726) & (g657) & (!g658) & (!g659)) + ((!g677) & (!sk[16]) & (g726) & (g657) & (!g658) & (g659)) + ((!g677) & (!sk[16]) & (g726) & (g657) & (g658) & (!g659)) + ((!g677) & (!sk[16]) & (g726) & (g657) & (g658) & (g659)) + ((!g677) & (sk[16]) & (g726) & (!g657) & (!g658) & (g659)) + ((!g677) & (sk[16]) & (g726) & (!g657) & (g658) & (g659)) + ((!g677) & (sk[16]) & (g726) & (g657) & (!g658) & (g659)) + ((!g677) & (sk[16]) & (g726) & (g657) & (g658) & (g659)) + ((g677) & (!sk[16]) & (!g726) & (!g657) & (g658) & (!g659)) + ((g677) & (!sk[16]) & (!g726) & (!g657) & (g658) & (g659)) + ((g677) & (!sk[16]) & (!g726) & (g657) & (!g658) & (!g659)) + ((g677) & (!sk[16]) & (!g726) & (g657) & (!g658) & (g659)) + ((g677) & (!sk[16]) & (!g726) & (g657) & (g658) & (!g659)) + ((g677) & (!sk[16]) & (!g726) & (g657) & (g658) & (g659)) + ((g677) & (!sk[16]) & (g726) & (!g657) & (!g658) & (!g659)) + ((g677) & (!sk[16]) & (g726) & (!g657) & (!g658) & (g659)) + ((g677) & (!sk[16]) & (g726) & (!g657) & (g658) & (!g659)) + ((g677) & (!sk[16]) & (g726) & (!g657) & (g658) & (g659)) + ((g677) & (!sk[16]) & (g726) & (g657) & (!g658) & (!g659)) + ((g677) & (!sk[16]) & (g726) & (g657) & (!g658) & (g659)) + ((g677) & (!sk[16]) & (g726) & (g657) & (g658) & (!g659)) + ((g677) & (!sk[16]) & (g726) & (g657) & (g658) & (g659)) + ((g677) & (sk[16]) & (!g726) & (g657) & (!g658) & (!g659)) + ((g677) & (sk[16]) & (!g726) & (g657) & (!g658) & (g659)) + ((g677) & (sk[16]) & (!g726) & (g657) & (g658) & (!g659)) + ((g677) & (sk[16]) & (!g726) & (g657) & (g658) & (g659)) + ((g677) & (sk[16]) & (g726) & (!g657) & (g658) & (!g659)) + ((g677) & (sk[16]) & (g726) & (!g657) & (g658) & (g659)) + ((g677) & (sk[16]) & (g726) & (g657) & (g658) & (!g659)) + ((g677) & (sk[16]) & (g726) & (g657) & (g658) & (g659)));
	assign g1743 = (((!g661) & (!g662) & (!g663) & (g664) & (g677) & (g726)) + ((!g661) & (!g662) & (g663) & (!g664) & (!g677) & (g726)) + ((!g661) & (!g662) & (g663) & (g664) & (!g677) & (g726)) + ((!g661) & (!g662) & (g663) & (g664) & (g677) & (g726)) + ((!g661) & (g662) & (!g663) & (!g664) & (g677) & (!g726)) + ((!g661) & (g662) & (!g663) & (g664) & (g677) & (!g726)) + ((!g661) & (g662) & (!g663) & (g664) & (g677) & (g726)) + ((!g661) & (g662) & (g663) & (!g664) & (!g677) & (g726)) + ((!g661) & (g662) & (g663) & (!g664) & (g677) & (!g726)) + ((!g661) & (g662) & (g663) & (g664) & (!g677) & (g726)) + ((!g661) & (g662) & (g663) & (g664) & (g677) & (!g726)) + ((!g661) & (g662) & (g663) & (g664) & (g677) & (g726)) + ((g661) & (!g662) & (!g663) & (!g664) & (!g677) & (!g726)) + ((g661) & (!g662) & (!g663) & (g664) & (!g677) & (!g726)) + ((g661) & (!g662) & (!g663) & (g664) & (g677) & (g726)) + ((g661) & (!g662) & (g663) & (!g664) & (!g677) & (!g726)) + ((g661) & (!g662) & (g663) & (!g664) & (!g677) & (g726)) + ((g661) & (!g662) & (g663) & (g664) & (!g677) & (!g726)) + ((g661) & (!g662) & (g663) & (g664) & (!g677) & (g726)) + ((g661) & (!g662) & (g663) & (g664) & (g677) & (g726)) + ((g661) & (g662) & (!g663) & (!g664) & (!g677) & (!g726)) + ((g661) & (g662) & (!g663) & (!g664) & (g677) & (!g726)) + ((g661) & (g662) & (!g663) & (g664) & (!g677) & (!g726)) + ((g661) & (g662) & (!g663) & (g664) & (g677) & (!g726)) + ((g661) & (g662) & (!g663) & (g664) & (g677) & (g726)) + ((g661) & (g662) & (g663) & (!g664) & (!g677) & (!g726)) + ((g661) & (g662) & (g663) & (!g664) & (!g677) & (g726)) + ((g661) & (g662) & (g663) & (!g664) & (g677) & (!g726)) + ((g661) & (g662) & (g663) & (g664) & (!g677) & (!g726)) + ((g661) & (g662) & (g663) & (g664) & (!g677) & (g726)) + ((g661) & (g662) & (g663) & (g664) & (g677) & (!g726)) + ((g661) & (g662) & (g663) & (g664) & (g677) & (g726)));
	assign g1744 = (((!g666) & (!g667) & (!g668) & (g669) & (g677) & (g726)) + ((!g666) & (!g667) & (g668) & (!g669) & (!g677) & (g726)) + ((!g666) & (!g667) & (g668) & (g669) & (!g677) & (g726)) + ((!g666) & (!g667) & (g668) & (g669) & (g677) & (g726)) + ((!g666) & (g667) & (!g668) & (!g669) & (g677) & (!g726)) + ((!g666) & (g667) & (!g668) & (g669) & (g677) & (!g726)) + ((!g666) & (g667) & (!g668) & (g669) & (g677) & (g726)) + ((!g666) & (g667) & (g668) & (!g669) & (!g677) & (g726)) + ((!g666) & (g667) & (g668) & (!g669) & (g677) & (!g726)) + ((!g666) & (g667) & (g668) & (g669) & (!g677) & (g726)) + ((!g666) & (g667) & (g668) & (g669) & (g677) & (!g726)) + ((!g666) & (g667) & (g668) & (g669) & (g677) & (g726)) + ((g666) & (!g667) & (!g668) & (!g669) & (!g677) & (!g726)) + ((g666) & (!g667) & (!g668) & (g669) & (!g677) & (!g726)) + ((g666) & (!g667) & (!g668) & (g669) & (g677) & (g726)) + ((g666) & (!g667) & (g668) & (!g669) & (!g677) & (!g726)) + ((g666) & (!g667) & (g668) & (!g669) & (!g677) & (g726)) + ((g666) & (!g667) & (g668) & (g669) & (!g677) & (!g726)) + ((g666) & (!g667) & (g668) & (g669) & (!g677) & (g726)) + ((g666) & (!g667) & (g668) & (g669) & (g677) & (g726)) + ((g666) & (g667) & (!g668) & (!g669) & (!g677) & (!g726)) + ((g666) & (g667) & (!g668) & (!g669) & (g677) & (!g726)) + ((g666) & (g667) & (!g668) & (g669) & (!g677) & (!g726)) + ((g666) & (g667) & (!g668) & (g669) & (g677) & (!g726)) + ((g666) & (g667) & (!g668) & (g669) & (g677) & (g726)) + ((g666) & (g667) & (g668) & (!g669) & (!g677) & (!g726)) + ((g666) & (g667) & (g668) & (!g669) & (!g677) & (g726)) + ((g666) & (g667) & (g668) & (!g669) & (g677) & (!g726)) + ((g666) & (g667) & (g668) & (g669) & (!g677) & (!g726)) + ((g666) & (g667) & (g668) & (g669) & (!g677) & (g726)) + ((g666) & (g667) & (g668) & (g669) & (g677) & (!g726)) + ((g666) & (g667) & (g668) & (g669) & (g677) & (g726)));
	assign g1745 = (((!g820) & (!g773) & (!g1741) & (g1742) & (!g1743) & (!g1744)) + ((!g820) & (!g773) & (!g1741) & (g1742) & (!g1743) & (g1744)) + ((!g820) & (!g773) & (!g1741) & (g1742) & (g1743) & (!g1744)) + ((!g820) & (!g773) & (!g1741) & (g1742) & (g1743) & (g1744)) + ((!g820) & (!g773) & (g1741) & (g1742) & (!g1743) & (!g1744)) + ((!g820) & (!g773) & (g1741) & (g1742) & (!g1743) & (g1744)) + ((!g820) & (!g773) & (g1741) & (g1742) & (g1743) & (!g1744)) + ((!g820) & (!g773) & (g1741) & (g1742) & (g1743) & (g1744)) + ((!g820) & (g773) & (!g1741) & (!g1742) & (!g1743) & (g1744)) + ((!g820) & (g773) & (!g1741) & (!g1742) & (g1743) & (g1744)) + ((!g820) & (g773) & (!g1741) & (g1742) & (!g1743) & (g1744)) + ((!g820) & (g773) & (!g1741) & (g1742) & (g1743) & (g1744)) + ((!g820) & (g773) & (g1741) & (!g1742) & (!g1743) & (g1744)) + ((!g820) & (g773) & (g1741) & (!g1742) & (g1743) & (g1744)) + ((!g820) & (g773) & (g1741) & (g1742) & (!g1743) & (g1744)) + ((!g820) & (g773) & (g1741) & (g1742) & (g1743) & (g1744)) + ((g820) & (!g773) & (g1741) & (!g1742) & (!g1743) & (!g1744)) + ((g820) & (!g773) & (g1741) & (!g1742) & (!g1743) & (g1744)) + ((g820) & (!g773) & (g1741) & (!g1742) & (g1743) & (!g1744)) + ((g820) & (!g773) & (g1741) & (!g1742) & (g1743) & (g1744)) + ((g820) & (!g773) & (g1741) & (g1742) & (!g1743) & (!g1744)) + ((g820) & (!g773) & (g1741) & (g1742) & (!g1743) & (g1744)) + ((g820) & (!g773) & (g1741) & (g1742) & (g1743) & (!g1744)) + ((g820) & (!g773) & (g1741) & (g1742) & (g1743) & (g1744)) + ((g820) & (g773) & (!g1741) & (!g1742) & (g1743) & (!g1744)) + ((g820) & (g773) & (!g1741) & (!g1742) & (g1743) & (g1744)) + ((g820) & (g773) & (!g1741) & (g1742) & (g1743) & (!g1744)) + ((g820) & (g773) & (!g1741) & (g1742) & (g1743) & (g1744)) + ((g820) & (g773) & (g1741) & (!g1742) & (g1743) & (!g1744)) + ((g820) & (g773) & (g1741) & (!g1742) & (g1743) & (g1744)) + ((g820) & (g773) & (g1741) & (g1742) & (g1743) & (!g1744)) + ((g820) & (g773) & (g1741) & (g1742) & (g1743) & (g1744)));
	assign g1746 = (((!sk[20]) & (!g867) & (!g1740) & (g1745)) + ((!sk[20]) & (!g867) & (g1740) & (!g1745)) + ((!sk[20]) & (!g867) & (g1740) & (g1745)) + ((!sk[20]) & (g867) & (!g1740) & (g1745)) + ((!sk[20]) & (g867) & (g1740) & (!g1745)) + ((!sk[20]) & (g867) & (g1740) & (g1745)) + ((sk[20]) & (!g867) & (!g1740) & (g1745)) + ((sk[20]) & (!g867) & (g1740) & (g1745)) + ((sk[20]) & (g867) & (g1740) & (!g1745)) + ((sk[20]) & (g867) & (g1740) & (g1745)));
	assign g1747 = (((!g132) & (!g1706) & (!g1707) & (g1735) & (!sk[21]) & (!g1746)) + ((!g132) & (!g1706) & (!g1707) & (g1735) & (!sk[21]) & (g1746)) + ((!g132) & (!g1706) & (g1707) & (!g1735) & (!sk[21]) & (!g1746)) + ((!g132) & (!g1706) & (g1707) & (!g1735) & (!sk[21]) & (g1746)) + ((!g132) & (!g1706) & (g1707) & (!g1735) & (sk[21]) & (g1746)) + ((!g132) & (!g1706) & (g1707) & (g1735) & (!sk[21]) & (!g1746)) + ((!g132) & (!g1706) & (g1707) & (g1735) & (!sk[21]) & (g1746)) + ((!g132) & (!g1706) & (g1707) & (g1735) & (sk[21]) & (!g1746)) + ((!g132) & (!g1706) & (g1707) & (g1735) & (sk[21]) & (g1746)) + ((!g132) & (g1706) & (!g1707) & (!g1735) & (!sk[21]) & (!g1746)) + ((!g132) & (g1706) & (!g1707) & (!g1735) & (!sk[21]) & (g1746)) + ((!g132) & (g1706) & (!g1707) & (g1735) & (!sk[21]) & (!g1746)) + ((!g132) & (g1706) & (!g1707) & (g1735) & (!sk[21]) & (g1746)) + ((!g132) & (g1706) & (g1707) & (!g1735) & (!sk[21]) & (!g1746)) + ((!g132) & (g1706) & (g1707) & (!g1735) & (!sk[21]) & (g1746)) + ((!g132) & (g1706) & (g1707) & (g1735) & (!sk[21]) & (!g1746)) + ((!g132) & (g1706) & (g1707) & (g1735) & (!sk[21]) & (g1746)) + ((!g132) & (g1706) & (g1707) & (g1735) & (sk[21]) & (!g1746)) + ((!g132) & (g1706) & (g1707) & (g1735) & (sk[21]) & (g1746)) + ((g132) & (!g1706) & (!g1707) & (g1735) & (!sk[21]) & (!g1746)) + ((g132) & (!g1706) & (!g1707) & (g1735) & (!sk[21]) & (g1746)) + ((g132) & (!g1706) & (g1707) & (!g1735) & (!sk[21]) & (!g1746)) + ((g132) & (!g1706) & (g1707) & (!g1735) & (!sk[21]) & (g1746)) + ((g132) & (!g1706) & (g1707) & (!g1735) & (sk[21]) & (g1746)) + ((g132) & (!g1706) & (g1707) & (g1735) & (!sk[21]) & (!g1746)) + ((g132) & (!g1706) & (g1707) & (g1735) & (!sk[21]) & (g1746)) + ((g132) & (!g1706) & (g1707) & (g1735) & (sk[21]) & (g1746)) + ((g132) & (g1706) & (!g1707) & (!g1735) & (!sk[21]) & (!g1746)) + ((g132) & (g1706) & (!g1707) & (!g1735) & (!sk[21]) & (g1746)) + ((g132) & (g1706) & (!g1707) & (g1735) & (!sk[21]) & (!g1746)) + ((g132) & (g1706) & (!g1707) & (g1735) & (!sk[21]) & (g1746)) + ((g132) & (g1706) & (g1707) & (!g1735) & (!sk[21]) & (!g1746)) + ((g132) & (g1706) & (g1707) & (!g1735) & (!sk[21]) & (g1746)) + ((g132) & (g1706) & (g1707) & (g1735) & (!sk[21]) & (!g1746)) + ((g132) & (g1706) & (g1707) & (g1735) & (!sk[21]) & (g1746)));
	assign g1748 = (((!g1592) & (!g1593) & (!g1656) & (!sk[22]) & (g47)) + ((!g1592) & (!g1593) & (g1656) & (!sk[22]) & (!g47)) + ((!g1592) & (!g1593) & (g1656) & (!sk[22]) & (g47)) + ((!g1592) & (!g1593) & (g1656) & (sk[22]) & (!g47)) + ((!g1592) & (!g1593) & (g1656) & (sk[22]) & (g47)) + ((!g1592) & (g1593) & (!g1656) & (!sk[22]) & (!g47)) + ((!g1592) & (g1593) & (!g1656) & (!sk[22]) & (g47)) + ((!g1592) & (g1593) & (g1656) & (!sk[22]) & (!g47)) + ((!g1592) & (g1593) & (g1656) & (!sk[22]) & (g47)) + ((!g1592) & (g1593) & (g1656) & (sk[22]) & (!g47)) + ((!g1592) & (g1593) & (g1656) & (sk[22]) & (g47)) + ((g1592) & (!g1593) & (!g1656) & (!sk[22]) & (g47)) + ((g1592) & (!g1593) & (g1656) & (!sk[22]) & (!g47)) + ((g1592) & (!g1593) & (g1656) & (!sk[22]) & (g47)) + ((g1592) & (g1593) & (!g1656) & (!sk[22]) & (!g47)) + ((g1592) & (g1593) & (!g1656) & (!sk[22]) & (g47)) + ((g1592) & (g1593) & (!g1656) & (sk[22]) & (g47)) + ((g1592) & (g1593) & (g1656) & (!sk[22]) & (!g47)) + ((g1592) & (g1593) & (g1656) & (!sk[22]) & (g47)) + ((g1592) & (g1593) & (g1656) & (sk[22]) & (g47)));
	assign g1749 = (((!g682) & (!g683) & (!g684) & (g685) & (g820) & (g773)) + ((!g682) & (!g683) & (g684) & (!g685) & (!g820) & (g773)) + ((!g682) & (!g683) & (g684) & (g685) & (!g820) & (g773)) + ((!g682) & (!g683) & (g684) & (g685) & (g820) & (g773)) + ((!g682) & (g683) & (!g684) & (!g685) & (g820) & (!g773)) + ((!g682) & (g683) & (!g684) & (g685) & (g820) & (!g773)) + ((!g682) & (g683) & (!g684) & (g685) & (g820) & (g773)) + ((!g682) & (g683) & (g684) & (!g685) & (!g820) & (g773)) + ((!g682) & (g683) & (g684) & (!g685) & (g820) & (!g773)) + ((!g682) & (g683) & (g684) & (g685) & (!g820) & (g773)) + ((!g682) & (g683) & (g684) & (g685) & (g820) & (!g773)) + ((!g682) & (g683) & (g684) & (g685) & (g820) & (g773)) + ((g682) & (!g683) & (!g684) & (!g685) & (!g820) & (!g773)) + ((g682) & (!g683) & (!g684) & (g685) & (!g820) & (!g773)) + ((g682) & (!g683) & (!g684) & (g685) & (g820) & (g773)) + ((g682) & (!g683) & (g684) & (!g685) & (!g820) & (!g773)) + ((g682) & (!g683) & (g684) & (!g685) & (!g820) & (g773)) + ((g682) & (!g683) & (g684) & (g685) & (!g820) & (!g773)) + ((g682) & (!g683) & (g684) & (g685) & (!g820) & (g773)) + ((g682) & (!g683) & (g684) & (g685) & (g820) & (g773)) + ((g682) & (g683) & (!g684) & (!g685) & (!g820) & (!g773)) + ((g682) & (g683) & (!g684) & (!g685) & (g820) & (!g773)) + ((g682) & (g683) & (!g684) & (g685) & (!g820) & (!g773)) + ((g682) & (g683) & (!g684) & (g685) & (g820) & (!g773)) + ((g682) & (g683) & (!g684) & (g685) & (g820) & (g773)) + ((g682) & (g683) & (g684) & (!g685) & (!g820) & (!g773)) + ((g682) & (g683) & (g684) & (!g685) & (!g820) & (g773)) + ((g682) & (g683) & (g684) & (!g685) & (g820) & (!g773)) + ((g682) & (g683) & (g684) & (g685) & (!g820) & (!g773)) + ((g682) & (g683) & (g684) & (g685) & (!g820) & (g773)) + ((g682) & (g683) & (g684) & (g685) & (g820) & (!g773)) + ((g682) & (g683) & (g684) & (g685) & (g820) & (g773)));
	assign g1750 = (((!g687) & (!g688) & (!g689) & (g690) & (g820) & (g773)) + ((!g687) & (!g688) & (g689) & (!g690) & (!g820) & (g773)) + ((!g687) & (!g688) & (g689) & (g690) & (!g820) & (g773)) + ((!g687) & (!g688) & (g689) & (g690) & (g820) & (g773)) + ((!g687) & (g688) & (!g689) & (!g690) & (g820) & (!g773)) + ((!g687) & (g688) & (!g689) & (g690) & (g820) & (!g773)) + ((!g687) & (g688) & (!g689) & (g690) & (g820) & (g773)) + ((!g687) & (g688) & (g689) & (!g690) & (!g820) & (g773)) + ((!g687) & (g688) & (g689) & (!g690) & (g820) & (!g773)) + ((!g687) & (g688) & (g689) & (g690) & (!g820) & (g773)) + ((!g687) & (g688) & (g689) & (g690) & (g820) & (!g773)) + ((!g687) & (g688) & (g689) & (g690) & (g820) & (g773)) + ((g687) & (!g688) & (!g689) & (!g690) & (!g820) & (!g773)) + ((g687) & (!g688) & (!g689) & (g690) & (!g820) & (!g773)) + ((g687) & (!g688) & (!g689) & (g690) & (g820) & (g773)) + ((g687) & (!g688) & (g689) & (!g690) & (!g820) & (!g773)) + ((g687) & (!g688) & (g689) & (!g690) & (!g820) & (g773)) + ((g687) & (!g688) & (g689) & (g690) & (!g820) & (!g773)) + ((g687) & (!g688) & (g689) & (g690) & (!g820) & (g773)) + ((g687) & (!g688) & (g689) & (g690) & (g820) & (g773)) + ((g687) & (g688) & (!g689) & (!g690) & (!g820) & (!g773)) + ((g687) & (g688) & (!g689) & (!g690) & (g820) & (!g773)) + ((g687) & (g688) & (!g689) & (g690) & (!g820) & (!g773)) + ((g687) & (g688) & (!g689) & (g690) & (g820) & (!g773)) + ((g687) & (g688) & (!g689) & (g690) & (g820) & (g773)) + ((g687) & (g688) & (g689) & (!g690) & (!g820) & (!g773)) + ((g687) & (g688) & (g689) & (!g690) & (!g820) & (g773)) + ((g687) & (g688) & (g689) & (!g690) & (g820) & (!g773)) + ((g687) & (g688) & (g689) & (g690) & (!g820) & (!g773)) + ((g687) & (g688) & (g689) & (g690) & (!g820) & (g773)) + ((g687) & (g688) & (g689) & (g690) & (g820) & (!g773)) + ((g687) & (g688) & (g689) & (g690) & (g820) & (g773)));
	assign g1751 = (((!g692) & (!g693) & (!g694) & (g695) & (g820) & (g773)) + ((!g692) & (!g693) & (g694) & (!g695) & (!g820) & (g773)) + ((!g692) & (!g693) & (g694) & (g695) & (!g820) & (g773)) + ((!g692) & (!g693) & (g694) & (g695) & (g820) & (g773)) + ((!g692) & (g693) & (!g694) & (!g695) & (g820) & (!g773)) + ((!g692) & (g693) & (!g694) & (g695) & (g820) & (!g773)) + ((!g692) & (g693) & (!g694) & (g695) & (g820) & (g773)) + ((!g692) & (g693) & (g694) & (!g695) & (!g820) & (g773)) + ((!g692) & (g693) & (g694) & (!g695) & (g820) & (!g773)) + ((!g692) & (g693) & (g694) & (g695) & (!g820) & (g773)) + ((!g692) & (g693) & (g694) & (g695) & (g820) & (!g773)) + ((!g692) & (g693) & (g694) & (g695) & (g820) & (g773)) + ((g692) & (!g693) & (!g694) & (!g695) & (!g820) & (!g773)) + ((g692) & (!g693) & (!g694) & (g695) & (!g820) & (!g773)) + ((g692) & (!g693) & (!g694) & (g695) & (g820) & (g773)) + ((g692) & (!g693) & (g694) & (!g695) & (!g820) & (!g773)) + ((g692) & (!g693) & (g694) & (!g695) & (!g820) & (g773)) + ((g692) & (!g693) & (g694) & (g695) & (!g820) & (!g773)) + ((g692) & (!g693) & (g694) & (g695) & (!g820) & (g773)) + ((g692) & (!g693) & (g694) & (g695) & (g820) & (g773)) + ((g692) & (g693) & (!g694) & (!g695) & (!g820) & (!g773)) + ((g692) & (g693) & (!g694) & (!g695) & (g820) & (!g773)) + ((g692) & (g693) & (!g694) & (g695) & (!g820) & (!g773)) + ((g692) & (g693) & (!g694) & (g695) & (g820) & (!g773)) + ((g692) & (g693) & (!g694) & (g695) & (g820) & (g773)) + ((g692) & (g693) & (g694) & (!g695) & (!g820) & (!g773)) + ((g692) & (g693) & (g694) & (!g695) & (!g820) & (g773)) + ((g692) & (g693) & (g694) & (!g695) & (g820) & (!g773)) + ((g692) & (g693) & (g694) & (g695) & (!g820) & (!g773)) + ((g692) & (g693) & (g694) & (g695) & (!g820) & (g773)) + ((g692) & (g693) & (g694) & (g695) & (g820) & (!g773)) + ((g692) & (g693) & (g694) & (g695) & (g820) & (g773)));
	assign g1752 = (((!g697) & (!g698) & (!g699) & (g700) & (g820) & (g773)) + ((!g697) & (!g698) & (g699) & (!g700) & (!g820) & (g773)) + ((!g697) & (!g698) & (g699) & (g700) & (!g820) & (g773)) + ((!g697) & (!g698) & (g699) & (g700) & (g820) & (g773)) + ((!g697) & (g698) & (!g699) & (!g700) & (g820) & (!g773)) + ((!g697) & (g698) & (!g699) & (g700) & (g820) & (!g773)) + ((!g697) & (g698) & (!g699) & (g700) & (g820) & (g773)) + ((!g697) & (g698) & (g699) & (!g700) & (!g820) & (g773)) + ((!g697) & (g698) & (g699) & (!g700) & (g820) & (!g773)) + ((!g697) & (g698) & (g699) & (g700) & (!g820) & (g773)) + ((!g697) & (g698) & (g699) & (g700) & (g820) & (!g773)) + ((!g697) & (g698) & (g699) & (g700) & (g820) & (g773)) + ((g697) & (!g698) & (!g699) & (!g700) & (!g820) & (!g773)) + ((g697) & (!g698) & (!g699) & (g700) & (!g820) & (!g773)) + ((g697) & (!g698) & (!g699) & (g700) & (g820) & (g773)) + ((g697) & (!g698) & (g699) & (!g700) & (!g820) & (!g773)) + ((g697) & (!g698) & (g699) & (!g700) & (!g820) & (g773)) + ((g697) & (!g698) & (g699) & (g700) & (!g820) & (!g773)) + ((g697) & (!g698) & (g699) & (g700) & (!g820) & (g773)) + ((g697) & (!g698) & (g699) & (g700) & (g820) & (g773)) + ((g697) & (g698) & (!g699) & (!g700) & (!g820) & (!g773)) + ((g697) & (g698) & (!g699) & (!g700) & (g820) & (!g773)) + ((g697) & (g698) & (!g699) & (g700) & (!g820) & (!g773)) + ((g697) & (g698) & (!g699) & (g700) & (g820) & (!g773)) + ((g697) & (g698) & (!g699) & (g700) & (g820) & (g773)) + ((g697) & (g698) & (g699) & (!g700) & (!g820) & (!g773)) + ((g697) & (g698) & (g699) & (!g700) & (!g820) & (g773)) + ((g697) & (g698) & (g699) & (!g700) & (g820) & (!g773)) + ((g697) & (g698) & (g699) & (g700) & (!g820) & (!g773)) + ((g697) & (g698) & (g699) & (g700) & (!g820) & (g773)) + ((g697) & (g698) & (g699) & (g700) & (g820) & (!g773)) + ((g697) & (g698) & (g699) & (g700) & (g820) & (g773)));
	assign g1753 = (((!g1749) & (!g1750) & (!g1751) & (g1752) & (g677) & (g726)) + ((!g1749) & (!g1750) & (g1751) & (!g1752) & (!g677) & (g726)) + ((!g1749) & (!g1750) & (g1751) & (g1752) & (!g677) & (g726)) + ((!g1749) & (!g1750) & (g1751) & (g1752) & (g677) & (g726)) + ((!g1749) & (g1750) & (!g1751) & (!g1752) & (g677) & (!g726)) + ((!g1749) & (g1750) & (!g1751) & (g1752) & (g677) & (!g726)) + ((!g1749) & (g1750) & (!g1751) & (g1752) & (g677) & (g726)) + ((!g1749) & (g1750) & (g1751) & (!g1752) & (!g677) & (g726)) + ((!g1749) & (g1750) & (g1751) & (!g1752) & (g677) & (!g726)) + ((!g1749) & (g1750) & (g1751) & (g1752) & (!g677) & (g726)) + ((!g1749) & (g1750) & (g1751) & (g1752) & (g677) & (!g726)) + ((!g1749) & (g1750) & (g1751) & (g1752) & (g677) & (g726)) + ((g1749) & (!g1750) & (!g1751) & (!g1752) & (!g677) & (!g726)) + ((g1749) & (!g1750) & (!g1751) & (g1752) & (!g677) & (!g726)) + ((g1749) & (!g1750) & (!g1751) & (g1752) & (g677) & (g726)) + ((g1749) & (!g1750) & (g1751) & (!g1752) & (!g677) & (!g726)) + ((g1749) & (!g1750) & (g1751) & (!g1752) & (!g677) & (g726)) + ((g1749) & (!g1750) & (g1751) & (g1752) & (!g677) & (!g726)) + ((g1749) & (!g1750) & (g1751) & (g1752) & (!g677) & (g726)) + ((g1749) & (!g1750) & (g1751) & (g1752) & (g677) & (g726)) + ((g1749) & (g1750) & (!g1751) & (!g1752) & (!g677) & (!g726)) + ((g1749) & (g1750) & (!g1751) & (!g1752) & (g677) & (!g726)) + ((g1749) & (g1750) & (!g1751) & (g1752) & (!g677) & (!g726)) + ((g1749) & (g1750) & (!g1751) & (g1752) & (g677) & (!g726)) + ((g1749) & (g1750) & (!g1751) & (g1752) & (g677) & (g726)) + ((g1749) & (g1750) & (g1751) & (!g1752) & (!g677) & (!g726)) + ((g1749) & (g1750) & (g1751) & (!g1752) & (!g677) & (g726)) + ((g1749) & (g1750) & (g1751) & (!g1752) & (g677) & (!g726)) + ((g1749) & (g1750) & (g1751) & (g1752) & (!g677) & (!g726)) + ((g1749) & (g1750) & (g1751) & (g1752) & (!g677) & (g726)) + ((g1749) & (g1750) & (g1751) & (g1752) & (g677) & (!g726)) + ((g1749) & (g1750) & (g1751) & (g1752) & (g677) & (g726)));
	assign g1754 = (((!g703) & (!g704) & (!g705) & (g706) & (g677) & (g726)) + ((!g703) & (!g704) & (g705) & (!g706) & (!g677) & (g726)) + ((!g703) & (!g704) & (g705) & (g706) & (!g677) & (g726)) + ((!g703) & (!g704) & (g705) & (g706) & (g677) & (g726)) + ((!g703) & (g704) & (!g705) & (!g706) & (g677) & (!g726)) + ((!g703) & (g704) & (!g705) & (g706) & (g677) & (!g726)) + ((!g703) & (g704) & (!g705) & (g706) & (g677) & (g726)) + ((!g703) & (g704) & (g705) & (!g706) & (!g677) & (g726)) + ((!g703) & (g704) & (g705) & (!g706) & (g677) & (!g726)) + ((!g703) & (g704) & (g705) & (g706) & (!g677) & (g726)) + ((!g703) & (g704) & (g705) & (g706) & (g677) & (!g726)) + ((!g703) & (g704) & (g705) & (g706) & (g677) & (g726)) + ((g703) & (!g704) & (!g705) & (!g706) & (!g677) & (!g726)) + ((g703) & (!g704) & (!g705) & (g706) & (!g677) & (!g726)) + ((g703) & (!g704) & (!g705) & (g706) & (g677) & (g726)) + ((g703) & (!g704) & (g705) & (!g706) & (!g677) & (!g726)) + ((g703) & (!g704) & (g705) & (!g706) & (!g677) & (g726)) + ((g703) & (!g704) & (g705) & (g706) & (!g677) & (!g726)) + ((g703) & (!g704) & (g705) & (g706) & (!g677) & (g726)) + ((g703) & (!g704) & (g705) & (g706) & (g677) & (g726)) + ((g703) & (g704) & (!g705) & (!g706) & (!g677) & (!g726)) + ((g703) & (g704) & (!g705) & (!g706) & (g677) & (!g726)) + ((g703) & (g704) & (!g705) & (g706) & (!g677) & (!g726)) + ((g703) & (g704) & (!g705) & (g706) & (g677) & (!g726)) + ((g703) & (g704) & (!g705) & (g706) & (g677) & (g726)) + ((g703) & (g704) & (g705) & (!g706) & (!g677) & (!g726)) + ((g703) & (g704) & (g705) & (!g706) & (!g677) & (g726)) + ((g703) & (g704) & (g705) & (!g706) & (g677) & (!g726)) + ((g703) & (g704) & (g705) & (g706) & (!g677) & (!g726)) + ((g703) & (g704) & (g705) & (g706) & (!g677) & (g726)) + ((g703) & (g704) & (g705) & (g706) & (g677) & (!g726)) + ((g703) & (g704) & (g705) & (g706) & (g677) & (g726)));
	assign g1755 = (((!g677) & (!g726) & (!sk[29]) & (!g708) & (g709) & (!g710)) + ((!g677) & (!g726) & (!sk[29]) & (!g708) & (g709) & (g710)) + ((!g677) & (!g726) & (!sk[29]) & (g708) & (!g709) & (!g710)) + ((!g677) & (!g726) & (!sk[29]) & (g708) & (!g709) & (g710)) + ((!g677) & (!g726) & (!sk[29]) & (g708) & (g709) & (!g710)) + ((!g677) & (!g726) & (!sk[29]) & (g708) & (g709) & (g710)) + ((!g677) & (g726) & (!sk[29]) & (!g708) & (!g709) & (!g710)) + ((!g677) & (g726) & (!sk[29]) & (!g708) & (!g709) & (g710)) + ((!g677) & (g726) & (!sk[29]) & (!g708) & (g709) & (!g710)) + ((!g677) & (g726) & (!sk[29]) & (!g708) & (g709) & (g710)) + ((!g677) & (g726) & (!sk[29]) & (g708) & (!g709) & (!g710)) + ((!g677) & (g726) & (!sk[29]) & (g708) & (!g709) & (g710)) + ((!g677) & (g726) & (!sk[29]) & (g708) & (g709) & (!g710)) + ((!g677) & (g726) & (!sk[29]) & (g708) & (g709) & (g710)) + ((!g677) & (g726) & (sk[29]) & (!g708) & (!g709) & (g710)) + ((!g677) & (g726) & (sk[29]) & (!g708) & (g709) & (g710)) + ((!g677) & (g726) & (sk[29]) & (g708) & (!g709) & (g710)) + ((!g677) & (g726) & (sk[29]) & (g708) & (g709) & (g710)) + ((g677) & (!g726) & (!sk[29]) & (!g708) & (g709) & (!g710)) + ((g677) & (!g726) & (!sk[29]) & (!g708) & (g709) & (g710)) + ((g677) & (!g726) & (!sk[29]) & (g708) & (!g709) & (!g710)) + ((g677) & (!g726) & (!sk[29]) & (g708) & (!g709) & (g710)) + ((g677) & (!g726) & (!sk[29]) & (g708) & (g709) & (!g710)) + ((g677) & (!g726) & (!sk[29]) & (g708) & (g709) & (g710)) + ((g677) & (!g726) & (sk[29]) & (g708) & (!g709) & (!g710)) + ((g677) & (!g726) & (sk[29]) & (g708) & (!g709) & (g710)) + ((g677) & (!g726) & (sk[29]) & (g708) & (g709) & (!g710)) + ((g677) & (!g726) & (sk[29]) & (g708) & (g709) & (g710)) + ((g677) & (g726) & (!sk[29]) & (!g708) & (!g709) & (!g710)) + ((g677) & (g726) & (!sk[29]) & (!g708) & (!g709) & (g710)) + ((g677) & (g726) & (!sk[29]) & (!g708) & (g709) & (!g710)) + ((g677) & (g726) & (!sk[29]) & (!g708) & (g709) & (g710)) + ((g677) & (g726) & (!sk[29]) & (g708) & (!g709) & (!g710)) + ((g677) & (g726) & (!sk[29]) & (g708) & (!g709) & (g710)) + ((g677) & (g726) & (!sk[29]) & (g708) & (g709) & (!g710)) + ((g677) & (g726) & (!sk[29]) & (g708) & (g709) & (g710)) + ((g677) & (g726) & (sk[29]) & (!g708) & (g709) & (!g710)) + ((g677) & (g726) & (sk[29]) & (!g708) & (g709) & (g710)) + ((g677) & (g726) & (sk[29]) & (g708) & (g709) & (!g710)) + ((g677) & (g726) & (sk[29]) & (g708) & (g709) & (g710)));
	assign g1756 = (((!g712) & (!g713) & (!g714) & (g715) & (g677) & (g726)) + ((!g712) & (!g713) & (g714) & (!g715) & (!g677) & (g726)) + ((!g712) & (!g713) & (g714) & (g715) & (!g677) & (g726)) + ((!g712) & (!g713) & (g714) & (g715) & (g677) & (g726)) + ((!g712) & (g713) & (!g714) & (!g715) & (g677) & (!g726)) + ((!g712) & (g713) & (!g714) & (g715) & (g677) & (!g726)) + ((!g712) & (g713) & (!g714) & (g715) & (g677) & (g726)) + ((!g712) & (g713) & (g714) & (!g715) & (!g677) & (g726)) + ((!g712) & (g713) & (g714) & (!g715) & (g677) & (!g726)) + ((!g712) & (g713) & (g714) & (g715) & (!g677) & (g726)) + ((!g712) & (g713) & (g714) & (g715) & (g677) & (!g726)) + ((!g712) & (g713) & (g714) & (g715) & (g677) & (g726)) + ((g712) & (!g713) & (!g714) & (!g715) & (!g677) & (!g726)) + ((g712) & (!g713) & (!g714) & (g715) & (!g677) & (!g726)) + ((g712) & (!g713) & (!g714) & (g715) & (g677) & (g726)) + ((g712) & (!g713) & (g714) & (!g715) & (!g677) & (!g726)) + ((g712) & (!g713) & (g714) & (!g715) & (!g677) & (g726)) + ((g712) & (!g713) & (g714) & (g715) & (!g677) & (!g726)) + ((g712) & (!g713) & (g714) & (g715) & (!g677) & (g726)) + ((g712) & (!g713) & (g714) & (g715) & (g677) & (g726)) + ((g712) & (g713) & (!g714) & (!g715) & (!g677) & (!g726)) + ((g712) & (g713) & (!g714) & (!g715) & (g677) & (!g726)) + ((g712) & (g713) & (!g714) & (g715) & (!g677) & (!g726)) + ((g712) & (g713) & (!g714) & (g715) & (g677) & (!g726)) + ((g712) & (g713) & (!g714) & (g715) & (g677) & (g726)) + ((g712) & (g713) & (g714) & (!g715) & (!g677) & (!g726)) + ((g712) & (g713) & (g714) & (!g715) & (!g677) & (g726)) + ((g712) & (g713) & (g714) & (!g715) & (g677) & (!g726)) + ((g712) & (g713) & (g714) & (g715) & (!g677) & (!g726)) + ((g712) & (g713) & (g714) & (g715) & (!g677) & (g726)) + ((g712) & (g713) & (g714) & (g715) & (g677) & (!g726)) + ((g712) & (g713) & (g714) & (g715) & (g677) & (g726)));
	assign g1757 = (((!g717) & (!g718) & (!g719) & (g720) & (g677) & (g726)) + ((!g717) & (!g718) & (g719) & (!g720) & (!g677) & (g726)) + ((!g717) & (!g718) & (g719) & (g720) & (!g677) & (g726)) + ((!g717) & (!g718) & (g719) & (g720) & (g677) & (g726)) + ((!g717) & (g718) & (!g719) & (!g720) & (g677) & (!g726)) + ((!g717) & (g718) & (!g719) & (g720) & (g677) & (!g726)) + ((!g717) & (g718) & (!g719) & (g720) & (g677) & (g726)) + ((!g717) & (g718) & (g719) & (!g720) & (!g677) & (g726)) + ((!g717) & (g718) & (g719) & (!g720) & (g677) & (!g726)) + ((!g717) & (g718) & (g719) & (g720) & (!g677) & (g726)) + ((!g717) & (g718) & (g719) & (g720) & (g677) & (!g726)) + ((!g717) & (g718) & (g719) & (g720) & (g677) & (g726)) + ((g717) & (!g718) & (!g719) & (!g720) & (!g677) & (!g726)) + ((g717) & (!g718) & (!g719) & (g720) & (!g677) & (!g726)) + ((g717) & (!g718) & (!g719) & (g720) & (g677) & (g726)) + ((g717) & (!g718) & (g719) & (!g720) & (!g677) & (!g726)) + ((g717) & (!g718) & (g719) & (!g720) & (!g677) & (g726)) + ((g717) & (!g718) & (g719) & (g720) & (!g677) & (!g726)) + ((g717) & (!g718) & (g719) & (g720) & (!g677) & (g726)) + ((g717) & (!g718) & (g719) & (g720) & (g677) & (g726)) + ((g717) & (g718) & (!g719) & (!g720) & (!g677) & (!g726)) + ((g717) & (g718) & (!g719) & (!g720) & (g677) & (!g726)) + ((g717) & (g718) & (!g719) & (g720) & (!g677) & (!g726)) + ((g717) & (g718) & (!g719) & (g720) & (g677) & (!g726)) + ((g717) & (g718) & (!g719) & (g720) & (g677) & (g726)) + ((g717) & (g718) & (g719) & (!g720) & (!g677) & (!g726)) + ((g717) & (g718) & (g719) & (!g720) & (!g677) & (g726)) + ((g717) & (g718) & (g719) & (!g720) & (g677) & (!g726)) + ((g717) & (g718) & (g719) & (g720) & (!g677) & (!g726)) + ((g717) & (g718) & (g719) & (g720) & (!g677) & (g726)) + ((g717) & (g718) & (g719) & (g720) & (g677) & (!g726)) + ((g717) & (g718) & (g719) & (g720) & (g677) & (g726)));
	assign g1758 = (((!g820) & (!g773) & (!g1754) & (g1755) & (!g1756) & (!g1757)) + ((!g820) & (!g773) & (!g1754) & (g1755) & (!g1756) & (g1757)) + ((!g820) & (!g773) & (!g1754) & (g1755) & (g1756) & (!g1757)) + ((!g820) & (!g773) & (!g1754) & (g1755) & (g1756) & (g1757)) + ((!g820) & (!g773) & (g1754) & (g1755) & (!g1756) & (!g1757)) + ((!g820) & (!g773) & (g1754) & (g1755) & (!g1756) & (g1757)) + ((!g820) & (!g773) & (g1754) & (g1755) & (g1756) & (!g1757)) + ((!g820) & (!g773) & (g1754) & (g1755) & (g1756) & (g1757)) + ((!g820) & (g773) & (!g1754) & (!g1755) & (!g1756) & (g1757)) + ((!g820) & (g773) & (!g1754) & (!g1755) & (g1756) & (g1757)) + ((!g820) & (g773) & (!g1754) & (g1755) & (!g1756) & (g1757)) + ((!g820) & (g773) & (!g1754) & (g1755) & (g1756) & (g1757)) + ((!g820) & (g773) & (g1754) & (!g1755) & (!g1756) & (g1757)) + ((!g820) & (g773) & (g1754) & (!g1755) & (g1756) & (g1757)) + ((!g820) & (g773) & (g1754) & (g1755) & (!g1756) & (g1757)) + ((!g820) & (g773) & (g1754) & (g1755) & (g1756) & (g1757)) + ((g820) & (!g773) & (g1754) & (!g1755) & (!g1756) & (!g1757)) + ((g820) & (!g773) & (g1754) & (!g1755) & (!g1756) & (g1757)) + ((g820) & (!g773) & (g1754) & (!g1755) & (g1756) & (!g1757)) + ((g820) & (!g773) & (g1754) & (!g1755) & (g1756) & (g1757)) + ((g820) & (!g773) & (g1754) & (g1755) & (!g1756) & (!g1757)) + ((g820) & (!g773) & (g1754) & (g1755) & (!g1756) & (g1757)) + ((g820) & (!g773) & (g1754) & (g1755) & (g1756) & (!g1757)) + ((g820) & (!g773) & (g1754) & (g1755) & (g1756) & (g1757)) + ((g820) & (g773) & (!g1754) & (!g1755) & (g1756) & (!g1757)) + ((g820) & (g773) & (!g1754) & (!g1755) & (g1756) & (g1757)) + ((g820) & (g773) & (!g1754) & (g1755) & (g1756) & (!g1757)) + ((g820) & (g773) & (!g1754) & (g1755) & (g1756) & (g1757)) + ((g820) & (g773) & (g1754) & (!g1755) & (g1756) & (!g1757)) + ((g820) & (g773) & (g1754) & (!g1755) & (g1756) & (g1757)) + ((g820) & (g773) & (g1754) & (g1755) & (g1756) & (!g1757)) + ((g820) & (g773) & (g1754) & (g1755) & (g1756) & (g1757)));
	assign g1759 = (((!sk[33]) & (!g867) & (!g1753) & (g1758)) + ((!sk[33]) & (!g867) & (g1753) & (!g1758)) + ((!sk[33]) & (!g867) & (g1753) & (g1758)) + ((!sk[33]) & (g867) & (!g1753) & (g1758)) + ((!sk[33]) & (g867) & (g1753) & (!g1758)) + ((!sk[33]) & (g867) & (g1753) & (g1758)) + ((sk[33]) & (!g867) & (!g1753) & (g1758)) + ((sk[33]) & (!g867) & (g1753) & (g1758)) + ((sk[33]) & (g867) & (g1753) & (!g1758)) + ((sk[33]) & (g867) & (g1753) & (g1758)));
	assign g1760 = (((!g132) & (!g1706) & (!g1707) & (!sk[34]) & (g1748) & (!g1759)) + ((!g132) & (!g1706) & (!g1707) & (!sk[34]) & (g1748) & (g1759)) + ((!g132) & (!g1706) & (g1707) & (!sk[34]) & (!g1748) & (!g1759)) + ((!g132) & (!g1706) & (g1707) & (!sk[34]) & (!g1748) & (g1759)) + ((!g132) & (!g1706) & (g1707) & (!sk[34]) & (g1748) & (!g1759)) + ((!g132) & (!g1706) & (g1707) & (!sk[34]) & (g1748) & (g1759)) + ((!g132) & (!g1706) & (g1707) & (sk[34]) & (!g1748) & (g1759)) + ((!g132) & (!g1706) & (g1707) & (sk[34]) & (g1748) & (!g1759)) + ((!g132) & (!g1706) & (g1707) & (sk[34]) & (g1748) & (g1759)) + ((!g132) & (g1706) & (!g1707) & (!sk[34]) & (!g1748) & (!g1759)) + ((!g132) & (g1706) & (!g1707) & (!sk[34]) & (!g1748) & (g1759)) + ((!g132) & (g1706) & (!g1707) & (!sk[34]) & (g1748) & (!g1759)) + ((!g132) & (g1706) & (!g1707) & (!sk[34]) & (g1748) & (g1759)) + ((!g132) & (g1706) & (g1707) & (!sk[34]) & (!g1748) & (!g1759)) + ((!g132) & (g1706) & (g1707) & (!sk[34]) & (!g1748) & (g1759)) + ((!g132) & (g1706) & (g1707) & (!sk[34]) & (g1748) & (!g1759)) + ((!g132) & (g1706) & (g1707) & (!sk[34]) & (g1748) & (g1759)) + ((!g132) & (g1706) & (g1707) & (sk[34]) & (g1748) & (!g1759)) + ((!g132) & (g1706) & (g1707) & (sk[34]) & (g1748) & (g1759)) + ((g132) & (!g1706) & (!g1707) & (!sk[34]) & (g1748) & (!g1759)) + ((g132) & (!g1706) & (!g1707) & (!sk[34]) & (g1748) & (g1759)) + ((g132) & (!g1706) & (g1707) & (!sk[34]) & (!g1748) & (!g1759)) + ((g132) & (!g1706) & (g1707) & (!sk[34]) & (!g1748) & (g1759)) + ((g132) & (!g1706) & (g1707) & (!sk[34]) & (g1748) & (!g1759)) + ((g132) & (!g1706) & (g1707) & (!sk[34]) & (g1748) & (g1759)) + ((g132) & (!g1706) & (g1707) & (sk[34]) & (!g1748) & (g1759)) + ((g132) & (!g1706) & (g1707) & (sk[34]) & (g1748) & (g1759)) + ((g132) & (g1706) & (!g1707) & (!sk[34]) & (!g1748) & (!g1759)) + ((g132) & (g1706) & (!g1707) & (!sk[34]) & (!g1748) & (g1759)) + ((g132) & (g1706) & (!g1707) & (!sk[34]) & (g1748) & (!g1759)) + ((g132) & (g1706) & (!g1707) & (!sk[34]) & (g1748) & (g1759)) + ((g132) & (g1706) & (g1707) & (!sk[34]) & (!g1748) & (!g1759)) + ((g132) & (g1706) & (g1707) & (!sk[34]) & (!g1748) & (g1759)) + ((g132) & (g1706) & (g1707) & (!sk[34]) & (g1748) & (!g1759)) + ((g132) & (g1706) & (g1707) & (!sk[34]) & (g1748) & (g1759)));
	assign g1761 = (((!g1592) & (!sk[35]) & (!g1593) & (!g1668) & (g48)) + ((!g1592) & (!sk[35]) & (!g1593) & (g1668) & (!g48)) + ((!g1592) & (!sk[35]) & (!g1593) & (g1668) & (g48)) + ((!g1592) & (!sk[35]) & (g1593) & (!g1668) & (!g48)) + ((!g1592) & (!sk[35]) & (g1593) & (!g1668) & (g48)) + ((!g1592) & (!sk[35]) & (g1593) & (g1668) & (!g48)) + ((!g1592) & (!sk[35]) & (g1593) & (g1668) & (g48)) + ((!g1592) & (sk[35]) & (!g1593) & (g1668) & (!g48)) + ((!g1592) & (sk[35]) & (!g1593) & (g1668) & (g48)) + ((!g1592) & (sk[35]) & (g1593) & (g1668) & (!g48)) + ((!g1592) & (sk[35]) & (g1593) & (g1668) & (g48)) + ((g1592) & (!sk[35]) & (!g1593) & (!g1668) & (g48)) + ((g1592) & (!sk[35]) & (!g1593) & (g1668) & (!g48)) + ((g1592) & (!sk[35]) & (!g1593) & (g1668) & (g48)) + ((g1592) & (!sk[35]) & (g1593) & (!g1668) & (!g48)) + ((g1592) & (!sk[35]) & (g1593) & (!g1668) & (g48)) + ((g1592) & (!sk[35]) & (g1593) & (g1668) & (!g48)) + ((g1592) & (!sk[35]) & (g1593) & (g1668) & (g48)) + ((g1592) & (sk[35]) & (g1593) & (!g1668) & (g48)) + ((g1592) & (sk[35]) & (g1593) & (g1668) & (g48)));
	assign g1762 = (((!g729) & (!g730) & (!g731) & (g732) & (g820) & (g773)) + ((!g729) & (!g730) & (g731) & (!g732) & (!g820) & (g773)) + ((!g729) & (!g730) & (g731) & (g732) & (!g820) & (g773)) + ((!g729) & (!g730) & (g731) & (g732) & (g820) & (g773)) + ((!g729) & (g730) & (!g731) & (!g732) & (g820) & (!g773)) + ((!g729) & (g730) & (!g731) & (g732) & (g820) & (!g773)) + ((!g729) & (g730) & (!g731) & (g732) & (g820) & (g773)) + ((!g729) & (g730) & (g731) & (!g732) & (!g820) & (g773)) + ((!g729) & (g730) & (g731) & (!g732) & (g820) & (!g773)) + ((!g729) & (g730) & (g731) & (g732) & (!g820) & (g773)) + ((!g729) & (g730) & (g731) & (g732) & (g820) & (!g773)) + ((!g729) & (g730) & (g731) & (g732) & (g820) & (g773)) + ((g729) & (!g730) & (!g731) & (!g732) & (!g820) & (!g773)) + ((g729) & (!g730) & (!g731) & (g732) & (!g820) & (!g773)) + ((g729) & (!g730) & (!g731) & (g732) & (g820) & (g773)) + ((g729) & (!g730) & (g731) & (!g732) & (!g820) & (!g773)) + ((g729) & (!g730) & (g731) & (!g732) & (!g820) & (g773)) + ((g729) & (!g730) & (g731) & (g732) & (!g820) & (!g773)) + ((g729) & (!g730) & (g731) & (g732) & (!g820) & (g773)) + ((g729) & (!g730) & (g731) & (g732) & (g820) & (g773)) + ((g729) & (g730) & (!g731) & (!g732) & (!g820) & (!g773)) + ((g729) & (g730) & (!g731) & (!g732) & (g820) & (!g773)) + ((g729) & (g730) & (!g731) & (g732) & (!g820) & (!g773)) + ((g729) & (g730) & (!g731) & (g732) & (g820) & (!g773)) + ((g729) & (g730) & (!g731) & (g732) & (g820) & (g773)) + ((g729) & (g730) & (g731) & (!g732) & (!g820) & (!g773)) + ((g729) & (g730) & (g731) & (!g732) & (!g820) & (g773)) + ((g729) & (g730) & (g731) & (!g732) & (g820) & (!g773)) + ((g729) & (g730) & (g731) & (g732) & (!g820) & (!g773)) + ((g729) & (g730) & (g731) & (g732) & (!g820) & (g773)) + ((g729) & (g730) & (g731) & (g732) & (g820) & (!g773)) + ((g729) & (g730) & (g731) & (g732) & (g820) & (g773)));
	assign g1763 = (((!g734) & (!g735) & (!g736) & (g737) & (g820) & (g773)) + ((!g734) & (!g735) & (g736) & (!g737) & (!g820) & (g773)) + ((!g734) & (!g735) & (g736) & (g737) & (!g820) & (g773)) + ((!g734) & (!g735) & (g736) & (g737) & (g820) & (g773)) + ((!g734) & (g735) & (!g736) & (!g737) & (g820) & (!g773)) + ((!g734) & (g735) & (!g736) & (g737) & (g820) & (!g773)) + ((!g734) & (g735) & (!g736) & (g737) & (g820) & (g773)) + ((!g734) & (g735) & (g736) & (!g737) & (!g820) & (g773)) + ((!g734) & (g735) & (g736) & (!g737) & (g820) & (!g773)) + ((!g734) & (g735) & (g736) & (g737) & (!g820) & (g773)) + ((!g734) & (g735) & (g736) & (g737) & (g820) & (!g773)) + ((!g734) & (g735) & (g736) & (g737) & (g820) & (g773)) + ((g734) & (!g735) & (!g736) & (!g737) & (!g820) & (!g773)) + ((g734) & (!g735) & (!g736) & (g737) & (!g820) & (!g773)) + ((g734) & (!g735) & (!g736) & (g737) & (g820) & (g773)) + ((g734) & (!g735) & (g736) & (!g737) & (!g820) & (!g773)) + ((g734) & (!g735) & (g736) & (!g737) & (!g820) & (g773)) + ((g734) & (!g735) & (g736) & (g737) & (!g820) & (!g773)) + ((g734) & (!g735) & (g736) & (g737) & (!g820) & (g773)) + ((g734) & (!g735) & (g736) & (g737) & (g820) & (g773)) + ((g734) & (g735) & (!g736) & (!g737) & (!g820) & (!g773)) + ((g734) & (g735) & (!g736) & (!g737) & (g820) & (!g773)) + ((g734) & (g735) & (!g736) & (g737) & (!g820) & (!g773)) + ((g734) & (g735) & (!g736) & (g737) & (g820) & (!g773)) + ((g734) & (g735) & (!g736) & (g737) & (g820) & (g773)) + ((g734) & (g735) & (g736) & (!g737) & (!g820) & (!g773)) + ((g734) & (g735) & (g736) & (!g737) & (!g820) & (g773)) + ((g734) & (g735) & (g736) & (!g737) & (g820) & (!g773)) + ((g734) & (g735) & (g736) & (g737) & (!g820) & (!g773)) + ((g734) & (g735) & (g736) & (g737) & (!g820) & (g773)) + ((g734) & (g735) & (g736) & (g737) & (g820) & (!g773)) + ((g734) & (g735) & (g736) & (g737) & (g820) & (g773)));
	assign g1764 = (((!g739) & (!g740) & (!g741) & (g742) & (g820) & (g773)) + ((!g739) & (!g740) & (g741) & (!g742) & (!g820) & (g773)) + ((!g739) & (!g740) & (g741) & (g742) & (!g820) & (g773)) + ((!g739) & (!g740) & (g741) & (g742) & (g820) & (g773)) + ((!g739) & (g740) & (!g741) & (!g742) & (g820) & (!g773)) + ((!g739) & (g740) & (!g741) & (g742) & (g820) & (!g773)) + ((!g739) & (g740) & (!g741) & (g742) & (g820) & (g773)) + ((!g739) & (g740) & (g741) & (!g742) & (!g820) & (g773)) + ((!g739) & (g740) & (g741) & (!g742) & (g820) & (!g773)) + ((!g739) & (g740) & (g741) & (g742) & (!g820) & (g773)) + ((!g739) & (g740) & (g741) & (g742) & (g820) & (!g773)) + ((!g739) & (g740) & (g741) & (g742) & (g820) & (g773)) + ((g739) & (!g740) & (!g741) & (!g742) & (!g820) & (!g773)) + ((g739) & (!g740) & (!g741) & (g742) & (!g820) & (!g773)) + ((g739) & (!g740) & (!g741) & (g742) & (g820) & (g773)) + ((g739) & (!g740) & (g741) & (!g742) & (!g820) & (!g773)) + ((g739) & (!g740) & (g741) & (!g742) & (!g820) & (g773)) + ((g739) & (!g740) & (g741) & (g742) & (!g820) & (!g773)) + ((g739) & (!g740) & (g741) & (g742) & (!g820) & (g773)) + ((g739) & (!g740) & (g741) & (g742) & (g820) & (g773)) + ((g739) & (g740) & (!g741) & (!g742) & (!g820) & (!g773)) + ((g739) & (g740) & (!g741) & (!g742) & (g820) & (!g773)) + ((g739) & (g740) & (!g741) & (g742) & (!g820) & (!g773)) + ((g739) & (g740) & (!g741) & (g742) & (g820) & (!g773)) + ((g739) & (g740) & (!g741) & (g742) & (g820) & (g773)) + ((g739) & (g740) & (g741) & (!g742) & (!g820) & (!g773)) + ((g739) & (g740) & (g741) & (!g742) & (!g820) & (g773)) + ((g739) & (g740) & (g741) & (!g742) & (g820) & (!g773)) + ((g739) & (g740) & (g741) & (g742) & (!g820) & (!g773)) + ((g739) & (g740) & (g741) & (g742) & (!g820) & (g773)) + ((g739) & (g740) & (g741) & (g742) & (g820) & (!g773)) + ((g739) & (g740) & (g741) & (g742) & (g820) & (g773)));
	assign g1765 = (((!g744) & (!g745) & (!g746) & (g747) & (g820) & (g773)) + ((!g744) & (!g745) & (g746) & (!g747) & (!g820) & (g773)) + ((!g744) & (!g745) & (g746) & (g747) & (!g820) & (g773)) + ((!g744) & (!g745) & (g746) & (g747) & (g820) & (g773)) + ((!g744) & (g745) & (!g746) & (!g747) & (g820) & (!g773)) + ((!g744) & (g745) & (!g746) & (g747) & (g820) & (!g773)) + ((!g744) & (g745) & (!g746) & (g747) & (g820) & (g773)) + ((!g744) & (g745) & (g746) & (!g747) & (!g820) & (g773)) + ((!g744) & (g745) & (g746) & (!g747) & (g820) & (!g773)) + ((!g744) & (g745) & (g746) & (g747) & (!g820) & (g773)) + ((!g744) & (g745) & (g746) & (g747) & (g820) & (!g773)) + ((!g744) & (g745) & (g746) & (g747) & (g820) & (g773)) + ((g744) & (!g745) & (!g746) & (!g747) & (!g820) & (!g773)) + ((g744) & (!g745) & (!g746) & (g747) & (!g820) & (!g773)) + ((g744) & (!g745) & (!g746) & (g747) & (g820) & (g773)) + ((g744) & (!g745) & (g746) & (!g747) & (!g820) & (!g773)) + ((g744) & (!g745) & (g746) & (!g747) & (!g820) & (g773)) + ((g744) & (!g745) & (g746) & (g747) & (!g820) & (!g773)) + ((g744) & (!g745) & (g746) & (g747) & (!g820) & (g773)) + ((g744) & (!g745) & (g746) & (g747) & (g820) & (g773)) + ((g744) & (g745) & (!g746) & (!g747) & (!g820) & (!g773)) + ((g744) & (g745) & (!g746) & (!g747) & (g820) & (!g773)) + ((g744) & (g745) & (!g746) & (g747) & (!g820) & (!g773)) + ((g744) & (g745) & (!g746) & (g747) & (g820) & (!g773)) + ((g744) & (g745) & (!g746) & (g747) & (g820) & (g773)) + ((g744) & (g745) & (g746) & (!g747) & (!g820) & (!g773)) + ((g744) & (g745) & (g746) & (!g747) & (!g820) & (g773)) + ((g744) & (g745) & (g746) & (!g747) & (g820) & (!g773)) + ((g744) & (g745) & (g746) & (g747) & (!g820) & (!g773)) + ((g744) & (g745) & (g746) & (g747) & (!g820) & (g773)) + ((g744) & (g745) & (g746) & (g747) & (g820) & (!g773)) + ((g744) & (g745) & (g746) & (g747) & (g820) & (g773)));
	assign g1766 = (((!g1762) & (!g1763) & (!g1764) & (g1765) & (g677) & (g726)) + ((!g1762) & (!g1763) & (g1764) & (!g1765) & (!g677) & (g726)) + ((!g1762) & (!g1763) & (g1764) & (g1765) & (!g677) & (g726)) + ((!g1762) & (!g1763) & (g1764) & (g1765) & (g677) & (g726)) + ((!g1762) & (g1763) & (!g1764) & (!g1765) & (g677) & (!g726)) + ((!g1762) & (g1763) & (!g1764) & (g1765) & (g677) & (!g726)) + ((!g1762) & (g1763) & (!g1764) & (g1765) & (g677) & (g726)) + ((!g1762) & (g1763) & (g1764) & (!g1765) & (!g677) & (g726)) + ((!g1762) & (g1763) & (g1764) & (!g1765) & (g677) & (!g726)) + ((!g1762) & (g1763) & (g1764) & (g1765) & (!g677) & (g726)) + ((!g1762) & (g1763) & (g1764) & (g1765) & (g677) & (!g726)) + ((!g1762) & (g1763) & (g1764) & (g1765) & (g677) & (g726)) + ((g1762) & (!g1763) & (!g1764) & (!g1765) & (!g677) & (!g726)) + ((g1762) & (!g1763) & (!g1764) & (g1765) & (!g677) & (!g726)) + ((g1762) & (!g1763) & (!g1764) & (g1765) & (g677) & (g726)) + ((g1762) & (!g1763) & (g1764) & (!g1765) & (!g677) & (!g726)) + ((g1762) & (!g1763) & (g1764) & (!g1765) & (!g677) & (g726)) + ((g1762) & (!g1763) & (g1764) & (g1765) & (!g677) & (!g726)) + ((g1762) & (!g1763) & (g1764) & (g1765) & (!g677) & (g726)) + ((g1762) & (!g1763) & (g1764) & (g1765) & (g677) & (g726)) + ((g1762) & (g1763) & (!g1764) & (!g1765) & (!g677) & (!g726)) + ((g1762) & (g1763) & (!g1764) & (!g1765) & (g677) & (!g726)) + ((g1762) & (g1763) & (!g1764) & (g1765) & (!g677) & (!g726)) + ((g1762) & (g1763) & (!g1764) & (g1765) & (g677) & (!g726)) + ((g1762) & (g1763) & (!g1764) & (g1765) & (g677) & (g726)) + ((g1762) & (g1763) & (g1764) & (!g1765) & (!g677) & (!g726)) + ((g1762) & (g1763) & (g1764) & (!g1765) & (!g677) & (g726)) + ((g1762) & (g1763) & (g1764) & (!g1765) & (g677) & (!g726)) + ((g1762) & (g1763) & (g1764) & (g1765) & (!g677) & (!g726)) + ((g1762) & (g1763) & (g1764) & (g1765) & (!g677) & (g726)) + ((g1762) & (g1763) & (g1764) & (g1765) & (g677) & (!g726)) + ((g1762) & (g1763) & (g1764) & (g1765) & (g677) & (g726)));
	assign g1767 = (((!g750) & (!g751) & (!g752) & (g753) & (g677) & (g726)) + ((!g750) & (!g751) & (g752) & (!g753) & (!g677) & (g726)) + ((!g750) & (!g751) & (g752) & (g753) & (!g677) & (g726)) + ((!g750) & (!g751) & (g752) & (g753) & (g677) & (g726)) + ((!g750) & (g751) & (!g752) & (!g753) & (g677) & (!g726)) + ((!g750) & (g751) & (!g752) & (g753) & (g677) & (!g726)) + ((!g750) & (g751) & (!g752) & (g753) & (g677) & (g726)) + ((!g750) & (g751) & (g752) & (!g753) & (!g677) & (g726)) + ((!g750) & (g751) & (g752) & (!g753) & (g677) & (!g726)) + ((!g750) & (g751) & (g752) & (g753) & (!g677) & (g726)) + ((!g750) & (g751) & (g752) & (g753) & (g677) & (!g726)) + ((!g750) & (g751) & (g752) & (g753) & (g677) & (g726)) + ((g750) & (!g751) & (!g752) & (!g753) & (!g677) & (!g726)) + ((g750) & (!g751) & (!g752) & (g753) & (!g677) & (!g726)) + ((g750) & (!g751) & (!g752) & (g753) & (g677) & (g726)) + ((g750) & (!g751) & (g752) & (!g753) & (!g677) & (!g726)) + ((g750) & (!g751) & (g752) & (!g753) & (!g677) & (g726)) + ((g750) & (!g751) & (g752) & (g753) & (!g677) & (!g726)) + ((g750) & (!g751) & (g752) & (g753) & (!g677) & (g726)) + ((g750) & (!g751) & (g752) & (g753) & (g677) & (g726)) + ((g750) & (g751) & (!g752) & (!g753) & (!g677) & (!g726)) + ((g750) & (g751) & (!g752) & (!g753) & (g677) & (!g726)) + ((g750) & (g751) & (!g752) & (g753) & (!g677) & (!g726)) + ((g750) & (g751) & (!g752) & (g753) & (g677) & (!g726)) + ((g750) & (g751) & (!g752) & (g753) & (g677) & (g726)) + ((g750) & (g751) & (g752) & (!g753) & (!g677) & (!g726)) + ((g750) & (g751) & (g752) & (!g753) & (!g677) & (g726)) + ((g750) & (g751) & (g752) & (!g753) & (g677) & (!g726)) + ((g750) & (g751) & (g752) & (g753) & (!g677) & (!g726)) + ((g750) & (g751) & (g752) & (g753) & (!g677) & (g726)) + ((g750) & (g751) & (g752) & (g753) & (g677) & (!g726)) + ((g750) & (g751) & (g752) & (g753) & (g677) & (g726)));
	assign g1768 = (((!g677) & (!g726) & (!g755) & (g756) & (!sk[42]) & (!g757)) + ((!g677) & (!g726) & (!g755) & (g756) & (!sk[42]) & (g757)) + ((!g677) & (!g726) & (g755) & (!g756) & (!sk[42]) & (!g757)) + ((!g677) & (!g726) & (g755) & (!g756) & (!sk[42]) & (g757)) + ((!g677) & (!g726) & (g755) & (g756) & (!sk[42]) & (!g757)) + ((!g677) & (!g726) & (g755) & (g756) & (!sk[42]) & (g757)) + ((!g677) & (g726) & (!g755) & (!g756) & (!sk[42]) & (!g757)) + ((!g677) & (g726) & (!g755) & (!g756) & (!sk[42]) & (g757)) + ((!g677) & (g726) & (!g755) & (!g756) & (sk[42]) & (g757)) + ((!g677) & (g726) & (!g755) & (g756) & (!sk[42]) & (!g757)) + ((!g677) & (g726) & (!g755) & (g756) & (!sk[42]) & (g757)) + ((!g677) & (g726) & (!g755) & (g756) & (sk[42]) & (g757)) + ((!g677) & (g726) & (g755) & (!g756) & (!sk[42]) & (!g757)) + ((!g677) & (g726) & (g755) & (!g756) & (!sk[42]) & (g757)) + ((!g677) & (g726) & (g755) & (!g756) & (sk[42]) & (g757)) + ((!g677) & (g726) & (g755) & (g756) & (!sk[42]) & (!g757)) + ((!g677) & (g726) & (g755) & (g756) & (!sk[42]) & (g757)) + ((!g677) & (g726) & (g755) & (g756) & (sk[42]) & (g757)) + ((g677) & (!g726) & (!g755) & (g756) & (!sk[42]) & (!g757)) + ((g677) & (!g726) & (!g755) & (g756) & (!sk[42]) & (g757)) + ((g677) & (!g726) & (g755) & (!g756) & (!sk[42]) & (!g757)) + ((g677) & (!g726) & (g755) & (!g756) & (!sk[42]) & (g757)) + ((g677) & (!g726) & (g755) & (!g756) & (sk[42]) & (!g757)) + ((g677) & (!g726) & (g755) & (!g756) & (sk[42]) & (g757)) + ((g677) & (!g726) & (g755) & (g756) & (!sk[42]) & (!g757)) + ((g677) & (!g726) & (g755) & (g756) & (!sk[42]) & (g757)) + ((g677) & (!g726) & (g755) & (g756) & (sk[42]) & (!g757)) + ((g677) & (!g726) & (g755) & (g756) & (sk[42]) & (g757)) + ((g677) & (g726) & (!g755) & (!g756) & (!sk[42]) & (!g757)) + ((g677) & (g726) & (!g755) & (!g756) & (!sk[42]) & (g757)) + ((g677) & (g726) & (!g755) & (g756) & (!sk[42]) & (!g757)) + ((g677) & (g726) & (!g755) & (g756) & (!sk[42]) & (g757)) + ((g677) & (g726) & (!g755) & (g756) & (sk[42]) & (!g757)) + ((g677) & (g726) & (!g755) & (g756) & (sk[42]) & (g757)) + ((g677) & (g726) & (g755) & (!g756) & (!sk[42]) & (!g757)) + ((g677) & (g726) & (g755) & (!g756) & (!sk[42]) & (g757)) + ((g677) & (g726) & (g755) & (g756) & (!sk[42]) & (!g757)) + ((g677) & (g726) & (g755) & (g756) & (!sk[42]) & (g757)) + ((g677) & (g726) & (g755) & (g756) & (sk[42]) & (!g757)) + ((g677) & (g726) & (g755) & (g756) & (sk[42]) & (g757)));
	assign g1769 = (((!g759) & (!g760) & (!g761) & (g762) & (g677) & (g726)) + ((!g759) & (!g760) & (g761) & (!g762) & (!g677) & (g726)) + ((!g759) & (!g760) & (g761) & (g762) & (!g677) & (g726)) + ((!g759) & (!g760) & (g761) & (g762) & (g677) & (g726)) + ((!g759) & (g760) & (!g761) & (!g762) & (g677) & (!g726)) + ((!g759) & (g760) & (!g761) & (g762) & (g677) & (!g726)) + ((!g759) & (g760) & (!g761) & (g762) & (g677) & (g726)) + ((!g759) & (g760) & (g761) & (!g762) & (!g677) & (g726)) + ((!g759) & (g760) & (g761) & (!g762) & (g677) & (!g726)) + ((!g759) & (g760) & (g761) & (g762) & (!g677) & (g726)) + ((!g759) & (g760) & (g761) & (g762) & (g677) & (!g726)) + ((!g759) & (g760) & (g761) & (g762) & (g677) & (g726)) + ((g759) & (!g760) & (!g761) & (!g762) & (!g677) & (!g726)) + ((g759) & (!g760) & (!g761) & (g762) & (!g677) & (!g726)) + ((g759) & (!g760) & (!g761) & (g762) & (g677) & (g726)) + ((g759) & (!g760) & (g761) & (!g762) & (!g677) & (!g726)) + ((g759) & (!g760) & (g761) & (!g762) & (!g677) & (g726)) + ((g759) & (!g760) & (g761) & (g762) & (!g677) & (!g726)) + ((g759) & (!g760) & (g761) & (g762) & (!g677) & (g726)) + ((g759) & (!g760) & (g761) & (g762) & (g677) & (g726)) + ((g759) & (g760) & (!g761) & (!g762) & (!g677) & (!g726)) + ((g759) & (g760) & (!g761) & (!g762) & (g677) & (!g726)) + ((g759) & (g760) & (!g761) & (g762) & (!g677) & (!g726)) + ((g759) & (g760) & (!g761) & (g762) & (g677) & (!g726)) + ((g759) & (g760) & (!g761) & (g762) & (g677) & (g726)) + ((g759) & (g760) & (g761) & (!g762) & (!g677) & (!g726)) + ((g759) & (g760) & (g761) & (!g762) & (!g677) & (g726)) + ((g759) & (g760) & (g761) & (!g762) & (g677) & (!g726)) + ((g759) & (g760) & (g761) & (g762) & (!g677) & (!g726)) + ((g759) & (g760) & (g761) & (g762) & (!g677) & (g726)) + ((g759) & (g760) & (g761) & (g762) & (g677) & (!g726)) + ((g759) & (g760) & (g761) & (g762) & (g677) & (g726)));
	assign g1770 = (((!g764) & (!g765) & (!g766) & (g767) & (g677) & (g726)) + ((!g764) & (!g765) & (g766) & (!g767) & (!g677) & (g726)) + ((!g764) & (!g765) & (g766) & (g767) & (!g677) & (g726)) + ((!g764) & (!g765) & (g766) & (g767) & (g677) & (g726)) + ((!g764) & (g765) & (!g766) & (!g767) & (g677) & (!g726)) + ((!g764) & (g765) & (!g766) & (g767) & (g677) & (!g726)) + ((!g764) & (g765) & (!g766) & (g767) & (g677) & (g726)) + ((!g764) & (g765) & (g766) & (!g767) & (!g677) & (g726)) + ((!g764) & (g765) & (g766) & (!g767) & (g677) & (!g726)) + ((!g764) & (g765) & (g766) & (g767) & (!g677) & (g726)) + ((!g764) & (g765) & (g766) & (g767) & (g677) & (!g726)) + ((!g764) & (g765) & (g766) & (g767) & (g677) & (g726)) + ((g764) & (!g765) & (!g766) & (!g767) & (!g677) & (!g726)) + ((g764) & (!g765) & (!g766) & (g767) & (!g677) & (!g726)) + ((g764) & (!g765) & (!g766) & (g767) & (g677) & (g726)) + ((g764) & (!g765) & (g766) & (!g767) & (!g677) & (!g726)) + ((g764) & (!g765) & (g766) & (!g767) & (!g677) & (g726)) + ((g764) & (!g765) & (g766) & (g767) & (!g677) & (!g726)) + ((g764) & (!g765) & (g766) & (g767) & (!g677) & (g726)) + ((g764) & (!g765) & (g766) & (g767) & (g677) & (g726)) + ((g764) & (g765) & (!g766) & (!g767) & (!g677) & (!g726)) + ((g764) & (g765) & (!g766) & (!g767) & (g677) & (!g726)) + ((g764) & (g765) & (!g766) & (g767) & (!g677) & (!g726)) + ((g764) & (g765) & (!g766) & (g767) & (g677) & (!g726)) + ((g764) & (g765) & (!g766) & (g767) & (g677) & (g726)) + ((g764) & (g765) & (g766) & (!g767) & (!g677) & (!g726)) + ((g764) & (g765) & (g766) & (!g767) & (!g677) & (g726)) + ((g764) & (g765) & (g766) & (!g767) & (g677) & (!g726)) + ((g764) & (g765) & (g766) & (g767) & (!g677) & (!g726)) + ((g764) & (g765) & (g766) & (g767) & (!g677) & (g726)) + ((g764) & (g765) & (g766) & (g767) & (g677) & (!g726)) + ((g764) & (g765) & (g766) & (g767) & (g677) & (g726)));
	assign g1771 = (((!g820) & (!g773) & (!g1767) & (g1768) & (!g1769) & (!g1770)) + ((!g820) & (!g773) & (!g1767) & (g1768) & (!g1769) & (g1770)) + ((!g820) & (!g773) & (!g1767) & (g1768) & (g1769) & (!g1770)) + ((!g820) & (!g773) & (!g1767) & (g1768) & (g1769) & (g1770)) + ((!g820) & (!g773) & (g1767) & (g1768) & (!g1769) & (!g1770)) + ((!g820) & (!g773) & (g1767) & (g1768) & (!g1769) & (g1770)) + ((!g820) & (!g773) & (g1767) & (g1768) & (g1769) & (!g1770)) + ((!g820) & (!g773) & (g1767) & (g1768) & (g1769) & (g1770)) + ((!g820) & (g773) & (!g1767) & (!g1768) & (!g1769) & (g1770)) + ((!g820) & (g773) & (!g1767) & (!g1768) & (g1769) & (g1770)) + ((!g820) & (g773) & (!g1767) & (g1768) & (!g1769) & (g1770)) + ((!g820) & (g773) & (!g1767) & (g1768) & (g1769) & (g1770)) + ((!g820) & (g773) & (g1767) & (!g1768) & (!g1769) & (g1770)) + ((!g820) & (g773) & (g1767) & (!g1768) & (g1769) & (g1770)) + ((!g820) & (g773) & (g1767) & (g1768) & (!g1769) & (g1770)) + ((!g820) & (g773) & (g1767) & (g1768) & (g1769) & (g1770)) + ((g820) & (!g773) & (g1767) & (!g1768) & (!g1769) & (!g1770)) + ((g820) & (!g773) & (g1767) & (!g1768) & (!g1769) & (g1770)) + ((g820) & (!g773) & (g1767) & (!g1768) & (g1769) & (!g1770)) + ((g820) & (!g773) & (g1767) & (!g1768) & (g1769) & (g1770)) + ((g820) & (!g773) & (g1767) & (g1768) & (!g1769) & (!g1770)) + ((g820) & (!g773) & (g1767) & (g1768) & (!g1769) & (g1770)) + ((g820) & (!g773) & (g1767) & (g1768) & (g1769) & (!g1770)) + ((g820) & (!g773) & (g1767) & (g1768) & (g1769) & (g1770)) + ((g820) & (g773) & (!g1767) & (!g1768) & (g1769) & (!g1770)) + ((g820) & (g773) & (!g1767) & (!g1768) & (g1769) & (g1770)) + ((g820) & (g773) & (!g1767) & (g1768) & (g1769) & (!g1770)) + ((g820) & (g773) & (!g1767) & (g1768) & (g1769) & (g1770)) + ((g820) & (g773) & (g1767) & (!g1768) & (g1769) & (!g1770)) + ((g820) & (g773) & (g1767) & (!g1768) & (g1769) & (g1770)) + ((g820) & (g773) & (g1767) & (g1768) & (g1769) & (!g1770)) + ((g820) & (g773) & (g1767) & (g1768) & (g1769) & (g1770)));
	assign g1772 = (((!sk[46]) & (!g867) & (!g1766) & (g1771)) + ((!sk[46]) & (!g867) & (g1766) & (!g1771)) + ((!sk[46]) & (!g867) & (g1766) & (g1771)) + ((!sk[46]) & (g867) & (!g1766) & (g1771)) + ((!sk[46]) & (g867) & (g1766) & (!g1771)) + ((!sk[46]) & (g867) & (g1766) & (g1771)) + ((sk[46]) & (!g867) & (!g1766) & (g1771)) + ((sk[46]) & (!g867) & (g1766) & (g1771)) + ((sk[46]) & (g867) & (g1766) & (!g1771)) + ((sk[46]) & (g867) & (g1766) & (g1771)));
	assign g1773 = (((!g132) & (!g1706) & (!g1707) & (g1761) & (!sk[47]) & (!g1772)) + ((!g132) & (!g1706) & (!g1707) & (g1761) & (!sk[47]) & (g1772)) + ((!g132) & (!g1706) & (g1707) & (!g1761) & (!sk[47]) & (!g1772)) + ((!g132) & (!g1706) & (g1707) & (!g1761) & (!sk[47]) & (g1772)) + ((!g132) & (!g1706) & (g1707) & (!g1761) & (sk[47]) & (g1772)) + ((!g132) & (!g1706) & (g1707) & (g1761) & (!sk[47]) & (!g1772)) + ((!g132) & (!g1706) & (g1707) & (g1761) & (!sk[47]) & (g1772)) + ((!g132) & (!g1706) & (g1707) & (g1761) & (sk[47]) & (!g1772)) + ((!g132) & (!g1706) & (g1707) & (g1761) & (sk[47]) & (g1772)) + ((!g132) & (g1706) & (!g1707) & (!g1761) & (!sk[47]) & (!g1772)) + ((!g132) & (g1706) & (!g1707) & (!g1761) & (!sk[47]) & (g1772)) + ((!g132) & (g1706) & (!g1707) & (g1761) & (!sk[47]) & (!g1772)) + ((!g132) & (g1706) & (!g1707) & (g1761) & (!sk[47]) & (g1772)) + ((!g132) & (g1706) & (g1707) & (!g1761) & (!sk[47]) & (!g1772)) + ((!g132) & (g1706) & (g1707) & (!g1761) & (!sk[47]) & (g1772)) + ((!g132) & (g1706) & (g1707) & (g1761) & (!sk[47]) & (!g1772)) + ((!g132) & (g1706) & (g1707) & (g1761) & (!sk[47]) & (g1772)) + ((!g132) & (g1706) & (g1707) & (g1761) & (sk[47]) & (!g1772)) + ((!g132) & (g1706) & (g1707) & (g1761) & (sk[47]) & (g1772)) + ((g132) & (!g1706) & (!g1707) & (g1761) & (!sk[47]) & (!g1772)) + ((g132) & (!g1706) & (!g1707) & (g1761) & (!sk[47]) & (g1772)) + ((g132) & (!g1706) & (g1707) & (!g1761) & (!sk[47]) & (!g1772)) + ((g132) & (!g1706) & (g1707) & (!g1761) & (!sk[47]) & (g1772)) + ((g132) & (!g1706) & (g1707) & (!g1761) & (sk[47]) & (g1772)) + ((g132) & (!g1706) & (g1707) & (g1761) & (!sk[47]) & (!g1772)) + ((g132) & (!g1706) & (g1707) & (g1761) & (!sk[47]) & (g1772)) + ((g132) & (!g1706) & (g1707) & (g1761) & (sk[47]) & (g1772)) + ((g132) & (g1706) & (!g1707) & (!g1761) & (!sk[47]) & (!g1772)) + ((g132) & (g1706) & (!g1707) & (!g1761) & (!sk[47]) & (g1772)) + ((g132) & (g1706) & (!g1707) & (g1761) & (!sk[47]) & (!g1772)) + ((g132) & (g1706) & (!g1707) & (g1761) & (!sk[47]) & (g1772)) + ((g132) & (g1706) & (g1707) & (!g1761) & (!sk[47]) & (!g1772)) + ((g132) & (g1706) & (g1707) & (!g1761) & (!sk[47]) & (g1772)) + ((g132) & (g1706) & (g1707) & (g1761) & (!sk[47]) & (!g1772)) + ((g132) & (g1706) & (g1707) & (g1761) & (!sk[47]) & (g1772)));
	assign g1774 = (((!sk[48]) & (!g1592) & (!g1593) & (!g1680) & (g49)) + ((!sk[48]) & (!g1592) & (!g1593) & (g1680) & (!g49)) + ((!sk[48]) & (!g1592) & (!g1593) & (g1680) & (g49)) + ((!sk[48]) & (!g1592) & (g1593) & (!g1680) & (!g49)) + ((!sk[48]) & (!g1592) & (g1593) & (!g1680) & (g49)) + ((!sk[48]) & (!g1592) & (g1593) & (g1680) & (!g49)) + ((!sk[48]) & (!g1592) & (g1593) & (g1680) & (g49)) + ((!sk[48]) & (g1592) & (!g1593) & (!g1680) & (g49)) + ((!sk[48]) & (g1592) & (!g1593) & (g1680) & (!g49)) + ((!sk[48]) & (g1592) & (!g1593) & (g1680) & (g49)) + ((!sk[48]) & (g1592) & (g1593) & (!g1680) & (!g49)) + ((!sk[48]) & (g1592) & (g1593) & (!g1680) & (g49)) + ((!sk[48]) & (g1592) & (g1593) & (g1680) & (!g49)) + ((!sk[48]) & (g1592) & (g1593) & (g1680) & (g49)) + ((sk[48]) & (!g1592) & (!g1593) & (g1680) & (!g49)) + ((sk[48]) & (!g1592) & (!g1593) & (g1680) & (g49)) + ((sk[48]) & (!g1592) & (g1593) & (g1680) & (!g49)) + ((sk[48]) & (!g1592) & (g1593) & (g1680) & (g49)) + ((sk[48]) & (g1592) & (g1593) & (!g1680) & (g49)) + ((sk[48]) & (g1592) & (g1593) & (g1680) & (g49)));
	assign g1775 = (((!g776) & (!g777) & (!g778) & (g779) & (g820) & (g773)) + ((!g776) & (!g777) & (g778) & (!g779) & (!g820) & (g773)) + ((!g776) & (!g777) & (g778) & (g779) & (!g820) & (g773)) + ((!g776) & (!g777) & (g778) & (g779) & (g820) & (g773)) + ((!g776) & (g777) & (!g778) & (!g779) & (g820) & (!g773)) + ((!g776) & (g777) & (!g778) & (g779) & (g820) & (!g773)) + ((!g776) & (g777) & (!g778) & (g779) & (g820) & (g773)) + ((!g776) & (g777) & (g778) & (!g779) & (!g820) & (g773)) + ((!g776) & (g777) & (g778) & (!g779) & (g820) & (!g773)) + ((!g776) & (g777) & (g778) & (g779) & (!g820) & (g773)) + ((!g776) & (g777) & (g778) & (g779) & (g820) & (!g773)) + ((!g776) & (g777) & (g778) & (g779) & (g820) & (g773)) + ((g776) & (!g777) & (!g778) & (!g779) & (!g820) & (!g773)) + ((g776) & (!g777) & (!g778) & (g779) & (!g820) & (!g773)) + ((g776) & (!g777) & (!g778) & (g779) & (g820) & (g773)) + ((g776) & (!g777) & (g778) & (!g779) & (!g820) & (!g773)) + ((g776) & (!g777) & (g778) & (!g779) & (!g820) & (g773)) + ((g776) & (!g777) & (g778) & (g779) & (!g820) & (!g773)) + ((g776) & (!g777) & (g778) & (g779) & (!g820) & (g773)) + ((g776) & (!g777) & (g778) & (g779) & (g820) & (g773)) + ((g776) & (g777) & (!g778) & (!g779) & (!g820) & (!g773)) + ((g776) & (g777) & (!g778) & (!g779) & (g820) & (!g773)) + ((g776) & (g777) & (!g778) & (g779) & (!g820) & (!g773)) + ((g776) & (g777) & (!g778) & (g779) & (g820) & (!g773)) + ((g776) & (g777) & (!g778) & (g779) & (g820) & (g773)) + ((g776) & (g777) & (g778) & (!g779) & (!g820) & (!g773)) + ((g776) & (g777) & (g778) & (!g779) & (!g820) & (g773)) + ((g776) & (g777) & (g778) & (!g779) & (g820) & (!g773)) + ((g776) & (g777) & (g778) & (g779) & (!g820) & (!g773)) + ((g776) & (g777) & (g778) & (g779) & (!g820) & (g773)) + ((g776) & (g777) & (g778) & (g779) & (g820) & (!g773)) + ((g776) & (g777) & (g778) & (g779) & (g820) & (g773)));
	assign g1776 = (((!g781) & (!g782) & (!g783) & (g784) & (g820) & (g773)) + ((!g781) & (!g782) & (g783) & (!g784) & (!g820) & (g773)) + ((!g781) & (!g782) & (g783) & (g784) & (!g820) & (g773)) + ((!g781) & (!g782) & (g783) & (g784) & (g820) & (g773)) + ((!g781) & (g782) & (!g783) & (!g784) & (g820) & (!g773)) + ((!g781) & (g782) & (!g783) & (g784) & (g820) & (!g773)) + ((!g781) & (g782) & (!g783) & (g784) & (g820) & (g773)) + ((!g781) & (g782) & (g783) & (!g784) & (!g820) & (g773)) + ((!g781) & (g782) & (g783) & (!g784) & (g820) & (!g773)) + ((!g781) & (g782) & (g783) & (g784) & (!g820) & (g773)) + ((!g781) & (g782) & (g783) & (g784) & (g820) & (!g773)) + ((!g781) & (g782) & (g783) & (g784) & (g820) & (g773)) + ((g781) & (!g782) & (!g783) & (!g784) & (!g820) & (!g773)) + ((g781) & (!g782) & (!g783) & (g784) & (!g820) & (!g773)) + ((g781) & (!g782) & (!g783) & (g784) & (g820) & (g773)) + ((g781) & (!g782) & (g783) & (!g784) & (!g820) & (!g773)) + ((g781) & (!g782) & (g783) & (!g784) & (!g820) & (g773)) + ((g781) & (!g782) & (g783) & (g784) & (!g820) & (!g773)) + ((g781) & (!g782) & (g783) & (g784) & (!g820) & (g773)) + ((g781) & (!g782) & (g783) & (g784) & (g820) & (g773)) + ((g781) & (g782) & (!g783) & (!g784) & (!g820) & (!g773)) + ((g781) & (g782) & (!g783) & (!g784) & (g820) & (!g773)) + ((g781) & (g782) & (!g783) & (g784) & (!g820) & (!g773)) + ((g781) & (g782) & (!g783) & (g784) & (g820) & (!g773)) + ((g781) & (g782) & (!g783) & (g784) & (g820) & (g773)) + ((g781) & (g782) & (g783) & (!g784) & (!g820) & (!g773)) + ((g781) & (g782) & (g783) & (!g784) & (!g820) & (g773)) + ((g781) & (g782) & (g783) & (!g784) & (g820) & (!g773)) + ((g781) & (g782) & (g783) & (g784) & (!g820) & (!g773)) + ((g781) & (g782) & (g783) & (g784) & (!g820) & (g773)) + ((g781) & (g782) & (g783) & (g784) & (g820) & (!g773)) + ((g781) & (g782) & (g783) & (g784) & (g820) & (g773)));
	assign g1777 = (((!g786) & (!g787) & (!g788) & (g789) & (g820) & (g773)) + ((!g786) & (!g787) & (g788) & (!g789) & (!g820) & (g773)) + ((!g786) & (!g787) & (g788) & (g789) & (!g820) & (g773)) + ((!g786) & (!g787) & (g788) & (g789) & (g820) & (g773)) + ((!g786) & (g787) & (!g788) & (!g789) & (g820) & (!g773)) + ((!g786) & (g787) & (!g788) & (g789) & (g820) & (!g773)) + ((!g786) & (g787) & (!g788) & (g789) & (g820) & (g773)) + ((!g786) & (g787) & (g788) & (!g789) & (!g820) & (g773)) + ((!g786) & (g787) & (g788) & (!g789) & (g820) & (!g773)) + ((!g786) & (g787) & (g788) & (g789) & (!g820) & (g773)) + ((!g786) & (g787) & (g788) & (g789) & (g820) & (!g773)) + ((!g786) & (g787) & (g788) & (g789) & (g820) & (g773)) + ((g786) & (!g787) & (!g788) & (!g789) & (!g820) & (!g773)) + ((g786) & (!g787) & (!g788) & (g789) & (!g820) & (!g773)) + ((g786) & (!g787) & (!g788) & (g789) & (g820) & (g773)) + ((g786) & (!g787) & (g788) & (!g789) & (!g820) & (!g773)) + ((g786) & (!g787) & (g788) & (!g789) & (!g820) & (g773)) + ((g786) & (!g787) & (g788) & (g789) & (!g820) & (!g773)) + ((g786) & (!g787) & (g788) & (g789) & (!g820) & (g773)) + ((g786) & (!g787) & (g788) & (g789) & (g820) & (g773)) + ((g786) & (g787) & (!g788) & (!g789) & (!g820) & (!g773)) + ((g786) & (g787) & (!g788) & (!g789) & (g820) & (!g773)) + ((g786) & (g787) & (!g788) & (g789) & (!g820) & (!g773)) + ((g786) & (g787) & (!g788) & (g789) & (g820) & (!g773)) + ((g786) & (g787) & (!g788) & (g789) & (g820) & (g773)) + ((g786) & (g787) & (g788) & (!g789) & (!g820) & (!g773)) + ((g786) & (g787) & (g788) & (!g789) & (!g820) & (g773)) + ((g786) & (g787) & (g788) & (!g789) & (g820) & (!g773)) + ((g786) & (g787) & (g788) & (g789) & (!g820) & (!g773)) + ((g786) & (g787) & (g788) & (g789) & (!g820) & (g773)) + ((g786) & (g787) & (g788) & (g789) & (g820) & (!g773)) + ((g786) & (g787) & (g788) & (g789) & (g820) & (g773)));
	assign g1778 = (((!g791) & (!g792) & (!g793) & (g794) & (g820) & (g773)) + ((!g791) & (!g792) & (g793) & (!g794) & (!g820) & (g773)) + ((!g791) & (!g792) & (g793) & (g794) & (!g820) & (g773)) + ((!g791) & (!g792) & (g793) & (g794) & (g820) & (g773)) + ((!g791) & (g792) & (!g793) & (!g794) & (g820) & (!g773)) + ((!g791) & (g792) & (!g793) & (g794) & (g820) & (!g773)) + ((!g791) & (g792) & (!g793) & (g794) & (g820) & (g773)) + ((!g791) & (g792) & (g793) & (!g794) & (!g820) & (g773)) + ((!g791) & (g792) & (g793) & (!g794) & (g820) & (!g773)) + ((!g791) & (g792) & (g793) & (g794) & (!g820) & (g773)) + ((!g791) & (g792) & (g793) & (g794) & (g820) & (!g773)) + ((!g791) & (g792) & (g793) & (g794) & (g820) & (g773)) + ((g791) & (!g792) & (!g793) & (!g794) & (!g820) & (!g773)) + ((g791) & (!g792) & (!g793) & (g794) & (!g820) & (!g773)) + ((g791) & (!g792) & (!g793) & (g794) & (g820) & (g773)) + ((g791) & (!g792) & (g793) & (!g794) & (!g820) & (!g773)) + ((g791) & (!g792) & (g793) & (!g794) & (!g820) & (g773)) + ((g791) & (!g792) & (g793) & (g794) & (!g820) & (!g773)) + ((g791) & (!g792) & (g793) & (g794) & (!g820) & (g773)) + ((g791) & (!g792) & (g793) & (g794) & (g820) & (g773)) + ((g791) & (g792) & (!g793) & (!g794) & (!g820) & (!g773)) + ((g791) & (g792) & (!g793) & (!g794) & (g820) & (!g773)) + ((g791) & (g792) & (!g793) & (g794) & (!g820) & (!g773)) + ((g791) & (g792) & (!g793) & (g794) & (g820) & (!g773)) + ((g791) & (g792) & (!g793) & (g794) & (g820) & (g773)) + ((g791) & (g792) & (g793) & (!g794) & (!g820) & (!g773)) + ((g791) & (g792) & (g793) & (!g794) & (!g820) & (g773)) + ((g791) & (g792) & (g793) & (!g794) & (g820) & (!g773)) + ((g791) & (g792) & (g793) & (g794) & (!g820) & (!g773)) + ((g791) & (g792) & (g793) & (g794) & (!g820) & (g773)) + ((g791) & (g792) & (g793) & (g794) & (g820) & (!g773)) + ((g791) & (g792) & (g793) & (g794) & (g820) & (g773)));
	assign g1779 = (((!g1775) & (!g1776) & (!g1777) & (g1778) & (g677) & (g726)) + ((!g1775) & (!g1776) & (g1777) & (!g1778) & (!g677) & (g726)) + ((!g1775) & (!g1776) & (g1777) & (g1778) & (!g677) & (g726)) + ((!g1775) & (!g1776) & (g1777) & (g1778) & (g677) & (g726)) + ((!g1775) & (g1776) & (!g1777) & (!g1778) & (g677) & (!g726)) + ((!g1775) & (g1776) & (!g1777) & (g1778) & (g677) & (!g726)) + ((!g1775) & (g1776) & (!g1777) & (g1778) & (g677) & (g726)) + ((!g1775) & (g1776) & (g1777) & (!g1778) & (!g677) & (g726)) + ((!g1775) & (g1776) & (g1777) & (!g1778) & (g677) & (!g726)) + ((!g1775) & (g1776) & (g1777) & (g1778) & (!g677) & (g726)) + ((!g1775) & (g1776) & (g1777) & (g1778) & (g677) & (!g726)) + ((!g1775) & (g1776) & (g1777) & (g1778) & (g677) & (g726)) + ((g1775) & (!g1776) & (!g1777) & (!g1778) & (!g677) & (!g726)) + ((g1775) & (!g1776) & (!g1777) & (g1778) & (!g677) & (!g726)) + ((g1775) & (!g1776) & (!g1777) & (g1778) & (g677) & (g726)) + ((g1775) & (!g1776) & (g1777) & (!g1778) & (!g677) & (!g726)) + ((g1775) & (!g1776) & (g1777) & (!g1778) & (!g677) & (g726)) + ((g1775) & (!g1776) & (g1777) & (g1778) & (!g677) & (!g726)) + ((g1775) & (!g1776) & (g1777) & (g1778) & (!g677) & (g726)) + ((g1775) & (!g1776) & (g1777) & (g1778) & (g677) & (g726)) + ((g1775) & (g1776) & (!g1777) & (!g1778) & (!g677) & (!g726)) + ((g1775) & (g1776) & (!g1777) & (!g1778) & (g677) & (!g726)) + ((g1775) & (g1776) & (!g1777) & (g1778) & (!g677) & (!g726)) + ((g1775) & (g1776) & (!g1777) & (g1778) & (g677) & (!g726)) + ((g1775) & (g1776) & (!g1777) & (g1778) & (g677) & (g726)) + ((g1775) & (g1776) & (g1777) & (!g1778) & (!g677) & (!g726)) + ((g1775) & (g1776) & (g1777) & (!g1778) & (!g677) & (g726)) + ((g1775) & (g1776) & (g1777) & (!g1778) & (g677) & (!g726)) + ((g1775) & (g1776) & (g1777) & (g1778) & (!g677) & (!g726)) + ((g1775) & (g1776) & (g1777) & (g1778) & (!g677) & (g726)) + ((g1775) & (g1776) & (g1777) & (g1778) & (g677) & (!g726)) + ((g1775) & (g1776) & (g1777) & (g1778) & (g677) & (g726)));
	assign g1780 = (((!g797) & (!g798) & (!g799) & (g800) & (g677) & (g726)) + ((!g797) & (!g798) & (g799) & (!g800) & (!g677) & (g726)) + ((!g797) & (!g798) & (g799) & (g800) & (!g677) & (g726)) + ((!g797) & (!g798) & (g799) & (g800) & (g677) & (g726)) + ((!g797) & (g798) & (!g799) & (!g800) & (g677) & (!g726)) + ((!g797) & (g798) & (!g799) & (g800) & (g677) & (!g726)) + ((!g797) & (g798) & (!g799) & (g800) & (g677) & (g726)) + ((!g797) & (g798) & (g799) & (!g800) & (!g677) & (g726)) + ((!g797) & (g798) & (g799) & (!g800) & (g677) & (!g726)) + ((!g797) & (g798) & (g799) & (g800) & (!g677) & (g726)) + ((!g797) & (g798) & (g799) & (g800) & (g677) & (!g726)) + ((!g797) & (g798) & (g799) & (g800) & (g677) & (g726)) + ((g797) & (!g798) & (!g799) & (!g800) & (!g677) & (!g726)) + ((g797) & (!g798) & (!g799) & (g800) & (!g677) & (!g726)) + ((g797) & (!g798) & (!g799) & (g800) & (g677) & (g726)) + ((g797) & (!g798) & (g799) & (!g800) & (!g677) & (!g726)) + ((g797) & (!g798) & (g799) & (!g800) & (!g677) & (g726)) + ((g797) & (!g798) & (g799) & (g800) & (!g677) & (!g726)) + ((g797) & (!g798) & (g799) & (g800) & (!g677) & (g726)) + ((g797) & (!g798) & (g799) & (g800) & (g677) & (g726)) + ((g797) & (g798) & (!g799) & (!g800) & (!g677) & (!g726)) + ((g797) & (g798) & (!g799) & (!g800) & (g677) & (!g726)) + ((g797) & (g798) & (!g799) & (g800) & (!g677) & (!g726)) + ((g797) & (g798) & (!g799) & (g800) & (g677) & (!g726)) + ((g797) & (g798) & (!g799) & (g800) & (g677) & (g726)) + ((g797) & (g798) & (g799) & (!g800) & (!g677) & (!g726)) + ((g797) & (g798) & (g799) & (!g800) & (!g677) & (g726)) + ((g797) & (g798) & (g799) & (!g800) & (g677) & (!g726)) + ((g797) & (g798) & (g799) & (g800) & (!g677) & (!g726)) + ((g797) & (g798) & (g799) & (g800) & (!g677) & (g726)) + ((g797) & (g798) & (g799) & (g800) & (g677) & (!g726)) + ((g797) & (g798) & (g799) & (g800) & (g677) & (g726)));
	assign g1781 = (((!g677) & (!g726) & (!g802) & (g803) & (!sk[55]) & (!g804)) + ((!g677) & (!g726) & (!g802) & (g803) & (!sk[55]) & (g804)) + ((!g677) & (!g726) & (g802) & (!g803) & (!sk[55]) & (!g804)) + ((!g677) & (!g726) & (g802) & (!g803) & (!sk[55]) & (g804)) + ((!g677) & (!g726) & (g802) & (g803) & (!sk[55]) & (!g804)) + ((!g677) & (!g726) & (g802) & (g803) & (!sk[55]) & (g804)) + ((!g677) & (g726) & (!g802) & (!g803) & (!sk[55]) & (!g804)) + ((!g677) & (g726) & (!g802) & (!g803) & (!sk[55]) & (g804)) + ((!g677) & (g726) & (!g802) & (!g803) & (sk[55]) & (g804)) + ((!g677) & (g726) & (!g802) & (g803) & (!sk[55]) & (!g804)) + ((!g677) & (g726) & (!g802) & (g803) & (!sk[55]) & (g804)) + ((!g677) & (g726) & (!g802) & (g803) & (sk[55]) & (g804)) + ((!g677) & (g726) & (g802) & (!g803) & (!sk[55]) & (!g804)) + ((!g677) & (g726) & (g802) & (!g803) & (!sk[55]) & (g804)) + ((!g677) & (g726) & (g802) & (!g803) & (sk[55]) & (g804)) + ((!g677) & (g726) & (g802) & (g803) & (!sk[55]) & (!g804)) + ((!g677) & (g726) & (g802) & (g803) & (!sk[55]) & (g804)) + ((!g677) & (g726) & (g802) & (g803) & (sk[55]) & (g804)) + ((g677) & (!g726) & (!g802) & (g803) & (!sk[55]) & (!g804)) + ((g677) & (!g726) & (!g802) & (g803) & (!sk[55]) & (g804)) + ((g677) & (!g726) & (g802) & (!g803) & (!sk[55]) & (!g804)) + ((g677) & (!g726) & (g802) & (!g803) & (!sk[55]) & (g804)) + ((g677) & (!g726) & (g802) & (!g803) & (sk[55]) & (!g804)) + ((g677) & (!g726) & (g802) & (!g803) & (sk[55]) & (g804)) + ((g677) & (!g726) & (g802) & (g803) & (!sk[55]) & (!g804)) + ((g677) & (!g726) & (g802) & (g803) & (!sk[55]) & (g804)) + ((g677) & (!g726) & (g802) & (g803) & (sk[55]) & (!g804)) + ((g677) & (!g726) & (g802) & (g803) & (sk[55]) & (g804)) + ((g677) & (g726) & (!g802) & (!g803) & (!sk[55]) & (!g804)) + ((g677) & (g726) & (!g802) & (!g803) & (!sk[55]) & (g804)) + ((g677) & (g726) & (!g802) & (g803) & (!sk[55]) & (!g804)) + ((g677) & (g726) & (!g802) & (g803) & (!sk[55]) & (g804)) + ((g677) & (g726) & (!g802) & (g803) & (sk[55]) & (!g804)) + ((g677) & (g726) & (!g802) & (g803) & (sk[55]) & (g804)) + ((g677) & (g726) & (g802) & (!g803) & (!sk[55]) & (!g804)) + ((g677) & (g726) & (g802) & (!g803) & (!sk[55]) & (g804)) + ((g677) & (g726) & (g802) & (g803) & (!sk[55]) & (!g804)) + ((g677) & (g726) & (g802) & (g803) & (!sk[55]) & (g804)) + ((g677) & (g726) & (g802) & (g803) & (sk[55]) & (!g804)) + ((g677) & (g726) & (g802) & (g803) & (sk[55]) & (g804)));
	assign g1782 = (((!g806) & (!g807) & (!g808) & (g809) & (g677) & (g726)) + ((!g806) & (!g807) & (g808) & (!g809) & (!g677) & (g726)) + ((!g806) & (!g807) & (g808) & (g809) & (!g677) & (g726)) + ((!g806) & (!g807) & (g808) & (g809) & (g677) & (g726)) + ((!g806) & (g807) & (!g808) & (!g809) & (g677) & (!g726)) + ((!g806) & (g807) & (!g808) & (g809) & (g677) & (!g726)) + ((!g806) & (g807) & (!g808) & (g809) & (g677) & (g726)) + ((!g806) & (g807) & (g808) & (!g809) & (!g677) & (g726)) + ((!g806) & (g807) & (g808) & (!g809) & (g677) & (!g726)) + ((!g806) & (g807) & (g808) & (g809) & (!g677) & (g726)) + ((!g806) & (g807) & (g808) & (g809) & (g677) & (!g726)) + ((!g806) & (g807) & (g808) & (g809) & (g677) & (g726)) + ((g806) & (!g807) & (!g808) & (!g809) & (!g677) & (!g726)) + ((g806) & (!g807) & (!g808) & (g809) & (!g677) & (!g726)) + ((g806) & (!g807) & (!g808) & (g809) & (g677) & (g726)) + ((g806) & (!g807) & (g808) & (!g809) & (!g677) & (!g726)) + ((g806) & (!g807) & (g808) & (!g809) & (!g677) & (g726)) + ((g806) & (!g807) & (g808) & (g809) & (!g677) & (!g726)) + ((g806) & (!g807) & (g808) & (g809) & (!g677) & (g726)) + ((g806) & (!g807) & (g808) & (g809) & (g677) & (g726)) + ((g806) & (g807) & (!g808) & (!g809) & (!g677) & (!g726)) + ((g806) & (g807) & (!g808) & (!g809) & (g677) & (!g726)) + ((g806) & (g807) & (!g808) & (g809) & (!g677) & (!g726)) + ((g806) & (g807) & (!g808) & (g809) & (g677) & (!g726)) + ((g806) & (g807) & (!g808) & (g809) & (g677) & (g726)) + ((g806) & (g807) & (g808) & (!g809) & (!g677) & (!g726)) + ((g806) & (g807) & (g808) & (!g809) & (!g677) & (g726)) + ((g806) & (g807) & (g808) & (!g809) & (g677) & (!g726)) + ((g806) & (g807) & (g808) & (g809) & (!g677) & (!g726)) + ((g806) & (g807) & (g808) & (g809) & (!g677) & (g726)) + ((g806) & (g807) & (g808) & (g809) & (g677) & (!g726)) + ((g806) & (g807) & (g808) & (g809) & (g677) & (g726)));
	assign g1783 = (((!g811) & (!g812) & (!g813) & (g814) & (g677) & (g726)) + ((!g811) & (!g812) & (g813) & (!g814) & (!g677) & (g726)) + ((!g811) & (!g812) & (g813) & (g814) & (!g677) & (g726)) + ((!g811) & (!g812) & (g813) & (g814) & (g677) & (g726)) + ((!g811) & (g812) & (!g813) & (!g814) & (g677) & (!g726)) + ((!g811) & (g812) & (!g813) & (g814) & (g677) & (!g726)) + ((!g811) & (g812) & (!g813) & (g814) & (g677) & (g726)) + ((!g811) & (g812) & (g813) & (!g814) & (!g677) & (g726)) + ((!g811) & (g812) & (g813) & (!g814) & (g677) & (!g726)) + ((!g811) & (g812) & (g813) & (g814) & (!g677) & (g726)) + ((!g811) & (g812) & (g813) & (g814) & (g677) & (!g726)) + ((!g811) & (g812) & (g813) & (g814) & (g677) & (g726)) + ((g811) & (!g812) & (!g813) & (!g814) & (!g677) & (!g726)) + ((g811) & (!g812) & (!g813) & (g814) & (!g677) & (!g726)) + ((g811) & (!g812) & (!g813) & (g814) & (g677) & (g726)) + ((g811) & (!g812) & (g813) & (!g814) & (!g677) & (!g726)) + ((g811) & (!g812) & (g813) & (!g814) & (!g677) & (g726)) + ((g811) & (!g812) & (g813) & (g814) & (!g677) & (!g726)) + ((g811) & (!g812) & (g813) & (g814) & (!g677) & (g726)) + ((g811) & (!g812) & (g813) & (g814) & (g677) & (g726)) + ((g811) & (g812) & (!g813) & (!g814) & (!g677) & (!g726)) + ((g811) & (g812) & (!g813) & (!g814) & (g677) & (!g726)) + ((g811) & (g812) & (!g813) & (g814) & (!g677) & (!g726)) + ((g811) & (g812) & (!g813) & (g814) & (g677) & (!g726)) + ((g811) & (g812) & (!g813) & (g814) & (g677) & (g726)) + ((g811) & (g812) & (g813) & (!g814) & (!g677) & (!g726)) + ((g811) & (g812) & (g813) & (!g814) & (!g677) & (g726)) + ((g811) & (g812) & (g813) & (!g814) & (g677) & (!g726)) + ((g811) & (g812) & (g813) & (g814) & (!g677) & (!g726)) + ((g811) & (g812) & (g813) & (g814) & (!g677) & (g726)) + ((g811) & (g812) & (g813) & (g814) & (g677) & (!g726)) + ((g811) & (g812) & (g813) & (g814) & (g677) & (g726)));
	assign g1784 = (((!g820) & (!g773) & (!g1780) & (g1781) & (!g1782) & (!g1783)) + ((!g820) & (!g773) & (!g1780) & (g1781) & (!g1782) & (g1783)) + ((!g820) & (!g773) & (!g1780) & (g1781) & (g1782) & (!g1783)) + ((!g820) & (!g773) & (!g1780) & (g1781) & (g1782) & (g1783)) + ((!g820) & (!g773) & (g1780) & (g1781) & (!g1782) & (!g1783)) + ((!g820) & (!g773) & (g1780) & (g1781) & (!g1782) & (g1783)) + ((!g820) & (!g773) & (g1780) & (g1781) & (g1782) & (!g1783)) + ((!g820) & (!g773) & (g1780) & (g1781) & (g1782) & (g1783)) + ((!g820) & (g773) & (!g1780) & (!g1781) & (!g1782) & (g1783)) + ((!g820) & (g773) & (!g1780) & (!g1781) & (g1782) & (g1783)) + ((!g820) & (g773) & (!g1780) & (g1781) & (!g1782) & (g1783)) + ((!g820) & (g773) & (!g1780) & (g1781) & (g1782) & (g1783)) + ((!g820) & (g773) & (g1780) & (!g1781) & (!g1782) & (g1783)) + ((!g820) & (g773) & (g1780) & (!g1781) & (g1782) & (g1783)) + ((!g820) & (g773) & (g1780) & (g1781) & (!g1782) & (g1783)) + ((!g820) & (g773) & (g1780) & (g1781) & (g1782) & (g1783)) + ((g820) & (!g773) & (g1780) & (!g1781) & (!g1782) & (!g1783)) + ((g820) & (!g773) & (g1780) & (!g1781) & (!g1782) & (g1783)) + ((g820) & (!g773) & (g1780) & (!g1781) & (g1782) & (!g1783)) + ((g820) & (!g773) & (g1780) & (!g1781) & (g1782) & (g1783)) + ((g820) & (!g773) & (g1780) & (g1781) & (!g1782) & (!g1783)) + ((g820) & (!g773) & (g1780) & (g1781) & (!g1782) & (g1783)) + ((g820) & (!g773) & (g1780) & (g1781) & (g1782) & (!g1783)) + ((g820) & (!g773) & (g1780) & (g1781) & (g1782) & (g1783)) + ((g820) & (g773) & (!g1780) & (!g1781) & (g1782) & (!g1783)) + ((g820) & (g773) & (!g1780) & (!g1781) & (g1782) & (g1783)) + ((g820) & (g773) & (!g1780) & (g1781) & (g1782) & (!g1783)) + ((g820) & (g773) & (!g1780) & (g1781) & (g1782) & (g1783)) + ((g820) & (g773) & (g1780) & (!g1781) & (g1782) & (!g1783)) + ((g820) & (g773) & (g1780) & (!g1781) & (g1782) & (g1783)) + ((g820) & (g773) & (g1780) & (g1781) & (g1782) & (!g1783)) + ((g820) & (g773) & (g1780) & (g1781) & (g1782) & (g1783)));
	assign g1785 = (((!sk[59]) & (!g867) & (!g1779) & (g1784)) + ((!sk[59]) & (!g867) & (g1779) & (!g1784)) + ((!sk[59]) & (!g867) & (g1779) & (g1784)) + ((!sk[59]) & (g867) & (!g1779) & (g1784)) + ((!sk[59]) & (g867) & (g1779) & (!g1784)) + ((!sk[59]) & (g867) & (g1779) & (g1784)) + ((sk[59]) & (!g867) & (!g1779) & (g1784)) + ((sk[59]) & (!g867) & (g1779) & (g1784)) + ((sk[59]) & (g867) & (g1779) & (!g1784)) + ((sk[59]) & (g867) & (g1779) & (g1784)));
	assign g1786 = (((!sk[60]) & (!g132) & (!g1706) & (!g1707) & (g1774) & (!g1785)) + ((!sk[60]) & (!g132) & (!g1706) & (!g1707) & (g1774) & (g1785)) + ((!sk[60]) & (!g132) & (!g1706) & (g1707) & (!g1774) & (!g1785)) + ((!sk[60]) & (!g132) & (!g1706) & (g1707) & (!g1774) & (g1785)) + ((!sk[60]) & (!g132) & (!g1706) & (g1707) & (g1774) & (!g1785)) + ((!sk[60]) & (!g132) & (!g1706) & (g1707) & (g1774) & (g1785)) + ((!sk[60]) & (!g132) & (g1706) & (!g1707) & (!g1774) & (!g1785)) + ((!sk[60]) & (!g132) & (g1706) & (!g1707) & (!g1774) & (g1785)) + ((!sk[60]) & (!g132) & (g1706) & (!g1707) & (g1774) & (!g1785)) + ((!sk[60]) & (!g132) & (g1706) & (!g1707) & (g1774) & (g1785)) + ((!sk[60]) & (!g132) & (g1706) & (g1707) & (!g1774) & (!g1785)) + ((!sk[60]) & (!g132) & (g1706) & (g1707) & (!g1774) & (g1785)) + ((!sk[60]) & (!g132) & (g1706) & (g1707) & (g1774) & (!g1785)) + ((!sk[60]) & (!g132) & (g1706) & (g1707) & (g1774) & (g1785)) + ((!sk[60]) & (g132) & (!g1706) & (!g1707) & (g1774) & (!g1785)) + ((!sk[60]) & (g132) & (!g1706) & (!g1707) & (g1774) & (g1785)) + ((!sk[60]) & (g132) & (!g1706) & (g1707) & (!g1774) & (!g1785)) + ((!sk[60]) & (g132) & (!g1706) & (g1707) & (!g1774) & (g1785)) + ((!sk[60]) & (g132) & (!g1706) & (g1707) & (g1774) & (!g1785)) + ((!sk[60]) & (g132) & (!g1706) & (g1707) & (g1774) & (g1785)) + ((!sk[60]) & (g132) & (g1706) & (!g1707) & (!g1774) & (!g1785)) + ((!sk[60]) & (g132) & (g1706) & (!g1707) & (!g1774) & (g1785)) + ((!sk[60]) & (g132) & (g1706) & (!g1707) & (g1774) & (!g1785)) + ((!sk[60]) & (g132) & (g1706) & (!g1707) & (g1774) & (g1785)) + ((!sk[60]) & (g132) & (g1706) & (g1707) & (!g1774) & (!g1785)) + ((!sk[60]) & (g132) & (g1706) & (g1707) & (!g1774) & (g1785)) + ((!sk[60]) & (g132) & (g1706) & (g1707) & (g1774) & (!g1785)) + ((!sk[60]) & (g132) & (g1706) & (g1707) & (g1774) & (g1785)) + ((sk[60]) & (!g132) & (!g1706) & (g1707) & (!g1774) & (g1785)) + ((sk[60]) & (!g132) & (!g1706) & (g1707) & (g1774) & (!g1785)) + ((sk[60]) & (!g132) & (!g1706) & (g1707) & (g1774) & (g1785)) + ((sk[60]) & (!g132) & (g1706) & (g1707) & (g1774) & (!g1785)) + ((sk[60]) & (!g132) & (g1706) & (g1707) & (g1774) & (g1785)) + ((sk[60]) & (g132) & (!g1706) & (g1707) & (!g1774) & (g1785)) + ((sk[60]) & (g132) & (!g1706) & (g1707) & (g1774) & (g1785)));
	assign g1787 = (((!g1592) & (!sk[61]) & (!g1593) & (!g1692) & (g50)) + ((!g1592) & (!sk[61]) & (!g1593) & (g1692) & (!g50)) + ((!g1592) & (!sk[61]) & (!g1593) & (g1692) & (g50)) + ((!g1592) & (!sk[61]) & (g1593) & (!g1692) & (!g50)) + ((!g1592) & (!sk[61]) & (g1593) & (!g1692) & (g50)) + ((!g1592) & (!sk[61]) & (g1593) & (g1692) & (!g50)) + ((!g1592) & (!sk[61]) & (g1593) & (g1692) & (g50)) + ((!g1592) & (sk[61]) & (!g1593) & (g1692) & (!g50)) + ((!g1592) & (sk[61]) & (!g1593) & (g1692) & (g50)) + ((!g1592) & (sk[61]) & (g1593) & (g1692) & (!g50)) + ((!g1592) & (sk[61]) & (g1593) & (g1692) & (g50)) + ((g1592) & (!sk[61]) & (!g1593) & (!g1692) & (g50)) + ((g1592) & (!sk[61]) & (!g1593) & (g1692) & (!g50)) + ((g1592) & (!sk[61]) & (!g1593) & (g1692) & (g50)) + ((g1592) & (!sk[61]) & (g1593) & (!g1692) & (!g50)) + ((g1592) & (!sk[61]) & (g1593) & (!g1692) & (g50)) + ((g1592) & (!sk[61]) & (g1593) & (g1692) & (!g50)) + ((g1592) & (!sk[61]) & (g1593) & (g1692) & (g50)) + ((g1592) & (sk[61]) & (g1593) & (!g1692) & (g50)) + ((g1592) & (sk[61]) & (g1593) & (g1692) & (g50)));
	assign g1788 = (((!g823) & (!g824) & (!g825) & (g826) & (g820) & (g773)) + ((!g823) & (!g824) & (g825) & (!g826) & (!g820) & (g773)) + ((!g823) & (!g824) & (g825) & (g826) & (!g820) & (g773)) + ((!g823) & (!g824) & (g825) & (g826) & (g820) & (g773)) + ((!g823) & (g824) & (!g825) & (!g826) & (g820) & (!g773)) + ((!g823) & (g824) & (!g825) & (g826) & (g820) & (!g773)) + ((!g823) & (g824) & (!g825) & (g826) & (g820) & (g773)) + ((!g823) & (g824) & (g825) & (!g826) & (!g820) & (g773)) + ((!g823) & (g824) & (g825) & (!g826) & (g820) & (!g773)) + ((!g823) & (g824) & (g825) & (g826) & (!g820) & (g773)) + ((!g823) & (g824) & (g825) & (g826) & (g820) & (!g773)) + ((!g823) & (g824) & (g825) & (g826) & (g820) & (g773)) + ((g823) & (!g824) & (!g825) & (!g826) & (!g820) & (!g773)) + ((g823) & (!g824) & (!g825) & (g826) & (!g820) & (!g773)) + ((g823) & (!g824) & (!g825) & (g826) & (g820) & (g773)) + ((g823) & (!g824) & (g825) & (!g826) & (!g820) & (!g773)) + ((g823) & (!g824) & (g825) & (!g826) & (!g820) & (g773)) + ((g823) & (!g824) & (g825) & (g826) & (!g820) & (!g773)) + ((g823) & (!g824) & (g825) & (g826) & (!g820) & (g773)) + ((g823) & (!g824) & (g825) & (g826) & (g820) & (g773)) + ((g823) & (g824) & (!g825) & (!g826) & (!g820) & (!g773)) + ((g823) & (g824) & (!g825) & (!g826) & (g820) & (!g773)) + ((g823) & (g824) & (!g825) & (g826) & (!g820) & (!g773)) + ((g823) & (g824) & (!g825) & (g826) & (g820) & (!g773)) + ((g823) & (g824) & (!g825) & (g826) & (g820) & (g773)) + ((g823) & (g824) & (g825) & (!g826) & (!g820) & (!g773)) + ((g823) & (g824) & (g825) & (!g826) & (!g820) & (g773)) + ((g823) & (g824) & (g825) & (!g826) & (g820) & (!g773)) + ((g823) & (g824) & (g825) & (g826) & (!g820) & (!g773)) + ((g823) & (g824) & (g825) & (g826) & (!g820) & (g773)) + ((g823) & (g824) & (g825) & (g826) & (g820) & (!g773)) + ((g823) & (g824) & (g825) & (g826) & (g820) & (g773)));
	assign g1789 = (((!g828) & (!g829) & (!g830) & (g831) & (g820) & (g773)) + ((!g828) & (!g829) & (g830) & (!g831) & (!g820) & (g773)) + ((!g828) & (!g829) & (g830) & (g831) & (!g820) & (g773)) + ((!g828) & (!g829) & (g830) & (g831) & (g820) & (g773)) + ((!g828) & (g829) & (!g830) & (!g831) & (g820) & (!g773)) + ((!g828) & (g829) & (!g830) & (g831) & (g820) & (!g773)) + ((!g828) & (g829) & (!g830) & (g831) & (g820) & (g773)) + ((!g828) & (g829) & (g830) & (!g831) & (!g820) & (g773)) + ((!g828) & (g829) & (g830) & (!g831) & (g820) & (!g773)) + ((!g828) & (g829) & (g830) & (g831) & (!g820) & (g773)) + ((!g828) & (g829) & (g830) & (g831) & (g820) & (!g773)) + ((!g828) & (g829) & (g830) & (g831) & (g820) & (g773)) + ((g828) & (!g829) & (!g830) & (!g831) & (!g820) & (!g773)) + ((g828) & (!g829) & (!g830) & (g831) & (!g820) & (!g773)) + ((g828) & (!g829) & (!g830) & (g831) & (g820) & (g773)) + ((g828) & (!g829) & (g830) & (!g831) & (!g820) & (!g773)) + ((g828) & (!g829) & (g830) & (!g831) & (!g820) & (g773)) + ((g828) & (!g829) & (g830) & (g831) & (!g820) & (!g773)) + ((g828) & (!g829) & (g830) & (g831) & (!g820) & (g773)) + ((g828) & (!g829) & (g830) & (g831) & (g820) & (g773)) + ((g828) & (g829) & (!g830) & (!g831) & (!g820) & (!g773)) + ((g828) & (g829) & (!g830) & (!g831) & (g820) & (!g773)) + ((g828) & (g829) & (!g830) & (g831) & (!g820) & (!g773)) + ((g828) & (g829) & (!g830) & (g831) & (g820) & (!g773)) + ((g828) & (g829) & (!g830) & (g831) & (g820) & (g773)) + ((g828) & (g829) & (g830) & (!g831) & (!g820) & (!g773)) + ((g828) & (g829) & (g830) & (!g831) & (!g820) & (g773)) + ((g828) & (g829) & (g830) & (!g831) & (g820) & (!g773)) + ((g828) & (g829) & (g830) & (g831) & (!g820) & (!g773)) + ((g828) & (g829) & (g830) & (g831) & (!g820) & (g773)) + ((g828) & (g829) & (g830) & (g831) & (g820) & (!g773)) + ((g828) & (g829) & (g830) & (g831) & (g820) & (g773)));
	assign g1790 = (((!g833) & (!g834) & (!g835) & (g836) & (g820) & (g773)) + ((!g833) & (!g834) & (g835) & (!g836) & (!g820) & (g773)) + ((!g833) & (!g834) & (g835) & (g836) & (!g820) & (g773)) + ((!g833) & (!g834) & (g835) & (g836) & (g820) & (g773)) + ((!g833) & (g834) & (!g835) & (!g836) & (g820) & (!g773)) + ((!g833) & (g834) & (!g835) & (g836) & (g820) & (!g773)) + ((!g833) & (g834) & (!g835) & (g836) & (g820) & (g773)) + ((!g833) & (g834) & (g835) & (!g836) & (!g820) & (g773)) + ((!g833) & (g834) & (g835) & (!g836) & (g820) & (!g773)) + ((!g833) & (g834) & (g835) & (g836) & (!g820) & (g773)) + ((!g833) & (g834) & (g835) & (g836) & (g820) & (!g773)) + ((!g833) & (g834) & (g835) & (g836) & (g820) & (g773)) + ((g833) & (!g834) & (!g835) & (!g836) & (!g820) & (!g773)) + ((g833) & (!g834) & (!g835) & (g836) & (!g820) & (!g773)) + ((g833) & (!g834) & (!g835) & (g836) & (g820) & (g773)) + ((g833) & (!g834) & (g835) & (!g836) & (!g820) & (!g773)) + ((g833) & (!g834) & (g835) & (!g836) & (!g820) & (g773)) + ((g833) & (!g834) & (g835) & (g836) & (!g820) & (!g773)) + ((g833) & (!g834) & (g835) & (g836) & (!g820) & (g773)) + ((g833) & (!g834) & (g835) & (g836) & (g820) & (g773)) + ((g833) & (g834) & (!g835) & (!g836) & (!g820) & (!g773)) + ((g833) & (g834) & (!g835) & (!g836) & (g820) & (!g773)) + ((g833) & (g834) & (!g835) & (g836) & (!g820) & (!g773)) + ((g833) & (g834) & (!g835) & (g836) & (g820) & (!g773)) + ((g833) & (g834) & (!g835) & (g836) & (g820) & (g773)) + ((g833) & (g834) & (g835) & (!g836) & (!g820) & (!g773)) + ((g833) & (g834) & (g835) & (!g836) & (!g820) & (g773)) + ((g833) & (g834) & (g835) & (!g836) & (g820) & (!g773)) + ((g833) & (g834) & (g835) & (g836) & (!g820) & (!g773)) + ((g833) & (g834) & (g835) & (g836) & (!g820) & (g773)) + ((g833) & (g834) & (g835) & (g836) & (g820) & (!g773)) + ((g833) & (g834) & (g835) & (g836) & (g820) & (g773)));
	assign g1791 = (((!g838) & (!g839) & (!g840) & (g841) & (g820) & (g773)) + ((!g838) & (!g839) & (g840) & (!g841) & (!g820) & (g773)) + ((!g838) & (!g839) & (g840) & (g841) & (!g820) & (g773)) + ((!g838) & (!g839) & (g840) & (g841) & (g820) & (g773)) + ((!g838) & (g839) & (!g840) & (!g841) & (g820) & (!g773)) + ((!g838) & (g839) & (!g840) & (g841) & (g820) & (!g773)) + ((!g838) & (g839) & (!g840) & (g841) & (g820) & (g773)) + ((!g838) & (g839) & (g840) & (!g841) & (!g820) & (g773)) + ((!g838) & (g839) & (g840) & (!g841) & (g820) & (!g773)) + ((!g838) & (g839) & (g840) & (g841) & (!g820) & (g773)) + ((!g838) & (g839) & (g840) & (g841) & (g820) & (!g773)) + ((!g838) & (g839) & (g840) & (g841) & (g820) & (g773)) + ((g838) & (!g839) & (!g840) & (!g841) & (!g820) & (!g773)) + ((g838) & (!g839) & (!g840) & (g841) & (!g820) & (!g773)) + ((g838) & (!g839) & (!g840) & (g841) & (g820) & (g773)) + ((g838) & (!g839) & (g840) & (!g841) & (!g820) & (!g773)) + ((g838) & (!g839) & (g840) & (!g841) & (!g820) & (g773)) + ((g838) & (!g839) & (g840) & (g841) & (!g820) & (!g773)) + ((g838) & (!g839) & (g840) & (g841) & (!g820) & (g773)) + ((g838) & (!g839) & (g840) & (g841) & (g820) & (g773)) + ((g838) & (g839) & (!g840) & (!g841) & (!g820) & (!g773)) + ((g838) & (g839) & (!g840) & (!g841) & (g820) & (!g773)) + ((g838) & (g839) & (!g840) & (g841) & (!g820) & (!g773)) + ((g838) & (g839) & (!g840) & (g841) & (g820) & (!g773)) + ((g838) & (g839) & (!g840) & (g841) & (g820) & (g773)) + ((g838) & (g839) & (g840) & (!g841) & (!g820) & (!g773)) + ((g838) & (g839) & (g840) & (!g841) & (!g820) & (g773)) + ((g838) & (g839) & (g840) & (!g841) & (g820) & (!g773)) + ((g838) & (g839) & (g840) & (g841) & (!g820) & (!g773)) + ((g838) & (g839) & (g840) & (g841) & (!g820) & (g773)) + ((g838) & (g839) & (g840) & (g841) & (g820) & (!g773)) + ((g838) & (g839) & (g840) & (g841) & (g820) & (g773)));
	assign g1792 = (((!g1788) & (!g1789) & (!g1790) & (g1791) & (g677) & (g726)) + ((!g1788) & (!g1789) & (g1790) & (!g1791) & (!g677) & (g726)) + ((!g1788) & (!g1789) & (g1790) & (g1791) & (!g677) & (g726)) + ((!g1788) & (!g1789) & (g1790) & (g1791) & (g677) & (g726)) + ((!g1788) & (g1789) & (!g1790) & (!g1791) & (g677) & (!g726)) + ((!g1788) & (g1789) & (!g1790) & (g1791) & (g677) & (!g726)) + ((!g1788) & (g1789) & (!g1790) & (g1791) & (g677) & (g726)) + ((!g1788) & (g1789) & (g1790) & (!g1791) & (!g677) & (g726)) + ((!g1788) & (g1789) & (g1790) & (!g1791) & (g677) & (!g726)) + ((!g1788) & (g1789) & (g1790) & (g1791) & (!g677) & (g726)) + ((!g1788) & (g1789) & (g1790) & (g1791) & (g677) & (!g726)) + ((!g1788) & (g1789) & (g1790) & (g1791) & (g677) & (g726)) + ((g1788) & (!g1789) & (!g1790) & (!g1791) & (!g677) & (!g726)) + ((g1788) & (!g1789) & (!g1790) & (g1791) & (!g677) & (!g726)) + ((g1788) & (!g1789) & (!g1790) & (g1791) & (g677) & (g726)) + ((g1788) & (!g1789) & (g1790) & (!g1791) & (!g677) & (!g726)) + ((g1788) & (!g1789) & (g1790) & (!g1791) & (!g677) & (g726)) + ((g1788) & (!g1789) & (g1790) & (g1791) & (!g677) & (!g726)) + ((g1788) & (!g1789) & (g1790) & (g1791) & (!g677) & (g726)) + ((g1788) & (!g1789) & (g1790) & (g1791) & (g677) & (g726)) + ((g1788) & (g1789) & (!g1790) & (!g1791) & (!g677) & (!g726)) + ((g1788) & (g1789) & (!g1790) & (!g1791) & (g677) & (!g726)) + ((g1788) & (g1789) & (!g1790) & (g1791) & (!g677) & (!g726)) + ((g1788) & (g1789) & (!g1790) & (g1791) & (g677) & (!g726)) + ((g1788) & (g1789) & (!g1790) & (g1791) & (g677) & (g726)) + ((g1788) & (g1789) & (g1790) & (!g1791) & (!g677) & (!g726)) + ((g1788) & (g1789) & (g1790) & (!g1791) & (!g677) & (g726)) + ((g1788) & (g1789) & (g1790) & (!g1791) & (g677) & (!g726)) + ((g1788) & (g1789) & (g1790) & (g1791) & (!g677) & (!g726)) + ((g1788) & (g1789) & (g1790) & (g1791) & (!g677) & (g726)) + ((g1788) & (g1789) & (g1790) & (g1791) & (g677) & (!g726)) + ((g1788) & (g1789) & (g1790) & (g1791) & (g677) & (g726)));
	assign g1793 = (((!g844) & (!g845) & (!g846) & (g847) & (g677) & (g726)) + ((!g844) & (!g845) & (g846) & (!g847) & (!g677) & (g726)) + ((!g844) & (!g845) & (g846) & (g847) & (!g677) & (g726)) + ((!g844) & (!g845) & (g846) & (g847) & (g677) & (g726)) + ((!g844) & (g845) & (!g846) & (!g847) & (g677) & (!g726)) + ((!g844) & (g845) & (!g846) & (g847) & (g677) & (!g726)) + ((!g844) & (g845) & (!g846) & (g847) & (g677) & (g726)) + ((!g844) & (g845) & (g846) & (!g847) & (!g677) & (g726)) + ((!g844) & (g845) & (g846) & (!g847) & (g677) & (!g726)) + ((!g844) & (g845) & (g846) & (g847) & (!g677) & (g726)) + ((!g844) & (g845) & (g846) & (g847) & (g677) & (!g726)) + ((!g844) & (g845) & (g846) & (g847) & (g677) & (g726)) + ((g844) & (!g845) & (!g846) & (!g847) & (!g677) & (!g726)) + ((g844) & (!g845) & (!g846) & (g847) & (!g677) & (!g726)) + ((g844) & (!g845) & (!g846) & (g847) & (g677) & (g726)) + ((g844) & (!g845) & (g846) & (!g847) & (!g677) & (!g726)) + ((g844) & (!g845) & (g846) & (!g847) & (!g677) & (g726)) + ((g844) & (!g845) & (g846) & (g847) & (!g677) & (!g726)) + ((g844) & (!g845) & (g846) & (g847) & (!g677) & (g726)) + ((g844) & (!g845) & (g846) & (g847) & (g677) & (g726)) + ((g844) & (g845) & (!g846) & (!g847) & (!g677) & (!g726)) + ((g844) & (g845) & (!g846) & (!g847) & (g677) & (!g726)) + ((g844) & (g845) & (!g846) & (g847) & (!g677) & (!g726)) + ((g844) & (g845) & (!g846) & (g847) & (g677) & (!g726)) + ((g844) & (g845) & (!g846) & (g847) & (g677) & (g726)) + ((g844) & (g845) & (g846) & (!g847) & (!g677) & (!g726)) + ((g844) & (g845) & (g846) & (!g847) & (!g677) & (g726)) + ((g844) & (g845) & (g846) & (!g847) & (g677) & (!g726)) + ((g844) & (g845) & (g846) & (g847) & (!g677) & (!g726)) + ((g844) & (g845) & (g846) & (g847) & (!g677) & (g726)) + ((g844) & (g845) & (g846) & (g847) & (g677) & (!g726)) + ((g844) & (g845) & (g846) & (g847) & (g677) & (g726)));
	assign g1794 = (((!g677) & (!g726) & (!sk[68]) & (!g849) & (g850) & (!g851)) + ((!g677) & (!g726) & (!sk[68]) & (!g849) & (g850) & (g851)) + ((!g677) & (!g726) & (!sk[68]) & (g849) & (!g850) & (!g851)) + ((!g677) & (!g726) & (!sk[68]) & (g849) & (!g850) & (g851)) + ((!g677) & (!g726) & (!sk[68]) & (g849) & (g850) & (!g851)) + ((!g677) & (!g726) & (!sk[68]) & (g849) & (g850) & (g851)) + ((!g677) & (g726) & (!sk[68]) & (!g849) & (!g850) & (!g851)) + ((!g677) & (g726) & (!sk[68]) & (!g849) & (!g850) & (g851)) + ((!g677) & (g726) & (!sk[68]) & (!g849) & (g850) & (!g851)) + ((!g677) & (g726) & (!sk[68]) & (!g849) & (g850) & (g851)) + ((!g677) & (g726) & (!sk[68]) & (g849) & (!g850) & (!g851)) + ((!g677) & (g726) & (!sk[68]) & (g849) & (!g850) & (g851)) + ((!g677) & (g726) & (!sk[68]) & (g849) & (g850) & (!g851)) + ((!g677) & (g726) & (!sk[68]) & (g849) & (g850) & (g851)) + ((!g677) & (g726) & (sk[68]) & (!g849) & (!g850) & (g851)) + ((!g677) & (g726) & (sk[68]) & (!g849) & (g850) & (g851)) + ((!g677) & (g726) & (sk[68]) & (g849) & (!g850) & (g851)) + ((!g677) & (g726) & (sk[68]) & (g849) & (g850) & (g851)) + ((g677) & (!g726) & (!sk[68]) & (!g849) & (g850) & (!g851)) + ((g677) & (!g726) & (!sk[68]) & (!g849) & (g850) & (g851)) + ((g677) & (!g726) & (!sk[68]) & (g849) & (!g850) & (!g851)) + ((g677) & (!g726) & (!sk[68]) & (g849) & (!g850) & (g851)) + ((g677) & (!g726) & (!sk[68]) & (g849) & (g850) & (!g851)) + ((g677) & (!g726) & (!sk[68]) & (g849) & (g850) & (g851)) + ((g677) & (!g726) & (sk[68]) & (g849) & (!g850) & (!g851)) + ((g677) & (!g726) & (sk[68]) & (g849) & (!g850) & (g851)) + ((g677) & (!g726) & (sk[68]) & (g849) & (g850) & (!g851)) + ((g677) & (!g726) & (sk[68]) & (g849) & (g850) & (g851)) + ((g677) & (g726) & (!sk[68]) & (!g849) & (!g850) & (!g851)) + ((g677) & (g726) & (!sk[68]) & (!g849) & (!g850) & (g851)) + ((g677) & (g726) & (!sk[68]) & (!g849) & (g850) & (!g851)) + ((g677) & (g726) & (!sk[68]) & (!g849) & (g850) & (g851)) + ((g677) & (g726) & (!sk[68]) & (g849) & (!g850) & (!g851)) + ((g677) & (g726) & (!sk[68]) & (g849) & (!g850) & (g851)) + ((g677) & (g726) & (!sk[68]) & (g849) & (g850) & (!g851)) + ((g677) & (g726) & (!sk[68]) & (g849) & (g850) & (g851)) + ((g677) & (g726) & (sk[68]) & (!g849) & (g850) & (!g851)) + ((g677) & (g726) & (sk[68]) & (!g849) & (g850) & (g851)) + ((g677) & (g726) & (sk[68]) & (g849) & (g850) & (!g851)) + ((g677) & (g726) & (sk[68]) & (g849) & (g850) & (g851)));
	assign g1795 = (((!g853) & (!g854) & (!g855) & (g856) & (g677) & (g726)) + ((!g853) & (!g854) & (g855) & (!g856) & (!g677) & (g726)) + ((!g853) & (!g854) & (g855) & (g856) & (!g677) & (g726)) + ((!g853) & (!g854) & (g855) & (g856) & (g677) & (g726)) + ((!g853) & (g854) & (!g855) & (!g856) & (g677) & (!g726)) + ((!g853) & (g854) & (!g855) & (g856) & (g677) & (!g726)) + ((!g853) & (g854) & (!g855) & (g856) & (g677) & (g726)) + ((!g853) & (g854) & (g855) & (!g856) & (!g677) & (g726)) + ((!g853) & (g854) & (g855) & (!g856) & (g677) & (!g726)) + ((!g853) & (g854) & (g855) & (g856) & (!g677) & (g726)) + ((!g853) & (g854) & (g855) & (g856) & (g677) & (!g726)) + ((!g853) & (g854) & (g855) & (g856) & (g677) & (g726)) + ((g853) & (!g854) & (!g855) & (!g856) & (!g677) & (!g726)) + ((g853) & (!g854) & (!g855) & (g856) & (!g677) & (!g726)) + ((g853) & (!g854) & (!g855) & (g856) & (g677) & (g726)) + ((g853) & (!g854) & (g855) & (!g856) & (!g677) & (!g726)) + ((g853) & (!g854) & (g855) & (!g856) & (!g677) & (g726)) + ((g853) & (!g854) & (g855) & (g856) & (!g677) & (!g726)) + ((g853) & (!g854) & (g855) & (g856) & (!g677) & (g726)) + ((g853) & (!g854) & (g855) & (g856) & (g677) & (g726)) + ((g853) & (g854) & (!g855) & (!g856) & (!g677) & (!g726)) + ((g853) & (g854) & (!g855) & (!g856) & (g677) & (!g726)) + ((g853) & (g854) & (!g855) & (g856) & (!g677) & (!g726)) + ((g853) & (g854) & (!g855) & (g856) & (g677) & (!g726)) + ((g853) & (g854) & (!g855) & (g856) & (g677) & (g726)) + ((g853) & (g854) & (g855) & (!g856) & (!g677) & (!g726)) + ((g853) & (g854) & (g855) & (!g856) & (!g677) & (g726)) + ((g853) & (g854) & (g855) & (!g856) & (g677) & (!g726)) + ((g853) & (g854) & (g855) & (g856) & (!g677) & (!g726)) + ((g853) & (g854) & (g855) & (g856) & (!g677) & (g726)) + ((g853) & (g854) & (g855) & (g856) & (g677) & (!g726)) + ((g853) & (g854) & (g855) & (g856) & (g677) & (g726)));
	assign g1796 = (((!g858) & (!g859) & (!g860) & (g861) & (g677) & (g726)) + ((!g858) & (!g859) & (g860) & (!g861) & (!g677) & (g726)) + ((!g858) & (!g859) & (g860) & (g861) & (!g677) & (g726)) + ((!g858) & (!g859) & (g860) & (g861) & (g677) & (g726)) + ((!g858) & (g859) & (!g860) & (!g861) & (g677) & (!g726)) + ((!g858) & (g859) & (!g860) & (g861) & (g677) & (!g726)) + ((!g858) & (g859) & (!g860) & (g861) & (g677) & (g726)) + ((!g858) & (g859) & (g860) & (!g861) & (!g677) & (g726)) + ((!g858) & (g859) & (g860) & (!g861) & (g677) & (!g726)) + ((!g858) & (g859) & (g860) & (g861) & (!g677) & (g726)) + ((!g858) & (g859) & (g860) & (g861) & (g677) & (!g726)) + ((!g858) & (g859) & (g860) & (g861) & (g677) & (g726)) + ((g858) & (!g859) & (!g860) & (!g861) & (!g677) & (!g726)) + ((g858) & (!g859) & (!g860) & (g861) & (!g677) & (!g726)) + ((g858) & (!g859) & (!g860) & (g861) & (g677) & (g726)) + ((g858) & (!g859) & (g860) & (!g861) & (!g677) & (!g726)) + ((g858) & (!g859) & (g860) & (!g861) & (!g677) & (g726)) + ((g858) & (!g859) & (g860) & (g861) & (!g677) & (!g726)) + ((g858) & (!g859) & (g860) & (g861) & (!g677) & (g726)) + ((g858) & (!g859) & (g860) & (g861) & (g677) & (g726)) + ((g858) & (g859) & (!g860) & (!g861) & (!g677) & (!g726)) + ((g858) & (g859) & (!g860) & (!g861) & (g677) & (!g726)) + ((g858) & (g859) & (!g860) & (g861) & (!g677) & (!g726)) + ((g858) & (g859) & (!g860) & (g861) & (g677) & (!g726)) + ((g858) & (g859) & (!g860) & (g861) & (g677) & (g726)) + ((g858) & (g859) & (g860) & (!g861) & (!g677) & (!g726)) + ((g858) & (g859) & (g860) & (!g861) & (!g677) & (g726)) + ((g858) & (g859) & (g860) & (!g861) & (g677) & (!g726)) + ((g858) & (g859) & (g860) & (g861) & (!g677) & (!g726)) + ((g858) & (g859) & (g860) & (g861) & (!g677) & (g726)) + ((g858) & (g859) & (g860) & (g861) & (g677) & (!g726)) + ((g858) & (g859) & (g860) & (g861) & (g677) & (g726)));
	assign g1797 = (((!g820) & (!g773) & (!g1793) & (g1794) & (!g1795) & (!g1796)) + ((!g820) & (!g773) & (!g1793) & (g1794) & (!g1795) & (g1796)) + ((!g820) & (!g773) & (!g1793) & (g1794) & (g1795) & (!g1796)) + ((!g820) & (!g773) & (!g1793) & (g1794) & (g1795) & (g1796)) + ((!g820) & (!g773) & (g1793) & (g1794) & (!g1795) & (!g1796)) + ((!g820) & (!g773) & (g1793) & (g1794) & (!g1795) & (g1796)) + ((!g820) & (!g773) & (g1793) & (g1794) & (g1795) & (!g1796)) + ((!g820) & (!g773) & (g1793) & (g1794) & (g1795) & (g1796)) + ((!g820) & (g773) & (!g1793) & (!g1794) & (!g1795) & (g1796)) + ((!g820) & (g773) & (!g1793) & (!g1794) & (g1795) & (g1796)) + ((!g820) & (g773) & (!g1793) & (g1794) & (!g1795) & (g1796)) + ((!g820) & (g773) & (!g1793) & (g1794) & (g1795) & (g1796)) + ((!g820) & (g773) & (g1793) & (!g1794) & (!g1795) & (g1796)) + ((!g820) & (g773) & (g1793) & (!g1794) & (g1795) & (g1796)) + ((!g820) & (g773) & (g1793) & (g1794) & (!g1795) & (g1796)) + ((!g820) & (g773) & (g1793) & (g1794) & (g1795) & (g1796)) + ((g820) & (!g773) & (g1793) & (!g1794) & (!g1795) & (!g1796)) + ((g820) & (!g773) & (g1793) & (!g1794) & (!g1795) & (g1796)) + ((g820) & (!g773) & (g1793) & (!g1794) & (g1795) & (!g1796)) + ((g820) & (!g773) & (g1793) & (!g1794) & (g1795) & (g1796)) + ((g820) & (!g773) & (g1793) & (g1794) & (!g1795) & (!g1796)) + ((g820) & (!g773) & (g1793) & (g1794) & (!g1795) & (g1796)) + ((g820) & (!g773) & (g1793) & (g1794) & (g1795) & (!g1796)) + ((g820) & (!g773) & (g1793) & (g1794) & (g1795) & (g1796)) + ((g820) & (g773) & (!g1793) & (!g1794) & (g1795) & (!g1796)) + ((g820) & (g773) & (!g1793) & (!g1794) & (g1795) & (g1796)) + ((g820) & (g773) & (!g1793) & (g1794) & (g1795) & (!g1796)) + ((g820) & (g773) & (!g1793) & (g1794) & (g1795) & (g1796)) + ((g820) & (g773) & (g1793) & (!g1794) & (g1795) & (!g1796)) + ((g820) & (g773) & (g1793) & (!g1794) & (g1795) & (g1796)) + ((g820) & (g773) & (g1793) & (g1794) & (g1795) & (!g1796)) + ((g820) & (g773) & (g1793) & (g1794) & (g1795) & (g1796)));
	assign g1798 = (((!g867) & (!g1792) & (!sk[72]) & (g1797)) + ((!g867) & (!g1792) & (sk[72]) & (g1797)) + ((!g867) & (g1792) & (!sk[72]) & (!g1797)) + ((!g867) & (g1792) & (!sk[72]) & (g1797)) + ((!g867) & (g1792) & (sk[72]) & (g1797)) + ((g867) & (!g1792) & (!sk[72]) & (g1797)) + ((g867) & (g1792) & (!sk[72]) & (!g1797)) + ((g867) & (g1792) & (!sk[72]) & (g1797)) + ((g867) & (g1792) & (sk[72]) & (!g1797)) + ((g867) & (g1792) & (sk[72]) & (g1797)));
	assign g1799 = (((!g132) & (!g1706) & (!g1707) & (!sk[73]) & (g1787) & (!g1798)) + ((!g132) & (!g1706) & (!g1707) & (!sk[73]) & (g1787) & (g1798)) + ((!g132) & (!g1706) & (g1707) & (!sk[73]) & (!g1787) & (!g1798)) + ((!g132) & (!g1706) & (g1707) & (!sk[73]) & (!g1787) & (g1798)) + ((!g132) & (!g1706) & (g1707) & (!sk[73]) & (g1787) & (!g1798)) + ((!g132) & (!g1706) & (g1707) & (!sk[73]) & (g1787) & (g1798)) + ((!g132) & (!g1706) & (g1707) & (sk[73]) & (!g1787) & (g1798)) + ((!g132) & (!g1706) & (g1707) & (sk[73]) & (g1787) & (!g1798)) + ((!g132) & (!g1706) & (g1707) & (sk[73]) & (g1787) & (g1798)) + ((!g132) & (g1706) & (!g1707) & (!sk[73]) & (!g1787) & (!g1798)) + ((!g132) & (g1706) & (!g1707) & (!sk[73]) & (!g1787) & (g1798)) + ((!g132) & (g1706) & (!g1707) & (!sk[73]) & (g1787) & (!g1798)) + ((!g132) & (g1706) & (!g1707) & (!sk[73]) & (g1787) & (g1798)) + ((!g132) & (g1706) & (g1707) & (!sk[73]) & (!g1787) & (!g1798)) + ((!g132) & (g1706) & (g1707) & (!sk[73]) & (!g1787) & (g1798)) + ((!g132) & (g1706) & (g1707) & (!sk[73]) & (g1787) & (!g1798)) + ((!g132) & (g1706) & (g1707) & (!sk[73]) & (g1787) & (g1798)) + ((!g132) & (g1706) & (g1707) & (sk[73]) & (g1787) & (!g1798)) + ((!g132) & (g1706) & (g1707) & (sk[73]) & (g1787) & (g1798)) + ((g132) & (!g1706) & (!g1707) & (!sk[73]) & (g1787) & (!g1798)) + ((g132) & (!g1706) & (!g1707) & (!sk[73]) & (g1787) & (g1798)) + ((g132) & (!g1706) & (g1707) & (!sk[73]) & (!g1787) & (!g1798)) + ((g132) & (!g1706) & (g1707) & (!sk[73]) & (!g1787) & (g1798)) + ((g132) & (!g1706) & (g1707) & (!sk[73]) & (g1787) & (!g1798)) + ((g132) & (!g1706) & (g1707) & (!sk[73]) & (g1787) & (g1798)) + ((g132) & (!g1706) & (g1707) & (sk[73]) & (!g1787) & (g1798)) + ((g132) & (!g1706) & (g1707) & (sk[73]) & (g1787) & (g1798)) + ((g132) & (g1706) & (!g1707) & (!sk[73]) & (!g1787) & (!g1798)) + ((g132) & (g1706) & (!g1707) & (!sk[73]) & (!g1787) & (g1798)) + ((g132) & (g1706) & (!g1707) & (!sk[73]) & (g1787) & (!g1798)) + ((g132) & (g1706) & (!g1707) & (!sk[73]) & (g1787) & (g1798)) + ((g132) & (g1706) & (g1707) & (!sk[73]) & (!g1787) & (!g1798)) + ((g132) & (g1706) & (g1707) & (!sk[73]) & (!g1787) & (g1798)) + ((g132) & (g1706) & (g1707) & (!sk[73]) & (g1787) & (!g1798)) + ((g132) & (g1706) & (g1707) & (!sk[73]) & (g1787) & (g1798)));
	assign g1800 = (((!g870) & (!g871) & (!g872) & (g873) & (g820) & (g773)) + ((!g870) & (!g871) & (g872) & (!g873) & (!g820) & (g773)) + ((!g870) & (!g871) & (g872) & (g873) & (!g820) & (g773)) + ((!g870) & (!g871) & (g872) & (g873) & (g820) & (g773)) + ((!g870) & (g871) & (!g872) & (!g873) & (g820) & (!g773)) + ((!g870) & (g871) & (!g872) & (g873) & (g820) & (!g773)) + ((!g870) & (g871) & (!g872) & (g873) & (g820) & (g773)) + ((!g870) & (g871) & (g872) & (!g873) & (!g820) & (g773)) + ((!g870) & (g871) & (g872) & (!g873) & (g820) & (!g773)) + ((!g870) & (g871) & (g872) & (g873) & (!g820) & (g773)) + ((!g870) & (g871) & (g872) & (g873) & (g820) & (!g773)) + ((!g870) & (g871) & (g872) & (g873) & (g820) & (g773)) + ((g870) & (!g871) & (!g872) & (!g873) & (!g820) & (!g773)) + ((g870) & (!g871) & (!g872) & (g873) & (!g820) & (!g773)) + ((g870) & (!g871) & (!g872) & (g873) & (g820) & (g773)) + ((g870) & (!g871) & (g872) & (!g873) & (!g820) & (!g773)) + ((g870) & (!g871) & (g872) & (!g873) & (!g820) & (g773)) + ((g870) & (!g871) & (g872) & (g873) & (!g820) & (!g773)) + ((g870) & (!g871) & (g872) & (g873) & (!g820) & (g773)) + ((g870) & (!g871) & (g872) & (g873) & (g820) & (g773)) + ((g870) & (g871) & (!g872) & (!g873) & (!g820) & (!g773)) + ((g870) & (g871) & (!g872) & (!g873) & (g820) & (!g773)) + ((g870) & (g871) & (!g872) & (g873) & (!g820) & (!g773)) + ((g870) & (g871) & (!g872) & (g873) & (g820) & (!g773)) + ((g870) & (g871) & (!g872) & (g873) & (g820) & (g773)) + ((g870) & (g871) & (g872) & (!g873) & (!g820) & (!g773)) + ((g870) & (g871) & (g872) & (!g873) & (!g820) & (g773)) + ((g870) & (g871) & (g872) & (!g873) & (g820) & (!g773)) + ((g870) & (g871) & (g872) & (g873) & (!g820) & (!g773)) + ((g870) & (g871) & (g872) & (g873) & (!g820) & (g773)) + ((g870) & (g871) & (g872) & (g873) & (g820) & (!g773)) + ((g870) & (g871) & (g872) & (g873) & (g820) & (g773)));
	assign g1801 = (((!g875) & (!g876) & (!g877) & (g878) & (g820) & (g773)) + ((!g875) & (!g876) & (g877) & (!g878) & (!g820) & (g773)) + ((!g875) & (!g876) & (g877) & (g878) & (!g820) & (g773)) + ((!g875) & (!g876) & (g877) & (g878) & (g820) & (g773)) + ((!g875) & (g876) & (!g877) & (!g878) & (g820) & (!g773)) + ((!g875) & (g876) & (!g877) & (g878) & (g820) & (!g773)) + ((!g875) & (g876) & (!g877) & (g878) & (g820) & (g773)) + ((!g875) & (g876) & (g877) & (!g878) & (!g820) & (g773)) + ((!g875) & (g876) & (g877) & (!g878) & (g820) & (!g773)) + ((!g875) & (g876) & (g877) & (g878) & (!g820) & (g773)) + ((!g875) & (g876) & (g877) & (g878) & (g820) & (!g773)) + ((!g875) & (g876) & (g877) & (g878) & (g820) & (g773)) + ((g875) & (!g876) & (!g877) & (!g878) & (!g820) & (!g773)) + ((g875) & (!g876) & (!g877) & (g878) & (!g820) & (!g773)) + ((g875) & (!g876) & (!g877) & (g878) & (g820) & (g773)) + ((g875) & (!g876) & (g877) & (!g878) & (!g820) & (!g773)) + ((g875) & (!g876) & (g877) & (!g878) & (!g820) & (g773)) + ((g875) & (!g876) & (g877) & (g878) & (!g820) & (!g773)) + ((g875) & (!g876) & (g877) & (g878) & (!g820) & (g773)) + ((g875) & (!g876) & (g877) & (g878) & (g820) & (g773)) + ((g875) & (g876) & (!g877) & (!g878) & (!g820) & (!g773)) + ((g875) & (g876) & (!g877) & (!g878) & (g820) & (!g773)) + ((g875) & (g876) & (!g877) & (g878) & (!g820) & (!g773)) + ((g875) & (g876) & (!g877) & (g878) & (g820) & (!g773)) + ((g875) & (g876) & (!g877) & (g878) & (g820) & (g773)) + ((g875) & (g876) & (g877) & (!g878) & (!g820) & (!g773)) + ((g875) & (g876) & (g877) & (!g878) & (!g820) & (g773)) + ((g875) & (g876) & (g877) & (!g878) & (g820) & (!g773)) + ((g875) & (g876) & (g877) & (g878) & (!g820) & (!g773)) + ((g875) & (g876) & (g877) & (g878) & (!g820) & (g773)) + ((g875) & (g876) & (g877) & (g878) & (g820) & (!g773)) + ((g875) & (g876) & (g877) & (g878) & (g820) & (g773)));
	assign g1802 = (((!g880) & (!g881) & (!g882) & (g883) & (g820) & (g773)) + ((!g880) & (!g881) & (g882) & (!g883) & (!g820) & (g773)) + ((!g880) & (!g881) & (g882) & (g883) & (!g820) & (g773)) + ((!g880) & (!g881) & (g882) & (g883) & (g820) & (g773)) + ((!g880) & (g881) & (!g882) & (!g883) & (g820) & (!g773)) + ((!g880) & (g881) & (!g882) & (g883) & (g820) & (!g773)) + ((!g880) & (g881) & (!g882) & (g883) & (g820) & (g773)) + ((!g880) & (g881) & (g882) & (!g883) & (!g820) & (g773)) + ((!g880) & (g881) & (g882) & (!g883) & (g820) & (!g773)) + ((!g880) & (g881) & (g882) & (g883) & (!g820) & (g773)) + ((!g880) & (g881) & (g882) & (g883) & (g820) & (!g773)) + ((!g880) & (g881) & (g882) & (g883) & (g820) & (g773)) + ((g880) & (!g881) & (!g882) & (!g883) & (!g820) & (!g773)) + ((g880) & (!g881) & (!g882) & (g883) & (!g820) & (!g773)) + ((g880) & (!g881) & (!g882) & (g883) & (g820) & (g773)) + ((g880) & (!g881) & (g882) & (!g883) & (!g820) & (!g773)) + ((g880) & (!g881) & (g882) & (!g883) & (!g820) & (g773)) + ((g880) & (!g881) & (g882) & (g883) & (!g820) & (!g773)) + ((g880) & (!g881) & (g882) & (g883) & (!g820) & (g773)) + ((g880) & (!g881) & (g882) & (g883) & (g820) & (g773)) + ((g880) & (g881) & (!g882) & (!g883) & (!g820) & (!g773)) + ((g880) & (g881) & (!g882) & (!g883) & (g820) & (!g773)) + ((g880) & (g881) & (!g882) & (g883) & (!g820) & (!g773)) + ((g880) & (g881) & (!g882) & (g883) & (g820) & (!g773)) + ((g880) & (g881) & (!g882) & (g883) & (g820) & (g773)) + ((g880) & (g881) & (g882) & (!g883) & (!g820) & (!g773)) + ((g880) & (g881) & (g882) & (!g883) & (!g820) & (g773)) + ((g880) & (g881) & (g882) & (!g883) & (g820) & (!g773)) + ((g880) & (g881) & (g882) & (g883) & (!g820) & (!g773)) + ((g880) & (g881) & (g882) & (g883) & (!g820) & (g773)) + ((g880) & (g881) & (g882) & (g883) & (g820) & (!g773)) + ((g880) & (g881) & (g882) & (g883) & (g820) & (g773)));
	assign g1803 = (((!g885) & (!g886) & (!g887) & (g888) & (g820) & (g773)) + ((!g885) & (!g886) & (g887) & (!g888) & (!g820) & (g773)) + ((!g885) & (!g886) & (g887) & (g888) & (!g820) & (g773)) + ((!g885) & (!g886) & (g887) & (g888) & (g820) & (g773)) + ((!g885) & (g886) & (!g887) & (!g888) & (g820) & (!g773)) + ((!g885) & (g886) & (!g887) & (g888) & (g820) & (!g773)) + ((!g885) & (g886) & (!g887) & (g888) & (g820) & (g773)) + ((!g885) & (g886) & (g887) & (!g888) & (!g820) & (g773)) + ((!g885) & (g886) & (g887) & (!g888) & (g820) & (!g773)) + ((!g885) & (g886) & (g887) & (g888) & (!g820) & (g773)) + ((!g885) & (g886) & (g887) & (g888) & (g820) & (!g773)) + ((!g885) & (g886) & (g887) & (g888) & (g820) & (g773)) + ((g885) & (!g886) & (!g887) & (!g888) & (!g820) & (!g773)) + ((g885) & (!g886) & (!g887) & (g888) & (!g820) & (!g773)) + ((g885) & (!g886) & (!g887) & (g888) & (g820) & (g773)) + ((g885) & (!g886) & (g887) & (!g888) & (!g820) & (!g773)) + ((g885) & (!g886) & (g887) & (!g888) & (!g820) & (g773)) + ((g885) & (!g886) & (g887) & (g888) & (!g820) & (!g773)) + ((g885) & (!g886) & (g887) & (g888) & (!g820) & (g773)) + ((g885) & (!g886) & (g887) & (g888) & (g820) & (g773)) + ((g885) & (g886) & (!g887) & (!g888) & (!g820) & (!g773)) + ((g885) & (g886) & (!g887) & (!g888) & (g820) & (!g773)) + ((g885) & (g886) & (!g887) & (g888) & (!g820) & (!g773)) + ((g885) & (g886) & (!g887) & (g888) & (g820) & (!g773)) + ((g885) & (g886) & (!g887) & (g888) & (g820) & (g773)) + ((g885) & (g886) & (g887) & (!g888) & (!g820) & (!g773)) + ((g885) & (g886) & (g887) & (!g888) & (!g820) & (g773)) + ((g885) & (g886) & (g887) & (!g888) & (g820) & (!g773)) + ((g885) & (g886) & (g887) & (g888) & (!g820) & (!g773)) + ((g885) & (g886) & (g887) & (g888) & (!g820) & (g773)) + ((g885) & (g886) & (g887) & (g888) & (g820) & (!g773)) + ((g885) & (g886) & (g887) & (g888) & (g820) & (g773)));
	assign g1804 = (((!g1800) & (!g1801) & (!g1802) & (g1803) & (g677) & (g726)) + ((!g1800) & (!g1801) & (g1802) & (!g1803) & (!g677) & (g726)) + ((!g1800) & (!g1801) & (g1802) & (g1803) & (!g677) & (g726)) + ((!g1800) & (!g1801) & (g1802) & (g1803) & (g677) & (g726)) + ((!g1800) & (g1801) & (!g1802) & (!g1803) & (g677) & (!g726)) + ((!g1800) & (g1801) & (!g1802) & (g1803) & (g677) & (!g726)) + ((!g1800) & (g1801) & (!g1802) & (g1803) & (g677) & (g726)) + ((!g1800) & (g1801) & (g1802) & (!g1803) & (!g677) & (g726)) + ((!g1800) & (g1801) & (g1802) & (!g1803) & (g677) & (!g726)) + ((!g1800) & (g1801) & (g1802) & (g1803) & (!g677) & (g726)) + ((!g1800) & (g1801) & (g1802) & (g1803) & (g677) & (!g726)) + ((!g1800) & (g1801) & (g1802) & (g1803) & (g677) & (g726)) + ((g1800) & (!g1801) & (!g1802) & (!g1803) & (!g677) & (!g726)) + ((g1800) & (!g1801) & (!g1802) & (g1803) & (!g677) & (!g726)) + ((g1800) & (!g1801) & (!g1802) & (g1803) & (g677) & (g726)) + ((g1800) & (!g1801) & (g1802) & (!g1803) & (!g677) & (!g726)) + ((g1800) & (!g1801) & (g1802) & (!g1803) & (!g677) & (g726)) + ((g1800) & (!g1801) & (g1802) & (g1803) & (!g677) & (!g726)) + ((g1800) & (!g1801) & (g1802) & (g1803) & (!g677) & (g726)) + ((g1800) & (!g1801) & (g1802) & (g1803) & (g677) & (g726)) + ((g1800) & (g1801) & (!g1802) & (!g1803) & (!g677) & (!g726)) + ((g1800) & (g1801) & (!g1802) & (!g1803) & (g677) & (!g726)) + ((g1800) & (g1801) & (!g1802) & (g1803) & (!g677) & (!g726)) + ((g1800) & (g1801) & (!g1802) & (g1803) & (g677) & (!g726)) + ((g1800) & (g1801) & (!g1802) & (g1803) & (g677) & (g726)) + ((g1800) & (g1801) & (g1802) & (!g1803) & (!g677) & (!g726)) + ((g1800) & (g1801) & (g1802) & (!g1803) & (!g677) & (g726)) + ((g1800) & (g1801) & (g1802) & (!g1803) & (g677) & (!g726)) + ((g1800) & (g1801) & (g1802) & (g1803) & (!g677) & (!g726)) + ((g1800) & (g1801) & (g1802) & (g1803) & (!g677) & (g726)) + ((g1800) & (g1801) & (g1802) & (g1803) & (g677) & (!g726)) + ((g1800) & (g1801) & (g1802) & (g1803) & (g677) & (g726)));
	assign g1805 = (((!g891) & (!g892) & (!g893) & (g894) & (g677) & (g726)) + ((!g891) & (!g892) & (g893) & (!g894) & (!g677) & (g726)) + ((!g891) & (!g892) & (g893) & (g894) & (!g677) & (g726)) + ((!g891) & (!g892) & (g893) & (g894) & (g677) & (g726)) + ((!g891) & (g892) & (!g893) & (!g894) & (g677) & (!g726)) + ((!g891) & (g892) & (!g893) & (g894) & (g677) & (!g726)) + ((!g891) & (g892) & (!g893) & (g894) & (g677) & (g726)) + ((!g891) & (g892) & (g893) & (!g894) & (!g677) & (g726)) + ((!g891) & (g892) & (g893) & (!g894) & (g677) & (!g726)) + ((!g891) & (g892) & (g893) & (g894) & (!g677) & (g726)) + ((!g891) & (g892) & (g893) & (g894) & (g677) & (!g726)) + ((!g891) & (g892) & (g893) & (g894) & (g677) & (g726)) + ((g891) & (!g892) & (!g893) & (!g894) & (!g677) & (!g726)) + ((g891) & (!g892) & (!g893) & (g894) & (!g677) & (!g726)) + ((g891) & (!g892) & (!g893) & (g894) & (g677) & (g726)) + ((g891) & (!g892) & (g893) & (!g894) & (!g677) & (!g726)) + ((g891) & (!g892) & (g893) & (!g894) & (!g677) & (g726)) + ((g891) & (!g892) & (g893) & (g894) & (!g677) & (!g726)) + ((g891) & (!g892) & (g893) & (g894) & (!g677) & (g726)) + ((g891) & (!g892) & (g893) & (g894) & (g677) & (g726)) + ((g891) & (g892) & (!g893) & (!g894) & (!g677) & (!g726)) + ((g891) & (g892) & (!g893) & (!g894) & (g677) & (!g726)) + ((g891) & (g892) & (!g893) & (g894) & (!g677) & (!g726)) + ((g891) & (g892) & (!g893) & (g894) & (g677) & (!g726)) + ((g891) & (g892) & (!g893) & (g894) & (g677) & (g726)) + ((g891) & (g892) & (g893) & (!g894) & (!g677) & (!g726)) + ((g891) & (g892) & (g893) & (!g894) & (!g677) & (g726)) + ((g891) & (g892) & (g893) & (!g894) & (g677) & (!g726)) + ((g891) & (g892) & (g893) & (g894) & (!g677) & (!g726)) + ((g891) & (g892) & (g893) & (g894) & (!g677) & (g726)) + ((g891) & (g892) & (g893) & (g894) & (g677) & (!g726)) + ((g891) & (g892) & (g893) & (g894) & (g677) & (g726)));
	assign g1806 = (((!sk[80]) & (!g677) & (!g726) & (!g896) & (g897) & (!g898)) + ((!sk[80]) & (!g677) & (!g726) & (!g896) & (g897) & (g898)) + ((!sk[80]) & (!g677) & (!g726) & (g896) & (!g897) & (!g898)) + ((!sk[80]) & (!g677) & (!g726) & (g896) & (!g897) & (g898)) + ((!sk[80]) & (!g677) & (!g726) & (g896) & (g897) & (!g898)) + ((!sk[80]) & (!g677) & (!g726) & (g896) & (g897) & (g898)) + ((!sk[80]) & (!g677) & (g726) & (!g896) & (!g897) & (!g898)) + ((!sk[80]) & (!g677) & (g726) & (!g896) & (!g897) & (g898)) + ((!sk[80]) & (!g677) & (g726) & (!g896) & (g897) & (!g898)) + ((!sk[80]) & (!g677) & (g726) & (!g896) & (g897) & (g898)) + ((!sk[80]) & (!g677) & (g726) & (g896) & (!g897) & (!g898)) + ((!sk[80]) & (!g677) & (g726) & (g896) & (!g897) & (g898)) + ((!sk[80]) & (!g677) & (g726) & (g896) & (g897) & (!g898)) + ((!sk[80]) & (!g677) & (g726) & (g896) & (g897) & (g898)) + ((!sk[80]) & (g677) & (!g726) & (!g896) & (g897) & (!g898)) + ((!sk[80]) & (g677) & (!g726) & (!g896) & (g897) & (g898)) + ((!sk[80]) & (g677) & (!g726) & (g896) & (!g897) & (!g898)) + ((!sk[80]) & (g677) & (!g726) & (g896) & (!g897) & (g898)) + ((!sk[80]) & (g677) & (!g726) & (g896) & (g897) & (!g898)) + ((!sk[80]) & (g677) & (!g726) & (g896) & (g897) & (g898)) + ((!sk[80]) & (g677) & (g726) & (!g896) & (!g897) & (!g898)) + ((!sk[80]) & (g677) & (g726) & (!g896) & (!g897) & (g898)) + ((!sk[80]) & (g677) & (g726) & (!g896) & (g897) & (!g898)) + ((!sk[80]) & (g677) & (g726) & (!g896) & (g897) & (g898)) + ((!sk[80]) & (g677) & (g726) & (g896) & (!g897) & (!g898)) + ((!sk[80]) & (g677) & (g726) & (g896) & (!g897) & (g898)) + ((!sk[80]) & (g677) & (g726) & (g896) & (g897) & (!g898)) + ((!sk[80]) & (g677) & (g726) & (g896) & (g897) & (g898)) + ((sk[80]) & (!g677) & (g726) & (!g896) & (!g897) & (g898)) + ((sk[80]) & (!g677) & (g726) & (!g896) & (g897) & (g898)) + ((sk[80]) & (!g677) & (g726) & (g896) & (!g897) & (g898)) + ((sk[80]) & (!g677) & (g726) & (g896) & (g897) & (g898)) + ((sk[80]) & (g677) & (!g726) & (g896) & (!g897) & (!g898)) + ((sk[80]) & (g677) & (!g726) & (g896) & (!g897) & (g898)) + ((sk[80]) & (g677) & (!g726) & (g896) & (g897) & (!g898)) + ((sk[80]) & (g677) & (!g726) & (g896) & (g897) & (g898)) + ((sk[80]) & (g677) & (g726) & (!g896) & (g897) & (!g898)) + ((sk[80]) & (g677) & (g726) & (!g896) & (g897) & (g898)) + ((sk[80]) & (g677) & (g726) & (g896) & (g897) & (!g898)) + ((sk[80]) & (g677) & (g726) & (g896) & (g897) & (g898)));
	assign g1807 = (((!g900) & (!g901) & (!g902) & (g903) & (g677) & (g726)) + ((!g900) & (!g901) & (g902) & (!g903) & (!g677) & (g726)) + ((!g900) & (!g901) & (g902) & (g903) & (!g677) & (g726)) + ((!g900) & (!g901) & (g902) & (g903) & (g677) & (g726)) + ((!g900) & (g901) & (!g902) & (!g903) & (g677) & (!g726)) + ((!g900) & (g901) & (!g902) & (g903) & (g677) & (!g726)) + ((!g900) & (g901) & (!g902) & (g903) & (g677) & (g726)) + ((!g900) & (g901) & (g902) & (!g903) & (!g677) & (g726)) + ((!g900) & (g901) & (g902) & (!g903) & (g677) & (!g726)) + ((!g900) & (g901) & (g902) & (g903) & (!g677) & (g726)) + ((!g900) & (g901) & (g902) & (g903) & (g677) & (!g726)) + ((!g900) & (g901) & (g902) & (g903) & (g677) & (g726)) + ((g900) & (!g901) & (!g902) & (!g903) & (!g677) & (!g726)) + ((g900) & (!g901) & (!g902) & (g903) & (!g677) & (!g726)) + ((g900) & (!g901) & (!g902) & (g903) & (g677) & (g726)) + ((g900) & (!g901) & (g902) & (!g903) & (!g677) & (!g726)) + ((g900) & (!g901) & (g902) & (!g903) & (!g677) & (g726)) + ((g900) & (!g901) & (g902) & (g903) & (!g677) & (!g726)) + ((g900) & (!g901) & (g902) & (g903) & (!g677) & (g726)) + ((g900) & (!g901) & (g902) & (g903) & (g677) & (g726)) + ((g900) & (g901) & (!g902) & (!g903) & (!g677) & (!g726)) + ((g900) & (g901) & (!g902) & (!g903) & (g677) & (!g726)) + ((g900) & (g901) & (!g902) & (g903) & (!g677) & (!g726)) + ((g900) & (g901) & (!g902) & (g903) & (g677) & (!g726)) + ((g900) & (g901) & (!g902) & (g903) & (g677) & (g726)) + ((g900) & (g901) & (g902) & (!g903) & (!g677) & (!g726)) + ((g900) & (g901) & (g902) & (!g903) & (!g677) & (g726)) + ((g900) & (g901) & (g902) & (!g903) & (g677) & (!g726)) + ((g900) & (g901) & (g902) & (g903) & (!g677) & (!g726)) + ((g900) & (g901) & (g902) & (g903) & (!g677) & (g726)) + ((g900) & (g901) & (g902) & (g903) & (g677) & (!g726)) + ((g900) & (g901) & (g902) & (g903) & (g677) & (g726)));
	assign g1808 = (((!g905) & (!g906) & (!g907) & (g908) & (g677) & (g726)) + ((!g905) & (!g906) & (g907) & (!g908) & (!g677) & (g726)) + ((!g905) & (!g906) & (g907) & (g908) & (!g677) & (g726)) + ((!g905) & (!g906) & (g907) & (g908) & (g677) & (g726)) + ((!g905) & (g906) & (!g907) & (!g908) & (g677) & (!g726)) + ((!g905) & (g906) & (!g907) & (g908) & (g677) & (!g726)) + ((!g905) & (g906) & (!g907) & (g908) & (g677) & (g726)) + ((!g905) & (g906) & (g907) & (!g908) & (!g677) & (g726)) + ((!g905) & (g906) & (g907) & (!g908) & (g677) & (!g726)) + ((!g905) & (g906) & (g907) & (g908) & (!g677) & (g726)) + ((!g905) & (g906) & (g907) & (g908) & (g677) & (!g726)) + ((!g905) & (g906) & (g907) & (g908) & (g677) & (g726)) + ((g905) & (!g906) & (!g907) & (!g908) & (!g677) & (!g726)) + ((g905) & (!g906) & (!g907) & (g908) & (!g677) & (!g726)) + ((g905) & (!g906) & (!g907) & (g908) & (g677) & (g726)) + ((g905) & (!g906) & (g907) & (!g908) & (!g677) & (!g726)) + ((g905) & (!g906) & (g907) & (!g908) & (!g677) & (g726)) + ((g905) & (!g906) & (g907) & (g908) & (!g677) & (!g726)) + ((g905) & (!g906) & (g907) & (g908) & (!g677) & (g726)) + ((g905) & (!g906) & (g907) & (g908) & (g677) & (g726)) + ((g905) & (g906) & (!g907) & (!g908) & (!g677) & (!g726)) + ((g905) & (g906) & (!g907) & (!g908) & (g677) & (!g726)) + ((g905) & (g906) & (!g907) & (g908) & (!g677) & (!g726)) + ((g905) & (g906) & (!g907) & (g908) & (g677) & (!g726)) + ((g905) & (g906) & (!g907) & (g908) & (g677) & (g726)) + ((g905) & (g906) & (g907) & (!g908) & (!g677) & (!g726)) + ((g905) & (g906) & (g907) & (!g908) & (!g677) & (g726)) + ((g905) & (g906) & (g907) & (!g908) & (g677) & (!g726)) + ((g905) & (g906) & (g907) & (g908) & (!g677) & (!g726)) + ((g905) & (g906) & (g907) & (g908) & (!g677) & (g726)) + ((g905) & (g906) & (g907) & (g908) & (g677) & (!g726)) + ((g905) & (g906) & (g907) & (g908) & (g677) & (g726)));
	assign g1809 = (((!g820) & (!g773) & (!g1805) & (g1806) & (!g1807) & (!g1808)) + ((!g820) & (!g773) & (!g1805) & (g1806) & (!g1807) & (g1808)) + ((!g820) & (!g773) & (!g1805) & (g1806) & (g1807) & (!g1808)) + ((!g820) & (!g773) & (!g1805) & (g1806) & (g1807) & (g1808)) + ((!g820) & (!g773) & (g1805) & (g1806) & (!g1807) & (!g1808)) + ((!g820) & (!g773) & (g1805) & (g1806) & (!g1807) & (g1808)) + ((!g820) & (!g773) & (g1805) & (g1806) & (g1807) & (!g1808)) + ((!g820) & (!g773) & (g1805) & (g1806) & (g1807) & (g1808)) + ((!g820) & (g773) & (!g1805) & (!g1806) & (!g1807) & (g1808)) + ((!g820) & (g773) & (!g1805) & (!g1806) & (g1807) & (g1808)) + ((!g820) & (g773) & (!g1805) & (g1806) & (!g1807) & (g1808)) + ((!g820) & (g773) & (!g1805) & (g1806) & (g1807) & (g1808)) + ((!g820) & (g773) & (g1805) & (!g1806) & (!g1807) & (g1808)) + ((!g820) & (g773) & (g1805) & (!g1806) & (g1807) & (g1808)) + ((!g820) & (g773) & (g1805) & (g1806) & (!g1807) & (g1808)) + ((!g820) & (g773) & (g1805) & (g1806) & (g1807) & (g1808)) + ((g820) & (!g773) & (g1805) & (!g1806) & (!g1807) & (!g1808)) + ((g820) & (!g773) & (g1805) & (!g1806) & (!g1807) & (g1808)) + ((g820) & (!g773) & (g1805) & (!g1806) & (g1807) & (!g1808)) + ((g820) & (!g773) & (g1805) & (!g1806) & (g1807) & (g1808)) + ((g820) & (!g773) & (g1805) & (g1806) & (!g1807) & (!g1808)) + ((g820) & (!g773) & (g1805) & (g1806) & (!g1807) & (g1808)) + ((g820) & (!g773) & (g1805) & (g1806) & (g1807) & (!g1808)) + ((g820) & (!g773) & (g1805) & (g1806) & (g1807) & (g1808)) + ((g820) & (g773) & (!g1805) & (!g1806) & (g1807) & (!g1808)) + ((g820) & (g773) & (!g1805) & (!g1806) & (g1807) & (g1808)) + ((g820) & (g773) & (!g1805) & (g1806) & (g1807) & (!g1808)) + ((g820) & (g773) & (!g1805) & (g1806) & (g1807) & (g1808)) + ((g820) & (g773) & (g1805) & (!g1806) & (g1807) & (!g1808)) + ((g820) & (g773) & (g1805) & (!g1806) & (g1807) & (g1808)) + ((g820) & (g773) & (g1805) & (g1806) & (g1807) & (!g1808)) + ((g820) & (g773) & (g1805) & (g1806) & (g1807) & (g1808)));
	assign g1810 = (((!g867) & (!g1804) & (!sk[84]) & (g1809)) + ((!g867) & (!g1804) & (sk[84]) & (g1809)) + ((!g867) & (g1804) & (!sk[84]) & (!g1809)) + ((!g867) & (g1804) & (!sk[84]) & (g1809)) + ((!g867) & (g1804) & (sk[84]) & (g1809)) + ((g867) & (!g1804) & (!sk[84]) & (g1809)) + ((g867) & (g1804) & (!sk[84]) & (!g1809)) + ((g867) & (g1804) & (!sk[84]) & (g1809)) + ((g867) & (g1804) & (sk[84]) & (!g1809)) + ((g867) & (g1804) & (sk[84]) & (g1809)));
	assign g1811 = (((!g1592) & (!sk[85]) & (!g1593) & (!g1604) & (g1605) & (!g51)) + ((!g1592) & (!sk[85]) & (!g1593) & (!g1604) & (g1605) & (g51)) + ((!g1592) & (!sk[85]) & (!g1593) & (g1604) & (!g1605) & (!g51)) + ((!g1592) & (!sk[85]) & (!g1593) & (g1604) & (!g1605) & (g51)) + ((!g1592) & (!sk[85]) & (!g1593) & (g1604) & (g1605) & (!g51)) + ((!g1592) & (!sk[85]) & (!g1593) & (g1604) & (g1605) & (g51)) + ((!g1592) & (!sk[85]) & (g1593) & (!g1604) & (!g1605) & (!g51)) + ((!g1592) & (!sk[85]) & (g1593) & (!g1604) & (!g1605) & (g51)) + ((!g1592) & (!sk[85]) & (g1593) & (!g1604) & (g1605) & (!g51)) + ((!g1592) & (!sk[85]) & (g1593) & (!g1604) & (g1605) & (g51)) + ((!g1592) & (!sk[85]) & (g1593) & (g1604) & (!g1605) & (!g51)) + ((!g1592) & (!sk[85]) & (g1593) & (g1604) & (!g1605) & (g51)) + ((!g1592) & (!sk[85]) & (g1593) & (g1604) & (g1605) & (!g51)) + ((!g1592) & (!sk[85]) & (g1593) & (g1604) & (g1605) & (g51)) + ((!g1592) & (sk[85]) & (!g1593) & (g1604) & (!g1605) & (!g51)) + ((!g1592) & (sk[85]) & (!g1593) & (g1604) & (!g1605) & (g51)) + ((!g1592) & (sk[85]) & (!g1593) & (g1604) & (g1605) & (!g51)) + ((!g1592) & (sk[85]) & (!g1593) & (g1604) & (g1605) & (g51)) + ((!g1592) & (sk[85]) & (g1593) & (g1604) & (!g1605) & (!g51)) + ((!g1592) & (sk[85]) & (g1593) & (g1604) & (!g1605) & (g51)) + ((!g1592) & (sk[85]) & (g1593) & (g1604) & (g1605) & (!g51)) + ((!g1592) & (sk[85]) & (g1593) & (g1604) & (g1605) & (g51)) + ((g1592) & (!sk[85]) & (!g1593) & (!g1604) & (g1605) & (!g51)) + ((g1592) & (!sk[85]) & (!g1593) & (!g1604) & (g1605) & (g51)) + ((g1592) & (!sk[85]) & (!g1593) & (g1604) & (!g1605) & (!g51)) + ((g1592) & (!sk[85]) & (!g1593) & (g1604) & (!g1605) & (g51)) + ((g1592) & (!sk[85]) & (!g1593) & (g1604) & (g1605) & (!g51)) + ((g1592) & (!sk[85]) & (!g1593) & (g1604) & (g1605) & (g51)) + ((g1592) & (!sk[85]) & (g1593) & (!g1604) & (!g1605) & (!g51)) + ((g1592) & (!sk[85]) & (g1593) & (!g1604) & (!g1605) & (g51)) + ((g1592) & (!sk[85]) & (g1593) & (!g1604) & (g1605) & (!g51)) + ((g1592) & (!sk[85]) & (g1593) & (!g1604) & (g1605) & (g51)) + ((g1592) & (!sk[85]) & (g1593) & (g1604) & (!g1605) & (!g51)) + ((g1592) & (!sk[85]) & (g1593) & (g1604) & (!g1605) & (g51)) + ((g1592) & (!sk[85]) & (g1593) & (g1604) & (g1605) & (!g51)) + ((g1592) & (!sk[85]) & (g1593) & (g1604) & (g1605) & (g51)) + ((g1592) & (sk[85]) & (!g1593) & (g1604) & (!g1605) & (!g51)) + ((g1592) & (sk[85]) & (!g1593) & (g1604) & (!g1605) & (g51)) + ((g1592) & (sk[85]) & (g1593) & (!g1604) & (!g1605) & (g51)) + ((g1592) & (sk[85]) & (g1593) & (!g1604) & (g1605) & (g51)) + ((g1592) & (sk[85]) & (g1593) & (g1604) & (!g1605) & (g51)) + ((g1592) & (sk[85]) & (g1593) & (g1604) & (g1605) & (g51)));
	assign g1812 = (((!g132) & (!g1592) & (g1606) & (!g136) & (g1593) & (!g1605)) + ((!g132) & (g1592) & (!g1606) & (!g136) & (!g1593) & (!g1605)) + ((!g132) & (g1592) & (!g1606) & (!g136) & (!g1593) & (g1605)) + ((!g132) & (g1592) & (!g1606) & (!g136) & (g1593) & (!g1605)) + ((!g132) & (g1592) & (!g1606) & (!g136) & (g1593) & (g1605)) + ((!g132) & (g1592) & (g1606) & (!g136) & (g1593) & (!g1605)) + ((g132) & (!g1592) & (!g1606) & (!g136) & (!g1593) & (!g1605)) + ((g132) & (!g1592) & (!g1606) & (!g136) & (!g1593) & (g1605)) + ((g132) & (!g1592) & (!g1606) & (!g136) & (g1593) & (!g1605)) + ((g132) & (!g1592) & (!g1606) & (!g136) & (g1593) & (g1605)) + ((g132) & (!g1592) & (g1606) & (!g136) & (g1593) & (!g1605)) + ((g132) & (g1592) & (!g1606) & (!g136) & (!g1593) & (!g1605)) + ((g132) & (g1592) & (!g1606) & (!g136) & (!g1593) & (g1605)) + ((g132) & (g1592) & (!g1606) & (!g136) & (g1593) & (!g1605)) + ((g132) & (g1592) & (!g1606) & (!g136) & (g1593) & (g1605)) + ((g132) & (g1592) & (g1606) & (!g136) & (g1593) & (!g1605)));
	assign g1813 = (((!g132) & (!g1810) & (!sk[87]) & (!g1811) & (g1812)) + ((!g132) & (!g1810) & (!sk[87]) & (g1811) & (!g1812)) + ((!g132) & (!g1810) & (!sk[87]) & (g1811) & (g1812)) + ((!g132) & (!g1810) & (sk[87]) & (g1811) & (g1812)) + ((!g132) & (g1810) & (!sk[87]) & (!g1811) & (!g1812)) + ((!g132) & (g1810) & (!sk[87]) & (!g1811) & (g1812)) + ((!g132) & (g1810) & (!sk[87]) & (g1811) & (!g1812)) + ((!g132) & (g1810) & (!sk[87]) & (g1811) & (g1812)) + ((!g132) & (g1810) & (sk[87]) & (g1811) & (g1812)) + ((g132) & (!g1810) & (!sk[87]) & (!g1811) & (g1812)) + ((g132) & (!g1810) & (!sk[87]) & (g1811) & (!g1812)) + ((g132) & (!g1810) & (!sk[87]) & (g1811) & (g1812)) + ((g132) & (g1810) & (!sk[87]) & (!g1811) & (!g1812)) + ((g132) & (g1810) & (!sk[87]) & (!g1811) & (g1812)) + ((g132) & (g1810) & (!sk[87]) & (g1811) & (!g1812)) + ((g132) & (g1810) & (!sk[87]) & (g1811) & (g1812)) + ((g132) & (g1810) & (sk[87]) & (!g1811) & (g1812)) + ((g132) & (g1810) & (sk[87]) & (g1811) & (g1812)));
	assign g1814 = (((!g918) & (!g919) & (!g920) & (g921) & (g820) & (g773)) + ((!g918) & (!g919) & (g920) & (!g921) & (!g820) & (g773)) + ((!g918) & (!g919) & (g920) & (g921) & (!g820) & (g773)) + ((!g918) & (!g919) & (g920) & (g921) & (g820) & (g773)) + ((!g918) & (g919) & (!g920) & (!g921) & (g820) & (!g773)) + ((!g918) & (g919) & (!g920) & (g921) & (g820) & (!g773)) + ((!g918) & (g919) & (!g920) & (g921) & (g820) & (g773)) + ((!g918) & (g919) & (g920) & (!g921) & (!g820) & (g773)) + ((!g918) & (g919) & (g920) & (!g921) & (g820) & (!g773)) + ((!g918) & (g919) & (g920) & (g921) & (!g820) & (g773)) + ((!g918) & (g919) & (g920) & (g921) & (g820) & (!g773)) + ((!g918) & (g919) & (g920) & (g921) & (g820) & (g773)) + ((g918) & (!g919) & (!g920) & (!g921) & (!g820) & (!g773)) + ((g918) & (!g919) & (!g920) & (g921) & (!g820) & (!g773)) + ((g918) & (!g919) & (!g920) & (g921) & (g820) & (g773)) + ((g918) & (!g919) & (g920) & (!g921) & (!g820) & (!g773)) + ((g918) & (!g919) & (g920) & (!g921) & (!g820) & (g773)) + ((g918) & (!g919) & (g920) & (g921) & (!g820) & (!g773)) + ((g918) & (!g919) & (g920) & (g921) & (!g820) & (g773)) + ((g918) & (!g919) & (g920) & (g921) & (g820) & (g773)) + ((g918) & (g919) & (!g920) & (!g921) & (!g820) & (!g773)) + ((g918) & (g919) & (!g920) & (!g921) & (g820) & (!g773)) + ((g918) & (g919) & (!g920) & (g921) & (!g820) & (!g773)) + ((g918) & (g919) & (!g920) & (g921) & (g820) & (!g773)) + ((g918) & (g919) & (!g920) & (g921) & (g820) & (g773)) + ((g918) & (g919) & (g920) & (!g921) & (!g820) & (!g773)) + ((g918) & (g919) & (g920) & (!g921) & (!g820) & (g773)) + ((g918) & (g919) & (g920) & (!g921) & (g820) & (!g773)) + ((g918) & (g919) & (g920) & (g921) & (!g820) & (!g773)) + ((g918) & (g919) & (g920) & (g921) & (!g820) & (g773)) + ((g918) & (g919) & (g920) & (g921) & (g820) & (!g773)) + ((g918) & (g919) & (g920) & (g921) & (g820) & (g773)));
	assign g1815 = (((!g923) & (!g924) & (!g925) & (g926) & (g820) & (g773)) + ((!g923) & (!g924) & (g925) & (!g926) & (!g820) & (g773)) + ((!g923) & (!g924) & (g925) & (g926) & (!g820) & (g773)) + ((!g923) & (!g924) & (g925) & (g926) & (g820) & (g773)) + ((!g923) & (g924) & (!g925) & (!g926) & (g820) & (!g773)) + ((!g923) & (g924) & (!g925) & (g926) & (g820) & (!g773)) + ((!g923) & (g924) & (!g925) & (g926) & (g820) & (g773)) + ((!g923) & (g924) & (g925) & (!g926) & (!g820) & (g773)) + ((!g923) & (g924) & (g925) & (!g926) & (g820) & (!g773)) + ((!g923) & (g924) & (g925) & (g926) & (!g820) & (g773)) + ((!g923) & (g924) & (g925) & (g926) & (g820) & (!g773)) + ((!g923) & (g924) & (g925) & (g926) & (g820) & (g773)) + ((g923) & (!g924) & (!g925) & (!g926) & (!g820) & (!g773)) + ((g923) & (!g924) & (!g925) & (g926) & (!g820) & (!g773)) + ((g923) & (!g924) & (!g925) & (g926) & (g820) & (g773)) + ((g923) & (!g924) & (g925) & (!g926) & (!g820) & (!g773)) + ((g923) & (!g924) & (g925) & (!g926) & (!g820) & (g773)) + ((g923) & (!g924) & (g925) & (g926) & (!g820) & (!g773)) + ((g923) & (!g924) & (g925) & (g926) & (!g820) & (g773)) + ((g923) & (!g924) & (g925) & (g926) & (g820) & (g773)) + ((g923) & (g924) & (!g925) & (!g926) & (!g820) & (!g773)) + ((g923) & (g924) & (!g925) & (!g926) & (g820) & (!g773)) + ((g923) & (g924) & (!g925) & (g926) & (!g820) & (!g773)) + ((g923) & (g924) & (!g925) & (g926) & (g820) & (!g773)) + ((g923) & (g924) & (!g925) & (g926) & (g820) & (g773)) + ((g923) & (g924) & (g925) & (!g926) & (!g820) & (!g773)) + ((g923) & (g924) & (g925) & (!g926) & (!g820) & (g773)) + ((g923) & (g924) & (g925) & (!g926) & (g820) & (!g773)) + ((g923) & (g924) & (g925) & (g926) & (!g820) & (!g773)) + ((g923) & (g924) & (g925) & (g926) & (!g820) & (g773)) + ((g923) & (g924) & (g925) & (g926) & (g820) & (!g773)) + ((g923) & (g924) & (g925) & (g926) & (g820) & (g773)));
	assign g1816 = (((!g928) & (!g929) & (!g930) & (g931) & (g820) & (g773)) + ((!g928) & (!g929) & (g930) & (!g931) & (!g820) & (g773)) + ((!g928) & (!g929) & (g930) & (g931) & (!g820) & (g773)) + ((!g928) & (!g929) & (g930) & (g931) & (g820) & (g773)) + ((!g928) & (g929) & (!g930) & (!g931) & (g820) & (!g773)) + ((!g928) & (g929) & (!g930) & (g931) & (g820) & (!g773)) + ((!g928) & (g929) & (!g930) & (g931) & (g820) & (g773)) + ((!g928) & (g929) & (g930) & (!g931) & (!g820) & (g773)) + ((!g928) & (g929) & (g930) & (!g931) & (g820) & (!g773)) + ((!g928) & (g929) & (g930) & (g931) & (!g820) & (g773)) + ((!g928) & (g929) & (g930) & (g931) & (g820) & (!g773)) + ((!g928) & (g929) & (g930) & (g931) & (g820) & (g773)) + ((g928) & (!g929) & (!g930) & (!g931) & (!g820) & (!g773)) + ((g928) & (!g929) & (!g930) & (g931) & (!g820) & (!g773)) + ((g928) & (!g929) & (!g930) & (g931) & (g820) & (g773)) + ((g928) & (!g929) & (g930) & (!g931) & (!g820) & (!g773)) + ((g928) & (!g929) & (g930) & (!g931) & (!g820) & (g773)) + ((g928) & (!g929) & (g930) & (g931) & (!g820) & (!g773)) + ((g928) & (!g929) & (g930) & (g931) & (!g820) & (g773)) + ((g928) & (!g929) & (g930) & (g931) & (g820) & (g773)) + ((g928) & (g929) & (!g930) & (!g931) & (!g820) & (!g773)) + ((g928) & (g929) & (!g930) & (!g931) & (g820) & (!g773)) + ((g928) & (g929) & (!g930) & (g931) & (!g820) & (!g773)) + ((g928) & (g929) & (!g930) & (g931) & (g820) & (!g773)) + ((g928) & (g929) & (!g930) & (g931) & (g820) & (g773)) + ((g928) & (g929) & (g930) & (!g931) & (!g820) & (!g773)) + ((g928) & (g929) & (g930) & (!g931) & (!g820) & (g773)) + ((g928) & (g929) & (g930) & (!g931) & (g820) & (!g773)) + ((g928) & (g929) & (g930) & (g931) & (!g820) & (!g773)) + ((g928) & (g929) & (g930) & (g931) & (!g820) & (g773)) + ((g928) & (g929) & (g930) & (g931) & (g820) & (!g773)) + ((g928) & (g929) & (g930) & (g931) & (g820) & (g773)));
	assign g1817 = (((!g933) & (!g934) & (!g935) & (g936) & (g820) & (g773)) + ((!g933) & (!g934) & (g935) & (!g936) & (!g820) & (g773)) + ((!g933) & (!g934) & (g935) & (g936) & (!g820) & (g773)) + ((!g933) & (!g934) & (g935) & (g936) & (g820) & (g773)) + ((!g933) & (g934) & (!g935) & (!g936) & (g820) & (!g773)) + ((!g933) & (g934) & (!g935) & (g936) & (g820) & (!g773)) + ((!g933) & (g934) & (!g935) & (g936) & (g820) & (g773)) + ((!g933) & (g934) & (g935) & (!g936) & (!g820) & (g773)) + ((!g933) & (g934) & (g935) & (!g936) & (g820) & (!g773)) + ((!g933) & (g934) & (g935) & (g936) & (!g820) & (g773)) + ((!g933) & (g934) & (g935) & (g936) & (g820) & (!g773)) + ((!g933) & (g934) & (g935) & (g936) & (g820) & (g773)) + ((g933) & (!g934) & (!g935) & (!g936) & (!g820) & (!g773)) + ((g933) & (!g934) & (!g935) & (g936) & (!g820) & (!g773)) + ((g933) & (!g934) & (!g935) & (g936) & (g820) & (g773)) + ((g933) & (!g934) & (g935) & (!g936) & (!g820) & (!g773)) + ((g933) & (!g934) & (g935) & (!g936) & (!g820) & (g773)) + ((g933) & (!g934) & (g935) & (g936) & (!g820) & (!g773)) + ((g933) & (!g934) & (g935) & (g936) & (!g820) & (g773)) + ((g933) & (!g934) & (g935) & (g936) & (g820) & (g773)) + ((g933) & (g934) & (!g935) & (!g936) & (!g820) & (!g773)) + ((g933) & (g934) & (!g935) & (!g936) & (g820) & (!g773)) + ((g933) & (g934) & (!g935) & (g936) & (!g820) & (!g773)) + ((g933) & (g934) & (!g935) & (g936) & (g820) & (!g773)) + ((g933) & (g934) & (!g935) & (g936) & (g820) & (g773)) + ((g933) & (g934) & (g935) & (!g936) & (!g820) & (!g773)) + ((g933) & (g934) & (g935) & (!g936) & (!g820) & (g773)) + ((g933) & (g934) & (g935) & (!g936) & (g820) & (!g773)) + ((g933) & (g934) & (g935) & (g936) & (!g820) & (!g773)) + ((g933) & (g934) & (g935) & (g936) & (!g820) & (g773)) + ((g933) & (g934) & (g935) & (g936) & (g820) & (!g773)) + ((g933) & (g934) & (g935) & (g936) & (g820) & (g773)));
	assign g1818 = (((!g1814) & (!g1815) & (!g1816) & (g1817) & (g677) & (g726)) + ((!g1814) & (!g1815) & (g1816) & (!g1817) & (!g677) & (g726)) + ((!g1814) & (!g1815) & (g1816) & (g1817) & (!g677) & (g726)) + ((!g1814) & (!g1815) & (g1816) & (g1817) & (g677) & (g726)) + ((!g1814) & (g1815) & (!g1816) & (!g1817) & (g677) & (!g726)) + ((!g1814) & (g1815) & (!g1816) & (g1817) & (g677) & (!g726)) + ((!g1814) & (g1815) & (!g1816) & (g1817) & (g677) & (g726)) + ((!g1814) & (g1815) & (g1816) & (!g1817) & (!g677) & (g726)) + ((!g1814) & (g1815) & (g1816) & (!g1817) & (g677) & (!g726)) + ((!g1814) & (g1815) & (g1816) & (g1817) & (!g677) & (g726)) + ((!g1814) & (g1815) & (g1816) & (g1817) & (g677) & (!g726)) + ((!g1814) & (g1815) & (g1816) & (g1817) & (g677) & (g726)) + ((g1814) & (!g1815) & (!g1816) & (!g1817) & (!g677) & (!g726)) + ((g1814) & (!g1815) & (!g1816) & (g1817) & (!g677) & (!g726)) + ((g1814) & (!g1815) & (!g1816) & (g1817) & (g677) & (g726)) + ((g1814) & (!g1815) & (g1816) & (!g1817) & (!g677) & (!g726)) + ((g1814) & (!g1815) & (g1816) & (!g1817) & (!g677) & (g726)) + ((g1814) & (!g1815) & (g1816) & (g1817) & (!g677) & (!g726)) + ((g1814) & (!g1815) & (g1816) & (g1817) & (!g677) & (g726)) + ((g1814) & (!g1815) & (g1816) & (g1817) & (g677) & (g726)) + ((g1814) & (g1815) & (!g1816) & (!g1817) & (!g677) & (!g726)) + ((g1814) & (g1815) & (!g1816) & (!g1817) & (g677) & (!g726)) + ((g1814) & (g1815) & (!g1816) & (g1817) & (!g677) & (!g726)) + ((g1814) & (g1815) & (!g1816) & (g1817) & (g677) & (!g726)) + ((g1814) & (g1815) & (!g1816) & (g1817) & (g677) & (g726)) + ((g1814) & (g1815) & (g1816) & (!g1817) & (!g677) & (!g726)) + ((g1814) & (g1815) & (g1816) & (!g1817) & (!g677) & (g726)) + ((g1814) & (g1815) & (g1816) & (!g1817) & (g677) & (!g726)) + ((g1814) & (g1815) & (g1816) & (g1817) & (!g677) & (!g726)) + ((g1814) & (g1815) & (g1816) & (g1817) & (!g677) & (g726)) + ((g1814) & (g1815) & (g1816) & (g1817) & (g677) & (!g726)) + ((g1814) & (g1815) & (g1816) & (g1817) & (g677) & (g726)));
	assign g1819 = (((!g939) & (!g940) & (!g941) & (g942) & (g677) & (g726)) + ((!g939) & (!g940) & (g941) & (!g942) & (!g677) & (g726)) + ((!g939) & (!g940) & (g941) & (g942) & (!g677) & (g726)) + ((!g939) & (!g940) & (g941) & (g942) & (g677) & (g726)) + ((!g939) & (g940) & (!g941) & (!g942) & (g677) & (!g726)) + ((!g939) & (g940) & (!g941) & (g942) & (g677) & (!g726)) + ((!g939) & (g940) & (!g941) & (g942) & (g677) & (g726)) + ((!g939) & (g940) & (g941) & (!g942) & (!g677) & (g726)) + ((!g939) & (g940) & (g941) & (!g942) & (g677) & (!g726)) + ((!g939) & (g940) & (g941) & (g942) & (!g677) & (g726)) + ((!g939) & (g940) & (g941) & (g942) & (g677) & (!g726)) + ((!g939) & (g940) & (g941) & (g942) & (g677) & (g726)) + ((g939) & (!g940) & (!g941) & (!g942) & (!g677) & (!g726)) + ((g939) & (!g940) & (!g941) & (g942) & (!g677) & (!g726)) + ((g939) & (!g940) & (!g941) & (g942) & (g677) & (g726)) + ((g939) & (!g940) & (g941) & (!g942) & (!g677) & (!g726)) + ((g939) & (!g940) & (g941) & (!g942) & (!g677) & (g726)) + ((g939) & (!g940) & (g941) & (g942) & (!g677) & (!g726)) + ((g939) & (!g940) & (g941) & (g942) & (!g677) & (g726)) + ((g939) & (!g940) & (g941) & (g942) & (g677) & (g726)) + ((g939) & (g940) & (!g941) & (!g942) & (!g677) & (!g726)) + ((g939) & (g940) & (!g941) & (!g942) & (g677) & (!g726)) + ((g939) & (g940) & (!g941) & (g942) & (!g677) & (!g726)) + ((g939) & (g940) & (!g941) & (g942) & (g677) & (!g726)) + ((g939) & (g940) & (!g941) & (g942) & (g677) & (g726)) + ((g939) & (g940) & (g941) & (!g942) & (!g677) & (!g726)) + ((g939) & (g940) & (g941) & (!g942) & (!g677) & (g726)) + ((g939) & (g940) & (g941) & (!g942) & (g677) & (!g726)) + ((g939) & (g940) & (g941) & (g942) & (!g677) & (!g726)) + ((g939) & (g940) & (g941) & (g942) & (!g677) & (g726)) + ((g939) & (g940) & (g941) & (g942) & (g677) & (!g726)) + ((g939) & (g940) & (g941) & (g942) & (g677) & (g726)));
	assign g1820 = (((!g677) & (!g726) & (!g944) & (g945) & (!sk[94]) & (!g946)) + ((!g677) & (!g726) & (!g944) & (g945) & (!sk[94]) & (g946)) + ((!g677) & (!g726) & (g944) & (!g945) & (!sk[94]) & (!g946)) + ((!g677) & (!g726) & (g944) & (!g945) & (!sk[94]) & (g946)) + ((!g677) & (!g726) & (g944) & (g945) & (!sk[94]) & (!g946)) + ((!g677) & (!g726) & (g944) & (g945) & (!sk[94]) & (g946)) + ((!g677) & (g726) & (!g944) & (!g945) & (!sk[94]) & (!g946)) + ((!g677) & (g726) & (!g944) & (!g945) & (!sk[94]) & (g946)) + ((!g677) & (g726) & (!g944) & (!g945) & (sk[94]) & (g946)) + ((!g677) & (g726) & (!g944) & (g945) & (!sk[94]) & (!g946)) + ((!g677) & (g726) & (!g944) & (g945) & (!sk[94]) & (g946)) + ((!g677) & (g726) & (!g944) & (g945) & (sk[94]) & (g946)) + ((!g677) & (g726) & (g944) & (!g945) & (!sk[94]) & (!g946)) + ((!g677) & (g726) & (g944) & (!g945) & (!sk[94]) & (g946)) + ((!g677) & (g726) & (g944) & (!g945) & (sk[94]) & (g946)) + ((!g677) & (g726) & (g944) & (g945) & (!sk[94]) & (!g946)) + ((!g677) & (g726) & (g944) & (g945) & (!sk[94]) & (g946)) + ((!g677) & (g726) & (g944) & (g945) & (sk[94]) & (g946)) + ((g677) & (!g726) & (!g944) & (g945) & (!sk[94]) & (!g946)) + ((g677) & (!g726) & (!g944) & (g945) & (!sk[94]) & (g946)) + ((g677) & (!g726) & (g944) & (!g945) & (!sk[94]) & (!g946)) + ((g677) & (!g726) & (g944) & (!g945) & (!sk[94]) & (g946)) + ((g677) & (!g726) & (g944) & (!g945) & (sk[94]) & (!g946)) + ((g677) & (!g726) & (g944) & (!g945) & (sk[94]) & (g946)) + ((g677) & (!g726) & (g944) & (g945) & (!sk[94]) & (!g946)) + ((g677) & (!g726) & (g944) & (g945) & (!sk[94]) & (g946)) + ((g677) & (!g726) & (g944) & (g945) & (sk[94]) & (!g946)) + ((g677) & (!g726) & (g944) & (g945) & (sk[94]) & (g946)) + ((g677) & (g726) & (!g944) & (!g945) & (!sk[94]) & (!g946)) + ((g677) & (g726) & (!g944) & (!g945) & (!sk[94]) & (g946)) + ((g677) & (g726) & (!g944) & (g945) & (!sk[94]) & (!g946)) + ((g677) & (g726) & (!g944) & (g945) & (!sk[94]) & (g946)) + ((g677) & (g726) & (!g944) & (g945) & (sk[94]) & (!g946)) + ((g677) & (g726) & (!g944) & (g945) & (sk[94]) & (g946)) + ((g677) & (g726) & (g944) & (!g945) & (!sk[94]) & (!g946)) + ((g677) & (g726) & (g944) & (!g945) & (!sk[94]) & (g946)) + ((g677) & (g726) & (g944) & (g945) & (!sk[94]) & (!g946)) + ((g677) & (g726) & (g944) & (g945) & (!sk[94]) & (g946)) + ((g677) & (g726) & (g944) & (g945) & (sk[94]) & (!g946)) + ((g677) & (g726) & (g944) & (g945) & (sk[94]) & (g946)));
	assign g1821 = (((!g948) & (!g949) & (!g950) & (g951) & (g677) & (g726)) + ((!g948) & (!g949) & (g950) & (!g951) & (!g677) & (g726)) + ((!g948) & (!g949) & (g950) & (g951) & (!g677) & (g726)) + ((!g948) & (!g949) & (g950) & (g951) & (g677) & (g726)) + ((!g948) & (g949) & (!g950) & (!g951) & (g677) & (!g726)) + ((!g948) & (g949) & (!g950) & (g951) & (g677) & (!g726)) + ((!g948) & (g949) & (!g950) & (g951) & (g677) & (g726)) + ((!g948) & (g949) & (g950) & (!g951) & (!g677) & (g726)) + ((!g948) & (g949) & (g950) & (!g951) & (g677) & (!g726)) + ((!g948) & (g949) & (g950) & (g951) & (!g677) & (g726)) + ((!g948) & (g949) & (g950) & (g951) & (g677) & (!g726)) + ((!g948) & (g949) & (g950) & (g951) & (g677) & (g726)) + ((g948) & (!g949) & (!g950) & (!g951) & (!g677) & (!g726)) + ((g948) & (!g949) & (!g950) & (g951) & (!g677) & (!g726)) + ((g948) & (!g949) & (!g950) & (g951) & (g677) & (g726)) + ((g948) & (!g949) & (g950) & (!g951) & (!g677) & (!g726)) + ((g948) & (!g949) & (g950) & (!g951) & (!g677) & (g726)) + ((g948) & (!g949) & (g950) & (g951) & (!g677) & (!g726)) + ((g948) & (!g949) & (g950) & (g951) & (!g677) & (g726)) + ((g948) & (!g949) & (g950) & (g951) & (g677) & (g726)) + ((g948) & (g949) & (!g950) & (!g951) & (!g677) & (!g726)) + ((g948) & (g949) & (!g950) & (!g951) & (g677) & (!g726)) + ((g948) & (g949) & (!g950) & (g951) & (!g677) & (!g726)) + ((g948) & (g949) & (!g950) & (g951) & (g677) & (!g726)) + ((g948) & (g949) & (!g950) & (g951) & (g677) & (g726)) + ((g948) & (g949) & (g950) & (!g951) & (!g677) & (!g726)) + ((g948) & (g949) & (g950) & (!g951) & (!g677) & (g726)) + ((g948) & (g949) & (g950) & (!g951) & (g677) & (!g726)) + ((g948) & (g949) & (g950) & (g951) & (!g677) & (!g726)) + ((g948) & (g949) & (g950) & (g951) & (!g677) & (g726)) + ((g948) & (g949) & (g950) & (g951) & (g677) & (!g726)) + ((g948) & (g949) & (g950) & (g951) & (g677) & (g726)));
	assign g1822 = (((!g953) & (!g954) & (!g955) & (g956) & (g677) & (g726)) + ((!g953) & (!g954) & (g955) & (!g956) & (!g677) & (g726)) + ((!g953) & (!g954) & (g955) & (g956) & (!g677) & (g726)) + ((!g953) & (!g954) & (g955) & (g956) & (g677) & (g726)) + ((!g953) & (g954) & (!g955) & (!g956) & (g677) & (!g726)) + ((!g953) & (g954) & (!g955) & (g956) & (g677) & (!g726)) + ((!g953) & (g954) & (!g955) & (g956) & (g677) & (g726)) + ((!g953) & (g954) & (g955) & (!g956) & (!g677) & (g726)) + ((!g953) & (g954) & (g955) & (!g956) & (g677) & (!g726)) + ((!g953) & (g954) & (g955) & (g956) & (!g677) & (g726)) + ((!g953) & (g954) & (g955) & (g956) & (g677) & (!g726)) + ((!g953) & (g954) & (g955) & (g956) & (g677) & (g726)) + ((g953) & (!g954) & (!g955) & (!g956) & (!g677) & (!g726)) + ((g953) & (!g954) & (!g955) & (g956) & (!g677) & (!g726)) + ((g953) & (!g954) & (!g955) & (g956) & (g677) & (g726)) + ((g953) & (!g954) & (g955) & (!g956) & (!g677) & (!g726)) + ((g953) & (!g954) & (g955) & (!g956) & (!g677) & (g726)) + ((g953) & (!g954) & (g955) & (g956) & (!g677) & (!g726)) + ((g953) & (!g954) & (g955) & (g956) & (!g677) & (g726)) + ((g953) & (!g954) & (g955) & (g956) & (g677) & (g726)) + ((g953) & (g954) & (!g955) & (!g956) & (!g677) & (!g726)) + ((g953) & (g954) & (!g955) & (!g956) & (g677) & (!g726)) + ((g953) & (g954) & (!g955) & (g956) & (!g677) & (!g726)) + ((g953) & (g954) & (!g955) & (g956) & (g677) & (!g726)) + ((g953) & (g954) & (!g955) & (g956) & (g677) & (g726)) + ((g953) & (g954) & (g955) & (!g956) & (!g677) & (!g726)) + ((g953) & (g954) & (g955) & (!g956) & (!g677) & (g726)) + ((g953) & (g954) & (g955) & (!g956) & (g677) & (!g726)) + ((g953) & (g954) & (g955) & (g956) & (!g677) & (!g726)) + ((g953) & (g954) & (g955) & (g956) & (!g677) & (g726)) + ((g953) & (g954) & (g955) & (g956) & (g677) & (!g726)) + ((g953) & (g954) & (g955) & (g956) & (g677) & (g726)));
	assign g1823 = (((!g820) & (!g773) & (!g1819) & (g1820) & (!g1821) & (!g1822)) + ((!g820) & (!g773) & (!g1819) & (g1820) & (!g1821) & (g1822)) + ((!g820) & (!g773) & (!g1819) & (g1820) & (g1821) & (!g1822)) + ((!g820) & (!g773) & (!g1819) & (g1820) & (g1821) & (g1822)) + ((!g820) & (!g773) & (g1819) & (g1820) & (!g1821) & (!g1822)) + ((!g820) & (!g773) & (g1819) & (g1820) & (!g1821) & (g1822)) + ((!g820) & (!g773) & (g1819) & (g1820) & (g1821) & (!g1822)) + ((!g820) & (!g773) & (g1819) & (g1820) & (g1821) & (g1822)) + ((!g820) & (g773) & (!g1819) & (!g1820) & (!g1821) & (g1822)) + ((!g820) & (g773) & (!g1819) & (!g1820) & (g1821) & (g1822)) + ((!g820) & (g773) & (!g1819) & (g1820) & (!g1821) & (g1822)) + ((!g820) & (g773) & (!g1819) & (g1820) & (g1821) & (g1822)) + ((!g820) & (g773) & (g1819) & (!g1820) & (!g1821) & (g1822)) + ((!g820) & (g773) & (g1819) & (!g1820) & (g1821) & (g1822)) + ((!g820) & (g773) & (g1819) & (g1820) & (!g1821) & (g1822)) + ((!g820) & (g773) & (g1819) & (g1820) & (g1821) & (g1822)) + ((g820) & (!g773) & (g1819) & (!g1820) & (!g1821) & (!g1822)) + ((g820) & (!g773) & (g1819) & (!g1820) & (!g1821) & (g1822)) + ((g820) & (!g773) & (g1819) & (!g1820) & (g1821) & (!g1822)) + ((g820) & (!g773) & (g1819) & (!g1820) & (g1821) & (g1822)) + ((g820) & (!g773) & (g1819) & (g1820) & (!g1821) & (!g1822)) + ((g820) & (!g773) & (g1819) & (g1820) & (!g1821) & (g1822)) + ((g820) & (!g773) & (g1819) & (g1820) & (g1821) & (!g1822)) + ((g820) & (!g773) & (g1819) & (g1820) & (g1821) & (g1822)) + ((g820) & (g773) & (!g1819) & (!g1820) & (g1821) & (!g1822)) + ((g820) & (g773) & (!g1819) & (!g1820) & (g1821) & (g1822)) + ((g820) & (g773) & (!g1819) & (g1820) & (g1821) & (!g1822)) + ((g820) & (g773) & (!g1819) & (g1820) & (g1821) & (g1822)) + ((g820) & (g773) & (g1819) & (!g1820) & (g1821) & (!g1822)) + ((g820) & (g773) & (g1819) & (!g1820) & (g1821) & (g1822)) + ((g820) & (g773) & (g1819) & (g1820) & (g1821) & (!g1822)) + ((g820) & (g773) & (g1819) & (g1820) & (g1821) & (g1822)));
	assign g1824 = (((!g867) & (!sk[98]) & (!g1818) & (g1823)) + ((!g867) & (!sk[98]) & (g1818) & (!g1823)) + ((!g867) & (!sk[98]) & (g1818) & (g1823)) + ((!g867) & (sk[98]) & (!g1818) & (g1823)) + ((!g867) & (sk[98]) & (g1818) & (g1823)) + ((g867) & (!sk[98]) & (!g1818) & (g1823)) + ((g867) & (!sk[98]) & (g1818) & (!g1823)) + ((g867) & (!sk[98]) & (g1818) & (g1823)) + ((g867) & (sk[98]) & (g1818) & (!g1823)) + ((g867) & (sk[98]) & (g1818) & (g1823)));
	assign g1825 = (((!g1592) & (!g1593) & (!g1605) & (g1620) & (!sk[99]) & (!g52)) + ((!g1592) & (!g1593) & (!g1605) & (g1620) & (!sk[99]) & (g52)) + ((!g1592) & (!g1593) & (!g1605) & (g1620) & (sk[99]) & (!g52)) + ((!g1592) & (!g1593) & (!g1605) & (g1620) & (sk[99]) & (g52)) + ((!g1592) & (!g1593) & (g1605) & (!g1620) & (!sk[99]) & (!g52)) + ((!g1592) & (!g1593) & (g1605) & (!g1620) & (!sk[99]) & (g52)) + ((!g1592) & (!g1593) & (g1605) & (g1620) & (!sk[99]) & (!g52)) + ((!g1592) & (!g1593) & (g1605) & (g1620) & (!sk[99]) & (g52)) + ((!g1592) & (!g1593) & (g1605) & (g1620) & (sk[99]) & (!g52)) + ((!g1592) & (!g1593) & (g1605) & (g1620) & (sk[99]) & (g52)) + ((!g1592) & (g1593) & (!g1605) & (!g1620) & (!sk[99]) & (!g52)) + ((!g1592) & (g1593) & (!g1605) & (!g1620) & (!sk[99]) & (g52)) + ((!g1592) & (g1593) & (!g1605) & (g1620) & (!sk[99]) & (!g52)) + ((!g1592) & (g1593) & (!g1605) & (g1620) & (!sk[99]) & (g52)) + ((!g1592) & (g1593) & (!g1605) & (g1620) & (sk[99]) & (!g52)) + ((!g1592) & (g1593) & (!g1605) & (g1620) & (sk[99]) & (g52)) + ((!g1592) & (g1593) & (g1605) & (!g1620) & (!sk[99]) & (!g52)) + ((!g1592) & (g1593) & (g1605) & (!g1620) & (!sk[99]) & (g52)) + ((!g1592) & (g1593) & (g1605) & (g1620) & (!sk[99]) & (!g52)) + ((!g1592) & (g1593) & (g1605) & (g1620) & (!sk[99]) & (g52)) + ((!g1592) & (g1593) & (g1605) & (g1620) & (sk[99]) & (!g52)) + ((!g1592) & (g1593) & (g1605) & (g1620) & (sk[99]) & (g52)) + ((g1592) & (!g1593) & (!g1605) & (g1620) & (!sk[99]) & (!g52)) + ((g1592) & (!g1593) & (!g1605) & (g1620) & (!sk[99]) & (g52)) + ((g1592) & (!g1593) & (!g1605) & (g1620) & (sk[99]) & (!g52)) + ((g1592) & (!g1593) & (!g1605) & (g1620) & (sk[99]) & (g52)) + ((g1592) & (!g1593) & (g1605) & (!g1620) & (!sk[99]) & (!g52)) + ((g1592) & (!g1593) & (g1605) & (!g1620) & (!sk[99]) & (g52)) + ((g1592) & (!g1593) & (g1605) & (g1620) & (!sk[99]) & (!g52)) + ((g1592) & (!g1593) & (g1605) & (g1620) & (!sk[99]) & (g52)) + ((g1592) & (g1593) & (!g1605) & (!g1620) & (!sk[99]) & (!g52)) + ((g1592) & (g1593) & (!g1605) & (!g1620) & (!sk[99]) & (g52)) + ((g1592) & (g1593) & (!g1605) & (!g1620) & (sk[99]) & (g52)) + ((g1592) & (g1593) & (!g1605) & (g1620) & (!sk[99]) & (!g52)) + ((g1592) & (g1593) & (!g1605) & (g1620) & (!sk[99]) & (g52)) + ((g1592) & (g1593) & (!g1605) & (g1620) & (sk[99]) & (g52)) + ((g1592) & (g1593) & (g1605) & (!g1620) & (!sk[99]) & (!g52)) + ((g1592) & (g1593) & (g1605) & (!g1620) & (!sk[99]) & (g52)) + ((g1592) & (g1593) & (g1605) & (!g1620) & (sk[99]) & (g52)) + ((g1592) & (g1593) & (g1605) & (g1620) & (!sk[99]) & (!g52)) + ((g1592) & (g1593) & (g1605) & (g1620) & (!sk[99]) & (g52)) + ((g1592) & (g1593) & (g1605) & (g1620) & (sk[99]) & (g52)));
	assign g1826 = (((!sk[100]) & (!g132) & (!g1812) & (!g1824) & (g1825)) + ((!sk[100]) & (!g132) & (!g1812) & (g1824) & (!g1825)) + ((!sk[100]) & (!g132) & (!g1812) & (g1824) & (g1825)) + ((!sk[100]) & (!g132) & (g1812) & (!g1824) & (!g1825)) + ((!sk[100]) & (!g132) & (g1812) & (!g1824) & (g1825)) + ((!sk[100]) & (!g132) & (g1812) & (g1824) & (!g1825)) + ((!sk[100]) & (!g132) & (g1812) & (g1824) & (g1825)) + ((!sk[100]) & (g132) & (!g1812) & (!g1824) & (g1825)) + ((!sk[100]) & (g132) & (!g1812) & (g1824) & (!g1825)) + ((!sk[100]) & (g132) & (!g1812) & (g1824) & (g1825)) + ((!sk[100]) & (g132) & (g1812) & (!g1824) & (!g1825)) + ((!sk[100]) & (g132) & (g1812) & (!g1824) & (g1825)) + ((!sk[100]) & (g132) & (g1812) & (g1824) & (!g1825)) + ((!sk[100]) & (g132) & (g1812) & (g1824) & (g1825)) + ((sk[100]) & (!g132) & (g1812) & (!g1824) & (g1825)) + ((sk[100]) & (!g132) & (g1812) & (g1824) & (g1825)) + ((sk[100]) & (g132) & (g1812) & (g1824) & (!g1825)) + ((sk[100]) & (g132) & (g1812) & (g1824) & (g1825)));
	assign g1827 = (((!g963) & (!g964) & (!g965) & (g966) & (g820) & (g773)) + ((!g963) & (!g964) & (g965) & (!g966) & (!g820) & (g773)) + ((!g963) & (!g964) & (g965) & (g966) & (!g820) & (g773)) + ((!g963) & (!g964) & (g965) & (g966) & (g820) & (g773)) + ((!g963) & (g964) & (!g965) & (!g966) & (g820) & (!g773)) + ((!g963) & (g964) & (!g965) & (g966) & (g820) & (!g773)) + ((!g963) & (g964) & (!g965) & (g966) & (g820) & (g773)) + ((!g963) & (g964) & (g965) & (!g966) & (!g820) & (g773)) + ((!g963) & (g964) & (g965) & (!g966) & (g820) & (!g773)) + ((!g963) & (g964) & (g965) & (g966) & (!g820) & (g773)) + ((!g963) & (g964) & (g965) & (g966) & (g820) & (!g773)) + ((!g963) & (g964) & (g965) & (g966) & (g820) & (g773)) + ((g963) & (!g964) & (!g965) & (!g966) & (!g820) & (!g773)) + ((g963) & (!g964) & (!g965) & (g966) & (!g820) & (!g773)) + ((g963) & (!g964) & (!g965) & (g966) & (g820) & (g773)) + ((g963) & (!g964) & (g965) & (!g966) & (!g820) & (!g773)) + ((g963) & (!g964) & (g965) & (!g966) & (!g820) & (g773)) + ((g963) & (!g964) & (g965) & (g966) & (!g820) & (!g773)) + ((g963) & (!g964) & (g965) & (g966) & (!g820) & (g773)) + ((g963) & (!g964) & (g965) & (g966) & (g820) & (g773)) + ((g963) & (g964) & (!g965) & (!g966) & (!g820) & (!g773)) + ((g963) & (g964) & (!g965) & (!g966) & (g820) & (!g773)) + ((g963) & (g964) & (!g965) & (g966) & (!g820) & (!g773)) + ((g963) & (g964) & (!g965) & (g966) & (g820) & (!g773)) + ((g963) & (g964) & (!g965) & (g966) & (g820) & (g773)) + ((g963) & (g964) & (g965) & (!g966) & (!g820) & (!g773)) + ((g963) & (g964) & (g965) & (!g966) & (!g820) & (g773)) + ((g963) & (g964) & (g965) & (!g966) & (g820) & (!g773)) + ((g963) & (g964) & (g965) & (g966) & (!g820) & (!g773)) + ((g963) & (g964) & (g965) & (g966) & (!g820) & (g773)) + ((g963) & (g964) & (g965) & (g966) & (g820) & (!g773)) + ((g963) & (g964) & (g965) & (g966) & (g820) & (g773)));
	assign g1828 = (((!g968) & (!g969) & (!g970) & (g971) & (g820) & (g773)) + ((!g968) & (!g969) & (g970) & (!g971) & (!g820) & (g773)) + ((!g968) & (!g969) & (g970) & (g971) & (!g820) & (g773)) + ((!g968) & (!g969) & (g970) & (g971) & (g820) & (g773)) + ((!g968) & (g969) & (!g970) & (!g971) & (g820) & (!g773)) + ((!g968) & (g969) & (!g970) & (g971) & (g820) & (!g773)) + ((!g968) & (g969) & (!g970) & (g971) & (g820) & (g773)) + ((!g968) & (g969) & (g970) & (!g971) & (!g820) & (g773)) + ((!g968) & (g969) & (g970) & (!g971) & (g820) & (!g773)) + ((!g968) & (g969) & (g970) & (g971) & (!g820) & (g773)) + ((!g968) & (g969) & (g970) & (g971) & (g820) & (!g773)) + ((!g968) & (g969) & (g970) & (g971) & (g820) & (g773)) + ((g968) & (!g969) & (!g970) & (!g971) & (!g820) & (!g773)) + ((g968) & (!g969) & (!g970) & (g971) & (!g820) & (!g773)) + ((g968) & (!g969) & (!g970) & (g971) & (g820) & (g773)) + ((g968) & (!g969) & (g970) & (!g971) & (!g820) & (!g773)) + ((g968) & (!g969) & (g970) & (!g971) & (!g820) & (g773)) + ((g968) & (!g969) & (g970) & (g971) & (!g820) & (!g773)) + ((g968) & (!g969) & (g970) & (g971) & (!g820) & (g773)) + ((g968) & (!g969) & (g970) & (g971) & (g820) & (g773)) + ((g968) & (g969) & (!g970) & (!g971) & (!g820) & (!g773)) + ((g968) & (g969) & (!g970) & (!g971) & (g820) & (!g773)) + ((g968) & (g969) & (!g970) & (g971) & (!g820) & (!g773)) + ((g968) & (g969) & (!g970) & (g971) & (g820) & (!g773)) + ((g968) & (g969) & (!g970) & (g971) & (g820) & (g773)) + ((g968) & (g969) & (g970) & (!g971) & (!g820) & (!g773)) + ((g968) & (g969) & (g970) & (!g971) & (!g820) & (g773)) + ((g968) & (g969) & (g970) & (!g971) & (g820) & (!g773)) + ((g968) & (g969) & (g970) & (g971) & (!g820) & (!g773)) + ((g968) & (g969) & (g970) & (g971) & (!g820) & (g773)) + ((g968) & (g969) & (g970) & (g971) & (g820) & (!g773)) + ((g968) & (g969) & (g970) & (g971) & (g820) & (g773)));
	assign g1829 = (((!g973) & (!g974) & (!g975) & (g976) & (g820) & (g773)) + ((!g973) & (!g974) & (g975) & (!g976) & (!g820) & (g773)) + ((!g973) & (!g974) & (g975) & (g976) & (!g820) & (g773)) + ((!g973) & (!g974) & (g975) & (g976) & (g820) & (g773)) + ((!g973) & (g974) & (!g975) & (!g976) & (g820) & (!g773)) + ((!g973) & (g974) & (!g975) & (g976) & (g820) & (!g773)) + ((!g973) & (g974) & (!g975) & (g976) & (g820) & (g773)) + ((!g973) & (g974) & (g975) & (!g976) & (!g820) & (g773)) + ((!g973) & (g974) & (g975) & (!g976) & (g820) & (!g773)) + ((!g973) & (g974) & (g975) & (g976) & (!g820) & (g773)) + ((!g973) & (g974) & (g975) & (g976) & (g820) & (!g773)) + ((!g973) & (g974) & (g975) & (g976) & (g820) & (g773)) + ((g973) & (!g974) & (!g975) & (!g976) & (!g820) & (!g773)) + ((g973) & (!g974) & (!g975) & (g976) & (!g820) & (!g773)) + ((g973) & (!g974) & (!g975) & (g976) & (g820) & (g773)) + ((g973) & (!g974) & (g975) & (!g976) & (!g820) & (!g773)) + ((g973) & (!g974) & (g975) & (!g976) & (!g820) & (g773)) + ((g973) & (!g974) & (g975) & (g976) & (!g820) & (!g773)) + ((g973) & (!g974) & (g975) & (g976) & (!g820) & (g773)) + ((g973) & (!g974) & (g975) & (g976) & (g820) & (g773)) + ((g973) & (g974) & (!g975) & (!g976) & (!g820) & (!g773)) + ((g973) & (g974) & (!g975) & (!g976) & (g820) & (!g773)) + ((g973) & (g974) & (!g975) & (g976) & (!g820) & (!g773)) + ((g973) & (g974) & (!g975) & (g976) & (g820) & (!g773)) + ((g973) & (g974) & (!g975) & (g976) & (g820) & (g773)) + ((g973) & (g974) & (g975) & (!g976) & (!g820) & (!g773)) + ((g973) & (g974) & (g975) & (!g976) & (!g820) & (g773)) + ((g973) & (g974) & (g975) & (!g976) & (g820) & (!g773)) + ((g973) & (g974) & (g975) & (g976) & (!g820) & (!g773)) + ((g973) & (g974) & (g975) & (g976) & (!g820) & (g773)) + ((g973) & (g974) & (g975) & (g976) & (g820) & (!g773)) + ((g973) & (g974) & (g975) & (g976) & (g820) & (g773)));
	assign g1830 = (((!g978) & (!g979) & (!g980) & (g981) & (g820) & (g773)) + ((!g978) & (!g979) & (g980) & (!g981) & (!g820) & (g773)) + ((!g978) & (!g979) & (g980) & (g981) & (!g820) & (g773)) + ((!g978) & (!g979) & (g980) & (g981) & (g820) & (g773)) + ((!g978) & (g979) & (!g980) & (!g981) & (g820) & (!g773)) + ((!g978) & (g979) & (!g980) & (g981) & (g820) & (!g773)) + ((!g978) & (g979) & (!g980) & (g981) & (g820) & (g773)) + ((!g978) & (g979) & (g980) & (!g981) & (!g820) & (g773)) + ((!g978) & (g979) & (g980) & (!g981) & (g820) & (!g773)) + ((!g978) & (g979) & (g980) & (g981) & (!g820) & (g773)) + ((!g978) & (g979) & (g980) & (g981) & (g820) & (!g773)) + ((!g978) & (g979) & (g980) & (g981) & (g820) & (g773)) + ((g978) & (!g979) & (!g980) & (!g981) & (!g820) & (!g773)) + ((g978) & (!g979) & (!g980) & (g981) & (!g820) & (!g773)) + ((g978) & (!g979) & (!g980) & (g981) & (g820) & (g773)) + ((g978) & (!g979) & (g980) & (!g981) & (!g820) & (!g773)) + ((g978) & (!g979) & (g980) & (!g981) & (!g820) & (g773)) + ((g978) & (!g979) & (g980) & (g981) & (!g820) & (!g773)) + ((g978) & (!g979) & (g980) & (g981) & (!g820) & (g773)) + ((g978) & (!g979) & (g980) & (g981) & (g820) & (g773)) + ((g978) & (g979) & (!g980) & (!g981) & (!g820) & (!g773)) + ((g978) & (g979) & (!g980) & (!g981) & (g820) & (!g773)) + ((g978) & (g979) & (!g980) & (g981) & (!g820) & (!g773)) + ((g978) & (g979) & (!g980) & (g981) & (g820) & (!g773)) + ((g978) & (g979) & (!g980) & (g981) & (g820) & (g773)) + ((g978) & (g979) & (g980) & (!g981) & (!g820) & (!g773)) + ((g978) & (g979) & (g980) & (!g981) & (!g820) & (g773)) + ((g978) & (g979) & (g980) & (!g981) & (g820) & (!g773)) + ((g978) & (g979) & (g980) & (g981) & (!g820) & (!g773)) + ((g978) & (g979) & (g980) & (g981) & (!g820) & (g773)) + ((g978) & (g979) & (g980) & (g981) & (g820) & (!g773)) + ((g978) & (g979) & (g980) & (g981) & (g820) & (g773)));
	assign g1831 = (((!g1827) & (!g1828) & (!g1829) & (g1830) & (g677) & (g726)) + ((!g1827) & (!g1828) & (g1829) & (!g1830) & (!g677) & (g726)) + ((!g1827) & (!g1828) & (g1829) & (g1830) & (!g677) & (g726)) + ((!g1827) & (!g1828) & (g1829) & (g1830) & (g677) & (g726)) + ((!g1827) & (g1828) & (!g1829) & (!g1830) & (g677) & (!g726)) + ((!g1827) & (g1828) & (!g1829) & (g1830) & (g677) & (!g726)) + ((!g1827) & (g1828) & (!g1829) & (g1830) & (g677) & (g726)) + ((!g1827) & (g1828) & (g1829) & (!g1830) & (!g677) & (g726)) + ((!g1827) & (g1828) & (g1829) & (!g1830) & (g677) & (!g726)) + ((!g1827) & (g1828) & (g1829) & (g1830) & (!g677) & (g726)) + ((!g1827) & (g1828) & (g1829) & (g1830) & (g677) & (!g726)) + ((!g1827) & (g1828) & (g1829) & (g1830) & (g677) & (g726)) + ((g1827) & (!g1828) & (!g1829) & (!g1830) & (!g677) & (!g726)) + ((g1827) & (!g1828) & (!g1829) & (g1830) & (!g677) & (!g726)) + ((g1827) & (!g1828) & (!g1829) & (g1830) & (g677) & (g726)) + ((g1827) & (!g1828) & (g1829) & (!g1830) & (!g677) & (!g726)) + ((g1827) & (!g1828) & (g1829) & (!g1830) & (!g677) & (g726)) + ((g1827) & (!g1828) & (g1829) & (g1830) & (!g677) & (!g726)) + ((g1827) & (!g1828) & (g1829) & (g1830) & (!g677) & (g726)) + ((g1827) & (!g1828) & (g1829) & (g1830) & (g677) & (g726)) + ((g1827) & (g1828) & (!g1829) & (!g1830) & (!g677) & (!g726)) + ((g1827) & (g1828) & (!g1829) & (!g1830) & (g677) & (!g726)) + ((g1827) & (g1828) & (!g1829) & (g1830) & (!g677) & (!g726)) + ((g1827) & (g1828) & (!g1829) & (g1830) & (g677) & (!g726)) + ((g1827) & (g1828) & (!g1829) & (g1830) & (g677) & (g726)) + ((g1827) & (g1828) & (g1829) & (!g1830) & (!g677) & (!g726)) + ((g1827) & (g1828) & (g1829) & (!g1830) & (!g677) & (g726)) + ((g1827) & (g1828) & (g1829) & (!g1830) & (g677) & (!g726)) + ((g1827) & (g1828) & (g1829) & (g1830) & (!g677) & (!g726)) + ((g1827) & (g1828) & (g1829) & (g1830) & (!g677) & (g726)) + ((g1827) & (g1828) & (g1829) & (g1830) & (g677) & (!g726)) + ((g1827) & (g1828) & (g1829) & (g1830) & (g677) & (g726)));
	assign g1832 = (((!g984) & (!g985) & (!g986) & (g987) & (g677) & (g726)) + ((!g984) & (!g985) & (g986) & (!g987) & (!g677) & (g726)) + ((!g984) & (!g985) & (g986) & (g987) & (!g677) & (g726)) + ((!g984) & (!g985) & (g986) & (g987) & (g677) & (g726)) + ((!g984) & (g985) & (!g986) & (!g987) & (g677) & (!g726)) + ((!g984) & (g985) & (!g986) & (g987) & (g677) & (!g726)) + ((!g984) & (g985) & (!g986) & (g987) & (g677) & (g726)) + ((!g984) & (g985) & (g986) & (!g987) & (!g677) & (g726)) + ((!g984) & (g985) & (g986) & (!g987) & (g677) & (!g726)) + ((!g984) & (g985) & (g986) & (g987) & (!g677) & (g726)) + ((!g984) & (g985) & (g986) & (g987) & (g677) & (!g726)) + ((!g984) & (g985) & (g986) & (g987) & (g677) & (g726)) + ((g984) & (!g985) & (!g986) & (!g987) & (!g677) & (!g726)) + ((g984) & (!g985) & (!g986) & (g987) & (!g677) & (!g726)) + ((g984) & (!g985) & (!g986) & (g987) & (g677) & (g726)) + ((g984) & (!g985) & (g986) & (!g987) & (!g677) & (!g726)) + ((g984) & (!g985) & (g986) & (!g987) & (!g677) & (g726)) + ((g984) & (!g985) & (g986) & (g987) & (!g677) & (!g726)) + ((g984) & (!g985) & (g986) & (g987) & (!g677) & (g726)) + ((g984) & (!g985) & (g986) & (g987) & (g677) & (g726)) + ((g984) & (g985) & (!g986) & (!g987) & (!g677) & (!g726)) + ((g984) & (g985) & (!g986) & (!g987) & (g677) & (!g726)) + ((g984) & (g985) & (!g986) & (g987) & (!g677) & (!g726)) + ((g984) & (g985) & (!g986) & (g987) & (g677) & (!g726)) + ((g984) & (g985) & (!g986) & (g987) & (g677) & (g726)) + ((g984) & (g985) & (g986) & (!g987) & (!g677) & (!g726)) + ((g984) & (g985) & (g986) & (!g987) & (!g677) & (g726)) + ((g984) & (g985) & (g986) & (!g987) & (g677) & (!g726)) + ((g984) & (g985) & (g986) & (g987) & (!g677) & (!g726)) + ((g984) & (g985) & (g986) & (g987) & (!g677) & (g726)) + ((g984) & (g985) & (g986) & (g987) & (g677) & (!g726)) + ((g984) & (g985) & (g986) & (g987) & (g677) & (g726)));
	assign g1833 = (((!g677) & (!g726) & (!sk[107]) & (!g989) & (g990) & (!g991)) + ((!g677) & (!g726) & (!sk[107]) & (!g989) & (g990) & (g991)) + ((!g677) & (!g726) & (!sk[107]) & (g989) & (!g990) & (!g991)) + ((!g677) & (!g726) & (!sk[107]) & (g989) & (!g990) & (g991)) + ((!g677) & (!g726) & (!sk[107]) & (g989) & (g990) & (!g991)) + ((!g677) & (!g726) & (!sk[107]) & (g989) & (g990) & (g991)) + ((!g677) & (g726) & (!sk[107]) & (!g989) & (!g990) & (!g991)) + ((!g677) & (g726) & (!sk[107]) & (!g989) & (!g990) & (g991)) + ((!g677) & (g726) & (!sk[107]) & (!g989) & (g990) & (!g991)) + ((!g677) & (g726) & (!sk[107]) & (!g989) & (g990) & (g991)) + ((!g677) & (g726) & (!sk[107]) & (g989) & (!g990) & (!g991)) + ((!g677) & (g726) & (!sk[107]) & (g989) & (!g990) & (g991)) + ((!g677) & (g726) & (!sk[107]) & (g989) & (g990) & (!g991)) + ((!g677) & (g726) & (!sk[107]) & (g989) & (g990) & (g991)) + ((!g677) & (g726) & (sk[107]) & (!g989) & (!g990) & (g991)) + ((!g677) & (g726) & (sk[107]) & (!g989) & (g990) & (g991)) + ((!g677) & (g726) & (sk[107]) & (g989) & (!g990) & (g991)) + ((!g677) & (g726) & (sk[107]) & (g989) & (g990) & (g991)) + ((g677) & (!g726) & (!sk[107]) & (!g989) & (g990) & (!g991)) + ((g677) & (!g726) & (!sk[107]) & (!g989) & (g990) & (g991)) + ((g677) & (!g726) & (!sk[107]) & (g989) & (!g990) & (!g991)) + ((g677) & (!g726) & (!sk[107]) & (g989) & (!g990) & (g991)) + ((g677) & (!g726) & (!sk[107]) & (g989) & (g990) & (!g991)) + ((g677) & (!g726) & (!sk[107]) & (g989) & (g990) & (g991)) + ((g677) & (!g726) & (sk[107]) & (g989) & (!g990) & (!g991)) + ((g677) & (!g726) & (sk[107]) & (g989) & (!g990) & (g991)) + ((g677) & (!g726) & (sk[107]) & (g989) & (g990) & (!g991)) + ((g677) & (!g726) & (sk[107]) & (g989) & (g990) & (g991)) + ((g677) & (g726) & (!sk[107]) & (!g989) & (!g990) & (!g991)) + ((g677) & (g726) & (!sk[107]) & (!g989) & (!g990) & (g991)) + ((g677) & (g726) & (!sk[107]) & (!g989) & (g990) & (!g991)) + ((g677) & (g726) & (!sk[107]) & (!g989) & (g990) & (g991)) + ((g677) & (g726) & (!sk[107]) & (g989) & (!g990) & (!g991)) + ((g677) & (g726) & (!sk[107]) & (g989) & (!g990) & (g991)) + ((g677) & (g726) & (!sk[107]) & (g989) & (g990) & (!g991)) + ((g677) & (g726) & (!sk[107]) & (g989) & (g990) & (g991)) + ((g677) & (g726) & (sk[107]) & (!g989) & (g990) & (!g991)) + ((g677) & (g726) & (sk[107]) & (!g989) & (g990) & (g991)) + ((g677) & (g726) & (sk[107]) & (g989) & (g990) & (!g991)) + ((g677) & (g726) & (sk[107]) & (g989) & (g990) & (g991)));
	assign g1834 = (((!g993) & (!g994) & (!g995) & (g996) & (g677) & (g726)) + ((!g993) & (!g994) & (g995) & (!g996) & (!g677) & (g726)) + ((!g993) & (!g994) & (g995) & (g996) & (!g677) & (g726)) + ((!g993) & (!g994) & (g995) & (g996) & (g677) & (g726)) + ((!g993) & (g994) & (!g995) & (!g996) & (g677) & (!g726)) + ((!g993) & (g994) & (!g995) & (g996) & (g677) & (!g726)) + ((!g993) & (g994) & (!g995) & (g996) & (g677) & (g726)) + ((!g993) & (g994) & (g995) & (!g996) & (!g677) & (g726)) + ((!g993) & (g994) & (g995) & (!g996) & (g677) & (!g726)) + ((!g993) & (g994) & (g995) & (g996) & (!g677) & (g726)) + ((!g993) & (g994) & (g995) & (g996) & (g677) & (!g726)) + ((!g993) & (g994) & (g995) & (g996) & (g677) & (g726)) + ((g993) & (!g994) & (!g995) & (!g996) & (!g677) & (!g726)) + ((g993) & (!g994) & (!g995) & (g996) & (!g677) & (!g726)) + ((g993) & (!g994) & (!g995) & (g996) & (g677) & (g726)) + ((g993) & (!g994) & (g995) & (!g996) & (!g677) & (!g726)) + ((g993) & (!g994) & (g995) & (!g996) & (!g677) & (g726)) + ((g993) & (!g994) & (g995) & (g996) & (!g677) & (!g726)) + ((g993) & (!g994) & (g995) & (g996) & (!g677) & (g726)) + ((g993) & (!g994) & (g995) & (g996) & (g677) & (g726)) + ((g993) & (g994) & (!g995) & (!g996) & (!g677) & (!g726)) + ((g993) & (g994) & (!g995) & (!g996) & (g677) & (!g726)) + ((g993) & (g994) & (!g995) & (g996) & (!g677) & (!g726)) + ((g993) & (g994) & (!g995) & (g996) & (g677) & (!g726)) + ((g993) & (g994) & (!g995) & (g996) & (g677) & (g726)) + ((g993) & (g994) & (g995) & (!g996) & (!g677) & (!g726)) + ((g993) & (g994) & (g995) & (!g996) & (!g677) & (g726)) + ((g993) & (g994) & (g995) & (!g996) & (g677) & (!g726)) + ((g993) & (g994) & (g995) & (g996) & (!g677) & (!g726)) + ((g993) & (g994) & (g995) & (g996) & (!g677) & (g726)) + ((g993) & (g994) & (g995) & (g996) & (g677) & (!g726)) + ((g993) & (g994) & (g995) & (g996) & (g677) & (g726)));
	assign g1835 = (((!g998) & (!g999) & (!g1000) & (g1001) & (g677) & (g726)) + ((!g998) & (!g999) & (g1000) & (!g1001) & (!g677) & (g726)) + ((!g998) & (!g999) & (g1000) & (g1001) & (!g677) & (g726)) + ((!g998) & (!g999) & (g1000) & (g1001) & (g677) & (g726)) + ((!g998) & (g999) & (!g1000) & (!g1001) & (g677) & (!g726)) + ((!g998) & (g999) & (!g1000) & (g1001) & (g677) & (!g726)) + ((!g998) & (g999) & (!g1000) & (g1001) & (g677) & (g726)) + ((!g998) & (g999) & (g1000) & (!g1001) & (!g677) & (g726)) + ((!g998) & (g999) & (g1000) & (!g1001) & (g677) & (!g726)) + ((!g998) & (g999) & (g1000) & (g1001) & (!g677) & (g726)) + ((!g998) & (g999) & (g1000) & (g1001) & (g677) & (!g726)) + ((!g998) & (g999) & (g1000) & (g1001) & (g677) & (g726)) + ((g998) & (!g999) & (!g1000) & (!g1001) & (!g677) & (!g726)) + ((g998) & (!g999) & (!g1000) & (g1001) & (!g677) & (!g726)) + ((g998) & (!g999) & (!g1000) & (g1001) & (g677) & (g726)) + ((g998) & (!g999) & (g1000) & (!g1001) & (!g677) & (!g726)) + ((g998) & (!g999) & (g1000) & (!g1001) & (!g677) & (g726)) + ((g998) & (!g999) & (g1000) & (g1001) & (!g677) & (!g726)) + ((g998) & (!g999) & (g1000) & (g1001) & (!g677) & (g726)) + ((g998) & (!g999) & (g1000) & (g1001) & (g677) & (g726)) + ((g998) & (g999) & (!g1000) & (!g1001) & (!g677) & (!g726)) + ((g998) & (g999) & (!g1000) & (!g1001) & (g677) & (!g726)) + ((g998) & (g999) & (!g1000) & (g1001) & (!g677) & (!g726)) + ((g998) & (g999) & (!g1000) & (g1001) & (g677) & (!g726)) + ((g998) & (g999) & (!g1000) & (g1001) & (g677) & (g726)) + ((g998) & (g999) & (g1000) & (!g1001) & (!g677) & (!g726)) + ((g998) & (g999) & (g1000) & (!g1001) & (!g677) & (g726)) + ((g998) & (g999) & (g1000) & (!g1001) & (g677) & (!g726)) + ((g998) & (g999) & (g1000) & (g1001) & (!g677) & (!g726)) + ((g998) & (g999) & (g1000) & (g1001) & (!g677) & (g726)) + ((g998) & (g999) & (g1000) & (g1001) & (g677) & (!g726)) + ((g998) & (g999) & (g1000) & (g1001) & (g677) & (g726)));
	assign g1836 = (((!g820) & (!g773) & (!g1832) & (g1833) & (!g1834) & (!g1835)) + ((!g820) & (!g773) & (!g1832) & (g1833) & (!g1834) & (g1835)) + ((!g820) & (!g773) & (!g1832) & (g1833) & (g1834) & (!g1835)) + ((!g820) & (!g773) & (!g1832) & (g1833) & (g1834) & (g1835)) + ((!g820) & (!g773) & (g1832) & (g1833) & (!g1834) & (!g1835)) + ((!g820) & (!g773) & (g1832) & (g1833) & (!g1834) & (g1835)) + ((!g820) & (!g773) & (g1832) & (g1833) & (g1834) & (!g1835)) + ((!g820) & (!g773) & (g1832) & (g1833) & (g1834) & (g1835)) + ((!g820) & (g773) & (!g1832) & (!g1833) & (!g1834) & (g1835)) + ((!g820) & (g773) & (!g1832) & (!g1833) & (g1834) & (g1835)) + ((!g820) & (g773) & (!g1832) & (g1833) & (!g1834) & (g1835)) + ((!g820) & (g773) & (!g1832) & (g1833) & (g1834) & (g1835)) + ((!g820) & (g773) & (g1832) & (!g1833) & (!g1834) & (g1835)) + ((!g820) & (g773) & (g1832) & (!g1833) & (g1834) & (g1835)) + ((!g820) & (g773) & (g1832) & (g1833) & (!g1834) & (g1835)) + ((!g820) & (g773) & (g1832) & (g1833) & (g1834) & (g1835)) + ((g820) & (!g773) & (g1832) & (!g1833) & (!g1834) & (!g1835)) + ((g820) & (!g773) & (g1832) & (!g1833) & (!g1834) & (g1835)) + ((g820) & (!g773) & (g1832) & (!g1833) & (g1834) & (!g1835)) + ((g820) & (!g773) & (g1832) & (!g1833) & (g1834) & (g1835)) + ((g820) & (!g773) & (g1832) & (g1833) & (!g1834) & (!g1835)) + ((g820) & (!g773) & (g1832) & (g1833) & (!g1834) & (g1835)) + ((g820) & (!g773) & (g1832) & (g1833) & (g1834) & (!g1835)) + ((g820) & (!g773) & (g1832) & (g1833) & (g1834) & (g1835)) + ((g820) & (g773) & (!g1832) & (!g1833) & (g1834) & (!g1835)) + ((g820) & (g773) & (!g1832) & (!g1833) & (g1834) & (g1835)) + ((g820) & (g773) & (!g1832) & (g1833) & (g1834) & (!g1835)) + ((g820) & (g773) & (!g1832) & (g1833) & (g1834) & (g1835)) + ((g820) & (g773) & (g1832) & (!g1833) & (g1834) & (!g1835)) + ((g820) & (g773) & (g1832) & (!g1833) & (g1834) & (g1835)) + ((g820) & (g773) & (g1832) & (g1833) & (g1834) & (!g1835)) + ((g820) & (g773) & (g1832) & (g1833) & (g1834) & (g1835)));
	assign g1837 = (((!sk[111]) & (!g867) & (!g1831) & (g1836)) + ((!sk[111]) & (!g867) & (g1831) & (!g1836)) + ((!sk[111]) & (!g867) & (g1831) & (g1836)) + ((!sk[111]) & (g867) & (!g1831) & (g1836)) + ((!sk[111]) & (g867) & (g1831) & (!g1836)) + ((!sk[111]) & (g867) & (g1831) & (g1836)) + ((sk[111]) & (!g867) & (!g1831) & (g1836)) + ((sk[111]) & (!g867) & (g1831) & (g1836)) + ((sk[111]) & (g867) & (g1831) & (!g1836)) + ((sk[111]) & (g867) & (g1831) & (g1836)));
	assign g1838 = (((!g1592) & (!sk[112]) & (!g1593) & (!g1605) & (g1632) & (!g53)) + ((!g1592) & (!sk[112]) & (!g1593) & (!g1605) & (g1632) & (g53)) + ((!g1592) & (!sk[112]) & (!g1593) & (g1605) & (!g1632) & (!g53)) + ((!g1592) & (!sk[112]) & (!g1593) & (g1605) & (!g1632) & (g53)) + ((!g1592) & (!sk[112]) & (!g1593) & (g1605) & (g1632) & (!g53)) + ((!g1592) & (!sk[112]) & (!g1593) & (g1605) & (g1632) & (g53)) + ((!g1592) & (!sk[112]) & (g1593) & (!g1605) & (!g1632) & (!g53)) + ((!g1592) & (!sk[112]) & (g1593) & (!g1605) & (!g1632) & (g53)) + ((!g1592) & (!sk[112]) & (g1593) & (!g1605) & (g1632) & (!g53)) + ((!g1592) & (!sk[112]) & (g1593) & (!g1605) & (g1632) & (g53)) + ((!g1592) & (!sk[112]) & (g1593) & (g1605) & (!g1632) & (!g53)) + ((!g1592) & (!sk[112]) & (g1593) & (g1605) & (!g1632) & (g53)) + ((!g1592) & (!sk[112]) & (g1593) & (g1605) & (g1632) & (!g53)) + ((!g1592) & (!sk[112]) & (g1593) & (g1605) & (g1632) & (g53)) + ((!g1592) & (sk[112]) & (!g1593) & (!g1605) & (g1632) & (!g53)) + ((!g1592) & (sk[112]) & (!g1593) & (!g1605) & (g1632) & (g53)) + ((!g1592) & (sk[112]) & (!g1593) & (g1605) & (g1632) & (!g53)) + ((!g1592) & (sk[112]) & (!g1593) & (g1605) & (g1632) & (g53)) + ((!g1592) & (sk[112]) & (g1593) & (!g1605) & (g1632) & (!g53)) + ((!g1592) & (sk[112]) & (g1593) & (!g1605) & (g1632) & (g53)) + ((!g1592) & (sk[112]) & (g1593) & (g1605) & (g1632) & (!g53)) + ((!g1592) & (sk[112]) & (g1593) & (g1605) & (g1632) & (g53)) + ((g1592) & (!sk[112]) & (!g1593) & (!g1605) & (g1632) & (!g53)) + ((g1592) & (!sk[112]) & (!g1593) & (!g1605) & (g1632) & (g53)) + ((g1592) & (!sk[112]) & (!g1593) & (g1605) & (!g1632) & (!g53)) + ((g1592) & (!sk[112]) & (!g1593) & (g1605) & (!g1632) & (g53)) + ((g1592) & (!sk[112]) & (!g1593) & (g1605) & (g1632) & (!g53)) + ((g1592) & (!sk[112]) & (!g1593) & (g1605) & (g1632) & (g53)) + ((g1592) & (!sk[112]) & (g1593) & (!g1605) & (!g1632) & (!g53)) + ((g1592) & (!sk[112]) & (g1593) & (!g1605) & (!g1632) & (g53)) + ((g1592) & (!sk[112]) & (g1593) & (!g1605) & (g1632) & (!g53)) + ((g1592) & (!sk[112]) & (g1593) & (!g1605) & (g1632) & (g53)) + ((g1592) & (!sk[112]) & (g1593) & (g1605) & (!g1632) & (!g53)) + ((g1592) & (!sk[112]) & (g1593) & (g1605) & (!g1632) & (g53)) + ((g1592) & (!sk[112]) & (g1593) & (g1605) & (g1632) & (!g53)) + ((g1592) & (!sk[112]) & (g1593) & (g1605) & (g1632) & (g53)) + ((g1592) & (sk[112]) & (!g1593) & (!g1605) & (g1632) & (!g53)) + ((g1592) & (sk[112]) & (!g1593) & (!g1605) & (g1632) & (g53)) + ((g1592) & (sk[112]) & (g1593) & (!g1605) & (!g1632) & (g53)) + ((g1592) & (sk[112]) & (g1593) & (!g1605) & (g1632) & (g53)) + ((g1592) & (sk[112]) & (g1593) & (g1605) & (!g1632) & (g53)) + ((g1592) & (sk[112]) & (g1593) & (g1605) & (g1632) & (g53)));
	assign g1839 = (((!g132) & (!g1812) & (!sk[113]) & (!g1837) & (g1838)) + ((!g132) & (!g1812) & (!sk[113]) & (g1837) & (!g1838)) + ((!g132) & (!g1812) & (!sk[113]) & (g1837) & (g1838)) + ((!g132) & (g1812) & (!sk[113]) & (!g1837) & (!g1838)) + ((!g132) & (g1812) & (!sk[113]) & (!g1837) & (g1838)) + ((!g132) & (g1812) & (!sk[113]) & (g1837) & (!g1838)) + ((!g132) & (g1812) & (!sk[113]) & (g1837) & (g1838)) + ((!g132) & (g1812) & (sk[113]) & (!g1837) & (g1838)) + ((!g132) & (g1812) & (sk[113]) & (g1837) & (g1838)) + ((g132) & (!g1812) & (!sk[113]) & (!g1837) & (g1838)) + ((g132) & (!g1812) & (!sk[113]) & (g1837) & (!g1838)) + ((g132) & (!g1812) & (!sk[113]) & (g1837) & (g1838)) + ((g132) & (g1812) & (!sk[113]) & (!g1837) & (!g1838)) + ((g132) & (g1812) & (!sk[113]) & (!g1837) & (g1838)) + ((g132) & (g1812) & (!sk[113]) & (g1837) & (!g1838)) + ((g132) & (g1812) & (!sk[113]) & (g1837) & (g1838)) + ((g132) & (g1812) & (sk[113]) & (g1837) & (!g1838)) + ((g132) & (g1812) & (sk[113]) & (g1837) & (g1838)));
	assign g1840 = (((!g1008) & (!g1009) & (!g1010) & (g1011) & (g820) & (g773)) + ((!g1008) & (!g1009) & (g1010) & (!g1011) & (!g820) & (g773)) + ((!g1008) & (!g1009) & (g1010) & (g1011) & (!g820) & (g773)) + ((!g1008) & (!g1009) & (g1010) & (g1011) & (g820) & (g773)) + ((!g1008) & (g1009) & (!g1010) & (!g1011) & (g820) & (!g773)) + ((!g1008) & (g1009) & (!g1010) & (g1011) & (g820) & (!g773)) + ((!g1008) & (g1009) & (!g1010) & (g1011) & (g820) & (g773)) + ((!g1008) & (g1009) & (g1010) & (!g1011) & (!g820) & (g773)) + ((!g1008) & (g1009) & (g1010) & (!g1011) & (g820) & (!g773)) + ((!g1008) & (g1009) & (g1010) & (g1011) & (!g820) & (g773)) + ((!g1008) & (g1009) & (g1010) & (g1011) & (g820) & (!g773)) + ((!g1008) & (g1009) & (g1010) & (g1011) & (g820) & (g773)) + ((g1008) & (!g1009) & (!g1010) & (!g1011) & (!g820) & (!g773)) + ((g1008) & (!g1009) & (!g1010) & (g1011) & (!g820) & (!g773)) + ((g1008) & (!g1009) & (!g1010) & (g1011) & (g820) & (g773)) + ((g1008) & (!g1009) & (g1010) & (!g1011) & (!g820) & (!g773)) + ((g1008) & (!g1009) & (g1010) & (!g1011) & (!g820) & (g773)) + ((g1008) & (!g1009) & (g1010) & (g1011) & (!g820) & (!g773)) + ((g1008) & (!g1009) & (g1010) & (g1011) & (!g820) & (g773)) + ((g1008) & (!g1009) & (g1010) & (g1011) & (g820) & (g773)) + ((g1008) & (g1009) & (!g1010) & (!g1011) & (!g820) & (!g773)) + ((g1008) & (g1009) & (!g1010) & (!g1011) & (g820) & (!g773)) + ((g1008) & (g1009) & (!g1010) & (g1011) & (!g820) & (!g773)) + ((g1008) & (g1009) & (!g1010) & (g1011) & (g820) & (!g773)) + ((g1008) & (g1009) & (!g1010) & (g1011) & (g820) & (g773)) + ((g1008) & (g1009) & (g1010) & (!g1011) & (!g820) & (!g773)) + ((g1008) & (g1009) & (g1010) & (!g1011) & (!g820) & (g773)) + ((g1008) & (g1009) & (g1010) & (!g1011) & (g820) & (!g773)) + ((g1008) & (g1009) & (g1010) & (g1011) & (!g820) & (!g773)) + ((g1008) & (g1009) & (g1010) & (g1011) & (!g820) & (g773)) + ((g1008) & (g1009) & (g1010) & (g1011) & (g820) & (!g773)) + ((g1008) & (g1009) & (g1010) & (g1011) & (g820) & (g773)));
	assign g1841 = (((!g1013) & (!g1014) & (!g1015) & (g1016) & (g820) & (g773)) + ((!g1013) & (!g1014) & (g1015) & (!g1016) & (!g820) & (g773)) + ((!g1013) & (!g1014) & (g1015) & (g1016) & (!g820) & (g773)) + ((!g1013) & (!g1014) & (g1015) & (g1016) & (g820) & (g773)) + ((!g1013) & (g1014) & (!g1015) & (!g1016) & (g820) & (!g773)) + ((!g1013) & (g1014) & (!g1015) & (g1016) & (g820) & (!g773)) + ((!g1013) & (g1014) & (!g1015) & (g1016) & (g820) & (g773)) + ((!g1013) & (g1014) & (g1015) & (!g1016) & (!g820) & (g773)) + ((!g1013) & (g1014) & (g1015) & (!g1016) & (g820) & (!g773)) + ((!g1013) & (g1014) & (g1015) & (g1016) & (!g820) & (g773)) + ((!g1013) & (g1014) & (g1015) & (g1016) & (g820) & (!g773)) + ((!g1013) & (g1014) & (g1015) & (g1016) & (g820) & (g773)) + ((g1013) & (!g1014) & (!g1015) & (!g1016) & (!g820) & (!g773)) + ((g1013) & (!g1014) & (!g1015) & (g1016) & (!g820) & (!g773)) + ((g1013) & (!g1014) & (!g1015) & (g1016) & (g820) & (g773)) + ((g1013) & (!g1014) & (g1015) & (!g1016) & (!g820) & (!g773)) + ((g1013) & (!g1014) & (g1015) & (!g1016) & (!g820) & (g773)) + ((g1013) & (!g1014) & (g1015) & (g1016) & (!g820) & (!g773)) + ((g1013) & (!g1014) & (g1015) & (g1016) & (!g820) & (g773)) + ((g1013) & (!g1014) & (g1015) & (g1016) & (g820) & (g773)) + ((g1013) & (g1014) & (!g1015) & (!g1016) & (!g820) & (!g773)) + ((g1013) & (g1014) & (!g1015) & (!g1016) & (g820) & (!g773)) + ((g1013) & (g1014) & (!g1015) & (g1016) & (!g820) & (!g773)) + ((g1013) & (g1014) & (!g1015) & (g1016) & (g820) & (!g773)) + ((g1013) & (g1014) & (!g1015) & (g1016) & (g820) & (g773)) + ((g1013) & (g1014) & (g1015) & (!g1016) & (!g820) & (!g773)) + ((g1013) & (g1014) & (g1015) & (!g1016) & (!g820) & (g773)) + ((g1013) & (g1014) & (g1015) & (!g1016) & (g820) & (!g773)) + ((g1013) & (g1014) & (g1015) & (g1016) & (!g820) & (!g773)) + ((g1013) & (g1014) & (g1015) & (g1016) & (!g820) & (g773)) + ((g1013) & (g1014) & (g1015) & (g1016) & (g820) & (!g773)) + ((g1013) & (g1014) & (g1015) & (g1016) & (g820) & (g773)));
	assign g1842 = (((!g1018) & (!g1019) & (!g1020) & (g1021) & (g820) & (g773)) + ((!g1018) & (!g1019) & (g1020) & (!g1021) & (!g820) & (g773)) + ((!g1018) & (!g1019) & (g1020) & (g1021) & (!g820) & (g773)) + ((!g1018) & (!g1019) & (g1020) & (g1021) & (g820) & (g773)) + ((!g1018) & (g1019) & (!g1020) & (!g1021) & (g820) & (!g773)) + ((!g1018) & (g1019) & (!g1020) & (g1021) & (g820) & (!g773)) + ((!g1018) & (g1019) & (!g1020) & (g1021) & (g820) & (g773)) + ((!g1018) & (g1019) & (g1020) & (!g1021) & (!g820) & (g773)) + ((!g1018) & (g1019) & (g1020) & (!g1021) & (g820) & (!g773)) + ((!g1018) & (g1019) & (g1020) & (g1021) & (!g820) & (g773)) + ((!g1018) & (g1019) & (g1020) & (g1021) & (g820) & (!g773)) + ((!g1018) & (g1019) & (g1020) & (g1021) & (g820) & (g773)) + ((g1018) & (!g1019) & (!g1020) & (!g1021) & (!g820) & (!g773)) + ((g1018) & (!g1019) & (!g1020) & (g1021) & (!g820) & (!g773)) + ((g1018) & (!g1019) & (!g1020) & (g1021) & (g820) & (g773)) + ((g1018) & (!g1019) & (g1020) & (!g1021) & (!g820) & (!g773)) + ((g1018) & (!g1019) & (g1020) & (!g1021) & (!g820) & (g773)) + ((g1018) & (!g1019) & (g1020) & (g1021) & (!g820) & (!g773)) + ((g1018) & (!g1019) & (g1020) & (g1021) & (!g820) & (g773)) + ((g1018) & (!g1019) & (g1020) & (g1021) & (g820) & (g773)) + ((g1018) & (g1019) & (!g1020) & (!g1021) & (!g820) & (!g773)) + ((g1018) & (g1019) & (!g1020) & (!g1021) & (g820) & (!g773)) + ((g1018) & (g1019) & (!g1020) & (g1021) & (!g820) & (!g773)) + ((g1018) & (g1019) & (!g1020) & (g1021) & (g820) & (!g773)) + ((g1018) & (g1019) & (!g1020) & (g1021) & (g820) & (g773)) + ((g1018) & (g1019) & (g1020) & (!g1021) & (!g820) & (!g773)) + ((g1018) & (g1019) & (g1020) & (!g1021) & (!g820) & (g773)) + ((g1018) & (g1019) & (g1020) & (!g1021) & (g820) & (!g773)) + ((g1018) & (g1019) & (g1020) & (g1021) & (!g820) & (!g773)) + ((g1018) & (g1019) & (g1020) & (g1021) & (!g820) & (g773)) + ((g1018) & (g1019) & (g1020) & (g1021) & (g820) & (!g773)) + ((g1018) & (g1019) & (g1020) & (g1021) & (g820) & (g773)));
	assign g1843 = (((!g1023) & (!g1024) & (!g1025) & (g1026) & (g820) & (g773)) + ((!g1023) & (!g1024) & (g1025) & (!g1026) & (!g820) & (g773)) + ((!g1023) & (!g1024) & (g1025) & (g1026) & (!g820) & (g773)) + ((!g1023) & (!g1024) & (g1025) & (g1026) & (g820) & (g773)) + ((!g1023) & (g1024) & (!g1025) & (!g1026) & (g820) & (!g773)) + ((!g1023) & (g1024) & (!g1025) & (g1026) & (g820) & (!g773)) + ((!g1023) & (g1024) & (!g1025) & (g1026) & (g820) & (g773)) + ((!g1023) & (g1024) & (g1025) & (!g1026) & (!g820) & (g773)) + ((!g1023) & (g1024) & (g1025) & (!g1026) & (g820) & (!g773)) + ((!g1023) & (g1024) & (g1025) & (g1026) & (!g820) & (g773)) + ((!g1023) & (g1024) & (g1025) & (g1026) & (g820) & (!g773)) + ((!g1023) & (g1024) & (g1025) & (g1026) & (g820) & (g773)) + ((g1023) & (!g1024) & (!g1025) & (!g1026) & (!g820) & (!g773)) + ((g1023) & (!g1024) & (!g1025) & (g1026) & (!g820) & (!g773)) + ((g1023) & (!g1024) & (!g1025) & (g1026) & (g820) & (g773)) + ((g1023) & (!g1024) & (g1025) & (!g1026) & (!g820) & (!g773)) + ((g1023) & (!g1024) & (g1025) & (!g1026) & (!g820) & (g773)) + ((g1023) & (!g1024) & (g1025) & (g1026) & (!g820) & (!g773)) + ((g1023) & (!g1024) & (g1025) & (g1026) & (!g820) & (g773)) + ((g1023) & (!g1024) & (g1025) & (g1026) & (g820) & (g773)) + ((g1023) & (g1024) & (!g1025) & (!g1026) & (!g820) & (!g773)) + ((g1023) & (g1024) & (!g1025) & (!g1026) & (g820) & (!g773)) + ((g1023) & (g1024) & (!g1025) & (g1026) & (!g820) & (!g773)) + ((g1023) & (g1024) & (!g1025) & (g1026) & (g820) & (!g773)) + ((g1023) & (g1024) & (!g1025) & (g1026) & (g820) & (g773)) + ((g1023) & (g1024) & (g1025) & (!g1026) & (!g820) & (!g773)) + ((g1023) & (g1024) & (g1025) & (!g1026) & (!g820) & (g773)) + ((g1023) & (g1024) & (g1025) & (!g1026) & (g820) & (!g773)) + ((g1023) & (g1024) & (g1025) & (g1026) & (!g820) & (!g773)) + ((g1023) & (g1024) & (g1025) & (g1026) & (!g820) & (g773)) + ((g1023) & (g1024) & (g1025) & (g1026) & (g820) & (!g773)) + ((g1023) & (g1024) & (g1025) & (g1026) & (g820) & (g773)));
	assign g1844 = (((!g1840) & (!g1841) & (!g1842) & (g1843) & (g677) & (g726)) + ((!g1840) & (!g1841) & (g1842) & (!g1843) & (!g677) & (g726)) + ((!g1840) & (!g1841) & (g1842) & (g1843) & (!g677) & (g726)) + ((!g1840) & (!g1841) & (g1842) & (g1843) & (g677) & (g726)) + ((!g1840) & (g1841) & (!g1842) & (!g1843) & (g677) & (!g726)) + ((!g1840) & (g1841) & (!g1842) & (g1843) & (g677) & (!g726)) + ((!g1840) & (g1841) & (!g1842) & (g1843) & (g677) & (g726)) + ((!g1840) & (g1841) & (g1842) & (!g1843) & (!g677) & (g726)) + ((!g1840) & (g1841) & (g1842) & (!g1843) & (g677) & (!g726)) + ((!g1840) & (g1841) & (g1842) & (g1843) & (!g677) & (g726)) + ((!g1840) & (g1841) & (g1842) & (g1843) & (g677) & (!g726)) + ((!g1840) & (g1841) & (g1842) & (g1843) & (g677) & (g726)) + ((g1840) & (!g1841) & (!g1842) & (!g1843) & (!g677) & (!g726)) + ((g1840) & (!g1841) & (!g1842) & (g1843) & (!g677) & (!g726)) + ((g1840) & (!g1841) & (!g1842) & (g1843) & (g677) & (g726)) + ((g1840) & (!g1841) & (g1842) & (!g1843) & (!g677) & (!g726)) + ((g1840) & (!g1841) & (g1842) & (!g1843) & (!g677) & (g726)) + ((g1840) & (!g1841) & (g1842) & (g1843) & (!g677) & (!g726)) + ((g1840) & (!g1841) & (g1842) & (g1843) & (!g677) & (g726)) + ((g1840) & (!g1841) & (g1842) & (g1843) & (g677) & (g726)) + ((g1840) & (g1841) & (!g1842) & (!g1843) & (!g677) & (!g726)) + ((g1840) & (g1841) & (!g1842) & (!g1843) & (g677) & (!g726)) + ((g1840) & (g1841) & (!g1842) & (g1843) & (!g677) & (!g726)) + ((g1840) & (g1841) & (!g1842) & (g1843) & (g677) & (!g726)) + ((g1840) & (g1841) & (!g1842) & (g1843) & (g677) & (g726)) + ((g1840) & (g1841) & (g1842) & (!g1843) & (!g677) & (!g726)) + ((g1840) & (g1841) & (g1842) & (!g1843) & (!g677) & (g726)) + ((g1840) & (g1841) & (g1842) & (!g1843) & (g677) & (!g726)) + ((g1840) & (g1841) & (g1842) & (g1843) & (!g677) & (!g726)) + ((g1840) & (g1841) & (g1842) & (g1843) & (!g677) & (g726)) + ((g1840) & (g1841) & (g1842) & (g1843) & (g677) & (!g726)) + ((g1840) & (g1841) & (g1842) & (g1843) & (g677) & (g726)));
	assign g1845 = (((!g1029) & (!g1030) & (!g1031) & (g1032) & (g677) & (g726)) + ((!g1029) & (!g1030) & (g1031) & (!g1032) & (!g677) & (g726)) + ((!g1029) & (!g1030) & (g1031) & (g1032) & (!g677) & (g726)) + ((!g1029) & (!g1030) & (g1031) & (g1032) & (g677) & (g726)) + ((!g1029) & (g1030) & (!g1031) & (!g1032) & (g677) & (!g726)) + ((!g1029) & (g1030) & (!g1031) & (g1032) & (g677) & (!g726)) + ((!g1029) & (g1030) & (!g1031) & (g1032) & (g677) & (g726)) + ((!g1029) & (g1030) & (g1031) & (!g1032) & (!g677) & (g726)) + ((!g1029) & (g1030) & (g1031) & (!g1032) & (g677) & (!g726)) + ((!g1029) & (g1030) & (g1031) & (g1032) & (!g677) & (g726)) + ((!g1029) & (g1030) & (g1031) & (g1032) & (g677) & (!g726)) + ((!g1029) & (g1030) & (g1031) & (g1032) & (g677) & (g726)) + ((g1029) & (!g1030) & (!g1031) & (!g1032) & (!g677) & (!g726)) + ((g1029) & (!g1030) & (!g1031) & (g1032) & (!g677) & (!g726)) + ((g1029) & (!g1030) & (!g1031) & (g1032) & (g677) & (g726)) + ((g1029) & (!g1030) & (g1031) & (!g1032) & (!g677) & (!g726)) + ((g1029) & (!g1030) & (g1031) & (!g1032) & (!g677) & (g726)) + ((g1029) & (!g1030) & (g1031) & (g1032) & (!g677) & (!g726)) + ((g1029) & (!g1030) & (g1031) & (g1032) & (!g677) & (g726)) + ((g1029) & (!g1030) & (g1031) & (g1032) & (g677) & (g726)) + ((g1029) & (g1030) & (!g1031) & (!g1032) & (!g677) & (!g726)) + ((g1029) & (g1030) & (!g1031) & (!g1032) & (g677) & (!g726)) + ((g1029) & (g1030) & (!g1031) & (g1032) & (!g677) & (!g726)) + ((g1029) & (g1030) & (!g1031) & (g1032) & (g677) & (!g726)) + ((g1029) & (g1030) & (!g1031) & (g1032) & (g677) & (g726)) + ((g1029) & (g1030) & (g1031) & (!g1032) & (!g677) & (!g726)) + ((g1029) & (g1030) & (g1031) & (!g1032) & (!g677) & (g726)) + ((g1029) & (g1030) & (g1031) & (!g1032) & (g677) & (!g726)) + ((g1029) & (g1030) & (g1031) & (g1032) & (!g677) & (!g726)) + ((g1029) & (g1030) & (g1031) & (g1032) & (!g677) & (g726)) + ((g1029) & (g1030) & (g1031) & (g1032) & (g677) & (!g726)) + ((g1029) & (g1030) & (g1031) & (g1032) & (g677) & (g726)));
	assign g1846 = (((!sk[120]) & (!g677) & (!g726) & (!g1034) & (g1035) & (!g1036)) + ((!sk[120]) & (!g677) & (!g726) & (!g1034) & (g1035) & (g1036)) + ((!sk[120]) & (!g677) & (!g726) & (g1034) & (!g1035) & (!g1036)) + ((!sk[120]) & (!g677) & (!g726) & (g1034) & (!g1035) & (g1036)) + ((!sk[120]) & (!g677) & (!g726) & (g1034) & (g1035) & (!g1036)) + ((!sk[120]) & (!g677) & (!g726) & (g1034) & (g1035) & (g1036)) + ((!sk[120]) & (!g677) & (g726) & (!g1034) & (!g1035) & (!g1036)) + ((!sk[120]) & (!g677) & (g726) & (!g1034) & (!g1035) & (g1036)) + ((!sk[120]) & (!g677) & (g726) & (!g1034) & (g1035) & (!g1036)) + ((!sk[120]) & (!g677) & (g726) & (!g1034) & (g1035) & (g1036)) + ((!sk[120]) & (!g677) & (g726) & (g1034) & (!g1035) & (!g1036)) + ((!sk[120]) & (!g677) & (g726) & (g1034) & (!g1035) & (g1036)) + ((!sk[120]) & (!g677) & (g726) & (g1034) & (g1035) & (!g1036)) + ((!sk[120]) & (!g677) & (g726) & (g1034) & (g1035) & (g1036)) + ((!sk[120]) & (g677) & (!g726) & (!g1034) & (g1035) & (!g1036)) + ((!sk[120]) & (g677) & (!g726) & (!g1034) & (g1035) & (g1036)) + ((!sk[120]) & (g677) & (!g726) & (g1034) & (!g1035) & (!g1036)) + ((!sk[120]) & (g677) & (!g726) & (g1034) & (!g1035) & (g1036)) + ((!sk[120]) & (g677) & (!g726) & (g1034) & (g1035) & (!g1036)) + ((!sk[120]) & (g677) & (!g726) & (g1034) & (g1035) & (g1036)) + ((!sk[120]) & (g677) & (g726) & (!g1034) & (!g1035) & (!g1036)) + ((!sk[120]) & (g677) & (g726) & (!g1034) & (!g1035) & (g1036)) + ((!sk[120]) & (g677) & (g726) & (!g1034) & (g1035) & (!g1036)) + ((!sk[120]) & (g677) & (g726) & (!g1034) & (g1035) & (g1036)) + ((!sk[120]) & (g677) & (g726) & (g1034) & (!g1035) & (!g1036)) + ((!sk[120]) & (g677) & (g726) & (g1034) & (!g1035) & (g1036)) + ((!sk[120]) & (g677) & (g726) & (g1034) & (g1035) & (!g1036)) + ((!sk[120]) & (g677) & (g726) & (g1034) & (g1035) & (g1036)) + ((sk[120]) & (!g677) & (g726) & (!g1034) & (!g1035) & (g1036)) + ((sk[120]) & (!g677) & (g726) & (!g1034) & (g1035) & (g1036)) + ((sk[120]) & (!g677) & (g726) & (g1034) & (!g1035) & (g1036)) + ((sk[120]) & (!g677) & (g726) & (g1034) & (g1035) & (g1036)) + ((sk[120]) & (g677) & (!g726) & (g1034) & (!g1035) & (!g1036)) + ((sk[120]) & (g677) & (!g726) & (g1034) & (!g1035) & (g1036)) + ((sk[120]) & (g677) & (!g726) & (g1034) & (g1035) & (!g1036)) + ((sk[120]) & (g677) & (!g726) & (g1034) & (g1035) & (g1036)) + ((sk[120]) & (g677) & (g726) & (!g1034) & (g1035) & (!g1036)) + ((sk[120]) & (g677) & (g726) & (!g1034) & (g1035) & (g1036)) + ((sk[120]) & (g677) & (g726) & (g1034) & (g1035) & (!g1036)) + ((sk[120]) & (g677) & (g726) & (g1034) & (g1035) & (g1036)));
	assign g1847 = (((!g1038) & (!g1039) & (!g1040) & (g1041) & (g677) & (g726)) + ((!g1038) & (!g1039) & (g1040) & (!g1041) & (!g677) & (g726)) + ((!g1038) & (!g1039) & (g1040) & (g1041) & (!g677) & (g726)) + ((!g1038) & (!g1039) & (g1040) & (g1041) & (g677) & (g726)) + ((!g1038) & (g1039) & (!g1040) & (!g1041) & (g677) & (!g726)) + ((!g1038) & (g1039) & (!g1040) & (g1041) & (g677) & (!g726)) + ((!g1038) & (g1039) & (!g1040) & (g1041) & (g677) & (g726)) + ((!g1038) & (g1039) & (g1040) & (!g1041) & (!g677) & (g726)) + ((!g1038) & (g1039) & (g1040) & (!g1041) & (g677) & (!g726)) + ((!g1038) & (g1039) & (g1040) & (g1041) & (!g677) & (g726)) + ((!g1038) & (g1039) & (g1040) & (g1041) & (g677) & (!g726)) + ((!g1038) & (g1039) & (g1040) & (g1041) & (g677) & (g726)) + ((g1038) & (!g1039) & (!g1040) & (!g1041) & (!g677) & (!g726)) + ((g1038) & (!g1039) & (!g1040) & (g1041) & (!g677) & (!g726)) + ((g1038) & (!g1039) & (!g1040) & (g1041) & (g677) & (g726)) + ((g1038) & (!g1039) & (g1040) & (!g1041) & (!g677) & (!g726)) + ((g1038) & (!g1039) & (g1040) & (!g1041) & (!g677) & (g726)) + ((g1038) & (!g1039) & (g1040) & (g1041) & (!g677) & (!g726)) + ((g1038) & (!g1039) & (g1040) & (g1041) & (!g677) & (g726)) + ((g1038) & (!g1039) & (g1040) & (g1041) & (g677) & (g726)) + ((g1038) & (g1039) & (!g1040) & (!g1041) & (!g677) & (!g726)) + ((g1038) & (g1039) & (!g1040) & (!g1041) & (g677) & (!g726)) + ((g1038) & (g1039) & (!g1040) & (g1041) & (!g677) & (!g726)) + ((g1038) & (g1039) & (!g1040) & (g1041) & (g677) & (!g726)) + ((g1038) & (g1039) & (!g1040) & (g1041) & (g677) & (g726)) + ((g1038) & (g1039) & (g1040) & (!g1041) & (!g677) & (!g726)) + ((g1038) & (g1039) & (g1040) & (!g1041) & (!g677) & (g726)) + ((g1038) & (g1039) & (g1040) & (!g1041) & (g677) & (!g726)) + ((g1038) & (g1039) & (g1040) & (g1041) & (!g677) & (!g726)) + ((g1038) & (g1039) & (g1040) & (g1041) & (!g677) & (g726)) + ((g1038) & (g1039) & (g1040) & (g1041) & (g677) & (!g726)) + ((g1038) & (g1039) & (g1040) & (g1041) & (g677) & (g726)));
	assign g1848 = (((!g1043) & (!g1044) & (!g1045) & (g1046) & (g677) & (g726)) + ((!g1043) & (!g1044) & (g1045) & (!g1046) & (!g677) & (g726)) + ((!g1043) & (!g1044) & (g1045) & (g1046) & (!g677) & (g726)) + ((!g1043) & (!g1044) & (g1045) & (g1046) & (g677) & (g726)) + ((!g1043) & (g1044) & (!g1045) & (!g1046) & (g677) & (!g726)) + ((!g1043) & (g1044) & (!g1045) & (g1046) & (g677) & (!g726)) + ((!g1043) & (g1044) & (!g1045) & (g1046) & (g677) & (g726)) + ((!g1043) & (g1044) & (g1045) & (!g1046) & (!g677) & (g726)) + ((!g1043) & (g1044) & (g1045) & (!g1046) & (g677) & (!g726)) + ((!g1043) & (g1044) & (g1045) & (g1046) & (!g677) & (g726)) + ((!g1043) & (g1044) & (g1045) & (g1046) & (g677) & (!g726)) + ((!g1043) & (g1044) & (g1045) & (g1046) & (g677) & (g726)) + ((g1043) & (!g1044) & (!g1045) & (!g1046) & (!g677) & (!g726)) + ((g1043) & (!g1044) & (!g1045) & (g1046) & (!g677) & (!g726)) + ((g1043) & (!g1044) & (!g1045) & (g1046) & (g677) & (g726)) + ((g1043) & (!g1044) & (g1045) & (!g1046) & (!g677) & (!g726)) + ((g1043) & (!g1044) & (g1045) & (!g1046) & (!g677) & (g726)) + ((g1043) & (!g1044) & (g1045) & (g1046) & (!g677) & (!g726)) + ((g1043) & (!g1044) & (g1045) & (g1046) & (!g677) & (g726)) + ((g1043) & (!g1044) & (g1045) & (g1046) & (g677) & (g726)) + ((g1043) & (g1044) & (!g1045) & (!g1046) & (!g677) & (!g726)) + ((g1043) & (g1044) & (!g1045) & (!g1046) & (g677) & (!g726)) + ((g1043) & (g1044) & (!g1045) & (g1046) & (!g677) & (!g726)) + ((g1043) & (g1044) & (!g1045) & (g1046) & (g677) & (!g726)) + ((g1043) & (g1044) & (!g1045) & (g1046) & (g677) & (g726)) + ((g1043) & (g1044) & (g1045) & (!g1046) & (!g677) & (!g726)) + ((g1043) & (g1044) & (g1045) & (!g1046) & (!g677) & (g726)) + ((g1043) & (g1044) & (g1045) & (!g1046) & (g677) & (!g726)) + ((g1043) & (g1044) & (g1045) & (g1046) & (!g677) & (!g726)) + ((g1043) & (g1044) & (g1045) & (g1046) & (!g677) & (g726)) + ((g1043) & (g1044) & (g1045) & (g1046) & (g677) & (!g726)) + ((g1043) & (g1044) & (g1045) & (g1046) & (g677) & (g726)));
	assign g1849 = (((!g820) & (!g773) & (!g1845) & (g1846) & (!g1847) & (!g1848)) + ((!g820) & (!g773) & (!g1845) & (g1846) & (!g1847) & (g1848)) + ((!g820) & (!g773) & (!g1845) & (g1846) & (g1847) & (!g1848)) + ((!g820) & (!g773) & (!g1845) & (g1846) & (g1847) & (g1848)) + ((!g820) & (!g773) & (g1845) & (g1846) & (!g1847) & (!g1848)) + ((!g820) & (!g773) & (g1845) & (g1846) & (!g1847) & (g1848)) + ((!g820) & (!g773) & (g1845) & (g1846) & (g1847) & (!g1848)) + ((!g820) & (!g773) & (g1845) & (g1846) & (g1847) & (g1848)) + ((!g820) & (g773) & (!g1845) & (!g1846) & (!g1847) & (g1848)) + ((!g820) & (g773) & (!g1845) & (!g1846) & (g1847) & (g1848)) + ((!g820) & (g773) & (!g1845) & (g1846) & (!g1847) & (g1848)) + ((!g820) & (g773) & (!g1845) & (g1846) & (g1847) & (g1848)) + ((!g820) & (g773) & (g1845) & (!g1846) & (!g1847) & (g1848)) + ((!g820) & (g773) & (g1845) & (!g1846) & (g1847) & (g1848)) + ((!g820) & (g773) & (g1845) & (g1846) & (!g1847) & (g1848)) + ((!g820) & (g773) & (g1845) & (g1846) & (g1847) & (g1848)) + ((g820) & (!g773) & (g1845) & (!g1846) & (!g1847) & (!g1848)) + ((g820) & (!g773) & (g1845) & (!g1846) & (!g1847) & (g1848)) + ((g820) & (!g773) & (g1845) & (!g1846) & (g1847) & (!g1848)) + ((g820) & (!g773) & (g1845) & (!g1846) & (g1847) & (g1848)) + ((g820) & (!g773) & (g1845) & (g1846) & (!g1847) & (!g1848)) + ((g820) & (!g773) & (g1845) & (g1846) & (!g1847) & (g1848)) + ((g820) & (!g773) & (g1845) & (g1846) & (g1847) & (!g1848)) + ((g820) & (!g773) & (g1845) & (g1846) & (g1847) & (g1848)) + ((g820) & (g773) & (!g1845) & (!g1846) & (g1847) & (!g1848)) + ((g820) & (g773) & (!g1845) & (!g1846) & (g1847) & (g1848)) + ((g820) & (g773) & (!g1845) & (g1846) & (g1847) & (!g1848)) + ((g820) & (g773) & (!g1845) & (g1846) & (g1847) & (g1848)) + ((g820) & (g773) & (g1845) & (!g1846) & (g1847) & (!g1848)) + ((g820) & (g773) & (g1845) & (!g1846) & (g1847) & (g1848)) + ((g820) & (g773) & (g1845) & (g1846) & (g1847) & (!g1848)) + ((g820) & (g773) & (g1845) & (g1846) & (g1847) & (g1848)));
	assign g1850 = (((!g867) & (!sk[124]) & (!g1844) & (g1849)) + ((!g867) & (!sk[124]) & (g1844) & (!g1849)) + ((!g867) & (!sk[124]) & (g1844) & (g1849)) + ((!g867) & (sk[124]) & (!g1844) & (g1849)) + ((!g867) & (sk[124]) & (g1844) & (g1849)) + ((g867) & (!sk[124]) & (!g1844) & (g1849)) + ((g867) & (!sk[124]) & (g1844) & (!g1849)) + ((g867) & (!sk[124]) & (g1844) & (g1849)) + ((g867) & (sk[124]) & (g1844) & (!g1849)) + ((g867) & (sk[124]) & (g1844) & (g1849)));
	assign g1851 = (((!g1592) & (!g1593) & (!sk[125]) & (!g1605) & (g1644) & (!g54)) + ((!g1592) & (!g1593) & (!sk[125]) & (!g1605) & (g1644) & (g54)) + ((!g1592) & (!g1593) & (!sk[125]) & (g1605) & (!g1644) & (!g54)) + ((!g1592) & (!g1593) & (!sk[125]) & (g1605) & (!g1644) & (g54)) + ((!g1592) & (!g1593) & (!sk[125]) & (g1605) & (g1644) & (!g54)) + ((!g1592) & (!g1593) & (!sk[125]) & (g1605) & (g1644) & (g54)) + ((!g1592) & (!g1593) & (sk[125]) & (!g1605) & (g1644) & (!g54)) + ((!g1592) & (!g1593) & (sk[125]) & (!g1605) & (g1644) & (g54)) + ((!g1592) & (!g1593) & (sk[125]) & (g1605) & (g1644) & (!g54)) + ((!g1592) & (!g1593) & (sk[125]) & (g1605) & (g1644) & (g54)) + ((!g1592) & (g1593) & (!sk[125]) & (!g1605) & (!g1644) & (!g54)) + ((!g1592) & (g1593) & (!sk[125]) & (!g1605) & (!g1644) & (g54)) + ((!g1592) & (g1593) & (!sk[125]) & (!g1605) & (g1644) & (!g54)) + ((!g1592) & (g1593) & (!sk[125]) & (!g1605) & (g1644) & (g54)) + ((!g1592) & (g1593) & (!sk[125]) & (g1605) & (!g1644) & (!g54)) + ((!g1592) & (g1593) & (!sk[125]) & (g1605) & (!g1644) & (g54)) + ((!g1592) & (g1593) & (!sk[125]) & (g1605) & (g1644) & (!g54)) + ((!g1592) & (g1593) & (!sk[125]) & (g1605) & (g1644) & (g54)) + ((!g1592) & (g1593) & (sk[125]) & (!g1605) & (g1644) & (!g54)) + ((!g1592) & (g1593) & (sk[125]) & (!g1605) & (g1644) & (g54)) + ((!g1592) & (g1593) & (sk[125]) & (g1605) & (g1644) & (!g54)) + ((!g1592) & (g1593) & (sk[125]) & (g1605) & (g1644) & (g54)) + ((g1592) & (!g1593) & (!sk[125]) & (!g1605) & (g1644) & (!g54)) + ((g1592) & (!g1593) & (!sk[125]) & (!g1605) & (g1644) & (g54)) + ((g1592) & (!g1593) & (!sk[125]) & (g1605) & (!g1644) & (!g54)) + ((g1592) & (!g1593) & (!sk[125]) & (g1605) & (!g1644) & (g54)) + ((g1592) & (!g1593) & (!sk[125]) & (g1605) & (g1644) & (!g54)) + ((g1592) & (!g1593) & (!sk[125]) & (g1605) & (g1644) & (g54)) + ((g1592) & (!g1593) & (sk[125]) & (!g1605) & (g1644) & (!g54)) + ((g1592) & (!g1593) & (sk[125]) & (!g1605) & (g1644) & (g54)) + ((g1592) & (g1593) & (!sk[125]) & (!g1605) & (!g1644) & (!g54)) + ((g1592) & (g1593) & (!sk[125]) & (!g1605) & (!g1644) & (g54)) + ((g1592) & (g1593) & (!sk[125]) & (!g1605) & (g1644) & (!g54)) + ((g1592) & (g1593) & (!sk[125]) & (!g1605) & (g1644) & (g54)) + ((g1592) & (g1593) & (!sk[125]) & (g1605) & (!g1644) & (!g54)) + ((g1592) & (g1593) & (!sk[125]) & (g1605) & (!g1644) & (g54)) + ((g1592) & (g1593) & (!sk[125]) & (g1605) & (g1644) & (!g54)) + ((g1592) & (g1593) & (!sk[125]) & (g1605) & (g1644) & (g54)) + ((g1592) & (g1593) & (sk[125]) & (!g1605) & (!g1644) & (g54)) + ((g1592) & (g1593) & (sk[125]) & (!g1605) & (g1644) & (g54)) + ((g1592) & (g1593) & (sk[125]) & (g1605) & (!g1644) & (g54)) + ((g1592) & (g1593) & (sk[125]) & (g1605) & (g1644) & (g54)));
	assign g1852 = (((!g132) & (!sk[126]) & (!g1812) & (!g1850) & (g1851)) + ((!g132) & (!sk[126]) & (!g1812) & (g1850) & (!g1851)) + ((!g132) & (!sk[126]) & (!g1812) & (g1850) & (g1851)) + ((!g132) & (!sk[126]) & (g1812) & (!g1850) & (!g1851)) + ((!g132) & (!sk[126]) & (g1812) & (!g1850) & (g1851)) + ((!g132) & (!sk[126]) & (g1812) & (g1850) & (!g1851)) + ((!g132) & (!sk[126]) & (g1812) & (g1850) & (g1851)) + ((!g132) & (sk[126]) & (g1812) & (!g1850) & (g1851)) + ((!g132) & (sk[126]) & (g1812) & (g1850) & (g1851)) + ((g132) & (!sk[126]) & (!g1812) & (!g1850) & (g1851)) + ((g132) & (!sk[126]) & (!g1812) & (g1850) & (!g1851)) + ((g132) & (!sk[126]) & (!g1812) & (g1850) & (g1851)) + ((g132) & (!sk[126]) & (g1812) & (!g1850) & (!g1851)) + ((g132) & (!sk[126]) & (g1812) & (!g1850) & (g1851)) + ((g132) & (!sk[126]) & (g1812) & (g1850) & (!g1851)) + ((g132) & (!sk[126]) & (g1812) & (g1850) & (g1851)) + ((g132) & (sk[126]) & (g1812) & (g1850) & (!g1851)) + ((g132) & (sk[126]) & (g1812) & (g1850) & (g1851)));
	assign g1853 = (((!g1053) & (!g1054) & (!g1055) & (g1056) & (g820) & (g773)) + ((!g1053) & (!g1054) & (g1055) & (!g1056) & (!g820) & (g773)) + ((!g1053) & (!g1054) & (g1055) & (g1056) & (!g820) & (g773)) + ((!g1053) & (!g1054) & (g1055) & (g1056) & (g820) & (g773)) + ((!g1053) & (g1054) & (!g1055) & (!g1056) & (g820) & (!g773)) + ((!g1053) & (g1054) & (!g1055) & (g1056) & (g820) & (!g773)) + ((!g1053) & (g1054) & (!g1055) & (g1056) & (g820) & (g773)) + ((!g1053) & (g1054) & (g1055) & (!g1056) & (!g820) & (g773)) + ((!g1053) & (g1054) & (g1055) & (!g1056) & (g820) & (!g773)) + ((!g1053) & (g1054) & (g1055) & (g1056) & (!g820) & (g773)) + ((!g1053) & (g1054) & (g1055) & (g1056) & (g820) & (!g773)) + ((!g1053) & (g1054) & (g1055) & (g1056) & (g820) & (g773)) + ((g1053) & (!g1054) & (!g1055) & (!g1056) & (!g820) & (!g773)) + ((g1053) & (!g1054) & (!g1055) & (g1056) & (!g820) & (!g773)) + ((g1053) & (!g1054) & (!g1055) & (g1056) & (g820) & (g773)) + ((g1053) & (!g1054) & (g1055) & (!g1056) & (!g820) & (!g773)) + ((g1053) & (!g1054) & (g1055) & (!g1056) & (!g820) & (g773)) + ((g1053) & (!g1054) & (g1055) & (g1056) & (!g820) & (!g773)) + ((g1053) & (!g1054) & (g1055) & (g1056) & (!g820) & (g773)) + ((g1053) & (!g1054) & (g1055) & (g1056) & (g820) & (g773)) + ((g1053) & (g1054) & (!g1055) & (!g1056) & (!g820) & (!g773)) + ((g1053) & (g1054) & (!g1055) & (!g1056) & (g820) & (!g773)) + ((g1053) & (g1054) & (!g1055) & (g1056) & (!g820) & (!g773)) + ((g1053) & (g1054) & (!g1055) & (g1056) & (g820) & (!g773)) + ((g1053) & (g1054) & (!g1055) & (g1056) & (g820) & (g773)) + ((g1053) & (g1054) & (g1055) & (!g1056) & (!g820) & (!g773)) + ((g1053) & (g1054) & (g1055) & (!g1056) & (!g820) & (g773)) + ((g1053) & (g1054) & (g1055) & (!g1056) & (g820) & (!g773)) + ((g1053) & (g1054) & (g1055) & (g1056) & (!g820) & (!g773)) + ((g1053) & (g1054) & (g1055) & (g1056) & (!g820) & (g773)) + ((g1053) & (g1054) & (g1055) & (g1056) & (g820) & (!g773)) + ((g1053) & (g1054) & (g1055) & (g1056) & (g820) & (g773)));
	assign g1854 = (((!g1058) & (!g1059) & (!g1060) & (g1061) & (g820) & (g773)) + ((!g1058) & (!g1059) & (g1060) & (!g1061) & (!g820) & (g773)) + ((!g1058) & (!g1059) & (g1060) & (g1061) & (!g820) & (g773)) + ((!g1058) & (!g1059) & (g1060) & (g1061) & (g820) & (g773)) + ((!g1058) & (g1059) & (!g1060) & (!g1061) & (g820) & (!g773)) + ((!g1058) & (g1059) & (!g1060) & (g1061) & (g820) & (!g773)) + ((!g1058) & (g1059) & (!g1060) & (g1061) & (g820) & (g773)) + ((!g1058) & (g1059) & (g1060) & (!g1061) & (!g820) & (g773)) + ((!g1058) & (g1059) & (g1060) & (!g1061) & (g820) & (!g773)) + ((!g1058) & (g1059) & (g1060) & (g1061) & (!g820) & (g773)) + ((!g1058) & (g1059) & (g1060) & (g1061) & (g820) & (!g773)) + ((!g1058) & (g1059) & (g1060) & (g1061) & (g820) & (g773)) + ((g1058) & (!g1059) & (!g1060) & (!g1061) & (!g820) & (!g773)) + ((g1058) & (!g1059) & (!g1060) & (g1061) & (!g820) & (!g773)) + ((g1058) & (!g1059) & (!g1060) & (g1061) & (g820) & (g773)) + ((g1058) & (!g1059) & (g1060) & (!g1061) & (!g820) & (!g773)) + ((g1058) & (!g1059) & (g1060) & (!g1061) & (!g820) & (g773)) + ((g1058) & (!g1059) & (g1060) & (g1061) & (!g820) & (!g773)) + ((g1058) & (!g1059) & (g1060) & (g1061) & (!g820) & (g773)) + ((g1058) & (!g1059) & (g1060) & (g1061) & (g820) & (g773)) + ((g1058) & (g1059) & (!g1060) & (!g1061) & (!g820) & (!g773)) + ((g1058) & (g1059) & (!g1060) & (!g1061) & (g820) & (!g773)) + ((g1058) & (g1059) & (!g1060) & (g1061) & (!g820) & (!g773)) + ((g1058) & (g1059) & (!g1060) & (g1061) & (g820) & (!g773)) + ((g1058) & (g1059) & (!g1060) & (g1061) & (g820) & (g773)) + ((g1058) & (g1059) & (g1060) & (!g1061) & (!g820) & (!g773)) + ((g1058) & (g1059) & (g1060) & (!g1061) & (!g820) & (g773)) + ((g1058) & (g1059) & (g1060) & (!g1061) & (g820) & (!g773)) + ((g1058) & (g1059) & (g1060) & (g1061) & (!g820) & (!g773)) + ((g1058) & (g1059) & (g1060) & (g1061) & (!g820) & (g773)) + ((g1058) & (g1059) & (g1060) & (g1061) & (g820) & (!g773)) + ((g1058) & (g1059) & (g1060) & (g1061) & (g820) & (g773)));
	assign g1855 = (((!g1063) & (!g1064) & (!g1065) & (g1066) & (g820) & (g773)) + ((!g1063) & (!g1064) & (g1065) & (!g1066) & (!g820) & (g773)) + ((!g1063) & (!g1064) & (g1065) & (g1066) & (!g820) & (g773)) + ((!g1063) & (!g1064) & (g1065) & (g1066) & (g820) & (g773)) + ((!g1063) & (g1064) & (!g1065) & (!g1066) & (g820) & (!g773)) + ((!g1063) & (g1064) & (!g1065) & (g1066) & (g820) & (!g773)) + ((!g1063) & (g1064) & (!g1065) & (g1066) & (g820) & (g773)) + ((!g1063) & (g1064) & (g1065) & (!g1066) & (!g820) & (g773)) + ((!g1063) & (g1064) & (g1065) & (!g1066) & (g820) & (!g773)) + ((!g1063) & (g1064) & (g1065) & (g1066) & (!g820) & (g773)) + ((!g1063) & (g1064) & (g1065) & (g1066) & (g820) & (!g773)) + ((!g1063) & (g1064) & (g1065) & (g1066) & (g820) & (g773)) + ((g1063) & (!g1064) & (!g1065) & (!g1066) & (!g820) & (!g773)) + ((g1063) & (!g1064) & (!g1065) & (g1066) & (!g820) & (!g773)) + ((g1063) & (!g1064) & (!g1065) & (g1066) & (g820) & (g773)) + ((g1063) & (!g1064) & (g1065) & (!g1066) & (!g820) & (!g773)) + ((g1063) & (!g1064) & (g1065) & (!g1066) & (!g820) & (g773)) + ((g1063) & (!g1064) & (g1065) & (g1066) & (!g820) & (!g773)) + ((g1063) & (!g1064) & (g1065) & (g1066) & (!g820) & (g773)) + ((g1063) & (!g1064) & (g1065) & (g1066) & (g820) & (g773)) + ((g1063) & (g1064) & (!g1065) & (!g1066) & (!g820) & (!g773)) + ((g1063) & (g1064) & (!g1065) & (!g1066) & (g820) & (!g773)) + ((g1063) & (g1064) & (!g1065) & (g1066) & (!g820) & (!g773)) + ((g1063) & (g1064) & (!g1065) & (g1066) & (g820) & (!g773)) + ((g1063) & (g1064) & (!g1065) & (g1066) & (g820) & (g773)) + ((g1063) & (g1064) & (g1065) & (!g1066) & (!g820) & (!g773)) + ((g1063) & (g1064) & (g1065) & (!g1066) & (!g820) & (g773)) + ((g1063) & (g1064) & (g1065) & (!g1066) & (g820) & (!g773)) + ((g1063) & (g1064) & (g1065) & (g1066) & (!g820) & (!g773)) + ((g1063) & (g1064) & (g1065) & (g1066) & (!g820) & (g773)) + ((g1063) & (g1064) & (g1065) & (g1066) & (g820) & (!g773)) + ((g1063) & (g1064) & (g1065) & (g1066) & (g820) & (g773)));
	assign g1856 = (((!g1068) & (!g1069) & (!g1070) & (g1071) & (g820) & (g773)) + ((!g1068) & (!g1069) & (g1070) & (!g1071) & (!g820) & (g773)) + ((!g1068) & (!g1069) & (g1070) & (g1071) & (!g820) & (g773)) + ((!g1068) & (!g1069) & (g1070) & (g1071) & (g820) & (g773)) + ((!g1068) & (g1069) & (!g1070) & (!g1071) & (g820) & (!g773)) + ((!g1068) & (g1069) & (!g1070) & (g1071) & (g820) & (!g773)) + ((!g1068) & (g1069) & (!g1070) & (g1071) & (g820) & (g773)) + ((!g1068) & (g1069) & (g1070) & (!g1071) & (!g820) & (g773)) + ((!g1068) & (g1069) & (g1070) & (!g1071) & (g820) & (!g773)) + ((!g1068) & (g1069) & (g1070) & (g1071) & (!g820) & (g773)) + ((!g1068) & (g1069) & (g1070) & (g1071) & (g820) & (!g773)) + ((!g1068) & (g1069) & (g1070) & (g1071) & (g820) & (g773)) + ((g1068) & (!g1069) & (!g1070) & (!g1071) & (!g820) & (!g773)) + ((g1068) & (!g1069) & (!g1070) & (g1071) & (!g820) & (!g773)) + ((g1068) & (!g1069) & (!g1070) & (g1071) & (g820) & (g773)) + ((g1068) & (!g1069) & (g1070) & (!g1071) & (!g820) & (!g773)) + ((g1068) & (!g1069) & (g1070) & (!g1071) & (!g820) & (g773)) + ((g1068) & (!g1069) & (g1070) & (g1071) & (!g820) & (!g773)) + ((g1068) & (!g1069) & (g1070) & (g1071) & (!g820) & (g773)) + ((g1068) & (!g1069) & (g1070) & (g1071) & (g820) & (g773)) + ((g1068) & (g1069) & (!g1070) & (!g1071) & (!g820) & (!g773)) + ((g1068) & (g1069) & (!g1070) & (!g1071) & (g820) & (!g773)) + ((g1068) & (g1069) & (!g1070) & (g1071) & (!g820) & (!g773)) + ((g1068) & (g1069) & (!g1070) & (g1071) & (g820) & (!g773)) + ((g1068) & (g1069) & (!g1070) & (g1071) & (g820) & (g773)) + ((g1068) & (g1069) & (g1070) & (!g1071) & (!g820) & (!g773)) + ((g1068) & (g1069) & (g1070) & (!g1071) & (!g820) & (g773)) + ((g1068) & (g1069) & (g1070) & (!g1071) & (g820) & (!g773)) + ((g1068) & (g1069) & (g1070) & (g1071) & (!g820) & (!g773)) + ((g1068) & (g1069) & (g1070) & (g1071) & (!g820) & (g773)) + ((g1068) & (g1069) & (g1070) & (g1071) & (g820) & (!g773)) + ((g1068) & (g1069) & (g1070) & (g1071) & (g820) & (g773)));
	assign g1857 = (((!g1853) & (!g1854) & (!g1855) & (g1856) & (g677) & (g726)) + ((!g1853) & (!g1854) & (g1855) & (!g1856) & (!g677) & (g726)) + ((!g1853) & (!g1854) & (g1855) & (g1856) & (!g677) & (g726)) + ((!g1853) & (!g1854) & (g1855) & (g1856) & (g677) & (g726)) + ((!g1853) & (g1854) & (!g1855) & (!g1856) & (g677) & (!g726)) + ((!g1853) & (g1854) & (!g1855) & (g1856) & (g677) & (!g726)) + ((!g1853) & (g1854) & (!g1855) & (g1856) & (g677) & (g726)) + ((!g1853) & (g1854) & (g1855) & (!g1856) & (!g677) & (g726)) + ((!g1853) & (g1854) & (g1855) & (!g1856) & (g677) & (!g726)) + ((!g1853) & (g1854) & (g1855) & (g1856) & (!g677) & (g726)) + ((!g1853) & (g1854) & (g1855) & (g1856) & (g677) & (!g726)) + ((!g1853) & (g1854) & (g1855) & (g1856) & (g677) & (g726)) + ((g1853) & (!g1854) & (!g1855) & (!g1856) & (!g677) & (!g726)) + ((g1853) & (!g1854) & (!g1855) & (g1856) & (!g677) & (!g726)) + ((g1853) & (!g1854) & (!g1855) & (g1856) & (g677) & (g726)) + ((g1853) & (!g1854) & (g1855) & (!g1856) & (!g677) & (!g726)) + ((g1853) & (!g1854) & (g1855) & (!g1856) & (!g677) & (g726)) + ((g1853) & (!g1854) & (g1855) & (g1856) & (!g677) & (!g726)) + ((g1853) & (!g1854) & (g1855) & (g1856) & (!g677) & (g726)) + ((g1853) & (!g1854) & (g1855) & (g1856) & (g677) & (g726)) + ((g1853) & (g1854) & (!g1855) & (!g1856) & (!g677) & (!g726)) + ((g1853) & (g1854) & (!g1855) & (!g1856) & (g677) & (!g726)) + ((g1853) & (g1854) & (!g1855) & (g1856) & (!g677) & (!g726)) + ((g1853) & (g1854) & (!g1855) & (g1856) & (g677) & (!g726)) + ((g1853) & (g1854) & (!g1855) & (g1856) & (g677) & (g726)) + ((g1853) & (g1854) & (g1855) & (!g1856) & (!g677) & (!g726)) + ((g1853) & (g1854) & (g1855) & (!g1856) & (!g677) & (g726)) + ((g1853) & (g1854) & (g1855) & (!g1856) & (g677) & (!g726)) + ((g1853) & (g1854) & (g1855) & (g1856) & (!g677) & (!g726)) + ((g1853) & (g1854) & (g1855) & (g1856) & (!g677) & (g726)) + ((g1853) & (g1854) & (g1855) & (g1856) & (g677) & (!g726)) + ((g1853) & (g1854) & (g1855) & (g1856) & (g677) & (g726)));
	assign g1858 = (((!g1074) & (!g1075) & (!g1076) & (g1077) & (g677) & (g726)) + ((!g1074) & (!g1075) & (g1076) & (!g1077) & (!g677) & (g726)) + ((!g1074) & (!g1075) & (g1076) & (g1077) & (!g677) & (g726)) + ((!g1074) & (!g1075) & (g1076) & (g1077) & (g677) & (g726)) + ((!g1074) & (g1075) & (!g1076) & (!g1077) & (g677) & (!g726)) + ((!g1074) & (g1075) & (!g1076) & (g1077) & (g677) & (!g726)) + ((!g1074) & (g1075) & (!g1076) & (g1077) & (g677) & (g726)) + ((!g1074) & (g1075) & (g1076) & (!g1077) & (!g677) & (g726)) + ((!g1074) & (g1075) & (g1076) & (!g1077) & (g677) & (!g726)) + ((!g1074) & (g1075) & (g1076) & (g1077) & (!g677) & (g726)) + ((!g1074) & (g1075) & (g1076) & (g1077) & (g677) & (!g726)) + ((!g1074) & (g1075) & (g1076) & (g1077) & (g677) & (g726)) + ((g1074) & (!g1075) & (!g1076) & (!g1077) & (!g677) & (!g726)) + ((g1074) & (!g1075) & (!g1076) & (g1077) & (!g677) & (!g726)) + ((g1074) & (!g1075) & (!g1076) & (g1077) & (g677) & (g726)) + ((g1074) & (!g1075) & (g1076) & (!g1077) & (!g677) & (!g726)) + ((g1074) & (!g1075) & (g1076) & (!g1077) & (!g677) & (g726)) + ((g1074) & (!g1075) & (g1076) & (g1077) & (!g677) & (!g726)) + ((g1074) & (!g1075) & (g1076) & (g1077) & (!g677) & (g726)) + ((g1074) & (!g1075) & (g1076) & (g1077) & (g677) & (g726)) + ((g1074) & (g1075) & (!g1076) & (!g1077) & (!g677) & (!g726)) + ((g1074) & (g1075) & (!g1076) & (!g1077) & (g677) & (!g726)) + ((g1074) & (g1075) & (!g1076) & (g1077) & (!g677) & (!g726)) + ((g1074) & (g1075) & (!g1076) & (g1077) & (g677) & (!g726)) + ((g1074) & (g1075) & (!g1076) & (g1077) & (g677) & (g726)) + ((g1074) & (g1075) & (g1076) & (!g1077) & (!g677) & (!g726)) + ((g1074) & (g1075) & (g1076) & (!g1077) & (!g677) & (g726)) + ((g1074) & (g1075) & (g1076) & (!g1077) & (g677) & (!g726)) + ((g1074) & (g1075) & (g1076) & (g1077) & (!g677) & (!g726)) + ((g1074) & (g1075) & (g1076) & (g1077) & (!g677) & (g726)) + ((g1074) & (g1075) & (g1076) & (g1077) & (g677) & (!g726)) + ((g1074) & (g1075) & (g1076) & (g1077) & (g677) & (g726)));
	assign g1859 = (((!g677) & (!sk[5]) & (!g726) & (!g1079) & (g1080) & (!g1081)) + ((!g677) & (!sk[5]) & (!g726) & (!g1079) & (g1080) & (g1081)) + ((!g677) & (!sk[5]) & (!g726) & (g1079) & (!g1080) & (!g1081)) + ((!g677) & (!sk[5]) & (!g726) & (g1079) & (!g1080) & (g1081)) + ((!g677) & (!sk[5]) & (!g726) & (g1079) & (g1080) & (!g1081)) + ((!g677) & (!sk[5]) & (!g726) & (g1079) & (g1080) & (g1081)) + ((!g677) & (!sk[5]) & (g726) & (!g1079) & (!g1080) & (!g1081)) + ((!g677) & (!sk[5]) & (g726) & (!g1079) & (!g1080) & (g1081)) + ((!g677) & (!sk[5]) & (g726) & (!g1079) & (g1080) & (!g1081)) + ((!g677) & (!sk[5]) & (g726) & (!g1079) & (g1080) & (g1081)) + ((!g677) & (!sk[5]) & (g726) & (g1079) & (!g1080) & (!g1081)) + ((!g677) & (!sk[5]) & (g726) & (g1079) & (!g1080) & (g1081)) + ((!g677) & (!sk[5]) & (g726) & (g1079) & (g1080) & (!g1081)) + ((!g677) & (!sk[5]) & (g726) & (g1079) & (g1080) & (g1081)) + ((!g677) & (sk[5]) & (g726) & (!g1079) & (!g1080) & (g1081)) + ((!g677) & (sk[5]) & (g726) & (!g1079) & (g1080) & (g1081)) + ((!g677) & (sk[5]) & (g726) & (g1079) & (!g1080) & (g1081)) + ((!g677) & (sk[5]) & (g726) & (g1079) & (g1080) & (g1081)) + ((g677) & (!sk[5]) & (!g726) & (!g1079) & (g1080) & (!g1081)) + ((g677) & (!sk[5]) & (!g726) & (!g1079) & (g1080) & (g1081)) + ((g677) & (!sk[5]) & (!g726) & (g1079) & (!g1080) & (!g1081)) + ((g677) & (!sk[5]) & (!g726) & (g1079) & (!g1080) & (g1081)) + ((g677) & (!sk[5]) & (!g726) & (g1079) & (g1080) & (!g1081)) + ((g677) & (!sk[5]) & (!g726) & (g1079) & (g1080) & (g1081)) + ((g677) & (!sk[5]) & (g726) & (!g1079) & (!g1080) & (!g1081)) + ((g677) & (!sk[5]) & (g726) & (!g1079) & (!g1080) & (g1081)) + ((g677) & (!sk[5]) & (g726) & (!g1079) & (g1080) & (!g1081)) + ((g677) & (!sk[5]) & (g726) & (!g1079) & (g1080) & (g1081)) + ((g677) & (!sk[5]) & (g726) & (g1079) & (!g1080) & (!g1081)) + ((g677) & (!sk[5]) & (g726) & (g1079) & (!g1080) & (g1081)) + ((g677) & (!sk[5]) & (g726) & (g1079) & (g1080) & (!g1081)) + ((g677) & (!sk[5]) & (g726) & (g1079) & (g1080) & (g1081)) + ((g677) & (sk[5]) & (!g726) & (g1079) & (!g1080) & (!g1081)) + ((g677) & (sk[5]) & (!g726) & (g1079) & (!g1080) & (g1081)) + ((g677) & (sk[5]) & (!g726) & (g1079) & (g1080) & (!g1081)) + ((g677) & (sk[5]) & (!g726) & (g1079) & (g1080) & (g1081)) + ((g677) & (sk[5]) & (g726) & (!g1079) & (g1080) & (!g1081)) + ((g677) & (sk[5]) & (g726) & (!g1079) & (g1080) & (g1081)) + ((g677) & (sk[5]) & (g726) & (g1079) & (g1080) & (!g1081)) + ((g677) & (sk[5]) & (g726) & (g1079) & (g1080) & (g1081)));
	assign g1860 = (((!g1083) & (!g1084) & (!g1085) & (g1086) & (g677) & (g726)) + ((!g1083) & (!g1084) & (g1085) & (!g1086) & (!g677) & (g726)) + ((!g1083) & (!g1084) & (g1085) & (g1086) & (!g677) & (g726)) + ((!g1083) & (!g1084) & (g1085) & (g1086) & (g677) & (g726)) + ((!g1083) & (g1084) & (!g1085) & (!g1086) & (g677) & (!g726)) + ((!g1083) & (g1084) & (!g1085) & (g1086) & (g677) & (!g726)) + ((!g1083) & (g1084) & (!g1085) & (g1086) & (g677) & (g726)) + ((!g1083) & (g1084) & (g1085) & (!g1086) & (!g677) & (g726)) + ((!g1083) & (g1084) & (g1085) & (!g1086) & (g677) & (!g726)) + ((!g1083) & (g1084) & (g1085) & (g1086) & (!g677) & (g726)) + ((!g1083) & (g1084) & (g1085) & (g1086) & (g677) & (!g726)) + ((!g1083) & (g1084) & (g1085) & (g1086) & (g677) & (g726)) + ((g1083) & (!g1084) & (!g1085) & (!g1086) & (!g677) & (!g726)) + ((g1083) & (!g1084) & (!g1085) & (g1086) & (!g677) & (!g726)) + ((g1083) & (!g1084) & (!g1085) & (g1086) & (g677) & (g726)) + ((g1083) & (!g1084) & (g1085) & (!g1086) & (!g677) & (!g726)) + ((g1083) & (!g1084) & (g1085) & (!g1086) & (!g677) & (g726)) + ((g1083) & (!g1084) & (g1085) & (g1086) & (!g677) & (!g726)) + ((g1083) & (!g1084) & (g1085) & (g1086) & (!g677) & (g726)) + ((g1083) & (!g1084) & (g1085) & (g1086) & (g677) & (g726)) + ((g1083) & (g1084) & (!g1085) & (!g1086) & (!g677) & (!g726)) + ((g1083) & (g1084) & (!g1085) & (!g1086) & (g677) & (!g726)) + ((g1083) & (g1084) & (!g1085) & (g1086) & (!g677) & (!g726)) + ((g1083) & (g1084) & (!g1085) & (g1086) & (g677) & (!g726)) + ((g1083) & (g1084) & (!g1085) & (g1086) & (g677) & (g726)) + ((g1083) & (g1084) & (g1085) & (!g1086) & (!g677) & (!g726)) + ((g1083) & (g1084) & (g1085) & (!g1086) & (!g677) & (g726)) + ((g1083) & (g1084) & (g1085) & (!g1086) & (g677) & (!g726)) + ((g1083) & (g1084) & (g1085) & (g1086) & (!g677) & (!g726)) + ((g1083) & (g1084) & (g1085) & (g1086) & (!g677) & (g726)) + ((g1083) & (g1084) & (g1085) & (g1086) & (g677) & (!g726)) + ((g1083) & (g1084) & (g1085) & (g1086) & (g677) & (g726)));
	assign g1861 = (((!g1088) & (!g1089) & (!g1090) & (g1091) & (g677) & (g726)) + ((!g1088) & (!g1089) & (g1090) & (!g1091) & (!g677) & (g726)) + ((!g1088) & (!g1089) & (g1090) & (g1091) & (!g677) & (g726)) + ((!g1088) & (!g1089) & (g1090) & (g1091) & (g677) & (g726)) + ((!g1088) & (g1089) & (!g1090) & (!g1091) & (g677) & (!g726)) + ((!g1088) & (g1089) & (!g1090) & (g1091) & (g677) & (!g726)) + ((!g1088) & (g1089) & (!g1090) & (g1091) & (g677) & (g726)) + ((!g1088) & (g1089) & (g1090) & (!g1091) & (!g677) & (g726)) + ((!g1088) & (g1089) & (g1090) & (!g1091) & (g677) & (!g726)) + ((!g1088) & (g1089) & (g1090) & (g1091) & (!g677) & (g726)) + ((!g1088) & (g1089) & (g1090) & (g1091) & (g677) & (!g726)) + ((!g1088) & (g1089) & (g1090) & (g1091) & (g677) & (g726)) + ((g1088) & (!g1089) & (!g1090) & (!g1091) & (!g677) & (!g726)) + ((g1088) & (!g1089) & (!g1090) & (g1091) & (!g677) & (!g726)) + ((g1088) & (!g1089) & (!g1090) & (g1091) & (g677) & (g726)) + ((g1088) & (!g1089) & (g1090) & (!g1091) & (!g677) & (!g726)) + ((g1088) & (!g1089) & (g1090) & (!g1091) & (!g677) & (g726)) + ((g1088) & (!g1089) & (g1090) & (g1091) & (!g677) & (!g726)) + ((g1088) & (!g1089) & (g1090) & (g1091) & (!g677) & (g726)) + ((g1088) & (!g1089) & (g1090) & (g1091) & (g677) & (g726)) + ((g1088) & (g1089) & (!g1090) & (!g1091) & (!g677) & (!g726)) + ((g1088) & (g1089) & (!g1090) & (!g1091) & (g677) & (!g726)) + ((g1088) & (g1089) & (!g1090) & (g1091) & (!g677) & (!g726)) + ((g1088) & (g1089) & (!g1090) & (g1091) & (g677) & (!g726)) + ((g1088) & (g1089) & (!g1090) & (g1091) & (g677) & (g726)) + ((g1088) & (g1089) & (g1090) & (!g1091) & (!g677) & (!g726)) + ((g1088) & (g1089) & (g1090) & (!g1091) & (!g677) & (g726)) + ((g1088) & (g1089) & (g1090) & (!g1091) & (g677) & (!g726)) + ((g1088) & (g1089) & (g1090) & (g1091) & (!g677) & (!g726)) + ((g1088) & (g1089) & (g1090) & (g1091) & (!g677) & (g726)) + ((g1088) & (g1089) & (g1090) & (g1091) & (g677) & (!g726)) + ((g1088) & (g1089) & (g1090) & (g1091) & (g677) & (g726)));
	assign g1862 = (((!g820) & (!g773) & (!g1858) & (g1859) & (!g1860) & (!g1861)) + ((!g820) & (!g773) & (!g1858) & (g1859) & (!g1860) & (g1861)) + ((!g820) & (!g773) & (!g1858) & (g1859) & (g1860) & (!g1861)) + ((!g820) & (!g773) & (!g1858) & (g1859) & (g1860) & (g1861)) + ((!g820) & (!g773) & (g1858) & (g1859) & (!g1860) & (!g1861)) + ((!g820) & (!g773) & (g1858) & (g1859) & (!g1860) & (g1861)) + ((!g820) & (!g773) & (g1858) & (g1859) & (g1860) & (!g1861)) + ((!g820) & (!g773) & (g1858) & (g1859) & (g1860) & (g1861)) + ((!g820) & (g773) & (!g1858) & (!g1859) & (!g1860) & (g1861)) + ((!g820) & (g773) & (!g1858) & (!g1859) & (g1860) & (g1861)) + ((!g820) & (g773) & (!g1858) & (g1859) & (!g1860) & (g1861)) + ((!g820) & (g773) & (!g1858) & (g1859) & (g1860) & (g1861)) + ((!g820) & (g773) & (g1858) & (!g1859) & (!g1860) & (g1861)) + ((!g820) & (g773) & (g1858) & (!g1859) & (g1860) & (g1861)) + ((!g820) & (g773) & (g1858) & (g1859) & (!g1860) & (g1861)) + ((!g820) & (g773) & (g1858) & (g1859) & (g1860) & (g1861)) + ((g820) & (!g773) & (g1858) & (!g1859) & (!g1860) & (!g1861)) + ((g820) & (!g773) & (g1858) & (!g1859) & (!g1860) & (g1861)) + ((g820) & (!g773) & (g1858) & (!g1859) & (g1860) & (!g1861)) + ((g820) & (!g773) & (g1858) & (!g1859) & (g1860) & (g1861)) + ((g820) & (!g773) & (g1858) & (g1859) & (!g1860) & (!g1861)) + ((g820) & (!g773) & (g1858) & (g1859) & (!g1860) & (g1861)) + ((g820) & (!g773) & (g1858) & (g1859) & (g1860) & (!g1861)) + ((g820) & (!g773) & (g1858) & (g1859) & (g1860) & (g1861)) + ((g820) & (g773) & (!g1858) & (!g1859) & (g1860) & (!g1861)) + ((g820) & (g773) & (!g1858) & (!g1859) & (g1860) & (g1861)) + ((g820) & (g773) & (!g1858) & (g1859) & (g1860) & (!g1861)) + ((g820) & (g773) & (!g1858) & (g1859) & (g1860) & (g1861)) + ((g820) & (g773) & (g1858) & (!g1859) & (g1860) & (!g1861)) + ((g820) & (g773) & (g1858) & (!g1859) & (g1860) & (g1861)) + ((g820) & (g773) & (g1858) & (g1859) & (g1860) & (!g1861)) + ((g820) & (g773) & (g1858) & (g1859) & (g1860) & (g1861)));
	assign g1863 = (((!sk[9]) & (!g867) & (!g1857) & (g1862)) + ((!sk[9]) & (!g867) & (g1857) & (!g1862)) + ((!sk[9]) & (!g867) & (g1857) & (g1862)) + ((!sk[9]) & (g867) & (!g1857) & (g1862)) + ((!sk[9]) & (g867) & (g1857) & (!g1862)) + ((!sk[9]) & (g867) & (g1857) & (g1862)) + ((sk[9]) & (!g867) & (!g1857) & (g1862)) + ((sk[9]) & (!g867) & (g1857) & (g1862)) + ((sk[9]) & (g867) & (g1857) & (!g1862)) + ((sk[9]) & (g867) & (g1857) & (g1862)));
	assign g1864 = (((!g1592) & (!g1593) & (!g1605) & (g1656) & (!sk[10]) & (!g55)) + ((!g1592) & (!g1593) & (!g1605) & (g1656) & (!sk[10]) & (g55)) + ((!g1592) & (!g1593) & (!g1605) & (g1656) & (sk[10]) & (!g55)) + ((!g1592) & (!g1593) & (!g1605) & (g1656) & (sk[10]) & (g55)) + ((!g1592) & (!g1593) & (g1605) & (!g1656) & (!sk[10]) & (!g55)) + ((!g1592) & (!g1593) & (g1605) & (!g1656) & (!sk[10]) & (g55)) + ((!g1592) & (!g1593) & (g1605) & (g1656) & (!sk[10]) & (!g55)) + ((!g1592) & (!g1593) & (g1605) & (g1656) & (!sk[10]) & (g55)) + ((!g1592) & (!g1593) & (g1605) & (g1656) & (sk[10]) & (!g55)) + ((!g1592) & (!g1593) & (g1605) & (g1656) & (sk[10]) & (g55)) + ((!g1592) & (g1593) & (!g1605) & (!g1656) & (!sk[10]) & (!g55)) + ((!g1592) & (g1593) & (!g1605) & (!g1656) & (!sk[10]) & (g55)) + ((!g1592) & (g1593) & (!g1605) & (g1656) & (!sk[10]) & (!g55)) + ((!g1592) & (g1593) & (!g1605) & (g1656) & (!sk[10]) & (g55)) + ((!g1592) & (g1593) & (!g1605) & (g1656) & (sk[10]) & (!g55)) + ((!g1592) & (g1593) & (!g1605) & (g1656) & (sk[10]) & (g55)) + ((!g1592) & (g1593) & (g1605) & (!g1656) & (!sk[10]) & (!g55)) + ((!g1592) & (g1593) & (g1605) & (!g1656) & (!sk[10]) & (g55)) + ((!g1592) & (g1593) & (g1605) & (g1656) & (!sk[10]) & (!g55)) + ((!g1592) & (g1593) & (g1605) & (g1656) & (!sk[10]) & (g55)) + ((!g1592) & (g1593) & (g1605) & (g1656) & (sk[10]) & (!g55)) + ((!g1592) & (g1593) & (g1605) & (g1656) & (sk[10]) & (g55)) + ((g1592) & (!g1593) & (!g1605) & (g1656) & (!sk[10]) & (!g55)) + ((g1592) & (!g1593) & (!g1605) & (g1656) & (!sk[10]) & (g55)) + ((g1592) & (!g1593) & (!g1605) & (g1656) & (sk[10]) & (!g55)) + ((g1592) & (!g1593) & (!g1605) & (g1656) & (sk[10]) & (g55)) + ((g1592) & (!g1593) & (g1605) & (!g1656) & (!sk[10]) & (!g55)) + ((g1592) & (!g1593) & (g1605) & (!g1656) & (!sk[10]) & (g55)) + ((g1592) & (!g1593) & (g1605) & (g1656) & (!sk[10]) & (!g55)) + ((g1592) & (!g1593) & (g1605) & (g1656) & (!sk[10]) & (g55)) + ((g1592) & (g1593) & (!g1605) & (!g1656) & (!sk[10]) & (!g55)) + ((g1592) & (g1593) & (!g1605) & (!g1656) & (!sk[10]) & (g55)) + ((g1592) & (g1593) & (!g1605) & (!g1656) & (sk[10]) & (g55)) + ((g1592) & (g1593) & (!g1605) & (g1656) & (!sk[10]) & (!g55)) + ((g1592) & (g1593) & (!g1605) & (g1656) & (!sk[10]) & (g55)) + ((g1592) & (g1593) & (!g1605) & (g1656) & (sk[10]) & (g55)) + ((g1592) & (g1593) & (g1605) & (!g1656) & (!sk[10]) & (!g55)) + ((g1592) & (g1593) & (g1605) & (!g1656) & (!sk[10]) & (g55)) + ((g1592) & (g1593) & (g1605) & (!g1656) & (sk[10]) & (g55)) + ((g1592) & (g1593) & (g1605) & (g1656) & (!sk[10]) & (!g55)) + ((g1592) & (g1593) & (g1605) & (g1656) & (!sk[10]) & (g55)) + ((g1592) & (g1593) & (g1605) & (g1656) & (sk[10]) & (g55)));
	assign g1865 = (((!g132) & (!sk[11]) & (!g1812) & (!g1863) & (g1864)) + ((!g132) & (!sk[11]) & (!g1812) & (g1863) & (!g1864)) + ((!g132) & (!sk[11]) & (!g1812) & (g1863) & (g1864)) + ((!g132) & (!sk[11]) & (g1812) & (!g1863) & (!g1864)) + ((!g132) & (!sk[11]) & (g1812) & (!g1863) & (g1864)) + ((!g132) & (!sk[11]) & (g1812) & (g1863) & (!g1864)) + ((!g132) & (!sk[11]) & (g1812) & (g1863) & (g1864)) + ((!g132) & (sk[11]) & (g1812) & (!g1863) & (g1864)) + ((!g132) & (sk[11]) & (g1812) & (g1863) & (g1864)) + ((g132) & (!sk[11]) & (!g1812) & (!g1863) & (g1864)) + ((g132) & (!sk[11]) & (!g1812) & (g1863) & (!g1864)) + ((g132) & (!sk[11]) & (!g1812) & (g1863) & (g1864)) + ((g132) & (!sk[11]) & (g1812) & (!g1863) & (!g1864)) + ((g132) & (!sk[11]) & (g1812) & (!g1863) & (g1864)) + ((g132) & (!sk[11]) & (g1812) & (g1863) & (!g1864)) + ((g132) & (!sk[11]) & (g1812) & (g1863) & (g1864)) + ((g132) & (sk[11]) & (g1812) & (g1863) & (!g1864)) + ((g132) & (sk[11]) & (g1812) & (g1863) & (g1864)));
	assign g1866 = (((!g1098) & (!g1099) & (!g1100) & (g1101) & (g820) & (g773)) + ((!g1098) & (!g1099) & (g1100) & (!g1101) & (!g820) & (g773)) + ((!g1098) & (!g1099) & (g1100) & (g1101) & (!g820) & (g773)) + ((!g1098) & (!g1099) & (g1100) & (g1101) & (g820) & (g773)) + ((!g1098) & (g1099) & (!g1100) & (!g1101) & (g820) & (!g773)) + ((!g1098) & (g1099) & (!g1100) & (g1101) & (g820) & (!g773)) + ((!g1098) & (g1099) & (!g1100) & (g1101) & (g820) & (g773)) + ((!g1098) & (g1099) & (g1100) & (!g1101) & (!g820) & (g773)) + ((!g1098) & (g1099) & (g1100) & (!g1101) & (g820) & (!g773)) + ((!g1098) & (g1099) & (g1100) & (g1101) & (!g820) & (g773)) + ((!g1098) & (g1099) & (g1100) & (g1101) & (g820) & (!g773)) + ((!g1098) & (g1099) & (g1100) & (g1101) & (g820) & (g773)) + ((g1098) & (!g1099) & (!g1100) & (!g1101) & (!g820) & (!g773)) + ((g1098) & (!g1099) & (!g1100) & (g1101) & (!g820) & (!g773)) + ((g1098) & (!g1099) & (!g1100) & (g1101) & (g820) & (g773)) + ((g1098) & (!g1099) & (g1100) & (!g1101) & (!g820) & (!g773)) + ((g1098) & (!g1099) & (g1100) & (!g1101) & (!g820) & (g773)) + ((g1098) & (!g1099) & (g1100) & (g1101) & (!g820) & (!g773)) + ((g1098) & (!g1099) & (g1100) & (g1101) & (!g820) & (g773)) + ((g1098) & (!g1099) & (g1100) & (g1101) & (g820) & (g773)) + ((g1098) & (g1099) & (!g1100) & (!g1101) & (!g820) & (!g773)) + ((g1098) & (g1099) & (!g1100) & (!g1101) & (g820) & (!g773)) + ((g1098) & (g1099) & (!g1100) & (g1101) & (!g820) & (!g773)) + ((g1098) & (g1099) & (!g1100) & (g1101) & (g820) & (!g773)) + ((g1098) & (g1099) & (!g1100) & (g1101) & (g820) & (g773)) + ((g1098) & (g1099) & (g1100) & (!g1101) & (!g820) & (!g773)) + ((g1098) & (g1099) & (g1100) & (!g1101) & (!g820) & (g773)) + ((g1098) & (g1099) & (g1100) & (!g1101) & (g820) & (!g773)) + ((g1098) & (g1099) & (g1100) & (g1101) & (!g820) & (!g773)) + ((g1098) & (g1099) & (g1100) & (g1101) & (!g820) & (g773)) + ((g1098) & (g1099) & (g1100) & (g1101) & (g820) & (!g773)) + ((g1098) & (g1099) & (g1100) & (g1101) & (g820) & (g773)));
	assign g1867 = (((!g1103) & (!g1104) & (!g1105) & (g1106) & (g820) & (g773)) + ((!g1103) & (!g1104) & (g1105) & (!g1106) & (!g820) & (g773)) + ((!g1103) & (!g1104) & (g1105) & (g1106) & (!g820) & (g773)) + ((!g1103) & (!g1104) & (g1105) & (g1106) & (g820) & (g773)) + ((!g1103) & (g1104) & (!g1105) & (!g1106) & (g820) & (!g773)) + ((!g1103) & (g1104) & (!g1105) & (g1106) & (g820) & (!g773)) + ((!g1103) & (g1104) & (!g1105) & (g1106) & (g820) & (g773)) + ((!g1103) & (g1104) & (g1105) & (!g1106) & (!g820) & (g773)) + ((!g1103) & (g1104) & (g1105) & (!g1106) & (g820) & (!g773)) + ((!g1103) & (g1104) & (g1105) & (g1106) & (!g820) & (g773)) + ((!g1103) & (g1104) & (g1105) & (g1106) & (g820) & (!g773)) + ((!g1103) & (g1104) & (g1105) & (g1106) & (g820) & (g773)) + ((g1103) & (!g1104) & (!g1105) & (!g1106) & (!g820) & (!g773)) + ((g1103) & (!g1104) & (!g1105) & (g1106) & (!g820) & (!g773)) + ((g1103) & (!g1104) & (!g1105) & (g1106) & (g820) & (g773)) + ((g1103) & (!g1104) & (g1105) & (!g1106) & (!g820) & (!g773)) + ((g1103) & (!g1104) & (g1105) & (!g1106) & (!g820) & (g773)) + ((g1103) & (!g1104) & (g1105) & (g1106) & (!g820) & (!g773)) + ((g1103) & (!g1104) & (g1105) & (g1106) & (!g820) & (g773)) + ((g1103) & (!g1104) & (g1105) & (g1106) & (g820) & (g773)) + ((g1103) & (g1104) & (!g1105) & (!g1106) & (!g820) & (!g773)) + ((g1103) & (g1104) & (!g1105) & (!g1106) & (g820) & (!g773)) + ((g1103) & (g1104) & (!g1105) & (g1106) & (!g820) & (!g773)) + ((g1103) & (g1104) & (!g1105) & (g1106) & (g820) & (!g773)) + ((g1103) & (g1104) & (!g1105) & (g1106) & (g820) & (g773)) + ((g1103) & (g1104) & (g1105) & (!g1106) & (!g820) & (!g773)) + ((g1103) & (g1104) & (g1105) & (!g1106) & (!g820) & (g773)) + ((g1103) & (g1104) & (g1105) & (!g1106) & (g820) & (!g773)) + ((g1103) & (g1104) & (g1105) & (g1106) & (!g820) & (!g773)) + ((g1103) & (g1104) & (g1105) & (g1106) & (!g820) & (g773)) + ((g1103) & (g1104) & (g1105) & (g1106) & (g820) & (!g773)) + ((g1103) & (g1104) & (g1105) & (g1106) & (g820) & (g773)));
	assign g1868 = (((!g1108) & (!g1109) & (!g1110) & (g1111) & (g820) & (g773)) + ((!g1108) & (!g1109) & (g1110) & (!g1111) & (!g820) & (g773)) + ((!g1108) & (!g1109) & (g1110) & (g1111) & (!g820) & (g773)) + ((!g1108) & (!g1109) & (g1110) & (g1111) & (g820) & (g773)) + ((!g1108) & (g1109) & (!g1110) & (!g1111) & (g820) & (!g773)) + ((!g1108) & (g1109) & (!g1110) & (g1111) & (g820) & (!g773)) + ((!g1108) & (g1109) & (!g1110) & (g1111) & (g820) & (g773)) + ((!g1108) & (g1109) & (g1110) & (!g1111) & (!g820) & (g773)) + ((!g1108) & (g1109) & (g1110) & (!g1111) & (g820) & (!g773)) + ((!g1108) & (g1109) & (g1110) & (g1111) & (!g820) & (g773)) + ((!g1108) & (g1109) & (g1110) & (g1111) & (g820) & (!g773)) + ((!g1108) & (g1109) & (g1110) & (g1111) & (g820) & (g773)) + ((g1108) & (!g1109) & (!g1110) & (!g1111) & (!g820) & (!g773)) + ((g1108) & (!g1109) & (!g1110) & (g1111) & (!g820) & (!g773)) + ((g1108) & (!g1109) & (!g1110) & (g1111) & (g820) & (g773)) + ((g1108) & (!g1109) & (g1110) & (!g1111) & (!g820) & (!g773)) + ((g1108) & (!g1109) & (g1110) & (!g1111) & (!g820) & (g773)) + ((g1108) & (!g1109) & (g1110) & (g1111) & (!g820) & (!g773)) + ((g1108) & (!g1109) & (g1110) & (g1111) & (!g820) & (g773)) + ((g1108) & (!g1109) & (g1110) & (g1111) & (g820) & (g773)) + ((g1108) & (g1109) & (!g1110) & (!g1111) & (!g820) & (!g773)) + ((g1108) & (g1109) & (!g1110) & (!g1111) & (g820) & (!g773)) + ((g1108) & (g1109) & (!g1110) & (g1111) & (!g820) & (!g773)) + ((g1108) & (g1109) & (!g1110) & (g1111) & (g820) & (!g773)) + ((g1108) & (g1109) & (!g1110) & (g1111) & (g820) & (g773)) + ((g1108) & (g1109) & (g1110) & (!g1111) & (!g820) & (!g773)) + ((g1108) & (g1109) & (g1110) & (!g1111) & (!g820) & (g773)) + ((g1108) & (g1109) & (g1110) & (!g1111) & (g820) & (!g773)) + ((g1108) & (g1109) & (g1110) & (g1111) & (!g820) & (!g773)) + ((g1108) & (g1109) & (g1110) & (g1111) & (!g820) & (g773)) + ((g1108) & (g1109) & (g1110) & (g1111) & (g820) & (!g773)) + ((g1108) & (g1109) & (g1110) & (g1111) & (g820) & (g773)));
	assign g1869 = (((!g1113) & (!g1114) & (!g1115) & (g1116) & (g820) & (g773)) + ((!g1113) & (!g1114) & (g1115) & (!g1116) & (!g820) & (g773)) + ((!g1113) & (!g1114) & (g1115) & (g1116) & (!g820) & (g773)) + ((!g1113) & (!g1114) & (g1115) & (g1116) & (g820) & (g773)) + ((!g1113) & (g1114) & (!g1115) & (!g1116) & (g820) & (!g773)) + ((!g1113) & (g1114) & (!g1115) & (g1116) & (g820) & (!g773)) + ((!g1113) & (g1114) & (!g1115) & (g1116) & (g820) & (g773)) + ((!g1113) & (g1114) & (g1115) & (!g1116) & (!g820) & (g773)) + ((!g1113) & (g1114) & (g1115) & (!g1116) & (g820) & (!g773)) + ((!g1113) & (g1114) & (g1115) & (g1116) & (!g820) & (g773)) + ((!g1113) & (g1114) & (g1115) & (g1116) & (g820) & (!g773)) + ((!g1113) & (g1114) & (g1115) & (g1116) & (g820) & (g773)) + ((g1113) & (!g1114) & (!g1115) & (!g1116) & (!g820) & (!g773)) + ((g1113) & (!g1114) & (!g1115) & (g1116) & (!g820) & (!g773)) + ((g1113) & (!g1114) & (!g1115) & (g1116) & (g820) & (g773)) + ((g1113) & (!g1114) & (g1115) & (!g1116) & (!g820) & (!g773)) + ((g1113) & (!g1114) & (g1115) & (!g1116) & (!g820) & (g773)) + ((g1113) & (!g1114) & (g1115) & (g1116) & (!g820) & (!g773)) + ((g1113) & (!g1114) & (g1115) & (g1116) & (!g820) & (g773)) + ((g1113) & (!g1114) & (g1115) & (g1116) & (g820) & (g773)) + ((g1113) & (g1114) & (!g1115) & (!g1116) & (!g820) & (!g773)) + ((g1113) & (g1114) & (!g1115) & (!g1116) & (g820) & (!g773)) + ((g1113) & (g1114) & (!g1115) & (g1116) & (!g820) & (!g773)) + ((g1113) & (g1114) & (!g1115) & (g1116) & (g820) & (!g773)) + ((g1113) & (g1114) & (!g1115) & (g1116) & (g820) & (g773)) + ((g1113) & (g1114) & (g1115) & (!g1116) & (!g820) & (!g773)) + ((g1113) & (g1114) & (g1115) & (!g1116) & (!g820) & (g773)) + ((g1113) & (g1114) & (g1115) & (!g1116) & (g820) & (!g773)) + ((g1113) & (g1114) & (g1115) & (g1116) & (!g820) & (!g773)) + ((g1113) & (g1114) & (g1115) & (g1116) & (!g820) & (g773)) + ((g1113) & (g1114) & (g1115) & (g1116) & (g820) & (!g773)) + ((g1113) & (g1114) & (g1115) & (g1116) & (g820) & (g773)));
	assign g1870 = (((!g1866) & (!g1867) & (!g1868) & (g1869) & (g677) & (g726)) + ((!g1866) & (!g1867) & (g1868) & (!g1869) & (!g677) & (g726)) + ((!g1866) & (!g1867) & (g1868) & (g1869) & (!g677) & (g726)) + ((!g1866) & (!g1867) & (g1868) & (g1869) & (g677) & (g726)) + ((!g1866) & (g1867) & (!g1868) & (!g1869) & (g677) & (!g726)) + ((!g1866) & (g1867) & (!g1868) & (g1869) & (g677) & (!g726)) + ((!g1866) & (g1867) & (!g1868) & (g1869) & (g677) & (g726)) + ((!g1866) & (g1867) & (g1868) & (!g1869) & (!g677) & (g726)) + ((!g1866) & (g1867) & (g1868) & (!g1869) & (g677) & (!g726)) + ((!g1866) & (g1867) & (g1868) & (g1869) & (!g677) & (g726)) + ((!g1866) & (g1867) & (g1868) & (g1869) & (g677) & (!g726)) + ((!g1866) & (g1867) & (g1868) & (g1869) & (g677) & (g726)) + ((g1866) & (!g1867) & (!g1868) & (!g1869) & (!g677) & (!g726)) + ((g1866) & (!g1867) & (!g1868) & (g1869) & (!g677) & (!g726)) + ((g1866) & (!g1867) & (!g1868) & (g1869) & (g677) & (g726)) + ((g1866) & (!g1867) & (g1868) & (!g1869) & (!g677) & (!g726)) + ((g1866) & (!g1867) & (g1868) & (!g1869) & (!g677) & (g726)) + ((g1866) & (!g1867) & (g1868) & (g1869) & (!g677) & (!g726)) + ((g1866) & (!g1867) & (g1868) & (g1869) & (!g677) & (g726)) + ((g1866) & (!g1867) & (g1868) & (g1869) & (g677) & (g726)) + ((g1866) & (g1867) & (!g1868) & (!g1869) & (!g677) & (!g726)) + ((g1866) & (g1867) & (!g1868) & (!g1869) & (g677) & (!g726)) + ((g1866) & (g1867) & (!g1868) & (g1869) & (!g677) & (!g726)) + ((g1866) & (g1867) & (!g1868) & (g1869) & (g677) & (!g726)) + ((g1866) & (g1867) & (!g1868) & (g1869) & (g677) & (g726)) + ((g1866) & (g1867) & (g1868) & (!g1869) & (!g677) & (!g726)) + ((g1866) & (g1867) & (g1868) & (!g1869) & (!g677) & (g726)) + ((g1866) & (g1867) & (g1868) & (!g1869) & (g677) & (!g726)) + ((g1866) & (g1867) & (g1868) & (g1869) & (!g677) & (!g726)) + ((g1866) & (g1867) & (g1868) & (g1869) & (!g677) & (g726)) + ((g1866) & (g1867) & (g1868) & (g1869) & (g677) & (!g726)) + ((g1866) & (g1867) & (g1868) & (g1869) & (g677) & (g726)));
	assign g1871 = (((!g1119) & (!g1120) & (!g1121) & (g1122) & (g677) & (g726)) + ((!g1119) & (!g1120) & (g1121) & (!g1122) & (!g677) & (g726)) + ((!g1119) & (!g1120) & (g1121) & (g1122) & (!g677) & (g726)) + ((!g1119) & (!g1120) & (g1121) & (g1122) & (g677) & (g726)) + ((!g1119) & (g1120) & (!g1121) & (!g1122) & (g677) & (!g726)) + ((!g1119) & (g1120) & (!g1121) & (g1122) & (g677) & (!g726)) + ((!g1119) & (g1120) & (!g1121) & (g1122) & (g677) & (g726)) + ((!g1119) & (g1120) & (g1121) & (!g1122) & (!g677) & (g726)) + ((!g1119) & (g1120) & (g1121) & (!g1122) & (g677) & (!g726)) + ((!g1119) & (g1120) & (g1121) & (g1122) & (!g677) & (g726)) + ((!g1119) & (g1120) & (g1121) & (g1122) & (g677) & (!g726)) + ((!g1119) & (g1120) & (g1121) & (g1122) & (g677) & (g726)) + ((g1119) & (!g1120) & (!g1121) & (!g1122) & (!g677) & (!g726)) + ((g1119) & (!g1120) & (!g1121) & (g1122) & (!g677) & (!g726)) + ((g1119) & (!g1120) & (!g1121) & (g1122) & (g677) & (g726)) + ((g1119) & (!g1120) & (g1121) & (!g1122) & (!g677) & (!g726)) + ((g1119) & (!g1120) & (g1121) & (!g1122) & (!g677) & (g726)) + ((g1119) & (!g1120) & (g1121) & (g1122) & (!g677) & (!g726)) + ((g1119) & (!g1120) & (g1121) & (g1122) & (!g677) & (g726)) + ((g1119) & (!g1120) & (g1121) & (g1122) & (g677) & (g726)) + ((g1119) & (g1120) & (!g1121) & (!g1122) & (!g677) & (!g726)) + ((g1119) & (g1120) & (!g1121) & (!g1122) & (g677) & (!g726)) + ((g1119) & (g1120) & (!g1121) & (g1122) & (!g677) & (!g726)) + ((g1119) & (g1120) & (!g1121) & (g1122) & (g677) & (!g726)) + ((g1119) & (g1120) & (!g1121) & (g1122) & (g677) & (g726)) + ((g1119) & (g1120) & (g1121) & (!g1122) & (!g677) & (!g726)) + ((g1119) & (g1120) & (g1121) & (!g1122) & (!g677) & (g726)) + ((g1119) & (g1120) & (g1121) & (!g1122) & (g677) & (!g726)) + ((g1119) & (g1120) & (g1121) & (g1122) & (!g677) & (!g726)) + ((g1119) & (g1120) & (g1121) & (g1122) & (!g677) & (g726)) + ((g1119) & (g1120) & (g1121) & (g1122) & (g677) & (!g726)) + ((g1119) & (g1120) & (g1121) & (g1122) & (g677) & (g726)));
	assign g1872 = (((!g677) & (!g726) & (!sk[18]) & (!g1124) & (g1125) & (!g1126)) + ((!g677) & (!g726) & (!sk[18]) & (!g1124) & (g1125) & (g1126)) + ((!g677) & (!g726) & (!sk[18]) & (g1124) & (!g1125) & (!g1126)) + ((!g677) & (!g726) & (!sk[18]) & (g1124) & (!g1125) & (g1126)) + ((!g677) & (!g726) & (!sk[18]) & (g1124) & (g1125) & (!g1126)) + ((!g677) & (!g726) & (!sk[18]) & (g1124) & (g1125) & (g1126)) + ((!g677) & (g726) & (!sk[18]) & (!g1124) & (!g1125) & (!g1126)) + ((!g677) & (g726) & (!sk[18]) & (!g1124) & (!g1125) & (g1126)) + ((!g677) & (g726) & (!sk[18]) & (!g1124) & (g1125) & (!g1126)) + ((!g677) & (g726) & (!sk[18]) & (!g1124) & (g1125) & (g1126)) + ((!g677) & (g726) & (!sk[18]) & (g1124) & (!g1125) & (!g1126)) + ((!g677) & (g726) & (!sk[18]) & (g1124) & (!g1125) & (g1126)) + ((!g677) & (g726) & (!sk[18]) & (g1124) & (g1125) & (!g1126)) + ((!g677) & (g726) & (!sk[18]) & (g1124) & (g1125) & (g1126)) + ((!g677) & (g726) & (sk[18]) & (!g1124) & (!g1125) & (g1126)) + ((!g677) & (g726) & (sk[18]) & (!g1124) & (g1125) & (g1126)) + ((!g677) & (g726) & (sk[18]) & (g1124) & (!g1125) & (g1126)) + ((!g677) & (g726) & (sk[18]) & (g1124) & (g1125) & (g1126)) + ((g677) & (!g726) & (!sk[18]) & (!g1124) & (g1125) & (!g1126)) + ((g677) & (!g726) & (!sk[18]) & (!g1124) & (g1125) & (g1126)) + ((g677) & (!g726) & (!sk[18]) & (g1124) & (!g1125) & (!g1126)) + ((g677) & (!g726) & (!sk[18]) & (g1124) & (!g1125) & (g1126)) + ((g677) & (!g726) & (!sk[18]) & (g1124) & (g1125) & (!g1126)) + ((g677) & (!g726) & (!sk[18]) & (g1124) & (g1125) & (g1126)) + ((g677) & (!g726) & (sk[18]) & (g1124) & (!g1125) & (!g1126)) + ((g677) & (!g726) & (sk[18]) & (g1124) & (!g1125) & (g1126)) + ((g677) & (!g726) & (sk[18]) & (g1124) & (g1125) & (!g1126)) + ((g677) & (!g726) & (sk[18]) & (g1124) & (g1125) & (g1126)) + ((g677) & (g726) & (!sk[18]) & (!g1124) & (!g1125) & (!g1126)) + ((g677) & (g726) & (!sk[18]) & (!g1124) & (!g1125) & (g1126)) + ((g677) & (g726) & (!sk[18]) & (!g1124) & (g1125) & (!g1126)) + ((g677) & (g726) & (!sk[18]) & (!g1124) & (g1125) & (g1126)) + ((g677) & (g726) & (!sk[18]) & (g1124) & (!g1125) & (!g1126)) + ((g677) & (g726) & (!sk[18]) & (g1124) & (!g1125) & (g1126)) + ((g677) & (g726) & (!sk[18]) & (g1124) & (g1125) & (!g1126)) + ((g677) & (g726) & (!sk[18]) & (g1124) & (g1125) & (g1126)) + ((g677) & (g726) & (sk[18]) & (!g1124) & (g1125) & (!g1126)) + ((g677) & (g726) & (sk[18]) & (!g1124) & (g1125) & (g1126)) + ((g677) & (g726) & (sk[18]) & (g1124) & (g1125) & (!g1126)) + ((g677) & (g726) & (sk[18]) & (g1124) & (g1125) & (g1126)));
	assign g1873 = (((!g1128) & (!g1129) & (!g1130) & (g1131) & (g677) & (g726)) + ((!g1128) & (!g1129) & (g1130) & (!g1131) & (!g677) & (g726)) + ((!g1128) & (!g1129) & (g1130) & (g1131) & (!g677) & (g726)) + ((!g1128) & (!g1129) & (g1130) & (g1131) & (g677) & (g726)) + ((!g1128) & (g1129) & (!g1130) & (!g1131) & (g677) & (!g726)) + ((!g1128) & (g1129) & (!g1130) & (g1131) & (g677) & (!g726)) + ((!g1128) & (g1129) & (!g1130) & (g1131) & (g677) & (g726)) + ((!g1128) & (g1129) & (g1130) & (!g1131) & (!g677) & (g726)) + ((!g1128) & (g1129) & (g1130) & (!g1131) & (g677) & (!g726)) + ((!g1128) & (g1129) & (g1130) & (g1131) & (!g677) & (g726)) + ((!g1128) & (g1129) & (g1130) & (g1131) & (g677) & (!g726)) + ((!g1128) & (g1129) & (g1130) & (g1131) & (g677) & (g726)) + ((g1128) & (!g1129) & (!g1130) & (!g1131) & (!g677) & (!g726)) + ((g1128) & (!g1129) & (!g1130) & (g1131) & (!g677) & (!g726)) + ((g1128) & (!g1129) & (!g1130) & (g1131) & (g677) & (g726)) + ((g1128) & (!g1129) & (g1130) & (!g1131) & (!g677) & (!g726)) + ((g1128) & (!g1129) & (g1130) & (!g1131) & (!g677) & (g726)) + ((g1128) & (!g1129) & (g1130) & (g1131) & (!g677) & (!g726)) + ((g1128) & (!g1129) & (g1130) & (g1131) & (!g677) & (g726)) + ((g1128) & (!g1129) & (g1130) & (g1131) & (g677) & (g726)) + ((g1128) & (g1129) & (!g1130) & (!g1131) & (!g677) & (!g726)) + ((g1128) & (g1129) & (!g1130) & (!g1131) & (g677) & (!g726)) + ((g1128) & (g1129) & (!g1130) & (g1131) & (!g677) & (!g726)) + ((g1128) & (g1129) & (!g1130) & (g1131) & (g677) & (!g726)) + ((g1128) & (g1129) & (!g1130) & (g1131) & (g677) & (g726)) + ((g1128) & (g1129) & (g1130) & (!g1131) & (!g677) & (!g726)) + ((g1128) & (g1129) & (g1130) & (!g1131) & (!g677) & (g726)) + ((g1128) & (g1129) & (g1130) & (!g1131) & (g677) & (!g726)) + ((g1128) & (g1129) & (g1130) & (g1131) & (!g677) & (!g726)) + ((g1128) & (g1129) & (g1130) & (g1131) & (!g677) & (g726)) + ((g1128) & (g1129) & (g1130) & (g1131) & (g677) & (!g726)) + ((g1128) & (g1129) & (g1130) & (g1131) & (g677) & (g726)));
	assign g1874 = (((!g1133) & (!g1134) & (!g1135) & (g1136) & (g677) & (g726)) + ((!g1133) & (!g1134) & (g1135) & (!g1136) & (!g677) & (g726)) + ((!g1133) & (!g1134) & (g1135) & (g1136) & (!g677) & (g726)) + ((!g1133) & (!g1134) & (g1135) & (g1136) & (g677) & (g726)) + ((!g1133) & (g1134) & (!g1135) & (!g1136) & (g677) & (!g726)) + ((!g1133) & (g1134) & (!g1135) & (g1136) & (g677) & (!g726)) + ((!g1133) & (g1134) & (!g1135) & (g1136) & (g677) & (g726)) + ((!g1133) & (g1134) & (g1135) & (!g1136) & (!g677) & (g726)) + ((!g1133) & (g1134) & (g1135) & (!g1136) & (g677) & (!g726)) + ((!g1133) & (g1134) & (g1135) & (g1136) & (!g677) & (g726)) + ((!g1133) & (g1134) & (g1135) & (g1136) & (g677) & (!g726)) + ((!g1133) & (g1134) & (g1135) & (g1136) & (g677) & (g726)) + ((g1133) & (!g1134) & (!g1135) & (!g1136) & (!g677) & (!g726)) + ((g1133) & (!g1134) & (!g1135) & (g1136) & (!g677) & (!g726)) + ((g1133) & (!g1134) & (!g1135) & (g1136) & (g677) & (g726)) + ((g1133) & (!g1134) & (g1135) & (!g1136) & (!g677) & (!g726)) + ((g1133) & (!g1134) & (g1135) & (!g1136) & (!g677) & (g726)) + ((g1133) & (!g1134) & (g1135) & (g1136) & (!g677) & (!g726)) + ((g1133) & (!g1134) & (g1135) & (g1136) & (!g677) & (g726)) + ((g1133) & (!g1134) & (g1135) & (g1136) & (g677) & (g726)) + ((g1133) & (g1134) & (!g1135) & (!g1136) & (!g677) & (!g726)) + ((g1133) & (g1134) & (!g1135) & (!g1136) & (g677) & (!g726)) + ((g1133) & (g1134) & (!g1135) & (g1136) & (!g677) & (!g726)) + ((g1133) & (g1134) & (!g1135) & (g1136) & (g677) & (!g726)) + ((g1133) & (g1134) & (!g1135) & (g1136) & (g677) & (g726)) + ((g1133) & (g1134) & (g1135) & (!g1136) & (!g677) & (!g726)) + ((g1133) & (g1134) & (g1135) & (!g1136) & (!g677) & (g726)) + ((g1133) & (g1134) & (g1135) & (!g1136) & (g677) & (!g726)) + ((g1133) & (g1134) & (g1135) & (g1136) & (!g677) & (!g726)) + ((g1133) & (g1134) & (g1135) & (g1136) & (!g677) & (g726)) + ((g1133) & (g1134) & (g1135) & (g1136) & (g677) & (!g726)) + ((g1133) & (g1134) & (g1135) & (g1136) & (g677) & (g726)));
	assign g1875 = (((!g820) & (!g773) & (!g1871) & (g1872) & (!g1873) & (!g1874)) + ((!g820) & (!g773) & (!g1871) & (g1872) & (!g1873) & (g1874)) + ((!g820) & (!g773) & (!g1871) & (g1872) & (g1873) & (!g1874)) + ((!g820) & (!g773) & (!g1871) & (g1872) & (g1873) & (g1874)) + ((!g820) & (!g773) & (g1871) & (g1872) & (!g1873) & (!g1874)) + ((!g820) & (!g773) & (g1871) & (g1872) & (!g1873) & (g1874)) + ((!g820) & (!g773) & (g1871) & (g1872) & (g1873) & (!g1874)) + ((!g820) & (!g773) & (g1871) & (g1872) & (g1873) & (g1874)) + ((!g820) & (g773) & (!g1871) & (!g1872) & (!g1873) & (g1874)) + ((!g820) & (g773) & (!g1871) & (!g1872) & (g1873) & (g1874)) + ((!g820) & (g773) & (!g1871) & (g1872) & (!g1873) & (g1874)) + ((!g820) & (g773) & (!g1871) & (g1872) & (g1873) & (g1874)) + ((!g820) & (g773) & (g1871) & (!g1872) & (!g1873) & (g1874)) + ((!g820) & (g773) & (g1871) & (!g1872) & (g1873) & (g1874)) + ((!g820) & (g773) & (g1871) & (g1872) & (!g1873) & (g1874)) + ((!g820) & (g773) & (g1871) & (g1872) & (g1873) & (g1874)) + ((g820) & (!g773) & (g1871) & (!g1872) & (!g1873) & (!g1874)) + ((g820) & (!g773) & (g1871) & (!g1872) & (!g1873) & (g1874)) + ((g820) & (!g773) & (g1871) & (!g1872) & (g1873) & (!g1874)) + ((g820) & (!g773) & (g1871) & (!g1872) & (g1873) & (g1874)) + ((g820) & (!g773) & (g1871) & (g1872) & (!g1873) & (!g1874)) + ((g820) & (!g773) & (g1871) & (g1872) & (!g1873) & (g1874)) + ((g820) & (!g773) & (g1871) & (g1872) & (g1873) & (!g1874)) + ((g820) & (!g773) & (g1871) & (g1872) & (g1873) & (g1874)) + ((g820) & (g773) & (!g1871) & (!g1872) & (g1873) & (!g1874)) + ((g820) & (g773) & (!g1871) & (!g1872) & (g1873) & (g1874)) + ((g820) & (g773) & (!g1871) & (g1872) & (g1873) & (!g1874)) + ((g820) & (g773) & (!g1871) & (g1872) & (g1873) & (g1874)) + ((g820) & (g773) & (g1871) & (!g1872) & (g1873) & (!g1874)) + ((g820) & (g773) & (g1871) & (!g1872) & (g1873) & (g1874)) + ((g820) & (g773) & (g1871) & (g1872) & (g1873) & (!g1874)) + ((g820) & (g773) & (g1871) & (g1872) & (g1873) & (g1874)));
	assign g1876 = (((!sk[22]) & (!g867) & (!g1870) & (g1875)) + ((!sk[22]) & (!g867) & (g1870) & (!g1875)) + ((!sk[22]) & (!g867) & (g1870) & (g1875)) + ((!sk[22]) & (g867) & (!g1870) & (g1875)) + ((!sk[22]) & (g867) & (g1870) & (!g1875)) + ((!sk[22]) & (g867) & (g1870) & (g1875)) + ((sk[22]) & (!g867) & (!g1870) & (g1875)) + ((sk[22]) & (!g867) & (g1870) & (g1875)) + ((sk[22]) & (g867) & (g1870) & (!g1875)) + ((sk[22]) & (g867) & (g1870) & (g1875)));
	assign g1877 = (((!sk[23]) & (!g1592) & (!g1593) & (!g1605) & (g1668) & (!g56)) + ((!sk[23]) & (!g1592) & (!g1593) & (!g1605) & (g1668) & (g56)) + ((!sk[23]) & (!g1592) & (!g1593) & (g1605) & (!g1668) & (!g56)) + ((!sk[23]) & (!g1592) & (!g1593) & (g1605) & (!g1668) & (g56)) + ((!sk[23]) & (!g1592) & (!g1593) & (g1605) & (g1668) & (!g56)) + ((!sk[23]) & (!g1592) & (!g1593) & (g1605) & (g1668) & (g56)) + ((!sk[23]) & (!g1592) & (g1593) & (!g1605) & (!g1668) & (!g56)) + ((!sk[23]) & (!g1592) & (g1593) & (!g1605) & (!g1668) & (g56)) + ((!sk[23]) & (!g1592) & (g1593) & (!g1605) & (g1668) & (!g56)) + ((!sk[23]) & (!g1592) & (g1593) & (!g1605) & (g1668) & (g56)) + ((!sk[23]) & (!g1592) & (g1593) & (g1605) & (!g1668) & (!g56)) + ((!sk[23]) & (!g1592) & (g1593) & (g1605) & (!g1668) & (g56)) + ((!sk[23]) & (!g1592) & (g1593) & (g1605) & (g1668) & (!g56)) + ((!sk[23]) & (!g1592) & (g1593) & (g1605) & (g1668) & (g56)) + ((!sk[23]) & (g1592) & (!g1593) & (!g1605) & (g1668) & (!g56)) + ((!sk[23]) & (g1592) & (!g1593) & (!g1605) & (g1668) & (g56)) + ((!sk[23]) & (g1592) & (!g1593) & (g1605) & (!g1668) & (!g56)) + ((!sk[23]) & (g1592) & (!g1593) & (g1605) & (!g1668) & (g56)) + ((!sk[23]) & (g1592) & (!g1593) & (g1605) & (g1668) & (!g56)) + ((!sk[23]) & (g1592) & (!g1593) & (g1605) & (g1668) & (g56)) + ((!sk[23]) & (g1592) & (g1593) & (!g1605) & (!g1668) & (!g56)) + ((!sk[23]) & (g1592) & (g1593) & (!g1605) & (!g1668) & (g56)) + ((!sk[23]) & (g1592) & (g1593) & (!g1605) & (g1668) & (!g56)) + ((!sk[23]) & (g1592) & (g1593) & (!g1605) & (g1668) & (g56)) + ((!sk[23]) & (g1592) & (g1593) & (g1605) & (!g1668) & (!g56)) + ((!sk[23]) & (g1592) & (g1593) & (g1605) & (!g1668) & (g56)) + ((!sk[23]) & (g1592) & (g1593) & (g1605) & (g1668) & (!g56)) + ((!sk[23]) & (g1592) & (g1593) & (g1605) & (g1668) & (g56)) + ((sk[23]) & (!g1592) & (!g1593) & (!g1605) & (g1668) & (!g56)) + ((sk[23]) & (!g1592) & (!g1593) & (!g1605) & (g1668) & (g56)) + ((sk[23]) & (!g1592) & (!g1593) & (g1605) & (g1668) & (!g56)) + ((sk[23]) & (!g1592) & (!g1593) & (g1605) & (g1668) & (g56)) + ((sk[23]) & (!g1592) & (g1593) & (!g1605) & (g1668) & (!g56)) + ((sk[23]) & (!g1592) & (g1593) & (!g1605) & (g1668) & (g56)) + ((sk[23]) & (!g1592) & (g1593) & (g1605) & (g1668) & (!g56)) + ((sk[23]) & (!g1592) & (g1593) & (g1605) & (g1668) & (g56)) + ((sk[23]) & (g1592) & (!g1593) & (!g1605) & (g1668) & (!g56)) + ((sk[23]) & (g1592) & (!g1593) & (!g1605) & (g1668) & (g56)) + ((sk[23]) & (g1592) & (g1593) & (!g1605) & (!g1668) & (g56)) + ((sk[23]) & (g1592) & (g1593) & (!g1605) & (g1668) & (g56)) + ((sk[23]) & (g1592) & (g1593) & (g1605) & (!g1668) & (g56)) + ((sk[23]) & (g1592) & (g1593) & (g1605) & (g1668) & (g56)));
	assign g1878 = (((!g132) & (!g1812) & (!g1876) & (!sk[24]) & (g1877)) + ((!g132) & (!g1812) & (g1876) & (!sk[24]) & (!g1877)) + ((!g132) & (!g1812) & (g1876) & (!sk[24]) & (g1877)) + ((!g132) & (g1812) & (!g1876) & (!sk[24]) & (!g1877)) + ((!g132) & (g1812) & (!g1876) & (!sk[24]) & (g1877)) + ((!g132) & (g1812) & (!g1876) & (sk[24]) & (g1877)) + ((!g132) & (g1812) & (g1876) & (!sk[24]) & (!g1877)) + ((!g132) & (g1812) & (g1876) & (!sk[24]) & (g1877)) + ((!g132) & (g1812) & (g1876) & (sk[24]) & (g1877)) + ((g132) & (!g1812) & (!g1876) & (!sk[24]) & (g1877)) + ((g132) & (!g1812) & (g1876) & (!sk[24]) & (!g1877)) + ((g132) & (!g1812) & (g1876) & (!sk[24]) & (g1877)) + ((g132) & (g1812) & (!g1876) & (!sk[24]) & (!g1877)) + ((g132) & (g1812) & (!g1876) & (!sk[24]) & (g1877)) + ((g132) & (g1812) & (g1876) & (!sk[24]) & (!g1877)) + ((g132) & (g1812) & (g1876) & (!sk[24]) & (g1877)) + ((g132) & (g1812) & (g1876) & (sk[24]) & (!g1877)) + ((g132) & (g1812) & (g1876) & (sk[24]) & (g1877)));
	assign g1879 = (((!g1143) & (!g1148) & (!g1153) & (g1158) & (g677) & (g726)) + ((!g1143) & (!g1148) & (g1153) & (!g1158) & (!g677) & (g726)) + ((!g1143) & (!g1148) & (g1153) & (g1158) & (!g677) & (g726)) + ((!g1143) & (!g1148) & (g1153) & (g1158) & (g677) & (g726)) + ((!g1143) & (g1148) & (!g1153) & (!g1158) & (g677) & (!g726)) + ((!g1143) & (g1148) & (!g1153) & (g1158) & (g677) & (!g726)) + ((!g1143) & (g1148) & (!g1153) & (g1158) & (g677) & (g726)) + ((!g1143) & (g1148) & (g1153) & (!g1158) & (!g677) & (g726)) + ((!g1143) & (g1148) & (g1153) & (!g1158) & (g677) & (!g726)) + ((!g1143) & (g1148) & (g1153) & (g1158) & (!g677) & (g726)) + ((!g1143) & (g1148) & (g1153) & (g1158) & (g677) & (!g726)) + ((!g1143) & (g1148) & (g1153) & (g1158) & (g677) & (g726)) + ((g1143) & (!g1148) & (!g1153) & (!g1158) & (!g677) & (!g726)) + ((g1143) & (!g1148) & (!g1153) & (g1158) & (!g677) & (!g726)) + ((g1143) & (!g1148) & (!g1153) & (g1158) & (g677) & (g726)) + ((g1143) & (!g1148) & (g1153) & (!g1158) & (!g677) & (!g726)) + ((g1143) & (!g1148) & (g1153) & (!g1158) & (!g677) & (g726)) + ((g1143) & (!g1148) & (g1153) & (g1158) & (!g677) & (!g726)) + ((g1143) & (!g1148) & (g1153) & (g1158) & (!g677) & (g726)) + ((g1143) & (!g1148) & (g1153) & (g1158) & (g677) & (g726)) + ((g1143) & (g1148) & (!g1153) & (!g1158) & (!g677) & (!g726)) + ((g1143) & (g1148) & (!g1153) & (!g1158) & (g677) & (!g726)) + ((g1143) & (g1148) & (!g1153) & (g1158) & (!g677) & (!g726)) + ((g1143) & (g1148) & (!g1153) & (g1158) & (g677) & (!g726)) + ((g1143) & (g1148) & (!g1153) & (g1158) & (g677) & (g726)) + ((g1143) & (g1148) & (g1153) & (!g1158) & (!g677) & (!g726)) + ((g1143) & (g1148) & (g1153) & (!g1158) & (!g677) & (g726)) + ((g1143) & (g1148) & (g1153) & (!g1158) & (g677) & (!g726)) + ((g1143) & (g1148) & (g1153) & (g1158) & (!g677) & (!g726)) + ((g1143) & (g1148) & (g1153) & (g1158) & (!g677) & (g726)) + ((g1143) & (g1148) & (g1153) & (g1158) & (g677) & (!g726)) + ((g1143) & (g1148) & (g1153) & (g1158) & (g677) & (g726)));
	assign g1880 = (((!g1144) & (!g1149) & (!g1154) & (g1159) & (g677) & (g726)) + ((!g1144) & (!g1149) & (g1154) & (!g1159) & (!g677) & (g726)) + ((!g1144) & (!g1149) & (g1154) & (g1159) & (!g677) & (g726)) + ((!g1144) & (!g1149) & (g1154) & (g1159) & (g677) & (g726)) + ((!g1144) & (g1149) & (!g1154) & (!g1159) & (g677) & (!g726)) + ((!g1144) & (g1149) & (!g1154) & (g1159) & (g677) & (!g726)) + ((!g1144) & (g1149) & (!g1154) & (g1159) & (g677) & (g726)) + ((!g1144) & (g1149) & (g1154) & (!g1159) & (!g677) & (g726)) + ((!g1144) & (g1149) & (g1154) & (!g1159) & (g677) & (!g726)) + ((!g1144) & (g1149) & (g1154) & (g1159) & (!g677) & (g726)) + ((!g1144) & (g1149) & (g1154) & (g1159) & (g677) & (!g726)) + ((!g1144) & (g1149) & (g1154) & (g1159) & (g677) & (g726)) + ((g1144) & (!g1149) & (!g1154) & (!g1159) & (!g677) & (!g726)) + ((g1144) & (!g1149) & (!g1154) & (g1159) & (!g677) & (!g726)) + ((g1144) & (!g1149) & (!g1154) & (g1159) & (g677) & (g726)) + ((g1144) & (!g1149) & (g1154) & (!g1159) & (!g677) & (!g726)) + ((g1144) & (!g1149) & (g1154) & (!g1159) & (!g677) & (g726)) + ((g1144) & (!g1149) & (g1154) & (g1159) & (!g677) & (!g726)) + ((g1144) & (!g1149) & (g1154) & (g1159) & (!g677) & (g726)) + ((g1144) & (!g1149) & (g1154) & (g1159) & (g677) & (g726)) + ((g1144) & (g1149) & (!g1154) & (!g1159) & (!g677) & (!g726)) + ((g1144) & (g1149) & (!g1154) & (!g1159) & (g677) & (!g726)) + ((g1144) & (g1149) & (!g1154) & (g1159) & (!g677) & (!g726)) + ((g1144) & (g1149) & (!g1154) & (g1159) & (g677) & (!g726)) + ((g1144) & (g1149) & (!g1154) & (g1159) & (g677) & (g726)) + ((g1144) & (g1149) & (g1154) & (!g1159) & (!g677) & (!g726)) + ((g1144) & (g1149) & (g1154) & (!g1159) & (!g677) & (g726)) + ((g1144) & (g1149) & (g1154) & (!g1159) & (g677) & (!g726)) + ((g1144) & (g1149) & (g1154) & (g1159) & (!g677) & (!g726)) + ((g1144) & (g1149) & (g1154) & (g1159) & (!g677) & (g726)) + ((g1144) & (g1149) & (g1154) & (g1159) & (g677) & (!g726)) + ((g1144) & (g1149) & (g1154) & (g1159) & (g677) & (g726)));
	assign g1881 = (((!g1145) & (!g1150) & (!g1155) & (g1160) & (g677) & (g726)) + ((!g1145) & (!g1150) & (g1155) & (!g1160) & (!g677) & (g726)) + ((!g1145) & (!g1150) & (g1155) & (g1160) & (!g677) & (g726)) + ((!g1145) & (!g1150) & (g1155) & (g1160) & (g677) & (g726)) + ((!g1145) & (g1150) & (!g1155) & (!g1160) & (g677) & (!g726)) + ((!g1145) & (g1150) & (!g1155) & (g1160) & (g677) & (!g726)) + ((!g1145) & (g1150) & (!g1155) & (g1160) & (g677) & (g726)) + ((!g1145) & (g1150) & (g1155) & (!g1160) & (!g677) & (g726)) + ((!g1145) & (g1150) & (g1155) & (!g1160) & (g677) & (!g726)) + ((!g1145) & (g1150) & (g1155) & (g1160) & (!g677) & (g726)) + ((!g1145) & (g1150) & (g1155) & (g1160) & (g677) & (!g726)) + ((!g1145) & (g1150) & (g1155) & (g1160) & (g677) & (g726)) + ((g1145) & (!g1150) & (!g1155) & (!g1160) & (!g677) & (!g726)) + ((g1145) & (!g1150) & (!g1155) & (g1160) & (!g677) & (!g726)) + ((g1145) & (!g1150) & (!g1155) & (g1160) & (g677) & (g726)) + ((g1145) & (!g1150) & (g1155) & (!g1160) & (!g677) & (!g726)) + ((g1145) & (!g1150) & (g1155) & (!g1160) & (!g677) & (g726)) + ((g1145) & (!g1150) & (g1155) & (g1160) & (!g677) & (!g726)) + ((g1145) & (!g1150) & (g1155) & (g1160) & (!g677) & (g726)) + ((g1145) & (!g1150) & (g1155) & (g1160) & (g677) & (g726)) + ((g1145) & (g1150) & (!g1155) & (!g1160) & (!g677) & (!g726)) + ((g1145) & (g1150) & (!g1155) & (!g1160) & (g677) & (!g726)) + ((g1145) & (g1150) & (!g1155) & (g1160) & (!g677) & (!g726)) + ((g1145) & (g1150) & (!g1155) & (g1160) & (g677) & (!g726)) + ((g1145) & (g1150) & (!g1155) & (g1160) & (g677) & (g726)) + ((g1145) & (g1150) & (g1155) & (!g1160) & (!g677) & (!g726)) + ((g1145) & (g1150) & (g1155) & (!g1160) & (!g677) & (g726)) + ((g1145) & (g1150) & (g1155) & (!g1160) & (g677) & (!g726)) + ((g1145) & (g1150) & (g1155) & (g1160) & (!g677) & (!g726)) + ((g1145) & (g1150) & (g1155) & (g1160) & (!g677) & (g726)) + ((g1145) & (g1150) & (g1155) & (g1160) & (g677) & (!g726)) + ((g1145) & (g1150) & (g1155) & (g1160) & (g677) & (g726)));
	assign g1882 = (((!g1146) & (!g1151) & (!g1156) & (g1161) & (g677) & (g726)) + ((!g1146) & (!g1151) & (g1156) & (!g1161) & (!g677) & (g726)) + ((!g1146) & (!g1151) & (g1156) & (g1161) & (!g677) & (g726)) + ((!g1146) & (!g1151) & (g1156) & (g1161) & (g677) & (g726)) + ((!g1146) & (g1151) & (!g1156) & (!g1161) & (g677) & (!g726)) + ((!g1146) & (g1151) & (!g1156) & (g1161) & (g677) & (!g726)) + ((!g1146) & (g1151) & (!g1156) & (g1161) & (g677) & (g726)) + ((!g1146) & (g1151) & (g1156) & (!g1161) & (!g677) & (g726)) + ((!g1146) & (g1151) & (g1156) & (!g1161) & (g677) & (!g726)) + ((!g1146) & (g1151) & (g1156) & (g1161) & (!g677) & (g726)) + ((!g1146) & (g1151) & (g1156) & (g1161) & (g677) & (!g726)) + ((!g1146) & (g1151) & (g1156) & (g1161) & (g677) & (g726)) + ((g1146) & (!g1151) & (!g1156) & (!g1161) & (!g677) & (!g726)) + ((g1146) & (!g1151) & (!g1156) & (g1161) & (!g677) & (!g726)) + ((g1146) & (!g1151) & (!g1156) & (g1161) & (g677) & (g726)) + ((g1146) & (!g1151) & (g1156) & (!g1161) & (!g677) & (!g726)) + ((g1146) & (!g1151) & (g1156) & (!g1161) & (!g677) & (g726)) + ((g1146) & (!g1151) & (g1156) & (g1161) & (!g677) & (!g726)) + ((g1146) & (!g1151) & (g1156) & (g1161) & (!g677) & (g726)) + ((g1146) & (!g1151) & (g1156) & (g1161) & (g677) & (g726)) + ((g1146) & (g1151) & (!g1156) & (!g1161) & (!g677) & (!g726)) + ((g1146) & (g1151) & (!g1156) & (!g1161) & (g677) & (!g726)) + ((g1146) & (g1151) & (!g1156) & (g1161) & (!g677) & (!g726)) + ((g1146) & (g1151) & (!g1156) & (g1161) & (g677) & (!g726)) + ((g1146) & (g1151) & (!g1156) & (g1161) & (g677) & (g726)) + ((g1146) & (g1151) & (g1156) & (!g1161) & (!g677) & (!g726)) + ((g1146) & (g1151) & (g1156) & (!g1161) & (!g677) & (g726)) + ((g1146) & (g1151) & (g1156) & (!g1161) & (g677) & (!g726)) + ((g1146) & (g1151) & (g1156) & (g1161) & (!g677) & (!g726)) + ((g1146) & (g1151) & (g1156) & (g1161) & (!g677) & (g726)) + ((g1146) & (g1151) & (g1156) & (g1161) & (g677) & (!g726)) + ((g1146) & (g1151) & (g1156) & (g1161) & (g677) & (g726)));
	assign g1883 = (((!g1879) & (!g1880) & (!g1881) & (g1882) & (g820) & (g773)) + ((!g1879) & (!g1880) & (g1881) & (!g1882) & (!g820) & (g773)) + ((!g1879) & (!g1880) & (g1881) & (g1882) & (!g820) & (g773)) + ((!g1879) & (!g1880) & (g1881) & (g1882) & (g820) & (g773)) + ((!g1879) & (g1880) & (!g1881) & (!g1882) & (g820) & (!g773)) + ((!g1879) & (g1880) & (!g1881) & (g1882) & (g820) & (!g773)) + ((!g1879) & (g1880) & (!g1881) & (g1882) & (g820) & (g773)) + ((!g1879) & (g1880) & (g1881) & (!g1882) & (!g820) & (g773)) + ((!g1879) & (g1880) & (g1881) & (!g1882) & (g820) & (!g773)) + ((!g1879) & (g1880) & (g1881) & (g1882) & (!g820) & (g773)) + ((!g1879) & (g1880) & (g1881) & (g1882) & (g820) & (!g773)) + ((!g1879) & (g1880) & (g1881) & (g1882) & (g820) & (g773)) + ((g1879) & (!g1880) & (!g1881) & (!g1882) & (!g820) & (!g773)) + ((g1879) & (!g1880) & (!g1881) & (g1882) & (!g820) & (!g773)) + ((g1879) & (!g1880) & (!g1881) & (g1882) & (g820) & (g773)) + ((g1879) & (!g1880) & (g1881) & (!g1882) & (!g820) & (!g773)) + ((g1879) & (!g1880) & (g1881) & (!g1882) & (!g820) & (g773)) + ((g1879) & (!g1880) & (g1881) & (g1882) & (!g820) & (!g773)) + ((g1879) & (!g1880) & (g1881) & (g1882) & (!g820) & (g773)) + ((g1879) & (!g1880) & (g1881) & (g1882) & (g820) & (g773)) + ((g1879) & (g1880) & (!g1881) & (!g1882) & (!g820) & (!g773)) + ((g1879) & (g1880) & (!g1881) & (!g1882) & (g820) & (!g773)) + ((g1879) & (g1880) & (!g1881) & (g1882) & (!g820) & (!g773)) + ((g1879) & (g1880) & (!g1881) & (g1882) & (g820) & (!g773)) + ((g1879) & (g1880) & (!g1881) & (g1882) & (g820) & (g773)) + ((g1879) & (g1880) & (g1881) & (!g1882) & (!g820) & (!g773)) + ((g1879) & (g1880) & (g1881) & (!g1882) & (!g820) & (g773)) + ((g1879) & (g1880) & (g1881) & (!g1882) & (g820) & (!g773)) + ((g1879) & (g1880) & (g1881) & (g1882) & (!g820) & (!g773)) + ((g1879) & (g1880) & (g1881) & (g1882) & (!g820) & (g773)) + ((g1879) & (g1880) & (g1881) & (g1882) & (g820) & (!g773)) + ((g1879) & (g1880) & (g1881) & (g1882) & (g820) & (g773)));
	assign g1884 = (((!g1164) & (!g1165) & (!g1166) & (g1167) & (g677) & (g726)) + ((!g1164) & (!g1165) & (g1166) & (!g1167) & (!g677) & (g726)) + ((!g1164) & (!g1165) & (g1166) & (g1167) & (!g677) & (g726)) + ((!g1164) & (!g1165) & (g1166) & (g1167) & (g677) & (g726)) + ((!g1164) & (g1165) & (!g1166) & (!g1167) & (g677) & (!g726)) + ((!g1164) & (g1165) & (!g1166) & (g1167) & (g677) & (!g726)) + ((!g1164) & (g1165) & (!g1166) & (g1167) & (g677) & (g726)) + ((!g1164) & (g1165) & (g1166) & (!g1167) & (!g677) & (g726)) + ((!g1164) & (g1165) & (g1166) & (!g1167) & (g677) & (!g726)) + ((!g1164) & (g1165) & (g1166) & (g1167) & (!g677) & (g726)) + ((!g1164) & (g1165) & (g1166) & (g1167) & (g677) & (!g726)) + ((!g1164) & (g1165) & (g1166) & (g1167) & (g677) & (g726)) + ((g1164) & (!g1165) & (!g1166) & (!g1167) & (!g677) & (!g726)) + ((g1164) & (!g1165) & (!g1166) & (g1167) & (!g677) & (!g726)) + ((g1164) & (!g1165) & (!g1166) & (g1167) & (g677) & (g726)) + ((g1164) & (!g1165) & (g1166) & (!g1167) & (!g677) & (!g726)) + ((g1164) & (!g1165) & (g1166) & (!g1167) & (!g677) & (g726)) + ((g1164) & (!g1165) & (g1166) & (g1167) & (!g677) & (!g726)) + ((g1164) & (!g1165) & (g1166) & (g1167) & (!g677) & (g726)) + ((g1164) & (!g1165) & (g1166) & (g1167) & (g677) & (g726)) + ((g1164) & (g1165) & (!g1166) & (!g1167) & (!g677) & (!g726)) + ((g1164) & (g1165) & (!g1166) & (!g1167) & (g677) & (!g726)) + ((g1164) & (g1165) & (!g1166) & (g1167) & (!g677) & (!g726)) + ((g1164) & (g1165) & (!g1166) & (g1167) & (g677) & (!g726)) + ((g1164) & (g1165) & (!g1166) & (g1167) & (g677) & (g726)) + ((g1164) & (g1165) & (g1166) & (!g1167) & (!g677) & (!g726)) + ((g1164) & (g1165) & (g1166) & (!g1167) & (!g677) & (g726)) + ((g1164) & (g1165) & (g1166) & (!g1167) & (g677) & (!g726)) + ((g1164) & (g1165) & (g1166) & (g1167) & (!g677) & (!g726)) + ((g1164) & (g1165) & (g1166) & (g1167) & (!g677) & (g726)) + ((g1164) & (g1165) & (g1166) & (g1167) & (g677) & (!g726)) + ((g1164) & (g1165) & (g1166) & (g1167) & (g677) & (g726)));
	assign g1885 = (((!g677) & (!sk[31]) & (!g726) & (!g1169) & (g1170) & (!g1171)) + ((!g677) & (!sk[31]) & (!g726) & (!g1169) & (g1170) & (g1171)) + ((!g677) & (!sk[31]) & (!g726) & (g1169) & (!g1170) & (!g1171)) + ((!g677) & (!sk[31]) & (!g726) & (g1169) & (!g1170) & (g1171)) + ((!g677) & (!sk[31]) & (!g726) & (g1169) & (g1170) & (!g1171)) + ((!g677) & (!sk[31]) & (!g726) & (g1169) & (g1170) & (g1171)) + ((!g677) & (!sk[31]) & (g726) & (!g1169) & (!g1170) & (!g1171)) + ((!g677) & (!sk[31]) & (g726) & (!g1169) & (!g1170) & (g1171)) + ((!g677) & (!sk[31]) & (g726) & (!g1169) & (g1170) & (!g1171)) + ((!g677) & (!sk[31]) & (g726) & (!g1169) & (g1170) & (g1171)) + ((!g677) & (!sk[31]) & (g726) & (g1169) & (!g1170) & (!g1171)) + ((!g677) & (!sk[31]) & (g726) & (g1169) & (!g1170) & (g1171)) + ((!g677) & (!sk[31]) & (g726) & (g1169) & (g1170) & (!g1171)) + ((!g677) & (!sk[31]) & (g726) & (g1169) & (g1170) & (g1171)) + ((!g677) & (sk[31]) & (g726) & (!g1169) & (!g1170) & (g1171)) + ((!g677) & (sk[31]) & (g726) & (!g1169) & (g1170) & (g1171)) + ((!g677) & (sk[31]) & (g726) & (g1169) & (!g1170) & (g1171)) + ((!g677) & (sk[31]) & (g726) & (g1169) & (g1170) & (g1171)) + ((g677) & (!sk[31]) & (!g726) & (!g1169) & (g1170) & (!g1171)) + ((g677) & (!sk[31]) & (!g726) & (!g1169) & (g1170) & (g1171)) + ((g677) & (!sk[31]) & (!g726) & (g1169) & (!g1170) & (!g1171)) + ((g677) & (!sk[31]) & (!g726) & (g1169) & (!g1170) & (g1171)) + ((g677) & (!sk[31]) & (!g726) & (g1169) & (g1170) & (!g1171)) + ((g677) & (!sk[31]) & (!g726) & (g1169) & (g1170) & (g1171)) + ((g677) & (!sk[31]) & (g726) & (!g1169) & (!g1170) & (!g1171)) + ((g677) & (!sk[31]) & (g726) & (!g1169) & (!g1170) & (g1171)) + ((g677) & (!sk[31]) & (g726) & (!g1169) & (g1170) & (!g1171)) + ((g677) & (!sk[31]) & (g726) & (!g1169) & (g1170) & (g1171)) + ((g677) & (!sk[31]) & (g726) & (g1169) & (!g1170) & (!g1171)) + ((g677) & (!sk[31]) & (g726) & (g1169) & (!g1170) & (g1171)) + ((g677) & (!sk[31]) & (g726) & (g1169) & (g1170) & (!g1171)) + ((g677) & (!sk[31]) & (g726) & (g1169) & (g1170) & (g1171)) + ((g677) & (sk[31]) & (!g726) & (g1169) & (!g1170) & (!g1171)) + ((g677) & (sk[31]) & (!g726) & (g1169) & (!g1170) & (g1171)) + ((g677) & (sk[31]) & (!g726) & (g1169) & (g1170) & (!g1171)) + ((g677) & (sk[31]) & (!g726) & (g1169) & (g1170) & (g1171)) + ((g677) & (sk[31]) & (g726) & (!g1169) & (g1170) & (!g1171)) + ((g677) & (sk[31]) & (g726) & (!g1169) & (g1170) & (g1171)) + ((g677) & (sk[31]) & (g726) & (g1169) & (g1170) & (!g1171)) + ((g677) & (sk[31]) & (g726) & (g1169) & (g1170) & (g1171)));
	assign g1886 = (((!g1173) & (!g1174) & (!g1175) & (g1176) & (g677) & (g726)) + ((!g1173) & (!g1174) & (g1175) & (!g1176) & (!g677) & (g726)) + ((!g1173) & (!g1174) & (g1175) & (g1176) & (!g677) & (g726)) + ((!g1173) & (!g1174) & (g1175) & (g1176) & (g677) & (g726)) + ((!g1173) & (g1174) & (!g1175) & (!g1176) & (g677) & (!g726)) + ((!g1173) & (g1174) & (!g1175) & (g1176) & (g677) & (!g726)) + ((!g1173) & (g1174) & (!g1175) & (g1176) & (g677) & (g726)) + ((!g1173) & (g1174) & (g1175) & (!g1176) & (!g677) & (g726)) + ((!g1173) & (g1174) & (g1175) & (!g1176) & (g677) & (!g726)) + ((!g1173) & (g1174) & (g1175) & (g1176) & (!g677) & (g726)) + ((!g1173) & (g1174) & (g1175) & (g1176) & (g677) & (!g726)) + ((!g1173) & (g1174) & (g1175) & (g1176) & (g677) & (g726)) + ((g1173) & (!g1174) & (!g1175) & (!g1176) & (!g677) & (!g726)) + ((g1173) & (!g1174) & (!g1175) & (g1176) & (!g677) & (!g726)) + ((g1173) & (!g1174) & (!g1175) & (g1176) & (g677) & (g726)) + ((g1173) & (!g1174) & (g1175) & (!g1176) & (!g677) & (!g726)) + ((g1173) & (!g1174) & (g1175) & (!g1176) & (!g677) & (g726)) + ((g1173) & (!g1174) & (g1175) & (g1176) & (!g677) & (!g726)) + ((g1173) & (!g1174) & (g1175) & (g1176) & (!g677) & (g726)) + ((g1173) & (!g1174) & (g1175) & (g1176) & (g677) & (g726)) + ((g1173) & (g1174) & (!g1175) & (!g1176) & (!g677) & (!g726)) + ((g1173) & (g1174) & (!g1175) & (!g1176) & (g677) & (!g726)) + ((g1173) & (g1174) & (!g1175) & (g1176) & (!g677) & (!g726)) + ((g1173) & (g1174) & (!g1175) & (g1176) & (g677) & (!g726)) + ((g1173) & (g1174) & (!g1175) & (g1176) & (g677) & (g726)) + ((g1173) & (g1174) & (g1175) & (!g1176) & (!g677) & (!g726)) + ((g1173) & (g1174) & (g1175) & (!g1176) & (!g677) & (g726)) + ((g1173) & (g1174) & (g1175) & (!g1176) & (g677) & (!g726)) + ((g1173) & (g1174) & (g1175) & (g1176) & (!g677) & (!g726)) + ((g1173) & (g1174) & (g1175) & (g1176) & (!g677) & (g726)) + ((g1173) & (g1174) & (g1175) & (g1176) & (g677) & (!g726)) + ((g1173) & (g1174) & (g1175) & (g1176) & (g677) & (g726)));
	assign g1887 = (((!g1178) & (!g1179) & (!g1180) & (g1181) & (g677) & (g726)) + ((!g1178) & (!g1179) & (g1180) & (!g1181) & (!g677) & (g726)) + ((!g1178) & (!g1179) & (g1180) & (g1181) & (!g677) & (g726)) + ((!g1178) & (!g1179) & (g1180) & (g1181) & (g677) & (g726)) + ((!g1178) & (g1179) & (!g1180) & (!g1181) & (g677) & (!g726)) + ((!g1178) & (g1179) & (!g1180) & (g1181) & (g677) & (!g726)) + ((!g1178) & (g1179) & (!g1180) & (g1181) & (g677) & (g726)) + ((!g1178) & (g1179) & (g1180) & (!g1181) & (!g677) & (g726)) + ((!g1178) & (g1179) & (g1180) & (!g1181) & (g677) & (!g726)) + ((!g1178) & (g1179) & (g1180) & (g1181) & (!g677) & (g726)) + ((!g1178) & (g1179) & (g1180) & (g1181) & (g677) & (!g726)) + ((!g1178) & (g1179) & (g1180) & (g1181) & (g677) & (g726)) + ((g1178) & (!g1179) & (!g1180) & (!g1181) & (!g677) & (!g726)) + ((g1178) & (!g1179) & (!g1180) & (g1181) & (!g677) & (!g726)) + ((g1178) & (!g1179) & (!g1180) & (g1181) & (g677) & (g726)) + ((g1178) & (!g1179) & (g1180) & (!g1181) & (!g677) & (!g726)) + ((g1178) & (!g1179) & (g1180) & (!g1181) & (!g677) & (g726)) + ((g1178) & (!g1179) & (g1180) & (g1181) & (!g677) & (!g726)) + ((g1178) & (!g1179) & (g1180) & (g1181) & (!g677) & (g726)) + ((g1178) & (!g1179) & (g1180) & (g1181) & (g677) & (g726)) + ((g1178) & (g1179) & (!g1180) & (!g1181) & (!g677) & (!g726)) + ((g1178) & (g1179) & (!g1180) & (!g1181) & (g677) & (!g726)) + ((g1178) & (g1179) & (!g1180) & (g1181) & (!g677) & (!g726)) + ((g1178) & (g1179) & (!g1180) & (g1181) & (g677) & (!g726)) + ((g1178) & (g1179) & (!g1180) & (g1181) & (g677) & (g726)) + ((g1178) & (g1179) & (g1180) & (!g1181) & (!g677) & (!g726)) + ((g1178) & (g1179) & (g1180) & (!g1181) & (!g677) & (g726)) + ((g1178) & (g1179) & (g1180) & (!g1181) & (g677) & (!g726)) + ((g1178) & (g1179) & (g1180) & (g1181) & (!g677) & (!g726)) + ((g1178) & (g1179) & (g1180) & (g1181) & (!g677) & (g726)) + ((g1178) & (g1179) & (g1180) & (g1181) & (g677) & (!g726)) + ((g1178) & (g1179) & (g1180) & (g1181) & (g677) & (g726)));
	assign g1888 = (((!g820) & (!g773) & (!g1884) & (g1885) & (!g1886) & (!g1887)) + ((!g820) & (!g773) & (!g1884) & (g1885) & (!g1886) & (g1887)) + ((!g820) & (!g773) & (!g1884) & (g1885) & (g1886) & (!g1887)) + ((!g820) & (!g773) & (!g1884) & (g1885) & (g1886) & (g1887)) + ((!g820) & (!g773) & (g1884) & (g1885) & (!g1886) & (!g1887)) + ((!g820) & (!g773) & (g1884) & (g1885) & (!g1886) & (g1887)) + ((!g820) & (!g773) & (g1884) & (g1885) & (g1886) & (!g1887)) + ((!g820) & (!g773) & (g1884) & (g1885) & (g1886) & (g1887)) + ((!g820) & (g773) & (!g1884) & (!g1885) & (!g1886) & (g1887)) + ((!g820) & (g773) & (!g1884) & (!g1885) & (g1886) & (g1887)) + ((!g820) & (g773) & (!g1884) & (g1885) & (!g1886) & (g1887)) + ((!g820) & (g773) & (!g1884) & (g1885) & (g1886) & (g1887)) + ((!g820) & (g773) & (g1884) & (!g1885) & (!g1886) & (g1887)) + ((!g820) & (g773) & (g1884) & (!g1885) & (g1886) & (g1887)) + ((!g820) & (g773) & (g1884) & (g1885) & (!g1886) & (g1887)) + ((!g820) & (g773) & (g1884) & (g1885) & (g1886) & (g1887)) + ((g820) & (!g773) & (g1884) & (!g1885) & (!g1886) & (!g1887)) + ((g820) & (!g773) & (g1884) & (!g1885) & (!g1886) & (g1887)) + ((g820) & (!g773) & (g1884) & (!g1885) & (g1886) & (!g1887)) + ((g820) & (!g773) & (g1884) & (!g1885) & (g1886) & (g1887)) + ((g820) & (!g773) & (g1884) & (g1885) & (!g1886) & (!g1887)) + ((g820) & (!g773) & (g1884) & (g1885) & (!g1886) & (g1887)) + ((g820) & (!g773) & (g1884) & (g1885) & (g1886) & (!g1887)) + ((g820) & (!g773) & (g1884) & (g1885) & (g1886) & (g1887)) + ((g820) & (g773) & (!g1884) & (!g1885) & (g1886) & (!g1887)) + ((g820) & (g773) & (!g1884) & (!g1885) & (g1886) & (g1887)) + ((g820) & (g773) & (!g1884) & (g1885) & (g1886) & (!g1887)) + ((g820) & (g773) & (!g1884) & (g1885) & (g1886) & (g1887)) + ((g820) & (g773) & (g1884) & (!g1885) & (g1886) & (!g1887)) + ((g820) & (g773) & (g1884) & (!g1885) & (g1886) & (g1887)) + ((g820) & (g773) & (g1884) & (g1885) & (g1886) & (!g1887)) + ((g820) & (g773) & (g1884) & (g1885) & (g1886) & (g1887)));
	assign g1889 = (((!sk[35]) & (!g867) & (!g1883) & (g1888)) + ((!sk[35]) & (!g867) & (g1883) & (!g1888)) + ((!sk[35]) & (!g867) & (g1883) & (g1888)) + ((!sk[35]) & (g867) & (!g1883) & (g1888)) + ((!sk[35]) & (g867) & (g1883) & (!g1888)) + ((!sk[35]) & (g867) & (g1883) & (g1888)) + ((sk[35]) & (!g867) & (!g1883) & (g1888)) + ((sk[35]) & (!g867) & (g1883) & (g1888)) + ((sk[35]) & (g867) & (g1883) & (!g1888)) + ((sk[35]) & (g867) & (g1883) & (g1888)));
	assign g1890 = (((!g1592) & (!g1593) & (!g1605) & (!sk[36]) & (g1680) & (!g57)) + ((!g1592) & (!g1593) & (!g1605) & (!sk[36]) & (g1680) & (g57)) + ((!g1592) & (!g1593) & (!g1605) & (sk[36]) & (g1680) & (!g57)) + ((!g1592) & (!g1593) & (!g1605) & (sk[36]) & (g1680) & (g57)) + ((!g1592) & (!g1593) & (g1605) & (!sk[36]) & (!g1680) & (!g57)) + ((!g1592) & (!g1593) & (g1605) & (!sk[36]) & (!g1680) & (g57)) + ((!g1592) & (!g1593) & (g1605) & (!sk[36]) & (g1680) & (!g57)) + ((!g1592) & (!g1593) & (g1605) & (!sk[36]) & (g1680) & (g57)) + ((!g1592) & (!g1593) & (g1605) & (sk[36]) & (g1680) & (!g57)) + ((!g1592) & (!g1593) & (g1605) & (sk[36]) & (g1680) & (g57)) + ((!g1592) & (g1593) & (!g1605) & (!sk[36]) & (!g1680) & (!g57)) + ((!g1592) & (g1593) & (!g1605) & (!sk[36]) & (!g1680) & (g57)) + ((!g1592) & (g1593) & (!g1605) & (!sk[36]) & (g1680) & (!g57)) + ((!g1592) & (g1593) & (!g1605) & (!sk[36]) & (g1680) & (g57)) + ((!g1592) & (g1593) & (!g1605) & (sk[36]) & (g1680) & (!g57)) + ((!g1592) & (g1593) & (!g1605) & (sk[36]) & (g1680) & (g57)) + ((!g1592) & (g1593) & (g1605) & (!sk[36]) & (!g1680) & (!g57)) + ((!g1592) & (g1593) & (g1605) & (!sk[36]) & (!g1680) & (g57)) + ((!g1592) & (g1593) & (g1605) & (!sk[36]) & (g1680) & (!g57)) + ((!g1592) & (g1593) & (g1605) & (!sk[36]) & (g1680) & (g57)) + ((!g1592) & (g1593) & (g1605) & (sk[36]) & (g1680) & (!g57)) + ((!g1592) & (g1593) & (g1605) & (sk[36]) & (g1680) & (g57)) + ((g1592) & (!g1593) & (!g1605) & (!sk[36]) & (g1680) & (!g57)) + ((g1592) & (!g1593) & (!g1605) & (!sk[36]) & (g1680) & (g57)) + ((g1592) & (!g1593) & (!g1605) & (sk[36]) & (g1680) & (!g57)) + ((g1592) & (!g1593) & (!g1605) & (sk[36]) & (g1680) & (g57)) + ((g1592) & (!g1593) & (g1605) & (!sk[36]) & (!g1680) & (!g57)) + ((g1592) & (!g1593) & (g1605) & (!sk[36]) & (!g1680) & (g57)) + ((g1592) & (!g1593) & (g1605) & (!sk[36]) & (g1680) & (!g57)) + ((g1592) & (!g1593) & (g1605) & (!sk[36]) & (g1680) & (g57)) + ((g1592) & (g1593) & (!g1605) & (!sk[36]) & (!g1680) & (!g57)) + ((g1592) & (g1593) & (!g1605) & (!sk[36]) & (!g1680) & (g57)) + ((g1592) & (g1593) & (!g1605) & (!sk[36]) & (g1680) & (!g57)) + ((g1592) & (g1593) & (!g1605) & (!sk[36]) & (g1680) & (g57)) + ((g1592) & (g1593) & (!g1605) & (sk[36]) & (!g1680) & (g57)) + ((g1592) & (g1593) & (!g1605) & (sk[36]) & (g1680) & (g57)) + ((g1592) & (g1593) & (g1605) & (!sk[36]) & (!g1680) & (!g57)) + ((g1592) & (g1593) & (g1605) & (!sk[36]) & (!g1680) & (g57)) + ((g1592) & (g1593) & (g1605) & (!sk[36]) & (g1680) & (!g57)) + ((g1592) & (g1593) & (g1605) & (!sk[36]) & (g1680) & (g57)) + ((g1592) & (g1593) & (g1605) & (sk[36]) & (!g1680) & (g57)) + ((g1592) & (g1593) & (g1605) & (sk[36]) & (g1680) & (g57)));
	assign g1891 = (((!g132) & (!g1812) & (!sk[37]) & (!g1889) & (g1890)) + ((!g132) & (!g1812) & (!sk[37]) & (g1889) & (!g1890)) + ((!g132) & (!g1812) & (!sk[37]) & (g1889) & (g1890)) + ((!g132) & (g1812) & (!sk[37]) & (!g1889) & (!g1890)) + ((!g132) & (g1812) & (!sk[37]) & (!g1889) & (g1890)) + ((!g132) & (g1812) & (!sk[37]) & (g1889) & (!g1890)) + ((!g132) & (g1812) & (!sk[37]) & (g1889) & (g1890)) + ((!g132) & (g1812) & (sk[37]) & (!g1889) & (g1890)) + ((!g132) & (g1812) & (sk[37]) & (g1889) & (g1890)) + ((g132) & (!g1812) & (!sk[37]) & (!g1889) & (g1890)) + ((g132) & (!g1812) & (!sk[37]) & (g1889) & (!g1890)) + ((g132) & (!g1812) & (!sk[37]) & (g1889) & (g1890)) + ((g132) & (g1812) & (!sk[37]) & (!g1889) & (!g1890)) + ((g132) & (g1812) & (!sk[37]) & (!g1889) & (g1890)) + ((g132) & (g1812) & (!sk[37]) & (g1889) & (!g1890)) + ((g132) & (g1812) & (!sk[37]) & (g1889) & (g1890)) + ((g132) & (g1812) & (sk[37]) & (g1889) & (!g1890)) + ((g132) & (g1812) & (sk[37]) & (g1889) & (g1890)));
	assign g1892 = (((!g1188) & (!g1189) & (!g1190) & (g1191) & (g820) & (g773)) + ((!g1188) & (!g1189) & (g1190) & (!g1191) & (!g820) & (g773)) + ((!g1188) & (!g1189) & (g1190) & (g1191) & (!g820) & (g773)) + ((!g1188) & (!g1189) & (g1190) & (g1191) & (g820) & (g773)) + ((!g1188) & (g1189) & (!g1190) & (!g1191) & (g820) & (!g773)) + ((!g1188) & (g1189) & (!g1190) & (g1191) & (g820) & (!g773)) + ((!g1188) & (g1189) & (!g1190) & (g1191) & (g820) & (g773)) + ((!g1188) & (g1189) & (g1190) & (!g1191) & (!g820) & (g773)) + ((!g1188) & (g1189) & (g1190) & (!g1191) & (g820) & (!g773)) + ((!g1188) & (g1189) & (g1190) & (g1191) & (!g820) & (g773)) + ((!g1188) & (g1189) & (g1190) & (g1191) & (g820) & (!g773)) + ((!g1188) & (g1189) & (g1190) & (g1191) & (g820) & (g773)) + ((g1188) & (!g1189) & (!g1190) & (!g1191) & (!g820) & (!g773)) + ((g1188) & (!g1189) & (!g1190) & (g1191) & (!g820) & (!g773)) + ((g1188) & (!g1189) & (!g1190) & (g1191) & (g820) & (g773)) + ((g1188) & (!g1189) & (g1190) & (!g1191) & (!g820) & (!g773)) + ((g1188) & (!g1189) & (g1190) & (!g1191) & (!g820) & (g773)) + ((g1188) & (!g1189) & (g1190) & (g1191) & (!g820) & (!g773)) + ((g1188) & (!g1189) & (g1190) & (g1191) & (!g820) & (g773)) + ((g1188) & (!g1189) & (g1190) & (g1191) & (g820) & (g773)) + ((g1188) & (g1189) & (!g1190) & (!g1191) & (!g820) & (!g773)) + ((g1188) & (g1189) & (!g1190) & (!g1191) & (g820) & (!g773)) + ((g1188) & (g1189) & (!g1190) & (g1191) & (!g820) & (!g773)) + ((g1188) & (g1189) & (!g1190) & (g1191) & (g820) & (!g773)) + ((g1188) & (g1189) & (!g1190) & (g1191) & (g820) & (g773)) + ((g1188) & (g1189) & (g1190) & (!g1191) & (!g820) & (!g773)) + ((g1188) & (g1189) & (g1190) & (!g1191) & (!g820) & (g773)) + ((g1188) & (g1189) & (g1190) & (!g1191) & (g820) & (!g773)) + ((g1188) & (g1189) & (g1190) & (g1191) & (!g820) & (!g773)) + ((g1188) & (g1189) & (g1190) & (g1191) & (!g820) & (g773)) + ((g1188) & (g1189) & (g1190) & (g1191) & (g820) & (!g773)) + ((g1188) & (g1189) & (g1190) & (g1191) & (g820) & (g773)));
	assign g1893 = (((!g1193) & (!g1194) & (!g1195) & (g1196) & (g820) & (g773)) + ((!g1193) & (!g1194) & (g1195) & (!g1196) & (!g820) & (g773)) + ((!g1193) & (!g1194) & (g1195) & (g1196) & (!g820) & (g773)) + ((!g1193) & (!g1194) & (g1195) & (g1196) & (g820) & (g773)) + ((!g1193) & (g1194) & (!g1195) & (!g1196) & (g820) & (!g773)) + ((!g1193) & (g1194) & (!g1195) & (g1196) & (g820) & (!g773)) + ((!g1193) & (g1194) & (!g1195) & (g1196) & (g820) & (g773)) + ((!g1193) & (g1194) & (g1195) & (!g1196) & (!g820) & (g773)) + ((!g1193) & (g1194) & (g1195) & (!g1196) & (g820) & (!g773)) + ((!g1193) & (g1194) & (g1195) & (g1196) & (!g820) & (g773)) + ((!g1193) & (g1194) & (g1195) & (g1196) & (g820) & (!g773)) + ((!g1193) & (g1194) & (g1195) & (g1196) & (g820) & (g773)) + ((g1193) & (!g1194) & (!g1195) & (!g1196) & (!g820) & (!g773)) + ((g1193) & (!g1194) & (!g1195) & (g1196) & (!g820) & (!g773)) + ((g1193) & (!g1194) & (!g1195) & (g1196) & (g820) & (g773)) + ((g1193) & (!g1194) & (g1195) & (!g1196) & (!g820) & (!g773)) + ((g1193) & (!g1194) & (g1195) & (!g1196) & (!g820) & (g773)) + ((g1193) & (!g1194) & (g1195) & (g1196) & (!g820) & (!g773)) + ((g1193) & (!g1194) & (g1195) & (g1196) & (!g820) & (g773)) + ((g1193) & (!g1194) & (g1195) & (g1196) & (g820) & (g773)) + ((g1193) & (g1194) & (!g1195) & (!g1196) & (!g820) & (!g773)) + ((g1193) & (g1194) & (!g1195) & (!g1196) & (g820) & (!g773)) + ((g1193) & (g1194) & (!g1195) & (g1196) & (!g820) & (!g773)) + ((g1193) & (g1194) & (!g1195) & (g1196) & (g820) & (!g773)) + ((g1193) & (g1194) & (!g1195) & (g1196) & (g820) & (g773)) + ((g1193) & (g1194) & (g1195) & (!g1196) & (!g820) & (!g773)) + ((g1193) & (g1194) & (g1195) & (!g1196) & (!g820) & (g773)) + ((g1193) & (g1194) & (g1195) & (!g1196) & (g820) & (!g773)) + ((g1193) & (g1194) & (g1195) & (g1196) & (!g820) & (!g773)) + ((g1193) & (g1194) & (g1195) & (g1196) & (!g820) & (g773)) + ((g1193) & (g1194) & (g1195) & (g1196) & (g820) & (!g773)) + ((g1193) & (g1194) & (g1195) & (g1196) & (g820) & (g773)));
	assign g1894 = (((!g1198) & (!g1199) & (!g1200) & (g1201) & (g820) & (g773)) + ((!g1198) & (!g1199) & (g1200) & (!g1201) & (!g820) & (g773)) + ((!g1198) & (!g1199) & (g1200) & (g1201) & (!g820) & (g773)) + ((!g1198) & (!g1199) & (g1200) & (g1201) & (g820) & (g773)) + ((!g1198) & (g1199) & (!g1200) & (!g1201) & (g820) & (!g773)) + ((!g1198) & (g1199) & (!g1200) & (g1201) & (g820) & (!g773)) + ((!g1198) & (g1199) & (!g1200) & (g1201) & (g820) & (g773)) + ((!g1198) & (g1199) & (g1200) & (!g1201) & (!g820) & (g773)) + ((!g1198) & (g1199) & (g1200) & (!g1201) & (g820) & (!g773)) + ((!g1198) & (g1199) & (g1200) & (g1201) & (!g820) & (g773)) + ((!g1198) & (g1199) & (g1200) & (g1201) & (g820) & (!g773)) + ((!g1198) & (g1199) & (g1200) & (g1201) & (g820) & (g773)) + ((g1198) & (!g1199) & (!g1200) & (!g1201) & (!g820) & (!g773)) + ((g1198) & (!g1199) & (!g1200) & (g1201) & (!g820) & (!g773)) + ((g1198) & (!g1199) & (!g1200) & (g1201) & (g820) & (g773)) + ((g1198) & (!g1199) & (g1200) & (!g1201) & (!g820) & (!g773)) + ((g1198) & (!g1199) & (g1200) & (!g1201) & (!g820) & (g773)) + ((g1198) & (!g1199) & (g1200) & (g1201) & (!g820) & (!g773)) + ((g1198) & (!g1199) & (g1200) & (g1201) & (!g820) & (g773)) + ((g1198) & (!g1199) & (g1200) & (g1201) & (g820) & (g773)) + ((g1198) & (g1199) & (!g1200) & (!g1201) & (!g820) & (!g773)) + ((g1198) & (g1199) & (!g1200) & (!g1201) & (g820) & (!g773)) + ((g1198) & (g1199) & (!g1200) & (g1201) & (!g820) & (!g773)) + ((g1198) & (g1199) & (!g1200) & (g1201) & (g820) & (!g773)) + ((g1198) & (g1199) & (!g1200) & (g1201) & (g820) & (g773)) + ((g1198) & (g1199) & (g1200) & (!g1201) & (!g820) & (!g773)) + ((g1198) & (g1199) & (g1200) & (!g1201) & (!g820) & (g773)) + ((g1198) & (g1199) & (g1200) & (!g1201) & (g820) & (!g773)) + ((g1198) & (g1199) & (g1200) & (g1201) & (!g820) & (!g773)) + ((g1198) & (g1199) & (g1200) & (g1201) & (!g820) & (g773)) + ((g1198) & (g1199) & (g1200) & (g1201) & (g820) & (!g773)) + ((g1198) & (g1199) & (g1200) & (g1201) & (g820) & (g773)));
	assign g1895 = (((!g1203) & (!g1204) & (!g1205) & (g1206) & (g820) & (g773)) + ((!g1203) & (!g1204) & (g1205) & (!g1206) & (!g820) & (g773)) + ((!g1203) & (!g1204) & (g1205) & (g1206) & (!g820) & (g773)) + ((!g1203) & (!g1204) & (g1205) & (g1206) & (g820) & (g773)) + ((!g1203) & (g1204) & (!g1205) & (!g1206) & (g820) & (!g773)) + ((!g1203) & (g1204) & (!g1205) & (g1206) & (g820) & (!g773)) + ((!g1203) & (g1204) & (!g1205) & (g1206) & (g820) & (g773)) + ((!g1203) & (g1204) & (g1205) & (!g1206) & (!g820) & (g773)) + ((!g1203) & (g1204) & (g1205) & (!g1206) & (g820) & (!g773)) + ((!g1203) & (g1204) & (g1205) & (g1206) & (!g820) & (g773)) + ((!g1203) & (g1204) & (g1205) & (g1206) & (g820) & (!g773)) + ((!g1203) & (g1204) & (g1205) & (g1206) & (g820) & (g773)) + ((g1203) & (!g1204) & (!g1205) & (!g1206) & (!g820) & (!g773)) + ((g1203) & (!g1204) & (!g1205) & (g1206) & (!g820) & (!g773)) + ((g1203) & (!g1204) & (!g1205) & (g1206) & (g820) & (g773)) + ((g1203) & (!g1204) & (g1205) & (!g1206) & (!g820) & (!g773)) + ((g1203) & (!g1204) & (g1205) & (!g1206) & (!g820) & (g773)) + ((g1203) & (!g1204) & (g1205) & (g1206) & (!g820) & (!g773)) + ((g1203) & (!g1204) & (g1205) & (g1206) & (!g820) & (g773)) + ((g1203) & (!g1204) & (g1205) & (g1206) & (g820) & (g773)) + ((g1203) & (g1204) & (!g1205) & (!g1206) & (!g820) & (!g773)) + ((g1203) & (g1204) & (!g1205) & (!g1206) & (g820) & (!g773)) + ((g1203) & (g1204) & (!g1205) & (g1206) & (!g820) & (!g773)) + ((g1203) & (g1204) & (!g1205) & (g1206) & (g820) & (!g773)) + ((g1203) & (g1204) & (!g1205) & (g1206) & (g820) & (g773)) + ((g1203) & (g1204) & (g1205) & (!g1206) & (!g820) & (!g773)) + ((g1203) & (g1204) & (g1205) & (!g1206) & (!g820) & (g773)) + ((g1203) & (g1204) & (g1205) & (!g1206) & (g820) & (!g773)) + ((g1203) & (g1204) & (g1205) & (g1206) & (!g820) & (!g773)) + ((g1203) & (g1204) & (g1205) & (g1206) & (!g820) & (g773)) + ((g1203) & (g1204) & (g1205) & (g1206) & (g820) & (!g773)) + ((g1203) & (g1204) & (g1205) & (g1206) & (g820) & (g773)));
	assign g1896 = (((!g1892) & (!g1893) & (!g1894) & (g1895) & (g677) & (g726)) + ((!g1892) & (!g1893) & (g1894) & (!g1895) & (!g677) & (g726)) + ((!g1892) & (!g1893) & (g1894) & (g1895) & (!g677) & (g726)) + ((!g1892) & (!g1893) & (g1894) & (g1895) & (g677) & (g726)) + ((!g1892) & (g1893) & (!g1894) & (!g1895) & (g677) & (!g726)) + ((!g1892) & (g1893) & (!g1894) & (g1895) & (g677) & (!g726)) + ((!g1892) & (g1893) & (!g1894) & (g1895) & (g677) & (g726)) + ((!g1892) & (g1893) & (g1894) & (!g1895) & (!g677) & (g726)) + ((!g1892) & (g1893) & (g1894) & (!g1895) & (g677) & (!g726)) + ((!g1892) & (g1893) & (g1894) & (g1895) & (!g677) & (g726)) + ((!g1892) & (g1893) & (g1894) & (g1895) & (g677) & (!g726)) + ((!g1892) & (g1893) & (g1894) & (g1895) & (g677) & (g726)) + ((g1892) & (!g1893) & (!g1894) & (!g1895) & (!g677) & (!g726)) + ((g1892) & (!g1893) & (!g1894) & (g1895) & (!g677) & (!g726)) + ((g1892) & (!g1893) & (!g1894) & (g1895) & (g677) & (g726)) + ((g1892) & (!g1893) & (g1894) & (!g1895) & (!g677) & (!g726)) + ((g1892) & (!g1893) & (g1894) & (!g1895) & (!g677) & (g726)) + ((g1892) & (!g1893) & (g1894) & (g1895) & (!g677) & (!g726)) + ((g1892) & (!g1893) & (g1894) & (g1895) & (!g677) & (g726)) + ((g1892) & (!g1893) & (g1894) & (g1895) & (g677) & (g726)) + ((g1892) & (g1893) & (!g1894) & (!g1895) & (!g677) & (!g726)) + ((g1892) & (g1893) & (!g1894) & (!g1895) & (g677) & (!g726)) + ((g1892) & (g1893) & (!g1894) & (g1895) & (!g677) & (!g726)) + ((g1892) & (g1893) & (!g1894) & (g1895) & (g677) & (!g726)) + ((g1892) & (g1893) & (!g1894) & (g1895) & (g677) & (g726)) + ((g1892) & (g1893) & (g1894) & (!g1895) & (!g677) & (!g726)) + ((g1892) & (g1893) & (g1894) & (!g1895) & (!g677) & (g726)) + ((g1892) & (g1893) & (g1894) & (!g1895) & (g677) & (!g726)) + ((g1892) & (g1893) & (g1894) & (g1895) & (!g677) & (!g726)) + ((g1892) & (g1893) & (g1894) & (g1895) & (!g677) & (g726)) + ((g1892) & (g1893) & (g1894) & (g1895) & (g677) & (!g726)) + ((g1892) & (g1893) & (g1894) & (g1895) & (g677) & (g726)));
	assign g1897 = (((!g1209) & (!g1210) & (!g1211) & (g1212) & (g677) & (g726)) + ((!g1209) & (!g1210) & (g1211) & (!g1212) & (!g677) & (g726)) + ((!g1209) & (!g1210) & (g1211) & (g1212) & (!g677) & (g726)) + ((!g1209) & (!g1210) & (g1211) & (g1212) & (g677) & (g726)) + ((!g1209) & (g1210) & (!g1211) & (!g1212) & (g677) & (!g726)) + ((!g1209) & (g1210) & (!g1211) & (g1212) & (g677) & (!g726)) + ((!g1209) & (g1210) & (!g1211) & (g1212) & (g677) & (g726)) + ((!g1209) & (g1210) & (g1211) & (!g1212) & (!g677) & (g726)) + ((!g1209) & (g1210) & (g1211) & (!g1212) & (g677) & (!g726)) + ((!g1209) & (g1210) & (g1211) & (g1212) & (!g677) & (g726)) + ((!g1209) & (g1210) & (g1211) & (g1212) & (g677) & (!g726)) + ((!g1209) & (g1210) & (g1211) & (g1212) & (g677) & (g726)) + ((g1209) & (!g1210) & (!g1211) & (!g1212) & (!g677) & (!g726)) + ((g1209) & (!g1210) & (!g1211) & (g1212) & (!g677) & (!g726)) + ((g1209) & (!g1210) & (!g1211) & (g1212) & (g677) & (g726)) + ((g1209) & (!g1210) & (g1211) & (!g1212) & (!g677) & (!g726)) + ((g1209) & (!g1210) & (g1211) & (!g1212) & (!g677) & (g726)) + ((g1209) & (!g1210) & (g1211) & (g1212) & (!g677) & (!g726)) + ((g1209) & (!g1210) & (g1211) & (g1212) & (!g677) & (g726)) + ((g1209) & (!g1210) & (g1211) & (g1212) & (g677) & (g726)) + ((g1209) & (g1210) & (!g1211) & (!g1212) & (!g677) & (!g726)) + ((g1209) & (g1210) & (!g1211) & (!g1212) & (g677) & (!g726)) + ((g1209) & (g1210) & (!g1211) & (g1212) & (!g677) & (!g726)) + ((g1209) & (g1210) & (!g1211) & (g1212) & (g677) & (!g726)) + ((g1209) & (g1210) & (!g1211) & (g1212) & (g677) & (g726)) + ((g1209) & (g1210) & (g1211) & (!g1212) & (!g677) & (!g726)) + ((g1209) & (g1210) & (g1211) & (!g1212) & (!g677) & (g726)) + ((g1209) & (g1210) & (g1211) & (!g1212) & (g677) & (!g726)) + ((g1209) & (g1210) & (g1211) & (g1212) & (!g677) & (!g726)) + ((g1209) & (g1210) & (g1211) & (g1212) & (!g677) & (g726)) + ((g1209) & (g1210) & (g1211) & (g1212) & (g677) & (!g726)) + ((g1209) & (g1210) & (g1211) & (g1212) & (g677) & (g726)));
	assign g1898 = (((!g677) & (!sk[44]) & (!g726) & (!g1214) & (g1215) & (!g1216)) + ((!g677) & (!sk[44]) & (!g726) & (!g1214) & (g1215) & (g1216)) + ((!g677) & (!sk[44]) & (!g726) & (g1214) & (!g1215) & (!g1216)) + ((!g677) & (!sk[44]) & (!g726) & (g1214) & (!g1215) & (g1216)) + ((!g677) & (!sk[44]) & (!g726) & (g1214) & (g1215) & (!g1216)) + ((!g677) & (!sk[44]) & (!g726) & (g1214) & (g1215) & (g1216)) + ((!g677) & (!sk[44]) & (g726) & (!g1214) & (!g1215) & (!g1216)) + ((!g677) & (!sk[44]) & (g726) & (!g1214) & (!g1215) & (g1216)) + ((!g677) & (!sk[44]) & (g726) & (!g1214) & (g1215) & (!g1216)) + ((!g677) & (!sk[44]) & (g726) & (!g1214) & (g1215) & (g1216)) + ((!g677) & (!sk[44]) & (g726) & (g1214) & (!g1215) & (!g1216)) + ((!g677) & (!sk[44]) & (g726) & (g1214) & (!g1215) & (g1216)) + ((!g677) & (!sk[44]) & (g726) & (g1214) & (g1215) & (!g1216)) + ((!g677) & (!sk[44]) & (g726) & (g1214) & (g1215) & (g1216)) + ((!g677) & (sk[44]) & (g726) & (!g1214) & (!g1215) & (g1216)) + ((!g677) & (sk[44]) & (g726) & (!g1214) & (g1215) & (g1216)) + ((!g677) & (sk[44]) & (g726) & (g1214) & (!g1215) & (g1216)) + ((!g677) & (sk[44]) & (g726) & (g1214) & (g1215) & (g1216)) + ((g677) & (!sk[44]) & (!g726) & (!g1214) & (g1215) & (!g1216)) + ((g677) & (!sk[44]) & (!g726) & (!g1214) & (g1215) & (g1216)) + ((g677) & (!sk[44]) & (!g726) & (g1214) & (!g1215) & (!g1216)) + ((g677) & (!sk[44]) & (!g726) & (g1214) & (!g1215) & (g1216)) + ((g677) & (!sk[44]) & (!g726) & (g1214) & (g1215) & (!g1216)) + ((g677) & (!sk[44]) & (!g726) & (g1214) & (g1215) & (g1216)) + ((g677) & (!sk[44]) & (g726) & (!g1214) & (!g1215) & (!g1216)) + ((g677) & (!sk[44]) & (g726) & (!g1214) & (!g1215) & (g1216)) + ((g677) & (!sk[44]) & (g726) & (!g1214) & (g1215) & (!g1216)) + ((g677) & (!sk[44]) & (g726) & (!g1214) & (g1215) & (g1216)) + ((g677) & (!sk[44]) & (g726) & (g1214) & (!g1215) & (!g1216)) + ((g677) & (!sk[44]) & (g726) & (g1214) & (!g1215) & (g1216)) + ((g677) & (!sk[44]) & (g726) & (g1214) & (g1215) & (!g1216)) + ((g677) & (!sk[44]) & (g726) & (g1214) & (g1215) & (g1216)) + ((g677) & (sk[44]) & (!g726) & (g1214) & (!g1215) & (!g1216)) + ((g677) & (sk[44]) & (!g726) & (g1214) & (!g1215) & (g1216)) + ((g677) & (sk[44]) & (!g726) & (g1214) & (g1215) & (!g1216)) + ((g677) & (sk[44]) & (!g726) & (g1214) & (g1215) & (g1216)) + ((g677) & (sk[44]) & (g726) & (!g1214) & (g1215) & (!g1216)) + ((g677) & (sk[44]) & (g726) & (!g1214) & (g1215) & (g1216)) + ((g677) & (sk[44]) & (g726) & (g1214) & (g1215) & (!g1216)) + ((g677) & (sk[44]) & (g726) & (g1214) & (g1215) & (g1216)));
	assign g1899 = (((!g1218) & (!g1219) & (!g1220) & (g1221) & (g677) & (g726)) + ((!g1218) & (!g1219) & (g1220) & (!g1221) & (!g677) & (g726)) + ((!g1218) & (!g1219) & (g1220) & (g1221) & (!g677) & (g726)) + ((!g1218) & (!g1219) & (g1220) & (g1221) & (g677) & (g726)) + ((!g1218) & (g1219) & (!g1220) & (!g1221) & (g677) & (!g726)) + ((!g1218) & (g1219) & (!g1220) & (g1221) & (g677) & (!g726)) + ((!g1218) & (g1219) & (!g1220) & (g1221) & (g677) & (g726)) + ((!g1218) & (g1219) & (g1220) & (!g1221) & (!g677) & (g726)) + ((!g1218) & (g1219) & (g1220) & (!g1221) & (g677) & (!g726)) + ((!g1218) & (g1219) & (g1220) & (g1221) & (!g677) & (g726)) + ((!g1218) & (g1219) & (g1220) & (g1221) & (g677) & (!g726)) + ((!g1218) & (g1219) & (g1220) & (g1221) & (g677) & (g726)) + ((g1218) & (!g1219) & (!g1220) & (!g1221) & (!g677) & (!g726)) + ((g1218) & (!g1219) & (!g1220) & (g1221) & (!g677) & (!g726)) + ((g1218) & (!g1219) & (!g1220) & (g1221) & (g677) & (g726)) + ((g1218) & (!g1219) & (g1220) & (!g1221) & (!g677) & (!g726)) + ((g1218) & (!g1219) & (g1220) & (!g1221) & (!g677) & (g726)) + ((g1218) & (!g1219) & (g1220) & (g1221) & (!g677) & (!g726)) + ((g1218) & (!g1219) & (g1220) & (g1221) & (!g677) & (g726)) + ((g1218) & (!g1219) & (g1220) & (g1221) & (g677) & (g726)) + ((g1218) & (g1219) & (!g1220) & (!g1221) & (!g677) & (!g726)) + ((g1218) & (g1219) & (!g1220) & (!g1221) & (g677) & (!g726)) + ((g1218) & (g1219) & (!g1220) & (g1221) & (!g677) & (!g726)) + ((g1218) & (g1219) & (!g1220) & (g1221) & (g677) & (!g726)) + ((g1218) & (g1219) & (!g1220) & (g1221) & (g677) & (g726)) + ((g1218) & (g1219) & (g1220) & (!g1221) & (!g677) & (!g726)) + ((g1218) & (g1219) & (g1220) & (!g1221) & (!g677) & (g726)) + ((g1218) & (g1219) & (g1220) & (!g1221) & (g677) & (!g726)) + ((g1218) & (g1219) & (g1220) & (g1221) & (!g677) & (!g726)) + ((g1218) & (g1219) & (g1220) & (g1221) & (!g677) & (g726)) + ((g1218) & (g1219) & (g1220) & (g1221) & (g677) & (!g726)) + ((g1218) & (g1219) & (g1220) & (g1221) & (g677) & (g726)));
	assign g1900 = (((!g1223) & (!g1224) & (!g1225) & (g1226) & (g677) & (g726)) + ((!g1223) & (!g1224) & (g1225) & (!g1226) & (!g677) & (g726)) + ((!g1223) & (!g1224) & (g1225) & (g1226) & (!g677) & (g726)) + ((!g1223) & (!g1224) & (g1225) & (g1226) & (g677) & (g726)) + ((!g1223) & (g1224) & (!g1225) & (!g1226) & (g677) & (!g726)) + ((!g1223) & (g1224) & (!g1225) & (g1226) & (g677) & (!g726)) + ((!g1223) & (g1224) & (!g1225) & (g1226) & (g677) & (g726)) + ((!g1223) & (g1224) & (g1225) & (!g1226) & (!g677) & (g726)) + ((!g1223) & (g1224) & (g1225) & (!g1226) & (g677) & (!g726)) + ((!g1223) & (g1224) & (g1225) & (g1226) & (!g677) & (g726)) + ((!g1223) & (g1224) & (g1225) & (g1226) & (g677) & (!g726)) + ((!g1223) & (g1224) & (g1225) & (g1226) & (g677) & (g726)) + ((g1223) & (!g1224) & (!g1225) & (!g1226) & (!g677) & (!g726)) + ((g1223) & (!g1224) & (!g1225) & (g1226) & (!g677) & (!g726)) + ((g1223) & (!g1224) & (!g1225) & (g1226) & (g677) & (g726)) + ((g1223) & (!g1224) & (g1225) & (!g1226) & (!g677) & (!g726)) + ((g1223) & (!g1224) & (g1225) & (!g1226) & (!g677) & (g726)) + ((g1223) & (!g1224) & (g1225) & (g1226) & (!g677) & (!g726)) + ((g1223) & (!g1224) & (g1225) & (g1226) & (!g677) & (g726)) + ((g1223) & (!g1224) & (g1225) & (g1226) & (g677) & (g726)) + ((g1223) & (g1224) & (!g1225) & (!g1226) & (!g677) & (!g726)) + ((g1223) & (g1224) & (!g1225) & (!g1226) & (g677) & (!g726)) + ((g1223) & (g1224) & (!g1225) & (g1226) & (!g677) & (!g726)) + ((g1223) & (g1224) & (!g1225) & (g1226) & (g677) & (!g726)) + ((g1223) & (g1224) & (!g1225) & (g1226) & (g677) & (g726)) + ((g1223) & (g1224) & (g1225) & (!g1226) & (!g677) & (!g726)) + ((g1223) & (g1224) & (g1225) & (!g1226) & (!g677) & (g726)) + ((g1223) & (g1224) & (g1225) & (!g1226) & (g677) & (!g726)) + ((g1223) & (g1224) & (g1225) & (g1226) & (!g677) & (!g726)) + ((g1223) & (g1224) & (g1225) & (g1226) & (!g677) & (g726)) + ((g1223) & (g1224) & (g1225) & (g1226) & (g677) & (!g726)) + ((g1223) & (g1224) & (g1225) & (g1226) & (g677) & (g726)));
	assign g1901 = (((!g820) & (!g773) & (!g1897) & (g1898) & (!g1899) & (!g1900)) + ((!g820) & (!g773) & (!g1897) & (g1898) & (!g1899) & (g1900)) + ((!g820) & (!g773) & (!g1897) & (g1898) & (g1899) & (!g1900)) + ((!g820) & (!g773) & (!g1897) & (g1898) & (g1899) & (g1900)) + ((!g820) & (!g773) & (g1897) & (g1898) & (!g1899) & (!g1900)) + ((!g820) & (!g773) & (g1897) & (g1898) & (!g1899) & (g1900)) + ((!g820) & (!g773) & (g1897) & (g1898) & (g1899) & (!g1900)) + ((!g820) & (!g773) & (g1897) & (g1898) & (g1899) & (g1900)) + ((!g820) & (g773) & (!g1897) & (!g1898) & (!g1899) & (g1900)) + ((!g820) & (g773) & (!g1897) & (!g1898) & (g1899) & (g1900)) + ((!g820) & (g773) & (!g1897) & (g1898) & (!g1899) & (g1900)) + ((!g820) & (g773) & (!g1897) & (g1898) & (g1899) & (g1900)) + ((!g820) & (g773) & (g1897) & (!g1898) & (!g1899) & (g1900)) + ((!g820) & (g773) & (g1897) & (!g1898) & (g1899) & (g1900)) + ((!g820) & (g773) & (g1897) & (g1898) & (!g1899) & (g1900)) + ((!g820) & (g773) & (g1897) & (g1898) & (g1899) & (g1900)) + ((g820) & (!g773) & (g1897) & (!g1898) & (!g1899) & (!g1900)) + ((g820) & (!g773) & (g1897) & (!g1898) & (!g1899) & (g1900)) + ((g820) & (!g773) & (g1897) & (!g1898) & (g1899) & (!g1900)) + ((g820) & (!g773) & (g1897) & (!g1898) & (g1899) & (g1900)) + ((g820) & (!g773) & (g1897) & (g1898) & (!g1899) & (!g1900)) + ((g820) & (!g773) & (g1897) & (g1898) & (!g1899) & (g1900)) + ((g820) & (!g773) & (g1897) & (g1898) & (g1899) & (!g1900)) + ((g820) & (!g773) & (g1897) & (g1898) & (g1899) & (g1900)) + ((g820) & (g773) & (!g1897) & (!g1898) & (g1899) & (!g1900)) + ((g820) & (g773) & (!g1897) & (!g1898) & (g1899) & (g1900)) + ((g820) & (g773) & (!g1897) & (g1898) & (g1899) & (!g1900)) + ((g820) & (g773) & (!g1897) & (g1898) & (g1899) & (g1900)) + ((g820) & (g773) & (g1897) & (!g1898) & (g1899) & (!g1900)) + ((g820) & (g773) & (g1897) & (!g1898) & (g1899) & (g1900)) + ((g820) & (g773) & (g1897) & (g1898) & (g1899) & (!g1900)) + ((g820) & (g773) & (g1897) & (g1898) & (g1899) & (g1900)));
	assign g1902 = (((!g867) & (!g1896) & (!sk[48]) & (g1901)) + ((!g867) & (!g1896) & (sk[48]) & (g1901)) + ((!g867) & (g1896) & (!sk[48]) & (!g1901)) + ((!g867) & (g1896) & (!sk[48]) & (g1901)) + ((!g867) & (g1896) & (sk[48]) & (g1901)) + ((g867) & (!g1896) & (!sk[48]) & (g1901)) + ((g867) & (g1896) & (!sk[48]) & (!g1901)) + ((g867) & (g1896) & (!sk[48]) & (g1901)) + ((g867) & (g1896) & (sk[48]) & (!g1901)) + ((g867) & (g1896) & (sk[48]) & (g1901)));
	assign g1903 = (((!g1592) & (!sk[49]) & (!g1593) & (!g1605) & (g1692) & (!g58)) + ((!g1592) & (!sk[49]) & (!g1593) & (!g1605) & (g1692) & (g58)) + ((!g1592) & (!sk[49]) & (!g1593) & (g1605) & (!g1692) & (!g58)) + ((!g1592) & (!sk[49]) & (!g1593) & (g1605) & (!g1692) & (g58)) + ((!g1592) & (!sk[49]) & (!g1593) & (g1605) & (g1692) & (!g58)) + ((!g1592) & (!sk[49]) & (!g1593) & (g1605) & (g1692) & (g58)) + ((!g1592) & (!sk[49]) & (g1593) & (!g1605) & (!g1692) & (!g58)) + ((!g1592) & (!sk[49]) & (g1593) & (!g1605) & (!g1692) & (g58)) + ((!g1592) & (!sk[49]) & (g1593) & (!g1605) & (g1692) & (!g58)) + ((!g1592) & (!sk[49]) & (g1593) & (!g1605) & (g1692) & (g58)) + ((!g1592) & (!sk[49]) & (g1593) & (g1605) & (!g1692) & (!g58)) + ((!g1592) & (!sk[49]) & (g1593) & (g1605) & (!g1692) & (g58)) + ((!g1592) & (!sk[49]) & (g1593) & (g1605) & (g1692) & (!g58)) + ((!g1592) & (!sk[49]) & (g1593) & (g1605) & (g1692) & (g58)) + ((!g1592) & (sk[49]) & (!g1593) & (!g1605) & (g1692) & (!g58)) + ((!g1592) & (sk[49]) & (!g1593) & (!g1605) & (g1692) & (g58)) + ((!g1592) & (sk[49]) & (!g1593) & (g1605) & (g1692) & (!g58)) + ((!g1592) & (sk[49]) & (!g1593) & (g1605) & (g1692) & (g58)) + ((!g1592) & (sk[49]) & (g1593) & (!g1605) & (g1692) & (!g58)) + ((!g1592) & (sk[49]) & (g1593) & (!g1605) & (g1692) & (g58)) + ((!g1592) & (sk[49]) & (g1593) & (g1605) & (g1692) & (!g58)) + ((!g1592) & (sk[49]) & (g1593) & (g1605) & (g1692) & (g58)) + ((g1592) & (!sk[49]) & (!g1593) & (!g1605) & (g1692) & (!g58)) + ((g1592) & (!sk[49]) & (!g1593) & (!g1605) & (g1692) & (g58)) + ((g1592) & (!sk[49]) & (!g1593) & (g1605) & (!g1692) & (!g58)) + ((g1592) & (!sk[49]) & (!g1593) & (g1605) & (!g1692) & (g58)) + ((g1592) & (!sk[49]) & (!g1593) & (g1605) & (g1692) & (!g58)) + ((g1592) & (!sk[49]) & (!g1593) & (g1605) & (g1692) & (g58)) + ((g1592) & (!sk[49]) & (g1593) & (!g1605) & (!g1692) & (!g58)) + ((g1592) & (!sk[49]) & (g1593) & (!g1605) & (!g1692) & (g58)) + ((g1592) & (!sk[49]) & (g1593) & (!g1605) & (g1692) & (!g58)) + ((g1592) & (!sk[49]) & (g1593) & (!g1605) & (g1692) & (g58)) + ((g1592) & (!sk[49]) & (g1593) & (g1605) & (!g1692) & (!g58)) + ((g1592) & (!sk[49]) & (g1593) & (g1605) & (!g1692) & (g58)) + ((g1592) & (!sk[49]) & (g1593) & (g1605) & (g1692) & (!g58)) + ((g1592) & (!sk[49]) & (g1593) & (g1605) & (g1692) & (g58)) + ((g1592) & (sk[49]) & (!g1593) & (!g1605) & (g1692) & (!g58)) + ((g1592) & (sk[49]) & (!g1593) & (!g1605) & (g1692) & (g58)) + ((g1592) & (sk[49]) & (g1593) & (!g1605) & (!g1692) & (g58)) + ((g1592) & (sk[49]) & (g1593) & (!g1605) & (g1692) & (g58)) + ((g1592) & (sk[49]) & (g1593) & (g1605) & (!g1692) & (g58)) + ((g1592) & (sk[49]) & (g1593) & (g1605) & (g1692) & (g58)));
	assign g1904 = (((!g132) & (!g1812) & (!sk[50]) & (!g1902) & (g1903)) + ((!g132) & (!g1812) & (!sk[50]) & (g1902) & (!g1903)) + ((!g132) & (!g1812) & (!sk[50]) & (g1902) & (g1903)) + ((!g132) & (g1812) & (!sk[50]) & (!g1902) & (!g1903)) + ((!g132) & (g1812) & (!sk[50]) & (!g1902) & (g1903)) + ((!g132) & (g1812) & (!sk[50]) & (g1902) & (!g1903)) + ((!g132) & (g1812) & (!sk[50]) & (g1902) & (g1903)) + ((!g132) & (g1812) & (sk[50]) & (!g1902) & (g1903)) + ((!g132) & (g1812) & (sk[50]) & (g1902) & (g1903)) + ((g132) & (!g1812) & (!sk[50]) & (!g1902) & (g1903)) + ((g132) & (!g1812) & (!sk[50]) & (g1902) & (!g1903)) + ((g132) & (!g1812) & (!sk[50]) & (g1902) & (g1903)) + ((g132) & (g1812) & (!sk[50]) & (!g1902) & (!g1903)) + ((g132) & (g1812) & (!sk[50]) & (!g1902) & (g1903)) + ((g132) & (g1812) & (!sk[50]) & (g1902) & (!g1903)) + ((g132) & (g1812) & (!sk[50]) & (g1902) & (g1903)) + ((g132) & (g1812) & (sk[50]) & (g1902) & (!g1903)) + ((g132) & (g1812) & (sk[50]) & (g1902) & (g1903)));
	assign g1905 = (((!g1233) & (!g1238) & (!g1243) & (g1248) & (g677) & (g726)) + ((!g1233) & (!g1238) & (g1243) & (!g1248) & (!g677) & (g726)) + ((!g1233) & (!g1238) & (g1243) & (g1248) & (!g677) & (g726)) + ((!g1233) & (!g1238) & (g1243) & (g1248) & (g677) & (g726)) + ((!g1233) & (g1238) & (!g1243) & (!g1248) & (g677) & (!g726)) + ((!g1233) & (g1238) & (!g1243) & (g1248) & (g677) & (!g726)) + ((!g1233) & (g1238) & (!g1243) & (g1248) & (g677) & (g726)) + ((!g1233) & (g1238) & (g1243) & (!g1248) & (!g677) & (g726)) + ((!g1233) & (g1238) & (g1243) & (!g1248) & (g677) & (!g726)) + ((!g1233) & (g1238) & (g1243) & (g1248) & (!g677) & (g726)) + ((!g1233) & (g1238) & (g1243) & (g1248) & (g677) & (!g726)) + ((!g1233) & (g1238) & (g1243) & (g1248) & (g677) & (g726)) + ((g1233) & (!g1238) & (!g1243) & (!g1248) & (!g677) & (!g726)) + ((g1233) & (!g1238) & (!g1243) & (g1248) & (!g677) & (!g726)) + ((g1233) & (!g1238) & (!g1243) & (g1248) & (g677) & (g726)) + ((g1233) & (!g1238) & (g1243) & (!g1248) & (!g677) & (!g726)) + ((g1233) & (!g1238) & (g1243) & (!g1248) & (!g677) & (g726)) + ((g1233) & (!g1238) & (g1243) & (g1248) & (!g677) & (!g726)) + ((g1233) & (!g1238) & (g1243) & (g1248) & (!g677) & (g726)) + ((g1233) & (!g1238) & (g1243) & (g1248) & (g677) & (g726)) + ((g1233) & (g1238) & (!g1243) & (!g1248) & (!g677) & (!g726)) + ((g1233) & (g1238) & (!g1243) & (!g1248) & (g677) & (!g726)) + ((g1233) & (g1238) & (!g1243) & (g1248) & (!g677) & (!g726)) + ((g1233) & (g1238) & (!g1243) & (g1248) & (g677) & (!g726)) + ((g1233) & (g1238) & (!g1243) & (g1248) & (g677) & (g726)) + ((g1233) & (g1238) & (g1243) & (!g1248) & (!g677) & (!g726)) + ((g1233) & (g1238) & (g1243) & (!g1248) & (!g677) & (g726)) + ((g1233) & (g1238) & (g1243) & (!g1248) & (g677) & (!g726)) + ((g1233) & (g1238) & (g1243) & (g1248) & (!g677) & (!g726)) + ((g1233) & (g1238) & (g1243) & (g1248) & (!g677) & (g726)) + ((g1233) & (g1238) & (g1243) & (g1248) & (g677) & (!g726)) + ((g1233) & (g1238) & (g1243) & (g1248) & (g677) & (g726)));
	assign g1906 = (((!g1234) & (!g1239) & (!g1244) & (g1249) & (g677) & (g726)) + ((!g1234) & (!g1239) & (g1244) & (!g1249) & (!g677) & (g726)) + ((!g1234) & (!g1239) & (g1244) & (g1249) & (!g677) & (g726)) + ((!g1234) & (!g1239) & (g1244) & (g1249) & (g677) & (g726)) + ((!g1234) & (g1239) & (!g1244) & (!g1249) & (g677) & (!g726)) + ((!g1234) & (g1239) & (!g1244) & (g1249) & (g677) & (!g726)) + ((!g1234) & (g1239) & (!g1244) & (g1249) & (g677) & (g726)) + ((!g1234) & (g1239) & (g1244) & (!g1249) & (!g677) & (g726)) + ((!g1234) & (g1239) & (g1244) & (!g1249) & (g677) & (!g726)) + ((!g1234) & (g1239) & (g1244) & (g1249) & (!g677) & (g726)) + ((!g1234) & (g1239) & (g1244) & (g1249) & (g677) & (!g726)) + ((!g1234) & (g1239) & (g1244) & (g1249) & (g677) & (g726)) + ((g1234) & (!g1239) & (!g1244) & (!g1249) & (!g677) & (!g726)) + ((g1234) & (!g1239) & (!g1244) & (g1249) & (!g677) & (!g726)) + ((g1234) & (!g1239) & (!g1244) & (g1249) & (g677) & (g726)) + ((g1234) & (!g1239) & (g1244) & (!g1249) & (!g677) & (!g726)) + ((g1234) & (!g1239) & (g1244) & (!g1249) & (!g677) & (g726)) + ((g1234) & (!g1239) & (g1244) & (g1249) & (!g677) & (!g726)) + ((g1234) & (!g1239) & (g1244) & (g1249) & (!g677) & (g726)) + ((g1234) & (!g1239) & (g1244) & (g1249) & (g677) & (g726)) + ((g1234) & (g1239) & (!g1244) & (!g1249) & (!g677) & (!g726)) + ((g1234) & (g1239) & (!g1244) & (!g1249) & (g677) & (!g726)) + ((g1234) & (g1239) & (!g1244) & (g1249) & (!g677) & (!g726)) + ((g1234) & (g1239) & (!g1244) & (g1249) & (g677) & (!g726)) + ((g1234) & (g1239) & (!g1244) & (g1249) & (g677) & (g726)) + ((g1234) & (g1239) & (g1244) & (!g1249) & (!g677) & (!g726)) + ((g1234) & (g1239) & (g1244) & (!g1249) & (!g677) & (g726)) + ((g1234) & (g1239) & (g1244) & (!g1249) & (g677) & (!g726)) + ((g1234) & (g1239) & (g1244) & (g1249) & (!g677) & (!g726)) + ((g1234) & (g1239) & (g1244) & (g1249) & (!g677) & (g726)) + ((g1234) & (g1239) & (g1244) & (g1249) & (g677) & (!g726)) + ((g1234) & (g1239) & (g1244) & (g1249) & (g677) & (g726)));
	assign g1907 = (((!g1235) & (!g1240) & (!g1245) & (g1250) & (g677) & (g726)) + ((!g1235) & (!g1240) & (g1245) & (!g1250) & (!g677) & (g726)) + ((!g1235) & (!g1240) & (g1245) & (g1250) & (!g677) & (g726)) + ((!g1235) & (!g1240) & (g1245) & (g1250) & (g677) & (g726)) + ((!g1235) & (g1240) & (!g1245) & (!g1250) & (g677) & (!g726)) + ((!g1235) & (g1240) & (!g1245) & (g1250) & (g677) & (!g726)) + ((!g1235) & (g1240) & (!g1245) & (g1250) & (g677) & (g726)) + ((!g1235) & (g1240) & (g1245) & (!g1250) & (!g677) & (g726)) + ((!g1235) & (g1240) & (g1245) & (!g1250) & (g677) & (!g726)) + ((!g1235) & (g1240) & (g1245) & (g1250) & (!g677) & (g726)) + ((!g1235) & (g1240) & (g1245) & (g1250) & (g677) & (!g726)) + ((!g1235) & (g1240) & (g1245) & (g1250) & (g677) & (g726)) + ((g1235) & (!g1240) & (!g1245) & (!g1250) & (!g677) & (!g726)) + ((g1235) & (!g1240) & (!g1245) & (g1250) & (!g677) & (!g726)) + ((g1235) & (!g1240) & (!g1245) & (g1250) & (g677) & (g726)) + ((g1235) & (!g1240) & (g1245) & (!g1250) & (!g677) & (!g726)) + ((g1235) & (!g1240) & (g1245) & (!g1250) & (!g677) & (g726)) + ((g1235) & (!g1240) & (g1245) & (g1250) & (!g677) & (!g726)) + ((g1235) & (!g1240) & (g1245) & (g1250) & (!g677) & (g726)) + ((g1235) & (!g1240) & (g1245) & (g1250) & (g677) & (g726)) + ((g1235) & (g1240) & (!g1245) & (!g1250) & (!g677) & (!g726)) + ((g1235) & (g1240) & (!g1245) & (!g1250) & (g677) & (!g726)) + ((g1235) & (g1240) & (!g1245) & (g1250) & (!g677) & (!g726)) + ((g1235) & (g1240) & (!g1245) & (g1250) & (g677) & (!g726)) + ((g1235) & (g1240) & (!g1245) & (g1250) & (g677) & (g726)) + ((g1235) & (g1240) & (g1245) & (!g1250) & (!g677) & (!g726)) + ((g1235) & (g1240) & (g1245) & (!g1250) & (!g677) & (g726)) + ((g1235) & (g1240) & (g1245) & (!g1250) & (g677) & (!g726)) + ((g1235) & (g1240) & (g1245) & (g1250) & (!g677) & (!g726)) + ((g1235) & (g1240) & (g1245) & (g1250) & (!g677) & (g726)) + ((g1235) & (g1240) & (g1245) & (g1250) & (g677) & (!g726)) + ((g1235) & (g1240) & (g1245) & (g1250) & (g677) & (g726)));
	assign g1908 = (((!g1236) & (!g1241) & (!g1246) & (g1251) & (g677) & (g726)) + ((!g1236) & (!g1241) & (g1246) & (!g1251) & (!g677) & (g726)) + ((!g1236) & (!g1241) & (g1246) & (g1251) & (!g677) & (g726)) + ((!g1236) & (!g1241) & (g1246) & (g1251) & (g677) & (g726)) + ((!g1236) & (g1241) & (!g1246) & (!g1251) & (g677) & (!g726)) + ((!g1236) & (g1241) & (!g1246) & (g1251) & (g677) & (!g726)) + ((!g1236) & (g1241) & (!g1246) & (g1251) & (g677) & (g726)) + ((!g1236) & (g1241) & (g1246) & (!g1251) & (!g677) & (g726)) + ((!g1236) & (g1241) & (g1246) & (!g1251) & (g677) & (!g726)) + ((!g1236) & (g1241) & (g1246) & (g1251) & (!g677) & (g726)) + ((!g1236) & (g1241) & (g1246) & (g1251) & (g677) & (!g726)) + ((!g1236) & (g1241) & (g1246) & (g1251) & (g677) & (g726)) + ((g1236) & (!g1241) & (!g1246) & (!g1251) & (!g677) & (!g726)) + ((g1236) & (!g1241) & (!g1246) & (g1251) & (!g677) & (!g726)) + ((g1236) & (!g1241) & (!g1246) & (g1251) & (g677) & (g726)) + ((g1236) & (!g1241) & (g1246) & (!g1251) & (!g677) & (!g726)) + ((g1236) & (!g1241) & (g1246) & (!g1251) & (!g677) & (g726)) + ((g1236) & (!g1241) & (g1246) & (g1251) & (!g677) & (!g726)) + ((g1236) & (!g1241) & (g1246) & (g1251) & (!g677) & (g726)) + ((g1236) & (!g1241) & (g1246) & (g1251) & (g677) & (g726)) + ((g1236) & (g1241) & (!g1246) & (!g1251) & (!g677) & (!g726)) + ((g1236) & (g1241) & (!g1246) & (!g1251) & (g677) & (!g726)) + ((g1236) & (g1241) & (!g1246) & (g1251) & (!g677) & (!g726)) + ((g1236) & (g1241) & (!g1246) & (g1251) & (g677) & (!g726)) + ((g1236) & (g1241) & (!g1246) & (g1251) & (g677) & (g726)) + ((g1236) & (g1241) & (g1246) & (!g1251) & (!g677) & (!g726)) + ((g1236) & (g1241) & (g1246) & (!g1251) & (!g677) & (g726)) + ((g1236) & (g1241) & (g1246) & (!g1251) & (g677) & (!g726)) + ((g1236) & (g1241) & (g1246) & (g1251) & (!g677) & (!g726)) + ((g1236) & (g1241) & (g1246) & (g1251) & (!g677) & (g726)) + ((g1236) & (g1241) & (g1246) & (g1251) & (g677) & (!g726)) + ((g1236) & (g1241) & (g1246) & (g1251) & (g677) & (g726)));
	assign g1909 = (((!g1905) & (!g1906) & (!g1907) & (g1908) & (g820) & (g773)) + ((!g1905) & (!g1906) & (g1907) & (!g1908) & (!g820) & (g773)) + ((!g1905) & (!g1906) & (g1907) & (g1908) & (!g820) & (g773)) + ((!g1905) & (!g1906) & (g1907) & (g1908) & (g820) & (g773)) + ((!g1905) & (g1906) & (!g1907) & (!g1908) & (g820) & (!g773)) + ((!g1905) & (g1906) & (!g1907) & (g1908) & (g820) & (!g773)) + ((!g1905) & (g1906) & (!g1907) & (g1908) & (g820) & (g773)) + ((!g1905) & (g1906) & (g1907) & (!g1908) & (!g820) & (g773)) + ((!g1905) & (g1906) & (g1907) & (!g1908) & (g820) & (!g773)) + ((!g1905) & (g1906) & (g1907) & (g1908) & (!g820) & (g773)) + ((!g1905) & (g1906) & (g1907) & (g1908) & (g820) & (!g773)) + ((!g1905) & (g1906) & (g1907) & (g1908) & (g820) & (g773)) + ((g1905) & (!g1906) & (!g1907) & (!g1908) & (!g820) & (!g773)) + ((g1905) & (!g1906) & (!g1907) & (g1908) & (!g820) & (!g773)) + ((g1905) & (!g1906) & (!g1907) & (g1908) & (g820) & (g773)) + ((g1905) & (!g1906) & (g1907) & (!g1908) & (!g820) & (!g773)) + ((g1905) & (!g1906) & (g1907) & (!g1908) & (!g820) & (g773)) + ((g1905) & (!g1906) & (g1907) & (g1908) & (!g820) & (!g773)) + ((g1905) & (!g1906) & (g1907) & (g1908) & (!g820) & (g773)) + ((g1905) & (!g1906) & (g1907) & (g1908) & (g820) & (g773)) + ((g1905) & (g1906) & (!g1907) & (!g1908) & (!g820) & (!g773)) + ((g1905) & (g1906) & (!g1907) & (!g1908) & (g820) & (!g773)) + ((g1905) & (g1906) & (!g1907) & (g1908) & (!g820) & (!g773)) + ((g1905) & (g1906) & (!g1907) & (g1908) & (g820) & (!g773)) + ((g1905) & (g1906) & (!g1907) & (g1908) & (g820) & (g773)) + ((g1905) & (g1906) & (g1907) & (!g1908) & (!g820) & (!g773)) + ((g1905) & (g1906) & (g1907) & (!g1908) & (!g820) & (g773)) + ((g1905) & (g1906) & (g1907) & (!g1908) & (g820) & (!g773)) + ((g1905) & (g1906) & (g1907) & (g1908) & (!g820) & (!g773)) + ((g1905) & (g1906) & (g1907) & (g1908) & (!g820) & (g773)) + ((g1905) & (g1906) & (g1907) & (g1908) & (g820) & (!g773)) + ((g1905) & (g1906) & (g1907) & (g1908) & (g820) & (g773)));
	assign g1910 = (((!g1254) & (!g1255) & (!g1256) & (g1257) & (g677) & (g726)) + ((!g1254) & (!g1255) & (g1256) & (!g1257) & (!g677) & (g726)) + ((!g1254) & (!g1255) & (g1256) & (g1257) & (!g677) & (g726)) + ((!g1254) & (!g1255) & (g1256) & (g1257) & (g677) & (g726)) + ((!g1254) & (g1255) & (!g1256) & (!g1257) & (g677) & (!g726)) + ((!g1254) & (g1255) & (!g1256) & (g1257) & (g677) & (!g726)) + ((!g1254) & (g1255) & (!g1256) & (g1257) & (g677) & (g726)) + ((!g1254) & (g1255) & (g1256) & (!g1257) & (!g677) & (g726)) + ((!g1254) & (g1255) & (g1256) & (!g1257) & (g677) & (!g726)) + ((!g1254) & (g1255) & (g1256) & (g1257) & (!g677) & (g726)) + ((!g1254) & (g1255) & (g1256) & (g1257) & (g677) & (!g726)) + ((!g1254) & (g1255) & (g1256) & (g1257) & (g677) & (g726)) + ((g1254) & (!g1255) & (!g1256) & (!g1257) & (!g677) & (!g726)) + ((g1254) & (!g1255) & (!g1256) & (g1257) & (!g677) & (!g726)) + ((g1254) & (!g1255) & (!g1256) & (g1257) & (g677) & (g726)) + ((g1254) & (!g1255) & (g1256) & (!g1257) & (!g677) & (!g726)) + ((g1254) & (!g1255) & (g1256) & (!g1257) & (!g677) & (g726)) + ((g1254) & (!g1255) & (g1256) & (g1257) & (!g677) & (!g726)) + ((g1254) & (!g1255) & (g1256) & (g1257) & (!g677) & (g726)) + ((g1254) & (!g1255) & (g1256) & (g1257) & (g677) & (g726)) + ((g1254) & (g1255) & (!g1256) & (!g1257) & (!g677) & (!g726)) + ((g1254) & (g1255) & (!g1256) & (!g1257) & (g677) & (!g726)) + ((g1254) & (g1255) & (!g1256) & (g1257) & (!g677) & (!g726)) + ((g1254) & (g1255) & (!g1256) & (g1257) & (g677) & (!g726)) + ((g1254) & (g1255) & (!g1256) & (g1257) & (g677) & (g726)) + ((g1254) & (g1255) & (g1256) & (!g1257) & (!g677) & (!g726)) + ((g1254) & (g1255) & (g1256) & (!g1257) & (!g677) & (g726)) + ((g1254) & (g1255) & (g1256) & (!g1257) & (g677) & (!g726)) + ((g1254) & (g1255) & (g1256) & (g1257) & (!g677) & (!g726)) + ((g1254) & (g1255) & (g1256) & (g1257) & (!g677) & (g726)) + ((g1254) & (g1255) & (g1256) & (g1257) & (g677) & (!g726)) + ((g1254) & (g1255) & (g1256) & (g1257) & (g677) & (g726)));
	assign g1911 = (((!sk[57]) & (!g677) & (!g726) & (!g1259) & (g1260) & (!g1261)) + ((!sk[57]) & (!g677) & (!g726) & (!g1259) & (g1260) & (g1261)) + ((!sk[57]) & (!g677) & (!g726) & (g1259) & (!g1260) & (!g1261)) + ((!sk[57]) & (!g677) & (!g726) & (g1259) & (!g1260) & (g1261)) + ((!sk[57]) & (!g677) & (!g726) & (g1259) & (g1260) & (!g1261)) + ((!sk[57]) & (!g677) & (!g726) & (g1259) & (g1260) & (g1261)) + ((!sk[57]) & (!g677) & (g726) & (!g1259) & (!g1260) & (!g1261)) + ((!sk[57]) & (!g677) & (g726) & (!g1259) & (!g1260) & (g1261)) + ((!sk[57]) & (!g677) & (g726) & (!g1259) & (g1260) & (!g1261)) + ((!sk[57]) & (!g677) & (g726) & (!g1259) & (g1260) & (g1261)) + ((!sk[57]) & (!g677) & (g726) & (g1259) & (!g1260) & (!g1261)) + ((!sk[57]) & (!g677) & (g726) & (g1259) & (!g1260) & (g1261)) + ((!sk[57]) & (!g677) & (g726) & (g1259) & (g1260) & (!g1261)) + ((!sk[57]) & (!g677) & (g726) & (g1259) & (g1260) & (g1261)) + ((!sk[57]) & (g677) & (!g726) & (!g1259) & (g1260) & (!g1261)) + ((!sk[57]) & (g677) & (!g726) & (!g1259) & (g1260) & (g1261)) + ((!sk[57]) & (g677) & (!g726) & (g1259) & (!g1260) & (!g1261)) + ((!sk[57]) & (g677) & (!g726) & (g1259) & (!g1260) & (g1261)) + ((!sk[57]) & (g677) & (!g726) & (g1259) & (g1260) & (!g1261)) + ((!sk[57]) & (g677) & (!g726) & (g1259) & (g1260) & (g1261)) + ((!sk[57]) & (g677) & (g726) & (!g1259) & (!g1260) & (!g1261)) + ((!sk[57]) & (g677) & (g726) & (!g1259) & (!g1260) & (g1261)) + ((!sk[57]) & (g677) & (g726) & (!g1259) & (g1260) & (!g1261)) + ((!sk[57]) & (g677) & (g726) & (!g1259) & (g1260) & (g1261)) + ((!sk[57]) & (g677) & (g726) & (g1259) & (!g1260) & (!g1261)) + ((!sk[57]) & (g677) & (g726) & (g1259) & (!g1260) & (g1261)) + ((!sk[57]) & (g677) & (g726) & (g1259) & (g1260) & (!g1261)) + ((!sk[57]) & (g677) & (g726) & (g1259) & (g1260) & (g1261)) + ((sk[57]) & (!g677) & (g726) & (!g1259) & (!g1260) & (g1261)) + ((sk[57]) & (!g677) & (g726) & (!g1259) & (g1260) & (g1261)) + ((sk[57]) & (!g677) & (g726) & (g1259) & (!g1260) & (g1261)) + ((sk[57]) & (!g677) & (g726) & (g1259) & (g1260) & (g1261)) + ((sk[57]) & (g677) & (!g726) & (g1259) & (!g1260) & (!g1261)) + ((sk[57]) & (g677) & (!g726) & (g1259) & (!g1260) & (g1261)) + ((sk[57]) & (g677) & (!g726) & (g1259) & (g1260) & (!g1261)) + ((sk[57]) & (g677) & (!g726) & (g1259) & (g1260) & (g1261)) + ((sk[57]) & (g677) & (g726) & (!g1259) & (g1260) & (!g1261)) + ((sk[57]) & (g677) & (g726) & (!g1259) & (g1260) & (g1261)) + ((sk[57]) & (g677) & (g726) & (g1259) & (g1260) & (!g1261)) + ((sk[57]) & (g677) & (g726) & (g1259) & (g1260) & (g1261)));
	assign g1912 = (((!g1263) & (!g1264) & (!g1265) & (g1266) & (g677) & (g726)) + ((!g1263) & (!g1264) & (g1265) & (!g1266) & (!g677) & (g726)) + ((!g1263) & (!g1264) & (g1265) & (g1266) & (!g677) & (g726)) + ((!g1263) & (!g1264) & (g1265) & (g1266) & (g677) & (g726)) + ((!g1263) & (g1264) & (!g1265) & (!g1266) & (g677) & (!g726)) + ((!g1263) & (g1264) & (!g1265) & (g1266) & (g677) & (!g726)) + ((!g1263) & (g1264) & (!g1265) & (g1266) & (g677) & (g726)) + ((!g1263) & (g1264) & (g1265) & (!g1266) & (!g677) & (g726)) + ((!g1263) & (g1264) & (g1265) & (!g1266) & (g677) & (!g726)) + ((!g1263) & (g1264) & (g1265) & (g1266) & (!g677) & (g726)) + ((!g1263) & (g1264) & (g1265) & (g1266) & (g677) & (!g726)) + ((!g1263) & (g1264) & (g1265) & (g1266) & (g677) & (g726)) + ((g1263) & (!g1264) & (!g1265) & (!g1266) & (!g677) & (!g726)) + ((g1263) & (!g1264) & (!g1265) & (g1266) & (!g677) & (!g726)) + ((g1263) & (!g1264) & (!g1265) & (g1266) & (g677) & (g726)) + ((g1263) & (!g1264) & (g1265) & (!g1266) & (!g677) & (!g726)) + ((g1263) & (!g1264) & (g1265) & (!g1266) & (!g677) & (g726)) + ((g1263) & (!g1264) & (g1265) & (g1266) & (!g677) & (!g726)) + ((g1263) & (!g1264) & (g1265) & (g1266) & (!g677) & (g726)) + ((g1263) & (!g1264) & (g1265) & (g1266) & (g677) & (g726)) + ((g1263) & (g1264) & (!g1265) & (!g1266) & (!g677) & (!g726)) + ((g1263) & (g1264) & (!g1265) & (!g1266) & (g677) & (!g726)) + ((g1263) & (g1264) & (!g1265) & (g1266) & (!g677) & (!g726)) + ((g1263) & (g1264) & (!g1265) & (g1266) & (g677) & (!g726)) + ((g1263) & (g1264) & (!g1265) & (g1266) & (g677) & (g726)) + ((g1263) & (g1264) & (g1265) & (!g1266) & (!g677) & (!g726)) + ((g1263) & (g1264) & (g1265) & (!g1266) & (!g677) & (g726)) + ((g1263) & (g1264) & (g1265) & (!g1266) & (g677) & (!g726)) + ((g1263) & (g1264) & (g1265) & (g1266) & (!g677) & (!g726)) + ((g1263) & (g1264) & (g1265) & (g1266) & (!g677) & (g726)) + ((g1263) & (g1264) & (g1265) & (g1266) & (g677) & (!g726)) + ((g1263) & (g1264) & (g1265) & (g1266) & (g677) & (g726)));
	assign g1913 = (((!g1268) & (!g1269) & (!g1270) & (g1271) & (g677) & (g726)) + ((!g1268) & (!g1269) & (g1270) & (!g1271) & (!g677) & (g726)) + ((!g1268) & (!g1269) & (g1270) & (g1271) & (!g677) & (g726)) + ((!g1268) & (!g1269) & (g1270) & (g1271) & (g677) & (g726)) + ((!g1268) & (g1269) & (!g1270) & (!g1271) & (g677) & (!g726)) + ((!g1268) & (g1269) & (!g1270) & (g1271) & (g677) & (!g726)) + ((!g1268) & (g1269) & (!g1270) & (g1271) & (g677) & (g726)) + ((!g1268) & (g1269) & (g1270) & (!g1271) & (!g677) & (g726)) + ((!g1268) & (g1269) & (g1270) & (!g1271) & (g677) & (!g726)) + ((!g1268) & (g1269) & (g1270) & (g1271) & (!g677) & (g726)) + ((!g1268) & (g1269) & (g1270) & (g1271) & (g677) & (!g726)) + ((!g1268) & (g1269) & (g1270) & (g1271) & (g677) & (g726)) + ((g1268) & (!g1269) & (!g1270) & (!g1271) & (!g677) & (!g726)) + ((g1268) & (!g1269) & (!g1270) & (g1271) & (!g677) & (!g726)) + ((g1268) & (!g1269) & (!g1270) & (g1271) & (g677) & (g726)) + ((g1268) & (!g1269) & (g1270) & (!g1271) & (!g677) & (!g726)) + ((g1268) & (!g1269) & (g1270) & (!g1271) & (!g677) & (g726)) + ((g1268) & (!g1269) & (g1270) & (g1271) & (!g677) & (!g726)) + ((g1268) & (!g1269) & (g1270) & (g1271) & (!g677) & (g726)) + ((g1268) & (!g1269) & (g1270) & (g1271) & (g677) & (g726)) + ((g1268) & (g1269) & (!g1270) & (!g1271) & (!g677) & (!g726)) + ((g1268) & (g1269) & (!g1270) & (!g1271) & (g677) & (!g726)) + ((g1268) & (g1269) & (!g1270) & (g1271) & (!g677) & (!g726)) + ((g1268) & (g1269) & (!g1270) & (g1271) & (g677) & (!g726)) + ((g1268) & (g1269) & (!g1270) & (g1271) & (g677) & (g726)) + ((g1268) & (g1269) & (g1270) & (!g1271) & (!g677) & (!g726)) + ((g1268) & (g1269) & (g1270) & (!g1271) & (!g677) & (g726)) + ((g1268) & (g1269) & (g1270) & (!g1271) & (g677) & (!g726)) + ((g1268) & (g1269) & (g1270) & (g1271) & (!g677) & (!g726)) + ((g1268) & (g1269) & (g1270) & (g1271) & (!g677) & (g726)) + ((g1268) & (g1269) & (g1270) & (g1271) & (g677) & (!g726)) + ((g1268) & (g1269) & (g1270) & (g1271) & (g677) & (g726)));
	assign g1914 = (((!g820) & (!g773) & (!g1910) & (g1911) & (!g1912) & (!g1913)) + ((!g820) & (!g773) & (!g1910) & (g1911) & (!g1912) & (g1913)) + ((!g820) & (!g773) & (!g1910) & (g1911) & (g1912) & (!g1913)) + ((!g820) & (!g773) & (!g1910) & (g1911) & (g1912) & (g1913)) + ((!g820) & (!g773) & (g1910) & (g1911) & (!g1912) & (!g1913)) + ((!g820) & (!g773) & (g1910) & (g1911) & (!g1912) & (g1913)) + ((!g820) & (!g773) & (g1910) & (g1911) & (g1912) & (!g1913)) + ((!g820) & (!g773) & (g1910) & (g1911) & (g1912) & (g1913)) + ((!g820) & (g773) & (!g1910) & (!g1911) & (!g1912) & (g1913)) + ((!g820) & (g773) & (!g1910) & (!g1911) & (g1912) & (g1913)) + ((!g820) & (g773) & (!g1910) & (g1911) & (!g1912) & (g1913)) + ((!g820) & (g773) & (!g1910) & (g1911) & (g1912) & (g1913)) + ((!g820) & (g773) & (g1910) & (!g1911) & (!g1912) & (g1913)) + ((!g820) & (g773) & (g1910) & (!g1911) & (g1912) & (g1913)) + ((!g820) & (g773) & (g1910) & (g1911) & (!g1912) & (g1913)) + ((!g820) & (g773) & (g1910) & (g1911) & (g1912) & (g1913)) + ((g820) & (!g773) & (g1910) & (!g1911) & (!g1912) & (!g1913)) + ((g820) & (!g773) & (g1910) & (!g1911) & (!g1912) & (g1913)) + ((g820) & (!g773) & (g1910) & (!g1911) & (g1912) & (!g1913)) + ((g820) & (!g773) & (g1910) & (!g1911) & (g1912) & (g1913)) + ((g820) & (!g773) & (g1910) & (g1911) & (!g1912) & (!g1913)) + ((g820) & (!g773) & (g1910) & (g1911) & (!g1912) & (g1913)) + ((g820) & (!g773) & (g1910) & (g1911) & (g1912) & (!g1913)) + ((g820) & (!g773) & (g1910) & (g1911) & (g1912) & (g1913)) + ((g820) & (g773) & (!g1910) & (!g1911) & (g1912) & (!g1913)) + ((g820) & (g773) & (!g1910) & (!g1911) & (g1912) & (g1913)) + ((g820) & (g773) & (!g1910) & (g1911) & (g1912) & (!g1913)) + ((g820) & (g773) & (!g1910) & (g1911) & (g1912) & (g1913)) + ((g820) & (g773) & (g1910) & (!g1911) & (g1912) & (!g1913)) + ((g820) & (g773) & (g1910) & (!g1911) & (g1912) & (g1913)) + ((g820) & (g773) & (g1910) & (g1911) & (g1912) & (!g1913)) + ((g820) & (g773) & (g1910) & (g1911) & (g1912) & (g1913)));
	assign g1915 = (((!sk[61]) & (!g867) & (!g1909) & (g1914)) + ((!sk[61]) & (!g867) & (g1909) & (!g1914)) + ((!sk[61]) & (!g867) & (g1909) & (g1914)) + ((!sk[61]) & (g867) & (!g1909) & (g1914)) + ((!sk[61]) & (g867) & (g1909) & (!g1914)) + ((!sk[61]) & (g867) & (g1909) & (g1914)) + ((sk[61]) & (!g867) & (!g1909) & (g1914)) + ((sk[61]) & (!g867) & (g1909) & (g1914)) + ((sk[61]) & (g867) & (g1909) & (!g1914)) + ((sk[61]) & (g867) & (g1909) & (g1914)));
	assign g1916 = (((!g1593) & (!sk[62]) & (!g1605) & (!g1705) & (g59)) + ((!g1593) & (!sk[62]) & (!g1605) & (g1705) & (!g59)) + ((!g1593) & (!sk[62]) & (!g1605) & (g1705) & (g59)) + ((!g1593) & (!sk[62]) & (g1605) & (!g1705) & (!g59)) + ((!g1593) & (!sk[62]) & (g1605) & (!g1705) & (g59)) + ((!g1593) & (!sk[62]) & (g1605) & (g1705) & (!g59)) + ((!g1593) & (!sk[62]) & (g1605) & (g1705) & (g59)) + ((!g1593) & (sk[62]) & (!g1605) & (g1705) & (!g59)) + ((!g1593) & (sk[62]) & (!g1605) & (g1705) & (g59)) + ((g1593) & (!sk[62]) & (!g1605) & (!g1705) & (g59)) + ((g1593) & (!sk[62]) & (!g1605) & (g1705) & (!g59)) + ((g1593) & (!sk[62]) & (!g1605) & (g1705) & (g59)) + ((g1593) & (!sk[62]) & (g1605) & (!g1705) & (!g59)) + ((g1593) & (!sk[62]) & (g1605) & (!g1705) & (g59)) + ((g1593) & (!sk[62]) & (g1605) & (g1705) & (!g59)) + ((g1593) & (!sk[62]) & (g1605) & (g1705) & (g59)) + ((g1593) & (sk[62]) & (!g1605) & (!g1705) & (g59)) + ((g1593) & (sk[62]) & (!g1605) & (g1705) & (g59)) + ((g1593) & (sk[62]) & (g1605) & (!g1705) & (g59)) + ((g1593) & (sk[62]) & (g1605) & (g1705) & (g59)));
	assign g1917 = (((!g132) & (!g1592) & (g1606) & (!g136) & (!g1593) & (!g1605)) + ((!g132) & (g1592) & (!g1606) & (!g136) & (!g1593) & (!g1605)) + ((!g132) & (g1592) & (!g1606) & (!g136) & (!g1593) & (g1605)) + ((!g132) & (g1592) & (!g1606) & (!g136) & (g1593) & (!g1605)) + ((!g132) & (g1592) & (!g1606) & (!g136) & (g1593) & (g1605)) + ((!g132) & (g1592) & (g1606) & (!g136) & (!g1593) & (!g1605)) + ((g132) & (!g1592) & (!g1606) & (!g136) & (!g1593) & (!g1605)) + ((g132) & (!g1592) & (!g1606) & (!g136) & (!g1593) & (g1605)) + ((g132) & (!g1592) & (!g1606) & (!g136) & (g1593) & (!g1605)) + ((g132) & (!g1592) & (!g1606) & (!g136) & (g1593) & (g1605)) + ((g132) & (!g1592) & (g1606) & (!g136) & (!g1593) & (!g1605)) + ((g132) & (g1592) & (!g1606) & (!g136) & (!g1593) & (!g1605)) + ((g132) & (g1592) & (!g1606) & (!g136) & (!g1593) & (g1605)) + ((g132) & (g1592) & (!g1606) & (!g136) & (g1593) & (!g1605)) + ((g132) & (g1592) & (!g1606) & (!g136) & (g1593) & (g1605)) + ((g132) & (g1592) & (g1606) & (!g136) & (!g1593) & (!g1605)));
	assign g1918 = (((!g132) & (!g1592) & (g1604) & (!g1915) & (!g1916) & (g1917)) + ((!g132) & (!g1592) & (g1604) & (!g1915) & (g1916) & (g1917)) + ((!g132) & (!g1592) & (g1604) & (g1915) & (!g1916) & (g1917)) + ((!g132) & (!g1592) & (g1604) & (g1915) & (g1916) & (g1917)) + ((!g132) & (g1592) & (!g1604) & (!g1915) & (g1916) & (g1917)) + ((!g132) & (g1592) & (!g1604) & (g1915) & (g1916) & (g1917)) + ((!g132) & (g1592) & (g1604) & (!g1915) & (g1916) & (g1917)) + ((!g132) & (g1592) & (g1604) & (g1915) & (g1916) & (g1917)) + ((g132) & (!g1592) & (!g1604) & (g1915) & (!g1916) & (g1917)) + ((g132) & (!g1592) & (!g1604) & (g1915) & (g1916) & (g1917)) + ((g132) & (!g1592) & (g1604) & (g1915) & (!g1916) & (g1917)) + ((g132) & (!g1592) & (g1604) & (g1915) & (g1916) & (g1917)) + ((g132) & (g1592) & (!g1604) & (g1915) & (!g1916) & (g1917)) + ((g132) & (g1592) & (!g1604) & (g1915) & (g1916) & (g1917)) + ((g132) & (g1592) & (g1604) & (g1915) & (!g1916) & (g1917)) + ((g132) & (g1592) & (g1604) & (g1915) & (g1916) & (g1917)));
	assign g1919 = (((!g1278) & (!g1279) & (!g1280) & (g1281) & (g820) & (g773)) + ((!g1278) & (!g1279) & (g1280) & (!g1281) & (!g820) & (g773)) + ((!g1278) & (!g1279) & (g1280) & (g1281) & (!g820) & (g773)) + ((!g1278) & (!g1279) & (g1280) & (g1281) & (g820) & (g773)) + ((!g1278) & (g1279) & (!g1280) & (!g1281) & (g820) & (!g773)) + ((!g1278) & (g1279) & (!g1280) & (g1281) & (g820) & (!g773)) + ((!g1278) & (g1279) & (!g1280) & (g1281) & (g820) & (g773)) + ((!g1278) & (g1279) & (g1280) & (!g1281) & (!g820) & (g773)) + ((!g1278) & (g1279) & (g1280) & (!g1281) & (g820) & (!g773)) + ((!g1278) & (g1279) & (g1280) & (g1281) & (!g820) & (g773)) + ((!g1278) & (g1279) & (g1280) & (g1281) & (g820) & (!g773)) + ((!g1278) & (g1279) & (g1280) & (g1281) & (g820) & (g773)) + ((g1278) & (!g1279) & (!g1280) & (!g1281) & (!g820) & (!g773)) + ((g1278) & (!g1279) & (!g1280) & (g1281) & (!g820) & (!g773)) + ((g1278) & (!g1279) & (!g1280) & (g1281) & (g820) & (g773)) + ((g1278) & (!g1279) & (g1280) & (!g1281) & (!g820) & (!g773)) + ((g1278) & (!g1279) & (g1280) & (!g1281) & (!g820) & (g773)) + ((g1278) & (!g1279) & (g1280) & (g1281) & (!g820) & (!g773)) + ((g1278) & (!g1279) & (g1280) & (g1281) & (!g820) & (g773)) + ((g1278) & (!g1279) & (g1280) & (g1281) & (g820) & (g773)) + ((g1278) & (g1279) & (!g1280) & (!g1281) & (!g820) & (!g773)) + ((g1278) & (g1279) & (!g1280) & (!g1281) & (g820) & (!g773)) + ((g1278) & (g1279) & (!g1280) & (g1281) & (!g820) & (!g773)) + ((g1278) & (g1279) & (!g1280) & (g1281) & (g820) & (!g773)) + ((g1278) & (g1279) & (!g1280) & (g1281) & (g820) & (g773)) + ((g1278) & (g1279) & (g1280) & (!g1281) & (!g820) & (!g773)) + ((g1278) & (g1279) & (g1280) & (!g1281) & (!g820) & (g773)) + ((g1278) & (g1279) & (g1280) & (!g1281) & (g820) & (!g773)) + ((g1278) & (g1279) & (g1280) & (g1281) & (!g820) & (!g773)) + ((g1278) & (g1279) & (g1280) & (g1281) & (!g820) & (g773)) + ((g1278) & (g1279) & (g1280) & (g1281) & (g820) & (!g773)) + ((g1278) & (g1279) & (g1280) & (g1281) & (g820) & (g773)));
	assign g1920 = (((!g1283) & (!g1284) & (!g1285) & (g1286) & (g820) & (g773)) + ((!g1283) & (!g1284) & (g1285) & (!g1286) & (!g820) & (g773)) + ((!g1283) & (!g1284) & (g1285) & (g1286) & (!g820) & (g773)) + ((!g1283) & (!g1284) & (g1285) & (g1286) & (g820) & (g773)) + ((!g1283) & (g1284) & (!g1285) & (!g1286) & (g820) & (!g773)) + ((!g1283) & (g1284) & (!g1285) & (g1286) & (g820) & (!g773)) + ((!g1283) & (g1284) & (!g1285) & (g1286) & (g820) & (g773)) + ((!g1283) & (g1284) & (g1285) & (!g1286) & (!g820) & (g773)) + ((!g1283) & (g1284) & (g1285) & (!g1286) & (g820) & (!g773)) + ((!g1283) & (g1284) & (g1285) & (g1286) & (!g820) & (g773)) + ((!g1283) & (g1284) & (g1285) & (g1286) & (g820) & (!g773)) + ((!g1283) & (g1284) & (g1285) & (g1286) & (g820) & (g773)) + ((g1283) & (!g1284) & (!g1285) & (!g1286) & (!g820) & (!g773)) + ((g1283) & (!g1284) & (!g1285) & (g1286) & (!g820) & (!g773)) + ((g1283) & (!g1284) & (!g1285) & (g1286) & (g820) & (g773)) + ((g1283) & (!g1284) & (g1285) & (!g1286) & (!g820) & (!g773)) + ((g1283) & (!g1284) & (g1285) & (!g1286) & (!g820) & (g773)) + ((g1283) & (!g1284) & (g1285) & (g1286) & (!g820) & (!g773)) + ((g1283) & (!g1284) & (g1285) & (g1286) & (!g820) & (g773)) + ((g1283) & (!g1284) & (g1285) & (g1286) & (g820) & (g773)) + ((g1283) & (g1284) & (!g1285) & (!g1286) & (!g820) & (!g773)) + ((g1283) & (g1284) & (!g1285) & (!g1286) & (g820) & (!g773)) + ((g1283) & (g1284) & (!g1285) & (g1286) & (!g820) & (!g773)) + ((g1283) & (g1284) & (!g1285) & (g1286) & (g820) & (!g773)) + ((g1283) & (g1284) & (!g1285) & (g1286) & (g820) & (g773)) + ((g1283) & (g1284) & (g1285) & (!g1286) & (!g820) & (!g773)) + ((g1283) & (g1284) & (g1285) & (!g1286) & (!g820) & (g773)) + ((g1283) & (g1284) & (g1285) & (!g1286) & (g820) & (!g773)) + ((g1283) & (g1284) & (g1285) & (g1286) & (!g820) & (!g773)) + ((g1283) & (g1284) & (g1285) & (g1286) & (!g820) & (g773)) + ((g1283) & (g1284) & (g1285) & (g1286) & (g820) & (!g773)) + ((g1283) & (g1284) & (g1285) & (g1286) & (g820) & (g773)));
	assign g1921 = (((!g1288) & (!g1289) & (!g1290) & (g1291) & (g820) & (g773)) + ((!g1288) & (!g1289) & (g1290) & (!g1291) & (!g820) & (g773)) + ((!g1288) & (!g1289) & (g1290) & (g1291) & (!g820) & (g773)) + ((!g1288) & (!g1289) & (g1290) & (g1291) & (g820) & (g773)) + ((!g1288) & (g1289) & (!g1290) & (!g1291) & (g820) & (!g773)) + ((!g1288) & (g1289) & (!g1290) & (g1291) & (g820) & (!g773)) + ((!g1288) & (g1289) & (!g1290) & (g1291) & (g820) & (g773)) + ((!g1288) & (g1289) & (g1290) & (!g1291) & (!g820) & (g773)) + ((!g1288) & (g1289) & (g1290) & (!g1291) & (g820) & (!g773)) + ((!g1288) & (g1289) & (g1290) & (g1291) & (!g820) & (g773)) + ((!g1288) & (g1289) & (g1290) & (g1291) & (g820) & (!g773)) + ((!g1288) & (g1289) & (g1290) & (g1291) & (g820) & (g773)) + ((g1288) & (!g1289) & (!g1290) & (!g1291) & (!g820) & (!g773)) + ((g1288) & (!g1289) & (!g1290) & (g1291) & (!g820) & (!g773)) + ((g1288) & (!g1289) & (!g1290) & (g1291) & (g820) & (g773)) + ((g1288) & (!g1289) & (g1290) & (!g1291) & (!g820) & (!g773)) + ((g1288) & (!g1289) & (g1290) & (!g1291) & (!g820) & (g773)) + ((g1288) & (!g1289) & (g1290) & (g1291) & (!g820) & (!g773)) + ((g1288) & (!g1289) & (g1290) & (g1291) & (!g820) & (g773)) + ((g1288) & (!g1289) & (g1290) & (g1291) & (g820) & (g773)) + ((g1288) & (g1289) & (!g1290) & (!g1291) & (!g820) & (!g773)) + ((g1288) & (g1289) & (!g1290) & (!g1291) & (g820) & (!g773)) + ((g1288) & (g1289) & (!g1290) & (g1291) & (!g820) & (!g773)) + ((g1288) & (g1289) & (!g1290) & (g1291) & (g820) & (!g773)) + ((g1288) & (g1289) & (!g1290) & (g1291) & (g820) & (g773)) + ((g1288) & (g1289) & (g1290) & (!g1291) & (!g820) & (!g773)) + ((g1288) & (g1289) & (g1290) & (!g1291) & (!g820) & (g773)) + ((g1288) & (g1289) & (g1290) & (!g1291) & (g820) & (!g773)) + ((g1288) & (g1289) & (g1290) & (g1291) & (!g820) & (!g773)) + ((g1288) & (g1289) & (g1290) & (g1291) & (!g820) & (g773)) + ((g1288) & (g1289) & (g1290) & (g1291) & (g820) & (!g773)) + ((g1288) & (g1289) & (g1290) & (g1291) & (g820) & (g773)));
	assign g1922 = (((!g1293) & (!g1294) & (!g1295) & (g1296) & (g820) & (g773)) + ((!g1293) & (!g1294) & (g1295) & (!g1296) & (!g820) & (g773)) + ((!g1293) & (!g1294) & (g1295) & (g1296) & (!g820) & (g773)) + ((!g1293) & (!g1294) & (g1295) & (g1296) & (g820) & (g773)) + ((!g1293) & (g1294) & (!g1295) & (!g1296) & (g820) & (!g773)) + ((!g1293) & (g1294) & (!g1295) & (g1296) & (g820) & (!g773)) + ((!g1293) & (g1294) & (!g1295) & (g1296) & (g820) & (g773)) + ((!g1293) & (g1294) & (g1295) & (!g1296) & (!g820) & (g773)) + ((!g1293) & (g1294) & (g1295) & (!g1296) & (g820) & (!g773)) + ((!g1293) & (g1294) & (g1295) & (g1296) & (!g820) & (g773)) + ((!g1293) & (g1294) & (g1295) & (g1296) & (g820) & (!g773)) + ((!g1293) & (g1294) & (g1295) & (g1296) & (g820) & (g773)) + ((g1293) & (!g1294) & (!g1295) & (!g1296) & (!g820) & (!g773)) + ((g1293) & (!g1294) & (!g1295) & (g1296) & (!g820) & (!g773)) + ((g1293) & (!g1294) & (!g1295) & (g1296) & (g820) & (g773)) + ((g1293) & (!g1294) & (g1295) & (!g1296) & (!g820) & (!g773)) + ((g1293) & (!g1294) & (g1295) & (!g1296) & (!g820) & (g773)) + ((g1293) & (!g1294) & (g1295) & (g1296) & (!g820) & (!g773)) + ((g1293) & (!g1294) & (g1295) & (g1296) & (!g820) & (g773)) + ((g1293) & (!g1294) & (g1295) & (g1296) & (g820) & (g773)) + ((g1293) & (g1294) & (!g1295) & (!g1296) & (!g820) & (!g773)) + ((g1293) & (g1294) & (!g1295) & (!g1296) & (g820) & (!g773)) + ((g1293) & (g1294) & (!g1295) & (g1296) & (!g820) & (!g773)) + ((g1293) & (g1294) & (!g1295) & (g1296) & (g820) & (!g773)) + ((g1293) & (g1294) & (!g1295) & (g1296) & (g820) & (g773)) + ((g1293) & (g1294) & (g1295) & (!g1296) & (!g820) & (!g773)) + ((g1293) & (g1294) & (g1295) & (!g1296) & (!g820) & (g773)) + ((g1293) & (g1294) & (g1295) & (!g1296) & (g820) & (!g773)) + ((g1293) & (g1294) & (g1295) & (g1296) & (!g820) & (!g773)) + ((g1293) & (g1294) & (g1295) & (g1296) & (!g820) & (g773)) + ((g1293) & (g1294) & (g1295) & (g1296) & (g820) & (!g773)) + ((g1293) & (g1294) & (g1295) & (g1296) & (g820) & (g773)));
	assign g1923 = (((!g1919) & (!g1920) & (!g1921) & (g1922) & (g677) & (g726)) + ((!g1919) & (!g1920) & (g1921) & (!g1922) & (!g677) & (g726)) + ((!g1919) & (!g1920) & (g1921) & (g1922) & (!g677) & (g726)) + ((!g1919) & (!g1920) & (g1921) & (g1922) & (g677) & (g726)) + ((!g1919) & (g1920) & (!g1921) & (!g1922) & (g677) & (!g726)) + ((!g1919) & (g1920) & (!g1921) & (g1922) & (g677) & (!g726)) + ((!g1919) & (g1920) & (!g1921) & (g1922) & (g677) & (g726)) + ((!g1919) & (g1920) & (g1921) & (!g1922) & (!g677) & (g726)) + ((!g1919) & (g1920) & (g1921) & (!g1922) & (g677) & (!g726)) + ((!g1919) & (g1920) & (g1921) & (g1922) & (!g677) & (g726)) + ((!g1919) & (g1920) & (g1921) & (g1922) & (g677) & (!g726)) + ((!g1919) & (g1920) & (g1921) & (g1922) & (g677) & (g726)) + ((g1919) & (!g1920) & (!g1921) & (!g1922) & (!g677) & (!g726)) + ((g1919) & (!g1920) & (!g1921) & (g1922) & (!g677) & (!g726)) + ((g1919) & (!g1920) & (!g1921) & (g1922) & (g677) & (g726)) + ((g1919) & (!g1920) & (g1921) & (!g1922) & (!g677) & (!g726)) + ((g1919) & (!g1920) & (g1921) & (!g1922) & (!g677) & (g726)) + ((g1919) & (!g1920) & (g1921) & (g1922) & (!g677) & (!g726)) + ((g1919) & (!g1920) & (g1921) & (g1922) & (!g677) & (g726)) + ((g1919) & (!g1920) & (g1921) & (g1922) & (g677) & (g726)) + ((g1919) & (g1920) & (!g1921) & (!g1922) & (!g677) & (!g726)) + ((g1919) & (g1920) & (!g1921) & (!g1922) & (g677) & (!g726)) + ((g1919) & (g1920) & (!g1921) & (g1922) & (!g677) & (!g726)) + ((g1919) & (g1920) & (!g1921) & (g1922) & (g677) & (!g726)) + ((g1919) & (g1920) & (!g1921) & (g1922) & (g677) & (g726)) + ((g1919) & (g1920) & (g1921) & (!g1922) & (!g677) & (!g726)) + ((g1919) & (g1920) & (g1921) & (!g1922) & (!g677) & (g726)) + ((g1919) & (g1920) & (g1921) & (!g1922) & (g677) & (!g726)) + ((g1919) & (g1920) & (g1921) & (g1922) & (!g677) & (!g726)) + ((g1919) & (g1920) & (g1921) & (g1922) & (!g677) & (g726)) + ((g1919) & (g1920) & (g1921) & (g1922) & (g677) & (!g726)) + ((g1919) & (g1920) & (g1921) & (g1922) & (g677) & (g726)));
	assign g1924 = (((!g1299) & (!g1300) & (!g1301) & (g1302) & (g677) & (g726)) + ((!g1299) & (!g1300) & (g1301) & (!g1302) & (!g677) & (g726)) + ((!g1299) & (!g1300) & (g1301) & (g1302) & (!g677) & (g726)) + ((!g1299) & (!g1300) & (g1301) & (g1302) & (g677) & (g726)) + ((!g1299) & (g1300) & (!g1301) & (!g1302) & (g677) & (!g726)) + ((!g1299) & (g1300) & (!g1301) & (g1302) & (g677) & (!g726)) + ((!g1299) & (g1300) & (!g1301) & (g1302) & (g677) & (g726)) + ((!g1299) & (g1300) & (g1301) & (!g1302) & (!g677) & (g726)) + ((!g1299) & (g1300) & (g1301) & (!g1302) & (g677) & (!g726)) + ((!g1299) & (g1300) & (g1301) & (g1302) & (!g677) & (g726)) + ((!g1299) & (g1300) & (g1301) & (g1302) & (g677) & (!g726)) + ((!g1299) & (g1300) & (g1301) & (g1302) & (g677) & (g726)) + ((g1299) & (!g1300) & (!g1301) & (!g1302) & (!g677) & (!g726)) + ((g1299) & (!g1300) & (!g1301) & (g1302) & (!g677) & (!g726)) + ((g1299) & (!g1300) & (!g1301) & (g1302) & (g677) & (g726)) + ((g1299) & (!g1300) & (g1301) & (!g1302) & (!g677) & (!g726)) + ((g1299) & (!g1300) & (g1301) & (!g1302) & (!g677) & (g726)) + ((g1299) & (!g1300) & (g1301) & (g1302) & (!g677) & (!g726)) + ((g1299) & (!g1300) & (g1301) & (g1302) & (!g677) & (g726)) + ((g1299) & (!g1300) & (g1301) & (g1302) & (g677) & (g726)) + ((g1299) & (g1300) & (!g1301) & (!g1302) & (!g677) & (!g726)) + ((g1299) & (g1300) & (!g1301) & (!g1302) & (g677) & (!g726)) + ((g1299) & (g1300) & (!g1301) & (g1302) & (!g677) & (!g726)) + ((g1299) & (g1300) & (!g1301) & (g1302) & (g677) & (!g726)) + ((g1299) & (g1300) & (!g1301) & (g1302) & (g677) & (g726)) + ((g1299) & (g1300) & (g1301) & (!g1302) & (!g677) & (!g726)) + ((g1299) & (g1300) & (g1301) & (!g1302) & (!g677) & (g726)) + ((g1299) & (g1300) & (g1301) & (!g1302) & (g677) & (!g726)) + ((g1299) & (g1300) & (g1301) & (g1302) & (!g677) & (!g726)) + ((g1299) & (g1300) & (g1301) & (g1302) & (!g677) & (g726)) + ((g1299) & (g1300) & (g1301) & (g1302) & (g677) & (!g726)) + ((g1299) & (g1300) & (g1301) & (g1302) & (g677) & (g726)));
	assign g1925 = (((!g677) & (!g726) & (!g1304) & (!sk[71]) & (g1305) & (!g1306)) + ((!g677) & (!g726) & (!g1304) & (!sk[71]) & (g1305) & (g1306)) + ((!g677) & (!g726) & (g1304) & (!sk[71]) & (!g1305) & (!g1306)) + ((!g677) & (!g726) & (g1304) & (!sk[71]) & (!g1305) & (g1306)) + ((!g677) & (!g726) & (g1304) & (!sk[71]) & (g1305) & (!g1306)) + ((!g677) & (!g726) & (g1304) & (!sk[71]) & (g1305) & (g1306)) + ((!g677) & (g726) & (!g1304) & (!sk[71]) & (!g1305) & (!g1306)) + ((!g677) & (g726) & (!g1304) & (!sk[71]) & (!g1305) & (g1306)) + ((!g677) & (g726) & (!g1304) & (!sk[71]) & (g1305) & (!g1306)) + ((!g677) & (g726) & (!g1304) & (!sk[71]) & (g1305) & (g1306)) + ((!g677) & (g726) & (!g1304) & (sk[71]) & (!g1305) & (g1306)) + ((!g677) & (g726) & (!g1304) & (sk[71]) & (g1305) & (g1306)) + ((!g677) & (g726) & (g1304) & (!sk[71]) & (!g1305) & (!g1306)) + ((!g677) & (g726) & (g1304) & (!sk[71]) & (!g1305) & (g1306)) + ((!g677) & (g726) & (g1304) & (!sk[71]) & (g1305) & (!g1306)) + ((!g677) & (g726) & (g1304) & (!sk[71]) & (g1305) & (g1306)) + ((!g677) & (g726) & (g1304) & (sk[71]) & (!g1305) & (g1306)) + ((!g677) & (g726) & (g1304) & (sk[71]) & (g1305) & (g1306)) + ((g677) & (!g726) & (!g1304) & (!sk[71]) & (g1305) & (!g1306)) + ((g677) & (!g726) & (!g1304) & (!sk[71]) & (g1305) & (g1306)) + ((g677) & (!g726) & (g1304) & (!sk[71]) & (!g1305) & (!g1306)) + ((g677) & (!g726) & (g1304) & (!sk[71]) & (!g1305) & (g1306)) + ((g677) & (!g726) & (g1304) & (!sk[71]) & (g1305) & (!g1306)) + ((g677) & (!g726) & (g1304) & (!sk[71]) & (g1305) & (g1306)) + ((g677) & (!g726) & (g1304) & (sk[71]) & (!g1305) & (!g1306)) + ((g677) & (!g726) & (g1304) & (sk[71]) & (!g1305) & (g1306)) + ((g677) & (!g726) & (g1304) & (sk[71]) & (g1305) & (!g1306)) + ((g677) & (!g726) & (g1304) & (sk[71]) & (g1305) & (g1306)) + ((g677) & (g726) & (!g1304) & (!sk[71]) & (!g1305) & (!g1306)) + ((g677) & (g726) & (!g1304) & (!sk[71]) & (!g1305) & (g1306)) + ((g677) & (g726) & (!g1304) & (!sk[71]) & (g1305) & (!g1306)) + ((g677) & (g726) & (!g1304) & (!sk[71]) & (g1305) & (g1306)) + ((g677) & (g726) & (!g1304) & (sk[71]) & (g1305) & (!g1306)) + ((g677) & (g726) & (!g1304) & (sk[71]) & (g1305) & (g1306)) + ((g677) & (g726) & (g1304) & (!sk[71]) & (!g1305) & (!g1306)) + ((g677) & (g726) & (g1304) & (!sk[71]) & (!g1305) & (g1306)) + ((g677) & (g726) & (g1304) & (!sk[71]) & (g1305) & (!g1306)) + ((g677) & (g726) & (g1304) & (!sk[71]) & (g1305) & (g1306)) + ((g677) & (g726) & (g1304) & (sk[71]) & (g1305) & (!g1306)) + ((g677) & (g726) & (g1304) & (sk[71]) & (g1305) & (g1306)));
	assign g1926 = (((!g1308) & (!g1309) & (!g1310) & (g1311) & (g677) & (g726)) + ((!g1308) & (!g1309) & (g1310) & (!g1311) & (!g677) & (g726)) + ((!g1308) & (!g1309) & (g1310) & (g1311) & (!g677) & (g726)) + ((!g1308) & (!g1309) & (g1310) & (g1311) & (g677) & (g726)) + ((!g1308) & (g1309) & (!g1310) & (!g1311) & (g677) & (!g726)) + ((!g1308) & (g1309) & (!g1310) & (g1311) & (g677) & (!g726)) + ((!g1308) & (g1309) & (!g1310) & (g1311) & (g677) & (g726)) + ((!g1308) & (g1309) & (g1310) & (!g1311) & (!g677) & (g726)) + ((!g1308) & (g1309) & (g1310) & (!g1311) & (g677) & (!g726)) + ((!g1308) & (g1309) & (g1310) & (g1311) & (!g677) & (g726)) + ((!g1308) & (g1309) & (g1310) & (g1311) & (g677) & (!g726)) + ((!g1308) & (g1309) & (g1310) & (g1311) & (g677) & (g726)) + ((g1308) & (!g1309) & (!g1310) & (!g1311) & (!g677) & (!g726)) + ((g1308) & (!g1309) & (!g1310) & (g1311) & (!g677) & (!g726)) + ((g1308) & (!g1309) & (!g1310) & (g1311) & (g677) & (g726)) + ((g1308) & (!g1309) & (g1310) & (!g1311) & (!g677) & (!g726)) + ((g1308) & (!g1309) & (g1310) & (!g1311) & (!g677) & (g726)) + ((g1308) & (!g1309) & (g1310) & (g1311) & (!g677) & (!g726)) + ((g1308) & (!g1309) & (g1310) & (g1311) & (!g677) & (g726)) + ((g1308) & (!g1309) & (g1310) & (g1311) & (g677) & (g726)) + ((g1308) & (g1309) & (!g1310) & (!g1311) & (!g677) & (!g726)) + ((g1308) & (g1309) & (!g1310) & (!g1311) & (g677) & (!g726)) + ((g1308) & (g1309) & (!g1310) & (g1311) & (!g677) & (!g726)) + ((g1308) & (g1309) & (!g1310) & (g1311) & (g677) & (!g726)) + ((g1308) & (g1309) & (!g1310) & (g1311) & (g677) & (g726)) + ((g1308) & (g1309) & (g1310) & (!g1311) & (!g677) & (!g726)) + ((g1308) & (g1309) & (g1310) & (!g1311) & (!g677) & (g726)) + ((g1308) & (g1309) & (g1310) & (!g1311) & (g677) & (!g726)) + ((g1308) & (g1309) & (g1310) & (g1311) & (!g677) & (!g726)) + ((g1308) & (g1309) & (g1310) & (g1311) & (!g677) & (g726)) + ((g1308) & (g1309) & (g1310) & (g1311) & (g677) & (!g726)) + ((g1308) & (g1309) & (g1310) & (g1311) & (g677) & (g726)));
	assign g1927 = (((!g1313) & (!g1314) & (!g1315) & (g1316) & (g677) & (g726)) + ((!g1313) & (!g1314) & (g1315) & (!g1316) & (!g677) & (g726)) + ((!g1313) & (!g1314) & (g1315) & (g1316) & (!g677) & (g726)) + ((!g1313) & (!g1314) & (g1315) & (g1316) & (g677) & (g726)) + ((!g1313) & (g1314) & (!g1315) & (!g1316) & (g677) & (!g726)) + ((!g1313) & (g1314) & (!g1315) & (g1316) & (g677) & (!g726)) + ((!g1313) & (g1314) & (!g1315) & (g1316) & (g677) & (g726)) + ((!g1313) & (g1314) & (g1315) & (!g1316) & (!g677) & (g726)) + ((!g1313) & (g1314) & (g1315) & (!g1316) & (g677) & (!g726)) + ((!g1313) & (g1314) & (g1315) & (g1316) & (!g677) & (g726)) + ((!g1313) & (g1314) & (g1315) & (g1316) & (g677) & (!g726)) + ((!g1313) & (g1314) & (g1315) & (g1316) & (g677) & (g726)) + ((g1313) & (!g1314) & (!g1315) & (!g1316) & (!g677) & (!g726)) + ((g1313) & (!g1314) & (!g1315) & (g1316) & (!g677) & (!g726)) + ((g1313) & (!g1314) & (!g1315) & (g1316) & (g677) & (g726)) + ((g1313) & (!g1314) & (g1315) & (!g1316) & (!g677) & (!g726)) + ((g1313) & (!g1314) & (g1315) & (!g1316) & (!g677) & (g726)) + ((g1313) & (!g1314) & (g1315) & (g1316) & (!g677) & (!g726)) + ((g1313) & (!g1314) & (g1315) & (g1316) & (!g677) & (g726)) + ((g1313) & (!g1314) & (g1315) & (g1316) & (g677) & (g726)) + ((g1313) & (g1314) & (!g1315) & (!g1316) & (!g677) & (!g726)) + ((g1313) & (g1314) & (!g1315) & (!g1316) & (g677) & (!g726)) + ((g1313) & (g1314) & (!g1315) & (g1316) & (!g677) & (!g726)) + ((g1313) & (g1314) & (!g1315) & (g1316) & (g677) & (!g726)) + ((g1313) & (g1314) & (!g1315) & (g1316) & (g677) & (g726)) + ((g1313) & (g1314) & (g1315) & (!g1316) & (!g677) & (!g726)) + ((g1313) & (g1314) & (g1315) & (!g1316) & (!g677) & (g726)) + ((g1313) & (g1314) & (g1315) & (!g1316) & (g677) & (!g726)) + ((g1313) & (g1314) & (g1315) & (g1316) & (!g677) & (!g726)) + ((g1313) & (g1314) & (g1315) & (g1316) & (!g677) & (g726)) + ((g1313) & (g1314) & (g1315) & (g1316) & (g677) & (!g726)) + ((g1313) & (g1314) & (g1315) & (g1316) & (g677) & (g726)));
	assign g1928 = (((!g820) & (!g773) & (!g1924) & (g1925) & (!g1926) & (!g1927)) + ((!g820) & (!g773) & (!g1924) & (g1925) & (!g1926) & (g1927)) + ((!g820) & (!g773) & (!g1924) & (g1925) & (g1926) & (!g1927)) + ((!g820) & (!g773) & (!g1924) & (g1925) & (g1926) & (g1927)) + ((!g820) & (!g773) & (g1924) & (g1925) & (!g1926) & (!g1927)) + ((!g820) & (!g773) & (g1924) & (g1925) & (!g1926) & (g1927)) + ((!g820) & (!g773) & (g1924) & (g1925) & (g1926) & (!g1927)) + ((!g820) & (!g773) & (g1924) & (g1925) & (g1926) & (g1927)) + ((!g820) & (g773) & (!g1924) & (!g1925) & (!g1926) & (g1927)) + ((!g820) & (g773) & (!g1924) & (!g1925) & (g1926) & (g1927)) + ((!g820) & (g773) & (!g1924) & (g1925) & (!g1926) & (g1927)) + ((!g820) & (g773) & (!g1924) & (g1925) & (g1926) & (g1927)) + ((!g820) & (g773) & (g1924) & (!g1925) & (!g1926) & (g1927)) + ((!g820) & (g773) & (g1924) & (!g1925) & (g1926) & (g1927)) + ((!g820) & (g773) & (g1924) & (g1925) & (!g1926) & (g1927)) + ((!g820) & (g773) & (g1924) & (g1925) & (g1926) & (g1927)) + ((g820) & (!g773) & (g1924) & (!g1925) & (!g1926) & (!g1927)) + ((g820) & (!g773) & (g1924) & (!g1925) & (!g1926) & (g1927)) + ((g820) & (!g773) & (g1924) & (!g1925) & (g1926) & (!g1927)) + ((g820) & (!g773) & (g1924) & (!g1925) & (g1926) & (g1927)) + ((g820) & (!g773) & (g1924) & (g1925) & (!g1926) & (!g1927)) + ((g820) & (!g773) & (g1924) & (g1925) & (!g1926) & (g1927)) + ((g820) & (!g773) & (g1924) & (g1925) & (g1926) & (!g1927)) + ((g820) & (!g773) & (g1924) & (g1925) & (g1926) & (g1927)) + ((g820) & (g773) & (!g1924) & (!g1925) & (g1926) & (!g1927)) + ((g820) & (g773) & (!g1924) & (!g1925) & (g1926) & (g1927)) + ((g820) & (g773) & (!g1924) & (g1925) & (g1926) & (!g1927)) + ((g820) & (g773) & (!g1924) & (g1925) & (g1926) & (g1927)) + ((g820) & (g773) & (g1924) & (!g1925) & (g1926) & (!g1927)) + ((g820) & (g773) & (g1924) & (!g1925) & (g1926) & (g1927)) + ((g820) & (g773) & (g1924) & (g1925) & (g1926) & (!g1927)) + ((g820) & (g773) & (g1924) & (g1925) & (g1926) & (g1927)));
	assign g1929 = (((!sk[75]) & (!g867) & (!g1923) & (g1928)) + ((!sk[75]) & (!g867) & (g1923) & (!g1928)) + ((!sk[75]) & (!g867) & (g1923) & (g1928)) + ((!sk[75]) & (g867) & (!g1923) & (g1928)) + ((!sk[75]) & (g867) & (g1923) & (!g1928)) + ((!sk[75]) & (g867) & (g1923) & (g1928)) + ((sk[75]) & (!g867) & (!g1923) & (g1928)) + ((sk[75]) & (!g867) & (g1923) & (g1928)) + ((sk[75]) & (g867) & (g1923) & (!g1928)) + ((sk[75]) & (g867) & (g1923) & (g1928)));
	assign g1930 = (((!g1593) & (!g1605) & (!sk[76]) & (!g1720) & (g60)) + ((!g1593) & (!g1605) & (!sk[76]) & (g1720) & (!g60)) + ((!g1593) & (!g1605) & (!sk[76]) & (g1720) & (g60)) + ((!g1593) & (!g1605) & (sk[76]) & (g1720) & (!g60)) + ((!g1593) & (!g1605) & (sk[76]) & (g1720) & (g60)) + ((!g1593) & (g1605) & (!sk[76]) & (!g1720) & (!g60)) + ((!g1593) & (g1605) & (!sk[76]) & (!g1720) & (g60)) + ((!g1593) & (g1605) & (!sk[76]) & (g1720) & (!g60)) + ((!g1593) & (g1605) & (!sk[76]) & (g1720) & (g60)) + ((g1593) & (!g1605) & (!sk[76]) & (!g1720) & (g60)) + ((g1593) & (!g1605) & (!sk[76]) & (g1720) & (!g60)) + ((g1593) & (!g1605) & (!sk[76]) & (g1720) & (g60)) + ((g1593) & (!g1605) & (sk[76]) & (!g1720) & (g60)) + ((g1593) & (!g1605) & (sk[76]) & (g1720) & (g60)) + ((g1593) & (g1605) & (!sk[76]) & (!g1720) & (!g60)) + ((g1593) & (g1605) & (!sk[76]) & (!g1720) & (g60)) + ((g1593) & (g1605) & (!sk[76]) & (g1720) & (!g60)) + ((g1593) & (g1605) & (!sk[76]) & (g1720) & (g60)) + ((g1593) & (g1605) & (sk[76]) & (!g1720) & (g60)) + ((g1593) & (g1605) & (sk[76]) & (g1720) & (g60)));
	assign g1931 = (((!g132) & (!g1592) & (g1620) & (g1917) & (!g1929) & (!g1930)) + ((!g132) & (!g1592) & (g1620) & (g1917) & (!g1929) & (g1930)) + ((!g132) & (!g1592) & (g1620) & (g1917) & (g1929) & (!g1930)) + ((!g132) & (!g1592) & (g1620) & (g1917) & (g1929) & (g1930)) + ((!g132) & (g1592) & (!g1620) & (g1917) & (!g1929) & (g1930)) + ((!g132) & (g1592) & (!g1620) & (g1917) & (g1929) & (g1930)) + ((!g132) & (g1592) & (g1620) & (g1917) & (!g1929) & (g1930)) + ((!g132) & (g1592) & (g1620) & (g1917) & (g1929) & (g1930)) + ((g132) & (!g1592) & (!g1620) & (g1917) & (g1929) & (!g1930)) + ((g132) & (!g1592) & (!g1620) & (g1917) & (g1929) & (g1930)) + ((g132) & (!g1592) & (g1620) & (g1917) & (g1929) & (!g1930)) + ((g132) & (!g1592) & (g1620) & (g1917) & (g1929) & (g1930)) + ((g132) & (g1592) & (!g1620) & (g1917) & (g1929) & (!g1930)) + ((g132) & (g1592) & (!g1620) & (g1917) & (g1929) & (g1930)) + ((g132) & (g1592) & (g1620) & (g1917) & (g1929) & (!g1930)) + ((g132) & (g1592) & (g1620) & (g1917) & (g1929) & (g1930)));
	assign g1932 = (((!g1323) & (!g1328) & (!g1333) & (g1338) & (g677) & (g726)) + ((!g1323) & (!g1328) & (g1333) & (!g1338) & (!g677) & (g726)) + ((!g1323) & (!g1328) & (g1333) & (g1338) & (!g677) & (g726)) + ((!g1323) & (!g1328) & (g1333) & (g1338) & (g677) & (g726)) + ((!g1323) & (g1328) & (!g1333) & (!g1338) & (g677) & (!g726)) + ((!g1323) & (g1328) & (!g1333) & (g1338) & (g677) & (!g726)) + ((!g1323) & (g1328) & (!g1333) & (g1338) & (g677) & (g726)) + ((!g1323) & (g1328) & (g1333) & (!g1338) & (!g677) & (g726)) + ((!g1323) & (g1328) & (g1333) & (!g1338) & (g677) & (!g726)) + ((!g1323) & (g1328) & (g1333) & (g1338) & (!g677) & (g726)) + ((!g1323) & (g1328) & (g1333) & (g1338) & (g677) & (!g726)) + ((!g1323) & (g1328) & (g1333) & (g1338) & (g677) & (g726)) + ((g1323) & (!g1328) & (!g1333) & (!g1338) & (!g677) & (!g726)) + ((g1323) & (!g1328) & (!g1333) & (g1338) & (!g677) & (!g726)) + ((g1323) & (!g1328) & (!g1333) & (g1338) & (g677) & (g726)) + ((g1323) & (!g1328) & (g1333) & (!g1338) & (!g677) & (!g726)) + ((g1323) & (!g1328) & (g1333) & (!g1338) & (!g677) & (g726)) + ((g1323) & (!g1328) & (g1333) & (g1338) & (!g677) & (!g726)) + ((g1323) & (!g1328) & (g1333) & (g1338) & (!g677) & (g726)) + ((g1323) & (!g1328) & (g1333) & (g1338) & (g677) & (g726)) + ((g1323) & (g1328) & (!g1333) & (!g1338) & (!g677) & (!g726)) + ((g1323) & (g1328) & (!g1333) & (!g1338) & (g677) & (!g726)) + ((g1323) & (g1328) & (!g1333) & (g1338) & (!g677) & (!g726)) + ((g1323) & (g1328) & (!g1333) & (g1338) & (g677) & (!g726)) + ((g1323) & (g1328) & (!g1333) & (g1338) & (g677) & (g726)) + ((g1323) & (g1328) & (g1333) & (!g1338) & (!g677) & (!g726)) + ((g1323) & (g1328) & (g1333) & (!g1338) & (!g677) & (g726)) + ((g1323) & (g1328) & (g1333) & (!g1338) & (g677) & (!g726)) + ((g1323) & (g1328) & (g1333) & (g1338) & (!g677) & (!g726)) + ((g1323) & (g1328) & (g1333) & (g1338) & (!g677) & (g726)) + ((g1323) & (g1328) & (g1333) & (g1338) & (g677) & (!g726)) + ((g1323) & (g1328) & (g1333) & (g1338) & (g677) & (g726)));
	assign g1933 = (((!g1324) & (!g1329) & (!g1334) & (g1339) & (g677) & (g726)) + ((!g1324) & (!g1329) & (g1334) & (!g1339) & (!g677) & (g726)) + ((!g1324) & (!g1329) & (g1334) & (g1339) & (!g677) & (g726)) + ((!g1324) & (!g1329) & (g1334) & (g1339) & (g677) & (g726)) + ((!g1324) & (g1329) & (!g1334) & (!g1339) & (g677) & (!g726)) + ((!g1324) & (g1329) & (!g1334) & (g1339) & (g677) & (!g726)) + ((!g1324) & (g1329) & (!g1334) & (g1339) & (g677) & (g726)) + ((!g1324) & (g1329) & (g1334) & (!g1339) & (!g677) & (g726)) + ((!g1324) & (g1329) & (g1334) & (!g1339) & (g677) & (!g726)) + ((!g1324) & (g1329) & (g1334) & (g1339) & (!g677) & (g726)) + ((!g1324) & (g1329) & (g1334) & (g1339) & (g677) & (!g726)) + ((!g1324) & (g1329) & (g1334) & (g1339) & (g677) & (g726)) + ((g1324) & (!g1329) & (!g1334) & (!g1339) & (!g677) & (!g726)) + ((g1324) & (!g1329) & (!g1334) & (g1339) & (!g677) & (!g726)) + ((g1324) & (!g1329) & (!g1334) & (g1339) & (g677) & (g726)) + ((g1324) & (!g1329) & (g1334) & (!g1339) & (!g677) & (!g726)) + ((g1324) & (!g1329) & (g1334) & (!g1339) & (!g677) & (g726)) + ((g1324) & (!g1329) & (g1334) & (g1339) & (!g677) & (!g726)) + ((g1324) & (!g1329) & (g1334) & (g1339) & (!g677) & (g726)) + ((g1324) & (!g1329) & (g1334) & (g1339) & (g677) & (g726)) + ((g1324) & (g1329) & (!g1334) & (!g1339) & (!g677) & (!g726)) + ((g1324) & (g1329) & (!g1334) & (!g1339) & (g677) & (!g726)) + ((g1324) & (g1329) & (!g1334) & (g1339) & (!g677) & (!g726)) + ((g1324) & (g1329) & (!g1334) & (g1339) & (g677) & (!g726)) + ((g1324) & (g1329) & (!g1334) & (g1339) & (g677) & (g726)) + ((g1324) & (g1329) & (g1334) & (!g1339) & (!g677) & (!g726)) + ((g1324) & (g1329) & (g1334) & (!g1339) & (!g677) & (g726)) + ((g1324) & (g1329) & (g1334) & (!g1339) & (g677) & (!g726)) + ((g1324) & (g1329) & (g1334) & (g1339) & (!g677) & (!g726)) + ((g1324) & (g1329) & (g1334) & (g1339) & (!g677) & (g726)) + ((g1324) & (g1329) & (g1334) & (g1339) & (g677) & (!g726)) + ((g1324) & (g1329) & (g1334) & (g1339) & (g677) & (g726)));
	assign g1934 = (((!g1325) & (!g1330) & (!g1335) & (g1340) & (g677) & (g726)) + ((!g1325) & (!g1330) & (g1335) & (!g1340) & (!g677) & (g726)) + ((!g1325) & (!g1330) & (g1335) & (g1340) & (!g677) & (g726)) + ((!g1325) & (!g1330) & (g1335) & (g1340) & (g677) & (g726)) + ((!g1325) & (g1330) & (!g1335) & (!g1340) & (g677) & (!g726)) + ((!g1325) & (g1330) & (!g1335) & (g1340) & (g677) & (!g726)) + ((!g1325) & (g1330) & (!g1335) & (g1340) & (g677) & (g726)) + ((!g1325) & (g1330) & (g1335) & (!g1340) & (!g677) & (g726)) + ((!g1325) & (g1330) & (g1335) & (!g1340) & (g677) & (!g726)) + ((!g1325) & (g1330) & (g1335) & (g1340) & (!g677) & (g726)) + ((!g1325) & (g1330) & (g1335) & (g1340) & (g677) & (!g726)) + ((!g1325) & (g1330) & (g1335) & (g1340) & (g677) & (g726)) + ((g1325) & (!g1330) & (!g1335) & (!g1340) & (!g677) & (!g726)) + ((g1325) & (!g1330) & (!g1335) & (g1340) & (!g677) & (!g726)) + ((g1325) & (!g1330) & (!g1335) & (g1340) & (g677) & (g726)) + ((g1325) & (!g1330) & (g1335) & (!g1340) & (!g677) & (!g726)) + ((g1325) & (!g1330) & (g1335) & (!g1340) & (!g677) & (g726)) + ((g1325) & (!g1330) & (g1335) & (g1340) & (!g677) & (!g726)) + ((g1325) & (!g1330) & (g1335) & (g1340) & (!g677) & (g726)) + ((g1325) & (!g1330) & (g1335) & (g1340) & (g677) & (g726)) + ((g1325) & (g1330) & (!g1335) & (!g1340) & (!g677) & (!g726)) + ((g1325) & (g1330) & (!g1335) & (!g1340) & (g677) & (!g726)) + ((g1325) & (g1330) & (!g1335) & (g1340) & (!g677) & (!g726)) + ((g1325) & (g1330) & (!g1335) & (g1340) & (g677) & (!g726)) + ((g1325) & (g1330) & (!g1335) & (g1340) & (g677) & (g726)) + ((g1325) & (g1330) & (g1335) & (!g1340) & (!g677) & (!g726)) + ((g1325) & (g1330) & (g1335) & (!g1340) & (!g677) & (g726)) + ((g1325) & (g1330) & (g1335) & (!g1340) & (g677) & (!g726)) + ((g1325) & (g1330) & (g1335) & (g1340) & (!g677) & (!g726)) + ((g1325) & (g1330) & (g1335) & (g1340) & (!g677) & (g726)) + ((g1325) & (g1330) & (g1335) & (g1340) & (g677) & (!g726)) + ((g1325) & (g1330) & (g1335) & (g1340) & (g677) & (g726)));
	assign g1935 = (((!g1326) & (!g1331) & (!g1336) & (g1341) & (g677) & (g726)) + ((!g1326) & (!g1331) & (g1336) & (!g1341) & (!g677) & (g726)) + ((!g1326) & (!g1331) & (g1336) & (g1341) & (!g677) & (g726)) + ((!g1326) & (!g1331) & (g1336) & (g1341) & (g677) & (g726)) + ((!g1326) & (g1331) & (!g1336) & (!g1341) & (g677) & (!g726)) + ((!g1326) & (g1331) & (!g1336) & (g1341) & (g677) & (!g726)) + ((!g1326) & (g1331) & (!g1336) & (g1341) & (g677) & (g726)) + ((!g1326) & (g1331) & (g1336) & (!g1341) & (!g677) & (g726)) + ((!g1326) & (g1331) & (g1336) & (!g1341) & (g677) & (!g726)) + ((!g1326) & (g1331) & (g1336) & (g1341) & (!g677) & (g726)) + ((!g1326) & (g1331) & (g1336) & (g1341) & (g677) & (!g726)) + ((!g1326) & (g1331) & (g1336) & (g1341) & (g677) & (g726)) + ((g1326) & (!g1331) & (!g1336) & (!g1341) & (!g677) & (!g726)) + ((g1326) & (!g1331) & (!g1336) & (g1341) & (!g677) & (!g726)) + ((g1326) & (!g1331) & (!g1336) & (g1341) & (g677) & (g726)) + ((g1326) & (!g1331) & (g1336) & (!g1341) & (!g677) & (!g726)) + ((g1326) & (!g1331) & (g1336) & (!g1341) & (!g677) & (g726)) + ((g1326) & (!g1331) & (g1336) & (g1341) & (!g677) & (!g726)) + ((g1326) & (!g1331) & (g1336) & (g1341) & (!g677) & (g726)) + ((g1326) & (!g1331) & (g1336) & (g1341) & (g677) & (g726)) + ((g1326) & (g1331) & (!g1336) & (!g1341) & (!g677) & (!g726)) + ((g1326) & (g1331) & (!g1336) & (!g1341) & (g677) & (!g726)) + ((g1326) & (g1331) & (!g1336) & (g1341) & (!g677) & (!g726)) + ((g1326) & (g1331) & (!g1336) & (g1341) & (g677) & (!g726)) + ((g1326) & (g1331) & (!g1336) & (g1341) & (g677) & (g726)) + ((g1326) & (g1331) & (g1336) & (!g1341) & (!g677) & (!g726)) + ((g1326) & (g1331) & (g1336) & (!g1341) & (!g677) & (g726)) + ((g1326) & (g1331) & (g1336) & (!g1341) & (g677) & (!g726)) + ((g1326) & (g1331) & (g1336) & (g1341) & (!g677) & (!g726)) + ((g1326) & (g1331) & (g1336) & (g1341) & (!g677) & (g726)) + ((g1326) & (g1331) & (g1336) & (g1341) & (g677) & (!g726)) + ((g1326) & (g1331) & (g1336) & (g1341) & (g677) & (g726)));
	assign g1936 = (((!g1932) & (!g1933) & (!g1934) & (g1935) & (g820) & (g773)) + ((!g1932) & (!g1933) & (g1934) & (!g1935) & (!g820) & (g773)) + ((!g1932) & (!g1933) & (g1934) & (g1935) & (!g820) & (g773)) + ((!g1932) & (!g1933) & (g1934) & (g1935) & (g820) & (g773)) + ((!g1932) & (g1933) & (!g1934) & (!g1935) & (g820) & (!g773)) + ((!g1932) & (g1933) & (!g1934) & (g1935) & (g820) & (!g773)) + ((!g1932) & (g1933) & (!g1934) & (g1935) & (g820) & (g773)) + ((!g1932) & (g1933) & (g1934) & (!g1935) & (!g820) & (g773)) + ((!g1932) & (g1933) & (g1934) & (!g1935) & (g820) & (!g773)) + ((!g1932) & (g1933) & (g1934) & (g1935) & (!g820) & (g773)) + ((!g1932) & (g1933) & (g1934) & (g1935) & (g820) & (!g773)) + ((!g1932) & (g1933) & (g1934) & (g1935) & (g820) & (g773)) + ((g1932) & (!g1933) & (!g1934) & (!g1935) & (!g820) & (!g773)) + ((g1932) & (!g1933) & (!g1934) & (g1935) & (!g820) & (!g773)) + ((g1932) & (!g1933) & (!g1934) & (g1935) & (g820) & (g773)) + ((g1932) & (!g1933) & (g1934) & (!g1935) & (!g820) & (!g773)) + ((g1932) & (!g1933) & (g1934) & (!g1935) & (!g820) & (g773)) + ((g1932) & (!g1933) & (g1934) & (g1935) & (!g820) & (!g773)) + ((g1932) & (!g1933) & (g1934) & (g1935) & (!g820) & (g773)) + ((g1932) & (!g1933) & (g1934) & (g1935) & (g820) & (g773)) + ((g1932) & (g1933) & (!g1934) & (!g1935) & (!g820) & (!g773)) + ((g1932) & (g1933) & (!g1934) & (!g1935) & (g820) & (!g773)) + ((g1932) & (g1933) & (!g1934) & (g1935) & (!g820) & (!g773)) + ((g1932) & (g1933) & (!g1934) & (g1935) & (g820) & (!g773)) + ((g1932) & (g1933) & (!g1934) & (g1935) & (g820) & (g773)) + ((g1932) & (g1933) & (g1934) & (!g1935) & (!g820) & (!g773)) + ((g1932) & (g1933) & (g1934) & (!g1935) & (!g820) & (g773)) + ((g1932) & (g1933) & (g1934) & (!g1935) & (g820) & (!g773)) + ((g1932) & (g1933) & (g1934) & (g1935) & (!g820) & (!g773)) + ((g1932) & (g1933) & (g1934) & (g1935) & (!g820) & (g773)) + ((g1932) & (g1933) & (g1934) & (g1935) & (g820) & (!g773)) + ((g1932) & (g1933) & (g1934) & (g1935) & (g820) & (g773)));
	assign g1937 = (((!g1344) & (!g1345) & (!g1346) & (g1347) & (g677) & (g726)) + ((!g1344) & (!g1345) & (g1346) & (!g1347) & (!g677) & (g726)) + ((!g1344) & (!g1345) & (g1346) & (g1347) & (!g677) & (g726)) + ((!g1344) & (!g1345) & (g1346) & (g1347) & (g677) & (g726)) + ((!g1344) & (g1345) & (!g1346) & (!g1347) & (g677) & (!g726)) + ((!g1344) & (g1345) & (!g1346) & (g1347) & (g677) & (!g726)) + ((!g1344) & (g1345) & (!g1346) & (g1347) & (g677) & (g726)) + ((!g1344) & (g1345) & (g1346) & (!g1347) & (!g677) & (g726)) + ((!g1344) & (g1345) & (g1346) & (!g1347) & (g677) & (!g726)) + ((!g1344) & (g1345) & (g1346) & (g1347) & (!g677) & (g726)) + ((!g1344) & (g1345) & (g1346) & (g1347) & (g677) & (!g726)) + ((!g1344) & (g1345) & (g1346) & (g1347) & (g677) & (g726)) + ((g1344) & (!g1345) & (!g1346) & (!g1347) & (!g677) & (!g726)) + ((g1344) & (!g1345) & (!g1346) & (g1347) & (!g677) & (!g726)) + ((g1344) & (!g1345) & (!g1346) & (g1347) & (g677) & (g726)) + ((g1344) & (!g1345) & (g1346) & (!g1347) & (!g677) & (!g726)) + ((g1344) & (!g1345) & (g1346) & (!g1347) & (!g677) & (g726)) + ((g1344) & (!g1345) & (g1346) & (g1347) & (!g677) & (!g726)) + ((g1344) & (!g1345) & (g1346) & (g1347) & (!g677) & (g726)) + ((g1344) & (!g1345) & (g1346) & (g1347) & (g677) & (g726)) + ((g1344) & (g1345) & (!g1346) & (!g1347) & (!g677) & (!g726)) + ((g1344) & (g1345) & (!g1346) & (!g1347) & (g677) & (!g726)) + ((g1344) & (g1345) & (!g1346) & (g1347) & (!g677) & (!g726)) + ((g1344) & (g1345) & (!g1346) & (g1347) & (g677) & (!g726)) + ((g1344) & (g1345) & (!g1346) & (g1347) & (g677) & (g726)) + ((g1344) & (g1345) & (g1346) & (!g1347) & (!g677) & (!g726)) + ((g1344) & (g1345) & (g1346) & (!g1347) & (!g677) & (g726)) + ((g1344) & (g1345) & (g1346) & (!g1347) & (g677) & (!g726)) + ((g1344) & (g1345) & (g1346) & (g1347) & (!g677) & (!g726)) + ((g1344) & (g1345) & (g1346) & (g1347) & (!g677) & (g726)) + ((g1344) & (g1345) & (g1346) & (g1347) & (g677) & (!g726)) + ((g1344) & (g1345) & (g1346) & (g1347) & (g677) & (g726)));
	assign g1938 = (((!g677) & (!g726) & (!g1349) & (g1350) & (!sk[84]) & (!g1351)) + ((!g677) & (!g726) & (!g1349) & (g1350) & (!sk[84]) & (g1351)) + ((!g677) & (!g726) & (g1349) & (!g1350) & (!sk[84]) & (!g1351)) + ((!g677) & (!g726) & (g1349) & (!g1350) & (!sk[84]) & (g1351)) + ((!g677) & (!g726) & (g1349) & (g1350) & (!sk[84]) & (!g1351)) + ((!g677) & (!g726) & (g1349) & (g1350) & (!sk[84]) & (g1351)) + ((!g677) & (g726) & (!g1349) & (!g1350) & (!sk[84]) & (!g1351)) + ((!g677) & (g726) & (!g1349) & (!g1350) & (!sk[84]) & (g1351)) + ((!g677) & (g726) & (!g1349) & (!g1350) & (sk[84]) & (g1351)) + ((!g677) & (g726) & (!g1349) & (g1350) & (!sk[84]) & (!g1351)) + ((!g677) & (g726) & (!g1349) & (g1350) & (!sk[84]) & (g1351)) + ((!g677) & (g726) & (!g1349) & (g1350) & (sk[84]) & (g1351)) + ((!g677) & (g726) & (g1349) & (!g1350) & (!sk[84]) & (!g1351)) + ((!g677) & (g726) & (g1349) & (!g1350) & (!sk[84]) & (g1351)) + ((!g677) & (g726) & (g1349) & (!g1350) & (sk[84]) & (g1351)) + ((!g677) & (g726) & (g1349) & (g1350) & (!sk[84]) & (!g1351)) + ((!g677) & (g726) & (g1349) & (g1350) & (!sk[84]) & (g1351)) + ((!g677) & (g726) & (g1349) & (g1350) & (sk[84]) & (g1351)) + ((g677) & (!g726) & (!g1349) & (g1350) & (!sk[84]) & (!g1351)) + ((g677) & (!g726) & (!g1349) & (g1350) & (!sk[84]) & (g1351)) + ((g677) & (!g726) & (g1349) & (!g1350) & (!sk[84]) & (!g1351)) + ((g677) & (!g726) & (g1349) & (!g1350) & (!sk[84]) & (g1351)) + ((g677) & (!g726) & (g1349) & (!g1350) & (sk[84]) & (!g1351)) + ((g677) & (!g726) & (g1349) & (!g1350) & (sk[84]) & (g1351)) + ((g677) & (!g726) & (g1349) & (g1350) & (!sk[84]) & (!g1351)) + ((g677) & (!g726) & (g1349) & (g1350) & (!sk[84]) & (g1351)) + ((g677) & (!g726) & (g1349) & (g1350) & (sk[84]) & (!g1351)) + ((g677) & (!g726) & (g1349) & (g1350) & (sk[84]) & (g1351)) + ((g677) & (g726) & (!g1349) & (!g1350) & (!sk[84]) & (!g1351)) + ((g677) & (g726) & (!g1349) & (!g1350) & (!sk[84]) & (g1351)) + ((g677) & (g726) & (!g1349) & (g1350) & (!sk[84]) & (!g1351)) + ((g677) & (g726) & (!g1349) & (g1350) & (!sk[84]) & (g1351)) + ((g677) & (g726) & (!g1349) & (g1350) & (sk[84]) & (!g1351)) + ((g677) & (g726) & (!g1349) & (g1350) & (sk[84]) & (g1351)) + ((g677) & (g726) & (g1349) & (!g1350) & (!sk[84]) & (!g1351)) + ((g677) & (g726) & (g1349) & (!g1350) & (!sk[84]) & (g1351)) + ((g677) & (g726) & (g1349) & (g1350) & (!sk[84]) & (!g1351)) + ((g677) & (g726) & (g1349) & (g1350) & (!sk[84]) & (g1351)) + ((g677) & (g726) & (g1349) & (g1350) & (sk[84]) & (!g1351)) + ((g677) & (g726) & (g1349) & (g1350) & (sk[84]) & (g1351)));
	assign g1939 = (((!g1353) & (!g1354) & (!g1355) & (g1356) & (g677) & (g726)) + ((!g1353) & (!g1354) & (g1355) & (!g1356) & (!g677) & (g726)) + ((!g1353) & (!g1354) & (g1355) & (g1356) & (!g677) & (g726)) + ((!g1353) & (!g1354) & (g1355) & (g1356) & (g677) & (g726)) + ((!g1353) & (g1354) & (!g1355) & (!g1356) & (g677) & (!g726)) + ((!g1353) & (g1354) & (!g1355) & (g1356) & (g677) & (!g726)) + ((!g1353) & (g1354) & (!g1355) & (g1356) & (g677) & (g726)) + ((!g1353) & (g1354) & (g1355) & (!g1356) & (!g677) & (g726)) + ((!g1353) & (g1354) & (g1355) & (!g1356) & (g677) & (!g726)) + ((!g1353) & (g1354) & (g1355) & (g1356) & (!g677) & (g726)) + ((!g1353) & (g1354) & (g1355) & (g1356) & (g677) & (!g726)) + ((!g1353) & (g1354) & (g1355) & (g1356) & (g677) & (g726)) + ((g1353) & (!g1354) & (!g1355) & (!g1356) & (!g677) & (!g726)) + ((g1353) & (!g1354) & (!g1355) & (g1356) & (!g677) & (!g726)) + ((g1353) & (!g1354) & (!g1355) & (g1356) & (g677) & (g726)) + ((g1353) & (!g1354) & (g1355) & (!g1356) & (!g677) & (!g726)) + ((g1353) & (!g1354) & (g1355) & (!g1356) & (!g677) & (g726)) + ((g1353) & (!g1354) & (g1355) & (g1356) & (!g677) & (!g726)) + ((g1353) & (!g1354) & (g1355) & (g1356) & (!g677) & (g726)) + ((g1353) & (!g1354) & (g1355) & (g1356) & (g677) & (g726)) + ((g1353) & (g1354) & (!g1355) & (!g1356) & (!g677) & (!g726)) + ((g1353) & (g1354) & (!g1355) & (!g1356) & (g677) & (!g726)) + ((g1353) & (g1354) & (!g1355) & (g1356) & (!g677) & (!g726)) + ((g1353) & (g1354) & (!g1355) & (g1356) & (g677) & (!g726)) + ((g1353) & (g1354) & (!g1355) & (g1356) & (g677) & (g726)) + ((g1353) & (g1354) & (g1355) & (!g1356) & (!g677) & (!g726)) + ((g1353) & (g1354) & (g1355) & (!g1356) & (!g677) & (g726)) + ((g1353) & (g1354) & (g1355) & (!g1356) & (g677) & (!g726)) + ((g1353) & (g1354) & (g1355) & (g1356) & (!g677) & (!g726)) + ((g1353) & (g1354) & (g1355) & (g1356) & (!g677) & (g726)) + ((g1353) & (g1354) & (g1355) & (g1356) & (g677) & (!g726)) + ((g1353) & (g1354) & (g1355) & (g1356) & (g677) & (g726)));
	assign g1940 = (((!g1358) & (!g1359) & (!g1360) & (g1361) & (g677) & (g726)) + ((!g1358) & (!g1359) & (g1360) & (!g1361) & (!g677) & (g726)) + ((!g1358) & (!g1359) & (g1360) & (g1361) & (!g677) & (g726)) + ((!g1358) & (!g1359) & (g1360) & (g1361) & (g677) & (g726)) + ((!g1358) & (g1359) & (!g1360) & (!g1361) & (g677) & (!g726)) + ((!g1358) & (g1359) & (!g1360) & (g1361) & (g677) & (!g726)) + ((!g1358) & (g1359) & (!g1360) & (g1361) & (g677) & (g726)) + ((!g1358) & (g1359) & (g1360) & (!g1361) & (!g677) & (g726)) + ((!g1358) & (g1359) & (g1360) & (!g1361) & (g677) & (!g726)) + ((!g1358) & (g1359) & (g1360) & (g1361) & (!g677) & (g726)) + ((!g1358) & (g1359) & (g1360) & (g1361) & (g677) & (!g726)) + ((!g1358) & (g1359) & (g1360) & (g1361) & (g677) & (g726)) + ((g1358) & (!g1359) & (!g1360) & (!g1361) & (!g677) & (!g726)) + ((g1358) & (!g1359) & (!g1360) & (g1361) & (!g677) & (!g726)) + ((g1358) & (!g1359) & (!g1360) & (g1361) & (g677) & (g726)) + ((g1358) & (!g1359) & (g1360) & (!g1361) & (!g677) & (!g726)) + ((g1358) & (!g1359) & (g1360) & (!g1361) & (!g677) & (g726)) + ((g1358) & (!g1359) & (g1360) & (g1361) & (!g677) & (!g726)) + ((g1358) & (!g1359) & (g1360) & (g1361) & (!g677) & (g726)) + ((g1358) & (!g1359) & (g1360) & (g1361) & (g677) & (g726)) + ((g1358) & (g1359) & (!g1360) & (!g1361) & (!g677) & (!g726)) + ((g1358) & (g1359) & (!g1360) & (!g1361) & (g677) & (!g726)) + ((g1358) & (g1359) & (!g1360) & (g1361) & (!g677) & (!g726)) + ((g1358) & (g1359) & (!g1360) & (g1361) & (g677) & (!g726)) + ((g1358) & (g1359) & (!g1360) & (g1361) & (g677) & (g726)) + ((g1358) & (g1359) & (g1360) & (!g1361) & (!g677) & (!g726)) + ((g1358) & (g1359) & (g1360) & (!g1361) & (!g677) & (g726)) + ((g1358) & (g1359) & (g1360) & (!g1361) & (g677) & (!g726)) + ((g1358) & (g1359) & (g1360) & (g1361) & (!g677) & (!g726)) + ((g1358) & (g1359) & (g1360) & (g1361) & (!g677) & (g726)) + ((g1358) & (g1359) & (g1360) & (g1361) & (g677) & (!g726)) + ((g1358) & (g1359) & (g1360) & (g1361) & (g677) & (g726)));
	assign g1941 = (((!g820) & (!g773) & (!g1937) & (g1938) & (!g1939) & (!g1940)) + ((!g820) & (!g773) & (!g1937) & (g1938) & (!g1939) & (g1940)) + ((!g820) & (!g773) & (!g1937) & (g1938) & (g1939) & (!g1940)) + ((!g820) & (!g773) & (!g1937) & (g1938) & (g1939) & (g1940)) + ((!g820) & (!g773) & (g1937) & (g1938) & (!g1939) & (!g1940)) + ((!g820) & (!g773) & (g1937) & (g1938) & (!g1939) & (g1940)) + ((!g820) & (!g773) & (g1937) & (g1938) & (g1939) & (!g1940)) + ((!g820) & (!g773) & (g1937) & (g1938) & (g1939) & (g1940)) + ((!g820) & (g773) & (!g1937) & (!g1938) & (!g1939) & (g1940)) + ((!g820) & (g773) & (!g1937) & (!g1938) & (g1939) & (g1940)) + ((!g820) & (g773) & (!g1937) & (g1938) & (!g1939) & (g1940)) + ((!g820) & (g773) & (!g1937) & (g1938) & (g1939) & (g1940)) + ((!g820) & (g773) & (g1937) & (!g1938) & (!g1939) & (g1940)) + ((!g820) & (g773) & (g1937) & (!g1938) & (g1939) & (g1940)) + ((!g820) & (g773) & (g1937) & (g1938) & (!g1939) & (g1940)) + ((!g820) & (g773) & (g1937) & (g1938) & (g1939) & (g1940)) + ((g820) & (!g773) & (g1937) & (!g1938) & (!g1939) & (!g1940)) + ((g820) & (!g773) & (g1937) & (!g1938) & (!g1939) & (g1940)) + ((g820) & (!g773) & (g1937) & (!g1938) & (g1939) & (!g1940)) + ((g820) & (!g773) & (g1937) & (!g1938) & (g1939) & (g1940)) + ((g820) & (!g773) & (g1937) & (g1938) & (!g1939) & (!g1940)) + ((g820) & (!g773) & (g1937) & (g1938) & (!g1939) & (g1940)) + ((g820) & (!g773) & (g1937) & (g1938) & (g1939) & (!g1940)) + ((g820) & (!g773) & (g1937) & (g1938) & (g1939) & (g1940)) + ((g820) & (g773) & (!g1937) & (!g1938) & (g1939) & (!g1940)) + ((g820) & (g773) & (!g1937) & (!g1938) & (g1939) & (g1940)) + ((g820) & (g773) & (!g1937) & (g1938) & (g1939) & (!g1940)) + ((g820) & (g773) & (!g1937) & (g1938) & (g1939) & (g1940)) + ((g820) & (g773) & (g1937) & (!g1938) & (g1939) & (!g1940)) + ((g820) & (g773) & (g1937) & (!g1938) & (g1939) & (g1940)) + ((g820) & (g773) & (g1937) & (g1938) & (g1939) & (!g1940)) + ((g820) & (g773) & (g1937) & (g1938) & (g1939) & (g1940)));
	assign g1942 = (((!g867) & (!sk[88]) & (!g1936) & (g1941)) + ((!g867) & (!sk[88]) & (g1936) & (!g1941)) + ((!g867) & (!sk[88]) & (g1936) & (g1941)) + ((!g867) & (sk[88]) & (!g1936) & (g1941)) + ((!g867) & (sk[88]) & (g1936) & (g1941)) + ((g867) & (!sk[88]) & (!g1936) & (g1941)) + ((g867) & (!sk[88]) & (g1936) & (!g1941)) + ((g867) & (!sk[88]) & (g1936) & (g1941)) + ((g867) & (sk[88]) & (g1936) & (!g1941)) + ((g867) & (sk[88]) & (g1936) & (g1941)));
	assign g1943 = (((!g1593) & (!g1605) & (!sk[89]) & (!g1733) & (g61)) + ((!g1593) & (!g1605) & (!sk[89]) & (g1733) & (!g61)) + ((!g1593) & (!g1605) & (!sk[89]) & (g1733) & (g61)) + ((!g1593) & (!g1605) & (sk[89]) & (g1733) & (!g61)) + ((!g1593) & (!g1605) & (sk[89]) & (g1733) & (g61)) + ((!g1593) & (g1605) & (!sk[89]) & (!g1733) & (!g61)) + ((!g1593) & (g1605) & (!sk[89]) & (!g1733) & (g61)) + ((!g1593) & (g1605) & (!sk[89]) & (g1733) & (!g61)) + ((!g1593) & (g1605) & (!sk[89]) & (g1733) & (g61)) + ((g1593) & (!g1605) & (!sk[89]) & (!g1733) & (g61)) + ((g1593) & (!g1605) & (!sk[89]) & (g1733) & (!g61)) + ((g1593) & (!g1605) & (!sk[89]) & (g1733) & (g61)) + ((g1593) & (!g1605) & (sk[89]) & (!g1733) & (g61)) + ((g1593) & (!g1605) & (sk[89]) & (g1733) & (g61)) + ((g1593) & (g1605) & (!sk[89]) & (!g1733) & (!g61)) + ((g1593) & (g1605) & (!sk[89]) & (!g1733) & (g61)) + ((g1593) & (g1605) & (!sk[89]) & (g1733) & (!g61)) + ((g1593) & (g1605) & (!sk[89]) & (g1733) & (g61)) + ((g1593) & (g1605) & (sk[89]) & (!g1733) & (g61)) + ((g1593) & (g1605) & (sk[89]) & (g1733) & (g61)));
	assign g1944 = (((!g132) & (!g1592) & (g1632) & (g1917) & (!g1942) & (!g1943)) + ((!g132) & (!g1592) & (g1632) & (g1917) & (!g1942) & (g1943)) + ((!g132) & (!g1592) & (g1632) & (g1917) & (g1942) & (!g1943)) + ((!g132) & (!g1592) & (g1632) & (g1917) & (g1942) & (g1943)) + ((!g132) & (g1592) & (!g1632) & (g1917) & (!g1942) & (g1943)) + ((!g132) & (g1592) & (!g1632) & (g1917) & (g1942) & (g1943)) + ((!g132) & (g1592) & (g1632) & (g1917) & (!g1942) & (g1943)) + ((!g132) & (g1592) & (g1632) & (g1917) & (g1942) & (g1943)) + ((g132) & (!g1592) & (!g1632) & (g1917) & (g1942) & (!g1943)) + ((g132) & (!g1592) & (!g1632) & (g1917) & (g1942) & (g1943)) + ((g132) & (!g1592) & (g1632) & (g1917) & (g1942) & (!g1943)) + ((g132) & (!g1592) & (g1632) & (g1917) & (g1942) & (g1943)) + ((g132) & (g1592) & (!g1632) & (g1917) & (g1942) & (!g1943)) + ((g132) & (g1592) & (!g1632) & (g1917) & (g1942) & (g1943)) + ((g132) & (g1592) & (g1632) & (g1917) & (g1942) & (!g1943)) + ((g132) & (g1592) & (g1632) & (g1917) & (g1942) & (g1943)));
	assign g1945 = (((!g1368) & (!g1369) & (!g1370) & (g1371) & (g820) & (g773)) + ((!g1368) & (!g1369) & (g1370) & (!g1371) & (!g820) & (g773)) + ((!g1368) & (!g1369) & (g1370) & (g1371) & (!g820) & (g773)) + ((!g1368) & (!g1369) & (g1370) & (g1371) & (g820) & (g773)) + ((!g1368) & (g1369) & (!g1370) & (!g1371) & (g820) & (!g773)) + ((!g1368) & (g1369) & (!g1370) & (g1371) & (g820) & (!g773)) + ((!g1368) & (g1369) & (!g1370) & (g1371) & (g820) & (g773)) + ((!g1368) & (g1369) & (g1370) & (!g1371) & (!g820) & (g773)) + ((!g1368) & (g1369) & (g1370) & (!g1371) & (g820) & (!g773)) + ((!g1368) & (g1369) & (g1370) & (g1371) & (!g820) & (g773)) + ((!g1368) & (g1369) & (g1370) & (g1371) & (g820) & (!g773)) + ((!g1368) & (g1369) & (g1370) & (g1371) & (g820) & (g773)) + ((g1368) & (!g1369) & (!g1370) & (!g1371) & (!g820) & (!g773)) + ((g1368) & (!g1369) & (!g1370) & (g1371) & (!g820) & (!g773)) + ((g1368) & (!g1369) & (!g1370) & (g1371) & (g820) & (g773)) + ((g1368) & (!g1369) & (g1370) & (!g1371) & (!g820) & (!g773)) + ((g1368) & (!g1369) & (g1370) & (!g1371) & (!g820) & (g773)) + ((g1368) & (!g1369) & (g1370) & (g1371) & (!g820) & (!g773)) + ((g1368) & (!g1369) & (g1370) & (g1371) & (!g820) & (g773)) + ((g1368) & (!g1369) & (g1370) & (g1371) & (g820) & (g773)) + ((g1368) & (g1369) & (!g1370) & (!g1371) & (!g820) & (!g773)) + ((g1368) & (g1369) & (!g1370) & (!g1371) & (g820) & (!g773)) + ((g1368) & (g1369) & (!g1370) & (g1371) & (!g820) & (!g773)) + ((g1368) & (g1369) & (!g1370) & (g1371) & (g820) & (!g773)) + ((g1368) & (g1369) & (!g1370) & (g1371) & (g820) & (g773)) + ((g1368) & (g1369) & (g1370) & (!g1371) & (!g820) & (!g773)) + ((g1368) & (g1369) & (g1370) & (!g1371) & (!g820) & (g773)) + ((g1368) & (g1369) & (g1370) & (!g1371) & (g820) & (!g773)) + ((g1368) & (g1369) & (g1370) & (g1371) & (!g820) & (!g773)) + ((g1368) & (g1369) & (g1370) & (g1371) & (!g820) & (g773)) + ((g1368) & (g1369) & (g1370) & (g1371) & (g820) & (!g773)) + ((g1368) & (g1369) & (g1370) & (g1371) & (g820) & (g773)));
	assign g1946 = (((!g1373) & (!g1374) & (!g1375) & (g1376) & (g820) & (g773)) + ((!g1373) & (!g1374) & (g1375) & (!g1376) & (!g820) & (g773)) + ((!g1373) & (!g1374) & (g1375) & (g1376) & (!g820) & (g773)) + ((!g1373) & (!g1374) & (g1375) & (g1376) & (g820) & (g773)) + ((!g1373) & (g1374) & (!g1375) & (!g1376) & (g820) & (!g773)) + ((!g1373) & (g1374) & (!g1375) & (g1376) & (g820) & (!g773)) + ((!g1373) & (g1374) & (!g1375) & (g1376) & (g820) & (g773)) + ((!g1373) & (g1374) & (g1375) & (!g1376) & (!g820) & (g773)) + ((!g1373) & (g1374) & (g1375) & (!g1376) & (g820) & (!g773)) + ((!g1373) & (g1374) & (g1375) & (g1376) & (!g820) & (g773)) + ((!g1373) & (g1374) & (g1375) & (g1376) & (g820) & (!g773)) + ((!g1373) & (g1374) & (g1375) & (g1376) & (g820) & (g773)) + ((g1373) & (!g1374) & (!g1375) & (!g1376) & (!g820) & (!g773)) + ((g1373) & (!g1374) & (!g1375) & (g1376) & (!g820) & (!g773)) + ((g1373) & (!g1374) & (!g1375) & (g1376) & (g820) & (g773)) + ((g1373) & (!g1374) & (g1375) & (!g1376) & (!g820) & (!g773)) + ((g1373) & (!g1374) & (g1375) & (!g1376) & (!g820) & (g773)) + ((g1373) & (!g1374) & (g1375) & (g1376) & (!g820) & (!g773)) + ((g1373) & (!g1374) & (g1375) & (g1376) & (!g820) & (g773)) + ((g1373) & (!g1374) & (g1375) & (g1376) & (g820) & (g773)) + ((g1373) & (g1374) & (!g1375) & (!g1376) & (!g820) & (!g773)) + ((g1373) & (g1374) & (!g1375) & (!g1376) & (g820) & (!g773)) + ((g1373) & (g1374) & (!g1375) & (g1376) & (!g820) & (!g773)) + ((g1373) & (g1374) & (!g1375) & (g1376) & (g820) & (!g773)) + ((g1373) & (g1374) & (!g1375) & (g1376) & (g820) & (g773)) + ((g1373) & (g1374) & (g1375) & (!g1376) & (!g820) & (!g773)) + ((g1373) & (g1374) & (g1375) & (!g1376) & (!g820) & (g773)) + ((g1373) & (g1374) & (g1375) & (!g1376) & (g820) & (!g773)) + ((g1373) & (g1374) & (g1375) & (g1376) & (!g820) & (!g773)) + ((g1373) & (g1374) & (g1375) & (g1376) & (!g820) & (g773)) + ((g1373) & (g1374) & (g1375) & (g1376) & (g820) & (!g773)) + ((g1373) & (g1374) & (g1375) & (g1376) & (g820) & (g773)));
	assign g1947 = (((!g1378) & (!g1379) & (!g1380) & (g1381) & (g820) & (g773)) + ((!g1378) & (!g1379) & (g1380) & (!g1381) & (!g820) & (g773)) + ((!g1378) & (!g1379) & (g1380) & (g1381) & (!g820) & (g773)) + ((!g1378) & (!g1379) & (g1380) & (g1381) & (g820) & (g773)) + ((!g1378) & (g1379) & (!g1380) & (!g1381) & (g820) & (!g773)) + ((!g1378) & (g1379) & (!g1380) & (g1381) & (g820) & (!g773)) + ((!g1378) & (g1379) & (!g1380) & (g1381) & (g820) & (g773)) + ((!g1378) & (g1379) & (g1380) & (!g1381) & (!g820) & (g773)) + ((!g1378) & (g1379) & (g1380) & (!g1381) & (g820) & (!g773)) + ((!g1378) & (g1379) & (g1380) & (g1381) & (!g820) & (g773)) + ((!g1378) & (g1379) & (g1380) & (g1381) & (g820) & (!g773)) + ((!g1378) & (g1379) & (g1380) & (g1381) & (g820) & (g773)) + ((g1378) & (!g1379) & (!g1380) & (!g1381) & (!g820) & (!g773)) + ((g1378) & (!g1379) & (!g1380) & (g1381) & (!g820) & (!g773)) + ((g1378) & (!g1379) & (!g1380) & (g1381) & (g820) & (g773)) + ((g1378) & (!g1379) & (g1380) & (!g1381) & (!g820) & (!g773)) + ((g1378) & (!g1379) & (g1380) & (!g1381) & (!g820) & (g773)) + ((g1378) & (!g1379) & (g1380) & (g1381) & (!g820) & (!g773)) + ((g1378) & (!g1379) & (g1380) & (g1381) & (!g820) & (g773)) + ((g1378) & (!g1379) & (g1380) & (g1381) & (g820) & (g773)) + ((g1378) & (g1379) & (!g1380) & (!g1381) & (!g820) & (!g773)) + ((g1378) & (g1379) & (!g1380) & (!g1381) & (g820) & (!g773)) + ((g1378) & (g1379) & (!g1380) & (g1381) & (!g820) & (!g773)) + ((g1378) & (g1379) & (!g1380) & (g1381) & (g820) & (!g773)) + ((g1378) & (g1379) & (!g1380) & (g1381) & (g820) & (g773)) + ((g1378) & (g1379) & (g1380) & (!g1381) & (!g820) & (!g773)) + ((g1378) & (g1379) & (g1380) & (!g1381) & (!g820) & (g773)) + ((g1378) & (g1379) & (g1380) & (!g1381) & (g820) & (!g773)) + ((g1378) & (g1379) & (g1380) & (g1381) & (!g820) & (!g773)) + ((g1378) & (g1379) & (g1380) & (g1381) & (!g820) & (g773)) + ((g1378) & (g1379) & (g1380) & (g1381) & (g820) & (!g773)) + ((g1378) & (g1379) & (g1380) & (g1381) & (g820) & (g773)));
	assign g1948 = (((!g1383) & (!g1384) & (!g1385) & (g1386) & (g820) & (g773)) + ((!g1383) & (!g1384) & (g1385) & (!g1386) & (!g820) & (g773)) + ((!g1383) & (!g1384) & (g1385) & (g1386) & (!g820) & (g773)) + ((!g1383) & (!g1384) & (g1385) & (g1386) & (g820) & (g773)) + ((!g1383) & (g1384) & (!g1385) & (!g1386) & (g820) & (!g773)) + ((!g1383) & (g1384) & (!g1385) & (g1386) & (g820) & (!g773)) + ((!g1383) & (g1384) & (!g1385) & (g1386) & (g820) & (g773)) + ((!g1383) & (g1384) & (g1385) & (!g1386) & (!g820) & (g773)) + ((!g1383) & (g1384) & (g1385) & (!g1386) & (g820) & (!g773)) + ((!g1383) & (g1384) & (g1385) & (g1386) & (!g820) & (g773)) + ((!g1383) & (g1384) & (g1385) & (g1386) & (g820) & (!g773)) + ((!g1383) & (g1384) & (g1385) & (g1386) & (g820) & (g773)) + ((g1383) & (!g1384) & (!g1385) & (!g1386) & (!g820) & (!g773)) + ((g1383) & (!g1384) & (!g1385) & (g1386) & (!g820) & (!g773)) + ((g1383) & (!g1384) & (!g1385) & (g1386) & (g820) & (g773)) + ((g1383) & (!g1384) & (g1385) & (!g1386) & (!g820) & (!g773)) + ((g1383) & (!g1384) & (g1385) & (!g1386) & (!g820) & (g773)) + ((g1383) & (!g1384) & (g1385) & (g1386) & (!g820) & (!g773)) + ((g1383) & (!g1384) & (g1385) & (g1386) & (!g820) & (g773)) + ((g1383) & (!g1384) & (g1385) & (g1386) & (g820) & (g773)) + ((g1383) & (g1384) & (!g1385) & (!g1386) & (!g820) & (!g773)) + ((g1383) & (g1384) & (!g1385) & (!g1386) & (g820) & (!g773)) + ((g1383) & (g1384) & (!g1385) & (g1386) & (!g820) & (!g773)) + ((g1383) & (g1384) & (!g1385) & (g1386) & (g820) & (!g773)) + ((g1383) & (g1384) & (!g1385) & (g1386) & (g820) & (g773)) + ((g1383) & (g1384) & (g1385) & (!g1386) & (!g820) & (!g773)) + ((g1383) & (g1384) & (g1385) & (!g1386) & (!g820) & (g773)) + ((g1383) & (g1384) & (g1385) & (!g1386) & (g820) & (!g773)) + ((g1383) & (g1384) & (g1385) & (g1386) & (!g820) & (!g773)) + ((g1383) & (g1384) & (g1385) & (g1386) & (!g820) & (g773)) + ((g1383) & (g1384) & (g1385) & (g1386) & (g820) & (!g773)) + ((g1383) & (g1384) & (g1385) & (g1386) & (g820) & (g773)));
	assign g1949 = (((!g1945) & (!g1946) & (!g1947) & (g1948) & (g677) & (g726)) + ((!g1945) & (!g1946) & (g1947) & (!g1948) & (!g677) & (g726)) + ((!g1945) & (!g1946) & (g1947) & (g1948) & (!g677) & (g726)) + ((!g1945) & (!g1946) & (g1947) & (g1948) & (g677) & (g726)) + ((!g1945) & (g1946) & (!g1947) & (!g1948) & (g677) & (!g726)) + ((!g1945) & (g1946) & (!g1947) & (g1948) & (g677) & (!g726)) + ((!g1945) & (g1946) & (!g1947) & (g1948) & (g677) & (g726)) + ((!g1945) & (g1946) & (g1947) & (!g1948) & (!g677) & (g726)) + ((!g1945) & (g1946) & (g1947) & (!g1948) & (g677) & (!g726)) + ((!g1945) & (g1946) & (g1947) & (g1948) & (!g677) & (g726)) + ((!g1945) & (g1946) & (g1947) & (g1948) & (g677) & (!g726)) + ((!g1945) & (g1946) & (g1947) & (g1948) & (g677) & (g726)) + ((g1945) & (!g1946) & (!g1947) & (!g1948) & (!g677) & (!g726)) + ((g1945) & (!g1946) & (!g1947) & (g1948) & (!g677) & (!g726)) + ((g1945) & (!g1946) & (!g1947) & (g1948) & (g677) & (g726)) + ((g1945) & (!g1946) & (g1947) & (!g1948) & (!g677) & (!g726)) + ((g1945) & (!g1946) & (g1947) & (!g1948) & (!g677) & (g726)) + ((g1945) & (!g1946) & (g1947) & (g1948) & (!g677) & (!g726)) + ((g1945) & (!g1946) & (g1947) & (g1948) & (!g677) & (g726)) + ((g1945) & (!g1946) & (g1947) & (g1948) & (g677) & (g726)) + ((g1945) & (g1946) & (!g1947) & (!g1948) & (!g677) & (!g726)) + ((g1945) & (g1946) & (!g1947) & (!g1948) & (g677) & (!g726)) + ((g1945) & (g1946) & (!g1947) & (g1948) & (!g677) & (!g726)) + ((g1945) & (g1946) & (!g1947) & (g1948) & (g677) & (!g726)) + ((g1945) & (g1946) & (!g1947) & (g1948) & (g677) & (g726)) + ((g1945) & (g1946) & (g1947) & (!g1948) & (!g677) & (!g726)) + ((g1945) & (g1946) & (g1947) & (!g1948) & (!g677) & (g726)) + ((g1945) & (g1946) & (g1947) & (!g1948) & (g677) & (!g726)) + ((g1945) & (g1946) & (g1947) & (g1948) & (!g677) & (!g726)) + ((g1945) & (g1946) & (g1947) & (g1948) & (!g677) & (g726)) + ((g1945) & (g1946) & (g1947) & (g1948) & (g677) & (!g726)) + ((g1945) & (g1946) & (g1947) & (g1948) & (g677) & (g726)));
	assign g1950 = (((!g1389) & (!g1390) & (!g1391) & (g1392) & (g677) & (g726)) + ((!g1389) & (!g1390) & (g1391) & (!g1392) & (!g677) & (g726)) + ((!g1389) & (!g1390) & (g1391) & (g1392) & (!g677) & (g726)) + ((!g1389) & (!g1390) & (g1391) & (g1392) & (g677) & (g726)) + ((!g1389) & (g1390) & (!g1391) & (!g1392) & (g677) & (!g726)) + ((!g1389) & (g1390) & (!g1391) & (g1392) & (g677) & (!g726)) + ((!g1389) & (g1390) & (!g1391) & (g1392) & (g677) & (g726)) + ((!g1389) & (g1390) & (g1391) & (!g1392) & (!g677) & (g726)) + ((!g1389) & (g1390) & (g1391) & (!g1392) & (g677) & (!g726)) + ((!g1389) & (g1390) & (g1391) & (g1392) & (!g677) & (g726)) + ((!g1389) & (g1390) & (g1391) & (g1392) & (g677) & (!g726)) + ((!g1389) & (g1390) & (g1391) & (g1392) & (g677) & (g726)) + ((g1389) & (!g1390) & (!g1391) & (!g1392) & (!g677) & (!g726)) + ((g1389) & (!g1390) & (!g1391) & (g1392) & (!g677) & (!g726)) + ((g1389) & (!g1390) & (!g1391) & (g1392) & (g677) & (g726)) + ((g1389) & (!g1390) & (g1391) & (!g1392) & (!g677) & (!g726)) + ((g1389) & (!g1390) & (g1391) & (!g1392) & (!g677) & (g726)) + ((g1389) & (!g1390) & (g1391) & (g1392) & (!g677) & (!g726)) + ((g1389) & (!g1390) & (g1391) & (g1392) & (!g677) & (g726)) + ((g1389) & (!g1390) & (g1391) & (g1392) & (g677) & (g726)) + ((g1389) & (g1390) & (!g1391) & (!g1392) & (!g677) & (!g726)) + ((g1389) & (g1390) & (!g1391) & (!g1392) & (g677) & (!g726)) + ((g1389) & (g1390) & (!g1391) & (g1392) & (!g677) & (!g726)) + ((g1389) & (g1390) & (!g1391) & (g1392) & (g677) & (!g726)) + ((g1389) & (g1390) & (!g1391) & (g1392) & (g677) & (g726)) + ((g1389) & (g1390) & (g1391) & (!g1392) & (!g677) & (!g726)) + ((g1389) & (g1390) & (g1391) & (!g1392) & (!g677) & (g726)) + ((g1389) & (g1390) & (g1391) & (!g1392) & (g677) & (!g726)) + ((g1389) & (g1390) & (g1391) & (g1392) & (!g677) & (!g726)) + ((g1389) & (g1390) & (g1391) & (g1392) & (!g677) & (g726)) + ((g1389) & (g1390) & (g1391) & (g1392) & (g677) & (!g726)) + ((g1389) & (g1390) & (g1391) & (g1392) & (g677) & (g726)));
	assign g1951 = (((!g677) & (!g726) & (!g1394) & (g1395) & (!sk[97]) & (!g1396)) + ((!g677) & (!g726) & (!g1394) & (g1395) & (!sk[97]) & (g1396)) + ((!g677) & (!g726) & (g1394) & (!g1395) & (!sk[97]) & (!g1396)) + ((!g677) & (!g726) & (g1394) & (!g1395) & (!sk[97]) & (g1396)) + ((!g677) & (!g726) & (g1394) & (g1395) & (!sk[97]) & (!g1396)) + ((!g677) & (!g726) & (g1394) & (g1395) & (!sk[97]) & (g1396)) + ((!g677) & (g726) & (!g1394) & (!g1395) & (!sk[97]) & (!g1396)) + ((!g677) & (g726) & (!g1394) & (!g1395) & (!sk[97]) & (g1396)) + ((!g677) & (g726) & (!g1394) & (!g1395) & (sk[97]) & (g1396)) + ((!g677) & (g726) & (!g1394) & (g1395) & (!sk[97]) & (!g1396)) + ((!g677) & (g726) & (!g1394) & (g1395) & (!sk[97]) & (g1396)) + ((!g677) & (g726) & (!g1394) & (g1395) & (sk[97]) & (g1396)) + ((!g677) & (g726) & (g1394) & (!g1395) & (!sk[97]) & (!g1396)) + ((!g677) & (g726) & (g1394) & (!g1395) & (!sk[97]) & (g1396)) + ((!g677) & (g726) & (g1394) & (!g1395) & (sk[97]) & (g1396)) + ((!g677) & (g726) & (g1394) & (g1395) & (!sk[97]) & (!g1396)) + ((!g677) & (g726) & (g1394) & (g1395) & (!sk[97]) & (g1396)) + ((!g677) & (g726) & (g1394) & (g1395) & (sk[97]) & (g1396)) + ((g677) & (!g726) & (!g1394) & (g1395) & (!sk[97]) & (!g1396)) + ((g677) & (!g726) & (!g1394) & (g1395) & (!sk[97]) & (g1396)) + ((g677) & (!g726) & (g1394) & (!g1395) & (!sk[97]) & (!g1396)) + ((g677) & (!g726) & (g1394) & (!g1395) & (!sk[97]) & (g1396)) + ((g677) & (!g726) & (g1394) & (!g1395) & (sk[97]) & (!g1396)) + ((g677) & (!g726) & (g1394) & (!g1395) & (sk[97]) & (g1396)) + ((g677) & (!g726) & (g1394) & (g1395) & (!sk[97]) & (!g1396)) + ((g677) & (!g726) & (g1394) & (g1395) & (!sk[97]) & (g1396)) + ((g677) & (!g726) & (g1394) & (g1395) & (sk[97]) & (!g1396)) + ((g677) & (!g726) & (g1394) & (g1395) & (sk[97]) & (g1396)) + ((g677) & (g726) & (!g1394) & (!g1395) & (!sk[97]) & (!g1396)) + ((g677) & (g726) & (!g1394) & (!g1395) & (!sk[97]) & (g1396)) + ((g677) & (g726) & (!g1394) & (g1395) & (!sk[97]) & (!g1396)) + ((g677) & (g726) & (!g1394) & (g1395) & (!sk[97]) & (g1396)) + ((g677) & (g726) & (!g1394) & (g1395) & (sk[97]) & (!g1396)) + ((g677) & (g726) & (!g1394) & (g1395) & (sk[97]) & (g1396)) + ((g677) & (g726) & (g1394) & (!g1395) & (!sk[97]) & (!g1396)) + ((g677) & (g726) & (g1394) & (!g1395) & (!sk[97]) & (g1396)) + ((g677) & (g726) & (g1394) & (g1395) & (!sk[97]) & (!g1396)) + ((g677) & (g726) & (g1394) & (g1395) & (!sk[97]) & (g1396)) + ((g677) & (g726) & (g1394) & (g1395) & (sk[97]) & (!g1396)) + ((g677) & (g726) & (g1394) & (g1395) & (sk[97]) & (g1396)));
	assign g1952 = (((!g1398) & (!g1399) & (!g1400) & (g1401) & (g677) & (g726)) + ((!g1398) & (!g1399) & (g1400) & (!g1401) & (!g677) & (g726)) + ((!g1398) & (!g1399) & (g1400) & (g1401) & (!g677) & (g726)) + ((!g1398) & (!g1399) & (g1400) & (g1401) & (g677) & (g726)) + ((!g1398) & (g1399) & (!g1400) & (!g1401) & (g677) & (!g726)) + ((!g1398) & (g1399) & (!g1400) & (g1401) & (g677) & (!g726)) + ((!g1398) & (g1399) & (!g1400) & (g1401) & (g677) & (g726)) + ((!g1398) & (g1399) & (g1400) & (!g1401) & (!g677) & (g726)) + ((!g1398) & (g1399) & (g1400) & (!g1401) & (g677) & (!g726)) + ((!g1398) & (g1399) & (g1400) & (g1401) & (!g677) & (g726)) + ((!g1398) & (g1399) & (g1400) & (g1401) & (g677) & (!g726)) + ((!g1398) & (g1399) & (g1400) & (g1401) & (g677) & (g726)) + ((g1398) & (!g1399) & (!g1400) & (!g1401) & (!g677) & (!g726)) + ((g1398) & (!g1399) & (!g1400) & (g1401) & (!g677) & (!g726)) + ((g1398) & (!g1399) & (!g1400) & (g1401) & (g677) & (g726)) + ((g1398) & (!g1399) & (g1400) & (!g1401) & (!g677) & (!g726)) + ((g1398) & (!g1399) & (g1400) & (!g1401) & (!g677) & (g726)) + ((g1398) & (!g1399) & (g1400) & (g1401) & (!g677) & (!g726)) + ((g1398) & (!g1399) & (g1400) & (g1401) & (!g677) & (g726)) + ((g1398) & (!g1399) & (g1400) & (g1401) & (g677) & (g726)) + ((g1398) & (g1399) & (!g1400) & (!g1401) & (!g677) & (!g726)) + ((g1398) & (g1399) & (!g1400) & (!g1401) & (g677) & (!g726)) + ((g1398) & (g1399) & (!g1400) & (g1401) & (!g677) & (!g726)) + ((g1398) & (g1399) & (!g1400) & (g1401) & (g677) & (!g726)) + ((g1398) & (g1399) & (!g1400) & (g1401) & (g677) & (g726)) + ((g1398) & (g1399) & (g1400) & (!g1401) & (!g677) & (!g726)) + ((g1398) & (g1399) & (g1400) & (!g1401) & (!g677) & (g726)) + ((g1398) & (g1399) & (g1400) & (!g1401) & (g677) & (!g726)) + ((g1398) & (g1399) & (g1400) & (g1401) & (!g677) & (!g726)) + ((g1398) & (g1399) & (g1400) & (g1401) & (!g677) & (g726)) + ((g1398) & (g1399) & (g1400) & (g1401) & (g677) & (!g726)) + ((g1398) & (g1399) & (g1400) & (g1401) & (g677) & (g726)));
	assign g1953 = (((!g1403) & (!g1404) & (!g1405) & (g1406) & (g677) & (g726)) + ((!g1403) & (!g1404) & (g1405) & (!g1406) & (!g677) & (g726)) + ((!g1403) & (!g1404) & (g1405) & (g1406) & (!g677) & (g726)) + ((!g1403) & (!g1404) & (g1405) & (g1406) & (g677) & (g726)) + ((!g1403) & (g1404) & (!g1405) & (!g1406) & (g677) & (!g726)) + ((!g1403) & (g1404) & (!g1405) & (g1406) & (g677) & (!g726)) + ((!g1403) & (g1404) & (!g1405) & (g1406) & (g677) & (g726)) + ((!g1403) & (g1404) & (g1405) & (!g1406) & (!g677) & (g726)) + ((!g1403) & (g1404) & (g1405) & (!g1406) & (g677) & (!g726)) + ((!g1403) & (g1404) & (g1405) & (g1406) & (!g677) & (g726)) + ((!g1403) & (g1404) & (g1405) & (g1406) & (g677) & (!g726)) + ((!g1403) & (g1404) & (g1405) & (g1406) & (g677) & (g726)) + ((g1403) & (!g1404) & (!g1405) & (!g1406) & (!g677) & (!g726)) + ((g1403) & (!g1404) & (!g1405) & (g1406) & (!g677) & (!g726)) + ((g1403) & (!g1404) & (!g1405) & (g1406) & (g677) & (g726)) + ((g1403) & (!g1404) & (g1405) & (!g1406) & (!g677) & (!g726)) + ((g1403) & (!g1404) & (g1405) & (!g1406) & (!g677) & (g726)) + ((g1403) & (!g1404) & (g1405) & (g1406) & (!g677) & (!g726)) + ((g1403) & (!g1404) & (g1405) & (g1406) & (!g677) & (g726)) + ((g1403) & (!g1404) & (g1405) & (g1406) & (g677) & (g726)) + ((g1403) & (g1404) & (!g1405) & (!g1406) & (!g677) & (!g726)) + ((g1403) & (g1404) & (!g1405) & (!g1406) & (g677) & (!g726)) + ((g1403) & (g1404) & (!g1405) & (g1406) & (!g677) & (!g726)) + ((g1403) & (g1404) & (!g1405) & (g1406) & (g677) & (!g726)) + ((g1403) & (g1404) & (!g1405) & (g1406) & (g677) & (g726)) + ((g1403) & (g1404) & (g1405) & (!g1406) & (!g677) & (!g726)) + ((g1403) & (g1404) & (g1405) & (!g1406) & (!g677) & (g726)) + ((g1403) & (g1404) & (g1405) & (!g1406) & (g677) & (!g726)) + ((g1403) & (g1404) & (g1405) & (g1406) & (!g677) & (!g726)) + ((g1403) & (g1404) & (g1405) & (g1406) & (!g677) & (g726)) + ((g1403) & (g1404) & (g1405) & (g1406) & (g677) & (!g726)) + ((g1403) & (g1404) & (g1405) & (g1406) & (g677) & (g726)));
	assign g1954 = (((!g820) & (!g773) & (!g1950) & (g1951) & (!g1952) & (!g1953)) + ((!g820) & (!g773) & (!g1950) & (g1951) & (!g1952) & (g1953)) + ((!g820) & (!g773) & (!g1950) & (g1951) & (g1952) & (!g1953)) + ((!g820) & (!g773) & (!g1950) & (g1951) & (g1952) & (g1953)) + ((!g820) & (!g773) & (g1950) & (g1951) & (!g1952) & (!g1953)) + ((!g820) & (!g773) & (g1950) & (g1951) & (!g1952) & (g1953)) + ((!g820) & (!g773) & (g1950) & (g1951) & (g1952) & (!g1953)) + ((!g820) & (!g773) & (g1950) & (g1951) & (g1952) & (g1953)) + ((!g820) & (g773) & (!g1950) & (!g1951) & (!g1952) & (g1953)) + ((!g820) & (g773) & (!g1950) & (!g1951) & (g1952) & (g1953)) + ((!g820) & (g773) & (!g1950) & (g1951) & (!g1952) & (g1953)) + ((!g820) & (g773) & (!g1950) & (g1951) & (g1952) & (g1953)) + ((!g820) & (g773) & (g1950) & (!g1951) & (!g1952) & (g1953)) + ((!g820) & (g773) & (g1950) & (!g1951) & (g1952) & (g1953)) + ((!g820) & (g773) & (g1950) & (g1951) & (!g1952) & (g1953)) + ((!g820) & (g773) & (g1950) & (g1951) & (g1952) & (g1953)) + ((g820) & (!g773) & (g1950) & (!g1951) & (!g1952) & (!g1953)) + ((g820) & (!g773) & (g1950) & (!g1951) & (!g1952) & (g1953)) + ((g820) & (!g773) & (g1950) & (!g1951) & (g1952) & (!g1953)) + ((g820) & (!g773) & (g1950) & (!g1951) & (g1952) & (g1953)) + ((g820) & (!g773) & (g1950) & (g1951) & (!g1952) & (!g1953)) + ((g820) & (!g773) & (g1950) & (g1951) & (!g1952) & (g1953)) + ((g820) & (!g773) & (g1950) & (g1951) & (g1952) & (!g1953)) + ((g820) & (!g773) & (g1950) & (g1951) & (g1952) & (g1953)) + ((g820) & (g773) & (!g1950) & (!g1951) & (g1952) & (!g1953)) + ((g820) & (g773) & (!g1950) & (!g1951) & (g1952) & (g1953)) + ((g820) & (g773) & (!g1950) & (g1951) & (g1952) & (!g1953)) + ((g820) & (g773) & (!g1950) & (g1951) & (g1952) & (g1953)) + ((g820) & (g773) & (g1950) & (!g1951) & (g1952) & (!g1953)) + ((g820) & (g773) & (g1950) & (!g1951) & (g1952) & (g1953)) + ((g820) & (g773) & (g1950) & (g1951) & (g1952) & (!g1953)) + ((g820) & (g773) & (g1950) & (g1951) & (g1952) & (g1953)));
	assign g1955 = (((!sk[101]) & (!g867) & (!g1949) & (g1954)) + ((!sk[101]) & (!g867) & (g1949) & (!g1954)) + ((!sk[101]) & (!g867) & (g1949) & (g1954)) + ((!sk[101]) & (g867) & (!g1949) & (g1954)) + ((!sk[101]) & (g867) & (g1949) & (!g1954)) + ((!sk[101]) & (g867) & (g1949) & (g1954)) + ((sk[101]) & (!g867) & (!g1949) & (g1954)) + ((sk[101]) & (!g867) & (g1949) & (g1954)) + ((sk[101]) & (g867) & (g1949) & (!g1954)) + ((sk[101]) & (g867) & (g1949) & (g1954)));
	assign g1956 = (((!g1593) & (!g1605) & (!g1746) & (!sk[102]) & (g62)) + ((!g1593) & (!g1605) & (g1746) & (!sk[102]) & (!g62)) + ((!g1593) & (!g1605) & (g1746) & (!sk[102]) & (g62)) + ((!g1593) & (!g1605) & (g1746) & (sk[102]) & (!g62)) + ((!g1593) & (!g1605) & (g1746) & (sk[102]) & (g62)) + ((!g1593) & (g1605) & (!g1746) & (!sk[102]) & (!g62)) + ((!g1593) & (g1605) & (!g1746) & (!sk[102]) & (g62)) + ((!g1593) & (g1605) & (g1746) & (!sk[102]) & (!g62)) + ((!g1593) & (g1605) & (g1746) & (!sk[102]) & (g62)) + ((g1593) & (!g1605) & (!g1746) & (!sk[102]) & (g62)) + ((g1593) & (!g1605) & (!g1746) & (sk[102]) & (g62)) + ((g1593) & (!g1605) & (g1746) & (!sk[102]) & (!g62)) + ((g1593) & (!g1605) & (g1746) & (!sk[102]) & (g62)) + ((g1593) & (!g1605) & (g1746) & (sk[102]) & (g62)) + ((g1593) & (g1605) & (!g1746) & (!sk[102]) & (!g62)) + ((g1593) & (g1605) & (!g1746) & (!sk[102]) & (g62)) + ((g1593) & (g1605) & (!g1746) & (sk[102]) & (g62)) + ((g1593) & (g1605) & (g1746) & (!sk[102]) & (!g62)) + ((g1593) & (g1605) & (g1746) & (!sk[102]) & (g62)) + ((g1593) & (g1605) & (g1746) & (sk[102]) & (g62)));
	assign g1957 = (((!g132) & (!g1592) & (g1644) & (g1917) & (!g1955) & (!g1956)) + ((!g132) & (!g1592) & (g1644) & (g1917) & (!g1955) & (g1956)) + ((!g132) & (!g1592) & (g1644) & (g1917) & (g1955) & (!g1956)) + ((!g132) & (!g1592) & (g1644) & (g1917) & (g1955) & (g1956)) + ((!g132) & (g1592) & (!g1644) & (g1917) & (!g1955) & (g1956)) + ((!g132) & (g1592) & (!g1644) & (g1917) & (g1955) & (g1956)) + ((!g132) & (g1592) & (g1644) & (g1917) & (!g1955) & (g1956)) + ((!g132) & (g1592) & (g1644) & (g1917) & (g1955) & (g1956)) + ((g132) & (!g1592) & (!g1644) & (g1917) & (g1955) & (!g1956)) + ((g132) & (!g1592) & (!g1644) & (g1917) & (g1955) & (g1956)) + ((g132) & (!g1592) & (g1644) & (g1917) & (g1955) & (!g1956)) + ((g132) & (!g1592) & (g1644) & (g1917) & (g1955) & (g1956)) + ((g132) & (g1592) & (!g1644) & (g1917) & (g1955) & (!g1956)) + ((g132) & (g1592) & (!g1644) & (g1917) & (g1955) & (g1956)) + ((g132) & (g1592) & (g1644) & (g1917) & (g1955) & (!g1956)) + ((g132) & (g1592) & (g1644) & (g1917) & (g1955) & (g1956)));
	assign g1958 = (((!g1413) & (!g1418) & (!g1423) & (g1428) & (g677) & (g726)) + ((!g1413) & (!g1418) & (g1423) & (!g1428) & (!g677) & (g726)) + ((!g1413) & (!g1418) & (g1423) & (g1428) & (!g677) & (g726)) + ((!g1413) & (!g1418) & (g1423) & (g1428) & (g677) & (g726)) + ((!g1413) & (g1418) & (!g1423) & (!g1428) & (g677) & (!g726)) + ((!g1413) & (g1418) & (!g1423) & (g1428) & (g677) & (!g726)) + ((!g1413) & (g1418) & (!g1423) & (g1428) & (g677) & (g726)) + ((!g1413) & (g1418) & (g1423) & (!g1428) & (!g677) & (g726)) + ((!g1413) & (g1418) & (g1423) & (!g1428) & (g677) & (!g726)) + ((!g1413) & (g1418) & (g1423) & (g1428) & (!g677) & (g726)) + ((!g1413) & (g1418) & (g1423) & (g1428) & (g677) & (!g726)) + ((!g1413) & (g1418) & (g1423) & (g1428) & (g677) & (g726)) + ((g1413) & (!g1418) & (!g1423) & (!g1428) & (!g677) & (!g726)) + ((g1413) & (!g1418) & (!g1423) & (g1428) & (!g677) & (!g726)) + ((g1413) & (!g1418) & (!g1423) & (g1428) & (g677) & (g726)) + ((g1413) & (!g1418) & (g1423) & (!g1428) & (!g677) & (!g726)) + ((g1413) & (!g1418) & (g1423) & (!g1428) & (!g677) & (g726)) + ((g1413) & (!g1418) & (g1423) & (g1428) & (!g677) & (!g726)) + ((g1413) & (!g1418) & (g1423) & (g1428) & (!g677) & (g726)) + ((g1413) & (!g1418) & (g1423) & (g1428) & (g677) & (g726)) + ((g1413) & (g1418) & (!g1423) & (!g1428) & (!g677) & (!g726)) + ((g1413) & (g1418) & (!g1423) & (!g1428) & (g677) & (!g726)) + ((g1413) & (g1418) & (!g1423) & (g1428) & (!g677) & (!g726)) + ((g1413) & (g1418) & (!g1423) & (g1428) & (g677) & (!g726)) + ((g1413) & (g1418) & (!g1423) & (g1428) & (g677) & (g726)) + ((g1413) & (g1418) & (g1423) & (!g1428) & (!g677) & (!g726)) + ((g1413) & (g1418) & (g1423) & (!g1428) & (!g677) & (g726)) + ((g1413) & (g1418) & (g1423) & (!g1428) & (g677) & (!g726)) + ((g1413) & (g1418) & (g1423) & (g1428) & (!g677) & (!g726)) + ((g1413) & (g1418) & (g1423) & (g1428) & (!g677) & (g726)) + ((g1413) & (g1418) & (g1423) & (g1428) & (g677) & (!g726)) + ((g1413) & (g1418) & (g1423) & (g1428) & (g677) & (g726)));
	assign g1959 = (((!g1414) & (!g1419) & (!g1424) & (g1429) & (g677) & (g726)) + ((!g1414) & (!g1419) & (g1424) & (!g1429) & (!g677) & (g726)) + ((!g1414) & (!g1419) & (g1424) & (g1429) & (!g677) & (g726)) + ((!g1414) & (!g1419) & (g1424) & (g1429) & (g677) & (g726)) + ((!g1414) & (g1419) & (!g1424) & (!g1429) & (g677) & (!g726)) + ((!g1414) & (g1419) & (!g1424) & (g1429) & (g677) & (!g726)) + ((!g1414) & (g1419) & (!g1424) & (g1429) & (g677) & (g726)) + ((!g1414) & (g1419) & (g1424) & (!g1429) & (!g677) & (g726)) + ((!g1414) & (g1419) & (g1424) & (!g1429) & (g677) & (!g726)) + ((!g1414) & (g1419) & (g1424) & (g1429) & (!g677) & (g726)) + ((!g1414) & (g1419) & (g1424) & (g1429) & (g677) & (!g726)) + ((!g1414) & (g1419) & (g1424) & (g1429) & (g677) & (g726)) + ((g1414) & (!g1419) & (!g1424) & (!g1429) & (!g677) & (!g726)) + ((g1414) & (!g1419) & (!g1424) & (g1429) & (!g677) & (!g726)) + ((g1414) & (!g1419) & (!g1424) & (g1429) & (g677) & (g726)) + ((g1414) & (!g1419) & (g1424) & (!g1429) & (!g677) & (!g726)) + ((g1414) & (!g1419) & (g1424) & (!g1429) & (!g677) & (g726)) + ((g1414) & (!g1419) & (g1424) & (g1429) & (!g677) & (!g726)) + ((g1414) & (!g1419) & (g1424) & (g1429) & (!g677) & (g726)) + ((g1414) & (!g1419) & (g1424) & (g1429) & (g677) & (g726)) + ((g1414) & (g1419) & (!g1424) & (!g1429) & (!g677) & (!g726)) + ((g1414) & (g1419) & (!g1424) & (!g1429) & (g677) & (!g726)) + ((g1414) & (g1419) & (!g1424) & (g1429) & (!g677) & (!g726)) + ((g1414) & (g1419) & (!g1424) & (g1429) & (g677) & (!g726)) + ((g1414) & (g1419) & (!g1424) & (g1429) & (g677) & (g726)) + ((g1414) & (g1419) & (g1424) & (!g1429) & (!g677) & (!g726)) + ((g1414) & (g1419) & (g1424) & (!g1429) & (!g677) & (g726)) + ((g1414) & (g1419) & (g1424) & (!g1429) & (g677) & (!g726)) + ((g1414) & (g1419) & (g1424) & (g1429) & (!g677) & (!g726)) + ((g1414) & (g1419) & (g1424) & (g1429) & (!g677) & (g726)) + ((g1414) & (g1419) & (g1424) & (g1429) & (g677) & (!g726)) + ((g1414) & (g1419) & (g1424) & (g1429) & (g677) & (g726)));
	assign g1960 = (((!g1415) & (!g1420) & (!g1425) & (g1430) & (g677) & (g726)) + ((!g1415) & (!g1420) & (g1425) & (!g1430) & (!g677) & (g726)) + ((!g1415) & (!g1420) & (g1425) & (g1430) & (!g677) & (g726)) + ((!g1415) & (!g1420) & (g1425) & (g1430) & (g677) & (g726)) + ((!g1415) & (g1420) & (!g1425) & (!g1430) & (g677) & (!g726)) + ((!g1415) & (g1420) & (!g1425) & (g1430) & (g677) & (!g726)) + ((!g1415) & (g1420) & (!g1425) & (g1430) & (g677) & (g726)) + ((!g1415) & (g1420) & (g1425) & (!g1430) & (!g677) & (g726)) + ((!g1415) & (g1420) & (g1425) & (!g1430) & (g677) & (!g726)) + ((!g1415) & (g1420) & (g1425) & (g1430) & (!g677) & (g726)) + ((!g1415) & (g1420) & (g1425) & (g1430) & (g677) & (!g726)) + ((!g1415) & (g1420) & (g1425) & (g1430) & (g677) & (g726)) + ((g1415) & (!g1420) & (!g1425) & (!g1430) & (!g677) & (!g726)) + ((g1415) & (!g1420) & (!g1425) & (g1430) & (!g677) & (!g726)) + ((g1415) & (!g1420) & (!g1425) & (g1430) & (g677) & (g726)) + ((g1415) & (!g1420) & (g1425) & (!g1430) & (!g677) & (!g726)) + ((g1415) & (!g1420) & (g1425) & (!g1430) & (!g677) & (g726)) + ((g1415) & (!g1420) & (g1425) & (g1430) & (!g677) & (!g726)) + ((g1415) & (!g1420) & (g1425) & (g1430) & (!g677) & (g726)) + ((g1415) & (!g1420) & (g1425) & (g1430) & (g677) & (g726)) + ((g1415) & (g1420) & (!g1425) & (!g1430) & (!g677) & (!g726)) + ((g1415) & (g1420) & (!g1425) & (!g1430) & (g677) & (!g726)) + ((g1415) & (g1420) & (!g1425) & (g1430) & (!g677) & (!g726)) + ((g1415) & (g1420) & (!g1425) & (g1430) & (g677) & (!g726)) + ((g1415) & (g1420) & (!g1425) & (g1430) & (g677) & (g726)) + ((g1415) & (g1420) & (g1425) & (!g1430) & (!g677) & (!g726)) + ((g1415) & (g1420) & (g1425) & (!g1430) & (!g677) & (g726)) + ((g1415) & (g1420) & (g1425) & (!g1430) & (g677) & (!g726)) + ((g1415) & (g1420) & (g1425) & (g1430) & (!g677) & (!g726)) + ((g1415) & (g1420) & (g1425) & (g1430) & (!g677) & (g726)) + ((g1415) & (g1420) & (g1425) & (g1430) & (g677) & (!g726)) + ((g1415) & (g1420) & (g1425) & (g1430) & (g677) & (g726)));
	assign g1961 = (((!g1416) & (!g1421) & (!g1426) & (g1431) & (g677) & (g726)) + ((!g1416) & (!g1421) & (g1426) & (!g1431) & (!g677) & (g726)) + ((!g1416) & (!g1421) & (g1426) & (g1431) & (!g677) & (g726)) + ((!g1416) & (!g1421) & (g1426) & (g1431) & (g677) & (g726)) + ((!g1416) & (g1421) & (!g1426) & (!g1431) & (g677) & (!g726)) + ((!g1416) & (g1421) & (!g1426) & (g1431) & (g677) & (!g726)) + ((!g1416) & (g1421) & (!g1426) & (g1431) & (g677) & (g726)) + ((!g1416) & (g1421) & (g1426) & (!g1431) & (!g677) & (g726)) + ((!g1416) & (g1421) & (g1426) & (!g1431) & (g677) & (!g726)) + ((!g1416) & (g1421) & (g1426) & (g1431) & (!g677) & (g726)) + ((!g1416) & (g1421) & (g1426) & (g1431) & (g677) & (!g726)) + ((!g1416) & (g1421) & (g1426) & (g1431) & (g677) & (g726)) + ((g1416) & (!g1421) & (!g1426) & (!g1431) & (!g677) & (!g726)) + ((g1416) & (!g1421) & (!g1426) & (g1431) & (!g677) & (!g726)) + ((g1416) & (!g1421) & (!g1426) & (g1431) & (g677) & (g726)) + ((g1416) & (!g1421) & (g1426) & (!g1431) & (!g677) & (!g726)) + ((g1416) & (!g1421) & (g1426) & (!g1431) & (!g677) & (g726)) + ((g1416) & (!g1421) & (g1426) & (g1431) & (!g677) & (!g726)) + ((g1416) & (!g1421) & (g1426) & (g1431) & (!g677) & (g726)) + ((g1416) & (!g1421) & (g1426) & (g1431) & (g677) & (g726)) + ((g1416) & (g1421) & (!g1426) & (!g1431) & (!g677) & (!g726)) + ((g1416) & (g1421) & (!g1426) & (!g1431) & (g677) & (!g726)) + ((g1416) & (g1421) & (!g1426) & (g1431) & (!g677) & (!g726)) + ((g1416) & (g1421) & (!g1426) & (g1431) & (g677) & (!g726)) + ((g1416) & (g1421) & (!g1426) & (g1431) & (g677) & (g726)) + ((g1416) & (g1421) & (g1426) & (!g1431) & (!g677) & (!g726)) + ((g1416) & (g1421) & (g1426) & (!g1431) & (!g677) & (g726)) + ((g1416) & (g1421) & (g1426) & (!g1431) & (g677) & (!g726)) + ((g1416) & (g1421) & (g1426) & (g1431) & (!g677) & (!g726)) + ((g1416) & (g1421) & (g1426) & (g1431) & (!g677) & (g726)) + ((g1416) & (g1421) & (g1426) & (g1431) & (g677) & (!g726)) + ((g1416) & (g1421) & (g1426) & (g1431) & (g677) & (g726)));
	assign g1962 = (((!g1958) & (!g1959) & (!g1960) & (g1961) & (g820) & (g773)) + ((!g1958) & (!g1959) & (g1960) & (!g1961) & (!g820) & (g773)) + ((!g1958) & (!g1959) & (g1960) & (g1961) & (!g820) & (g773)) + ((!g1958) & (!g1959) & (g1960) & (g1961) & (g820) & (g773)) + ((!g1958) & (g1959) & (!g1960) & (!g1961) & (g820) & (!g773)) + ((!g1958) & (g1959) & (!g1960) & (g1961) & (g820) & (!g773)) + ((!g1958) & (g1959) & (!g1960) & (g1961) & (g820) & (g773)) + ((!g1958) & (g1959) & (g1960) & (!g1961) & (!g820) & (g773)) + ((!g1958) & (g1959) & (g1960) & (!g1961) & (g820) & (!g773)) + ((!g1958) & (g1959) & (g1960) & (g1961) & (!g820) & (g773)) + ((!g1958) & (g1959) & (g1960) & (g1961) & (g820) & (!g773)) + ((!g1958) & (g1959) & (g1960) & (g1961) & (g820) & (g773)) + ((g1958) & (!g1959) & (!g1960) & (!g1961) & (!g820) & (!g773)) + ((g1958) & (!g1959) & (!g1960) & (g1961) & (!g820) & (!g773)) + ((g1958) & (!g1959) & (!g1960) & (g1961) & (g820) & (g773)) + ((g1958) & (!g1959) & (g1960) & (!g1961) & (!g820) & (!g773)) + ((g1958) & (!g1959) & (g1960) & (!g1961) & (!g820) & (g773)) + ((g1958) & (!g1959) & (g1960) & (g1961) & (!g820) & (!g773)) + ((g1958) & (!g1959) & (g1960) & (g1961) & (!g820) & (g773)) + ((g1958) & (!g1959) & (g1960) & (g1961) & (g820) & (g773)) + ((g1958) & (g1959) & (!g1960) & (!g1961) & (!g820) & (!g773)) + ((g1958) & (g1959) & (!g1960) & (!g1961) & (g820) & (!g773)) + ((g1958) & (g1959) & (!g1960) & (g1961) & (!g820) & (!g773)) + ((g1958) & (g1959) & (!g1960) & (g1961) & (g820) & (!g773)) + ((g1958) & (g1959) & (!g1960) & (g1961) & (g820) & (g773)) + ((g1958) & (g1959) & (g1960) & (!g1961) & (!g820) & (!g773)) + ((g1958) & (g1959) & (g1960) & (!g1961) & (!g820) & (g773)) + ((g1958) & (g1959) & (g1960) & (!g1961) & (g820) & (!g773)) + ((g1958) & (g1959) & (g1960) & (g1961) & (!g820) & (!g773)) + ((g1958) & (g1959) & (g1960) & (g1961) & (!g820) & (g773)) + ((g1958) & (g1959) & (g1960) & (g1961) & (g820) & (!g773)) + ((g1958) & (g1959) & (g1960) & (g1961) & (g820) & (g773)));
	assign g1963 = (((!g1434) & (!g1435) & (!g1436) & (g1437) & (g677) & (g726)) + ((!g1434) & (!g1435) & (g1436) & (!g1437) & (!g677) & (g726)) + ((!g1434) & (!g1435) & (g1436) & (g1437) & (!g677) & (g726)) + ((!g1434) & (!g1435) & (g1436) & (g1437) & (g677) & (g726)) + ((!g1434) & (g1435) & (!g1436) & (!g1437) & (g677) & (!g726)) + ((!g1434) & (g1435) & (!g1436) & (g1437) & (g677) & (!g726)) + ((!g1434) & (g1435) & (!g1436) & (g1437) & (g677) & (g726)) + ((!g1434) & (g1435) & (g1436) & (!g1437) & (!g677) & (g726)) + ((!g1434) & (g1435) & (g1436) & (!g1437) & (g677) & (!g726)) + ((!g1434) & (g1435) & (g1436) & (g1437) & (!g677) & (g726)) + ((!g1434) & (g1435) & (g1436) & (g1437) & (g677) & (!g726)) + ((!g1434) & (g1435) & (g1436) & (g1437) & (g677) & (g726)) + ((g1434) & (!g1435) & (!g1436) & (!g1437) & (!g677) & (!g726)) + ((g1434) & (!g1435) & (!g1436) & (g1437) & (!g677) & (!g726)) + ((g1434) & (!g1435) & (!g1436) & (g1437) & (g677) & (g726)) + ((g1434) & (!g1435) & (g1436) & (!g1437) & (!g677) & (!g726)) + ((g1434) & (!g1435) & (g1436) & (!g1437) & (!g677) & (g726)) + ((g1434) & (!g1435) & (g1436) & (g1437) & (!g677) & (!g726)) + ((g1434) & (!g1435) & (g1436) & (g1437) & (!g677) & (g726)) + ((g1434) & (!g1435) & (g1436) & (g1437) & (g677) & (g726)) + ((g1434) & (g1435) & (!g1436) & (!g1437) & (!g677) & (!g726)) + ((g1434) & (g1435) & (!g1436) & (!g1437) & (g677) & (!g726)) + ((g1434) & (g1435) & (!g1436) & (g1437) & (!g677) & (!g726)) + ((g1434) & (g1435) & (!g1436) & (g1437) & (g677) & (!g726)) + ((g1434) & (g1435) & (!g1436) & (g1437) & (g677) & (g726)) + ((g1434) & (g1435) & (g1436) & (!g1437) & (!g677) & (!g726)) + ((g1434) & (g1435) & (g1436) & (!g1437) & (!g677) & (g726)) + ((g1434) & (g1435) & (g1436) & (!g1437) & (g677) & (!g726)) + ((g1434) & (g1435) & (g1436) & (g1437) & (!g677) & (!g726)) + ((g1434) & (g1435) & (g1436) & (g1437) & (!g677) & (g726)) + ((g1434) & (g1435) & (g1436) & (g1437) & (g677) & (!g726)) + ((g1434) & (g1435) & (g1436) & (g1437) & (g677) & (g726)));
	assign g1964 = (((!g677) & (!g726) & (!g1439) & (!sk[110]) & (g1440) & (!g1441)) + ((!g677) & (!g726) & (!g1439) & (!sk[110]) & (g1440) & (g1441)) + ((!g677) & (!g726) & (g1439) & (!sk[110]) & (!g1440) & (!g1441)) + ((!g677) & (!g726) & (g1439) & (!sk[110]) & (!g1440) & (g1441)) + ((!g677) & (!g726) & (g1439) & (!sk[110]) & (g1440) & (!g1441)) + ((!g677) & (!g726) & (g1439) & (!sk[110]) & (g1440) & (g1441)) + ((!g677) & (g726) & (!g1439) & (!sk[110]) & (!g1440) & (!g1441)) + ((!g677) & (g726) & (!g1439) & (!sk[110]) & (!g1440) & (g1441)) + ((!g677) & (g726) & (!g1439) & (!sk[110]) & (g1440) & (!g1441)) + ((!g677) & (g726) & (!g1439) & (!sk[110]) & (g1440) & (g1441)) + ((!g677) & (g726) & (!g1439) & (sk[110]) & (!g1440) & (g1441)) + ((!g677) & (g726) & (!g1439) & (sk[110]) & (g1440) & (g1441)) + ((!g677) & (g726) & (g1439) & (!sk[110]) & (!g1440) & (!g1441)) + ((!g677) & (g726) & (g1439) & (!sk[110]) & (!g1440) & (g1441)) + ((!g677) & (g726) & (g1439) & (!sk[110]) & (g1440) & (!g1441)) + ((!g677) & (g726) & (g1439) & (!sk[110]) & (g1440) & (g1441)) + ((!g677) & (g726) & (g1439) & (sk[110]) & (!g1440) & (g1441)) + ((!g677) & (g726) & (g1439) & (sk[110]) & (g1440) & (g1441)) + ((g677) & (!g726) & (!g1439) & (!sk[110]) & (g1440) & (!g1441)) + ((g677) & (!g726) & (!g1439) & (!sk[110]) & (g1440) & (g1441)) + ((g677) & (!g726) & (g1439) & (!sk[110]) & (!g1440) & (!g1441)) + ((g677) & (!g726) & (g1439) & (!sk[110]) & (!g1440) & (g1441)) + ((g677) & (!g726) & (g1439) & (!sk[110]) & (g1440) & (!g1441)) + ((g677) & (!g726) & (g1439) & (!sk[110]) & (g1440) & (g1441)) + ((g677) & (!g726) & (g1439) & (sk[110]) & (!g1440) & (!g1441)) + ((g677) & (!g726) & (g1439) & (sk[110]) & (!g1440) & (g1441)) + ((g677) & (!g726) & (g1439) & (sk[110]) & (g1440) & (!g1441)) + ((g677) & (!g726) & (g1439) & (sk[110]) & (g1440) & (g1441)) + ((g677) & (g726) & (!g1439) & (!sk[110]) & (!g1440) & (!g1441)) + ((g677) & (g726) & (!g1439) & (!sk[110]) & (!g1440) & (g1441)) + ((g677) & (g726) & (!g1439) & (!sk[110]) & (g1440) & (!g1441)) + ((g677) & (g726) & (!g1439) & (!sk[110]) & (g1440) & (g1441)) + ((g677) & (g726) & (!g1439) & (sk[110]) & (g1440) & (!g1441)) + ((g677) & (g726) & (!g1439) & (sk[110]) & (g1440) & (g1441)) + ((g677) & (g726) & (g1439) & (!sk[110]) & (!g1440) & (!g1441)) + ((g677) & (g726) & (g1439) & (!sk[110]) & (!g1440) & (g1441)) + ((g677) & (g726) & (g1439) & (!sk[110]) & (g1440) & (!g1441)) + ((g677) & (g726) & (g1439) & (!sk[110]) & (g1440) & (g1441)) + ((g677) & (g726) & (g1439) & (sk[110]) & (g1440) & (!g1441)) + ((g677) & (g726) & (g1439) & (sk[110]) & (g1440) & (g1441)));
	assign g1965 = (((!g1443) & (!g1444) & (!g1445) & (g1446) & (g677) & (g726)) + ((!g1443) & (!g1444) & (g1445) & (!g1446) & (!g677) & (g726)) + ((!g1443) & (!g1444) & (g1445) & (g1446) & (!g677) & (g726)) + ((!g1443) & (!g1444) & (g1445) & (g1446) & (g677) & (g726)) + ((!g1443) & (g1444) & (!g1445) & (!g1446) & (g677) & (!g726)) + ((!g1443) & (g1444) & (!g1445) & (g1446) & (g677) & (!g726)) + ((!g1443) & (g1444) & (!g1445) & (g1446) & (g677) & (g726)) + ((!g1443) & (g1444) & (g1445) & (!g1446) & (!g677) & (g726)) + ((!g1443) & (g1444) & (g1445) & (!g1446) & (g677) & (!g726)) + ((!g1443) & (g1444) & (g1445) & (g1446) & (!g677) & (g726)) + ((!g1443) & (g1444) & (g1445) & (g1446) & (g677) & (!g726)) + ((!g1443) & (g1444) & (g1445) & (g1446) & (g677) & (g726)) + ((g1443) & (!g1444) & (!g1445) & (!g1446) & (!g677) & (!g726)) + ((g1443) & (!g1444) & (!g1445) & (g1446) & (!g677) & (!g726)) + ((g1443) & (!g1444) & (!g1445) & (g1446) & (g677) & (g726)) + ((g1443) & (!g1444) & (g1445) & (!g1446) & (!g677) & (!g726)) + ((g1443) & (!g1444) & (g1445) & (!g1446) & (!g677) & (g726)) + ((g1443) & (!g1444) & (g1445) & (g1446) & (!g677) & (!g726)) + ((g1443) & (!g1444) & (g1445) & (g1446) & (!g677) & (g726)) + ((g1443) & (!g1444) & (g1445) & (g1446) & (g677) & (g726)) + ((g1443) & (g1444) & (!g1445) & (!g1446) & (!g677) & (!g726)) + ((g1443) & (g1444) & (!g1445) & (!g1446) & (g677) & (!g726)) + ((g1443) & (g1444) & (!g1445) & (g1446) & (!g677) & (!g726)) + ((g1443) & (g1444) & (!g1445) & (g1446) & (g677) & (!g726)) + ((g1443) & (g1444) & (!g1445) & (g1446) & (g677) & (g726)) + ((g1443) & (g1444) & (g1445) & (!g1446) & (!g677) & (!g726)) + ((g1443) & (g1444) & (g1445) & (!g1446) & (!g677) & (g726)) + ((g1443) & (g1444) & (g1445) & (!g1446) & (g677) & (!g726)) + ((g1443) & (g1444) & (g1445) & (g1446) & (!g677) & (!g726)) + ((g1443) & (g1444) & (g1445) & (g1446) & (!g677) & (g726)) + ((g1443) & (g1444) & (g1445) & (g1446) & (g677) & (!g726)) + ((g1443) & (g1444) & (g1445) & (g1446) & (g677) & (g726)));
	assign g1966 = (((!g1448) & (!g1449) & (!g1450) & (g1451) & (g677) & (g726)) + ((!g1448) & (!g1449) & (g1450) & (!g1451) & (!g677) & (g726)) + ((!g1448) & (!g1449) & (g1450) & (g1451) & (!g677) & (g726)) + ((!g1448) & (!g1449) & (g1450) & (g1451) & (g677) & (g726)) + ((!g1448) & (g1449) & (!g1450) & (!g1451) & (g677) & (!g726)) + ((!g1448) & (g1449) & (!g1450) & (g1451) & (g677) & (!g726)) + ((!g1448) & (g1449) & (!g1450) & (g1451) & (g677) & (g726)) + ((!g1448) & (g1449) & (g1450) & (!g1451) & (!g677) & (g726)) + ((!g1448) & (g1449) & (g1450) & (!g1451) & (g677) & (!g726)) + ((!g1448) & (g1449) & (g1450) & (g1451) & (!g677) & (g726)) + ((!g1448) & (g1449) & (g1450) & (g1451) & (g677) & (!g726)) + ((!g1448) & (g1449) & (g1450) & (g1451) & (g677) & (g726)) + ((g1448) & (!g1449) & (!g1450) & (!g1451) & (!g677) & (!g726)) + ((g1448) & (!g1449) & (!g1450) & (g1451) & (!g677) & (!g726)) + ((g1448) & (!g1449) & (!g1450) & (g1451) & (g677) & (g726)) + ((g1448) & (!g1449) & (g1450) & (!g1451) & (!g677) & (!g726)) + ((g1448) & (!g1449) & (g1450) & (!g1451) & (!g677) & (g726)) + ((g1448) & (!g1449) & (g1450) & (g1451) & (!g677) & (!g726)) + ((g1448) & (!g1449) & (g1450) & (g1451) & (!g677) & (g726)) + ((g1448) & (!g1449) & (g1450) & (g1451) & (g677) & (g726)) + ((g1448) & (g1449) & (!g1450) & (!g1451) & (!g677) & (!g726)) + ((g1448) & (g1449) & (!g1450) & (!g1451) & (g677) & (!g726)) + ((g1448) & (g1449) & (!g1450) & (g1451) & (!g677) & (!g726)) + ((g1448) & (g1449) & (!g1450) & (g1451) & (g677) & (!g726)) + ((g1448) & (g1449) & (!g1450) & (g1451) & (g677) & (g726)) + ((g1448) & (g1449) & (g1450) & (!g1451) & (!g677) & (!g726)) + ((g1448) & (g1449) & (g1450) & (!g1451) & (!g677) & (g726)) + ((g1448) & (g1449) & (g1450) & (!g1451) & (g677) & (!g726)) + ((g1448) & (g1449) & (g1450) & (g1451) & (!g677) & (!g726)) + ((g1448) & (g1449) & (g1450) & (g1451) & (!g677) & (g726)) + ((g1448) & (g1449) & (g1450) & (g1451) & (g677) & (!g726)) + ((g1448) & (g1449) & (g1450) & (g1451) & (g677) & (g726)));
	assign g1967 = (((!g820) & (!g773) & (!g1963) & (g1964) & (!g1965) & (!g1966)) + ((!g820) & (!g773) & (!g1963) & (g1964) & (!g1965) & (g1966)) + ((!g820) & (!g773) & (!g1963) & (g1964) & (g1965) & (!g1966)) + ((!g820) & (!g773) & (!g1963) & (g1964) & (g1965) & (g1966)) + ((!g820) & (!g773) & (g1963) & (g1964) & (!g1965) & (!g1966)) + ((!g820) & (!g773) & (g1963) & (g1964) & (!g1965) & (g1966)) + ((!g820) & (!g773) & (g1963) & (g1964) & (g1965) & (!g1966)) + ((!g820) & (!g773) & (g1963) & (g1964) & (g1965) & (g1966)) + ((!g820) & (g773) & (!g1963) & (!g1964) & (!g1965) & (g1966)) + ((!g820) & (g773) & (!g1963) & (!g1964) & (g1965) & (g1966)) + ((!g820) & (g773) & (!g1963) & (g1964) & (!g1965) & (g1966)) + ((!g820) & (g773) & (!g1963) & (g1964) & (g1965) & (g1966)) + ((!g820) & (g773) & (g1963) & (!g1964) & (!g1965) & (g1966)) + ((!g820) & (g773) & (g1963) & (!g1964) & (g1965) & (g1966)) + ((!g820) & (g773) & (g1963) & (g1964) & (!g1965) & (g1966)) + ((!g820) & (g773) & (g1963) & (g1964) & (g1965) & (g1966)) + ((g820) & (!g773) & (g1963) & (!g1964) & (!g1965) & (!g1966)) + ((g820) & (!g773) & (g1963) & (!g1964) & (!g1965) & (g1966)) + ((g820) & (!g773) & (g1963) & (!g1964) & (g1965) & (!g1966)) + ((g820) & (!g773) & (g1963) & (!g1964) & (g1965) & (g1966)) + ((g820) & (!g773) & (g1963) & (g1964) & (!g1965) & (!g1966)) + ((g820) & (!g773) & (g1963) & (g1964) & (!g1965) & (g1966)) + ((g820) & (!g773) & (g1963) & (g1964) & (g1965) & (!g1966)) + ((g820) & (!g773) & (g1963) & (g1964) & (g1965) & (g1966)) + ((g820) & (g773) & (!g1963) & (!g1964) & (g1965) & (!g1966)) + ((g820) & (g773) & (!g1963) & (!g1964) & (g1965) & (g1966)) + ((g820) & (g773) & (!g1963) & (g1964) & (g1965) & (!g1966)) + ((g820) & (g773) & (!g1963) & (g1964) & (g1965) & (g1966)) + ((g820) & (g773) & (g1963) & (!g1964) & (g1965) & (!g1966)) + ((g820) & (g773) & (g1963) & (!g1964) & (g1965) & (g1966)) + ((g820) & (g773) & (g1963) & (g1964) & (g1965) & (!g1966)) + ((g820) & (g773) & (g1963) & (g1964) & (g1965) & (g1966)));
	assign g1968 = (((!g867) & (!sk[114]) & (!g1962) & (g1967)) + ((!g867) & (!sk[114]) & (g1962) & (!g1967)) + ((!g867) & (!sk[114]) & (g1962) & (g1967)) + ((!g867) & (sk[114]) & (!g1962) & (g1967)) + ((!g867) & (sk[114]) & (g1962) & (g1967)) + ((g867) & (!sk[114]) & (!g1962) & (g1967)) + ((g867) & (!sk[114]) & (g1962) & (!g1967)) + ((g867) & (!sk[114]) & (g1962) & (g1967)) + ((g867) & (sk[114]) & (g1962) & (!g1967)) + ((g867) & (sk[114]) & (g1962) & (g1967)));
	assign g1969 = (((!g1593) & (!g1605) & (!sk[115]) & (!g1759) & (g63)) + ((!g1593) & (!g1605) & (!sk[115]) & (g1759) & (!g63)) + ((!g1593) & (!g1605) & (!sk[115]) & (g1759) & (g63)) + ((!g1593) & (!g1605) & (sk[115]) & (g1759) & (!g63)) + ((!g1593) & (!g1605) & (sk[115]) & (g1759) & (g63)) + ((!g1593) & (g1605) & (!sk[115]) & (!g1759) & (!g63)) + ((!g1593) & (g1605) & (!sk[115]) & (!g1759) & (g63)) + ((!g1593) & (g1605) & (!sk[115]) & (g1759) & (!g63)) + ((!g1593) & (g1605) & (!sk[115]) & (g1759) & (g63)) + ((g1593) & (!g1605) & (!sk[115]) & (!g1759) & (g63)) + ((g1593) & (!g1605) & (!sk[115]) & (g1759) & (!g63)) + ((g1593) & (!g1605) & (!sk[115]) & (g1759) & (g63)) + ((g1593) & (!g1605) & (sk[115]) & (!g1759) & (g63)) + ((g1593) & (!g1605) & (sk[115]) & (g1759) & (g63)) + ((g1593) & (g1605) & (!sk[115]) & (!g1759) & (!g63)) + ((g1593) & (g1605) & (!sk[115]) & (!g1759) & (g63)) + ((g1593) & (g1605) & (!sk[115]) & (g1759) & (!g63)) + ((g1593) & (g1605) & (!sk[115]) & (g1759) & (g63)) + ((g1593) & (g1605) & (sk[115]) & (!g1759) & (g63)) + ((g1593) & (g1605) & (sk[115]) & (g1759) & (g63)));
	assign g1970 = (((!g132) & (!g1592) & (g1656) & (g1917) & (!g1968) & (!g1969)) + ((!g132) & (!g1592) & (g1656) & (g1917) & (!g1968) & (g1969)) + ((!g132) & (!g1592) & (g1656) & (g1917) & (g1968) & (!g1969)) + ((!g132) & (!g1592) & (g1656) & (g1917) & (g1968) & (g1969)) + ((!g132) & (g1592) & (!g1656) & (g1917) & (!g1968) & (g1969)) + ((!g132) & (g1592) & (!g1656) & (g1917) & (g1968) & (g1969)) + ((!g132) & (g1592) & (g1656) & (g1917) & (!g1968) & (g1969)) + ((!g132) & (g1592) & (g1656) & (g1917) & (g1968) & (g1969)) + ((g132) & (!g1592) & (!g1656) & (g1917) & (g1968) & (!g1969)) + ((g132) & (!g1592) & (!g1656) & (g1917) & (g1968) & (g1969)) + ((g132) & (!g1592) & (g1656) & (g1917) & (g1968) & (!g1969)) + ((g132) & (!g1592) & (g1656) & (g1917) & (g1968) & (g1969)) + ((g132) & (g1592) & (!g1656) & (g1917) & (g1968) & (!g1969)) + ((g132) & (g1592) & (!g1656) & (g1917) & (g1968) & (g1969)) + ((g132) & (g1592) & (g1656) & (g1917) & (g1968) & (!g1969)) + ((g132) & (g1592) & (g1656) & (g1917) & (g1968) & (g1969)));
	assign g1971 = (((!g1458) & (!g1459) & (!g1460) & (g1461) & (g820) & (g773)) + ((!g1458) & (!g1459) & (g1460) & (!g1461) & (!g820) & (g773)) + ((!g1458) & (!g1459) & (g1460) & (g1461) & (!g820) & (g773)) + ((!g1458) & (!g1459) & (g1460) & (g1461) & (g820) & (g773)) + ((!g1458) & (g1459) & (!g1460) & (!g1461) & (g820) & (!g773)) + ((!g1458) & (g1459) & (!g1460) & (g1461) & (g820) & (!g773)) + ((!g1458) & (g1459) & (!g1460) & (g1461) & (g820) & (g773)) + ((!g1458) & (g1459) & (g1460) & (!g1461) & (!g820) & (g773)) + ((!g1458) & (g1459) & (g1460) & (!g1461) & (g820) & (!g773)) + ((!g1458) & (g1459) & (g1460) & (g1461) & (!g820) & (g773)) + ((!g1458) & (g1459) & (g1460) & (g1461) & (g820) & (!g773)) + ((!g1458) & (g1459) & (g1460) & (g1461) & (g820) & (g773)) + ((g1458) & (!g1459) & (!g1460) & (!g1461) & (!g820) & (!g773)) + ((g1458) & (!g1459) & (!g1460) & (g1461) & (!g820) & (!g773)) + ((g1458) & (!g1459) & (!g1460) & (g1461) & (g820) & (g773)) + ((g1458) & (!g1459) & (g1460) & (!g1461) & (!g820) & (!g773)) + ((g1458) & (!g1459) & (g1460) & (!g1461) & (!g820) & (g773)) + ((g1458) & (!g1459) & (g1460) & (g1461) & (!g820) & (!g773)) + ((g1458) & (!g1459) & (g1460) & (g1461) & (!g820) & (g773)) + ((g1458) & (!g1459) & (g1460) & (g1461) & (g820) & (g773)) + ((g1458) & (g1459) & (!g1460) & (!g1461) & (!g820) & (!g773)) + ((g1458) & (g1459) & (!g1460) & (!g1461) & (g820) & (!g773)) + ((g1458) & (g1459) & (!g1460) & (g1461) & (!g820) & (!g773)) + ((g1458) & (g1459) & (!g1460) & (g1461) & (g820) & (!g773)) + ((g1458) & (g1459) & (!g1460) & (g1461) & (g820) & (g773)) + ((g1458) & (g1459) & (g1460) & (!g1461) & (!g820) & (!g773)) + ((g1458) & (g1459) & (g1460) & (!g1461) & (!g820) & (g773)) + ((g1458) & (g1459) & (g1460) & (!g1461) & (g820) & (!g773)) + ((g1458) & (g1459) & (g1460) & (g1461) & (!g820) & (!g773)) + ((g1458) & (g1459) & (g1460) & (g1461) & (!g820) & (g773)) + ((g1458) & (g1459) & (g1460) & (g1461) & (g820) & (!g773)) + ((g1458) & (g1459) & (g1460) & (g1461) & (g820) & (g773)));
	assign g1972 = (((!g1463) & (!g1464) & (!g1465) & (g1466) & (g820) & (g773)) + ((!g1463) & (!g1464) & (g1465) & (!g1466) & (!g820) & (g773)) + ((!g1463) & (!g1464) & (g1465) & (g1466) & (!g820) & (g773)) + ((!g1463) & (!g1464) & (g1465) & (g1466) & (g820) & (g773)) + ((!g1463) & (g1464) & (!g1465) & (!g1466) & (g820) & (!g773)) + ((!g1463) & (g1464) & (!g1465) & (g1466) & (g820) & (!g773)) + ((!g1463) & (g1464) & (!g1465) & (g1466) & (g820) & (g773)) + ((!g1463) & (g1464) & (g1465) & (!g1466) & (!g820) & (g773)) + ((!g1463) & (g1464) & (g1465) & (!g1466) & (g820) & (!g773)) + ((!g1463) & (g1464) & (g1465) & (g1466) & (!g820) & (g773)) + ((!g1463) & (g1464) & (g1465) & (g1466) & (g820) & (!g773)) + ((!g1463) & (g1464) & (g1465) & (g1466) & (g820) & (g773)) + ((g1463) & (!g1464) & (!g1465) & (!g1466) & (!g820) & (!g773)) + ((g1463) & (!g1464) & (!g1465) & (g1466) & (!g820) & (!g773)) + ((g1463) & (!g1464) & (!g1465) & (g1466) & (g820) & (g773)) + ((g1463) & (!g1464) & (g1465) & (!g1466) & (!g820) & (!g773)) + ((g1463) & (!g1464) & (g1465) & (!g1466) & (!g820) & (g773)) + ((g1463) & (!g1464) & (g1465) & (g1466) & (!g820) & (!g773)) + ((g1463) & (!g1464) & (g1465) & (g1466) & (!g820) & (g773)) + ((g1463) & (!g1464) & (g1465) & (g1466) & (g820) & (g773)) + ((g1463) & (g1464) & (!g1465) & (!g1466) & (!g820) & (!g773)) + ((g1463) & (g1464) & (!g1465) & (!g1466) & (g820) & (!g773)) + ((g1463) & (g1464) & (!g1465) & (g1466) & (!g820) & (!g773)) + ((g1463) & (g1464) & (!g1465) & (g1466) & (g820) & (!g773)) + ((g1463) & (g1464) & (!g1465) & (g1466) & (g820) & (g773)) + ((g1463) & (g1464) & (g1465) & (!g1466) & (!g820) & (!g773)) + ((g1463) & (g1464) & (g1465) & (!g1466) & (!g820) & (g773)) + ((g1463) & (g1464) & (g1465) & (!g1466) & (g820) & (!g773)) + ((g1463) & (g1464) & (g1465) & (g1466) & (!g820) & (!g773)) + ((g1463) & (g1464) & (g1465) & (g1466) & (!g820) & (g773)) + ((g1463) & (g1464) & (g1465) & (g1466) & (g820) & (!g773)) + ((g1463) & (g1464) & (g1465) & (g1466) & (g820) & (g773)));
	assign g1973 = (((!g1468) & (!g1469) & (!g1470) & (g1471) & (g820) & (g773)) + ((!g1468) & (!g1469) & (g1470) & (!g1471) & (!g820) & (g773)) + ((!g1468) & (!g1469) & (g1470) & (g1471) & (!g820) & (g773)) + ((!g1468) & (!g1469) & (g1470) & (g1471) & (g820) & (g773)) + ((!g1468) & (g1469) & (!g1470) & (!g1471) & (g820) & (!g773)) + ((!g1468) & (g1469) & (!g1470) & (g1471) & (g820) & (!g773)) + ((!g1468) & (g1469) & (!g1470) & (g1471) & (g820) & (g773)) + ((!g1468) & (g1469) & (g1470) & (!g1471) & (!g820) & (g773)) + ((!g1468) & (g1469) & (g1470) & (!g1471) & (g820) & (!g773)) + ((!g1468) & (g1469) & (g1470) & (g1471) & (!g820) & (g773)) + ((!g1468) & (g1469) & (g1470) & (g1471) & (g820) & (!g773)) + ((!g1468) & (g1469) & (g1470) & (g1471) & (g820) & (g773)) + ((g1468) & (!g1469) & (!g1470) & (!g1471) & (!g820) & (!g773)) + ((g1468) & (!g1469) & (!g1470) & (g1471) & (!g820) & (!g773)) + ((g1468) & (!g1469) & (!g1470) & (g1471) & (g820) & (g773)) + ((g1468) & (!g1469) & (g1470) & (!g1471) & (!g820) & (!g773)) + ((g1468) & (!g1469) & (g1470) & (!g1471) & (!g820) & (g773)) + ((g1468) & (!g1469) & (g1470) & (g1471) & (!g820) & (!g773)) + ((g1468) & (!g1469) & (g1470) & (g1471) & (!g820) & (g773)) + ((g1468) & (!g1469) & (g1470) & (g1471) & (g820) & (g773)) + ((g1468) & (g1469) & (!g1470) & (!g1471) & (!g820) & (!g773)) + ((g1468) & (g1469) & (!g1470) & (!g1471) & (g820) & (!g773)) + ((g1468) & (g1469) & (!g1470) & (g1471) & (!g820) & (!g773)) + ((g1468) & (g1469) & (!g1470) & (g1471) & (g820) & (!g773)) + ((g1468) & (g1469) & (!g1470) & (g1471) & (g820) & (g773)) + ((g1468) & (g1469) & (g1470) & (!g1471) & (!g820) & (!g773)) + ((g1468) & (g1469) & (g1470) & (!g1471) & (!g820) & (g773)) + ((g1468) & (g1469) & (g1470) & (!g1471) & (g820) & (!g773)) + ((g1468) & (g1469) & (g1470) & (g1471) & (!g820) & (!g773)) + ((g1468) & (g1469) & (g1470) & (g1471) & (!g820) & (g773)) + ((g1468) & (g1469) & (g1470) & (g1471) & (g820) & (!g773)) + ((g1468) & (g1469) & (g1470) & (g1471) & (g820) & (g773)));
	assign g1974 = (((!g1473) & (!g1474) & (!g1475) & (g1476) & (g820) & (g773)) + ((!g1473) & (!g1474) & (g1475) & (!g1476) & (!g820) & (g773)) + ((!g1473) & (!g1474) & (g1475) & (g1476) & (!g820) & (g773)) + ((!g1473) & (!g1474) & (g1475) & (g1476) & (g820) & (g773)) + ((!g1473) & (g1474) & (!g1475) & (!g1476) & (g820) & (!g773)) + ((!g1473) & (g1474) & (!g1475) & (g1476) & (g820) & (!g773)) + ((!g1473) & (g1474) & (!g1475) & (g1476) & (g820) & (g773)) + ((!g1473) & (g1474) & (g1475) & (!g1476) & (!g820) & (g773)) + ((!g1473) & (g1474) & (g1475) & (!g1476) & (g820) & (!g773)) + ((!g1473) & (g1474) & (g1475) & (g1476) & (!g820) & (g773)) + ((!g1473) & (g1474) & (g1475) & (g1476) & (g820) & (!g773)) + ((!g1473) & (g1474) & (g1475) & (g1476) & (g820) & (g773)) + ((g1473) & (!g1474) & (!g1475) & (!g1476) & (!g820) & (!g773)) + ((g1473) & (!g1474) & (!g1475) & (g1476) & (!g820) & (!g773)) + ((g1473) & (!g1474) & (!g1475) & (g1476) & (g820) & (g773)) + ((g1473) & (!g1474) & (g1475) & (!g1476) & (!g820) & (!g773)) + ((g1473) & (!g1474) & (g1475) & (!g1476) & (!g820) & (g773)) + ((g1473) & (!g1474) & (g1475) & (g1476) & (!g820) & (!g773)) + ((g1473) & (!g1474) & (g1475) & (g1476) & (!g820) & (g773)) + ((g1473) & (!g1474) & (g1475) & (g1476) & (g820) & (g773)) + ((g1473) & (g1474) & (!g1475) & (!g1476) & (!g820) & (!g773)) + ((g1473) & (g1474) & (!g1475) & (!g1476) & (g820) & (!g773)) + ((g1473) & (g1474) & (!g1475) & (g1476) & (!g820) & (!g773)) + ((g1473) & (g1474) & (!g1475) & (g1476) & (g820) & (!g773)) + ((g1473) & (g1474) & (!g1475) & (g1476) & (g820) & (g773)) + ((g1473) & (g1474) & (g1475) & (!g1476) & (!g820) & (!g773)) + ((g1473) & (g1474) & (g1475) & (!g1476) & (!g820) & (g773)) + ((g1473) & (g1474) & (g1475) & (!g1476) & (g820) & (!g773)) + ((g1473) & (g1474) & (g1475) & (g1476) & (!g820) & (!g773)) + ((g1473) & (g1474) & (g1475) & (g1476) & (!g820) & (g773)) + ((g1473) & (g1474) & (g1475) & (g1476) & (g820) & (!g773)) + ((g1473) & (g1474) & (g1475) & (g1476) & (g820) & (g773)));
	assign g1975 = (((!g1971) & (!g1972) & (!g1973) & (g1974) & (g677) & (g726)) + ((!g1971) & (!g1972) & (g1973) & (!g1974) & (!g677) & (g726)) + ((!g1971) & (!g1972) & (g1973) & (g1974) & (!g677) & (g726)) + ((!g1971) & (!g1972) & (g1973) & (g1974) & (g677) & (g726)) + ((!g1971) & (g1972) & (!g1973) & (!g1974) & (g677) & (!g726)) + ((!g1971) & (g1972) & (!g1973) & (g1974) & (g677) & (!g726)) + ((!g1971) & (g1972) & (!g1973) & (g1974) & (g677) & (g726)) + ((!g1971) & (g1972) & (g1973) & (!g1974) & (!g677) & (g726)) + ((!g1971) & (g1972) & (g1973) & (!g1974) & (g677) & (!g726)) + ((!g1971) & (g1972) & (g1973) & (g1974) & (!g677) & (g726)) + ((!g1971) & (g1972) & (g1973) & (g1974) & (g677) & (!g726)) + ((!g1971) & (g1972) & (g1973) & (g1974) & (g677) & (g726)) + ((g1971) & (!g1972) & (!g1973) & (!g1974) & (!g677) & (!g726)) + ((g1971) & (!g1972) & (!g1973) & (g1974) & (!g677) & (!g726)) + ((g1971) & (!g1972) & (!g1973) & (g1974) & (g677) & (g726)) + ((g1971) & (!g1972) & (g1973) & (!g1974) & (!g677) & (!g726)) + ((g1971) & (!g1972) & (g1973) & (!g1974) & (!g677) & (g726)) + ((g1971) & (!g1972) & (g1973) & (g1974) & (!g677) & (!g726)) + ((g1971) & (!g1972) & (g1973) & (g1974) & (!g677) & (g726)) + ((g1971) & (!g1972) & (g1973) & (g1974) & (g677) & (g726)) + ((g1971) & (g1972) & (!g1973) & (!g1974) & (!g677) & (!g726)) + ((g1971) & (g1972) & (!g1973) & (!g1974) & (g677) & (!g726)) + ((g1971) & (g1972) & (!g1973) & (g1974) & (!g677) & (!g726)) + ((g1971) & (g1972) & (!g1973) & (g1974) & (g677) & (!g726)) + ((g1971) & (g1972) & (!g1973) & (g1974) & (g677) & (g726)) + ((g1971) & (g1972) & (g1973) & (!g1974) & (!g677) & (!g726)) + ((g1971) & (g1972) & (g1973) & (!g1974) & (!g677) & (g726)) + ((g1971) & (g1972) & (g1973) & (!g1974) & (g677) & (!g726)) + ((g1971) & (g1972) & (g1973) & (g1974) & (!g677) & (!g726)) + ((g1971) & (g1972) & (g1973) & (g1974) & (!g677) & (g726)) + ((g1971) & (g1972) & (g1973) & (g1974) & (g677) & (!g726)) + ((g1971) & (g1972) & (g1973) & (g1974) & (g677) & (g726)));
	assign g1976 = (((!g1479) & (!g1480) & (!g1481) & (g1482) & (g677) & (g726)) + ((!g1479) & (!g1480) & (g1481) & (!g1482) & (!g677) & (g726)) + ((!g1479) & (!g1480) & (g1481) & (g1482) & (!g677) & (g726)) + ((!g1479) & (!g1480) & (g1481) & (g1482) & (g677) & (g726)) + ((!g1479) & (g1480) & (!g1481) & (!g1482) & (g677) & (!g726)) + ((!g1479) & (g1480) & (!g1481) & (g1482) & (g677) & (!g726)) + ((!g1479) & (g1480) & (!g1481) & (g1482) & (g677) & (g726)) + ((!g1479) & (g1480) & (g1481) & (!g1482) & (!g677) & (g726)) + ((!g1479) & (g1480) & (g1481) & (!g1482) & (g677) & (!g726)) + ((!g1479) & (g1480) & (g1481) & (g1482) & (!g677) & (g726)) + ((!g1479) & (g1480) & (g1481) & (g1482) & (g677) & (!g726)) + ((!g1479) & (g1480) & (g1481) & (g1482) & (g677) & (g726)) + ((g1479) & (!g1480) & (!g1481) & (!g1482) & (!g677) & (!g726)) + ((g1479) & (!g1480) & (!g1481) & (g1482) & (!g677) & (!g726)) + ((g1479) & (!g1480) & (!g1481) & (g1482) & (g677) & (g726)) + ((g1479) & (!g1480) & (g1481) & (!g1482) & (!g677) & (!g726)) + ((g1479) & (!g1480) & (g1481) & (!g1482) & (!g677) & (g726)) + ((g1479) & (!g1480) & (g1481) & (g1482) & (!g677) & (!g726)) + ((g1479) & (!g1480) & (g1481) & (g1482) & (!g677) & (g726)) + ((g1479) & (!g1480) & (g1481) & (g1482) & (g677) & (g726)) + ((g1479) & (g1480) & (!g1481) & (!g1482) & (!g677) & (!g726)) + ((g1479) & (g1480) & (!g1481) & (!g1482) & (g677) & (!g726)) + ((g1479) & (g1480) & (!g1481) & (g1482) & (!g677) & (!g726)) + ((g1479) & (g1480) & (!g1481) & (g1482) & (g677) & (!g726)) + ((g1479) & (g1480) & (!g1481) & (g1482) & (g677) & (g726)) + ((g1479) & (g1480) & (g1481) & (!g1482) & (!g677) & (!g726)) + ((g1479) & (g1480) & (g1481) & (!g1482) & (!g677) & (g726)) + ((g1479) & (g1480) & (g1481) & (!g1482) & (g677) & (!g726)) + ((g1479) & (g1480) & (g1481) & (g1482) & (!g677) & (!g726)) + ((g1479) & (g1480) & (g1481) & (g1482) & (!g677) & (g726)) + ((g1479) & (g1480) & (g1481) & (g1482) & (g677) & (!g726)) + ((g1479) & (g1480) & (g1481) & (g1482) & (g677) & (g726)));
	assign g1977 = (((!g677) & (!g726) & (!sk[123]) & (!g1484) & (g1485) & (!g1486)) + ((!g677) & (!g726) & (!sk[123]) & (!g1484) & (g1485) & (g1486)) + ((!g677) & (!g726) & (!sk[123]) & (g1484) & (!g1485) & (!g1486)) + ((!g677) & (!g726) & (!sk[123]) & (g1484) & (!g1485) & (g1486)) + ((!g677) & (!g726) & (!sk[123]) & (g1484) & (g1485) & (!g1486)) + ((!g677) & (!g726) & (!sk[123]) & (g1484) & (g1485) & (g1486)) + ((!g677) & (g726) & (!sk[123]) & (!g1484) & (!g1485) & (!g1486)) + ((!g677) & (g726) & (!sk[123]) & (!g1484) & (!g1485) & (g1486)) + ((!g677) & (g726) & (!sk[123]) & (!g1484) & (g1485) & (!g1486)) + ((!g677) & (g726) & (!sk[123]) & (!g1484) & (g1485) & (g1486)) + ((!g677) & (g726) & (!sk[123]) & (g1484) & (!g1485) & (!g1486)) + ((!g677) & (g726) & (!sk[123]) & (g1484) & (!g1485) & (g1486)) + ((!g677) & (g726) & (!sk[123]) & (g1484) & (g1485) & (!g1486)) + ((!g677) & (g726) & (!sk[123]) & (g1484) & (g1485) & (g1486)) + ((!g677) & (g726) & (sk[123]) & (!g1484) & (!g1485) & (g1486)) + ((!g677) & (g726) & (sk[123]) & (!g1484) & (g1485) & (g1486)) + ((!g677) & (g726) & (sk[123]) & (g1484) & (!g1485) & (g1486)) + ((!g677) & (g726) & (sk[123]) & (g1484) & (g1485) & (g1486)) + ((g677) & (!g726) & (!sk[123]) & (!g1484) & (g1485) & (!g1486)) + ((g677) & (!g726) & (!sk[123]) & (!g1484) & (g1485) & (g1486)) + ((g677) & (!g726) & (!sk[123]) & (g1484) & (!g1485) & (!g1486)) + ((g677) & (!g726) & (!sk[123]) & (g1484) & (!g1485) & (g1486)) + ((g677) & (!g726) & (!sk[123]) & (g1484) & (g1485) & (!g1486)) + ((g677) & (!g726) & (!sk[123]) & (g1484) & (g1485) & (g1486)) + ((g677) & (!g726) & (sk[123]) & (g1484) & (!g1485) & (!g1486)) + ((g677) & (!g726) & (sk[123]) & (g1484) & (!g1485) & (g1486)) + ((g677) & (!g726) & (sk[123]) & (g1484) & (g1485) & (!g1486)) + ((g677) & (!g726) & (sk[123]) & (g1484) & (g1485) & (g1486)) + ((g677) & (g726) & (!sk[123]) & (!g1484) & (!g1485) & (!g1486)) + ((g677) & (g726) & (!sk[123]) & (!g1484) & (!g1485) & (g1486)) + ((g677) & (g726) & (!sk[123]) & (!g1484) & (g1485) & (!g1486)) + ((g677) & (g726) & (!sk[123]) & (!g1484) & (g1485) & (g1486)) + ((g677) & (g726) & (!sk[123]) & (g1484) & (!g1485) & (!g1486)) + ((g677) & (g726) & (!sk[123]) & (g1484) & (!g1485) & (g1486)) + ((g677) & (g726) & (!sk[123]) & (g1484) & (g1485) & (!g1486)) + ((g677) & (g726) & (!sk[123]) & (g1484) & (g1485) & (g1486)) + ((g677) & (g726) & (sk[123]) & (!g1484) & (g1485) & (!g1486)) + ((g677) & (g726) & (sk[123]) & (!g1484) & (g1485) & (g1486)) + ((g677) & (g726) & (sk[123]) & (g1484) & (g1485) & (!g1486)) + ((g677) & (g726) & (sk[123]) & (g1484) & (g1485) & (g1486)));
	assign g1978 = (((!g1488) & (!g1489) & (!g1490) & (g1491) & (g677) & (g726)) + ((!g1488) & (!g1489) & (g1490) & (!g1491) & (!g677) & (g726)) + ((!g1488) & (!g1489) & (g1490) & (g1491) & (!g677) & (g726)) + ((!g1488) & (!g1489) & (g1490) & (g1491) & (g677) & (g726)) + ((!g1488) & (g1489) & (!g1490) & (!g1491) & (g677) & (!g726)) + ((!g1488) & (g1489) & (!g1490) & (g1491) & (g677) & (!g726)) + ((!g1488) & (g1489) & (!g1490) & (g1491) & (g677) & (g726)) + ((!g1488) & (g1489) & (g1490) & (!g1491) & (!g677) & (g726)) + ((!g1488) & (g1489) & (g1490) & (!g1491) & (g677) & (!g726)) + ((!g1488) & (g1489) & (g1490) & (g1491) & (!g677) & (g726)) + ((!g1488) & (g1489) & (g1490) & (g1491) & (g677) & (!g726)) + ((!g1488) & (g1489) & (g1490) & (g1491) & (g677) & (g726)) + ((g1488) & (!g1489) & (!g1490) & (!g1491) & (!g677) & (!g726)) + ((g1488) & (!g1489) & (!g1490) & (g1491) & (!g677) & (!g726)) + ((g1488) & (!g1489) & (!g1490) & (g1491) & (g677) & (g726)) + ((g1488) & (!g1489) & (g1490) & (!g1491) & (!g677) & (!g726)) + ((g1488) & (!g1489) & (g1490) & (!g1491) & (!g677) & (g726)) + ((g1488) & (!g1489) & (g1490) & (g1491) & (!g677) & (!g726)) + ((g1488) & (!g1489) & (g1490) & (g1491) & (!g677) & (g726)) + ((g1488) & (!g1489) & (g1490) & (g1491) & (g677) & (g726)) + ((g1488) & (g1489) & (!g1490) & (!g1491) & (!g677) & (!g726)) + ((g1488) & (g1489) & (!g1490) & (!g1491) & (g677) & (!g726)) + ((g1488) & (g1489) & (!g1490) & (g1491) & (!g677) & (!g726)) + ((g1488) & (g1489) & (!g1490) & (g1491) & (g677) & (!g726)) + ((g1488) & (g1489) & (!g1490) & (g1491) & (g677) & (g726)) + ((g1488) & (g1489) & (g1490) & (!g1491) & (!g677) & (!g726)) + ((g1488) & (g1489) & (g1490) & (!g1491) & (!g677) & (g726)) + ((g1488) & (g1489) & (g1490) & (!g1491) & (g677) & (!g726)) + ((g1488) & (g1489) & (g1490) & (g1491) & (!g677) & (!g726)) + ((g1488) & (g1489) & (g1490) & (g1491) & (!g677) & (g726)) + ((g1488) & (g1489) & (g1490) & (g1491) & (g677) & (!g726)) + ((g1488) & (g1489) & (g1490) & (g1491) & (g677) & (g726)));
	assign g1979 = (((!g1493) & (!g1494) & (!g1495) & (g1496) & (g677) & (g726)) + ((!g1493) & (!g1494) & (g1495) & (!g1496) & (!g677) & (g726)) + ((!g1493) & (!g1494) & (g1495) & (g1496) & (!g677) & (g726)) + ((!g1493) & (!g1494) & (g1495) & (g1496) & (g677) & (g726)) + ((!g1493) & (g1494) & (!g1495) & (!g1496) & (g677) & (!g726)) + ((!g1493) & (g1494) & (!g1495) & (g1496) & (g677) & (!g726)) + ((!g1493) & (g1494) & (!g1495) & (g1496) & (g677) & (g726)) + ((!g1493) & (g1494) & (g1495) & (!g1496) & (!g677) & (g726)) + ((!g1493) & (g1494) & (g1495) & (!g1496) & (g677) & (!g726)) + ((!g1493) & (g1494) & (g1495) & (g1496) & (!g677) & (g726)) + ((!g1493) & (g1494) & (g1495) & (g1496) & (g677) & (!g726)) + ((!g1493) & (g1494) & (g1495) & (g1496) & (g677) & (g726)) + ((g1493) & (!g1494) & (!g1495) & (!g1496) & (!g677) & (!g726)) + ((g1493) & (!g1494) & (!g1495) & (g1496) & (!g677) & (!g726)) + ((g1493) & (!g1494) & (!g1495) & (g1496) & (g677) & (g726)) + ((g1493) & (!g1494) & (g1495) & (!g1496) & (!g677) & (!g726)) + ((g1493) & (!g1494) & (g1495) & (!g1496) & (!g677) & (g726)) + ((g1493) & (!g1494) & (g1495) & (g1496) & (!g677) & (!g726)) + ((g1493) & (!g1494) & (g1495) & (g1496) & (!g677) & (g726)) + ((g1493) & (!g1494) & (g1495) & (g1496) & (g677) & (g726)) + ((g1493) & (g1494) & (!g1495) & (!g1496) & (!g677) & (!g726)) + ((g1493) & (g1494) & (!g1495) & (!g1496) & (g677) & (!g726)) + ((g1493) & (g1494) & (!g1495) & (g1496) & (!g677) & (!g726)) + ((g1493) & (g1494) & (!g1495) & (g1496) & (g677) & (!g726)) + ((g1493) & (g1494) & (!g1495) & (g1496) & (g677) & (g726)) + ((g1493) & (g1494) & (g1495) & (!g1496) & (!g677) & (!g726)) + ((g1493) & (g1494) & (g1495) & (!g1496) & (!g677) & (g726)) + ((g1493) & (g1494) & (g1495) & (!g1496) & (g677) & (!g726)) + ((g1493) & (g1494) & (g1495) & (g1496) & (!g677) & (!g726)) + ((g1493) & (g1494) & (g1495) & (g1496) & (!g677) & (g726)) + ((g1493) & (g1494) & (g1495) & (g1496) & (g677) & (!g726)) + ((g1493) & (g1494) & (g1495) & (g1496) & (g677) & (g726)));
	assign g1980 = (((!g820) & (!g773) & (!g1976) & (g1977) & (!g1978) & (!g1979)) + ((!g820) & (!g773) & (!g1976) & (g1977) & (!g1978) & (g1979)) + ((!g820) & (!g773) & (!g1976) & (g1977) & (g1978) & (!g1979)) + ((!g820) & (!g773) & (!g1976) & (g1977) & (g1978) & (g1979)) + ((!g820) & (!g773) & (g1976) & (g1977) & (!g1978) & (!g1979)) + ((!g820) & (!g773) & (g1976) & (g1977) & (!g1978) & (g1979)) + ((!g820) & (!g773) & (g1976) & (g1977) & (g1978) & (!g1979)) + ((!g820) & (!g773) & (g1976) & (g1977) & (g1978) & (g1979)) + ((!g820) & (g773) & (!g1976) & (!g1977) & (!g1978) & (g1979)) + ((!g820) & (g773) & (!g1976) & (!g1977) & (g1978) & (g1979)) + ((!g820) & (g773) & (!g1976) & (g1977) & (!g1978) & (g1979)) + ((!g820) & (g773) & (!g1976) & (g1977) & (g1978) & (g1979)) + ((!g820) & (g773) & (g1976) & (!g1977) & (!g1978) & (g1979)) + ((!g820) & (g773) & (g1976) & (!g1977) & (g1978) & (g1979)) + ((!g820) & (g773) & (g1976) & (g1977) & (!g1978) & (g1979)) + ((!g820) & (g773) & (g1976) & (g1977) & (g1978) & (g1979)) + ((g820) & (!g773) & (g1976) & (!g1977) & (!g1978) & (!g1979)) + ((g820) & (!g773) & (g1976) & (!g1977) & (!g1978) & (g1979)) + ((g820) & (!g773) & (g1976) & (!g1977) & (g1978) & (!g1979)) + ((g820) & (!g773) & (g1976) & (!g1977) & (g1978) & (g1979)) + ((g820) & (!g773) & (g1976) & (g1977) & (!g1978) & (!g1979)) + ((g820) & (!g773) & (g1976) & (g1977) & (!g1978) & (g1979)) + ((g820) & (!g773) & (g1976) & (g1977) & (g1978) & (!g1979)) + ((g820) & (!g773) & (g1976) & (g1977) & (g1978) & (g1979)) + ((g820) & (g773) & (!g1976) & (!g1977) & (g1978) & (!g1979)) + ((g820) & (g773) & (!g1976) & (!g1977) & (g1978) & (g1979)) + ((g820) & (g773) & (!g1976) & (g1977) & (g1978) & (!g1979)) + ((g820) & (g773) & (!g1976) & (g1977) & (g1978) & (g1979)) + ((g820) & (g773) & (g1976) & (!g1977) & (g1978) & (!g1979)) + ((g820) & (g773) & (g1976) & (!g1977) & (g1978) & (g1979)) + ((g820) & (g773) & (g1976) & (g1977) & (g1978) & (!g1979)) + ((g820) & (g773) & (g1976) & (g1977) & (g1978) & (g1979)));
	assign g1981 = (((!g867) & (!sk[127]) & (!g1975) & (g1980)) + ((!g867) & (!sk[127]) & (g1975) & (!g1980)) + ((!g867) & (!sk[127]) & (g1975) & (g1980)) + ((!g867) & (sk[127]) & (!g1975) & (g1980)) + ((!g867) & (sk[127]) & (g1975) & (g1980)) + ((g867) & (!sk[127]) & (!g1975) & (g1980)) + ((g867) & (!sk[127]) & (g1975) & (!g1980)) + ((g867) & (!sk[127]) & (g1975) & (g1980)) + ((g867) & (sk[127]) & (g1975) & (!g1980)) + ((g867) & (sk[127]) & (g1975) & (g1980)));
	assign g1982 = (((!g1593) & (!g1605) & (!sk[0]) & (!g1772) & (g64)) + ((!g1593) & (!g1605) & (!sk[0]) & (g1772) & (!g64)) + ((!g1593) & (!g1605) & (!sk[0]) & (g1772) & (g64)) + ((!g1593) & (!g1605) & (sk[0]) & (g1772) & (!g64)) + ((!g1593) & (!g1605) & (sk[0]) & (g1772) & (g64)) + ((!g1593) & (g1605) & (!sk[0]) & (!g1772) & (!g64)) + ((!g1593) & (g1605) & (!sk[0]) & (!g1772) & (g64)) + ((!g1593) & (g1605) & (!sk[0]) & (g1772) & (!g64)) + ((!g1593) & (g1605) & (!sk[0]) & (g1772) & (g64)) + ((g1593) & (!g1605) & (!sk[0]) & (!g1772) & (g64)) + ((g1593) & (!g1605) & (!sk[0]) & (g1772) & (!g64)) + ((g1593) & (!g1605) & (!sk[0]) & (g1772) & (g64)) + ((g1593) & (!g1605) & (sk[0]) & (!g1772) & (g64)) + ((g1593) & (!g1605) & (sk[0]) & (g1772) & (g64)) + ((g1593) & (g1605) & (!sk[0]) & (!g1772) & (!g64)) + ((g1593) & (g1605) & (!sk[0]) & (!g1772) & (g64)) + ((g1593) & (g1605) & (!sk[0]) & (g1772) & (!g64)) + ((g1593) & (g1605) & (!sk[0]) & (g1772) & (g64)) + ((g1593) & (g1605) & (sk[0]) & (!g1772) & (g64)) + ((g1593) & (g1605) & (sk[0]) & (g1772) & (g64)));
	assign g1983 = (((!g132) & (!g1592) & (g1668) & (g1917) & (!g1981) & (!g1982)) + ((!g132) & (!g1592) & (g1668) & (g1917) & (!g1981) & (g1982)) + ((!g132) & (!g1592) & (g1668) & (g1917) & (g1981) & (!g1982)) + ((!g132) & (!g1592) & (g1668) & (g1917) & (g1981) & (g1982)) + ((!g132) & (g1592) & (!g1668) & (g1917) & (!g1981) & (g1982)) + ((!g132) & (g1592) & (!g1668) & (g1917) & (g1981) & (g1982)) + ((!g132) & (g1592) & (g1668) & (g1917) & (!g1981) & (g1982)) + ((!g132) & (g1592) & (g1668) & (g1917) & (g1981) & (g1982)) + ((g132) & (!g1592) & (!g1668) & (g1917) & (g1981) & (!g1982)) + ((g132) & (!g1592) & (!g1668) & (g1917) & (g1981) & (g1982)) + ((g132) & (!g1592) & (g1668) & (g1917) & (g1981) & (!g1982)) + ((g132) & (!g1592) & (g1668) & (g1917) & (g1981) & (g1982)) + ((g132) & (g1592) & (!g1668) & (g1917) & (g1981) & (!g1982)) + ((g132) & (g1592) & (!g1668) & (g1917) & (g1981) & (g1982)) + ((g132) & (g1592) & (g1668) & (g1917) & (g1981) & (!g1982)) + ((g132) & (g1592) & (g1668) & (g1917) & (g1981) & (g1982)));
	assign g1984 = (((!g1502) & (!g1507) & (!g1512) & (g1517) & (g677) & (g726)) + ((!g1502) & (!g1507) & (g1512) & (!g1517) & (!g677) & (g726)) + ((!g1502) & (!g1507) & (g1512) & (g1517) & (!g677) & (g726)) + ((!g1502) & (!g1507) & (g1512) & (g1517) & (g677) & (g726)) + ((!g1502) & (g1507) & (!g1512) & (!g1517) & (g677) & (!g726)) + ((!g1502) & (g1507) & (!g1512) & (g1517) & (g677) & (!g726)) + ((!g1502) & (g1507) & (!g1512) & (g1517) & (g677) & (g726)) + ((!g1502) & (g1507) & (g1512) & (!g1517) & (!g677) & (g726)) + ((!g1502) & (g1507) & (g1512) & (!g1517) & (g677) & (!g726)) + ((!g1502) & (g1507) & (g1512) & (g1517) & (!g677) & (g726)) + ((!g1502) & (g1507) & (g1512) & (g1517) & (g677) & (!g726)) + ((!g1502) & (g1507) & (g1512) & (g1517) & (g677) & (g726)) + ((g1502) & (!g1507) & (!g1512) & (!g1517) & (!g677) & (!g726)) + ((g1502) & (!g1507) & (!g1512) & (g1517) & (!g677) & (!g726)) + ((g1502) & (!g1507) & (!g1512) & (g1517) & (g677) & (g726)) + ((g1502) & (!g1507) & (g1512) & (!g1517) & (!g677) & (!g726)) + ((g1502) & (!g1507) & (g1512) & (!g1517) & (!g677) & (g726)) + ((g1502) & (!g1507) & (g1512) & (g1517) & (!g677) & (!g726)) + ((g1502) & (!g1507) & (g1512) & (g1517) & (!g677) & (g726)) + ((g1502) & (!g1507) & (g1512) & (g1517) & (g677) & (g726)) + ((g1502) & (g1507) & (!g1512) & (!g1517) & (!g677) & (!g726)) + ((g1502) & (g1507) & (!g1512) & (!g1517) & (g677) & (!g726)) + ((g1502) & (g1507) & (!g1512) & (g1517) & (!g677) & (!g726)) + ((g1502) & (g1507) & (!g1512) & (g1517) & (g677) & (!g726)) + ((g1502) & (g1507) & (!g1512) & (g1517) & (g677) & (g726)) + ((g1502) & (g1507) & (g1512) & (!g1517) & (!g677) & (!g726)) + ((g1502) & (g1507) & (g1512) & (!g1517) & (!g677) & (g726)) + ((g1502) & (g1507) & (g1512) & (!g1517) & (g677) & (!g726)) + ((g1502) & (g1507) & (g1512) & (g1517) & (!g677) & (!g726)) + ((g1502) & (g1507) & (g1512) & (g1517) & (!g677) & (g726)) + ((g1502) & (g1507) & (g1512) & (g1517) & (g677) & (!g726)) + ((g1502) & (g1507) & (g1512) & (g1517) & (g677) & (g726)));
	assign g1985 = (((!g1503) & (!g1508) & (!g1513) & (g1518) & (g677) & (g726)) + ((!g1503) & (!g1508) & (g1513) & (!g1518) & (!g677) & (g726)) + ((!g1503) & (!g1508) & (g1513) & (g1518) & (!g677) & (g726)) + ((!g1503) & (!g1508) & (g1513) & (g1518) & (g677) & (g726)) + ((!g1503) & (g1508) & (!g1513) & (!g1518) & (g677) & (!g726)) + ((!g1503) & (g1508) & (!g1513) & (g1518) & (g677) & (!g726)) + ((!g1503) & (g1508) & (!g1513) & (g1518) & (g677) & (g726)) + ((!g1503) & (g1508) & (g1513) & (!g1518) & (!g677) & (g726)) + ((!g1503) & (g1508) & (g1513) & (!g1518) & (g677) & (!g726)) + ((!g1503) & (g1508) & (g1513) & (g1518) & (!g677) & (g726)) + ((!g1503) & (g1508) & (g1513) & (g1518) & (g677) & (!g726)) + ((!g1503) & (g1508) & (g1513) & (g1518) & (g677) & (g726)) + ((g1503) & (!g1508) & (!g1513) & (!g1518) & (!g677) & (!g726)) + ((g1503) & (!g1508) & (!g1513) & (g1518) & (!g677) & (!g726)) + ((g1503) & (!g1508) & (!g1513) & (g1518) & (g677) & (g726)) + ((g1503) & (!g1508) & (g1513) & (!g1518) & (!g677) & (!g726)) + ((g1503) & (!g1508) & (g1513) & (!g1518) & (!g677) & (g726)) + ((g1503) & (!g1508) & (g1513) & (g1518) & (!g677) & (!g726)) + ((g1503) & (!g1508) & (g1513) & (g1518) & (!g677) & (g726)) + ((g1503) & (!g1508) & (g1513) & (g1518) & (g677) & (g726)) + ((g1503) & (g1508) & (!g1513) & (!g1518) & (!g677) & (!g726)) + ((g1503) & (g1508) & (!g1513) & (!g1518) & (g677) & (!g726)) + ((g1503) & (g1508) & (!g1513) & (g1518) & (!g677) & (!g726)) + ((g1503) & (g1508) & (!g1513) & (g1518) & (g677) & (!g726)) + ((g1503) & (g1508) & (!g1513) & (g1518) & (g677) & (g726)) + ((g1503) & (g1508) & (g1513) & (!g1518) & (!g677) & (!g726)) + ((g1503) & (g1508) & (g1513) & (!g1518) & (!g677) & (g726)) + ((g1503) & (g1508) & (g1513) & (!g1518) & (g677) & (!g726)) + ((g1503) & (g1508) & (g1513) & (g1518) & (!g677) & (!g726)) + ((g1503) & (g1508) & (g1513) & (g1518) & (!g677) & (g726)) + ((g1503) & (g1508) & (g1513) & (g1518) & (g677) & (!g726)) + ((g1503) & (g1508) & (g1513) & (g1518) & (g677) & (g726)));
	assign g1986 = (((!g1504) & (!g1509) & (!g1514) & (g1519) & (g677) & (g726)) + ((!g1504) & (!g1509) & (g1514) & (!g1519) & (!g677) & (g726)) + ((!g1504) & (!g1509) & (g1514) & (g1519) & (!g677) & (g726)) + ((!g1504) & (!g1509) & (g1514) & (g1519) & (g677) & (g726)) + ((!g1504) & (g1509) & (!g1514) & (!g1519) & (g677) & (!g726)) + ((!g1504) & (g1509) & (!g1514) & (g1519) & (g677) & (!g726)) + ((!g1504) & (g1509) & (!g1514) & (g1519) & (g677) & (g726)) + ((!g1504) & (g1509) & (g1514) & (!g1519) & (!g677) & (g726)) + ((!g1504) & (g1509) & (g1514) & (!g1519) & (g677) & (!g726)) + ((!g1504) & (g1509) & (g1514) & (g1519) & (!g677) & (g726)) + ((!g1504) & (g1509) & (g1514) & (g1519) & (g677) & (!g726)) + ((!g1504) & (g1509) & (g1514) & (g1519) & (g677) & (g726)) + ((g1504) & (!g1509) & (!g1514) & (!g1519) & (!g677) & (!g726)) + ((g1504) & (!g1509) & (!g1514) & (g1519) & (!g677) & (!g726)) + ((g1504) & (!g1509) & (!g1514) & (g1519) & (g677) & (g726)) + ((g1504) & (!g1509) & (g1514) & (!g1519) & (!g677) & (!g726)) + ((g1504) & (!g1509) & (g1514) & (!g1519) & (!g677) & (g726)) + ((g1504) & (!g1509) & (g1514) & (g1519) & (!g677) & (!g726)) + ((g1504) & (!g1509) & (g1514) & (g1519) & (!g677) & (g726)) + ((g1504) & (!g1509) & (g1514) & (g1519) & (g677) & (g726)) + ((g1504) & (g1509) & (!g1514) & (!g1519) & (!g677) & (!g726)) + ((g1504) & (g1509) & (!g1514) & (!g1519) & (g677) & (!g726)) + ((g1504) & (g1509) & (!g1514) & (g1519) & (!g677) & (!g726)) + ((g1504) & (g1509) & (!g1514) & (g1519) & (g677) & (!g726)) + ((g1504) & (g1509) & (!g1514) & (g1519) & (g677) & (g726)) + ((g1504) & (g1509) & (g1514) & (!g1519) & (!g677) & (!g726)) + ((g1504) & (g1509) & (g1514) & (!g1519) & (!g677) & (g726)) + ((g1504) & (g1509) & (g1514) & (!g1519) & (g677) & (!g726)) + ((g1504) & (g1509) & (g1514) & (g1519) & (!g677) & (!g726)) + ((g1504) & (g1509) & (g1514) & (g1519) & (!g677) & (g726)) + ((g1504) & (g1509) & (g1514) & (g1519) & (g677) & (!g726)) + ((g1504) & (g1509) & (g1514) & (g1519) & (g677) & (g726)));
	assign g1987 = (((!g1505) & (!g1510) & (!g1515) & (g1520) & (g677) & (g726)) + ((!g1505) & (!g1510) & (g1515) & (!g1520) & (!g677) & (g726)) + ((!g1505) & (!g1510) & (g1515) & (g1520) & (!g677) & (g726)) + ((!g1505) & (!g1510) & (g1515) & (g1520) & (g677) & (g726)) + ((!g1505) & (g1510) & (!g1515) & (!g1520) & (g677) & (!g726)) + ((!g1505) & (g1510) & (!g1515) & (g1520) & (g677) & (!g726)) + ((!g1505) & (g1510) & (!g1515) & (g1520) & (g677) & (g726)) + ((!g1505) & (g1510) & (g1515) & (!g1520) & (!g677) & (g726)) + ((!g1505) & (g1510) & (g1515) & (!g1520) & (g677) & (!g726)) + ((!g1505) & (g1510) & (g1515) & (g1520) & (!g677) & (g726)) + ((!g1505) & (g1510) & (g1515) & (g1520) & (g677) & (!g726)) + ((!g1505) & (g1510) & (g1515) & (g1520) & (g677) & (g726)) + ((g1505) & (!g1510) & (!g1515) & (!g1520) & (!g677) & (!g726)) + ((g1505) & (!g1510) & (!g1515) & (g1520) & (!g677) & (!g726)) + ((g1505) & (!g1510) & (!g1515) & (g1520) & (g677) & (g726)) + ((g1505) & (!g1510) & (g1515) & (!g1520) & (!g677) & (!g726)) + ((g1505) & (!g1510) & (g1515) & (!g1520) & (!g677) & (g726)) + ((g1505) & (!g1510) & (g1515) & (g1520) & (!g677) & (!g726)) + ((g1505) & (!g1510) & (g1515) & (g1520) & (!g677) & (g726)) + ((g1505) & (!g1510) & (g1515) & (g1520) & (g677) & (g726)) + ((g1505) & (g1510) & (!g1515) & (!g1520) & (!g677) & (!g726)) + ((g1505) & (g1510) & (!g1515) & (!g1520) & (g677) & (!g726)) + ((g1505) & (g1510) & (!g1515) & (g1520) & (!g677) & (!g726)) + ((g1505) & (g1510) & (!g1515) & (g1520) & (g677) & (!g726)) + ((g1505) & (g1510) & (!g1515) & (g1520) & (g677) & (g726)) + ((g1505) & (g1510) & (g1515) & (!g1520) & (!g677) & (!g726)) + ((g1505) & (g1510) & (g1515) & (!g1520) & (!g677) & (g726)) + ((g1505) & (g1510) & (g1515) & (!g1520) & (g677) & (!g726)) + ((g1505) & (g1510) & (g1515) & (g1520) & (!g677) & (!g726)) + ((g1505) & (g1510) & (g1515) & (g1520) & (!g677) & (g726)) + ((g1505) & (g1510) & (g1515) & (g1520) & (g677) & (!g726)) + ((g1505) & (g1510) & (g1515) & (g1520) & (g677) & (g726)));
	assign g1988 = (((!g1984) & (!g1985) & (!g1986) & (g1987) & (g820) & (g773)) + ((!g1984) & (!g1985) & (g1986) & (!g1987) & (!g820) & (g773)) + ((!g1984) & (!g1985) & (g1986) & (g1987) & (!g820) & (g773)) + ((!g1984) & (!g1985) & (g1986) & (g1987) & (g820) & (g773)) + ((!g1984) & (g1985) & (!g1986) & (!g1987) & (g820) & (!g773)) + ((!g1984) & (g1985) & (!g1986) & (g1987) & (g820) & (!g773)) + ((!g1984) & (g1985) & (!g1986) & (g1987) & (g820) & (g773)) + ((!g1984) & (g1985) & (g1986) & (!g1987) & (!g820) & (g773)) + ((!g1984) & (g1985) & (g1986) & (!g1987) & (g820) & (!g773)) + ((!g1984) & (g1985) & (g1986) & (g1987) & (!g820) & (g773)) + ((!g1984) & (g1985) & (g1986) & (g1987) & (g820) & (!g773)) + ((!g1984) & (g1985) & (g1986) & (g1987) & (g820) & (g773)) + ((g1984) & (!g1985) & (!g1986) & (!g1987) & (!g820) & (!g773)) + ((g1984) & (!g1985) & (!g1986) & (g1987) & (!g820) & (!g773)) + ((g1984) & (!g1985) & (!g1986) & (g1987) & (g820) & (g773)) + ((g1984) & (!g1985) & (g1986) & (!g1987) & (!g820) & (!g773)) + ((g1984) & (!g1985) & (g1986) & (!g1987) & (!g820) & (g773)) + ((g1984) & (!g1985) & (g1986) & (g1987) & (!g820) & (!g773)) + ((g1984) & (!g1985) & (g1986) & (g1987) & (!g820) & (g773)) + ((g1984) & (!g1985) & (g1986) & (g1987) & (g820) & (g773)) + ((g1984) & (g1985) & (!g1986) & (!g1987) & (!g820) & (!g773)) + ((g1984) & (g1985) & (!g1986) & (!g1987) & (g820) & (!g773)) + ((g1984) & (g1985) & (!g1986) & (g1987) & (!g820) & (!g773)) + ((g1984) & (g1985) & (!g1986) & (g1987) & (g820) & (!g773)) + ((g1984) & (g1985) & (!g1986) & (g1987) & (g820) & (g773)) + ((g1984) & (g1985) & (g1986) & (!g1987) & (!g820) & (!g773)) + ((g1984) & (g1985) & (g1986) & (!g1987) & (!g820) & (g773)) + ((g1984) & (g1985) & (g1986) & (!g1987) & (g820) & (!g773)) + ((g1984) & (g1985) & (g1986) & (g1987) & (!g820) & (!g773)) + ((g1984) & (g1985) & (g1986) & (g1987) & (!g820) & (g773)) + ((g1984) & (g1985) & (g1986) & (g1987) & (g820) & (!g773)) + ((g1984) & (g1985) & (g1986) & (g1987) & (g820) & (g773)));
	assign g1989 = (((!g1523) & (!g1524) & (!g1525) & (g1526) & (g677) & (g726)) + ((!g1523) & (!g1524) & (g1525) & (!g1526) & (!g677) & (g726)) + ((!g1523) & (!g1524) & (g1525) & (g1526) & (!g677) & (g726)) + ((!g1523) & (!g1524) & (g1525) & (g1526) & (g677) & (g726)) + ((!g1523) & (g1524) & (!g1525) & (!g1526) & (g677) & (!g726)) + ((!g1523) & (g1524) & (!g1525) & (g1526) & (g677) & (!g726)) + ((!g1523) & (g1524) & (!g1525) & (g1526) & (g677) & (g726)) + ((!g1523) & (g1524) & (g1525) & (!g1526) & (!g677) & (g726)) + ((!g1523) & (g1524) & (g1525) & (!g1526) & (g677) & (!g726)) + ((!g1523) & (g1524) & (g1525) & (g1526) & (!g677) & (g726)) + ((!g1523) & (g1524) & (g1525) & (g1526) & (g677) & (!g726)) + ((!g1523) & (g1524) & (g1525) & (g1526) & (g677) & (g726)) + ((g1523) & (!g1524) & (!g1525) & (!g1526) & (!g677) & (!g726)) + ((g1523) & (!g1524) & (!g1525) & (g1526) & (!g677) & (!g726)) + ((g1523) & (!g1524) & (!g1525) & (g1526) & (g677) & (g726)) + ((g1523) & (!g1524) & (g1525) & (!g1526) & (!g677) & (!g726)) + ((g1523) & (!g1524) & (g1525) & (!g1526) & (!g677) & (g726)) + ((g1523) & (!g1524) & (g1525) & (g1526) & (!g677) & (!g726)) + ((g1523) & (!g1524) & (g1525) & (g1526) & (!g677) & (g726)) + ((g1523) & (!g1524) & (g1525) & (g1526) & (g677) & (g726)) + ((g1523) & (g1524) & (!g1525) & (!g1526) & (!g677) & (!g726)) + ((g1523) & (g1524) & (!g1525) & (!g1526) & (g677) & (!g726)) + ((g1523) & (g1524) & (!g1525) & (g1526) & (!g677) & (!g726)) + ((g1523) & (g1524) & (!g1525) & (g1526) & (g677) & (!g726)) + ((g1523) & (g1524) & (!g1525) & (g1526) & (g677) & (g726)) + ((g1523) & (g1524) & (g1525) & (!g1526) & (!g677) & (!g726)) + ((g1523) & (g1524) & (g1525) & (!g1526) & (!g677) & (g726)) + ((g1523) & (g1524) & (g1525) & (!g1526) & (g677) & (!g726)) + ((g1523) & (g1524) & (g1525) & (g1526) & (!g677) & (!g726)) + ((g1523) & (g1524) & (g1525) & (g1526) & (!g677) & (g726)) + ((g1523) & (g1524) & (g1525) & (g1526) & (g677) & (!g726)) + ((g1523) & (g1524) & (g1525) & (g1526) & (g677) & (g726)));
	assign g1990 = (((!g677) & (!g726) & (!g1528) & (g1529) & (!sk[8]) & (!g1530)) + ((!g677) & (!g726) & (!g1528) & (g1529) & (!sk[8]) & (g1530)) + ((!g677) & (!g726) & (g1528) & (!g1529) & (!sk[8]) & (!g1530)) + ((!g677) & (!g726) & (g1528) & (!g1529) & (!sk[8]) & (g1530)) + ((!g677) & (!g726) & (g1528) & (g1529) & (!sk[8]) & (!g1530)) + ((!g677) & (!g726) & (g1528) & (g1529) & (!sk[8]) & (g1530)) + ((!g677) & (g726) & (!g1528) & (!g1529) & (!sk[8]) & (!g1530)) + ((!g677) & (g726) & (!g1528) & (!g1529) & (!sk[8]) & (g1530)) + ((!g677) & (g726) & (!g1528) & (!g1529) & (sk[8]) & (g1530)) + ((!g677) & (g726) & (!g1528) & (g1529) & (!sk[8]) & (!g1530)) + ((!g677) & (g726) & (!g1528) & (g1529) & (!sk[8]) & (g1530)) + ((!g677) & (g726) & (!g1528) & (g1529) & (sk[8]) & (g1530)) + ((!g677) & (g726) & (g1528) & (!g1529) & (!sk[8]) & (!g1530)) + ((!g677) & (g726) & (g1528) & (!g1529) & (!sk[8]) & (g1530)) + ((!g677) & (g726) & (g1528) & (!g1529) & (sk[8]) & (g1530)) + ((!g677) & (g726) & (g1528) & (g1529) & (!sk[8]) & (!g1530)) + ((!g677) & (g726) & (g1528) & (g1529) & (!sk[8]) & (g1530)) + ((!g677) & (g726) & (g1528) & (g1529) & (sk[8]) & (g1530)) + ((g677) & (!g726) & (!g1528) & (g1529) & (!sk[8]) & (!g1530)) + ((g677) & (!g726) & (!g1528) & (g1529) & (!sk[8]) & (g1530)) + ((g677) & (!g726) & (g1528) & (!g1529) & (!sk[8]) & (!g1530)) + ((g677) & (!g726) & (g1528) & (!g1529) & (!sk[8]) & (g1530)) + ((g677) & (!g726) & (g1528) & (!g1529) & (sk[8]) & (!g1530)) + ((g677) & (!g726) & (g1528) & (!g1529) & (sk[8]) & (g1530)) + ((g677) & (!g726) & (g1528) & (g1529) & (!sk[8]) & (!g1530)) + ((g677) & (!g726) & (g1528) & (g1529) & (!sk[8]) & (g1530)) + ((g677) & (!g726) & (g1528) & (g1529) & (sk[8]) & (!g1530)) + ((g677) & (!g726) & (g1528) & (g1529) & (sk[8]) & (g1530)) + ((g677) & (g726) & (!g1528) & (!g1529) & (!sk[8]) & (!g1530)) + ((g677) & (g726) & (!g1528) & (!g1529) & (!sk[8]) & (g1530)) + ((g677) & (g726) & (!g1528) & (g1529) & (!sk[8]) & (!g1530)) + ((g677) & (g726) & (!g1528) & (g1529) & (!sk[8]) & (g1530)) + ((g677) & (g726) & (!g1528) & (g1529) & (sk[8]) & (!g1530)) + ((g677) & (g726) & (!g1528) & (g1529) & (sk[8]) & (g1530)) + ((g677) & (g726) & (g1528) & (!g1529) & (!sk[8]) & (!g1530)) + ((g677) & (g726) & (g1528) & (!g1529) & (!sk[8]) & (g1530)) + ((g677) & (g726) & (g1528) & (g1529) & (!sk[8]) & (!g1530)) + ((g677) & (g726) & (g1528) & (g1529) & (!sk[8]) & (g1530)) + ((g677) & (g726) & (g1528) & (g1529) & (sk[8]) & (!g1530)) + ((g677) & (g726) & (g1528) & (g1529) & (sk[8]) & (g1530)));
	assign g1991 = (((!g1532) & (!g1533) & (!g1534) & (g1535) & (g677) & (g726)) + ((!g1532) & (!g1533) & (g1534) & (!g1535) & (!g677) & (g726)) + ((!g1532) & (!g1533) & (g1534) & (g1535) & (!g677) & (g726)) + ((!g1532) & (!g1533) & (g1534) & (g1535) & (g677) & (g726)) + ((!g1532) & (g1533) & (!g1534) & (!g1535) & (g677) & (!g726)) + ((!g1532) & (g1533) & (!g1534) & (g1535) & (g677) & (!g726)) + ((!g1532) & (g1533) & (!g1534) & (g1535) & (g677) & (g726)) + ((!g1532) & (g1533) & (g1534) & (!g1535) & (!g677) & (g726)) + ((!g1532) & (g1533) & (g1534) & (!g1535) & (g677) & (!g726)) + ((!g1532) & (g1533) & (g1534) & (g1535) & (!g677) & (g726)) + ((!g1532) & (g1533) & (g1534) & (g1535) & (g677) & (!g726)) + ((!g1532) & (g1533) & (g1534) & (g1535) & (g677) & (g726)) + ((g1532) & (!g1533) & (!g1534) & (!g1535) & (!g677) & (!g726)) + ((g1532) & (!g1533) & (!g1534) & (g1535) & (!g677) & (!g726)) + ((g1532) & (!g1533) & (!g1534) & (g1535) & (g677) & (g726)) + ((g1532) & (!g1533) & (g1534) & (!g1535) & (!g677) & (!g726)) + ((g1532) & (!g1533) & (g1534) & (!g1535) & (!g677) & (g726)) + ((g1532) & (!g1533) & (g1534) & (g1535) & (!g677) & (!g726)) + ((g1532) & (!g1533) & (g1534) & (g1535) & (!g677) & (g726)) + ((g1532) & (!g1533) & (g1534) & (g1535) & (g677) & (g726)) + ((g1532) & (g1533) & (!g1534) & (!g1535) & (!g677) & (!g726)) + ((g1532) & (g1533) & (!g1534) & (!g1535) & (g677) & (!g726)) + ((g1532) & (g1533) & (!g1534) & (g1535) & (!g677) & (!g726)) + ((g1532) & (g1533) & (!g1534) & (g1535) & (g677) & (!g726)) + ((g1532) & (g1533) & (!g1534) & (g1535) & (g677) & (g726)) + ((g1532) & (g1533) & (g1534) & (!g1535) & (!g677) & (!g726)) + ((g1532) & (g1533) & (g1534) & (!g1535) & (!g677) & (g726)) + ((g1532) & (g1533) & (g1534) & (!g1535) & (g677) & (!g726)) + ((g1532) & (g1533) & (g1534) & (g1535) & (!g677) & (!g726)) + ((g1532) & (g1533) & (g1534) & (g1535) & (!g677) & (g726)) + ((g1532) & (g1533) & (g1534) & (g1535) & (g677) & (!g726)) + ((g1532) & (g1533) & (g1534) & (g1535) & (g677) & (g726)));
	assign g1992 = (((!g1537) & (!g1538) & (!g1539) & (g1540) & (g677) & (g726)) + ((!g1537) & (!g1538) & (g1539) & (!g1540) & (!g677) & (g726)) + ((!g1537) & (!g1538) & (g1539) & (g1540) & (!g677) & (g726)) + ((!g1537) & (!g1538) & (g1539) & (g1540) & (g677) & (g726)) + ((!g1537) & (g1538) & (!g1539) & (!g1540) & (g677) & (!g726)) + ((!g1537) & (g1538) & (!g1539) & (g1540) & (g677) & (!g726)) + ((!g1537) & (g1538) & (!g1539) & (g1540) & (g677) & (g726)) + ((!g1537) & (g1538) & (g1539) & (!g1540) & (!g677) & (g726)) + ((!g1537) & (g1538) & (g1539) & (!g1540) & (g677) & (!g726)) + ((!g1537) & (g1538) & (g1539) & (g1540) & (!g677) & (g726)) + ((!g1537) & (g1538) & (g1539) & (g1540) & (g677) & (!g726)) + ((!g1537) & (g1538) & (g1539) & (g1540) & (g677) & (g726)) + ((g1537) & (!g1538) & (!g1539) & (!g1540) & (!g677) & (!g726)) + ((g1537) & (!g1538) & (!g1539) & (g1540) & (!g677) & (!g726)) + ((g1537) & (!g1538) & (!g1539) & (g1540) & (g677) & (g726)) + ((g1537) & (!g1538) & (g1539) & (!g1540) & (!g677) & (!g726)) + ((g1537) & (!g1538) & (g1539) & (!g1540) & (!g677) & (g726)) + ((g1537) & (!g1538) & (g1539) & (g1540) & (!g677) & (!g726)) + ((g1537) & (!g1538) & (g1539) & (g1540) & (!g677) & (g726)) + ((g1537) & (!g1538) & (g1539) & (g1540) & (g677) & (g726)) + ((g1537) & (g1538) & (!g1539) & (!g1540) & (!g677) & (!g726)) + ((g1537) & (g1538) & (!g1539) & (!g1540) & (g677) & (!g726)) + ((g1537) & (g1538) & (!g1539) & (g1540) & (!g677) & (!g726)) + ((g1537) & (g1538) & (!g1539) & (g1540) & (g677) & (!g726)) + ((g1537) & (g1538) & (!g1539) & (g1540) & (g677) & (g726)) + ((g1537) & (g1538) & (g1539) & (!g1540) & (!g677) & (!g726)) + ((g1537) & (g1538) & (g1539) & (!g1540) & (!g677) & (g726)) + ((g1537) & (g1538) & (g1539) & (!g1540) & (g677) & (!g726)) + ((g1537) & (g1538) & (g1539) & (g1540) & (!g677) & (!g726)) + ((g1537) & (g1538) & (g1539) & (g1540) & (!g677) & (g726)) + ((g1537) & (g1538) & (g1539) & (g1540) & (g677) & (!g726)) + ((g1537) & (g1538) & (g1539) & (g1540) & (g677) & (g726)));
	assign g1993 = (((!g820) & (!g773) & (!g1989) & (g1990) & (!g1991) & (!g1992)) + ((!g820) & (!g773) & (!g1989) & (g1990) & (!g1991) & (g1992)) + ((!g820) & (!g773) & (!g1989) & (g1990) & (g1991) & (!g1992)) + ((!g820) & (!g773) & (!g1989) & (g1990) & (g1991) & (g1992)) + ((!g820) & (!g773) & (g1989) & (g1990) & (!g1991) & (!g1992)) + ((!g820) & (!g773) & (g1989) & (g1990) & (!g1991) & (g1992)) + ((!g820) & (!g773) & (g1989) & (g1990) & (g1991) & (!g1992)) + ((!g820) & (!g773) & (g1989) & (g1990) & (g1991) & (g1992)) + ((!g820) & (g773) & (!g1989) & (!g1990) & (!g1991) & (g1992)) + ((!g820) & (g773) & (!g1989) & (!g1990) & (g1991) & (g1992)) + ((!g820) & (g773) & (!g1989) & (g1990) & (!g1991) & (g1992)) + ((!g820) & (g773) & (!g1989) & (g1990) & (g1991) & (g1992)) + ((!g820) & (g773) & (g1989) & (!g1990) & (!g1991) & (g1992)) + ((!g820) & (g773) & (g1989) & (!g1990) & (g1991) & (g1992)) + ((!g820) & (g773) & (g1989) & (g1990) & (!g1991) & (g1992)) + ((!g820) & (g773) & (g1989) & (g1990) & (g1991) & (g1992)) + ((g820) & (!g773) & (g1989) & (!g1990) & (!g1991) & (!g1992)) + ((g820) & (!g773) & (g1989) & (!g1990) & (!g1991) & (g1992)) + ((g820) & (!g773) & (g1989) & (!g1990) & (g1991) & (!g1992)) + ((g820) & (!g773) & (g1989) & (!g1990) & (g1991) & (g1992)) + ((g820) & (!g773) & (g1989) & (g1990) & (!g1991) & (!g1992)) + ((g820) & (!g773) & (g1989) & (g1990) & (!g1991) & (g1992)) + ((g820) & (!g773) & (g1989) & (g1990) & (g1991) & (!g1992)) + ((g820) & (!g773) & (g1989) & (g1990) & (g1991) & (g1992)) + ((g820) & (g773) & (!g1989) & (!g1990) & (g1991) & (!g1992)) + ((g820) & (g773) & (!g1989) & (!g1990) & (g1991) & (g1992)) + ((g820) & (g773) & (!g1989) & (g1990) & (g1991) & (!g1992)) + ((g820) & (g773) & (!g1989) & (g1990) & (g1991) & (g1992)) + ((g820) & (g773) & (g1989) & (!g1990) & (g1991) & (!g1992)) + ((g820) & (g773) & (g1989) & (!g1990) & (g1991) & (g1992)) + ((g820) & (g773) & (g1989) & (g1990) & (g1991) & (!g1992)) + ((g820) & (g773) & (g1989) & (g1990) & (g1991) & (g1992)));
	assign g1994 = (((!sk[12]) & (!g867) & (!g1988) & (g1993)) + ((!sk[12]) & (!g867) & (g1988) & (!g1993)) + ((!sk[12]) & (!g867) & (g1988) & (g1993)) + ((!sk[12]) & (g867) & (!g1988) & (g1993)) + ((!sk[12]) & (g867) & (g1988) & (!g1993)) + ((!sk[12]) & (g867) & (g1988) & (g1993)) + ((sk[12]) & (!g867) & (!g1988) & (g1993)) + ((sk[12]) & (!g867) & (g1988) & (g1993)) + ((sk[12]) & (g867) & (g1988) & (!g1993)) + ((sk[12]) & (g867) & (g1988) & (g1993)));
	assign g1995 = (((!g1593) & (!sk[13]) & (!g1605) & (!g1785) & (g65)) + ((!g1593) & (!sk[13]) & (!g1605) & (g1785) & (!g65)) + ((!g1593) & (!sk[13]) & (!g1605) & (g1785) & (g65)) + ((!g1593) & (!sk[13]) & (g1605) & (!g1785) & (!g65)) + ((!g1593) & (!sk[13]) & (g1605) & (!g1785) & (g65)) + ((!g1593) & (!sk[13]) & (g1605) & (g1785) & (!g65)) + ((!g1593) & (!sk[13]) & (g1605) & (g1785) & (g65)) + ((!g1593) & (sk[13]) & (!g1605) & (g1785) & (!g65)) + ((!g1593) & (sk[13]) & (!g1605) & (g1785) & (g65)) + ((g1593) & (!sk[13]) & (!g1605) & (!g1785) & (g65)) + ((g1593) & (!sk[13]) & (!g1605) & (g1785) & (!g65)) + ((g1593) & (!sk[13]) & (!g1605) & (g1785) & (g65)) + ((g1593) & (!sk[13]) & (g1605) & (!g1785) & (!g65)) + ((g1593) & (!sk[13]) & (g1605) & (!g1785) & (g65)) + ((g1593) & (!sk[13]) & (g1605) & (g1785) & (!g65)) + ((g1593) & (!sk[13]) & (g1605) & (g1785) & (g65)) + ((g1593) & (sk[13]) & (!g1605) & (!g1785) & (g65)) + ((g1593) & (sk[13]) & (!g1605) & (g1785) & (g65)) + ((g1593) & (sk[13]) & (g1605) & (!g1785) & (g65)) + ((g1593) & (sk[13]) & (g1605) & (g1785) & (g65)));
	assign g1996 = (((!g132) & (!g1592) & (g1680) & (g1917) & (!g1994) & (!g1995)) + ((!g132) & (!g1592) & (g1680) & (g1917) & (!g1994) & (g1995)) + ((!g132) & (!g1592) & (g1680) & (g1917) & (g1994) & (!g1995)) + ((!g132) & (!g1592) & (g1680) & (g1917) & (g1994) & (g1995)) + ((!g132) & (g1592) & (!g1680) & (g1917) & (!g1994) & (g1995)) + ((!g132) & (g1592) & (!g1680) & (g1917) & (g1994) & (g1995)) + ((!g132) & (g1592) & (g1680) & (g1917) & (!g1994) & (g1995)) + ((!g132) & (g1592) & (g1680) & (g1917) & (g1994) & (g1995)) + ((g132) & (!g1592) & (!g1680) & (g1917) & (g1994) & (!g1995)) + ((g132) & (!g1592) & (!g1680) & (g1917) & (g1994) & (g1995)) + ((g132) & (!g1592) & (g1680) & (g1917) & (g1994) & (!g1995)) + ((g132) & (!g1592) & (g1680) & (g1917) & (g1994) & (g1995)) + ((g132) & (g1592) & (!g1680) & (g1917) & (g1994) & (!g1995)) + ((g132) & (g1592) & (!g1680) & (g1917) & (g1994) & (g1995)) + ((g132) & (g1592) & (g1680) & (g1917) & (g1994) & (!g1995)) + ((g132) & (g1592) & (g1680) & (g1917) & (g1994) & (g1995)));
	assign g1997 = (((!g1548) & (!g1549) & (!g1550) & (g1551) & (g820) & (g773)) + ((!g1548) & (!g1549) & (g1550) & (!g1551) & (!g820) & (g773)) + ((!g1548) & (!g1549) & (g1550) & (g1551) & (!g820) & (g773)) + ((!g1548) & (!g1549) & (g1550) & (g1551) & (g820) & (g773)) + ((!g1548) & (g1549) & (!g1550) & (!g1551) & (g820) & (!g773)) + ((!g1548) & (g1549) & (!g1550) & (g1551) & (g820) & (!g773)) + ((!g1548) & (g1549) & (!g1550) & (g1551) & (g820) & (g773)) + ((!g1548) & (g1549) & (g1550) & (!g1551) & (!g820) & (g773)) + ((!g1548) & (g1549) & (g1550) & (!g1551) & (g820) & (!g773)) + ((!g1548) & (g1549) & (g1550) & (g1551) & (!g820) & (g773)) + ((!g1548) & (g1549) & (g1550) & (g1551) & (g820) & (!g773)) + ((!g1548) & (g1549) & (g1550) & (g1551) & (g820) & (g773)) + ((g1548) & (!g1549) & (!g1550) & (!g1551) & (!g820) & (!g773)) + ((g1548) & (!g1549) & (!g1550) & (g1551) & (!g820) & (!g773)) + ((g1548) & (!g1549) & (!g1550) & (g1551) & (g820) & (g773)) + ((g1548) & (!g1549) & (g1550) & (!g1551) & (!g820) & (!g773)) + ((g1548) & (!g1549) & (g1550) & (!g1551) & (!g820) & (g773)) + ((g1548) & (!g1549) & (g1550) & (g1551) & (!g820) & (!g773)) + ((g1548) & (!g1549) & (g1550) & (g1551) & (!g820) & (g773)) + ((g1548) & (!g1549) & (g1550) & (g1551) & (g820) & (g773)) + ((g1548) & (g1549) & (!g1550) & (!g1551) & (!g820) & (!g773)) + ((g1548) & (g1549) & (!g1550) & (!g1551) & (g820) & (!g773)) + ((g1548) & (g1549) & (!g1550) & (g1551) & (!g820) & (!g773)) + ((g1548) & (g1549) & (!g1550) & (g1551) & (g820) & (!g773)) + ((g1548) & (g1549) & (!g1550) & (g1551) & (g820) & (g773)) + ((g1548) & (g1549) & (g1550) & (!g1551) & (!g820) & (!g773)) + ((g1548) & (g1549) & (g1550) & (!g1551) & (!g820) & (g773)) + ((g1548) & (g1549) & (g1550) & (!g1551) & (g820) & (!g773)) + ((g1548) & (g1549) & (g1550) & (g1551) & (!g820) & (!g773)) + ((g1548) & (g1549) & (g1550) & (g1551) & (!g820) & (g773)) + ((g1548) & (g1549) & (g1550) & (g1551) & (g820) & (!g773)) + ((g1548) & (g1549) & (g1550) & (g1551) & (g820) & (g773)));
	assign g1998 = (((!g1553) & (!g1554) & (!g1555) & (g1556) & (g820) & (g773)) + ((!g1553) & (!g1554) & (g1555) & (!g1556) & (!g820) & (g773)) + ((!g1553) & (!g1554) & (g1555) & (g1556) & (!g820) & (g773)) + ((!g1553) & (!g1554) & (g1555) & (g1556) & (g820) & (g773)) + ((!g1553) & (g1554) & (!g1555) & (!g1556) & (g820) & (!g773)) + ((!g1553) & (g1554) & (!g1555) & (g1556) & (g820) & (!g773)) + ((!g1553) & (g1554) & (!g1555) & (g1556) & (g820) & (g773)) + ((!g1553) & (g1554) & (g1555) & (!g1556) & (!g820) & (g773)) + ((!g1553) & (g1554) & (g1555) & (!g1556) & (g820) & (!g773)) + ((!g1553) & (g1554) & (g1555) & (g1556) & (!g820) & (g773)) + ((!g1553) & (g1554) & (g1555) & (g1556) & (g820) & (!g773)) + ((!g1553) & (g1554) & (g1555) & (g1556) & (g820) & (g773)) + ((g1553) & (!g1554) & (!g1555) & (!g1556) & (!g820) & (!g773)) + ((g1553) & (!g1554) & (!g1555) & (g1556) & (!g820) & (!g773)) + ((g1553) & (!g1554) & (!g1555) & (g1556) & (g820) & (g773)) + ((g1553) & (!g1554) & (g1555) & (!g1556) & (!g820) & (!g773)) + ((g1553) & (!g1554) & (g1555) & (!g1556) & (!g820) & (g773)) + ((g1553) & (!g1554) & (g1555) & (g1556) & (!g820) & (!g773)) + ((g1553) & (!g1554) & (g1555) & (g1556) & (!g820) & (g773)) + ((g1553) & (!g1554) & (g1555) & (g1556) & (g820) & (g773)) + ((g1553) & (g1554) & (!g1555) & (!g1556) & (!g820) & (!g773)) + ((g1553) & (g1554) & (!g1555) & (!g1556) & (g820) & (!g773)) + ((g1553) & (g1554) & (!g1555) & (g1556) & (!g820) & (!g773)) + ((g1553) & (g1554) & (!g1555) & (g1556) & (g820) & (!g773)) + ((g1553) & (g1554) & (!g1555) & (g1556) & (g820) & (g773)) + ((g1553) & (g1554) & (g1555) & (!g1556) & (!g820) & (!g773)) + ((g1553) & (g1554) & (g1555) & (!g1556) & (!g820) & (g773)) + ((g1553) & (g1554) & (g1555) & (!g1556) & (g820) & (!g773)) + ((g1553) & (g1554) & (g1555) & (g1556) & (!g820) & (!g773)) + ((g1553) & (g1554) & (g1555) & (g1556) & (!g820) & (g773)) + ((g1553) & (g1554) & (g1555) & (g1556) & (g820) & (!g773)) + ((g1553) & (g1554) & (g1555) & (g1556) & (g820) & (g773)));
	assign g1999 = (((!g1558) & (!g1559) & (!g1560) & (g1561) & (g820) & (g773)) + ((!g1558) & (!g1559) & (g1560) & (!g1561) & (!g820) & (g773)) + ((!g1558) & (!g1559) & (g1560) & (g1561) & (!g820) & (g773)) + ((!g1558) & (!g1559) & (g1560) & (g1561) & (g820) & (g773)) + ((!g1558) & (g1559) & (!g1560) & (!g1561) & (g820) & (!g773)) + ((!g1558) & (g1559) & (!g1560) & (g1561) & (g820) & (!g773)) + ((!g1558) & (g1559) & (!g1560) & (g1561) & (g820) & (g773)) + ((!g1558) & (g1559) & (g1560) & (!g1561) & (!g820) & (g773)) + ((!g1558) & (g1559) & (g1560) & (!g1561) & (g820) & (!g773)) + ((!g1558) & (g1559) & (g1560) & (g1561) & (!g820) & (g773)) + ((!g1558) & (g1559) & (g1560) & (g1561) & (g820) & (!g773)) + ((!g1558) & (g1559) & (g1560) & (g1561) & (g820) & (g773)) + ((g1558) & (!g1559) & (!g1560) & (!g1561) & (!g820) & (!g773)) + ((g1558) & (!g1559) & (!g1560) & (g1561) & (!g820) & (!g773)) + ((g1558) & (!g1559) & (!g1560) & (g1561) & (g820) & (g773)) + ((g1558) & (!g1559) & (g1560) & (!g1561) & (!g820) & (!g773)) + ((g1558) & (!g1559) & (g1560) & (!g1561) & (!g820) & (g773)) + ((g1558) & (!g1559) & (g1560) & (g1561) & (!g820) & (!g773)) + ((g1558) & (!g1559) & (g1560) & (g1561) & (!g820) & (g773)) + ((g1558) & (!g1559) & (g1560) & (g1561) & (g820) & (g773)) + ((g1558) & (g1559) & (!g1560) & (!g1561) & (!g820) & (!g773)) + ((g1558) & (g1559) & (!g1560) & (!g1561) & (g820) & (!g773)) + ((g1558) & (g1559) & (!g1560) & (g1561) & (!g820) & (!g773)) + ((g1558) & (g1559) & (!g1560) & (g1561) & (g820) & (!g773)) + ((g1558) & (g1559) & (!g1560) & (g1561) & (g820) & (g773)) + ((g1558) & (g1559) & (g1560) & (!g1561) & (!g820) & (!g773)) + ((g1558) & (g1559) & (g1560) & (!g1561) & (!g820) & (g773)) + ((g1558) & (g1559) & (g1560) & (!g1561) & (g820) & (!g773)) + ((g1558) & (g1559) & (g1560) & (g1561) & (!g820) & (!g773)) + ((g1558) & (g1559) & (g1560) & (g1561) & (!g820) & (g773)) + ((g1558) & (g1559) & (g1560) & (g1561) & (g820) & (!g773)) + ((g1558) & (g1559) & (g1560) & (g1561) & (g820) & (g773)));
	assign g2000 = (((!g1563) & (!g1564) & (!g1565) & (g1566) & (g820) & (g773)) + ((!g1563) & (!g1564) & (g1565) & (!g1566) & (!g820) & (g773)) + ((!g1563) & (!g1564) & (g1565) & (g1566) & (!g820) & (g773)) + ((!g1563) & (!g1564) & (g1565) & (g1566) & (g820) & (g773)) + ((!g1563) & (g1564) & (!g1565) & (!g1566) & (g820) & (!g773)) + ((!g1563) & (g1564) & (!g1565) & (g1566) & (g820) & (!g773)) + ((!g1563) & (g1564) & (!g1565) & (g1566) & (g820) & (g773)) + ((!g1563) & (g1564) & (g1565) & (!g1566) & (!g820) & (g773)) + ((!g1563) & (g1564) & (g1565) & (!g1566) & (g820) & (!g773)) + ((!g1563) & (g1564) & (g1565) & (g1566) & (!g820) & (g773)) + ((!g1563) & (g1564) & (g1565) & (g1566) & (g820) & (!g773)) + ((!g1563) & (g1564) & (g1565) & (g1566) & (g820) & (g773)) + ((g1563) & (!g1564) & (!g1565) & (!g1566) & (!g820) & (!g773)) + ((g1563) & (!g1564) & (!g1565) & (g1566) & (!g820) & (!g773)) + ((g1563) & (!g1564) & (!g1565) & (g1566) & (g820) & (g773)) + ((g1563) & (!g1564) & (g1565) & (!g1566) & (!g820) & (!g773)) + ((g1563) & (!g1564) & (g1565) & (!g1566) & (!g820) & (g773)) + ((g1563) & (!g1564) & (g1565) & (g1566) & (!g820) & (!g773)) + ((g1563) & (!g1564) & (g1565) & (g1566) & (!g820) & (g773)) + ((g1563) & (!g1564) & (g1565) & (g1566) & (g820) & (g773)) + ((g1563) & (g1564) & (!g1565) & (!g1566) & (!g820) & (!g773)) + ((g1563) & (g1564) & (!g1565) & (!g1566) & (g820) & (!g773)) + ((g1563) & (g1564) & (!g1565) & (g1566) & (!g820) & (!g773)) + ((g1563) & (g1564) & (!g1565) & (g1566) & (g820) & (!g773)) + ((g1563) & (g1564) & (!g1565) & (g1566) & (g820) & (g773)) + ((g1563) & (g1564) & (g1565) & (!g1566) & (!g820) & (!g773)) + ((g1563) & (g1564) & (g1565) & (!g1566) & (!g820) & (g773)) + ((g1563) & (g1564) & (g1565) & (!g1566) & (g820) & (!g773)) + ((g1563) & (g1564) & (g1565) & (g1566) & (!g820) & (!g773)) + ((g1563) & (g1564) & (g1565) & (g1566) & (!g820) & (g773)) + ((g1563) & (g1564) & (g1565) & (g1566) & (g820) & (!g773)) + ((g1563) & (g1564) & (g1565) & (g1566) & (g820) & (g773)));
	assign g2001 = (((!g1997) & (!g1998) & (!g1999) & (g2000) & (g677) & (g726)) + ((!g1997) & (!g1998) & (g1999) & (!g2000) & (!g677) & (g726)) + ((!g1997) & (!g1998) & (g1999) & (g2000) & (!g677) & (g726)) + ((!g1997) & (!g1998) & (g1999) & (g2000) & (g677) & (g726)) + ((!g1997) & (g1998) & (!g1999) & (!g2000) & (g677) & (!g726)) + ((!g1997) & (g1998) & (!g1999) & (g2000) & (g677) & (!g726)) + ((!g1997) & (g1998) & (!g1999) & (g2000) & (g677) & (g726)) + ((!g1997) & (g1998) & (g1999) & (!g2000) & (!g677) & (g726)) + ((!g1997) & (g1998) & (g1999) & (!g2000) & (g677) & (!g726)) + ((!g1997) & (g1998) & (g1999) & (g2000) & (!g677) & (g726)) + ((!g1997) & (g1998) & (g1999) & (g2000) & (g677) & (!g726)) + ((!g1997) & (g1998) & (g1999) & (g2000) & (g677) & (g726)) + ((g1997) & (!g1998) & (!g1999) & (!g2000) & (!g677) & (!g726)) + ((g1997) & (!g1998) & (!g1999) & (g2000) & (!g677) & (!g726)) + ((g1997) & (!g1998) & (!g1999) & (g2000) & (g677) & (g726)) + ((g1997) & (!g1998) & (g1999) & (!g2000) & (!g677) & (!g726)) + ((g1997) & (!g1998) & (g1999) & (!g2000) & (!g677) & (g726)) + ((g1997) & (!g1998) & (g1999) & (g2000) & (!g677) & (!g726)) + ((g1997) & (!g1998) & (g1999) & (g2000) & (!g677) & (g726)) + ((g1997) & (!g1998) & (g1999) & (g2000) & (g677) & (g726)) + ((g1997) & (g1998) & (!g1999) & (!g2000) & (!g677) & (!g726)) + ((g1997) & (g1998) & (!g1999) & (!g2000) & (g677) & (!g726)) + ((g1997) & (g1998) & (!g1999) & (g2000) & (!g677) & (!g726)) + ((g1997) & (g1998) & (!g1999) & (g2000) & (g677) & (!g726)) + ((g1997) & (g1998) & (!g1999) & (g2000) & (g677) & (g726)) + ((g1997) & (g1998) & (g1999) & (!g2000) & (!g677) & (!g726)) + ((g1997) & (g1998) & (g1999) & (!g2000) & (!g677) & (g726)) + ((g1997) & (g1998) & (g1999) & (!g2000) & (g677) & (!g726)) + ((g1997) & (g1998) & (g1999) & (g2000) & (!g677) & (!g726)) + ((g1997) & (g1998) & (g1999) & (g2000) & (!g677) & (g726)) + ((g1997) & (g1998) & (g1999) & (g2000) & (g677) & (!g726)) + ((g1997) & (g1998) & (g1999) & (g2000) & (g677) & (g726)));
	assign g2002 = (((!g1569) & (!g1570) & (!g1571) & (g1572) & (g677) & (g726)) + ((!g1569) & (!g1570) & (g1571) & (!g1572) & (!g677) & (g726)) + ((!g1569) & (!g1570) & (g1571) & (g1572) & (!g677) & (g726)) + ((!g1569) & (!g1570) & (g1571) & (g1572) & (g677) & (g726)) + ((!g1569) & (g1570) & (!g1571) & (!g1572) & (g677) & (!g726)) + ((!g1569) & (g1570) & (!g1571) & (g1572) & (g677) & (!g726)) + ((!g1569) & (g1570) & (!g1571) & (g1572) & (g677) & (g726)) + ((!g1569) & (g1570) & (g1571) & (!g1572) & (!g677) & (g726)) + ((!g1569) & (g1570) & (g1571) & (!g1572) & (g677) & (!g726)) + ((!g1569) & (g1570) & (g1571) & (g1572) & (!g677) & (g726)) + ((!g1569) & (g1570) & (g1571) & (g1572) & (g677) & (!g726)) + ((!g1569) & (g1570) & (g1571) & (g1572) & (g677) & (g726)) + ((g1569) & (!g1570) & (!g1571) & (!g1572) & (!g677) & (!g726)) + ((g1569) & (!g1570) & (!g1571) & (g1572) & (!g677) & (!g726)) + ((g1569) & (!g1570) & (!g1571) & (g1572) & (g677) & (g726)) + ((g1569) & (!g1570) & (g1571) & (!g1572) & (!g677) & (!g726)) + ((g1569) & (!g1570) & (g1571) & (!g1572) & (!g677) & (g726)) + ((g1569) & (!g1570) & (g1571) & (g1572) & (!g677) & (!g726)) + ((g1569) & (!g1570) & (g1571) & (g1572) & (!g677) & (g726)) + ((g1569) & (!g1570) & (g1571) & (g1572) & (g677) & (g726)) + ((g1569) & (g1570) & (!g1571) & (!g1572) & (!g677) & (!g726)) + ((g1569) & (g1570) & (!g1571) & (!g1572) & (g677) & (!g726)) + ((g1569) & (g1570) & (!g1571) & (g1572) & (!g677) & (!g726)) + ((g1569) & (g1570) & (!g1571) & (g1572) & (g677) & (!g726)) + ((g1569) & (g1570) & (!g1571) & (g1572) & (g677) & (g726)) + ((g1569) & (g1570) & (g1571) & (!g1572) & (!g677) & (!g726)) + ((g1569) & (g1570) & (g1571) & (!g1572) & (!g677) & (g726)) + ((g1569) & (g1570) & (g1571) & (!g1572) & (g677) & (!g726)) + ((g1569) & (g1570) & (g1571) & (g1572) & (!g677) & (!g726)) + ((g1569) & (g1570) & (g1571) & (g1572) & (!g677) & (g726)) + ((g1569) & (g1570) & (g1571) & (g1572) & (g677) & (!g726)) + ((g1569) & (g1570) & (g1571) & (g1572) & (g677) & (g726)));
	assign g2003 = (((!g677) & (!g726) & (!sk[21]) & (!g1574) & (g1575) & (!g1576)) + ((!g677) & (!g726) & (!sk[21]) & (!g1574) & (g1575) & (g1576)) + ((!g677) & (!g726) & (!sk[21]) & (g1574) & (!g1575) & (!g1576)) + ((!g677) & (!g726) & (!sk[21]) & (g1574) & (!g1575) & (g1576)) + ((!g677) & (!g726) & (!sk[21]) & (g1574) & (g1575) & (!g1576)) + ((!g677) & (!g726) & (!sk[21]) & (g1574) & (g1575) & (g1576)) + ((!g677) & (g726) & (!sk[21]) & (!g1574) & (!g1575) & (!g1576)) + ((!g677) & (g726) & (!sk[21]) & (!g1574) & (!g1575) & (g1576)) + ((!g677) & (g726) & (!sk[21]) & (!g1574) & (g1575) & (!g1576)) + ((!g677) & (g726) & (!sk[21]) & (!g1574) & (g1575) & (g1576)) + ((!g677) & (g726) & (!sk[21]) & (g1574) & (!g1575) & (!g1576)) + ((!g677) & (g726) & (!sk[21]) & (g1574) & (!g1575) & (g1576)) + ((!g677) & (g726) & (!sk[21]) & (g1574) & (g1575) & (!g1576)) + ((!g677) & (g726) & (!sk[21]) & (g1574) & (g1575) & (g1576)) + ((!g677) & (g726) & (sk[21]) & (!g1574) & (!g1575) & (g1576)) + ((!g677) & (g726) & (sk[21]) & (!g1574) & (g1575) & (g1576)) + ((!g677) & (g726) & (sk[21]) & (g1574) & (!g1575) & (g1576)) + ((!g677) & (g726) & (sk[21]) & (g1574) & (g1575) & (g1576)) + ((g677) & (!g726) & (!sk[21]) & (!g1574) & (g1575) & (!g1576)) + ((g677) & (!g726) & (!sk[21]) & (!g1574) & (g1575) & (g1576)) + ((g677) & (!g726) & (!sk[21]) & (g1574) & (!g1575) & (!g1576)) + ((g677) & (!g726) & (!sk[21]) & (g1574) & (!g1575) & (g1576)) + ((g677) & (!g726) & (!sk[21]) & (g1574) & (g1575) & (!g1576)) + ((g677) & (!g726) & (!sk[21]) & (g1574) & (g1575) & (g1576)) + ((g677) & (!g726) & (sk[21]) & (g1574) & (!g1575) & (!g1576)) + ((g677) & (!g726) & (sk[21]) & (g1574) & (!g1575) & (g1576)) + ((g677) & (!g726) & (sk[21]) & (g1574) & (g1575) & (!g1576)) + ((g677) & (!g726) & (sk[21]) & (g1574) & (g1575) & (g1576)) + ((g677) & (g726) & (!sk[21]) & (!g1574) & (!g1575) & (!g1576)) + ((g677) & (g726) & (!sk[21]) & (!g1574) & (!g1575) & (g1576)) + ((g677) & (g726) & (!sk[21]) & (!g1574) & (g1575) & (!g1576)) + ((g677) & (g726) & (!sk[21]) & (!g1574) & (g1575) & (g1576)) + ((g677) & (g726) & (!sk[21]) & (g1574) & (!g1575) & (!g1576)) + ((g677) & (g726) & (!sk[21]) & (g1574) & (!g1575) & (g1576)) + ((g677) & (g726) & (!sk[21]) & (g1574) & (g1575) & (!g1576)) + ((g677) & (g726) & (!sk[21]) & (g1574) & (g1575) & (g1576)) + ((g677) & (g726) & (sk[21]) & (!g1574) & (g1575) & (!g1576)) + ((g677) & (g726) & (sk[21]) & (!g1574) & (g1575) & (g1576)) + ((g677) & (g726) & (sk[21]) & (g1574) & (g1575) & (!g1576)) + ((g677) & (g726) & (sk[21]) & (g1574) & (g1575) & (g1576)));
	assign g2004 = (((!g1578) & (!g1579) & (!g1580) & (g1581) & (g677) & (g726)) + ((!g1578) & (!g1579) & (g1580) & (!g1581) & (!g677) & (g726)) + ((!g1578) & (!g1579) & (g1580) & (g1581) & (!g677) & (g726)) + ((!g1578) & (!g1579) & (g1580) & (g1581) & (g677) & (g726)) + ((!g1578) & (g1579) & (!g1580) & (!g1581) & (g677) & (!g726)) + ((!g1578) & (g1579) & (!g1580) & (g1581) & (g677) & (!g726)) + ((!g1578) & (g1579) & (!g1580) & (g1581) & (g677) & (g726)) + ((!g1578) & (g1579) & (g1580) & (!g1581) & (!g677) & (g726)) + ((!g1578) & (g1579) & (g1580) & (!g1581) & (g677) & (!g726)) + ((!g1578) & (g1579) & (g1580) & (g1581) & (!g677) & (g726)) + ((!g1578) & (g1579) & (g1580) & (g1581) & (g677) & (!g726)) + ((!g1578) & (g1579) & (g1580) & (g1581) & (g677) & (g726)) + ((g1578) & (!g1579) & (!g1580) & (!g1581) & (!g677) & (!g726)) + ((g1578) & (!g1579) & (!g1580) & (g1581) & (!g677) & (!g726)) + ((g1578) & (!g1579) & (!g1580) & (g1581) & (g677) & (g726)) + ((g1578) & (!g1579) & (g1580) & (!g1581) & (!g677) & (!g726)) + ((g1578) & (!g1579) & (g1580) & (!g1581) & (!g677) & (g726)) + ((g1578) & (!g1579) & (g1580) & (g1581) & (!g677) & (!g726)) + ((g1578) & (!g1579) & (g1580) & (g1581) & (!g677) & (g726)) + ((g1578) & (!g1579) & (g1580) & (g1581) & (g677) & (g726)) + ((g1578) & (g1579) & (!g1580) & (!g1581) & (!g677) & (!g726)) + ((g1578) & (g1579) & (!g1580) & (!g1581) & (g677) & (!g726)) + ((g1578) & (g1579) & (!g1580) & (g1581) & (!g677) & (!g726)) + ((g1578) & (g1579) & (!g1580) & (g1581) & (g677) & (!g726)) + ((g1578) & (g1579) & (!g1580) & (g1581) & (g677) & (g726)) + ((g1578) & (g1579) & (g1580) & (!g1581) & (!g677) & (!g726)) + ((g1578) & (g1579) & (g1580) & (!g1581) & (!g677) & (g726)) + ((g1578) & (g1579) & (g1580) & (!g1581) & (g677) & (!g726)) + ((g1578) & (g1579) & (g1580) & (g1581) & (!g677) & (!g726)) + ((g1578) & (g1579) & (g1580) & (g1581) & (!g677) & (g726)) + ((g1578) & (g1579) & (g1580) & (g1581) & (g677) & (!g726)) + ((g1578) & (g1579) & (g1580) & (g1581) & (g677) & (g726)));
	assign g2005 = (((!g1583) & (!g1584) & (!g1585) & (g1586) & (g677) & (g726)) + ((!g1583) & (!g1584) & (g1585) & (!g1586) & (!g677) & (g726)) + ((!g1583) & (!g1584) & (g1585) & (g1586) & (!g677) & (g726)) + ((!g1583) & (!g1584) & (g1585) & (g1586) & (g677) & (g726)) + ((!g1583) & (g1584) & (!g1585) & (!g1586) & (g677) & (!g726)) + ((!g1583) & (g1584) & (!g1585) & (g1586) & (g677) & (!g726)) + ((!g1583) & (g1584) & (!g1585) & (g1586) & (g677) & (g726)) + ((!g1583) & (g1584) & (g1585) & (!g1586) & (!g677) & (g726)) + ((!g1583) & (g1584) & (g1585) & (!g1586) & (g677) & (!g726)) + ((!g1583) & (g1584) & (g1585) & (g1586) & (!g677) & (g726)) + ((!g1583) & (g1584) & (g1585) & (g1586) & (g677) & (!g726)) + ((!g1583) & (g1584) & (g1585) & (g1586) & (g677) & (g726)) + ((g1583) & (!g1584) & (!g1585) & (!g1586) & (!g677) & (!g726)) + ((g1583) & (!g1584) & (!g1585) & (g1586) & (!g677) & (!g726)) + ((g1583) & (!g1584) & (!g1585) & (g1586) & (g677) & (g726)) + ((g1583) & (!g1584) & (g1585) & (!g1586) & (!g677) & (!g726)) + ((g1583) & (!g1584) & (g1585) & (!g1586) & (!g677) & (g726)) + ((g1583) & (!g1584) & (g1585) & (g1586) & (!g677) & (!g726)) + ((g1583) & (!g1584) & (g1585) & (g1586) & (!g677) & (g726)) + ((g1583) & (!g1584) & (g1585) & (g1586) & (g677) & (g726)) + ((g1583) & (g1584) & (!g1585) & (!g1586) & (!g677) & (!g726)) + ((g1583) & (g1584) & (!g1585) & (!g1586) & (g677) & (!g726)) + ((g1583) & (g1584) & (!g1585) & (g1586) & (!g677) & (!g726)) + ((g1583) & (g1584) & (!g1585) & (g1586) & (g677) & (!g726)) + ((g1583) & (g1584) & (!g1585) & (g1586) & (g677) & (g726)) + ((g1583) & (g1584) & (g1585) & (!g1586) & (!g677) & (!g726)) + ((g1583) & (g1584) & (g1585) & (!g1586) & (!g677) & (g726)) + ((g1583) & (g1584) & (g1585) & (!g1586) & (g677) & (!g726)) + ((g1583) & (g1584) & (g1585) & (g1586) & (!g677) & (!g726)) + ((g1583) & (g1584) & (g1585) & (g1586) & (!g677) & (g726)) + ((g1583) & (g1584) & (g1585) & (g1586) & (g677) & (!g726)) + ((g1583) & (g1584) & (g1585) & (g1586) & (g677) & (g726)));
	assign g2006 = (((!g820) & (!g773) & (!g2002) & (g2003) & (!g2004) & (!g2005)) + ((!g820) & (!g773) & (!g2002) & (g2003) & (!g2004) & (g2005)) + ((!g820) & (!g773) & (!g2002) & (g2003) & (g2004) & (!g2005)) + ((!g820) & (!g773) & (!g2002) & (g2003) & (g2004) & (g2005)) + ((!g820) & (!g773) & (g2002) & (g2003) & (!g2004) & (!g2005)) + ((!g820) & (!g773) & (g2002) & (g2003) & (!g2004) & (g2005)) + ((!g820) & (!g773) & (g2002) & (g2003) & (g2004) & (!g2005)) + ((!g820) & (!g773) & (g2002) & (g2003) & (g2004) & (g2005)) + ((!g820) & (g773) & (!g2002) & (!g2003) & (!g2004) & (g2005)) + ((!g820) & (g773) & (!g2002) & (!g2003) & (g2004) & (g2005)) + ((!g820) & (g773) & (!g2002) & (g2003) & (!g2004) & (g2005)) + ((!g820) & (g773) & (!g2002) & (g2003) & (g2004) & (g2005)) + ((!g820) & (g773) & (g2002) & (!g2003) & (!g2004) & (g2005)) + ((!g820) & (g773) & (g2002) & (!g2003) & (g2004) & (g2005)) + ((!g820) & (g773) & (g2002) & (g2003) & (!g2004) & (g2005)) + ((!g820) & (g773) & (g2002) & (g2003) & (g2004) & (g2005)) + ((g820) & (!g773) & (g2002) & (!g2003) & (!g2004) & (!g2005)) + ((g820) & (!g773) & (g2002) & (!g2003) & (!g2004) & (g2005)) + ((g820) & (!g773) & (g2002) & (!g2003) & (g2004) & (!g2005)) + ((g820) & (!g773) & (g2002) & (!g2003) & (g2004) & (g2005)) + ((g820) & (!g773) & (g2002) & (g2003) & (!g2004) & (!g2005)) + ((g820) & (!g773) & (g2002) & (g2003) & (!g2004) & (g2005)) + ((g820) & (!g773) & (g2002) & (g2003) & (g2004) & (!g2005)) + ((g820) & (!g773) & (g2002) & (g2003) & (g2004) & (g2005)) + ((g820) & (g773) & (!g2002) & (!g2003) & (g2004) & (!g2005)) + ((g820) & (g773) & (!g2002) & (!g2003) & (g2004) & (g2005)) + ((g820) & (g773) & (!g2002) & (g2003) & (g2004) & (!g2005)) + ((g820) & (g773) & (!g2002) & (g2003) & (g2004) & (g2005)) + ((g820) & (g773) & (g2002) & (!g2003) & (g2004) & (!g2005)) + ((g820) & (g773) & (g2002) & (!g2003) & (g2004) & (g2005)) + ((g820) & (g773) & (g2002) & (g2003) & (g2004) & (!g2005)) + ((g820) & (g773) & (g2002) & (g2003) & (g2004) & (g2005)));
	assign g2007 = (((!sk[25]) & (!g867) & (!g2001) & (g2006)) + ((!sk[25]) & (!g867) & (g2001) & (!g2006)) + ((!sk[25]) & (!g867) & (g2001) & (g2006)) + ((!sk[25]) & (g867) & (!g2001) & (g2006)) + ((!sk[25]) & (g867) & (g2001) & (!g2006)) + ((!sk[25]) & (g867) & (g2001) & (g2006)) + ((sk[25]) & (!g867) & (!g2001) & (g2006)) + ((sk[25]) & (!g867) & (g2001) & (g2006)) + ((sk[25]) & (g867) & (g2001) & (!g2006)) + ((sk[25]) & (g867) & (g2001) & (g2006)));
	assign g2008 = (((!g1593) & (!g1605) & (!g1798) & (!sk[26]) & (g66)) + ((!g1593) & (!g1605) & (g1798) & (!sk[26]) & (!g66)) + ((!g1593) & (!g1605) & (g1798) & (!sk[26]) & (g66)) + ((!g1593) & (!g1605) & (g1798) & (sk[26]) & (!g66)) + ((!g1593) & (!g1605) & (g1798) & (sk[26]) & (g66)) + ((!g1593) & (g1605) & (!g1798) & (!sk[26]) & (!g66)) + ((!g1593) & (g1605) & (!g1798) & (!sk[26]) & (g66)) + ((!g1593) & (g1605) & (g1798) & (!sk[26]) & (!g66)) + ((!g1593) & (g1605) & (g1798) & (!sk[26]) & (g66)) + ((g1593) & (!g1605) & (!g1798) & (!sk[26]) & (g66)) + ((g1593) & (!g1605) & (!g1798) & (sk[26]) & (g66)) + ((g1593) & (!g1605) & (g1798) & (!sk[26]) & (!g66)) + ((g1593) & (!g1605) & (g1798) & (!sk[26]) & (g66)) + ((g1593) & (!g1605) & (g1798) & (sk[26]) & (g66)) + ((g1593) & (g1605) & (!g1798) & (!sk[26]) & (!g66)) + ((g1593) & (g1605) & (!g1798) & (!sk[26]) & (g66)) + ((g1593) & (g1605) & (!g1798) & (sk[26]) & (g66)) + ((g1593) & (g1605) & (g1798) & (!sk[26]) & (!g66)) + ((g1593) & (g1605) & (g1798) & (!sk[26]) & (g66)) + ((g1593) & (g1605) & (g1798) & (sk[26]) & (g66)));
	assign g2009 = (((!g132) & (!g1592) & (g1692) & (g1917) & (!g2007) & (!g2008)) + ((!g132) & (!g1592) & (g1692) & (g1917) & (!g2007) & (g2008)) + ((!g132) & (!g1592) & (g1692) & (g1917) & (g2007) & (!g2008)) + ((!g132) & (!g1592) & (g1692) & (g1917) & (g2007) & (g2008)) + ((!g132) & (g1592) & (!g1692) & (g1917) & (!g2007) & (g2008)) + ((!g132) & (g1592) & (!g1692) & (g1917) & (g2007) & (g2008)) + ((!g132) & (g1592) & (g1692) & (g1917) & (!g2007) & (g2008)) + ((!g132) & (g1592) & (g1692) & (g1917) & (g2007) & (g2008)) + ((g132) & (!g1592) & (!g1692) & (g1917) & (g2007) & (!g2008)) + ((g132) & (!g1592) & (!g1692) & (g1917) & (g2007) & (g2008)) + ((g132) & (!g1592) & (g1692) & (g1917) & (g2007) & (!g2008)) + ((g132) & (!g1592) & (g1692) & (g1917) & (g2007) & (g2008)) + ((g132) & (g1592) & (!g1692) & (g1917) & (g2007) & (!g2008)) + ((g132) & (g1592) & (!g1692) & (g1917) & (g2007) & (g2008)) + ((g132) & (g1592) & (g1692) & (g1917) & (g2007) & (!g2008)) + ((g132) & (g1592) & (g1692) & (g1917) & (g2007) & (g2008)));
	assign g2010 = (((!g1592) & (!g137) & (!sk[28]) & (!g126) & (g1593)) + ((!g1592) & (!g137) & (!sk[28]) & (g126) & (!g1593)) + ((!g1592) & (!g137) & (!sk[28]) & (g126) & (g1593)) + ((!g1592) & (!g137) & (sk[28]) & (!g126) & (!g1593)) + ((!g1592) & (!g137) & (sk[28]) & (!g126) & (g1593)) + ((!g1592) & (!g137) & (sk[28]) & (g126) & (!g1593)) + ((!g1592) & (!g137) & (sk[28]) & (g126) & (g1593)) + ((!g1592) & (g137) & (!sk[28]) & (!g126) & (!g1593)) + ((!g1592) & (g137) & (!sk[28]) & (!g126) & (g1593)) + ((!g1592) & (g137) & (!sk[28]) & (g126) & (!g1593)) + ((!g1592) & (g137) & (!sk[28]) & (g126) & (g1593)) + ((!g1592) & (g137) & (sk[28]) & (!g126) & (!g1593)) + ((!g1592) & (g137) & (sk[28]) & (!g126) & (g1593)) + ((g1592) & (!g137) & (!sk[28]) & (!g126) & (g1593)) + ((g1592) & (!g137) & (!sk[28]) & (g126) & (!g1593)) + ((g1592) & (!g137) & (!sk[28]) & (g126) & (g1593)) + ((g1592) & (!g137) & (sk[28]) & (!g126) & (!g1593)) + ((g1592) & (!g137) & (sk[28]) & (!g126) & (g1593)) + ((g1592) & (!g137) & (sk[28]) & (g126) & (!g1593)) + ((g1592) & (g137) & (!sk[28]) & (!g126) & (!g1593)) + ((g1592) & (g137) & (!sk[28]) & (!g126) & (g1593)) + ((g1592) & (g137) & (!sk[28]) & (g126) & (!g1593)) + ((g1592) & (g137) & (!sk[28]) & (g126) & (g1593)) + ((g1592) & (g137) & (sk[28]) & (!g126) & (!g1593)) + ((g1592) & (g137) & (sk[28]) & (!g126) & (g1593)));
	assign g2011 = (((!g68) & (!g130) & (!sk[29]) & (!g2010) & (dmem_stall_i)) + ((!g68) & (!g130) & (!sk[29]) & (g2010) & (!dmem_stall_i)) + ((!g68) & (!g130) & (!sk[29]) & (g2010) & (dmem_stall_i)) + ((!g68) & (g130) & (!sk[29]) & (!g2010) & (!dmem_stall_i)) + ((!g68) & (g130) & (!sk[29]) & (!g2010) & (dmem_stall_i)) + ((!g68) & (g130) & (!sk[29]) & (g2010) & (!dmem_stall_i)) + ((!g68) & (g130) & (!sk[29]) & (g2010) & (dmem_stall_i)) + ((!g68) & (g130) & (sk[29]) & (g2010) & (!dmem_stall_i)) + ((!g68) & (g130) & (sk[29]) & (g2010) & (dmem_stall_i)) + ((g68) & (!g130) & (!sk[29]) & (!g2010) & (dmem_stall_i)) + ((g68) & (!g130) & (!sk[29]) & (g2010) & (!dmem_stall_i)) + ((g68) & (!g130) & (!sk[29]) & (g2010) & (dmem_stall_i)) + ((g68) & (!g130) & (sk[29]) & (!g2010) & (dmem_stall_i)) + ((g68) & (!g130) & (sk[29]) & (g2010) & (dmem_stall_i)) + ((g68) & (g130) & (!sk[29]) & (!g2010) & (!dmem_stall_i)) + ((g68) & (g130) & (!sk[29]) & (!g2010) & (dmem_stall_i)) + ((g68) & (g130) & (!sk[29]) & (g2010) & (!dmem_stall_i)) + ((g68) & (g130) & (!sk[29]) & (g2010) & (dmem_stall_i)) + ((g68) & (g130) & (sk[29]) & (!g2010) & (dmem_stall_i)) + ((g68) & (g130) & (sk[29]) & (g2010) & (!dmem_stall_i)) + ((g68) & (g130) & (sk[29]) & (g2010) & (dmem_stall_i)));
	assign g2012 = (((!g69) & (!g132) & (!g1592) & (!g1606) & (!g136) & (!g1593)) + ((!g69) & (!g132) & (!g1592) & (!g1606) & (!g136) & (g1593)) + ((!g69) & (!g132) & (!g1592) & (!g1606) & (g136) & (!g1593)) + ((!g69) & (!g132) & (!g1592) & (!g1606) & (g136) & (g1593)) + ((!g69) & (!g132) & (g1592) & (!g1606) & (!g136) & (g1593)) + ((!g69) & (!g132) & (g1592) & (!g1606) & (g136) & (g1593)) + ((g69) & (!g132) & (!g1592) & (!g1606) & (g136) & (!g1593)) + ((g69) & (!g132) & (!g1592) & (!g1606) & (g136) & (g1593)));
	assign g2013 = (((!g69) & (!sk[31]) & (!g126) & (!g130) & (g2012)) + ((!g69) & (!sk[31]) & (!g126) & (g130) & (!g2012)) + ((!g69) & (!sk[31]) & (!g126) & (g130) & (g2012)) + ((!g69) & (!sk[31]) & (g126) & (!g130) & (!g2012)) + ((!g69) & (!sk[31]) & (g126) & (!g130) & (g2012)) + ((!g69) & (!sk[31]) & (g126) & (g130) & (!g2012)) + ((!g69) & (!sk[31]) & (g126) & (g130) & (g2012)) + ((!g69) & (sk[31]) & (g126) & (!g130) & (!g2012)) + ((!g69) & (sk[31]) & (g126) & (g130) & (!g2012)) + ((g69) & (!sk[31]) & (!g126) & (!g130) & (g2012)) + ((g69) & (!sk[31]) & (!g126) & (g130) & (!g2012)) + ((g69) & (!sk[31]) & (!g126) & (g130) & (g2012)) + ((g69) & (!sk[31]) & (g126) & (!g130) & (!g2012)) + ((g69) & (!sk[31]) & (g126) & (!g130) & (g2012)) + ((g69) & (!sk[31]) & (g126) & (g130) & (!g2012)) + ((g69) & (!sk[31]) & (g126) & (g130) & (g2012)) + ((g69) & (sk[31]) & (!g126) & (!g130) & (!g2012)) + ((g69) & (sk[31]) & (!g126) & (!g130) & (g2012)) + ((g69) & (sk[31]) & (g126) & (!g130) & (!g2012)) + ((g69) & (sk[31]) & (g126) & (!g130) & (g2012)) + ((g69) & (sk[31]) & (g126) & (g130) & (!g2012)));
	assign g2014 = (((!g1592) & (!g1606) & (!sk[32]) & (!g1593) & (g1605)) + ((!g1592) & (!g1606) & (!sk[32]) & (g1593) & (!g1605)) + ((!g1592) & (!g1606) & (!sk[32]) & (g1593) & (g1605)) + ((!g1592) & (!g1606) & (sk[32]) & (!g1593) & (!g1605)) + ((!g1592) & (!g1606) & (sk[32]) & (!g1593) & (g1605)) + ((!g1592) & (!g1606) & (sk[32]) & (g1593) & (!g1605)) + ((!g1592) & (!g1606) & (sk[32]) & (g1593) & (g1605)) + ((!g1592) & (g1606) & (!sk[32]) & (!g1593) & (!g1605)) + ((!g1592) & (g1606) & (!sk[32]) & (!g1593) & (g1605)) + ((!g1592) & (g1606) & (!sk[32]) & (g1593) & (!g1605)) + ((!g1592) & (g1606) & (!sk[32]) & (g1593) & (g1605)) + ((!g1592) & (g1606) & (sk[32]) & (g1593) & (g1605)) + ((g1592) & (!g1606) & (!sk[32]) & (!g1593) & (g1605)) + ((g1592) & (!g1606) & (!sk[32]) & (g1593) & (!g1605)) + ((g1592) & (!g1606) & (!sk[32]) & (g1593) & (g1605)) + ((g1592) & (!g1606) & (sk[32]) & (!g1593) & (g1605)) + ((g1592) & (!g1606) & (sk[32]) & (g1593) & (g1605)) + ((g1592) & (g1606) & (!sk[32]) & (!g1593) & (!g1605)) + ((g1592) & (g1606) & (!sk[32]) & (!g1593) & (g1605)) + ((g1592) & (g1606) & (!sk[32]) & (g1593) & (!g1605)) + ((g1592) & (g1606) & (!sk[32]) & (g1593) & (g1605)) + ((g1592) & (g1606) & (sk[32]) & (!g1593) & (g1605)) + ((g1592) & (g1606) & (sk[32]) & (g1593) & (g1605)));
	assign g2015 = (((!g1592) & (!g1593) & (!sk[33]) & (g1609)) + ((!g1592) & (!g1593) & (sk[33]) & (g1609)) + ((!g1592) & (g1593) & (!sk[33]) & (!g1609)) + ((!g1592) & (g1593) & (!sk[33]) & (g1609)) + ((!g1592) & (g1593) & (sk[33]) & (g1609)) + ((g1592) & (!g1593) & (!sk[33]) & (g1609)) + ((g1592) & (!g1593) & (sk[33]) & (g1609)) + ((g1592) & (g1593) & (!sk[33]) & (!g1609)) + ((g1592) & (g1593) & (!sk[33]) & (g1609)));
	assign g2016 = (((!g1592) & (!sk[34]) & (!g1606) & (!g1593) & (g1605)) + ((!g1592) & (!sk[34]) & (!g1606) & (g1593) & (!g1605)) + ((!g1592) & (!sk[34]) & (!g1606) & (g1593) & (g1605)) + ((!g1592) & (!sk[34]) & (g1606) & (!g1593) & (!g1605)) + ((!g1592) & (!sk[34]) & (g1606) & (!g1593) & (g1605)) + ((!g1592) & (!sk[34]) & (g1606) & (g1593) & (!g1605)) + ((!g1592) & (!sk[34]) & (g1606) & (g1593) & (g1605)) + ((!g1592) & (sk[34]) & (!g1606) & (!g1593) & (!g1605)) + ((!g1592) & (sk[34]) & (!g1606) & (!g1593) & (g1605)) + ((!g1592) & (sk[34]) & (!g1606) & (g1593) & (!g1605)) + ((!g1592) & (sk[34]) & (!g1606) & (g1593) & (g1605)) + ((!g1592) & (sk[34]) & (g1606) & (!g1593) & (g1605)) + ((g1592) & (!sk[34]) & (!g1606) & (!g1593) & (g1605)) + ((g1592) & (!sk[34]) & (!g1606) & (g1593) & (!g1605)) + ((g1592) & (!sk[34]) & (!g1606) & (g1593) & (g1605)) + ((g1592) & (!sk[34]) & (g1606) & (!g1593) & (!g1605)) + ((g1592) & (!sk[34]) & (g1606) & (!g1593) & (g1605)) + ((g1592) & (!sk[34]) & (g1606) & (g1593) & (!g1605)) + ((g1592) & (!sk[34]) & (g1606) & (g1593) & (g1605)) + ((g1592) & (sk[34]) & (!g1606) & (!g1593) & (g1605)) + ((g1592) & (sk[34]) & (!g1606) & (g1593) & (g1605)) + ((g1592) & (sk[34]) & (g1606) & (!g1593) & (g1605)) + ((g1592) & (sk[34]) & (g1606) & (g1593) & (g1605)));
	assign g2017 = (((!g1592) & (!g1606) & (!g1593) & (!sk[35]) & (g1605)) + ((!g1592) & (!g1606) & (!g1593) & (sk[35]) & (!g1605)) + ((!g1592) & (!g1606) & (!g1593) & (sk[35]) & (g1605)) + ((!g1592) & (!g1606) & (g1593) & (!sk[35]) & (!g1605)) + ((!g1592) & (!g1606) & (g1593) & (!sk[35]) & (g1605)) + ((!g1592) & (!g1606) & (g1593) & (sk[35]) & (!g1605)) + ((!g1592) & (!g1606) & (g1593) & (sk[35]) & (g1605)) + ((!g1592) & (g1606) & (!g1593) & (!sk[35]) & (!g1605)) + ((!g1592) & (g1606) & (!g1593) & (!sk[35]) & (g1605)) + ((!g1592) & (g1606) & (g1593) & (!sk[35]) & (!g1605)) + ((!g1592) & (g1606) & (g1593) & (!sk[35]) & (g1605)) + ((!g1592) & (g1606) & (g1593) & (sk[35]) & (!g1605)) + ((g1592) & (!g1606) & (!g1593) & (!sk[35]) & (g1605)) + ((g1592) & (!g1606) & (!g1593) & (sk[35]) & (!g1605)) + ((g1592) & (!g1606) & (g1593) & (!sk[35]) & (!g1605)) + ((g1592) & (!g1606) & (g1593) & (!sk[35]) & (g1605)) + ((g1592) & (!g1606) & (g1593) & (sk[35]) & (!g1605)) + ((g1592) & (g1606) & (!g1593) & (!sk[35]) & (!g1605)) + ((g1592) & (g1606) & (!g1593) & (!sk[35]) & (g1605)) + ((g1592) & (g1606) & (!g1593) & (sk[35]) & (!g1605)) + ((g1592) & (g1606) & (g1593) & (!sk[35]) & (!g1605)) + ((g1592) & (g1606) & (g1593) & (!sk[35]) & (g1605)) + ((g1592) & (g1606) & (g1593) & (sk[35]) & (!g1605)));
	assign g2018 = (((!g1592) & (!g1606) & (!sk[36]) & (!g1593) & (g1605)) + ((!g1592) & (!g1606) & (!sk[36]) & (g1593) & (!g1605)) + ((!g1592) & (!g1606) & (!sk[36]) & (g1593) & (g1605)) + ((!g1592) & (!g1606) & (sk[36]) & (!g1593) & (!g1605)) + ((!g1592) & (!g1606) & (sk[36]) & (!g1593) & (g1605)) + ((!g1592) & (!g1606) & (sk[36]) & (g1593) & (!g1605)) + ((!g1592) & (!g1606) & (sk[36]) & (g1593) & (g1605)) + ((!g1592) & (g1606) & (!sk[36]) & (!g1593) & (!g1605)) + ((!g1592) & (g1606) & (!sk[36]) & (!g1593) & (g1605)) + ((!g1592) & (g1606) & (!sk[36]) & (g1593) & (!g1605)) + ((!g1592) & (g1606) & (!sk[36]) & (g1593) & (g1605)) + ((!g1592) & (g1606) & (sk[36]) & (!g1593) & (!g1605)) + ((g1592) & (!g1606) & (!sk[36]) & (!g1593) & (g1605)) + ((g1592) & (!g1606) & (!sk[36]) & (g1593) & (!g1605)) + ((g1592) & (!g1606) & (!sk[36]) & (g1593) & (g1605)) + ((g1592) & (!g1606) & (sk[36]) & (!g1593) & (!g1605)) + ((g1592) & (!g1606) & (sk[36]) & (g1593) & (!g1605)) + ((g1592) & (g1606) & (!sk[36]) & (!g1593) & (!g1605)) + ((g1592) & (g1606) & (!sk[36]) & (!g1593) & (g1605)) + ((g1592) & (g1606) & (!sk[36]) & (g1593) & (!g1605)) + ((g1592) & (g1606) & (!sk[36]) & (g1593) & (g1605)) + ((g1592) & (g1606) & (sk[36]) & (!g1593) & (!g1605)) + ((g1592) & (g1606) & (sk[36]) & (g1593) & (!g1605)));
	assign g2020 = (((!dmem_ack_i) & (!g75) & (!g126) & (g128) & (!sk[37]) & (!g2019)) + ((!dmem_ack_i) & (!g75) & (!g126) & (g128) & (!sk[37]) & (g2019)) + ((!dmem_ack_i) & (!g75) & (g126) & (!g128) & (!sk[37]) & (!g2019)) + ((!dmem_ack_i) & (!g75) & (g126) & (!g128) & (!sk[37]) & (g2019)) + ((!dmem_ack_i) & (!g75) & (g126) & (g128) & (!sk[37]) & (!g2019)) + ((!dmem_ack_i) & (!g75) & (g126) & (g128) & (!sk[37]) & (g2019)) + ((!dmem_ack_i) & (g75) & (!g126) & (!g128) & (!sk[37]) & (!g2019)) + ((!dmem_ack_i) & (g75) & (!g126) & (!g128) & (!sk[37]) & (g2019)) + ((!dmem_ack_i) & (g75) & (!g126) & (g128) & (!sk[37]) & (!g2019)) + ((!dmem_ack_i) & (g75) & (!g126) & (g128) & (!sk[37]) & (g2019)) + ((!dmem_ack_i) & (g75) & (!g126) & (g128) & (sk[37]) & (!g2019)) + ((!dmem_ack_i) & (g75) & (g126) & (!g128) & (!sk[37]) & (!g2019)) + ((!dmem_ack_i) & (g75) & (g126) & (!g128) & (!sk[37]) & (g2019)) + ((!dmem_ack_i) & (g75) & (g126) & (g128) & (!sk[37]) & (!g2019)) + ((!dmem_ack_i) & (g75) & (g126) & (g128) & (!sk[37]) & (g2019)) + ((dmem_ack_i) & (!g75) & (!g126) & (g128) & (!sk[37]) & (!g2019)) + ((dmem_ack_i) & (!g75) & (!g126) & (g128) & (!sk[37]) & (g2019)) + ((dmem_ack_i) & (!g75) & (g126) & (!g128) & (!sk[37]) & (!g2019)) + ((dmem_ack_i) & (!g75) & (g126) & (!g128) & (!sk[37]) & (g2019)) + ((dmem_ack_i) & (!g75) & (g126) & (g128) & (!sk[37]) & (!g2019)) + ((dmem_ack_i) & (!g75) & (g126) & (g128) & (!sk[37]) & (g2019)) + ((dmem_ack_i) & (g75) & (!g126) & (!g128) & (!sk[37]) & (!g2019)) + ((dmem_ack_i) & (g75) & (!g126) & (!g128) & (!sk[37]) & (g2019)) + ((dmem_ack_i) & (g75) & (!g126) & (g128) & (!sk[37]) & (!g2019)) + ((dmem_ack_i) & (g75) & (!g126) & (g128) & (!sk[37]) & (g2019)) + ((dmem_ack_i) & (g75) & (g126) & (!g128) & (!sk[37]) & (!g2019)) + ((dmem_ack_i) & (g75) & (g126) & (!g128) & (!sk[37]) & (g2019)) + ((dmem_ack_i) & (g75) & (g126) & (g128) & (!sk[37]) & (!g2019)) + ((dmem_ack_i) & (g75) & (g126) & (g128) & (!sk[37]) & (g2019)));
	assign g2021 = (((!g74) & (!g132) & (!g134) & (!g136) & (!g126) & (g2020)) + ((!g74) & (!g132) & (!g134) & (!g136) & (g126) & (g2020)) + ((!g74) & (!g132) & (!g134) & (g136) & (!g126) & (g2020)) + ((!g74) & (!g132) & (!g134) & (g136) & (g126) & (!g2020)) + ((!g74) & (!g132) & (!g134) & (g136) & (g126) & (g2020)) + ((!g74) & (!g132) & (g134) & (!g136) & (!g126) & (g2020)) + ((!g74) & (!g132) & (g134) & (!g136) & (g126) & (!g2020)) + ((!g74) & (!g132) & (g134) & (!g136) & (g126) & (g2020)) + ((!g74) & (!g132) & (g134) & (g136) & (!g126) & (g2020)) + ((!g74) & (!g132) & (g134) & (g136) & (g126) & (!g2020)) + ((!g74) & (!g132) & (g134) & (g136) & (g126) & (g2020)) + ((!g74) & (g132) & (!g134) & (!g136) & (!g126) & (g2020)) + ((!g74) & (g132) & (!g134) & (!g136) & (g126) & (!g2020)) + ((!g74) & (g132) & (!g134) & (!g136) & (g126) & (g2020)) + ((!g74) & (g132) & (!g134) & (g136) & (!g126) & (g2020)) + ((!g74) & (g132) & (!g134) & (g136) & (g126) & (!g2020)) + ((!g74) & (g132) & (!g134) & (g136) & (g126) & (g2020)) + ((!g74) & (g132) & (g134) & (!g136) & (!g126) & (g2020)) + ((!g74) & (g132) & (g134) & (!g136) & (g126) & (!g2020)) + ((!g74) & (g132) & (g134) & (!g136) & (g126) & (g2020)) + ((!g74) & (g132) & (g134) & (g136) & (!g126) & (g2020)) + ((!g74) & (g132) & (g134) & (g136) & (g126) & (!g2020)) + ((!g74) & (g132) & (g134) & (g136) & (g126) & (g2020)));
	assign g2022 = (((!g114) & (sk[39]) & (!g115)) + ((!g114) & (sk[39]) & (g115)) + ((g114) & (!sk[39]) & (!g115)) + ((g114) & (!sk[39]) & (g115)) + ((g114) & (sk[39]) & (!g115)));
	assign g2024 = (((!g78) & (!g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((!g78) & (g79) & (!g80) & (g81) & (!g82) & (!g83)));
	assign g2025 = (((!g78) & (g79) & (!g80) & (!g81) & (!g82) & (g83)));
	assign g5018 = (((!g2059) & (!sk[42]) & (!g2917) & (g2026)) + ((!g2059) & (!sk[42]) & (g2917) & (!g2026)) + ((!g2059) & (!sk[42]) & (g2917) & (g2026)) + ((!g2059) & (sk[42]) & (!g2917) & (g2026)) + ((!g2059) & (sk[42]) & (g2917) & (g2026)) + ((g2059) & (!sk[42]) & (!g2917) & (g2026)) + ((g2059) & (!sk[42]) & (g2917) & (!g2026)) + ((g2059) & (!sk[42]) & (g2917) & (g2026)) + ((g2059) & (sk[42]) & (g2917) & (!g2026)) + ((g2059) & (sk[42]) & (g2917) & (g2026)));
	assign g2027 = (((!sk[43]) & (!g79) & (!g80) & (!g81) & (g133) & (!g2026)) + ((!sk[43]) & (!g79) & (!g80) & (!g81) & (g133) & (g2026)) + ((!sk[43]) & (!g79) & (!g80) & (g81) & (!g133) & (!g2026)) + ((!sk[43]) & (!g79) & (!g80) & (g81) & (!g133) & (g2026)) + ((!sk[43]) & (!g79) & (!g80) & (g81) & (g133) & (!g2026)) + ((!sk[43]) & (!g79) & (!g80) & (g81) & (g133) & (g2026)) + ((!sk[43]) & (!g79) & (g80) & (!g81) & (!g133) & (!g2026)) + ((!sk[43]) & (!g79) & (g80) & (!g81) & (!g133) & (g2026)) + ((!sk[43]) & (!g79) & (g80) & (!g81) & (g133) & (!g2026)) + ((!sk[43]) & (!g79) & (g80) & (!g81) & (g133) & (g2026)) + ((!sk[43]) & (!g79) & (g80) & (g81) & (!g133) & (!g2026)) + ((!sk[43]) & (!g79) & (g80) & (g81) & (!g133) & (g2026)) + ((!sk[43]) & (!g79) & (g80) & (g81) & (g133) & (!g2026)) + ((!sk[43]) & (!g79) & (g80) & (g81) & (g133) & (g2026)) + ((!sk[43]) & (g79) & (!g80) & (!g81) & (g133) & (!g2026)) + ((!sk[43]) & (g79) & (!g80) & (!g81) & (g133) & (g2026)) + ((!sk[43]) & (g79) & (!g80) & (g81) & (!g133) & (!g2026)) + ((!sk[43]) & (g79) & (!g80) & (g81) & (!g133) & (g2026)) + ((!sk[43]) & (g79) & (!g80) & (g81) & (g133) & (!g2026)) + ((!sk[43]) & (g79) & (!g80) & (g81) & (g133) & (g2026)) + ((!sk[43]) & (g79) & (g80) & (!g81) & (!g133) & (!g2026)) + ((!sk[43]) & (g79) & (g80) & (!g81) & (!g133) & (g2026)) + ((!sk[43]) & (g79) & (g80) & (!g81) & (g133) & (!g2026)) + ((!sk[43]) & (g79) & (g80) & (!g81) & (g133) & (g2026)) + ((!sk[43]) & (g79) & (g80) & (g81) & (!g133) & (!g2026)) + ((!sk[43]) & (g79) & (g80) & (g81) & (!g133) & (g2026)) + ((!sk[43]) & (g79) & (g80) & (g81) & (g133) & (!g2026)) + ((!sk[43]) & (g79) & (g80) & (g81) & (g133) & (g2026)) + ((sk[43]) & (!g79) & (!g80) & (!g81) & (g133) & (g2026)));
	assign g2028 = (((!sk[44]) & (!g2024) & (!g2025) & (!g117) & (g2026) & (!g2027)) + ((!sk[44]) & (!g2024) & (!g2025) & (!g117) & (g2026) & (g2027)) + ((!sk[44]) & (!g2024) & (!g2025) & (g117) & (!g2026) & (!g2027)) + ((!sk[44]) & (!g2024) & (!g2025) & (g117) & (!g2026) & (g2027)) + ((!sk[44]) & (!g2024) & (!g2025) & (g117) & (g2026) & (!g2027)) + ((!sk[44]) & (!g2024) & (!g2025) & (g117) & (g2026) & (g2027)) + ((!sk[44]) & (!g2024) & (g2025) & (!g117) & (!g2026) & (!g2027)) + ((!sk[44]) & (!g2024) & (g2025) & (!g117) & (!g2026) & (g2027)) + ((!sk[44]) & (!g2024) & (g2025) & (!g117) & (g2026) & (!g2027)) + ((!sk[44]) & (!g2024) & (g2025) & (!g117) & (g2026) & (g2027)) + ((!sk[44]) & (!g2024) & (g2025) & (g117) & (!g2026) & (!g2027)) + ((!sk[44]) & (!g2024) & (g2025) & (g117) & (!g2026) & (g2027)) + ((!sk[44]) & (!g2024) & (g2025) & (g117) & (g2026) & (!g2027)) + ((!sk[44]) & (!g2024) & (g2025) & (g117) & (g2026) & (g2027)) + ((!sk[44]) & (g2024) & (!g2025) & (!g117) & (g2026) & (!g2027)) + ((!sk[44]) & (g2024) & (!g2025) & (!g117) & (g2026) & (g2027)) + ((!sk[44]) & (g2024) & (!g2025) & (g117) & (!g2026) & (!g2027)) + ((!sk[44]) & (g2024) & (!g2025) & (g117) & (!g2026) & (g2027)) + ((!sk[44]) & (g2024) & (!g2025) & (g117) & (g2026) & (!g2027)) + ((!sk[44]) & (g2024) & (!g2025) & (g117) & (g2026) & (g2027)) + ((!sk[44]) & (g2024) & (g2025) & (!g117) & (!g2026) & (!g2027)) + ((!sk[44]) & (g2024) & (g2025) & (!g117) & (!g2026) & (g2027)) + ((!sk[44]) & (g2024) & (g2025) & (!g117) & (g2026) & (!g2027)) + ((!sk[44]) & (g2024) & (g2025) & (!g117) & (g2026) & (g2027)) + ((!sk[44]) & (g2024) & (g2025) & (g117) & (!g2026) & (!g2027)) + ((!sk[44]) & (g2024) & (g2025) & (g117) & (!g2026) & (g2027)) + ((!sk[44]) & (g2024) & (g2025) & (g117) & (g2026) & (!g2027)) + ((!sk[44]) & (g2024) & (g2025) & (g117) & (g2026) & (g2027)) + ((sk[44]) & (!g2024) & (!g2025) & (!g117) & (!g2026) & (!g2027)) + ((sk[44]) & (!g2024) & (!g2025) & (!g117) & (!g2026) & (g2027)) + ((sk[44]) & (!g2024) & (!g2025) & (!g117) & (g2026) & (!g2027)) + ((sk[44]) & (!g2024) & (!g2025) & (!g117) & (g2026) & (g2027)) + ((sk[44]) & (!g2024) & (!g2025) & (g117) & (!g2026) & (g2027)) + ((sk[44]) & (!g2024) & (!g2025) & (g117) & (g2026) & (g2027)) + ((sk[44]) & (!g2024) & (g2025) & (!g117) & (!g2026) & (!g2027)) + ((sk[44]) & (!g2024) & (g2025) & (!g117) & (!g2026) & (g2027)) + ((sk[44]) & (!g2024) & (g2025) & (!g117) & (g2026) & (!g2027)) + ((sk[44]) & (!g2024) & (g2025) & (!g117) & (g2026) & (g2027)) + ((sk[44]) & (!g2024) & (g2025) & (g117) & (!g2026) & (!g2027)) + ((sk[44]) & (!g2024) & (g2025) & (g117) & (!g2026) & (g2027)) + ((sk[44]) & (!g2024) & (g2025) & (g117) & (g2026) & (g2027)) + ((sk[44]) & (g2024) & (!g2025) & (!g117) & (!g2026) & (!g2027)) + ((sk[44]) & (g2024) & (!g2025) & (!g117) & (!g2026) & (g2027)) + ((sk[44]) & (g2024) & (!g2025) & (!g117) & (g2026) & (!g2027)) + ((sk[44]) & (g2024) & (!g2025) & (!g117) & (g2026) & (g2027)) + ((sk[44]) & (g2024) & (!g2025) & (g117) & (!g2026) & (!g2027)) + ((sk[44]) & (g2024) & (!g2025) & (g117) & (!g2026) & (g2027)) + ((sk[44]) & (g2024) & (!g2025) & (g117) & (g2026) & (!g2027)) + ((sk[44]) & (g2024) & (!g2025) & (g117) & (g2026) & (g2027)) + ((sk[44]) & (g2024) & (g2025) & (!g117) & (!g2026) & (!g2027)) + ((sk[44]) & (g2024) & (g2025) & (!g117) & (!g2026) & (g2027)) + ((sk[44]) & (g2024) & (g2025) & (!g117) & (g2026) & (!g2027)) + ((sk[44]) & (g2024) & (g2025) & (!g117) & (g2026) & (g2027)) + ((sk[44]) & (g2024) & (g2025) & (g117) & (!g2026) & (!g2027)) + ((sk[44]) & (g2024) & (g2025) & (g117) & (!g2026) & (g2027)) + ((sk[44]) & (g2024) & (g2025) & (g117) & (g2026) & (!g2027)) + ((sk[44]) & (g2024) & (g2025) & (g117) & (g2026) & (g2027)));
	assign g2029 = (((g2022) & (!sk[45]) & (!g2028)) + ((g2022) & (!sk[45]) & (g2028)) + ((g2022) & (sk[45]) & (!g2028)));
	assign g2030 = (((!g82) & (!sk[46]) & (!g83) & (g114)) + ((!g82) & (!sk[46]) & (g83) & (!g114)) + ((!g82) & (!sk[46]) & (g83) & (g114)) + ((g82) & (!sk[46]) & (!g83) & (g114)) + ((g82) & (!sk[46]) & (g83) & (!g114)) + ((g82) & (!sk[46]) & (g83) & (g114)) + ((g82) & (sk[46]) & (g83) & (g114)));
	assign g2031 = (((!g78) & (!g79) & (!g80) & (g81) & (!g82) & (g83)) + ((!g78) & (g79) & (!g80) & (g81) & (!g82) & (!g83)));
	assign g2032 = (((!g78) & (!g79) & (!g80) & (!g81) & (!g82) & (!g83)) + ((!g78) & (!g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((!g78) & (g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((g78) & (!g79) & (!g80) & (!g81) & (!g82) & (!g83)));
	assign g2033 = (((!g2030) & (!g2031) & (!sk[49]) & (g2032)) + ((!g2030) & (!g2031) & (sk[49]) & (!g2032)) + ((!g2030) & (!g2031) & (sk[49]) & (g2032)) + ((!g2030) & (g2031) & (!sk[49]) & (!g2032)) + ((!g2030) & (g2031) & (!sk[49]) & (g2032)) + ((!g2030) & (g2031) & (sk[49]) & (g2032)) + ((g2030) & (!g2031) & (!sk[49]) & (g2032)) + ((g2030) & (!g2031) & (sk[49]) & (g2032)) + ((g2030) & (g2031) & (!sk[49]) & (!g2032)) + ((g2030) & (g2031) & (!sk[49]) & (g2032)) + ((g2030) & (g2031) & (sk[49]) & (g2032)));
	assign g2034 = (((!sk[50]) & (g2022) & (!g2031)) + ((!sk[50]) & (g2022) & (g2031)) + ((sk[50]) & (!g2022) & (!g2031)) + ((sk[50]) & (!g2022) & (g2031)) + ((sk[50]) & (g2022) & (g2031)));
	assign g5019 = (((!g2921) & (!sk[51]) & (!g2918) & (g2035)) + ((!g2921) & (!sk[51]) & (g2918) & (!g2035)) + ((!g2921) & (!sk[51]) & (g2918) & (g2035)) + ((!g2921) & (sk[51]) & (!g2918) & (g2035)) + ((!g2921) & (sk[51]) & (g2918) & (g2035)) + ((g2921) & (!sk[51]) & (!g2918) & (g2035)) + ((g2921) & (!sk[51]) & (g2918) & (!g2035)) + ((g2921) & (!sk[51]) & (g2918) & (g2035)) + ((g2921) & (sk[51]) & (g2918) & (!g2035)) + ((g2921) & (sk[51]) & (g2918) & (g2035)));
	assign g2036 = (((!g76) & (!g1620) & (!g2033) & (!sk[52]) & (g2034) & (!g2035)) + ((!g76) & (!g1620) & (!g2033) & (!sk[52]) & (g2034) & (g2035)) + ((!g76) & (!g1620) & (!g2033) & (sk[52]) & (!g2034) & (g2035)) + ((!g76) & (!g1620) & (g2033) & (!sk[52]) & (!g2034) & (!g2035)) + ((!g76) & (!g1620) & (g2033) & (!sk[52]) & (!g2034) & (g2035)) + ((!g76) & (!g1620) & (g2033) & (!sk[52]) & (g2034) & (!g2035)) + ((!g76) & (!g1620) & (g2033) & (!sk[52]) & (g2034) & (g2035)) + ((!g76) & (g1620) & (!g2033) & (!sk[52]) & (!g2034) & (!g2035)) + ((!g76) & (g1620) & (!g2033) & (!sk[52]) & (!g2034) & (g2035)) + ((!g76) & (g1620) & (!g2033) & (!sk[52]) & (g2034) & (!g2035)) + ((!g76) & (g1620) & (!g2033) & (!sk[52]) & (g2034) & (g2035)) + ((!g76) & (g1620) & (!g2033) & (sk[52]) & (!g2034) & (g2035)) + ((!g76) & (g1620) & (!g2033) & (sk[52]) & (g2034) & (!g2035)) + ((!g76) & (g1620) & (!g2033) & (sk[52]) & (g2034) & (g2035)) + ((!g76) & (g1620) & (g2033) & (!sk[52]) & (!g2034) & (!g2035)) + ((!g76) & (g1620) & (g2033) & (!sk[52]) & (!g2034) & (g2035)) + ((!g76) & (g1620) & (g2033) & (!sk[52]) & (g2034) & (!g2035)) + ((!g76) & (g1620) & (g2033) & (!sk[52]) & (g2034) & (g2035)) + ((g76) & (!g1620) & (!g2033) & (!sk[52]) & (g2034) & (!g2035)) + ((g76) & (!g1620) & (!g2033) & (!sk[52]) & (g2034) & (g2035)) + ((g76) & (!g1620) & (!g2033) & (sk[52]) & (!g2034) & (g2035)) + ((g76) & (!g1620) & (g2033) & (!sk[52]) & (!g2034) & (!g2035)) + ((g76) & (!g1620) & (g2033) & (!sk[52]) & (!g2034) & (g2035)) + ((g76) & (!g1620) & (g2033) & (!sk[52]) & (g2034) & (!g2035)) + ((g76) & (!g1620) & (g2033) & (!sk[52]) & (g2034) & (g2035)) + ((g76) & (!g1620) & (g2033) & (sk[52]) & (!g2034) & (!g2035)) + ((g76) & (!g1620) & (g2033) & (sk[52]) & (!g2034) & (g2035)) + ((g76) & (g1620) & (!g2033) & (!sk[52]) & (!g2034) & (!g2035)) + ((g76) & (g1620) & (!g2033) & (!sk[52]) & (!g2034) & (g2035)) + ((g76) & (g1620) & (!g2033) & (!sk[52]) & (g2034) & (!g2035)) + ((g76) & (g1620) & (!g2033) & (!sk[52]) & (g2034) & (g2035)) + ((g76) & (g1620) & (!g2033) & (sk[52]) & (!g2034) & (g2035)) + ((g76) & (g1620) & (!g2033) & (sk[52]) & (g2034) & (!g2035)) + ((g76) & (g1620) & (!g2033) & (sk[52]) & (g2034) & (g2035)) + ((g76) & (g1620) & (g2033) & (!sk[52]) & (!g2034) & (!g2035)) + ((g76) & (g1620) & (g2033) & (!sk[52]) & (!g2034) & (g2035)) + ((g76) & (g1620) & (g2033) & (!sk[52]) & (g2034) & (!g2035)) + ((g76) & (g1620) & (g2033) & (!sk[52]) & (g2034) & (g2035)) + ((g76) & (g1620) & (g2033) & (sk[52]) & (!g2034) & (!g2035)) + ((g76) & (g1620) & (g2033) & (sk[52]) & (!g2034) & (g2035)));
	assign g2037 = (((!g2022) & (!g76) & (!nmi_i) & (!g2023) & (!g2029) & (g2036)) + ((!g2022) & (!g76) & (!nmi_i) & (g2023) & (!g2029) & (g2036)) + ((!g2022) & (!g76) & (nmi_i) & (!g2023) & (!g2029) & (g2036)) + ((!g2022) & (!g76) & (nmi_i) & (g2023) & (!g2029) & (g2036)) + ((!g2022) & (g76) & (!nmi_i) & (!g2023) & (!g2029) & (g2036)) + ((!g2022) & (g76) & (!nmi_i) & (!g2023) & (g2029) & (!g2036)) + ((!g2022) & (g76) & (!nmi_i) & (!g2023) & (g2029) & (g2036)) + ((!g2022) & (g76) & (!nmi_i) & (g2023) & (!g2029) & (g2036)) + ((!g2022) & (g76) & (!nmi_i) & (g2023) & (g2029) & (!g2036)) + ((!g2022) & (g76) & (!nmi_i) & (g2023) & (g2029) & (g2036)) + ((!g2022) & (g76) & (nmi_i) & (!g2023) & (!g2029) & (g2036)) + ((!g2022) & (g76) & (nmi_i) & (!g2023) & (g2029) & (!g2036)) + ((!g2022) & (g76) & (nmi_i) & (!g2023) & (g2029) & (g2036)) + ((!g2022) & (g76) & (nmi_i) & (g2023) & (!g2029) & (g2036)) + ((!g2022) & (g76) & (nmi_i) & (g2023) & (g2029) & (!g2036)) + ((!g2022) & (g76) & (nmi_i) & (g2023) & (g2029) & (g2036)) + ((g2022) & (!g76) & (!nmi_i) & (!g2023) & (!g2029) & (g2036)) + ((g2022) & (g76) & (!nmi_i) & (!g2023) & (!g2029) & (g2036)) + ((g2022) & (g76) & (!nmi_i) & (!g2023) & (g2029) & (!g2036)) + ((g2022) & (g76) & (!nmi_i) & (!g2023) & (g2029) & (g2036)));
	assign g5020 = (((!g2924) & (!sk[54]) & (!g2922) & (g2038)) + ((!g2924) & (!sk[54]) & (g2922) & (!g2038)) + ((!g2924) & (!sk[54]) & (g2922) & (g2038)) + ((!g2924) & (sk[54]) & (!g2922) & (g2038)) + ((!g2924) & (sk[54]) & (g2922) & (g2038)) + ((g2924) & (!sk[54]) & (!g2922) & (g2038)) + ((g2924) & (!sk[54]) & (g2922) & (!g2038)) + ((g2924) & (!sk[54]) & (g2922) & (g2038)) + ((g2924) & (sk[54]) & (g2922) & (!g2038)) + ((g2924) & (sk[54]) & (g2922) & (g2038)));
	assign g2039 = (((g2030) & (!sk[55]) & (!g2038)) + ((g2030) & (!sk[55]) & (g2038)) + ((g2030) & (sk[55]) & (g2038)));
	assign g2040 = (((!g78) & (!g79) & (g80) & (g81) & (!g82) & (!g83)));
	assign g2041 = (((!g142) & (!sk[57]) & (!g702) & (!g722) & (g651) & (!g671)) + ((!g142) & (!sk[57]) & (!g702) & (!g722) & (g651) & (g671)) + ((!g142) & (!sk[57]) & (!g702) & (g722) & (!g651) & (!g671)) + ((!g142) & (!sk[57]) & (!g702) & (g722) & (!g651) & (g671)) + ((!g142) & (!sk[57]) & (!g702) & (g722) & (g651) & (!g671)) + ((!g142) & (!sk[57]) & (!g702) & (g722) & (g651) & (g671)) + ((!g142) & (!sk[57]) & (g702) & (!g722) & (!g651) & (!g671)) + ((!g142) & (!sk[57]) & (g702) & (!g722) & (!g651) & (g671)) + ((!g142) & (!sk[57]) & (g702) & (!g722) & (g651) & (!g671)) + ((!g142) & (!sk[57]) & (g702) & (!g722) & (g651) & (g671)) + ((!g142) & (!sk[57]) & (g702) & (g722) & (!g651) & (!g671)) + ((!g142) & (!sk[57]) & (g702) & (g722) & (!g651) & (g671)) + ((!g142) & (!sk[57]) & (g702) & (g722) & (g651) & (!g671)) + ((!g142) & (!sk[57]) & (g702) & (g722) & (g651) & (g671)) + ((!g142) & (sk[57]) & (!g702) & (!g722) & (!g651) & (!g671)) + ((!g142) & (sk[57]) & (!g702) & (!g722) & (g651) & (!g671)) + ((!g142) & (sk[57]) & (g702) & (!g722) & (!g651) & (!g671)) + ((!g142) & (sk[57]) & (g702) & (!g722) & (g651) & (!g671)) + ((g142) & (!sk[57]) & (!g702) & (!g722) & (g651) & (!g671)) + ((g142) & (!sk[57]) & (!g702) & (!g722) & (g651) & (g671)) + ((g142) & (!sk[57]) & (!g702) & (g722) & (!g651) & (!g671)) + ((g142) & (!sk[57]) & (!g702) & (g722) & (!g651) & (g671)) + ((g142) & (!sk[57]) & (!g702) & (g722) & (g651) & (!g671)) + ((g142) & (!sk[57]) & (!g702) & (g722) & (g651) & (g671)) + ((g142) & (!sk[57]) & (g702) & (!g722) & (!g651) & (!g671)) + ((g142) & (!sk[57]) & (g702) & (!g722) & (!g651) & (g671)) + ((g142) & (!sk[57]) & (g702) & (!g722) & (g651) & (!g671)) + ((g142) & (!sk[57]) & (g702) & (!g722) & (g651) & (g671)) + ((g142) & (!sk[57]) & (g702) & (g722) & (!g651) & (!g671)) + ((g142) & (!sk[57]) & (g702) & (g722) & (!g651) & (g671)) + ((g142) & (!sk[57]) & (g702) & (g722) & (g651) & (!g671)) + ((g142) & (!sk[57]) & (g702) & (g722) & (g651) & (g671)) + ((g142) & (sk[57]) & (!g702) & (!g722) & (!g651) & (!g671)) + ((g142) & (sk[57]) & (!g702) & (!g722) & (!g651) & (g671)) + ((g142) & (sk[57]) & (!g702) & (g722) & (!g651) & (!g671)) + ((g142) & (sk[57]) & (!g702) & (g722) & (!g651) & (g671)));
	assign g2042 = (((!sk[58]) & (!g142) & (!g796) & (!g816) & (g749) & (!g769)) + ((!sk[58]) & (!g142) & (!g796) & (!g816) & (g749) & (g769)) + ((!sk[58]) & (!g142) & (!g796) & (g816) & (!g749) & (!g769)) + ((!sk[58]) & (!g142) & (!g796) & (g816) & (!g749) & (g769)) + ((!sk[58]) & (!g142) & (!g796) & (g816) & (g749) & (!g769)) + ((!sk[58]) & (!g142) & (!g796) & (g816) & (g749) & (g769)) + ((!sk[58]) & (!g142) & (g796) & (!g816) & (!g749) & (!g769)) + ((!sk[58]) & (!g142) & (g796) & (!g816) & (!g749) & (g769)) + ((!sk[58]) & (!g142) & (g796) & (!g816) & (g749) & (!g769)) + ((!sk[58]) & (!g142) & (g796) & (!g816) & (g749) & (g769)) + ((!sk[58]) & (!g142) & (g796) & (g816) & (!g749) & (!g769)) + ((!sk[58]) & (!g142) & (g796) & (g816) & (!g749) & (g769)) + ((!sk[58]) & (!g142) & (g796) & (g816) & (g749) & (!g769)) + ((!sk[58]) & (!g142) & (g796) & (g816) & (g749) & (g769)) + ((!sk[58]) & (g142) & (!g796) & (!g816) & (g749) & (!g769)) + ((!sk[58]) & (g142) & (!g796) & (!g816) & (g749) & (g769)) + ((!sk[58]) & (g142) & (!g796) & (g816) & (!g749) & (!g769)) + ((!sk[58]) & (g142) & (!g796) & (g816) & (!g749) & (g769)) + ((!sk[58]) & (g142) & (!g796) & (g816) & (g749) & (!g769)) + ((!sk[58]) & (g142) & (!g796) & (g816) & (g749) & (g769)) + ((!sk[58]) & (g142) & (g796) & (!g816) & (!g749) & (!g769)) + ((!sk[58]) & (g142) & (g796) & (!g816) & (!g749) & (g769)) + ((!sk[58]) & (g142) & (g796) & (!g816) & (g749) & (!g769)) + ((!sk[58]) & (g142) & (g796) & (!g816) & (g749) & (g769)) + ((!sk[58]) & (g142) & (g796) & (g816) & (!g749) & (!g769)) + ((!sk[58]) & (g142) & (g796) & (g816) & (!g749) & (g769)) + ((!sk[58]) & (g142) & (g796) & (g816) & (g749) & (!g769)) + ((!sk[58]) & (g142) & (g796) & (g816) & (g749) & (g769)) + ((sk[58]) & (!g142) & (!g796) & (!g816) & (!g749) & (!g769)) + ((sk[58]) & (!g142) & (!g796) & (!g816) & (g749) & (!g769)) + ((sk[58]) & (!g142) & (g796) & (!g816) & (!g749) & (!g769)) + ((sk[58]) & (!g142) & (g796) & (!g816) & (g749) & (!g769)) + ((sk[58]) & (g142) & (!g796) & (!g816) & (!g749) & (!g769)) + ((sk[58]) & (g142) & (!g796) & (!g816) & (!g749) & (g769)) + ((sk[58]) & (g142) & (!g796) & (g816) & (!g749) & (!g769)) + ((sk[58]) & (g142) & (!g796) & (g816) & (!g749) & (g769)));
	assign g2043 = (((!g142) & (!g608) & (!g628) & (!sk[59]) & (g843) & (!g863)) + ((!g142) & (!g608) & (!g628) & (!sk[59]) & (g843) & (g863)) + ((!g142) & (!g608) & (!g628) & (sk[59]) & (!g843) & (!g863)) + ((!g142) & (!g608) & (!g628) & (sk[59]) & (g843) & (!g863)) + ((!g142) & (!g608) & (g628) & (!sk[59]) & (!g843) & (!g863)) + ((!g142) & (!g608) & (g628) & (!sk[59]) & (!g843) & (g863)) + ((!g142) & (!g608) & (g628) & (!sk[59]) & (g843) & (!g863)) + ((!g142) & (!g608) & (g628) & (!sk[59]) & (g843) & (g863)) + ((!g142) & (g608) & (!g628) & (!sk[59]) & (!g843) & (!g863)) + ((!g142) & (g608) & (!g628) & (!sk[59]) & (!g843) & (g863)) + ((!g142) & (g608) & (!g628) & (!sk[59]) & (g843) & (!g863)) + ((!g142) & (g608) & (!g628) & (!sk[59]) & (g843) & (g863)) + ((!g142) & (g608) & (!g628) & (sk[59]) & (!g843) & (!g863)) + ((!g142) & (g608) & (!g628) & (sk[59]) & (g843) & (!g863)) + ((!g142) & (g608) & (g628) & (!sk[59]) & (!g843) & (!g863)) + ((!g142) & (g608) & (g628) & (!sk[59]) & (!g843) & (g863)) + ((!g142) & (g608) & (g628) & (!sk[59]) & (g843) & (!g863)) + ((!g142) & (g608) & (g628) & (!sk[59]) & (g843) & (g863)) + ((g142) & (!g608) & (!g628) & (!sk[59]) & (g843) & (!g863)) + ((g142) & (!g608) & (!g628) & (!sk[59]) & (g843) & (g863)) + ((g142) & (!g608) & (!g628) & (sk[59]) & (!g843) & (!g863)) + ((g142) & (!g608) & (!g628) & (sk[59]) & (!g843) & (g863)) + ((g142) & (!g608) & (g628) & (!sk[59]) & (!g843) & (!g863)) + ((g142) & (!g608) & (g628) & (!sk[59]) & (!g843) & (g863)) + ((g142) & (!g608) & (g628) & (!sk[59]) & (g843) & (!g863)) + ((g142) & (!g608) & (g628) & (!sk[59]) & (g843) & (g863)) + ((g142) & (!g608) & (g628) & (sk[59]) & (!g843) & (!g863)) + ((g142) & (!g608) & (g628) & (sk[59]) & (!g843) & (g863)) + ((g142) & (g608) & (!g628) & (!sk[59]) & (!g843) & (!g863)) + ((g142) & (g608) & (!g628) & (!sk[59]) & (!g843) & (g863)) + ((g142) & (g608) & (!g628) & (!sk[59]) & (g843) & (!g863)) + ((g142) & (g608) & (!g628) & (!sk[59]) & (g843) & (g863)) + ((g142) & (g608) & (g628) & (!sk[59]) & (!g843) & (!g863)) + ((g142) & (g608) & (g628) & (!sk[59]) & (!g843) & (g863)) + ((g142) & (g608) & (g628) & (!sk[59]) & (g843) & (!g863)) + ((g142) & (g608) & (g628) & (!sk[59]) & (g843) & (g863)));
	assign g2044 = (((!g142) & (!g518) & (!g538) & (!sk[60]) & (g563) & (!g583)) + ((!g142) & (!g518) & (!g538) & (!sk[60]) & (g563) & (g583)) + ((!g142) & (!g518) & (!g538) & (sk[60]) & (!g563) & (!g583)) + ((!g142) & (!g518) & (!g538) & (sk[60]) & (g563) & (!g583)) + ((!g142) & (!g518) & (g538) & (!sk[60]) & (!g563) & (!g583)) + ((!g142) & (!g518) & (g538) & (!sk[60]) & (!g563) & (g583)) + ((!g142) & (!g518) & (g538) & (!sk[60]) & (g563) & (!g583)) + ((!g142) & (!g518) & (g538) & (!sk[60]) & (g563) & (g583)) + ((!g142) & (g518) & (!g538) & (!sk[60]) & (!g563) & (!g583)) + ((!g142) & (g518) & (!g538) & (!sk[60]) & (!g563) & (g583)) + ((!g142) & (g518) & (!g538) & (!sk[60]) & (g563) & (!g583)) + ((!g142) & (g518) & (!g538) & (!sk[60]) & (g563) & (g583)) + ((!g142) & (g518) & (!g538) & (sk[60]) & (!g563) & (!g583)) + ((!g142) & (g518) & (!g538) & (sk[60]) & (g563) & (!g583)) + ((!g142) & (g518) & (g538) & (!sk[60]) & (!g563) & (!g583)) + ((!g142) & (g518) & (g538) & (!sk[60]) & (!g563) & (g583)) + ((!g142) & (g518) & (g538) & (!sk[60]) & (g563) & (!g583)) + ((!g142) & (g518) & (g538) & (!sk[60]) & (g563) & (g583)) + ((g142) & (!g518) & (!g538) & (!sk[60]) & (g563) & (!g583)) + ((g142) & (!g518) & (!g538) & (!sk[60]) & (g563) & (g583)) + ((g142) & (!g518) & (!g538) & (sk[60]) & (!g563) & (!g583)) + ((g142) & (!g518) & (!g538) & (sk[60]) & (!g563) & (g583)) + ((g142) & (!g518) & (g538) & (!sk[60]) & (!g563) & (!g583)) + ((g142) & (!g518) & (g538) & (!sk[60]) & (!g563) & (g583)) + ((g142) & (!g518) & (g538) & (!sk[60]) & (g563) & (!g583)) + ((g142) & (!g518) & (g538) & (!sk[60]) & (g563) & (g583)) + ((g142) & (!g518) & (g538) & (sk[60]) & (!g563) & (!g583)) + ((g142) & (!g518) & (g538) & (sk[60]) & (!g563) & (g583)) + ((g142) & (g518) & (!g538) & (!sk[60]) & (!g563) & (!g583)) + ((g142) & (g518) & (!g538) & (!sk[60]) & (!g563) & (g583)) + ((g142) & (g518) & (!g538) & (!sk[60]) & (g563) & (!g583)) + ((g142) & (g518) & (!g538) & (!sk[60]) & (g563) & (g583)) + ((g142) & (g518) & (g538) & (!sk[60]) & (!g563) & (!g583)) + ((g142) & (g518) & (g538) & (!sk[60]) & (!g563) & (g583)) + ((g142) & (g518) & (g538) & (!sk[60]) & (g563) & (!g583)) + ((g142) & (g518) & (g538) & (!sk[60]) & (g563) & (g583)));
	assign g2045 = (((!g87) & (!sk[61]) & (!g88) & (!g91) & (g92)) + ((!g87) & (!sk[61]) & (!g88) & (g91) & (!g92)) + ((!g87) & (!sk[61]) & (!g88) & (g91) & (g92)) + ((!g87) & (!sk[61]) & (g88) & (!g91) & (!g92)) + ((!g87) & (!sk[61]) & (g88) & (!g91) & (g92)) + ((!g87) & (!sk[61]) & (g88) & (g91) & (!g92)) + ((!g87) & (!sk[61]) & (g88) & (g91) & (g92)) + ((!g87) & (sk[61]) & (!g88) & (!g91) & (!g92)) + ((g87) & (!sk[61]) & (!g88) & (!g91) & (g92)) + ((g87) & (!sk[61]) & (!g88) & (g91) & (!g92)) + ((g87) & (!sk[61]) & (!g88) & (g91) & (g92)) + ((g87) & (!sk[61]) & (g88) & (!g91) & (!g92)) + ((g87) & (!sk[61]) & (g88) & (!g91) & (g92)) + ((g87) & (!sk[61]) & (g88) & (g91) & (!g92)) + ((g87) & (!sk[61]) & (g88) & (g91) & (g92)));
	assign g2046 = (((!sk[62]) & (!g85) & (!g90) & (!g2045) & (g586)) + ((!sk[62]) & (!g85) & (!g90) & (g2045) & (!g586)) + ((!sk[62]) & (!g85) & (!g90) & (g2045) & (g586)) + ((!sk[62]) & (!g85) & (g90) & (!g2045) & (!g586)) + ((!sk[62]) & (!g85) & (g90) & (!g2045) & (g586)) + ((!sk[62]) & (!g85) & (g90) & (g2045) & (!g586)) + ((!sk[62]) & (!g85) & (g90) & (g2045) & (g586)) + ((!sk[62]) & (g85) & (!g90) & (!g2045) & (g586)) + ((!sk[62]) & (g85) & (!g90) & (g2045) & (!g586)) + ((!sk[62]) & (g85) & (!g90) & (g2045) & (g586)) + ((!sk[62]) & (g85) & (g90) & (!g2045) & (!g586)) + ((!sk[62]) & (g85) & (g90) & (!g2045) & (g586)) + ((!sk[62]) & (g85) & (g90) & (g2045) & (!g586)) + ((!sk[62]) & (g85) & (g90) & (g2045) & (g586)) + ((sk[62]) & (!g85) & (!g90) & (g2045) & (!g586)));
	assign g2047 = (((!g142) & (!g209) & (!g229) & (!g252) & (!g272) & (g2046)) + ((!g142) & (!g209) & (!g229) & (g252) & (!g272) & (g2046)) + ((!g142) & (g209) & (!g229) & (!g252) & (!g272) & (g2046)) + ((!g142) & (g209) & (!g229) & (g252) & (!g272) & (g2046)) + ((g142) & (!g209) & (!g229) & (!g252) & (!g272) & (g2046)) + ((g142) & (!g209) & (!g229) & (!g252) & (g272) & (g2046)) + ((g142) & (!g209) & (g229) & (!g252) & (!g272) & (g2046)) + ((g142) & (!g209) & (g229) & (!g252) & (g272) & (g2046)));
	assign g2048 = (((!g142) & (!g296) & (!sk[64]) & (!g316) & (g474) & (!g494)) + ((!g142) & (!g296) & (!sk[64]) & (!g316) & (g474) & (g494)) + ((!g142) & (!g296) & (!sk[64]) & (g316) & (!g474) & (!g494)) + ((!g142) & (!g296) & (!sk[64]) & (g316) & (!g474) & (g494)) + ((!g142) & (!g296) & (!sk[64]) & (g316) & (g474) & (!g494)) + ((!g142) & (!g296) & (!sk[64]) & (g316) & (g474) & (g494)) + ((!g142) & (!g296) & (sk[64]) & (!g316) & (!g474) & (!g494)) + ((!g142) & (!g296) & (sk[64]) & (!g316) & (g474) & (!g494)) + ((!g142) & (g296) & (!sk[64]) & (!g316) & (!g474) & (!g494)) + ((!g142) & (g296) & (!sk[64]) & (!g316) & (!g474) & (g494)) + ((!g142) & (g296) & (!sk[64]) & (!g316) & (g474) & (!g494)) + ((!g142) & (g296) & (!sk[64]) & (!g316) & (g474) & (g494)) + ((!g142) & (g296) & (!sk[64]) & (g316) & (!g474) & (!g494)) + ((!g142) & (g296) & (!sk[64]) & (g316) & (!g474) & (g494)) + ((!g142) & (g296) & (!sk[64]) & (g316) & (g474) & (!g494)) + ((!g142) & (g296) & (!sk[64]) & (g316) & (g474) & (g494)) + ((!g142) & (g296) & (sk[64]) & (!g316) & (!g474) & (!g494)) + ((!g142) & (g296) & (sk[64]) & (!g316) & (g474) & (!g494)) + ((g142) & (!g296) & (!sk[64]) & (!g316) & (g474) & (!g494)) + ((g142) & (!g296) & (!sk[64]) & (!g316) & (g474) & (g494)) + ((g142) & (!g296) & (!sk[64]) & (g316) & (!g474) & (!g494)) + ((g142) & (!g296) & (!sk[64]) & (g316) & (!g474) & (g494)) + ((g142) & (!g296) & (!sk[64]) & (g316) & (g474) & (!g494)) + ((g142) & (!g296) & (!sk[64]) & (g316) & (g474) & (g494)) + ((g142) & (!g296) & (sk[64]) & (!g316) & (!g474) & (!g494)) + ((g142) & (!g296) & (sk[64]) & (!g316) & (!g474) & (g494)) + ((g142) & (!g296) & (sk[64]) & (g316) & (!g474) & (!g494)) + ((g142) & (!g296) & (sk[64]) & (g316) & (!g474) & (g494)) + ((g142) & (g296) & (!sk[64]) & (!g316) & (!g474) & (!g494)) + ((g142) & (g296) & (!sk[64]) & (!g316) & (!g474) & (g494)) + ((g142) & (g296) & (!sk[64]) & (!g316) & (g474) & (!g494)) + ((g142) & (g296) & (!sk[64]) & (!g316) & (g474) & (g494)) + ((g142) & (g296) & (!sk[64]) & (g316) & (!g474) & (!g494)) + ((g142) & (g296) & (!sk[64]) & (g316) & (!g474) & (g494)) + ((g142) & (g296) & (!sk[64]) & (g316) & (g474) & (!g494)) + ((g142) & (g296) & (!sk[64]) & (g316) & (g474) & (g494)));
	assign g2049 = (((g2041) & (g2042) & (g2043) & (g2044) & (g2047) & (g2048)));
	assign g2050 = (((!g89) & (!g142) & (!g167) & (!sk[66]) & (g187)) + ((!g89) & (!g142) & (!g167) & (sk[66]) & (!g187)) + ((!g89) & (!g142) & (g167) & (!sk[66]) & (!g187)) + ((!g89) & (!g142) & (g167) & (!sk[66]) & (g187)) + ((!g89) & (!g142) & (g167) & (sk[66]) & (!g187)) + ((!g89) & (g142) & (!g167) & (!sk[66]) & (!g187)) + ((!g89) & (g142) & (!g167) & (!sk[66]) & (g187)) + ((!g89) & (g142) & (!g167) & (sk[66]) & (!g187)) + ((!g89) & (g142) & (!g167) & (sk[66]) & (g187)) + ((!g89) & (g142) & (g167) & (!sk[66]) & (!g187)) + ((!g89) & (g142) & (g167) & (!sk[66]) & (g187)) + ((g89) & (!g142) & (!g167) & (!sk[66]) & (g187)) + ((g89) & (!g142) & (g167) & (!sk[66]) & (!g187)) + ((g89) & (!g142) & (g167) & (!sk[66]) & (g187)) + ((g89) & (g142) & (!g167) & (!sk[66]) & (!g187)) + ((g89) & (g142) & (!g167) & (!sk[66]) & (g187)) + ((g89) & (g142) & (g167) & (!sk[66]) & (!g187)) + ((g89) & (g142) & (g167) & (!sk[66]) & (g187)));
	assign g2051 = (((!sk[67]) & (!g142) & (!g318) & (!g341) & (g361)) + ((!sk[67]) & (!g142) & (!g318) & (g341) & (!g361)) + ((!sk[67]) & (!g142) & (!g318) & (g341) & (g361)) + ((!sk[67]) & (!g142) & (g318) & (!g341) & (!g361)) + ((!sk[67]) & (!g142) & (g318) & (!g341) & (g361)) + ((!sk[67]) & (!g142) & (g318) & (g341) & (!g361)) + ((!sk[67]) & (!g142) & (g318) & (g341) & (g361)) + ((!sk[67]) & (g142) & (!g318) & (!g341) & (g361)) + ((!sk[67]) & (g142) & (!g318) & (g341) & (!g361)) + ((!sk[67]) & (g142) & (!g318) & (g341) & (g361)) + ((!sk[67]) & (g142) & (g318) & (!g341) & (!g361)) + ((!sk[67]) & (g142) & (g318) & (!g341) & (g361)) + ((!sk[67]) & (g142) & (g318) & (g341) & (!g361)) + ((!sk[67]) & (g142) & (g318) & (g341) & (g361)) + ((sk[67]) & (!g142) & (!g318) & (!g341) & (!g361)) + ((sk[67]) & (!g142) & (!g318) & (g341) & (!g361)) + ((sk[67]) & (g142) & (!g318) & (!g341) & (!g361)) + ((sk[67]) & (g142) & (!g318) & (!g341) & (g361)));
	assign g2052 = (((!sk[68]) & (!g86) & (!g142) & (!g430) & (g450)) + ((!sk[68]) & (!g86) & (!g142) & (g430) & (!g450)) + ((!sk[68]) & (!g86) & (!g142) & (g430) & (g450)) + ((!sk[68]) & (!g86) & (g142) & (!g430) & (!g450)) + ((!sk[68]) & (!g86) & (g142) & (!g430) & (g450)) + ((!sk[68]) & (!g86) & (g142) & (g430) & (!g450)) + ((!sk[68]) & (!g86) & (g142) & (g430) & (g450)) + ((!sk[68]) & (g86) & (!g142) & (!g430) & (g450)) + ((!sk[68]) & (g86) & (!g142) & (g430) & (!g450)) + ((!sk[68]) & (g86) & (!g142) & (g430) & (g450)) + ((!sk[68]) & (g86) & (g142) & (!g430) & (!g450)) + ((!sk[68]) & (g86) & (g142) & (!g430) & (g450)) + ((!sk[68]) & (g86) & (g142) & (g430) & (!g450)) + ((!sk[68]) & (g86) & (g142) & (g430) & (g450)) + ((sk[68]) & (!g86) & (!g142) & (!g430) & (!g450)) + ((sk[68]) & (!g86) & (!g142) & (g430) & (!g450)) + ((sk[68]) & (!g86) & (g142) & (!g430) & (!g450)) + ((sk[68]) & (!g86) & (g142) & (!g430) & (g450)));
	assign g2053 = (((!g142) & (!g364) & (!sk[69]) & (!g386) & (g406)) + ((!g142) & (!g364) & (!sk[69]) & (g386) & (!g406)) + ((!g142) & (!g364) & (!sk[69]) & (g386) & (g406)) + ((!g142) & (!g364) & (sk[69]) & (!g386) & (!g406)) + ((!g142) & (!g364) & (sk[69]) & (g386) & (!g406)) + ((!g142) & (g364) & (!sk[69]) & (!g386) & (!g406)) + ((!g142) & (g364) & (!sk[69]) & (!g386) & (g406)) + ((!g142) & (g364) & (!sk[69]) & (g386) & (!g406)) + ((!g142) & (g364) & (!sk[69]) & (g386) & (g406)) + ((g142) & (!g364) & (!sk[69]) & (!g386) & (g406)) + ((g142) & (!g364) & (!sk[69]) & (g386) & (!g406)) + ((g142) & (!g364) & (!sk[69]) & (g386) & (g406)) + ((g142) & (!g364) & (sk[69]) & (!g386) & (!g406)) + ((g142) & (!g364) & (sk[69]) & (!g386) & (g406)) + ((g142) & (g364) & (!sk[69]) & (!g386) & (!g406)) + ((g142) & (g364) & (!sk[69]) & (!g386) & (g406)) + ((g142) & (g364) & (!sk[69]) & (g386) & (!g406)) + ((g142) & (g364) & (!sk[69]) & (g386) & (g406)));
	assign g2054 = (((!g2050) & (!g2051) & (!g2052) & (!sk[70]) & (g2053)) + ((!g2050) & (!g2051) & (g2052) & (!sk[70]) & (!g2053)) + ((!g2050) & (!g2051) & (g2052) & (!sk[70]) & (g2053)) + ((!g2050) & (!g2051) & (g2052) & (sk[70]) & (g2053)) + ((!g2050) & (g2051) & (!g2052) & (!sk[70]) & (!g2053)) + ((!g2050) & (g2051) & (!g2052) & (!sk[70]) & (g2053)) + ((!g2050) & (g2051) & (g2052) & (!sk[70]) & (!g2053)) + ((!g2050) & (g2051) & (g2052) & (!sk[70]) & (g2053)) + ((g2050) & (!g2051) & (!g2052) & (!sk[70]) & (g2053)) + ((g2050) & (!g2051) & (g2052) & (!sk[70]) & (!g2053)) + ((g2050) & (!g2051) & (g2052) & (!sk[70]) & (g2053)) + ((g2050) & (g2051) & (!g2052) & (!sk[70]) & (!g2053)) + ((g2050) & (g2051) & (!g2052) & (!sk[70]) & (g2053)) + ((g2050) & (g2051) & (g2052) & (!sk[70]) & (!g2053)) + ((g2050) & (g2051) & (g2052) & (!sk[70]) & (g2053)));
	assign g5021 = (((!g2059) & (!sk[71]) & (!g2925) & (g2055)) + ((!g2059) & (!sk[71]) & (g2925) & (!g2055)) + ((!g2059) & (!sk[71]) & (g2925) & (g2055)) + ((!g2059) & (sk[71]) & (!g2925) & (g2055)) + ((!g2059) & (sk[71]) & (g2925) & (g2055)) + ((g2059) & (!sk[71]) & (!g2925) & (g2055)) + ((g2059) & (!sk[71]) & (g2925) & (!g2055)) + ((g2059) & (!sk[71]) & (g2925) & (g2055)) + ((g2059) & (sk[71]) & (g2925) & (!g2055)) + ((g2059) & (sk[71]) & (g2925) & (g2055)));
	assign g2056 = (((!g2040) & (!g2030) & (!g1632) & (!g2049) & (!g2054) & (g2055)) + ((!g2040) & (!g2030) & (!g1632) & (!g2049) & (g2054) & (g2055)) + ((!g2040) & (!g2030) & (!g1632) & (g2049) & (!g2054) & (g2055)) + ((!g2040) & (!g2030) & (!g1632) & (g2049) & (g2054) & (g2055)) + ((!g2040) & (!g2030) & (g1632) & (!g2049) & (!g2054) & (g2055)) + ((!g2040) & (!g2030) & (g1632) & (!g2049) & (g2054) & (g2055)) + ((!g2040) & (!g2030) & (g1632) & (g2049) & (!g2054) & (g2055)) + ((!g2040) & (!g2030) & (g1632) & (g2049) & (g2054) & (g2055)) + ((g2040) & (!g2030) & (!g1632) & (!g2049) & (!g2054) & (g2055)) + ((g2040) & (!g2030) & (!g1632) & (!g2049) & (g2054) & (g2055)) + ((g2040) & (!g2030) & (!g1632) & (g2049) & (!g2054) & (g2055)) + ((g2040) & (!g2030) & (g1632) & (!g2049) & (!g2054) & (g2055)) + ((g2040) & (!g2030) & (g1632) & (!g2049) & (g2054) & (g2055)) + ((g2040) & (!g2030) & (g1632) & (g2049) & (!g2054) & (g2055)) + ((g2040) & (!g2030) & (g1632) & (g2049) & (g2054) & (!g2055)) + ((g2040) & (!g2030) & (g1632) & (g2049) & (g2054) & (g2055)));
	assign g2057 = (((!sk[73]) & (!g114) & (!g115) & (!nmi_i) & (g2023)) + ((!sk[73]) & (!g114) & (!g115) & (nmi_i) & (!g2023)) + ((!sk[73]) & (!g114) & (!g115) & (nmi_i) & (g2023)) + ((!sk[73]) & (!g114) & (g115) & (!nmi_i) & (!g2023)) + ((!sk[73]) & (!g114) & (g115) & (!nmi_i) & (g2023)) + ((!sk[73]) & (!g114) & (g115) & (nmi_i) & (!g2023)) + ((!sk[73]) & (!g114) & (g115) & (nmi_i) & (g2023)) + ((!sk[73]) & (g114) & (!g115) & (!nmi_i) & (g2023)) + ((!sk[73]) & (g114) & (!g115) & (nmi_i) & (!g2023)) + ((!sk[73]) & (g114) & (!g115) & (nmi_i) & (g2023)) + ((!sk[73]) & (g114) & (g115) & (!nmi_i) & (!g2023)) + ((!sk[73]) & (g114) & (g115) & (!nmi_i) & (g2023)) + ((!sk[73]) & (g114) & (g115) & (nmi_i) & (!g2023)) + ((!sk[73]) & (g114) & (g115) & (nmi_i) & (g2023)) + ((sk[73]) & (!g114) & (!g115) & (!nmi_i) & (!g2023)) + ((sk[73]) & (!g114) & (g115) & (!nmi_i) & (!g2023)) + ((sk[73]) & (g114) & (!g115) & (!nmi_i) & (!g2023)));
	assign g2058 = (((!g123) & (g2037) & (!intr_i) & (!g2039) & (!g2056) & (!g2057)) + ((!g123) & (g2037) & (!intr_i) & (!g2039) & (!g2056) & (g2057)) + ((!g123) & (g2037) & (!intr_i) & (!g2039) & (g2056) & (!g2057)) + ((!g123) & (g2037) & (!intr_i) & (!g2039) & (g2056) & (g2057)) + ((!g123) & (g2037) & (!intr_i) & (g2039) & (!g2056) & (!g2057)) + ((!g123) & (g2037) & (!intr_i) & (g2039) & (!g2056) & (g2057)) + ((!g123) & (g2037) & (!intr_i) & (g2039) & (g2056) & (!g2057)) + ((!g123) & (g2037) & (!intr_i) & (g2039) & (g2056) & (g2057)) + ((!g123) & (g2037) & (intr_i) & (!g2039) & (!g2056) & (!g2057)) + ((!g123) & (g2037) & (intr_i) & (!g2039) & (!g2056) & (g2057)) + ((!g123) & (g2037) & (intr_i) & (!g2039) & (g2056) & (!g2057)) + ((!g123) & (g2037) & (intr_i) & (g2039) & (!g2056) & (!g2057)) + ((!g123) & (g2037) & (intr_i) & (g2039) & (g2056) & (!g2057)));
	assign g2059 = (((!g74) & (!sk[75]) & (!dmem_ack_i) & (g75)) + ((!g74) & (!sk[75]) & (dmem_ack_i) & (!g75)) + ((!g74) & (!sk[75]) & (dmem_ack_i) & (g75)) + ((!g74) & (sk[75]) & (dmem_ack_i) & (g75)) + ((g74) & (!sk[75]) & (!dmem_ack_i) & (g75)) + ((g74) & (!sk[75]) & (dmem_ack_i) & (!g75)) + ((g74) & (!sk[75]) & (dmem_ack_i) & (g75)) + ((g74) & (sk[75]) & (!dmem_ack_i) & (!g75)) + ((g74) & (sk[75]) & (!dmem_ack_i) & (g75)) + ((g74) & (sk[75]) & (dmem_ack_i) & (!g75)) + ((g74) & (sk[75]) & (dmem_ack_i) & (g75)));
	assign g5022 = (((!sk[76]) & (!g2921) & (!g2926) & (g2060)) + ((!sk[76]) & (!g2921) & (g2926) & (!g2060)) + ((!sk[76]) & (!g2921) & (g2926) & (g2060)) + ((!sk[76]) & (g2921) & (!g2926) & (g2060)) + ((!sk[76]) & (g2921) & (g2926) & (!g2060)) + ((!sk[76]) & (g2921) & (g2926) & (g2060)) + ((sk[76]) & (!g2921) & (!g2926) & (g2060)) + ((sk[76]) & (!g2921) & (g2926) & (g2060)) + ((sk[76]) & (g2921) & (g2926) & (!g2060)) + ((sk[76]) & (g2921) & (g2926) & (g2060)));
	assign g2061 = (((!g77) & (!sk[77]) & (!g1604) & (!g2033) & (g2034) & (!g2060)) + ((!g77) & (!sk[77]) & (!g1604) & (!g2033) & (g2034) & (g2060)) + ((!g77) & (!sk[77]) & (!g1604) & (g2033) & (!g2034) & (!g2060)) + ((!g77) & (!sk[77]) & (!g1604) & (g2033) & (!g2034) & (g2060)) + ((!g77) & (!sk[77]) & (!g1604) & (g2033) & (g2034) & (!g2060)) + ((!g77) & (!sk[77]) & (!g1604) & (g2033) & (g2034) & (g2060)) + ((!g77) & (!sk[77]) & (g1604) & (!g2033) & (!g2034) & (!g2060)) + ((!g77) & (!sk[77]) & (g1604) & (!g2033) & (!g2034) & (g2060)) + ((!g77) & (!sk[77]) & (g1604) & (!g2033) & (g2034) & (!g2060)) + ((!g77) & (!sk[77]) & (g1604) & (!g2033) & (g2034) & (g2060)) + ((!g77) & (!sk[77]) & (g1604) & (g2033) & (!g2034) & (!g2060)) + ((!g77) & (!sk[77]) & (g1604) & (g2033) & (!g2034) & (g2060)) + ((!g77) & (!sk[77]) & (g1604) & (g2033) & (g2034) & (!g2060)) + ((!g77) & (!sk[77]) & (g1604) & (g2033) & (g2034) & (g2060)) + ((!g77) & (sk[77]) & (!g1604) & (!g2033) & (!g2034) & (g2060)) + ((!g77) & (sk[77]) & (g1604) & (!g2033) & (!g2034) & (g2060)) + ((!g77) & (sk[77]) & (g1604) & (!g2033) & (g2034) & (!g2060)) + ((!g77) & (sk[77]) & (g1604) & (!g2033) & (g2034) & (g2060)) + ((g77) & (!sk[77]) & (!g1604) & (!g2033) & (g2034) & (!g2060)) + ((g77) & (!sk[77]) & (!g1604) & (!g2033) & (g2034) & (g2060)) + ((g77) & (!sk[77]) & (!g1604) & (g2033) & (!g2034) & (!g2060)) + ((g77) & (!sk[77]) & (!g1604) & (g2033) & (!g2034) & (g2060)) + ((g77) & (!sk[77]) & (!g1604) & (g2033) & (g2034) & (!g2060)) + ((g77) & (!sk[77]) & (!g1604) & (g2033) & (g2034) & (g2060)) + ((g77) & (!sk[77]) & (g1604) & (!g2033) & (!g2034) & (!g2060)) + ((g77) & (!sk[77]) & (g1604) & (!g2033) & (!g2034) & (g2060)) + ((g77) & (!sk[77]) & (g1604) & (!g2033) & (g2034) & (!g2060)) + ((g77) & (!sk[77]) & (g1604) & (!g2033) & (g2034) & (g2060)) + ((g77) & (!sk[77]) & (g1604) & (g2033) & (!g2034) & (!g2060)) + ((g77) & (!sk[77]) & (g1604) & (g2033) & (!g2034) & (g2060)) + ((g77) & (!sk[77]) & (g1604) & (g2033) & (g2034) & (!g2060)) + ((g77) & (!sk[77]) & (g1604) & (g2033) & (g2034) & (g2060)) + ((g77) & (sk[77]) & (!g1604) & (!g2033) & (!g2034) & (g2060)) + ((g77) & (sk[77]) & (!g1604) & (g2033) & (!g2034) & (!g2060)) + ((g77) & (sk[77]) & (!g1604) & (g2033) & (!g2034) & (g2060)) + ((g77) & (sk[77]) & (g1604) & (!g2033) & (!g2034) & (g2060)) + ((g77) & (sk[77]) & (g1604) & (!g2033) & (g2034) & (!g2060)) + ((g77) & (sk[77]) & (g1604) & (!g2033) & (g2034) & (g2060)) + ((g77) & (sk[77]) & (g1604) & (g2033) & (!g2034) & (!g2060)) + ((g77) & (sk[77]) & (g1604) & (g2033) & (!g2034) & (g2060)));
	assign g2062 = (((!g2022) & (!g77) & (!nmi_i) & (!g2023) & (!g2029) & (g2061)) + ((!g2022) & (!g77) & (!nmi_i) & (g2023) & (!g2029) & (g2061)) + ((!g2022) & (!g77) & (nmi_i) & (!g2023) & (!g2029) & (g2061)) + ((!g2022) & (!g77) & (nmi_i) & (g2023) & (!g2029) & (g2061)) + ((!g2022) & (g77) & (!nmi_i) & (!g2023) & (!g2029) & (g2061)) + ((!g2022) & (g77) & (!nmi_i) & (!g2023) & (g2029) & (!g2061)) + ((!g2022) & (g77) & (!nmi_i) & (!g2023) & (g2029) & (g2061)) + ((!g2022) & (g77) & (!nmi_i) & (g2023) & (!g2029) & (g2061)) + ((!g2022) & (g77) & (!nmi_i) & (g2023) & (g2029) & (!g2061)) + ((!g2022) & (g77) & (!nmi_i) & (g2023) & (g2029) & (g2061)) + ((!g2022) & (g77) & (nmi_i) & (!g2023) & (!g2029) & (g2061)) + ((!g2022) & (g77) & (nmi_i) & (!g2023) & (g2029) & (!g2061)) + ((!g2022) & (g77) & (nmi_i) & (!g2023) & (g2029) & (g2061)) + ((!g2022) & (g77) & (nmi_i) & (g2023) & (!g2029) & (g2061)) + ((!g2022) & (g77) & (nmi_i) & (g2023) & (g2029) & (!g2061)) + ((!g2022) & (g77) & (nmi_i) & (g2023) & (g2029) & (g2061)) + ((g2022) & (!g77) & (!nmi_i) & (!g2023) & (!g2029) & (g2061)) + ((g2022) & (g77) & (!nmi_i) & (!g2023) & (!g2029) & (g2061)) + ((g2022) & (g77) & (!nmi_i) & (!g2023) & (g2029) & (!g2061)) + ((g2022) & (g77) & (!nmi_i) & (!g2023) & (g2029) & (g2061)));
	assign g2063 = (((!g123) & (!intr_i) & (!g2039) & (!g2056) & (!g2057) & (g2062)) + ((!g123) & (!intr_i) & (!g2039) & (!g2056) & (g2057) & (g2062)) + ((!g123) & (!intr_i) & (!g2039) & (g2056) & (!g2057) & (g2062)) + ((!g123) & (!intr_i) & (!g2039) & (g2056) & (g2057) & (g2062)) + ((!g123) & (!intr_i) & (g2039) & (!g2056) & (!g2057) & (g2062)) + ((!g123) & (!intr_i) & (g2039) & (!g2056) & (g2057) & (g2062)) + ((!g123) & (!intr_i) & (g2039) & (g2056) & (!g2057) & (g2062)) + ((!g123) & (!intr_i) & (g2039) & (g2056) & (g2057) & (g2062)) + ((!g123) & (intr_i) & (!g2039) & (!g2056) & (!g2057) & (g2062)) + ((!g123) & (intr_i) & (!g2039) & (!g2056) & (g2057) & (g2062)) + ((!g123) & (intr_i) & (!g2039) & (g2056) & (!g2057) & (g2062)) + ((!g123) & (intr_i) & (g2039) & (!g2056) & (!g2057) & (g2062)) + ((!g123) & (intr_i) & (g2039) & (g2056) & (!g2057) & (g2062)));
	assign g2064 = (((dmem_ack_i) & (!sk[80]) & (!g129)) + ((dmem_ack_i) & (!sk[80]) & (g129)) + ((dmem_ack_i) & (sk[80]) & (g129)));
	assign g2065 = (((!sk[81]) & (!dmem_ack_i) & (!g129) & (g2019)) + ((!sk[81]) & (!dmem_ack_i) & (g129) & (!g2019)) + ((!sk[81]) & (!dmem_ack_i) & (g129) & (g2019)) + ((!sk[81]) & (dmem_ack_i) & (!g129) & (g2019)) + ((!sk[81]) & (dmem_ack_i) & (g129) & (!g2019)) + ((!sk[81]) & (dmem_ack_i) & (g129) & (g2019)) + ((sk[81]) & (!dmem_ack_i) & (!g129) & (g2019)) + ((sk[81]) & (!dmem_ack_i) & (g129) & (!g2019)) + ((sk[81]) & (!dmem_ack_i) & (g129) & (g2019)) + ((sk[81]) & (dmem_ack_i) & (!g129) & (g2019)) + ((sk[81]) & (dmem_ack_i) & (g129) & (g2019)));
	assign g5023 = (((!g2921) & (!g2927) & (!sk[82]) & (g2066)) + ((!g2921) & (!g2927) & (sk[82]) & (g2066)) + ((!g2921) & (g2927) & (!sk[82]) & (!g2066)) + ((!g2921) & (g2927) & (!sk[82]) & (g2066)) + ((!g2921) & (g2927) & (sk[82]) & (g2066)) + ((g2921) & (!g2927) & (!sk[82]) & (g2066)) + ((g2921) & (g2927) & (!sk[82]) & (!g2066)) + ((g2921) & (g2927) & (!sk[82]) & (g2066)) + ((g2921) & (g2927) & (sk[82]) & (!g2066)) + ((g2921) & (g2927) & (sk[82]) & (g2066)));
	assign g2067 = (((!g89) & (!g1632) & (!g2033) & (!g2034) & (!g141) & (g2066)) + ((!g89) & (!g1632) & (!g2033) & (!g2034) & (g141) & (g2066)) + ((!g89) & (!g1632) & (g2033) & (!g2034) & (g141) & (!g2066)) + ((!g89) & (!g1632) & (g2033) & (!g2034) & (g141) & (g2066)) + ((!g89) & (g1632) & (!g2033) & (!g2034) & (!g141) & (g2066)) + ((!g89) & (g1632) & (!g2033) & (!g2034) & (g141) & (g2066)) + ((!g89) & (g1632) & (!g2033) & (g2034) & (!g141) & (!g2066)) + ((!g89) & (g1632) & (!g2033) & (g2034) & (!g141) & (g2066)) + ((!g89) & (g1632) & (!g2033) & (g2034) & (g141) & (!g2066)) + ((!g89) & (g1632) & (!g2033) & (g2034) & (g141) & (g2066)) + ((!g89) & (g1632) & (g2033) & (!g2034) & (g141) & (!g2066)) + ((!g89) & (g1632) & (g2033) & (!g2034) & (g141) & (g2066)) + ((g89) & (!g1632) & (!g2033) & (!g2034) & (!g141) & (g2066)) + ((g89) & (!g1632) & (!g2033) & (!g2034) & (g141) & (g2066)) + ((g89) & (!g1632) & (g2033) & (!g2034) & (!g141) & (!g2066)) + ((g89) & (!g1632) & (g2033) & (!g2034) & (!g141) & (g2066)) + ((g89) & (g1632) & (!g2033) & (!g2034) & (!g141) & (g2066)) + ((g89) & (g1632) & (!g2033) & (!g2034) & (g141) & (g2066)) + ((g89) & (g1632) & (!g2033) & (g2034) & (!g141) & (!g2066)) + ((g89) & (g1632) & (!g2033) & (g2034) & (!g141) & (g2066)) + ((g89) & (g1632) & (!g2033) & (g2034) & (g141) & (!g2066)) + ((g89) & (g1632) & (!g2033) & (g2034) & (g141) & (g2066)) + ((g89) & (g1632) & (g2033) & (!g2034) & (!g141) & (!g2066)) + ((g89) & (g1632) & (g2033) & (!g2034) & (!g141) & (g2066)));
	assign g2068 = (((!g2022) & (!nmi_i) & (!g2023) & (!g2029) & (!g141) & (g2067)) + ((!g2022) & (!nmi_i) & (!g2023) & (!g2029) & (g141) & (g2067)) + ((!g2022) & (!nmi_i) & (!g2023) & (g2029) & (!g141) & (!g2067)) + ((!g2022) & (!nmi_i) & (!g2023) & (g2029) & (!g141) & (g2067)) + ((!g2022) & (!nmi_i) & (g2023) & (!g2029) & (!g141) & (g2067)) + ((!g2022) & (!nmi_i) & (g2023) & (!g2029) & (g141) & (g2067)) + ((!g2022) & (!nmi_i) & (g2023) & (g2029) & (!g141) & (!g2067)) + ((!g2022) & (!nmi_i) & (g2023) & (g2029) & (!g141) & (g2067)) + ((!g2022) & (nmi_i) & (!g2023) & (!g2029) & (!g141) & (g2067)) + ((!g2022) & (nmi_i) & (!g2023) & (!g2029) & (g141) & (g2067)) + ((!g2022) & (nmi_i) & (!g2023) & (g2029) & (!g141) & (!g2067)) + ((!g2022) & (nmi_i) & (!g2023) & (g2029) & (!g141) & (g2067)) + ((!g2022) & (nmi_i) & (g2023) & (!g2029) & (!g141) & (g2067)) + ((!g2022) & (nmi_i) & (g2023) & (!g2029) & (g141) & (g2067)) + ((!g2022) & (nmi_i) & (g2023) & (g2029) & (!g141) & (!g2067)) + ((!g2022) & (nmi_i) & (g2023) & (g2029) & (!g141) & (g2067)) + ((g2022) & (!nmi_i) & (!g2023) & (!g2029) & (!g141) & (g2067)) + ((g2022) & (!nmi_i) & (!g2023) & (!g2029) & (g141) & (g2067)) + ((g2022) & (!nmi_i) & (!g2023) & (g2029) & (!g141) & (!g2067)) + ((g2022) & (!nmi_i) & (!g2023) & (g2029) & (!g141) & (g2067)));
	assign g2069 = (((!g123) & (!intr_i) & (!g2039) & (!g2056) & (!g2057) & (g2068)) + ((!g123) & (!intr_i) & (!g2039) & (!g2056) & (g2057) & (g2068)) + ((!g123) & (!intr_i) & (!g2039) & (g2056) & (!g2057) & (g2068)) + ((!g123) & (!intr_i) & (!g2039) & (g2056) & (g2057) & (g2068)) + ((!g123) & (!intr_i) & (g2039) & (!g2056) & (!g2057) & (g2068)) + ((!g123) & (!intr_i) & (g2039) & (!g2056) & (g2057) & (g2068)) + ((!g123) & (!intr_i) & (g2039) & (g2056) & (!g2057) & (g2068)) + ((!g123) & (!intr_i) & (g2039) & (g2056) & (g2057) & (g2068)) + ((!g123) & (intr_i) & (!g2039) & (!g2056) & (!g2057) & (g2068)) + ((!g123) & (intr_i) & (!g2039) & (!g2056) & (g2057) & (g2068)) + ((!g123) & (intr_i) & (!g2039) & (g2056) & (!g2057) & (g2068)) + ((!g123) & (intr_i) & (g2039) & (!g2056) & (!g2057) & (g2068)) + ((!g123) & (intr_i) & (g2039) & (g2056) & (!g2057) & (g2068)));
	assign g2072 = (((!sk[86]) & (g2071) & (!g2070)) + ((!sk[86]) & (g2071) & (g2070)) + ((sk[86]) & (!g2071) & (g2070)) + ((sk[86]) & (g2071) & (!g2070)));
	assign g2075 = (((!sk[87]) & (!g2074) & (!g2071) & (g2070)) + ((!sk[87]) & (!g2074) & (g2071) & (!g2070)) + ((!sk[87]) & (!g2074) & (g2071) & (g2070)) + ((!sk[87]) & (g2074) & (!g2071) & (g2070)) + ((!sk[87]) & (g2074) & (g2071) & (!g2070)) + ((!sk[87]) & (g2074) & (g2071) & (g2070)) + ((sk[87]) & (!g2074) & (!g2071) & (g2070)));
	assign g2078 = (((!g2075) & (!g2076) & (!sk[88]) & (g2077)) + ((!g2075) & (g2076) & (!sk[88]) & (!g2077)) + ((!g2075) & (g2076) & (!sk[88]) & (g2077)) + ((g2075) & (!g2076) & (!sk[88]) & (g2077)) + ((g2075) & (!g2076) & (sk[88]) & (!g2077)) + ((g2075) & (g2076) & (!sk[88]) & (!g2077)) + ((g2075) & (g2076) & (!sk[88]) & (g2077)));
	assign g5024 = (((!sk[89]) & (!g2059) & (!g2973) & (g2079)) + ((!sk[89]) & (!g2059) & (g2973) & (!g2079)) + ((!sk[89]) & (!g2059) & (g2973) & (g2079)) + ((!sk[89]) & (g2059) & (!g2973) & (g2079)) + ((!sk[89]) & (g2059) & (g2973) & (!g2079)) + ((!sk[89]) & (g2059) & (g2973) & (g2079)) + ((sk[89]) & (!g2059) & (!g2973) & (g2079)) + ((sk[89]) & (!g2059) & (g2973) & (g2079)) + ((sk[89]) & (g2059) & (g2973) & (!g2079)) + ((sk[89]) & (g2059) & (g2973) & (g2079)));
	assign g2082 = (((!g2071) & (!g2070) & (!sk[90]) & (!g2080) & (g2081)) + ((!g2071) & (!g2070) & (!sk[90]) & (g2080) & (!g2081)) + ((!g2071) & (!g2070) & (!sk[90]) & (g2080) & (g2081)) + ((!g2071) & (!g2070) & (sk[90]) & (!g2080) & (!g2081)) + ((!g2071) & (!g2070) & (sk[90]) & (!g2080) & (g2081)) + ((!g2071) & (!g2070) & (sk[90]) & (g2080) & (!g2081)) + ((!g2071) & (!g2070) & (sk[90]) & (g2080) & (g2081)) + ((!g2071) & (g2070) & (!sk[90]) & (!g2080) & (!g2081)) + ((!g2071) & (g2070) & (!sk[90]) & (!g2080) & (g2081)) + ((!g2071) & (g2070) & (!sk[90]) & (g2080) & (!g2081)) + ((!g2071) & (g2070) & (!sk[90]) & (g2080) & (g2081)) + ((g2071) & (!g2070) & (!sk[90]) & (!g2080) & (g2081)) + ((g2071) & (!g2070) & (!sk[90]) & (g2080) & (!g2081)) + ((g2071) & (!g2070) & (!sk[90]) & (g2080) & (g2081)) + ((g2071) & (!g2070) & (sk[90]) & (g2080) & (!g2081)) + ((g2071) & (!g2070) & (sk[90]) & (g2080) & (g2081)) + ((g2071) & (g2070) & (!sk[90]) & (!g2080) & (!g2081)) + ((g2071) & (g2070) & (!sk[90]) & (!g2080) & (g2081)) + ((g2071) & (g2070) & (!sk[90]) & (g2080) & (!g2081)) + ((g2071) & (g2070) & (!sk[90]) & (g2080) & (g2081)) + ((g2071) & (g2070) & (sk[90]) & (!g2080) & (g2081)));
	assign g2087 = (((!g2083) & (!g2084) & (!g2085) & (g2086) & (g2071) & (g2074)) + ((!g2083) & (!g2084) & (g2085) & (!g2086) & (!g2071) & (g2074)) + ((!g2083) & (!g2084) & (g2085) & (g2086) & (!g2071) & (g2074)) + ((!g2083) & (!g2084) & (g2085) & (g2086) & (g2071) & (g2074)) + ((!g2083) & (g2084) & (!g2085) & (!g2086) & (g2071) & (!g2074)) + ((!g2083) & (g2084) & (!g2085) & (g2086) & (g2071) & (!g2074)) + ((!g2083) & (g2084) & (!g2085) & (g2086) & (g2071) & (g2074)) + ((!g2083) & (g2084) & (g2085) & (!g2086) & (!g2071) & (g2074)) + ((!g2083) & (g2084) & (g2085) & (!g2086) & (g2071) & (!g2074)) + ((!g2083) & (g2084) & (g2085) & (g2086) & (!g2071) & (g2074)) + ((!g2083) & (g2084) & (g2085) & (g2086) & (g2071) & (!g2074)) + ((!g2083) & (g2084) & (g2085) & (g2086) & (g2071) & (g2074)) + ((g2083) & (!g2084) & (!g2085) & (!g2086) & (!g2071) & (!g2074)) + ((g2083) & (!g2084) & (!g2085) & (g2086) & (!g2071) & (!g2074)) + ((g2083) & (!g2084) & (!g2085) & (g2086) & (g2071) & (g2074)) + ((g2083) & (!g2084) & (g2085) & (!g2086) & (!g2071) & (!g2074)) + ((g2083) & (!g2084) & (g2085) & (!g2086) & (!g2071) & (g2074)) + ((g2083) & (!g2084) & (g2085) & (g2086) & (!g2071) & (!g2074)) + ((g2083) & (!g2084) & (g2085) & (g2086) & (!g2071) & (g2074)) + ((g2083) & (!g2084) & (g2085) & (g2086) & (g2071) & (g2074)) + ((g2083) & (g2084) & (!g2085) & (!g2086) & (!g2071) & (!g2074)) + ((g2083) & (g2084) & (!g2085) & (!g2086) & (g2071) & (!g2074)) + ((g2083) & (g2084) & (!g2085) & (g2086) & (!g2071) & (!g2074)) + ((g2083) & (g2084) & (!g2085) & (g2086) & (g2071) & (!g2074)) + ((g2083) & (g2084) & (!g2085) & (g2086) & (g2071) & (g2074)) + ((g2083) & (g2084) & (g2085) & (!g2086) & (!g2071) & (!g2074)) + ((g2083) & (g2084) & (g2085) & (!g2086) & (!g2071) & (g2074)) + ((g2083) & (g2084) & (g2085) & (!g2086) & (g2071) & (!g2074)) + ((g2083) & (g2084) & (g2085) & (g2086) & (!g2071) & (!g2074)) + ((g2083) & (g2084) & (g2085) & (g2086) & (!g2071) & (g2074)) + ((g2083) & (g2084) & (g2085) & (g2086) & (g2071) & (!g2074)) + ((g2083) & (g2084) & (g2085) & (g2086) & (g2071) & (g2074)));
	assign g2092 = (((!g2088) & (!g2089) & (!g2090) & (g2091) & (g2071) & (g2074)) + ((!g2088) & (!g2089) & (g2090) & (!g2091) & (!g2071) & (g2074)) + ((!g2088) & (!g2089) & (g2090) & (g2091) & (!g2071) & (g2074)) + ((!g2088) & (!g2089) & (g2090) & (g2091) & (g2071) & (g2074)) + ((!g2088) & (g2089) & (!g2090) & (!g2091) & (g2071) & (!g2074)) + ((!g2088) & (g2089) & (!g2090) & (g2091) & (g2071) & (!g2074)) + ((!g2088) & (g2089) & (!g2090) & (g2091) & (g2071) & (g2074)) + ((!g2088) & (g2089) & (g2090) & (!g2091) & (!g2071) & (g2074)) + ((!g2088) & (g2089) & (g2090) & (!g2091) & (g2071) & (!g2074)) + ((!g2088) & (g2089) & (g2090) & (g2091) & (!g2071) & (g2074)) + ((!g2088) & (g2089) & (g2090) & (g2091) & (g2071) & (!g2074)) + ((!g2088) & (g2089) & (g2090) & (g2091) & (g2071) & (g2074)) + ((g2088) & (!g2089) & (!g2090) & (!g2091) & (!g2071) & (!g2074)) + ((g2088) & (!g2089) & (!g2090) & (g2091) & (!g2071) & (!g2074)) + ((g2088) & (!g2089) & (!g2090) & (g2091) & (g2071) & (g2074)) + ((g2088) & (!g2089) & (g2090) & (!g2091) & (!g2071) & (!g2074)) + ((g2088) & (!g2089) & (g2090) & (!g2091) & (!g2071) & (g2074)) + ((g2088) & (!g2089) & (g2090) & (g2091) & (!g2071) & (!g2074)) + ((g2088) & (!g2089) & (g2090) & (g2091) & (!g2071) & (g2074)) + ((g2088) & (!g2089) & (g2090) & (g2091) & (g2071) & (g2074)) + ((g2088) & (g2089) & (!g2090) & (!g2091) & (!g2071) & (!g2074)) + ((g2088) & (g2089) & (!g2090) & (!g2091) & (g2071) & (!g2074)) + ((g2088) & (g2089) & (!g2090) & (g2091) & (!g2071) & (!g2074)) + ((g2088) & (g2089) & (!g2090) & (g2091) & (g2071) & (!g2074)) + ((g2088) & (g2089) & (!g2090) & (g2091) & (g2071) & (g2074)) + ((g2088) & (g2089) & (g2090) & (!g2091) & (!g2071) & (!g2074)) + ((g2088) & (g2089) & (g2090) & (!g2091) & (!g2071) & (g2074)) + ((g2088) & (g2089) & (g2090) & (!g2091) & (g2071) & (!g2074)) + ((g2088) & (g2089) & (g2090) & (g2091) & (!g2071) & (!g2074)) + ((g2088) & (g2089) & (g2090) & (g2091) & (!g2071) & (g2074)) + ((g2088) & (g2089) & (g2090) & (g2091) & (g2071) & (!g2074)) + ((g2088) & (g2089) & (g2090) & (g2091) & (g2071) & (g2074)));
	assign g2097 = (((!g2093) & (!g2094) & (!g2095) & (g2096) & (g2071) & (g2074)) + ((!g2093) & (!g2094) & (g2095) & (!g2096) & (!g2071) & (g2074)) + ((!g2093) & (!g2094) & (g2095) & (g2096) & (!g2071) & (g2074)) + ((!g2093) & (!g2094) & (g2095) & (g2096) & (g2071) & (g2074)) + ((!g2093) & (g2094) & (!g2095) & (!g2096) & (g2071) & (!g2074)) + ((!g2093) & (g2094) & (!g2095) & (g2096) & (g2071) & (!g2074)) + ((!g2093) & (g2094) & (!g2095) & (g2096) & (g2071) & (g2074)) + ((!g2093) & (g2094) & (g2095) & (!g2096) & (!g2071) & (g2074)) + ((!g2093) & (g2094) & (g2095) & (!g2096) & (g2071) & (!g2074)) + ((!g2093) & (g2094) & (g2095) & (g2096) & (!g2071) & (g2074)) + ((!g2093) & (g2094) & (g2095) & (g2096) & (g2071) & (!g2074)) + ((!g2093) & (g2094) & (g2095) & (g2096) & (g2071) & (g2074)) + ((g2093) & (!g2094) & (!g2095) & (!g2096) & (!g2071) & (!g2074)) + ((g2093) & (!g2094) & (!g2095) & (g2096) & (!g2071) & (!g2074)) + ((g2093) & (!g2094) & (!g2095) & (g2096) & (g2071) & (g2074)) + ((g2093) & (!g2094) & (g2095) & (!g2096) & (!g2071) & (!g2074)) + ((g2093) & (!g2094) & (g2095) & (!g2096) & (!g2071) & (g2074)) + ((g2093) & (!g2094) & (g2095) & (g2096) & (!g2071) & (!g2074)) + ((g2093) & (!g2094) & (g2095) & (g2096) & (!g2071) & (g2074)) + ((g2093) & (!g2094) & (g2095) & (g2096) & (g2071) & (g2074)) + ((g2093) & (g2094) & (!g2095) & (!g2096) & (!g2071) & (!g2074)) + ((g2093) & (g2094) & (!g2095) & (!g2096) & (g2071) & (!g2074)) + ((g2093) & (g2094) & (!g2095) & (g2096) & (!g2071) & (!g2074)) + ((g2093) & (g2094) & (!g2095) & (g2096) & (g2071) & (!g2074)) + ((g2093) & (g2094) & (!g2095) & (g2096) & (g2071) & (g2074)) + ((g2093) & (g2094) & (g2095) & (!g2096) & (!g2071) & (!g2074)) + ((g2093) & (g2094) & (g2095) & (!g2096) & (!g2071) & (g2074)) + ((g2093) & (g2094) & (g2095) & (!g2096) & (g2071) & (!g2074)) + ((g2093) & (g2094) & (g2095) & (g2096) & (!g2071) & (!g2074)) + ((g2093) & (g2094) & (g2095) & (g2096) & (!g2071) & (g2074)) + ((g2093) & (g2094) & (g2095) & (g2096) & (g2071) & (!g2074)) + ((g2093) & (g2094) & (g2095) & (g2096) & (g2071) & (g2074)));
	assign g2102 = (((!g2098) & (!g2099) & (!g2100) & (g2101) & (g2071) & (g2074)) + ((!g2098) & (!g2099) & (g2100) & (!g2101) & (!g2071) & (g2074)) + ((!g2098) & (!g2099) & (g2100) & (g2101) & (!g2071) & (g2074)) + ((!g2098) & (!g2099) & (g2100) & (g2101) & (g2071) & (g2074)) + ((!g2098) & (g2099) & (!g2100) & (!g2101) & (g2071) & (!g2074)) + ((!g2098) & (g2099) & (!g2100) & (g2101) & (g2071) & (!g2074)) + ((!g2098) & (g2099) & (!g2100) & (g2101) & (g2071) & (g2074)) + ((!g2098) & (g2099) & (g2100) & (!g2101) & (!g2071) & (g2074)) + ((!g2098) & (g2099) & (g2100) & (!g2101) & (g2071) & (!g2074)) + ((!g2098) & (g2099) & (g2100) & (g2101) & (!g2071) & (g2074)) + ((!g2098) & (g2099) & (g2100) & (g2101) & (g2071) & (!g2074)) + ((!g2098) & (g2099) & (g2100) & (g2101) & (g2071) & (g2074)) + ((g2098) & (!g2099) & (!g2100) & (!g2101) & (!g2071) & (!g2074)) + ((g2098) & (!g2099) & (!g2100) & (g2101) & (!g2071) & (!g2074)) + ((g2098) & (!g2099) & (!g2100) & (g2101) & (g2071) & (g2074)) + ((g2098) & (!g2099) & (g2100) & (!g2101) & (!g2071) & (!g2074)) + ((g2098) & (!g2099) & (g2100) & (!g2101) & (!g2071) & (g2074)) + ((g2098) & (!g2099) & (g2100) & (g2101) & (!g2071) & (!g2074)) + ((g2098) & (!g2099) & (g2100) & (g2101) & (!g2071) & (g2074)) + ((g2098) & (!g2099) & (g2100) & (g2101) & (g2071) & (g2074)) + ((g2098) & (g2099) & (!g2100) & (!g2101) & (!g2071) & (!g2074)) + ((g2098) & (g2099) & (!g2100) & (!g2101) & (g2071) & (!g2074)) + ((g2098) & (g2099) & (!g2100) & (g2101) & (!g2071) & (!g2074)) + ((g2098) & (g2099) & (!g2100) & (g2101) & (g2071) & (!g2074)) + ((g2098) & (g2099) & (!g2100) & (g2101) & (g2071) & (g2074)) + ((g2098) & (g2099) & (g2100) & (!g2101) & (!g2071) & (!g2074)) + ((g2098) & (g2099) & (g2100) & (!g2101) & (!g2071) & (g2074)) + ((g2098) & (g2099) & (g2100) & (!g2101) & (g2071) & (!g2074)) + ((g2098) & (g2099) & (g2100) & (g2101) & (!g2071) & (!g2074)) + ((g2098) & (g2099) & (g2100) & (g2101) & (!g2071) & (g2074)) + ((g2098) & (g2099) & (g2100) & (g2101) & (g2071) & (!g2074)) + ((g2098) & (g2099) & (g2100) & (g2101) & (g2071) & (g2074)));
	assign g2103 = (((!g2087) & (!g2092) & (!g2097) & (g2102) & (g2076) & (g2077)) + ((!g2087) & (!g2092) & (g2097) & (!g2102) & (!g2076) & (g2077)) + ((!g2087) & (!g2092) & (g2097) & (g2102) & (!g2076) & (g2077)) + ((!g2087) & (!g2092) & (g2097) & (g2102) & (g2076) & (g2077)) + ((!g2087) & (g2092) & (!g2097) & (!g2102) & (g2076) & (!g2077)) + ((!g2087) & (g2092) & (!g2097) & (g2102) & (g2076) & (!g2077)) + ((!g2087) & (g2092) & (!g2097) & (g2102) & (g2076) & (g2077)) + ((!g2087) & (g2092) & (g2097) & (!g2102) & (!g2076) & (g2077)) + ((!g2087) & (g2092) & (g2097) & (!g2102) & (g2076) & (!g2077)) + ((!g2087) & (g2092) & (g2097) & (g2102) & (!g2076) & (g2077)) + ((!g2087) & (g2092) & (g2097) & (g2102) & (g2076) & (!g2077)) + ((!g2087) & (g2092) & (g2097) & (g2102) & (g2076) & (g2077)) + ((g2087) & (!g2092) & (!g2097) & (!g2102) & (!g2076) & (!g2077)) + ((g2087) & (!g2092) & (!g2097) & (g2102) & (!g2076) & (!g2077)) + ((g2087) & (!g2092) & (!g2097) & (g2102) & (g2076) & (g2077)) + ((g2087) & (!g2092) & (g2097) & (!g2102) & (!g2076) & (!g2077)) + ((g2087) & (!g2092) & (g2097) & (!g2102) & (!g2076) & (g2077)) + ((g2087) & (!g2092) & (g2097) & (g2102) & (!g2076) & (!g2077)) + ((g2087) & (!g2092) & (g2097) & (g2102) & (!g2076) & (g2077)) + ((g2087) & (!g2092) & (g2097) & (g2102) & (g2076) & (g2077)) + ((g2087) & (g2092) & (!g2097) & (!g2102) & (!g2076) & (!g2077)) + ((g2087) & (g2092) & (!g2097) & (!g2102) & (g2076) & (!g2077)) + ((g2087) & (g2092) & (!g2097) & (g2102) & (!g2076) & (!g2077)) + ((g2087) & (g2092) & (!g2097) & (g2102) & (g2076) & (!g2077)) + ((g2087) & (g2092) & (!g2097) & (g2102) & (g2076) & (g2077)) + ((g2087) & (g2092) & (g2097) & (!g2102) & (!g2076) & (!g2077)) + ((g2087) & (g2092) & (g2097) & (!g2102) & (!g2076) & (g2077)) + ((g2087) & (g2092) & (g2097) & (!g2102) & (g2076) & (!g2077)) + ((g2087) & (g2092) & (g2097) & (g2102) & (!g2076) & (!g2077)) + ((g2087) & (g2092) & (g2097) & (g2102) & (!g2076) & (g2077)) + ((g2087) & (g2092) & (g2097) & (g2102) & (g2076) & (!g2077)) + ((g2087) & (g2092) & (g2097) & (g2102) & (g2076) & (g2077)));
	assign g2107 = (((!g2070) & (!g2104) & (!g2105) & (g2106) & (g2071) & (g2074)) + ((!g2070) & (!g2104) & (g2105) & (!g2106) & (!g2071) & (g2074)) + ((!g2070) & (!g2104) & (g2105) & (g2106) & (!g2071) & (g2074)) + ((!g2070) & (!g2104) & (g2105) & (g2106) & (g2071) & (g2074)) + ((!g2070) & (g2104) & (!g2105) & (!g2106) & (g2071) & (!g2074)) + ((!g2070) & (g2104) & (!g2105) & (g2106) & (g2071) & (!g2074)) + ((!g2070) & (g2104) & (!g2105) & (g2106) & (g2071) & (g2074)) + ((!g2070) & (g2104) & (g2105) & (!g2106) & (!g2071) & (g2074)) + ((!g2070) & (g2104) & (g2105) & (!g2106) & (g2071) & (!g2074)) + ((!g2070) & (g2104) & (g2105) & (g2106) & (!g2071) & (g2074)) + ((!g2070) & (g2104) & (g2105) & (g2106) & (g2071) & (!g2074)) + ((!g2070) & (g2104) & (g2105) & (g2106) & (g2071) & (g2074)) + ((g2070) & (!g2104) & (!g2105) & (!g2106) & (!g2071) & (!g2074)) + ((g2070) & (!g2104) & (!g2105) & (g2106) & (!g2071) & (!g2074)) + ((g2070) & (!g2104) & (!g2105) & (g2106) & (g2071) & (g2074)) + ((g2070) & (!g2104) & (g2105) & (!g2106) & (!g2071) & (!g2074)) + ((g2070) & (!g2104) & (g2105) & (!g2106) & (!g2071) & (g2074)) + ((g2070) & (!g2104) & (g2105) & (g2106) & (!g2071) & (!g2074)) + ((g2070) & (!g2104) & (g2105) & (g2106) & (!g2071) & (g2074)) + ((g2070) & (!g2104) & (g2105) & (g2106) & (g2071) & (g2074)) + ((g2070) & (g2104) & (!g2105) & (!g2106) & (!g2071) & (!g2074)) + ((g2070) & (g2104) & (!g2105) & (!g2106) & (g2071) & (!g2074)) + ((g2070) & (g2104) & (!g2105) & (g2106) & (!g2071) & (!g2074)) + ((g2070) & (g2104) & (!g2105) & (g2106) & (g2071) & (!g2074)) + ((g2070) & (g2104) & (!g2105) & (g2106) & (g2071) & (g2074)) + ((g2070) & (g2104) & (g2105) & (!g2106) & (!g2071) & (!g2074)) + ((g2070) & (g2104) & (g2105) & (!g2106) & (!g2071) & (g2074)) + ((g2070) & (g2104) & (g2105) & (!g2106) & (g2071) & (!g2074)) + ((g2070) & (g2104) & (g2105) & (g2106) & (!g2071) & (!g2074)) + ((g2070) & (g2104) & (g2105) & (g2106) & (!g2071) & (g2074)) + ((g2070) & (g2104) & (g2105) & (g2106) & (g2071) & (!g2074)) + ((g2070) & (g2104) & (g2105) & (g2106) & (g2071) & (g2074)));
	assign g2112 = (((!g2108) & (!g2109) & (!g2110) & (g2111) & (g2071) & (g2074)) + ((!g2108) & (!g2109) & (g2110) & (!g2111) & (!g2071) & (g2074)) + ((!g2108) & (!g2109) & (g2110) & (g2111) & (!g2071) & (g2074)) + ((!g2108) & (!g2109) & (g2110) & (g2111) & (g2071) & (g2074)) + ((!g2108) & (g2109) & (!g2110) & (!g2111) & (g2071) & (!g2074)) + ((!g2108) & (g2109) & (!g2110) & (g2111) & (g2071) & (!g2074)) + ((!g2108) & (g2109) & (!g2110) & (g2111) & (g2071) & (g2074)) + ((!g2108) & (g2109) & (g2110) & (!g2111) & (!g2071) & (g2074)) + ((!g2108) & (g2109) & (g2110) & (!g2111) & (g2071) & (!g2074)) + ((!g2108) & (g2109) & (g2110) & (g2111) & (!g2071) & (g2074)) + ((!g2108) & (g2109) & (g2110) & (g2111) & (g2071) & (!g2074)) + ((!g2108) & (g2109) & (g2110) & (g2111) & (g2071) & (g2074)) + ((g2108) & (!g2109) & (!g2110) & (!g2111) & (!g2071) & (!g2074)) + ((g2108) & (!g2109) & (!g2110) & (g2111) & (!g2071) & (!g2074)) + ((g2108) & (!g2109) & (!g2110) & (g2111) & (g2071) & (g2074)) + ((g2108) & (!g2109) & (g2110) & (!g2111) & (!g2071) & (!g2074)) + ((g2108) & (!g2109) & (g2110) & (!g2111) & (!g2071) & (g2074)) + ((g2108) & (!g2109) & (g2110) & (g2111) & (!g2071) & (!g2074)) + ((g2108) & (!g2109) & (g2110) & (g2111) & (!g2071) & (g2074)) + ((g2108) & (!g2109) & (g2110) & (g2111) & (g2071) & (g2074)) + ((g2108) & (g2109) & (!g2110) & (!g2111) & (!g2071) & (!g2074)) + ((g2108) & (g2109) & (!g2110) & (!g2111) & (g2071) & (!g2074)) + ((g2108) & (g2109) & (!g2110) & (g2111) & (!g2071) & (!g2074)) + ((g2108) & (g2109) & (!g2110) & (g2111) & (g2071) & (!g2074)) + ((g2108) & (g2109) & (!g2110) & (g2111) & (g2071) & (g2074)) + ((g2108) & (g2109) & (g2110) & (!g2111) & (!g2071) & (!g2074)) + ((g2108) & (g2109) & (g2110) & (!g2111) & (!g2071) & (g2074)) + ((g2108) & (g2109) & (g2110) & (!g2111) & (g2071) & (!g2074)) + ((g2108) & (g2109) & (g2110) & (g2111) & (!g2071) & (!g2074)) + ((g2108) & (g2109) & (g2110) & (g2111) & (!g2071) & (g2074)) + ((g2108) & (g2109) & (g2110) & (g2111) & (g2071) & (!g2074)) + ((g2108) & (g2109) & (g2110) & (g2111) & (g2071) & (g2074)));
	assign g2117 = (((!g2113) & (!g2114) & (!g2115) & (g2116) & (g2071) & (g2074)) + ((!g2113) & (!g2114) & (g2115) & (!g2116) & (!g2071) & (g2074)) + ((!g2113) & (!g2114) & (g2115) & (g2116) & (!g2071) & (g2074)) + ((!g2113) & (!g2114) & (g2115) & (g2116) & (g2071) & (g2074)) + ((!g2113) & (g2114) & (!g2115) & (!g2116) & (g2071) & (!g2074)) + ((!g2113) & (g2114) & (!g2115) & (g2116) & (g2071) & (!g2074)) + ((!g2113) & (g2114) & (!g2115) & (g2116) & (g2071) & (g2074)) + ((!g2113) & (g2114) & (g2115) & (!g2116) & (!g2071) & (g2074)) + ((!g2113) & (g2114) & (g2115) & (!g2116) & (g2071) & (!g2074)) + ((!g2113) & (g2114) & (g2115) & (g2116) & (!g2071) & (g2074)) + ((!g2113) & (g2114) & (g2115) & (g2116) & (g2071) & (!g2074)) + ((!g2113) & (g2114) & (g2115) & (g2116) & (g2071) & (g2074)) + ((g2113) & (!g2114) & (!g2115) & (!g2116) & (!g2071) & (!g2074)) + ((g2113) & (!g2114) & (!g2115) & (g2116) & (!g2071) & (!g2074)) + ((g2113) & (!g2114) & (!g2115) & (g2116) & (g2071) & (g2074)) + ((g2113) & (!g2114) & (g2115) & (!g2116) & (!g2071) & (!g2074)) + ((g2113) & (!g2114) & (g2115) & (!g2116) & (!g2071) & (g2074)) + ((g2113) & (!g2114) & (g2115) & (g2116) & (!g2071) & (!g2074)) + ((g2113) & (!g2114) & (g2115) & (g2116) & (!g2071) & (g2074)) + ((g2113) & (!g2114) & (g2115) & (g2116) & (g2071) & (g2074)) + ((g2113) & (g2114) & (!g2115) & (!g2116) & (!g2071) & (!g2074)) + ((g2113) & (g2114) & (!g2115) & (!g2116) & (g2071) & (!g2074)) + ((g2113) & (g2114) & (!g2115) & (g2116) & (!g2071) & (!g2074)) + ((g2113) & (g2114) & (!g2115) & (g2116) & (g2071) & (!g2074)) + ((g2113) & (g2114) & (!g2115) & (g2116) & (g2071) & (g2074)) + ((g2113) & (g2114) & (g2115) & (!g2116) & (!g2071) & (!g2074)) + ((g2113) & (g2114) & (g2115) & (!g2116) & (!g2071) & (g2074)) + ((g2113) & (g2114) & (g2115) & (!g2116) & (g2071) & (!g2074)) + ((g2113) & (g2114) & (g2115) & (g2116) & (!g2071) & (!g2074)) + ((g2113) & (g2114) & (g2115) & (g2116) & (!g2071) & (g2074)) + ((g2113) & (g2114) & (g2115) & (g2116) & (g2071) & (!g2074)) + ((g2113) & (g2114) & (g2115) & (g2116) & (g2071) & (g2074)));
	assign g2122 = (((!g2118) & (!g2119) & (!g2120) & (g2121) & (g2071) & (g2074)) + ((!g2118) & (!g2119) & (g2120) & (!g2121) & (!g2071) & (g2074)) + ((!g2118) & (!g2119) & (g2120) & (g2121) & (!g2071) & (g2074)) + ((!g2118) & (!g2119) & (g2120) & (g2121) & (g2071) & (g2074)) + ((!g2118) & (g2119) & (!g2120) & (!g2121) & (g2071) & (!g2074)) + ((!g2118) & (g2119) & (!g2120) & (g2121) & (g2071) & (!g2074)) + ((!g2118) & (g2119) & (!g2120) & (g2121) & (g2071) & (g2074)) + ((!g2118) & (g2119) & (g2120) & (!g2121) & (!g2071) & (g2074)) + ((!g2118) & (g2119) & (g2120) & (!g2121) & (g2071) & (!g2074)) + ((!g2118) & (g2119) & (g2120) & (g2121) & (!g2071) & (g2074)) + ((!g2118) & (g2119) & (g2120) & (g2121) & (g2071) & (!g2074)) + ((!g2118) & (g2119) & (g2120) & (g2121) & (g2071) & (g2074)) + ((g2118) & (!g2119) & (!g2120) & (!g2121) & (!g2071) & (!g2074)) + ((g2118) & (!g2119) & (!g2120) & (g2121) & (!g2071) & (!g2074)) + ((g2118) & (!g2119) & (!g2120) & (g2121) & (g2071) & (g2074)) + ((g2118) & (!g2119) & (g2120) & (!g2121) & (!g2071) & (!g2074)) + ((g2118) & (!g2119) & (g2120) & (!g2121) & (!g2071) & (g2074)) + ((g2118) & (!g2119) & (g2120) & (g2121) & (!g2071) & (!g2074)) + ((g2118) & (!g2119) & (g2120) & (g2121) & (!g2071) & (g2074)) + ((g2118) & (!g2119) & (g2120) & (g2121) & (g2071) & (g2074)) + ((g2118) & (g2119) & (!g2120) & (!g2121) & (!g2071) & (!g2074)) + ((g2118) & (g2119) & (!g2120) & (!g2121) & (g2071) & (!g2074)) + ((g2118) & (g2119) & (!g2120) & (g2121) & (!g2071) & (!g2074)) + ((g2118) & (g2119) & (!g2120) & (g2121) & (g2071) & (!g2074)) + ((g2118) & (g2119) & (!g2120) & (g2121) & (g2071) & (g2074)) + ((g2118) & (g2119) & (g2120) & (!g2121) & (!g2071) & (!g2074)) + ((g2118) & (g2119) & (g2120) & (!g2121) & (!g2071) & (g2074)) + ((g2118) & (g2119) & (g2120) & (!g2121) & (g2071) & (!g2074)) + ((g2118) & (g2119) & (g2120) & (g2121) & (!g2071) & (!g2074)) + ((g2118) & (g2119) & (g2120) & (g2121) & (!g2071) & (g2074)) + ((g2118) & (g2119) & (g2120) & (g2121) & (g2071) & (!g2074)) + ((g2118) & (g2119) & (g2120) & (g2121) & (g2071) & (g2074)));
	assign g2123 = (((!g2107) & (!g2112) & (!g2117) & (g2122) & (g2076) & (g2077)) + ((!g2107) & (!g2112) & (g2117) & (!g2122) & (!g2076) & (g2077)) + ((!g2107) & (!g2112) & (g2117) & (g2122) & (!g2076) & (g2077)) + ((!g2107) & (!g2112) & (g2117) & (g2122) & (g2076) & (g2077)) + ((!g2107) & (g2112) & (!g2117) & (!g2122) & (g2076) & (!g2077)) + ((!g2107) & (g2112) & (!g2117) & (g2122) & (g2076) & (!g2077)) + ((!g2107) & (g2112) & (!g2117) & (g2122) & (g2076) & (g2077)) + ((!g2107) & (g2112) & (g2117) & (!g2122) & (!g2076) & (g2077)) + ((!g2107) & (g2112) & (g2117) & (!g2122) & (g2076) & (!g2077)) + ((!g2107) & (g2112) & (g2117) & (g2122) & (!g2076) & (g2077)) + ((!g2107) & (g2112) & (g2117) & (g2122) & (g2076) & (!g2077)) + ((!g2107) & (g2112) & (g2117) & (g2122) & (g2076) & (g2077)) + ((g2107) & (!g2112) & (!g2117) & (!g2122) & (!g2076) & (!g2077)) + ((g2107) & (!g2112) & (!g2117) & (g2122) & (!g2076) & (!g2077)) + ((g2107) & (!g2112) & (!g2117) & (g2122) & (g2076) & (g2077)) + ((g2107) & (!g2112) & (g2117) & (!g2122) & (!g2076) & (!g2077)) + ((g2107) & (!g2112) & (g2117) & (!g2122) & (!g2076) & (g2077)) + ((g2107) & (!g2112) & (g2117) & (g2122) & (!g2076) & (!g2077)) + ((g2107) & (!g2112) & (g2117) & (g2122) & (!g2076) & (g2077)) + ((g2107) & (!g2112) & (g2117) & (g2122) & (g2076) & (g2077)) + ((g2107) & (g2112) & (!g2117) & (!g2122) & (!g2076) & (!g2077)) + ((g2107) & (g2112) & (!g2117) & (!g2122) & (g2076) & (!g2077)) + ((g2107) & (g2112) & (!g2117) & (g2122) & (!g2076) & (!g2077)) + ((g2107) & (g2112) & (!g2117) & (g2122) & (g2076) & (!g2077)) + ((g2107) & (g2112) & (!g2117) & (g2122) & (g2076) & (g2077)) + ((g2107) & (g2112) & (g2117) & (!g2122) & (!g2076) & (!g2077)) + ((g2107) & (g2112) & (g2117) & (!g2122) & (!g2076) & (g2077)) + ((g2107) & (g2112) & (g2117) & (!g2122) & (g2076) & (!g2077)) + ((g2107) & (g2112) & (g2117) & (g2122) & (!g2076) & (!g2077)) + ((g2107) & (g2112) & (g2117) & (g2122) & (!g2076) & (g2077)) + ((g2107) & (g2112) & (g2117) & (g2122) & (g2076) & (!g2077)) + ((g2107) & (g2112) & (g2117) & (g2122) & (g2076) & (g2077)));
	assign g2126 = (((!g3801) & (!g2082) & (!g3788) & (!g2070) & (g2124) & (!g2125)) + ((!g3801) & (!g2082) & (!g3788) & (g2070) & (g2124) & (!g2125)) + ((!g3801) & (!g2082) & (!g3788) & (g2070) & (g2124) & (g2125)) + ((!g3801) & (!g2082) & (g3788) & (!g2070) & (!g2124) & (g2125)) + ((!g3801) & (!g2082) & (g3788) & (!g2070) & (g2124) & (!g2125)) + ((!g3801) & (!g2082) & (g3788) & (g2070) & (!g2124) & (g2125)) + ((!g3801) & (!g2082) & (g3788) & (g2070) & (g2124) & (!g2125)) + ((!g3801) & (!g2082) & (g3788) & (g2070) & (g2124) & (g2125)) + ((!g3801) & (g2082) & (!g3788) & (g2070) & (g2124) & (g2125)) + ((!g3801) & (g2082) & (g3788) & (!g2070) & (!g2124) & (g2125)) + ((!g3801) & (g2082) & (g3788) & (g2070) & (!g2124) & (g2125)) + ((!g3801) & (g2082) & (g3788) & (g2070) & (g2124) & (g2125)) + ((g3801) & (!g2082) & (!g3788) & (!g2070) & (!g2124) & (!g2125)) + ((g3801) & (!g2082) & (!g3788) & (!g2070) & (g2124) & (!g2125)) + ((g3801) & (!g2082) & (!g3788) & (g2070) & (!g2124) & (!g2125)) + ((g3801) & (!g2082) & (!g3788) & (g2070) & (g2124) & (!g2125)) + ((g3801) & (!g2082) & (!g3788) & (g2070) & (g2124) & (g2125)) + ((g3801) & (!g2082) & (g3788) & (!g2070) & (!g2124) & (!g2125)) + ((g3801) & (!g2082) & (g3788) & (!g2070) & (!g2124) & (g2125)) + ((g3801) & (!g2082) & (g3788) & (!g2070) & (g2124) & (!g2125)) + ((g3801) & (!g2082) & (g3788) & (g2070) & (!g2124) & (!g2125)) + ((g3801) & (!g2082) & (g3788) & (g2070) & (!g2124) & (g2125)) + ((g3801) & (!g2082) & (g3788) & (g2070) & (g2124) & (!g2125)) + ((g3801) & (!g2082) & (g3788) & (g2070) & (g2124) & (g2125)) + ((g3801) & (g2082) & (!g3788) & (!g2070) & (!g2124) & (!g2125)) + ((g3801) & (g2082) & (!g3788) & (g2070) & (!g2124) & (!g2125)) + ((g3801) & (g2082) & (!g3788) & (g2070) & (g2124) & (g2125)) + ((g3801) & (g2082) & (g3788) & (!g2070) & (!g2124) & (!g2125)) + ((g3801) & (g2082) & (g3788) & (!g2070) & (!g2124) & (g2125)) + ((g3801) & (g2082) & (g3788) & (g2070) & (!g2124) & (!g2125)) + ((g3801) & (g2082) & (g3788) & (g2070) & (!g2124) & (g2125)) + ((g3801) & (g2082) & (g3788) & (g2070) & (g2124) & (g2125)));
	assign g2127 = (((!g78) & (!g79) & (!g80) & (!g81) & (!g82) & (!g83)) + ((!g78) & (!g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((!g78) & (!g79) & (!g80) & (!g81) & (g82) & (!g83)) + ((!g78) & (!g79) & (!g80) & (!g81) & (g82) & (g83)) + ((!g78) & (!g79) & (!g80) & (g81) & (!g82) & (!g83)) + ((!g78) & (!g79) & (!g80) & (g81) & (!g82) & (g83)) + ((!g78) & (!g79) & (!g80) & (g81) & (g82) & (!g83)) + ((!g78) & (!g79) & (!g80) & (g81) & (g82) & (g83)) + ((!g78) & (!g79) & (g80) & (!g81) & (!g82) & (!g83)) + ((!g78) & (!g79) & (g80) & (!g81) & (!g82) & (g83)) + ((!g78) & (!g79) & (g80) & (!g81) & (g82) & (!g83)) + ((!g78) & (!g79) & (g80) & (!g81) & (g82) & (g83)) + ((!g78) & (!g79) & (g80) & (g81) & (!g82) & (!g83)) + ((!g78) & (!g79) & (g80) & (g81) & (!g82) & (g83)) + ((!g78) & (!g79) & (g80) & (g81) & (g82) & (!g83)) + ((!g78) & (!g79) & (g80) & (g81) & (g82) & (g83)) + ((!g78) & (g79) & (!g80) & (!g81) & (!g82) & (!g83)) + ((!g78) & (g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((!g78) & (g79) & (!g80) & (!g81) & (g82) & (!g83)) + ((!g78) & (g79) & (!g80) & (!g81) & (g82) & (g83)) + ((!g78) & (g79) & (!g80) & (g81) & (!g82) & (!g83)) + ((!g78) & (g79) & (!g80) & (g81) & (!g82) & (g83)) + ((!g78) & (g79) & (!g80) & (g81) & (g82) & (!g83)) + ((!g78) & (g79) & (!g80) & (g81) & (g82) & (g83)) + ((!g78) & (g79) & (g80) & (!g81) & (!g82) & (!g83)) + ((!g78) & (g79) & (g80) & (!g81) & (g82) & (!g83)) + ((!g78) & (g79) & (g80) & (!g81) & (g82) & (g83)) + ((!g78) & (g79) & (g80) & (g81) & (!g82) & (!g83)) + ((!g78) & (g79) & (g80) & (g81) & (!g82) & (g83)) + ((!g78) & (g79) & (g80) & (g81) & (g82) & (!g83)) + ((!g78) & (g79) & (g80) & (g81) & (g82) & (g83)) + ((g78) & (!g79) & (!g80) & (!g81) & (!g82) & (!g83)) + ((g78) & (!g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((g78) & (!g79) & (!g80) & (!g81) & (g82) & (!g83)) + ((g78) & (!g79) & (!g80) & (!g81) & (g82) & (g83)) + ((g78) & (!g79) & (!g80) & (g81) & (!g82) & (!g83)) + ((g78) & (!g79) & (!g80) & (g81) & (!g82) & (g83)) + ((g78) & (!g79) & (!g80) & (g81) & (g82) & (!g83)) + ((g78) & (!g79) & (!g80) & (g81) & (g82) & (g83)) + ((g78) & (!g79) & (g80) & (!g81) & (g82) & (!g83)) + ((g78) & (!g79) & (g80) & (!g81) & (g82) & (g83)) + ((g78) & (!g79) & (g80) & (g81) & (!g82) & (!g83)) + ((g78) & (!g79) & (g80) & (g81) & (!g82) & (g83)) + ((g78) & (!g79) & (g80) & (g81) & (g82) & (!g83)) + ((g78) & (!g79) & (g80) & (g81) & (g82) & (g83)) + ((g78) & (g79) & (!g80) & (!g81) & (!g82) & (!g83)) + ((g78) & (g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((g78) & (g79) & (!g80) & (!g81) & (g82) & (!g83)) + ((g78) & (g79) & (!g80) & (!g81) & (g82) & (g83)) + ((g78) & (g79) & (!g80) & (g81) & (!g82) & (!g83)) + ((g78) & (g79) & (!g80) & (g81) & (!g82) & (g83)) + ((g78) & (g79) & (!g80) & (g81) & (g82) & (!g83)) + ((g78) & (g79) & (!g80) & (g81) & (g82) & (g83)) + ((g78) & (g79) & (g80) & (!g81) & (!g82) & (g83)) + ((g78) & (g79) & (g80) & (!g81) & (g82) & (!g83)) + ((g78) & (g79) & (g80) & (!g81) & (g82) & (g83)) + ((g78) & (g79) & (g80) & (g81) & (!g82) & (!g83)) + ((g78) & (g79) & (g80) & (g81) & (!g82) & (g83)) + ((g78) & (g79) & (g80) & (g81) & (g82) & (!g83)) + ((g78) & (g79) & (g80) & (g81) & (g82) & (g83)));
	assign g5025 = (((!sk[103]) & (!g1609) & (!g1593) & (g2128)) + ((!sk[103]) & (!g1609) & (g1593) & (!g2128)) + ((!sk[103]) & (!g1609) & (g1593) & (g2128)) + ((!sk[103]) & (g1609) & (!g1593) & (g2128)) + ((!sk[103]) & (g1609) & (g1593) & (!g2128)) + ((!sk[103]) & (g1609) & (g1593) & (g2128)) + ((sk[103]) & (!g1609) & (!g1593) & (g2128)) + ((sk[103]) & (!g1609) & (g1593) & (g2128)) + ((sk[103]) & (g1609) & (g1593) & (!g2128)) + ((sk[103]) & (g1609) & (g1593) & (g2128)));
	assign g5026 = (((!g1609) & (!g1605) & (!sk[104]) & (g2129)) + ((!g1609) & (!g1605) & (sk[104]) & (g2129)) + ((!g1609) & (g1605) & (!sk[104]) & (!g2129)) + ((!g1609) & (g1605) & (!sk[104]) & (g2129)) + ((!g1609) & (g1605) & (sk[104]) & (g2129)) + ((g1609) & (!g1605) & (!sk[104]) & (g2129)) + ((g1609) & (g1605) & (!sk[104]) & (!g2129)) + ((g1609) & (g1605) & (!sk[104]) & (g2129)) + ((g1609) & (g1605) & (sk[104]) & (!g2129)) + ((g1609) & (g1605) & (sk[104]) & (g2129)));
	assign g2130 = (((!dmem_dat_ix24x) & (!dmem_dat_ix16x) & (!dmem_dat_ix8x) & (dmem_dat_ix0x) & (g2128) & (g2129)) + ((!dmem_dat_ix24x) & (!dmem_dat_ix16x) & (dmem_dat_ix8x) & (!dmem_dat_ix0x) & (!g2128) & (g2129)) + ((!dmem_dat_ix24x) & (!dmem_dat_ix16x) & (dmem_dat_ix8x) & (dmem_dat_ix0x) & (!g2128) & (g2129)) + ((!dmem_dat_ix24x) & (!dmem_dat_ix16x) & (dmem_dat_ix8x) & (dmem_dat_ix0x) & (g2128) & (g2129)) + ((!dmem_dat_ix24x) & (dmem_dat_ix16x) & (!dmem_dat_ix8x) & (!dmem_dat_ix0x) & (g2128) & (!g2129)) + ((!dmem_dat_ix24x) & (dmem_dat_ix16x) & (!dmem_dat_ix8x) & (dmem_dat_ix0x) & (g2128) & (!g2129)) + ((!dmem_dat_ix24x) & (dmem_dat_ix16x) & (!dmem_dat_ix8x) & (dmem_dat_ix0x) & (g2128) & (g2129)) + ((!dmem_dat_ix24x) & (dmem_dat_ix16x) & (dmem_dat_ix8x) & (!dmem_dat_ix0x) & (!g2128) & (g2129)) + ((!dmem_dat_ix24x) & (dmem_dat_ix16x) & (dmem_dat_ix8x) & (!dmem_dat_ix0x) & (g2128) & (!g2129)) + ((!dmem_dat_ix24x) & (dmem_dat_ix16x) & (dmem_dat_ix8x) & (dmem_dat_ix0x) & (!g2128) & (g2129)) + ((!dmem_dat_ix24x) & (dmem_dat_ix16x) & (dmem_dat_ix8x) & (dmem_dat_ix0x) & (g2128) & (!g2129)) + ((!dmem_dat_ix24x) & (dmem_dat_ix16x) & (dmem_dat_ix8x) & (dmem_dat_ix0x) & (g2128) & (g2129)) + ((dmem_dat_ix24x) & (!dmem_dat_ix16x) & (!dmem_dat_ix8x) & (!dmem_dat_ix0x) & (!g2128) & (!g2129)) + ((dmem_dat_ix24x) & (!dmem_dat_ix16x) & (!dmem_dat_ix8x) & (dmem_dat_ix0x) & (!g2128) & (!g2129)) + ((dmem_dat_ix24x) & (!dmem_dat_ix16x) & (!dmem_dat_ix8x) & (dmem_dat_ix0x) & (g2128) & (g2129)) + ((dmem_dat_ix24x) & (!dmem_dat_ix16x) & (dmem_dat_ix8x) & (!dmem_dat_ix0x) & (!g2128) & (!g2129)) + ((dmem_dat_ix24x) & (!dmem_dat_ix16x) & (dmem_dat_ix8x) & (!dmem_dat_ix0x) & (!g2128) & (g2129)) + ((dmem_dat_ix24x) & (!dmem_dat_ix16x) & (dmem_dat_ix8x) & (dmem_dat_ix0x) & (!g2128) & (!g2129)) + ((dmem_dat_ix24x) & (!dmem_dat_ix16x) & (dmem_dat_ix8x) & (dmem_dat_ix0x) & (!g2128) & (g2129)) + ((dmem_dat_ix24x) & (!dmem_dat_ix16x) & (dmem_dat_ix8x) & (dmem_dat_ix0x) & (g2128) & (g2129)) + ((dmem_dat_ix24x) & (dmem_dat_ix16x) & (!dmem_dat_ix8x) & (!dmem_dat_ix0x) & (!g2128) & (!g2129)) + ((dmem_dat_ix24x) & (dmem_dat_ix16x) & (!dmem_dat_ix8x) & (!dmem_dat_ix0x) & (g2128) & (!g2129)) + ((dmem_dat_ix24x) & (dmem_dat_ix16x) & (!dmem_dat_ix8x) & (dmem_dat_ix0x) & (!g2128) & (!g2129)) + ((dmem_dat_ix24x) & (dmem_dat_ix16x) & (!dmem_dat_ix8x) & (dmem_dat_ix0x) & (g2128) & (!g2129)) + ((dmem_dat_ix24x) & (dmem_dat_ix16x) & (!dmem_dat_ix8x) & (dmem_dat_ix0x) & (g2128) & (g2129)) + ((dmem_dat_ix24x) & (dmem_dat_ix16x) & (dmem_dat_ix8x) & (!dmem_dat_ix0x) & (!g2128) & (!g2129)) + ((dmem_dat_ix24x) & (dmem_dat_ix16x) & (dmem_dat_ix8x) & (!dmem_dat_ix0x) & (!g2128) & (g2129)) + ((dmem_dat_ix24x) & (dmem_dat_ix16x) & (dmem_dat_ix8x) & (!dmem_dat_ix0x) & (g2128) & (!g2129)) + ((dmem_dat_ix24x) & (dmem_dat_ix16x) & (dmem_dat_ix8x) & (dmem_dat_ix0x) & (!g2128) & (!g2129)) + ((dmem_dat_ix24x) & (dmem_dat_ix16x) & (dmem_dat_ix8x) & (dmem_dat_ix0x) & (!g2128) & (g2129)) + ((dmem_dat_ix24x) & (dmem_dat_ix16x) & (dmem_dat_ix8x) & (dmem_dat_ix0x) & (g2128) & (!g2129)) + ((dmem_dat_ix24x) & (dmem_dat_ix16x) & (dmem_dat_ix8x) & (dmem_dat_ix0x) & (g2128) & (g2129)));
	assign g2131 = (((!g78) & (!g79) & (!g80) & (!g81) & (!g82) & (!g83)) + ((!g78) & (!g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((!g78) & (!g79) & (!g80) & (!g81) & (g82) & (!g83)) + ((!g78) & (!g79) & (!g80) & (!g81) & (g82) & (g83)) + ((!g78) & (!g79) & (!g80) & (g81) & (!g82) & (!g83)) + ((!g78) & (!g79) & (!g80) & (g81) & (!g82) & (g83)) + ((!g78) & (!g79) & (!g80) & (g81) & (g82) & (!g83)) + ((!g78) & (!g79) & (!g80) & (g81) & (g82) & (g83)) + ((!g78) & (!g79) & (g80) & (!g81) & (!g82) & (!g83)) + ((!g78) & (!g79) & (g80) & (!g81) & (!g82) & (g83)) + ((!g78) & (!g79) & (g80) & (!g81) & (g82) & (!g83)) + ((!g78) & (!g79) & (g80) & (!g81) & (g82) & (g83)) + ((!g78) & (!g79) & (g80) & (g81) & (!g82) & (!g83)) + ((!g78) & (!g79) & (g80) & (g81) & (!g82) & (g83)) + ((!g78) & (!g79) & (g80) & (g81) & (g82) & (!g83)) + ((!g78) & (!g79) & (g80) & (g81) & (g82) & (g83)) + ((!g78) & (g79) & (!g80) & (!g81) & (!g82) & (!g83)) + ((!g78) & (g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((!g78) & (g79) & (!g80) & (!g81) & (g82) & (!g83)) + ((!g78) & (g79) & (!g80) & (!g81) & (g82) & (g83)) + ((!g78) & (g79) & (!g80) & (g81) & (!g82) & (!g83)) + ((!g78) & (g79) & (!g80) & (g81) & (!g82) & (g83)) + ((!g78) & (g79) & (!g80) & (g81) & (g82) & (!g83)) + ((!g78) & (g79) & (!g80) & (g81) & (g82) & (g83)) + ((!g78) & (g79) & (g80) & (!g81) & (!g82) & (!g83)) + ((!g78) & (g79) & (g80) & (!g81) & (g82) & (!g83)) + ((!g78) & (g79) & (g80) & (!g81) & (g82) & (g83)) + ((!g78) & (g79) & (g80) & (g81) & (!g82) & (!g83)) + ((!g78) & (g79) & (g80) & (g81) & (!g82) & (g83)) + ((!g78) & (g79) & (g80) & (g81) & (g82) & (!g83)) + ((!g78) & (g79) & (g80) & (g81) & (g82) & (g83)) + ((g78) & (!g79) & (!g80) & (!g81) & (!g82) & (!g83)) + ((g78) & (!g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((g78) & (!g79) & (!g80) & (!g81) & (g82) & (!g83)) + ((g78) & (!g79) & (!g80) & (!g81) & (g82) & (g83)) + ((g78) & (!g79) & (!g80) & (g81) & (!g82) & (!g83)) + ((g78) & (!g79) & (!g80) & (g81) & (!g82) & (g83)) + ((g78) & (!g79) & (!g80) & (g81) & (g82) & (!g83)) + ((g78) & (!g79) & (!g80) & (g81) & (g82) & (g83)) + ((g78) & (!g79) & (g80) & (!g81) & (!g82) & (g83)) + ((g78) & (!g79) & (g80) & (!g81) & (g82) & (!g83)) + ((g78) & (!g79) & (g80) & (!g81) & (g82) & (g83)) + ((g78) & (!g79) & (g80) & (g81) & (!g82) & (!g83)) + ((g78) & (!g79) & (g80) & (g81) & (!g82) & (g83)) + ((g78) & (!g79) & (g80) & (g81) & (g82) & (!g83)) + ((g78) & (!g79) & (g80) & (g81) & (g82) & (g83)) + ((g78) & (g79) & (!g80) & (!g81) & (!g82) & (!g83)) + ((g78) & (g79) & (!g80) & (!g81) & (!g82) & (g83)) + ((g78) & (g79) & (!g80) & (!g81) & (g82) & (!g83)) + ((g78) & (g79) & (!g80) & (!g81) & (g82) & (g83)) + ((g78) & (g79) & (!g80) & (g81) & (!g82) & (!g83)) + ((g78) & (g79) & (!g80) & (g81) & (!g82) & (g83)) + ((g78) & (g79) & (!g80) & (g81) & (g82) & (!g83)) + ((g78) & (g79) & (!g80) & (g81) & (g82) & (g83)) + ((g78) & (g79) & (g80) & (!g81) & (!g82) & (!g83)) + ((g78) & (g79) & (g80) & (!g81) & (!g82) & (g83)) + ((g78) & (g79) & (g80) & (!g81) & (g82) & (!g83)) + ((g78) & (g79) & (g80) & (!g81) & (g82) & (g83)) + ((g78) & (g79) & (g80) & (g81) & (!g82) & (!g83)) + ((g78) & (g79) & (g80) & (g81) & (!g82) & (g83)) + ((g78) & (g79) & (g80) & (g81) & (g82) & (!g83)) + ((g78) & (g79) & (g80) & (g81) & (g82) & (g83)));
	assign g2132 = (((g78) & (!g79) & (g80) & (!g81) & (!g82) & (g83)) + ((g78) & (g79) & (g80) & (!g81) & (!g82) & (!g83)));
	assign g2133 = (((g2131) & (g2132) & (!dmem_dat_ix0x) & (dmem_dat_ix16x) & (!g2128) & (!g2129)) + ((g2131) & (g2132) & (dmem_dat_ix0x) & (!dmem_dat_ix16x) & (!g2128) & (g2129)) + ((g2131) & (g2132) & (dmem_dat_ix0x) & (dmem_dat_ix16x) & (!g2128) & (!g2129)) + ((g2131) & (g2132) & (dmem_dat_ix0x) & (dmem_dat_ix16x) & (!g2128) & (g2129)));
	assign g2139 = (((!g2136) & (!sk[109]) & (!g2137) & (g2138)) + ((!g2136) & (!sk[109]) & (g2137) & (!g2138)) + ((!g2136) & (!sk[109]) & (g2137) & (g2138)) + ((!g2136) & (sk[109]) & (g2137) & (!g2138)) + ((g2136) & (!sk[109]) & (!g2137) & (g2138)) + ((g2136) & (!sk[109]) & (g2137) & (!g2138)) + ((g2136) & (!sk[109]) & (g2137) & (g2138)));
	assign g2140 = (((!g74) & (dmem_ack_i) & (g75) & (!g2134) & (!g2135) & (g2139)) + ((g74) & (!dmem_ack_i) & (!g75) & (!g2134) & (!g2135) & (g2139)) + ((g74) & (!dmem_ack_i) & (g75) & (!g2134) & (!g2135) & (g2139)) + ((g74) & (dmem_ack_i) & (!g75) & (!g2134) & (!g2135) & (g2139)) + ((g74) & (dmem_ack_i) & (g75) & (!g2134) & (!g2135) & (g2139)));
	assign g2141 = (((!sk[111]) & (!g74) & (!dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((!sk[111]) & (!g74) & (!dmem_ack_i) & (!g75) & (g2134) & (g2135)) + ((!sk[111]) & (!g74) & (!dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((!sk[111]) & (!g74) & (!dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((!sk[111]) & (!g74) & (!dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((!sk[111]) & (!g74) & (!dmem_ack_i) & (g75) & (g2134) & (g2135)) + ((!sk[111]) & (!g74) & (dmem_ack_i) & (!g75) & (!g2134) & (!g2135)) + ((!sk[111]) & (!g74) & (dmem_ack_i) & (!g75) & (!g2134) & (g2135)) + ((!sk[111]) & (!g74) & (dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((!sk[111]) & (!g74) & (dmem_ack_i) & (!g75) & (g2134) & (g2135)) + ((!sk[111]) & (!g74) & (dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((!sk[111]) & (!g74) & (dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((!sk[111]) & (!g74) & (dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((!sk[111]) & (!g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135)) + ((!sk[111]) & (g74) & (!dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((!sk[111]) & (g74) & (!dmem_ack_i) & (!g75) & (g2134) & (g2135)) + ((!sk[111]) & (g74) & (!dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((!sk[111]) & (g74) & (!dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((!sk[111]) & (g74) & (!dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((!sk[111]) & (g74) & (!dmem_ack_i) & (g75) & (g2134) & (g2135)) + ((!sk[111]) & (g74) & (dmem_ack_i) & (!g75) & (!g2134) & (!g2135)) + ((!sk[111]) & (g74) & (dmem_ack_i) & (!g75) & (!g2134) & (g2135)) + ((!sk[111]) & (g74) & (dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((!sk[111]) & (g74) & (dmem_ack_i) & (!g75) & (g2134) & (g2135)) + ((!sk[111]) & (g74) & (dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((!sk[111]) & (g74) & (dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((!sk[111]) & (g74) & (dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((!sk[111]) & (g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135)) + ((sk[111]) & (!g74) & (dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((sk[111]) & (g74) & (!dmem_ack_i) & (!g75) & (!g2134) & (!g2135)) + ((sk[111]) & (g74) & (!dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((sk[111]) & (g74) & (dmem_ack_i) & (!g75) & (!g2134) & (!g2135)) + ((sk[111]) & (g74) & (dmem_ack_i) & (g75) & (!g2134) & (!g2135)));
	assign g2142 = (((!sk[112]) & (!g2141) & (!g2136) & (!g2137) & (g2138)) + ((!sk[112]) & (!g2141) & (!g2136) & (g2137) & (!g2138)) + ((!sk[112]) & (!g2141) & (!g2136) & (g2137) & (g2138)) + ((!sk[112]) & (!g2141) & (g2136) & (!g2137) & (!g2138)) + ((!sk[112]) & (!g2141) & (g2136) & (!g2137) & (g2138)) + ((!sk[112]) & (!g2141) & (g2136) & (g2137) & (!g2138)) + ((!sk[112]) & (!g2141) & (g2136) & (g2137) & (g2138)) + ((!sk[112]) & (g2141) & (!g2136) & (!g2137) & (g2138)) + ((!sk[112]) & (g2141) & (!g2136) & (g2137) & (!g2138)) + ((!sk[112]) & (g2141) & (!g2136) & (g2137) & (g2138)) + ((!sk[112]) & (g2141) & (g2136) & (!g2137) & (!g2138)) + ((!sk[112]) & (g2141) & (g2136) & (!g2137) & (g2138)) + ((!sk[112]) & (g2141) & (g2136) & (g2137) & (!g2138)) + ((!sk[112]) & (g2141) & (g2136) & (g2137) & (g2138)) + ((sk[112]) & (g2141) & (!g2136) & (g2137) & (g2138)));
	assign g2143 = (((!g74) & (dmem_ack_i) & (g75) & (!g2134) & (!g2135) & (g2136)) + ((g74) & (!dmem_ack_i) & (!g75) & (!g2134) & (!g2135) & (g2136)) + ((g74) & (!dmem_ack_i) & (g75) & (!g2134) & (!g2135) & (g2136)) + ((g74) & (dmem_ack_i) & (!g75) & (!g2134) & (!g2135) & (g2136)) + ((g74) & (dmem_ack_i) & (g75) & (!g2134) & (!g2135) & (g2136)));
	assign g2144 = (((!g2137) & (!g2138) & (!sk[114]) & (g2143)) + ((!g2137) & (g2138) & (!sk[114]) & (!g2143)) + ((!g2137) & (g2138) & (!sk[114]) & (g2143)) + ((g2137) & (!g2138) & (!sk[114]) & (g2143)) + ((g2137) & (!g2138) & (sk[114]) & (g2143)) + ((g2137) & (g2138) & (!sk[114]) & (!g2143)) + ((g2137) & (g2138) & (!sk[114]) & (g2143)));
	assign g2145 = (((!g2137) & (!g2138) & (!sk[115]) & (g2143)) + ((!g2137) & (g2138) & (!sk[115]) & (!g2143)) + ((!g2137) & (g2138) & (!sk[115]) & (g2143)) + ((g2137) & (!g2138) & (!sk[115]) & (g2143)) + ((g2137) & (g2138) & (!sk[115]) & (!g2143)) + ((g2137) & (g2138) & (!sk[115]) & (g2143)) + ((g2137) & (g2138) & (sk[115]) & (g2143)));
	assign g2146 = (((!g74) & (dmem_ack_i) & (g75) & (!g2134) & (g2135) & (g2139)) + ((g74) & (!dmem_ack_i) & (!g75) & (!g2134) & (g2135) & (g2139)) + ((g74) & (!dmem_ack_i) & (g75) & (!g2134) & (g2135) & (g2139)) + ((g74) & (dmem_ack_i) & (!g75) & (!g2134) & (g2135) & (g2139)) + ((g74) & (dmem_ack_i) & (g75) & (!g2134) & (g2135) & (g2139)));
	assign g2147 = (((!g2136) & (!sk[117]) & (!g2137) & (g2138)) + ((!g2136) & (!sk[117]) & (g2137) & (!g2138)) + ((!g2136) & (!sk[117]) & (g2137) & (g2138)) + ((!g2136) & (sk[117]) & (g2137) & (g2138)) + ((g2136) & (!sk[117]) & (!g2137) & (g2138)) + ((g2136) & (!sk[117]) & (g2137) & (!g2138)) + ((g2136) & (!sk[117]) & (g2137) & (g2138)));
	assign g2148 = (((!g74) & (dmem_ack_i) & (g75) & (!g2134) & (g2135) & (g2147)) + ((g74) & (!dmem_ack_i) & (!g75) & (!g2134) & (g2135) & (g2147)) + ((g74) & (!dmem_ack_i) & (g75) & (!g2134) & (g2135) & (g2147)) + ((g74) & (dmem_ack_i) & (!g75) & (!g2134) & (g2135) & (g2147)) + ((g74) & (dmem_ack_i) & (g75) & (!g2134) & (g2135) & (g2147)));
	assign g2149 = (((!sk[119]) & (!g74) & (!dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((!sk[119]) & (!g74) & (!dmem_ack_i) & (!g75) & (g2134) & (g2135)) + ((!sk[119]) & (!g74) & (!dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((!sk[119]) & (!g74) & (!dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((!sk[119]) & (!g74) & (!dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((!sk[119]) & (!g74) & (!dmem_ack_i) & (g75) & (g2134) & (g2135)) + ((!sk[119]) & (!g74) & (dmem_ack_i) & (!g75) & (!g2134) & (!g2135)) + ((!sk[119]) & (!g74) & (dmem_ack_i) & (!g75) & (!g2134) & (g2135)) + ((!sk[119]) & (!g74) & (dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((!sk[119]) & (!g74) & (dmem_ack_i) & (!g75) & (g2134) & (g2135)) + ((!sk[119]) & (!g74) & (dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((!sk[119]) & (!g74) & (dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((!sk[119]) & (!g74) & (dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((!sk[119]) & (!g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135)) + ((!sk[119]) & (g74) & (!dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((!sk[119]) & (g74) & (!dmem_ack_i) & (!g75) & (g2134) & (g2135)) + ((!sk[119]) & (g74) & (!dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((!sk[119]) & (g74) & (!dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((!sk[119]) & (g74) & (!dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((!sk[119]) & (g74) & (!dmem_ack_i) & (g75) & (g2134) & (g2135)) + ((!sk[119]) & (g74) & (dmem_ack_i) & (!g75) & (!g2134) & (!g2135)) + ((!sk[119]) & (g74) & (dmem_ack_i) & (!g75) & (!g2134) & (g2135)) + ((!sk[119]) & (g74) & (dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((!sk[119]) & (g74) & (dmem_ack_i) & (!g75) & (g2134) & (g2135)) + ((!sk[119]) & (g74) & (dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((!sk[119]) & (g74) & (dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((!sk[119]) & (g74) & (dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((!sk[119]) & (g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135)) + ((sk[119]) & (!g74) & (dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((sk[119]) & (g74) & (!dmem_ack_i) & (!g75) & (!g2134) & (g2135)) + ((sk[119]) & (g74) & (!dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((sk[119]) & (g74) & (dmem_ack_i) & (!g75) & (!g2134) & (g2135)) + ((sk[119]) & (g74) & (dmem_ack_i) & (g75) & (!g2134) & (g2135)));
	assign g2150 = (((!g2136) & (!sk[120]) & (!g2137) & (!g2138) & (g2149)) + ((!g2136) & (!sk[120]) & (!g2137) & (g2138) & (!g2149)) + ((!g2136) & (!sk[120]) & (!g2137) & (g2138) & (g2149)) + ((!g2136) & (!sk[120]) & (g2137) & (!g2138) & (!g2149)) + ((!g2136) & (!sk[120]) & (g2137) & (!g2138) & (g2149)) + ((!g2136) & (!sk[120]) & (g2137) & (g2138) & (!g2149)) + ((!g2136) & (!sk[120]) & (g2137) & (g2138) & (g2149)) + ((g2136) & (!sk[120]) & (!g2137) & (!g2138) & (g2149)) + ((g2136) & (!sk[120]) & (!g2137) & (g2138) & (!g2149)) + ((g2136) & (!sk[120]) & (!g2137) & (g2138) & (g2149)) + ((g2136) & (!sk[120]) & (g2137) & (!g2138) & (!g2149)) + ((g2136) & (!sk[120]) & (g2137) & (!g2138) & (g2149)) + ((g2136) & (!sk[120]) & (g2137) & (g2138) & (!g2149)) + ((g2136) & (!sk[120]) & (g2137) & (g2138) & (g2149)) + ((g2136) & (sk[120]) & (g2137) & (!g2138) & (g2149)));
	assign g2151 = (((!g2136) & (!sk[121]) & (!g2137) & (!g2138) & (g2149)) + ((!g2136) & (!sk[121]) & (!g2137) & (g2138) & (!g2149)) + ((!g2136) & (!sk[121]) & (!g2137) & (g2138) & (g2149)) + ((!g2136) & (!sk[121]) & (g2137) & (!g2138) & (!g2149)) + ((!g2136) & (!sk[121]) & (g2137) & (!g2138) & (g2149)) + ((!g2136) & (!sk[121]) & (g2137) & (g2138) & (!g2149)) + ((!g2136) & (!sk[121]) & (g2137) & (g2138) & (g2149)) + ((g2136) & (!sk[121]) & (!g2137) & (!g2138) & (g2149)) + ((g2136) & (!sk[121]) & (!g2137) & (g2138) & (!g2149)) + ((g2136) & (!sk[121]) & (!g2137) & (g2138) & (g2149)) + ((g2136) & (!sk[121]) & (g2137) & (!g2138) & (!g2149)) + ((g2136) & (!sk[121]) & (g2137) & (!g2138) & (g2149)) + ((g2136) & (!sk[121]) & (g2137) & (g2138) & (!g2149)) + ((g2136) & (!sk[121]) & (g2137) & (g2138) & (g2149)) + ((g2136) & (sk[121]) & (g2137) & (g2138) & (g2149)));
	assign g2152 = (((!g74) & (dmem_ack_i) & (g75) & (g2134) & (!g2135) & (g2139)) + ((g74) & (!dmem_ack_i) & (!g75) & (g2134) & (!g2135) & (g2139)) + ((g74) & (!dmem_ack_i) & (g75) & (g2134) & (!g2135) & (g2139)) + ((g74) & (dmem_ack_i) & (!g75) & (g2134) & (!g2135) & (g2139)) + ((g74) & (dmem_ack_i) & (g75) & (g2134) & (!g2135) & (g2139)));
	assign g2153 = (((!g74) & (dmem_ack_i) & (g75) & (g2134) & (!g2135) & (g2147)) + ((g74) & (!dmem_ack_i) & (!g75) & (g2134) & (!g2135) & (g2147)) + ((g74) & (!dmem_ack_i) & (g75) & (g2134) & (!g2135) & (g2147)) + ((g74) & (dmem_ack_i) & (!g75) & (g2134) & (!g2135) & (g2147)) + ((g74) & (dmem_ack_i) & (g75) & (g2134) & (!g2135) & (g2147)));
	assign g2154 = (((!g2136) & (!g2137) & (!sk[124]) & (g2138)) + ((!g2136) & (g2137) & (!sk[124]) & (!g2138)) + ((!g2136) & (g2137) & (!sk[124]) & (g2138)) + ((g2136) & (!g2137) & (!sk[124]) & (g2138)) + ((g2136) & (g2137) & (!sk[124]) & (!g2138)) + ((g2136) & (g2137) & (!sk[124]) & (g2138)) + ((g2136) & (g2137) & (sk[124]) & (!g2138)));
	assign g2155 = (((!g74) & (dmem_ack_i) & (g75) & (g2134) & (!g2135) & (g2154)) + ((g74) & (!dmem_ack_i) & (!g75) & (g2134) & (!g2135) & (g2154)) + ((g74) & (!dmem_ack_i) & (g75) & (g2134) & (!g2135) & (g2154)) + ((g74) & (dmem_ack_i) & (!g75) & (g2134) & (!g2135) & (g2154)) + ((g74) & (dmem_ack_i) & (g75) & (g2134) & (!g2135) & (g2154)));
	assign g2156 = (((!g2136) & (!g2137) & (!sk[126]) & (g2138)) + ((!g2136) & (g2137) & (!sk[126]) & (!g2138)) + ((!g2136) & (g2137) & (!sk[126]) & (g2138)) + ((g2136) & (!g2137) & (!sk[126]) & (g2138)) + ((g2136) & (g2137) & (!sk[126]) & (!g2138)) + ((g2136) & (g2137) & (!sk[126]) & (g2138)) + ((g2136) & (g2137) & (sk[126]) & (g2138)));
	assign g2157 = (((!g74) & (dmem_ack_i) & (g75) & (g2134) & (!g2135) & (g2156)) + ((g74) & (!dmem_ack_i) & (!g75) & (g2134) & (!g2135) & (g2156)) + ((g74) & (!dmem_ack_i) & (g75) & (g2134) & (!g2135) & (g2156)) + ((g74) & (dmem_ack_i) & (!g75) & (g2134) & (!g2135) & (g2156)) + ((g74) & (dmem_ack_i) & (g75) & (g2134) & (!g2135) & (g2156)));
	assign g2158 = (((!g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135) & (g2139)) + ((g74) & (!dmem_ack_i) & (!g75) & (g2134) & (g2135) & (g2139)) + ((g74) & (!dmem_ack_i) & (g75) & (g2134) & (g2135) & (g2139)) + ((g74) & (dmem_ack_i) & (!g75) & (g2134) & (g2135) & (g2139)) + ((g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135) & (g2139)));
	assign g2159 = (((!g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135) & (g2147)) + ((g74) & (!dmem_ack_i) & (!g75) & (g2134) & (g2135) & (g2147)) + ((g74) & (!dmem_ack_i) & (g75) & (g2134) & (g2135) & (g2147)) + ((g74) & (dmem_ack_i) & (!g75) & (g2134) & (g2135) & (g2147)) + ((g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135) & (g2147)));
	assign g2160 = (((!g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135) & (g2154)) + ((g74) & (!dmem_ack_i) & (!g75) & (g2134) & (g2135) & (g2154)) + ((g74) & (!dmem_ack_i) & (g75) & (g2134) & (g2135) & (g2154)) + ((g74) & (dmem_ack_i) & (!g75) & (g2134) & (g2135) & (g2154)) + ((g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135) & (g2154)));
	assign g2161 = (((!g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135) & (g2156)) + ((g74) & (!dmem_ack_i) & (!g75) & (g2134) & (g2135) & (g2156)) + ((g74) & (!dmem_ack_i) & (g75) & (g2134) & (g2135) & (g2156)) + ((g74) & (dmem_ack_i) & (!g75) & (g2134) & (g2135) & (g2156)) + ((g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135) & (g2156)));
	assign g2162 = (((!g2137) & (!sk[4]) & (!g2138) & (g2143)) + ((!g2137) & (!sk[4]) & (g2138) & (!g2143)) + ((!g2137) & (!sk[4]) & (g2138) & (g2143)) + ((!g2137) & (sk[4]) & (g2138) & (g2143)) + ((g2137) & (!sk[4]) & (!g2138) & (g2143)) + ((g2137) & (!sk[4]) & (g2138) & (!g2143)) + ((g2137) & (!sk[4]) & (g2138) & (g2143)));
	assign g2163 = (((!g74) & (dmem_ack_i) & (g75) & (!g2134) & (g2135) & (!g2137)) + ((g74) & (!dmem_ack_i) & (!g75) & (!g2134) & (g2135) & (!g2137)) + ((g74) & (!dmem_ack_i) & (g75) & (!g2134) & (g2135) & (!g2137)) + ((g74) & (dmem_ack_i) & (!g75) & (!g2134) & (g2135) & (!g2137)) + ((g74) & (dmem_ack_i) & (g75) & (!g2134) & (g2135) & (!g2137)));
	assign g2164 = (((!g2136) & (!sk[6]) & (!g2138) & (g2163)) + ((!g2136) & (!sk[6]) & (g2138) & (!g2163)) + ((!g2136) & (!sk[6]) & (g2138) & (g2163)) + ((g2136) & (!sk[6]) & (!g2138) & (g2163)) + ((g2136) & (!sk[6]) & (g2138) & (!g2163)) + ((g2136) & (!sk[6]) & (g2138) & (g2163)) + ((g2136) & (sk[6]) & (g2138) & (g2163)));
	assign g2165 = (((!g74) & (!sk[7]) & (!dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((!g74) & (!sk[7]) & (!dmem_ack_i) & (!g75) & (g2134) & (g2135)) + ((!g74) & (!sk[7]) & (!dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((!g74) & (!sk[7]) & (!dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((!g74) & (!sk[7]) & (!dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((!g74) & (!sk[7]) & (!dmem_ack_i) & (g75) & (g2134) & (g2135)) + ((!g74) & (!sk[7]) & (dmem_ack_i) & (!g75) & (!g2134) & (!g2135)) + ((!g74) & (!sk[7]) & (dmem_ack_i) & (!g75) & (!g2134) & (g2135)) + ((!g74) & (!sk[7]) & (dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((!g74) & (!sk[7]) & (dmem_ack_i) & (!g75) & (g2134) & (g2135)) + ((!g74) & (!sk[7]) & (dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((!g74) & (!sk[7]) & (dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((!g74) & (!sk[7]) & (dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((!g74) & (!sk[7]) & (dmem_ack_i) & (g75) & (g2134) & (g2135)) + ((!g74) & (sk[7]) & (dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((g74) & (!sk[7]) & (!dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((g74) & (!sk[7]) & (!dmem_ack_i) & (!g75) & (g2134) & (g2135)) + ((g74) & (!sk[7]) & (!dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((g74) & (!sk[7]) & (!dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((g74) & (!sk[7]) & (!dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((g74) & (!sk[7]) & (!dmem_ack_i) & (g75) & (g2134) & (g2135)) + ((g74) & (!sk[7]) & (dmem_ack_i) & (!g75) & (!g2134) & (!g2135)) + ((g74) & (!sk[7]) & (dmem_ack_i) & (!g75) & (!g2134) & (g2135)) + ((g74) & (!sk[7]) & (dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((g74) & (!sk[7]) & (dmem_ack_i) & (!g75) & (g2134) & (g2135)) + ((g74) & (!sk[7]) & (dmem_ack_i) & (g75) & (!g2134) & (!g2135)) + ((g74) & (!sk[7]) & (dmem_ack_i) & (g75) & (!g2134) & (g2135)) + ((g74) & (!sk[7]) & (dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((g74) & (!sk[7]) & (dmem_ack_i) & (g75) & (g2134) & (g2135)) + ((g74) & (sk[7]) & (!dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((g74) & (sk[7]) & (!dmem_ack_i) & (g75) & (g2134) & (!g2135)) + ((g74) & (sk[7]) & (dmem_ack_i) & (!g75) & (g2134) & (!g2135)) + ((g74) & (sk[7]) & (dmem_ack_i) & (g75) & (g2134) & (!g2135)));
	assign g2166 = (((!g2136) & (!g2137) & (!g2138) & (!sk[8]) & (g2165)) + ((!g2136) & (!g2137) & (g2138) & (!sk[8]) & (!g2165)) + ((!g2136) & (!g2137) & (g2138) & (!sk[8]) & (g2165)) + ((!g2136) & (g2137) & (!g2138) & (!sk[8]) & (!g2165)) + ((!g2136) & (g2137) & (!g2138) & (!sk[8]) & (g2165)) + ((!g2136) & (g2137) & (g2138) & (!sk[8]) & (!g2165)) + ((!g2136) & (g2137) & (g2138) & (!sk[8]) & (g2165)) + ((g2136) & (!g2137) & (!g2138) & (!sk[8]) & (g2165)) + ((g2136) & (!g2137) & (g2138) & (!sk[8]) & (!g2165)) + ((g2136) & (!g2137) & (g2138) & (!sk[8]) & (g2165)) + ((g2136) & (!g2137) & (g2138) & (sk[8]) & (g2165)) + ((g2136) & (g2137) & (!g2138) & (!sk[8]) & (!g2165)) + ((g2136) & (g2137) & (!g2138) & (!sk[8]) & (g2165)) + ((g2136) & (g2137) & (g2138) & (!sk[8]) & (!g2165)) + ((g2136) & (g2137) & (g2138) & (!sk[8]) & (g2165)));
	assign g2167 = (((!g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135) & (!g2137)) + ((g74) & (!dmem_ack_i) & (!g75) & (g2134) & (g2135) & (!g2137)) + ((g74) & (!dmem_ack_i) & (g75) & (g2134) & (g2135) & (!g2137)) + ((g74) & (dmem_ack_i) & (!g75) & (g2134) & (g2135) & (!g2137)) + ((g74) & (dmem_ack_i) & (g75) & (g2134) & (g2135) & (!g2137)));
	assign g2168 = (((!g2136) & (!g2138) & (!sk[10]) & (g2167)) + ((!g2136) & (g2138) & (!sk[10]) & (!g2167)) + ((!g2136) & (g2138) & (!sk[10]) & (g2167)) + ((g2136) & (!g2138) & (!sk[10]) & (g2167)) + ((g2136) & (g2138) & (!sk[10]) & (!g2167)) + ((g2136) & (g2138) & (!sk[10]) & (g2167)) + ((g2136) & (g2138) & (sk[10]) & (g2167)));
	assign g2169 = (((!g2137) & (!sk[11]) & (!g2138) & (g2143)) + ((!g2137) & (!sk[11]) & (g2138) & (!g2143)) + ((!g2137) & (!sk[11]) & (g2138) & (g2143)) + ((!g2137) & (sk[11]) & (!g2138) & (g2143)) + ((g2137) & (!sk[11]) & (!g2138) & (g2143)) + ((g2137) & (!sk[11]) & (g2138) & (!g2143)) + ((g2137) & (!sk[11]) & (g2138) & (g2143)));
	assign g2170 = (((!g2136) & (!g2138) & (!sk[12]) & (g2163)) + ((!g2136) & (g2138) & (!sk[12]) & (!g2163)) + ((!g2136) & (g2138) & (!sk[12]) & (g2163)) + ((g2136) & (!g2138) & (!sk[12]) & (g2163)) + ((g2136) & (!g2138) & (sk[12]) & (g2163)) + ((g2136) & (g2138) & (!sk[12]) & (!g2163)) + ((g2136) & (g2138) & (!sk[12]) & (g2163)));
	assign g2171 = (((!sk[13]) & (!g2136) & (!g2137) & (!g2138) & (g2165)) + ((!sk[13]) & (!g2136) & (!g2137) & (g2138) & (!g2165)) + ((!sk[13]) & (!g2136) & (!g2137) & (g2138) & (g2165)) + ((!sk[13]) & (!g2136) & (g2137) & (!g2138) & (!g2165)) + ((!sk[13]) & (!g2136) & (g2137) & (!g2138) & (g2165)) + ((!sk[13]) & (!g2136) & (g2137) & (g2138) & (!g2165)) + ((!sk[13]) & (!g2136) & (g2137) & (g2138) & (g2165)) + ((!sk[13]) & (g2136) & (!g2137) & (!g2138) & (g2165)) + ((!sk[13]) & (g2136) & (!g2137) & (g2138) & (!g2165)) + ((!sk[13]) & (g2136) & (!g2137) & (g2138) & (g2165)) + ((!sk[13]) & (g2136) & (g2137) & (!g2138) & (!g2165)) + ((!sk[13]) & (g2136) & (g2137) & (!g2138) & (g2165)) + ((!sk[13]) & (g2136) & (g2137) & (g2138) & (!g2165)) + ((!sk[13]) & (g2136) & (g2137) & (g2138) & (g2165)) + ((sk[13]) & (g2136) & (!g2137) & (!g2138) & (g2165)));
	assign g2172 = (((!g2136) & (!sk[14]) & (!g2138) & (g2167)) + ((!g2136) & (!sk[14]) & (g2138) & (!g2167)) + ((!g2136) & (!sk[14]) & (g2138) & (g2167)) + ((g2136) & (!sk[14]) & (!g2138) & (g2167)) + ((g2136) & (!sk[14]) & (g2138) & (!g2167)) + ((g2136) & (!sk[14]) & (g2138) & (g2167)) + ((g2136) & (sk[14]) & (!g2138) & (g2167)));
	assign g2173 = (((!g2141) & (!g2136) & (!sk[15]) & (!g2137) & (g2138)) + ((!g2141) & (!g2136) & (!sk[15]) & (g2137) & (!g2138)) + ((!g2141) & (!g2136) & (!sk[15]) & (g2137) & (g2138)) + ((!g2141) & (g2136) & (!sk[15]) & (!g2137) & (!g2138)) + ((!g2141) & (g2136) & (!sk[15]) & (!g2137) & (g2138)) + ((!g2141) & (g2136) & (!sk[15]) & (g2137) & (!g2138)) + ((!g2141) & (g2136) & (!sk[15]) & (g2137) & (g2138)) + ((g2141) & (!g2136) & (!sk[15]) & (!g2137) & (g2138)) + ((g2141) & (!g2136) & (!sk[15]) & (g2137) & (!g2138)) + ((g2141) & (!g2136) & (!sk[15]) & (g2137) & (g2138)) + ((g2141) & (!g2136) & (sk[15]) & (!g2137) & (g2138)) + ((g2141) & (g2136) & (!sk[15]) & (!g2137) & (!g2138)) + ((g2141) & (g2136) & (!sk[15]) & (!g2137) & (g2138)) + ((g2141) & (g2136) & (!sk[15]) & (g2137) & (!g2138)) + ((g2141) & (g2136) & (!sk[15]) & (g2137) & (g2138)));
	assign g2174 = (((!g2136) & (!g2138) & (!sk[16]) & (g2163)) + ((!g2136) & (g2138) & (!sk[16]) & (!g2163)) + ((!g2136) & (g2138) & (!sk[16]) & (g2163)) + ((!g2136) & (g2138) & (sk[16]) & (g2163)) + ((g2136) & (!g2138) & (!sk[16]) & (g2163)) + ((g2136) & (g2138) & (!sk[16]) & (!g2163)) + ((g2136) & (g2138) & (!sk[16]) & (g2163)));
	assign g2175 = (((!g2136) & (!g2137) & (!sk[17]) & (!g2138) & (g2165)) + ((!g2136) & (!g2137) & (!sk[17]) & (g2138) & (!g2165)) + ((!g2136) & (!g2137) & (!sk[17]) & (g2138) & (g2165)) + ((!g2136) & (!g2137) & (sk[17]) & (g2138) & (g2165)) + ((!g2136) & (g2137) & (!sk[17]) & (!g2138) & (!g2165)) + ((!g2136) & (g2137) & (!sk[17]) & (!g2138) & (g2165)) + ((!g2136) & (g2137) & (!sk[17]) & (g2138) & (!g2165)) + ((!g2136) & (g2137) & (!sk[17]) & (g2138) & (g2165)) + ((g2136) & (!g2137) & (!sk[17]) & (!g2138) & (g2165)) + ((g2136) & (!g2137) & (!sk[17]) & (g2138) & (!g2165)) + ((g2136) & (!g2137) & (!sk[17]) & (g2138) & (g2165)) + ((g2136) & (g2137) & (!sk[17]) & (!g2138) & (!g2165)) + ((g2136) & (g2137) & (!sk[17]) & (!g2138) & (g2165)) + ((g2136) & (g2137) & (!sk[17]) & (g2138) & (!g2165)) + ((g2136) & (g2137) & (!sk[17]) & (g2138) & (g2165)));
	assign g2176 = (((!g2136) & (!g2138) & (!sk[18]) & (g2167)) + ((!g2136) & (g2138) & (!sk[18]) & (!g2167)) + ((!g2136) & (g2138) & (!sk[18]) & (g2167)) + ((!g2136) & (g2138) & (sk[18]) & (g2167)) + ((g2136) & (!g2138) & (!sk[18]) & (g2167)) + ((g2136) & (g2138) & (!sk[18]) & (!g2167)) + ((g2136) & (g2138) & (!sk[18]) & (g2167)));
	assign g2177 = (((!sk[19]) & (!g2136) & (!g2138) & (g2163)) + ((!sk[19]) & (!g2136) & (g2138) & (!g2163)) + ((!sk[19]) & (!g2136) & (g2138) & (g2163)) + ((!sk[19]) & (g2136) & (!g2138) & (g2163)) + ((!sk[19]) & (g2136) & (g2138) & (!g2163)) + ((!sk[19]) & (g2136) & (g2138) & (g2163)) + ((sk[19]) & (!g2136) & (!g2138) & (g2163)));
	assign g2178 = (((!g2136) & (!sk[20]) & (!g2138) & (g2167)) + ((!g2136) & (!sk[20]) & (g2138) & (!g2167)) + ((!g2136) & (!sk[20]) & (g2138) & (g2167)) + ((!g2136) & (sk[20]) & (!g2138) & (g2167)) + ((g2136) & (!sk[20]) & (!g2138) & (g2167)) + ((g2136) & (!sk[20]) & (g2138) & (!g2167)) + ((g2136) & (!sk[20]) & (g2138) & (g2167)));
	assign g2179 = (((!g2136) & (!g2137) & (!sk[21]) & (!g2138) & (g2165)) + ((!g2136) & (!g2137) & (!sk[21]) & (g2138) & (!g2165)) + ((!g2136) & (!g2137) & (!sk[21]) & (g2138) & (g2165)) + ((!g2136) & (!g2137) & (sk[21]) & (!g2138) & (g2165)) + ((!g2136) & (g2137) & (!sk[21]) & (!g2138) & (!g2165)) + ((!g2136) & (g2137) & (!sk[21]) & (!g2138) & (g2165)) + ((!g2136) & (g2137) & (!sk[21]) & (g2138) & (!g2165)) + ((!g2136) & (g2137) & (!sk[21]) & (g2138) & (g2165)) + ((g2136) & (!g2137) & (!sk[21]) & (!g2138) & (g2165)) + ((g2136) & (!g2137) & (!sk[21]) & (g2138) & (!g2165)) + ((g2136) & (!g2137) & (!sk[21]) & (g2138) & (g2165)) + ((g2136) & (g2137) & (!sk[21]) & (!g2138) & (!g2165)) + ((g2136) & (g2137) & (!sk[21]) & (!g2138) & (g2165)) + ((g2136) & (g2137) & (!sk[21]) & (g2138) & (!g2165)) + ((g2136) & (g2137) & (!sk[21]) & (g2138) & (g2165)));
	assign g2180 = (((g2131) & (!sk[22]) & (!g2132)) + ((g2131) & (!sk[22]) & (g2132)) + ((g2131) & (sk[22]) & (g2132)));
	assign g2181 = (((!sk[23]) & (!g2073) & (!g2074) & (!g2071) & (g2076) & (!g2077)) + ((!sk[23]) & (!g2073) & (!g2074) & (!g2071) & (g2076) & (g2077)) + ((!sk[23]) & (!g2073) & (!g2074) & (g2071) & (!g2076) & (!g2077)) + ((!sk[23]) & (!g2073) & (!g2074) & (g2071) & (!g2076) & (g2077)) + ((!sk[23]) & (!g2073) & (!g2074) & (g2071) & (g2076) & (!g2077)) + ((!sk[23]) & (!g2073) & (!g2074) & (g2071) & (g2076) & (g2077)) + ((!sk[23]) & (!g2073) & (g2074) & (!g2071) & (!g2076) & (!g2077)) + ((!sk[23]) & (!g2073) & (g2074) & (!g2071) & (!g2076) & (g2077)) + ((!sk[23]) & (!g2073) & (g2074) & (!g2071) & (g2076) & (!g2077)) + ((!sk[23]) & (!g2073) & (g2074) & (!g2071) & (g2076) & (g2077)) + ((!sk[23]) & (!g2073) & (g2074) & (g2071) & (!g2076) & (!g2077)) + ((!sk[23]) & (!g2073) & (g2074) & (g2071) & (!g2076) & (g2077)) + ((!sk[23]) & (!g2073) & (g2074) & (g2071) & (g2076) & (!g2077)) + ((!sk[23]) & (!g2073) & (g2074) & (g2071) & (g2076) & (g2077)) + ((!sk[23]) & (g2073) & (!g2074) & (!g2071) & (g2076) & (!g2077)) + ((!sk[23]) & (g2073) & (!g2074) & (!g2071) & (g2076) & (g2077)) + ((!sk[23]) & (g2073) & (!g2074) & (g2071) & (!g2076) & (!g2077)) + ((!sk[23]) & (g2073) & (!g2074) & (g2071) & (!g2076) & (g2077)) + ((!sk[23]) & (g2073) & (!g2074) & (g2071) & (g2076) & (!g2077)) + ((!sk[23]) & (g2073) & (!g2074) & (g2071) & (g2076) & (g2077)) + ((!sk[23]) & (g2073) & (g2074) & (!g2071) & (!g2076) & (!g2077)) + ((!sk[23]) & (g2073) & (g2074) & (!g2071) & (!g2076) & (g2077)) + ((!sk[23]) & (g2073) & (g2074) & (!g2071) & (g2076) & (!g2077)) + ((!sk[23]) & (g2073) & (g2074) & (!g2071) & (g2076) & (g2077)) + ((!sk[23]) & (g2073) & (g2074) & (g2071) & (!g2076) & (!g2077)) + ((!sk[23]) & (g2073) & (g2074) & (g2071) & (!g2076) & (g2077)) + ((!sk[23]) & (g2073) & (g2074) & (g2071) & (g2076) & (!g2077)) + ((!sk[23]) & (g2073) & (g2074) & (g2071) & (g2076) & (g2077)) + ((sk[23]) & (!g2073) & (!g2074) & (!g2071) & (!g2076) & (!g2077)));
	assign g2182 = (((!g2080) & (!sk[24]) & (!g2081) & (!g2124) & (g2125) & (!g2181)) + ((!g2080) & (!sk[24]) & (!g2081) & (!g2124) & (g2125) & (g2181)) + ((!g2080) & (!sk[24]) & (!g2081) & (g2124) & (!g2125) & (!g2181)) + ((!g2080) & (!sk[24]) & (!g2081) & (g2124) & (!g2125) & (g2181)) + ((!g2080) & (!sk[24]) & (!g2081) & (g2124) & (g2125) & (!g2181)) + ((!g2080) & (!sk[24]) & (!g2081) & (g2124) & (g2125) & (g2181)) + ((!g2080) & (!sk[24]) & (g2081) & (!g2124) & (!g2125) & (!g2181)) + ((!g2080) & (!sk[24]) & (g2081) & (!g2124) & (!g2125) & (g2181)) + ((!g2080) & (!sk[24]) & (g2081) & (!g2124) & (g2125) & (!g2181)) + ((!g2080) & (!sk[24]) & (g2081) & (!g2124) & (g2125) & (g2181)) + ((!g2080) & (!sk[24]) & (g2081) & (g2124) & (!g2125) & (!g2181)) + ((!g2080) & (!sk[24]) & (g2081) & (g2124) & (!g2125) & (g2181)) + ((!g2080) & (!sk[24]) & (g2081) & (g2124) & (g2125) & (!g2181)) + ((!g2080) & (!sk[24]) & (g2081) & (g2124) & (g2125) & (g2181)) + ((!g2080) & (sk[24]) & (!g2081) & (!g2124) & (!g2125) & (!g2181)) + ((!g2080) & (sk[24]) & (!g2081) & (!g2124) & (!g2125) & (g2181)) + ((!g2080) & (sk[24]) & (!g2081) & (!g2124) & (g2125) & (g2181)) + ((!g2080) & (sk[24]) & (!g2081) & (g2124) & (g2125) & (!g2181)) + ((!g2080) & (sk[24]) & (!g2081) & (g2124) & (g2125) & (g2181)) + ((!g2080) & (sk[24]) & (g2081) & (!g2124) & (g2125) & (g2181)) + ((!g2080) & (sk[24]) & (g2081) & (g2124) & (g2125) & (!g2181)) + ((!g2080) & (sk[24]) & (g2081) & (g2124) & (g2125) & (g2181)) + ((g2080) & (!sk[24]) & (!g2081) & (!g2124) & (g2125) & (!g2181)) + ((g2080) & (!sk[24]) & (!g2081) & (!g2124) & (g2125) & (g2181)) + ((g2080) & (!sk[24]) & (!g2081) & (g2124) & (!g2125) & (!g2181)) + ((g2080) & (!sk[24]) & (!g2081) & (g2124) & (!g2125) & (g2181)) + ((g2080) & (!sk[24]) & (!g2081) & (g2124) & (g2125) & (!g2181)) + ((g2080) & (!sk[24]) & (!g2081) & (g2124) & (g2125) & (g2181)) + ((g2080) & (!sk[24]) & (g2081) & (!g2124) & (!g2125) & (!g2181)) + ((g2080) & (!sk[24]) & (g2081) & (!g2124) & (!g2125) & (g2181)) + ((g2080) & (!sk[24]) & (g2081) & (!g2124) & (g2125) & (!g2181)) + ((g2080) & (!sk[24]) & (g2081) & (!g2124) & (g2125) & (g2181)) + ((g2080) & (!sk[24]) & (g2081) & (g2124) & (!g2125) & (!g2181)) + ((g2080) & (!sk[24]) & (g2081) & (g2124) & (!g2125) & (g2181)) + ((g2080) & (!sk[24]) & (g2081) & (g2124) & (g2125) & (!g2181)) + ((g2080) & (!sk[24]) & (g2081) & (g2124) & (g2125) & (g2181)) + ((g2080) & (sk[24]) & (!g2081) & (g2124) & (!g2125) & (!g2181)) + ((g2080) & (sk[24]) & (!g2081) & (g2124) & (!g2125) & (g2181)) + ((g2080) & (sk[24]) & (!g2081) & (g2124) & (g2125) & (!g2181)) + ((g2080) & (sk[24]) & (!g2081) & (g2124) & (g2125) & (g2181)) + ((g2080) & (sk[24]) & (g2081) & (g2124) & (!g2125) & (!g2181)) + ((g2080) & (sk[24]) & (g2081) & (g2124) & (!g2125) & (g2181)) + ((g2080) & (sk[24]) & (g2081) & (g2124) & (g2125) & (!g2181)) + ((g2080) & (sk[24]) & (g2081) & (g2124) & (g2125) & (g2181)));
	assign g2183 = (((!g2074) & (!sk[25]) & (!g2071) & (!g2070) & (g2104)) + ((!g2074) & (!sk[25]) & (!g2071) & (g2070) & (!g2104)) + ((!g2074) & (!sk[25]) & (!g2071) & (g2070) & (g2104)) + ((!g2074) & (!sk[25]) & (g2071) & (!g2070) & (!g2104)) + ((!g2074) & (!sk[25]) & (g2071) & (!g2070) & (g2104)) + ((!g2074) & (!sk[25]) & (g2071) & (g2070) & (!g2104)) + ((!g2074) & (!sk[25]) & (g2071) & (g2070) & (g2104)) + ((!g2074) & (sk[25]) & (!g2071) & (!g2070) & (g2104)) + ((!g2074) & (sk[25]) & (!g2071) & (g2070) & (g2104)) + ((!g2074) & (sk[25]) & (g2071) & (g2070) & (!g2104)) + ((!g2074) & (sk[25]) & (g2071) & (g2070) & (g2104)) + ((g2074) & (!sk[25]) & (!g2071) & (!g2070) & (g2104)) + ((g2074) & (!sk[25]) & (!g2071) & (g2070) & (!g2104)) + ((g2074) & (!sk[25]) & (!g2071) & (g2070) & (g2104)) + ((g2074) & (!sk[25]) & (g2071) & (!g2070) & (!g2104)) + ((g2074) & (!sk[25]) & (g2071) & (!g2070) & (g2104)) + ((g2074) & (!sk[25]) & (g2071) & (g2070) & (!g2104)) + ((g2074) & (!sk[25]) & (g2071) & (g2070) & (g2104)));
	assign g2184 = (((!g2076) & (!g2077) & (!sk[26]) & (g2183)) + ((!g2076) & (!g2077) & (sk[26]) & (g2183)) + ((!g2076) & (g2077) & (!sk[26]) & (!g2183)) + ((!g2076) & (g2077) & (!sk[26]) & (g2183)) + ((g2076) & (!g2077) & (!sk[26]) & (g2183)) + ((g2076) & (g2077) & (!sk[26]) & (!g2183)) + ((g2076) & (g2077) & (!sk[26]) & (g2183)));
	assign g2185 = (((!sk[27]) & (!g2074) & (!g2071) & (!g2070) & (g2104)) + ((!sk[27]) & (!g2074) & (!g2071) & (g2070) & (!g2104)) + ((!sk[27]) & (!g2074) & (!g2071) & (g2070) & (g2104)) + ((!sk[27]) & (!g2074) & (g2071) & (!g2070) & (!g2104)) + ((!sk[27]) & (!g2074) & (g2071) & (!g2070) & (g2104)) + ((!sk[27]) & (!g2074) & (g2071) & (g2070) & (!g2104)) + ((!sk[27]) & (!g2074) & (g2071) & (g2070) & (g2104)) + ((!sk[27]) & (g2074) & (!g2071) & (!g2070) & (g2104)) + ((!sk[27]) & (g2074) & (!g2071) & (g2070) & (!g2104)) + ((!sk[27]) & (g2074) & (!g2071) & (g2070) & (g2104)) + ((!sk[27]) & (g2074) & (g2071) & (!g2070) & (!g2104)) + ((!sk[27]) & (g2074) & (g2071) & (!g2070) & (g2104)) + ((!sk[27]) & (g2074) & (g2071) & (g2070) & (!g2104)) + ((!sk[27]) & (g2074) & (g2071) & (g2070) & (g2104)) + ((sk[27]) & (!g2074) & (!g2071) & (!g2070) & (g2104)) + ((sk[27]) & (!g2074) & (!g2071) & (g2070) & (g2104)) + ((sk[27]) & (!g2074) & (g2071) & (!g2070) & (g2104)) + ((sk[27]) & (!g2074) & (g2071) & (g2070) & (!g2104)) + ((sk[27]) & (g2074) & (!g2071) & (!g2070) & (!g2104)) + ((sk[27]) & (g2074) & (!g2071) & (g2070) & (!g2104)) + ((sk[27]) & (g2074) & (g2071) & (!g2070) & (!g2104)) + ((sk[27]) & (g2074) & (g2071) & (g2070) & (g2104)));
	assign g2186 = (((!sk[28]) & (g2071) & (!g2070)) + ((!sk[28]) & (g2071) & (g2070)) + ((sk[28]) & (g2071) & (!g2070)));
	assign g2187 = (((!g2084) & (!g2085) & (!g2086) & (g2093) & (g2071) & (g2074)) + ((!g2084) & (!g2085) & (g2086) & (!g2093) & (!g2071) & (g2074)) + ((!g2084) & (!g2085) & (g2086) & (g2093) & (!g2071) & (g2074)) + ((!g2084) & (!g2085) & (g2086) & (g2093) & (g2071) & (g2074)) + ((!g2084) & (g2085) & (!g2086) & (!g2093) & (g2071) & (!g2074)) + ((!g2084) & (g2085) & (!g2086) & (g2093) & (g2071) & (!g2074)) + ((!g2084) & (g2085) & (!g2086) & (g2093) & (g2071) & (g2074)) + ((!g2084) & (g2085) & (g2086) & (!g2093) & (!g2071) & (g2074)) + ((!g2084) & (g2085) & (g2086) & (!g2093) & (g2071) & (!g2074)) + ((!g2084) & (g2085) & (g2086) & (g2093) & (!g2071) & (g2074)) + ((!g2084) & (g2085) & (g2086) & (g2093) & (g2071) & (!g2074)) + ((!g2084) & (g2085) & (g2086) & (g2093) & (g2071) & (g2074)) + ((g2084) & (!g2085) & (!g2086) & (!g2093) & (!g2071) & (!g2074)) + ((g2084) & (!g2085) & (!g2086) & (g2093) & (!g2071) & (!g2074)) + ((g2084) & (!g2085) & (!g2086) & (g2093) & (g2071) & (g2074)) + ((g2084) & (!g2085) & (g2086) & (!g2093) & (!g2071) & (!g2074)) + ((g2084) & (!g2085) & (g2086) & (!g2093) & (!g2071) & (g2074)) + ((g2084) & (!g2085) & (g2086) & (g2093) & (!g2071) & (!g2074)) + ((g2084) & (!g2085) & (g2086) & (g2093) & (!g2071) & (g2074)) + ((g2084) & (!g2085) & (g2086) & (g2093) & (g2071) & (g2074)) + ((g2084) & (g2085) & (!g2086) & (!g2093) & (!g2071) & (!g2074)) + ((g2084) & (g2085) & (!g2086) & (!g2093) & (g2071) & (!g2074)) + ((g2084) & (g2085) & (!g2086) & (g2093) & (!g2071) & (!g2074)) + ((g2084) & (g2085) & (!g2086) & (g2093) & (g2071) & (!g2074)) + ((g2084) & (g2085) & (!g2086) & (g2093) & (g2071) & (g2074)) + ((g2084) & (g2085) & (g2086) & (!g2093) & (!g2071) & (!g2074)) + ((g2084) & (g2085) & (g2086) & (!g2093) & (!g2071) & (g2074)) + ((g2084) & (g2085) & (g2086) & (!g2093) & (g2071) & (!g2074)) + ((g2084) & (g2085) & (g2086) & (g2093) & (!g2071) & (!g2074)) + ((g2084) & (g2085) & (g2086) & (g2093) & (!g2071) & (g2074)) + ((g2084) & (g2085) & (g2086) & (g2093) & (g2071) & (!g2074)) + ((g2084) & (g2085) & (g2086) & (g2093) & (g2071) & (g2074)));
	assign g2188 = (((!g2089) & (!g2090) & (!g2091) & (g2098) & (g2071) & (g2074)) + ((!g2089) & (!g2090) & (g2091) & (!g2098) & (!g2071) & (g2074)) + ((!g2089) & (!g2090) & (g2091) & (g2098) & (!g2071) & (g2074)) + ((!g2089) & (!g2090) & (g2091) & (g2098) & (g2071) & (g2074)) + ((!g2089) & (g2090) & (!g2091) & (!g2098) & (g2071) & (!g2074)) + ((!g2089) & (g2090) & (!g2091) & (g2098) & (g2071) & (!g2074)) + ((!g2089) & (g2090) & (!g2091) & (g2098) & (g2071) & (g2074)) + ((!g2089) & (g2090) & (g2091) & (!g2098) & (!g2071) & (g2074)) + ((!g2089) & (g2090) & (g2091) & (!g2098) & (g2071) & (!g2074)) + ((!g2089) & (g2090) & (g2091) & (g2098) & (!g2071) & (g2074)) + ((!g2089) & (g2090) & (g2091) & (g2098) & (g2071) & (!g2074)) + ((!g2089) & (g2090) & (g2091) & (g2098) & (g2071) & (g2074)) + ((g2089) & (!g2090) & (!g2091) & (!g2098) & (!g2071) & (!g2074)) + ((g2089) & (!g2090) & (!g2091) & (g2098) & (!g2071) & (!g2074)) + ((g2089) & (!g2090) & (!g2091) & (g2098) & (g2071) & (g2074)) + ((g2089) & (!g2090) & (g2091) & (!g2098) & (!g2071) & (!g2074)) + ((g2089) & (!g2090) & (g2091) & (!g2098) & (!g2071) & (g2074)) + ((g2089) & (!g2090) & (g2091) & (g2098) & (!g2071) & (!g2074)) + ((g2089) & (!g2090) & (g2091) & (g2098) & (!g2071) & (g2074)) + ((g2089) & (!g2090) & (g2091) & (g2098) & (g2071) & (g2074)) + ((g2089) & (g2090) & (!g2091) & (!g2098) & (!g2071) & (!g2074)) + ((g2089) & (g2090) & (!g2091) & (!g2098) & (g2071) & (!g2074)) + ((g2089) & (g2090) & (!g2091) & (g2098) & (!g2071) & (!g2074)) + ((g2089) & (g2090) & (!g2091) & (g2098) & (g2071) & (!g2074)) + ((g2089) & (g2090) & (!g2091) & (g2098) & (g2071) & (g2074)) + ((g2089) & (g2090) & (g2091) & (!g2098) & (!g2071) & (!g2074)) + ((g2089) & (g2090) & (g2091) & (!g2098) & (!g2071) & (g2074)) + ((g2089) & (g2090) & (g2091) & (!g2098) & (g2071) & (!g2074)) + ((g2089) & (g2090) & (g2091) & (g2098) & (!g2071) & (!g2074)) + ((g2089) & (g2090) & (g2091) & (g2098) & (!g2071) & (g2074)) + ((g2089) & (g2090) & (g2091) & (g2098) & (g2071) & (!g2074)) + ((g2089) & (g2090) & (g2091) & (g2098) & (g2071) & (g2074)));
	assign g2189 = (((!g2094) & (!g2095) & (!g2096) & (g2088) & (g2071) & (g2074)) + ((!g2094) & (!g2095) & (g2096) & (!g2088) & (!g2071) & (g2074)) + ((!g2094) & (!g2095) & (g2096) & (g2088) & (!g2071) & (g2074)) + ((!g2094) & (!g2095) & (g2096) & (g2088) & (g2071) & (g2074)) + ((!g2094) & (g2095) & (!g2096) & (!g2088) & (g2071) & (!g2074)) + ((!g2094) & (g2095) & (!g2096) & (g2088) & (g2071) & (!g2074)) + ((!g2094) & (g2095) & (!g2096) & (g2088) & (g2071) & (g2074)) + ((!g2094) & (g2095) & (g2096) & (!g2088) & (!g2071) & (g2074)) + ((!g2094) & (g2095) & (g2096) & (!g2088) & (g2071) & (!g2074)) + ((!g2094) & (g2095) & (g2096) & (g2088) & (!g2071) & (g2074)) + ((!g2094) & (g2095) & (g2096) & (g2088) & (g2071) & (!g2074)) + ((!g2094) & (g2095) & (g2096) & (g2088) & (g2071) & (g2074)) + ((g2094) & (!g2095) & (!g2096) & (!g2088) & (!g2071) & (!g2074)) + ((g2094) & (!g2095) & (!g2096) & (g2088) & (!g2071) & (!g2074)) + ((g2094) & (!g2095) & (!g2096) & (g2088) & (g2071) & (g2074)) + ((g2094) & (!g2095) & (g2096) & (!g2088) & (!g2071) & (!g2074)) + ((g2094) & (!g2095) & (g2096) & (!g2088) & (!g2071) & (g2074)) + ((g2094) & (!g2095) & (g2096) & (g2088) & (!g2071) & (!g2074)) + ((g2094) & (!g2095) & (g2096) & (g2088) & (!g2071) & (g2074)) + ((g2094) & (!g2095) & (g2096) & (g2088) & (g2071) & (g2074)) + ((g2094) & (g2095) & (!g2096) & (!g2088) & (!g2071) & (!g2074)) + ((g2094) & (g2095) & (!g2096) & (!g2088) & (g2071) & (!g2074)) + ((g2094) & (g2095) & (!g2096) & (g2088) & (!g2071) & (!g2074)) + ((g2094) & (g2095) & (!g2096) & (g2088) & (g2071) & (!g2074)) + ((g2094) & (g2095) & (!g2096) & (g2088) & (g2071) & (g2074)) + ((g2094) & (g2095) & (g2096) & (!g2088) & (!g2071) & (!g2074)) + ((g2094) & (g2095) & (g2096) & (!g2088) & (!g2071) & (g2074)) + ((g2094) & (g2095) & (g2096) & (!g2088) & (g2071) & (!g2074)) + ((g2094) & (g2095) & (g2096) & (g2088) & (!g2071) & (!g2074)) + ((g2094) & (g2095) & (g2096) & (g2088) & (!g2071) & (g2074)) + ((g2094) & (g2095) & (g2096) & (g2088) & (g2071) & (!g2074)) + ((g2094) & (g2095) & (g2096) & (g2088) & (g2071) & (g2074)));
	assign g2190 = (((!sk[32]) & (g2080) & (!g2125)) + ((!sk[32]) & (g2080) & (g2125)) + ((sk[32]) & (!g2080) & (g2125)));
	assign g2191 = (((g2081) & (!sk[33]) & (!g2101)) + ((g2081) & (!sk[33]) & (g2101)) + ((g2081) & (sk[33]) & (g2101)));
	assign g2192 = (((!g2124) & (!g2190) & (!sk[34]) & (g2191)) + ((!g2124) & (g2190) & (!sk[34]) & (!g2191)) + ((!g2124) & (g2190) & (!sk[34]) & (g2191)) + ((!g2124) & (g2190) & (sk[34]) & (g2191)) + ((g2124) & (!g2190) & (!sk[34]) & (g2191)) + ((g2124) & (g2190) & (!sk[34]) & (!g2191)) + ((g2124) & (g2190) & (!sk[34]) & (g2191)));
	assign g2193 = (((!g2099) & (!g2100) & (!g2101) & (g2192) & (g2071) & (g2074)) + ((!g2099) & (!g2100) & (g2101) & (!g2192) & (!g2071) & (g2074)) + ((!g2099) & (!g2100) & (g2101) & (g2192) & (!g2071) & (g2074)) + ((!g2099) & (!g2100) & (g2101) & (g2192) & (g2071) & (g2074)) + ((!g2099) & (g2100) & (!g2101) & (!g2192) & (g2071) & (!g2074)) + ((!g2099) & (g2100) & (!g2101) & (g2192) & (g2071) & (!g2074)) + ((!g2099) & (g2100) & (!g2101) & (g2192) & (g2071) & (g2074)) + ((!g2099) & (g2100) & (g2101) & (!g2192) & (!g2071) & (g2074)) + ((!g2099) & (g2100) & (g2101) & (!g2192) & (g2071) & (!g2074)) + ((!g2099) & (g2100) & (g2101) & (g2192) & (!g2071) & (g2074)) + ((!g2099) & (g2100) & (g2101) & (g2192) & (g2071) & (!g2074)) + ((!g2099) & (g2100) & (g2101) & (g2192) & (g2071) & (g2074)) + ((g2099) & (!g2100) & (!g2101) & (!g2192) & (!g2071) & (!g2074)) + ((g2099) & (!g2100) & (!g2101) & (g2192) & (!g2071) & (!g2074)) + ((g2099) & (!g2100) & (!g2101) & (g2192) & (g2071) & (g2074)) + ((g2099) & (!g2100) & (g2101) & (!g2192) & (!g2071) & (!g2074)) + ((g2099) & (!g2100) & (g2101) & (!g2192) & (!g2071) & (g2074)) + ((g2099) & (!g2100) & (g2101) & (g2192) & (!g2071) & (!g2074)) + ((g2099) & (!g2100) & (g2101) & (g2192) & (!g2071) & (g2074)) + ((g2099) & (!g2100) & (g2101) & (g2192) & (g2071) & (g2074)) + ((g2099) & (g2100) & (!g2101) & (!g2192) & (!g2071) & (!g2074)) + ((g2099) & (g2100) & (!g2101) & (!g2192) & (g2071) & (!g2074)) + ((g2099) & (g2100) & (!g2101) & (g2192) & (!g2071) & (!g2074)) + ((g2099) & (g2100) & (!g2101) & (g2192) & (g2071) & (!g2074)) + ((g2099) & (g2100) & (!g2101) & (g2192) & (g2071) & (g2074)) + ((g2099) & (g2100) & (g2101) & (!g2192) & (!g2071) & (!g2074)) + ((g2099) & (g2100) & (g2101) & (!g2192) & (!g2071) & (g2074)) + ((g2099) & (g2100) & (g2101) & (!g2192) & (g2071) & (!g2074)) + ((g2099) & (g2100) & (g2101) & (g2192) & (!g2071) & (!g2074)) + ((g2099) & (g2100) & (g2101) & (g2192) & (!g2071) & (g2074)) + ((g2099) & (g2100) & (g2101) & (g2192) & (g2071) & (!g2074)) + ((g2099) & (g2100) & (g2101) & (g2192) & (g2071) & (g2074)));
	assign g2194 = (((!g2187) & (!g2188) & (!g2189) & (g2193) & (g2076) & (g2077)) + ((!g2187) & (!g2188) & (g2189) & (!g2193) & (!g2076) & (g2077)) + ((!g2187) & (!g2188) & (g2189) & (g2193) & (!g2076) & (g2077)) + ((!g2187) & (!g2188) & (g2189) & (g2193) & (g2076) & (g2077)) + ((!g2187) & (g2188) & (!g2189) & (!g2193) & (g2076) & (!g2077)) + ((!g2187) & (g2188) & (!g2189) & (g2193) & (g2076) & (!g2077)) + ((!g2187) & (g2188) & (!g2189) & (g2193) & (g2076) & (g2077)) + ((!g2187) & (g2188) & (g2189) & (!g2193) & (!g2076) & (g2077)) + ((!g2187) & (g2188) & (g2189) & (!g2193) & (g2076) & (!g2077)) + ((!g2187) & (g2188) & (g2189) & (g2193) & (!g2076) & (g2077)) + ((!g2187) & (g2188) & (g2189) & (g2193) & (g2076) & (!g2077)) + ((!g2187) & (g2188) & (g2189) & (g2193) & (g2076) & (g2077)) + ((g2187) & (!g2188) & (!g2189) & (!g2193) & (!g2076) & (!g2077)) + ((g2187) & (!g2188) & (!g2189) & (g2193) & (!g2076) & (!g2077)) + ((g2187) & (!g2188) & (!g2189) & (g2193) & (g2076) & (g2077)) + ((g2187) & (!g2188) & (g2189) & (!g2193) & (!g2076) & (!g2077)) + ((g2187) & (!g2188) & (g2189) & (!g2193) & (!g2076) & (g2077)) + ((g2187) & (!g2188) & (g2189) & (g2193) & (!g2076) & (!g2077)) + ((g2187) & (!g2188) & (g2189) & (g2193) & (!g2076) & (g2077)) + ((g2187) & (!g2188) & (g2189) & (g2193) & (g2076) & (g2077)) + ((g2187) & (g2188) & (!g2189) & (!g2193) & (!g2076) & (!g2077)) + ((g2187) & (g2188) & (!g2189) & (!g2193) & (g2076) & (!g2077)) + ((g2187) & (g2188) & (!g2189) & (g2193) & (!g2076) & (!g2077)) + ((g2187) & (g2188) & (!g2189) & (g2193) & (g2076) & (!g2077)) + ((g2187) & (g2188) & (!g2189) & (g2193) & (g2076) & (g2077)) + ((g2187) & (g2188) & (g2189) & (!g2193) & (!g2076) & (!g2077)) + ((g2187) & (g2188) & (g2189) & (!g2193) & (!g2076) & (g2077)) + ((g2187) & (g2188) & (g2189) & (!g2193) & (g2076) & (!g2077)) + ((g2187) & (g2188) & (g2189) & (g2193) & (!g2076) & (!g2077)) + ((g2187) & (g2188) & (g2189) & (g2193) & (!g2076) & (g2077)) + ((g2187) & (g2188) & (g2189) & (g2193) & (g2076) & (!g2077)) + ((g2187) & (g2188) & (g2189) & (g2193) & (g2076) & (g2077)));
	assign g2195 = (((!g2114) & (!g2115) & (!g2116) & (g2108) & (g2071) & (g2074)) + ((!g2114) & (!g2115) & (g2116) & (!g2108) & (!g2071) & (g2074)) + ((!g2114) & (!g2115) & (g2116) & (g2108) & (!g2071) & (g2074)) + ((!g2114) & (!g2115) & (g2116) & (g2108) & (g2071) & (g2074)) + ((!g2114) & (g2115) & (!g2116) & (!g2108) & (g2071) & (!g2074)) + ((!g2114) & (g2115) & (!g2116) & (g2108) & (g2071) & (!g2074)) + ((!g2114) & (g2115) & (!g2116) & (g2108) & (g2071) & (g2074)) + ((!g2114) & (g2115) & (g2116) & (!g2108) & (!g2071) & (g2074)) + ((!g2114) & (g2115) & (g2116) & (!g2108) & (g2071) & (!g2074)) + ((!g2114) & (g2115) & (g2116) & (g2108) & (!g2071) & (g2074)) + ((!g2114) & (g2115) & (g2116) & (g2108) & (g2071) & (!g2074)) + ((!g2114) & (g2115) & (g2116) & (g2108) & (g2071) & (g2074)) + ((g2114) & (!g2115) & (!g2116) & (!g2108) & (!g2071) & (!g2074)) + ((g2114) & (!g2115) & (!g2116) & (g2108) & (!g2071) & (!g2074)) + ((g2114) & (!g2115) & (!g2116) & (g2108) & (g2071) & (g2074)) + ((g2114) & (!g2115) & (g2116) & (!g2108) & (!g2071) & (!g2074)) + ((g2114) & (!g2115) & (g2116) & (!g2108) & (!g2071) & (g2074)) + ((g2114) & (!g2115) & (g2116) & (g2108) & (!g2071) & (!g2074)) + ((g2114) & (!g2115) & (g2116) & (g2108) & (!g2071) & (g2074)) + ((g2114) & (!g2115) & (g2116) & (g2108) & (g2071) & (g2074)) + ((g2114) & (g2115) & (!g2116) & (!g2108) & (!g2071) & (!g2074)) + ((g2114) & (g2115) & (!g2116) & (!g2108) & (g2071) & (!g2074)) + ((g2114) & (g2115) & (!g2116) & (g2108) & (!g2071) & (!g2074)) + ((g2114) & (g2115) & (!g2116) & (g2108) & (g2071) & (!g2074)) + ((g2114) & (g2115) & (!g2116) & (g2108) & (g2071) & (g2074)) + ((g2114) & (g2115) & (g2116) & (!g2108) & (!g2071) & (!g2074)) + ((g2114) & (g2115) & (g2116) & (!g2108) & (!g2071) & (g2074)) + ((g2114) & (g2115) & (g2116) & (!g2108) & (g2071) & (!g2074)) + ((g2114) & (g2115) & (g2116) & (g2108) & (!g2071) & (!g2074)) + ((g2114) & (g2115) & (g2116) & (g2108) & (!g2071) & (g2074)) + ((g2114) & (g2115) & (g2116) & (g2108) & (g2071) & (!g2074)) + ((g2114) & (g2115) & (g2116) & (g2108) & (g2071) & (g2074)));
	assign g2196 = (((!g2074) & (!sk[38]) & (!g2071) & (g2077)) + ((!g2074) & (!sk[38]) & (g2071) & (!g2077)) + ((!g2074) & (!sk[38]) & (g2071) & (g2077)) + ((!g2074) & (sk[38]) & (!g2071) & (!g2077)) + ((!g2074) & (sk[38]) & (g2071) & (!g2077)) + ((g2074) & (!sk[38]) & (!g2071) & (g2077)) + ((g2074) & (!sk[38]) & (g2071) & (!g2077)) + ((g2074) & (!sk[38]) & (g2071) & (g2077)) + ((g2074) & (sk[38]) & (g2071) & (!g2077)));
	assign g2197 = (((g2074) & (!sk[39]) & (!g2077)) + ((g2074) & (!sk[39]) & (g2077)) + ((g2074) & (sk[39]) & (!g2077)));
	assign g2198 = (((!g2195) & (!g2105) & (!g2106) & (g2113) & (g2196) & (g2197)) + ((!g2195) & (!g2105) & (g2106) & (!g2113) & (!g2196) & (g2197)) + ((!g2195) & (!g2105) & (g2106) & (g2113) & (!g2196) & (g2197)) + ((!g2195) & (!g2105) & (g2106) & (g2113) & (g2196) & (g2197)) + ((!g2195) & (g2105) & (!g2106) & (!g2113) & (g2196) & (!g2197)) + ((!g2195) & (g2105) & (!g2106) & (g2113) & (g2196) & (!g2197)) + ((!g2195) & (g2105) & (!g2106) & (g2113) & (g2196) & (g2197)) + ((!g2195) & (g2105) & (g2106) & (!g2113) & (!g2196) & (g2197)) + ((!g2195) & (g2105) & (g2106) & (!g2113) & (g2196) & (!g2197)) + ((!g2195) & (g2105) & (g2106) & (g2113) & (!g2196) & (g2197)) + ((!g2195) & (g2105) & (g2106) & (g2113) & (g2196) & (!g2197)) + ((!g2195) & (g2105) & (g2106) & (g2113) & (g2196) & (g2197)) + ((g2195) & (!g2105) & (!g2106) & (!g2113) & (!g2196) & (!g2197)) + ((g2195) & (!g2105) & (!g2106) & (g2113) & (!g2196) & (!g2197)) + ((g2195) & (!g2105) & (!g2106) & (g2113) & (g2196) & (g2197)) + ((g2195) & (!g2105) & (g2106) & (!g2113) & (!g2196) & (!g2197)) + ((g2195) & (!g2105) & (g2106) & (!g2113) & (!g2196) & (g2197)) + ((g2195) & (!g2105) & (g2106) & (g2113) & (!g2196) & (!g2197)) + ((g2195) & (!g2105) & (g2106) & (g2113) & (!g2196) & (g2197)) + ((g2195) & (!g2105) & (g2106) & (g2113) & (g2196) & (g2197)) + ((g2195) & (g2105) & (!g2106) & (!g2113) & (!g2196) & (!g2197)) + ((g2195) & (g2105) & (!g2106) & (!g2113) & (g2196) & (!g2197)) + ((g2195) & (g2105) & (!g2106) & (g2113) & (!g2196) & (!g2197)) + ((g2195) & (g2105) & (!g2106) & (g2113) & (g2196) & (!g2197)) + ((g2195) & (g2105) & (!g2106) & (g2113) & (g2196) & (g2197)) + ((g2195) & (g2105) & (g2106) & (!g2113) & (!g2196) & (!g2197)) + ((g2195) & (g2105) & (g2106) & (!g2113) & (!g2196) & (g2197)) + ((g2195) & (g2105) & (g2106) & (!g2113) & (g2196) & (!g2197)) + ((g2195) & (g2105) & (g2106) & (g2113) & (!g2196) & (!g2197)) + ((g2195) & (g2105) & (g2106) & (g2113) & (!g2196) & (g2197)) + ((g2195) & (g2105) & (g2106) & (g2113) & (g2196) & (!g2197)) + ((g2195) & (g2105) & (g2106) & (g2113) & (g2196) & (g2197)));
	assign g2199 = (((!g2109) & (!g2110) & (!g2111) & (g2118) & (g2071) & (g2074)) + ((!g2109) & (!g2110) & (g2111) & (!g2118) & (!g2071) & (g2074)) + ((!g2109) & (!g2110) & (g2111) & (g2118) & (!g2071) & (g2074)) + ((!g2109) & (!g2110) & (g2111) & (g2118) & (g2071) & (g2074)) + ((!g2109) & (g2110) & (!g2111) & (!g2118) & (g2071) & (!g2074)) + ((!g2109) & (g2110) & (!g2111) & (g2118) & (g2071) & (!g2074)) + ((!g2109) & (g2110) & (!g2111) & (g2118) & (g2071) & (g2074)) + ((!g2109) & (g2110) & (g2111) & (!g2118) & (!g2071) & (g2074)) + ((!g2109) & (g2110) & (g2111) & (!g2118) & (g2071) & (!g2074)) + ((!g2109) & (g2110) & (g2111) & (g2118) & (!g2071) & (g2074)) + ((!g2109) & (g2110) & (g2111) & (g2118) & (g2071) & (!g2074)) + ((!g2109) & (g2110) & (g2111) & (g2118) & (g2071) & (g2074)) + ((g2109) & (!g2110) & (!g2111) & (!g2118) & (!g2071) & (!g2074)) + ((g2109) & (!g2110) & (!g2111) & (g2118) & (!g2071) & (!g2074)) + ((g2109) & (!g2110) & (!g2111) & (g2118) & (g2071) & (g2074)) + ((g2109) & (!g2110) & (g2111) & (!g2118) & (!g2071) & (!g2074)) + ((g2109) & (!g2110) & (g2111) & (!g2118) & (!g2071) & (g2074)) + ((g2109) & (!g2110) & (g2111) & (g2118) & (!g2071) & (!g2074)) + ((g2109) & (!g2110) & (g2111) & (g2118) & (!g2071) & (g2074)) + ((g2109) & (!g2110) & (g2111) & (g2118) & (g2071) & (g2074)) + ((g2109) & (g2110) & (!g2111) & (!g2118) & (!g2071) & (!g2074)) + ((g2109) & (g2110) & (!g2111) & (!g2118) & (g2071) & (!g2074)) + ((g2109) & (g2110) & (!g2111) & (g2118) & (!g2071) & (!g2074)) + ((g2109) & (g2110) & (!g2111) & (g2118) & (g2071) & (!g2074)) + ((g2109) & (g2110) & (!g2111) & (g2118) & (g2071) & (g2074)) + ((g2109) & (g2110) & (g2111) & (!g2118) & (!g2071) & (!g2074)) + ((g2109) & (g2110) & (g2111) & (!g2118) & (!g2071) & (g2074)) + ((g2109) & (g2110) & (g2111) & (!g2118) & (g2071) & (!g2074)) + ((g2109) & (g2110) & (g2111) & (g2118) & (!g2071) & (!g2074)) + ((g2109) & (g2110) & (g2111) & (g2118) & (!g2071) & (g2074)) + ((g2109) & (g2110) & (g2111) & (g2118) & (g2071) & (!g2074)) + ((g2109) & (g2110) & (g2111) & (g2118) & (g2071) & (g2074)));
	assign g2200 = (((!g2119) & (!g2120) & (!g2121) & (g2083) & (g2071) & (g2074)) + ((!g2119) & (!g2120) & (g2121) & (!g2083) & (!g2071) & (g2074)) + ((!g2119) & (!g2120) & (g2121) & (g2083) & (!g2071) & (g2074)) + ((!g2119) & (!g2120) & (g2121) & (g2083) & (g2071) & (g2074)) + ((!g2119) & (g2120) & (!g2121) & (!g2083) & (g2071) & (!g2074)) + ((!g2119) & (g2120) & (!g2121) & (g2083) & (g2071) & (!g2074)) + ((!g2119) & (g2120) & (!g2121) & (g2083) & (g2071) & (g2074)) + ((!g2119) & (g2120) & (g2121) & (!g2083) & (!g2071) & (g2074)) + ((!g2119) & (g2120) & (g2121) & (!g2083) & (g2071) & (!g2074)) + ((!g2119) & (g2120) & (g2121) & (g2083) & (!g2071) & (g2074)) + ((!g2119) & (g2120) & (g2121) & (g2083) & (g2071) & (!g2074)) + ((!g2119) & (g2120) & (g2121) & (g2083) & (g2071) & (g2074)) + ((g2119) & (!g2120) & (!g2121) & (!g2083) & (!g2071) & (!g2074)) + ((g2119) & (!g2120) & (!g2121) & (g2083) & (!g2071) & (!g2074)) + ((g2119) & (!g2120) & (!g2121) & (g2083) & (g2071) & (g2074)) + ((g2119) & (!g2120) & (g2121) & (!g2083) & (!g2071) & (!g2074)) + ((g2119) & (!g2120) & (g2121) & (!g2083) & (!g2071) & (g2074)) + ((g2119) & (!g2120) & (g2121) & (g2083) & (!g2071) & (!g2074)) + ((g2119) & (!g2120) & (g2121) & (g2083) & (!g2071) & (g2074)) + ((g2119) & (!g2120) & (g2121) & (g2083) & (g2071) & (g2074)) + ((g2119) & (g2120) & (!g2121) & (!g2083) & (!g2071) & (!g2074)) + ((g2119) & (g2120) & (!g2121) & (!g2083) & (g2071) & (!g2074)) + ((g2119) & (g2120) & (!g2121) & (g2083) & (!g2071) & (!g2074)) + ((g2119) & (g2120) & (!g2121) & (g2083) & (g2071) & (!g2074)) + ((g2119) & (g2120) & (!g2121) & (g2083) & (g2071) & (g2074)) + ((g2119) & (g2120) & (g2121) & (!g2083) & (!g2071) & (!g2074)) + ((g2119) & (g2120) & (g2121) & (!g2083) & (!g2071) & (g2074)) + ((g2119) & (g2120) & (g2121) & (!g2083) & (g2071) & (!g2074)) + ((g2119) & (g2120) & (g2121) & (g2083) & (!g2071) & (!g2074)) + ((g2119) & (g2120) & (g2121) & (g2083) & (!g2071) & (g2074)) + ((g2119) & (g2120) & (g2121) & (g2083) & (g2071) & (!g2074)) + ((g2119) & (g2120) & (g2121) & (g2083) & (g2071) & (g2074)));
	assign g2201 = (((!g2073) & (!sk[43]) & (!g2076) & (g2077)) + ((!g2073) & (!sk[43]) & (g2076) & (!g2077)) + ((!g2073) & (!sk[43]) & (g2076) & (g2077)) + ((!g2073) & (sk[43]) & (!g2076) & (!g2077)) + ((!g2073) & (sk[43]) & (!g2076) & (g2077)) + ((!g2073) & (sk[43]) & (g2076) & (g2077)) + ((g2073) & (!sk[43]) & (!g2076) & (g2077)) + ((g2073) & (!sk[43]) & (g2076) & (!g2077)) + ((g2073) & (!sk[43]) & (g2076) & (g2077)));
	assign g2202 = (((!g2073) & (sk[44]) & (g2076)) + ((g2073) & (!sk[44]) & (!g2076)) + ((g2073) & (!sk[44]) & (g2076)));
	assign g2203 = (((!g2194) & (!g2198) & (!g2199) & (g2200) & (g2201) & (g2202)) + ((!g2194) & (!g2198) & (g2199) & (!g2200) & (!g2201) & (g2202)) + ((!g2194) & (!g2198) & (g2199) & (g2200) & (!g2201) & (g2202)) + ((!g2194) & (!g2198) & (g2199) & (g2200) & (g2201) & (g2202)) + ((!g2194) & (g2198) & (!g2199) & (!g2200) & (g2201) & (!g2202)) + ((!g2194) & (g2198) & (!g2199) & (g2200) & (g2201) & (!g2202)) + ((!g2194) & (g2198) & (!g2199) & (g2200) & (g2201) & (g2202)) + ((!g2194) & (g2198) & (g2199) & (!g2200) & (!g2201) & (g2202)) + ((!g2194) & (g2198) & (g2199) & (!g2200) & (g2201) & (!g2202)) + ((!g2194) & (g2198) & (g2199) & (g2200) & (!g2201) & (g2202)) + ((!g2194) & (g2198) & (g2199) & (g2200) & (g2201) & (!g2202)) + ((!g2194) & (g2198) & (g2199) & (g2200) & (g2201) & (g2202)) + ((g2194) & (!g2198) & (!g2199) & (!g2200) & (!g2201) & (!g2202)) + ((g2194) & (!g2198) & (!g2199) & (g2200) & (!g2201) & (!g2202)) + ((g2194) & (!g2198) & (!g2199) & (g2200) & (g2201) & (g2202)) + ((g2194) & (!g2198) & (g2199) & (!g2200) & (!g2201) & (!g2202)) + ((g2194) & (!g2198) & (g2199) & (!g2200) & (!g2201) & (g2202)) + ((g2194) & (!g2198) & (g2199) & (g2200) & (!g2201) & (!g2202)) + ((g2194) & (!g2198) & (g2199) & (g2200) & (!g2201) & (g2202)) + ((g2194) & (!g2198) & (g2199) & (g2200) & (g2201) & (g2202)) + ((g2194) & (g2198) & (!g2199) & (!g2200) & (!g2201) & (!g2202)) + ((g2194) & (g2198) & (!g2199) & (!g2200) & (g2201) & (!g2202)) + ((g2194) & (g2198) & (!g2199) & (g2200) & (!g2201) & (!g2202)) + ((g2194) & (g2198) & (!g2199) & (g2200) & (g2201) & (!g2202)) + ((g2194) & (g2198) & (!g2199) & (g2200) & (g2201) & (g2202)) + ((g2194) & (g2198) & (g2199) & (!g2200) & (!g2201) & (!g2202)) + ((g2194) & (g2198) & (g2199) & (!g2200) & (!g2201) & (g2202)) + ((g2194) & (g2198) & (g2199) & (!g2200) & (g2201) & (!g2202)) + ((g2194) & (g2198) & (g2199) & (g2200) & (!g2201) & (!g2202)) + ((g2194) & (g2198) & (g2199) & (g2200) & (!g2201) & (g2202)) + ((g2194) & (g2198) & (g2199) & (g2200) & (g2201) & (!g2202)) + ((g2194) & (g2198) & (g2199) & (g2200) & (g2201) & (g2202)));
	assign g2204 = (((!g2073) & (!g2080) & (!g2125) & (g2184) & (!g3147) & (!g2203)) + ((!g2073) & (!g2080) & (!g2125) & (g2184) & (!g3147) & (g2203)) + ((!g2073) & (!g2080) & (!g2125) & (g2184) & (g3147) & (!g2203)) + ((!g2073) & (!g2080) & (!g2125) & (g2184) & (g3147) & (g2203)) + ((!g2073) & (!g2080) & (g2125) & (!g2184) & (!g3147) & (g2203)) + ((!g2073) & (!g2080) & (g2125) & (!g2184) & (g3147) & (g2203)) + ((!g2073) & (!g2080) & (g2125) & (g2184) & (!g3147) & (g2203)) + ((!g2073) & (!g2080) & (g2125) & (g2184) & (g3147) & (g2203)) + ((!g2073) & (g2080) & (!g2125) & (!g2184) & (g3147) & (!g2203)) + ((!g2073) & (g2080) & (!g2125) & (!g2184) & (g3147) & (g2203)) + ((!g2073) & (g2080) & (!g2125) & (g2184) & (g3147) & (!g2203)) + ((!g2073) & (g2080) & (!g2125) & (g2184) & (g3147) & (g2203)) + ((!g2073) & (g2080) & (g2125) & (!g2184) & (g3147) & (!g2203)) + ((!g2073) & (g2080) & (g2125) & (!g2184) & (g3147) & (g2203)) + ((!g2073) & (g2080) & (g2125) & (g2184) & (g3147) & (!g2203)) + ((!g2073) & (g2080) & (g2125) & (g2184) & (g3147) & (g2203)) + ((g2073) & (!g2080) & (g2125) & (!g2184) & (!g3147) & (g2203)) + ((g2073) & (!g2080) & (g2125) & (!g2184) & (g3147) & (g2203)) + ((g2073) & (!g2080) & (g2125) & (g2184) & (!g3147) & (g2203)) + ((g2073) & (!g2080) & (g2125) & (g2184) & (g3147) & (g2203)) + ((g2073) & (g2080) & (!g2125) & (!g2184) & (g3147) & (!g2203)) + ((g2073) & (g2080) & (!g2125) & (!g2184) & (g3147) & (g2203)) + ((g2073) & (g2080) & (!g2125) & (g2184) & (g3147) & (!g2203)) + ((g2073) & (g2080) & (!g2125) & (g2184) & (g3147) & (g2203)) + ((g2073) & (g2080) & (g2125) & (!g2184) & (g3147) & (!g2203)) + ((g2073) & (g2080) & (g2125) & (!g2184) & (g3147) & (g2203)) + ((g2073) & (g2080) & (g2125) & (g2184) & (g3147) & (!g2203)) + ((g2073) & (g2080) & (g2125) & (g2184) & (g3147) & (g2203)));
	assign g2205 = (((!g2081) & (!g2124) & (!g2182) & (!g2074) & (!g2204) & (!g2104)) + ((!g2081) & (!g2124) & (!g2182) & (!g2074) & (!g2204) & (g2104)) + ((!g2081) & (!g2124) & (!g2182) & (g2074) & (!g2204) & (!g2104)) + ((!g2081) & (!g2124) & (!g2182) & (g2074) & (!g2204) & (g2104)) + ((!g2081) & (!g2124) & (g2182) & (!g2074) & (!g2204) & (!g2104)) + ((!g2081) & (!g2124) & (g2182) & (!g2074) & (g2204) & (!g2104)) + ((!g2081) & (!g2124) & (g2182) & (g2074) & (!g2204) & (!g2104)) + ((!g2081) & (!g2124) & (g2182) & (g2074) & (g2204) & (!g2104)) + ((!g2081) & (g2124) & (!g2182) & (!g2074) & (!g2204) & (!g2104)) + ((!g2081) & (g2124) & (!g2182) & (!g2074) & (g2204) & (!g2104)) + ((!g2081) & (g2124) & (g2182) & (!g2074) & (!g2204) & (!g2104)) + ((!g2081) & (g2124) & (g2182) & (!g2074) & (g2204) & (!g2104)) + ((!g2081) & (g2124) & (g2182) & (g2074) & (!g2204) & (!g2104)) + ((!g2081) & (g2124) & (g2182) & (g2074) & (g2204) & (!g2104)) + ((g2081) & (!g2124) & (!g2182) & (!g2074) & (!g2204) & (!g2104)) + ((g2081) & (!g2124) & (!g2182) & (!g2074) & (!g2204) & (g2104)) + ((g2081) & (!g2124) & (!g2182) & (g2074) & (!g2204) & (!g2104)) + ((g2081) & (!g2124) & (!g2182) & (g2074) & (!g2204) & (g2104)) + ((g2081) & (!g2124) & (g2182) & (!g2074) & (!g2204) & (!g2104)) + ((g2081) & (!g2124) & (g2182) & (!g2074) & (g2204) & (!g2104)) + ((g2081) & (!g2124) & (g2182) & (g2074) & (!g2204) & (!g2104)) + ((g2081) & (!g2124) & (g2182) & (g2074) & (g2204) & (!g2104)) + ((g2081) & (g2124) & (!g2182) & (!g2074) & (!g2204) & (!g2104)) + ((g2081) & (g2124) & (!g2182) & (!g2074) & (g2204) & (!g2104)) + ((g2081) & (g2124) & (!g2182) & (g2074) & (!g2204) & (g2104)) + ((g2081) & (g2124) & (!g2182) & (g2074) & (g2204) & (g2104)) + ((g2081) & (g2124) & (g2182) & (!g2074) & (!g2204) & (!g2104)) + ((g2081) & (g2124) & (g2182) & (!g2074) & (g2204) & (!g2104)) + ((g2081) & (g2124) & (g2182) & (g2074) & (!g2204) & (!g2104)) + ((g2081) & (g2124) & (g2182) & (g2074) & (g2204) & (!g2104)));
	assign g2206 = (((!g2131) & (!g2128) & (!sk[48]) & (g2129)) + ((!g2131) & (!g2128) & (sk[48]) & (g2129)) + ((!g2131) & (g2128) & (!sk[48]) & (!g2129)) + ((!g2131) & (g2128) & (!sk[48]) & (g2129)) + ((!g2131) & (g2128) & (sk[48]) & (!g2129)) + ((g2131) & (!g2128) & (!sk[48]) & (g2129)) + ((g2131) & (g2128) & (!sk[48]) & (!g2129)) + ((g2131) & (g2128) & (!sk[48]) & (g2129)));
	assign g2207 = (((!sk[49]) & (g2131) & (!g2129)) + ((!sk[49]) & (g2131) & (g2129)) + ((sk[49]) & (!g2131) & (!g2129)));
	assign g2208 = (((!dmem_dat_ix1x) & (!dmem_dat_ix9x) & (!dmem_dat_ix25x) & (dmem_dat_ix17x) & (g2206) & (g2207)) + ((!dmem_dat_ix1x) & (!dmem_dat_ix9x) & (dmem_dat_ix25x) & (!dmem_dat_ix17x) & (!g2206) & (g2207)) + ((!dmem_dat_ix1x) & (!dmem_dat_ix9x) & (dmem_dat_ix25x) & (dmem_dat_ix17x) & (!g2206) & (g2207)) + ((!dmem_dat_ix1x) & (!dmem_dat_ix9x) & (dmem_dat_ix25x) & (dmem_dat_ix17x) & (g2206) & (g2207)) + ((!dmem_dat_ix1x) & (dmem_dat_ix9x) & (!dmem_dat_ix25x) & (!dmem_dat_ix17x) & (g2206) & (!g2207)) + ((!dmem_dat_ix1x) & (dmem_dat_ix9x) & (!dmem_dat_ix25x) & (dmem_dat_ix17x) & (g2206) & (!g2207)) + ((!dmem_dat_ix1x) & (dmem_dat_ix9x) & (!dmem_dat_ix25x) & (dmem_dat_ix17x) & (g2206) & (g2207)) + ((!dmem_dat_ix1x) & (dmem_dat_ix9x) & (dmem_dat_ix25x) & (!dmem_dat_ix17x) & (!g2206) & (g2207)) + ((!dmem_dat_ix1x) & (dmem_dat_ix9x) & (dmem_dat_ix25x) & (!dmem_dat_ix17x) & (g2206) & (!g2207)) + ((!dmem_dat_ix1x) & (dmem_dat_ix9x) & (dmem_dat_ix25x) & (dmem_dat_ix17x) & (!g2206) & (g2207)) + ((!dmem_dat_ix1x) & (dmem_dat_ix9x) & (dmem_dat_ix25x) & (dmem_dat_ix17x) & (g2206) & (!g2207)) + ((!dmem_dat_ix1x) & (dmem_dat_ix9x) & (dmem_dat_ix25x) & (dmem_dat_ix17x) & (g2206) & (g2207)) + ((dmem_dat_ix1x) & (!dmem_dat_ix9x) & (!dmem_dat_ix25x) & (!dmem_dat_ix17x) & (!g2206) & (!g2207)) + ((dmem_dat_ix1x) & (!dmem_dat_ix9x) & (!dmem_dat_ix25x) & (dmem_dat_ix17x) & (!g2206) & (!g2207)) + ((dmem_dat_ix1x) & (!dmem_dat_ix9x) & (!dmem_dat_ix25x) & (dmem_dat_ix17x) & (g2206) & (g2207)) + ((dmem_dat_ix1x) & (!dmem_dat_ix9x) & (dmem_dat_ix25x) & (!dmem_dat_ix17x) & (!g2206) & (!g2207)) + ((dmem_dat_ix1x) & (!dmem_dat_ix9x) & (dmem_dat_ix25x) & (!dmem_dat_ix17x) & (!g2206) & (g2207)) + ((dmem_dat_ix1x) & (!dmem_dat_ix9x) & (dmem_dat_ix25x) & (dmem_dat_ix17x) & (!g2206) & (!g2207)) + ((dmem_dat_ix1x) & (!dmem_dat_ix9x) & (dmem_dat_ix25x) & (dmem_dat_ix17x) & (!g2206) & (g2207)) + ((dmem_dat_ix1x) & (!dmem_dat_ix9x) & (dmem_dat_ix25x) & (dmem_dat_ix17x) & (g2206) & (g2207)) + ((dmem_dat_ix1x) & (dmem_dat_ix9x) & (!dmem_dat_ix25x) & (!dmem_dat_ix17x) & (!g2206) & (!g2207)) + ((dmem_dat_ix1x) & (dmem_dat_ix9x) & (!dmem_dat_ix25x) & (!dmem_dat_ix17x) & (g2206) & (!g2207)) + ((dmem_dat_ix1x) & (dmem_dat_ix9x) & (!dmem_dat_ix25x) & (dmem_dat_ix17x) & (!g2206) & (!g2207)) + ((dmem_dat_ix1x) & (dmem_dat_ix9x) & (!dmem_dat_ix25x) & (dmem_dat_ix17x) & (g2206) & (!g2207)) + ((dmem_dat_ix1x) & (dmem_dat_ix9x) & (!dmem_dat_ix25x) & (dmem_dat_ix17x) & (g2206) & (g2207)) + ((dmem_dat_ix1x) & (dmem_dat_ix9x) & (dmem_dat_ix25x) & (!dmem_dat_ix17x) & (!g2206) & (!g2207)) + ((dmem_dat_ix1x) & (dmem_dat_ix9x) & (dmem_dat_ix25x) & (!dmem_dat_ix17x) & (!g2206) & (g2207)) + ((dmem_dat_ix1x) & (dmem_dat_ix9x) & (dmem_dat_ix25x) & (!dmem_dat_ix17x) & (g2206) & (!g2207)) + ((dmem_dat_ix1x) & (dmem_dat_ix9x) & (dmem_dat_ix25x) & (dmem_dat_ix17x) & (!g2206) & (!g2207)) + ((dmem_dat_ix1x) & (dmem_dat_ix9x) & (dmem_dat_ix25x) & (dmem_dat_ix17x) & (!g2206) & (g2207)) + ((dmem_dat_ix1x) & (dmem_dat_ix9x) & (dmem_dat_ix25x) & (dmem_dat_ix17x) & (g2206) & (!g2207)) + ((dmem_dat_ix1x) & (dmem_dat_ix9x) & (dmem_dat_ix25x) & (dmem_dat_ix17x) & (g2206) & (g2207)));
	assign g2209 = (((!dmem_dat_ix1x) & (!sk[51]) & (!g2129) & (dmem_dat_ix17x)) + ((!dmem_dat_ix1x) & (!sk[51]) & (g2129) & (!dmem_dat_ix17x)) + ((!dmem_dat_ix1x) & (!sk[51]) & (g2129) & (dmem_dat_ix17x)) + ((!dmem_dat_ix1x) & (sk[51]) & (!g2129) & (dmem_dat_ix17x)) + ((dmem_dat_ix1x) & (!sk[51]) & (!g2129) & (dmem_dat_ix17x)) + ((dmem_dat_ix1x) & (!sk[51]) & (g2129) & (!dmem_dat_ix17x)) + ((dmem_dat_ix1x) & (!sk[51]) & (g2129) & (dmem_dat_ix17x)) + ((dmem_dat_ix1x) & (sk[51]) & (!g2129) & (dmem_dat_ix17x)) + ((dmem_dat_ix1x) & (sk[51]) & (g2129) & (!dmem_dat_ix17x)) + ((dmem_dat_ix1x) & (sk[51]) & (g2129) & (dmem_dat_ix17x)));
	assign g2210 = (((!g75) & (!g2128) & (!g2180) & (!g2205) & (!g2208) & (!g2209)) + ((!g75) & (!g2128) & (!g2180) & (!g2205) & (!g2208) & (g2209)) + ((!g75) & (!g2128) & (!g2180) & (!g2205) & (g2208) & (!g2209)) + ((!g75) & (!g2128) & (!g2180) & (!g2205) & (g2208) & (g2209)) + ((!g75) & (!g2128) & (g2180) & (!g2205) & (!g2208) & (!g2209)) + ((!g75) & (!g2128) & (g2180) & (!g2205) & (!g2208) & (g2209)) + ((!g75) & (!g2128) & (g2180) & (!g2205) & (g2208) & (!g2209)) + ((!g75) & (!g2128) & (g2180) & (!g2205) & (g2208) & (g2209)) + ((!g75) & (g2128) & (!g2180) & (!g2205) & (!g2208) & (!g2209)) + ((!g75) & (g2128) & (!g2180) & (!g2205) & (!g2208) & (g2209)) + ((!g75) & (g2128) & (!g2180) & (!g2205) & (g2208) & (!g2209)) + ((!g75) & (g2128) & (!g2180) & (!g2205) & (g2208) & (g2209)) + ((!g75) & (g2128) & (g2180) & (!g2205) & (!g2208) & (!g2209)) + ((!g75) & (g2128) & (g2180) & (!g2205) & (!g2208) & (g2209)) + ((!g75) & (g2128) & (g2180) & (!g2205) & (g2208) & (!g2209)) + ((!g75) & (g2128) & (g2180) & (!g2205) & (g2208) & (g2209)) + ((g75) & (!g2128) & (!g2180) & (!g2205) & (g2208) & (!g2209)) + ((g75) & (!g2128) & (!g2180) & (!g2205) & (g2208) & (g2209)) + ((g75) & (!g2128) & (!g2180) & (g2205) & (g2208) & (!g2209)) + ((g75) & (!g2128) & (!g2180) & (g2205) & (g2208) & (g2209)) + ((g75) & (!g2128) & (g2180) & (!g2205) & (!g2208) & (g2209)) + ((g75) & (!g2128) & (g2180) & (!g2205) & (g2208) & (g2209)) + ((g75) & (!g2128) & (g2180) & (g2205) & (!g2208) & (g2209)) + ((g75) & (!g2128) & (g2180) & (g2205) & (g2208) & (g2209)) + ((g75) & (g2128) & (!g2180) & (!g2205) & (g2208) & (!g2209)) + ((g75) & (g2128) & (!g2180) & (!g2205) & (g2208) & (g2209)) + ((g75) & (g2128) & (!g2180) & (g2205) & (g2208) & (!g2209)) + ((g75) & (g2128) & (!g2180) & (g2205) & (g2208) & (g2209)));
	assign g2211 = (((!g2074) & (!g2071) & (!sk[53]) & (!g2070) & (g2105) & (!g2104)) + ((!g2074) & (!g2071) & (!sk[53]) & (!g2070) & (g2105) & (g2104)) + ((!g2074) & (!g2071) & (!sk[53]) & (g2070) & (!g2105) & (!g2104)) + ((!g2074) & (!g2071) & (!sk[53]) & (g2070) & (!g2105) & (g2104)) + ((!g2074) & (!g2071) & (!sk[53]) & (g2070) & (g2105) & (!g2104)) + ((!g2074) & (!g2071) & (!sk[53]) & (g2070) & (g2105) & (g2104)) + ((!g2074) & (!g2071) & (sk[53]) & (!g2070) & (g2105) & (!g2104)) + ((!g2074) & (!g2071) & (sk[53]) & (!g2070) & (g2105) & (g2104)) + ((!g2074) & (!g2071) & (sk[53]) & (g2070) & (g2105) & (!g2104)) + ((!g2074) & (!g2071) & (sk[53]) & (g2070) & (g2105) & (g2104)) + ((!g2074) & (g2071) & (!sk[53]) & (!g2070) & (!g2105) & (!g2104)) + ((!g2074) & (g2071) & (!sk[53]) & (!g2070) & (!g2105) & (g2104)) + ((!g2074) & (g2071) & (!sk[53]) & (!g2070) & (g2105) & (!g2104)) + ((!g2074) & (g2071) & (!sk[53]) & (!g2070) & (g2105) & (g2104)) + ((!g2074) & (g2071) & (!sk[53]) & (g2070) & (!g2105) & (!g2104)) + ((!g2074) & (g2071) & (!sk[53]) & (g2070) & (!g2105) & (g2104)) + ((!g2074) & (g2071) & (!sk[53]) & (g2070) & (g2105) & (!g2104)) + ((!g2074) & (g2071) & (!sk[53]) & (g2070) & (g2105) & (g2104)) + ((!g2074) & (g2071) & (sk[53]) & (!g2070) & (!g2105) & (g2104)) + ((!g2074) & (g2071) & (sk[53]) & (!g2070) & (g2105) & (g2104)) + ((!g2074) & (g2071) & (sk[53]) & (g2070) & (!g2105) & (g2104)) + ((!g2074) & (g2071) & (sk[53]) & (g2070) & (g2105) & (g2104)) + ((g2074) & (!g2071) & (!sk[53]) & (!g2070) & (g2105) & (!g2104)) + ((g2074) & (!g2071) & (!sk[53]) & (!g2070) & (g2105) & (g2104)) + ((g2074) & (!g2071) & (!sk[53]) & (g2070) & (!g2105) & (!g2104)) + ((g2074) & (!g2071) & (!sk[53]) & (g2070) & (!g2105) & (g2104)) + ((g2074) & (!g2071) & (!sk[53]) & (g2070) & (g2105) & (!g2104)) + ((g2074) & (!g2071) & (!sk[53]) & (g2070) & (g2105) & (g2104)) + ((g2074) & (!g2071) & (sk[53]) & (g2070) & (!g2105) & (!g2104)) + ((g2074) & (!g2071) & (sk[53]) & (g2070) & (!g2105) & (g2104)) + ((g2074) & (!g2071) & (sk[53]) & (g2070) & (g2105) & (!g2104)) + ((g2074) & (!g2071) & (sk[53]) & (g2070) & (g2105) & (g2104)) + ((g2074) & (g2071) & (!sk[53]) & (!g2070) & (!g2105) & (!g2104)) + ((g2074) & (g2071) & (!sk[53]) & (!g2070) & (!g2105) & (g2104)) + ((g2074) & (g2071) & (!sk[53]) & (!g2070) & (g2105) & (!g2104)) + ((g2074) & (g2071) & (!sk[53]) & (!g2070) & (g2105) & (g2104)) + ((g2074) & (g2071) & (!sk[53]) & (g2070) & (!g2105) & (!g2104)) + ((g2074) & (g2071) & (!sk[53]) & (g2070) & (!g2105) & (g2104)) + ((g2074) & (g2071) & (!sk[53]) & (g2070) & (g2105) & (!g2104)) + ((g2074) & (g2071) & (!sk[53]) & (g2070) & (g2105) & (g2104)));
	assign g2212 = (((!sk[54]) & (!g2076) & (!g2077) & (g2211)) + ((!sk[54]) & (!g2076) & (g2077) & (!g2211)) + ((!sk[54]) & (!g2076) & (g2077) & (g2211)) + ((!sk[54]) & (g2076) & (!g2077) & (g2211)) + ((!sk[54]) & (g2076) & (g2077) & (!g2211)) + ((!sk[54]) & (g2076) & (g2077) & (g2211)) + ((sk[54]) & (!g2076) & (!g2077) & (g2211)));
	assign g2213 = (((!g2074) & (!g2071) & (!g2070) & (!g2077) & (g2105) & (!g2104)) + ((!g2074) & (!g2071) & (!g2070) & (!g2077) & (g2105) & (g2104)) + ((!g2074) & (!g2071) & (!g2070) & (g2077) & (!g2105) & (!g2104)) + ((!g2074) & (!g2071) & (!g2070) & (g2077) & (!g2105) & (g2104)) + ((!g2074) & (!g2071) & (g2070) & (!g2077) & (g2105) & (!g2104)) + ((!g2074) & (!g2071) & (g2070) & (!g2077) & (g2105) & (g2104)) + ((!g2074) & (!g2071) & (g2070) & (g2077) & (!g2105) & (!g2104)) + ((!g2074) & (!g2071) & (g2070) & (g2077) & (!g2105) & (g2104)) + ((!g2074) & (g2071) & (!g2070) & (!g2077) & (g2105) & (!g2104)) + ((!g2074) & (g2071) & (!g2070) & (!g2077) & (g2105) & (g2104)) + ((!g2074) & (g2071) & (!g2070) & (g2077) & (!g2105) & (!g2104)) + ((!g2074) & (g2071) & (!g2070) & (g2077) & (!g2105) & (g2104)) + ((!g2074) & (g2071) & (g2070) & (!g2077) & (!g2105) & (g2104)) + ((!g2074) & (g2071) & (g2070) & (!g2077) & (g2105) & (!g2104)) + ((!g2074) & (g2071) & (g2070) & (g2077) & (!g2105) & (!g2104)) + ((!g2074) & (g2071) & (g2070) & (g2077) & (g2105) & (g2104)) + ((g2074) & (!g2071) & (!g2070) & (!g2077) & (!g2105) & (g2104)) + ((g2074) & (!g2071) & (!g2070) & (!g2077) & (g2105) & (!g2104)) + ((g2074) & (!g2071) & (!g2070) & (g2077) & (!g2105) & (!g2104)) + ((g2074) & (!g2071) & (!g2070) & (g2077) & (g2105) & (g2104)) + ((g2074) & (!g2071) & (g2070) & (!g2077) & (!g2105) & (g2104)) + ((g2074) & (!g2071) & (g2070) & (!g2077) & (g2105) & (!g2104)) + ((g2074) & (!g2071) & (g2070) & (g2077) & (!g2105) & (!g2104)) + ((g2074) & (!g2071) & (g2070) & (g2077) & (g2105) & (g2104)) + ((g2074) & (g2071) & (!g2070) & (!g2077) & (!g2105) & (g2104)) + ((g2074) & (g2071) & (!g2070) & (!g2077) & (g2105) & (!g2104)) + ((g2074) & (g2071) & (!g2070) & (g2077) & (!g2105) & (!g2104)) + ((g2074) & (g2071) & (!g2070) & (g2077) & (g2105) & (g2104)) + ((g2074) & (g2071) & (g2070) & (!g2077) & (!g2105) & (!g2104)) + ((g2074) & (g2071) & (g2070) & (!g2077) & (!g2105) & (g2104)) + ((g2074) & (g2071) & (g2070) & (g2077) & (g2105) & (!g2104)) + ((g2074) & (g2071) & (g2070) & (g2077) & (g2105) & (g2104)));
	assign g2214 = (((!g2072) & (!g2079) & (!g2185) & (!sk[56]) & (g2213)) + ((!g2072) & (!g2079) & (!g2185) & (sk[56]) & (g2213)) + ((!g2072) & (!g2079) & (g2185) & (!sk[56]) & (!g2213)) + ((!g2072) & (!g2079) & (g2185) & (!sk[56]) & (g2213)) + ((!g2072) & (!g2079) & (g2185) & (sk[56]) & (g2213)) + ((!g2072) & (g2079) & (!g2185) & (!sk[56]) & (!g2213)) + ((!g2072) & (g2079) & (!g2185) & (!sk[56]) & (g2213)) + ((!g2072) & (g2079) & (!g2185) & (sk[56]) & (g2213)) + ((!g2072) & (g2079) & (g2185) & (!sk[56]) & (!g2213)) + ((!g2072) & (g2079) & (g2185) & (!sk[56]) & (g2213)) + ((!g2072) & (g2079) & (g2185) & (sk[56]) & (g2213)) + ((g2072) & (!g2079) & (!g2185) & (!sk[56]) & (g2213)) + ((g2072) & (!g2079) & (!g2185) & (sk[56]) & (g2213)) + ((g2072) & (!g2079) & (g2185) & (!sk[56]) & (!g2213)) + ((g2072) & (!g2079) & (g2185) & (!sk[56]) & (g2213)) + ((g2072) & (!g2079) & (g2185) & (sk[56]) & (g2213)) + ((g2072) & (g2079) & (!g2185) & (!sk[56]) & (!g2213)) + ((g2072) & (g2079) & (!g2185) & (!sk[56]) & (g2213)) + ((g2072) & (g2079) & (!g2185) & (sk[56]) & (g2213)) + ((g2072) & (g2079) & (g2185) & (!sk[56]) & (!g2213)) + ((g2072) & (g2079) & (g2185) & (!sk[56]) & (g2213)) + ((g2072) & (g2079) & (g2185) & (sk[56]) & (!g2213)));
	assign g2215 = (((!g2085) & (!g2086) & (!g2093) & (g2094) & (g2071) & (g2074)) + ((!g2085) & (!g2086) & (g2093) & (!g2094) & (!g2071) & (g2074)) + ((!g2085) & (!g2086) & (g2093) & (g2094) & (!g2071) & (g2074)) + ((!g2085) & (!g2086) & (g2093) & (g2094) & (g2071) & (g2074)) + ((!g2085) & (g2086) & (!g2093) & (!g2094) & (g2071) & (!g2074)) + ((!g2085) & (g2086) & (!g2093) & (g2094) & (g2071) & (!g2074)) + ((!g2085) & (g2086) & (!g2093) & (g2094) & (g2071) & (g2074)) + ((!g2085) & (g2086) & (g2093) & (!g2094) & (!g2071) & (g2074)) + ((!g2085) & (g2086) & (g2093) & (!g2094) & (g2071) & (!g2074)) + ((!g2085) & (g2086) & (g2093) & (g2094) & (!g2071) & (g2074)) + ((!g2085) & (g2086) & (g2093) & (g2094) & (g2071) & (!g2074)) + ((!g2085) & (g2086) & (g2093) & (g2094) & (g2071) & (g2074)) + ((g2085) & (!g2086) & (!g2093) & (!g2094) & (!g2071) & (!g2074)) + ((g2085) & (!g2086) & (!g2093) & (g2094) & (!g2071) & (!g2074)) + ((g2085) & (!g2086) & (!g2093) & (g2094) & (g2071) & (g2074)) + ((g2085) & (!g2086) & (g2093) & (!g2094) & (!g2071) & (!g2074)) + ((g2085) & (!g2086) & (g2093) & (!g2094) & (!g2071) & (g2074)) + ((g2085) & (!g2086) & (g2093) & (g2094) & (!g2071) & (!g2074)) + ((g2085) & (!g2086) & (g2093) & (g2094) & (!g2071) & (g2074)) + ((g2085) & (!g2086) & (g2093) & (g2094) & (g2071) & (g2074)) + ((g2085) & (g2086) & (!g2093) & (!g2094) & (!g2071) & (!g2074)) + ((g2085) & (g2086) & (!g2093) & (!g2094) & (g2071) & (!g2074)) + ((g2085) & (g2086) & (!g2093) & (g2094) & (!g2071) & (!g2074)) + ((g2085) & (g2086) & (!g2093) & (g2094) & (g2071) & (!g2074)) + ((g2085) & (g2086) & (!g2093) & (g2094) & (g2071) & (g2074)) + ((g2085) & (g2086) & (g2093) & (!g2094) & (!g2071) & (!g2074)) + ((g2085) & (g2086) & (g2093) & (!g2094) & (!g2071) & (g2074)) + ((g2085) & (g2086) & (g2093) & (!g2094) & (g2071) & (!g2074)) + ((g2085) & (g2086) & (g2093) & (g2094) & (!g2071) & (!g2074)) + ((g2085) & (g2086) & (g2093) & (g2094) & (!g2071) & (g2074)) + ((g2085) & (g2086) & (g2093) & (g2094) & (g2071) & (!g2074)) + ((g2085) & (g2086) & (g2093) & (g2094) & (g2071) & (g2074)));
	assign g2216 = (((!g2090) & (!g2091) & (!g2098) & (g2099) & (g2071) & (g2074)) + ((!g2090) & (!g2091) & (g2098) & (!g2099) & (!g2071) & (g2074)) + ((!g2090) & (!g2091) & (g2098) & (g2099) & (!g2071) & (g2074)) + ((!g2090) & (!g2091) & (g2098) & (g2099) & (g2071) & (g2074)) + ((!g2090) & (g2091) & (!g2098) & (!g2099) & (g2071) & (!g2074)) + ((!g2090) & (g2091) & (!g2098) & (g2099) & (g2071) & (!g2074)) + ((!g2090) & (g2091) & (!g2098) & (g2099) & (g2071) & (g2074)) + ((!g2090) & (g2091) & (g2098) & (!g2099) & (!g2071) & (g2074)) + ((!g2090) & (g2091) & (g2098) & (!g2099) & (g2071) & (!g2074)) + ((!g2090) & (g2091) & (g2098) & (g2099) & (!g2071) & (g2074)) + ((!g2090) & (g2091) & (g2098) & (g2099) & (g2071) & (!g2074)) + ((!g2090) & (g2091) & (g2098) & (g2099) & (g2071) & (g2074)) + ((g2090) & (!g2091) & (!g2098) & (!g2099) & (!g2071) & (!g2074)) + ((g2090) & (!g2091) & (!g2098) & (g2099) & (!g2071) & (!g2074)) + ((g2090) & (!g2091) & (!g2098) & (g2099) & (g2071) & (g2074)) + ((g2090) & (!g2091) & (g2098) & (!g2099) & (!g2071) & (!g2074)) + ((g2090) & (!g2091) & (g2098) & (!g2099) & (!g2071) & (g2074)) + ((g2090) & (!g2091) & (g2098) & (g2099) & (!g2071) & (!g2074)) + ((g2090) & (!g2091) & (g2098) & (g2099) & (!g2071) & (g2074)) + ((g2090) & (!g2091) & (g2098) & (g2099) & (g2071) & (g2074)) + ((g2090) & (g2091) & (!g2098) & (!g2099) & (!g2071) & (!g2074)) + ((g2090) & (g2091) & (!g2098) & (!g2099) & (g2071) & (!g2074)) + ((g2090) & (g2091) & (!g2098) & (g2099) & (!g2071) & (!g2074)) + ((g2090) & (g2091) & (!g2098) & (g2099) & (g2071) & (!g2074)) + ((g2090) & (g2091) & (!g2098) & (g2099) & (g2071) & (g2074)) + ((g2090) & (g2091) & (g2098) & (!g2099) & (!g2071) & (!g2074)) + ((g2090) & (g2091) & (g2098) & (!g2099) & (!g2071) & (g2074)) + ((g2090) & (g2091) & (g2098) & (!g2099) & (g2071) & (!g2074)) + ((g2090) & (g2091) & (g2098) & (g2099) & (!g2071) & (!g2074)) + ((g2090) & (g2091) & (g2098) & (g2099) & (!g2071) & (g2074)) + ((g2090) & (g2091) & (g2098) & (g2099) & (g2071) & (!g2074)) + ((g2090) & (g2091) & (g2098) & (g2099) & (g2071) & (g2074)));
	assign g2217 = (((!g2095) & (!g2096) & (!g2088) & (g2089) & (g2071) & (g2074)) + ((!g2095) & (!g2096) & (g2088) & (!g2089) & (!g2071) & (g2074)) + ((!g2095) & (!g2096) & (g2088) & (g2089) & (!g2071) & (g2074)) + ((!g2095) & (!g2096) & (g2088) & (g2089) & (g2071) & (g2074)) + ((!g2095) & (g2096) & (!g2088) & (!g2089) & (g2071) & (!g2074)) + ((!g2095) & (g2096) & (!g2088) & (g2089) & (g2071) & (!g2074)) + ((!g2095) & (g2096) & (!g2088) & (g2089) & (g2071) & (g2074)) + ((!g2095) & (g2096) & (g2088) & (!g2089) & (!g2071) & (g2074)) + ((!g2095) & (g2096) & (g2088) & (!g2089) & (g2071) & (!g2074)) + ((!g2095) & (g2096) & (g2088) & (g2089) & (!g2071) & (g2074)) + ((!g2095) & (g2096) & (g2088) & (g2089) & (g2071) & (!g2074)) + ((!g2095) & (g2096) & (g2088) & (g2089) & (g2071) & (g2074)) + ((g2095) & (!g2096) & (!g2088) & (!g2089) & (!g2071) & (!g2074)) + ((g2095) & (!g2096) & (!g2088) & (g2089) & (!g2071) & (!g2074)) + ((g2095) & (!g2096) & (!g2088) & (g2089) & (g2071) & (g2074)) + ((g2095) & (!g2096) & (g2088) & (!g2089) & (!g2071) & (!g2074)) + ((g2095) & (!g2096) & (g2088) & (!g2089) & (!g2071) & (g2074)) + ((g2095) & (!g2096) & (g2088) & (g2089) & (!g2071) & (!g2074)) + ((g2095) & (!g2096) & (g2088) & (g2089) & (!g2071) & (g2074)) + ((g2095) & (!g2096) & (g2088) & (g2089) & (g2071) & (g2074)) + ((g2095) & (g2096) & (!g2088) & (!g2089) & (!g2071) & (!g2074)) + ((g2095) & (g2096) & (!g2088) & (!g2089) & (g2071) & (!g2074)) + ((g2095) & (g2096) & (!g2088) & (g2089) & (!g2071) & (!g2074)) + ((g2095) & (g2096) & (!g2088) & (g2089) & (g2071) & (!g2074)) + ((g2095) & (g2096) & (!g2088) & (g2089) & (g2071) & (g2074)) + ((g2095) & (g2096) & (g2088) & (!g2089) & (!g2071) & (!g2074)) + ((g2095) & (g2096) & (g2088) & (!g2089) & (!g2071) & (g2074)) + ((g2095) & (g2096) & (g2088) & (!g2089) & (g2071) & (!g2074)) + ((g2095) & (g2096) & (g2088) & (g2089) & (!g2071) & (!g2074)) + ((g2095) & (g2096) & (g2088) & (g2089) & (!g2071) & (g2074)) + ((g2095) & (g2096) & (g2088) & (g2089) & (g2071) & (!g2074)) + ((g2095) & (g2096) & (g2088) & (g2089) & (g2071) & (g2074)));
	assign g2218 = (((!g2074) & (!g2071) & (!g2100) & (!sk[60]) & (g2101) & (!g2192)) + ((!g2074) & (!g2071) & (!g2100) & (!sk[60]) & (g2101) & (g2192)) + ((!g2074) & (!g2071) & (g2100) & (!sk[60]) & (!g2101) & (!g2192)) + ((!g2074) & (!g2071) & (g2100) & (!sk[60]) & (!g2101) & (g2192)) + ((!g2074) & (!g2071) & (g2100) & (!sk[60]) & (g2101) & (!g2192)) + ((!g2074) & (!g2071) & (g2100) & (!sk[60]) & (g2101) & (g2192)) + ((!g2074) & (!g2071) & (g2100) & (sk[60]) & (!g2101) & (!g2192)) + ((!g2074) & (!g2071) & (g2100) & (sk[60]) & (!g2101) & (g2192)) + ((!g2074) & (!g2071) & (g2100) & (sk[60]) & (g2101) & (!g2192)) + ((!g2074) & (!g2071) & (g2100) & (sk[60]) & (g2101) & (g2192)) + ((!g2074) & (g2071) & (!g2100) & (!sk[60]) & (!g2101) & (!g2192)) + ((!g2074) & (g2071) & (!g2100) & (!sk[60]) & (!g2101) & (g2192)) + ((!g2074) & (g2071) & (!g2100) & (!sk[60]) & (g2101) & (!g2192)) + ((!g2074) & (g2071) & (!g2100) & (!sk[60]) & (g2101) & (g2192)) + ((!g2074) & (g2071) & (!g2100) & (sk[60]) & (g2101) & (!g2192)) + ((!g2074) & (g2071) & (!g2100) & (sk[60]) & (g2101) & (g2192)) + ((!g2074) & (g2071) & (g2100) & (!sk[60]) & (!g2101) & (!g2192)) + ((!g2074) & (g2071) & (g2100) & (!sk[60]) & (!g2101) & (g2192)) + ((!g2074) & (g2071) & (g2100) & (!sk[60]) & (g2101) & (!g2192)) + ((!g2074) & (g2071) & (g2100) & (!sk[60]) & (g2101) & (g2192)) + ((!g2074) & (g2071) & (g2100) & (sk[60]) & (g2101) & (!g2192)) + ((!g2074) & (g2071) & (g2100) & (sk[60]) & (g2101) & (g2192)) + ((g2074) & (!g2071) & (!g2100) & (!sk[60]) & (g2101) & (!g2192)) + ((g2074) & (!g2071) & (!g2100) & (!sk[60]) & (g2101) & (g2192)) + ((g2074) & (!g2071) & (!g2100) & (sk[60]) & (!g2101) & (g2192)) + ((g2074) & (!g2071) & (!g2100) & (sk[60]) & (g2101) & (g2192)) + ((g2074) & (!g2071) & (g2100) & (!sk[60]) & (!g2101) & (!g2192)) + ((g2074) & (!g2071) & (g2100) & (!sk[60]) & (!g2101) & (g2192)) + ((g2074) & (!g2071) & (g2100) & (!sk[60]) & (g2101) & (!g2192)) + ((g2074) & (!g2071) & (g2100) & (!sk[60]) & (g2101) & (g2192)) + ((g2074) & (!g2071) & (g2100) & (sk[60]) & (!g2101) & (g2192)) + ((g2074) & (!g2071) & (g2100) & (sk[60]) & (g2101) & (g2192)) + ((g2074) & (g2071) & (!g2100) & (!sk[60]) & (!g2101) & (!g2192)) + ((g2074) & (g2071) & (!g2100) & (!sk[60]) & (!g2101) & (g2192)) + ((g2074) & (g2071) & (!g2100) & (!sk[60]) & (g2101) & (!g2192)) + ((g2074) & (g2071) & (!g2100) & (!sk[60]) & (g2101) & (g2192)) + ((g2074) & (g2071) & (!g2100) & (sk[60]) & (!g2101) & (g2192)) + ((g2074) & (g2071) & (!g2100) & (sk[60]) & (g2101) & (g2192)) + ((g2074) & (g2071) & (g2100) & (!sk[60]) & (!g2101) & (!g2192)) + ((g2074) & (g2071) & (g2100) & (!sk[60]) & (!g2101) & (g2192)) + ((g2074) & (g2071) & (g2100) & (!sk[60]) & (g2101) & (!g2192)) + ((g2074) & (g2071) & (g2100) & (!sk[60]) & (g2101) & (g2192)) + ((g2074) & (g2071) & (g2100) & (sk[60]) & (!g2101) & (g2192)) + ((g2074) & (g2071) & (g2100) & (sk[60]) & (g2101) & (g2192)));
	assign g2219 = (((!g2215) & (!g2216) & (!g2217) & (g2218) & (g2076) & (g2077)) + ((!g2215) & (!g2216) & (g2217) & (!g2218) & (!g2076) & (g2077)) + ((!g2215) & (!g2216) & (g2217) & (g2218) & (!g2076) & (g2077)) + ((!g2215) & (!g2216) & (g2217) & (g2218) & (g2076) & (g2077)) + ((!g2215) & (g2216) & (!g2217) & (!g2218) & (g2076) & (!g2077)) + ((!g2215) & (g2216) & (!g2217) & (g2218) & (g2076) & (!g2077)) + ((!g2215) & (g2216) & (!g2217) & (g2218) & (g2076) & (g2077)) + ((!g2215) & (g2216) & (g2217) & (!g2218) & (!g2076) & (g2077)) + ((!g2215) & (g2216) & (g2217) & (!g2218) & (g2076) & (!g2077)) + ((!g2215) & (g2216) & (g2217) & (g2218) & (!g2076) & (g2077)) + ((!g2215) & (g2216) & (g2217) & (g2218) & (g2076) & (!g2077)) + ((!g2215) & (g2216) & (g2217) & (g2218) & (g2076) & (g2077)) + ((g2215) & (!g2216) & (!g2217) & (!g2218) & (!g2076) & (!g2077)) + ((g2215) & (!g2216) & (!g2217) & (g2218) & (!g2076) & (!g2077)) + ((g2215) & (!g2216) & (!g2217) & (g2218) & (g2076) & (g2077)) + ((g2215) & (!g2216) & (g2217) & (!g2218) & (!g2076) & (!g2077)) + ((g2215) & (!g2216) & (g2217) & (!g2218) & (!g2076) & (g2077)) + ((g2215) & (!g2216) & (g2217) & (g2218) & (!g2076) & (!g2077)) + ((g2215) & (!g2216) & (g2217) & (g2218) & (!g2076) & (g2077)) + ((g2215) & (!g2216) & (g2217) & (g2218) & (g2076) & (g2077)) + ((g2215) & (g2216) & (!g2217) & (!g2218) & (!g2076) & (!g2077)) + ((g2215) & (g2216) & (!g2217) & (!g2218) & (g2076) & (!g2077)) + ((g2215) & (g2216) & (!g2217) & (g2218) & (!g2076) & (!g2077)) + ((g2215) & (g2216) & (!g2217) & (g2218) & (g2076) & (!g2077)) + ((g2215) & (g2216) & (!g2217) & (g2218) & (g2076) & (g2077)) + ((g2215) & (g2216) & (g2217) & (!g2218) & (!g2076) & (!g2077)) + ((g2215) & (g2216) & (g2217) & (!g2218) & (!g2076) & (g2077)) + ((g2215) & (g2216) & (g2217) & (!g2218) & (g2076) & (!g2077)) + ((g2215) & (g2216) & (g2217) & (g2218) & (!g2076) & (!g2077)) + ((g2215) & (g2216) & (g2217) & (g2218) & (!g2076) & (g2077)) + ((g2215) & (g2216) & (g2217) & (g2218) & (g2076) & (!g2077)) + ((g2215) & (g2216) & (g2217) & (g2218) & (g2076) & (g2077)));
	assign g2220 = (((!g2115) & (!g2116) & (!g2108) & (g2109) & (g2071) & (g2074)) + ((!g2115) & (!g2116) & (g2108) & (!g2109) & (!g2071) & (g2074)) + ((!g2115) & (!g2116) & (g2108) & (g2109) & (!g2071) & (g2074)) + ((!g2115) & (!g2116) & (g2108) & (g2109) & (g2071) & (g2074)) + ((!g2115) & (g2116) & (!g2108) & (!g2109) & (g2071) & (!g2074)) + ((!g2115) & (g2116) & (!g2108) & (g2109) & (g2071) & (!g2074)) + ((!g2115) & (g2116) & (!g2108) & (g2109) & (g2071) & (g2074)) + ((!g2115) & (g2116) & (g2108) & (!g2109) & (!g2071) & (g2074)) + ((!g2115) & (g2116) & (g2108) & (!g2109) & (g2071) & (!g2074)) + ((!g2115) & (g2116) & (g2108) & (g2109) & (!g2071) & (g2074)) + ((!g2115) & (g2116) & (g2108) & (g2109) & (g2071) & (!g2074)) + ((!g2115) & (g2116) & (g2108) & (g2109) & (g2071) & (g2074)) + ((g2115) & (!g2116) & (!g2108) & (!g2109) & (!g2071) & (!g2074)) + ((g2115) & (!g2116) & (!g2108) & (g2109) & (!g2071) & (!g2074)) + ((g2115) & (!g2116) & (!g2108) & (g2109) & (g2071) & (g2074)) + ((g2115) & (!g2116) & (g2108) & (!g2109) & (!g2071) & (!g2074)) + ((g2115) & (!g2116) & (g2108) & (!g2109) & (!g2071) & (g2074)) + ((g2115) & (!g2116) & (g2108) & (g2109) & (!g2071) & (!g2074)) + ((g2115) & (!g2116) & (g2108) & (g2109) & (!g2071) & (g2074)) + ((g2115) & (!g2116) & (g2108) & (g2109) & (g2071) & (g2074)) + ((g2115) & (g2116) & (!g2108) & (!g2109) & (!g2071) & (!g2074)) + ((g2115) & (g2116) & (!g2108) & (!g2109) & (g2071) & (!g2074)) + ((g2115) & (g2116) & (!g2108) & (g2109) & (!g2071) & (!g2074)) + ((g2115) & (g2116) & (!g2108) & (g2109) & (g2071) & (!g2074)) + ((g2115) & (g2116) & (!g2108) & (g2109) & (g2071) & (g2074)) + ((g2115) & (g2116) & (g2108) & (!g2109) & (!g2071) & (!g2074)) + ((g2115) & (g2116) & (g2108) & (!g2109) & (!g2071) & (g2074)) + ((g2115) & (g2116) & (g2108) & (!g2109) & (g2071) & (!g2074)) + ((g2115) & (g2116) & (g2108) & (g2109) & (!g2071) & (!g2074)) + ((g2115) & (g2116) & (g2108) & (g2109) & (!g2071) & (g2074)) + ((g2115) & (g2116) & (g2108) & (g2109) & (g2071) & (!g2074)) + ((g2115) & (g2116) & (g2108) & (g2109) & (g2071) & (g2074)));
	assign g2221 = (((!g2220) & (!g2106) & (!g2113) & (g2114) & (g2196) & (g2197)) + ((!g2220) & (!g2106) & (g2113) & (!g2114) & (!g2196) & (g2197)) + ((!g2220) & (!g2106) & (g2113) & (g2114) & (!g2196) & (g2197)) + ((!g2220) & (!g2106) & (g2113) & (g2114) & (g2196) & (g2197)) + ((!g2220) & (g2106) & (!g2113) & (!g2114) & (g2196) & (!g2197)) + ((!g2220) & (g2106) & (!g2113) & (g2114) & (g2196) & (!g2197)) + ((!g2220) & (g2106) & (!g2113) & (g2114) & (g2196) & (g2197)) + ((!g2220) & (g2106) & (g2113) & (!g2114) & (!g2196) & (g2197)) + ((!g2220) & (g2106) & (g2113) & (!g2114) & (g2196) & (!g2197)) + ((!g2220) & (g2106) & (g2113) & (g2114) & (!g2196) & (g2197)) + ((!g2220) & (g2106) & (g2113) & (g2114) & (g2196) & (!g2197)) + ((!g2220) & (g2106) & (g2113) & (g2114) & (g2196) & (g2197)) + ((g2220) & (!g2106) & (!g2113) & (!g2114) & (!g2196) & (!g2197)) + ((g2220) & (!g2106) & (!g2113) & (g2114) & (!g2196) & (!g2197)) + ((g2220) & (!g2106) & (!g2113) & (g2114) & (g2196) & (g2197)) + ((g2220) & (!g2106) & (g2113) & (!g2114) & (!g2196) & (!g2197)) + ((g2220) & (!g2106) & (g2113) & (!g2114) & (!g2196) & (g2197)) + ((g2220) & (!g2106) & (g2113) & (g2114) & (!g2196) & (!g2197)) + ((g2220) & (!g2106) & (g2113) & (g2114) & (!g2196) & (g2197)) + ((g2220) & (!g2106) & (g2113) & (g2114) & (g2196) & (g2197)) + ((g2220) & (g2106) & (!g2113) & (!g2114) & (!g2196) & (!g2197)) + ((g2220) & (g2106) & (!g2113) & (!g2114) & (g2196) & (!g2197)) + ((g2220) & (g2106) & (!g2113) & (g2114) & (!g2196) & (!g2197)) + ((g2220) & (g2106) & (!g2113) & (g2114) & (g2196) & (!g2197)) + ((g2220) & (g2106) & (!g2113) & (g2114) & (g2196) & (g2197)) + ((g2220) & (g2106) & (g2113) & (!g2114) & (!g2196) & (!g2197)) + ((g2220) & (g2106) & (g2113) & (!g2114) & (!g2196) & (g2197)) + ((g2220) & (g2106) & (g2113) & (!g2114) & (g2196) & (!g2197)) + ((g2220) & (g2106) & (g2113) & (g2114) & (!g2196) & (!g2197)) + ((g2220) & (g2106) & (g2113) & (g2114) & (!g2196) & (g2197)) + ((g2220) & (g2106) & (g2113) & (g2114) & (g2196) & (!g2197)) + ((g2220) & (g2106) & (g2113) & (g2114) & (g2196) & (g2197)));
	assign g2222 = (((!g2110) & (!g2111) & (!g2118) & (g2119) & (g2071) & (g2074)) + ((!g2110) & (!g2111) & (g2118) & (!g2119) & (!g2071) & (g2074)) + ((!g2110) & (!g2111) & (g2118) & (g2119) & (!g2071) & (g2074)) + ((!g2110) & (!g2111) & (g2118) & (g2119) & (g2071) & (g2074)) + ((!g2110) & (g2111) & (!g2118) & (!g2119) & (g2071) & (!g2074)) + ((!g2110) & (g2111) & (!g2118) & (g2119) & (g2071) & (!g2074)) + ((!g2110) & (g2111) & (!g2118) & (g2119) & (g2071) & (g2074)) + ((!g2110) & (g2111) & (g2118) & (!g2119) & (!g2071) & (g2074)) + ((!g2110) & (g2111) & (g2118) & (!g2119) & (g2071) & (!g2074)) + ((!g2110) & (g2111) & (g2118) & (g2119) & (!g2071) & (g2074)) + ((!g2110) & (g2111) & (g2118) & (g2119) & (g2071) & (!g2074)) + ((!g2110) & (g2111) & (g2118) & (g2119) & (g2071) & (g2074)) + ((g2110) & (!g2111) & (!g2118) & (!g2119) & (!g2071) & (!g2074)) + ((g2110) & (!g2111) & (!g2118) & (g2119) & (!g2071) & (!g2074)) + ((g2110) & (!g2111) & (!g2118) & (g2119) & (g2071) & (g2074)) + ((g2110) & (!g2111) & (g2118) & (!g2119) & (!g2071) & (!g2074)) + ((g2110) & (!g2111) & (g2118) & (!g2119) & (!g2071) & (g2074)) + ((g2110) & (!g2111) & (g2118) & (g2119) & (!g2071) & (!g2074)) + ((g2110) & (!g2111) & (g2118) & (g2119) & (!g2071) & (g2074)) + ((g2110) & (!g2111) & (g2118) & (g2119) & (g2071) & (g2074)) + ((g2110) & (g2111) & (!g2118) & (!g2119) & (!g2071) & (!g2074)) + ((g2110) & (g2111) & (!g2118) & (!g2119) & (g2071) & (!g2074)) + ((g2110) & (g2111) & (!g2118) & (g2119) & (!g2071) & (!g2074)) + ((g2110) & (g2111) & (!g2118) & (g2119) & (g2071) & (!g2074)) + ((g2110) & (g2111) & (!g2118) & (g2119) & (g2071) & (g2074)) + ((g2110) & (g2111) & (g2118) & (!g2119) & (!g2071) & (!g2074)) + ((g2110) & (g2111) & (g2118) & (!g2119) & (!g2071) & (g2074)) + ((g2110) & (g2111) & (g2118) & (!g2119) & (g2071) & (!g2074)) + ((g2110) & (g2111) & (g2118) & (g2119) & (!g2071) & (!g2074)) + ((g2110) & (g2111) & (g2118) & (g2119) & (!g2071) & (g2074)) + ((g2110) & (g2111) & (g2118) & (g2119) & (g2071) & (!g2074)) + ((g2110) & (g2111) & (g2118) & (g2119) & (g2071) & (g2074)));
	assign g2223 = (((!g2120) & (!g2121) & (!g2083) & (g2084) & (g2071) & (g2074)) + ((!g2120) & (!g2121) & (g2083) & (!g2084) & (!g2071) & (g2074)) + ((!g2120) & (!g2121) & (g2083) & (g2084) & (!g2071) & (g2074)) + ((!g2120) & (!g2121) & (g2083) & (g2084) & (g2071) & (g2074)) + ((!g2120) & (g2121) & (!g2083) & (!g2084) & (g2071) & (!g2074)) + ((!g2120) & (g2121) & (!g2083) & (g2084) & (g2071) & (!g2074)) + ((!g2120) & (g2121) & (!g2083) & (g2084) & (g2071) & (g2074)) + ((!g2120) & (g2121) & (g2083) & (!g2084) & (!g2071) & (g2074)) + ((!g2120) & (g2121) & (g2083) & (!g2084) & (g2071) & (!g2074)) + ((!g2120) & (g2121) & (g2083) & (g2084) & (!g2071) & (g2074)) + ((!g2120) & (g2121) & (g2083) & (g2084) & (g2071) & (!g2074)) + ((!g2120) & (g2121) & (g2083) & (g2084) & (g2071) & (g2074)) + ((g2120) & (!g2121) & (!g2083) & (!g2084) & (!g2071) & (!g2074)) + ((g2120) & (!g2121) & (!g2083) & (g2084) & (!g2071) & (!g2074)) + ((g2120) & (!g2121) & (!g2083) & (g2084) & (g2071) & (g2074)) + ((g2120) & (!g2121) & (g2083) & (!g2084) & (!g2071) & (!g2074)) + ((g2120) & (!g2121) & (g2083) & (!g2084) & (!g2071) & (g2074)) + ((g2120) & (!g2121) & (g2083) & (g2084) & (!g2071) & (!g2074)) + ((g2120) & (!g2121) & (g2083) & (g2084) & (!g2071) & (g2074)) + ((g2120) & (!g2121) & (g2083) & (g2084) & (g2071) & (g2074)) + ((g2120) & (g2121) & (!g2083) & (!g2084) & (!g2071) & (!g2074)) + ((g2120) & (g2121) & (!g2083) & (!g2084) & (g2071) & (!g2074)) + ((g2120) & (g2121) & (!g2083) & (g2084) & (!g2071) & (!g2074)) + ((g2120) & (g2121) & (!g2083) & (g2084) & (g2071) & (!g2074)) + ((g2120) & (g2121) & (!g2083) & (g2084) & (g2071) & (g2074)) + ((g2120) & (g2121) & (g2083) & (!g2084) & (!g2071) & (!g2074)) + ((g2120) & (g2121) & (g2083) & (!g2084) & (!g2071) & (g2074)) + ((g2120) & (g2121) & (g2083) & (!g2084) & (g2071) & (!g2074)) + ((g2120) & (g2121) & (g2083) & (g2084) & (!g2071) & (!g2074)) + ((g2120) & (g2121) & (g2083) & (g2084) & (!g2071) & (g2074)) + ((g2120) & (g2121) & (g2083) & (g2084) & (g2071) & (!g2074)) + ((g2120) & (g2121) & (g2083) & (g2084) & (g2071) & (g2074)));
	assign g2224 = (((!g2219) & (!g2221) & (!g2222) & (g2223) & (g2201) & (g2202)) + ((!g2219) & (!g2221) & (g2222) & (!g2223) & (!g2201) & (g2202)) + ((!g2219) & (!g2221) & (g2222) & (g2223) & (!g2201) & (g2202)) + ((!g2219) & (!g2221) & (g2222) & (g2223) & (g2201) & (g2202)) + ((!g2219) & (g2221) & (!g2222) & (!g2223) & (g2201) & (!g2202)) + ((!g2219) & (g2221) & (!g2222) & (g2223) & (g2201) & (!g2202)) + ((!g2219) & (g2221) & (!g2222) & (g2223) & (g2201) & (g2202)) + ((!g2219) & (g2221) & (g2222) & (!g2223) & (!g2201) & (g2202)) + ((!g2219) & (g2221) & (g2222) & (!g2223) & (g2201) & (!g2202)) + ((!g2219) & (g2221) & (g2222) & (g2223) & (!g2201) & (g2202)) + ((!g2219) & (g2221) & (g2222) & (g2223) & (g2201) & (!g2202)) + ((!g2219) & (g2221) & (g2222) & (g2223) & (g2201) & (g2202)) + ((g2219) & (!g2221) & (!g2222) & (!g2223) & (!g2201) & (!g2202)) + ((g2219) & (!g2221) & (!g2222) & (g2223) & (!g2201) & (!g2202)) + ((g2219) & (!g2221) & (!g2222) & (g2223) & (g2201) & (g2202)) + ((g2219) & (!g2221) & (g2222) & (!g2223) & (!g2201) & (!g2202)) + ((g2219) & (!g2221) & (g2222) & (!g2223) & (!g2201) & (g2202)) + ((g2219) & (!g2221) & (g2222) & (g2223) & (!g2201) & (!g2202)) + ((g2219) & (!g2221) & (g2222) & (g2223) & (!g2201) & (g2202)) + ((g2219) & (!g2221) & (g2222) & (g2223) & (g2201) & (g2202)) + ((g2219) & (g2221) & (!g2222) & (!g2223) & (!g2201) & (!g2202)) + ((g2219) & (g2221) & (!g2222) & (!g2223) & (g2201) & (!g2202)) + ((g2219) & (g2221) & (!g2222) & (g2223) & (!g2201) & (!g2202)) + ((g2219) & (g2221) & (!g2222) & (g2223) & (g2201) & (!g2202)) + ((g2219) & (g2221) & (!g2222) & (g2223) & (g2201) & (g2202)) + ((g2219) & (g2221) & (g2222) & (!g2223) & (!g2201) & (!g2202)) + ((g2219) & (g2221) & (g2222) & (!g2223) & (!g2201) & (g2202)) + ((g2219) & (g2221) & (g2222) & (!g2223) & (g2201) & (!g2202)) + ((g2219) & (g2221) & (g2222) & (g2223) & (!g2201) & (!g2202)) + ((g2219) & (g2221) & (g2222) & (g2223) & (!g2201) & (g2202)) + ((g2219) & (g2221) & (g2222) & (g2223) & (g2201) & (!g2202)) + ((g2219) & (g2221) & (g2222) & (g2223) & (g2201) & (g2202)));
	assign g2225 = (((!g2073) & (!g2080) & (!g2125) & (g2212) & (!g3764) & (!g2224)) + ((!g2073) & (!g2080) & (!g2125) & (g2212) & (!g3764) & (g2224)) + ((!g2073) & (!g2080) & (!g2125) & (g2212) & (g3764) & (!g2224)) + ((!g2073) & (!g2080) & (!g2125) & (g2212) & (g3764) & (g2224)) + ((!g2073) & (!g2080) & (g2125) & (!g2212) & (!g3764) & (g2224)) + ((!g2073) & (!g2080) & (g2125) & (!g2212) & (g3764) & (g2224)) + ((!g2073) & (!g2080) & (g2125) & (g2212) & (!g3764) & (g2224)) + ((!g2073) & (!g2080) & (g2125) & (g2212) & (g3764) & (g2224)) + ((!g2073) & (g2080) & (!g2125) & (!g2212) & (g3764) & (!g2224)) + ((!g2073) & (g2080) & (!g2125) & (!g2212) & (g3764) & (g2224)) + ((!g2073) & (g2080) & (!g2125) & (g2212) & (g3764) & (!g2224)) + ((!g2073) & (g2080) & (!g2125) & (g2212) & (g3764) & (g2224)) + ((!g2073) & (g2080) & (g2125) & (!g2212) & (g3764) & (!g2224)) + ((!g2073) & (g2080) & (g2125) & (!g2212) & (g3764) & (g2224)) + ((!g2073) & (g2080) & (g2125) & (g2212) & (g3764) & (!g2224)) + ((!g2073) & (g2080) & (g2125) & (g2212) & (g3764) & (g2224)) + ((g2073) & (!g2080) & (g2125) & (!g2212) & (!g3764) & (g2224)) + ((g2073) & (!g2080) & (g2125) & (!g2212) & (g3764) & (g2224)) + ((g2073) & (!g2080) & (g2125) & (g2212) & (!g3764) & (g2224)) + ((g2073) & (!g2080) & (g2125) & (g2212) & (g3764) & (g2224)) + ((g2073) & (g2080) & (!g2125) & (!g2212) & (g3764) & (!g2224)) + ((g2073) & (g2080) & (!g2125) & (!g2212) & (g3764) & (g2224)) + ((g2073) & (g2080) & (!g2125) & (g2212) & (g3764) & (!g2224)) + ((g2073) & (g2080) & (!g2125) & (g2212) & (g3764) & (g2224)) + ((g2073) & (g2080) & (g2125) & (!g2212) & (g3764) & (!g2224)) + ((g2073) & (g2080) & (g2125) & (!g2212) & (g3764) & (g2224)) + ((g2073) & (g2080) & (g2125) & (g2212) & (g3764) & (!g2224)) + ((g2073) & (g2080) & (g2125) & (g2212) & (g3764) & (g2224)));
	assign g2226 = (((!g2081) & (!g2124) & (!g2182) & (!g2077) & (!g2225) & (!g2105)) + ((!g2081) & (!g2124) & (!g2182) & (!g2077) & (!g2225) & (g2105)) + ((!g2081) & (!g2124) & (!g2182) & (g2077) & (!g2225) & (!g2105)) + ((!g2081) & (!g2124) & (!g2182) & (g2077) & (!g2225) & (g2105)) + ((!g2081) & (!g2124) & (g2182) & (!g2077) & (!g2225) & (!g2105)) + ((!g2081) & (!g2124) & (g2182) & (!g2077) & (g2225) & (!g2105)) + ((!g2081) & (!g2124) & (g2182) & (g2077) & (!g2225) & (!g2105)) + ((!g2081) & (!g2124) & (g2182) & (g2077) & (g2225) & (!g2105)) + ((!g2081) & (g2124) & (!g2182) & (!g2077) & (!g2225) & (!g2105)) + ((!g2081) & (g2124) & (!g2182) & (!g2077) & (g2225) & (!g2105)) + ((!g2081) & (g2124) & (g2182) & (!g2077) & (!g2225) & (!g2105)) + ((!g2081) & (g2124) & (g2182) & (!g2077) & (g2225) & (!g2105)) + ((!g2081) & (g2124) & (g2182) & (g2077) & (!g2225) & (!g2105)) + ((!g2081) & (g2124) & (g2182) & (g2077) & (g2225) & (!g2105)) + ((g2081) & (!g2124) & (!g2182) & (!g2077) & (!g2225) & (!g2105)) + ((g2081) & (!g2124) & (!g2182) & (!g2077) & (!g2225) & (g2105)) + ((g2081) & (!g2124) & (!g2182) & (g2077) & (!g2225) & (!g2105)) + ((g2081) & (!g2124) & (!g2182) & (g2077) & (!g2225) & (g2105)) + ((g2081) & (!g2124) & (g2182) & (!g2077) & (!g2225) & (!g2105)) + ((g2081) & (!g2124) & (g2182) & (!g2077) & (g2225) & (!g2105)) + ((g2081) & (!g2124) & (g2182) & (g2077) & (!g2225) & (!g2105)) + ((g2081) & (!g2124) & (g2182) & (g2077) & (g2225) & (!g2105)) + ((g2081) & (g2124) & (!g2182) & (!g2077) & (!g2225) & (!g2105)) + ((g2081) & (g2124) & (!g2182) & (!g2077) & (g2225) & (!g2105)) + ((g2081) & (g2124) & (!g2182) & (g2077) & (!g2225) & (g2105)) + ((g2081) & (g2124) & (!g2182) & (g2077) & (g2225) & (g2105)) + ((g2081) & (g2124) & (g2182) & (!g2077) & (!g2225) & (!g2105)) + ((g2081) & (g2124) & (g2182) & (!g2077) & (g2225) & (!g2105)) + ((g2081) & (g2124) & (g2182) & (g2077) & (!g2225) & (!g2105)) + ((g2081) & (g2124) & (g2182) & (g2077) & (g2225) & (!g2105)));
	assign g2227 = (((!dmem_dat_ix2x) & (!dmem_dat_ix10x) & (!dmem_dat_ix26x) & (dmem_dat_ix18x) & (g2206) & (g2207)) + ((!dmem_dat_ix2x) & (!dmem_dat_ix10x) & (dmem_dat_ix26x) & (!dmem_dat_ix18x) & (!g2206) & (g2207)) + ((!dmem_dat_ix2x) & (!dmem_dat_ix10x) & (dmem_dat_ix26x) & (dmem_dat_ix18x) & (!g2206) & (g2207)) + ((!dmem_dat_ix2x) & (!dmem_dat_ix10x) & (dmem_dat_ix26x) & (dmem_dat_ix18x) & (g2206) & (g2207)) + ((!dmem_dat_ix2x) & (dmem_dat_ix10x) & (!dmem_dat_ix26x) & (!dmem_dat_ix18x) & (g2206) & (!g2207)) + ((!dmem_dat_ix2x) & (dmem_dat_ix10x) & (!dmem_dat_ix26x) & (dmem_dat_ix18x) & (g2206) & (!g2207)) + ((!dmem_dat_ix2x) & (dmem_dat_ix10x) & (!dmem_dat_ix26x) & (dmem_dat_ix18x) & (g2206) & (g2207)) + ((!dmem_dat_ix2x) & (dmem_dat_ix10x) & (dmem_dat_ix26x) & (!dmem_dat_ix18x) & (!g2206) & (g2207)) + ((!dmem_dat_ix2x) & (dmem_dat_ix10x) & (dmem_dat_ix26x) & (!dmem_dat_ix18x) & (g2206) & (!g2207)) + ((!dmem_dat_ix2x) & (dmem_dat_ix10x) & (dmem_dat_ix26x) & (dmem_dat_ix18x) & (!g2206) & (g2207)) + ((!dmem_dat_ix2x) & (dmem_dat_ix10x) & (dmem_dat_ix26x) & (dmem_dat_ix18x) & (g2206) & (!g2207)) + ((!dmem_dat_ix2x) & (dmem_dat_ix10x) & (dmem_dat_ix26x) & (dmem_dat_ix18x) & (g2206) & (g2207)) + ((dmem_dat_ix2x) & (!dmem_dat_ix10x) & (!dmem_dat_ix26x) & (!dmem_dat_ix18x) & (!g2206) & (!g2207)) + ((dmem_dat_ix2x) & (!dmem_dat_ix10x) & (!dmem_dat_ix26x) & (dmem_dat_ix18x) & (!g2206) & (!g2207)) + ((dmem_dat_ix2x) & (!dmem_dat_ix10x) & (!dmem_dat_ix26x) & (dmem_dat_ix18x) & (g2206) & (g2207)) + ((dmem_dat_ix2x) & (!dmem_dat_ix10x) & (dmem_dat_ix26x) & (!dmem_dat_ix18x) & (!g2206) & (!g2207)) + ((dmem_dat_ix2x) & (!dmem_dat_ix10x) & (dmem_dat_ix26x) & (!dmem_dat_ix18x) & (!g2206) & (g2207)) + ((dmem_dat_ix2x) & (!dmem_dat_ix10x) & (dmem_dat_ix26x) & (dmem_dat_ix18x) & (!g2206) & (!g2207)) + ((dmem_dat_ix2x) & (!dmem_dat_ix10x) & (dmem_dat_ix26x) & (dmem_dat_ix18x) & (!g2206) & (g2207)) + ((dmem_dat_ix2x) & (!dmem_dat_ix10x) & (dmem_dat_ix26x) & (dmem_dat_ix18x) & (g2206) & (g2207)) + ((dmem_dat_ix2x) & (dmem_dat_ix10x) & (!dmem_dat_ix26x) & (!dmem_dat_ix18x) & (!g2206) & (!g2207)) + ((dmem_dat_ix2x) & (dmem_dat_ix10x) & (!dmem_dat_ix26x) & (!dmem_dat_ix18x) & (g2206) & (!g2207)) + ((dmem_dat_ix2x) & (dmem_dat_ix10x) & (!dmem_dat_ix26x) & (dmem_dat_ix18x) & (!g2206) & (!g2207)) + ((dmem_dat_ix2x) & (dmem_dat_ix10x) & (!dmem_dat_ix26x) & (dmem_dat_ix18x) & (g2206) & (!g2207)) + ((dmem_dat_ix2x) & (dmem_dat_ix10x) & (!dmem_dat_ix26x) & (dmem_dat_ix18x) & (g2206) & (g2207)) + ((dmem_dat_ix2x) & (dmem_dat_ix10x) & (dmem_dat_ix26x) & (!dmem_dat_ix18x) & (!g2206) & (!g2207)) + ((dmem_dat_ix2x) & (dmem_dat_ix10x) & (dmem_dat_ix26x) & (!dmem_dat_ix18x) & (!g2206) & (g2207)) + ((dmem_dat_ix2x) & (dmem_dat_ix10x) & (dmem_dat_ix26x) & (!dmem_dat_ix18x) & (g2206) & (!g2207)) + ((dmem_dat_ix2x) & (dmem_dat_ix10x) & (dmem_dat_ix26x) & (dmem_dat_ix18x) & (!g2206) & (!g2207)) + ((dmem_dat_ix2x) & (dmem_dat_ix10x) & (dmem_dat_ix26x) & (dmem_dat_ix18x) & (!g2206) & (g2207)) + ((dmem_dat_ix2x) & (dmem_dat_ix10x) & (dmem_dat_ix26x) & (dmem_dat_ix18x) & (g2206) & (!g2207)) + ((dmem_dat_ix2x) & (dmem_dat_ix10x) & (dmem_dat_ix26x) & (dmem_dat_ix18x) & (g2206) & (g2207)));
	assign g2228 = (((!dmem_dat_ix2x) & (!sk[70]) & (!g2129) & (dmem_dat_ix18x)) + ((!dmem_dat_ix2x) & (!sk[70]) & (g2129) & (!dmem_dat_ix18x)) + ((!dmem_dat_ix2x) & (!sk[70]) & (g2129) & (dmem_dat_ix18x)) + ((!dmem_dat_ix2x) & (sk[70]) & (!g2129) & (dmem_dat_ix18x)) + ((dmem_dat_ix2x) & (!sk[70]) & (!g2129) & (dmem_dat_ix18x)) + ((dmem_dat_ix2x) & (!sk[70]) & (g2129) & (!dmem_dat_ix18x)) + ((dmem_dat_ix2x) & (!sk[70]) & (g2129) & (dmem_dat_ix18x)) + ((dmem_dat_ix2x) & (sk[70]) & (!g2129) & (dmem_dat_ix18x)) + ((dmem_dat_ix2x) & (sk[70]) & (g2129) & (!dmem_dat_ix18x)) + ((dmem_dat_ix2x) & (sk[70]) & (g2129) & (dmem_dat_ix18x)));
	assign g2229 = (((!g75) & (!g2128) & (!g2180) & (!g2226) & (!g2227) & (!g2228)) + ((!g75) & (!g2128) & (!g2180) & (!g2226) & (!g2227) & (g2228)) + ((!g75) & (!g2128) & (!g2180) & (!g2226) & (g2227) & (!g2228)) + ((!g75) & (!g2128) & (!g2180) & (!g2226) & (g2227) & (g2228)) + ((!g75) & (!g2128) & (g2180) & (!g2226) & (!g2227) & (!g2228)) + ((!g75) & (!g2128) & (g2180) & (!g2226) & (!g2227) & (g2228)) + ((!g75) & (!g2128) & (g2180) & (!g2226) & (g2227) & (!g2228)) + ((!g75) & (!g2128) & (g2180) & (!g2226) & (g2227) & (g2228)) + ((!g75) & (g2128) & (!g2180) & (!g2226) & (!g2227) & (!g2228)) + ((!g75) & (g2128) & (!g2180) & (!g2226) & (!g2227) & (g2228)) + ((!g75) & (g2128) & (!g2180) & (!g2226) & (g2227) & (!g2228)) + ((!g75) & (g2128) & (!g2180) & (!g2226) & (g2227) & (g2228)) + ((!g75) & (g2128) & (g2180) & (!g2226) & (!g2227) & (!g2228)) + ((!g75) & (g2128) & (g2180) & (!g2226) & (!g2227) & (g2228)) + ((!g75) & (g2128) & (g2180) & (!g2226) & (g2227) & (!g2228)) + ((!g75) & (g2128) & (g2180) & (!g2226) & (g2227) & (g2228)) + ((g75) & (!g2128) & (!g2180) & (!g2226) & (g2227) & (!g2228)) + ((g75) & (!g2128) & (!g2180) & (!g2226) & (g2227) & (g2228)) + ((g75) & (!g2128) & (!g2180) & (g2226) & (g2227) & (!g2228)) + ((g75) & (!g2128) & (!g2180) & (g2226) & (g2227) & (g2228)) + ((g75) & (!g2128) & (g2180) & (!g2226) & (!g2227) & (g2228)) + ((g75) & (!g2128) & (g2180) & (!g2226) & (g2227) & (g2228)) + ((g75) & (!g2128) & (g2180) & (g2226) & (!g2227) & (g2228)) + ((g75) & (!g2128) & (g2180) & (g2226) & (g2227) & (g2228)) + ((g75) & (g2128) & (!g2180) & (!g2226) & (g2227) & (!g2228)) + ((g75) & (g2128) & (!g2180) & (!g2226) & (g2227) & (g2228)) + ((g75) & (g2128) & (!g2180) & (g2226) & (g2227) & (!g2228)) + ((g75) & (g2128) & (!g2180) & (g2226) & (g2227) & (g2228)));
	assign g2230 = (((!sk[72]) & (g141) & (!g275)) + ((!sk[72]) & (g141) & (g275)) + ((sk[72]) & (!g141) & (g275)) + ((sk[72]) & (g141) & (!g275)));
	assign g5027 = (((!g2921) & (!sk[73]) & (!g3056) & (g2231)) + ((!g2921) & (!sk[73]) & (g3056) & (!g2231)) + ((!g2921) & (!sk[73]) & (g3056) & (g2231)) + ((!g2921) & (sk[73]) & (!g3056) & (g2231)) + ((!g2921) & (sk[73]) & (g3056) & (g2231)) + ((g2921) & (!sk[73]) & (!g3056) & (g2231)) + ((g2921) & (!sk[73]) & (g3056) & (!g2231)) + ((g2921) & (!sk[73]) & (g3056) & (g2231)) + ((g2921) & (sk[73]) & (g3056) & (!g2231)) + ((g2921) & (sk[73]) & (g3056) & (g2231)));
	assign g2232 = (((!sk[74]) & (!g88) & (!g89) & (!g141) & (g275)) + ((!sk[74]) & (!g88) & (!g89) & (g141) & (!g275)) + ((!sk[74]) & (!g88) & (!g89) & (g141) & (g275)) + ((!sk[74]) & (!g88) & (g89) & (!g141) & (!g275)) + ((!sk[74]) & (!g88) & (g89) & (!g141) & (g275)) + ((!sk[74]) & (!g88) & (g89) & (g141) & (!g275)) + ((!sk[74]) & (!g88) & (g89) & (g141) & (g275)) + ((!sk[74]) & (g88) & (!g89) & (!g141) & (g275)) + ((!sk[74]) & (g88) & (!g89) & (g141) & (!g275)) + ((!sk[74]) & (g88) & (!g89) & (g141) & (g275)) + ((!sk[74]) & (g88) & (g89) & (!g141) & (!g275)) + ((!sk[74]) & (g88) & (g89) & (!g141) & (g275)) + ((!sk[74]) & (g88) & (g89) & (g141) & (!g275)) + ((!sk[74]) & (g88) & (g89) & (g141) & (g275)) + ((sk[74]) & (!g88) & (!g89) & (!g141) & (g275)) + ((sk[74]) & (!g88) & (!g89) & (g141) & (g275)) + ((sk[74]) & (!g88) & (g89) & (!g141) & (g275)) + ((sk[74]) & (!g88) & (g89) & (g141) & (!g275)) + ((sk[74]) & (g88) & (!g89) & (!g141) & (!g275)) + ((sk[74]) & (g88) & (!g89) & (g141) & (!g275)) + ((sk[74]) & (g88) & (g89) & (!g141) & (!g275)) + ((sk[74]) & (g88) & (g89) & (g141) & (g275)));
	assign g2233 = (((!g1644) & (!g2033) & (!sk[75]) & (!g2034) & (g2231) & (!g2232)) + ((!g1644) & (!g2033) & (!sk[75]) & (!g2034) & (g2231) & (g2232)) + ((!g1644) & (!g2033) & (!sk[75]) & (g2034) & (!g2231) & (!g2232)) + ((!g1644) & (!g2033) & (!sk[75]) & (g2034) & (!g2231) & (g2232)) + ((!g1644) & (!g2033) & (!sk[75]) & (g2034) & (g2231) & (!g2232)) + ((!g1644) & (!g2033) & (!sk[75]) & (g2034) & (g2231) & (g2232)) + ((!g1644) & (!g2033) & (sk[75]) & (!g2034) & (g2231) & (!g2232)) + ((!g1644) & (!g2033) & (sk[75]) & (!g2034) & (g2231) & (g2232)) + ((!g1644) & (g2033) & (!sk[75]) & (!g2034) & (!g2231) & (!g2232)) + ((!g1644) & (g2033) & (!sk[75]) & (!g2034) & (!g2231) & (g2232)) + ((!g1644) & (g2033) & (!sk[75]) & (!g2034) & (g2231) & (!g2232)) + ((!g1644) & (g2033) & (!sk[75]) & (!g2034) & (g2231) & (g2232)) + ((!g1644) & (g2033) & (!sk[75]) & (g2034) & (!g2231) & (!g2232)) + ((!g1644) & (g2033) & (!sk[75]) & (g2034) & (!g2231) & (g2232)) + ((!g1644) & (g2033) & (!sk[75]) & (g2034) & (g2231) & (!g2232)) + ((!g1644) & (g2033) & (!sk[75]) & (g2034) & (g2231) & (g2232)) + ((!g1644) & (g2033) & (sk[75]) & (!g2034) & (!g2231) & (g2232)) + ((!g1644) & (g2033) & (sk[75]) & (!g2034) & (g2231) & (g2232)) + ((g1644) & (!g2033) & (!sk[75]) & (!g2034) & (g2231) & (!g2232)) + ((g1644) & (!g2033) & (!sk[75]) & (!g2034) & (g2231) & (g2232)) + ((g1644) & (!g2033) & (!sk[75]) & (g2034) & (!g2231) & (!g2232)) + ((g1644) & (!g2033) & (!sk[75]) & (g2034) & (!g2231) & (g2232)) + ((g1644) & (!g2033) & (!sk[75]) & (g2034) & (g2231) & (!g2232)) + ((g1644) & (!g2033) & (!sk[75]) & (g2034) & (g2231) & (g2232)) + ((g1644) & (!g2033) & (sk[75]) & (!g2034) & (g2231) & (!g2232)) + ((g1644) & (!g2033) & (sk[75]) & (!g2034) & (g2231) & (g2232)) + ((g1644) & (!g2033) & (sk[75]) & (g2034) & (!g2231) & (!g2232)) + ((g1644) & (!g2033) & (sk[75]) & (g2034) & (!g2231) & (g2232)) + ((g1644) & (!g2033) & (sk[75]) & (g2034) & (g2231) & (!g2232)) + ((g1644) & (!g2033) & (sk[75]) & (g2034) & (g2231) & (g2232)) + ((g1644) & (g2033) & (!sk[75]) & (!g2034) & (!g2231) & (!g2232)) + ((g1644) & (g2033) & (!sk[75]) & (!g2034) & (!g2231) & (g2232)) + ((g1644) & (g2033) & (!sk[75]) & (!g2034) & (g2231) & (!g2232)) + ((g1644) & (g2033) & (!sk[75]) & (!g2034) & (g2231) & (g2232)) + ((g1644) & (g2033) & (!sk[75]) & (g2034) & (!g2231) & (!g2232)) + ((g1644) & (g2033) & (!sk[75]) & (g2034) & (!g2231) & (g2232)) + ((g1644) & (g2033) & (!sk[75]) & (g2034) & (g2231) & (!g2232)) + ((g1644) & (g2033) & (!sk[75]) & (g2034) & (g2231) & (g2232)) + ((g1644) & (g2033) & (sk[75]) & (!g2034) & (!g2231) & (g2232)) + ((g1644) & (g2033) & (sk[75]) & (!g2034) & (g2231) & (g2232)));
	assign g2234 = (((!g2022) & (!nmi_i) & (!g2023) & (!g2029) & (!g2230) & (g2233)) + ((!g2022) & (!nmi_i) & (!g2023) & (!g2029) & (g2230) & (g2233)) + ((!g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2230) & (!g2233)) + ((!g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2230) & (g2233)) + ((!g2022) & (!nmi_i) & (g2023) & (!g2029) & (!g2230) & (g2233)) + ((!g2022) & (!nmi_i) & (g2023) & (!g2029) & (g2230) & (g2233)) + ((!g2022) & (!nmi_i) & (g2023) & (g2029) & (g2230) & (!g2233)) + ((!g2022) & (!nmi_i) & (g2023) & (g2029) & (g2230) & (g2233)) + ((!g2022) & (nmi_i) & (!g2023) & (!g2029) & (!g2230) & (g2233)) + ((!g2022) & (nmi_i) & (!g2023) & (!g2029) & (g2230) & (g2233)) + ((!g2022) & (nmi_i) & (!g2023) & (g2029) & (g2230) & (!g2233)) + ((!g2022) & (nmi_i) & (!g2023) & (g2029) & (g2230) & (g2233)) + ((!g2022) & (nmi_i) & (g2023) & (!g2029) & (!g2230) & (g2233)) + ((!g2022) & (nmi_i) & (g2023) & (!g2029) & (g2230) & (g2233)) + ((!g2022) & (nmi_i) & (g2023) & (g2029) & (g2230) & (!g2233)) + ((!g2022) & (nmi_i) & (g2023) & (g2029) & (g2230) & (g2233)) + ((g2022) & (!nmi_i) & (!g2023) & (!g2029) & (!g2230) & (g2233)) + ((g2022) & (!nmi_i) & (!g2023) & (!g2029) & (g2230) & (g2233)) + ((g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2230) & (!g2233)) + ((g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2230) & (g2233)));
	assign g2235 = (((!g123) & (!intr_i) & (!g2039) & (!g2056) & (!g2057) & (g2234)) + ((!g123) & (!intr_i) & (!g2039) & (!g2056) & (g2057) & (g2234)) + ((!g123) & (!intr_i) & (!g2039) & (g2056) & (!g2057) & (g2234)) + ((!g123) & (!intr_i) & (!g2039) & (g2056) & (g2057) & (g2234)) + ((!g123) & (!intr_i) & (g2039) & (!g2056) & (!g2057) & (g2234)) + ((!g123) & (!intr_i) & (g2039) & (!g2056) & (g2057) & (g2234)) + ((!g123) & (!intr_i) & (g2039) & (g2056) & (!g2057) & (g2234)) + ((!g123) & (!intr_i) & (g2039) & (g2056) & (g2057) & (g2234)) + ((!g123) & (intr_i) & (!g2039) & (!g2056) & (!g2057) & (g2234)) + ((!g123) & (intr_i) & (!g2039) & (!g2056) & (g2057) & (g2234)) + ((!g123) & (intr_i) & (!g2039) & (g2056) & (!g2057) & (g2234)) + ((!g123) & (intr_i) & (g2039) & (!g2056) & (!g2057) & (g2234)) + ((!g123) & (intr_i) & (g2039) & (g2056) & (!g2057) & (g2234)));
	assign g2236 = (((!g2106) & (!g2105) & (!g2104) & (g2070) & (g2071) & (g2074)) + ((!g2106) & (!g2105) & (g2104) & (!g2070) & (!g2071) & (g2074)) + ((!g2106) & (!g2105) & (g2104) & (g2070) & (!g2071) & (g2074)) + ((!g2106) & (!g2105) & (g2104) & (g2070) & (g2071) & (g2074)) + ((!g2106) & (g2105) & (!g2104) & (!g2070) & (g2071) & (!g2074)) + ((!g2106) & (g2105) & (!g2104) & (g2070) & (g2071) & (!g2074)) + ((!g2106) & (g2105) & (!g2104) & (g2070) & (g2071) & (g2074)) + ((!g2106) & (g2105) & (g2104) & (!g2070) & (!g2071) & (g2074)) + ((!g2106) & (g2105) & (g2104) & (!g2070) & (g2071) & (!g2074)) + ((!g2106) & (g2105) & (g2104) & (g2070) & (!g2071) & (g2074)) + ((!g2106) & (g2105) & (g2104) & (g2070) & (g2071) & (!g2074)) + ((!g2106) & (g2105) & (g2104) & (g2070) & (g2071) & (g2074)) + ((g2106) & (!g2105) & (!g2104) & (!g2070) & (!g2071) & (!g2074)) + ((g2106) & (!g2105) & (!g2104) & (g2070) & (!g2071) & (!g2074)) + ((g2106) & (!g2105) & (!g2104) & (g2070) & (g2071) & (g2074)) + ((g2106) & (!g2105) & (g2104) & (!g2070) & (!g2071) & (!g2074)) + ((g2106) & (!g2105) & (g2104) & (!g2070) & (!g2071) & (g2074)) + ((g2106) & (!g2105) & (g2104) & (g2070) & (!g2071) & (!g2074)) + ((g2106) & (!g2105) & (g2104) & (g2070) & (!g2071) & (g2074)) + ((g2106) & (!g2105) & (g2104) & (g2070) & (g2071) & (g2074)) + ((g2106) & (g2105) & (!g2104) & (!g2070) & (!g2071) & (!g2074)) + ((g2106) & (g2105) & (!g2104) & (!g2070) & (g2071) & (!g2074)) + ((g2106) & (g2105) & (!g2104) & (g2070) & (!g2071) & (!g2074)) + ((g2106) & (g2105) & (!g2104) & (g2070) & (g2071) & (!g2074)) + ((g2106) & (g2105) & (!g2104) & (g2070) & (g2071) & (g2074)) + ((g2106) & (g2105) & (g2104) & (!g2070) & (!g2071) & (!g2074)) + ((g2106) & (g2105) & (g2104) & (!g2070) & (!g2071) & (g2074)) + ((g2106) & (g2105) & (g2104) & (!g2070) & (g2071) & (!g2074)) + ((g2106) & (g2105) & (g2104) & (g2070) & (!g2071) & (!g2074)) + ((g2106) & (g2105) & (g2104) & (g2070) & (!g2071) & (g2074)) + ((g2106) & (g2105) & (g2104) & (g2070) & (g2071) & (!g2074)) + ((g2106) & (g2105) & (g2104) & (g2070) & (g2071) & (g2074)));
	assign g2237 = (((!g2076) & (!g2077) & (!sk[79]) & (g2236)) + ((!g2076) & (!g2077) & (sk[79]) & (g2236)) + ((!g2076) & (g2077) & (!sk[79]) & (!g2236)) + ((!g2076) & (g2077) & (!sk[79]) & (g2236)) + ((g2076) & (!g2077) & (!sk[79]) & (g2236)) + ((g2076) & (g2077) & (!sk[79]) & (!g2236)) + ((g2076) & (g2077) & (!sk[79]) & (g2236)));
	assign g2238 = (((!g2074) & (!g2071) & (!g2070) & (g2077) & (g2105) & (!g2104)) + ((!g2074) & (!g2071) & (!g2070) & (g2077) & (g2105) & (g2104)) + ((!g2074) & (!g2071) & (g2070) & (g2077) & (g2105) & (!g2104)) + ((!g2074) & (!g2071) & (g2070) & (g2077) & (g2105) & (g2104)) + ((!g2074) & (g2071) & (!g2070) & (g2077) & (g2105) & (!g2104)) + ((!g2074) & (g2071) & (!g2070) & (g2077) & (g2105) & (g2104)) + ((!g2074) & (g2071) & (g2070) & (!g2077) & (g2105) & (g2104)) + ((!g2074) & (g2071) & (g2070) & (g2077) & (!g2105) & (g2104)) + ((!g2074) & (g2071) & (g2070) & (g2077) & (g2105) & (!g2104)) + ((!g2074) & (g2071) & (g2070) & (g2077) & (g2105) & (g2104)) + ((g2074) & (!g2071) & (!g2070) & (!g2077) & (g2105) & (g2104)) + ((g2074) & (!g2071) & (!g2070) & (g2077) & (!g2105) & (g2104)) + ((g2074) & (!g2071) & (!g2070) & (g2077) & (g2105) & (!g2104)) + ((g2074) & (!g2071) & (!g2070) & (g2077) & (g2105) & (g2104)) + ((g2074) & (!g2071) & (g2070) & (!g2077) & (g2105) & (g2104)) + ((g2074) & (!g2071) & (g2070) & (g2077) & (!g2105) & (g2104)) + ((g2074) & (!g2071) & (g2070) & (g2077) & (g2105) & (!g2104)) + ((g2074) & (!g2071) & (g2070) & (g2077) & (g2105) & (g2104)) + ((g2074) & (g2071) & (!g2070) & (!g2077) & (g2105) & (g2104)) + ((g2074) & (g2071) & (!g2070) & (g2077) & (!g2105) & (g2104)) + ((g2074) & (g2071) & (!g2070) & (g2077) & (g2105) & (!g2104)) + ((g2074) & (g2071) & (!g2070) & (g2077) & (g2105) & (g2104)) + ((g2074) & (g2071) & (g2070) & (!g2077) & (g2105) & (!g2104)) + ((g2074) & (g2071) & (g2070) & (!g2077) & (g2105) & (g2104)) + ((g2074) & (g2071) & (g2070) & (g2077) & (!g2105) & (!g2104)) + ((g2074) & (g2071) & (g2070) & (g2077) & (!g2105) & (g2104)) + ((g2074) & (g2071) & (g2070) & (g2077) & (g2105) & (!g2104)) + ((g2074) & (g2071) & (g2070) & (g2077) & (g2105) & (g2104)));
	assign g2239 = (((!sk[81]) & (!g2076) & (!g2106) & (g2238)) + ((!sk[81]) & (!g2076) & (g2106) & (!g2238)) + ((!sk[81]) & (!g2076) & (g2106) & (g2238)) + ((!sk[81]) & (g2076) & (!g2106) & (g2238)) + ((!sk[81]) & (g2076) & (g2106) & (!g2238)) + ((!sk[81]) & (g2076) & (g2106) & (g2238)) + ((sk[81]) & (!g2076) & (!g2106) & (g2238)) + ((sk[81]) & (!g2076) & (g2106) & (!g2238)) + ((sk[81]) & (g2076) & (!g2106) & (!g2238)) + ((sk[81]) & (g2076) & (g2106) & (g2238)));
	assign g2240 = (((!g2072) & (!g2079) & (!sk[82]) & (!g2185) & (g2213)) + ((!g2072) & (!g2079) & (!sk[82]) & (g2185) & (!g2213)) + ((!g2072) & (!g2079) & (!sk[82]) & (g2185) & (g2213)) + ((!g2072) & (g2079) & (!sk[82]) & (!g2185) & (!g2213)) + ((!g2072) & (g2079) & (!sk[82]) & (!g2185) & (g2213)) + ((!g2072) & (g2079) & (!sk[82]) & (g2185) & (!g2213)) + ((!g2072) & (g2079) & (!sk[82]) & (g2185) & (g2213)) + ((g2072) & (!g2079) & (!sk[82]) & (!g2185) & (g2213)) + ((g2072) & (!g2079) & (!sk[82]) & (g2185) & (!g2213)) + ((g2072) & (!g2079) & (!sk[82]) & (g2185) & (g2213)) + ((g2072) & (g2079) & (!sk[82]) & (!g2185) & (!g2213)) + ((g2072) & (g2079) & (!sk[82]) & (!g2185) & (g2213)) + ((g2072) & (g2079) & (!sk[82]) & (g2185) & (!g2213)) + ((g2072) & (g2079) & (!sk[82]) & (g2185) & (g2213)) + ((g2072) & (g2079) & (sk[82]) & (g2185) & (g2213)));
	assign g2241 = (((!g2076) & (sk[83]) & (!g2106)) + ((g2076) & (!sk[83]) & (!g2106)) + ((g2076) & (!sk[83]) & (g2106)) + ((g2076) & (sk[83]) & (g2106)));
	assign g2242 = (((!g2086) & (!g2093) & (!g2094) & (g2095) & (g2071) & (g2074)) + ((!g2086) & (!g2093) & (g2094) & (!g2095) & (!g2071) & (g2074)) + ((!g2086) & (!g2093) & (g2094) & (g2095) & (!g2071) & (g2074)) + ((!g2086) & (!g2093) & (g2094) & (g2095) & (g2071) & (g2074)) + ((!g2086) & (g2093) & (!g2094) & (!g2095) & (g2071) & (!g2074)) + ((!g2086) & (g2093) & (!g2094) & (g2095) & (g2071) & (!g2074)) + ((!g2086) & (g2093) & (!g2094) & (g2095) & (g2071) & (g2074)) + ((!g2086) & (g2093) & (g2094) & (!g2095) & (!g2071) & (g2074)) + ((!g2086) & (g2093) & (g2094) & (!g2095) & (g2071) & (!g2074)) + ((!g2086) & (g2093) & (g2094) & (g2095) & (!g2071) & (g2074)) + ((!g2086) & (g2093) & (g2094) & (g2095) & (g2071) & (!g2074)) + ((!g2086) & (g2093) & (g2094) & (g2095) & (g2071) & (g2074)) + ((g2086) & (!g2093) & (!g2094) & (!g2095) & (!g2071) & (!g2074)) + ((g2086) & (!g2093) & (!g2094) & (g2095) & (!g2071) & (!g2074)) + ((g2086) & (!g2093) & (!g2094) & (g2095) & (g2071) & (g2074)) + ((g2086) & (!g2093) & (g2094) & (!g2095) & (!g2071) & (!g2074)) + ((g2086) & (!g2093) & (g2094) & (!g2095) & (!g2071) & (g2074)) + ((g2086) & (!g2093) & (g2094) & (g2095) & (!g2071) & (!g2074)) + ((g2086) & (!g2093) & (g2094) & (g2095) & (!g2071) & (g2074)) + ((g2086) & (!g2093) & (g2094) & (g2095) & (g2071) & (g2074)) + ((g2086) & (g2093) & (!g2094) & (!g2095) & (!g2071) & (!g2074)) + ((g2086) & (g2093) & (!g2094) & (!g2095) & (g2071) & (!g2074)) + ((g2086) & (g2093) & (!g2094) & (g2095) & (!g2071) & (!g2074)) + ((g2086) & (g2093) & (!g2094) & (g2095) & (g2071) & (!g2074)) + ((g2086) & (g2093) & (!g2094) & (g2095) & (g2071) & (g2074)) + ((g2086) & (g2093) & (g2094) & (!g2095) & (!g2071) & (!g2074)) + ((g2086) & (g2093) & (g2094) & (!g2095) & (!g2071) & (g2074)) + ((g2086) & (g2093) & (g2094) & (!g2095) & (g2071) & (!g2074)) + ((g2086) & (g2093) & (g2094) & (g2095) & (!g2071) & (!g2074)) + ((g2086) & (g2093) & (g2094) & (g2095) & (!g2071) & (g2074)) + ((g2086) & (g2093) & (g2094) & (g2095) & (g2071) & (!g2074)) + ((g2086) & (g2093) & (g2094) & (g2095) & (g2071) & (g2074)));
	assign g2243 = (((!g2091) & (!g2098) & (!g2099) & (g2100) & (g2071) & (g2074)) + ((!g2091) & (!g2098) & (g2099) & (!g2100) & (!g2071) & (g2074)) + ((!g2091) & (!g2098) & (g2099) & (g2100) & (!g2071) & (g2074)) + ((!g2091) & (!g2098) & (g2099) & (g2100) & (g2071) & (g2074)) + ((!g2091) & (g2098) & (!g2099) & (!g2100) & (g2071) & (!g2074)) + ((!g2091) & (g2098) & (!g2099) & (g2100) & (g2071) & (!g2074)) + ((!g2091) & (g2098) & (!g2099) & (g2100) & (g2071) & (g2074)) + ((!g2091) & (g2098) & (g2099) & (!g2100) & (!g2071) & (g2074)) + ((!g2091) & (g2098) & (g2099) & (!g2100) & (g2071) & (!g2074)) + ((!g2091) & (g2098) & (g2099) & (g2100) & (!g2071) & (g2074)) + ((!g2091) & (g2098) & (g2099) & (g2100) & (g2071) & (!g2074)) + ((!g2091) & (g2098) & (g2099) & (g2100) & (g2071) & (g2074)) + ((g2091) & (!g2098) & (!g2099) & (!g2100) & (!g2071) & (!g2074)) + ((g2091) & (!g2098) & (!g2099) & (g2100) & (!g2071) & (!g2074)) + ((g2091) & (!g2098) & (!g2099) & (g2100) & (g2071) & (g2074)) + ((g2091) & (!g2098) & (g2099) & (!g2100) & (!g2071) & (!g2074)) + ((g2091) & (!g2098) & (g2099) & (!g2100) & (!g2071) & (g2074)) + ((g2091) & (!g2098) & (g2099) & (g2100) & (!g2071) & (!g2074)) + ((g2091) & (!g2098) & (g2099) & (g2100) & (!g2071) & (g2074)) + ((g2091) & (!g2098) & (g2099) & (g2100) & (g2071) & (g2074)) + ((g2091) & (g2098) & (!g2099) & (!g2100) & (!g2071) & (!g2074)) + ((g2091) & (g2098) & (!g2099) & (!g2100) & (g2071) & (!g2074)) + ((g2091) & (g2098) & (!g2099) & (g2100) & (!g2071) & (!g2074)) + ((g2091) & (g2098) & (!g2099) & (g2100) & (g2071) & (!g2074)) + ((g2091) & (g2098) & (!g2099) & (g2100) & (g2071) & (g2074)) + ((g2091) & (g2098) & (g2099) & (!g2100) & (!g2071) & (!g2074)) + ((g2091) & (g2098) & (g2099) & (!g2100) & (!g2071) & (g2074)) + ((g2091) & (g2098) & (g2099) & (!g2100) & (g2071) & (!g2074)) + ((g2091) & (g2098) & (g2099) & (g2100) & (!g2071) & (!g2074)) + ((g2091) & (g2098) & (g2099) & (g2100) & (!g2071) & (g2074)) + ((g2091) & (g2098) & (g2099) & (g2100) & (g2071) & (!g2074)) + ((g2091) & (g2098) & (g2099) & (g2100) & (g2071) & (g2074)));
	assign g2244 = (((!g2096) & (!g2088) & (!g2089) & (g2090) & (g2071) & (g2074)) + ((!g2096) & (!g2088) & (g2089) & (!g2090) & (!g2071) & (g2074)) + ((!g2096) & (!g2088) & (g2089) & (g2090) & (!g2071) & (g2074)) + ((!g2096) & (!g2088) & (g2089) & (g2090) & (g2071) & (g2074)) + ((!g2096) & (g2088) & (!g2089) & (!g2090) & (g2071) & (!g2074)) + ((!g2096) & (g2088) & (!g2089) & (g2090) & (g2071) & (!g2074)) + ((!g2096) & (g2088) & (!g2089) & (g2090) & (g2071) & (g2074)) + ((!g2096) & (g2088) & (g2089) & (!g2090) & (!g2071) & (g2074)) + ((!g2096) & (g2088) & (g2089) & (!g2090) & (g2071) & (!g2074)) + ((!g2096) & (g2088) & (g2089) & (g2090) & (!g2071) & (g2074)) + ((!g2096) & (g2088) & (g2089) & (g2090) & (g2071) & (!g2074)) + ((!g2096) & (g2088) & (g2089) & (g2090) & (g2071) & (g2074)) + ((g2096) & (!g2088) & (!g2089) & (!g2090) & (!g2071) & (!g2074)) + ((g2096) & (!g2088) & (!g2089) & (g2090) & (!g2071) & (!g2074)) + ((g2096) & (!g2088) & (!g2089) & (g2090) & (g2071) & (g2074)) + ((g2096) & (!g2088) & (g2089) & (!g2090) & (!g2071) & (!g2074)) + ((g2096) & (!g2088) & (g2089) & (!g2090) & (!g2071) & (g2074)) + ((g2096) & (!g2088) & (g2089) & (g2090) & (!g2071) & (!g2074)) + ((g2096) & (!g2088) & (g2089) & (g2090) & (!g2071) & (g2074)) + ((g2096) & (!g2088) & (g2089) & (g2090) & (g2071) & (g2074)) + ((g2096) & (g2088) & (!g2089) & (!g2090) & (!g2071) & (!g2074)) + ((g2096) & (g2088) & (!g2089) & (!g2090) & (g2071) & (!g2074)) + ((g2096) & (g2088) & (!g2089) & (g2090) & (!g2071) & (!g2074)) + ((g2096) & (g2088) & (!g2089) & (g2090) & (g2071) & (!g2074)) + ((g2096) & (g2088) & (!g2089) & (g2090) & (g2071) & (g2074)) + ((g2096) & (g2088) & (g2089) & (!g2090) & (!g2071) & (!g2074)) + ((g2096) & (g2088) & (g2089) & (!g2090) & (!g2071) & (g2074)) + ((g2096) & (g2088) & (g2089) & (!g2090) & (g2071) & (!g2074)) + ((g2096) & (g2088) & (g2089) & (g2090) & (!g2071) & (!g2074)) + ((g2096) & (g2088) & (g2089) & (g2090) & (!g2071) & (g2074)) + ((g2096) & (g2088) & (g2089) & (g2090) & (g2071) & (!g2074)) + ((g2096) & (g2088) & (g2089) & (g2090) & (g2071) & (g2074)));
	assign g2245 = (((!g2074) & (!g2071) & (!sk[87]) & (!g2101) & (g2192)) + ((!g2074) & (!g2071) & (!sk[87]) & (g2101) & (!g2192)) + ((!g2074) & (!g2071) & (!sk[87]) & (g2101) & (g2192)) + ((!g2074) & (!g2071) & (sk[87]) & (g2101) & (!g2192)) + ((!g2074) & (!g2071) & (sk[87]) & (g2101) & (g2192)) + ((!g2074) & (g2071) & (!sk[87]) & (!g2101) & (!g2192)) + ((!g2074) & (g2071) & (!sk[87]) & (!g2101) & (g2192)) + ((!g2074) & (g2071) & (!sk[87]) & (g2101) & (!g2192)) + ((!g2074) & (g2071) & (!sk[87]) & (g2101) & (g2192)) + ((!g2074) & (g2071) & (sk[87]) & (!g2101) & (g2192)) + ((!g2074) & (g2071) & (sk[87]) & (g2101) & (g2192)) + ((g2074) & (!g2071) & (!sk[87]) & (!g2101) & (g2192)) + ((g2074) & (!g2071) & (!sk[87]) & (g2101) & (!g2192)) + ((g2074) & (!g2071) & (!sk[87]) & (g2101) & (g2192)) + ((g2074) & (!g2071) & (sk[87]) & (!g2101) & (g2192)) + ((g2074) & (!g2071) & (sk[87]) & (g2101) & (g2192)) + ((g2074) & (g2071) & (!sk[87]) & (!g2101) & (!g2192)) + ((g2074) & (g2071) & (!sk[87]) & (!g2101) & (g2192)) + ((g2074) & (g2071) & (!sk[87]) & (g2101) & (!g2192)) + ((g2074) & (g2071) & (!sk[87]) & (g2101) & (g2192)) + ((g2074) & (g2071) & (sk[87]) & (!g2101) & (g2192)) + ((g2074) & (g2071) & (sk[87]) & (g2101) & (g2192)));
	assign g2246 = (((!g2242) & (!g2243) & (!g2244) & (g2245) & (g2076) & (g2077)) + ((!g2242) & (!g2243) & (g2244) & (!g2245) & (!g2076) & (g2077)) + ((!g2242) & (!g2243) & (g2244) & (g2245) & (!g2076) & (g2077)) + ((!g2242) & (!g2243) & (g2244) & (g2245) & (g2076) & (g2077)) + ((!g2242) & (g2243) & (!g2244) & (!g2245) & (g2076) & (!g2077)) + ((!g2242) & (g2243) & (!g2244) & (g2245) & (g2076) & (!g2077)) + ((!g2242) & (g2243) & (!g2244) & (g2245) & (g2076) & (g2077)) + ((!g2242) & (g2243) & (g2244) & (!g2245) & (!g2076) & (g2077)) + ((!g2242) & (g2243) & (g2244) & (!g2245) & (g2076) & (!g2077)) + ((!g2242) & (g2243) & (g2244) & (g2245) & (!g2076) & (g2077)) + ((!g2242) & (g2243) & (g2244) & (g2245) & (g2076) & (!g2077)) + ((!g2242) & (g2243) & (g2244) & (g2245) & (g2076) & (g2077)) + ((g2242) & (!g2243) & (!g2244) & (!g2245) & (!g2076) & (!g2077)) + ((g2242) & (!g2243) & (!g2244) & (g2245) & (!g2076) & (!g2077)) + ((g2242) & (!g2243) & (!g2244) & (g2245) & (g2076) & (g2077)) + ((g2242) & (!g2243) & (g2244) & (!g2245) & (!g2076) & (!g2077)) + ((g2242) & (!g2243) & (g2244) & (!g2245) & (!g2076) & (g2077)) + ((g2242) & (!g2243) & (g2244) & (g2245) & (!g2076) & (!g2077)) + ((g2242) & (!g2243) & (g2244) & (g2245) & (!g2076) & (g2077)) + ((g2242) & (!g2243) & (g2244) & (g2245) & (g2076) & (g2077)) + ((g2242) & (g2243) & (!g2244) & (!g2245) & (!g2076) & (!g2077)) + ((g2242) & (g2243) & (!g2244) & (!g2245) & (g2076) & (!g2077)) + ((g2242) & (g2243) & (!g2244) & (g2245) & (!g2076) & (!g2077)) + ((g2242) & (g2243) & (!g2244) & (g2245) & (g2076) & (!g2077)) + ((g2242) & (g2243) & (!g2244) & (g2245) & (g2076) & (g2077)) + ((g2242) & (g2243) & (g2244) & (!g2245) & (!g2076) & (!g2077)) + ((g2242) & (g2243) & (g2244) & (!g2245) & (!g2076) & (g2077)) + ((g2242) & (g2243) & (g2244) & (!g2245) & (g2076) & (!g2077)) + ((g2242) & (g2243) & (g2244) & (g2245) & (!g2076) & (!g2077)) + ((g2242) & (g2243) & (g2244) & (g2245) & (!g2076) & (g2077)) + ((g2242) & (g2243) & (g2244) & (g2245) & (g2076) & (!g2077)) + ((g2242) & (g2243) & (g2244) & (g2245) & (g2076) & (g2077)));
	assign g2247 = (((!g2116) & (!g2108) & (!g2109) & (g2110) & (g2071) & (g2074)) + ((!g2116) & (!g2108) & (g2109) & (!g2110) & (!g2071) & (g2074)) + ((!g2116) & (!g2108) & (g2109) & (g2110) & (!g2071) & (g2074)) + ((!g2116) & (!g2108) & (g2109) & (g2110) & (g2071) & (g2074)) + ((!g2116) & (g2108) & (!g2109) & (!g2110) & (g2071) & (!g2074)) + ((!g2116) & (g2108) & (!g2109) & (g2110) & (g2071) & (!g2074)) + ((!g2116) & (g2108) & (!g2109) & (g2110) & (g2071) & (g2074)) + ((!g2116) & (g2108) & (g2109) & (!g2110) & (!g2071) & (g2074)) + ((!g2116) & (g2108) & (g2109) & (!g2110) & (g2071) & (!g2074)) + ((!g2116) & (g2108) & (g2109) & (g2110) & (!g2071) & (g2074)) + ((!g2116) & (g2108) & (g2109) & (g2110) & (g2071) & (!g2074)) + ((!g2116) & (g2108) & (g2109) & (g2110) & (g2071) & (g2074)) + ((g2116) & (!g2108) & (!g2109) & (!g2110) & (!g2071) & (!g2074)) + ((g2116) & (!g2108) & (!g2109) & (g2110) & (!g2071) & (!g2074)) + ((g2116) & (!g2108) & (!g2109) & (g2110) & (g2071) & (g2074)) + ((g2116) & (!g2108) & (g2109) & (!g2110) & (!g2071) & (!g2074)) + ((g2116) & (!g2108) & (g2109) & (!g2110) & (!g2071) & (g2074)) + ((g2116) & (!g2108) & (g2109) & (g2110) & (!g2071) & (!g2074)) + ((g2116) & (!g2108) & (g2109) & (g2110) & (!g2071) & (g2074)) + ((g2116) & (!g2108) & (g2109) & (g2110) & (g2071) & (g2074)) + ((g2116) & (g2108) & (!g2109) & (!g2110) & (!g2071) & (!g2074)) + ((g2116) & (g2108) & (!g2109) & (!g2110) & (g2071) & (!g2074)) + ((g2116) & (g2108) & (!g2109) & (g2110) & (!g2071) & (!g2074)) + ((g2116) & (g2108) & (!g2109) & (g2110) & (g2071) & (!g2074)) + ((g2116) & (g2108) & (!g2109) & (g2110) & (g2071) & (g2074)) + ((g2116) & (g2108) & (g2109) & (!g2110) & (!g2071) & (!g2074)) + ((g2116) & (g2108) & (g2109) & (!g2110) & (!g2071) & (g2074)) + ((g2116) & (g2108) & (g2109) & (!g2110) & (g2071) & (!g2074)) + ((g2116) & (g2108) & (g2109) & (g2110) & (!g2071) & (!g2074)) + ((g2116) & (g2108) & (g2109) & (g2110) & (!g2071) & (g2074)) + ((g2116) & (g2108) & (g2109) & (g2110) & (g2071) & (!g2074)) + ((g2116) & (g2108) & (g2109) & (g2110) & (g2071) & (g2074)));
	assign g2248 = (((!g2247) & (!g2113) & (!g2114) & (g2115) & (g2196) & (g2197)) + ((!g2247) & (!g2113) & (g2114) & (!g2115) & (!g2196) & (g2197)) + ((!g2247) & (!g2113) & (g2114) & (g2115) & (!g2196) & (g2197)) + ((!g2247) & (!g2113) & (g2114) & (g2115) & (g2196) & (g2197)) + ((!g2247) & (g2113) & (!g2114) & (!g2115) & (g2196) & (!g2197)) + ((!g2247) & (g2113) & (!g2114) & (g2115) & (g2196) & (!g2197)) + ((!g2247) & (g2113) & (!g2114) & (g2115) & (g2196) & (g2197)) + ((!g2247) & (g2113) & (g2114) & (!g2115) & (!g2196) & (g2197)) + ((!g2247) & (g2113) & (g2114) & (!g2115) & (g2196) & (!g2197)) + ((!g2247) & (g2113) & (g2114) & (g2115) & (!g2196) & (g2197)) + ((!g2247) & (g2113) & (g2114) & (g2115) & (g2196) & (!g2197)) + ((!g2247) & (g2113) & (g2114) & (g2115) & (g2196) & (g2197)) + ((g2247) & (!g2113) & (!g2114) & (!g2115) & (!g2196) & (!g2197)) + ((g2247) & (!g2113) & (!g2114) & (g2115) & (!g2196) & (!g2197)) + ((g2247) & (!g2113) & (!g2114) & (g2115) & (g2196) & (g2197)) + ((g2247) & (!g2113) & (g2114) & (!g2115) & (!g2196) & (!g2197)) + ((g2247) & (!g2113) & (g2114) & (!g2115) & (!g2196) & (g2197)) + ((g2247) & (!g2113) & (g2114) & (g2115) & (!g2196) & (!g2197)) + ((g2247) & (!g2113) & (g2114) & (g2115) & (!g2196) & (g2197)) + ((g2247) & (!g2113) & (g2114) & (g2115) & (g2196) & (g2197)) + ((g2247) & (g2113) & (!g2114) & (!g2115) & (!g2196) & (!g2197)) + ((g2247) & (g2113) & (!g2114) & (!g2115) & (g2196) & (!g2197)) + ((g2247) & (g2113) & (!g2114) & (g2115) & (!g2196) & (!g2197)) + ((g2247) & (g2113) & (!g2114) & (g2115) & (g2196) & (!g2197)) + ((g2247) & (g2113) & (!g2114) & (g2115) & (g2196) & (g2197)) + ((g2247) & (g2113) & (g2114) & (!g2115) & (!g2196) & (!g2197)) + ((g2247) & (g2113) & (g2114) & (!g2115) & (!g2196) & (g2197)) + ((g2247) & (g2113) & (g2114) & (!g2115) & (g2196) & (!g2197)) + ((g2247) & (g2113) & (g2114) & (g2115) & (!g2196) & (!g2197)) + ((g2247) & (g2113) & (g2114) & (g2115) & (!g2196) & (g2197)) + ((g2247) & (g2113) & (g2114) & (g2115) & (g2196) & (!g2197)) + ((g2247) & (g2113) & (g2114) & (g2115) & (g2196) & (g2197)));
	assign g2249 = (((!g2111) & (!g2118) & (!g2119) & (g2120) & (g2071) & (g2074)) + ((!g2111) & (!g2118) & (g2119) & (!g2120) & (!g2071) & (g2074)) + ((!g2111) & (!g2118) & (g2119) & (g2120) & (!g2071) & (g2074)) + ((!g2111) & (!g2118) & (g2119) & (g2120) & (g2071) & (g2074)) + ((!g2111) & (g2118) & (!g2119) & (!g2120) & (g2071) & (!g2074)) + ((!g2111) & (g2118) & (!g2119) & (g2120) & (g2071) & (!g2074)) + ((!g2111) & (g2118) & (!g2119) & (g2120) & (g2071) & (g2074)) + ((!g2111) & (g2118) & (g2119) & (!g2120) & (!g2071) & (g2074)) + ((!g2111) & (g2118) & (g2119) & (!g2120) & (g2071) & (!g2074)) + ((!g2111) & (g2118) & (g2119) & (g2120) & (!g2071) & (g2074)) + ((!g2111) & (g2118) & (g2119) & (g2120) & (g2071) & (!g2074)) + ((!g2111) & (g2118) & (g2119) & (g2120) & (g2071) & (g2074)) + ((g2111) & (!g2118) & (!g2119) & (!g2120) & (!g2071) & (!g2074)) + ((g2111) & (!g2118) & (!g2119) & (g2120) & (!g2071) & (!g2074)) + ((g2111) & (!g2118) & (!g2119) & (g2120) & (g2071) & (g2074)) + ((g2111) & (!g2118) & (g2119) & (!g2120) & (!g2071) & (!g2074)) + ((g2111) & (!g2118) & (g2119) & (!g2120) & (!g2071) & (g2074)) + ((g2111) & (!g2118) & (g2119) & (g2120) & (!g2071) & (!g2074)) + ((g2111) & (!g2118) & (g2119) & (g2120) & (!g2071) & (g2074)) + ((g2111) & (!g2118) & (g2119) & (g2120) & (g2071) & (g2074)) + ((g2111) & (g2118) & (!g2119) & (!g2120) & (!g2071) & (!g2074)) + ((g2111) & (g2118) & (!g2119) & (!g2120) & (g2071) & (!g2074)) + ((g2111) & (g2118) & (!g2119) & (g2120) & (!g2071) & (!g2074)) + ((g2111) & (g2118) & (!g2119) & (g2120) & (g2071) & (!g2074)) + ((g2111) & (g2118) & (!g2119) & (g2120) & (g2071) & (g2074)) + ((g2111) & (g2118) & (g2119) & (!g2120) & (!g2071) & (!g2074)) + ((g2111) & (g2118) & (g2119) & (!g2120) & (!g2071) & (g2074)) + ((g2111) & (g2118) & (g2119) & (!g2120) & (g2071) & (!g2074)) + ((g2111) & (g2118) & (g2119) & (g2120) & (!g2071) & (!g2074)) + ((g2111) & (g2118) & (g2119) & (g2120) & (!g2071) & (g2074)) + ((g2111) & (g2118) & (g2119) & (g2120) & (g2071) & (!g2074)) + ((g2111) & (g2118) & (g2119) & (g2120) & (g2071) & (g2074)));
	assign g2250 = (((!g2121) & (!g2083) & (!g2084) & (g2085) & (g2071) & (g2074)) + ((!g2121) & (!g2083) & (g2084) & (!g2085) & (!g2071) & (g2074)) + ((!g2121) & (!g2083) & (g2084) & (g2085) & (!g2071) & (g2074)) + ((!g2121) & (!g2083) & (g2084) & (g2085) & (g2071) & (g2074)) + ((!g2121) & (g2083) & (!g2084) & (!g2085) & (g2071) & (!g2074)) + ((!g2121) & (g2083) & (!g2084) & (g2085) & (g2071) & (!g2074)) + ((!g2121) & (g2083) & (!g2084) & (g2085) & (g2071) & (g2074)) + ((!g2121) & (g2083) & (g2084) & (!g2085) & (!g2071) & (g2074)) + ((!g2121) & (g2083) & (g2084) & (!g2085) & (g2071) & (!g2074)) + ((!g2121) & (g2083) & (g2084) & (g2085) & (!g2071) & (g2074)) + ((!g2121) & (g2083) & (g2084) & (g2085) & (g2071) & (!g2074)) + ((!g2121) & (g2083) & (g2084) & (g2085) & (g2071) & (g2074)) + ((g2121) & (!g2083) & (!g2084) & (!g2085) & (!g2071) & (!g2074)) + ((g2121) & (!g2083) & (!g2084) & (g2085) & (!g2071) & (!g2074)) + ((g2121) & (!g2083) & (!g2084) & (g2085) & (g2071) & (g2074)) + ((g2121) & (!g2083) & (g2084) & (!g2085) & (!g2071) & (!g2074)) + ((g2121) & (!g2083) & (g2084) & (!g2085) & (!g2071) & (g2074)) + ((g2121) & (!g2083) & (g2084) & (g2085) & (!g2071) & (!g2074)) + ((g2121) & (!g2083) & (g2084) & (g2085) & (!g2071) & (g2074)) + ((g2121) & (!g2083) & (g2084) & (g2085) & (g2071) & (g2074)) + ((g2121) & (g2083) & (!g2084) & (!g2085) & (!g2071) & (!g2074)) + ((g2121) & (g2083) & (!g2084) & (!g2085) & (g2071) & (!g2074)) + ((g2121) & (g2083) & (!g2084) & (g2085) & (!g2071) & (!g2074)) + ((g2121) & (g2083) & (!g2084) & (g2085) & (g2071) & (!g2074)) + ((g2121) & (g2083) & (!g2084) & (g2085) & (g2071) & (g2074)) + ((g2121) & (g2083) & (g2084) & (!g2085) & (!g2071) & (!g2074)) + ((g2121) & (g2083) & (g2084) & (!g2085) & (!g2071) & (g2074)) + ((g2121) & (g2083) & (g2084) & (!g2085) & (g2071) & (!g2074)) + ((g2121) & (g2083) & (g2084) & (g2085) & (!g2071) & (!g2074)) + ((g2121) & (g2083) & (g2084) & (g2085) & (!g2071) & (g2074)) + ((g2121) & (g2083) & (g2084) & (g2085) & (g2071) & (!g2074)) + ((g2121) & (g2083) & (g2084) & (g2085) & (g2071) & (g2074)));
	assign g2251 = (((!g2246) & (!g2248) & (!g2249) & (g2250) & (g2201) & (g2202)) + ((!g2246) & (!g2248) & (g2249) & (!g2250) & (!g2201) & (g2202)) + ((!g2246) & (!g2248) & (g2249) & (g2250) & (!g2201) & (g2202)) + ((!g2246) & (!g2248) & (g2249) & (g2250) & (g2201) & (g2202)) + ((!g2246) & (g2248) & (!g2249) & (!g2250) & (g2201) & (!g2202)) + ((!g2246) & (g2248) & (!g2249) & (g2250) & (g2201) & (!g2202)) + ((!g2246) & (g2248) & (!g2249) & (g2250) & (g2201) & (g2202)) + ((!g2246) & (g2248) & (g2249) & (!g2250) & (!g2201) & (g2202)) + ((!g2246) & (g2248) & (g2249) & (!g2250) & (g2201) & (!g2202)) + ((!g2246) & (g2248) & (g2249) & (g2250) & (!g2201) & (g2202)) + ((!g2246) & (g2248) & (g2249) & (g2250) & (g2201) & (!g2202)) + ((!g2246) & (g2248) & (g2249) & (g2250) & (g2201) & (g2202)) + ((g2246) & (!g2248) & (!g2249) & (!g2250) & (!g2201) & (!g2202)) + ((g2246) & (!g2248) & (!g2249) & (g2250) & (!g2201) & (!g2202)) + ((g2246) & (!g2248) & (!g2249) & (g2250) & (g2201) & (g2202)) + ((g2246) & (!g2248) & (g2249) & (!g2250) & (!g2201) & (!g2202)) + ((g2246) & (!g2248) & (g2249) & (!g2250) & (!g2201) & (g2202)) + ((g2246) & (!g2248) & (g2249) & (g2250) & (!g2201) & (!g2202)) + ((g2246) & (!g2248) & (g2249) & (g2250) & (!g2201) & (g2202)) + ((g2246) & (!g2248) & (g2249) & (g2250) & (g2201) & (g2202)) + ((g2246) & (g2248) & (!g2249) & (!g2250) & (!g2201) & (!g2202)) + ((g2246) & (g2248) & (!g2249) & (!g2250) & (g2201) & (!g2202)) + ((g2246) & (g2248) & (!g2249) & (g2250) & (!g2201) & (!g2202)) + ((g2246) & (g2248) & (!g2249) & (g2250) & (g2201) & (!g2202)) + ((g2246) & (g2248) & (!g2249) & (g2250) & (g2201) & (g2202)) + ((g2246) & (g2248) & (g2249) & (!g2250) & (!g2201) & (!g2202)) + ((g2246) & (g2248) & (g2249) & (!g2250) & (!g2201) & (g2202)) + ((g2246) & (g2248) & (g2249) & (!g2250) & (g2201) & (!g2202)) + ((g2246) & (g2248) & (g2249) & (g2250) & (!g2201) & (!g2202)) + ((g2246) & (g2248) & (g2249) & (g2250) & (!g2201) & (g2202)) + ((g2246) & (g2248) & (g2249) & (g2250) & (g2201) & (!g2202)) + ((g2246) & (g2248) & (g2249) & (g2250) & (g2201) & (g2202)));
	assign g2252 = (((!g2073) & (!g2080) & (!g2125) & (g2237) & (!g3751) & (!g2251)) + ((!g2073) & (!g2080) & (!g2125) & (g2237) & (!g3751) & (g2251)) + ((!g2073) & (!g2080) & (!g2125) & (g2237) & (g3751) & (!g2251)) + ((!g2073) & (!g2080) & (!g2125) & (g2237) & (g3751) & (g2251)) + ((!g2073) & (!g2080) & (g2125) & (!g2237) & (!g3751) & (g2251)) + ((!g2073) & (!g2080) & (g2125) & (!g2237) & (g3751) & (g2251)) + ((!g2073) & (!g2080) & (g2125) & (g2237) & (!g3751) & (g2251)) + ((!g2073) & (!g2080) & (g2125) & (g2237) & (g3751) & (g2251)) + ((!g2073) & (g2080) & (!g2125) & (!g2237) & (g3751) & (!g2251)) + ((!g2073) & (g2080) & (!g2125) & (!g2237) & (g3751) & (g2251)) + ((!g2073) & (g2080) & (!g2125) & (g2237) & (g3751) & (!g2251)) + ((!g2073) & (g2080) & (!g2125) & (g2237) & (g3751) & (g2251)) + ((!g2073) & (g2080) & (g2125) & (!g2237) & (g3751) & (!g2251)) + ((!g2073) & (g2080) & (g2125) & (!g2237) & (g3751) & (g2251)) + ((!g2073) & (g2080) & (g2125) & (g2237) & (g3751) & (!g2251)) + ((!g2073) & (g2080) & (g2125) & (g2237) & (g3751) & (g2251)) + ((g2073) & (!g2080) & (g2125) & (!g2237) & (!g3751) & (g2251)) + ((g2073) & (!g2080) & (g2125) & (!g2237) & (g3751) & (g2251)) + ((g2073) & (!g2080) & (g2125) & (g2237) & (!g3751) & (g2251)) + ((g2073) & (!g2080) & (g2125) & (g2237) & (g3751) & (g2251)) + ((g2073) & (g2080) & (!g2125) & (!g2237) & (g3751) & (!g2251)) + ((g2073) & (g2080) & (!g2125) & (!g2237) & (g3751) & (g2251)) + ((g2073) & (g2080) & (!g2125) & (g2237) & (g3751) & (!g2251)) + ((g2073) & (g2080) & (!g2125) & (g2237) & (g3751) & (g2251)) + ((g2073) & (g2080) & (g2125) & (!g2237) & (g3751) & (!g2251)) + ((g2073) & (g2080) & (g2125) & (!g2237) & (g3751) & (g2251)) + ((g2073) & (g2080) & (g2125) & (g2237) & (g3751) & (!g2251)) + ((g2073) & (g2080) & (g2125) & (g2237) & (g3751) & (g2251)));
	assign g2253 = (((!g2081) & (!g2124) & (!g2182) & (!g2076) & (!g2252) & (!g2106)) + ((!g2081) & (!g2124) & (!g2182) & (!g2076) & (!g2252) & (g2106)) + ((!g2081) & (!g2124) & (!g2182) & (g2076) & (!g2252) & (!g2106)) + ((!g2081) & (!g2124) & (!g2182) & (g2076) & (!g2252) & (g2106)) + ((!g2081) & (!g2124) & (g2182) & (!g2076) & (!g2252) & (!g2106)) + ((!g2081) & (!g2124) & (g2182) & (!g2076) & (g2252) & (!g2106)) + ((!g2081) & (!g2124) & (g2182) & (g2076) & (!g2252) & (!g2106)) + ((!g2081) & (!g2124) & (g2182) & (g2076) & (g2252) & (!g2106)) + ((!g2081) & (g2124) & (!g2182) & (!g2076) & (!g2252) & (!g2106)) + ((!g2081) & (g2124) & (!g2182) & (!g2076) & (g2252) & (!g2106)) + ((!g2081) & (g2124) & (g2182) & (!g2076) & (!g2252) & (!g2106)) + ((!g2081) & (g2124) & (g2182) & (!g2076) & (g2252) & (!g2106)) + ((!g2081) & (g2124) & (g2182) & (g2076) & (!g2252) & (!g2106)) + ((!g2081) & (g2124) & (g2182) & (g2076) & (g2252) & (!g2106)) + ((g2081) & (!g2124) & (!g2182) & (!g2076) & (!g2252) & (!g2106)) + ((g2081) & (!g2124) & (!g2182) & (!g2076) & (!g2252) & (g2106)) + ((g2081) & (!g2124) & (!g2182) & (g2076) & (!g2252) & (!g2106)) + ((g2081) & (!g2124) & (!g2182) & (g2076) & (!g2252) & (g2106)) + ((g2081) & (!g2124) & (g2182) & (!g2076) & (!g2252) & (!g2106)) + ((g2081) & (!g2124) & (g2182) & (!g2076) & (g2252) & (!g2106)) + ((g2081) & (!g2124) & (g2182) & (g2076) & (!g2252) & (!g2106)) + ((g2081) & (!g2124) & (g2182) & (g2076) & (g2252) & (!g2106)) + ((g2081) & (g2124) & (!g2182) & (!g2076) & (!g2252) & (!g2106)) + ((g2081) & (g2124) & (!g2182) & (!g2076) & (g2252) & (!g2106)) + ((g2081) & (g2124) & (!g2182) & (g2076) & (!g2252) & (g2106)) + ((g2081) & (g2124) & (!g2182) & (g2076) & (g2252) & (g2106)) + ((g2081) & (g2124) & (g2182) & (!g2076) & (!g2252) & (!g2106)) + ((g2081) & (g2124) & (g2182) & (!g2076) & (g2252) & (!g2106)) + ((g2081) & (g2124) & (g2182) & (g2076) & (!g2252) & (!g2106)) + ((g2081) & (g2124) & (g2182) & (g2076) & (g2252) & (!g2106)));
	assign g2254 = (((!dmem_dat_ix3x) & (!dmem_dat_ix11x) & (!dmem_dat_ix27x) & (dmem_dat_ix19x) & (g2206) & (g2207)) + ((!dmem_dat_ix3x) & (!dmem_dat_ix11x) & (dmem_dat_ix27x) & (!dmem_dat_ix19x) & (!g2206) & (g2207)) + ((!dmem_dat_ix3x) & (!dmem_dat_ix11x) & (dmem_dat_ix27x) & (dmem_dat_ix19x) & (!g2206) & (g2207)) + ((!dmem_dat_ix3x) & (!dmem_dat_ix11x) & (dmem_dat_ix27x) & (dmem_dat_ix19x) & (g2206) & (g2207)) + ((!dmem_dat_ix3x) & (dmem_dat_ix11x) & (!dmem_dat_ix27x) & (!dmem_dat_ix19x) & (g2206) & (!g2207)) + ((!dmem_dat_ix3x) & (dmem_dat_ix11x) & (!dmem_dat_ix27x) & (dmem_dat_ix19x) & (g2206) & (!g2207)) + ((!dmem_dat_ix3x) & (dmem_dat_ix11x) & (!dmem_dat_ix27x) & (dmem_dat_ix19x) & (g2206) & (g2207)) + ((!dmem_dat_ix3x) & (dmem_dat_ix11x) & (dmem_dat_ix27x) & (!dmem_dat_ix19x) & (!g2206) & (g2207)) + ((!dmem_dat_ix3x) & (dmem_dat_ix11x) & (dmem_dat_ix27x) & (!dmem_dat_ix19x) & (g2206) & (!g2207)) + ((!dmem_dat_ix3x) & (dmem_dat_ix11x) & (dmem_dat_ix27x) & (dmem_dat_ix19x) & (!g2206) & (g2207)) + ((!dmem_dat_ix3x) & (dmem_dat_ix11x) & (dmem_dat_ix27x) & (dmem_dat_ix19x) & (g2206) & (!g2207)) + ((!dmem_dat_ix3x) & (dmem_dat_ix11x) & (dmem_dat_ix27x) & (dmem_dat_ix19x) & (g2206) & (g2207)) + ((dmem_dat_ix3x) & (!dmem_dat_ix11x) & (!dmem_dat_ix27x) & (!dmem_dat_ix19x) & (!g2206) & (!g2207)) + ((dmem_dat_ix3x) & (!dmem_dat_ix11x) & (!dmem_dat_ix27x) & (dmem_dat_ix19x) & (!g2206) & (!g2207)) + ((dmem_dat_ix3x) & (!dmem_dat_ix11x) & (!dmem_dat_ix27x) & (dmem_dat_ix19x) & (g2206) & (g2207)) + ((dmem_dat_ix3x) & (!dmem_dat_ix11x) & (dmem_dat_ix27x) & (!dmem_dat_ix19x) & (!g2206) & (!g2207)) + ((dmem_dat_ix3x) & (!dmem_dat_ix11x) & (dmem_dat_ix27x) & (!dmem_dat_ix19x) & (!g2206) & (g2207)) + ((dmem_dat_ix3x) & (!dmem_dat_ix11x) & (dmem_dat_ix27x) & (dmem_dat_ix19x) & (!g2206) & (!g2207)) + ((dmem_dat_ix3x) & (!dmem_dat_ix11x) & (dmem_dat_ix27x) & (dmem_dat_ix19x) & (!g2206) & (g2207)) + ((dmem_dat_ix3x) & (!dmem_dat_ix11x) & (dmem_dat_ix27x) & (dmem_dat_ix19x) & (g2206) & (g2207)) + ((dmem_dat_ix3x) & (dmem_dat_ix11x) & (!dmem_dat_ix27x) & (!dmem_dat_ix19x) & (!g2206) & (!g2207)) + ((dmem_dat_ix3x) & (dmem_dat_ix11x) & (!dmem_dat_ix27x) & (!dmem_dat_ix19x) & (g2206) & (!g2207)) + ((dmem_dat_ix3x) & (dmem_dat_ix11x) & (!dmem_dat_ix27x) & (dmem_dat_ix19x) & (!g2206) & (!g2207)) + ((dmem_dat_ix3x) & (dmem_dat_ix11x) & (!dmem_dat_ix27x) & (dmem_dat_ix19x) & (g2206) & (!g2207)) + ((dmem_dat_ix3x) & (dmem_dat_ix11x) & (!dmem_dat_ix27x) & (dmem_dat_ix19x) & (g2206) & (g2207)) + ((dmem_dat_ix3x) & (dmem_dat_ix11x) & (dmem_dat_ix27x) & (!dmem_dat_ix19x) & (!g2206) & (!g2207)) + ((dmem_dat_ix3x) & (dmem_dat_ix11x) & (dmem_dat_ix27x) & (!dmem_dat_ix19x) & (!g2206) & (g2207)) + ((dmem_dat_ix3x) & (dmem_dat_ix11x) & (dmem_dat_ix27x) & (!dmem_dat_ix19x) & (g2206) & (!g2207)) + ((dmem_dat_ix3x) & (dmem_dat_ix11x) & (dmem_dat_ix27x) & (dmem_dat_ix19x) & (!g2206) & (!g2207)) + ((dmem_dat_ix3x) & (dmem_dat_ix11x) & (dmem_dat_ix27x) & (dmem_dat_ix19x) & (!g2206) & (g2207)) + ((dmem_dat_ix3x) & (dmem_dat_ix11x) & (dmem_dat_ix27x) & (dmem_dat_ix19x) & (g2206) & (!g2207)) + ((dmem_dat_ix3x) & (dmem_dat_ix11x) & (dmem_dat_ix27x) & (dmem_dat_ix19x) & (g2206) & (g2207)));
	assign g2255 = (((!dmem_dat_ix3x) & (!g2129) & (!sk[97]) & (dmem_dat_ix19x)) + ((!dmem_dat_ix3x) & (!g2129) & (sk[97]) & (dmem_dat_ix19x)) + ((!dmem_dat_ix3x) & (g2129) & (!sk[97]) & (!dmem_dat_ix19x)) + ((!dmem_dat_ix3x) & (g2129) & (!sk[97]) & (dmem_dat_ix19x)) + ((dmem_dat_ix3x) & (!g2129) & (!sk[97]) & (dmem_dat_ix19x)) + ((dmem_dat_ix3x) & (!g2129) & (sk[97]) & (dmem_dat_ix19x)) + ((dmem_dat_ix3x) & (g2129) & (!sk[97]) & (!dmem_dat_ix19x)) + ((dmem_dat_ix3x) & (g2129) & (!sk[97]) & (dmem_dat_ix19x)) + ((dmem_dat_ix3x) & (g2129) & (sk[97]) & (!dmem_dat_ix19x)) + ((dmem_dat_ix3x) & (g2129) & (sk[97]) & (dmem_dat_ix19x)));
	assign g2256 = (((!g75) & (!g2128) & (!g2180) & (!g2253) & (!g2254) & (!g2255)) + ((!g75) & (!g2128) & (!g2180) & (!g2253) & (!g2254) & (g2255)) + ((!g75) & (!g2128) & (!g2180) & (!g2253) & (g2254) & (!g2255)) + ((!g75) & (!g2128) & (!g2180) & (!g2253) & (g2254) & (g2255)) + ((!g75) & (!g2128) & (g2180) & (!g2253) & (!g2254) & (!g2255)) + ((!g75) & (!g2128) & (g2180) & (!g2253) & (!g2254) & (g2255)) + ((!g75) & (!g2128) & (g2180) & (!g2253) & (g2254) & (!g2255)) + ((!g75) & (!g2128) & (g2180) & (!g2253) & (g2254) & (g2255)) + ((!g75) & (g2128) & (!g2180) & (!g2253) & (!g2254) & (!g2255)) + ((!g75) & (g2128) & (!g2180) & (!g2253) & (!g2254) & (g2255)) + ((!g75) & (g2128) & (!g2180) & (!g2253) & (g2254) & (!g2255)) + ((!g75) & (g2128) & (!g2180) & (!g2253) & (g2254) & (g2255)) + ((!g75) & (g2128) & (g2180) & (!g2253) & (!g2254) & (!g2255)) + ((!g75) & (g2128) & (g2180) & (!g2253) & (!g2254) & (g2255)) + ((!g75) & (g2128) & (g2180) & (!g2253) & (g2254) & (!g2255)) + ((!g75) & (g2128) & (g2180) & (!g2253) & (g2254) & (g2255)) + ((g75) & (!g2128) & (!g2180) & (!g2253) & (g2254) & (!g2255)) + ((g75) & (!g2128) & (!g2180) & (!g2253) & (g2254) & (g2255)) + ((g75) & (!g2128) & (!g2180) & (g2253) & (g2254) & (!g2255)) + ((g75) & (!g2128) & (!g2180) & (g2253) & (g2254) & (g2255)) + ((g75) & (!g2128) & (g2180) & (!g2253) & (!g2254) & (g2255)) + ((g75) & (!g2128) & (g2180) & (!g2253) & (g2254) & (g2255)) + ((g75) & (!g2128) & (g2180) & (g2253) & (!g2254) & (g2255)) + ((g75) & (!g2128) & (g2180) & (g2253) & (g2254) & (g2255)) + ((g75) & (g2128) & (!g2180) & (!g2253) & (g2254) & (!g2255)) + ((g75) & (g2128) & (!g2180) & (!g2253) & (g2254) & (g2255)) + ((g75) & (g2128) & (!g2180) & (g2253) & (g2254) & (!g2255)) + ((g75) & (g2128) & (!g2180) & (g2253) & (g2254) & (g2255)));
	assign g2257 = (((!g141) & (!sk[99]) & (!g275) & (g319)) + ((!g141) & (!sk[99]) & (g275) & (!g319)) + ((!g141) & (!sk[99]) & (g275) & (g319)) + ((!g141) & (sk[99]) & (!g275) & (g319)) + ((!g141) & (sk[99]) & (g275) & (g319)) + ((g141) & (!sk[99]) & (!g275) & (g319)) + ((g141) & (!sk[99]) & (g275) & (!g319)) + ((g141) & (!sk[99]) & (g275) & (g319)) + ((g141) & (sk[99]) & (!g275) & (g319)) + ((g141) & (sk[99]) & (g275) & (!g319)));
	assign g5028 = (((!g2921) & (!g3057) & (!sk[100]) & (g2258)) + ((!g2921) & (!g3057) & (sk[100]) & (g2258)) + ((!g2921) & (g3057) & (!sk[100]) & (!g2258)) + ((!g2921) & (g3057) & (!sk[100]) & (g2258)) + ((!g2921) & (g3057) & (sk[100]) & (g2258)) + ((g2921) & (!g3057) & (!sk[100]) & (g2258)) + ((g2921) & (g3057) & (!sk[100]) & (!g2258)) + ((g2921) & (g3057) & (!sk[100]) & (g2258)) + ((g2921) & (g3057) & (sk[100]) & (!g2258)) + ((g2921) & (g3057) & (sk[100]) & (g2258)));
	assign g2259 = (((!g88) & (!g89) & (!sk[101]) & (!g141) & (g275)) + ((!g88) & (!g89) & (!sk[101]) & (g141) & (!g275)) + ((!g88) & (!g89) & (!sk[101]) & (g141) & (g275)) + ((!g88) & (g89) & (!sk[101]) & (!g141) & (!g275)) + ((!g88) & (g89) & (!sk[101]) & (!g141) & (g275)) + ((!g88) & (g89) & (!sk[101]) & (g141) & (!g275)) + ((!g88) & (g89) & (!sk[101]) & (g141) & (g275)) + ((!g88) & (g89) & (sk[101]) & (g141) & (g275)) + ((g88) & (!g89) & (!sk[101]) & (!g141) & (g275)) + ((g88) & (!g89) & (!sk[101]) & (g141) & (!g275)) + ((g88) & (!g89) & (!sk[101]) & (g141) & (g275)) + ((g88) & (!g89) & (sk[101]) & (!g141) & (g275)) + ((g88) & (!g89) & (sk[101]) & (g141) & (g275)) + ((g88) & (g89) & (!sk[101]) & (!g141) & (!g275)) + ((g88) & (g89) & (!sk[101]) & (!g141) & (g275)) + ((g88) & (g89) & (!sk[101]) & (g141) & (!g275)) + ((g88) & (g89) & (!sk[101]) & (g141) & (g275)) + ((g88) & (g89) & (sk[101]) & (!g141) & (g275)) + ((g88) & (g89) & (sk[101]) & (g141) & (!g275)) + ((g88) & (g89) & (sk[101]) & (g141) & (g275)));
	assign g2260 = (((!sk[102]) & (!g87) & (!g319) & (g2259)) + ((!sk[102]) & (!g87) & (g319) & (!g2259)) + ((!sk[102]) & (!g87) & (g319) & (g2259)) + ((!sk[102]) & (g87) & (!g319) & (g2259)) + ((!sk[102]) & (g87) & (g319) & (!g2259)) + ((!sk[102]) & (g87) & (g319) & (g2259)) + ((sk[102]) & (!g87) & (!g319) & (g2259)) + ((sk[102]) & (!g87) & (g319) & (!g2259)) + ((sk[102]) & (g87) & (!g319) & (!g2259)) + ((sk[102]) & (g87) & (g319) & (g2259)));
	assign g2261 = (((!sk[103]) & (!g1656) & (!g2033) & (!g2034) & (g2258) & (!g2260)) + ((!sk[103]) & (!g1656) & (!g2033) & (!g2034) & (g2258) & (g2260)) + ((!sk[103]) & (!g1656) & (!g2033) & (g2034) & (!g2258) & (!g2260)) + ((!sk[103]) & (!g1656) & (!g2033) & (g2034) & (!g2258) & (g2260)) + ((!sk[103]) & (!g1656) & (!g2033) & (g2034) & (g2258) & (!g2260)) + ((!sk[103]) & (!g1656) & (!g2033) & (g2034) & (g2258) & (g2260)) + ((!sk[103]) & (!g1656) & (g2033) & (!g2034) & (!g2258) & (!g2260)) + ((!sk[103]) & (!g1656) & (g2033) & (!g2034) & (!g2258) & (g2260)) + ((!sk[103]) & (!g1656) & (g2033) & (!g2034) & (g2258) & (!g2260)) + ((!sk[103]) & (!g1656) & (g2033) & (!g2034) & (g2258) & (g2260)) + ((!sk[103]) & (!g1656) & (g2033) & (g2034) & (!g2258) & (!g2260)) + ((!sk[103]) & (!g1656) & (g2033) & (g2034) & (!g2258) & (g2260)) + ((!sk[103]) & (!g1656) & (g2033) & (g2034) & (g2258) & (!g2260)) + ((!sk[103]) & (!g1656) & (g2033) & (g2034) & (g2258) & (g2260)) + ((!sk[103]) & (g1656) & (!g2033) & (!g2034) & (g2258) & (!g2260)) + ((!sk[103]) & (g1656) & (!g2033) & (!g2034) & (g2258) & (g2260)) + ((!sk[103]) & (g1656) & (!g2033) & (g2034) & (!g2258) & (!g2260)) + ((!sk[103]) & (g1656) & (!g2033) & (g2034) & (!g2258) & (g2260)) + ((!sk[103]) & (g1656) & (!g2033) & (g2034) & (g2258) & (!g2260)) + ((!sk[103]) & (g1656) & (!g2033) & (g2034) & (g2258) & (g2260)) + ((!sk[103]) & (g1656) & (g2033) & (!g2034) & (!g2258) & (!g2260)) + ((!sk[103]) & (g1656) & (g2033) & (!g2034) & (!g2258) & (g2260)) + ((!sk[103]) & (g1656) & (g2033) & (!g2034) & (g2258) & (!g2260)) + ((!sk[103]) & (g1656) & (g2033) & (!g2034) & (g2258) & (g2260)) + ((!sk[103]) & (g1656) & (g2033) & (g2034) & (!g2258) & (!g2260)) + ((!sk[103]) & (g1656) & (g2033) & (g2034) & (!g2258) & (g2260)) + ((!sk[103]) & (g1656) & (g2033) & (g2034) & (g2258) & (!g2260)) + ((!sk[103]) & (g1656) & (g2033) & (g2034) & (g2258) & (g2260)) + ((sk[103]) & (!g1656) & (!g2033) & (!g2034) & (g2258) & (!g2260)) + ((sk[103]) & (!g1656) & (!g2033) & (!g2034) & (g2258) & (g2260)) + ((sk[103]) & (!g1656) & (g2033) & (!g2034) & (!g2258) & (g2260)) + ((sk[103]) & (!g1656) & (g2033) & (!g2034) & (g2258) & (g2260)) + ((sk[103]) & (g1656) & (!g2033) & (!g2034) & (g2258) & (!g2260)) + ((sk[103]) & (g1656) & (!g2033) & (!g2034) & (g2258) & (g2260)) + ((sk[103]) & (g1656) & (!g2033) & (g2034) & (!g2258) & (!g2260)) + ((sk[103]) & (g1656) & (!g2033) & (g2034) & (!g2258) & (g2260)) + ((sk[103]) & (g1656) & (!g2033) & (g2034) & (g2258) & (!g2260)) + ((sk[103]) & (g1656) & (!g2033) & (g2034) & (g2258) & (g2260)) + ((sk[103]) & (g1656) & (g2033) & (!g2034) & (!g2258) & (g2260)) + ((sk[103]) & (g1656) & (g2033) & (!g2034) & (g2258) & (g2260)));
	assign g2262 = (((!g2022) & (!nmi_i) & (!g2023) & (!g2029) & (!g2257) & (g2261)) + ((!g2022) & (!nmi_i) & (!g2023) & (!g2029) & (g2257) & (g2261)) + ((!g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2257) & (!g2261)) + ((!g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2257) & (g2261)) + ((!g2022) & (!nmi_i) & (g2023) & (!g2029) & (!g2257) & (g2261)) + ((!g2022) & (!nmi_i) & (g2023) & (!g2029) & (g2257) & (g2261)) + ((!g2022) & (!nmi_i) & (g2023) & (g2029) & (g2257) & (!g2261)) + ((!g2022) & (!nmi_i) & (g2023) & (g2029) & (g2257) & (g2261)) + ((!g2022) & (nmi_i) & (!g2023) & (!g2029) & (!g2257) & (g2261)) + ((!g2022) & (nmi_i) & (!g2023) & (!g2029) & (g2257) & (g2261)) + ((!g2022) & (nmi_i) & (!g2023) & (g2029) & (g2257) & (!g2261)) + ((!g2022) & (nmi_i) & (!g2023) & (g2029) & (g2257) & (g2261)) + ((!g2022) & (nmi_i) & (g2023) & (!g2029) & (!g2257) & (g2261)) + ((!g2022) & (nmi_i) & (g2023) & (!g2029) & (g2257) & (g2261)) + ((!g2022) & (nmi_i) & (g2023) & (g2029) & (g2257) & (!g2261)) + ((!g2022) & (nmi_i) & (g2023) & (g2029) & (g2257) & (g2261)) + ((g2022) & (!nmi_i) & (!g2023) & (!g2029) & (!g2257) & (g2261)) + ((g2022) & (!nmi_i) & (!g2023) & (!g2029) & (g2257) & (g2261)) + ((g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2257) & (!g2261)) + ((g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2257) & (g2261)));
	assign g2263 = (((!g123) & (!intr_i) & (!g2039) & (!g2056) & (!g2057) & (g2262)) + ((!g123) & (!intr_i) & (!g2039) & (!g2056) & (g2057) & (g2262)) + ((!g123) & (!intr_i) & (!g2039) & (g2056) & (!g2057) & (g2262)) + ((!g123) & (!intr_i) & (!g2039) & (g2056) & (g2057) & (g2262)) + ((!g123) & (!intr_i) & (g2039) & (!g2056) & (!g2057) & (g2262)) + ((!g123) & (!intr_i) & (g2039) & (!g2056) & (g2057) & (g2262)) + ((!g123) & (!intr_i) & (g2039) & (g2056) & (!g2057) & (g2262)) + ((!g123) & (!intr_i) & (g2039) & (g2056) & (g2057) & (g2262)) + ((!g123) & (intr_i) & (!g2039) & (!g2056) & (!g2057) & (g2262)) + ((!g123) & (intr_i) & (!g2039) & (!g2056) & (g2057) & (g2262)) + ((!g123) & (intr_i) & (!g2039) & (g2056) & (!g2057) & (g2262)) + ((!g123) & (intr_i) & (g2039) & (!g2056) & (!g2057) & (g2262)) + ((!g123) & (intr_i) & (g2039) & (g2056) & (!g2057) & (g2262)));
	assign g2264 = (((!sk[106]) & (!g2080) & (!g2081) & (g2124)) + ((!sk[106]) & (!g2080) & (g2081) & (!g2124)) + ((!sk[106]) & (!g2080) & (g2081) & (g2124)) + ((!sk[106]) & (g2080) & (!g2081) & (g2124)) + ((!sk[106]) & (g2080) & (g2081) & (!g2124)) + ((!sk[106]) & (g2080) & (g2081) & (g2124)) + ((sk[106]) & (!g2080) & (g2081) & (g2124)) + ((sk[106]) & (g2080) & (!g2081) & (!g2124)) + ((sk[106]) & (g2080) & (g2081) & (!g2124)) + ((sk[106]) & (g2080) & (g2081) & (g2124)));
	assign g2265 = (((!sk[107]) & (!g2076) & (!g2106) & (g2238)) + ((!sk[107]) & (!g2076) & (g2106) & (!g2238)) + ((!sk[107]) & (!g2076) & (g2106) & (g2238)) + ((!sk[107]) & (g2076) & (!g2106) & (g2238)) + ((!sk[107]) & (g2076) & (g2106) & (!g2238)) + ((!sk[107]) & (g2076) & (g2106) & (g2238)) + ((sk[107]) & (!g2076) & (g2106) & (g2238)) + ((sk[107]) & (g2076) & (!g2106) & (g2238)) + ((sk[107]) & (g2076) & (g2106) & (!g2238)) + ((sk[107]) & (g2076) & (g2106) & (g2238)));
	assign g2266 = (((!sk[108]) & (!g2073) & (!g2113) & (g2265)) + ((!sk[108]) & (!g2073) & (g2113) & (!g2265)) + ((!sk[108]) & (!g2073) & (g2113) & (g2265)) + ((!sk[108]) & (g2073) & (!g2113) & (g2265)) + ((!sk[108]) & (g2073) & (g2113) & (!g2265)) + ((!sk[108]) & (g2073) & (g2113) & (g2265)) + ((sk[108]) & (!g2073) & (!g2113) & (g2265)) + ((sk[108]) & (!g2073) & (g2113) & (!g2265)) + ((sk[108]) & (g2073) & (!g2113) & (!g2265)) + ((sk[108]) & (g2073) & (g2113) & (g2265)));
	assign g2267 = (((!sk[109]) & (g2239) & (!g2240)) + ((!sk[109]) & (g2239) & (g2240)) + ((sk[109]) & (g2239) & (g2240)));
	assign g2268 = (((!sk[110]) & (!g2076) & (!g2106) & (g3125)) + ((!sk[110]) & (!g2076) & (g2106) & (!g3125)) + ((!sk[110]) & (!g2076) & (g2106) & (g3125)) + ((!sk[110]) & (g2076) & (!g2106) & (g3125)) + ((!sk[110]) & (g2076) & (g2106) & (!g3125)) + ((!sk[110]) & (g2076) & (g2106) & (g3125)) + ((sk[110]) & (!g2076) & (!g2106) & (!g3125)) + ((sk[110]) & (g2076) & (g2106) & (!g3125)));
	assign g2269 = (((!sk[111]) & (g2076) & (!g2106)) + ((!sk[111]) & (g2076) & (g2106)) + ((sk[111]) & (!g2076) & (g2106)));
	assign g2270 = (((!g2073) & (sk[112]) & (!g2113)) + ((g2073) & (!sk[112]) & (!g2113)) + ((g2073) & (!sk[112]) & (g2113)) + ((g2073) & (sk[112]) & (g2113)));
	assign g2271 = (((!sk[113]) & (!g2268) & (!g2269) & (g2270)) + ((!sk[113]) & (!g2268) & (g2269) & (!g2270)) + ((!sk[113]) & (!g2268) & (g2269) & (g2270)) + ((!sk[113]) & (g2268) & (!g2269) & (g2270)) + ((!sk[113]) & (g2268) & (g2269) & (!g2270)) + ((!sk[113]) & (g2268) & (g2269) & (g2270)) + ((sk[113]) & (!g2268) & (!g2269) & (g2270)) + ((sk[113]) & (!g2268) & (g2269) & (!g2270)) + ((sk[113]) & (g2268) & (!g2269) & (!g2270)) + ((sk[113]) & (g2268) & (g2269) & (g2270)));
	assign g2272 = (((!g2113) & (!g2106) & (!g2105) & (g2104) & (g2071) & (g2074)) + ((!g2113) & (!g2106) & (g2105) & (!g2104) & (!g2071) & (g2074)) + ((!g2113) & (!g2106) & (g2105) & (g2104) & (!g2071) & (g2074)) + ((!g2113) & (!g2106) & (g2105) & (g2104) & (g2071) & (g2074)) + ((!g2113) & (g2106) & (!g2105) & (!g2104) & (g2071) & (!g2074)) + ((!g2113) & (g2106) & (!g2105) & (g2104) & (g2071) & (!g2074)) + ((!g2113) & (g2106) & (!g2105) & (g2104) & (g2071) & (g2074)) + ((!g2113) & (g2106) & (g2105) & (!g2104) & (!g2071) & (g2074)) + ((!g2113) & (g2106) & (g2105) & (!g2104) & (g2071) & (!g2074)) + ((!g2113) & (g2106) & (g2105) & (g2104) & (!g2071) & (g2074)) + ((!g2113) & (g2106) & (g2105) & (g2104) & (g2071) & (!g2074)) + ((!g2113) & (g2106) & (g2105) & (g2104) & (g2071) & (g2074)) + ((g2113) & (!g2106) & (!g2105) & (!g2104) & (!g2071) & (!g2074)) + ((g2113) & (!g2106) & (!g2105) & (g2104) & (!g2071) & (!g2074)) + ((g2113) & (!g2106) & (!g2105) & (g2104) & (g2071) & (g2074)) + ((g2113) & (!g2106) & (g2105) & (!g2104) & (!g2071) & (!g2074)) + ((g2113) & (!g2106) & (g2105) & (!g2104) & (!g2071) & (g2074)) + ((g2113) & (!g2106) & (g2105) & (g2104) & (!g2071) & (!g2074)) + ((g2113) & (!g2106) & (g2105) & (g2104) & (!g2071) & (g2074)) + ((g2113) & (!g2106) & (g2105) & (g2104) & (g2071) & (g2074)) + ((g2113) & (g2106) & (!g2105) & (!g2104) & (!g2071) & (!g2074)) + ((g2113) & (g2106) & (!g2105) & (!g2104) & (g2071) & (!g2074)) + ((g2113) & (g2106) & (!g2105) & (g2104) & (!g2071) & (!g2074)) + ((g2113) & (g2106) & (!g2105) & (g2104) & (g2071) & (!g2074)) + ((g2113) & (g2106) & (!g2105) & (g2104) & (g2071) & (g2074)) + ((g2113) & (g2106) & (g2105) & (!g2104) & (!g2071) & (!g2074)) + ((g2113) & (g2106) & (g2105) & (!g2104) & (!g2071) & (g2074)) + ((g2113) & (g2106) & (g2105) & (!g2104) & (g2071) & (!g2074)) + ((g2113) & (g2106) & (g2105) & (g2104) & (!g2071) & (!g2074)) + ((g2113) & (g2106) & (g2105) & (g2104) & (!g2071) & (g2074)) + ((g2113) & (g2106) & (g2105) & (g2104) & (g2071) & (!g2074)) + ((g2113) & (g2106) & (g2105) & (g2104) & (g2071) & (g2074)));
	assign g2273 = (((!sk[115]) & (!g2075) & (!g2076) & (!g2077) & (g2272)) + ((!sk[115]) & (!g2075) & (!g2076) & (g2077) & (!g2272)) + ((!sk[115]) & (!g2075) & (!g2076) & (g2077) & (g2272)) + ((!sk[115]) & (!g2075) & (g2076) & (!g2077) & (!g2272)) + ((!sk[115]) & (!g2075) & (g2076) & (!g2077) & (g2272)) + ((!sk[115]) & (!g2075) & (g2076) & (g2077) & (!g2272)) + ((!sk[115]) & (!g2075) & (g2076) & (g2077) & (g2272)) + ((!sk[115]) & (g2075) & (!g2076) & (!g2077) & (g2272)) + ((!sk[115]) & (g2075) & (!g2076) & (g2077) & (!g2272)) + ((!sk[115]) & (g2075) & (!g2076) & (g2077) & (g2272)) + ((!sk[115]) & (g2075) & (g2076) & (!g2077) & (!g2272)) + ((!sk[115]) & (g2075) & (g2076) & (!g2077) & (g2272)) + ((!sk[115]) & (g2075) & (g2076) & (g2077) & (!g2272)) + ((!sk[115]) & (g2075) & (g2076) & (g2077) & (g2272)) + ((sk[115]) & (!g2075) & (!g2076) & (!g2077) & (g2272)) + ((sk[115]) & (g2075) & (!g2076) & (!g2077) & (g2272)) + ((sk[115]) & (g2075) & (!g2076) & (g2077) & (!g2272)) + ((sk[115]) & (g2075) & (!g2076) & (g2077) & (g2272)));
	assign g2274 = (((!g2097) & (!g2102) & (!g2092) & (g2192) & (g2076) & (g2077)) + ((!g2097) & (!g2102) & (g2092) & (!g2192) & (!g2076) & (g2077)) + ((!g2097) & (!g2102) & (g2092) & (g2192) & (!g2076) & (g2077)) + ((!g2097) & (!g2102) & (g2092) & (g2192) & (g2076) & (g2077)) + ((!g2097) & (g2102) & (!g2092) & (!g2192) & (g2076) & (!g2077)) + ((!g2097) & (g2102) & (!g2092) & (g2192) & (g2076) & (!g2077)) + ((!g2097) & (g2102) & (!g2092) & (g2192) & (g2076) & (g2077)) + ((!g2097) & (g2102) & (g2092) & (!g2192) & (!g2076) & (g2077)) + ((!g2097) & (g2102) & (g2092) & (!g2192) & (g2076) & (!g2077)) + ((!g2097) & (g2102) & (g2092) & (g2192) & (!g2076) & (g2077)) + ((!g2097) & (g2102) & (g2092) & (g2192) & (g2076) & (!g2077)) + ((!g2097) & (g2102) & (g2092) & (g2192) & (g2076) & (g2077)) + ((g2097) & (!g2102) & (!g2092) & (!g2192) & (!g2076) & (!g2077)) + ((g2097) & (!g2102) & (!g2092) & (g2192) & (!g2076) & (!g2077)) + ((g2097) & (!g2102) & (!g2092) & (g2192) & (g2076) & (g2077)) + ((g2097) & (!g2102) & (g2092) & (!g2192) & (!g2076) & (!g2077)) + ((g2097) & (!g2102) & (g2092) & (!g2192) & (!g2076) & (g2077)) + ((g2097) & (!g2102) & (g2092) & (g2192) & (!g2076) & (!g2077)) + ((g2097) & (!g2102) & (g2092) & (g2192) & (!g2076) & (g2077)) + ((g2097) & (!g2102) & (g2092) & (g2192) & (g2076) & (g2077)) + ((g2097) & (g2102) & (!g2092) & (!g2192) & (!g2076) & (!g2077)) + ((g2097) & (g2102) & (!g2092) & (!g2192) & (g2076) & (!g2077)) + ((g2097) & (g2102) & (!g2092) & (g2192) & (!g2076) & (!g2077)) + ((g2097) & (g2102) & (!g2092) & (g2192) & (g2076) & (!g2077)) + ((g2097) & (g2102) & (!g2092) & (g2192) & (g2076) & (g2077)) + ((g2097) & (g2102) & (g2092) & (!g2192) & (!g2076) & (!g2077)) + ((g2097) & (g2102) & (g2092) & (!g2192) & (!g2076) & (g2077)) + ((g2097) & (g2102) & (g2092) & (!g2192) & (g2076) & (!g2077)) + ((g2097) & (g2102) & (g2092) & (g2192) & (!g2076) & (!g2077)) + ((g2097) & (g2102) & (g2092) & (g2192) & (!g2076) & (g2077)) + ((g2097) & (g2102) & (g2092) & (g2192) & (g2076) & (!g2077)) + ((g2097) & (g2102) & (g2092) & (g2192) & (g2076) & (g2077)));
	assign g2275 = (((!g2117) & (!g2122) & (!g2112) & (g2087) & (g2076) & (g2077)) + ((!g2117) & (!g2122) & (g2112) & (!g2087) & (!g2076) & (g2077)) + ((!g2117) & (!g2122) & (g2112) & (g2087) & (!g2076) & (g2077)) + ((!g2117) & (!g2122) & (g2112) & (g2087) & (g2076) & (g2077)) + ((!g2117) & (g2122) & (!g2112) & (!g2087) & (g2076) & (!g2077)) + ((!g2117) & (g2122) & (!g2112) & (g2087) & (g2076) & (!g2077)) + ((!g2117) & (g2122) & (!g2112) & (g2087) & (g2076) & (g2077)) + ((!g2117) & (g2122) & (g2112) & (!g2087) & (!g2076) & (g2077)) + ((!g2117) & (g2122) & (g2112) & (!g2087) & (g2076) & (!g2077)) + ((!g2117) & (g2122) & (g2112) & (g2087) & (!g2076) & (g2077)) + ((!g2117) & (g2122) & (g2112) & (g2087) & (g2076) & (!g2077)) + ((!g2117) & (g2122) & (g2112) & (g2087) & (g2076) & (g2077)) + ((g2117) & (!g2122) & (!g2112) & (!g2087) & (!g2076) & (!g2077)) + ((g2117) & (!g2122) & (!g2112) & (g2087) & (!g2076) & (!g2077)) + ((g2117) & (!g2122) & (!g2112) & (g2087) & (g2076) & (g2077)) + ((g2117) & (!g2122) & (g2112) & (!g2087) & (!g2076) & (!g2077)) + ((g2117) & (!g2122) & (g2112) & (!g2087) & (!g2076) & (g2077)) + ((g2117) & (!g2122) & (g2112) & (g2087) & (!g2076) & (!g2077)) + ((g2117) & (!g2122) & (g2112) & (g2087) & (!g2076) & (g2077)) + ((g2117) & (!g2122) & (g2112) & (g2087) & (g2076) & (g2077)) + ((g2117) & (g2122) & (!g2112) & (!g2087) & (!g2076) & (!g2077)) + ((g2117) & (g2122) & (!g2112) & (!g2087) & (g2076) & (!g2077)) + ((g2117) & (g2122) & (!g2112) & (g2087) & (!g2076) & (!g2077)) + ((g2117) & (g2122) & (!g2112) & (g2087) & (g2076) & (!g2077)) + ((g2117) & (g2122) & (!g2112) & (g2087) & (g2076) & (g2077)) + ((g2117) & (g2122) & (g2112) & (!g2087) & (!g2076) & (!g2077)) + ((g2117) & (g2122) & (g2112) & (!g2087) & (!g2076) & (g2077)) + ((g2117) & (g2122) & (g2112) & (!g2087) & (g2076) & (!g2077)) + ((g2117) & (g2122) & (g2112) & (g2087) & (!g2076) & (!g2077)) + ((g2117) & (g2122) & (g2112) & (g2087) & (!g2076) & (g2077)) + ((g2117) & (g2122) & (g2112) & (g2087) & (g2076) & (!g2077)) + ((g2117) & (g2122) & (g2112) & (g2087) & (g2076) & (g2077)));
	assign g2276 = (((!g2073) & (!g2080) & (!g2125) & (g2273) & (!g2274) & (!g2275)) + ((!g2073) & (!g2080) & (!g2125) & (g2273) & (!g2274) & (g2275)) + ((!g2073) & (!g2080) & (!g2125) & (g2273) & (g2274) & (!g2275)) + ((!g2073) & (!g2080) & (!g2125) & (g2273) & (g2274) & (g2275)) + ((!g2073) & (!g2080) & (g2125) & (!g2273) & (!g2274) & (g2275)) + ((!g2073) & (!g2080) & (g2125) & (!g2273) & (g2274) & (g2275)) + ((!g2073) & (!g2080) & (g2125) & (g2273) & (!g2274) & (g2275)) + ((!g2073) & (!g2080) & (g2125) & (g2273) & (g2274) & (g2275)) + ((!g2073) & (g2080) & (!g2125) & (g2273) & (!g2274) & (!g2275)) + ((!g2073) & (g2080) & (!g2125) & (g2273) & (!g2274) & (g2275)) + ((!g2073) & (g2080) & (!g2125) & (g2273) & (g2274) & (!g2275)) + ((!g2073) & (g2080) & (!g2125) & (g2273) & (g2274) & (g2275)) + ((!g2073) & (g2080) & (g2125) & (!g2273) & (!g2274) & (g2275)) + ((!g2073) & (g2080) & (g2125) & (!g2273) & (g2274) & (g2275)) + ((!g2073) & (g2080) & (g2125) & (g2273) & (!g2274) & (g2275)) + ((!g2073) & (g2080) & (g2125) & (g2273) & (g2274) & (g2275)) + ((g2073) & (!g2080) & (g2125) & (!g2273) & (g2274) & (!g2275)) + ((g2073) & (!g2080) & (g2125) & (!g2273) & (g2274) & (g2275)) + ((g2073) & (!g2080) & (g2125) & (g2273) & (g2274) & (!g2275)) + ((g2073) & (!g2080) & (g2125) & (g2273) & (g2274) & (g2275)) + ((g2073) & (g2080) & (!g2125) & (g2273) & (!g2274) & (!g2275)) + ((g2073) & (g2080) & (!g2125) & (g2273) & (!g2274) & (g2275)) + ((g2073) & (g2080) & (!g2125) & (g2273) & (g2274) & (!g2275)) + ((g2073) & (g2080) & (!g2125) & (g2273) & (g2274) & (g2275)) + ((g2073) & (g2080) & (g2125) & (!g2273) & (g2274) & (!g2275)) + ((g2073) & (g2080) & (g2125) & (!g2273) & (g2274) & (g2275)) + ((g2073) & (g2080) & (g2125) & (g2273) & (g2274) & (!g2275)) + ((g2073) & (g2080) & (g2125) & (g2273) & (g2274) & (g2275)));
	assign g2277 = (((!g2113) & (!g2073) & (!g2124) & (!g2264) & (!g3738) & (!g2276)) + ((!g2113) & (!g2073) & (!g2124) & (!g2264) & (g3738) & (!g2276)) + ((!g2113) & (!g2073) & (!g2124) & (g2264) & (!g3738) & (!g2276)) + ((!g2113) & (!g2073) & (!g2124) & (g2264) & (!g3738) & (g2276)) + ((!g2113) & (!g2073) & (g2124) & (!g2264) & (!g3738) & (!g2276)) + ((!g2113) & (!g2073) & (g2124) & (!g2264) & (!g3738) & (g2276)) + ((!g2113) & (!g2073) & (g2124) & (!g2264) & (g3738) & (!g2276)) + ((!g2113) & (!g2073) & (g2124) & (!g2264) & (g3738) & (g2276)) + ((!g2113) & (!g2073) & (g2124) & (g2264) & (!g3738) & (!g2276)) + ((!g2113) & (!g2073) & (g2124) & (g2264) & (!g3738) & (g2276)) + ((!g2113) & (!g2073) & (g2124) & (g2264) & (g3738) & (!g2276)) + ((!g2113) & (!g2073) & (g2124) & (g2264) & (g3738) & (g2276)) + ((!g2113) & (g2073) & (!g2124) & (!g2264) & (!g3738) & (!g2276)) + ((!g2113) & (g2073) & (!g2124) & (!g2264) & (g3738) & (!g2276)) + ((!g2113) & (g2073) & (!g2124) & (g2264) & (!g3738) & (!g2276)) + ((!g2113) & (g2073) & (!g2124) & (g2264) & (!g3738) & (g2276)) + ((g2113) & (!g2073) & (!g2124) & (!g2264) & (!g3738) & (!g2276)) + ((g2113) & (!g2073) & (!g2124) & (!g2264) & (g3738) & (!g2276)) + ((g2113) & (!g2073) & (!g2124) & (g2264) & (!g3738) & (!g2276)) + ((g2113) & (!g2073) & (!g2124) & (g2264) & (!g3738) & (g2276)) + ((g2113) & (g2073) & (!g2124) & (!g2264) & (!g3738) & (!g2276)) + ((g2113) & (g2073) & (!g2124) & (!g2264) & (g3738) & (!g2276)) + ((g2113) & (g2073) & (!g2124) & (g2264) & (!g3738) & (!g2276)) + ((g2113) & (g2073) & (!g2124) & (g2264) & (!g3738) & (g2276)) + ((g2113) & (g2073) & (g2124) & (g2264) & (!g3738) & (!g2276)) + ((g2113) & (g2073) & (g2124) & (g2264) & (!g3738) & (g2276)) + ((g2113) & (g2073) & (g2124) & (g2264) & (g3738) & (!g2276)) + ((g2113) & (g2073) & (g2124) & (g2264) & (g3738) & (g2276)));
	assign g2278 = (((!dmem_dat_ix4x) & (!dmem_dat_ix12x) & (!dmem_dat_ix28x) & (dmem_dat_ix20x) & (g2206) & (g2207)) + ((!dmem_dat_ix4x) & (!dmem_dat_ix12x) & (dmem_dat_ix28x) & (!dmem_dat_ix20x) & (!g2206) & (g2207)) + ((!dmem_dat_ix4x) & (!dmem_dat_ix12x) & (dmem_dat_ix28x) & (dmem_dat_ix20x) & (!g2206) & (g2207)) + ((!dmem_dat_ix4x) & (!dmem_dat_ix12x) & (dmem_dat_ix28x) & (dmem_dat_ix20x) & (g2206) & (g2207)) + ((!dmem_dat_ix4x) & (dmem_dat_ix12x) & (!dmem_dat_ix28x) & (!dmem_dat_ix20x) & (g2206) & (!g2207)) + ((!dmem_dat_ix4x) & (dmem_dat_ix12x) & (!dmem_dat_ix28x) & (dmem_dat_ix20x) & (g2206) & (!g2207)) + ((!dmem_dat_ix4x) & (dmem_dat_ix12x) & (!dmem_dat_ix28x) & (dmem_dat_ix20x) & (g2206) & (g2207)) + ((!dmem_dat_ix4x) & (dmem_dat_ix12x) & (dmem_dat_ix28x) & (!dmem_dat_ix20x) & (!g2206) & (g2207)) + ((!dmem_dat_ix4x) & (dmem_dat_ix12x) & (dmem_dat_ix28x) & (!dmem_dat_ix20x) & (g2206) & (!g2207)) + ((!dmem_dat_ix4x) & (dmem_dat_ix12x) & (dmem_dat_ix28x) & (dmem_dat_ix20x) & (!g2206) & (g2207)) + ((!dmem_dat_ix4x) & (dmem_dat_ix12x) & (dmem_dat_ix28x) & (dmem_dat_ix20x) & (g2206) & (!g2207)) + ((!dmem_dat_ix4x) & (dmem_dat_ix12x) & (dmem_dat_ix28x) & (dmem_dat_ix20x) & (g2206) & (g2207)) + ((dmem_dat_ix4x) & (!dmem_dat_ix12x) & (!dmem_dat_ix28x) & (!dmem_dat_ix20x) & (!g2206) & (!g2207)) + ((dmem_dat_ix4x) & (!dmem_dat_ix12x) & (!dmem_dat_ix28x) & (dmem_dat_ix20x) & (!g2206) & (!g2207)) + ((dmem_dat_ix4x) & (!dmem_dat_ix12x) & (!dmem_dat_ix28x) & (dmem_dat_ix20x) & (g2206) & (g2207)) + ((dmem_dat_ix4x) & (!dmem_dat_ix12x) & (dmem_dat_ix28x) & (!dmem_dat_ix20x) & (!g2206) & (!g2207)) + ((dmem_dat_ix4x) & (!dmem_dat_ix12x) & (dmem_dat_ix28x) & (!dmem_dat_ix20x) & (!g2206) & (g2207)) + ((dmem_dat_ix4x) & (!dmem_dat_ix12x) & (dmem_dat_ix28x) & (dmem_dat_ix20x) & (!g2206) & (!g2207)) + ((dmem_dat_ix4x) & (!dmem_dat_ix12x) & (dmem_dat_ix28x) & (dmem_dat_ix20x) & (!g2206) & (g2207)) + ((dmem_dat_ix4x) & (!dmem_dat_ix12x) & (dmem_dat_ix28x) & (dmem_dat_ix20x) & (g2206) & (g2207)) + ((dmem_dat_ix4x) & (dmem_dat_ix12x) & (!dmem_dat_ix28x) & (!dmem_dat_ix20x) & (!g2206) & (!g2207)) + ((dmem_dat_ix4x) & (dmem_dat_ix12x) & (!dmem_dat_ix28x) & (!dmem_dat_ix20x) & (g2206) & (!g2207)) + ((dmem_dat_ix4x) & (dmem_dat_ix12x) & (!dmem_dat_ix28x) & (dmem_dat_ix20x) & (!g2206) & (!g2207)) + ((dmem_dat_ix4x) & (dmem_dat_ix12x) & (!dmem_dat_ix28x) & (dmem_dat_ix20x) & (g2206) & (!g2207)) + ((dmem_dat_ix4x) & (dmem_dat_ix12x) & (!dmem_dat_ix28x) & (dmem_dat_ix20x) & (g2206) & (g2207)) + ((dmem_dat_ix4x) & (dmem_dat_ix12x) & (dmem_dat_ix28x) & (!dmem_dat_ix20x) & (!g2206) & (!g2207)) + ((dmem_dat_ix4x) & (dmem_dat_ix12x) & (dmem_dat_ix28x) & (!dmem_dat_ix20x) & (!g2206) & (g2207)) + ((dmem_dat_ix4x) & (dmem_dat_ix12x) & (dmem_dat_ix28x) & (!dmem_dat_ix20x) & (g2206) & (!g2207)) + ((dmem_dat_ix4x) & (dmem_dat_ix12x) & (dmem_dat_ix28x) & (dmem_dat_ix20x) & (!g2206) & (!g2207)) + ((dmem_dat_ix4x) & (dmem_dat_ix12x) & (dmem_dat_ix28x) & (dmem_dat_ix20x) & (!g2206) & (g2207)) + ((dmem_dat_ix4x) & (dmem_dat_ix12x) & (dmem_dat_ix28x) & (dmem_dat_ix20x) & (g2206) & (!g2207)) + ((dmem_dat_ix4x) & (dmem_dat_ix12x) & (dmem_dat_ix28x) & (dmem_dat_ix20x) & (g2206) & (g2207)));
	assign g2279 = (((!g2128) & (!g2129) & (!sk[121]) & (!dmem_dat_ix4x) & (dmem_dat_ix20x)) + ((!g2128) & (!g2129) & (!sk[121]) & (dmem_dat_ix4x) & (!dmem_dat_ix20x)) + ((!g2128) & (!g2129) & (!sk[121]) & (dmem_dat_ix4x) & (dmem_dat_ix20x)) + ((!g2128) & (!g2129) & (sk[121]) & (!dmem_dat_ix4x) & (dmem_dat_ix20x)) + ((!g2128) & (!g2129) & (sk[121]) & (dmem_dat_ix4x) & (dmem_dat_ix20x)) + ((!g2128) & (g2129) & (!sk[121]) & (!dmem_dat_ix4x) & (!dmem_dat_ix20x)) + ((!g2128) & (g2129) & (!sk[121]) & (!dmem_dat_ix4x) & (dmem_dat_ix20x)) + ((!g2128) & (g2129) & (!sk[121]) & (dmem_dat_ix4x) & (!dmem_dat_ix20x)) + ((!g2128) & (g2129) & (!sk[121]) & (dmem_dat_ix4x) & (dmem_dat_ix20x)) + ((!g2128) & (g2129) & (sk[121]) & (dmem_dat_ix4x) & (!dmem_dat_ix20x)) + ((!g2128) & (g2129) & (sk[121]) & (dmem_dat_ix4x) & (dmem_dat_ix20x)) + ((g2128) & (!g2129) & (!sk[121]) & (!dmem_dat_ix4x) & (dmem_dat_ix20x)) + ((g2128) & (!g2129) & (!sk[121]) & (dmem_dat_ix4x) & (!dmem_dat_ix20x)) + ((g2128) & (!g2129) & (!sk[121]) & (dmem_dat_ix4x) & (dmem_dat_ix20x)) + ((g2128) & (g2129) & (!sk[121]) & (!dmem_dat_ix4x) & (!dmem_dat_ix20x)) + ((g2128) & (g2129) & (!sk[121]) & (!dmem_dat_ix4x) & (dmem_dat_ix20x)) + ((g2128) & (g2129) & (!sk[121]) & (dmem_dat_ix4x) & (!dmem_dat_ix20x)) + ((g2128) & (g2129) & (!sk[121]) & (dmem_dat_ix4x) & (dmem_dat_ix20x)));
	assign g2280 = (((!sk[122]) & (!g2080) & (!g2081) & (!g2124) & (g2125)) + ((!sk[122]) & (!g2080) & (!g2081) & (g2124) & (!g2125)) + ((!sk[122]) & (!g2080) & (!g2081) & (g2124) & (g2125)) + ((!sk[122]) & (!g2080) & (g2081) & (!g2124) & (!g2125)) + ((!sk[122]) & (!g2080) & (g2081) & (!g2124) & (g2125)) + ((!sk[122]) & (!g2080) & (g2081) & (g2124) & (!g2125)) + ((!sk[122]) & (!g2080) & (g2081) & (g2124) & (g2125)) + ((!sk[122]) & (g2080) & (!g2081) & (!g2124) & (g2125)) + ((!sk[122]) & (g2080) & (!g2081) & (g2124) & (!g2125)) + ((!sk[122]) & (g2080) & (!g2081) & (g2124) & (g2125)) + ((!sk[122]) & (g2080) & (g2081) & (!g2124) & (!g2125)) + ((!sk[122]) & (g2080) & (g2081) & (!g2124) & (g2125)) + ((!sk[122]) & (g2080) & (g2081) & (g2124) & (!g2125)) + ((!sk[122]) & (g2080) & (g2081) & (g2124) & (g2125)) + ((sk[122]) & (!g2080) & (!g2081) & (!g2124) & (!g2125)) + ((sk[122]) & (!g2080) & (!g2081) & (g2124) & (g2125)) + ((sk[122]) & (!g2080) & (g2081) & (g2124) & (g2125)) + ((sk[122]) & (g2080) & (!g2081) & (g2124) & (!g2125)) + ((sk[122]) & (g2080) & (!g2081) & (g2124) & (g2125)) + ((sk[122]) & (g2080) & (g2081) & (g2124) & (!g2125)) + ((sk[122]) & (g2080) & (g2081) & (g2124) & (g2125)));
	assign g2281 = (((!g75) & (!g2180) & (!sk[123]) & (g2280)) + ((!g75) & (!g2180) & (sk[123]) & (g2280)) + ((!g75) & (g2180) & (!sk[123]) & (!g2280)) + ((!g75) & (g2180) & (!sk[123]) & (g2280)) + ((!g75) & (g2180) & (sk[123]) & (g2280)) + ((g75) & (!g2180) & (!sk[123]) & (g2280)) + ((g75) & (g2180) & (!sk[123]) & (!g2280)) + ((g75) & (g2180) & (!sk[123]) & (g2280)) + ((g75) & (g2180) & (sk[123]) & (!g2280)) + ((g75) & (g2180) & (sk[123]) & (g2280)));
	assign g2282 = (((!g2277) & (!g2113) & (!g2278) & (!g2279) & (!g2281) & (!g75)) + ((!g2277) & (!g2113) & (!g2278) & (g2279) & (!g2281) & (!g75)) + ((!g2277) & (!g2113) & (!g2278) & (g2279) & (g2281) & (g75)) + ((!g2277) & (!g2113) & (g2278) & (!g2279) & (!g2281) & (!g75)) + ((!g2277) & (!g2113) & (g2278) & (!g2279) & (!g2281) & (g75)) + ((!g2277) & (!g2113) & (g2278) & (g2279) & (!g2281) & (!g75)) + ((!g2277) & (!g2113) & (g2278) & (g2279) & (!g2281) & (g75)) + ((!g2277) & (!g2113) & (g2278) & (g2279) & (g2281) & (g75)) + ((!g2277) & (g2113) & (!g2278) & (!g2279) & (!g2281) & (!g75)) + ((!g2277) & (g2113) & (!g2278) & (!g2279) & (g2281) & (!g75)) + ((!g2277) & (g2113) & (!g2278) & (g2279) & (!g2281) & (!g75)) + ((!g2277) & (g2113) & (!g2278) & (g2279) & (g2281) & (!g75)) + ((!g2277) & (g2113) & (!g2278) & (g2279) & (g2281) & (g75)) + ((!g2277) & (g2113) & (g2278) & (!g2279) & (!g2281) & (!g75)) + ((!g2277) & (g2113) & (g2278) & (!g2279) & (!g2281) & (g75)) + ((!g2277) & (g2113) & (g2278) & (!g2279) & (g2281) & (!g75)) + ((!g2277) & (g2113) & (g2278) & (g2279) & (!g2281) & (!g75)) + ((!g2277) & (g2113) & (g2278) & (g2279) & (!g2281) & (g75)) + ((!g2277) & (g2113) & (g2278) & (g2279) & (g2281) & (!g75)) + ((!g2277) & (g2113) & (g2278) & (g2279) & (g2281) & (g75)) + ((g2277) & (!g2113) & (!g2278) & (g2279) & (g2281) & (g75)) + ((g2277) & (!g2113) & (g2278) & (!g2279) & (!g2281) & (g75)) + ((g2277) & (!g2113) & (g2278) & (g2279) & (!g2281) & (g75)) + ((g2277) & (!g2113) & (g2278) & (g2279) & (g2281) & (g75)) + ((g2277) & (g2113) & (!g2278) & (!g2279) & (g2281) & (!g75)) + ((g2277) & (g2113) & (!g2278) & (g2279) & (g2281) & (!g75)) + ((g2277) & (g2113) & (!g2278) & (g2279) & (g2281) & (g75)) + ((g2277) & (g2113) & (g2278) & (!g2279) & (!g2281) & (g75)) + ((g2277) & (g2113) & (g2278) & (!g2279) & (g2281) & (!g75)) + ((g2277) & (g2113) & (g2278) & (g2279) & (!g2281) & (g75)) + ((g2277) & (g2113) & (g2278) & (g2279) & (g2281) & (!g75)) + ((g2277) & (g2113) & (g2278) & (g2279) & (g2281) & (g75)));
	assign g2283 = (((!g141) & (!g275) & (!g319) & (!sk[125]) & (g365)) + ((!g141) & (!g275) & (!g319) & (sk[125]) & (g365)) + ((!g141) & (!g275) & (g319) & (!sk[125]) & (!g365)) + ((!g141) & (!g275) & (g319) & (!sk[125]) & (g365)) + ((!g141) & (!g275) & (g319) & (sk[125]) & (g365)) + ((!g141) & (g275) & (!g319) & (!sk[125]) & (!g365)) + ((!g141) & (g275) & (!g319) & (!sk[125]) & (g365)) + ((!g141) & (g275) & (!g319) & (sk[125]) & (g365)) + ((!g141) & (g275) & (g319) & (!sk[125]) & (!g365)) + ((!g141) & (g275) & (g319) & (!sk[125]) & (g365)) + ((!g141) & (g275) & (g319) & (sk[125]) & (g365)) + ((g141) & (!g275) & (!g319) & (!sk[125]) & (g365)) + ((g141) & (!g275) & (!g319) & (sk[125]) & (g365)) + ((g141) & (!g275) & (g319) & (!sk[125]) & (!g365)) + ((g141) & (!g275) & (g319) & (!sk[125]) & (g365)) + ((g141) & (!g275) & (g319) & (sk[125]) & (g365)) + ((g141) & (g275) & (!g319) & (!sk[125]) & (!g365)) + ((g141) & (g275) & (!g319) & (!sk[125]) & (g365)) + ((g141) & (g275) & (!g319) & (sk[125]) & (g365)) + ((g141) & (g275) & (g319) & (!sk[125]) & (!g365)) + ((g141) & (g275) & (g319) & (!sk[125]) & (g365)) + ((g141) & (g275) & (g319) & (sk[125]) & (!g365)));
	assign g5029 = (((!sk[126]) & (!g2921) & (!g3058) & (g2284)) + ((!sk[126]) & (!g2921) & (g3058) & (!g2284)) + ((!sk[126]) & (!g2921) & (g3058) & (g2284)) + ((!sk[126]) & (g2921) & (!g3058) & (g2284)) + ((!sk[126]) & (g2921) & (g3058) & (!g2284)) + ((!sk[126]) & (g2921) & (g3058) & (g2284)) + ((sk[126]) & (!g2921) & (!g3058) & (g2284)) + ((sk[126]) & (!g2921) & (g3058) & (g2284)) + ((sk[126]) & (g2921) & (g3058) & (!g2284)) + ((sk[126]) & (g2921) & (g3058) & (g2284)));
	assign g2285 = (((!g87) & (!sk[127]) & (!g90) & (!g319) & (g2259) & (!g365)) + ((!g87) & (!sk[127]) & (!g90) & (!g319) & (g2259) & (g365)) + ((!g87) & (!sk[127]) & (!g90) & (g319) & (!g2259) & (!g365)) + ((!g87) & (!sk[127]) & (!g90) & (g319) & (!g2259) & (g365)) + ((!g87) & (!sk[127]) & (!g90) & (g319) & (g2259) & (!g365)) + ((!g87) & (!sk[127]) & (!g90) & (g319) & (g2259) & (g365)) + ((!g87) & (!sk[127]) & (g90) & (!g319) & (!g2259) & (!g365)) + ((!g87) & (!sk[127]) & (g90) & (!g319) & (!g2259) & (g365)) + ((!g87) & (!sk[127]) & (g90) & (!g319) & (g2259) & (!g365)) + ((!g87) & (!sk[127]) & (g90) & (!g319) & (g2259) & (g365)) + ((!g87) & (!sk[127]) & (g90) & (g319) & (!g2259) & (!g365)) + ((!g87) & (!sk[127]) & (g90) & (g319) & (!g2259) & (g365)) + ((!g87) & (!sk[127]) & (g90) & (g319) & (g2259) & (!g365)) + ((!g87) & (!sk[127]) & (g90) & (g319) & (g2259) & (g365)) + ((!g87) & (sk[127]) & (!g90) & (!g319) & (!g2259) & (g365)) + ((!g87) & (sk[127]) & (!g90) & (!g319) & (g2259) & (g365)) + ((!g87) & (sk[127]) & (!g90) & (g319) & (!g2259) & (g365)) + ((!g87) & (sk[127]) & (!g90) & (g319) & (g2259) & (!g365)) + ((!g87) & (sk[127]) & (g90) & (!g319) & (!g2259) & (!g365)) + ((!g87) & (sk[127]) & (g90) & (!g319) & (g2259) & (!g365)) + ((!g87) & (sk[127]) & (g90) & (g319) & (!g2259) & (!g365)) + ((!g87) & (sk[127]) & (g90) & (g319) & (g2259) & (g365)) + ((g87) & (!sk[127]) & (!g90) & (!g319) & (g2259) & (!g365)) + ((g87) & (!sk[127]) & (!g90) & (!g319) & (g2259) & (g365)) + ((g87) & (!sk[127]) & (!g90) & (g319) & (!g2259) & (!g365)) + ((g87) & (!sk[127]) & (!g90) & (g319) & (!g2259) & (g365)) + ((g87) & (!sk[127]) & (!g90) & (g319) & (g2259) & (!g365)) + ((g87) & (!sk[127]) & (!g90) & (g319) & (g2259) & (g365)) + ((g87) & (!sk[127]) & (g90) & (!g319) & (!g2259) & (!g365)) + ((g87) & (!sk[127]) & (g90) & (!g319) & (!g2259) & (g365)) + ((g87) & (!sk[127]) & (g90) & (!g319) & (g2259) & (!g365)) + ((g87) & (!sk[127]) & (g90) & (!g319) & (g2259) & (g365)) + ((g87) & (!sk[127]) & (g90) & (g319) & (!g2259) & (!g365)) + ((g87) & (!sk[127]) & (g90) & (g319) & (!g2259) & (g365)) + ((g87) & (!sk[127]) & (g90) & (g319) & (g2259) & (!g365)) + ((g87) & (!sk[127]) & (g90) & (g319) & (g2259) & (g365)) + ((g87) & (sk[127]) & (!g90) & (!g319) & (!g2259) & (g365)) + ((g87) & (sk[127]) & (!g90) & (!g319) & (g2259) & (!g365)) + ((g87) & (sk[127]) & (!g90) & (g319) & (!g2259) & (!g365)) + ((g87) & (sk[127]) & (!g90) & (g319) & (g2259) & (!g365)) + ((g87) & (sk[127]) & (g90) & (!g319) & (!g2259) & (!g365)) + ((g87) & (sk[127]) & (g90) & (!g319) & (g2259) & (g365)) + ((g87) & (sk[127]) & (g90) & (g319) & (!g2259) & (g365)) + ((g87) & (sk[127]) & (g90) & (g319) & (g2259) & (g365)));
	assign g2286 = (((!g1668) & (!g2033) & (!g2034) & (!sk[0]) & (g2284) & (!g2285)) + ((!g1668) & (!g2033) & (!g2034) & (!sk[0]) & (g2284) & (g2285)) + ((!g1668) & (!g2033) & (!g2034) & (sk[0]) & (g2284) & (!g2285)) + ((!g1668) & (!g2033) & (!g2034) & (sk[0]) & (g2284) & (g2285)) + ((!g1668) & (!g2033) & (g2034) & (!sk[0]) & (!g2284) & (!g2285)) + ((!g1668) & (!g2033) & (g2034) & (!sk[0]) & (!g2284) & (g2285)) + ((!g1668) & (!g2033) & (g2034) & (!sk[0]) & (g2284) & (!g2285)) + ((!g1668) & (!g2033) & (g2034) & (!sk[0]) & (g2284) & (g2285)) + ((!g1668) & (g2033) & (!g2034) & (!sk[0]) & (!g2284) & (!g2285)) + ((!g1668) & (g2033) & (!g2034) & (!sk[0]) & (!g2284) & (g2285)) + ((!g1668) & (g2033) & (!g2034) & (!sk[0]) & (g2284) & (!g2285)) + ((!g1668) & (g2033) & (!g2034) & (!sk[0]) & (g2284) & (g2285)) + ((!g1668) & (g2033) & (!g2034) & (sk[0]) & (!g2284) & (g2285)) + ((!g1668) & (g2033) & (!g2034) & (sk[0]) & (g2284) & (g2285)) + ((!g1668) & (g2033) & (g2034) & (!sk[0]) & (!g2284) & (!g2285)) + ((!g1668) & (g2033) & (g2034) & (!sk[0]) & (!g2284) & (g2285)) + ((!g1668) & (g2033) & (g2034) & (!sk[0]) & (g2284) & (!g2285)) + ((!g1668) & (g2033) & (g2034) & (!sk[0]) & (g2284) & (g2285)) + ((g1668) & (!g2033) & (!g2034) & (!sk[0]) & (g2284) & (!g2285)) + ((g1668) & (!g2033) & (!g2034) & (!sk[0]) & (g2284) & (g2285)) + ((g1668) & (!g2033) & (!g2034) & (sk[0]) & (g2284) & (!g2285)) + ((g1668) & (!g2033) & (!g2034) & (sk[0]) & (g2284) & (g2285)) + ((g1668) & (!g2033) & (g2034) & (!sk[0]) & (!g2284) & (!g2285)) + ((g1668) & (!g2033) & (g2034) & (!sk[0]) & (!g2284) & (g2285)) + ((g1668) & (!g2033) & (g2034) & (!sk[0]) & (g2284) & (!g2285)) + ((g1668) & (!g2033) & (g2034) & (!sk[0]) & (g2284) & (g2285)) + ((g1668) & (!g2033) & (g2034) & (sk[0]) & (!g2284) & (!g2285)) + ((g1668) & (!g2033) & (g2034) & (sk[0]) & (!g2284) & (g2285)) + ((g1668) & (!g2033) & (g2034) & (sk[0]) & (g2284) & (!g2285)) + ((g1668) & (!g2033) & (g2034) & (sk[0]) & (g2284) & (g2285)) + ((g1668) & (g2033) & (!g2034) & (!sk[0]) & (!g2284) & (!g2285)) + ((g1668) & (g2033) & (!g2034) & (!sk[0]) & (!g2284) & (g2285)) + ((g1668) & (g2033) & (!g2034) & (!sk[0]) & (g2284) & (!g2285)) + ((g1668) & (g2033) & (!g2034) & (!sk[0]) & (g2284) & (g2285)) + ((g1668) & (g2033) & (!g2034) & (sk[0]) & (!g2284) & (g2285)) + ((g1668) & (g2033) & (!g2034) & (sk[0]) & (g2284) & (g2285)) + ((g1668) & (g2033) & (g2034) & (!sk[0]) & (!g2284) & (!g2285)) + ((g1668) & (g2033) & (g2034) & (!sk[0]) & (!g2284) & (g2285)) + ((g1668) & (g2033) & (g2034) & (!sk[0]) & (g2284) & (!g2285)) + ((g1668) & (g2033) & (g2034) & (!sk[0]) & (g2284) & (g2285)));
	assign g2287 = (((!g2022) & (!nmi_i) & (!g2023) & (!g2029) & (!g2283) & (g2286)) + ((!g2022) & (!nmi_i) & (!g2023) & (!g2029) & (g2283) & (g2286)) + ((!g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2283) & (!g2286)) + ((!g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2283) & (g2286)) + ((!g2022) & (!nmi_i) & (g2023) & (!g2029) & (!g2283) & (g2286)) + ((!g2022) & (!nmi_i) & (g2023) & (!g2029) & (g2283) & (g2286)) + ((!g2022) & (!nmi_i) & (g2023) & (g2029) & (g2283) & (!g2286)) + ((!g2022) & (!nmi_i) & (g2023) & (g2029) & (g2283) & (g2286)) + ((!g2022) & (nmi_i) & (!g2023) & (!g2029) & (!g2283) & (g2286)) + ((!g2022) & (nmi_i) & (!g2023) & (!g2029) & (g2283) & (g2286)) + ((!g2022) & (nmi_i) & (!g2023) & (g2029) & (g2283) & (!g2286)) + ((!g2022) & (nmi_i) & (!g2023) & (g2029) & (g2283) & (g2286)) + ((!g2022) & (nmi_i) & (g2023) & (!g2029) & (!g2283) & (g2286)) + ((!g2022) & (nmi_i) & (g2023) & (!g2029) & (g2283) & (g2286)) + ((!g2022) & (nmi_i) & (g2023) & (g2029) & (g2283) & (!g2286)) + ((!g2022) & (nmi_i) & (g2023) & (g2029) & (g2283) & (g2286)) + ((g2022) & (!nmi_i) & (!g2023) & (!g2029) & (!g2283) & (g2286)) + ((g2022) & (!nmi_i) & (!g2023) & (!g2029) & (g2283) & (g2286)) + ((g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2283) & (!g2286)) + ((g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2283) & (g2286)));
	assign g2288 = (((!g123) & (!intr_i) & (!g2039) & (!g2056) & (!g2057) & (g2287)) + ((!g123) & (!intr_i) & (!g2039) & (!g2056) & (g2057) & (g2287)) + ((!g123) & (!intr_i) & (!g2039) & (g2056) & (!g2057) & (g2287)) + ((!g123) & (!intr_i) & (!g2039) & (g2056) & (g2057) & (g2287)) + ((!g123) & (!intr_i) & (g2039) & (!g2056) & (!g2057) & (g2287)) + ((!g123) & (!intr_i) & (g2039) & (!g2056) & (g2057) & (g2287)) + ((!g123) & (!intr_i) & (g2039) & (g2056) & (!g2057) & (g2287)) + ((!g123) & (!intr_i) & (g2039) & (g2056) & (g2057) & (g2287)) + ((!g123) & (intr_i) & (!g2039) & (!g2056) & (!g2057) & (g2287)) + ((!g123) & (intr_i) & (!g2039) & (!g2056) & (g2057) & (g2287)) + ((!g123) & (intr_i) & (!g2039) & (g2056) & (!g2057) & (g2287)) + ((!g123) & (intr_i) & (g2039) & (!g2056) & (!g2057) & (g2287)) + ((!g123) & (intr_i) & (g2039) & (g2056) & (!g2057) & (g2287)));
	assign g2290 = (((!g2073) & (!g2113) & (!g2114) & (!sk[3]) & (g2265) & (!g2289)) + ((!g2073) & (!g2113) & (!g2114) & (!sk[3]) & (g2265) & (g2289)) + ((!g2073) & (!g2113) & (!g2114) & (sk[3]) & (!g2265) & (g2289)) + ((!g2073) & (!g2113) & (!g2114) & (sk[3]) & (g2265) & (g2289)) + ((!g2073) & (!g2113) & (g2114) & (!sk[3]) & (!g2265) & (!g2289)) + ((!g2073) & (!g2113) & (g2114) & (!sk[3]) & (!g2265) & (g2289)) + ((!g2073) & (!g2113) & (g2114) & (!sk[3]) & (g2265) & (!g2289)) + ((!g2073) & (!g2113) & (g2114) & (!sk[3]) & (g2265) & (g2289)) + ((!g2073) & (!g2113) & (g2114) & (sk[3]) & (!g2265) & (!g2289)) + ((!g2073) & (!g2113) & (g2114) & (sk[3]) & (g2265) & (!g2289)) + ((!g2073) & (g2113) & (!g2114) & (!sk[3]) & (!g2265) & (!g2289)) + ((!g2073) & (g2113) & (!g2114) & (!sk[3]) & (!g2265) & (g2289)) + ((!g2073) & (g2113) & (!g2114) & (!sk[3]) & (g2265) & (!g2289)) + ((!g2073) & (g2113) & (!g2114) & (!sk[3]) & (g2265) & (g2289)) + ((!g2073) & (g2113) & (!g2114) & (sk[3]) & (!g2265) & (g2289)) + ((!g2073) & (g2113) & (!g2114) & (sk[3]) & (g2265) & (!g2289)) + ((!g2073) & (g2113) & (g2114) & (!sk[3]) & (!g2265) & (!g2289)) + ((!g2073) & (g2113) & (g2114) & (!sk[3]) & (!g2265) & (g2289)) + ((!g2073) & (g2113) & (g2114) & (!sk[3]) & (g2265) & (!g2289)) + ((!g2073) & (g2113) & (g2114) & (!sk[3]) & (g2265) & (g2289)) + ((!g2073) & (g2113) & (g2114) & (sk[3]) & (!g2265) & (!g2289)) + ((!g2073) & (g2113) & (g2114) & (sk[3]) & (g2265) & (g2289)) + ((g2073) & (!g2113) & (!g2114) & (!sk[3]) & (g2265) & (!g2289)) + ((g2073) & (!g2113) & (!g2114) & (!sk[3]) & (g2265) & (g2289)) + ((g2073) & (!g2113) & (!g2114) & (sk[3]) & (!g2265) & (g2289)) + ((g2073) & (!g2113) & (!g2114) & (sk[3]) & (g2265) & (!g2289)) + ((g2073) & (!g2113) & (g2114) & (!sk[3]) & (!g2265) & (!g2289)) + ((g2073) & (!g2113) & (g2114) & (!sk[3]) & (!g2265) & (g2289)) + ((g2073) & (!g2113) & (g2114) & (!sk[3]) & (g2265) & (!g2289)) + ((g2073) & (!g2113) & (g2114) & (!sk[3]) & (g2265) & (g2289)) + ((g2073) & (!g2113) & (g2114) & (sk[3]) & (!g2265) & (!g2289)) + ((g2073) & (!g2113) & (g2114) & (sk[3]) & (g2265) & (g2289)) + ((g2073) & (g2113) & (!g2114) & (!sk[3]) & (!g2265) & (!g2289)) + ((g2073) & (g2113) & (!g2114) & (!sk[3]) & (!g2265) & (g2289)) + ((g2073) & (g2113) & (!g2114) & (!sk[3]) & (g2265) & (!g2289)) + ((g2073) & (g2113) & (!g2114) & (!sk[3]) & (g2265) & (g2289)) + ((g2073) & (g2113) & (!g2114) & (sk[3]) & (!g2265) & (!g2289)) + ((g2073) & (g2113) & (!g2114) & (sk[3]) & (g2265) & (!g2289)) + ((g2073) & (g2113) & (g2114) & (!sk[3]) & (!g2265) & (!g2289)) + ((g2073) & (g2113) & (g2114) & (!sk[3]) & (!g2265) & (g2289)) + ((g2073) & (g2113) & (g2114) & (!sk[3]) & (g2265) & (!g2289)) + ((g2073) & (g2113) & (g2114) & (!sk[3]) & (g2265) & (g2289)) + ((g2073) & (g2113) & (g2114) & (sk[3]) & (!g2265) & (g2289)) + ((g2073) & (g2113) & (g2114) & (sk[3]) & (g2265) & (g2289)));
	assign g2291 = (((!sk[4]) & (!g2268) & (!g2269) & (g2270)) + ((!sk[4]) & (!g2268) & (g2269) & (!g2270)) + ((!sk[4]) & (!g2268) & (g2269) & (g2270)) + ((!sk[4]) & (g2268) & (!g2269) & (g2270)) + ((!sk[4]) & (g2268) & (g2269) & (!g2270)) + ((!sk[4]) & (g2268) & (g2269) & (g2270)) + ((sk[4]) & (!g2268) & (g2269) & (g2270)) + ((sk[4]) & (g2268) & (!g2269) & (g2270)) + ((sk[4]) & (g2268) & (g2269) & (!g2270)) + ((sk[4]) & (g2268) & (g2269) & (g2270)));
	assign g2292 = (((!g2073) & (sk[5]) & (g2113)) + ((g2073) & (!sk[5]) & (!g2113)) + ((g2073) & (!sk[5]) & (g2113)));
	assign g2293 = (((!g2289) & (sk[6]) & (!g2114)) + ((g2289) & (!sk[6]) & (!g2114)) + ((g2289) & (!sk[6]) & (g2114)) + ((g2289) & (sk[6]) & (g2114)));
	assign g2294 = (((!g2291) & (!g2292) & (!sk[7]) & (g2293)) + ((!g2291) & (!g2292) & (sk[7]) & (g2293)) + ((!g2291) & (g2292) & (!sk[7]) & (!g2293)) + ((!g2291) & (g2292) & (!sk[7]) & (g2293)) + ((!g2291) & (g2292) & (sk[7]) & (!g2293)) + ((g2291) & (!g2292) & (!sk[7]) & (g2293)) + ((g2291) & (!g2292) & (sk[7]) & (!g2293)) + ((g2291) & (g2292) & (!sk[7]) & (!g2293)) + ((g2291) & (g2292) & (!sk[7]) & (g2293)) + ((g2291) & (g2292) & (sk[7]) & (g2293)));
	assign g2295 = (((!sk[8]) & (g2114) & (!g2289)) + ((!sk[8]) & (g2114) & (g2289)) + ((sk[8]) & (g2114) & (g2289)));
	assign g2296 = (((!g2114) & (!g2113) & (!g2106) & (g2105) & (g2071) & (g2074)) + ((!g2114) & (!g2113) & (g2106) & (!g2105) & (!g2071) & (g2074)) + ((!g2114) & (!g2113) & (g2106) & (g2105) & (!g2071) & (g2074)) + ((!g2114) & (!g2113) & (g2106) & (g2105) & (g2071) & (g2074)) + ((!g2114) & (g2113) & (!g2106) & (!g2105) & (g2071) & (!g2074)) + ((!g2114) & (g2113) & (!g2106) & (g2105) & (g2071) & (!g2074)) + ((!g2114) & (g2113) & (!g2106) & (g2105) & (g2071) & (g2074)) + ((!g2114) & (g2113) & (g2106) & (!g2105) & (!g2071) & (g2074)) + ((!g2114) & (g2113) & (g2106) & (!g2105) & (g2071) & (!g2074)) + ((!g2114) & (g2113) & (g2106) & (g2105) & (!g2071) & (g2074)) + ((!g2114) & (g2113) & (g2106) & (g2105) & (g2071) & (!g2074)) + ((!g2114) & (g2113) & (g2106) & (g2105) & (g2071) & (g2074)) + ((g2114) & (!g2113) & (!g2106) & (!g2105) & (!g2071) & (!g2074)) + ((g2114) & (!g2113) & (!g2106) & (g2105) & (!g2071) & (!g2074)) + ((g2114) & (!g2113) & (!g2106) & (g2105) & (g2071) & (g2074)) + ((g2114) & (!g2113) & (g2106) & (!g2105) & (!g2071) & (!g2074)) + ((g2114) & (!g2113) & (g2106) & (!g2105) & (!g2071) & (g2074)) + ((g2114) & (!g2113) & (g2106) & (g2105) & (!g2071) & (!g2074)) + ((g2114) & (!g2113) & (g2106) & (g2105) & (!g2071) & (g2074)) + ((g2114) & (!g2113) & (g2106) & (g2105) & (g2071) & (g2074)) + ((g2114) & (g2113) & (!g2106) & (!g2105) & (!g2071) & (!g2074)) + ((g2114) & (g2113) & (!g2106) & (!g2105) & (g2071) & (!g2074)) + ((g2114) & (g2113) & (!g2106) & (g2105) & (!g2071) & (!g2074)) + ((g2114) & (g2113) & (!g2106) & (g2105) & (g2071) & (!g2074)) + ((g2114) & (g2113) & (!g2106) & (g2105) & (g2071) & (g2074)) + ((g2114) & (g2113) & (g2106) & (!g2105) & (!g2071) & (!g2074)) + ((g2114) & (g2113) & (g2106) & (!g2105) & (!g2071) & (g2074)) + ((g2114) & (g2113) & (g2106) & (!g2105) & (g2071) & (!g2074)) + ((g2114) & (g2113) & (g2106) & (g2105) & (!g2071) & (!g2074)) + ((g2114) & (g2113) & (g2106) & (g2105) & (!g2071) & (g2074)) + ((g2114) & (g2113) & (g2106) & (g2105) & (g2071) & (!g2074)) + ((g2114) & (g2113) & (g2106) & (g2105) & (g2071) & (g2074)));
	assign g2297 = (((!g2076) & (!sk[10]) & (!g2077) & (!g2183) & (g2296)) + ((!g2076) & (!sk[10]) & (!g2077) & (g2183) & (!g2296)) + ((!g2076) & (!sk[10]) & (!g2077) & (g2183) & (g2296)) + ((!g2076) & (!sk[10]) & (g2077) & (!g2183) & (!g2296)) + ((!g2076) & (!sk[10]) & (g2077) & (!g2183) & (g2296)) + ((!g2076) & (!sk[10]) & (g2077) & (g2183) & (!g2296)) + ((!g2076) & (!sk[10]) & (g2077) & (g2183) & (g2296)) + ((!g2076) & (sk[10]) & (!g2077) & (!g2183) & (g2296)) + ((!g2076) & (sk[10]) & (!g2077) & (g2183) & (g2296)) + ((!g2076) & (sk[10]) & (g2077) & (g2183) & (!g2296)) + ((!g2076) & (sk[10]) & (g2077) & (g2183) & (g2296)) + ((g2076) & (!sk[10]) & (!g2077) & (!g2183) & (g2296)) + ((g2076) & (!sk[10]) & (!g2077) & (g2183) & (!g2296)) + ((g2076) & (!sk[10]) & (!g2077) & (g2183) & (g2296)) + ((g2076) & (!sk[10]) & (g2077) & (!g2183) & (!g2296)) + ((g2076) & (!sk[10]) & (g2077) & (!g2183) & (g2296)) + ((g2076) & (!sk[10]) & (g2077) & (g2183) & (!g2296)) + ((g2076) & (!sk[10]) & (g2077) & (g2183) & (g2296)));
	assign g2298 = (((!g2195) & (!g2200) & (!g2199) & (g2187) & (g2076) & (g2077)) + ((!g2195) & (!g2200) & (g2199) & (!g2187) & (!g2076) & (g2077)) + ((!g2195) & (!g2200) & (g2199) & (g2187) & (!g2076) & (g2077)) + ((!g2195) & (!g2200) & (g2199) & (g2187) & (g2076) & (g2077)) + ((!g2195) & (g2200) & (!g2199) & (!g2187) & (g2076) & (!g2077)) + ((!g2195) & (g2200) & (!g2199) & (g2187) & (g2076) & (!g2077)) + ((!g2195) & (g2200) & (!g2199) & (g2187) & (g2076) & (g2077)) + ((!g2195) & (g2200) & (g2199) & (!g2187) & (!g2076) & (g2077)) + ((!g2195) & (g2200) & (g2199) & (!g2187) & (g2076) & (!g2077)) + ((!g2195) & (g2200) & (g2199) & (g2187) & (!g2076) & (g2077)) + ((!g2195) & (g2200) & (g2199) & (g2187) & (g2076) & (!g2077)) + ((!g2195) & (g2200) & (g2199) & (g2187) & (g2076) & (g2077)) + ((g2195) & (!g2200) & (!g2199) & (!g2187) & (!g2076) & (!g2077)) + ((g2195) & (!g2200) & (!g2199) & (g2187) & (!g2076) & (!g2077)) + ((g2195) & (!g2200) & (!g2199) & (g2187) & (g2076) & (g2077)) + ((g2195) & (!g2200) & (g2199) & (!g2187) & (!g2076) & (!g2077)) + ((g2195) & (!g2200) & (g2199) & (!g2187) & (!g2076) & (g2077)) + ((g2195) & (!g2200) & (g2199) & (g2187) & (!g2076) & (!g2077)) + ((g2195) & (!g2200) & (g2199) & (g2187) & (!g2076) & (g2077)) + ((g2195) & (!g2200) & (g2199) & (g2187) & (g2076) & (g2077)) + ((g2195) & (g2200) & (!g2199) & (!g2187) & (!g2076) & (!g2077)) + ((g2195) & (g2200) & (!g2199) & (!g2187) & (g2076) & (!g2077)) + ((g2195) & (g2200) & (!g2199) & (g2187) & (!g2076) & (!g2077)) + ((g2195) & (g2200) & (!g2199) & (g2187) & (g2076) & (!g2077)) + ((g2195) & (g2200) & (!g2199) & (g2187) & (g2076) & (g2077)) + ((g2195) & (g2200) & (g2199) & (!g2187) & (!g2076) & (!g2077)) + ((g2195) & (g2200) & (g2199) & (!g2187) & (!g2076) & (g2077)) + ((g2195) & (g2200) & (g2199) & (!g2187) & (g2076) & (!g2077)) + ((g2195) & (g2200) & (g2199) & (g2187) & (!g2076) & (!g2077)) + ((g2195) & (g2200) & (g2199) & (g2187) & (!g2076) & (g2077)) + ((g2195) & (g2200) & (g2199) & (g2187) & (g2076) & (!g2077)) + ((g2195) & (g2200) & (g2199) & (g2187) & (g2076) & (g2077)));
	assign g2299 = (((!g2189) & (!g2193) & (!g2188) & (g2192) & (g2076) & (g2077)) + ((!g2189) & (!g2193) & (g2188) & (!g2192) & (!g2076) & (g2077)) + ((!g2189) & (!g2193) & (g2188) & (g2192) & (!g2076) & (g2077)) + ((!g2189) & (!g2193) & (g2188) & (g2192) & (g2076) & (g2077)) + ((!g2189) & (g2193) & (!g2188) & (!g2192) & (g2076) & (!g2077)) + ((!g2189) & (g2193) & (!g2188) & (g2192) & (g2076) & (!g2077)) + ((!g2189) & (g2193) & (!g2188) & (g2192) & (g2076) & (g2077)) + ((!g2189) & (g2193) & (g2188) & (!g2192) & (!g2076) & (g2077)) + ((!g2189) & (g2193) & (g2188) & (!g2192) & (g2076) & (!g2077)) + ((!g2189) & (g2193) & (g2188) & (g2192) & (!g2076) & (g2077)) + ((!g2189) & (g2193) & (g2188) & (g2192) & (g2076) & (!g2077)) + ((!g2189) & (g2193) & (g2188) & (g2192) & (g2076) & (g2077)) + ((g2189) & (!g2193) & (!g2188) & (!g2192) & (!g2076) & (!g2077)) + ((g2189) & (!g2193) & (!g2188) & (g2192) & (!g2076) & (!g2077)) + ((g2189) & (!g2193) & (!g2188) & (g2192) & (g2076) & (g2077)) + ((g2189) & (!g2193) & (g2188) & (!g2192) & (!g2076) & (!g2077)) + ((g2189) & (!g2193) & (g2188) & (!g2192) & (!g2076) & (g2077)) + ((g2189) & (!g2193) & (g2188) & (g2192) & (!g2076) & (!g2077)) + ((g2189) & (!g2193) & (g2188) & (g2192) & (!g2076) & (g2077)) + ((g2189) & (!g2193) & (g2188) & (g2192) & (g2076) & (g2077)) + ((g2189) & (g2193) & (!g2188) & (!g2192) & (!g2076) & (!g2077)) + ((g2189) & (g2193) & (!g2188) & (!g2192) & (g2076) & (!g2077)) + ((g2189) & (g2193) & (!g2188) & (g2192) & (!g2076) & (!g2077)) + ((g2189) & (g2193) & (!g2188) & (g2192) & (g2076) & (!g2077)) + ((g2189) & (g2193) & (!g2188) & (g2192) & (g2076) & (g2077)) + ((g2189) & (g2193) & (g2188) & (!g2192) & (!g2076) & (!g2077)) + ((g2189) & (g2193) & (g2188) & (!g2192) & (!g2076) & (g2077)) + ((g2189) & (g2193) & (g2188) & (!g2192) & (g2076) & (!g2077)) + ((g2189) & (g2193) & (g2188) & (g2192) & (!g2076) & (!g2077)) + ((g2189) & (g2193) & (g2188) & (g2192) & (!g2076) & (g2077)) + ((g2189) & (g2193) & (g2188) & (g2192) & (g2076) & (!g2077)) + ((g2189) & (g2193) & (g2188) & (g2192) & (g2076) & (g2077)));
	assign g2300 = (((!g2073) & (!g2080) & (!g2125) & (g2297) & (!g2298) & (!g2299)) + ((!g2073) & (!g2080) & (!g2125) & (g2297) & (!g2298) & (g2299)) + ((!g2073) & (!g2080) & (!g2125) & (g2297) & (g2298) & (!g2299)) + ((!g2073) & (!g2080) & (!g2125) & (g2297) & (g2298) & (g2299)) + ((!g2073) & (!g2080) & (g2125) & (!g2297) & (g2298) & (!g2299)) + ((!g2073) & (!g2080) & (g2125) & (!g2297) & (g2298) & (g2299)) + ((!g2073) & (!g2080) & (g2125) & (g2297) & (g2298) & (!g2299)) + ((!g2073) & (!g2080) & (g2125) & (g2297) & (g2298) & (g2299)) + ((!g2073) & (g2080) & (!g2125) & (g2297) & (!g2298) & (!g2299)) + ((!g2073) & (g2080) & (!g2125) & (g2297) & (!g2298) & (g2299)) + ((!g2073) & (g2080) & (!g2125) & (g2297) & (g2298) & (!g2299)) + ((!g2073) & (g2080) & (!g2125) & (g2297) & (g2298) & (g2299)) + ((!g2073) & (g2080) & (g2125) & (!g2297) & (g2298) & (!g2299)) + ((!g2073) & (g2080) & (g2125) & (!g2297) & (g2298) & (g2299)) + ((!g2073) & (g2080) & (g2125) & (g2297) & (g2298) & (!g2299)) + ((!g2073) & (g2080) & (g2125) & (g2297) & (g2298) & (g2299)) + ((g2073) & (!g2080) & (g2125) & (!g2297) & (!g2298) & (g2299)) + ((g2073) & (!g2080) & (g2125) & (!g2297) & (g2298) & (g2299)) + ((g2073) & (!g2080) & (g2125) & (g2297) & (!g2298) & (g2299)) + ((g2073) & (!g2080) & (g2125) & (g2297) & (g2298) & (g2299)) + ((g2073) & (g2080) & (!g2125) & (g2297) & (!g2298) & (!g2299)) + ((g2073) & (g2080) & (!g2125) & (g2297) & (!g2298) & (g2299)) + ((g2073) & (g2080) & (!g2125) & (g2297) & (g2298) & (!g2299)) + ((g2073) & (g2080) & (!g2125) & (g2297) & (g2298) & (g2299)) + ((g2073) & (g2080) & (g2125) & (!g2297) & (!g2298) & (g2299)) + ((g2073) & (g2080) & (g2125) & (!g2297) & (g2298) & (g2299)) + ((g2073) & (g2080) & (g2125) & (g2297) & (!g2298) & (g2299)) + ((g2073) & (g2080) & (g2125) & (g2297) & (g2298) & (g2299)));
	assign g2301 = (((!g2114) & (!g2289) & (!g2124) & (!g2264) & (!g3725) & (!g2300)) + ((!g2114) & (!g2289) & (!g2124) & (!g2264) & (g3725) & (!g2300)) + ((!g2114) & (!g2289) & (!g2124) & (g2264) & (!g3725) & (!g2300)) + ((!g2114) & (!g2289) & (!g2124) & (g2264) & (!g3725) & (g2300)) + ((!g2114) & (!g2289) & (g2124) & (!g2264) & (!g3725) & (!g2300)) + ((!g2114) & (!g2289) & (g2124) & (!g2264) & (!g3725) & (g2300)) + ((!g2114) & (!g2289) & (g2124) & (!g2264) & (g3725) & (!g2300)) + ((!g2114) & (!g2289) & (g2124) & (!g2264) & (g3725) & (g2300)) + ((!g2114) & (!g2289) & (g2124) & (g2264) & (!g3725) & (!g2300)) + ((!g2114) & (!g2289) & (g2124) & (g2264) & (!g3725) & (g2300)) + ((!g2114) & (!g2289) & (g2124) & (g2264) & (g3725) & (!g2300)) + ((!g2114) & (!g2289) & (g2124) & (g2264) & (g3725) & (g2300)) + ((!g2114) & (g2289) & (!g2124) & (!g2264) & (!g3725) & (!g2300)) + ((!g2114) & (g2289) & (!g2124) & (!g2264) & (g3725) & (!g2300)) + ((!g2114) & (g2289) & (!g2124) & (g2264) & (!g3725) & (!g2300)) + ((!g2114) & (g2289) & (!g2124) & (g2264) & (!g3725) & (g2300)) + ((g2114) & (!g2289) & (!g2124) & (!g2264) & (!g3725) & (!g2300)) + ((g2114) & (!g2289) & (!g2124) & (!g2264) & (g3725) & (!g2300)) + ((g2114) & (!g2289) & (!g2124) & (g2264) & (!g3725) & (!g2300)) + ((g2114) & (!g2289) & (!g2124) & (g2264) & (!g3725) & (g2300)) + ((g2114) & (g2289) & (!g2124) & (!g2264) & (!g3725) & (!g2300)) + ((g2114) & (g2289) & (!g2124) & (!g2264) & (g3725) & (!g2300)) + ((g2114) & (g2289) & (!g2124) & (g2264) & (!g3725) & (!g2300)) + ((g2114) & (g2289) & (!g2124) & (g2264) & (!g3725) & (g2300)) + ((g2114) & (g2289) & (g2124) & (g2264) & (!g3725) & (!g2300)) + ((g2114) & (g2289) & (g2124) & (g2264) & (!g3725) & (g2300)) + ((g2114) & (g2289) & (g2124) & (g2264) & (g3725) & (!g2300)) + ((g2114) & (g2289) & (g2124) & (g2264) & (g3725) & (g2300)));
	assign g2302 = (((!dmem_dat_ix5x) & (!dmem_dat_ix13x) & (!dmem_dat_ix29x) & (dmem_dat_ix21x) & (g2206) & (g2207)) + ((!dmem_dat_ix5x) & (!dmem_dat_ix13x) & (dmem_dat_ix29x) & (!dmem_dat_ix21x) & (!g2206) & (g2207)) + ((!dmem_dat_ix5x) & (!dmem_dat_ix13x) & (dmem_dat_ix29x) & (dmem_dat_ix21x) & (!g2206) & (g2207)) + ((!dmem_dat_ix5x) & (!dmem_dat_ix13x) & (dmem_dat_ix29x) & (dmem_dat_ix21x) & (g2206) & (g2207)) + ((!dmem_dat_ix5x) & (dmem_dat_ix13x) & (!dmem_dat_ix29x) & (!dmem_dat_ix21x) & (g2206) & (!g2207)) + ((!dmem_dat_ix5x) & (dmem_dat_ix13x) & (!dmem_dat_ix29x) & (dmem_dat_ix21x) & (g2206) & (!g2207)) + ((!dmem_dat_ix5x) & (dmem_dat_ix13x) & (!dmem_dat_ix29x) & (dmem_dat_ix21x) & (g2206) & (g2207)) + ((!dmem_dat_ix5x) & (dmem_dat_ix13x) & (dmem_dat_ix29x) & (!dmem_dat_ix21x) & (!g2206) & (g2207)) + ((!dmem_dat_ix5x) & (dmem_dat_ix13x) & (dmem_dat_ix29x) & (!dmem_dat_ix21x) & (g2206) & (!g2207)) + ((!dmem_dat_ix5x) & (dmem_dat_ix13x) & (dmem_dat_ix29x) & (dmem_dat_ix21x) & (!g2206) & (g2207)) + ((!dmem_dat_ix5x) & (dmem_dat_ix13x) & (dmem_dat_ix29x) & (dmem_dat_ix21x) & (g2206) & (!g2207)) + ((!dmem_dat_ix5x) & (dmem_dat_ix13x) & (dmem_dat_ix29x) & (dmem_dat_ix21x) & (g2206) & (g2207)) + ((dmem_dat_ix5x) & (!dmem_dat_ix13x) & (!dmem_dat_ix29x) & (!dmem_dat_ix21x) & (!g2206) & (!g2207)) + ((dmem_dat_ix5x) & (!dmem_dat_ix13x) & (!dmem_dat_ix29x) & (dmem_dat_ix21x) & (!g2206) & (!g2207)) + ((dmem_dat_ix5x) & (!dmem_dat_ix13x) & (!dmem_dat_ix29x) & (dmem_dat_ix21x) & (g2206) & (g2207)) + ((dmem_dat_ix5x) & (!dmem_dat_ix13x) & (dmem_dat_ix29x) & (!dmem_dat_ix21x) & (!g2206) & (!g2207)) + ((dmem_dat_ix5x) & (!dmem_dat_ix13x) & (dmem_dat_ix29x) & (!dmem_dat_ix21x) & (!g2206) & (g2207)) + ((dmem_dat_ix5x) & (!dmem_dat_ix13x) & (dmem_dat_ix29x) & (dmem_dat_ix21x) & (!g2206) & (!g2207)) + ((dmem_dat_ix5x) & (!dmem_dat_ix13x) & (dmem_dat_ix29x) & (dmem_dat_ix21x) & (!g2206) & (g2207)) + ((dmem_dat_ix5x) & (!dmem_dat_ix13x) & (dmem_dat_ix29x) & (dmem_dat_ix21x) & (g2206) & (g2207)) + ((dmem_dat_ix5x) & (dmem_dat_ix13x) & (!dmem_dat_ix29x) & (!dmem_dat_ix21x) & (!g2206) & (!g2207)) + ((dmem_dat_ix5x) & (dmem_dat_ix13x) & (!dmem_dat_ix29x) & (!dmem_dat_ix21x) & (g2206) & (!g2207)) + ((dmem_dat_ix5x) & (dmem_dat_ix13x) & (!dmem_dat_ix29x) & (dmem_dat_ix21x) & (!g2206) & (!g2207)) + ((dmem_dat_ix5x) & (dmem_dat_ix13x) & (!dmem_dat_ix29x) & (dmem_dat_ix21x) & (g2206) & (!g2207)) + ((dmem_dat_ix5x) & (dmem_dat_ix13x) & (!dmem_dat_ix29x) & (dmem_dat_ix21x) & (g2206) & (g2207)) + ((dmem_dat_ix5x) & (dmem_dat_ix13x) & (dmem_dat_ix29x) & (!dmem_dat_ix21x) & (!g2206) & (!g2207)) + ((dmem_dat_ix5x) & (dmem_dat_ix13x) & (dmem_dat_ix29x) & (!dmem_dat_ix21x) & (!g2206) & (g2207)) + ((dmem_dat_ix5x) & (dmem_dat_ix13x) & (dmem_dat_ix29x) & (!dmem_dat_ix21x) & (g2206) & (!g2207)) + ((dmem_dat_ix5x) & (dmem_dat_ix13x) & (dmem_dat_ix29x) & (dmem_dat_ix21x) & (!g2206) & (!g2207)) + ((dmem_dat_ix5x) & (dmem_dat_ix13x) & (dmem_dat_ix29x) & (dmem_dat_ix21x) & (!g2206) & (g2207)) + ((dmem_dat_ix5x) & (dmem_dat_ix13x) & (dmem_dat_ix29x) & (dmem_dat_ix21x) & (g2206) & (!g2207)) + ((dmem_dat_ix5x) & (dmem_dat_ix13x) & (dmem_dat_ix29x) & (dmem_dat_ix21x) & (g2206) & (g2207)));
	assign g2303 = (((!g2128) & (!sk[16]) & (!g2129) & (!dmem_dat_ix5x) & (dmem_dat_ix21x)) + ((!g2128) & (!sk[16]) & (!g2129) & (dmem_dat_ix5x) & (!dmem_dat_ix21x)) + ((!g2128) & (!sk[16]) & (!g2129) & (dmem_dat_ix5x) & (dmem_dat_ix21x)) + ((!g2128) & (!sk[16]) & (g2129) & (!dmem_dat_ix5x) & (!dmem_dat_ix21x)) + ((!g2128) & (!sk[16]) & (g2129) & (!dmem_dat_ix5x) & (dmem_dat_ix21x)) + ((!g2128) & (!sk[16]) & (g2129) & (dmem_dat_ix5x) & (!dmem_dat_ix21x)) + ((!g2128) & (!sk[16]) & (g2129) & (dmem_dat_ix5x) & (dmem_dat_ix21x)) + ((!g2128) & (sk[16]) & (!g2129) & (!dmem_dat_ix5x) & (dmem_dat_ix21x)) + ((!g2128) & (sk[16]) & (!g2129) & (dmem_dat_ix5x) & (dmem_dat_ix21x)) + ((!g2128) & (sk[16]) & (g2129) & (dmem_dat_ix5x) & (!dmem_dat_ix21x)) + ((!g2128) & (sk[16]) & (g2129) & (dmem_dat_ix5x) & (dmem_dat_ix21x)) + ((g2128) & (!sk[16]) & (!g2129) & (!dmem_dat_ix5x) & (dmem_dat_ix21x)) + ((g2128) & (!sk[16]) & (!g2129) & (dmem_dat_ix5x) & (!dmem_dat_ix21x)) + ((g2128) & (!sk[16]) & (!g2129) & (dmem_dat_ix5x) & (dmem_dat_ix21x)) + ((g2128) & (!sk[16]) & (g2129) & (!dmem_dat_ix5x) & (!dmem_dat_ix21x)) + ((g2128) & (!sk[16]) & (g2129) & (!dmem_dat_ix5x) & (dmem_dat_ix21x)) + ((g2128) & (!sk[16]) & (g2129) & (dmem_dat_ix5x) & (!dmem_dat_ix21x)) + ((g2128) & (!sk[16]) & (g2129) & (dmem_dat_ix5x) & (dmem_dat_ix21x)));
	assign g2304 = (((!g2301) & (!g2114) & (!g2302) & (!g2303) & (!g2281) & (!g75)) + ((!g2301) & (!g2114) & (!g2302) & (g2303) & (!g2281) & (!g75)) + ((!g2301) & (!g2114) & (!g2302) & (g2303) & (g2281) & (g75)) + ((!g2301) & (!g2114) & (g2302) & (!g2303) & (!g2281) & (!g75)) + ((!g2301) & (!g2114) & (g2302) & (!g2303) & (!g2281) & (g75)) + ((!g2301) & (!g2114) & (g2302) & (g2303) & (!g2281) & (!g75)) + ((!g2301) & (!g2114) & (g2302) & (g2303) & (!g2281) & (g75)) + ((!g2301) & (!g2114) & (g2302) & (g2303) & (g2281) & (g75)) + ((!g2301) & (g2114) & (!g2302) & (!g2303) & (!g2281) & (!g75)) + ((!g2301) & (g2114) & (!g2302) & (!g2303) & (g2281) & (!g75)) + ((!g2301) & (g2114) & (!g2302) & (g2303) & (!g2281) & (!g75)) + ((!g2301) & (g2114) & (!g2302) & (g2303) & (g2281) & (!g75)) + ((!g2301) & (g2114) & (!g2302) & (g2303) & (g2281) & (g75)) + ((!g2301) & (g2114) & (g2302) & (!g2303) & (!g2281) & (!g75)) + ((!g2301) & (g2114) & (g2302) & (!g2303) & (!g2281) & (g75)) + ((!g2301) & (g2114) & (g2302) & (!g2303) & (g2281) & (!g75)) + ((!g2301) & (g2114) & (g2302) & (g2303) & (!g2281) & (!g75)) + ((!g2301) & (g2114) & (g2302) & (g2303) & (!g2281) & (g75)) + ((!g2301) & (g2114) & (g2302) & (g2303) & (g2281) & (!g75)) + ((!g2301) & (g2114) & (g2302) & (g2303) & (g2281) & (g75)) + ((g2301) & (!g2114) & (!g2302) & (g2303) & (g2281) & (g75)) + ((g2301) & (!g2114) & (g2302) & (!g2303) & (!g2281) & (g75)) + ((g2301) & (!g2114) & (g2302) & (g2303) & (!g2281) & (g75)) + ((g2301) & (!g2114) & (g2302) & (g2303) & (g2281) & (g75)) + ((g2301) & (g2114) & (!g2302) & (!g2303) & (g2281) & (!g75)) + ((g2301) & (g2114) & (!g2302) & (g2303) & (g2281) & (!g75)) + ((g2301) & (g2114) & (!g2302) & (g2303) & (g2281) & (g75)) + ((g2301) & (g2114) & (g2302) & (!g2303) & (!g2281) & (g75)) + ((g2301) & (g2114) & (g2302) & (!g2303) & (g2281) & (!g75)) + ((g2301) & (g2114) & (g2302) & (g2303) & (!g2281) & (g75)) + ((g2301) & (g2114) & (g2302) & (g2303) & (g2281) & (!g75)) + ((g2301) & (g2114) & (g2302) & (g2303) & (g2281) & (g75)));
	assign g2305 = (((!g141) & (!sk[18]) & (!g275) & (!g319) & (g365) & (!g408)) + ((!g141) & (!sk[18]) & (!g275) & (!g319) & (g365) & (g408)) + ((!g141) & (!sk[18]) & (!g275) & (g319) & (!g365) & (!g408)) + ((!g141) & (!sk[18]) & (!g275) & (g319) & (!g365) & (g408)) + ((!g141) & (!sk[18]) & (!g275) & (g319) & (g365) & (!g408)) + ((!g141) & (!sk[18]) & (!g275) & (g319) & (g365) & (g408)) + ((!g141) & (!sk[18]) & (g275) & (!g319) & (!g365) & (!g408)) + ((!g141) & (!sk[18]) & (g275) & (!g319) & (!g365) & (g408)) + ((!g141) & (!sk[18]) & (g275) & (!g319) & (g365) & (!g408)) + ((!g141) & (!sk[18]) & (g275) & (!g319) & (g365) & (g408)) + ((!g141) & (!sk[18]) & (g275) & (g319) & (!g365) & (!g408)) + ((!g141) & (!sk[18]) & (g275) & (g319) & (!g365) & (g408)) + ((!g141) & (!sk[18]) & (g275) & (g319) & (g365) & (!g408)) + ((!g141) & (!sk[18]) & (g275) & (g319) & (g365) & (g408)) + ((!g141) & (sk[18]) & (!g275) & (!g319) & (!g365) & (g408)) + ((!g141) & (sk[18]) & (!g275) & (!g319) & (g365) & (g408)) + ((!g141) & (sk[18]) & (!g275) & (g319) & (!g365) & (g408)) + ((!g141) & (sk[18]) & (!g275) & (g319) & (g365) & (g408)) + ((!g141) & (sk[18]) & (g275) & (!g319) & (!g365) & (g408)) + ((!g141) & (sk[18]) & (g275) & (!g319) & (g365) & (g408)) + ((!g141) & (sk[18]) & (g275) & (g319) & (!g365) & (g408)) + ((!g141) & (sk[18]) & (g275) & (g319) & (g365) & (g408)) + ((g141) & (!sk[18]) & (!g275) & (!g319) & (g365) & (!g408)) + ((g141) & (!sk[18]) & (!g275) & (!g319) & (g365) & (g408)) + ((g141) & (!sk[18]) & (!g275) & (g319) & (!g365) & (!g408)) + ((g141) & (!sk[18]) & (!g275) & (g319) & (!g365) & (g408)) + ((g141) & (!sk[18]) & (!g275) & (g319) & (g365) & (!g408)) + ((g141) & (!sk[18]) & (!g275) & (g319) & (g365) & (g408)) + ((g141) & (!sk[18]) & (g275) & (!g319) & (!g365) & (!g408)) + ((g141) & (!sk[18]) & (g275) & (!g319) & (!g365) & (g408)) + ((g141) & (!sk[18]) & (g275) & (!g319) & (g365) & (!g408)) + ((g141) & (!sk[18]) & (g275) & (!g319) & (g365) & (g408)) + ((g141) & (!sk[18]) & (g275) & (g319) & (!g365) & (!g408)) + ((g141) & (!sk[18]) & (g275) & (g319) & (!g365) & (g408)) + ((g141) & (!sk[18]) & (g275) & (g319) & (g365) & (!g408)) + ((g141) & (!sk[18]) & (g275) & (g319) & (g365) & (g408)) + ((g141) & (sk[18]) & (!g275) & (!g319) & (!g365) & (g408)) + ((g141) & (sk[18]) & (!g275) & (!g319) & (g365) & (g408)) + ((g141) & (sk[18]) & (!g275) & (g319) & (!g365) & (g408)) + ((g141) & (sk[18]) & (!g275) & (g319) & (g365) & (g408)) + ((g141) & (sk[18]) & (g275) & (!g319) & (!g365) & (g408)) + ((g141) & (sk[18]) & (g275) & (!g319) & (g365) & (g408)) + ((g141) & (sk[18]) & (g275) & (g319) & (!g365) & (g408)) + ((g141) & (sk[18]) & (g275) & (g319) & (g365) & (!g408)));
	assign g5030 = (((!g2921) & (!sk[19]) & (!g3060) & (g2306)) + ((!g2921) & (!sk[19]) & (g3060) & (!g2306)) + ((!g2921) & (!sk[19]) & (g3060) & (g2306)) + ((!g2921) & (sk[19]) & (!g3060) & (g2306)) + ((!g2921) & (sk[19]) & (g3060) & (g2306)) + ((g2921) & (!sk[19]) & (!g3060) & (g2306)) + ((g2921) & (!sk[19]) & (g3060) & (!g2306)) + ((g2921) & (!sk[19]) & (g3060) & (g2306)) + ((g2921) & (sk[19]) & (g3060) & (!g2306)) + ((g2921) & (sk[19]) & (g3060) & (g2306)));
	assign g2307 = (((!sk[20]) & (!g87) & (!g90) & (!g319) & (g2259) & (!g365)) + ((!sk[20]) & (!g87) & (!g90) & (!g319) & (g2259) & (g365)) + ((!sk[20]) & (!g87) & (!g90) & (g319) & (!g2259) & (!g365)) + ((!sk[20]) & (!g87) & (!g90) & (g319) & (!g2259) & (g365)) + ((!sk[20]) & (!g87) & (!g90) & (g319) & (g2259) & (!g365)) + ((!sk[20]) & (!g87) & (!g90) & (g319) & (g2259) & (g365)) + ((!sk[20]) & (!g87) & (g90) & (!g319) & (!g2259) & (!g365)) + ((!sk[20]) & (!g87) & (g90) & (!g319) & (!g2259) & (g365)) + ((!sk[20]) & (!g87) & (g90) & (!g319) & (g2259) & (!g365)) + ((!sk[20]) & (!g87) & (g90) & (!g319) & (g2259) & (g365)) + ((!sk[20]) & (!g87) & (g90) & (g319) & (!g2259) & (!g365)) + ((!sk[20]) & (!g87) & (g90) & (g319) & (!g2259) & (g365)) + ((!sk[20]) & (!g87) & (g90) & (g319) & (g2259) & (!g365)) + ((!sk[20]) & (!g87) & (g90) & (g319) & (g2259) & (g365)) + ((!sk[20]) & (g87) & (!g90) & (!g319) & (g2259) & (!g365)) + ((!sk[20]) & (g87) & (!g90) & (!g319) & (g2259) & (g365)) + ((!sk[20]) & (g87) & (!g90) & (g319) & (!g2259) & (!g365)) + ((!sk[20]) & (g87) & (!g90) & (g319) & (!g2259) & (g365)) + ((!sk[20]) & (g87) & (!g90) & (g319) & (g2259) & (!g365)) + ((!sk[20]) & (g87) & (!g90) & (g319) & (g2259) & (g365)) + ((!sk[20]) & (g87) & (g90) & (!g319) & (!g2259) & (!g365)) + ((!sk[20]) & (g87) & (g90) & (!g319) & (!g2259) & (g365)) + ((!sk[20]) & (g87) & (g90) & (!g319) & (g2259) & (!g365)) + ((!sk[20]) & (g87) & (g90) & (!g319) & (g2259) & (g365)) + ((!sk[20]) & (g87) & (g90) & (g319) & (!g2259) & (!g365)) + ((!sk[20]) & (g87) & (g90) & (g319) & (!g2259) & (g365)) + ((!sk[20]) & (g87) & (g90) & (g319) & (g2259) & (!g365)) + ((!sk[20]) & (g87) & (g90) & (g319) & (g2259) & (g365)) + ((sk[20]) & (!g87) & (!g90) & (g319) & (g2259) & (g365)) + ((sk[20]) & (!g87) & (g90) & (!g319) & (!g2259) & (g365)) + ((sk[20]) & (!g87) & (g90) & (!g319) & (g2259) & (g365)) + ((sk[20]) & (!g87) & (g90) & (g319) & (!g2259) & (g365)) + ((sk[20]) & (!g87) & (g90) & (g319) & (g2259) & (!g365)) + ((sk[20]) & (!g87) & (g90) & (g319) & (g2259) & (g365)) + ((sk[20]) & (g87) & (!g90) & (!g319) & (g2259) & (g365)) + ((sk[20]) & (g87) & (!g90) & (g319) & (!g2259) & (g365)) + ((sk[20]) & (g87) & (!g90) & (g319) & (g2259) & (g365)) + ((sk[20]) & (g87) & (g90) & (!g319) & (!g2259) & (g365)) + ((sk[20]) & (g87) & (g90) & (!g319) & (g2259) & (!g365)) + ((sk[20]) & (g87) & (g90) & (!g319) & (g2259) & (g365)) + ((sk[20]) & (g87) & (g90) & (g319) & (!g2259) & (!g365)) + ((sk[20]) & (g87) & (g90) & (g319) & (!g2259) & (g365)) + ((sk[20]) & (g87) & (g90) & (g319) & (g2259) & (!g365)) + ((sk[20]) & (g87) & (g90) & (g319) & (g2259) & (g365)));
	assign g2308 = (((!g318) & (!sk[21]) & (!g408) & (g2307)) + ((!g318) & (!sk[21]) & (g408) & (!g2307)) + ((!g318) & (!sk[21]) & (g408) & (g2307)) + ((!g318) & (sk[21]) & (!g408) & (g2307)) + ((!g318) & (sk[21]) & (g408) & (!g2307)) + ((g318) & (!sk[21]) & (!g408) & (g2307)) + ((g318) & (!sk[21]) & (g408) & (!g2307)) + ((g318) & (!sk[21]) & (g408) & (g2307)) + ((g318) & (sk[21]) & (!g408) & (!g2307)) + ((g318) & (sk[21]) & (g408) & (g2307)));
	assign g2309 = (((!g1680) & (!g2033) & (!sk[22]) & (!g2034) & (g2306) & (!g2308)) + ((!g1680) & (!g2033) & (!sk[22]) & (!g2034) & (g2306) & (g2308)) + ((!g1680) & (!g2033) & (!sk[22]) & (g2034) & (!g2306) & (!g2308)) + ((!g1680) & (!g2033) & (!sk[22]) & (g2034) & (!g2306) & (g2308)) + ((!g1680) & (!g2033) & (!sk[22]) & (g2034) & (g2306) & (!g2308)) + ((!g1680) & (!g2033) & (!sk[22]) & (g2034) & (g2306) & (g2308)) + ((!g1680) & (!g2033) & (sk[22]) & (!g2034) & (g2306) & (!g2308)) + ((!g1680) & (!g2033) & (sk[22]) & (!g2034) & (g2306) & (g2308)) + ((!g1680) & (g2033) & (!sk[22]) & (!g2034) & (!g2306) & (!g2308)) + ((!g1680) & (g2033) & (!sk[22]) & (!g2034) & (!g2306) & (g2308)) + ((!g1680) & (g2033) & (!sk[22]) & (!g2034) & (g2306) & (!g2308)) + ((!g1680) & (g2033) & (!sk[22]) & (!g2034) & (g2306) & (g2308)) + ((!g1680) & (g2033) & (!sk[22]) & (g2034) & (!g2306) & (!g2308)) + ((!g1680) & (g2033) & (!sk[22]) & (g2034) & (!g2306) & (g2308)) + ((!g1680) & (g2033) & (!sk[22]) & (g2034) & (g2306) & (!g2308)) + ((!g1680) & (g2033) & (!sk[22]) & (g2034) & (g2306) & (g2308)) + ((!g1680) & (g2033) & (sk[22]) & (!g2034) & (!g2306) & (g2308)) + ((!g1680) & (g2033) & (sk[22]) & (!g2034) & (g2306) & (g2308)) + ((g1680) & (!g2033) & (!sk[22]) & (!g2034) & (g2306) & (!g2308)) + ((g1680) & (!g2033) & (!sk[22]) & (!g2034) & (g2306) & (g2308)) + ((g1680) & (!g2033) & (!sk[22]) & (g2034) & (!g2306) & (!g2308)) + ((g1680) & (!g2033) & (!sk[22]) & (g2034) & (!g2306) & (g2308)) + ((g1680) & (!g2033) & (!sk[22]) & (g2034) & (g2306) & (!g2308)) + ((g1680) & (!g2033) & (!sk[22]) & (g2034) & (g2306) & (g2308)) + ((g1680) & (!g2033) & (sk[22]) & (!g2034) & (g2306) & (!g2308)) + ((g1680) & (!g2033) & (sk[22]) & (!g2034) & (g2306) & (g2308)) + ((g1680) & (!g2033) & (sk[22]) & (g2034) & (!g2306) & (!g2308)) + ((g1680) & (!g2033) & (sk[22]) & (g2034) & (!g2306) & (g2308)) + ((g1680) & (!g2033) & (sk[22]) & (g2034) & (g2306) & (!g2308)) + ((g1680) & (!g2033) & (sk[22]) & (g2034) & (g2306) & (g2308)) + ((g1680) & (g2033) & (!sk[22]) & (!g2034) & (!g2306) & (!g2308)) + ((g1680) & (g2033) & (!sk[22]) & (!g2034) & (!g2306) & (g2308)) + ((g1680) & (g2033) & (!sk[22]) & (!g2034) & (g2306) & (!g2308)) + ((g1680) & (g2033) & (!sk[22]) & (!g2034) & (g2306) & (g2308)) + ((g1680) & (g2033) & (!sk[22]) & (g2034) & (!g2306) & (!g2308)) + ((g1680) & (g2033) & (!sk[22]) & (g2034) & (!g2306) & (g2308)) + ((g1680) & (g2033) & (!sk[22]) & (g2034) & (g2306) & (!g2308)) + ((g1680) & (g2033) & (!sk[22]) & (g2034) & (g2306) & (g2308)) + ((g1680) & (g2033) & (sk[22]) & (!g2034) & (!g2306) & (g2308)) + ((g1680) & (g2033) & (sk[22]) & (!g2034) & (g2306) & (g2308)));
	assign g2310 = (((!g2022) & (!nmi_i) & (!g2023) & (!g2029) & (!g2305) & (g2309)) + ((!g2022) & (!nmi_i) & (!g2023) & (!g2029) & (g2305) & (g2309)) + ((!g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2305) & (!g2309)) + ((!g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2305) & (g2309)) + ((!g2022) & (!nmi_i) & (g2023) & (!g2029) & (!g2305) & (g2309)) + ((!g2022) & (!nmi_i) & (g2023) & (!g2029) & (g2305) & (g2309)) + ((!g2022) & (!nmi_i) & (g2023) & (g2029) & (g2305) & (!g2309)) + ((!g2022) & (!nmi_i) & (g2023) & (g2029) & (g2305) & (g2309)) + ((!g2022) & (nmi_i) & (!g2023) & (!g2029) & (!g2305) & (g2309)) + ((!g2022) & (nmi_i) & (!g2023) & (!g2029) & (g2305) & (g2309)) + ((!g2022) & (nmi_i) & (!g2023) & (g2029) & (g2305) & (!g2309)) + ((!g2022) & (nmi_i) & (!g2023) & (g2029) & (g2305) & (g2309)) + ((!g2022) & (nmi_i) & (g2023) & (!g2029) & (!g2305) & (g2309)) + ((!g2022) & (nmi_i) & (g2023) & (!g2029) & (g2305) & (g2309)) + ((!g2022) & (nmi_i) & (g2023) & (g2029) & (g2305) & (!g2309)) + ((!g2022) & (nmi_i) & (g2023) & (g2029) & (g2305) & (g2309)) + ((g2022) & (!nmi_i) & (!g2023) & (!g2029) & (!g2305) & (g2309)) + ((g2022) & (!nmi_i) & (!g2023) & (!g2029) & (g2305) & (g2309)) + ((g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2305) & (!g2309)) + ((g2022) & (!nmi_i) & (!g2023) & (g2029) & (g2305) & (g2309)));
	assign g2311 = (((!g123) & (!intr_i) & (!g2039) & (!g2056) & (!g2057) & (g2310)) + ((!g123) & (!intr_i) & (!g2039) & (!g2056) & (g2057) & (g2310)) + ((!g123) & (!intr_i) & (!g2039) & (g2056) & (!g2057) & (g2310)) + ((!g123) & (!intr_i) & (!g2039) & (g2056) & (g2057) & (g2310)) + ((!g123) & (!intr_i) & (g2039) & (!g2056) & (!g2057) & (g2310)) + ((!g123) & (!intr_i) & (g2039) & (!g2056) & (g2057) & (g2310)) + ((!g123) & (!intr_i) & (g2039) & (g2056) & (!g2057) & (g2310)) + ((!g123) & (!intr_i) & (g2039) & (g2056) & (g2057) & (g2310)) + ((!g123) & (intr_i) & (!g2039) & (!g2056) & (!g2057) & (g2310)) + ((!g123) & (intr_i) & (!g2039) & (!g2056) & (g2057) & (g2310)) + ((!g123) & (intr_i) & (!g2039) & (g2056) & (!g2057) & (g2310)) + ((!g123) & (intr_i) & (g2039) & (!g2056) & (!g2057) & (g2310)) + ((!g123) & (intr_i) & (g2039) & (g2056) & (!g2057) & (g2310)));
	assign g2313 = (((!sk[25]) & (g2114) & (!g2289)) + ((!sk[25]) & (g2114) & (g2289)) + ((sk[25]) & (!g2114) & (g2289)) + ((sk[25]) & (g2114) & (!g2289)));
	assign g2314 = (((!g2073) & (!g2076) & (g2106) & (g2113) & (g2238) & (g2313)) + ((!g2073) & (g2076) & (!g2106) & (g2113) & (g2238) & (g2313)) + ((!g2073) & (g2076) & (g2106) & (g2113) & (!g2238) & (g2313)) + ((!g2073) & (g2076) & (g2106) & (g2113) & (g2238) & (g2313)) + ((g2073) & (!g2076) & (!g2106) & (g2113) & (!g2238) & (g2313)) + ((g2073) & (!g2076) & (!g2106) & (g2113) & (g2238) & (g2313)) + ((g2073) & (!g2076) & (g2106) & (!g2113) & (g2238) & (g2313)) + ((g2073) & (!g2076) & (g2106) & (g2113) & (!g2238) & (g2313)) + ((g2073) & (!g2076) & (g2106) & (g2113) & (g2238) & (g2313)) + ((g2073) & (g2076) & (!g2106) & (!g2113) & (g2238) & (g2313)) + ((g2073) & (g2076) & (!g2106) & (g2113) & (!g2238) & (g2313)) + ((g2073) & (g2076) & (!g2106) & (g2113) & (g2238) & (g2313)) + ((g2073) & (g2076) & (g2106) & (!g2113) & (!g2238) & (g2313)) + ((g2073) & (g2076) & (g2106) & (!g2113) & (g2238) & (g2313)) + ((g2073) & (g2076) & (g2106) & (g2113) & (!g2238) & (g2313)) + ((g2073) & (g2076) & (g2106) & (g2113) & (g2238) & (g2313)));
	assign g2315 = (((!g2115) & (!g2312) & (!sk[27]) & (!g2314) & (g2295)) + ((!g2115) & (!g2312) & (!sk[27]) & (g2314) & (!g2295)) + ((!g2115) & (!g2312) & (!sk[27]) & (g2314) & (g2295)) + ((!g2115) & (!g2312) & (sk[27]) & (!g2314) & (g2295)) + ((!g2115) & (!g2312) & (sk[27]) & (g2314) & (!g2295)) + ((!g2115) & (!g2312) & (sk[27]) & (g2314) & (g2295)) + ((!g2115) & (g2312) & (!sk[27]) & (!g2314) & (!g2295)) + ((!g2115) & (g2312) & (!sk[27]) & (!g2314) & (g2295)) + ((!g2115) & (g2312) & (!sk[27]) & (g2314) & (!g2295)) + ((!g2115) & (g2312) & (!sk[27]) & (g2314) & (g2295)) + ((!g2115) & (g2312) & (sk[27]) & (!g2314) & (!g2295)) + ((g2115) & (!g2312) & (!sk[27]) & (!g2314) & (g2295)) + ((g2115) & (!g2312) & (!sk[27]) & (g2314) & (!g2295)) + ((g2115) & (!g2312) & (!sk[27]) & (g2314) & (g2295)) + ((g2115) & (!g2312) & (sk[27]) & (!g2314) & (!g2295)) + ((g2115) & (g2312) & (!sk[27]) & (!g2314) & (!g2295)) + ((g2115) & (g2312) & (!sk[27]) & (!g2314) & (g2295)) + ((g2115) & (g2312) & (!sk[27]) & (g2314) & (!g2295)) + ((g2115) & (g2312) & (!sk[27]) & (g2314) & (g2295)) + ((g2115) & (g2312) & (sk[27]) & (!g2314) & (g2295)) + ((g2115) & (g2312) & (sk[27]) & (g2314) & (!g2295)) + ((g2115) & (g2312) & (sk[27]) & (g2314) & (g2295)));
	assign g2316 = (((!sk[28]) & (!g2266) & (!g2267) & (!g2290) & (g2315)) + ((!sk[28]) & (!g2266) & (!g2267) & (g2290) & (!g2315)) + ((!sk[28]) & (!g2266) & (!g2267) & (g2290) & (g2315)) + ((!sk[28]) & (!g2266) & (g2267) & (!g2290) & (!g2315)) + ((!sk[28]) & (!g2266) & (g2267) & (!g2290) & (g2315)) + ((!sk[28]) & (!g2266) & (g2267) & (g2290) & (!g2315)) + ((!sk[28]) & (!g2266) & (g2267) & (g2290) & (g2315)) + ((!sk[28]) & (g2266) & (!g2267) & (!g2290) & (g2315)) + ((!sk[28]) & (g2266) & (!g2267) & (g2290) & (!g2315)) + ((!sk[28]) & (g2266) & (!g2267) & (g2290) & (g2315)) + ((!sk[28]) & (g2266) & (g2267) & (!g2290) & (!g2315)) + ((!sk[28]) & (g2266) & (g2267) & (!g2290) & (g2315)) + ((!sk[28]) & (g2266) & (g2267) & (g2290) & (!g2315)) + ((!sk[28]) & (g2266) & (g2267) & (g2290) & (g2315)) + ((sk[28]) & (!g2266) & (!g2267) & (!g2290) & (g2315)) + ((sk[28]) & (!g2266) & (!g2267) & (g2290) & (g2315)) + ((sk[28]) & (!g2266) & (g2267) & (!g2290) & (g2315)) + ((sk[28]) & (!g2266) & (g2267) & (g2290) & (g2315)) + ((sk[28]) & (g2266) & (!g2267) & (!g2290) & (g2315)) + ((sk[28]) & (g2266) & (!g2267) & (g2290) & (g2315)) + ((sk[28]) & (g2266) & (g2267) & (!g2290) & (g2315)) + ((sk[28]) & (g2266) & (g2267) & (g2290) & (!g2315)));
	assign g2317 = (((!g2289) & (sk[29]) & (g2114)) + ((g2289) & (!sk[29]) & (!g2114)) + ((g2289) & (!sk[29]) & (g2114)));
	assign g2318 = (((!g2115) & (sk[30]) & (!g2312)) + ((g2115) & (!sk[30]) & (!g2312)) + ((g2115) & (!sk[30]) & (g2312)) + ((g2115) & (sk[30]) & (g2312)));
	assign g2319 = (((!g2291) & (!sk[31]) & (!g2292) & (!g2293) & (g2317) & (!g2318)) + ((!g2291) & (!sk[31]) & (!g2292) & (!g2293) & (g2317) & (g2318)) + ((!g2291) & (!sk[31]) & (!g2292) & (g2293) & (!g2317) & (!g2318)) + ((!g2291) & (!sk[31]) & (!g2292) & (g2293) & (!g2317) & (g2318)) + ((!g2291) & (!sk[31]) & (!g2292) & (g2293) & (g2317) & (!g2318)) + ((!g2291) & (!sk[31]) & (!g2292) & (g2293) & (g2317) & (g2318)) + ((!g2291) & (!sk[31]) & (g2292) & (!g2293) & (!g2317) & (!g2318)) + ((!g2291) & (!sk[31]) & (g2292) & (!g2293) & (!g2317) & (g2318)) + ((!g2291) & (!sk[31]) & (g2292) & (!g2293) & (g2317) & (!g2318)) + ((!g2291) & (!sk[31]) & (g2292) & (!g2293) & (g2317) & (g2318)) + ((!g2291) & (!sk[31]) & (g2292) & (g2293) & (!g2317) & (!g2318)) + ((!g2291) & (!sk[31]) & (g2292) & (g2293) & (!g2317) & (g2318)) + ((!g2291) & (!sk[31]) & (g2292) & (g2293) & (g2317) & (!g2318)) + ((!g2291) & (!sk[31]) & (g2292) & (g2293) & (g2317) & (g2318)) + ((!g2291) & (sk[31]) & (!g2292) & (!g2293) & (!g2317) & (g2318)) + ((!g2291) & (sk[31]) & (!g2292) & (!g2293) & (g2317) & (!g2318)) + ((!g2291) & (sk[31]) & (!g2292) & (g2293) & (!g2317) & (g2318)) + ((!g2291) & (sk[31]) & (!g2292) & (g2293) & (g2317) & (!g2318)) + ((!g2291) & (sk[31]) & (g2292) & (!g2293) & (!g2317) & (g2318)) + ((!g2291) & (sk[31]) & (g2292) & (!g2293) & (g2317) & (!g2318)) + ((!g2291) & (sk[31]) & (g2292) & (g2293) & (!g2317) & (!g2318)) + ((!g2291) & (sk[31]) & (g2292) & (g2293) & (g2317) & (g2318)) + ((g2291) & (!sk[31]) & (!g2292) & (!g2293) & (g2317) & (!g2318)) + ((g2291) & (!sk[31]) & (!g2292) & (!g2293) & (g2317) & (g2318)) + ((g2291) & (!sk[31]) & (!g2292) & (g2293) & (!g2317) & (!g2318)) + ((g2291) & (!sk[31]) & (!g2292) & (g2293) & (!g2317) & (g2318)) + ((g2291) & (!sk[31]) & (!g2292) & (g2293) & (g2317) & (!g2318)) + ((g2291) & (!sk[31]) & (!g2292) & (g2293) & (g2317) & (g2318)) + ((g2291) & (!sk[31]) & (g2292) & (!g2293) & (!g2317) & (!g2318)) + ((g2291) & (!sk[31]) & (g2292) & (!g2293) & (!g2317) & (g2318)) + ((g2291) & (!sk[31]) & (g2292) & (!g2293) & (g2317) & (!g2318)) + ((g2291) & (!sk[31]) & (g2292) & (!g2293) & (g2317) & (g2318)) + ((g2291) & (!sk[31]) & (g2292) & (g2293) & (!g2317) & (!g2318)) + ((g2291) & (!sk[31]) & (g2292) & (g2293) & (!g2317) & (g2318)) + ((g2291) & (!sk[31]) & (g2292) & (g2293) & (g2317) & (!g2318)) + ((g2291) & (!sk[31]) & (g2292) & (g2293) & (g2317) & (g2318)) + ((g2291) & (sk[31]) & (!g2292) & (!g2293) & (!g2317) & (g2318)) + ((g2291) & (sk[31]) & (!g2292) & (!g2293) & (g2317) & (!g2318)) + ((g2291) & (sk[31]) & (!g2292) & (g2293) & (!g2317) & (!g2318)) + ((g2291) & (sk[31]) & (!g2292) & (g2293) & (g2317) & (g2318)) + ((g2291) & (sk[31]) & (g2292) & (!g2293) & (!g2317) & (!g2318)) + ((g2291) & (sk[31]) & (g2292) & (!g2293) & (g2317) & (g2318)) + ((g2291) & (sk[31]) & (g2292) & (g2293) & (!g2317) & (!g2318)) + ((g2291) & (sk[31]) & (g2292) & (g2293) & (g2317) & (g2318)));
	assign g2320 = (((!g2115) & (!g2114) & (!g2113) & (g2106) & (g2071) & (g2074)) + ((!g2115) & (!g2114) & (g2113) & (!g2106) & (!g2071) & (g2074)) + ((!g2115) & (!g2114) & (g2113) & (g2106) & (!g2071) & (g2074)) + ((!g2115) & (!g2114) & (g2113) & (g2106) & (g2071) & (g2074)) + ((!g2115) & (g2114) & (!g2113) & (!g2106) & (g2071) & (!g2074)) + ((!g2115) & (g2114) & (!g2113) & (g2106) & (g2071) & (!g2074)) + ((!g2115) & (g2114) & (!g2113) & (g2106) & (g2071) & (g2074)) + ((!g2115) & (g2114) & (g2113) & (!g2106) & (!g2071) & (g2074)) + ((!g2115) & (g2114) & (g2113) & (!g2106) & (g2071) & (!g2074)) + ((!g2115) & (g2114) & (g2113) & (g2106) & (!g2071) & (g2074)) + ((!g2115) & (g2114) & (g2113) & (g2106) & (g2071) & (!g2074)) + ((!g2115) & (g2114) & (g2113) & (g2106) & (g2071) & (g2074)) + ((g2115) & (!g2114) & (!g2113) & (!g2106) & (!g2071) & (!g2074)) + ((g2115) & (!g2114) & (!g2113) & (g2106) & (!g2071) & (!g2074)) + ((g2115) & (!g2114) & (!g2113) & (g2106) & (g2071) & (g2074)) + ((g2115) & (!g2114) & (g2113) & (!g2106) & (!g2071) & (!g2074)) + ((g2115) & (!g2114) & (g2113) & (!g2106) & (!g2071) & (g2074)) + ((g2115) & (!g2114) & (g2113) & (g2106) & (!g2071) & (!g2074)) + ((g2115) & (!g2114) & (g2113) & (g2106) & (!g2071) & (g2074)) + ((g2115) & (!g2114) & (g2113) & (g2106) & (g2071) & (g2074)) + ((g2115) & (g2114) & (!g2113) & (!g2106) & (!g2071) & (!g2074)) + ((g2115) & (g2114) & (!g2113) & (!g2106) & (g2071) & (!g2074)) + ((g2115) & (g2114) & (!g2113) & (g2106) & (!g2071) & (!g2074)) + ((g2115) & (g2114) & (!g2113) & (g2106) & (g2071) & (!g2074)) + ((g2115) & (g2114) & (!g2113) & (g2106) & (g2071) & (g2074)) + ((g2115) & (g2114) & (g2113) & (!g2106) & (!g2071) & (!g2074)) + ((g2115) & (g2114) & (g2113) & (!g2106) & (!g2071) & (g2074)) + ((g2115) & (g2114) & (g2113) & (!g2106) & (g2071) & (!g2074)) + ((g2115) & (g2114) & (g2113) & (g2106) & (!g2071) & (!g2074)) + ((g2115) & (g2114) & (g2113) & (g2106) & (!g2071) & (g2074)) + ((g2115) & (g2114) & (g2113) & (g2106) & (g2071) & (!g2074)) + ((g2115) & (g2114) & (g2113) & (g2106) & (g2071) & (g2074)));
	assign g2321 = (((!g2076) & (!sk[33]) & (!g2077) & (!g2211) & (g2320)) + ((!g2076) & (!sk[33]) & (!g2077) & (g2211) & (!g2320)) + ((!g2076) & (!sk[33]) & (!g2077) & (g2211) & (g2320)) + ((!g2076) & (!sk[33]) & (g2077) & (!g2211) & (!g2320)) + ((!g2076) & (!sk[33]) & (g2077) & (!g2211) & (g2320)) + ((!g2076) & (!sk[33]) & (g2077) & (g2211) & (!g2320)) + ((!g2076) & (!sk[33]) & (g2077) & (g2211) & (g2320)) + ((!g2076) & (sk[33]) & (!g2077) & (!g2211) & (g2320)) + ((!g2076) & (sk[33]) & (!g2077) & (g2211) & (g2320)) + ((!g2076) & (sk[33]) & (g2077) & (g2211) & (!g2320)) + ((!g2076) & (sk[33]) & (g2077) & (g2211) & (g2320)) + ((g2076) & (!sk[33]) & (!g2077) & (!g2211) & (g2320)) + ((g2076) & (!sk[33]) & (!g2077) & (g2211) & (!g2320)) + ((g2076) & (!sk[33]) & (!g2077) & (g2211) & (g2320)) + ((g2076) & (!sk[33]) & (g2077) & (!g2211) & (!g2320)) + ((g2076) & (!sk[33]) & (g2077) & (!g2211) & (g2320)) + ((g2076) & (!sk[33]) & (g2077) & (g2211) & (!g2320)) + ((g2076) & (!sk[33]) & (g2077) & (g2211) & (g2320)));
	assign g2322 = (((!g2220) & (!g2223) & (!g2222) & (g2215) & (g2076) & (g2077)) + ((!g2220) & (!g2223) & (g2222) & (!g2215) & (!g2076) & (g2077)) + ((!g2220) & (!g2223) & (g2222) & (g2215) & (!g2076) & (g2077)) + ((!g2220) & (!g2223) & (g2222) & (g2215) & (g2076) & (g2077)) + ((!g2220) & (g2223) & (!g2222) & (!g2215) & (g2076) & (!g2077)) + ((!g2220) & (g2223) & (!g2222) & (g2215) & (g2076) & (!g2077)) + ((!g2220) & (g2223) & (!g2222) & (g2215) & (g2076) & (g2077)) + ((!g2220) & (g2223) & (g2222) & (!g2215) & (!g2076) & (g2077)) + ((!g2220) & (g2223) & (g2222) & (!g2215) & (g2076) & (!g2077)) + ((!g2220) & (g2223) & (g2222) & (g2215) & (!g2076) & (g2077)) + ((!g2220) & (g2223) & (g2222) & (g2215) & (g2076) & (!g2077)) + ((!g2220) & (g2223) & (g2222) & (g2215) & (g2076) & (g2077)) + ((g2220) & (!g2223) & (!g2222) & (!g2215) & (!g2076) & (!g2077)) + ((g2220) & (!g2223) & (!g2222) & (g2215) & (!g2076) & (!g2077)) + ((g2220) & (!g2223) & (!g2222) & (g2215) & (g2076) & (g2077)) + ((g2220) & (!g2223) & (g2222) & (!g2215) & (!g2076) & (!g2077)) + ((g2220) & (!g2223) & (g2222) & (!g2215) & (!g2076) & (g2077)) + ((g2220) & (!g2223) & (g2222) & (g2215) & (!g2076) & (!g2077)) + ((g2220) & (!g2223) & (g2222) & (g2215) & (!g2076) & (g2077)) + ((g2220) & (!g2223) & (g2222) & (g2215) & (g2076) & (g2077)) + ((g2220) & (g2223) & (!g2222) & (!g2215) & (!g2076) & (!g2077)) + ((g2220) & (g2223) & (!g2222) & (!g2215) & (g2076) & (!g2077)) + ((g2220) & (g2223) & (!g2222) & (g2215) & (!g2076) & (!g2077)) + ((g2220) & (g2223) & (!g2222) & (g2215) & (g2076) & (!g2077)) + ((g2220) & (g2223) & (!g2222) & (g2215) & (g2076) & (g2077)) + ((g2220) & (g2223) & (g2222) & (!g2215) & (!g2076) & (!g2077)) + ((g2220) & (g2223) & (g2222) & (!g2215) & (!g2076) & (g2077)) + ((g2220) & (g2223) & (g2222) & (!g2215) & (g2076) & (!g2077)) + ((g2220) & (g2223) & (g2222) & (g2215) & (!g2076) & (!g2077)) + ((g2220) & (g2223) & (g2222) & (g2215) & (!g2076) & (g2077)) + ((g2220) & (g2223) & (g2222) & (g2215) & (g2076) & (!g2077)) + ((g2220) & (g2223) & (g2222) & (g2215) & (g2076) & (g2077)));
	assign g2323 = (((!g2217) & (!g2218) & (!g2216) & (g2192) & (g2076) & (g2077)) + ((!g2217) & (!g2218) & (g2216) & (!g2192) & (!g2076) & (g2077)) + ((!g2217) & (!g2218) & (g2216) & (g2192) & (!g2076) & (g2077)) + ((!g2217) & (!g2218) & (g2216) & (g2192) & (g2076) & (g2077)) + ((!g2217) & (g2218) & (!g2216) & (!g2192) & (g2076) & (!g2077)) + ((!g2217) & (g2218) & (!g2216) & (g2192) & (g2076) & (!g2077)) + ((!g2217) & (g2218) & (!g2216) & (g2192) & (g2076) & (g2077)) + ((!g2217) & (g2218) & (g2216) & (!g2192) & (!g2076) & (g2077)) + ((!g2217) & (g2218) & (g2216) & (!g2192) & (g2076) & (!g2077)) + ((!g2217) & (g2218) & (g2216) & (g2192) & (!g2076) & (g2077)) + ((!g2217) & (g2218) & (g2216) & (g2192) & (g2076) & (!g2077)) + ((!g2217) & (g2218) & (g2216) & (g2192) & (g2076) & (g2077)) + ((g2217) & (!g2218) & (!g2216) & (!g2192) & (!g2076) & (!g2077)) + ((g2217) & (!g2218) & (!g2216) & (g2192) & (!g2076) & (!g2077)) + ((g2217) & (!g2218) & (!g2216) & (g2192) & (g2076) & (g2077)) + ((g2217) & (!g2218) & (g2216) & (!g2192) & (!g2076) & (!g2077)) + ((g2217) & (!g2218) & (g2216) & (!g2192) & (!g2076) & (g2077)) + ((g2217) & (!g2218) & (g2216) & (g2192) & (!g2076) & (!g2077)) + ((g2217) & (!g2218) & (g2216) & (g2192) & (!g2076) & (g2077)) + ((g2217) & (!g2218) & (g2216) & (g2192) & (g2076) & (g2077)) + ((g2217) & (g2218) & (!g2216) & (!g2192) & (!g2076) & (!g2077)) + ((g2217) & (g2218) & (!g2216) & (!g2192) & (g2076) & (!g2077)) + ((g2217) & (g2218) & (!g2216) & (g2192) & (!g2076) & (!g2077)) + ((g2217) & (g2218) & (!g2216) & (g2192) & (g2076) & (!g2077)) + ((g2217) & (g2218) & (!g2216) & (g2192) & (g2076) & (g2077)) + ((g2217) & (g2218) & (g2216) & (!g2192) & (!g2076) & (!g2077)) + ((g2217) & (g2218) & (g2216) & (!g2192) & (!g2076) & (g2077)) + ((g2217) & (g2218) & (g2216) & (!g2192) & (g2076) & (!g2077)) + ((g2217) & (g2218) & (g2216) & (g2192) & (!g2076) & (!g2077)) + ((g2217) & (g2218) & (g2216) & (g2192) & (!g2076) & (g2077)) + ((g2217) & (g2218) & (g2216) & (g2192) & (g2076) & (!g2077)) + ((g2217) & (g2218) & (g2216) & (g2192) & (g2076) & (g2077)));
	assign g2324 = (((!g2073) & (!g2080) & (!g2125) & (g2321) & (!g2322) & (!g2323)) + ((!g2073) & (!g2080) & (!g2125) & (g2321) & (!g2322) & (g2323)) + ((!g2073) & (!g2080) & (!g2125) & (g2321) & (g2322) & (!g2323)) + ((!g2073) & (!g2080) & (!g2125) & (g2321) & (g2322) & (g2323)) + ((!g2073) & (!g2080) & (g2125) & (!g2321) & (g2322) & (!g2323)) + ((!g2073) & (!g2080) & (g2125) & (!g2321) & (g2322) & (g2323)) + ((!g2073) & (!g2080) & (g2125) & (g2321) & (g2322) & (!g2323)) + ((!g2073) & (!g2080) & (g2125) & (g2321) & (g2322) & (g2323)) + ((!g2073) & (g2080) & (!g2125) & (g2321) & (!g2322) & (!g2323)) + ((!g2073) & (g2080) & (!g2125) & (g2321) & (!g2322) & (g2323)) + ((!g2073) & (g2080) & (!g2125) & (g2321) & (g2322) & (!g2323)) + ((!g2073) & (g2080) & (!g2125) & (g2321) & (g2322) & (g2323)) + ((!g2073) & (g2080) & (g2125) & (!g2321) & (g2322) & (!g2323)) + ((!g2073) & (g2080) & (g2125) & (!g2321) & (g2322) & (g2323)) + ((!g2073) & (g2080) & (g2125) & (g2321) & (g2322) & (!g2323)) + ((!g2073) & (g2080) & (g2125) & (g2321) & (g2322) & (g2323)) + ((g2073) & (!g2080) & (g2125) & (!g2321) & (!g2322) & (g2323)) + ((g2073) & (!g2080) & (g2125) & (!g2321) & (g2322) & (g2323)) + ((g2073) & (!g2080) & (g2125) & (g2321) & (!g2322) & (g2323)) + ((g2073) & (!g2080) & (g2125) & (g2321) & (g2322) & (g2323)) + ((g2073) & (g2080) & (!g2125) & (g2321) & (!g2322) & (!g2323)) + ((g2073) & (g2080) & (!g2125) & (g2321) & (!g2322) & (g2323)) + ((g2073) & (g2080) & (!g2125) & (g2321) & (g2322) & (!g2323)) + ((g2073) & (g2080) & (!g2125) & (g2321) & (g2322) & (g2323)) + ((g2073) & (g2080) & (g2125) & (!g2321) & (!g2322) & (g2323)) + ((g2073) & (g2080) & (g2125) & (!g2321) & (g2322) & (g2323)) + ((g2073) & (g2080) & (g2125) & (g2321) & (!g2322) & (g2323)) + ((g2073) & (g2080) & (g2125) & (g2321) & (g2322) & (g2323)));
	assign g2325 = (((!g2312) & (!g2115) & (!g2124) & (!g2264) & (!g3712) & (!g2324)) + ((!g2312) & (!g2115) & (!g2124) & (!g2264) & (g3712) & (!g2324)) + ((!g2312) & (!g2115) & (!g2124) & (g2264) & (!g3712) & (!g2324)) + ((!g2312) & (!g2115) & (!g2124) & (g2264) & (!g3712) & (g2324)) + ((!g2312) & (!g2115) & (g2124) & (!g2264) & (!g3712) & (!g2324)) + ((!g2312) & (!g2115) & (g2124) & (!g2264) & (!g3712) & (g2324)) + ((!g2312) & (!g2115) & (g2124) & (!g2264) & (g3712) & (!g2324)) + ((!g2312) & (!g2115) & (g2124) & (!g2264) & (g3712) & (g2324)) + ((!g2312) & (!g2115) & (g2124) & (g2264) & (!g3712) & (!g2324)) + ((!g2312) & (!g2115) & (g2124) & (g2264) & (!g3712) & (g2324)) + ((!g2312) & (!g2115) & (g2124) & (g2264) & (g3712) & (!g2324)) + ((!g2312) & (!g2115) & (g2124) & (g2264) & (g3712) & (g2324)) + ((!g2312) & (g2115) & (!g2124) & (!g2264) & (!g3712) & (!g2324)) + ((!g2312) & (g2115) & (!g2124) & (!g2264) & (g3712) & (!g2324)) + ((!g2312) & (g2115) & (!g2124) & (g2264) & (!g3712) & (!g2324)) + ((!g2312) & (g2115) & (!g2124) & (g2264) & (!g3712) & (g2324)) + ((g2312) & (!g2115) & (!g2124) & (!g2264) & (!g3712) & (!g2324)) + ((g2312) & (!g2115) & (!g2124) & (!g2264) & (g3712) & (!g2324)) + ((g2312) & (!g2115) & (!g2124) & (g2264) & (!g3712) & (!g2324)) + ((g2312) & (!g2115) & (!g2124) & (g2264) & (!g3712) & (g2324)) + ((g2312) & (g2115) & (!g2124) & (!g2264) & (!g3712) & (!g2324)) + ((g2312) & (g2115) & (!g2124) & (!g2264) & (g3712) & (!g2324)) + ((g2312) & (g2115) & (!g2124) & (g2264) & (!g3712) & (!g2324)) + ((g2312) & (g2115) & (!g2124) & (g2264) & (!g3712) & (g2324)) + ((g2312) & (g2115) & (g2124) & (g2264) & (!g3712) & (!g2324)) + ((g2312) & (g2115) & (g2124) & (g2264) & (!g3712) & (g2324)) + ((g2312) & (g2115) & (g2124) & (g2264) & (g3712) & (!g2324)) + ((g2312) & (g2115) & (g2124) & (g2264) & (g3712) & (g2324)));
	assign g2326 = (((!dmem_dat_ix6x) & (!dmem_dat_ix14x) & (!dmem_dat_ix30x) & (dmem_dat_ix22x) & (g2206) & (g2207)) + ((!dmem_dat_ix6x) & (!dmem_dat_ix14x) & (dmem_dat_ix30x) & (!dmem_dat_ix22x) & (!g2206) & (g2207)) + ((!dmem_dat_ix6x) & (!dmem_dat_ix14x) & (dmem_dat_ix30x) & (dmem_dat_ix22x) & (!g2206) & (g2207)) + ((!dmem_dat_ix6x) & (!dmem_dat_ix14x) & (dmem_dat_ix30x) & (dmem_dat_ix22x) & (g2206) & (g2207)) + ((!dmem_dat_ix6x) & (dmem_dat_ix14x) & (!dmem_dat_ix30x) & (!dmem_dat_ix22x) & (g2206) & (!g2207)) + ((!dmem_dat_ix6x) & (dmem_dat_ix14x) & (!dmem_dat_ix30x) & (dmem_dat_ix22x) & (g2206) & (!g2207)) + ((!dmem_dat_ix6x) & (dmem_dat_ix14x) & (!dmem_dat_ix30x) & (dmem_dat_ix22x) & (g2206) & (g2207)) + ((!dmem_dat_ix6x) & (dmem_dat_ix14x) & (dmem_dat_ix30x) & (!dmem_dat_ix22x) & (!g2206) & (g2207)) + ((!dmem_dat_ix6x) & (dmem_dat_ix14x) & (dmem_dat_ix30x) & (!dmem_dat_ix22x) & (g2206) & (!g2207)) + ((!dmem_dat_ix6x) & (dmem_dat_ix14x) & (dmem_dat_ix30x) & (dmem_dat_ix22x) & (!g2206) & (g2207)) + ((!dmem_dat_ix6x) & (dmem_dat_ix14x) & (dmem_dat_ix30x) & (dmem_dat_ix22x) & (g2206) & (!g2207)) + ((!dmem_dat_ix6x) & (dmem_dat_ix14x) & (dmem_dat_ix30x) & (dmem_dat_ix22x) & (g2206) & (g2207)) + ((dmem_dat_ix6x) & (!dmem_dat_ix14x) & (!dmem_dat_ix30x) & (!dmem_dat_ix22x) & (!g2206) & (!g2207)) + ((dmem_dat_ix6x) & (!dmem_dat_ix14x) & (!dmem_dat_ix30x) & (dmem_dat_ix22x) & (!g2206) & (!g2207)) + ((dmem_dat_ix6x) & (!dmem_dat_ix14x) & (!dmem_dat_ix30x) & (dmem_dat_ix22x) & (g2206) & (g2207)) + ((dmem_dat_ix6x) & (!dmem_dat_ix14x) & (dmem_dat_ix30x) & (!dmem_dat_ix22x) & (!g2206) & (!g2207)) + ((dmem_dat_ix6x) & (!dmem_dat_ix14x) & (dmem_dat_ix30x) & (!dmem_dat_ix22x) & (!g2206) & (g2207)) + ((dmem_dat_ix6x) & (!dmem_dat_ix14x) & (dmem_dat_ix30x) & (dmem_dat_ix22x) & (!g2206) & (!g2207)) + ((dmem_dat_ix6x) & (!dmem_dat_ix14x) & (dmem_dat_ix30x) & (dmem_dat_ix22x) & (!g2206) & (g2207)) + ((dmem_dat_ix6x) & (!dmem_dat_ix14x) & (dmem_dat_ix30x) & (dmem_dat_ix22x) & (g2206) & (g2207)) + ((dmem_dat_ix6x) & (dmem_dat_ix14x) & (!dmem_dat_ix30x) & (!dmem_dat_ix22x) & (!g2206) & (!g2207)) + ((dmem_dat_ix6x) & (dmem_dat_ix14x) & (!dmem_dat_ix30x) & (!dmem_dat_ix22x) & (g2206) & (!g2207)) + ((dmem_dat_ix6x) & (dmem_dat_ix14x) & (!dmem_dat_ix30x) & (dmem_dat_ix22x) & (!g2206) & (!g2207)) + ((dmem_dat_ix6x) & (dmem_dat_ix14x) & (!dmem_dat_ix30x) & (dmem_dat_ix22x) & (g2206) & (!g2207)) + ((dmem_dat_ix6x) & (dmem_dat_ix14x) & (!dmem_dat_ix30x) & (dmem_dat_ix22x) & (g2206) & (g2207)) + ((dmem_dat_ix6x) & (dmem_dat_ix14x) & (dmem_dat_ix30x) & (!dmem_dat_ix22x) & (!g2206) & (!g2207)) + ((dmem_dat_ix6x) & (dmem_dat_ix14x) & (dmem_dat_ix30x) & (!dmem_dat_ix22x) & (!g2206) & (g2207)) + ((dmem_dat_ix6x) & (dmem_dat_ix14x) & (dmem_dat_ix30x) & (!dmem_dat_ix22x) & (g2206) & (!g2207)) + ((dmem_dat_ix6x) & (dmem_dat_ix14x) & (dmem_dat_ix30x) & (dmem_dat_ix22x) & (!g2206) & (!g2207)) + ((dmem_dat_ix6x) & (dmem_dat_ix14x) & (dmem_dat_ix30x) & (dmem_dat_ix22x) & (!g2206) & (g2207)) + ((dmem_dat_ix6x) & (dmem_dat_ix14x) & (dmem_dat_ix30x) & (dmem_dat_ix22x) & (g2206) & (!g2207)) + ((dmem_dat_ix6x) & (dmem_dat_ix14x) & (dmem_dat_ix30x) & (dmem_dat_ix22x) & (g2206) & (g2207)));
	assign g2327 = (((!dmem_dat_ix6x) & (!dmem_dat_ix22x) & (!g2128) & (!sk[39]) & (g2129)) + ((!dmem_dat_ix6x) & (!dmem_dat_ix22x) & (g2128) & (!sk[39]) & (!g2129)) + ((!dmem_dat_ix6x) & (!dmem_dat_ix22x) & (g2128) & (!sk[39]) & (g2129)) + ((!dmem_dat_ix6x) & (dmem_dat_ix22x) & (!g2128) & (!sk[39]) & (!g2129)) + ((!dmem_dat_ix6x) & (dmem_dat_ix22x) & (!g2128) & (!sk[39]) & (g2129)) + ((!dmem_dat_ix6x) & (dmem_dat_ix22x) & (!g2128) & (sk[39]) & (!g2129)) + ((!dmem_dat_ix6x) & (dmem_dat_ix22x) & (g2128) & (!sk[39]) & (!g2129)) + ((!dmem_dat_ix6x) & (dmem_dat_ix22x) & (g2128) & (!sk[39]) & (g2129)) + ((dmem_dat_ix6x) & (!dmem_dat_ix22x) & (!g2128) & (!sk[39]) & (g2129)) + ((dmem_dat_ix6x) & (!dmem_dat_ix22x) & (!g2128) & (sk[39]) & (g2129)) + ((dmem_dat_ix6x) & (!dmem_dat_ix22x) & (g2128) & (!sk[39]) & (!g2129)) + ((dmem_dat_ix6x) & (!dmem_dat_ix22x) & (g2128) & (!sk[39]) & (g2129)) + ((dmem_dat_ix6x) & (dmem_dat_ix22x) & (!g2128) & (!sk[39]) & (!g2129)) + ((dmem_dat_ix6x) & (dmem_dat_ix22x) & (!g2128) & (!sk[39]) & (g2129)) + ((dmem_dat_ix6x) & (dmem_dat_ix22x) & (!g2128) & (sk[39]) & (!g2129)) + ((dmem_dat_ix6x) & (dmem_dat_ix22x) & (!g2128) & (sk[39]) & (g2129)) + ((dmem_dat_ix6x) & (dmem_dat_ix22x) & (g2128) & (!sk[39]) & (!g2129)) + ((dmem_dat_ix6x) & (dmem_dat_ix22x) & (g2128) & (!sk[39]) & (g2129)));
	assign g2328 = (((!g2325) & (!g2115) & (!g2326) & (!g2327) & (!g2281) & (!g75)) + ((!g2325) & (!g2115) & (!g2326) & (g2327) & (!g2281) & (!g75)) + ((!g2325) & (!g2115) & (!g2326) & (g2327) & (g2281) & (g75)) + ((!g2325) & (!g2115) & (g2326) & (!g2327) & (!g2281) & (!g75)) + ((!g2325) & (!g2115) & (g2326) & (!g2327) & (!g2281) & (g75)) + ((!g2325) & (!g2115) & (g2326) & (g2327) & (!g2281) & (!g75)) + ((!g2325) & (!g2115) & (g2326) & (g2327) & (!g2281) & (g75)) + ((!g2325) & (!g2115) & (g2326) & (g2327) & (g2281) & (g75)) + ((!g2325) & (g2115) & (!g2326) & (!g2327) & (!g2281) & (!g75)) + ((!g2325) & (g2115) & (!g2326) & (!g2327) & (g2281) & (!g75)) + ((!g2325) & (g2115) & (!g2326) & (g2327) & (!g2281) & (!g75)) + ((!g2325) & (g2115) & (!g2326) & (g2327) & (g2281) & (!g75)) + ((!g2325) & (g2115) & (!g2326) & (g2327) & (g2281) & (g75)) + ((!g2325) & (g2115) & (g2326) & (!g2327) & (!g2281) & (!g75)) + ((!g2325) & (g2115) & (g2326) & (!g2327) & (!g2281) & (g75)) + ((!g2325) & (g2115) & (g2326) & (!g2327) & (g2281) & (!g75)) + ((!g2325) & (g2115) & (g2326) & (g2327) & (!g2281) & (!g75)) + ((!g2325) & (g2115) & (g2326) & (g2327) & (!g2281) & (g75)) + ((!g2325) & (g2115) & (g2326) & (g2327) & (g2281) & (!g75)) + ((!g2325) & (g2115) & (g2326) & (g2327) & (g2281) & (g75)) + ((g2325) & (!g2115) & (!g2326) & (g2327) & (g2281) & (g75)) + ((g2325) & (!g2115) & (g2326) & (!g2327) & (!g2281) & (g75)) + ((g2325) & (!g2115) & (g2326) & (g2327) & (!g2281) & (g75)) + ((g2325) & (!g2115) & (g2326) & (g2327) & (g2281) & (g75)) + ((g2325) & (g2115) & (!g2326) & (!g2327) & (g2281) & (!g75)) + ((g2325) & (g2115) & (!g2326) & (g2327) & (g2281) & (!g75)) + ((g2325) & (g2115) & (!g2326) & (g2327) & (g2281) & (g75)) + ((g2325) & (g2115) & (g2326) & (!g2327) & (!g2281) & (g75)) + ((g2325) & (g2115) & (g2326) & (!g2327) & (g2281) & (!g75)) + ((g2325) & (g2115) & (g2326) & (g2327) & (!g2281) & (g75)) + ((g2325) & (g2115) & (g2326) & (g2327) & (g2281) & (!g75)) + ((g2325) & (g2115) & (g2326) & (g2327) & (g2281) & (g75)));
	assign g2329 = (((!g114) & (!g115) & (!sk[41]) & (!nmi_i) & (g2023)) + ((!g114) & (!g115) & (!sk[41]) & (nmi_i) & (!g2023)) + ((!g114) & (!g115) & (!sk[41]) & (nmi_i) & (g2023)) + ((!g114) & (!g115) & (sk[41]) & (!nmi_i) & (!g2023)) + ((!g114) & (g115) & (!sk[41]) & (!nmi_i) & (!g2023)) + ((!g114) & (g115) & (!sk[41]) & (!nmi_i) & (g2023)) + ((!g114) & (g115) & (!sk[41]) & (nmi_i) & (!g2023)) + ((!g114) & (g115) & (!sk[41]) & (nmi_i) & (g2023)) + ((!g114) & (g115) & (sk[41]) & (!nmi_i) & (!g2023)) + ((g114) & (!g115) & (!sk[41]) & (!nmi_i) & (g2023)) + ((g114) & (!g115) & (!sk[41]) & (nmi_i) & (!g2023)) + ((g114) & (!g115) & (!sk[41]) & (nmi_i) & (g2023)) + ((g114) & (!g115) & (sk[41]) & (!nmi_i) & (!g2023)) + ((g114) & (g115) & (!sk[41]) & (!nmi_i) & (!g2023)) + ((g114) & (g115) & (!sk[41]) & (!nmi_i) & (g2023)) + ((g114) & (g115) & (!sk[41]) & (nmi_i) & (!g2023)) + ((g114) & (g115) & (!sk[41]) & (nmi_i) & (g2023)) + ((g114) & (g115) & (sk[41]) & (!nmi_i) & (!g2023)) + ((g114) & (g115) & (sk[41]) & (!nmi_i) & (g2023)) + ((g114) & (g115) & (sk[41]) & (nmi_i) & (!g2023)) + ((g114) & (g115) & (sk[41]) & (nmi_i) & (g2023)));
	assign g2330 = (((!sk[42]) & (g2039) & (!g2056)) + ((!sk[42]) & (g2039) & (g2056)) + ((sk[42]) & (!g2039) & (!g2056)));
	assign g2331 = (((!g141) & (!g275) & (!sk[43]) & (!g319) & (g365) & (!g408)) + ((!g141) & (!g275) & (!sk[43]) & (!g319) & (g365) & (g408)) + ((!g141) & (!g275) & (!sk[43]) & (g319) & (!g365) & (!g408)) + ((!g141) & (!g275) & (!sk[43]) & (g319) & (!g365) & (g408)) + ((!g141) & (!g275) & (!sk[43]) & (g319) & (g365) & (!g408)) + ((!g141) & (!g275) & (!sk[43]) & (g319) & (g365) & (g408)) + ((!g141) & (g275) & (!sk[43]) & (!g319) & (!g365) & (!g408)) + ((!g141) & (g275) & (!sk[43]) & (!g319) & (!g365) & (g408)) + ((!g141) & (g275) & (!sk[43]) & (!g319) & (g365) & (!g408)) + ((!g141) & (g275) & (!sk[43]) & (!g319) & (g365) & (g408)) + ((!g141) & (g275) & (!sk[43]) & (g319) & (!g365) & (!g408)) + ((!g141) & (g275) & (!sk[43]) & (g319) & (!g365) & (g408)) + ((!g141) & (g275) & (!sk[43]) & (g319) & (g365) & (!g408)) + ((!g141) & (g275) & (!sk[43]) & (g319) & (g365) & (g408)) + ((g141) & (!g275) & (!sk[43]) & (!g319) & (g365) & (!g408)) + ((g141) & (!g275) & (!sk[43]) & (!g319) & (g365) & (g408)) + ((g141) & (!g275) & (!sk[43]) & (g319) & (!g365) & (!g408)) + ((g141) & (!g275) & (!sk[43]) & (g319) & (!g365) & (g408)) + ((g141) & (!g275) & (!sk[43]) & (g319) & (g365) & (!g408)) + ((g141) & (!g275) & (!sk[43]) & (g319) & (g365) & (g408)) + ((g141) & (g275) & (!sk[43]) & (!g319) & (!g365) & (!g408)) + ((g141) & (g275) & (!sk[43]) & (!g319) & (!g365) & (g408)) + ((g141) & (g275) & (!sk[43]) & (!g319) & (g365) & (!g408)) + ((g141) & (g275) & (!sk[43]) & (!g319) & (g365) & (g408)) + ((g141) & (g275) & (!sk[43]) & (g319) & (!g365) & (!g408)) + ((g141) & (g275) & (!sk[43]) & (g319) & (!g365) & (g408)) + ((g141) & (g275) & (!sk[43]) & (g319) & (g365) & (!g408)) + ((g141) & (g275) & (!sk[43]) & (g319) & (g365) & (g408)) + ((g141) & (g275) & (sk[43]) & (g319) & (g365) & (g408)));
	assign g2332 = (((!sk[44]) & (g453) & (!g2331)) + ((!sk[44]) & (g453) & (g2331)) + ((sk[44]) & (!g453) & (g2331)) + ((sk[44]) & (g453) & (!g2331)));
	assign g5031 = (((!sk[45]) & (!g2921) & (!g3066) & (g2333)) + ((!sk[45]) & (!g2921) & (g3066) & (!g2333)) + ((!sk[45]) & (!g2921) & (g3066) & (g2333)) + ((!sk[45]) & (g2921) & (!g3066) & (g2333)) + ((!sk[45]) & (g2921) & (g3066) & (!g2333)) + ((!sk[45]) & (g2921) & (g3066) & (g2333)) + ((sk[45]) & (!g2921) & (!g3066) & (g2333)) + ((sk[45]) & (!g2921) & (g3066) & (g2333)) + ((sk[45]) & (g2921) & (g3066) & (!g2333)) + ((sk[45]) & (g2921) & (g3066) & (g2333)));
	assign g2334 = (((!sk[46]) & (!g318) & (!g408) & (!g2307) & (g364) & (!g453)) + ((!sk[46]) & (!g318) & (!g408) & (!g2307) & (g364) & (g453)) + ((!sk[46]) & (!g318) & (!g408) & (g2307) & (!g364) & (!g453)) + ((!sk[46]) & (!g318) & (!g408) & (g2307) & (!g364) & (g453)) + ((!sk[46]) & (!g318) & (!g408) & (g2307) & (g364) & (!g453)) + ((!sk[46]) & (!g318) & (!g408) & (g2307) & (g364) & (g453)) + ((!sk[46]) & (!g318) & (g408) & (!g2307) & (!g364) & (!g453)) + ((!sk[46]) & (!g318) & (g408) & (!g2307) & (!g364) & (g453)) + ((!sk[46]) & (!g318) & (g408) & (!g2307) & (g364) & (!g453)) + ((!sk[46]) & (!g318) & (g408) & (!g2307) & (g364) & (g453)) + ((!sk[46]) & (!g318) & (g408) & (g2307) & (!g364) & (!g453)) + ((!sk[46]) & (!g318) & (g408) & (g2307) & (!g364) & (g453)) + ((!sk[46]) & (!g318) & (g408) & (g2307) & (g364) & (!g453)) + ((!sk[46]) & (!g318) & (g408) & (g2307) & (g364) & (g453)) + ((!sk[46]) & (g318) & (!g408) & (!g2307) & (g364) & (!g453)) + ((!sk[46]) & (g318) & (!g408) & (!g2307) & (g364) & (g453)) + ((!sk[46]) & (g318) & (!g408) & (g2307) & (!g364) & (!g453)) + ((!sk[46]) & (g318) & (!g408) & (g2307) & (!g364) & (g453)) + ((!sk[46]) & (g318) & (!g408) & (g2307) & (g364) & (!g453)) + ((!sk[46]) & (g318) & (!g408) & (g2307) & (g364) & (g453)) + ((!sk[46]) & (g318) & (g408) & (!g2307) & (!g364) & (!g453)) + ((!sk[46]) & (g318) & (g408) & (!g2307) & (!g364) & (g453)) + ((!sk[46]) & (g318) & (g408) & (!g2307) & (g364) & (!g453)) + ((!sk[46]) & (g318) & (g408) & (!g2307) & (g364) & (g453)) + ((!sk[46]) & (g318) & (g408) & (g2307) & (!g364) & (!g453)) + ((!sk[46]) & (g318) & (g408) & (g2307) & (!g364) & (g453)) + ((!sk[46]) & (g318) & (g408) & (g2307) & (g364) & (!g453)) + ((!sk[46]) & (g318) & (g408) & (g2307) & (g364) & (g453)) + ((sk[46]) & (!g318) & (!g408) & (!g2307) & (!g364) & (g453)) + ((sk[46]) & (!g318) & (!g408) & (!g2307) & (g364) & (!g453)) + ((sk[46]) & (!g318) & (!g408) & (g2307) & (!g364) & (g453)) + ((sk[46]) & (!g318) & (!g408) & (g2307) & (g364) & (!g453)) + ((sk[46]) & (!g318) & (g408) & (!g2307) & (!g364) & (g453)) + ((sk[46]) & (!g318) & (g408) & (!g2307) & (g364) & (!g453)) + ((sk[46]) & (!g318) & (g408) & (g2307) & (!g364) & (!g453)) + ((sk[46]) & (!g318) & (g408) & (g2307) & (g364) & (g453)) + ((sk[46]) & (g318) & (!g408) & (!g2307) & (!g364) & (g453)) + ((sk[46]) & (g318) & (!g408) & (!g2307) & (g364) & (!g453)) + ((sk[46]) & (g318) & (!g408) & (g2307) & (!g364) & (!g453)) + ((sk[46]) & (g318) & (!g408) & (g2307) & (g364) & (g453)) + ((sk[46]) & (g318) & (g408) & (!g2307) & (!g364) & (!g453)) + ((sk[46]) & (g318) & (g408) & (!g2307) & (g364) & (g453)) + ((sk[46]) & (g318) & (g408) & (g2307) & (!g364) & (!g453)) + ((sk[46]) & (g318) & (g408) & (g2307) & (g364) & (g453)));
	assign g2335 = (((!g1692) & (!g2033) & (!g2034) & (g2333) & (!sk[47]) & (!g2334)) + ((!g1692) & (!g2033) & (!g2034) & (g2333) & (!sk[47]) & (g2334)) + ((!g1692) & (!g2033) & (!g2034) & (g2333) & (sk[47]) & (!g2334)) + ((!g1692) & (!g2033) & (!g2034) & (g2333) & (sk[47]) & (g2334)) + ((!g1692) & (!g2033) & (g2034) & (!g2333) & (!sk[47]) & (!g2334)) + ((!g1692) & (!g2033) & (g2034) & (!g2333) & (!sk[47]) & (g2334)) + ((!g1692) & (!g2033) & (g2034) & (g2333) & (!sk[47]) & (!g2334)) + ((!g1692) & (!g2033) & (g2034) & (g2333) & (!sk[47]) & (g2334)) + ((!g1692) & (g2033) & (!g2034) & (!g2333) & (!sk[47]) & (!g2334)) + ((!g1692) & (g2033) & (!g2034) & (!g2333) & (!sk[47]) & (g2334)) + ((!g1692) & (g2033) & (!g2034) & (!g2333) & (sk[47]) & (g2334)) + ((!g1692) & (g2033) & (!g2034) & (g2333) & (!sk[47]) & (!g2334)) + ((!g1692) & (g2033) & (!g2034) & (g2333) & (!sk[47]) & (g2334)) + ((!g1692) & (g2033) & (!g2034) & (g2333) & (sk[47]) & (g2334)) + ((!g1692) & (g2033) & (g2034) & (!g2333) & (!sk[47]) & (!g2334)) + ((!g1692) & (g2033) & (g2034) & (!g2333) & (!sk[47]) & (g2334)) + ((!g1692) & (g2033) & (g2034) & (g2333) & (!sk[47]) & (!g2334)) + ((!g1692) & (g2033) & (g2034) & (g2333) & (!sk[47]) & (g2334)) + ((g1692) & (!g2033) & (!g2034) & (g2333) & (!sk[47]) & (!g2334)) + ((g1692) & (!g2033) & (!g2034) & (g2333) & (!sk[47]) & (g2334)) + ((g1692) & (!g2033) & (!g2034) & (g2333) & (sk[47]) & (!g2334)) + ((g1692) & (!g2033) & (!g2034) & (g2333) & (sk[47]) & (g2334)) + ((g1692) & (!g2033) & (g2034) & (!g2333) & (!sk[47]) & (!g2334)) + ((g1692) & (!g2033) & (g2034) & (!g2333) & (!sk[47]) & (g2334)) + ((g1692) & (!g2033) & (g2034) & (!g2333) & (sk[47]) & (!g2334)) + ((g1692) & (!g2033) & (g2034) & (!g2333) & (sk[47]) & (g2334)) + ((g1692) & (!g2033) & (g2034) & (g2333) & (!sk[47]) & (!g2334)) + ((g1692) & (!g2033) & (g2034) & (g2333) & (!sk[47]) & (g2334)) + ((g1692) & (!g2033) & (g2034) & (g2333) & (sk[47]) & (!g2334)) + ((g1692) & (!g2033) & (g2034) & (g2333) & (sk[47]) & (g2334)) + ((g1692) & (g2033) & (!g2034) & (!g2333) & (!sk[47]) & (!g2334)) + ((g1692) & (g2033) & (!g2034) & (!g2333) & (!sk[47]) & (g2334)) + ((g1692) & (g2033) & (!g2034) & (!g2333) & (sk[47]) & (g2334)) + ((g1692) & (g2033) & (!g2034) & (g2333) & (!sk[47]) & (!g2334)) + ((g1692) & (g2033) & (!g2034) & (g2333) & (!sk[47]) & (g2334)) + ((g1692) & (g2033) & (!g2034) & (g2333) & (sk[47]) & (g2334)) + ((g1692) & (g2033) & (g2034) & (!g2333) & (!sk[47]) & (!g2334)) + ((g1692) & (g2033) & (g2034) & (!g2333) & (!sk[47]) & (g2334)) + ((g1692) & (g2033) & (g2034) & (g2333) & (!sk[47]) & (!g2334)) + ((g1692) & (g2033) & (g2034) & (g2333) & (!sk[47]) & (g2334)));
	assign g2336 = (((!g2029) & (!g2332) & (!sk[48]) & (g2335)) + ((!g2029) & (!g2332) & (sk[48]) & (g2335)) + ((!g2029) & (g2332) & (!sk[48]) & (!g2335)) + ((!g2029) & (g2332) & (!sk[48]) & (g2335)) + ((!g2029) & (g2332) & (sk[48]) & (g2335)) + ((g2029) & (!g2332) & (!sk[48]) & (g2335)) + ((g2029) & (g2332) & (!sk[48]) & (!g2335)) + ((g2029) & (g2332) & (!sk[48]) & (g2335)) + ((g2029) & (g2332) & (sk[48]) & (!g2335)) + ((g2029) & (g2332) & (sk[48]) & (g2335)));
	assign g2337 = (((!g123) & (g2329) & (!intr_i) & (!g2330) & (!g2057) & (g2336)) + ((!g123) & (g2329) & (!intr_i) & (!g2330) & (g2057) & (g2336)) + ((!g123) & (g2329) & (!intr_i) & (g2330) & (!g2057) & (g2336)) + ((!g123) & (g2329) & (!intr_i) & (g2330) & (g2057) & (g2336)) + ((!g123) & (g2329) & (intr_i) & (!g2330) & (!g2057) & (g2336)) + ((!g123) & (g2329) & (intr_i) & (g2330) & (!g2057) & (g2336)) + ((!g123) & (g2329) & (intr_i) & (g2330) & (g2057) & (g2336)));
	assign g2338 = (((!dmem_dat_ix31x) & (!dmem_dat_ix23x) & (!dmem_dat_ix15x) & (dmem_dat_ix7x) & (g2128) & (g2129)) + ((!dmem_dat_ix31x) & (!dmem_dat_ix23x) & (dmem_dat_ix15x) & (!dmem_dat_ix7x) & (!g2128) & (g2129)) + ((!dmem_dat_ix31x) & (!dmem_dat_ix23x) & (dmem_dat_ix15x) & (dmem_dat_ix7x) & (!g2128) & (g2129)) + ((!dmem_dat_ix31x) & (!dmem_dat_ix23x) & (dmem_dat_ix15x) & (dmem_dat_ix7x) & (g2128) & (g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix23x) & (!dmem_dat_ix15x) & (!dmem_dat_ix7x) & (g2128) & (!g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix23x) & (!dmem_dat_ix15x) & (dmem_dat_ix7x) & (g2128) & (!g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix23x) & (!dmem_dat_ix15x) & (dmem_dat_ix7x) & (g2128) & (g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix23x) & (dmem_dat_ix15x) & (!dmem_dat_ix7x) & (!g2128) & (g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix23x) & (dmem_dat_ix15x) & (!dmem_dat_ix7x) & (g2128) & (!g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix23x) & (dmem_dat_ix15x) & (dmem_dat_ix7x) & (!g2128) & (g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix23x) & (dmem_dat_ix15x) & (dmem_dat_ix7x) & (g2128) & (!g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix23x) & (dmem_dat_ix15x) & (dmem_dat_ix7x) & (g2128) & (g2129)) + ((dmem_dat_ix31x) & (!dmem_dat_ix23x) & (!dmem_dat_ix15x) & (!dmem_dat_ix7x) & (!g2128) & (!g2129)) + ((dmem_dat_ix31x) & (!dmem_dat_ix23x) & (!dmem_dat_ix15x) & (dmem_dat_ix7x) & (!g2128) & (!g2129)) + ((dmem_dat_ix31x) & (!dmem_dat_ix23x) & (!dmem_dat_ix15x) & (dmem_dat_ix7x) & (g2128) & (g2129)) + ((dmem_dat_ix31x) & (!dmem_dat_ix23x) & (dmem_dat_ix15x) & (!dmem_dat_ix7x) & (!g2128) & (!g2129)) + ((dmem_dat_ix31x) & (!dmem_dat_ix23x) & (dmem_dat_ix15x) & (!dmem_dat_ix7x) & (!g2128) & (g2129)) + ((dmem_dat_ix31x) & (!dmem_dat_ix23x) & (dmem_dat_ix15x) & (dmem_dat_ix7x) & (!g2128) & (!g2129)) + ((dmem_dat_ix31x) & (!dmem_dat_ix23x) & (dmem_dat_ix15x) & (dmem_dat_ix7x) & (!g2128) & (g2129)) + ((dmem_dat_ix31x) & (!dmem_dat_ix23x) & (dmem_dat_ix15x) & (dmem_dat_ix7x) & (g2128) & (g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix23x) & (!dmem_dat_ix15x) & (!dmem_dat_ix7x) & (!g2128) & (!g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix23x) & (!dmem_dat_ix15x) & (!dmem_dat_ix7x) & (g2128) & (!g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix23x) & (!dmem_dat_ix15x) & (dmem_dat_ix7x) & (!g2128) & (!g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix23x) & (!dmem_dat_ix15x) & (dmem_dat_ix7x) & (g2128) & (!g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix23x) & (!dmem_dat_ix15x) & (dmem_dat_ix7x) & (g2128) & (g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix23x) & (dmem_dat_ix15x) & (!dmem_dat_ix7x) & (!g2128) & (!g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix23x) & (dmem_dat_ix15x) & (!dmem_dat_ix7x) & (!g2128) & (g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix23x) & (dmem_dat_ix15x) & (!dmem_dat_ix7x) & (g2128) & (!g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix23x) & (dmem_dat_ix15x) & (dmem_dat_ix7x) & (!g2128) & (!g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix23x) & (dmem_dat_ix15x) & (dmem_dat_ix7x) & (!g2128) & (g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix23x) & (dmem_dat_ix15x) & (dmem_dat_ix7x) & (g2128) & (!g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix23x) & (dmem_dat_ix15x) & (dmem_dat_ix7x) & (g2128) & (g2129)));
	assign g2339 = (((g2131) & (g2132) & (!dmem_dat_ix7x) & (dmem_dat_ix23x) & (!g2128) & (!g2129)) + ((g2131) & (g2132) & (dmem_dat_ix7x) & (!dmem_dat_ix23x) & (!g2128) & (g2129)) + ((g2131) & (g2132) & (dmem_dat_ix7x) & (dmem_dat_ix23x) & (!g2128) & (!g2129)) + ((g2131) & (g2132) & (dmem_dat_ix7x) & (dmem_dat_ix23x) & (!g2128) & (g2129)));
	assign g2341 = (((!g2115) & (!g2116) & (!g2312) & (!g2314) & (!g2295) & (g2340)) + ((!g2115) & (!g2116) & (!g2312) & (!g2314) & (g2295) & (g2340)) + ((!g2115) & (!g2116) & (!g2312) & (g2314) & (!g2295) & (g2340)) + ((!g2115) & (!g2116) & (!g2312) & (g2314) & (g2295) & (g2340)) + ((!g2115) & (!g2116) & (g2312) & (!g2314) & (!g2295) & (g2340)) + ((!g2115) & (!g2116) & (g2312) & (!g2314) & (g2295) & (!g2340)) + ((!g2115) & (!g2116) & (g2312) & (g2314) & (!g2295) & (!g2340)) + ((!g2115) & (!g2116) & (g2312) & (g2314) & (g2295) & (!g2340)) + ((!g2115) & (g2116) & (!g2312) & (!g2314) & (!g2295) & (!g2340)) + ((!g2115) & (g2116) & (!g2312) & (!g2314) & (g2295) & (!g2340)) + ((!g2115) & (g2116) & (!g2312) & (g2314) & (!g2295) & (!g2340)) + ((!g2115) & (g2116) & (!g2312) & (g2314) & (g2295) & (!g2340)) + ((!g2115) & (g2116) & (g2312) & (!g2314) & (!g2295) & (!g2340)) + ((!g2115) & (g2116) & (g2312) & (!g2314) & (g2295) & (g2340)) + ((!g2115) & (g2116) & (g2312) & (g2314) & (!g2295) & (g2340)) + ((!g2115) & (g2116) & (g2312) & (g2314) & (g2295) & (g2340)) + ((g2115) & (!g2116) & (!g2312) & (!g2314) & (!g2295) & (g2340)) + ((g2115) & (!g2116) & (!g2312) & (!g2314) & (g2295) & (!g2340)) + ((g2115) & (!g2116) & (!g2312) & (g2314) & (!g2295) & (!g2340)) + ((g2115) & (!g2116) & (!g2312) & (g2314) & (g2295) & (!g2340)) + ((g2115) & (!g2116) & (g2312) & (!g2314) & (!g2295) & (!g2340)) + ((g2115) & (!g2116) & (g2312) & (!g2314) & (g2295) & (!g2340)) + ((g2115) & (!g2116) & (g2312) & (g2314) & (!g2295) & (!g2340)) + ((g2115) & (!g2116) & (g2312) & (g2314) & (g2295) & (!g2340)) + ((g2115) & (g2116) & (!g2312) & (!g2314) & (!g2295) & (!g2340)) + ((g2115) & (g2116) & (!g2312) & (!g2314) & (g2295) & (g2340)) + ((g2115) & (g2116) & (!g2312) & (g2314) & (!g2295) & (g2340)) + ((g2115) & (g2116) & (!g2312) & (g2314) & (g2295) & (g2340)) + ((g2115) & (g2116) & (g2312) & (!g2314) & (!g2295) & (g2340)) + ((g2115) & (g2116) & (g2312) & (!g2314) & (g2295) & (g2340)) + ((g2115) & (g2116) & (g2312) & (g2314) & (!g2295) & (g2340)) + ((g2115) & (g2116) & (g2312) & (g2314) & (g2295) & (g2340)));
	assign g2342 = (((!g2266) & (!sk[53]) & (!g2267) & (!g2290) & (g2315)) + ((!g2266) & (!sk[53]) & (!g2267) & (g2290) & (!g2315)) + ((!g2266) & (!sk[53]) & (!g2267) & (g2290) & (g2315)) + ((!g2266) & (!sk[53]) & (g2267) & (!g2290) & (!g2315)) + ((!g2266) & (!sk[53]) & (g2267) & (!g2290) & (g2315)) + ((!g2266) & (!sk[53]) & (g2267) & (g2290) & (!g2315)) + ((!g2266) & (!sk[53]) & (g2267) & (g2290) & (g2315)) + ((g2266) & (!sk[53]) & (!g2267) & (!g2290) & (g2315)) + ((g2266) & (!sk[53]) & (!g2267) & (g2290) & (!g2315)) + ((g2266) & (!sk[53]) & (!g2267) & (g2290) & (g2315)) + ((g2266) & (!sk[53]) & (g2267) & (!g2290) & (!g2315)) + ((g2266) & (!sk[53]) & (g2267) & (!g2290) & (g2315)) + ((g2266) & (!sk[53]) & (g2267) & (g2290) & (!g2315)) + ((g2266) & (!sk[53]) & (g2267) & (g2290) & (g2315)) + ((g2266) & (sk[53]) & (g2267) & (g2290) & (g2315)));
	assign g2343 = (((!g2289) & (!g2114) & (!sk[54]) & (!g2115) & (g2312)) + ((!g2289) & (!g2114) & (!sk[54]) & (g2115) & (!g2312)) + ((!g2289) & (!g2114) & (!sk[54]) & (g2115) & (g2312)) + ((!g2289) & (!g2114) & (sk[54]) & (!g2115) & (!g2312)) + ((!g2289) & (!g2114) & (sk[54]) & (g2115) & (g2312)) + ((!g2289) & (g2114) & (!sk[54]) & (!g2115) & (!g2312)) + ((!g2289) & (g2114) & (!sk[54]) & (!g2115) & (g2312)) + ((!g2289) & (g2114) & (!sk[54]) & (g2115) & (!g2312)) + ((!g2289) & (g2114) & (!sk[54]) & (g2115) & (g2312)) + ((!g2289) & (g2114) & (sk[54]) & (!g2115) & (g2312)) + ((!g2289) & (g2114) & (sk[54]) & (g2115) & (!g2312)) + ((g2289) & (!g2114) & (!sk[54]) & (!g2115) & (g2312)) + ((g2289) & (!g2114) & (!sk[54]) & (g2115) & (!g2312)) + ((g2289) & (!g2114) & (!sk[54]) & (g2115) & (g2312)) + ((g2289) & (!g2114) & (sk[54]) & (!g2115) & (!g2312)) + ((g2289) & (!g2114) & (sk[54]) & (g2115) & (g2312)) + ((g2289) & (g2114) & (!sk[54]) & (!g2115) & (!g2312)) + ((g2289) & (g2114) & (!sk[54]) & (!g2115) & (g2312)) + ((g2289) & (g2114) & (!sk[54]) & (g2115) & (!g2312)) + ((g2289) & (g2114) & (!sk[54]) & (g2115) & (g2312)) + ((g2289) & (g2114) & (sk[54]) & (!g2115) & (!g2312)) + ((g2289) & (g2114) & (sk[54]) & (g2115) & (g2312)));
	assign g2344 = (((!g2268) & (!g2269) & (!g2270) & (g2292) & (g2293) & (g2343)) + ((!g2268) & (!g2269) & (g2270) & (g2292) & (g2293) & (g2343)) + ((!g2268) & (g2269) & (!g2270) & (g2292) & (g2293) & (g2343)) + ((!g2268) & (g2269) & (g2270) & (!g2292) & (g2293) & (g2343)) + ((!g2268) & (g2269) & (g2270) & (g2292) & (!g2293) & (g2343)) + ((!g2268) & (g2269) & (g2270) & (g2292) & (g2293) & (g2343)) + ((g2268) & (!g2269) & (!g2270) & (g2292) & (g2293) & (g2343)) + ((g2268) & (!g2269) & (g2270) & (!g2292) & (g2293) & (g2343)) + ((g2268) & (!g2269) & (g2270) & (g2292) & (!g2293) & (g2343)) + ((g2268) & (!g2269) & (g2270) & (g2292) & (g2293) & (g2343)) + ((g2268) & (g2269) & (!g2270) & (!g2292) & (g2293) & (g2343)) + ((g2268) & (g2269) & (!g2270) & (g2292) & (!g2293) & (g2343)) + ((g2268) & (g2269) & (!g2270) & (g2292) & (g2293) & (g2343)) + ((g2268) & (g2269) & (g2270) & (!g2292) & (g2293) & (g2343)) + ((g2268) & (g2269) & (g2270) & (g2292) & (!g2293) & (g2343)) + ((g2268) & (g2269) & (g2270) & (g2292) & (g2293) & (g2343)));
	assign g2345 = (((!sk[56]) & (g2317) & (!g2318)) + ((!sk[56]) & (g2317) & (g2318)) + ((sk[56]) & (g2317) & (g2318)));
	assign g2346 = (((!sk[57]) & (g2344) & (!g2345)) + ((!sk[57]) & (g2344) & (g2345)) + ((sk[57]) & (!g2344) & (!g2345)));
	assign g2347 = (((!sk[58]) & (g2115) & (!g2312)) + ((!sk[58]) & (g2115) & (g2312)) + ((sk[58]) & (g2115) & (!g2312)));
	assign g2348 = (((!g2116) & (sk[59]) & (!g2340)) + ((g2116) & (!sk[59]) & (!g2340)) + ((g2116) & (!sk[59]) & (g2340)) + ((g2116) & (sk[59]) & (g2340)));
	assign g2349 = (((!g2346) & (!g2347) & (!sk[60]) & (g2348)) + ((!g2346) & (!g2347) & (sk[60]) & (!g2348)) + ((!g2346) & (g2347) & (!sk[60]) & (!g2348)) + ((!g2346) & (g2347) & (!sk[60]) & (g2348)) + ((!g2346) & (g2347) & (sk[60]) & (g2348)) + ((g2346) & (!g2347) & (!sk[60]) & (g2348)) + ((g2346) & (!g2347) & (sk[60]) & (g2348)) + ((g2346) & (g2347) & (!sk[60]) & (!g2348)) + ((g2346) & (g2347) & (!sk[60]) & (g2348)) + ((g2346) & (g2347) & (sk[60]) & (!g2348)));
	assign g2350 = (((!g2116) & (!g2115) & (!g2114) & (g2113) & (g2071) & (g2074)) + ((!g2116) & (!g2115) & (g2114) & (!g2113) & (!g2071) & (g2074)) + ((!g2116) & (!g2115) & (g2114) & (g2113) & (!g2071) & (g2074)) + ((!g2116) & (!g2115) & (g2114) & (g2113) & (g2071) & (g2074)) + ((!g2116) & (g2115) & (!g2114) & (!g2113) & (g2071) & (!g2074)) + ((!g2116) & (g2115) & (!g2114) & (g2113) & (g2071) & (!g2074)) + ((!g2116) & (g2115) & (!g2114) & (g2113) & (g2071) & (g2074)) + ((!g2116) & (g2115) & (g2114) & (!g2113) & (!g2071) & (g2074)) + ((!g2116) & (g2115) & (g2114) & (!g2113) & (g2071) & (!g2074)) + ((!g2116) & (g2115) & (g2114) & (g2113) & (!g2071) & (g2074)) + ((!g2116) & (g2115) & (g2114) & (g2113) & (g2071) & (!g2074)) + ((!g2116) & (g2115) & (g2114) & (g2113) & (g2071) & (g2074)) + ((g2116) & (!g2115) & (!g2114) & (!g2113) & (!g2071) & (!g2074)) + ((g2116) & (!g2115) & (!g2114) & (g2113) & (!g2071) & (!g2074)) + ((g2116) & (!g2115) & (!g2114) & (g2113) & (g2071) & (g2074)) + ((g2116) & (!g2115) & (g2114) & (!g2113) & (!g2071) & (!g2074)) + ((g2116) & (!g2115) & (g2114) & (!g2113) & (!g2071) & (g2074)) + ((g2116) & (!g2115) & (g2114) & (g2113) & (!g2071) & (!g2074)) + ((g2116) & (!g2115) & (g2114) & (g2113) & (!g2071) & (g2074)) + ((g2116) & (!g2115) & (g2114) & (g2113) & (g2071) & (g2074)) + ((g2116) & (g2115) & (!g2114) & (!g2113) & (!g2071) & (!g2074)) + ((g2116) & (g2115) & (!g2114) & (!g2113) & (g2071) & (!g2074)) + ((g2116) & (g2115) & (!g2114) & (g2113) & (!g2071) & (!g2074)) + ((g2116) & (g2115) & (!g2114) & (g2113) & (g2071) & (!g2074)) + ((g2116) & (g2115) & (!g2114) & (g2113) & (g2071) & (g2074)) + ((g2116) & (g2115) & (g2114) & (!g2113) & (!g2071) & (!g2074)) + ((g2116) & (g2115) & (g2114) & (!g2113) & (!g2071) & (g2074)) + ((g2116) & (g2115) & (g2114) & (!g2113) & (g2071) & (!g2074)) + ((g2116) & (g2115) & (g2114) & (g2113) & (!g2071) & (!g2074)) + ((g2116) & (g2115) & (g2114) & (g2113) & (!g2071) & (g2074)) + ((g2116) & (g2115) & (g2114) & (g2113) & (g2071) & (!g2074)) + ((g2116) & (g2115) & (g2114) & (g2113) & (g2071) & (g2074)));
	assign g2351 = (((!g2076) & (!g2077) & (!sk[62]) & (!g2236) & (g2350)) + ((!g2076) & (!g2077) & (!sk[62]) & (g2236) & (!g2350)) + ((!g2076) & (!g2077) & (!sk[62]) & (g2236) & (g2350)) + ((!g2076) & (!g2077) & (sk[62]) & (!g2236) & (g2350)) + ((!g2076) & (!g2077) & (sk[62]) & (g2236) & (g2350)) + ((!g2076) & (g2077) & (!sk[62]) & (!g2236) & (!g2350)) + ((!g2076) & (g2077) & (!sk[62]) & (!g2236) & (g2350)) + ((!g2076) & (g2077) & (!sk[62]) & (g2236) & (!g2350)) + ((!g2076) & (g2077) & (!sk[62]) & (g2236) & (g2350)) + ((!g2076) & (g2077) & (sk[62]) & (g2236) & (!g2350)) + ((!g2076) & (g2077) & (sk[62]) & (g2236) & (g2350)) + ((g2076) & (!g2077) & (!sk[62]) & (!g2236) & (g2350)) + ((g2076) & (!g2077) & (!sk[62]) & (g2236) & (!g2350)) + ((g2076) & (!g2077) & (!sk[62]) & (g2236) & (g2350)) + ((g2076) & (g2077) & (!sk[62]) & (!g2236) & (!g2350)) + ((g2076) & (g2077) & (!sk[62]) & (!g2236) & (g2350)) + ((g2076) & (g2077) & (!sk[62]) & (g2236) & (!g2350)) + ((g2076) & (g2077) & (!sk[62]) & (g2236) & (g2350)));
	assign g2352 = (((!g2247) & (!g2250) & (!g2249) & (g2242) & (g2076) & (g2077)) + ((!g2247) & (!g2250) & (g2249) & (!g2242) & (!g2076) & (g2077)) + ((!g2247) & (!g2250) & (g2249) & (g2242) & (!g2076) & (g2077)) + ((!g2247) & (!g2250) & (g2249) & (g2242) & (g2076) & (g2077)) + ((!g2247) & (g2250) & (!g2249) & (!g2242) & (g2076) & (!g2077)) + ((!g2247) & (g2250) & (!g2249) & (g2242) & (g2076) & (!g2077)) + ((!g2247) & (g2250) & (!g2249) & (g2242) & (g2076) & (g2077)) + ((!g2247) & (g2250) & (g2249) & (!g2242) & (!g2076) & (g2077)) + ((!g2247) & (g2250) & (g2249) & (!g2242) & (g2076) & (!g2077)) + ((!g2247) & (g2250) & (g2249) & (g2242) & (!g2076) & (g2077)) + ((!g2247) & (g2250) & (g2249) & (g2242) & (g2076) & (!g2077)) + ((!g2247) & (g2250) & (g2249) & (g2242) & (g2076) & (g2077)) + ((g2247) & (!g2250) & (!g2249) & (!g2242) & (!g2076) & (!g2077)) + ((g2247) & (!g2250) & (!g2249) & (g2242) & (!g2076) & (!g2077)) + ((g2247) & (!g2250) & (!g2249) & (g2242) & (g2076) & (g2077)) + ((g2247) & (!g2250) & (g2249) & (!g2242) & (!g2076) & (!g2077)) + ((g2247) & (!g2250) & (g2249) & (!g2242) & (!g2076) & (g2077)) + ((g2247) & (!g2250) & (g2249) & (g2242) & (!g2076) & (!g2077)) + ((g2247) & (!g2250) & (g2249) & (g2242) & (!g2076) & (g2077)) + ((g2247) & (!g2250) & (g2249) & (g2242) & (g2076) & (g2077)) + ((g2247) & (g2250) & (!g2249) & (!g2242) & (!g2076) & (!g2077)) + ((g2247) & (g2250) & (!g2249) & (!g2242) & (g2076) & (!g2077)) + ((g2247) & (g2250) & (!g2249) & (g2242) & (!g2076) & (!g2077)) + ((g2247) & (g2250) & (!g2249) & (g2242) & (g2076) & (!g2077)) + ((g2247) & (g2250) & (!g2249) & (g2242) & (g2076) & (g2077)) + ((g2247) & (g2250) & (g2249) & (!g2242) & (!g2076) & (!g2077)) + ((g2247) & (g2250) & (g2249) & (!g2242) & (!g2076) & (g2077)) + ((g2247) & (g2250) & (g2249) & (!g2242) & (g2076) & (!g2077)) + ((g2247) & (g2250) & (g2249) & (g2242) & (!g2076) & (!g2077)) + ((g2247) & (g2250) & (g2249) & (g2242) & (!g2076) & (g2077)) + ((g2247) & (g2250) & (g2249) & (g2242) & (g2076) & (!g2077)) + ((g2247) & (g2250) & (g2249) & (g2242) & (g2076) & (g2077)));
	assign g2353 = (((!g2244) & (!g2245) & (!g2243) & (g2192) & (g2076) & (g2077)) + ((!g2244) & (!g2245) & (g2243) & (!g2192) & (!g2076) & (g2077)) + ((!g2244) & (!g2245) & (g2243) & (g2192) & (!g2076) & (g2077)) + ((!g2244) & (!g2245) & (g2243) & (g2192) & (g2076) & (g2077)) + ((!g2244) & (g2245) & (!g2243) & (!g2192) & (g2076) & (!g2077)) + ((!g2244) & (g2245) & (!g2243) & (g2192) & (g2076) & (!g2077)) + ((!g2244) & (g2245) & (!g2243) & (g2192) & (g2076) & (g2077)) + ((!g2244) & (g2245) & (g2243) & (!g2192) & (!g2076) & (g2077)) + ((!g2244) & (g2245) & (g2243) & (!g2192) & (g2076) & (!g2077)) + ((!g2244) & (g2245) & (g2243) & (g2192) & (!g2076) & (g2077)) + ((!g2244) & (g2245) & (g2243) & (g2192) & (g2076) & (!g2077)) + ((!g2244) & (g2245) & (g2243) & (g2192) & (g2076) & (g2077)) + ((g2244) & (!g2245) & (!g2243) & (!g2192) & (!g2076) & (!g2077)) + ((g2244) & (!g2245) & (!g2243) & (g2192) & (!g2076) & (!g2077)) + ((g2244) & (!g2245) & (!g2243) & (g2192) & (g2076) & (g2077)) + ((g2244) & (!g2245) & (g2243) & (!g2192) & (!g2076) & (!g2077)) + ((g2244) & (!g2245) & (g2243) & (!g2192) & (!g2076) & (g2077)) + ((g2244) & (!g2245) & (g2243) & (g2192) & (!g2076) & (!g2077)) + ((g2244) & (!g2245) & (g2243) & (g2192) & (!g2076) & (g2077)) + ((g2244) & (!g2245) & (g2243) & (g2192) & (g2076) & (g2077)) + ((g2244) & (g2245) & (!g2243) & (!g2192) & (!g2076) & (!g2077)) + ((g2244) & (g2245) & (!g2243) & (!g2192) & (g2076) & (!g2077)) + ((g2244) & (g2245) & (!g2243) & (g2192) & (!g2076) & (!g2077)) + ((g2244) & (g2245) & (!g2243) & (g2192) & (g2076) & (!g2077)) + ((g2244) & (g2245) & (!g2243) & (g2192) & (g2076) & (g2077)) + ((g2244) & (g2245) & (g2243) & (!g2192) & (!g2076) & (!g2077)) + ((g2244) & (g2245) & (g2243) & (!g2192) & (!g2076) & (g2077)) + ((g2244) & (g2245) & (g2243) & (!g2192) & (g2076) & (!g2077)) + ((g2244) & (g2245) & (g2243) & (g2192) & (!g2076) & (!g2077)) + ((g2244) & (g2245) & (g2243) & (g2192) & (!g2076) & (g2077)) + ((g2244) & (g2245) & (g2243) & (g2192) & (g2076) & (!g2077)) + ((g2244) & (g2245) & (g2243) & (g2192) & (g2076) & (g2077)));
	assign g2354 = (((!g2073) & (!g2080) & (!g2125) & (g2351) & (!g2352) & (!g2353)) + ((!g2073) & (!g2080) & (!g2125) & (g2351) & (!g2352) & (g2353)) + ((!g2073) & (!g2080) & (!g2125) & (g2351) & (g2352) & (!g2353)) + ((!g2073) & (!g2080) & (!g2125) & (g2351) & (g2352) & (g2353)) + ((!g2073) & (!g2080) & (g2125) & (!g2351) & (g2352) & (!g2353)) + ((!g2073) & (!g2080) & (g2125) & (!g2351) & (g2352) & (g2353)) + ((!g2073) & (!g2080) & (g2125) & (g2351) & (g2352) & (!g2353)) + ((!g2073) & (!g2080) & (g2125) & (g2351) & (g2352) & (g2353)) + ((!g2073) & (g2080) & (!g2125) & (g2351) & (!g2352) & (!g2353)) + ((!g2073) & (g2080) & (!g2125) & (g2351) & (!g2352) & (g2353)) + ((!g2073) & (g2080) & (!g2125) & (g2351) & (g2352) & (!g2353)) + ((!g2073) & (g2080) & (!g2125) & (g2351) & (g2352) & (g2353)) + ((!g2073) & (g2080) & (g2125) & (!g2351) & (g2352) & (!g2353)) + ((!g2073) & (g2080) & (g2125) & (!g2351) & (g2352) & (g2353)) + ((!g2073) & (g2080) & (g2125) & (g2351) & (g2352) & (!g2353)) + ((!g2073) & (g2080) & (g2125) & (g2351) & (g2352) & (g2353)) + ((g2073) & (!g2080) & (g2125) & (!g2351) & (!g2352) & (g2353)) + ((g2073) & (!g2080) & (g2125) & (!g2351) & (g2352) & (g2353)) + ((g2073) & (!g2080) & (g2125) & (g2351) & (!g2352) & (g2353)) + ((g2073) & (!g2080) & (g2125) & (g2351) & (g2352) & (g2353)) + ((g2073) & (g2080) & (!g2125) & (g2351) & (!g2352) & (!g2353)) + ((g2073) & (g2080) & (!g2125) & (g2351) & (!g2352) & (g2353)) + ((g2073) & (g2080) & (!g2125) & (g2351) & (g2352) & (!g2353)) + ((g2073) & (g2080) & (!g2125) & (g2351) & (g2352) & (g2353)) + ((g2073) & (g2080) & (g2125) & (!g2351) & (!g2352) & (g2353)) + ((g2073) & (g2080) & (g2125) & (!g2351) & (g2352) & (g2353)) + ((g2073) & (g2080) & (g2125) & (g2351) & (!g2352) & (g2353)) + ((g2073) & (g2080) & (g2125) & (g2351) & (g2352) & (g2353)));
	assign g2355 = (((!sk[66]) & (!g496) & (!g453) & (g2331)) + ((!sk[66]) & (!g496) & (g453) & (!g2331)) + ((!sk[66]) & (!g496) & (g453) & (g2331)) + ((!sk[66]) & (g496) & (!g453) & (g2331)) + ((!sk[66]) & (g496) & (g453) & (!g2331)) + ((!sk[66]) & (g496) & (g453) & (g2331)) + ((sk[66]) & (!g496) & (!g453) & (!g2331)) + ((sk[66]) & (!g496) & (!g453) & (g2331)) + ((sk[66]) & (!g496) & (g453) & (!g2331)) + ((sk[66]) & (g496) & (g453) & (g2331)));
	assign g2356 = (((!nmi_i) & (!sk[67]) & (!g2023) & (!intr_i) & (g2039) & (!g2056)) + ((!nmi_i) & (!sk[67]) & (!g2023) & (!intr_i) & (g2039) & (g2056)) + ((!nmi_i) & (!sk[67]) & (!g2023) & (intr_i) & (!g2039) & (!g2056)) + ((!nmi_i) & (!sk[67]) & (!g2023) & (intr_i) & (!g2039) & (g2056)) + ((!nmi_i) & (!sk[67]) & (!g2023) & (intr_i) & (g2039) & (!g2056)) + ((!nmi_i) & (!sk[67]) & (!g2023) & (intr_i) & (g2039) & (g2056)) + ((!nmi_i) & (!sk[67]) & (g2023) & (!intr_i) & (!g2039) & (!g2056)) + ((!nmi_i) & (!sk[67]) & (g2023) & (!intr_i) & (!g2039) & (g2056)) + ((!nmi_i) & (!sk[67]) & (g2023) & (!intr_i) & (g2039) & (!g2056)) + ((!nmi_i) & (!sk[67]) & (g2023) & (!intr_i) & (g2039) & (g2056)) + ((!nmi_i) & (!sk[67]) & (g2023) & (intr_i) & (!g2039) & (!g2056)) + ((!nmi_i) & (!sk[67]) & (g2023) & (intr_i) & (!g2039) & (g2056)) + ((!nmi_i) & (!sk[67]) & (g2023) & (intr_i) & (g2039) & (!g2056)) + ((!nmi_i) & (!sk[67]) & (g2023) & (intr_i) & (g2039) & (g2056)) + ((!nmi_i) & (sk[67]) & (!g2023) & (!intr_i) & (!g2039) & (!g2056)) + ((!nmi_i) & (sk[67]) & (!g2023) & (!intr_i) & (!g2039) & (g2056)) + ((!nmi_i) & (sk[67]) & (!g2023) & (!intr_i) & (g2039) & (!g2056)) + ((!nmi_i) & (sk[67]) & (!g2023) & (!intr_i) & (g2039) & (g2056)) + ((!nmi_i) & (sk[67]) & (!g2023) & (intr_i) & (!g2039) & (!g2056)) + ((nmi_i) & (!sk[67]) & (!g2023) & (!intr_i) & (g2039) & (!g2056)) + ((nmi_i) & (!sk[67]) & (!g2023) & (!intr_i) & (g2039) & (g2056)) + ((nmi_i) & (!sk[67]) & (!g2023) & (intr_i) & (!g2039) & (!g2056)) + ((nmi_i) & (!sk[67]) & (!g2023) & (intr_i) & (!g2039) & (g2056)) + ((nmi_i) & (!sk[67]) & (!g2023) & (intr_i) & (g2039) & (!g2056)) + ((nmi_i) & (!sk[67]) & (!g2023) & (intr_i) & (g2039) & (g2056)) + ((nmi_i) & (!sk[67]) & (g2023) & (!intr_i) & (!g2039) & (!g2056)) + ((nmi_i) & (!sk[67]) & (g2023) & (!intr_i) & (!g2039) & (g2056)) + ((nmi_i) & (!sk[67]) & (g2023) & (!intr_i) & (g2039) & (!g2056)) + ((nmi_i) & (!sk[67]) & (g2023) & (!intr_i) & (g2039) & (g2056)) + ((nmi_i) & (!sk[67]) & (g2023) & (intr_i) & (!g2039) & (!g2056)) + ((nmi_i) & (!sk[67]) & (g2023) & (intr_i) & (!g2039) & (g2056)) + ((nmi_i) & (!sk[67]) & (g2023) & (intr_i) & (g2039) & (!g2056)) + ((nmi_i) & (!sk[67]) & (g2023) & (intr_i) & (g2039) & (g2056)));
	assign g5032 = (((!sk[68]) & (!g2921) & (!g3068) & (g2357)) + ((!sk[68]) & (!g2921) & (g3068) & (!g2357)) + ((!sk[68]) & (!g2921) & (g3068) & (g2357)) + ((!sk[68]) & (g2921) & (!g3068) & (g2357)) + ((!sk[68]) & (g2921) & (g3068) & (!g2357)) + ((!sk[68]) & (g2921) & (g3068) & (g2357)) + ((sk[68]) & (!g2921) & (!g3068) & (g2357)) + ((sk[68]) & (!g2921) & (g3068) & (g2357)) + ((sk[68]) & (g2921) & (g3068) & (!g2357)) + ((sk[68]) & (g2921) & (g3068) & (g2357)));
	assign g2358 = (((!g364) & (!g453) & (!g318) & (!sk[69]) & (g408) & (!g2307)) + ((!g364) & (!g453) & (!g318) & (!sk[69]) & (g408) & (g2307)) + ((!g364) & (!g453) & (g318) & (!sk[69]) & (!g408) & (!g2307)) + ((!g364) & (!g453) & (g318) & (!sk[69]) & (!g408) & (g2307)) + ((!g364) & (!g453) & (g318) & (!sk[69]) & (g408) & (!g2307)) + ((!g364) & (!g453) & (g318) & (!sk[69]) & (g408) & (g2307)) + ((!g364) & (g453) & (!g318) & (!sk[69]) & (!g408) & (!g2307)) + ((!g364) & (g453) & (!g318) & (!sk[69]) & (!g408) & (g2307)) + ((!g364) & (g453) & (!g318) & (!sk[69]) & (g408) & (!g2307)) + ((!g364) & (g453) & (!g318) & (!sk[69]) & (g408) & (g2307)) + ((!g364) & (g453) & (!g318) & (sk[69]) & (g408) & (g2307)) + ((!g364) & (g453) & (g318) & (!sk[69]) & (!g408) & (!g2307)) + ((!g364) & (g453) & (g318) & (!sk[69]) & (!g408) & (g2307)) + ((!g364) & (g453) & (g318) & (!sk[69]) & (g408) & (!g2307)) + ((!g364) & (g453) & (g318) & (!sk[69]) & (g408) & (g2307)) + ((!g364) & (g453) & (g318) & (sk[69]) & (!g408) & (g2307)) + ((!g364) & (g453) & (g318) & (sk[69]) & (g408) & (!g2307)) + ((!g364) & (g453) & (g318) & (sk[69]) & (g408) & (g2307)) + ((g364) & (!g453) & (!g318) & (!sk[69]) & (g408) & (!g2307)) + ((g364) & (!g453) & (!g318) & (!sk[69]) & (g408) & (g2307)) + ((g364) & (!g453) & (!g318) & (sk[69]) & (g408) & (g2307)) + ((g364) & (!g453) & (g318) & (!sk[69]) & (!g408) & (!g2307)) + ((g364) & (!g453) & (g318) & (!sk[69]) & (!g408) & (g2307)) + ((g364) & (!g453) & (g318) & (!sk[69]) & (g408) & (!g2307)) + ((g364) & (!g453) & (g318) & (!sk[69]) & (g408) & (g2307)) + ((g364) & (!g453) & (g318) & (sk[69]) & (!g408) & (g2307)) + ((g364) & (!g453) & (g318) & (sk[69]) & (g408) & (!g2307)) + ((g364) & (!g453) & (g318) & (sk[69]) & (g408) & (g2307)) + ((g364) & (g453) & (!g318) & (!sk[69]) & (!g408) & (!g2307)) + ((g364) & (g453) & (!g318) & (!sk[69]) & (!g408) & (g2307)) + ((g364) & (g453) & (!g318) & (!sk[69]) & (g408) & (!g2307)) + ((g364) & (g453) & (!g318) & (!sk[69]) & (g408) & (g2307)) + ((g364) & (g453) & (!g318) & (sk[69]) & (!g408) & (!g2307)) + ((g364) & (g453) & (!g318) & (sk[69]) & (!g408) & (g2307)) + ((g364) & (g453) & (!g318) & (sk[69]) & (g408) & (!g2307)) + ((g364) & (g453) & (!g318) & (sk[69]) & (g408) & (g2307)) + ((g364) & (g453) & (g318) & (!sk[69]) & (!g408) & (!g2307)) + ((g364) & (g453) & (g318) & (!sk[69]) & (!g408) & (g2307)) + ((g364) & (g453) & (g318) & (!sk[69]) & (g408) & (!g2307)) + ((g364) & (g453) & (g318) & (!sk[69]) & (g408) & (g2307)) + ((g364) & (g453) & (g318) & (sk[69]) & (!g408) & (!g2307)) + ((g364) & (g453) & (g318) & (sk[69]) & (!g408) & (g2307)) + ((g364) & (g453) & (g318) & (sk[69]) & (g408) & (!g2307)) + ((g364) & (g453) & (g318) & (sk[69]) & (g408) & (g2307)));
	assign g2359 = (((!g86) & (!g496) & (!sk[70]) & (g2358)) + ((!g86) & (!g496) & (sk[70]) & (!g2358)) + ((!g86) & (g496) & (!sk[70]) & (!g2358)) + ((!g86) & (g496) & (!sk[70]) & (g2358)) + ((!g86) & (g496) & (sk[70]) & (g2358)) + ((g86) & (!g496) & (!sk[70]) & (g2358)) + ((g86) & (!g496) & (sk[70]) & (g2358)) + ((g86) & (g496) & (!sk[70]) & (!g2358)) + ((g86) & (g496) & (!sk[70]) & (g2358)) + ((g86) & (g496) & (sk[70]) & (!g2358)));
	assign g2360 = (((!g1705) & (!g2033) & (!g2034) & (g2357) & (!sk[71]) & (!g2359)) + ((!g1705) & (!g2033) & (!g2034) & (g2357) & (!sk[71]) & (g2359)) + ((!g1705) & (!g2033) & (!g2034) & (g2357) & (sk[71]) & (!g2359)) + ((!g1705) & (!g2033) & (!g2034) & (g2357) & (sk[71]) & (g2359)) + ((!g1705) & (!g2033) & (g2034) & (!g2357) & (!sk[71]) & (!g2359)) + ((!g1705) & (!g2033) & (g2034) & (!g2357) & (!sk[71]) & (g2359)) + ((!g1705) & (!g2033) & (g2034) & (g2357) & (!sk[71]) & (!g2359)) + ((!g1705) & (!g2033) & (g2034) & (g2357) & (!sk[71]) & (g2359)) + ((!g1705) & (g2033) & (!g2034) & (!g2357) & (!sk[71]) & (!g2359)) + ((!g1705) & (g2033) & (!g2034) & (!g2357) & (!sk[71]) & (g2359)) + ((!g1705) & (g2033) & (!g2034) & (!g2357) & (sk[71]) & (g2359)) + ((!g1705) & (g2033) & (!g2034) & (g2357) & (!sk[71]) & (!g2359)) + ((!g1705) & (g2033) & (!g2034) & (g2357) & (!sk[71]) & (g2359)) + ((!g1705) & (g2033) & (!g2034) & (g2357) & (sk[71]) & (g2359)) + ((!g1705) & (g2033) & (g2034) & (!g2357) & (!sk[71]) & (!g2359)) + ((!g1705) & (g2033) & (g2034) & (!g2357) & (!sk[71]) & (g2359)) + ((!g1705) & (g2033) & (g2034) & (g2357) & (!sk[71]) & (!g2359)) + ((!g1705) & (g2033) & (g2034) & (g2357) & (!sk[71]) & (g2359)) + ((g1705) & (!g2033) & (!g2034) & (g2357) & (!sk[71]) & (!g2359)) + ((g1705) & (!g2033) & (!g2034) & (g2357) & (!sk[71]) & (g2359)) + ((g1705) & (!g2033) & (!g2034) & (g2357) & (sk[71]) & (!g2359)) + ((g1705) & (!g2033) & (!g2034) & (g2357) & (sk[71]) & (g2359)) + ((g1705) & (!g2033) & (g2034) & (!g2357) & (!sk[71]) & (!g2359)) + ((g1705) & (!g2033) & (g2034) & (!g2357) & (!sk[71]) & (g2359)) + ((g1705) & (!g2033) & (g2034) & (!g2357) & (sk[71]) & (!g2359)) + ((g1705) & (!g2033) & (g2034) & (!g2357) & (sk[71]) & (g2359)) + ((g1705) & (!g2033) & (g2034) & (g2357) & (!sk[71]) & (!g2359)) + ((g1705) & (!g2033) & (g2034) & (g2357) & (!sk[71]) & (g2359)) + ((g1705) & (!g2033) & (g2034) & (g2357) & (sk[71]) & (!g2359)) + ((g1705) & (!g2033) & (g2034) & (g2357) & (sk[71]) & (g2359)) + ((g1705) & (g2033) & (!g2034) & (!g2357) & (!sk[71]) & (!g2359)) + ((g1705) & (g2033) & (!g2034) & (!g2357) & (!sk[71]) & (g2359)) + ((g1705) & (g2033) & (!g2034) & (!g2357) & (sk[71]) & (g2359)) + ((g1705) & (g2033) & (!g2034) & (g2357) & (!sk[71]) & (!g2359)) + ((g1705) & (g2033) & (!g2034) & (g2357) & (!sk[71]) & (g2359)) + ((g1705) & (g2033) & (!g2034) & (g2357) & (sk[71]) & (g2359)) + ((g1705) & (g2033) & (g2034) & (!g2357) & (!sk[71]) & (!g2359)) + ((g1705) & (g2033) & (g2034) & (!g2357) & (!sk[71]) & (g2359)) + ((g1705) & (g2033) & (g2034) & (g2357) & (!sk[71]) & (!g2359)) + ((g1705) & (g2033) & (g2034) & (g2357) & (!sk[71]) & (g2359)));
	assign g2361 = (((!g2022) & (!g123) & (!g2028) & (!g2355) & (!g2356) & (g2360)) + ((!g2022) & (!g123) & (!g2028) & (!g2355) & (g2356) & (g2360)) + ((!g2022) & (!g123) & (!g2028) & (g2355) & (!g2356) & (g2360)) + ((!g2022) & (!g123) & (!g2028) & (g2355) & (g2356) & (g2360)) + ((!g2022) & (!g123) & (g2028) & (!g2355) & (!g2356) & (g2360)) + ((!g2022) & (!g123) & (g2028) & (!g2355) & (g2356) & (g2360)) + ((!g2022) & (!g123) & (g2028) & (g2355) & (!g2356) & (g2360)) + ((!g2022) & (!g123) & (g2028) & (g2355) & (g2356) & (g2360)) + ((g2022) & (!g123) & (!g2028) & (!g2355) & (!g2356) & (!g2360)) + ((g2022) & (!g123) & (!g2028) & (!g2355) & (!g2356) & (g2360)) + ((g2022) & (!g123) & (!g2028) & (g2355) & (!g2356) & (!g2360)) + ((g2022) & (!g123) & (!g2028) & (g2355) & (!g2356) & (g2360)) + ((g2022) & (!g123) & (!g2028) & (g2355) & (g2356) & (!g2360)) + ((g2022) & (!g123) & (!g2028) & (g2355) & (g2356) & (g2360)) + ((g2022) & (!g123) & (g2028) & (!g2355) & (!g2356) & (!g2360)) + ((g2022) & (!g123) & (g2028) & (!g2355) & (!g2356) & (g2360)) + ((g2022) & (!g123) & (g2028) & (!g2355) & (g2356) & (g2360)) + ((g2022) & (!g123) & (g2028) & (g2355) & (!g2356) & (!g2360)) + ((g2022) & (!g123) & (g2028) & (g2355) & (!g2356) & (g2360)) + ((g2022) & (!g123) & (g2028) & (g2355) & (g2356) & (g2360)));
	assign g2362 = (((g2131) & (g2132) & (!dmem_dat_ix24x) & (dmem_dat_ix8x) & (!g2128) & (g2129)) + ((g2131) & (g2132) & (dmem_dat_ix24x) & (!dmem_dat_ix8x) & (!g2128) & (!g2129)) + ((g2131) & (g2132) & (dmem_dat_ix24x) & (dmem_dat_ix8x) & (!g2128) & (!g2129)) + ((g2131) & (g2132) & (dmem_dat_ix24x) & (dmem_dat_ix8x) & (!g2128) & (g2129)));
	assign g2363 = (((g78) & (!g79) & (g80) & (!g81) & (!g82) & (!g83)));
	assign g2364 = (((!g2363) & (!g2131) & (!sk[75]) & (!g2132) & (dmem_dat_ix8x) & (!g2338)) + ((!g2363) & (!g2131) & (!sk[75]) & (!g2132) & (dmem_dat_ix8x) & (g2338)) + ((!g2363) & (!g2131) & (!sk[75]) & (g2132) & (!dmem_dat_ix8x) & (!g2338)) + ((!g2363) & (!g2131) & (!sk[75]) & (g2132) & (!dmem_dat_ix8x) & (g2338)) + ((!g2363) & (!g2131) & (!sk[75]) & (g2132) & (dmem_dat_ix8x) & (!g2338)) + ((!g2363) & (!g2131) & (!sk[75]) & (g2132) & (dmem_dat_ix8x) & (g2338)) + ((!g2363) & (g2131) & (!sk[75]) & (!g2132) & (!dmem_dat_ix8x) & (!g2338)) + ((!g2363) & (g2131) & (!sk[75]) & (!g2132) & (!dmem_dat_ix8x) & (g2338)) + ((!g2363) & (g2131) & (!sk[75]) & (!g2132) & (dmem_dat_ix8x) & (!g2338)) + ((!g2363) & (g2131) & (!sk[75]) & (!g2132) & (dmem_dat_ix8x) & (g2338)) + ((!g2363) & (g2131) & (!sk[75]) & (g2132) & (!dmem_dat_ix8x) & (!g2338)) + ((!g2363) & (g2131) & (!sk[75]) & (g2132) & (!dmem_dat_ix8x) & (g2338)) + ((!g2363) & (g2131) & (!sk[75]) & (g2132) & (dmem_dat_ix8x) & (!g2338)) + ((!g2363) & (g2131) & (!sk[75]) & (g2132) & (dmem_dat_ix8x) & (g2338)) + ((!g2363) & (g2131) & (sk[75]) & (!g2132) & (dmem_dat_ix8x) & (!g2338)) + ((!g2363) & (g2131) & (sk[75]) & (!g2132) & (dmem_dat_ix8x) & (g2338)) + ((g2363) & (!g2131) & (!sk[75]) & (!g2132) & (dmem_dat_ix8x) & (!g2338)) + ((g2363) & (!g2131) & (!sk[75]) & (!g2132) & (dmem_dat_ix8x) & (g2338)) + ((g2363) & (!g2131) & (!sk[75]) & (g2132) & (!dmem_dat_ix8x) & (!g2338)) + ((g2363) & (!g2131) & (!sk[75]) & (g2132) & (!dmem_dat_ix8x) & (g2338)) + ((g2363) & (!g2131) & (!sk[75]) & (g2132) & (dmem_dat_ix8x) & (!g2338)) + ((g2363) & (!g2131) & (!sk[75]) & (g2132) & (dmem_dat_ix8x) & (g2338)) + ((g2363) & (!g2131) & (sk[75]) & (!g2132) & (!dmem_dat_ix8x) & (g2338)) + ((g2363) & (!g2131) & (sk[75]) & (!g2132) & (dmem_dat_ix8x) & (g2338)) + ((g2363) & (!g2131) & (sk[75]) & (g2132) & (!dmem_dat_ix8x) & (g2338)) + ((g2363) & (!g2131) & (sk[75]) & (g2132) & (dmem_dat_ix8x) & (g2338)) + ((g2363) & (g2131) & (!sk[75]) & (!g2132) & (!dmem_dat_ix8x) & (!g2338)) + ((g2363) & (g2131) & (!sk[75]) & (!g2132) & (!dmem_dat_ix8x) & (g2338)) + ((g2363) & (g2131) & (!sk[75]) & (!g2132) & (dmem_dat_ix8x) & (!g2338)) + ((g2363) & (g2131) & (!sk[75]) & (!g2132) & (dmem_dat_ix8x) & (g2338)) + ((g2363) & (g2131) & (!sk[75]) & (g2132) & (!dmem_dat_ix8x) & (!g2338)) + ((g2363) & (g2131) & (!sk[75]) & (g2132) & (!dmem_dat_ix8x) & (g2338)) + ((g2363) & (g2131) & (!sk[75]) & (g2132) & (dmem_dat_ix8x) & (!g2338)) + ((g2363) & (g2131) & (!sk[75]) & (g2132) & (dmem_dat_ix8x) & (g2338)) + ((g2363) & (g2131) & (sk[75]) & (!g2132) & (dmem_dat_ix8x) & (!g2338)) + ((g2363) & (g2131) & (sk[75]) & (!g2132) & (dmem_dat_ix8x) & (g2338)));
	assign g2366 = (((!g2115) & (!g2116) & (g2312) & (!g2314) & (g2295) & (g2340)) + ((!g2115) & (!g2116) & (g2312) & (g2314) & (!g2295) & (g2340)) + ((!g2115) & (!g2116) & (g2312) & (g2314) & (g2295) & (g2340)) + ((!g2115) & (g2116) & (!g2312) & (!g2314) & (!g2295) & (g2340)) + ((!g2115) & (g2116) & (!g2312) & (!g2314) & (g2295) & (g2340)) + ((!g2115) & (g2116) & (!g2312) & (g2314) & (!g2295) & (g2340)) + ((!g2115) & (g2116) & (!g2312) & (g2314) & (g2295) & (g2340)) + ((!g2115) & (g2116) & (g2312) & (!g2314) & (!g2295) & (g2340)) + ((!g2115) & (g2116) & (g2312) & (!g2314) & (g2295) & (!g2340)) + ((!g2115) & (g2116) & (g2312) & (!g2314) & (g2295) & (g2340)) + ((!g2115) & (g2116) & (g2312) & (g2314) & (!g2295) & (!g2340)) + ((!g2115) & (g2116) & (g2312) & (g2314) & (!g2295) & (g2340)) + ((!g2115) & (g2116) & (g2312) & (g2314) & (g2295) & (!g2340)) + ((!g2115) & (g2116) & (g2312) & (g2314) & (g2295) & (g2340)) + ((g2115) & (!g2116) & (!g2312) & (!g2314) & (g2295) & (g2340)) + ((g2115) & (!g2116) & (!g2312) & (g2314) & (!g2295) & (g2340)) + ((g2115) & (!g2116) & (!g2312) & (g2314) & (g2295) & (g2340)) + ((g2115) & (!g2116) & (g2312) & (!g2314) & (!g2295) & (g2340)) + ((g2115) & (!g2116) & (g2312) & (!g2314) & (g2295) & (g2340)) + ((g2115) & (!g2116) & (g2312) & (g2314) & (!g2295) & (g2340)) + ((g2115) & (!g2116) & (g2312) & (g2314) & (g2295) & (g2340)) + ((g2115) & (g2116) & (!g2312) & (!g2314) & (!g2295) & (g2340)) + ((g2115) & (g2116) & (!g2312) & (!g2314) & (g2295) & (!g2340)) + ((g2115) & (g2116) & (!g2312) & (!g2314) & (g2295) & (g2340)) + ((g2115) & (g2116) & (!g2312) & (g2314) & (!g2295) & (!g2340)) + ((g2115) & (g2116) & (!g2312) & (g2314) & (!g2295) & (g2340)) + ((g2115) & (g2116) & (!g2312) & (g2314) & (g2295) & (!g2340)) + ((g2115) & (g2116) & (!g2312) & (g2314) & (g2295) & (g2340)) + ((g2115) & (g2116) & (g2312) & (!g2314) & (!g2295) & (!g2340)) + ((g2115) & (g2116) & (g2312) & (!g2314) & (!g2295) & (g2340)) + ((g2115) & (g2116) & (g2312) & (!g2314) & (g2295) & (!g2340)) + ((g2115) & (g2116) & (g2312) & (!g2314) & (g2295) & (g2340)) + ((g2115) & (g2116) & (g2312) & (g2314) & (!g2295) & (!g2340)) + ((g2115) & (g2116) & (g2312) & (g2314) & (!g2295) & (g2340)) + ((g2115) & (g2116) & (g2312) & (g2314) & (g2295) & (!g2340)) + ((g2115) & (g2116) & (g2312) & (g2314) & (g2295) & (g2340)));
	assign g2367 = (((!sk[77]) & (!g2108) & (!g2365) & (g2366)) + ((!sk[77]) & (!g2108) & (g2365) & (!g2366)) + ((!sk[77]) & (!g2108) & (g2365) & (g2366)) + ((!sk[77]) & (g2108) & (!g2365) & (g2366)) + ((!sk[77]) & (g2108) & (g2365) & (!g2366)) + ((!sk[77]) & (g2108) & (g2365) & (g2366)) + ((sk[77]) & (!g2108) & (!g2365) & (g2366)) + ((sk[77]) & (!g2108) & (g2365) & (!g2366)) + ((sk[77]) & (g2108) & (!g2365) & (!g2366)) + ((sk[77]) & (g2108) & (g2365) & (g2366)));
	assign g2368 = (((!g2341) & (!sk[78]) & (!g2342) & (g2367)) + ((!g2341) & (!sk[78]) & (g2342) & (!g2367)) + ((!g2341) & (!sk[78]) & (g2342) & (g2367)) + ((!g2341) & (sk[78]) & (!g2342) & (g2367)) + ((!g2341) & (sk[78]) & (g2342) & (g2367)) + ((g2341) & (!sk[78]) & (!g2342) & (g2367)) + ((g2341) & (!sk[78]) & (g2342) & (!g2367)) + ((g2341) & (!sk[78]) & (g2342) & (g2367)) + ((g2341) & (sk[78]) & (!g2342) & (g2367)) + ((g2341) & (sk[78]) & (g2342) & (!g2367)));
	assign g2369 = (((g2116) & (!sk[79]) & (!g2340)) + ((g2116) & (!sk[79]) & (g2340)) + ((g2116) & (sk[79]) & (!g2340)));
	assign g2370 = (((!g2108) & (sk[80]) & (!g2365)) + ((g2108) & (!sk[80]) & (!g2365)) + ((g2108) & (!sk[80]) & (g2365)) + ((g2108) & (sk[80]) & (g2365)));
	assign g2371 = (((!g2346) & (!sk[81]) & (!g2347) & (!g2348) & (g2369) & (!g2370)) + ((!g2346) & (!sk[81]) & (!g2347) & (!g2348) & (g2369) & (g2370)) + ((!g2346) & (!sk[81]) & (!g2347) & (g2348) & (!g2369) & (!g2370)) + ((!g2346) & (!sk[81]) & (!g2347) & (g2348) & (!g2369) & (g2370)) + ((!g2346) & (!sk[81]) & (!g2347) & (g2348) & (g2369) & (!g2370)) + ((!g2346) & (!sk[81]) & (!g2347) & (g2348) & (g2369) & (g2370)) + ((!g2346) & (!sk[81]) & (g2347) & (!g2348) & (!g2369) & (!g2370)) + ((!g2346) & (!sk[81]) & (g2347) & (!g2348) & (!g2369) & (g2370)) + ((!g2346) & (!sk[81]) & (g2347) & (!g2348) & (g2369) & (!g2370)) + ((!g2346) & (!sk[81]) & (g2347) & (!g2348) & (g2369) & (g2370)) + ((!g2346) & (!sk[81]) & (g2347) & (g2348) & (!g2369) & (!g2370)) + ((!g2346) & (!sk[81]) & (g2347) & (g2348) & (!g2369) & (g2370)) + ((!g2346) & (!sk[81]) & (g2347) & (g2348) & (g2369) & (!g2370)) + ((!g2346) & (!sk[81]) & (g2347) & (g2348) & (g2369) & (g2370)) + ((!g2346) & (sk[81]) & (!g2347) & (!g2348) & (!g2369) & (g2370)) + ((!g2346) & (sk[81]) & (!g2347) & (!g2348) & (g2369) & (!g2370)) + ((!g2346) & (sk[81]) & (!g2347) & (g2348) & (!g2369) & (!g2370)) + ((!g2346) & (sk[81]) & (!g2347) & (g2348) & (g2369) & (g2370)) + ((!g2346) & (sk[81]) & (g2347) & (!g2348) & (!g2369) & (!g2370)) + ((!g2346) & (sk[81]) & (g2347) & (!g2348) & (g2369) & (g2370)) + ((!g2346) & (sk[81]) & (g2347) & (g2348) & (!g2369) & (!g2370)) + ((!g2346) & (sk[81]) & (g2347) & (g2348) & (g2369) & (g2370)) + ((g2346) & (!sk[81]) & (!g2347) & (!g2348) & (g2369) & (!g2370)) + ((g2346) & (!sk[81]) & (!g2347) & (!g2348) & (g2369) & (g2370)) + ((g2346) & (!sk[81]) & (!g2347) & (g2348) & (!g2369) & (!g2370)) + ((g2346) & (!sk[81]) & (!g2347) & (g2348) & (!g2369) & (g2370)) + ((g2346) & (!sk[81]) & (!g2347) & (g2348) & (g2369) & (!g2370)) + ((g2346) & (!sk[81]) & (!g2347) & (g2348) & (g2369) & (g2370)) + ((g2346) & (!sk[81]) & (g2347) & (!g2348) & (!g2369) & (!g2370)) + ((g2346) & (!sk[81]) & (g2347) & (!g2348) & (!g2369) & (g2370)) + ((g2346) & (!sk[81]) & (g2347) & (!g2348) & (g2369) & (!g2370)) + ((g2346) & (!sk[81]) & (g2347) & (!g2348) & (g2369) & (g2370)) + ((g2346) & (!sk[81]) & (g2347) & (g2348) & (!g2369) & (!g2370)) + ((g2346) & (!sk[81]) & (g2347) & (g2348) & (!g2369) & (g2370)) + ((g2346) & (!sk[81]) & (g2347) & (g2348) & (g2369) & (!g2370)) + ((g2346) & (!sk[81]) & (g2347) & (g2348) & (g2369) & (g2370)) + ((g2346) & (sk[81]) & (!g2347) & (!g2348) & (!g2369) & (g2370)) + ((g2346) & (sk[81]) & (!g2347) & (!g2348) & (g2369) & (!g2370)) + ((g2346) & (sk[81]) & (!g2347) & (g2348) & (!g2369) & (g2370)) + ((g2346) & (sk[81]) & (!g2347) & (g2348) & (g2369) & (!g2370)) + ((g2346) & (sk[81]) & (g2347) & (!g2348) & (!g2369) & (g2370)) + ((g2346) & (sk[81]) & (g2347) & (!g2348) & (g2369) & (!g2370)) + ((g2346) & (sk[81]) & (g2347) & (g2348) & (!g2369) & (!g2370)) + ((g2346) & (sk[81]) & (g2347) & (g2348) & (g2369) & (g2370)));
	assign g2372 = (((!g2108) & (!g2116) & (!g2115) & (g2114) & (g2071) & (g2074)) + ((!g2108) & (!g2116) & (g2115) & (!g2114) & (!g2071) & (g2074)) + ((!g2108) & (!g2116) & (g2115) & (g2114) & (!g2071) & (g2074)) + ((!g2108) & (!g2116) & (g2115) & (g2114) & (g2071) & (g2074)) + ((!g2108) & (g2116) & (!g2115) & (!g2114) & (g2071) & (!g2074)) + ((!g2108) & (g2116) & (!g2115) & (g2114) & (g2071) & (!g2074)) + ((!g2108) & (g2116) & (!g2115) & (g2114) & (g2071) & (g2074)) + ((!g2108) & (g2116) & (g2115) & (!g2114) & (!g2071) & (g2074)) + ((!g2108) & (g2116) & (g2115) & (!g2114) & (g2071) & (!g2074)) + ((!g2108) & (g2116) & (g2115) & (g2114) & (!g2071) & (g2074)) + ((!g2108) & (g2116) & (g2115) & (g2114) & (g2071) & (!g2074)) + ((!g2108) & (g2116) & (g2115) & (g2114) & (g2071) & (g2074)) + ((g2108) & (!g2116) & (!g2115) & (!g2114) & (!g2071) & (!g2074)) + ((g2108) & (!g2116) & (!g2115) & (g2114) & (!g2071) & (!g2074)) + ((g2108) & (!g2116) & (!g2115) & (g2114) & (g2071) & (g2074)) + ((g2108) & (!g2116) & (g2115) & (!g2114) & (!g2071) & (!g2074)) + ((g2108) & (!g2116) & (g2115) & (!g2114) & (!g2071) & (g2074)) + ((g2108) & (!g2116) & (g2115) & (g2114) & (!g2071) & (!g2074)) + ((g2108) & (!g2116) & (g2115) & (g2114) & (!g2071) & (g2074)) + ((g2108) & (!g2116) & (g2115) & (g2114) & (g2071) & (g2074)) + ((g2108) & (g2116) & (!g2115) & (!g2114) & (!g2071) & (!g2074)) + ((g2108) & (g2116) & (!g2115) & (!g2114) & (g2071) & (!g2074)) + ((g2108) & (g2116) & (!g2115) & (g2114) & (!g2071) & (!g2074)) + ((g2108) & (g2116) & (!g2115) & (g2114) & (g2071) & (!g2074)) + ((g2108) & (g2116) & (!g2115) & (g2114) & (g2071) & (g2074)) + ((g2108) & (g2116) & (g2115) & (!g2114) & (!g2071) & (!g2074)) + ((g2108) & (g2116) & (g2115) & (!g2114) & (!g2071) & (g2074)) + ((g2108) & (g2116) & (g2115) & (!g2114) & (g2071) & (!g2074)) + ((g2108) & (g2116) & (g2115) & (g2114) & (!g2071) & (!g2074)) + ((g2108) & (g2116) & (g2115) & (g2114) & (!g2071) & (g2074)) + ((g2108) & (g2116) & (g2115) & (g2114) & (g2071) & (!g2074)) + ((g2108) & (g2116) & (g2115) & (g2114) & (g2071) & (g2074)));
	assign g2373 = (((!sk[83]) & (!g2075) & (!g2076) & (!g2077) & (g2272) & (!g2372)) + ((!sk[83]) & (!g2075) & (!g2076) & (!g2077) & (g2272) & (g2372)) + ((!sk[83]) & (!g2075) & (!g2076) & (g2077) & (!g2272) & (!g2372)) + ((!sk[83]) & (!g2075) & (!g2076) & (g2077) & (!g2272) & (g2372)) + ((!sk[83]) & (!g2075) & (!g2076) & (g2077) & (g2272) & (!g2372)) + ((!sk[83]) & (!g2075) & (!g2076) & (g2077) & (g2272) & (g2372)) + ((!sk[83]) & (!g2075) & (g2076) & (!g2077) & (!g2272) & (!g2372)) + ((!sk[83]) & (!g2075) & (g2076) & (!g2077) & (!g2272) & (g2372)) + ((!sk[83]) & (!g2075) & (g2076) & (!g2077) & (g2272) & (!g2372)) + ((!sk[83]) & (!g2075) & (g2076) & (!g2077) & (g2272) & (g2372)) + ((!sk[83]) & (!g2075) & (g2076) & (g2077) & (!g2272) & (!g2372)) + ((!sk[83]) & (!g2075) & (g2076) & (g2077) & (!g2272) & (g2372)) + ((!sk[83]) & (!g2075) & (g2076) & (g2077) & (g2272) & (!g2372)) + ((!sk[83]) & (!g2075) & (g2076) & (g2077) & (g2272) & (g2372)) + ((!sk[83]) & (g2075) & (!g2076) & (!g2077) & (g2272) & (!g2372)) + ((!sk[83]) & (g2075) & (!g2076) & (!g2077) & (g2272) & (g2372)) + ((!sk[83]) & (g2075) & (!g2076) & (g2077) & (!g2272) & (!g2372)) + ((!sk[83]) & (g2075) & (!g2076) & (g2077) & (!g2272) & (g2372)) + ((!sk[83]) & (g2075) & (!g2076) & (g2077) & (g2272) & (!g2372)) + ((!sk[83]) & (g2075) & (!g2076) & (g2077) & (g2272) & (g2372)) + ((!sk[83]) & (g2075) & (g2076) & (!g2077) & (!g2272) & (!g2372)) + ((!sk[83]) & (g2075) & (g2076) & (!g2077) & (!g2272) & (g2372)) + ((!sk[83]) & (g2075) & (g2076) & (!g2077) & (g2272) & (!g2372)) + ((!sk[83]) & (g2075) & (g2076) & (!g2077) & (g2272) & (g2372)) + ((!sk[83]) & (g2075) & (g2076) & (g2077) & (!g2272) & (!g2372)) + ((!sk[83]) & (g2075) & (g2076) & (g2077) & (!g2272) & (g2372)) + ((!sk[83]) & (g2075) & (g2076) & (g2077) & (g2272) & (!g2372)) + ((!sk[83]) & (g2075) & (g2076) & (g2077) & (g2272) & (g2372)) + ((sk[83]) & (!g2075) & (!g2076) & (!g2077) & (!g2272) & (g2372)) + ((sk[83]) & (!g2075) & (!g2076) & (!g2077) & (g2272) & (g2372)) + ((sk[83]) & (!g2075) & (!g2076) & (g2077) & (g2272) & (!g2372)) + ((sk[83]) & (!g2075) & (!g2076) & (g2077) & (g2272) & (g2372)) + ((sk[83]) & (g2075) & (!g2076) & (!g2077) & (!g2272) & (g2372)) + ((sk[83]) & (g2075) & (!g2076) & (!g2077) & (g2272) & (g2372)) + ((sk[83]) & (g2075) & (!g2076) & (g2077) & (g2272) & (!g2372)) + ((sk[83]) & (g2075) & (!g2076) & (g2077) & (g2272) & (g2372)) + ((sk[83]) & (g2075) & (g2076) & (!g2077) & (!g2272) & (!g2372)) + ((sk[83]) & (g2075) & (g2076) & (!g2077) & (!g2272) & (g2372)) + ((sk[83]) & (g2075) & (g2076) & (!g2077) & (g2272) & (!g2372)) + ((sk[83]) & (g2075) & (g2076) & (!g2077) & (g2272) & (g2372)));
	assign g2374 = (((!sk[84]) & (!g2076) & (!g2077) & (!g2092) & (g2102) & (!g2192)) + ((!sk[84]) & (!g2076) & (!g2077) & (!g2092) & (g2102) & (g2192)) + ((!sk[84]) & (!g2076) & (!g2077) & (g2092) & (!g2102) & (!g2192)) + ((!sk[84]) & (!g2076) & (!g2077) & (g2092) & (!g2102) & (g2192)) + ((!sk[84]) & (!g2076) & (!g2077) & (g2092) & (g2102) & (!g2192)) + ((!sk[84]) & (!g2076) & (!g2077) & (g2092) & (g2102) & (g2192)) + ((!sk[84]) & (!g2076) & (g2077) & (!g2092) & (!g2102) & (!g2192)) + ((!sk[84]) & (!g2076) & (g2077) & (!g2092) & (!g2102) & (g2192)) + ((!sk[84]) & (!g2076) & (g2077) & (!g2092) & (g2102) & (!g2192)) + ((!sk[84]) & (!g2076) & (g2077) & (!g2092) & (g2102) & (g2192)) + ((!sk[84]) & (!g2076) & (g2077) & (g2092) & (!g2102) & (!g2192)) + ((!sk[84]) & (!g2076) & (g2077) & (g2092) & (!g2102) & (g2192)) + ((!sk[84]) & (!g2076) & (g2077) & (g2092) & (g2102) & (!g2192)) + ((!sk[84]) & (!g2076) & (g2077) & (g2092) & (g2102) & (g2192)) + ((!sk[84]) & (g2076) & (!g2077) & (!g2092) & (g2102) & (!g2192)) + ((!sk[84]) & (g2076) & (!g2077) & (!g2092) & (g2102) & (g2192)) + ((!sk[84]) & (g2076) & (!g2077) & (g2092) & (!g2102) & (!g2192)) + ((!sk[84]) & (g2076) & (!g2077) & (g2092) & (!g2102) & (g2192)) + ((!sk[84]) & (g2076) & (!g2077) & (g2092) & (g2102) & (!g2192)) + ((!sk[84]) & (g2076) & (!g2077) & (g2092) & (g2102) & (g2192)) + ((!sk[84]) & (g2076) & (g2077) & (!g2092) & (!g2102) & (!g2192)) + ((!sk[84]) & (g2076) & (g2077) & (!g2092) & (!g2102) & (g2192)) + ((!sk[84]) & (g2076) & (g2077) & (!g2092) & (g2102) & (!g2192)) + ((!sk[84]) & (g2076) & (g2077) & (!g2092) & (g2102) & (g2192)) + ((!sk[84]) & (g2076) & (g2077) & (g2092) & (!g2102) & (!g2192)) + ((!sk[84]) & (g2076) & (g2077) & (g2092) & (!g2102) & (g2192)) + ((!sk[84]) & (g2076) & (g2077) & (g2092) & (g2102) & (!g2192)) + ((!sk[84]) & (g2076) & (g2077) & (g2092) & (g2102) & (g2192)) + ((sk[84]) & (!g2076) & (!g2077) & (g2092) & (!g2102) & (!g2192)) + ((sk[84]) & (!g2076) & (!g2077) & (g2092) & (!g2102) & (g2192)) + ((sk[84]) & (!g2076) & (!g2077) & (g2092) & (g2102) & (!g2192)) + ((sk[84]) & (!g2076) & (!g2077) & (g2092) & (g2102) & (g2192)) + ((sk[84]) & (!g2076) & (g2077) & (!g2092) & (g2102) & (!g2192)) + ((sk[84]) & (!g2076) & (g2077) & (!g2092) & (g2102) & (g2192)) + ((sk[84]) & (!g2076) & (g2077) & (g2092) & (g2102) & (!g2192)) + ((sk[84]) & (!g2076) & (g2077) & (g2092) & (g2102) & (g2192)) + ((sk[84]) & (g2076) & (!g2077) & (!g2092) & (!g2102) & (g2192)) + ((sk[84]) & (g2076) & (!g2077) & (!g2092) & (g2102) & (g2192)) + ((sk[84]) & (g2076) & (!g2077) & (g2092) & (!g2102) & (g2192)) + ((sk[84]) & (g2076) & (!g2077) & (g2092) & (g2102) & (g2192)) + ((sk[84]) & (g2076) & (g2077) & (!g2092) & (!g2102) & (g2192)) + ((sk[84]) & (g2076) & (g2077) & (!g2092) & (g2102) & (g2192)) + ((sk[84]) & (g2076) & (g2077) & (g2092) & (!g2102) & (g2192)) + ((sk[84]) & (g2076) & (g2077) & (g2092) & (g2102) & (g2192)));
	assign g2375 = (((!g2112) & (!g2087) & (!g2122) & (g2097) & (g2076) & (g2077)) + ((!g2112) & (!g2087) & (g2122) & (!g2097) & (!g2076) & (g2077)) + ((!g2112) & (!g2087) & (g2122) & (g2097) & (!g2076) & (g2077)) + ((!g2112) & (!g2087) & (g2122) & (g2097) & (g2076) & (g2077)) + ((!g2112) & (g2087) & (!g2122) & (!g2097) & (g2076) & (!g2077)) + ((!g2112) & (g2087) & (!g2122) & (g2097) & (g2076) & (!g2077)) + ((!g2112) & (g2087) & (!g2122) & (g2097) & (g2076) & (g2077)) + ((!g2112) & (g2087) & (g2122) & (!g2097) & (!g2076) & (g2077)) + ((!g2112) & (g2087) & (g2122) & (!g2097) & (g2076) & (!g2077)) + ((!g2112) & (g2087) & (g2122) & (g2097) & (!g2076) & (g2077)) + ((!g2112) & (g2087) & (g2122) & (g2097) & (g2076) & (!g2077)) + ((!g2112) & (g2087) & (g2122) & (g2097) & (g2076) & (g2077)) + ((g2112) & (!g2087) & (!g2122) & (!g2097) & (!g2076) & (!g2077)) + ((g2112) & (!g2087) & (!g2122) & (g2097) & (!g2076) & (!g2077)) + ((g2112) & (!g2087) & (!g2122) & (g2097) & (g2076) & (g2077)) + ((g2112) & (!g2087) & (g2122) & (!g2097) & (!g2076) & (!g2077)) + ((g2112) & (!g2087) & (g2122) & (!g2097) & (!g2076) & (g2077)) + ((g2112) & (!g2087) & (g2122) & (g2097) & (!g2076) & (!g2077)) + ((g2112) & (!g2087) & (g2122) & (g2097) & (!g2076) & (g2077)) + ((g2112) & (!g2087) & (g2122) & (g2097) & (g2076) & (g2077)) + ((g2112) & (g2087) & (!g2122) & (!g2097) & (!g2076) & (!g2077)) + ((g2112) & (g2087) & (!g2122) & (!g2097) & (g2076) & (!g2077)) + ((g2112) & (g2087) & (!g2122) & (g2097) & (!g2076) & (!g2077)) + ((g2112) & (g2087) & (!g2122) & (g2097) & (g2076) & (!g2077)) + ((g2112) & (g2087) & (!g2122) & (g2097) & (g2076) & (g2077)) + ((g2112) & (g2087) & (g2122) & (!g2097) & (!g2076) & (!g2077)) + ((g2112) & (g2087) & (g2122) & (!g2097) & (!g2076) & (g2077)) + ((g2112) & (g2087) & (g2122) & (!g2097) & (g2076) & (!g2077)) + ((g2112) & (g2087) & (g2122) & (g2097) & (!g2076) & (!g2077)) + ((g2112) & (g2087) & (g2122) & (g2097) & (!g2076) & (g2077)) + ((g2112) & (g2087) & (g2122) & (g2097) & (g2076) & (!g2077)) + ((g2112) & (g2087) & (g2122) & (g2097) & (g2076) & (g2077)));
	assign g2376 = (((!g2073) & (!g2080) & (!g2125) & (g2373) & (!g2374) & (!g2375)) + ((!g2073) & (!g2080) & (!g2125) & (g2373) & (!g2374) & (g2375)) + ((!g2073) & (!g2080) & (!g2125) & (g2373) & (g2374) & (!g2375)) + ((!g2073) & (!g2080) & (!g2125) & (g2373) & (g2374) & (g2375)) + ((!g2073) & (!g2080) & (g2125) & (!g2373) & (!g2374) & (g2375)) + ((!g2073) & (!g2080) & (g2125) & (!g2373) & (g2374) & (g2375)) + ((!g2073) & (!g2080) & (g2125) & (g2373) & (!g2374) & (g2375)) + ((!g2073) & (!g2080) & (g2125) & (g2373) & (g2374) & (g2375)) + ((!g2073) & (g2080) & (!g2125) & (g2373) & (!g2374) & (!g2375)) + ((!g2073) & (g2080) & (!g2125) & (g2373) & (!g2374) & (g2375)) + ((!g2073) & (g2080) & (!g2125) & (g2373) & (g2374) & (!g2375)) + ((!g2073) & (g2080) & (!g2125) & (g2373) & (g2374) & (g2375)) + ((!g2073) & (g2080) & (g2125) & (!g2373) & (!g2374) & (g2375)) + ((!g2073) & (g2080) & (g2125) & (!g2373) & (g2374) & (g2375)) + ((!g2073) & (g2080) & (g2125) & (g2373) & (!g2374) & (g2375)) + ((!g2073) & (g2080) & (g2125) & (g2373) & (g2374) & (g2375)) + ((g2073) & (!g2080) & (g2125) & (!g2373) & (g2374) & (!g2375)) + ((g2073) & (!g2080) & (g2125) & (!g2373) & (g2374) & (g2375)) + ((g2073) & (!g2080) & (g2125) & (g2373) & (g2374) & (!g2375)) + ((g2073) & (!g2080) & (g2125) & (g2373) & (g2374) & (g2375)) + ((g2073) & (g2080) & (!g2125) & (g2373) & (!g2374) & (!g2375)) + ((g2073) & (g2080) & (!g2125) & (g2373) & (!g2374) & (g2375)) + ((g2073) & (g2080) & (!g2125) & (g2373) & (g2374) & (!g2375)) + ((g2073) & (g2080) & (!g2125) & (g2373) & (g2374) & (g2375)) + ((g2073) & (g2080) & (g2125) & (!g2373) & (g2374) & (!g2375)) + ((g2073) & (g2080) & (g2125) & (!g2373) & (g2374) & (g2375)) + ((g2073) & (g2080) & (g2125) & (g2373) & (g2374) & (!g2375)) + ((g2073) & (g2080) & (g2125) & (g2373) & (g2374) & (g2375)));
	assign g2377 = (((!g2365) & (!g2108) & (!g2124) & (!g2264) & (!g3663) & (!g2376)) + ((!g2365) & (!g2108) & (!g2124) & (!g2264) & (g3663) & (!g2376)) + ((!g2365) & (!g2108) & (!g2124) & (g2264) & (!g3663) & (!g2376)) + ((!g2365) & (!g2108) & (!g2124) & (g2264) & (!g3663) & (g2376)) + ((!g2365) & (!g2108) & (g2124) & (!g2264) & (!g3663) & (!g2376)) + ((!g2365) & (!g2108) & (g2124) & (!g2264) & (!g3663) & (g2376)) + ((!g2365) & (!g2108) & (g2124) & (!g2264) & (g3663) & (!g2376)) + ((!g2365) & (!g2108) & (g2124) & (!g2264) & (g3663) & (g2376)) + ((!g2365) & (!g2108) & (g2124) & (g2264) & (!g3663) & (!g2376)) + ((!g2365) & (!g2108) & (g2124) & (g2264) & (!g3663) & (g2376)) + ((!g2365) & (!g2108) & (g2124) & (g2264) & (g3663) & (!g2376)) + ((!g2365) & (!g2108) & (g2124) & (g2264) & (g3663) & (g2376)) + ((!g2365) & (g2108) & (!g2124) & (!g2264) & (!g3663) & (!g2376)) + ((!g2365) & (g2108) & (!g2124) & (!g2264) & (g3663) & (!g2376)) + ((!g2365) & (g2108) & (!g2124) & (g2264) & (!g3663) & (!g2376)) + ((!g2365) & (g2108) & (!g2124) & (g2264) & (!g3663) & (g2376)) + ((g2365) & (!g2108) & (!g2124) & (!g2264) & (!g3663) & (!g2376)) + ((g2365) & (!g2108) & (!g2124) & (!g2264) & (g3663) & (!g2376)) + ((g2365) & (!g2108) & (!g2124) & (g2264) & (!g3663) & (!g2376)) + ((g2365) & (!g2108) & (!g2124) & (g2264) & (!g3663) & (g2376)) + ((g2365) & (g2108) & (!g2124) & (!g2264) & (!g3663) & (!g2376)) + ((g2365) & (g2108) & (!g2124) & (!g2264) & (g3663) & (!g2376)) + ((g2365) & (g2108) & (!g2124) & (g2264) & (!g3663) & (!g2376)) + ((g2365) & (g2108) & (!g2124) & (g2264) & (!g3663) & (g2376)) + ((g2365) & (g2108) & (g2124) & (g2264) & (!g3663) & (!g2376)) + ((g2365) & (g2108) & (g2124) & (g2264) & (!g3663) & (g2376)) + ((g2365) & (g2108) & (g2124) & (g2264) & (g3663) & (!g2376)) + ((g2365) & (g2108) & (g2124) & (g2264) & (g3663) & (g2376)));
	assign g2378 = (((!g75) & (!g2108) & (!g2280) & (!g2362) & (!g2364) & (!g2377)) + ((!g75) & (!g2108) & (!g2280) & (!g2362) & (g2364) & (!g2377)) + ((!g75) & (!g2108) & (!g2280) & (g2362) & (!g2364) & (!g2377)) + ((!g75) & (!g2108) & (!g2280) & (g2362) & (g2364) & (!g2377)) + ((!g75) & (g2108) & (!g2280) & (!g2362) & (!g2364) & (!g2377)) + ((!g75) & (g2108) & (!g2280) & (!g2362) & (g2364) & (!g2377)) + ((!g75) & (g2108) & (!g2280) & (g2362) & (!g2364) & (!g2377)) + ((!g75) & (g2108) & (!g2280) & (g2362) & (g2364) & (!g2377)) + ((!g75) & (g2108) & (g2280) & (!g2362) & (!g2364) & (!g2377)) + ((!g75) & (g2108) & (g2280) & (!g2362) & (!g2364) & (g2377)) + ((!g75) & (g2108) & (g2280) & (!g2362) & (g2364) & (!g2377)) + ((!g75) & (g2108) & (g2280) & (!g2362) & (g2364) & (g2377)) + ((!g75) & (g2108) & (g2280) & (g2362) & (!g2364) & (!g2377)) + ((!g75) & (g2108) & (g2280) & (g2362) & (!g2364) & (g2377)) + ((!g75) & (g2108) & (g2280) & (g2362) & (g2364) & (!g2377)) + ((!g75) & (g2108) & (g2280) & (g2362) & (g2364) & (g2377)) + ((g75) & (!g2108) & (!g2280) & (!g2362) & (g2364) & (!g2377)) + ((g75) & (!g2108) & (!g2280) & (!g2362) & (g2364) & (g2377)) + ((g75) & (!g2108) & (!g2280) & (g2362) & (!g2364) & (!g2377)) + ((g75) & (!g2108) & (!g2280) & (g2362) & (!g2364) & (g2377)) + ((g75) & (!g2108) & (!g2280) & (g2362) & (g2364) & (!g2377)) + ((g75) & (!g2108) & (!g2280) & (g2362) & (g2364) & (g2377)) + ((g75) & (!g2108) & (g2280) & (!g2362) & (g2364) & (!g2377)) + ((g75) & (!g2108) & (g2280) & (!g2362) & (g2364) & (g2377)) + ((g75) & (!g2108) & (g2280) & (g2362) & (!g2364) & (!g2377)) + ((g75) & (!g2108) & (g2280) & (g2362) & (!g2364) & (g2377)) + ((g75) & (!g2108) & (g2280) & (g2362) & (g2364) & (!g2377)) + ((g75) & (!g2108) & (g2280) & (g2362) & (g2364) & (g2377)) + ((g75) & (g2108) & (!g2280) & (!g2362) & (g2364) & (!g2377)) + ((g75) & (g2108) & (!g2280) & (!g2362) & (g2364) & (g2377)) + ((g75) & (g2108) & (!g2280) & (g2362) & (!g2364) & (!g2377)) + ((g75) & (g2108) & (!g2280) & (g2362) & (!g2364) & (g2377)) + ((g75) & (g2108) & (!g2280) & (g2362) & (g2364) & (!g2377)) + ((g75) & (g2108) & (!g2280) & (g2362) & (g2364) & (g2377)) + ((g75) & (g2108) & (g2280) & (!g2362) & (g2364) & (!g2377)) + ((g75) & (g2108) & (g2280) & (!g2362) & (g2364) & (g2377)) + ((g75) & (g2108) & (g2280) & (g2362) & (!g2364) & (!g2377)) + ((g75) & (g2108) & (g2280) & (g2362) & (!g2364) & (g2377)) + ((g75) & (g2108) & (g2280) & (g2362) & (g2364) & (!g2377)) + ((g75) & (g2108) & (g2280) & (g2362) & (g2364) & (g2377)));
	assign g2379 = (((!g104) & (sk[89]) & (!g122)) + ((!g104) & (sk[89]) & (g122)) + ((g104) & (!sk[89]) & (!g122)) + ((g104) & (!sk[89]) & (g122)) + ((g104) & (sk[89]) & (!g122)));
	assign g2380 = (((!g496) & (!g541) & (!g453) & (!sk[90]) & (g2331)) + ((!g496) & (!g541) & (g453) & (!sk[90]) & (!g2331)) + ((!g496) & (!g541) & (g453) & (!sk[90]) & (g2331)) + ((!g496) & (!g541) & (g453) & (sk[90]) & (g2331)) + ((!g496) & (g541) & (!g453) & (!sk[90]) & (!g2331)) + ((!g496) & (g541) & (!g453) & (!sk[90]) & (g2331)) + ((!g496) & (g541) & (!g453) & (sk[90]) & (!g2331)) + ((!g496) & (g541) & (!g453) & (sk[90]) & (g2331)) + ((!g496) & (g541) & (g453) & (!sk[90]) & (!g2331)) + ((!g496) & (g541) & (g453) & (!sk[90]) & (g2331)) + ((!g496) & (g541) & (g453) & (sk[90]) & (!g2331)) + ((g496) & (!g541) & (!g453) & (!sk[90]) & (g2331)) + ((g496) & (!g541) & (g453) & (!sk[90]) & (!g2331)) + ((g496) & (!g541) & (g453) & (!sk[90]) & (g2331)) + ((g496) & (g541) & (!g453) & (!sk[90]) & (!g2331)) + ((g496) & (g541) & (!g453) & (!sk[90]) & (g2331)) + ((g496) & (g541) & (!g453) & (sk[90]) & (!g2331)) + ((g496) & (g541) & (!g453) & (sk[90]) & (g2331)) + ((g496) & (g541) & (g453) & (!sk[90]) & (!g2331)) + ((g496) & (g541) & (g453) & (!sk[90]) & (g2331)) + ((g496) & (g541) & (g453) & (sk[90]) & (!g2331)) + ((g496) & (g541) & (g453) & (sk[90]) & (g2331)));
	assign g2381 = (((!g2028) & (sk[91]) & (g2380)) + ((g2028) & (!sk[91]) & (!g2380)) + ((g2028) & (!sk[91]) & (g2380)));
	assign g2382 = (((g2022) & (!nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (g2381)) + ((g2022) & (!nmi_i) & (!g2023) & (!intr_i) & (g2330) & (g2381)) + ((g2022) & (!nmi_i) & (!g2023) & (intr_i) & (!g2330) & (!g2381)) + ((g2022) & (!nmi_i) & (!g2023) & (intr_i) & (!g2330) & (g2381)) + ((g2022) & (!nmi_i) & (!g2023) & (intr_i) & (g2330) & (g2381)) + ((g2022) & (!nmi_i) & (g2023) & (!intr_i) & (!g2330) & (!g2381)) + ((g2022) & (!nmi_i) & (g2023) & (!intr_i) & (!g2330) & (g2381)) + ((g2022) & (!nmi_i) & (g2023) & (!intr_i) & (g2330) & (!g2381)) + ((g2022) & (!nmi_i) & (g2023) & (!intr_i) & (g2330) & (g2381)) + ((g2022) & (!nmi_i) & (g2023) & (intr_i) & (!g2330) & (!g2381)) + ((g2022) & (!nmi_i) & (g2023) & (intr_i) & (!g2330) & (g2381)) + ((g2022) & (!nmi_i) & (g2023) & (intr_i) & (g2330) & (!g2381)) + ((g2022) & (!nmi_i) & (g2023) & (intr_i) & (g2330) & (g2381)) + ((g2022) & (nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (!g2381)) + ((g2022) & (nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (g2381)) + ((g2022) & (nmi_i) & (!g2023) & (!intr_i) & (g2330) & (!g2381)) + ((g2022) & (nmi_i) & (!g2023) & (!intr_i) & (g2330) & (g2381)) + ((g2022) & (nmi_i) & (!g2023) & (intr_i) & (!g2330) & (!g2381)) + ((g2022) & (nmi_i) & (!g2023) & (intr_i) & (!g2330) & (g2381)) + ((g2022) & (nmi_i) & (!g2023) & (intr_i) & (g2330) & (!g2381)) + ((g2022) & (nmi_i) & (!g2023) & (intr_i) & (g2330) & (g2381)) + ((g2022) & (nmi_i) & (g2023) & (!intr_i) & (!g2330) & (!g2381)) + ((g2022) & (nmi_i) & (g2023) & (!intr_i) & (!g2330) & (g2381)) + ((g2022) & (nmi_i) & (g2023) & (!intr_i) & (g2330) & (!g2381)) + ((g2022) & (nmi_i) & (g2023) & (!intr_i) & (g2330) & (g2381)) + ((g2022) & (nmi_i) & (g2023) & (intr_i) & (!g2330) & (!g2381)) + ((g2022) & (nmi_i) & (g2023) & (intr_i) & (!g2330) & (g2381)) + ((g2022) & (nmi_i) & (g2023) & (intr_i) & (g2330) & (!g2381)) + ((g2022) & (nmi_i) & (g2023) & (intr_i) & (g2330) & (g2381)));
	assign g5033 = (((!g2921) & (!g3070) & (!sk[93]) & (g2383)) + ((!g2921) & (!g3070) & (sk[93]) & (g2383)) + ((!g2921) & (g3070) & (!sk[93]) & (!g2383)) + ((!g2921) & (g3070) & (!sk[93]) & (g2383)) + ((!g2921) & (g3070) & (sk[93]) & (g2383)) + ((g2921) & (!g3070) & (!sk[93]) & (g2383)) + ((g2921) & (g3070) & (!sk[93]) & (!g2383)) + ((g2921) & (g3070) & (!sk[93]) & (g2383)) + ((g2921) & (g3070) & (sk[93]) & (!g2383)) + ((g2921) & (g3070) & (sk[93]) & (g2383)));
	assign g2384 = (((!g110) & (!g114) & (!g2030) & (!g115) & (sk[94]) & (!g2031)) + ((!g110) & (!g114) & (!g2030) & (g115) & (!sk[94]) & (!g2031)) + ((!g110) & (!g114) & (!g2030) & (g115) & (!sk[94]) & (g2031)) + ((!g110) & (!g114) & (!g2030) & (g115) & (sk[94]) & (!g2031)) + ((!g110) & (!g114) & (g2030) & (!g115) & (!sk[94]) & (!g2031)) + ((!g110) & (!g114) & (g2030) & (!g115) & (!sk[94]) & (g2031)) + ((!g110) & (!g114) & (g2030) & (g115) & (!sk[94]) & (!g2031)) + ((!g110) & (!g114) & (g2030) & (g115) & (!sk[94]) & (g2031)) + ((!g110) & (g114) & (!g2030) & (!g115) & (!sk[94]) & (!g2031)) + ((!g110) & (g114) & (!g2030) & (!g115) & (!sk[94]) & (g2031)) + ((!g110) & (g114) & (!g2030) & (!g115) & (sk[94]) & (!g2031)) + ((!g110) & (g114) & (!g2030) & (g115) & (!sk[94]) & (!g2031)) + ((!g110) & (g114) & (!g2030) & (g115) & (!sk[94]) & (g2031)) + ((!g110) & (g114) & (g2030) & (!g115) & (!sk[94]) & (!g2031)) + ((!g110) & (g114) & (g2030) & (!g115) & (!sk[94]) & (g2031)) + ((!g110) & (g114) & (g2030) & (g115) & (!sk[94]) & (!g2031)) + ((!g110) & (g114) & (g2030) & (g115) & (!sk[94]) & (g2031)) + ((g110) & (!g114) & (!g2030) & (!g115) & (sk[94]) & (!g2031)) + ((g110) & (!g114) & (!g2030) & (g115) & (!sk[94]) & (!g2031)) + ((g110) & (!g114) & (!g2030) & (g115) & (!sk[94]) & (g2031)) + ((g110) & (!g114) & (!g2030) & (g115) & (sk[94]) & (!g2031)) + ((g110) & (!g114) & (g2030) & (!g115) & (!sk[94]) & (!g2031)) + ((g110) & (!g114) & (g2030) & (!g115) & (!sk[94]) & (g2031)) + ((g110) & (!g114) & (g2030) & (g115) & (!sk[94]) & (!g2031)) + ((g110) & (!g114) & (g2030) & (g115) & (!sk[94]) & (g2031)) + ((g110) & (g114) & (!g2030) & (!g115) & (!sk[94]) & (!g2031)) + ((g110) & (g114) & (!g2030) & (!g115) & (!sk[94]) & (g2031)) + ((g110) & (g114) & (!g2030) & (!g115) & (sk[94]) & (!g2031)) + ((g110) & (g114) & (!g2030) & (g115) & (!sk[94]) & (!g2031)) + ((g110) & (g114) & (!g2030) & (g115) & (!sk[94]) & (g2031)) + ((g110) & (g114) & (!g2030) & (g115) & (sk[94]) & (!g2031)) + ((g110) & (g114) & (g2030) & (!g115) & (!sk[94]) & (!g2031)) + ((g110) & (g114) & (g2030) & (!g115) & (!sk[94]) & (g2031)) + ((g110) & (g114) & (g2030) & (g115) & (!sk[94]) & (!g2031)) + ((g110) & (g114) & (g2030) & (g115) & (!sk[94]) & (g2031)));
	assign g2385 = (((!g86) & (!sk[95]) & (!g496) & (g2358)) + ((!g86) & (!sk[95]) & (g496) & (!g2358)) + ((!g86) & (!sk[95]) & (g496) & (g2358)) + ((!g86) & (sk[95]) & (!g496) & (g2358)) + ((g86) & (!sk[95]) & (!g496) & (g2358)) + ((g86) & (!sk[95]) & (g496) & (!g2358)) + ((g86) & (!sk[95]) & (g496) & (g2358)) + ((g86) & (sk[95]) & (!g496) & (!g2358)) + ((g86) & (sk[95]) & (!g496) & (g2358)) + ((g86) & (sk[95]) & (g496) & (g2358)));
	assign g2386 = (((!g85) & (!g541) & (!sk[96]) & (!g2032) & (g2384) & (!g2385)) + ((!g85) & (!g541) & (!sk[96]) & (!g2032) & (g2384) & (g2385)) + ((!g85) & (!g541) & (!sk[96]) & (g2032) & (!g2384) & (!g2385)) + ((!g85) & (!g541) & (!sk[96]) & (g2032) & (!g2384) & (g2385)) + ((!g85) & (!g541) & (!sk[96]) & (g2032) & (g2384) & (!g2385)) + ((!g85) & (!g541) & (!sk[96]) & (g2032) & (g2384) & (g2385)) + ((!g85) & (!g541) & (sk[96]) & (!g2032) & (g2384) & (g2385)) + ((!g85) & (!g541) & (sk[96]) & (g2032) & (!g2384) & (g2385)) + ((!g85) & (!g541) & (sk[96]) & (g2032) & (g2384) & (g2385)) + ((!g85) & (g541) & (!sk[96]) & (!g2032) & (!g2384) & (!g2385)) + ((!g85) & (g541) & (!sk[96]) & (!g2032) & (!g2384) & (g2385)) + ((!g85) & (g541) & (!sk[96]) & (!g2032) & (g2384) & (!g2385)) + ((!g85) & (g541) & (!sk[96]) & (!g2032) & (g2384) & (g2385)) + ((!g85) & (g541) & (!sk[96]) & (g2032) & (!g2384) & (!g2385)) + ((!g85) & (g541) & (!sk[96]) & (g2032) & (!g2384) & (g2385)) + ((!g85) & (g541) & (!sk[96]) & (g2032) & (g2384) & (!g2385)) + ((!g85) & (g541) & (!sk[96]) & (g2032) & (g2384) & (g2385)) + ((!g85) & (g541) & (sk[96]) & (!g2032) & (g2384) & (!g2385)) + ((!g85) & (g541) & (sk[96]) & (g2032) & (!g2384) & (!g2385)) + ((!g85) & (g541) & (sk[96]) & (g2032) & (g2384) & (!g2385)) + ((g85) & (!g541) & (!sk[96]) & (!g2032) & (g2384) & (!g2385)) + ((g85) & (!g541) & (!sk[96]) & (!g2032) & (g2384) & (g2385)) + ((g85) & (!g541) & (!sk[96]) & (g2032) & (!g2384) & (!g2385)) + ((g85) & (!g541) & (!sk[96]) & (g2032) & (!g2384) & (g2385)) + ((g85) & (!g541) & (!sk[96]) & (g2032) & (g2384) & (!g2385)) + ((g85) & (!g541) & (!sk[96]) & (g2032) & (g2384) & (g2385)) + ((g85) & (!g541) & (sk[96]) & (!g2032) & (g2384) & (!g2385)) + ((g85) & (!g541) & (sk[96]) & (g2032) & (!g2384) & (!g2385)) + ((g85) & (!g541) & (sk[96]) & (g2032) & (g2384) & (!g2385)) + ((g85) & (g541) & (!sk[96]) & (!g2032) & (!g2384) & (!g2385)) + ((g85) & (g541) & (!sk[96]) & (!g2032) & (!g2384) & (g2385)) + ((g85) & (g541) & (!sk[96]) & (!g2032) & (g2384) & (!g2385)) + ((g85) & (g541) & (!sk[96]) & (!g2032) & (g2384) & (g2385)) + ((g85) & (g541) & (!sk[96]) & (g2032) & (!g2384) & (!g2385)) + ((g85) & (g541) & (!sk[96]) & (g2032) & (!g2384) & (g2385)) + ((g85) & (g541) & (!sk[96]) & (g2032) & (g2384) & (!g2385)) + ((g85) & (g541) & (!sk[96]) & (g2032) & (g2384) & (g2385)) + ((g85) & (g541) & (sk[96]) & (!g2032) & (g2384) & (g2385)) + ((g85) & (g541) & (sk[96]) & (g2032) & (!g2384) & (g2385)) + ((g85) & (g541) & (sk[96]) & (g2032) & (g2384) & (g2385)));
	assign g2387 = (((!g2030) & (!g125) & (!g1720) & (!g2031) & (!g2383) & (!g2386)) + ((!g2030) & (!g125) & (!g1720) & (!g2031) & (g2383) & (!g2386)) + ((!g2030) & (!g125) & (!g1720) & (g2031) & (!g2383) & (!g2386)) + ((!g2030) & (!g125) & (!g1720) & (g2031) & (g2383) & (!g2386)) + ((!g2030) & (!g125) & (g1720) & (!g2031) & (!g2383) & (!g2386)) + ((!g2030) & (!g125) & (g1720) & (!g2031) & (g2383) & (!g2386)) + ((g2030) & (!g125) & (!g1720) & (!g2031) & (!g2383) & (!g2386)) + ((g2030) & (!g125) & (!g1720) & (g2031) & (!g2383) & (!g2386)) + ((g2030) & (!g125) & (g1720) & (!g2031) & (!g2383) & (!g2386)));
	assign g2388 = (((!g76) & (!g77) & (!g2379) & (!g2029) & (!g2382) & (!g2387)) + ((!g76) & (!g77) & (!g2379) & (!g2029) & (!g2382) & (g2387)) + ((!g76) & (!g77) & (!g2379) & (!g2029) & (g2382) & (!g2387)) + ((!g76) & (!g77) & (!g2379) & (!g2029) & (g2382) & (g2387)) + ((!g76) & (!g77) & (!g2379) & (g2029) & (!g2382) & (!g2387)) + ((!g76) & (!g77) & (!g2379) & (g2029) & (!g2382) & (g2387)) + ((!g76) & (!g77) & (!g2379) & (g2029) & (g2382) & (!g2387)) + ((!g76) & (!g77) & (!g2379) & (g2029) & (g2382) & (g2387)) + ((!g76) & (!g77) & (g2379) & (!g2029) & (!g2382) & (!g2387)) + ((!g76) & (!g77) & (g2379) & (!g2029) & (g2382) & (!g2387)) + ((!g76) & (!g77) & (g2379) & (!g2029) & (g2382) & (g2387)) + ((!g76) & (!g77) & (g2379) & (g2029) & (g2382) & (!g2387)) + ((!g76) & (!g77) & (g2379) & (g2029) & (g2382) & (g2387)) + ((!g76) & (g77) & (!g2379) & (!g2029) & (!g2382) & (!g2387)) + ((!g76) & (g77) & (!g2379) & (!g2029) & (!g2382) & (g2387)) + ((!g76) & (g77) & (!g2379) & (!g2029) & (g2382) & (!g2387)) + ((!g76) & (g77) & (!g2379) & (!g2029) & (g2382) & (g2387)) + ((!g76) & (g77) & (!g2379) & (g2029) & (!g2382) & (!g2387)) + ((!g76) & (g77) & (!g2379) & (g2029) & (!g2382) & (g2387)) + ((!g76) & (g77) & (!g2379) & (g2029) & (g2382) & (!g2387)) + ((!g76) & (g77) & (!g2379) & (g2029) & (g2382) & (g2387)) + ((g76) & (!g77) & (!g2379) & (!g2029) & (!g2382) & (!g2387)) + ((g76) & (!g77) & (!g2379) & (!g2029) & (!g2382) & (g2387)) + ((g76) & (!g77) & (!g2379) & (!g2029) & (g2382) & (!g2387)) + ((g76) & (!g77) & (!g2379) & (!g2029) & (g2382) & (g2387)) + ((g76) & (!g77) & (!g2379) & (g2029) & (!g2382) & (!g2387)) + ((g76) & (!g77) & (!g2379) & (g2029) & (!g2382) & (g2387)) + ((g76) & (!g77) & (!g2379) & (g2029) & (g2382) & (!g2387)) + ((g76) & (!g77) & (!g2379) & (g2029) & (g2382) & (g2387)) + ((g76) & (g77) & (!g2379) & (!g2029) & (!g2382) & (!g2387)) + ((g76) & (g77) & (!g2379) & (!g2029) & (!g2382) & (g2387)) + ((g76) & (g77) & (!g2379) & (!g2029) & (g2382) & (!g2387)) + ((g76) & (g77) & (!g2379) & (!g2029) & (g2382) & (g2387)) + ((g76) & (g77) & (!g2379) & (g2029) & (!g2382) & (!g2387)) + ((g76) & (g77) & (!g2379) & (g2029) & (!g2382) & (g2387)) + ((g76) & (g77) & (!g2379) & (g2029) & (g2382) & (!g2387)) + ((g76) & (g77) & (!g2379) & (g2029) & (g2382) & (g2387)));
	assign g2389 = (((g2131) & (g2132) & (!dmem_dat_ix25x) & (dmem_dat_ix9x) & (!g2128) & (g2129)) + ((g2131) & (g2132) & (dmem_dat_ix25x) & (!dmem_dat_ix9x) & (!g2128) & (!g2129)) + ((g2131) & (g2132) & (dmem_dat_ix25x) & (dmem_dat_ix9x) & (!g2128) & (!g2129)) + ((g2131) & (g2132) & (dmem_dat_ix25x) & (dmem_dat_ix9x) & (!g2128) & (g2129)));
	assign g2390 = (((!g2363) & (!g2131) & (!g2132) & (!sk[100]) & (dmem_dat_ix9x) & (!g2338)) + ((!g2363) & (!g2131) & (!g2132) & (!sk[100]) & (dmem_dat_ix9x) & (g2338)) + ((!g2363) & (!g2131) & (g2132) & (!sk[100]) & (!dmem_dat_ix9x) & (!g2338)) + ((!g2363) & (!g2131) & (g2132) & (!sk[100]) & (!dmem_dat_ix9x) & (g2338)) + ((!g2363) & (!g2131) & (g2132) & (!sk[100]) & (dmem_dat_ix9x) & (!g2338)) + ((!g2363) & (!g2131) & (g2132) & (!sk[100]) & (dmem_dat_ix9x) & (g2338)) + ((!g2363) & (g2131) & (!g2132) & (!sk[100]) & (!dmem_dat_ix9x) & (!g2338)) + ((!g2363) & (g2131) & (!g2132) & (!sk[100]) & (!dmem_dat_ix9x) & (g2338)) + ((!g2363) & (g2131) & (!g2132) & (!sk[100]) & (dmem_dat_ix9x) & (!g2338)) + ((!g2363) & (g2131) & (!g2132) & (!sk[100]) & (dmem_dat_ix9x) & (g2338)) + ((!g2363) & (g2131) & (!g2132) & (sk[100]) & (dmem_dat_ix9x) & (!g2338)) + ((!g2363) & (g2131) & (!g2132) & (sk[100]) & (dmem_dat_ix9x) & (g2338)) + ((!g2363) & (g2131) & (g2132) & (!sk[100]) & (!dmem_dat_ix9x) & (!g2338)) + ((!g2363) & (g2131) & (g2132) & (!sk[100]) & (!dmem_dat_ix9x) & (g2338)) + ((!g2363) & (g2131) & (g2132) & (!sk[100]) & (dmem_dat_ix9x) & (!g2338)) + ((!g2363) & (g2131) & (g2132) & (!sk[100]) & (dmem_dat_ix9x) & (g2338)) + ((g2363) & (!g2131) & (!g2132) & (!sk[100]) & (dmem_dat_ix9x) & (!g2338)) + ((g2363) & (!g2131) & (!g2132) & (!sk[100]) & (dmem_dat_ix9x) & (g2338)) + ((g2363) & (!g2131) & (!g2132) & (sk[100]) & (!dmem_dat_ix9x) & (g2338)) + ((g2363) & (!g2131) & (!g2132) & (sk[100]) & (dmem_dat_ix9x) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (!sk[100]) & (!dmem_dat_ix9x) & (!g2338)) + ((g2363) & (!g2131) & (g2132) & (!sk[100]) & (!dmem_dat_ix9x) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (!sk[100]) & (dmem_dat_ix9x) & (!g2338)) + ((g2363) & (!g2131) & (g2132) & (!sk[100]) & (dmem_dat_ix9x) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (sk[100]) & (!dmem_dat_ix9x) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (sk[100]) & (dmem_dat_ix9x) & (g2338)) + ((g2363) & (g2131) & (!g2132) & (!sk[100]) & (!dmem_dat_ix9x) & (!g2338)) + ((g2363) & (g2131) & (!g2132) & (!sk[100]) & (!dmem_dat_ix9x) & (g2338)) + ((g2363) & (g2131) & (!g2132) & (!sk[100]) & (dmem_dat_ix9x) & (!g2338)) + ((g2363) & (g2131) & (!g2132) & (!sk[100]) & (dmem_dat_ix9x) & (g2338)) + ((g2363) & (g2131) & (!g2132) & (sk[100]) & (dmem_dat_ix9x) & (!g2338)) + ((g2363) & (g2131) & (!g2132) & (sk[100]) & (dmem_dat_ix9x) & (g2338)) + ((g2363) & (g2131) & (g2132) & (!sk[100]) & (!dmem_dat_ix9x) & (!g2338)) + ((g2363) & (g2131) & (g2132) & (!sk[100]) & (!dmem_dat_ix9x) & (g2338)) + ((g2363) & (g2131) & (g2132) & (!sk[100]) & (dmem_dat_ix9x) & (!g2338)) + ((g2363) & (g2131) & (g2132) & (!sk[100]) & (dmem_dat_ix9x) & (g2338)));
	assign g2392 = (((!g2108) & (!sk[101]) & (!g2365) & (g2366)) + ((!g2108) & (!sk[101]) & (g2365) & (!g2366)) + ((!g2108) & (!sk[101]) & (g2365) & (g2366)) + ((!g2108) & (sk[101]) & (g2365) & (g2366)) + ((g2108) & (!sk[101]) & (!g2365) & (g2366)) + ((g2108) & (!sk[101]) & (g2365) & (!g2366)) + ((g2108) & (!sk[101]) & (g2365) & (g2366)) + ((g2108) & (sk[101]) & (!g2365) & (g2366)) + ((g2108) & (sk[101]) & (g2365) & (!g2366)) + ((g2108) & (sk[101]) & (g2365) & (g2366)));
	assign g2393 = (((!g2109) & (!sk[102]) & (!g2391) & (!g2108) & (g2365) & (!g2366)) + ((!g2109) & (!sk[102]) & (!g2391) & (!g2108) & (g2365) & (g2366)) + ((!g2109) & (!sk[102]) & (!g2391) & (g2108) & (!g2365) & (!g2366)) + ((!g2109) & (!sk[102]) & (!g2391) & (g2108) & (!g2365) & (g2366)) + ((!g2109) & (!sk[102]) & (!g2391) & (g2108) & (g2365) & (!g2366)) + ((!g2109) & (!sk[102]) & (!g2391) & (g2108) & (g2365) & (g2366)) + ((!g2109) & (!sk[102]) & (g2391) & (!g2108) & (!g2365) & (!g2366)) + ((!g2109) & (!sk[102]) & (g2391) & (!g2108) & (!g2365) & (g2366)) + ((!g2109) & (!sk[102]) & (g2391) & (!g2108) & (g2365) & (!g2366)) + ((!g2109) & (!sk[102]) & (g2391) & (!g2108) & (g2365) & (g2366)) + ((!g2109) & (!sk[102]) & (g2391) & (g2108) & (!g2365) & (!g2366)) + ((!g2109) & (!sk[102]) & (g2391) & (g2108) & (!g2365) & (g2366)) + ((!g2109) & (!sk[102]) & (g2391) & (g2108) & (g2365) & (!g2366)) + ((!g2109) & (!sk[102]) & (g2391) & (g2108) & (g2365) & (g2366)) + ((!g2109) & (sk[102]) & (!g2391) & (!g2108) & (g2365) & (g2366)) + ((!g2109) & (sk[102]) & (!g2391) & (g2108) & (!g2365) & (g2366)) + ((!g2109) & (sk[102]) & (!g2391) & (g2108) & (g2365) & (!g2366)) + ((!g2109) & (sk[102]) & (!g2391) & (g2108) & (g2365) & (g2366)) + ((!g2109) & (sk[102]) & (g2391) & (!g2108) & (!g2365) & (!g2366)) + ((!g2109) & (sk[102]) & (g2391) & (!g2108) & (!g2365) & (g2366)) + ((!g2109) & (sk[102]) & (g2391) & (!g2108) & (g2365) & (!g2366)) + ((!g2109) & (sk[102]) & (g2391) & (g2108) & (!g2365) & (!g2366)) + ((g2109) & (!sk[102]) & (!g2391) & (!g2108) & (g2365) & (!g2366)) + ((g2109) & (!sk[102]) & (!g2391) & (!g2108) & (g2365) & (g2366)) + ((g2109) & (!sk[102]) & (!g2391) & (g2108) & (!g2365) & (!g2366)) + ((g2109) & (!sk[102]) & (!g2391) & (g2108) & (!g2365) & (g2366)) + ((g2109) & (!sk[102]) & (!g2391) & (g2108) & (g2365) & (!g2366)) + ((g2109) & (!sk[102]) & (!g2391) & (g2108) & (g2365) & (g2366)) + ((g2109) & (!sk[102]) & (g2391) & (!g2108) & (!g2365) & (!g2366)) + ((g2109) & (!sk[102]) & (g2391) & (!g2108) & (!g2365) & (g2366)) + ((g2109) & (!sk[102]) & (g2391) & (!g2108) & (g2365) & (!g2366)) + ((g2109) & (!sk[102]) & (g2391) & (!g2108) & (g2365) & (g2366)) + ((g2109) & (!sk[102]) & (g2391) & (g2108) & (!g2365) & (!g2366)) + ((g2109) & (!sk[102]) & (g2391) & (g2108) & (!g2365) & (g2366)) + ((g2109) & (!sk[102]) & (g2391) & (g2108) & (g2365) & (!g2366)) + ((g2109) & (!sk[102]) & (g2391) & (g2108) & (g2365) & (g2366)) + ((g2109) & (sk[102]) & (!g2391) & (!g2108) & (!g2365) & (!g2366)) + ((g2109) & (sk[102]) & (!g2391) & (!g2108) & (!g2365) & (g2366)) + ((g2109) & (sk[102]) & (!g2391) & (!g2108) & (g2365) & (!g2366)) + ((g2109) & (sk[102]) & (!g2391) & (g2108) & (!g2365) & (!g2366)) + ((g2109) & (sk[102]) & (g2391) & (!g2108) & (g2365) & (g2366)) + ((g2109) & (sk[102]) & (g2391) & (g2108) & (!g2365) & (g2366)) + ((g2109) & (sk[102]) & (g2391) & (g2108) & (g2365) & (!g2366)) + ((g2109) & (sk[102]) & (g2391) & (g2108) & (g2365) & (g2366)));
	assign g2394 = (((!g2341) & (!g2342) & (!sk[103]) & (!g2367) & (g2393)) + ((!g2341) & (!g2342) & (!sk[103]) & (g2367) & (!g2393)) + ((!g2341) & (!g2342) & (!sk[103]) & (g2367) & (g2393)) + ((!g2341) & (!g2342) & (sk[103]) & (!g2367) & (g2393)) + ((!g2341) & (!g2342) & (sk[103]) & (g2367) & (g2393)) + ((!g2341) & (g2342) & (!sk[103]) & (!g2367) & (!g2393)) + ((!g2341) & (g2342) & (!sk[103]) & (!g2367) & (g2393)) + ((!g2341) & (g2342) & (!sk[103]) & (g2367) & (!g2393)) + ((!g2341) & (g2342) & (!sk[103]) & (g2367) & (g2393)) + ((!g2341) & (g2342) & (sk[103]) & (!g2367) & (g2393)) + ((!g2341) & (g2342) & (sk[103]) & (g2367) & (g2393)) + ((g2341) & (!g2342) & (!sk[103]) & (!g2367) & (g2393)) + ((g2341) & (!g2342) & (!sk[103]) & (g2367) & (!g2393)) + ((g2341) & (!g2342) & (!sk[103]) & (g2367) & (g2393)) + ((g2341) & (!g2342) & (sk[103]) & (!g2367) & (g2393)) + ((g2341) & (!g2342) & (sk[103]) & (g2367) & (g2393)) + ((g2341) & (g2342) & (!sk[103]) & (!g2367) & (!g2393)) + ((g2341) & (g2342) & (!sk[103]) & (!g2367) & (g2393)) + ((g2341) & (g2342) & (!sk[103]) & (g2367) & (!g2393)) + ((g2341) & (g2342) & (!sk[103]) & (g2367) & (g2393)) + ((g2341) & (g2342) & (sk[103]) & (!g2367) & (g2393)) + ((g2341) & (g2342) & (sk[103]) & (g2367) & (!g2393)));
	assign g2395 = (((!g2344) & (!g2345) & (!g2347) & (!g2348) & (!g2369) & (!g2370)) + ((!g2344) & (!g2345) & (!g2347) & (!g2348) & (!g2369) & (g2370)) + ((!g2344) & (!g2345) & (!g2347) & (!g2348) & (g2369) & (!g2370)) + ((!g2344) & (!g2345) & (!g2347) & (g2348) & (!g2369) & (!g2370)) + ((!g2344) & (!g2345) & (!g2347) & (g2348) & (!g2369) & (g2370)) + ((!g2344) & (!g2345) & (!g2347) & (g2348) & (g2369) & (!g2370)) + ((!g2344) & (!g2345) & (g2347) & (!g2348) & (!g2369) & (!g2370)) + ((!g2344) & (!g2345) & (g2347) & (!g2348) & (!g2369) & (g2370)) + ((!g2344) & (!g2345) & (g2347) & (!g2348) & (g2369) & (!g2370)) + ((!g2344) & (!g2345) & (g2347) & (g2348) & (!g2369) & (!g2370)) + ((!g2344) & (g2345) & (!g2347) & (!g2348) & (!g2369) & (!g2370)) + ((!g2344) & (g2345) & (!g2347) & (!g2348) & (!g2369) & (g2370)) + ((!g2344) & (g2345) & (!g2347) & (!g2348) & (g2369) & (!g2370)) + ((!g2344) & (g2345) & (!g2347) & (g2348) & (!g2369) & (!g2370)) + ((!g2344) & (g2345) & (g2347) & (!g2348) & (!g2369) & (!g2370)) + ((!g2344) & (g2345) & (g2347) & (g2348) & (!g2369) & (!g2370)) + ((g2344) & (!g2345) & (!g2347) & (!g2348) & (!g2369) & (!g2370)) + ((g2344) & (!g2345) & (!g2347) & (!g2348) & (!g2369) & (g2370)) + ((g2344) & (!g2345) & (!g2347) & (!g2348) & (g2369) & (!g2370)) + ((g2344) & (!g2345) & (!g2347) & (g2348) & (!g2369) & (!g2370)) + ((g2344) & (!g2345) & (g2347) & (!g2348) & (!g2369) & (!g2370)) + ((g2344) & (!g2345) & (g2347) & (g2348) & (!g2369) & (!g2370)) + ((g2344) & (g2345) & (!g2347) & (!g2348) & (!g2369) & (!g2370)) + ((g2344) & (g2345) & (!g2347) & (!g2348) & (!g2369) & (g2370)) + ((g2344) & (g2345) & (!g2347) & (!g2348) & (g2369) & (!g2370)) + ((g2344) & (g2345) & (!g2347) & (g2348) & (!g2369) & (!g2370)) + ((g2344) & (g2345) & (g2347) & (!g2348) & (!g2369) & (!g2370)) + ((g2344) & (g2345) & (g2347) & (g2348) & (!g2369) & (!g2370)));
	assign g2396 = (((g2108) & (!sk[105]) & (!g2365)) + ((g2108) & (!sk[105]) & (g2365)) + ((g2108) & (sk[105]) & (!g2365)));
	assign g2397 = (((!g2109) & (sk[106]) & (!g2391)) + ((g2109) & (!sk[106]) & (!g2391)) + ((g2109) & (!sk[106]) & (g2391)) + ((g2109) & (sk[106]) & (g2391)));
	assign g2398 = (((!g2395) & (!g2396) & (!sk[107]) & (g2397)) + ((!g2395) & (!g2396) & (sk[107]) & (!g2397)) + ((!g2395) & (g2396) & (!sk[107]) & (!g2397)) + ((!g2395) & (g2396) & (!sk[107]) & (g2397)) + ((!g2395) & (g2396) & (sk[107]) & (g2397)) + ((g2395) & (!g2396) & (!sk[107]) & (g2397)) + ((g2395) & (!g2396) & (sk[107]) & (g2397)) + ((g2395) & (g2396) & (!sk[107]) & (!g2397)) + ((g2395) & (g2396) & (!sk[107]) & (g2397)) + ((g2395) & (g2396) & (sk[107]) & (!g2397)));
	assign g2399 = (((!g2073) & (!sk[108]) & (!g2080) & (g2125)) + ((!g2073) & (!sk[108]) & (g2080) & (!g2125)) + ((!g2073) & (!sk[108]) & (g2080) & (g2125)) + ((!g2073) & (sk[108]) & (!g2080) & (g2125)) + ((!g2073) & (sk[108]) & (g2080) & (g2125)) + ((g2073) & (!sk[108]) & (!g2080) & (g2125)) + ((g2073) & (!sk[108]) & (g2080) & (!g2125)) + ((g2073) & (!sk[108]) & (g2080) & (g2125)) + ((g2073) & (sk[108]) & (!g2080) & (!g2125)));
	assign g2400 = (((!sk[109]) & (!g2073) & (!g2080) & (g2125)) + ((!sk[109]) & (!g2073) & (g2080) & (!g2125)) + ((!sk[109]) & (!g2073) & (g2080) & (g2125)) + ((!sk[109]) & (g2073) & (!g2080) & (g2125)) + ((!sk[109]) & (g2073) & (g2080) & (!g2125)) + ((!sk[109]) & (g2073) & (g2080) & (g2125)) + ((sk[109]) & (g2073) & (!g2080) & (!g2125)) + ((sk[109]) & (g2073) & (!g2080) & (g2125)) + ((sk[109]) & (g2073) & (g2080) & (g2125)));
	assign g2401 = (((!g2076) & (!g2077) & (!sk[110]) & (!g2188) & (g2192) & (!g2193)) + ((!g2076) & (!g2077) & (!sk[110]) & (!g2188) & (g2192) & (g2193)) + ((!g2076) & (!g2077) & (!sk[110]) & (g2188) & (!g2192) & (!g2193)) + ((!g2076) & (!g2077) & (!sk[110]) & (g2188) & (!g2192) & (g2193)) + ((!g2076) & (!g2077) & (!sk[110]) & (g2188) & (g2192) & (!g2193)) + ((!g2076) & (!g2077) & (!sk[110]) & (g2188) & (g2192) & (g2193)) + ((!g2076) & (!g2077) & (sk[110]) & (g2188) & (!g2192) & (!g2193)) + ((!g2076) & (!g2077) & (sk[110]) & (g2188) & (!g2192) & (g2193)) + ((!g2076) & (!g2077) & (sk[110]) & (g2188) & (g2192) & (!g2193)) + ((!g2076) & (!g2077) & (sk[110]) & (g2188) & (g2192) & (g2193)) + ((!g2076) & (g2077) & (!sk[110]) & (!g2188) & (!g2192) & (!g2193)) + ((!g2076) & (g2077) & (!sk[110]) & (!g2188) & (!g2192) & (g2193)) + ((!g2076) & (g2077) & (!sk[110]) & (!g2188) & (g2192) & (!g2193)) + ((!g2076) & (g2077) & (!sk[110]) & (!g2188) & (g2192) & (g2193)) + ((!g2076) & (g2077) & (!sk[110]) & (g2188) & (!g2192) & (!g2193)) + ((!g2076) & (g2077) & (!sk[110]) & (g2188) & (!g2192) & (g2193)) + ((!g2076) & (g2077) & (!sk[110]) & (g2188) & (g2192) & (!g2193)) + ((!g2076) & (g2077) & (!sk[110]) & (g2188) & (g2192) & (g2193)) + ((!g2076) & (g2077) & (sk[110]) & (!g2188) & (!g2192) & (g2193)) + ((!g2076) & (g2077) & (sk[110]) & (!g2188) & (g2192) & (g2193)) + ((!g2076) & (g2077) & (sk[110]) & (g2188) & (!g2192) & (g2193)) + ((!g2076) & (g2077) & (sk[110]) & (g2188) & (g2192) & (g2193)) + ((g2076) & (!g2077) & (!sk[110]) & (!g2188) & (g2192) & (!g2193)) + ((g2076) & (!g2077) & (!sk[110]) & (!g2188) & (g2192) & (g2193)) + ((g2076) & (!g2077) & (!sk[110]) & (g2188) & (!g2192) & (!g2193)) + ((g2076) & (!g2077) & (!sk[110]) & (g2188) & (!g2192) & (g2193)) + ((g2076) & (!g2077) & (!sk[110]) & (g2188) & (g2192) & (!g2193)) + ((g2076) & (!g2077) & (!sk[110]) & (g2188) & (g2192) & (g2193)) + ((g2076) & (!g2077) & (sk[110]) & (!g2188) & (g2192) & (!g2193)) + ((g2076) & (!g2077) & (sk[110]) & (!g2188) & (g2192) & (g2193)) + ((g2076) & (!g2077) & (sk[110]) & (g2188) & (g2192) & (!g2193)) + ((g2076) & (!g2077) & (sk[110]) & (g2188) & (g2192) & (g2193)) + ((g2076) & (g2077) & (!sk[110]) & (!g2188) & (!g2192) & (!g2193)) + ((g2076) & (g2077) & (!sk[110]) & (!g2188) & (!g2192) & (g2193)) + ((g2076) & (g2077) & (!sk[110]) & (!g2188) & (g2192) & (!g2193)) + ((g2076) & (g2077) & (!sk[110]) & (!g2188) & (g2192) & (g2193)) + ((g2076) & (g2077) & (!sk[110]) & (g2188) & (!g2192) & (!g2193)) + ((g2076) & (g2077) & (!sk[110]) & (g2188) & (!g2192) & (g2193)) + ((g2076) & (g2077) & (!sk[110]) & (g2188) & (g2192) & (!g2193)) + ((g2076) & (g2077) & (!sk[110]) & (g2188) & (g2192) & (g2193)) + ((g2076) & (g2077) & (sk[110]) & (!g2188) & (g2192) & (!g2193)) + ((g2076) & (g2077) & (sk[110]) & (!g2188) & (g2192) & (g2193)) + ((g2076) & (g2077) & (sk[110]) & (g2188) & (g2192) & (!g2193)) + ((g2076) & (g2077) & (sk[110]) & (g2188) & (g2192) & (g2193)));
	assign g2402 = (((!g2109) & (!g2108) & (!g2116) & (g2115) & (g2071) & (g2074)) + ((!g2109) & (!g2108) & (g2116) & (!g2115) & (!g2071) & (g2074)) + ((!g2109) & (!g2108) & (g2116) & (g2115) & (!g2071) & (g2074)) + ((!g2109) & (!g2108) & (g2116) & (g2115) & (g2071) & (g2074)) + ((!g2109) & (g2108) & (!g2116) & (!g2115) & (g2071) & (!g2074)) + ((!g2109) & (g2108) & (!g2116) & (g2115) & (g2071) & (!g2074)) + ((!g2109) & (g2108) & (!g2116) & (g2115) & (g2071) & (g2074)) + ((!g2109) & (g2108) & (g2116) & (!g2115) & (!g2071) & (g2074)) + ((!g2109) & (g2108) & (g2116) & (!g2115) & (g2071) & (!g2074)) + ((!g2109) & (g2108) & (g2116) & (g2115) & (!g2071) & (g2074)) + ((!g2109) & (g2108) & (g2116) & (g2115) & (g2071) & (!g2074)) + ((!g2109) & (g2108) & (g2116) & (g2115) & (g2071) & (g2074)) + ((g2109) & (!g2108) & (!g2116) & (!g2115) & (!g2071) & (!g2074)) + ((g2109) & (!g2108) & (!g2116) & (g2115) & (!g2071) & (!g2074)) + ((g2109) & (!g2108) & (!g2116) & (g2115) & (g2071) & (g2074)) + ((g2109) & (!g2108) & (g2116) & (!g2115) & (!g2071) & (!g2074)) + ((g2109) & (!g2108) & (g2116) & (!g2115) & (!g2071) & (g2074)) + ((g2109) & (!g2108) & (g2116) & (g2115) & (!g2071) & (!g2074)) + ((g2109) & (!g2108) & (g2116) & (g2115) & (!g2071) & (g2074)) + ((g2109) & (!g2108) & (g2116) & (g2115) & (g2071) & (g2074)) + ((g2109) & (g2108) & (!g2116) & (!g2115) & (!g2071) & (!g2074)) + ((g2109) & (g2108) & (!g2116) & (!g2115) & (g2071) & (!g2074)) + ((g2109) & (g2108) & (!g2116) & (g2115) & (!g2071) & (!g2074)) + ((g2109) & (g2108) & (!g2116) & (g2115) & (g2071) & (!g2074)) + ((g2109) & (g2108) & (!g2116) & (g2115) & (g2071) & (g2074)) + ((g2109) & (g2108) & (g2116) & (!g2115) & (!g2071) & (!g2074)) + ((g2109) & (g2108) & (g2116) & (!g2115) & (!g2071) & (g2074)) + ((g2109) & (g2108) & (g2116) & (!g2115) & (g2071) & (!g2074)) + ((g2109) & (g2108) & (g2116) & (g2115) & (!g2071) & (!g2074)) + ((g2109) & (g2108) & (g2116) & (g2115) & (!g2071) & (g2074)) + ((g2109) & (g2108) & (g2116) & (g2115) & (g2071) & (!g2074)) + ((g2109) & (g2108) & (g2116) & (g2115) & (g2071) & (g2074)));
	assign g2403 = (((!g2076) & (!g2077) & (!sk[112]) & (!g2183) & (g2296) & (!g2402)) + ((!g2076) & (!g2077) & (!sk[112]) & (!g2183) & (g2296) & (g2402)) + ((!g2076) & (!g2077) & (!sk[112]) & (g2183) & (!g2296) & (!g2402)) + ((!g2076) & (!g2077) & (!sk[112]) & (g2183) & (!g2296) & (g2402)) + ((!g2076) & (!g2077) & (!sk[112]) & (g2183) & (g2296) & (!g2402)) + ((!g2076) & (!g2077) & (!sk[112]) & (g2183) & (g2296) & (g2402)) + ((!g2076) & (!g2077) & (sk[112]) & (!g2183) & (!g2296) & (g2402)) + ((!g2076) & (!g2077) & (sk[112]) & (!g2183) & (g2296) & (g2402)) + ((!g2076) & (!g2077) & (sk[112]) & (g2183) & (!g2296) & (g2402)) + ((!g2076) & (!g2077) & (sk[112]) & (g2183) & (g2296) & (g2402)) + ((!g2076) & (g2077) & (!sk[112]) & (!g2183) & (!g2296) & (!g2402)) + ((!g2076) & (g2077) & (!sk[112]) & (!g2183) & (!g2296) & (g2402)) + ((!g2076) & (g2077) & (!sk[112]) & (!g2183) & (g2296) & (!g2402)) + ((!g2076) & (g2077) & (!sk[112]) & (!g2183) & (g2296) & (g2402)) + ((!g2076) & (g2077) & (!sk[112]) & (g2183) & (!g2296) & (!g2402)) + ((!g2076) & (g2077) & (!sk[112]) & (g2183) & (!g2296) & (g2402)) + ((!g2076) & (g2077) & (!sk[112]) & (g2183) & (g2296) & (!g2402)) + ((!g2076) & (g2077) & (!sk[112]) & (g2183) & (g2296) & (g2402)) + ((!g2076) & (g2077) & (sk[112]) & (!g2183) & (g2296) & (!g2402)) + ((!g2076) & (g2077) & (sk[112]) & (!g2183) & (g2296) & (g2402)) + ((!g2076) & (g2077) & (sk[112]) & (g2183) & (g2296) & (!g2402)) + ((!g2076) & (g2077) & (sk[112]) & (g2183) & (g2296) & (g2402)) + ((g2076) & (!g2077) & (!sk[112]) & (!g2183) & (g2296) & (!g2402)) + ((g2076) & (!g2077) & (!sk[112]) & (!g2183) & (g2296) & (g2402)) + ((g2076) & (!g2077) & (!sk[112]) & (g2183) & (!g2296) & (!g2402)) + ((g2076) & (!g2077) & (!sk[112]) & (g2183) & (!g2296) & (g2402)) + ((g2076) & (!g2077) & (!sk[112]) & (g2183) & (g2296) & (!g2402)) + ((g2076) & (!g2077) & (!sk[112]) & (g2183) & (g2296) & (g2402)) + ((g2076) & (!g2077) & (sk[112]) & (g2183) & (!g2296) & (!g2402)) + ((g2076) & (!g2077) & (sk[112]) & (g2183) & (!g2296) & (g2402)) + ((g2076) & (!g2077) & (sk[112]) & (g2183) & (g2296) & (!g2402)) + ((g2076) & (!g2077) & (sk[112]) & (g2183) & (g2296) & (g2402)) + ((g2076) & (g2077) & (!sk[112]) & (!g2183) & (!g2296) & (!g2402)) + ((g2076) & (g2077) & (!sk[112]) & (!g2183) & (!g2296) & (g2402)) + ((g2076) & (g2077) & (!sk[112]) & (!g2183) & (g2296) & (!g2402)) + ((g2076) & (g2077) & (!sk[112]) & (!g2183) & (g2296) & (g2402)) + ((g2076) & (g2077) & (!sk[112]) & (g2183) & (!g2296) & (!g2402)) + ((g2076) & (g2077) & (!sk[112]) & (g2183) & (!g2296) & (g2402)) + ((g2076) & (g2077) & (!sk[112]) & (g2183) & (g2296) & (!g2402)) + ((g2076) & (g2077) & (!sk[112]) & (g2183) & (g2296) & (g2402)));
	assign g2404 = (((!g2199) & (!g2187) & (!g2200) & (g2189) & (g2076) & (g2077)) + ((!g2199) & (!g2187) & (g2200) & (!g2189) & (!g2076) & (g2077)) + ((!g2199) & (!g2187) & (g2200) & (g2189) & (!g2076) & (g2077)) + ((!g2199) & (!g2187) & (g2200) & (g2189) & (g2076) & (g2077)) + ((!g2199) & (g2187) & (!g2200) & (!g2189) & (g2076) & (!g2077)) + ((!g2199) & (g2187) & (!g2200) & (g2189) & (g2076) & (!g2077)) + ((!g2199) & (g2187) & (!g2200) & (g2189) & (g2076) & (g2077)) + ((!g2199) & (g2187) & (g2200) & (!g2189) & (!g2076) & (g2077)) + ((!g2199) & (g2187) & (g2200) & (!g2189) & (g2076) & (!g2077)) + ((!g2199) & (g2187) & (g2200) & (g2189) & (!g2076) & (g2077)) + ((!g2199) & (g2187) & (g2200) & (g2189) & (g2076) & (!g2077)) + ((!g2199) & (g2187) & (g2200) & (g2189) & (g2076) & (g2077)) + ((g2199) & (!g2187) & (!g2200) & (!g2189) & (!g2076) & (!g2077)) + ((g2199) & (!g2187) & (!g2200) & (g2189) & (!g2076) & (!g2077)) + ((g2199) & (!g2187) & (!g2200) & (g2189) & (g2076) & (g2077)) + ((g2199) & (!g2187) & (g2200) & (!g2189) & (!g2076) & (!g2077)) + ((g2199) & (!g2187) & (g2200) & (!g2189) & (!g2076) & (g2077)) + ((g2199) & (!g2187) & (g2200) & (g2189) & (!g2076) & (!g2077)) + ((g2199) & (!g2187) & (g2200) & (g2189) & (!g2076) & (g2077)) + ((g2199) & (!g2187) & (g2200) & (g2189) & (g2076) & (g2077)) + ((g2199) & (g2187) & (!g2200) & (!g2189) & (!g2076) & (!g2077)) + ((g2199) & (g2187) & (!g2200) & (!g2189) & (g2076) & (!g2077)) + ((g2199) & (g2187) & (!g2200) & (g2189) & (!g2076) & (!g2077)) + ((g2199) & (g2187) & (!g2200) & (g2189) & (g2076) & (!g2077)) + ((g2199) & (g2187) & (!g2200) & (g2189) & (g2076) & (g2077)) + ((g2199) & (g2187) & (g2200) & (!g2189) & (!g2076) & (!g2077)) + ((g2199) & (g2187) & (g2200) & (!g2189) & (!g2076) & (g2077)) + ((g2199) & (g2187) & (g2200) & (!g2189) & (g2076) & (!g2077)) + ((g2199) & (g2187) & (g2200) & (g2189) & (!g2076) & (!g2077)) + ((g2199) & (g2187) & (g2200) & (g2189) & (!g2076) & (g2077)) + ((g2199) & (g2187) & (g2200) & (g2189) & (g2076) & (!g2077)) + ((g2199) & (g2187) & (g2200) & (g2189) & (g2076) & (g2077)));
	assign g2405 = (((!g2399) & (!g2400) & (!g2401) & (!sk[114]) & (g2403) & (!g2404)) + ((!g2399) & (!g2400) & (!g2401) & (!sk[114]) & (g2403) & (g2404)) + ((!g2399) & (!g2400) & (!g2401) & (sk[114]) & (g2403) & (!g2404)) + ((!g2399) & (!g2400) & (!g2401) & (sk[114]) & (g2403) & (g2404)) + ((!g2399) & (!g2400) & (g2401) & (!sk[114]) & (!g2403) & (!g2404)) + ((!g2399) & (!g2400) & (g2401) & (!sk[114]) & (!g2403) & (g2404)) + ((!g2399) & (!g2400) & (g2401) & (!sk[114]) & (g2403) & (!g2404)) + ((!g2399) & (!g2400) & (g2401) & (!sk[114]) & (g2403) & (g2404)) + ((!g2399) & (!g2400) & (g2401) & (sk[114]) & (g2403) & (!g2404)) + ((!g2399) & (!g2400) & (g2401) & (sk[114]) & (g2403) & (g2404)) + ((!g2399) & (g2400) & (!g2401) & (!sk[114]) & (!g2403) & (!g2404)) + ((!g2399) & (g2400) & (!g2401) & (!sk[114]) & (!g2403) & (g2404)) + ((!g2399) & (g2400) & (!g2401) & (!sk[114]) & (g2403) & (!g2404)) + ((!g2399) & (g2400) & (!g2401) & (!sk[114]) & (g2403) & (g2404)) + ((!g2399) & (g2400) & (g2401) & (!sk[114]) & (!g2403) & (!g2404)) + ((!g2399) & (g2400) & (g2401) & (!sk[114]) & (!g2403) & (g2404)) + ((!g2399) & (g2400) & (g2401) & (!sk[114]) & (g2403) & (!g2404)) + ((!g2399) & (g2400) & (g2401) & (!sk[114]) & (g2403) & (g2404)) + ((!g2399) & (g2400) & (g2401) & (sk[114]) & (!g2403) & (!g2404)) + ((!g2399) & (g2400) & (g2401) & (sk[114]) & (!g2403) & (g2404)) + ((!g2399) & (g2400) & (g2401) & (sk[114]) & (g2403) & (!g2404)) + ((!g2399) & (g2400) & (g2401) & (sk[114]) & (g2403) & (g2404)) + ((g2399) & (!g2400) & (!g2401) & (!sk[114]) & (g2403) & (!g2404)) + ((g2399) & (!g2400) & (!g2401) & (!sk[114]) & (g2403) & (g2404)) + ((g2399) & (!g2400) & (!g2401) & (sk[114]) & (!g2403) & (g2404)) + ((g2399) & (!g2400) & (!g2401) & (sk[114]) & (g2403) & (g2404)) + ((g2399) & (!g2400) & (g2401) & (!sk[114]) & (!g2403) & (!g2404)) + ((g2399) & (!g2400) & (g2401) & (!sk[114]) & (!g2403) & (g2404)) + ((g2399) & (!g2400) & (g2401) & (!sk[114]) & (g2403) & (!g2404)) + ((g2399) & (!g2400) & (g2401) & (!sk[114]) & (g2403) & (g2404)) + ((g2399) & (!g2400) & (g2401) & (sk[114]) & (!g2403) & (g2404)) + ((g2399) & (!g2400) & (g2401) & (sk[114]) & (g2403) & (g2404)) + ((g2399) & (g2400) & (!g2401) & (!sk[114]) & (!g2403) & (!g2404)) + ((g2399) & (g2400) & (!g2401) & (!sk[114]) & (!g2403) & (g2404)) + ((g2399) & (g2400) & (!g2401) & (!sk[114]) & (g2403) & (!g2404)) + ((g2399) & (g2400) & (!g2401) & (!sk[114]) & (g2403) & (g2404)) + ((g2399) & (g2400) & (g2401) & (!sk[114]) & (!g2403) & (!g2404)) + ((g2399) & (g2400) & (g2401) & (!sk[114]) & (!g2403) & (g2404)) + ((g2399) & (g2400) & (g2401) & (!sk[114]) & (g2403) & (!g2404)) + ((g2399) & (g2400) & (g2401) & (!sk[114]) & (g2403) & (g2404)));
	assign g2406 = (((!g2391) & (!g2109) & (!g2124) & (!g2264) & (!g3650) & (!g2405)) + ((!g2391) & (!g2109) & (!g2124) & (!g2264) & (g3650) & (!g2405)) + ((!g2391) & (!g2109) & (!g2124) & (g2264) & (!g3650) & (!g2405)) + ((!g2391) & (!g2109) & (!g2124) & (g2264) & (!g3650) & (g2405)) + ((!g2391) & (!g2109) & (g2124) & (!g2264) & (!g3650) & (!g2405)) + ((!g2391) & (!g2109) & (g2124) & (!g2264) & (!g3650) & (g2405)) + ((!g2391) & (!g2109) & (g2124) & (!g2264) & (g3650) & (!g2405)) + ((!g2391) & (!g2109) & (g2124) & (!g2264) & (g3650) & (g2405)) + ((!g2391) & (!g2109) & (g2124) & (g2264) & (!g3650) & (!g2405)) + ((!g2391) & (!g2109) & (g2124) & (g2264) & (!g3650) & (g2405)) + ((!g2391) & (!g2109) & (g2124) & (g2264) & (g3650) & (!g2405)) + ((!g2391) & (!g2109) & (g2124) & (g2264) & (g3650) & (g2405)) + ((!g2391) & (g2109) & (!g2124) & (!g2264) & (!g3650) & (!g2405)) + ((!g2391) & (g2109) & (!g2124) & (!g2264) & (g3650) & (!g2405)) + ((!g2391) & (g2109) & (!g2124) & (g2264) & (!g3650) & (!g2405)) + ((!g2391) & (g2109) & (!g2124) & (g2264) & (!g3650) & (g2405)) + ((g2391) & (!g2109) & (!g2124) & (!g2264) & (!g3650) & (!g2405)) + ((g2391) & (!g2109) & (!g2124) & (!g2264) & (g3650) & (!g2405)) + ((g2391) & (!g2109) & (!g2124) & (g2264) & (!g3650) & (!g2405)) + ((g2391) & (!g2109) & (!g2124) & (g2264) & (!g3650) & (g2405)) + ((g2391) & (g2109) & (!g2124) & (!g2264) & (!g3650) & (!g2405)) + ((g2391) & (g2109) & (!g2124) & (!g2264) & (g3650) & (!g2405)) + ((g2391) & (g2109) & (!g2124) & (g2264) & (!g3650) & (!g2405)) + ((g2391) & (g2109) & (!g2124) & (g2264) & (!g3650) & (g2405)) + ((g2391) & (g2109) & (g2124) & (g2264) & (!g3650) & (!g2405)) + ((g2391) & (g2109) & (g2124) & (g2264) & (!g3650) & (g2405)) + ((g2391) & (g2109) & (g2124) & (g2264) & (g3650) & (!g2405)) + ((g2391) & (g2109) & (g2124) & (g2264) & (g3650) & (g2405)));
	assign g2407 = (((!g75) & (!g2109) & (!g2280) & (!g2389) & (!g2390) & (!g2406)) + ((!g75) & (!g2109) & (!g2280) & (!g2389) & (g2390) & (!g2406)) + ((!g75) & (!g2109) & (!g2280) & (g2389) & (!g2390) & (!g2406)) + ((!g75) & (!g2109) & (!g2280) & (g2389) & (g2390) & (!g2406)) + ((!g75) & (g2109) & (!g2280) & (!g2389) & (!g2390) & (!g2406)) + ((!g75) & (g2109) & (!g2280) & (!g2389) & (g2390) & (!g2406)) + ((!g75) & (g2109) & (!g2280) & (g2389) & (!g2390) & (!g2406)) + ((!g75) & (g2109) & (!g2280) & (g2389) & (g2390) & (!g2406)) + ((!g75) & (g2109) & (g2280) & (!g2389) & (!g2390) & (!g2406)) + ((!g75) & (g2109) & (g2280) & (!g2389) & (!g2390) & (g2406)) + ((!g75) & (g2109) & (g2280) & (!g2389) & (g2390) & (!g2406)) + ((!g75) & (g2109) & (g2280) & (!g2389) & (g2390) & (g2406)) + ((!g75) & (g2109) & (g2280) & (g2389) & (!g2390) & (!g2406)) + ((!g75) & (g2109) & (g2280) & (g2389) & (!g2390) & (g2406)) + ((!g75) & (g2109) & (g2280) & (g2389) & (g2390) & (!g2406)) + ((!g75) & (g2109) & (g2280) & (g2389) & (g2390) & (g2406)) + ((g75) & (!g2109) & (!g2280) & (!g2389) & (g2390) & (!g2406)) + ((g75) & (!g2109) & (!g2280) & (!g2389) & (g2390) & (g2406)) + ((g75) & (!g2109) & (!g2280) & (g2389) & (!g2390) & (!g2406)) + ((g75) & (!g2109) & (!g2280) & (g2389) & (!g2390) & (g2406)) + ((g75) & (!g2109) & (!g2280) & (g2389) & (g2390) & (!g2406)) + ((g75) & (!g2109) & (!g2280) & (g2389) & (g2390) & (g2406)) + ((g75) & (!g2109) & (g2280) & (!g2389) & (g2390) & (!g2406)) + ((g75) & (!g2109) & (g2280) & (!g2389) & (g2390) & (g2406)) + ((g75) & (!g2109) & (g2280) & (g2389) & (!g2390) & (!g2406)) + ((g75) & (!g2109) & (g2280) & (g2389) & (!g2390) & (g2406)) + ((g75) & (!g2109) & (g2280) & (g2389) & (g2390) & (!g2406)) + ((g75) & (!g2109) & (g2280) & (g2389) & (g2390) & (g2406)) + ((g75) & (g2109) & (!g2280) & (!g2389) & (g2390) & (!g2406)) + ((g75) & (g2109) & (!g2280) & (!g2389) & (g2390) & (g2406)) + ((g75) & (g2109) & (!g2280) & (g2389) & (!g2390) & (!g2406)) + ((g75) & (g2109) & (!g2280) & (g2389) & (!g2390) & (g2406)) + ((g75) & (g2109) & (!g2280) & (g2389) & (g2390) & (!g2406)) + ((g75) & (g2109) & (!g2280) & (g2389) & (g2390) & (g2406)) + ((g75) & (g2109) & (g2280) & (!g2389) & (g2390) & (!g2406)) + ((g75) & (g2109) & (g2280) & (!g2389) & (g2390) & (g2406)) + ((g75) & (g2109) & (g2280) & (g2389) & (!g2390) & (!g2406)) + ((g75) & (g2109) & (g2280) & (g2389) & (!g2390) & (g2406)) + ((g75) & (g2109) & (g2280) & (g2389) & (g2390) & (!g2406)) + ((g75) & (g2109) & (g2280) & (g2389) & (g2390) & (g2406)));
	assign g2408 = (((!g2022) & (!g123) & (!nmi_i) & (!g2023) & (!intr_i) & (!g2330)) + ((!g2022) & (!g123) & (!nmi_i) & (!g2023) & (!intr_i) & (g2330)) + ((!g2022) & (!g123) & (!nmi_i) & (!g2023) & (intr_i) & (!g2330)) + ((!g2022) & (!g123) & (!nmi_i) & (!g2023) & (intr_i) & (g2330)) + ((!g2022) & (!g123) & (!nmi_i) & (g2023) & (!intr_i) & (!g2330)) + ((!g2022) & (!g123) & (!nmi_i) & (g2023) & (!intr_i) & (g2330)) + ((!g2022) & (!g123) & (!nmi_i) & (g2023) & (intr_i) & (!g2330)) + ((!g2022) & (!g123) & (!nmi_i) & (g2023) & (intr_i) & (g2330)) + ((!g2022) & (!g123) & (nmi_i) & (!g2023) & (!intr_i) & (!g2330)) + ((!g2022) & (!g123) & (nmi_i) & (!g2023) & (!intr_i) & (g2330)) + ((!g2022) & (!g123) & (nmi_i) & (!g2023) & (intr_i) & (!g2330)) + ((!g2022) & (!g123) & (nmi_i) & (!g2023) & (intr_i) & (g2330)) + ((!g2022) & (!g123) & (nmi_i) & (g2023) & (!intr_i) & (!g2330)) + ((!g2022) & (!g123) & (nmi_i) & (g2023) & (!intr_i) & (g2330)) + ((!g2022) & (!g123) & (nmi_i) & (g2023) & (intr_i) & (!g2330)) + ((!g2022) & (!g123) & (nmi_i) & (g2023) & (intr_i) & (g2330)) + ((g2022) & (!g123) & (!nmi_i) & (!g2023) & (!intr_i) & (!g2330)) + ((g2022) & (!g123) & (!nmi_i) & (!g2023) & (!intr_i) & (g2330)) + ((g2022) & (!g123) & (!nmi_i) & (!g2023) & (intr_i) & (g2330)) + ((g2022) & (!g123) & (!nmi_i) & (g2023) & (!intr_i) & (!g2330)) + ((g2022) & (!g123) & (!nmi_i) & (g2023) & (!intr_i) & (g2330)) + ((g2022) & (!g123) & (!nmi_i) & (g2023) & (intr_i) & (!g2330)) + ((g2022) & (!g123) & (!nmi_i) & (g2023) & (intr_i) & (g2330)) + ((g2022) & (!g123) & (nmi_i) & (!g2023) & (!intr_i) & (!g2330)) + ((g2022) & (!g123) & (nmi_i) & (!g2023) & (!intr_i) & (g2330)) + ((g2022) & (!g123) & (nmi_i) & (!g2023) & (intr_i) & (!g2330)) + ((g2022) & (!g123) & (nmi_i) & (!g2023) & (intr_i) & (g2330)) + ((g2022) & (!g123) & (nmi_i) & (g2023) & (!intr_i) & (!g2330)) + ((g2022) & (!g123) & (nmi_i) & (g2023) & (!intr_i) & (g2330)) + ((g2022) & (!g123) & (nmi_i) & (g2023) & (intr_i) & (!g2330)) + ((g2022) & (!g123) & (nmi_i) & (g2023) & (intr_i) & (g2330)));
	assign g2409 = (((!g496) & (!sk[118]) & (!g541) & (!g453) & (g2331)) + ((!g496) & (!sk[118]) & (!g541) & (g453) & (!g2331)) + ((!g496) & (!sk[118]) & (!g541) & (g453) & (g2331)) + ((!g496) & (!sk[118]) & (g541) & (!g453) & (!g2331)) + ((!g496) & (!sk[118]) & (g541) & (!g453) & (g2331)) + ((!g496) & (!sk[118]) & (g541) & (g453) & (!g2331)) + ((!g496) & (!sk[118]) & (g541) & (g453) & (g2331)) + ((!g496) & (sk[118]) & (g541) & (g453) & (g2331)) + ((g496) & (!sk[118]) & (!g541) & (!g453) & (g2331)) + ((g496) & (!sk[118]) & (!g541) & (g453) & (!g2331)) + ((g496) & (!sk[118]) & (!g541) & (g453) & (g2331)) + ((g496) & (!sk[118]) & (g541) & (!g453) & (!g2331)) + ((g496) & (!sk[118]) & (g541) & (!g453) & (g2331)) + ((g496) & (!sk[118]) & (g541) & (g453) & (!g2331)) + ((g496) & (!sk[118]) & (g541) & (g453) & (g2331)));
	assign g2410 = (((!g587) & (sk[119]) & (g2409)) + ((g587) & (!sk[119]) & (!g2409)) + ((g587) & (!sk[119]) & (g2409)) + ((g587) & (sk[119]) & (!g2409)));
	assign g2411 = (((!g85) & (!sk[120]) & (!g541) & (g2385)) + ((!g85) & (!sk[120]) & (g541) & (!g2385)) + ((!g85) & (!sk[120]) & (g541) & (g2385)) + ((!g85) & (sk[120]) & (g541) & (g2385)) + ((g85) & (!sk[120]) & (!g541) & (g2385)) + ((g85) & (!sk[120]) & (g541) & (!g2385)) + ((g85) & (!sk[120]) & (g541) & (g2385)) + ((g85) & (sk[120]) & (!g541) & (g2385)) + ((g85) & (sk[120]) & (g541) & (!g2385)) + ((g85) & (sk[120]) & (g541) & (g2385)));
	assign g2412 = (((!g92) & (!sk[121]) & (!g2033) & (!g2034) & (g587) & (!g2411)) + ((!g92) & (!sk[121]) & (!g2033) & (!g2034) & (g587) & (g2411)) + ((!g92) & (!sk[121]) & (!g2033) & (g2034) & (!g587) & (!g2411)) + ((!g92) & (!sk[121]) & (!g2033) & (g2034) & (!g587) & (g2411)) + ((!g92) & (!sk[121]) & (!g2033) & (g2034) & (g587) & (!g2411)) + ((!g92) & (!sk[121]) & (!g2033) & (g2034) & (g587) & (g2411)) + ((!g92) & (!sk[121]) & (g2033) & (!g2034) & (!g587) & (!g2411)) + ((!g92) & (!sk[121]) & (g2033) & (!g2034) & (!g587) & (g2411)) + ((!g92) & (!sk[121]) & (g2033) & (!g2034) & (g587) & (!g2411)) + ((!g92) & (!sk[121]) & (g2033) & (!g2034) & (g587) & (g2411)) + ((!g92) & (!sk[121]) & (g2033) & (g2034) & (!g587) & (!g2411)) + ((!g92) & (!sk[121]) & (g2033) & (g2034) & (!g587) & (g2411)) + ((!g92) & (!sk[121]) & (g2033) & (g2034) & (g587) & (!g2411)) + ((!g92) & (!sk[121]) & (g2033) & (g2034) & (g587) & (g2411)) + ((!g92) & (sk[121]) & (g2033) & (!g2034) & (!g587) & (g2411)) + ((!g92) & (sk[121]) & (g2033) & (!g2034) & (g587) & (!g2411)) + ((!g92) & (sk[121]) & (g2033) & (g2034) & (!g587) & (!g2411)) + ((!g92) & (sk[121]) & (g2033) & (g2034) & (!g587) & (g2411)) + ((!g92) & (sk[121]) & (g2033) & (g2034) & (g587) & (!g2411)) + ((!g92) & (sk[121]) & (g2033) & (g2034) & (g587) & (g2411)) + ((g92) & (!sk[121]) & (!g2033) & (!g2034) & (g587) & (!g2411)) + ((g92) & (!sk[121]) & (!g2033) & (!g2034) & (g587) & (g2411)) + ((g92) & (!sk[121]) & (!g2033) & (g2034) & (!g587) & (!g2411)) + ((g92) & (!sk[121]) & (!g2033) & (g2034) & (!g587) & (g2411)) + ((g92) & (!sk[121]) & (!g2033) & (g2034) & (g587) & (!g2411)) + ((g92) & (!sk[121]) & (!g2033) & (g2034) & (g587) & (g2411)) + ((g92) & (!sk[121]) & (g2033) & (!g2034) & (!g587) & (!g2411)) + ((g92) & (!sk[121]) & (g2033) & (!g2034) & (!g587) & (g2411)) + ((g92) & (!sk[121]) & (g2033) & (!g2034) & (g587) & (!g2411)) + ((g92) & (!sk[121]) & (g2033) & (!g2034) & (g587) & (g2411)) + ((g92) & (!sk[121]) & (g2033) & (g2034) & (!g587) & (!g2411)) + ((g92) & (!sk[121]) & (g2033) & (g2034) & (!g587) & (g2411)) + ((g92) & (!sk[121]) & (g2033) & (g2034) & (g587) & (!g2411)) + ((g92) & (!sk[121]) & (g2033) & (g2034) & (g587) & (g2411)) + ((g92) & (sk[121]) & (g2033) & (!g2034) & (!g587) & (!g2411)) + ((g92) & (sk[121]) & (g2033) & (!g2034) & (g587) & (g2411)) + ((g92) & (sk[121]) & (g2033) & (g2034) & (!g587) & (!g2411)) + ((g92) & (sk[121]) & (g2033) & (g2034) & (!g587) & (g2411)) + ((g92) & (sk[121]) & (g2033) & (g2034) & (g587) & (!g2411)) + ((g92) & (sk[121]) & (g2033) & (g2034) & (g587) & (g2411)));
	assign g5034 = (((!g2921) & (!g3073) & (!sk[122]) & (g2413)) + ((!g2921) & (!g3073) & (sk[122]) & (g2413)) + ((!g2921) & (g3073) & (!sk[122]) & (!g2413)) + ((!g2921) & (g3073) & (!sk[122]) & (g2413)) + ((!g2921) & (g3073) & (sk[122]) & (g2413)) + ((g2921) & (!g3073) & (!sk[122]) & (g2413)) + ((g2921) & (g3073) & (!sk[122]) & (!g2413)) + ((g2921) & (g3073) & (!sk[122]) & (g2413)) + ((g2921) & (g3073) & (sk[122]) & (!g2413)) + ((g2921) & (g3073) & (sk[122]) & (g2413)));
	assign g2414 = (((!sk[123]) & (!g1733) & (!g2033) & (!g2034) & (g2413)) + ((!sk[123]) & (!g1733) & (!g2033) & (g2034) & (!g2413)) + ((!sk[123]) & (!g1733) & (!g2033) & (g2034) & (g2413)) + ((!sk[123]) & (!g1733) & (g2033) & (!g2034) & (!g2413)) + ((!sk[123]) & (!g1733) & (g2033) & (!g2034) & (g2413)) + ((!sk[123]) & (!g1733) & (g2033) & (g2034) & (!g2413)) + ((!sk[123]) & (!g1733) & (g2033) & (g2034) & (g2413)) + ((!sk[123]) & (g1733) & (!g2033) & (!g2034) & (g2413)) + ((!sk[123]) & (g1733) & (!g2033) & (g2034) & (!g2413)) + ((!sk[123]) & (g1733) & (!g2033) & (g2034) & (g2413)) + ((!sk[123]) & (g1733) & (g2033) & (!g2034) & (!g2413)) + ((!sk[123]) & (g1733) & (g2033) & (!g2034) & (g2413)) + ((!sk[123]) & (g1733) & (g2033) & (g2034) & (!g2413)) + ((!sk[123]) & (g1733) & (g2033) & (g2034) & (g2413)) + ((sk[123]) & (!g1733) & (!g2033) & (!g2034) & (g2413)) + ((sk[123]) & (g1733) & (!g2033) & (!g2034) & (g2413)) + ((sk[123]) & (g1733) & (!g2033) & (g2034) & (!g2413)) + ((sk[123]) & (g1733) & (!g2033) & (g2034) & (g2413)) + ((sk[123]) & (g1733) & (g2033) & (g2034) & (!g2413)) + ((sk[123]) & (g1733) & (g2033) & (g2034) & (g2413)));
	assign g2415 = (((!g2329) & (!g2029) & (g2408) & (!g2410) & (!g2412) & (!g2414)) + ((!g2329) & (!g2029) & (g2408) & (!g2410) & (!g2412) & (g2414)) + ((!g2329) & (!g2029) & (g2408) & (!g2410) & (g2412) & (!g2414)) + ((!g2329) & (!g2029) & (g2408) & (!g2410) & (g2412) & (g2414)) + ((!g2329) & (!g2029) & (g2408) & (g2410) & (!g2412) & (!g2414)) + ((!g2329) & (!g2029) & (g2408) & (g2410) & (!g2412) & (g2414)) + ((!g2329) & (!g2029) & (g2408) & (g2410) & (g2412) & (!g2414)) + ((!g2329) & (!g2029) & (g2408) & (g2410) & (g2412) & (g2414)) + ((!g2329) & (g2029) & (g2408) & (!g2410) & (!g2412) & (!g2414)) + ((!g2329) & (g2029) & (g2408) & (!g2410) & (!g2412) & (g2414)) + ((!g2329) & (g2029) & (g2408) & (!g2410) & (g2412) & (!g2414)) + ((!g2329) & (g2029) & (g2408) & (!g2410) & (g2412) & (g2414)) + ((!g2329) & (g2029) & (g2408) & (g2410) & (!g2412) & (!g2414)) + ((!g2329) & (g2029) & (g2408) & (g2410) & (!g2412) & (g2414)) + ((!g2329) & (g2029) & (g2408) & (g2410) & (g2412) & (!g2414)) + ((!g2329) & (g2029) & (g2408) & (g2410) & (g2412) & (g2414)) + ((g2329) & (!g2029) & (g2408) & (!g2410) & (!g2412) & (g2414)) + ((g2329) & (!g2029) & (g2408) & (!g2410) & (g2412) & (!g2414)) + ((g2329) & (!g2029) & (g2408) & (!g2410) & (g2412) & (g2414)) + ((g2329) & (!g2029) & (g2408) & (g2410) & (!g2412) & (g2414)) + ((g2329) & (!g2029) & (g2408) & (g2410) & (g2412) & (!g2414)) + ((g2329) & (!g2029) & (g2408) & (g2410) & (g2412) & (g2414)) + ((g2329) & (g2029) & (g2408) & (g2410) & (!g2412) & (!g2414)) + ((g2329) & (g2029) & (g2408) & (g2410) & (!g2412) & (g2414)) + ((g2329) & (g2029) & (g2408) & (g2410) & (g2412) & (!g2414)) + ((g2329) & (g2029) & (g2408) & (g2410) & (g2412) & (g2414)));
	assign g2416 = (((g2131) & (g2132) & (!dmem_dat_ix26x) & (!g2128) & (g2129) & (dmem_dat_ix10x)) + ((g2131) & (g2132) & (dmem_dat_ix26x) & (!g2128) & (!g2129) & (!dmem_dat_ix10x)) + ((g2131) & (g2132) & (dmem_dat_ix26x) & (!g2128) & (!g2129) & (dmem_dat_ix10x)) + ((g2131) & (g2132) & (dmem_dat_ix26x) & (!g2128) & (g2129) & (dmem_dat_ix10x)));
	assign g2417 = (((!g2363) & (!g2131) & (!g2132) & (!sk[126]) & (dmem_dat_ix10x) & (!g2338)) + ((!g2363) & (!g2131) & (!g2132) & (!sk[126]) & (dmem_dat_ix10x) & (g2338)) + ((!g2363) & (!g2131) & (g2132) & (!sk[126]) & (!dmem_dat_ix10x) & (!g2338)) + ((!g2363) & (!g2131) & (g2132) & (!sk[126]) & (!dmem_dat_ix10x) & (g2338)) + ((!g2363) & (!g2131) & (g2132) & (!sk[126]) & (dmem_dat_ix10x) & (!g2338)) + ((!g2363) & (!g2131) & (g2132) & (!sk[126]) & (dmem_dat_ix10x) & (g2338)) + ((!g2363) & (g2131) & (!g2132) & (!sk[126]) & (!dmem_dat_ix10x) & (!g2338)) + ((!g2363) & (g2131) & (!g2132) & (!sk[126]) & (!dmem_dat_ix10x) & (g2338)) + ((!g2363) & (g2131) & (!g2132) & (!sk[126]) & (dmem_dat_ix10x) & (!g2338)) + ((!g2363) & (g2131) & (!g2132) & (!sk[126]) & (dmem_dat_ix10x) & (g2338)) + ((!g2363) & (g2131) & (!g2132) & (sk[126]) & (dmem_dat_ix10x) & (!g2338)) + ((!g2363) & (g2131) & (!g2132) & (sk[126]) & (dmem_dat_ix10x) & (g2338)) + ((!g2363) & (g2131) & (g2132) & (!sk[126]) & (!dmem_dat_ix10x) & (!g2338)) + ((!g2363) & (g2131) & (g2132) & (!sk[126]) & (!dmem_dat_ix10x) & (g2338)) + ((!g2363) & (g2131) & (g2132) & (!sk[126]) & (dmem_dat_ix10x) & (!g2338)) + ((!g2363) & (g2131) & (g2132) & (!sk[126]) & (dmem_dat_ix10x) & (g2338)) + ((g2363) & (!g2131) & (!g2132) & (!sk[126]) & (dmem_dat_ix10x) & (!g2338)) + ((g2363) & (!g2131) & (!g2132) & (!sk[126]) & (dmem_dat_ix10x) & (g2338)) + ((g2363) & (!g2131) & (!g2132) & (sk[126]) & (!dmem_dat_ix10x) & (g2338)) + ((g2363) & (!g2131) & (!g2132) & (sk[126]) & (dmem_dat_ix10x) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (!sk[126]) & (!dmem_dat_ix10x) & (!g2338)) + ((g2363) & (!g2131) & (g2132) & (!sk[126]) & (!dmem_dat_ix10x) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (!sk[126]) & (dmem_dat_ix10x) & (!g2338)) + ((g2363) & (!g2131) & (g2132) & (!sk[126]) & (dmem_dat_ix10x) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (sk[126]) & (!dmem_dat_ix10x) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (sk[126]) & (dmem_dat_ix10x) & (g2338)) + ((g2363) & (g2131) & (!g2132) & (!sk[126]) & (!dmem_dat_ix10x) & (!g2338)) + ((g2363) & (g2131) & (!g2132) & (!sk[126]) & (!dmem_dat_ix10x) & (g2338)) + ((g2363) & (g2131) & (!g2132) & (!sk[126]) & (dmem_dat_ix10x) & (!g2338)) + ((g2363) & (g2131) & (!g2132) & (!sk[126]) & (dmem_dat_ix10x) & (g2338)) + ((g2363) & (g2131) & (!g2132) & (sk[126]) & (dmem_dat_ix10x) & (!g2338)) + ((g2363) & (g2131) & (!g2132) & (sk[126]) & (dmem_dat_ix10x) & (g2338)) + ((g2363) & (g2131) & (g2132) & (!sk[126]) & (!dmem_dat_ix10x) & (!g2338)) + ((g2363) & (g2131) & (g2132) & (!sk[126]) & (!dmem_dat_ix10x) & (g2338)) + ((g2363) & (g2131) & (g2132) & (!sk[126]) & (dmem_dat_ix10x) & (!g2338)) + ((g2363) & (g2131) & (g2132) & (!sk[126]) & (dmem_dat_ix10x) & (g2338)));
	assign g2419 = (((!sk[127]) & (!g2109) & (!g2110) & (!g2391) & (g2392) & (!g2418)) + ((!sk[127]) & (!g2109) & (!g2110) & (!g2391) & (g2392) & (g2418)) + ((!sk[127]) & (!g2109) & (!g2110) & (g2391) & (!g2392) & (!g2418)) + ((!sk[127]) & (!g2109) & (!g2110) & (g2391) & (!g2392) & (g2418)) + ((!sk[127]) & (!g2109) & (!g2110) & (g2391) & (g2392) & (!g2418)) + ((!sk[127]) & (!g2109) & (!g2110) & (g2391) & (g2392) & (g2418)) + ((!sk[127]) & (!g2109) & (g2110) & (!g2391) & (!g2392) & (!g2418)) + ((!sk[127]) & (!g2109) & (g2110) & (!g2391) & (!g2392) & (g2418)) + ((!sk[127]) & (!g2109) & (g2110) & (!g2391) & (g2392) & (!g2418)) + ((!sk[127]) & (!g2109) & (g2110) & (!g2391) & (g2392) & (g2418)) + ((!sk[127]) & (!g2109) & (g2110) & (g2391) & (!g2392) & (!g2418)) + ((!sk[127]) & (!g2109) & (g2110) & (g2391) & (!g2392) & (g2418)) + ((!sk[127]) & (!g2109) & (g2110) & (g2391) & (g2392) & (!g2418)) + ((!sk[127]) & (!g2109) & (g2110) & (g2391) & (g2392) & (g2418)) + ((!sk[127]) & (g2109) & (!g2110) & (!g2391) & (g2392) & (!g2418)) + ((!sk[127]) & (g2109) & (!g2110) & (!g2391) & (g2392) & (g2418)) + ((!sk[127]) & (g2109) & (!g2110) & (g2391) & (!g2392) & (!g2418)) + ((!sk[127]) & (g2109) & (!g2110) & (g2391) & (!g2392) & (g2418)) + ((!sk[127]) & (g2109) & (!g2110) & (g2391) & (g2392) & (!g2418)) + ((!sk[127]) & (g2109) & (!g2110) & (g2391) & (g2392) & (g2418)) + ((!sk[127]) & (g2109) & (g2110) & (!g2391) & (!g2392) & (!g2418)) + ((!sk[127]) & (g2109) & (g2110) & (!g2391) & (!g2392) & (g2418)) + ((!sk[127]) & (g2109) & (g2110) & (!g2391) & (g2392) & (!g2418)) + ((!sk[127]) & (g2109) & (g2110) & (!g2391) & (g2392) & (g2418)) + ((!sk[127]) & (g2109) & (g2110) & (g2391) & (!g2392) & (!g2418)) + ((!sk[127]) & (g2109) & (g2110) & (g2391) & (!g2392) & (g2418)) + ((!sk[127]) & (g2109) & (g2110) & (g2391) & (g2392) & (!g2418)) + ((!sk[127]) & (g2109) & (g2110) & (g2391) & (g2392) & (g2418)) + ((sk[127]) & (!g2109) & (!g2110) & (!g2391) & (!g2392) & (g2418)) + ((sk[127]) & (!g2109) & (!g2110) & (!g2391) & (g2392) & (g2418)) + ((sk[127]) & (!g2109) & (!g2110) & (g2391) & (!g2392) & (g2418)) + ((sk[127]) & (!g2109) & (!g2110) & (g2391) & (g2392) & (!g2418)) + ((sk[127]) & (!g2109) & (g2110) & (!g2391) & (!g2392) & (!g2418)) + ((sk[127]) & (!g2109) & (g2110) & (!g2391) & (g2392) & (!g2418)) + ((sk[127]) & (!g2109) & (g2110) & (g2391) & (!g2392) & (!g2418)) + ((sk[127]) & (!g2109) & (g2110) & (g2391) & (g2392) & (g2418)) + ((sk[127]) & (g2109) & (!g2110) & (!g2391) & (!g2392) & (g2418)) + ((sk[127]) & (g2109) & (!g2110) & (!g2391) & (g2392) & (!g2418)) + ((sk[127]) & (g2109) & (!g2110) & (g2391) & (!g2392) & (!g2418)) + ((sk[127]) & (g2109) & (!g2110) & (g2391) & (g2392) & (!g2418)) + ((sk[127]) & (g2109) & (g2110) & (!g2391) & (!g2392) & (!g2418)) + ((sk[127]) & (g2109) & (g2110) & (!g2391) & (g2392) & (g2418)) + ((sk[127]) & (g2109) & (g2110) & (g2391) & (!g2392) & (g2418)) + ((sk[127]) & (g2109) & (g2110) & (g2391) & (g2392) & (g2418)));
	assign g2420 = (((!g2341) & (!sk[0]) & (!g2342) & (!g2367) & (g2393)) + ((!g2341) & (!sk[0]) & (!g2342) & (g2367) & (!g2393)) + ((!g2341) & (!sk[0]) & (!g2342) & (g2367) & (g2393)) + ((!g2341) & (!sk[0]) & (g2342) & (!g2367) & (!g2393)) + ((!g2341) & (!sk[0]) & (g2342) & (!g2367) & (g2393)) + ((!g2341) & (!sk[0]) & (g2342) & (g2367) & (!g2393)) + ((!g2341) & (!sk[0]) & (g2342) & (g2367) & (g2393)) + ((g2341) & (!sk[0]) & (!g2342) & (!g2367) & (g2393)) + ((g2341) & (!sk[0]) & (!g2342) & (g2367) & (!g2393)) + ((g2341) & (!sk[0]) & (!g2342) & (g2367) & (g2393)) + ((g2341) & (!sk[0]) & (g2342) & (!g2367) & (!g2393)) + ((g2341) & (!sk[0]) & (g2342) & (!g2367) & (g2393)) + ((g2341) & (!sk[0]) & (g2342) & (g2367) & (!g2393)) + ((g2341) & (!sk[0]) & (g2342) & (g2367) & (g2393)) + ((g2341) & (sk[0]) & (g2342) & (g2367) & (g2393)));
	assign g2421 = (((!g2395) & (!sk[1]) & (!g2396) & (g2397)) + ((!g2395) & (!sk[1]) & (g2396) & (!g2397)) + ((!g2395) & (!sk[1]) & (g2396) & (g2397)) + ((!g2395) & (sk[1]) & (!g2396) & (g2397)) + ((!g2395) & (sk[1]) & (g2396) & (!g2397)) + ((!g2395) & (sk[1]) & (g2396) & (g2397)) + ((g2395) & (!sk[1]) & (!g2396) & (g2397)) + ((g2395) & (!sk[1]) & (g2396) & (!g2397)) + ((g2395) & (!sk[1]) & (g2396) & (g2397)) + ((g2395) & (sk[1]) & (g2396) & (g2397)));
	assign g2422 = (((g2109) & (!sk[2]) & (!g2391)) + ((g2109) & (!sk[2]) & (g2391)) + ((g2109) & (sk[2]) & (!g2391)));
	assign g2423 = (((!sk[3]) & (g2110) & (!g2418)) + ((!sk[3]) & (g2110) & (g2418)) + ((sk[3]) & (!g2110) & (!g2418)) + ((sk[3]) & (g2110) & (g2418)));
	assign g2424 = (((!g2421) & (!sk[4]) & (!g2422) & (g2423)) + ((!g2421) & (!sk[4]) & (g2422) & (!g2423)) + ((!g2421) & (!sk[4]) & (g2422) & (g2423)) + ((!g2421) & (sk[4]) & (!g2422) & (g2423)) + ((!g2421) & (sk[4]) & (g2422) & (!g2423)) + ((g2421) & (!sk[4]) & (!g2422) & (g2423)) + ((g2421) & (!sk[4]) & (g2422) & (!g2423)) + ((g2421) & (!sk[4]) & (g2422) & (g2423)) + ((g2421) & (sk[4]) & (!g2422) & (!g2423)) + ((g2421) & (sk[4]) & (g2422) & (g2423)));
	assign g2425 = (((!g2076) & (!g2077) & (!g2192) & (!sk[5]) & (g2216) & (!g2218)) + ((!g2076) & (!g2077) & (!g2192) & (!sk[5]) & (g2216) & (g2218)) + ((!g2076) & (!g2077) & (!g2192) & (sk[5]) & (g2216) & (!g2218)) + ((!g2076) & (!g2077) & (!g2192) & (sk[5]) & (g2216) & (g2218)) + ((!g2076) & (!g2077) & (g2192) & (!sk[5]) & (!g2216) & (!g2218)) + ((!g2076) & (!g2077) & (g2192) & (!sk[5]) & (!g2216) & (g2218)) + ((!g2076) & (!g2077) & (g2192) & (!sk[5]) & (g2216) & (!g2218)) + ((!g2076) & (!g2077) & (g2192) & (!sk[5]) & (g2216) & (g2218)) + ((!g2076) & (!g2077) & (g2192) & (sk[5]) & (g2216) & (!g2218)) + ((!g2076) & (!g2077) & (g2192) & (sk[5]) & (g2216) & (g2218)) + ((!g2076) & (g2077) & (!g2192) & (!sk[5]) & (!g2216) & (!g2218)) + ((!g2076) & (g2077) & (!g2192) & (!sk[5]) & (!g2216) & (g2218)) + ((!g2076) & (g2077) & (!g2192) & (!sk[5]) & (g2216) & (!g2218)) + ((!g2076) & (g2077) & (!g2192) & (!sk[5]) & (g2216) & (g2218)) + ((!g2076) & (g2077) & (!g2192) & (sk[5]) & (!g2216) & (g2218)) + ((!g2076) & (g2077) & (!g2192) & (sk[5]) & (g2216) & (g2218)) + ((!g2076) & (g2077) & (g2192) & (!sk[5]) & (!g2216) & (!g2218)) + ((!g2076) & (g2077) & (g2192) & (!sk[5]) & (!g2216) & (g2218)) + ((!g2076) & (g2077) & (g2192) & (!sk[5]) & (g2216) & (!g2218)) + ((!g2076) & (g2077) & (g2192) & (!sk[5]) & (g2216) & (g2218)) + ((!g2076) & (g2077) & (g2192) & (sk[5]) & (!g2216) & (g2218)) + ((!g2076) & (g2077) & (g2192) & (sk[5]) & (g2216) & (g2218)) + ((g2076) & (!g2077) & (!g2192) & (!sk[5]) & (g2216) & (!g2218)) + ((g2076) & (!g2077) & (!g2192) & (!sk[5]) & (g2216) & (g2218)) + ((g2076) & (!g2077) & (g2192) & (!sk[5]) & (!g2216) & (!g2218)) + ((g2076) & (!g2077) & (g2192) & (!sk[5]) & (!g2216) & (g2218)) + ((g2076) & (!g2077) & (g2192) & (!sk[5]) & (g2216) & (!g2218)) + ((g2076) & (!g2077) & (g2192) & (!sk[5]) & (g2216) & (g2218)) + ((g2076) & (!g2077) & (g2192) & (sk[5]) & (!g2216) & (!g2218)) + ((g2076) & (!g2077) & (g2192) & (sk[5]) & (!g2216) & (g2218)) + ((g2076) & (!g2077) & (g2192) & (sk[5]) & (g2216) & (!g2218)) + ((g2076) & (!g2077) & (g2192) & (sk[5]) & (g2216) & (g2218)) + ((g2076) & (g2077) & (!g2192) & (!sk[5]) & (!g2216) & (!g2218)) + ((g2076) & (g2077) & (!g2192) & (!sk[5]) & (!g2216) & (g2218)) + ((g2076) & (g2077) & (!g2192) & (!sk[5]) & (g2216) & (!g2218)) + ((g2076) & (g2077) & (!g2192) & (!sk[5]) & (g2216) & (g2218)) + ((g2076) & (g2077) & (g2192) & (!sk[5]) & (!g2216) & (!g2218)) + ((g2076) & (g2077) & (g2192) & (!sk[5]) & (!g2216) & (g2218)) + ((g2076) & (g2077) & (g2192) & (!sk[5]) & (g2216) & (!g2218)) + ((g2076) & (g2077) & (g2192) & (!sk[5]) & (g2216) & (g2218)) + ((g2076) & (g2077) & (g2192) & (sk[5]) & (!g2216) & (!g2218)) + ((g2076) & (g2077) & (g2192) & (sk[5]) & (!g2216) & (g2218)) + ((g2076) & (g2077) & (g2192) & (sk[5]) & (g2216) & (!g2218)) + ((g2076) & (g2077) & (g2192) & (sk[5]) & (g2216) & (g2218)));
	assign g2426 = (((!g2110) & (!g2109) & (!g2108) & (g2116) & (g2071) & (g2074)) + ((!g2110) & (!g2109) & (g2108) & (!g2116) & (!g2071) & (g2074)) + ((!g2110) & (!g2109) & (g2108) & (g2116) & (!g2071) & (g2074)) + ((!g2110) & (!g2109) & (g2108) & (g2116) & (g2071) & (g2074)) + ((!g2110) & (g2109) & (!g2108) & (!g2116) & (g2071) & (!g2074)) + ((!g2110) & (g2109) & (!g2108) & (g2116) & (g2071) & (!g2074)) + ((!g2110) & (g2109) & (!g2108) & (g2116) & (g2071) & (g2074)) + ((!g2110) & (g2109) & (g2108) & (!g2116) & (!g2071) & (g2074)) + ((!g2110) & (g2109) & (g2108) & (!g2116) & (g2071) & (!g2074)) + ((!g2110) & (g2109) & (g2108) & (g2116) & (!g2071) & (g2074)) + ((!g2110) & (g2109) & (g2108) & (g2116) & (g2071) & (!g2074)) + ((!g2110) & (g2109) & (g2108) & (g2116) & (g2071) & (g2074)) + ((g2110) & (!g2109) & (!g2108) & (!g2116) & (!g2071) & (!g2074)) + ((g2110) & (!g2109) & (!g2108) & (g2116) & (!g2071) & (!g2074)) + ((g2110) & (!g2109) & (!g2108) & (g2116) & (g2071) & (g2074)) + ((g2110) & (!g2109) & (g2108) & (!g2116) & (!g2071) & (!g2074)) + ((g2110) & (!g2109) & (g2108) & (!g2116) & (!g2071) & (g2074)) + ((g2110) & (!g2109) & (g2108) & (g2116) & (!g2071) & (!g2074)) + ((g2110) & (!g2109) & (g2108) & (g2116) & (!g2071) & (g2074)) + ((g2110) & (!g2109) & (g2108) & (g2116) & (g2071) & (g2074)) + ((g2110) & (g2109) & (!g2108) & (!g2116) & (!g2071) & (!g2074)) + ((g2110) & (g2109) & (!g2108) & (!g2116) & (g2071) & (!g2074)) + ((g2110) & (g2109) & (!g2108) & (g2116) & (!g2071) & (!g2074)) + ((g2110) & (g2109) & (!g2108) & (g2116) & (g2071) & (!g2074)) + ((g2110) & (g2109) & (!g2108) & (g2116) & (g2071) & (g2074)) + ((g2110) & (g2109) & (g2108) & (!g2116) & (!g2071) & (!g2074)) + ((g2110) & (g2109) & (g2108) & (!g2116) & (!g2071) & (g2074)) + ((g2110) & (g2109) & (g2108) & (!g2116) & (g2071) & (!g2074)) + ((g2110) & (g2109) & (g2108) & (g2116) & (!g2071) & (!g2074)) + ((g2110) & (g2109) & (g2108) & (g2116) & (!g2071) & (g2074)) + ((g2110) & (g2109) & (g2108) & (g2116) & (g2071) & (!g2074)) + ((g2110) & (g2109) & (g2108) & (g2116) & (g2071) & (g2074)));
	assign g2427 = (((!sk[7]) & (!g2076) & (!g2077) & (!g2211) & (g2320) & (!g2426)) + ((!sk[7]) & (!g2076) & (!g2077) & (!g2211) & (g2320) & (g2426)) + ((!sk[7]) & (!g2076) & (!g2077) & (g2211) & (!g2320) & (!g2426)) + ((!sk[7]) & (!g2076) & (!g2077) & (g2211) & (!g2320) & (g2426)) + ((!sk[7]) & (!g2076) & (!g2077) & (g2211) & (g2320) & (!g2426)) + ((!sk[7]) & (!g2076) & (!g2077) & (g2211) & (g2320) & (g2426)) + ((!sk[7]) & (!g2076) & (g2077) & (!g2211) & (!g2320) & (!g2426)) + ((!sk[7]) & (!g2076) & (g2077) & (!g2211) & (!g2320) & (g2426)) + ((!sk[7]) & (!g2076) & (g2077) & (!g2211) & (g2320) & (!g2426)) + ((!sk[7]) & (!g2076) & (g2077) & (!g2211) & (g2320) & (g2426)) + ((!sk[7]) & (!g2076) & (g2077) & (g2211) & (!g2320) & (!g2426)) + ((!sk[7]) & (!g2076) & (g2077) & (g2211) & (!g2320) & (g2426)) + ((!sk[7]) & (!g2076) & (g2077) & (g2211) & (g2320) & (!g2426)) + ((!sk[7]) & (!g2076) & (g2077) & (g2211) & (g2320) & (g2426)) + ((!sk[7]) & (g2076) & (!g2077) & (!g2211) & (g2320) & (!g2426)) + ((!sk[7]) & (g2076) & (!g2077) & (!g2211) & (g2320) & (g2426)) + ((!sk[7]) & (g2076) & (!g2077) & (g2211) & (!g2320) & (!g2426)) + ((!sk[7]) & (g2076) & (!g2077) & (g2211) & (!g2320) & (g2426)) + ((!sk[7]) & (g2076) & (!g2077) & (g2211) & (g2320) & (!g2426)) + ((!sk[7]) & (g2076) & (!g2077) & (g2211) & (g2320) & (g2426)) + ((!sk[7]) & (g2076) & (g2077) & (!g2211) & (!g2320) & (!g2426)) + ((!sk[7]) & (g2076) & (g2077) & (!g2211) & (!g2320) & (g2426)) + ((!sk[7]) & (g2076) & (g2077) & (!g2211) & (g2320) & (!g2426)) + ((!sk[7]) & (g2076) & (g2077) & (!g2211) & (g2320) & (g2426)) + ((!sk[7]) & (g2076) & (g2077) & (g2211) & (!g2320) & (!g2426)) + ((!sk[7]) & (g2076) & (g2077) & (g2211) & (!g2320) & (g2426)) + ((!sk[7]) & (g2076) & (g2077) & (g2211) & (g2320) & (!g2426)) + ((!sk[7]) & (g2076) & (g2077) & (g2211) & (g2320) & (g2426)) + ((sk[7]) & (!g2076) & (!g2077) & (!g2211) & (!g2320) & (g2426)) + ((sk[7]) & (!g2076) & (!g2077) & (!g2211) & (g2320) & (g2426)) + ((sk[7]) & (!g2076) & (!g2077) & (g2211) & (!g2320) & (g2426)) + ((sk[7]) & (!g2076) & (!g2077) & (g2211) & (g2320) & (g2426)) + ((sk[7]) & (!g2076) & (g2077) & (!g2211) & (g2320) & (!g2426)) + ((sk[7]) & (!g2076) & (g2077) & (!g2211) & (g2320) & (g2426)) + ((sk[7]) & (!g2076) & (g2077) & (g2211) & (g2320) & (!g2426)) + ((sk[7]) & (!g2076) & (g2077) & (g2211) & (g2320) & (g2426)) + ((sk[7]) & (g2076) & (!g2077) & (g2211) & (!g2320) & (!g2426)) + ((sk[7]) & (g2076) & (!g2077) & (g2211) & (!g2320) & (g2426)) + ((sk[7]) & (g2076) & (!g2077) & (g2211) & (g2320) & (!g2426)) + ((sk[7]) & (g2076) & (!g2077) & (g2211) & (g2320) & (g2426)));
	assign g2428 = (((!g2222) & (!g2215) & (!g2223) & (g2217) & (g2076) & (g2077)) + ((!g2222) & (!g2215) & (g2223) & (!g2217) & (!g2076) & (g2077)) + ((!g2222) & (!g2215) & (g2223) & (g2217) & (!g2076) & (g2077)) + ((!g2222) & (!g2215) & (g2223) & (g2217) & (g2076) & (g2077)) + ((!g2222) & (g2215) & (!g2223) & (!g2217) & (g2076) & (!g2077)) + ((!g2222) & (g2215) & (!g2223) & (g2217) & (g2076) & (!g2077)) + ((!g2222) & (g2215) & (!g2223) & (g2217) & (g2076) & (g2077)) + ((!g2222) & (g2215) & (g2223) & (!g2217) & (!g2076) & (g2077)) + ((!g2222) & (g2215) & (g2223) & (!g2217) & (g2076) & (!g2077)) + ((!g2222) & (g2215) & (g2223) & (g2217) & (!g2076) & (g2077)) + ((!g2222) & (g2215) & (g2223) & (g2217) & (g2076) & (!g2077)) + ((!g2222) & (g2215) & (g2223) & (g2217) & (g2076) & (g2077)) + ((g2222) & (!g2215) & (!g2223) & (!g2217) & (!g2076) & (!g2077)) + ((g2222) & (!g2215) & (!g2223) & (g2217) & (!g2076) & (!g2077)) + ((g2222) & (!g2215) & (!g2223) & (g2217) & (g2076) & (g2077)) + ((g2222) & (!g2215) & (g2223) & (!g2217) & (!g2076) & (!g2077)) + ((g2222) & (!g2215) & (g2223) & (!g2217) & (!g2076) & (g2077)) + ((g2222) & (!g2215) & (g2223) & (g2217) & (!g2076) & (!g2077)) + ((g2222) & (!g2215) & (g2223) & (g2217) & (!g2076) & (g2077)) + ((g2222) & (!g2215) & (g2223) & (g2217) & (g2076) & (g2077)) + ((g2222) & (g2215) & (!g2223) & (!g2217) & (!g2076) & (!g2077)) + ((g2222) & (g2215) & (!g2223) & (!g2217) & (g2076) & (!g2077)) + ((g2222) & (g2215) & (!g2223) & (g2217) & (!g2076) & (!g2077)) + ((g2222) & (g2215) & (!g2223) & (g2217) & (g2076) & (!g2077)) + ((g2222) & (g2215) & (!g2223) & (g2217) & (g2076) & (g2077)) + ((g2222) & (g2215) & (g2223) & (!g2217) & (!g2076) & (!g2077)) + ((g2222) & (g2215) & (g2223) & (!g2217) & (!g2076) & (g2077)) + ((g2222) & (g2215) & (g2223) & (!g2217) & (g2076) & (!g2077)) + ((g2222) & (g2215) & (g2223) & (g2217) & (!g2076) & (!g2077)) + ((g2222) & (g2215) & (g2223) & (g2217) & (!g2076) & (g2077)) + ((g2222) & (g2215) & (g2223) & (g2217) & (g2076) & (!g2077)) + ((g2222) & (g2215) & (g2223) & (g2217) & (g2076) & (g2077)));
	assign g2429 = (((!g2399) & (!g2400) & (!g2425) & (g2427) & (!sk[9]) & (!g2428)) + ((!g2399) & (!g2400) & (!g2425) & (g2427) & (!sk[9]) & (g2428)) + ((!g2399) & (!g2400) & (!g2425) & (g2427) & (sk[9]) & (!g2428)) + ((!g2399) & (!g2400) & (!g2425) & (g2427) & (sk[9]) & (g2428)) + ((!g2399) & (!g2400) & (g2425) & (!g2427) & (!sk[9]) & (!g2428)) + ((!g2399) & (!g2400) & (g2425) & (!g2427) & (!sk[9]) & (g2428)) + ((!g2399) & (!g2400) & (g2425) & (g2427) & (!sk[9]) & (!g2428)) + ((!g2399) & (!g2400) & (g2425) & (g2427) & (!sk[9]) & (g2428)) + ((!g2399) & (!g2400) & (g2425) & (g2427) & (sk[9]) & (!g2428)) + ((!g2399) & (!g2400) & (g2425) & (g2427) & (sk[9]) & (g2428)) + ((!g2399) & (g2400) & (!g2425) & (!g2427) & (!sk[9]) & (!g2428)) + ((!g2399) & (g2400) & (!g2425) & (!g2427) & (!sk[9]) & (g2428)) + ((!g2399) & (g2400) & (!g2425) & (g2427) & (!sk[9]) & (!g2428)) + ((!g2399) & (g2400) & (!g2425) & (g2427) & (!sk[9]) & (g2428)) + ((!g2399) & (g2400) & (g2425) & (!g2427) & (!sk[9]) & (!g2428)) + ((!g2399) & (g2400) & (g2425) & (!g2427) & (!sk[9]) & (g2428)) + ((!g2399) & (g2400) & (g2425) & (!g2427) & (sk[9]) & (!g2428)) + ((!g2399) & (g2400) & (g2425) & (!g2427) & (sk[9]) & (g2428)) + ((!g2399) & (g2400) & (g2425) & (g2427) & (!sk[9]) & (!g2428)) + ((!g2399) & (g2400) & (g2425) & (g2427) & (!sk[9]) & (g2428)) + ((!g2399) & (g2400) & (g2425) & (g2427) & (sk[9]) & (!g2428)) + ((!g2399) & (g2400) & (g2425) & (g2427) & (sk[9]) & (g2428)) + ((g2399) & (!g2400) & (!g2425) & (!g2427) & (sk[9]) & (g2428)) + ((g2399) & (!g2400) & (!g2425) & (g2427) & (!sk[9]) & (!g2428)) + ((g2399) & (!g2400) & (!g2425) & (g2427) & (!sk[9]) & (g2428)) + ((g2399) & (!g2400) & (!g2425) & (g2427) & (sk[9]) & (g2428)) + ((g2399) & (!g2400) & (g2425) & (!g2427) & (!sk[9]) & (!g2428)) + ((g2399) & (!g2400) & (g2425) & (!g2427) & (!sk[9]) & (g2428)) + ((g2399) & (!g2400) & (g2425) & (!g2427) & (sk[9]) & (g2428)) + ((g2399) & (!g2400) & (g2425) & (g2427) & (!sk[9]) & (!g2428)) + ((g2399) & (!g2400) & (g2425) & (g2427) & (!sk[9]) & (g2428)) + ((g2399) & (!g2400) & (g2425) & (g2427) & (sk[9]) & (g2428)) + ((g2399) & (g2400) & (!g2425) & (!g2427) & (!sk[9]) & (!g2428)) + ((g2399) & (g2400) & (!g2425) & (!g2427) & (!sk[9]) & (g2428)) + ((g2399) & (g2400) & (!g2425) & (g2427) & (!sk[9]) & (!g2428)) + ((g2399) & (g2400) & (!g2425) & (g2427) & (!sk[9]) & (g2428)) + ((g2399) & (g2400) & (g2425) & (!g2427) & (!sk[9]) & (!g2428)) + ((g2399) & (g2400) & (g2425) & (!g2427) & (!sk[9]) & (g2428)) + ((g2399) & (g2400) & (g2425) & (g2427) & (!sk[9]) & (!g2428)) + ((g2399) & (g2400) & (g2425) & (g2427) & (!sk[9]) & (g2428)));
	assign g2430 = (((!g2418) & (!g2110) & (!g2124) & (!g2264) & (!g3638) & (!g2429)) + ((!g2418) & (!g2110) & (!g2124) & (!g2264) & (g3638) & (!g2429)) + ((!g2418) & (!g2110) & (!g2124) & (g2264) & (!g3638) & (!g2429)) + ((!g2418) & (!g2110) & (!g2124) & (g2264) & (!g3638) & (g2429)) + ((!g2418) & (!g2110) & (g2124) & (!g2264) & (!g3638) & (!g2429)) + ((!g2418) & (!g2110) & (g2124) & (!g2264) & (!g3638) & (g2429)) + ((!g2418) & (!g2110) & (g2124) & (!g2264) & (g3638) & (!g2429)) + ((!g2418) & (!g2110) & (g2124) & (!g2264) & (g3638) & (g2429)) + ((!g2418) & (!g2110) & (g2124) & (g2264) & (!g3638) & (!g2429)) + ((!g2418) & (!g2110) & (g2124) & (g2264) & (!g3638) & (g2429)) + ((!g2418) & (!g2110) & (g2124) & (g2264) & (g3638) & (!g2429)) + ((!g2418) & (!g2110) & (g2124) & (g2264) & (g3638) & (g2429)) + ((!g2418) & (g2110) & (!g2124) & (!g2264) & (!g3638) & (!g2429)) + ((!g2418) & (g2110) & (!g2124) & (!g2264) & (g3638) & (!g2429)) + ((!g2418) & (g2110) & (!g2124) & (g2264) & (!g3638) & (!g2429)) + ((!g2418) & (g2110) & (!g2124) & (g2264) & (!g3638) & (g2429)) + ((g2418) & (!g2110) & (!g2124) & (!g2264) & (!g3638) & (!g2429)) + ((g2418) & (!g2110) & (!g2124) & (!g2264) & (g3638) & (!g2429)) + ((g2418) & (!g2110) & (!g2124) & (g2264) & (!g3638) & (!g2429)) + ((g2418) & (!g2110) & (!g2124) & (g2264) & (!g3638) & (g2429)) + ((g2418) & (g2110) & (!g2124) & (!g2264) & (!g3638) & (!g2429)) + ((g2418) & (g2110) & (!g2124) & (!g2264) & (g3638) & (!g2429)) + ((g2418) & (g2110) & (!g2124) & (g2264) & (!g3638) & (!g2429)) + ((g2418) & (g2110) & (!g2124) & (g2264) & (!g3638) & (g2429)) + ((g2418) & (g2110) & (g2124) & (g2264) & (!g3638) & (!g2429)) + ((g2418) & (g2110) & (g2124) & (g2264) & (!g3638) & (g2429)) + ((g2418) & (g2110) & (g2124) & (g2264) & (g3638) & (!g2429)) + ((g2418) & (g2110) & (g2124) & (g2264) & (g3638) & (g2429)));
	assign g2431 = (((!g75) & (!g2110) & (!g2280) & (!g2416) & (!g2417) & (!g2430)) + ((!g75) & (!g2110) & (!g2280) & (!g2416) & (g2417) & (!g2430)) + ((!g75) & (!g2110) & (!g2280) & (g2416) & (!g2417) & (!g2430)) + ((!g75) & (!g2110) & (!g2280) & (g2416) & (g2417) & (!g2430)) + ((!g75) & (g2110) & (!g2280) & (!g2416) & (!g2417) & (!g2430)) + ((!g75) & (g2110) & (!g2280) & (!g2416) & (g2417) & (!g2430)) + ((!g75) & (g2110) & (!g2280) & (g2416) & (!g2417) & (!g2430)) + ((!g75) & (g2110) & (!g2280) & (g2416) & (g2417) & (!g2430)) + ((!g75) & (g2110) & (g2280) & (!g2416) & (!g2417) & (!g2430)) + ((!g75) & (g2110) & (g2280) & (!g2416) & (!g2417) & (g2430)) + ((!g75) & (g2110) & (g2280) & (!g2416) & (g2417) & (!g2430)) + ((!g75) & (g2110) & (g2280) & (!g2416) & (g2417) & (g2430)) + ((!g75) & (g2110) & (g2280) & (g2416) & (!g2417) & (!g2430)) + ((!g75) & (g2110) & (g2280) & (g2416) & (!g2417) & (g2430)) + ((!g75) & (g2110) & (g2280) & (g2416) & (g2417) & (!g2430)) + ((!g75) & (g2110) & (g2280) & (g2416) & (g2417) & (g2430)) + ((g75) & (!g2110) & (!g2280) & (!g2416) & (g2417) & (!g2430)) + ((g75) & (!g2110) & (!g2280) & (!g2416) & (g2417) & (g2430)) + ((g75) & (!g2110) & (!g2280) & (g2416) & (!g2417) & (!g2430)) + ((g75) & (!g2110) & (!g2280) & (g2416) & (!g2417) & (g2430)) + ((g75) & (!g2110) & (!g2280) & (g2416) & (g2417) & (!g2430)) + ((g75) & (!g2110) & (!g2280) & (g2416) & (g2417) & (g2430)) + ((g75) & (!g2110) & (g2280) & (!g2416) & (g2417) & (!g2430)) + ((g75) & (!g2110) & (g2280) & (!g2416) & (g2417) & (g2430)) + ((g75) & (!g2110) & (g2280) & (g2416) & (!g2417) & (!g2430)) + ((g75) & (!g2110) & (g2280) & (g2416) & (!g2417) & (g2430)) + ((g75) & (!g2110) & (g2280) & (g2416) & (g2417) & (!g2430)) + ((g75) & (!g2110) & (g2280) & (g2416) & (g2417) & (g2430)) + ((g75) & (g2110) & (!g2280) & (!g2416) & (g2417) & (!g2430)) + ((g75) & (g2110) & (!g2280) & (!g2416) & (g2417) & (g2430)) + ((g75) & (g2110) & (!g2280) & (g2416) & (!g2417) & (!g2430)) + ((g75) & (g2110) & (!g2280) & (g2416) & (!g2417) & (g2430)) + ((g75) & (g2110) & (!g2280) & (g2416) & (g2417) & (!g2430)) + ((g75) & (g2110) & (!g2280) & (g2416) & (g2417) & (g2430)) + ((g75) & (g2110) & (g2280) & (!g2416) & (g2417) & (!g2430)) + ((g75) & (g2110) & (g2280) & (!g2416) & (g2417) & (g2430)) + ((g75) & (g2110) & (g2280) & (g2416) & (!g2417) & (!g2430)) + ((g75) & (g2110) & (g2280) & (g2416) & (!g2417) & (g2430)) + ((g75) & (g2110) & (g2280) & (g2416) & (g2417) & (!g2430)) + ((g75) & (g2110) & (g2280) & (g2416) & (g2417) & (g2430)));
	assign g5035 = (((!g2921) & (!sk[12]) & (!g3075) & (g2432)) + ((!g2921) & (!sk[12]) & (g3075) & (!g2432)) + ((!g2921) & (!sk[12]) & (g3075) & (g2432)) + ((!g2921) & (sk[12]) & (!g3075) & (g2432)) + ((!g2921) & (sk[12]) & (g3075) & (g2432)) + ((g2921) & (!sk[12]) & (!g3075) & (g2432)) + ((g2921) & (!sk[12]) & (g3075) & (!g2432)) + ((g2921) & (!sk[12]) & (g3075) & (g2432)) + ((g2921) & (sk[12]) & (g3075) & (!g2432)) + ((g2921) & (sk[12]) & (g3075) & (g2432)));
	assign g2433 = (((!g92) & (!sk[13]) & (!g587) & (g2411)) + ((!g92) & (!sk[13]) & (g587) & (!g2411)) + ((!g92) & (!sk[13]) & (g587) & (g2411)) + ((!g92) & (sk[13]) & (g587) & (g2411)) + ((g92) & (!sk[13]) & (!g587) & (g2411)) + ((g92) & (!sk[13]) & (g587) & (!g2411)) + ((g92) & (!sk[13]) & (g587) & (g2411)) + ((g92) & (sk[13]) & (!g587) & (g2411)) + ((g92) & (sk[13]) & (g587) & (!g2411)) + ((g92) & (sk[13]) & (g587) & (g2411)));
	assign g2434 = (((!sk[14]) & (!g91) & (!g630) & (g2433)) + ((!sk[14]) & (!g91) & (g630) & (!g2433)) + ((!sk[14]) & (!g91) & (g630) & (g2433)) + ((!sk[14]) & (g91) & (!g630) & (g2433)) + ((!sk[14]) & (g91) & (g630) & (!g2433)) + ((!sk[14]) & (g91) & (g630) & (g2433)) + ((sk[14]) & (!g91) & (!g630) & (g2433)) + ((sk[14]) & (!g91) & (g630) & (!g2433)) + ((sk[14]) & (g91) & (!g630) & (!g2433)) + ((sk[14]) & (g91) & (g630) & (g2433)));
	assign g2435 = (((!g1746) & (!g2033) & (!g2034) & (g2432) & (!sk[15]) & (!g2434)) + ((!g1746) & (!g2033) & (!g2034) & (g2432) & (!sk[15]) & (g2434)) + ((!g1746) & (!g2033) & (!g2034) & (g2432) & (sk[15]) & (!g2434)) + ((!g1746) & (!g2033) & (!g2034) & (g2432) & (sk[15]) & (g2434)) + ((!g1746) & (!g2033) & (g2034) & (!g2432) & (!sk[15]) & (!g2434)) + ((!g1746) & (!g2033) & (g2034) & (!g2432) & (!sk[15]) & (g2434)) + ((!g1746) & (!g2033) & (g2034) & (g2432) & (!sk[15]) & (!g2434)) + ((!g1746) & (!g2033) & (g2034) & (g2432) & (!sk[15]) & (g2434)) + ((!g1746) & (g2033) & (!g2034) & (!g2432) & (!sk[15]) & (!g2434)) + ((!g1746) & (g2033) & (!g2034) & (!g2432) & (!sk[15]) & (g2434)) + ((!g1746) & (g2033) & (!g2034) & (!g2432) & (sk[15]) & (g2434)) + ((!g1746) & (g2033) & (!g2034) & (g2432) & (!sk[15]) & (!g2434)) + ((!g1746) & (g2033) & (!g2034) & (g2432) & (!sk[15]) & (g2434)) + ((!g1746) & (g2033) & (!g2034) & (g2432) & (sk[15]) & (g2434)) + ((!g1746) & (g2033) & (g2034) & (!g2432) & (!sk[15]) & (!g2434)) + ((!g1746) & (g2033) & (g2034) & (!g2432) & (!sk[15]) & (g2434)) + ((!g1746) & (g2033) & (g2034) & (g2432) & (!sk[15]) & (!g2434)) + ((!g1746) & (g2033) & (g2034) & (g2432) & (!sk[15]) & (g2434)) + ((g1746) & (!g2033) & (!g2034) & (g2432) & (!sk[15]) & (!g2434)) + ((g1746) & (!g2033) & (!g2034) & (g2432) & (!sk[15]) & (g2434)) + ((g1746) & (!g2033) & (!g2034) & (g2432) & (sk[15]) & (!g2434)) + ((g1746) & (!g2033) & (!g2034) & (g2432) & (sk[15]) & (g2434)) + ((g1746) & (!g2033) & (g2034) & (!g2432) & (!sk[15]) & (!g2434)) + ((g1746) & (!g2033) & (g2034) & (!g2432) & (!sk[15]) & (g2434)) + ((g1746) & (!g2033) & (g2034) & (!g2432) & (sk[15]) & (!g2434)) + ((g1746) & (!g2033) & (g2034) & (!g2432) & (sk[15]) & (g2434)) + ((g1746) & (!g2033) & (g2034) & (g2432) & (!sk[15]) & (!g2434)) + ((g1746) & (!g2033) & (g2034) & (g2432) & (!sk[15]) & (g2434)) + ((g1746) & (!g2033) & (g2034) & (g2432) & (sk[15]) & (!g2434)) + ((g1746) & (!g2033) & (g2034) & (g2432) & (sk[15]) & (g2434)) + ((g1746) & (g2033) & (!g2034) & (!g2432) & (!sk[15]) & (!g2434)) + ((g1746) & (g2033) & (!g2034) & (!g2432) & (!sk[15]) & (g2434)) + ((g1746) & (g2033) & (!g2034) & (!g2432) & (sk[15]) & (g2434)) + ((g1746) & (g2033) & (!g2034) & (g2432) & (!sk[15]) & (!g2434)) + ((g1746) & (g2033) & (!g2034) & (g2432) & (!sk[15]) & (g2434)) + ((g1746) & (g2033) & (!g2034) & (g2432) & (sk[15]) & (g2434)) + ((g1746) & (g2033) & (g2034) & (!g2432) & (!sk[15]) & (!g2434)) + ((g1746) & (g2033) & (g2034) & (!g2432) & (!sk[15]) & (g2434)) + ((g1746) & (g2033) & (g2034) & (g2432) & (!sk[15]) & (!g2434)) + ((g1746) & (g2033) & (g2034) & (g2432) & (!sk[15]) & (g2434)));
	assign g2436 = (((!sk[16]) & (!g630) & (!g587) & (g2409)) + ((!sk[16]) & (!g630) & (g587) & (!g2409)) + ((!sk[16]) & (!g630) & (g587) & (g2409)) + ((!sk[16]) & (g630) & (!g587) & (g2409)) + ((!sk[16]) & (g630) & (g587) & (!g2409)) + ((!sk[16]) & (g630) & (g587) & (g2409)) + ((sk[16]) & (!g630) & (g587) & (g2409)) + ((sk[16]) & (g630) & (!g587) & (!g2409)) + ((sk[16]) & (g630) & (!g587) & (g2409)) + ((sk[16]) & (g630) & (g587) & (!g2409)));
	assign g2437 = (((g2131) & (g2132) & (!dmem_dat_ix27x) & (!g2128) & (g2129) & (dmem_dat_ix11x)) + ((g2131) & (g2132) & (dmem_dat_ix27x) & (!g2128) & (!g2129) & (!dmem_dat_ix11x)) + ((g2131) & (g2132) & (dmem_dat_ix27x) & (!g2128) & (!g2129) & (dmem_dat_ix11x)) + ((g2131) & (g2132) & (dmem_dat_ix27x) & (!g2128) & (g2129) & (dmem_dat_ix11x)));
	assign g2438 = (((!sk[18]) & (!g2363) & (!g2131) & (!g2132) & (dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (!g2363) & (!g2131) & (!g2132) & (dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (!g2363) & (!g2131) & (g2132) & (!dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (!g2363) & (!g2131) & (g2132) & (!dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (!g2363) & (!g2131) & (g2132) & (dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (!g2363) & (!g2131) & (g2132) & (dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (!g2363) & (g2131) & (!g2132) & (!dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (!g2363) & (g2131) & (!g2132) & (!dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (!g2363) & (g2131) & (!g2132) & (dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (!g2363) & (g2131) & (!g2132) & (dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (!g2363) & (g2131) & (g2132) & (!dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (!g2363) & (g2131) & (g2132) & (!dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (!g2363) & (g2131) & (g2132) & (dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (!g2363) & (g2131) & (g2132) & (dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (g2363) & (!g2131) & (!g2132) & (dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (g2363) & (!g2131) & (!g2132) & (dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (g2363) & (!g2131) & (g2132) & (!dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (g2363) & (!g2131) & (g2132) & (!dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (g2363) & (!g2131) & (g2132) & (dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (g2363) & (!g2131) & (g2132) & (dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (g2363) & (g2131) & (!g2132) & (!dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (g2363) & (g2131) & (!g2132) & (!dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (g2363) & (g2131) & (!g2132) & (dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (g2363) & (g2131) & (!g2132) & (dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (g2363) & (g2131) & (g2132) & (!dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (g2363) & (g2131) & (g2132) & (!dmem_dat_ix11x) & (g2338)) + ((!sk[18]) & (g2363) & (g2131) & (g2132) & (dmem_dat_ix11x) & (!g2338)) + ((!sk[18]) & (g2363) & (g2131) & (g2132) & (dmem_dat_ix11x) & (g2338)) + ((sk[18]) & (!g2363) & (g2131) & (!g2132) & (dmem_dat_ix11x) & (!g2338)) + ((sk[18]) & (!g2363) & (g2131) & (!g2132) & (dmem_dat_ix11x) & (g2338)) + ((sk[18]) & (g2363) & (!g2131) & (!g2132) & (!dmem_dat_ix11x) & (g2338)) + ((sk[18]) & (g2363) & (!g2131) & (!g2132) & (dmem_dat_ix11x) & (g2338)) + ((sk[18]) & (g2363) & (!g2131) & (g2132) & (!dmem_dat_ix11x) & (g2338)) + ((sk[18]) & (g2363) & (!g2131) & (g2132) & (dmem_dat_ix11x) & (g2338)) + ((sk[18]) & (g2363) & (g2131) & (!g2132) & (dmem_dat_ix11x) & (!g2338)) + ((sk[18]) & (g2363) & (g2131) & (!g2132) & (dmem_dat_ix11x) & (g2338)));
	assign g2440 = (((!sk[19]) & (g2110) & (!g2418)) + ((!sk[19]) & (g2110) & (g2418)) + ((sk[19]) & (!g2110) & (g2418)) + ((sk[19]) & (g2110) & (!g2418)));
	assign g2441 = (((!g2109) & (!g2108) & (g2365) & (g2366) & (g2391) & (g2440)) + ((!g2109) & (g2108) & (!g2365) & (g2366) & (g2391) & (g2440)) + ((!g2109) & (g2108) & (g2365) & (!g2366) & (g2391) & (g2440)) + ((!g2109) & (g2108) & (g2365) & (g2366) & (g2391) & (g2440)) + ((g2109) & (!g2108) & (!g2365) & (!g2366) & (g2391) & (g2440)) + ((g2109) & (!g2108) & (!g2365) & (g2366) & (g2391) & (g2440)) + ((g2109) & (!g2108) & (g2365) & (!g2366) & (g2391) & (g2440)) + ((g2109) & (!g2108) & (g2365) & (g2366) & (!g2391) & (g2440)) + ((g2109) & (!g2108) & (g2365) & (g2366) & (g2391) & (g2440)) + ((g2109) & (g2108) & (!g2365) & (!g2366) & (g2391) & (g2440)) + ((g2109) & (g2108) & (!g2365) & (g2366) & (!g2391) & (g2440)) + ((g2109) & (g2108) & (!g2365) & (g2366) & (g2391) & (g2440)) + ((g2109) & (g2108) & (g2365) & (!g2366) & (!g2391) & (g2440)) + ((g2109) & (g2108) & (g2365) & (!g2366) & (g2391) & (g2440)) + ((g2109) & (g2108) & (g2365) & (g2366) & (!g2391) & (g2440)) + ((g2109) & (g2108) & (g2365) & (g2366) & (g2391) & (g2440)));
	assign g2442 = (((g2110) & (!sk[21]) & (!g2418)) + ((g2110) & (!sk[21]) & (g2418)) + ((g2110) & (sk[21]) & (g2418)));
	assign g2443 = (((!g2111) & (!g2439) & (!g2441) & (!sk[22]) & (g2442)) + ((!g2111) & (!g2439) & (!g2441) & (sk[22]) & (g2442)) + ((!g2111) & (!g2439) & (g2441) & (!sk[22]) & (!g2442)) + ((!g2111) & (!g2439) & (g2441) & (!sk[22]) & (g2442)) + ((!g2111) & (!g2439) & (g2441) & (sk[22]) & (!g2442)) + ((!g2111) & (!g2439) & (g2441) & (sk[22]) & (g2442)) + ((!g2111) & (g2439) & (!g2441) & (!sk[22]) & (!g2442)) + ((!g2111) & (g2439) & (!g2441) & (!sk[22]) & (g2442)) + ((!g2111) & (g2439) & (!g2441) & (sk[22]) & (!g2442)) + ((!g2111) & (g2439) & (g2441) & (!sk[22]) & (!g2442)) + ((!g2111) & (g2439) & (g2441) & (!sk[22]) & (g2442)) + ((g2111) & (!g2439) & (!g2441) & (!sk[22]) & (g2442)) + ((g2111) & (!g2439) & (!g2441) & (sk[22]) & (!g2442)) + ((g2111) & (!g2439) & (g2441) & (!sk[22]) & (!g2442)) + ((g2111) & (!g2439) & (g2441) & (!sk[22]) & (g2442)) + ((g2111) & (g2439) & (!g2441) & (!sk[22]) & (!g2442)) + ((g2111) & (g2439) & (!g2441) & (!sk[22]) & (g2442)) + ((g2111) & (g2439) & (!g2441) & (sk[22]) & (g2442)) + ((g2111) & (g2439) & (g2441) & (!sk[22]) & (!g2442)) + ((g2111) & (g2439) & (g2441) & (!sk[22]) & (g2442)) + ((g2111) & (g2439) & (g2441) & (sk[22]) & (!g2442)) + ((g2111) & (g2439) & (g2441) & (sk[22]) & (g2442)));
	assign g2444 = (((!sk[23]) & (g2110) & (!g2418)) + ((!sk[23]) & (g2110) & (g2418)) + ((sk[23]) & (g2110) & (!g2418)));
	assign g2445 = (((!sk[24]) & (g2111) & (!g2439)) + ((!sk[24]) & (g2111) & (g2439)) + ((sk[24]) & (!g2111) & (!g2439)) + ((sk[24]) & (g2111) & (g2439)));
	assign g2446 = (((!g2421) & (!g2422) & (!g2423) & (!g2444) & (sk[25]) & (g2445)) + ((!g2421) & (!g2422) & (!g2423) & (g2444) & (!sk[25]) & (!g2445)) + ((!g2421) & (!g2422) & (!g2423) & (g2444) & (!sk[25]) & (g2445)) + ((!g2421) & (!g2422) & (!g2423) & (g2444) & (sk[25]) & (!g2445)) + ((!g2421) & (!g2422) & (g2423) & (!g2444) & (!sk[25]) & (!g2445)) + ((!g2421) & (!g2422) & (g2423) & (!g2444) & (!sk[25]) & (g2445)) + ((!g2421) & (!g2422) & (g2423) & (!g2444) & (sk[25]) & (g2445)) + ((!g2421) & (!g2422) & (g2423) & (g2444) & (!sk[25]) & (!g2445)) + ((!g2421) & (!g2422) & (g2423) & (g2444) & (!sk[25]) & (g2445)) + ((!g2421) & (!g2422) & (g2423) & (g2444) & (sk[25]) & (!g2445)) + ((!g2421) & (g2422) & (!g2423) & (!g2444) & (!sk[25]) & (!g2445)) + ((!g2421) & (g2422) & (!g2423) & (!g2444) & (!sk[25]) & (g2445)) + ((!g2421) & (g2422) & (!g2423) & (!g2444) & (sk[25]) & (g2445)) + ((!g2421) & (g2422) & (!g2423) & (g2444) & (!sk[25]) & (!g2445)) + ((!g2421) & (g2422) & (!g2423) & (g2444) & (!sk[25]) & (g2445)) + ((!g2421) & (g2422) & (!g2423) & (g2444) & (sk[25]) & (!g2445)) + ((!g2421) & (g2422) & (g2423) & (!g2444) & (!sk[25]) & (!g2445)) + ((!g2421) & (g2422) & (g2423) & (!g2444) & (!sk[25]) & (g2445)) + ((!g2421) & (g2422) & (g2423) & (!g2444) & (sk[25]) & (!g2445)) + ((!g2421) & (g2422) & (g2423) & (g2444) & (!sk[25]) & (!g2445)) + ((!g2421) & (g2422) & (g2423) & (g2444) & (!sk[25]) & (g2445)) + ((!g2421) & (g2422) & (g2423) & (g2444) & (sk[25]) & (g2445)) + ((g2421) & (!g2422) & (!g2423) & (!g2444) & (sk[25]) & (g2445)) + ((g2421) & (!g2422) & (!g2423) & (g2444) & (!sk[25]) & (!g2445)) + ((g2421) & (!g2422) & (!g2423) & (g2444) & (!sk[25]) & (g2445)) + ((g2421) & (!g2422) & (!g2423) & (g2444) & (sk[25]) & (!g2445)) + ((g2421) & (!g2422) & (g2423) & (!g2444) & (!sk[25]) & (!g2445)) + ((g2421) & (!g2422) & (g2423) & (!g2444) & (!sk[25]) & (g2445)) + ((g2421) & (!g2422) & (g2423) & (!g2444) & (sk[25]) & (!g2445)) + ((g2421) & (!g2422) & (g2423) & (g2444) & (!sk[25]) & (!g2445)) + ((g2421) & (!g2422) & (g2423) & (g2444) & (!sk[25]) & (g2445)) + ((g2421) & (!g2422) & (g2423) & (g2444) & (sk[25]) & (g2445)) + ((g2421) & (g2422) & (!g2423) & (!g2444) & (!sk[25]) & (!g2445)) + ((g2421) & (g2422) & (!g2423) & (!g2444) & (!sk[25]) & (g2445)) + ((g2421) & (g2422) & (!g2423) & (!g2444) & (sk[25]) & (!g2445)) + ((g2421) & (g2422) & (!g2423) & (g2444) & (!sk[25]) & (!g2445)) + ((g2421) & (g2422) & (!g2423) & (g2444) & (!sk[25]) & (g2445)) + ((g2421) & (g2422) & (!g2423) & (g2444) & (sk[25]) & (g2445)) + ((g2421) & (g2422) & (g2423) & (!g2444) & (!sk[25]) & (!g2445)) + ((g2421) & (g2422) & (g2423) & (!g2444) & (!sk[25]) & (g2445)) + ((g2421) & (g2422) & (g2423) & (!g2444) & (sk[25]) & (!g2445)) + ((g2421) & (g2422) & (g2423) & (g2444) & (!sk[25]) & (!g2445)) + ((g2421) & (g2422) & (g2423) & (g2444) & (!sk[25]) & (g2445)) + ((g2421) & (g2422) & (g2423) & (g2444) & (sk[25]) & (g2445)));
	assign g2447 = (((g2111) & (!sk[26]) & (!g2439)) + ((g2111) & (!sk[26]) & (g2439)) + ((g2111) & (sk[26]) & (g2439)));
	assign g2448 = (((!g2076) & (!g2077) & (!sk[27]) & (!g2192) & (g2243) & (!g2245)) + ((!g2076) & (!g2077) & (!sk[27]) & (!g2192) & (g2243) & (g2245)) + ((!g2076) & (!g2077) & (!sk[27]) & (g2192) & (!g2243) & (!g2245)) + ((!g2076) & (!g2077) & (!sk[27]) & (g2192) & (!g2243) & (g2245)) + ((!g2076) & (!g2077) & (!sk[27]) & (g2192) & (g2243) & (!g2245)) + ((!g2076) & (!g2077) & (!sk[27]) & (g2192) & (g2243) & (g2245)) + ((!g2076) & (!g2077) & (sk[27]) & (!g2192) & (g2243) & (!g2245)) + ((!g2076) & (!g2077) & (sk[27]) & (!g2192) & (g2243) & (g2245)) + ((!g2076) & (!g2077) & (sk[27]) & (g2192) & (g2243) & (!g2245)) + ((!g2076) & (!g2077) & (sk[27]) & (g2192) & (g2243) & (g2245)) + ((!g2076) & (g2077) & (!sk[27]) & (!g2192) & (!g2243) & (!g2245)) + ((!g2076) & (g2077) & (!sk[27]) & (!g2192) & (!g2243) & (g2245)) + ((!g2076) & (g2077) & (!sk[27]) & (!g2192) & (g2243) & (!g2245)) + ((!g2076) & (g2077) & (!sk[27]) & (!g2192) & (g2243) & (g2245)) + ((!g2076) & (g2077) & (!sk[27]) & (g2192) & (!g2243) & (!g2245)) + ((!g2076) & (g2077) & (!sk[27]) & (g2192) & (!g2243) & (g2245)) + ((!g2076) & (g2077) & (!sk[27]) & (g2192) & (g2243) & (!g2245)) + ((!g2076) & (g2077) & (!sk[27]) & (g2192) & (g2243) & (g2245)) + ((!g2076) & (g2077) & (sk[27]) & (!g2192) & (!g2243) & (g2245)) + ((!g2076) & (g2077) & (sk[27]) & (!g2192) & (g2243) & (g2245)) + ((!g2076) & (g2077) & (sk[27]) & (g2192) & (!g2243) & (g2245)) + ((!g2076) & (g2077) & (sk[27]) & (g2192) & (g2243) & (g2245)) + ((g2076) & (!g2077) & (!sk[27]) & (!g2192) & (g2243) & (!g2245)) + ((g2076) & (!g2077) & (!sk[27]) & (!g2192) & (g2243) & (g2245)) + ((g2076) & (!g2077) & (!sk[27]) & (g2192) & (!g2243) & (!g2245)) + ((g2076) & (!g2077) & (!sk[27]) & (g2192) & (!g2243) & (g2245)) + ((g2076) & (!g2077) & (!sk[27]) & (g2192) & (g2243) & (!g2245)) + ((g2076) & (!g2077) & (!sk[27]) & (g2192) & (g2243) & (g2245)) + ((g2076) & (!g2077) & (sk[27]) & (g2192) & (!g2243) & (!g2245)) + ((g2076) & (!g2077) & (sk[27]) & (g2192) & (!g2243) & (g2245)) + ((g2076) & (!g2077) & (sk[27]) & (g2192) & (g2243) & (!g2245)) + ((g2076) & (!g2077) & (sk[27]) & (g2192) & (g2243) & (g2245)) + ((g2076) & (g2077) & (!sk[27]) & (!g2192) & (!g2243) & (!g2245)) + ((g2076) & (g2077) & (!sk[27]) & (!g2192) & (!g2243) & (g2245)) + ((g2076) & (g2077) & (!sk[27]) & (!g2192) & (g2243) & (!g2245)) + ((g2076) & (g2077) & (!sk[27]) & (!g2192) & (g2243) & (g2245)) + ((g2076) & (g2077) & (!sk[27]) & (g2192) & (!g2243) & (!g2245)) + ((g2076) & (g2077) & (!sk[27]) & (g2192) & (!g2243) & (g2245)) + ((g2076) & (g2077) & (!sk[27]) & (g2192) & (g2243) & (!g2245)) + ((g2076) & (g2077) & (!sk[27]) & (g2192) & (g2243) & (g2245)) + ((g2076) & (g2077) & (sk[27]) & (g2192) & (!g2243) & (!g2245)) + ((g2076) & (g2077) & (sk[27]) & (g2192) & (!g2243) & (g2245)) + ((g2076) & (g2077) & (sk[27]) & (g2192) & (g2243) & (!g2245)) + ((g2076) & (g2077) & (sk[27]) & (g2192) & (g2243) & (g2245)));
	assign g2449 = (((!g2111) & (!g2110) & (!g2109) & (g2108) & (g2071) & (g2074)) + ((!g2111) & (!g2110) & (g2109) & (!g2108) & (!g2071) & (g2074)) + ((!g2111) & (!g2110) & (g2109) & (g2108) & (!g2071) & (g2074)) + ((!g2111) & (!g2110) & (g2109) & (g2108) & (g2071) & (g2074)) + ((!g2111) & (g2110) & (!g2109) & (!g2108) & (g2071) & (!g2074)) + ((!g2111) & (g2110) & (!g2109) & (g2108) & (g2071) & (!g2074)) + ((!g2111) & (g2110) & (!g2109) & (g2108) & (g2071) & (g2074)) + ((!g2111) & (g2110) & (g2109) & (!g2108) & (!g2071) & (g2074)) + ((!g2111) & (g2110) & (g2109) & (!g2108) & (g2071) & (!g2074)) + ((!g2111) & (g2110) & (g2109) & (g2108) & (!g2071) & (g2074)) + ((!g2111) & (g2110) & (g2109) & (g2108) & (g2071) & (!g2074)) + ((!g2111) & (g2110) & (g2109) & (g2108) & (g2071) & (g2074)) + ((g2111) & (!g2110) & (!g2109) & (!g2108) & (!g2071) & (!g2074)) + ((g2111) & (!g2110) & (!g2109) & (g2108) & (!g2071) & (!g2074)) + ((g2111) & (!g2110) & (!g2109) & (g2108) & (g2071) & (g2074)) + ((g2111) & (!g2110) & (g2109) & (!g2108) & (!g2071) & (!g2074)) + ((g2111) & (!g2110) & (g2109) & (!g2108) & (!g2071) & (g2074)) + ((g2111) & (!g2110) & (g2109) & (g2108) & (!g2071) & (!g2074)) + ((g2111) & (!g2110) & (g2109) & (g2108) & (!g2071) & (g2074)) + ((g2111) & (!g2110) & (g2109) & (g2108) & (g2071) & (g2074)) + ((g2111) & (g2110) & (!g2109) & (!g2108) & (!g2071) & (!g2074)) + ((g2111) & (g2110) & (!g2109) & (!g2108) & (g2071) & (!g2074)) + ((g2111) & (g2110) & (!g2109) & (g2108) & (!g2071) & (!g2074)) + ((g2111) & (g2110) & (!g2109) & (g2108) & (g2071) & (!g2074)) + ((g2111) & (g2110) & (!g2109) & (g2108) & (g2071) & (g2074)) + ((g2111) & (g2110) & (g2109) & (!g2108) & (!g2071) & (!g2074)) + ((g2111) & (g2110) & (g2109) & (!g2108) & (!g2071) & (g2074)) + ((g2111) & (g2110) & (g2109) & (!g2108) & (g2071) & (!g2074)) + ((g2111) & (g2110) & (g2109) & (g2108) & (!g2071) & (!g2074)) + ((g2111) & (g2110) & (g2109) & (g2108) & (!g2071) & (g2074)) + ((g2111) & (g2110) & (g2109) & (g2108) & (g2071) & (!g2074)) + ((g2111) & (g2110) & (g2109) & (g2108) & (g2071) & (g2074)));
	assign g2450 = (((!g2076) & (!g2077) & (!sk[29]) & (!g2236) & (g2350) & (!g2449)) + ((!g2076) & (!g2077) & (!sk[29]) & (!g2236) & (g2350) & (g2449)) + ((!g2076) & (!g2077) & (!sk[29]) & (g2236) & (!g2350) & (!g2449)) + ((!g2076) & (!g2077) & (!sk[29]) & (g2236) & (!g2350) & (g2449)) + ((!g2076) & (!g2077) & (!sk[29]) & (g2236) & (g2350) & (!g2449)) + ((!g2076) & (!g2077) & (!sk[29]) & (g2236) & (g2350) & (g2449)) + ((!g2076) & (!g2077) & (sk[29]) & (!g2236) & (!g2350) & (g2449)) + ((!g2076) & (!g2077) & (sk[29]) & (!g2236) & (g2350) & (g2449)) + ((!g2076) & (!g2077) & (sk[29]) & (g2236) & (!g2350) & (g2449)) + ((!g2076) & (!g2077) & (sk[29]) & (g2236) & (g2350) & (g2449)) + ((!g2076) & (g2077) & (!sk[29]) & (!g2236) & (!g2350) & (!g2449)) + ((!g2076) & (g2077) & (!sk[29]) & (!g2236) & (!g2350) & (g2449)) + ((!g2076) & (g2077) & (!sk[29]) & (!g2236) & (g2350) & (!g2449)) + ((!g2076) & (g2077) & (!sk[29]) & (!g2236) & (g2350) & (g2449)) + ((!g2076) & (g2077) & (!sk[29]) & (g2236) & (!g2350) & (!g2449)) + ((!g2076) & (g2077) & (!sk[29]) & (g2236) & (!g2350) & (g2449)) + ((!g2076) & (g2077) & (!sk[29]) & (g2236) & (g2350) & (!g2449)) + ((!g2076) & (g2077) & (!sk[29]) & (g2236) & (g2350) & (g2449)) + ((!g2076) & (g2077) & (sk[29]) & (!g2236) & (g2350) & (!g2449)) + ((!g2076) & (g2077) & (sk[29]) & (!g2236) & (g2350) & (g2449)) + ((!g2076) & (g2077) & (sk[29]) & (g2236) & (g2350) & (!g2449)) + ((!g2076) & (g2077) & (sk[29]) & (g2236) & (g2350) & (g2449)) + ((g2076) & (!g2077) & (!sk[29]) & (!g2236) & (g2350) & (!g2449)) + ((g2076) & (!g2077) & (!sk[29]) & (!g2236) & (g2350) & (g2449)) + ((g2076) & (!g2077) & (!sk[29]) & (g2236) & (!g2350) & (!g2449)) + ((g2076) & (!g2077) & (!sk[29]) & (g2236) & (!g2350) & (g2449)) + ((g2076) & (!g2077) & (!sk[29]) & (g2236) & (g2350) & (!g2449)) + ((g2076) & (!g2077) & (!sk[29]) & (g2236) & (g2350) & (g2449)) + ((g2076) & (!g2077) & (sk[29]) & (g2236) & (!g2350) & (!g2449)) + ((g2076) & (!g2077) & (sk[29]) & (g2236) & (!g2350) & (g2449)) + ((g2076) & (!g2077) & (sk[29]) & (g2236) & (g2350) & (!g2449)) + ((g2076) & (!g2077) & (sk[29]) & (g2236) & (g2350) & (g2449)) + ((g2076) & (g2077) & (!sk[29]) & (!g2236) & (!g2350) & (!g2449)) + ((g2076) & (g2077) & (!sk[29]) & (!g2236) & (!g2350) & (g2449)) + ((g2076) & (g2077) & (!sk[29]) & (!g2236) & (g2350) & (!g2449)) + ((g2076) & (g2077) & (!sk[29]) & (!g2236) & (g2350) & (g2449)) + ((g2076) & (g2077) & (!sk[29]) & (g2236) & (!g2350) & (!g2449)) + ((g2076) & (g2077) & (!sk[29]) & (g2236) & (!g2350) & (g2449)) + ((g2076) & (g2077) & (!sk[29]) & (g2236) & (g2350) & (!g2449)) + ((g2076) & (g2077) & (!sk[29]) & (g2236) & (g2350) & (g2449)));
	assign g2451 = (((!g2249) & (!g2242) & (!g2250) & (g2244) & (g2076) & (g2077)) + ((!g2249) & (!g2242) & (g2250) & (!g2244) & (!g2076) & (g2077)) + ((!g2249) & (!g2242) & (g2250) & (g2244) & (!g2076) & (g2077)) + ((!g2249) & (!g2242) & (g2250) & (g2244) & (g2076) & (g2077)) + ((!g2249) & (g2242) & (!g2250) & (!g2244) & (g2076) & (!g2077)) + ((!g2249) & (g2242) & (!g2250) & (g2244) & (g2076) & (!g2077)) + ((!g2249) & (g2242) & (!g2250) & (g2244) & (g2076) & (g2077)) + ((!g2249) & (g2242) & (g2250) & (!g2244) & (!g2076) & (g2077)) + ((!g2249) & (g2242) & (g2250) & (!g2244) & (g2076) & (!g2077)) + ((!g2249) & (g2242) & (g2250) & (g2244) & (!g2076) & (g2077)) + ((!g2249) & (g2242) & (g2250) & (g2244) & (g2076) & (!g2077)) + ((!g2249) & (g2242) & (g2250) & (g2244) & (g2076) & (g2077)) + ((g2249) & (!g2242) & (!g2250) & (!g2244) & (!g2076) & (!g2077)) + ((g2249) & (!g2242) & (!g2250) & (g2244) & (!g2076) & (!g2077)) + ((g2249) & (!g2242) & (!g2250) & (g2244) & (g2076) & (g2077)) + ((g2249) & (!g2242) & (g2250) & (!g2244) & (!g2076) & (!g2077)) + ((g2249) & (!g2242) & (g2250) & (!g2244) & (!g2076) & (g2077)) + ((g2249) & (!g2242) & (g2250) & (g2244) & (!g2076) & (!g2077)) + ((g2249) & (!g2242) & (g2250) & (g2244) & (!g2076) & (g2077)) + ((g2249) & (!g2242) & (g2250) & (g2244) & (g2076) & (g2077)) + ((g2249) & (g2242) & (!g2250) & (!g2244) & (!g2076) & (!g2077)) + ((g2249) & (g2242) & (!g2250) & (!g2244) & (g2076) & (!g2077)) + ((g2249) & (g2242) & (!g2250) & (g2244) & (!g2076) & (!g2077)) + ((g2249) & (g2242) & (!g2250) & (g2244) & (g2076) & (!g2077)) + ((g2249) & (g2242) & (!g2250) & (g2244) & (g2076) & (g2077)) + ((g2249) & (g2242) & (g2250) & (!g2244) & (!g2076) & (!g2077)) + ((g2249) & (g2242) & (g2250) & (!g2244) & (!g2076) & (g2077)) + ((g2249) & (g2242) & (g2250) & (!g2244) & (g2076) & (!g2077)) + ((g2249) & (g2242) & (g2250) & (g2244) & (!g2076) & (!g2077)) + ((g2249) & (g2242) & (g2250) & (g2244) & (!g2076) & (g2077)) + ((g2249) & (g2242) & (g2250) & (g2244) & (g2076) & (!g2077)) + ((g2249) & (g2242) & (g2250) & (g2244) & (g2076) & (g2077)));
	assign g2452 = (((!sk[31]) & (!g2399) & (!g2400) & (!g2448) & (g2450) & (!g2451)) + ((!sk[31]) & (!g2399) & (!g2400) & (!g2448) & (g2450) & (g2451)) + ((!sk[31]) & (!g2399) & (!g2400) & (g2448) & (!g2450) & (!g2451)) + ((!sk[31]) & (!g2399) & (!g2400) & (g2448) & (!g2450) & (g2451)) + ((!sk[31]) & (!g2399) & (!g2400) & (g2448) & (g2450) & (!g2451)) + ((!sk[31]) & (!g2399) & (!g2400) & (g2448) & (g2450) & (g2451)) + ((!sk[31]) & (!g2399) & (g2400) & (!g2448) & (!g2450) & (!g2451)) + ((!sk[31]) & (!g2399) & (g2400) & (!g2448) & (!g2450) & (g2451)) + ((!sk[31]) & (!g2399) & (g2400) & (!g2448) & (g2450) & (!g2451)) + ((!sk[31]) & (!g2399) & (g2400) & (!g2448) & (g2450) & (g2451)) + ((!sk[31]) & (!g2399) & (g2400) & (g2448) & (!g2450) & (!g2451)) + ((!sk[31]) & (!g2399) & (g2400) & (g2448) & (!g2450) & (g2451)) + ((!sk[31]) & (!g2399) & (g2400) & (g2448) & (g2450) & (!g2451)) + ((!sk[31]) & (!g2399) & (g2400) & (g2448) & (g2450) & (g2451)) + ((!sk[31]) & (g2399) & (!g2400) & (!g2448) & (g2450) & (!g2451)) + ((!sk[31]) & (g2399) & (!g2400) & (!g2448) & (g2450) & (g2451)) + ((!sk[31]) & (g2399) & (!g2400) & (g2448) & (!g2450) & (!g2451)) + ((!sk[31]) & (g2399) & (!g2400) & (g2448) & (!g2450) & (g2451)) + ((!sk[31]) & (g2399) & (!g2400) & (g2448) & (g2450) & (!g2451)) + ((!sk[31]) & (g2399) & (!g2400) & (g2448) & (g2450) & (g2451)) + ((!sk[31]) & (g2399) & (g2400) & (!g2448) & (!g2450) & (!g2451)) + ((!sk[31]) & (g2399) & (g2400) & (!g2448) & (!g2450) & (g2451)) + ((!sk[31]) & (g2399) & (g2400) & (!g2448) & (g2450) & (!g2451)) + ((!sk[31]) & (g2399) & (g2400) & (!g2448) & (g2450) & (g2451)) + ((!sk[31]) & (g2399) & (g2400) & (g2448) & (!g2450) & (!g2451)) + ((!sk[31]) & (g2399) & (g2400) & (g2448) & (!g2450) & (g2451)) + ((!sk[31]) & (g2399) & (g2400) & (g2448) & (g2450) & (!g2451)) + ((!sk[31]) & (g2399) & (g2400) & (g2448) & (g2450) & (g2451)) + ((sk[31]) & (!g2399) & (!g2400) & (!g2448) & (g2450) & (!g2451)) + ((sk[31]) & (!g2399) & (!g2400) & (!g2448) & (g2450) & (g2451)) + ((sk[31]) & (!g2399) & (!g2400) & (g2448) & (g2450) & (!g2451)) + ((sk[31]) & (!g2399) & (!g2400) & (g2448) & (g2450) & (g2451)) + ((sk[31]) & (!g2399) & (g2400) & (g2448) & (!g2450) & (!g2451)) + ((sk[31]) & (!g2399) & (g2400) & (g2448) & (!g2450) & (g2451)) + ((sk[31]) & (!g2399) & (g2400) & (g2448) & (g2450) & (!g2451)) + ((sk[31]) & (!g2399) & (g2400) & (g2448) & (g2450) & (g2451)) + ((sk[31]) & (g2399) & (!g2400) & (!g2448) & (!g2450) & (g2451)) + ((sk[31]) & (g2399) & (!g2400) & (!g2448) & (g2450) & (g2451)) + ((sk[31]) & (g2399) & (!g2400) & (g2448) & (!g2450) & (g2451)) + ((sk[31]) & (g2399) & (!g2400) & (g2448) & (g2450) & (g2451)));
	assign g2453 = (((!g2439) & (!g2111) & (!g2124) & (!g2264) & (!g3614) & (!g2452)) + ((!g2439) & (!g2111) & (!g2124) & (!g2264) & (g3614) & (!g2452)) + ((!g2439) & (!g2111) & (!g2124) & (g2264) & (!g3614) & (!g2452)) + ((!g2439) & (!g2111) & (!g2124) & (g2264) & (!g3614) & (g2452)) + ((!g2439) & (!g2111) & (g2124) & (!g2264) & (!g3614) & (!g2452)) + ((!g2439) & (!g2111) & (g2124) & (!g2264) & (!g3614) & (g2452)) + ((!g2439) & (!g2111) & (g2124) & (!g2264) & (g3614) & (!g2452)) + ((!g2439) & (!g2111) & (g2124) & (!g2264) & (g3614) & (g2452)) + ((!g2439) & (!g2111) & (g2124) & (g2264) & (!g3614) & (!g2452)) + ((!g2439) & (!g2111) & (g2124) & (g2264) & (!g3614) & (g2452)) + ((!g2439) & (!g2111) & (g2124) & (g2264) & (g3614) & (!g2452)) + ((!g2439) & (!g2111) & (g2124) & (g2264) & (g3614) & (g2452)) + ((!g2439) & (g2111) & (!g2124) & (!g2264) & (!g3614) & (!g2452)) + ((!g2439) & (g2111) & (!g2124) & (!g2264) & (g3614) & (!g2452)) + ((!g2439) & (g2111) & (!g2124) & (g2264) & (!g3614) & (!g2452)) + ((!g2439) & (g2111) & (!g2124) & (g2264) & (!g3614) & (g2452)) + ((g2439) & (!g2111) & (!g2124) & (!g2264) & (!g3614) & (!g2452)) + ((g2439) & (!g2111) & (!g2124) & (!g2264) & (g3614) & (!g2452)) + ((g2439) & (!g2111) & (!g2124) & (g2264) & (!g3614) & (!g2452)) + ((g2439) & (!g2111) & (!g2124) & (g2264) & (!g3614) & (g2452)) + ((g2439) & (g2111) & (!g2124) & (!g2264) & (!g3614) & (!g2452)) + ((g2439) & (g2111) & (!g2124) & (!g2264) & (g3614) & (!g2452)) + ((g2439) & (g2111) & (!g2124) & (g2264) & (!g3614) & (!g2452)) + ((g2439) & (g2111) & (!g2124) & (g2264) & (!g3614) & (g2452)) + ((g2439) & (g2111) & (g2124) & (g2264) & (!g3614) & (!g2452)) + ((g2439) & (g2111) & (g2124) & (g2264) & (!g3614) & (g2452)) + ((g2439) & (g2111) & (g2124) & (g2264) & (g3614) & (!g2452)) + ((g2439) & (g2111) & (g2124) & (g2264) & (g3614) & (g2452)));
	assign g2454 = (((!g75) & (!g2111) & (!g2280) & (!g2437) & (!g2438) & (!g2453)) + ((!g75) & (!g2111) & (!g2280) & (!g2437) & (g2438) & (!g2453)) + ((!g75) & (!g2111) & (!g2280) & (g2437) & (!g2438) & (!g2453)) + ((!g75) & (!g2111) & (!g2280) & (g2437) & (g2438) & (!g2453)) + ((!g75) & (g2111) & (!g2280) & (!g2437) & (!g2438) & (!g2453)) + ((!g75) & (g2111) & (!g2280) & (!g2437) & (g2438) & (!g2453)) + ((!g75) & (g2111) & (!g2280) & (g2437) & (!g2438) & (!g2453)) + ((!g75) & (g2111) & (!g2280) & (g2437) & (g2438) & (!g2453)) + ((!g75) & (g2111) & (g2280) & (!g2437) & (!g2438) & (!g2453)) + ((!g75) & (g2111) & (g2280) & (!g2437) & (!g2438) & (g2453)) + ((!g75) & (g2111) & (g2280) & (!g2437) & (g2438) & (!g2453)) + ((!g75) & (g2111) & (g2280) & (!g2437) & (g2438) & (g2453)) + ((!g75) & (g2111) & (g2280) & (g2437) & (!g2438) & (!g2453)) + ((!g75) & (g2111) & (g2280) & (g2437) & (!g2438) & (g2453)) + ((!g75) & (g2111) & (g2280) & (g2437) & (g2438) & (!g2453)) + ((!g75) & (g2111) & (g2280) & (g2437) & (g2438) & (g2453)) + ((g75) & (!g2111) & (!g2280) & (!g2437) & (g2438) & (!g2453)) + ((g75) & (!g2111) & (!g2280) & (!g2437) & (g2438) & (g2453)) + ((g75) & (!g2111) & (!g2280) & (g2437) & (!g2438) & (!g2453)) + ((g75) & (!g2111) & (!g2280) & (g2437) & (!g2438) & (g2453)) + ((g75) & (!g2111) & (!g2280) & (g2437) & (g2438) & (!g2453)) + ((g75) & (!g2111) & (!g2280) & (g2437) & (g2438) & (g2453)) + ((g75) & (!g2111) & (g2280) & (!g2437) & (g2438) & (!g2453)) + ((g75) & (!g2111) & (g2280) & (!g2437) & (g2438) & (g2453)) + ((g75) & (!g2111) & (g2280) & (g2437) & (!g2438) & (!g2453)) + ((g75) & (!g2111) & (g2280) & (g2437) & (!g2438) & (g2453)) + ((g75) & (!g2111) & (g2280) & (g2437) & (g2438) & (!g2453)) + ((g75) & (!g2111) & (g2280) & (g2437) & (g2438) & (g2453)) + ((g75) & (g2111) & (!g2280) & (!g2437) & (g2438) & (!g2453)) + ((g75) & (g2111) & (!g2280) & (!g2437) & (g2438) & (g2453)) + ((g75) & (g2111) & (!g2280) & (g2437) & (!g2438) & (!g2453)) + ((g75) & (g2111) & (!g2280) & (g2437) & (!g2438) & (g2453)) + ((g75) & (g2111) & (!g2280) & (g2437) & (g2438) & (!g2453)) + ((g75) & (g2111) & (!g2280) & (g2437) & (g2438) & (g2453)) + ((g75) & (g2111) & (g2280) & (!g2437) & (g2438) & (!g2453)) + ((g75) & (g2111) & (g2280) & (!g2437) & (g2438) & (g2453)) + ((g75) & (g2111) & (g2280) & (g2437) & (!g2438) & (!g2453)) + ((g75) & (g2111) & (g2280) & (g2437) & (!g2438) & (g2453)) + ((g75) & (g2111) & (g2280) & (g2437) & (g2438) & (!g2453)) + ((g75) & (g2111) & (g2280) & (g2437) & (g2438) & (g2453)));
	assign g2455 = (((g2131) & (g2132) & (!dmem_dat_ix28x) & (!g2128) & (g2129) & (dmem_dat_ix12x)) + ((g2131) & (g2132) & (dmem_dat_ix28x) & (!g2128) & (!g2129) & (!dmem_dat_ix12x)) + ((g2131) & (g2132) & (dmem_dat_ix28x) & (!g2128) & (!g2129) & (dmem_dat_ix12x)) + ((g2131) & (g2132) & (dmem_dat_ix28x) & (!g2128) & (g2129) & (dmem_dat_ix12x)));
	assign g2456 = (((!g2363) & (!g2131) & (!sk[35]) & (!g2132) & (dmem_dat_ix12x) & (!g2338)) + ((!g2363) & (!g2131) & (!sk[35]) & (!g2132) & (dmem_dat_ix12x) & (g2338)) + ((!g2363) & (!g2131) & (!sk[35]) & (g2132) & (!dmem_dat_ix12x) & (!g2338)) + ((!g2363) & (!g2131) & (!sk[35]) & (g2132) & (!dmem_dat_ix12x) & (g2338)) + ((!g2363) & (!g2131) & (!sk[35]) & (g2132) & (dmem_dat_ix12x) & (!g2338)) + ((!g2363) & (!g2131) & (!sk[35]) & (g2132) & (dmem_dat_ix12x) & (g2338)) + ((!g2363) & (g2131) & (!sk[35]) & (!g2132) & (!dmem_dat_ix12x) & (!g2338)) + ((!g2363) & (g2131) & (!sk[35]) & (!g2132) & (!dmem_dat_ix12x) & (g2338)) + ((!g2363) & (g2131) & (!sk[35]) & (!g2132) & (dmem_dat_ix12x) & (!g2338)) + ((!g2363) & (g2131) & (!sk[35]) & (!g2132) & (dmem_dat_ix12x) & (g2338)) + ((!g2363) & (g2131) & (!sk[35]) & (g2132) & (!dmem_dat_ix12x) & (!g2338)) + ((!g2363) & (g2131) & (!sk[35]) & (g2132) & (!dmem_dat_ix12x) & (g2338)) + ((!g2363) & (g2131) & (!sk[35]) & (g2132) & (dmem_dat_ix12x) & (!g2338)) + ((!g2363) & (g2131) & (!sk[35]) & (g2132) & (dmem_dat_ix12x) & (g2338)) + ((!g2363) & (g2131) & (sk[35]) & (!g2132) & (dmem_dat_ix12x) & (!g2338)) + ((!g2363) & (g2131) & (sk[35]) & (!g2132) & (dmem_dat_ix12x) & (g2338)) + ((g2363) & (!g2131) & (!sk[35]) & (!g2132) & (dmem_dat_ix12x) & (!g2338)) + ((g2363) & (!g2131) & (!sk[35]) & (!g2132) & (dmem_dat_ix12x) & (g2338)) + ((g2363) & (!g2131) & (!sk[35]) & (g2132) & (!dmem_dat_ix12x) & (!g2338)) + ((g2363) & (!g2131) & (!sk[35]) & (g2132) & (!dmem_dat_ix12x) & (g2338)) + ((g2363) & (!g2131) & (!sk[35]) & (g2132) & (dmem_dat_ix12x) & (!g2338)) + ((g2363) & (!g2131) & (!sk[35]) & (g2132) & (dmem_dat_ix12x) & (g2338)) + ((g2363) & (!g2131) & (sk[35]) & (!g2132) & (!dmem_dat_ix12x) & (g2338)) + ((g2363) & (!g2131) & (sk[35]) & (!g2132) & (dmem_dat_ix12x) & (g2338)) + ((g2363) & (!g2131) & (sk[35]) & (g2132) & (!dmem_dat_ix12x) & (g2338)) + ((g2363) & (!g2131) & (sk[35]) & (g2132) & (dmem_dat_ix12x) & (g2338)) + ((g2363) & (g2131) & (!sk[35]) & (!g2132) & (!dmem_dat_ix12x) & (!g2338)) + ((g2363) & (g2131) & (!sk[35]) & (!g2132) & (!dmem_dat_ix12x) & (g2338)) + ((g2363) & (g2131) & (!sk[35]) & (!g2132) & (dmem_dat_ix12x) & (!g2338)) + ((g2363) & (g2131) & (!sk[35]) & (!g2132) & (dmem_dat_ix12x) & (g2338)) + ((g2363) & (g2131) & (!sk[35]) & (g2132) & (!dmem_dat_ix12x) & (!g2338)) + ((g2363) & (g2131) & (!sk[35]) & (g2132) & (!dmem_dat_ix12x) & (g2338)) + ((g2363) & (g2131) & (!sk[35]) & (g2132) & (dmem_dat_ix12x) & (!g2338)) + ((g2363) & (g2131) & (!sk[35]) & (g2132) & (dmem_dat_ix12x) & (g2338)) + ((g2363) & (g2131) & (sk[35]) & (!g2132) & (dmem_dat_ix12x) & (!g2338)) + ((g2363) & (g2131) & (sk[35]) & (!g2132) & (dmem_dat_ix12x) & (g2338)));
	assign g2458 = (((!g2111) & (!g2118) & (!g2439) & (g2457) & (!g2441) & (!g2442)) + ((!g2111) & (!g2118) & (!g2439) & (g2457) & (!g2441) & (g2442)) + ((!g2111) & (!g2118) & (!g2439) & (g2457) & (g2441) & (!g2442)) + ((!g2111) & (!g2118) & (!g2439) & (g2457) & (g2441) & (g2442)) + ((!g2111) & (!g2118) & (g2439) & (!g2457) & (!g2441) & (g2442)) + ((!g2111) & (!g2118) & (g2439) & (!g2457) & (g2441) & (!g2442)) + ((!g2111) & (!g2118) & (g2439) & (!g2457) & (g2441) & (g2442)) + ((!g2111) & (!g2118) & (g2439) & (g2457) & (!g2441) & (!g2442)) + ((!g2111) & (g2118) & (!g2439) & (!g2457) & (!g2441) & (!g2442)) + ((!g2111) & (g2118) & (!g2439) & (!g2457) & (!g2441) & (g2442)) + ((!g2111) & (g2118) & (!g2439) & (!g2457) & (g2441) & (!g2442)) + ((!g2111) & (g2118) & (!g2439) & (!g2457) & (g2441) & (g2442)) + ((!g2111) & (g2118) & (g2439) & (!g2457) & (!g2441) & (!g2442)) + ((!g2111) & (g2118) & (g2439) & (g2457) & (!g2441) & (g2442)) + ((!g2111) & (g2118) & (g2439) & (g2457) & (g2441) & (!g2442)) + ((!g2111) & (g2118) & (g2439) & (g2457) & (g2441) & (g2442)) + ((g2111) & (!g2118) & (!g2439) & (!g2457) & (!g2441) & (g2442)) + ((g2111) & (!g2118) & (!g2439) & (!g2457) & (g2441) & (!g2442)) + ((g2111) & (!g2118) & (!g2439) & (!g2457) & (g2441) & (g2442)) + ((g2111) & (!g2118) & (!g2439) & (g2457) & (!g2441) & (!g2442)) + ((g2111) & (!g2118) & (g2439) & (!g2457) & (!g2441) & (!g2442)) + ((g2111) & (!g2118) & (g2439) & (!g2457) & (!g2441) & (g2442)) + ((g2111) & (!g2118) & (g2439) & (!g2457) & (g2441) & (!g2442)) + ((g2111) & (!g2118) & (g2439) & (!g2457) & (g2441) & (g2442)) + ((g2111) & (g2118) & (!g2439) & (!g2457) & (!g2441) & (!g2442)) + ((g2111) & (g2118) & (!g2439) & (g2457) & (!g2441) & (g2442)) + ((g2111) & (g2118) & (!g2439) & (g2457) & (g2441) & (!g2442)) + ((g2111) & (g2118) & (!g2439) & (g2457) & (g2441) & (g2442)) + ((g2111) & (g2118) & (g2439) & (g2457) & (!g2441) & (!g2442)) + ((g2111) & (g2118) & (g2439) & (g2457) & (!g2441) & (g2442)) + ((g2111) & (g2118) & (g2439) & (g2457) & (g2441) & (!g2442)) + ((g2111) & (g2118) & (g2439) & (g2457) & (g2441) & (g2442)));
	assign g2459 = (((!g2419) & (!sk[37]) & (!g2420) & (!g2443) & (g2458)) + ((!g2419) & (!sk[37]) & (!g2420) & (g2443) & (!g2458)) + ((!g2419) & (!sk[37]) & (!g2420) & (g2443) & (g2458)) + ((!g2419) & (!sk[37]) & (g2420) & (!g2443) & (!g2458)) + ((!g2419) & (!sk[37]) & (g2420) & (!g2443) & (g2458)) + ((!g2419) & (!sk[37]) & (g2420) & (g2443) & (!g2458)) + ((!g2419) & (!sk[37]) & (g2420) & (g2443) & (g2458)) + ((!g2419) & (sk[37]) & (!g2420) & (!g2443) & (g2458)) + ((!g2419) & (sk[37]) & (!g2420) & (g2443) & (g2458)) + ((!g2419) & (sk[37]) & (g2420) & (!g2443) & (g2458)) + ((!g2419) & (sk[37]) & (g2420) & (g2443) & (g2458)) + ((g2419) & (!sk[37]) & (!g2420) & (!g2443) & (g2458)) + ((g2419) & (!sk[37]) & (!g2420) & (g2443) & (!g2458)) + ((g2419) & (!sk[37]) & (!g2420) & (g2443) & (g2458)) + ((g2419) & (!sk[37]) & (g2420) & (!g2443) & (!g2458)) + ((g2419) & (!sk[37]) & (g2420) & (!g2443) & (g2458)) + ((g2419) & (!sk[37]) & (g2420) & (g2443) & (!g2458)) + ((g2419) & (!sk[37]) & (g2420) & (g2443) & (g2458)) + ((g2419) & (sk[37]) & (!g2420) & (!g2443) & (g2458)) + ((g2419) & (sk[37]) & (!g2420) & (g2443) & (g2458)) + ((g2419) & (sk[37]) & (g2420) & (!g2443) & (g2458)) + ((g2419) & (sk[37]) & (g2420) & (g2443) & (!g2458)));
	assign g2460 = (((!g2444) & (sk[38]) & (g2445)) + ((g2444) & (!sk[38]) & (!g2445)) + ((g2444) & (!sk[38]) & (g2445)) + ((g2444) & (sk[38]) & (!g2445)));
	assign g2461 = (((!g2395) & (!g2396) & (!g2397) & (g2422) & (g2423) & (g2460)) + ((!g2395) & (!g2396) & (g2397) & (!g2422) & (g2423) & (g2460)) + ((!g2395) & (!g2396) & (g2397) & (g2422) & (!g2423) & (g2460)) + ((!g2395) & (!g2396) & (g2397) & (g2422) & (g2423) & (g2460)) + ((!g2395) & (g2396) & (!g2397) & (!g2422) & (g2423) & (g2460)) + ((!g2395) & (g2396) & (!g2397) & (g2422) & (!g2423) & (g2460)) + ((!g2395) & (g2396) & (!g2397) & (g2422) & (g2423) & (g2460)) + ((!g2395) & (g2396) & (g2397) & (!g2422) & (g2423) & (g2460)) + ((!g2395) & (g2396) & (g2397) & (g2422) & (!g2423) & (g2460)) + ((!g2395) & (g2396) & (g2397) & (g2422) & (g2423) & (g2460)) + ((g2395) & (!g2396) & (!g2397) & (g2422) & (g2423) & (g2460)) + ((g2395) & (!g2396) & (g2397) & (g2422) & (g2423) & (g2460)) + ((g2395) & (g2396) & (!g2397) & (g2422) & (g2423) & (g2460)) + ((g2395) & (g2396) & (g2397) & (!g2422) & (g2423) & (g2460)) + ((g2395) & (g2396) & (g2397) & (g2422) & (!g2423) & (g2460)) + ((g2395) & (g2396) & (g2397) & (g2422) & (g2423) & (g2460)));
	assign g2462 = (((g2444) & (!sk[40]) & (!g2445)) + ((g2444) & (!sk[40]) & (g2445)) + ((g2444) & (sk[40]) & (g2445)));
	assign g2463 = (((!sk[41]) & (g2461) & (!g2462)) + ((!sk[41]) & (g2461) & (g2462)) + ((sk[41]) & (!g2461) & (!g2462)));
	assign g2464 = (((g2111) & (!sk[42]) & (!g2439)) + ((g2111) & (!sk[42]) & (g2439)) + ((g2111) & (sk[42]) & (!g2439)));
	assign g2465 = (((!sk[43]) & (g2118) & (!g2457)) + ((!sk[43]) & (g2118) & (g2457)) + ((sk[43]) & (!g2118) & (!g2457)) + ((sk[43]) & (g2118) & (g2457)));
	assign g2466 = (((!g2463) & (!g2464) & (!sk[44]) & (g2465)) + ((!g2463) & (!g2464) & (sk[44]) & (!g2465)) + ((!g2463) & (g2464) & (!sk[44]) & (!g2465)) + ((!g2463) & (g2464) & (!sk[44]) & (g2465)) + ((!g2463) & (g2464) & (sk[44]) & (g2465)) + ((g2463) & (!g2464) & (!sk[44]) & (g2465)) + ((g2463) & (!g2464) & (sk[44]) & (g2465)) + ((g2463) & (g2464) & (!sk[44]) & (!g2465)) + ((g2463) & (g2464) & (!sk[44]) & (g2465)) + ((g2463) & (g2464) & (sk[44]) & (!g2465)));
	assign g2467 = (((!g2118) & (!g2111) & (!g2110) & (g2109) & (g2071) & (g2074)) + ((!g2118) & (!g2111) & (g2110) & (!g2109) & (!g2071) & (g2074)) + ((!g2118) & (!g2111) & (g2110) & (g2109) & (!g2071) & (g2074)) + ((!g2118) & (!g2111) & (g2110) & (g2109) & (g2071) & (g2074)) + ((!g2118) & (g2111) & (!g2110) & (!g2109) & (g2071) & (!g2074)) + ((!g2118) & (g2111) & (!g2110) & (g2109) & (g2071) & (!g2074)) + ((!g2118) & (g2111) & (!g2110) & (g2109) & (g2071) & (g2074)) + ((!g2118) & (g2111) & (g2110) & (!g2109) & (!g2071) & (g2074)) + ((!g2118) & (g2111) & (g2110) & (!g2109) & (g2071) & (!g2074)) + ((!g2118) & (g2111) & (g2110) & (g2109) & (!g2071) & (g2074)) + ((!g2118) & (g2111) & (g2110) & (g2109) & (g2071) & (!g2074)) + ((!g2118) & (g2111) & (g2110) & (g2109) & (g2071) & (g2074)) + ((g2118) & (!g2111) & (!g2110) & (!g2109) & (!g2071) & (!g2074)) + ((g2118) & (!g2111) & (!g2110) & (g2109) & (!g2071) & (!g2074)) + ((g2118) & (!g2111) & (!g2110) & (g2109) & (g2071) & (g2074)) + ((g2118) & (!g2111) & (g2110) & (!g2109) & (!g2071) & (!g2074)) + ((g2118) & (!g2111) & (g2110) & (!g2109) & (!g2071) & (g2074)) + ((g2118) & (!g2111) & (g2110) & (g2109) & (!g2071) & (!g2074)) + ((g2118) & (!g2111) & (g2110) & (g2109) & (!g2071) & (g2074)) + ((g2118) & (!g2111) & (g2110) & (g2109) & (g2071) & (g2074)) + ((g2118) & (g2111) & (!g2110) & (!g2109) & (!g2071) & (!g2074)) + ((g2118) & (g2111) & (!g2110) & (!g2109) & (g2071) & (!g2074)) + ((g2118) & (g2111) & (!g2110) & (g2109) & (!g2071) & (!g2074)) + ((g2118) & (g2111) & (!g2110) & (g2109) & (g2071) & (!g2074)) + ((g2118) & (g2111) & (!g2110) & (g2109) & (g2071) & (g2074)) + ((g2118) & (g2111) & (g2110) & (!g2109) & (!g2071) & (!g2074)) + ((g2118) & (g2111) & (g2110) & (!g2109) & (!g2071) & (g2074)) + ((g2118) & (g2111) & (g2110) & (!g2109) & (g2071) & (!g2074)) + ((g2118) & (g2111) & (g2110) & (g2109) & (!g2071) & (!g2074)) + ((g2118) & (g2111) & (g2110) & (g2109) & (!g2071) & (g2074)) + ((g2118) & (g2111) & (g2110) & (g2109) & (g2071) & (!g2074)) + ((g2118) & (g2111) & (g2110) & (g2109) & (g2071) & (g2074)));
	assign g2468 = (((!g2467) & (!g2272) & (!g2372) & (g2075) & (g2076) & (g2077)) + ((!g2467) & (!g2272) & (g2372) & (!g2075) & (!g2076) & (g2077)) + ((!g2467) & (!g2272) & (g2372) & (g2075) & (!g2076) & (g2077)) + ((!g2467) & (!g2272) & (g2372) & (g2075) & (g2076) & (g2077)) + ((!g2467) & (g2272) & (!g2372) & (!g2075) & (g2076) & (!g2077)) + ((!g2467) & (g2272) & (!g2372) & (g2075) & (g2076) & (!g2077)) + ((!g2467) & (g2272) & (!g2372) & (g2075) & (g2076) & (g2077)) + ((!g2467) & (g2272) & (g2372) & (!g2075) & (!g2076) & (g2077)) + ((!g2467) & (g2272) & (g2372) & (!g2075) & (g2076) & (!g2077)) + ((!g2467) & (g2272) & (g2372) & (g2075) & (!g2076) & (g2077)) + ((!g2467) & (g2272) & (g2372) & (g2075) & (g2076) & (!g2077)) + ((!g2467) & (g2272) & (g2372) & (g2075) & (g2076) & (g2077)) + ((g2467) & (!g2272) & (!g2372) & (!g2075) & (!g2076) & (!g2077)) + ((g2467) & (!g2272) & (!g2372) & (g2075) & (!g2076) & (!g2077)) + ((g2467) & (!g2272) & (!g2372) & (g2075) & (g2076) & (g2077)) + ((g2467) & (!g2272) & (g2372) & (!g2075) & (!g2076) & (!g2077)) + ((g2467) & (!g2272) & (g2372) & (!g2075) & (!g2076) & (g2077)) + ((g2467) & (!g2272) & (g2372) & (g2075) & (!g2076) & (!g2077)) + ((g2467) & (!g2272) & (g2372) & (g2075) & (!g2076) & (g2077)) + ((g2467) & (!g2272) & (g2372) & (g2075) & (g2076) & (g2077)) + ((g2467) & (g2272) & (!g2372) & (!g2075) & (!g2076) & (!g2077)) + ((g2467) & (g2272) & (!g2372) & (!g2075) & (g2076) & (!g2077)) + ((g2467) & (g2272) & (!g2372) & (g2075) & (!g2076) & (!g2077)) + ((g2467) & (g2272) & (!g2372) & (g2075) & (g2076) & (!g2077)) + ((g2467) & (g2272) & (!g2372) & (g2075) & (g2076) & (g2077)) + ((g2467) & (g2272) & (g2372) & (!g2075) & (!g2076) & (!g2077)) + ((g2467) & (g2272) & (g2372) & (!g2075) & (!g2076) & (g2077)) + ((g2467) & (g2272) & (g2372) & (!g2075) & (g2076) & (!g2077)) + ((g2467) & (g2272) & (g2372) & (g2075) & (!g2076) & (!g2077)) + ((g2467) & (g2272) & (g2372) & (g2075) & (!g2076) & (g2077)) + ((g2467) & (g2272) & (g2372) & (g2075) & (g2076) & (!g2077)) + ((g2467) & (g2272) & (g2372) & (g2075) & (g2076) & (g2077)));
	assign g2469 = (((!sk[47]) & (!g2076) & (!g2077) & (!g2102) & (g2192)) + ((!sk[47]) & (!g2076) & (!g2077) & (g2102) & (!g2192)) + ((!sk[47]) & (!g2076) & (!g2077) & (g2102) & (g2192)) + ((!sk[47]) & (!g2076) & (g2077) & (!g2102) & (!g2192)) + ((!sk[47]) & (!g2076) & (g2077) & (!g2102) & (g2192)) + ((!sk[47]) & (!g2076) & (g2077) & (g2102) & (!g2192)) + ((!sk[47]) & (!g2076) & (g2077) & (g2102) & (g2192)) + ((!sk[47]) & (g2076) & (!g2077) & (!g2102) & (g2192)) + ((!sk[47]) & (g2076) & (!g2077) & (g2102) & (!g2192)) + ((!sk[47]) & (g2076) & (!g2077) & (g2102) & (g2192)) + ((!sk[47]) & (g2076) & (g2077) & (!g2102) & (!g2192)) + ((!sk[47]) & (g2076) & (g2077) & (!g2102) & (g2192)) + ((!sk[47]) & (g2076) & (g2077) & (g2102) & (!g2192)) + ((!sk[47]) & (g2076) & (g2077) & (g2102) & (g2192)) + ((sk[47]) & (!g2076) & (!g2077) & (g2102) & (!g2192)) + ((sk[47]) & (!g2076) & (!g2077) & (g2102) & (g2192)) + ((sk[47]) & (!g2076) & (g2077) & (!g2102) & (g2192)) + ((sk[47]) & (!g2076) & (g2077) & (g2102) & (g2192)) + ((sk[47]) & (g2076) & (!g2077) & (!g2102) & (g2192)) + ((sk[47]) & (g2076) & (!g2077) & (g2102) & (g2192)) + ((sk[47]) & (g2076) & (g2077) & (!g2102) & (g2192)) + ((sk[47]) & (g2076) & (g2077) & (g2102) & (g2192)));
	assign g2470 = (((!g2122) & (!g2097) & (!g2087) & (g2092) & (g2076) & (g2077)) + ((!g2122) & (!g2097) & (g2087) & (!g2092) & (!g2076) & (g2077)) + ((!g2122) & (!g2097) & (g2087) & (g2092) & (!g2076) & (g2077)) + ((!g2122) & (!g2097) & (g2087) & (g2092) & (g2076) & (g2077)) + ((!g2122) & (g2097) & (!g2087) & (!g2092) & (g2076) & (!g2077)) + ((!g2122) & (g2097) & (!g2087) & (g2092) & (g2076) & (!g2077)) + ((!g2122) & (g2097) & (!g2087) & (g2092) & (g2076) & (g2077)) + ((!g2122) & (g2097) & (g2087) & (!g2092) & (!g2076) & (g2077)) + ((!g2122) & (g2097) & (g2087) & (!g2092) & (g2076) & (!g2077)) + ((!g2122) & (g2097) & (g2087) & (g2092) & (!g2076) & (g2077)) + ((!g2122) & (g2097) & (g2087) & (g2092) & (g2076) & (!g2077)) + ((!g2122) & (g2097) & (g2087) & (g2092) & (g2076) & (g2077)) + ((g2122) & (!g2097) & (!g2087) & (!g2092) & (!g2076) & (!g2077)) + ((g2122) & (!g2097) & (!g2087) & (g2092) & (!g2076) & (!g2077)) + ((g2122) & (!g2097) & (!g2087) & (g2092) & (g2076) & (g2077)) + ((g2122) & (!g2097) & (g2087) & (!g2092) & (!g2076) & (!g2077)) + ((g2122) & (!g2097) & (g2087) & (!g2092) & (!g2076) & (g2077)) + ((g2122) & (!g2097) & (g2087) & (g2092) & (!g2076) & (!g2077)) + ((g2122) & (!g2097) & (g2087) & (g2092) & (!g2076) & (g2077)) + ((g2122) & (!g2097) & (g2087) & (g2092) & (g2076) & (g2077)) + ((g2122) & (g2097) & (!g2087) & (!g2092) & (!g2076) & (!g2077)) + ((g2122) & (g2097) & (!g2087) & (!g2092) & (g2076) & (!g2077)) + ((g2122) & (g2097) & (!g2087) & (g2092) & (!g2076) & (!g2077)) + ((g2122) & (g2097) & (!g2087) & (g2092) & (g2076) & (!g2077)) + ((g2122) & (g2097) & (!g2087) & (g2092) & (g2076) & (g2077)) + ((g2122) & (g2097) & (g2087) & (!g2092) & (!g2076) & (!g2077)) + ((g2122) & (g2097) & (g2087) & (!g2092) & (!g2076) & (g2077)) + ((g2122) & (g2097) & (g2087) & (!g2092) & (g2076) & (!g2077)) + ((g2122) & (g2097) & (g2087) & (g2092) & (!g2076) & (!g2077)) + ((g2122) & (g2097) & (g2087) & (g2092) & (!g2076) & (g2077)) + ((g2122) & (g2097) & (g2087) & (g2092) & (g2076) & (!g2077)) + ((g2122) & (g2097) & (g2087) & (g2092) & (g2076) & (g2077)));
	assign g2471 = (((!g2073) & (!g2080) & (!g2125) & (g2468) & (!g2469) & (!g2470)) + ((!g2073) & (!g2080) & (!g2125) & (g2468) & (!g2469) & (g2470)) + ((!g2073) & (!g2080) & (!g2125) & (g2468) & (g2469) & (!g2470)) + ((!g2073) & (!g2080) & (!g2125) & (g2468) & (g2469) & (g2470)) + ((!g2073) & (!g2080) & (g2125) & (!g2468) & (!g2469) & (g2470)) + ((!g2073) & (!g2080) & (g2125) & (!g2468) & (g2469) & (g2470)) + ((!g2073) & (!g2080) & (g2125) & (g2468) & (!g2469) & (g2470)) + ((!g2073) & (!g2080) & (g2125) & (g2468) & (g2469) & (g2470)) + ((!g2073) & (g2080) & (!g2125) & (g2468) & (!g2469) & (!g2470)) + ((!g2073) & (g2080) & (!g2125) & (g2468) & (!g2469) & (g2470)) + ((!g2073) & (g2080) & (!g2125) & (g2468) & (g2469) & (!g2470)) + ((!g2073) & (g2080) & (!g2125) & (g2468) & (g2469) & (g2470)) + ((!g2073) & (g2080) & (g2125) & (!g2468) & (!g2469) & (g2470)) + ((!g2073) & (g2080) & (g2125) & (!g2468) & (g2469) & (g2470)) + ((!g2073) & (g2080) & (g2125) & (g2468) & (!g2469) & (g2470)) + ((!g2073) & (g2080) & (g2125) & (g2468) & (g2469) & (g2470)) + ((g2073) & (!g2080) & (g2125) & (!g2468) & (g2469) & (!g2470)) + ((g2073) & (!g2080) & (g2125) & (!g2468) & (g2469) & (g2470)) + ((g2073) & (!g2080) & (g2125) & (g2468) & (g2469) & (!g2470)) + ((g2073) & (!g2080) & (g2125) & (g2468) & (g2469) & (g2470)) + ((g2073) & (g2080) & (!g2125) & (g2468) & (!g2469) & (!g2470)) + ((g2073) & (g2080) & (!g2125) & (g2468) & (!g2469) & (g2470)) + ((g2073) & (g2080) & (!g2125) & (g2468) & (g2469) & (!g2470)) + ((g2073) & (g2080) & (!g2125) & (g2468) & (g2469) & (g2470)) + ((g2073) & (g2080) & (g2125) & (!g2468) & (g2469) & (!g2470)) + ((g2073) & (g2080) & (g2125) & (!g2468) & (g2469) & (g2470)) + ((g2073) & (g2080) & (g2125) & (g2468) & (g2469) & (!g2470)) + ((g2073) & (g2080) & (g2125) & (g2468) & (g2469) & (g2470)));
	assign g2472 = (((!g2457) & (!g2118) & (!g2124) & (!g2264) & (!g3601) & (!g2471)) + ((!g2457) & (!g2118) & (!g2124) & (!g2264) & (g3601) & (!g2471)) + ((!g2457) & (!g2118) & (!g2124) & (g2264) & (!g3601) & (!g2471)) + ((!g2457) & (!g2118) & (!g2124) & (g2264) & (!g3601) & (g2471)) + ((!g2457) & (!g2118) & (g2124) & (!g2264) & (!g3601) & (!g2471)) + ((!g2457) & (!g2118) & (g2124) & (!g2264) & (!g3601) & (g2471)) + ((!g2457) & (!g2118) & (g2124) & (!g2264) & (g3601) & (!g2471)) + ((!g2457) & (!g2118) & (g2124) & (!g2264) & (g3601) & (g2471)) + ((!g2457) & (!g2118) & (g2124) & (g2264) & (!g3601) & (!g2471)) + ((!g2457) & (!g2118) & (g2124) & (g2264) & (!g3601) & (g2471)) + ((!g2457) & (!g2118) & (g2124) & (g2264) & (g3601) & (!g2471)) + ((!g2457) & (!g2118) & (g2124) & (g2264) & (g3601) & (g2471)) + ((!g2457) & (g2118) & (!g2124) & (!g2264) & (!g3601) & (!g2471)) + ((!g2457) & (g2118) & (!g2124) & (!g2264) & (g3601) & (!g2471)) + ((!g2457) & (g2118) & (!g2124) & (g2264) & (!g3601) & (!g2471)) + ((!g2457) & (g2118) & (!g2124) & (g2264) & (!g3601) & (g2471)) + ((g2457) & (!g2118) & (!g2124) & (!g2264) & (!g3601) & (!g2471)) + ((g2457) & (!g2118) & (!g2124) & (!g2264) & (g3601) & (!g2471)) + ((g2457) & (!g2118) & (!g2124) & (g2264) & (!g3601) & (!g2471)) + ((g2457) & (!g2118) & (!g2124) & (g2264) & (!g3601) & (g2471)) + ((g2457) & (g2118) & (!g2124) & (!g2264) & (!g3601) & (!g2471)) + ((g2457) & (g2118) & (!g2124) & (!g2264) & (g3601) & (!g2471)) + ((g2457) & (g2118) & (!g2124) & (g2264) & (!g3601) & (!g2471)) + ((g2457) & (g2118) & (!g2124) & (g2264) & (!g3601) & (g2471)) + ((g2457) & (g2118) & (g2124) & (g2264) & (!g3601) & (!g2471)) + ((g2457) & (g2118) & (g2124) & (g2264) & (!g3601) & (g2471)) + ((g2457) & (g2118) & (g2124) & (g2264) & (g3601) & (!g2471)) + ((g2457) & (g2118) & (g2124) & (g2264) & (g3601) & (g2471)));
	assign g2473 = (((!g75) & (!g2118) & (!g2280) & (!g2455) & (!g2456) & (!g2472)) + ((!g75) & (!g2118) & (!g2280) & (!g2455) & (g2456) & (!g2472)) + ((!g75) & (!g2118) & (!g2280) & (g2455) & (!g2456) & (!g2472)) + ((!g75) & (!g2118) & (!g2280) & (g2455) & (g2456) & (!g2472)) + ((!g75) & (g2118) & (!g2280) & (!g2455) & (!g2456) & (!g2472)) + ((!g75) & (g2118) & (!g2280) & (!g2455) & (g2456) & (!g2472)) + ((!g75) & (g2118) & (!g2280) & (g2455) & (!g2456) & (!g2472)) + ((!g75) & (g2118) & (!g2280) & (g2455) & (g2456) & (!g2472)) + ((!g75) & (g2118) & (g2280) & (!g2455) & (!g2456) & (!g2472)) + ((!g75) & (g2118) & (g2280) & (!g2455) & (!g2456) & (g2472)) + ((!g75) & (g2118) & (g2280) & (!g2455) & (g2456) & (!g2472)) + ((!g75) & (g2118) & (g2280) & (!g2455) & (g2456) & (g2472)) + ((!g75) & (g2118) & (g2280) & (g2455) & (!g2456) & (!g2472)) + ((!g75) & (g2118) & (g2280) & (g2455) & (!g2456) & (g2472)) + ((!g75) & (g2118) & (g2280) & (g2455) & (g2456) & (!g2472)) + ((!g75) & (g2118) & (g2280) & (g2455) & (g2456) & (g2472)) + ((g75) & (!g2118) & (!g2280) & (!g2455) & (g2456) & (!g2472)) + ((g75) & (!g2118) & (!g2280) & (!g2455) & (g2456) & (g2472)) + ((g75) & (!g2118) & (!g2280) & (g2455) & (!g2456) & (!g2472)) + ((g75) & (!g2118) & (!g2280) & (g2455) & (!g2456) & (g2472)) + ((g75) & (!g2118) & (!g2280) & (g2455) & (g2456) & (!g2472)) + ((g75) & (!g2118) & (!g2280) & (g2455) & (g2456) & (g2472)) + ((g75) & (!g2118) & (g2280) & (!g2455) & (g2456) & (!g2472)) + ((g75) & (!g2118) & (g2280) & (!g2455) & (g2456) & (g2472)) + ((g75) & (!g2118) & (g2280) & (g2455) & (!g2456) & (!g2472)) + ((g75) & (!g2118) & (g2280) & (g2455) & (!g2456) & (g2472)) + ((g75) & (!g2118) & (g2280) & (g2455) & (g2456) & (!g2472)) + ((g75) & (!g2118) & (g2280) & (g2455) & (g2456) & (g2472)) + ((g75) & (g2118) & (!g2280) & (!g2455) & (g2456) & (!g2472)) + ((g75) & (g2118) & (!g2280) & (!g2455) & (g2456) & (g2472)) + ((g75) & (g2118) & (!g2280) & (g2455) & (!g2456) & (!g2472)) + ((g75) & (g2118) & (!g2280) & (g2455) & (!g2456) & (g2472)) + ((g75) & (g2118) & (!g2280) & (g2455) & (g2456) & (!g2472)) + ((g75) & (g2118) & (!g2280) & (g2455) & (g2456) & (g2472)) + ((g75) & (g2118) & (g2280) & (!g2455) & (g2456) & (!g2472)) + ((g75) & (g2118) & (g2280) & (!g2455) & (g2456) & (g2472)) + ((g75) & (g2118) & (g2280) & (g2455) & (!g2456) & (!g2472)) + ((g75) & (g2118) & (g2280) & (g2455) & (!g2456) & (g2472)) + ((g75) & (g2118) & (g2280) & (g2455) & (g2456) & (!g2472)) + ((g75) & (g2118) & (g2280) & (g2455) & (g2456) & (g2472)));
	assign g2474 = (((!g630) & (!g587) & (!sk[52]) & (!g2409) & (g724)) + ((!g630) & (!g587) & (!sk[52]) & (g2409) & (!g724)) + ((!g630) & (!g587) & (!sk[52]) & (g2409) & (g724)) + ((!g630) & (!g587) & (sk[52]) & (!g2409) & (g724)) + ((!g630) & (!g587) & (sk[52]) & (g2409) & (g724)) + ((!g630) & (g587) & (!sk[52]) & (!g2409) & (!g724)) + ((!g630) & (g587) & (!sk[52]) & (!g2409) & (g724)) + ((!g630) & (g587) & (!sk[52]) & (g2409) & (!g724)) + ((!g630) & (g587) & (!sk[52]) & (g2409) & (g724)) + ((!g630) & (g587) & (sk[52]) & (!g2409) & (g724)) + ((!g630) & (g587) & (sk[52]) & (g2409) & (g724)) + ((g630) & (!g587) & (!sk[52]) & (!g2409) & (g724)) + ((g630) & (!g587) & (!sk[52]) & (g2409) & (!g724)) + ((g630) & (!g587) & (!sk[52]) & (g2409) & (g724)) + ((g630) & (!g587) & (sk[52]) & (!g2409) & (g724)) + ((g630) & (!g587) & (sk[52]) & (g2409) & (g724)) + ((g630) & (g587) & (!sk[52]) & (!g2409) & (!g724)) + ((g630) & (g587) & (!sk[52]) & (!g2409) & (g724)) + ((g630) & (g587) & (!sk[52]) & (g2409) & (!g724)) + ((g630) & (g587) & (!sk[52]) & (g2409) & (g724)) + ((g630) & (g587) & (sk[52]) & (!g2409) & (g724)) + ((g630) & (g587) & (sk[52]) & (g2409) & (!g724)));
	assign g2475 = (((!sk[53]) & (!g1759) & (!g2033) & (g2034)) + ((!sk[53]) & (!g1759) & (g2033) & (!g2034)) + ((!sk[53]) & (!g1759) & (g2033) & (g2034)) + ((!sk[53]) & (g1759) & (!g2033) & (g2034)) + ((!sk[53]) & (g1759) & (g2033) & (!g2034)) + ((!sk[53]) & (g1759) & (g2033) & (g2034)) + ((sk[53]) & (g1759) & (!g2033) & (g2034)));
	assign g5036 = (((!sk[54]) & (!g2921) & (!g3239) & (g2476)) + ((!sk[54]) & (!g2921) & (g3239) & (!g2476)) + ((!sk[54]) & (!g2921) & (g3239) & (g2476)) + ((!sk[54]) & (g2921) & (!g3239) & (g2476)) + ((!sk[54]) & (g2921) & (g3239) & (!g2476)) + ((!sk[54]) & (g2921) & (g3239) & (g2476)) + ((sk[54]) & (!g2921) & (!g3239) & (g2476)) + ((sk[54]) & (!g2921) & (g3239) & (g2476)) + ((sk[54]) & (g2921) & (g3239) & (!g2476)) + ((sk[54]) & (g2921) & (g3239) & (g2476)));
	assign g2477 = (((!g91) & (!g630) & (!g586) & (!sk[55]) & (g2433) & (!g724)) + ((!g91) & (!g630) & (!g586) & (!sk[55]) & (g2433) & (g724)) + ((!g91) & (!g630) & (!g586) & (sk[55]) & (!g2433) & (g724)) + ((!g91) & (!g630) & (!g586) & (sk[55]) & (g2433) & (g724)) + ((!g91) & (!g630) & (g586) & (!sk[55]) & (!g2433) & (!g724)) + ((!g91) & (!g630) & (g586) & (!sk[55]) & (!g2433) & (g724)) + ((!g91) & (!g630) & (g586) & (!sk[55]) & (g2433) & (!g724)) + ((!g91) & (!g630) & (g586) & (!sk[55]) & (g2433) & (g724)) + ((!g91) & (!g630) & (g586) & (sk[55]) & (!g2433) & (!g724)) + ((!g91) & (!g630) & (g586) & (sk[55]) & (g2433) & (!g724)) + ((!g91) & (g630) & (!g586) & (!sk[55]) & (!g2433) & (!g724)) + ((!g91) & (g630) & (!g586) & (!sk[55]) & (!g2433) & (g724)) + ((!g91) & (g630) & (!g586) & (!sk[55]) & (g2433) & (!g724)) + ((!g91) & (g630) & (!g586) & (!sk[55]) & (g2433) & (g724)) + ((!g91) & (g630) & (!g586) & (sk[55]) & (!g2433) & (g724)) + ((!g91) & (g630) & (!g586) & (sk[55]) & (g2433) & (!g724)) + ((!g91) & (g630) & (g586) & (!sk[55]) & (!g2433) & (!g724)) + ((!g91) & (g630) & (g586) & (!sk[55]) & (!g2433) & (g724)) + ((!g91) & (g630) & (g586) & (!sk[55]) & (g2433) & (!g724)) + ((!g91) & (g630) & (g586) & (!sk[55]) & (g2433) & (g724)) + ((!g91) & (g630) & (g586) & (sk[55]) & (!g2433) & (!g724)) + ((!g91) & (g630) & (g586) & (sk[55]) & (g2433) & (g724)) + ((g91) & (!g630) & (!g586) & (!sk[55]) & (g2433) & (!g724)) + ((g91) & (!g630) & (!g586) & (!sk[55]) & (g2433) & (g724)) + ((g91) & (!g630) & (!g586) & (sk[55]) & (!g2433) & (g724)) + ((g91) & (!g630) & (!g586) & (sk[55]) & (g2433) & (!g724)) + ((g91) & (!g630) & (g586) & (!sk[55]) & (!g2433) & (!g724)) + ((g91) & (!g630) & (g586) & (!sk[55]) & (!g2433) & (g724)) + ((g91) & (!g630) & (g586) & (!sk[55]) & (g2433) & (!g724)) + ((g91) & (!g630) & (g586) & (!sk[55]) & (g2433) & (g724)) + ((g91) & (!g630) & (g586) & (sk[55]) & (!g2433) & (!g724)) + ((g91) & (!g630) & (g586) & (sk[55]) & (g2433) & (g724)) + ((g91) & (g630) & (!g586) & (!sk[55]) & (!g2433) & (!g724)) + ((g91) & (g630) & (!g586) & (!sk[55]) & (!g2433) & (g724)) + ((g91) & (g630) & (!g586) & (!sk[55]) & (g2433) & (!g724)) + ((g91) & (g630) & (!g586) & (!sk[55]) & (g2433) & (g724)) + ((g91) & (g630) & (!g586) & (sk[55]) & (!g2433) & (!g724)) + ((g91) & (g630) & (!g586) & (sk[55]) & (g2433) & (!g724)) + ((g91) & (g630) & (g586) & (!sk[55]) & (!g2433) & (!g724)) + ((g91) & (g630) & (g586) & (!sk[55]) & (!g2433) & (g724)) + ((g91) & (g630) & (g586) & (!sk[55]) & (g2433) & (!g724)) + ((g91) & (g630) & (g586) & (!sk[55]) & (g2433) & (g724)) + ((g91) & (g630) & (g586) & (sk[55]) & (!g2433) & (g724)) + ((g91) & (g630) & (g586) & (sk[55]) & (g2433) & (g724)));
	assign g2478 = (((!sk[56]) & (!g2033) & (!g2034) & (!g2476) & (g2477)) + ((!sk[56]) & (!g2033) & (!g2034) & (g2476) & (!g2477)) + ((!sk[56]) & (!g2033) & (!g2034) & (g2476) & (g2477)) + ((!sk[56]) & (!g2033) & (g2034) & (!g2476) & (!g2477)) + ((!sk[56]) & (!g2033) & (g2034) & (!g2476) & (g2477)) + ((!sk[56]) & (!g2033) & (g2034) & (g2476) & (!g2477)) + ((!sk[56]) & (!g2033) & (g2034) & (g2476) & (g2477)) + ((!sk[56]) & (g2033) & (!g2034) & (!g2476) & (g2477)) + ((!sk[56]) & (g2033) & (!g2034) & (g2476) & (!g2477)) + ((!sk[56]) & (g2033) & (!g2034) & (g2476) & (g2477)) + ((!sk[56]) & (g2033) & (g2034) & (!g2476) & (!g2477)) + ((!sk[56]) & (g2033) & (g2034) & (!g2476) & (g2477)) + ((!sk[56]) & (g2033) & (g2034) & (g2476) & (!g2477)) + ((!sk[56]) & (g2033) & (g2034) & (g2476) & (g2477)) + ((sk[56]) & (!g2033) & (!g2034) & (g2476) & (!g2477)) + ((sk[56]) & (!g2033) & (!g2034) & (g2476) & (g2477)) + ((sk[56]) & (g2033) & (!g2034) & (!g2476) & (g2477)) + ((sk[56]) & (g2033) & (!g2034) & (g2476) & (g2477)));
	assign g2479 = (((g2329) & (!g2029) & (g2408) & (!g2474) & (!g2475) & (g2478)) + ((g2329) & (!g2029) & (g2408) & (!g2474) & (g2475) & (!g2478)) + ((g2329) & (!g2029) & (g2408) & (!g2474) & (g2475) & (g2478)) + ((g2329) & (!g2029) & (g2408) & (g2474) & (!g2475) & (g2478)) + ((g2329) & (!g2029) & (g2408) & (g2474) & (g2475) & (!g2478)) + ((g2329) & (!g2029) & (g2408) & (g2474) & (g2475) & (g2478)) + ((g2329) & (g2029) & (g2408) & (g2474) & (!g2475) & (!g2478)) + ((g2329) & (g2029) & (g2408) & (g2474) & (!g2475) & (g2478)) + ((g2329) & (g2029) & (g2408) & (g2474) & (g2475) & (!g2478)) + ((g2329) & (g2029) & (g2408) & (g2474) & (g2475) & (g2478)));
	assign g2480 = (((g2131) & (g2132) & (!dmem_dat_ix29x) & (!g2128) & (g2129) & (dmem_dat_ix13x)) + ((g2131) & (g2132) & (dmem_dat_ix29x) & (!g2128) & (!g2129) & (!dmem_dat_ix13x)) + ((g2131) & (g2132) & (dmem_dat_ix29x) & (!g2128) & (!g2129) & (dmem_dat_ix13x)) + ((g2131) & (g2132) & (dmem_dat_ix29x) & (!g2128) & (g2129) & (dmem_dat_ix13x)));
	assign g2481 = (((!g2363) & (!g2131) & (!g2132) & (dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((!g2363) & (!g2131) & (!g2132) & (dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((!g2363) & (!g2131) & (g2132) & (!dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((!g2363) & (!g2131) & (g2132) & (!dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((!g2363) & (!g2131) & (g2132) & (dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((!g2363) & (!g2131) & (g2132) & (dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((!g2363) & (g2131) & (!g2132) & (!dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((!g2363) & (g2131) & (!g2132) & (!dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((!g2363) & (g2131) & (!g2132) & (dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((!g2363) & (g2131) & (!g2132) & (dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((!g2363) & (g2131) & (!g2132) & (dmem_dat_ix13x) & (sk[59]) & (!g2338)) + ((!g2363) & (g2131) & (!g2132) & (dmem_dat_ix13x) & (sk[59]) & (g2338)) + ((!g2363) & (g2131) & (g2132) & (!dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((!g2363) & (g2131) & (g2132) & (!dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((!g2363) & (g2131) & (g2132) & (dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((!g2363) & (g2131) & (g2132) & (dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((g2363) & (!g2131) & (!g2132) & (!dmem_dat_ix13x) & (sk[59]) & (g2338)) + ((g2363) & (!g2131) & (!g2132) & (dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((g2363) & (!g2131) & (!g2132) & (dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((g2363) & (!g2131) & (!g2132) & (dmem_dat_ix13x) & (sk[59]) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (!dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((g2363) & (!g2131) & (g2132) & (!dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (!dmem_dat_ix13x) & (sk[59]) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((g2363) & (!g2131) & (g2132) & (dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (dmem_dat_ix13x) & (sk[59]) & (g2338)) + ((g2363) & (g2131) & (!g2132) & (!dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((g2363) & (g2131) & (!g2132) & (!dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((g2363) & (g2131) & (!g2132) & (dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((g2363) & (g2131) & (!g2132) & (dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((g2363) & (g2131) & (!g2132) & (dmem_dat_ix13x) & (sk[59]) & (!g2338)) + ((g2363) & (g2131) & (!g2132) & (dmem_dat_ix13x) & (sk[59]) & (g2338)) + ((g2363) & (g2131) & (g2132) & (!dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((g2363) & (g2131) & (g2132) & (!dmem_dat_ix13x) & (!sk[59]) & (g2338)) + ((g2363) & (g2131) & (g2132) & (dmem_dat_ix13x) & (!sk[59]) & (!g2338)) + ((g2363) & (g2131) & (g2132) & (dmem_dat_ix13x) & (!sk[59]) & (g2338)));
	assign g2483 = (((!g2111) & (!g2118) & (g2439) & (!g2441) & (g2442) & (g2457)) + ((!g2111) & (!g2118) & (g2439) & (g2441) & (!g2442) & (g2457)) + ((!g2111) & (!g2118) & (g2439) & (g2441) & (g2442) & (g2457)) + ((!g2111) & (g2118) & (!g2439) & (!g2441) & (!g2442) & (g2457)) + ((!g2111) & (g2118) & (!g2439) & (!g2441) & (g2442) & (g2457)) + ((!g2111) & (g2118) & (!g2439) & (g2441) & (!g2442) & (g2457)) + ((!g2111) & (g2118) & (!g2439) & (g2441) & (g2442) & (g2457)) + ((!g2111) & (g2118) & (g2439) & (!g2441) & (!g2442) & (g2457)) + ((!g2111) & (g2118) & (g2439) & (!g2441) & (g2442) & (!g2457)) + ((!g2111) & (g2118) & (g2439) & (!g2441) & (g2442) & (g2457)) + ((!g2111) & (g2118) & (g2439) & (g2441) & (!g2442) & (!g2457)) + ((!g2111) & (g2118) & (g2439) & (g2441) & (!g2442) & (g2457)) + ((!g2111) & (g2118) & (g2439) & (g2441) & (g2442) & (!g2457)) + ((!g2111) & (g2118) & (g2439) & (g2441) & (g2442) & (g2457)) + ((g2111) & (!g2118) & (!g2439) & (!g2441) & (g2442) & (g2457)) + ((g2111) & (!g2118) & (!g2439) & (g2441) & (!g2442) & (g2457)) + ((g2111) & (!g2118) & (!g2439) & (g2441) & (g2442) & (g2457)) + ((g2111) & (!g2118) & (g2439) & (!g2441) & (!g2442) & (g2457)) + ((g2111) & (!g2118) & (g2439) & (!g2441) & (g2442) & (g2457)) + ((g2111) & (!g2118) & (g2439) & (g2441) & (!g2442) & (g2457)) + ((g2111) & (!g2118) & (g2439) & (g2441) & (g2442) & (g2457)) + ((g2111) & (g2118) & (!g2439) & (!g2441) & (!g2442) & (g2457)) + ((g2111) & (g2118) & (!g2439) & (!g2441) & (g2442) & (!g2457)) + ((g2111) & (g2118) & (!g2439) & (!g2441) & (g2442) & (g2457)) + ((g2111) & (g2118) & (!g2439) & (g2441) & (!g2442) & (!g2457)) + ((g2111) & (g2118) & (!g2439) & (g2441) & (!g2442) & (g2457)) + ((g2111) & (g2118) & (!g2439) & (g2441) & (g2442) & (!g2457)) + ((g2111) & (g2118) & (!g2439) & (g2441) & (g2442) & (g2457)) + ((g2111) & (g2118) & (g2439) & (!g2441) & (!g2442) & (!g2457)) + ((g2111) & (g2118) & (g2439) & (!g2441) & (!g2442) & (g2457)) + ((g2111) & (g2118) & (g2439) & (!g2441) & (g2442) & (!g2457)) + ((g2111) & (g2118) & (g2439) & (!g2441) & (g2442) & (g2457)) + ((g2111) & (g2118) & (g2439) & (g2441) & (!g2442) & (!g2457)) + ((g2111) & (g2118) & (g2439) & (g2441) & (!g2442) & (g2457)) + ((g2111) & (g2118) & (g2439) & (g2441) & (g2442) & (!g2457)) + ((g2111) & (g2118) & (g2439) & (g2441) & (g2442) & (g2457)));
	assign g2484 = (((!g2119) & (!g2482) & (!sk[61]) & (g2483)) + ((!g2119) & (!g2482) & (sk[61]) & (g2483)) + ((!g2119) & (g2482) & (!sk[61]) & (!g2483)) + ((!g2119) & (g2482) & (!sk[61]) & (g2483)) + ((!g2119) & (g2482) & (sk[61]) & (!g2483)) + ((g2119) & (!g2482) & (!sk[61]) & (g2483)) + ((g2119) & (!g2482) & (sk[61]) & (!g2483)) + ((g2119) & (g2482) & (!sk[61]) & (!g2483)) + ((g2119) & (g2482) & (!sk[61]) & (g2483)) + ((g2119) & (g2482) & (sk[61]) & (g2483)));
	assign g2485 = (((!g2419) & (!g2420) & (!g2443) & (!sk[62]) & (g2458)) + ((!g2419) & (!g2420) & (g2443) & (!sk[62]) & (!g2458)) + ((!g2419) & (!g2420) & (g2443) & (!sk[62]) & (g2458)) + ((!g2419) & (g2420) & (!g2443) & (!sk[62]) & (!g2458)) + ((!g2419) & (g2420) & (!g2443) & (!sk[62]) & (g2458)) + ((!g2419) & (g2420) & (g2443) & (!sk[62]) & (!g2458)) + ((!g2419) & (g2420) & (g2443) & (!sk[62]) & (g2458)) + ((g2419) & (!g2420) & (!g2443) & (!sk[62]) & (g2458)) + ((g2419) & (!g2420) & (g2443) & (!sk[62]) & (!g2458)) + ((g2419) & (!g2420) & (g2443) & (!sk[62]) & (g2458)) + ((g2419) & (g2420) & (!g2443) & (!sk[62]) & (!g2458)) + ((g2419) & (g2420) & (!g2443) & (!sk[62]) & (g2458)) + ((g2419) & (g2420) & (g2443) & (!sk[62]) & (!g2458)) + ((g2419) & (g2420) & (g2443) & (!sk[62]) & (g2458)) + ((g2419) & (g2420) & (g2443) & (sk[62]) & (g2458)));
	assign g2486 = (((!sk[63]) & (g2118) & (!g2457)) + ((!sk[63]) & (g2118) & (g2457)) + ((sk[63]) & (g2118) & (!g2457)));
	assign g2487 = (((!sk[64]) & (g2119) & (!g2482)) + ((!sk[64]) & (g2119) & (g2482)) + ((sk[64]) & (!g2119) & (!g2482)) + ((sk[64]) & (g2119) & (g2482)));
	assign g2488 = (((!g2463) & (!g2464) & (!g2465) & (!sk[65]) & (g2486) & (!g2487)) + ((!g2463) & (!g2464) & (!g2465) & (!sk[65]) & (g2486) & (g2487)) + ((!g2463) & (!g2464) & (!g2465) & (sk[65]) & (!g2486) & (g2487)) + ((!g2463) & (!g2464) & (!g2465) & (sk[65]) & (g2486) & (!g2487)) + ((!g2463) & (!g2464) & (g2465) & (!sk[65]) & (!g2486) & (!g2487)) + ((!g2463) & (!g2464) & (g2465) & (!sk[65]) & (!g2486) & (g2487)) + ((!g2463) & (!g2464) & (g2465) & (!sk[65]) & (g2486) & (!g2487)) + ((!g2463) & (!g2464) & (g2465) & (!sk[65]) & (g2486) & (g2487)) + ((!g2463) & (!g2464) & (g2465) & (sk[65]) & (!g2486) & (!g2487)) + ((!g2463) & (!g2464) & (g2465) & (sk[65]) & (g2486) & (g2487)) + ((!g2463) & (g2464) & (!g2465) & (!sk[65]) & (!g2486) & (!g2487)) + ((!g2463) & (g2464) & (!g2465) & (!sk[65]) & (!g2486) & (g2487)) + ((!g2463) & (g2464) & (!g2465) & (!sk[65]) & (g2486) & (!g2487)) + ((!g2463) & (g2464) & (!g2465) & (!sk[65]) & (g2486) & (g2487)) + ((!g2463) & (g2464) & (!g2465) & (sk[65]) & (!g2486) & (!g2487)) + ((!g2463) & (g2464) & (!g2465) & (sk[65]) & (g2486) & (g2487)) + ((!g2463) & (g2464) & (g2465) & (!sk[65]) & (!g2486) & (!g2487)) + ((!g2463) & (g2464) & (g2465) & (!sk[65]) & (!g2486) & (g2487)) + ((!g2463) & (g2464) & (g2465) & (!sk[65]) & (g2486) & (!g2487)) + ((!g2463) & (g2464) & (g2465) & (!sk[65]) & (g2486) & (g2487)) + ((!g2463) & (g2464) & (g2465) & (sk[65]) & (!g2486) & (!g2487)) + ((!g2463) & (g2464) & (g2465) & (sk[65]) & (g2486) & (g2487)) + ((g2463) & (!g2464) & (!g2465) & (!sk[65]) & (g2486) & (!g2487)) + ((g2463) & (!g2464) & (!g2465) & (!sk[65]) & (g2486) & (g2487)) + ((g2463) & (!g2464) & (!g2465) & (sk[65]) & (!g2486) & (g2487)) + ((g2463) & (!g2464) & (!g2465) & (sk[65]) & (g2486) & (!g2487)) + ((g2463) & (!g2464) & (g2465) & (!sk[65]) & (!g2486) & (!g2487)) + ((g2463) & (!g2464) & (g2465) & (!sk[65]) & (!g2486) & (g2487)) + ((g2463) & (!g2464) & (g2465) & (!sk[65]) & (g2486) & (!g2487)) + ((g2463) & (!g2464) & (g2465) & (!sk[65]) & (g2486) & (g2487)) + ((g2463) & (!g2464) & (g2465) & (sk[65]) & (!g2486) & (g2487)) + ((g2463) & (!g2464) & (g2465) & (sk[65]) & (g2486) & (!g2487)) + ((g2463) & (g2464) & (!g2465) & (!sk[65]) & (!g2486) & (!g2487)) + ((g2463) & (g2464) & (!g2465) & (!sk[65]) & (!g2486) & (g2487)) + ((g2463) & (g2464) & (!g2465) & (!sk[65]) & (g2486) & (!g2487)) + ((g2463) & (g2464) & (!g2465) & (!sk[65]) & (g2486) & (g2487)) + ((g2463) & (g2464) & (!g2465) & (sk[65]) & (!g2486) & (g2487)) + ((g2463) & (g2464) & (!g2465) & (sk[65]) & (g2486) & (!g2487)) + ((g2463) & (g2464) & (g2465) & (!sk[65]) & (!g2486) & (!g2487)) + ((g2463) & (g2464) & (g2465) & (!sk[65]) & (!g2486) & (g2487)) + ((g2463) & (g2464) & (g2465) & (!sk[65]) & (g2486) & (!g2487)) + ((g2463) & (g2464) & (g2465) & (!sk[65]) & (g2486) & (g2487)) + ((g2463) & (g2464) & (g2465) & (sk[65]) & (!g2486) & (!g2487)) + ((g2463) & (g2464) & (g2465) & (sk[65]) & (g2486) & (g2487)));
	assign g2489 = (((!sk[66]) & (!g2076) & (!g2077) & (!g2192) & (g2193)) + ((!sk[66]) & (!g2076) & (!g2077) & (g2192) & (!g2193)) + ((!sk[66]) & (!g2076) & (!g2077) & (g2192) & (g2193)) + ((!sk[66]) & (!g2076) & (g2077) & (!g2192) & (!g2193)) + ((!sk[66]) & (!g2076) & (g2077) & (!g2192) & (g2193)) + ((!sk[66]) & (!g2076) & (g2077) & (g2192) & (!g2193)) + ((!sk[66]) & (!g2076) & (g2077) & (g2192) & (g2193)) + ((!sk[66]) & (g2076) & (!g2077) & (!g2192) & (g2193)) + ((!sk[66]) & (g2076) & (!g2077) & (g2192) & (!g2193)) + ((!sk[66]) & (g2076) & (!g2077) & (g2192) & (g2193)) + ((!sk[66]) & (g2076) & (g2077) & (!g2192) & (!g2193)) + ((!sk[66]) & (g2076) & (g2077) & (!g2192) & (g2193)) + ((!sk[66]) & (g2076) & (g2077) & (g2192) & (!g2193)) + ((!sk[66]) & (g2076) & (g2077) & (g2192) & (g2193)) + ((sk[66]) & (!g2076) & (!g2077) & (!g2192) & (g2193)) + ((sk[66]) & (!g2076) & (!g2077) & (g2192) & (g2193)) + ((sk[66]) & (!g2076) & (g2077) & (g2192) & (!g2193)) + ((sk[66]) & (!g2076) & (g2077) & (g2192) & (g2193)) + ((sk[66]) & (g2076) & (!g2077) & (g2192) & (!g2193)) + ((sk[66]) & (g2076) & (!g2077) & (g2192) & (g2193)) + ((sk[66]) & (g2076) & (g2077) & (g2192) & (!g2193)) + ((sk[66]) & (g2076) & (g2077) & (g2192) & (g2193)));
	assign g2490 = (((!g2119) & (!g2118) & (!g2111) & (g2110) & (g2071) & (g2074)) + ((!g2119) & (!g2118) & (g2111) & (!g2110) & (!g2071) & (g2074)) + ((!g2119) & (!g2118) & (g2111) & (g2110) & (!g2071) & (g2074)) + ((!g2119) & (!g2118) & (g2111) & (g2110) & (g2071) & (g2074)) + ((!g2119) & (g2118) & (!g2111) & (!g2110) & (g2071) & (!g2074)) + ((!g2119) & (g2118) & (!g2111) & (g2110) & (g2071) & (!g2074)) + ((!g2119) & (g2118) & (!g2111) & (g2110) & (g2071) & (g2074)) + ((!g2119) & (g2118) & (g2111) & (!g2110) & (!g2071) & (g2074)) + ((!g2119) & (g2118) & (g2111) & (!g2110) & (g2071) & (!g2074)) + ((!g2119) & (g2118) & (g2111) & (g2110) & (!g2071) & (g2074)) + ((!g2119) & (g2118) & (g2111) & (g2110) & (g2071) & (!g2074)) + ((!g2119) & (g2118) & (g2111) & (g2110) & (g2071) & (g2074)) + ((g2119) & (!g2118) & (!g2111) & (!g2110) & (!g2071) & (!g2074)) + ((g2119) & (!g2118) & (!g2111) & (g2110) & (!g2071) & (!g2074)) + ((g2119) & (!g2118) & (!g2111) & (g2110) & (g2071) & (g2074)) + ((g2119) & (!g2118) & (g2111) & (!g2110) & (!g2071) & (!g2074)) + ((g2119) & (!g2118) & (g2111) & (!g2110) & (!g2071) & (g2074)) + ((g2119) & (!g2118) & (g2111) & (g2110) & (!g2071) & (!g2074)) + ((g2119) & (!g2118) & (g2111) & (g2110) & (!g2071) & (g2074)) + ((g2119) & (!g2118) & (g2111) & (g2110) & (g2071) & (g2074)) + ((g2119) & (g2118) & (!g2111) & (!g2110) & (!g2071) & (!g2074)) + ((g2119) & (g2118) & (!g2111) & (!g2110) & (g2071) & (!g2074)) + ((g2119) & (g2118) & (!g2111) & (g2110) & (!g2071) & (!g2074)) + ((g2119) & (g2118) & (!g2111) & (g2110) & (g2071) & (!g2074)) + ((g2119) & (g2118) & (!g2111) & (g2110) & (g2071) & (g2074)) + ((g2119) & (g2118) & (g2111) & (!g2110) & (!g2071) & (!g2074)) + ((g2119) & (g2118) & (g2111) & (!g2110) & (!g2071) & (g2074)) + ((g2119) & (g2118) & (g2111) & (!g2110) & (g2071) & (!g2074)) + ((g2119) & (g2118) & (g2111) & (g2110) & (!g2071) & (!g2074)) + ((g2119) & (g2118) & (g2111) & (g2110) & (!g2071) & (g2074)) + ((g2119) & (g2118) & (g2111) & (g2110) & (g2071) & (!g2074)) + ((g2119) & (g2118) & (g2111) & (g2110) & (g2071) & (g2074)));
	assign g2491 = (((!g2490) & (!g2296) & (!g2402) & (g2183) & (g2076) & (g2077)) + ((!g2490) & (!g2296) & (g2402) & (!g2183) & (!g2076) & (g2077)) + ((!g2490) & (!g2296) & (g2402) & (g2183) & (!g2076) & (g2077)) + ((!g2490) & (!g2296) & (g2402) & (g2183) & (g2076) & (g2077)) + ((!g2490) & (g2296) & (!g2402) & (!g2183) & (g2076) & (!g2077)) + ((!g2490) & (g2296) & (!g2402) & (g2183) & (g2076) & (!g2077)) + ((!g2490) & (g2296) & (!g2402) & (g2183) & (g2076) & (g2077)) + ((!g2490) & (g2296) & (g2402) & (!g2183) & (!g2076) & (g2077)) + ((!g2490) & (g2296) & (g2402) & (!g2183) & (g2076) & (!g2077)) + ((!g2490) & (g2296) & (g2402) & (g2183) & (!g2076) & (g2077)) + ((!g2490) & (g2296) & (g2402) & (g2183) & (g2076) & (!g2077)) + ((!g2490) & (g2296) & (g2402) & (g2183) & (g2076) & (g2077)) + ((g2490) & (!g2296) & (!g2402) & (!g2183) & (!g2076) & (!g2077)) + ((g2490) & (!g2296) & (!g2402) & (g2183) & (!g2076) & (!g2077)) + ((g2490) & (!g2296) & (!g2402) & (g2183) & (g2076) & (g2077)) + ((g2490) & (!g2296) & (g2402) & (!g2183) & (!g2076) & (!g2077)) + ((g2490) & (!g2296) & (g2402) & (!g2183) & (!g2076) & (g2077)) + ((g2490) & (!g2296) & (g2402) & (g2183) & (!g2076) & (!g2077)) + ((g2490) & (!g2296) & (g2402) & (g2183) & (!g2076) & (g2077)) + ((g2490) & (!g2296) & (g2402) & (g2183) & (g2076) & (g2077)) + ((g2490) & (g2296) & (!g2402) & (!g2183) & (!g2076) & (!g2077)) + ((g2490) & (g2296) & (!g2402) & (!g2183) & (g2076) & (!g2077)) + ((g2490) & (g2296) & (!g2402) & (g2183) & (!g2076) & (!g2077)) + ((g2490) & (g2296) & (!g2402) & (g2183) & (g2076) & (!g2077)) + ((g2490) & (g2296) & (!g2402) & (g2183) & (g2076) & (g2077)) + ((g2490) & (g2296) & (g2402) & (!g2183) & (!g2076) & (!g2077)) + ((g2490) & (g2296) & (g2402) & (!g2183) & (!g2076) & (g2077)) + ((g2490) & (g2296) & (g2402) & (!g2183) & (g2076) & (!g2077)) + ((g2490) & (g2296) & (g2402) & (g2183) & (!g2076) & (!g2077)) + ((g2490) & (g2296) & (g2402) & (g2183) & (!g2076) & (g2077)) + ((g2490) & (g2296) & (g2402) & (g2183) & (g2076) & (!g2077)) + ((g2490) & (g2296) & (g2402) & (g2183) & (g2076) & (g2077)));
	assign g2492 = (((!g2200) & (!g2189) & (!g2187) & (g2188) & (g2076) & (g2077)) + ((!g2200) & (!g2189) & (g2187) & (!g2188) & (!g2076) & (g2077)) + ((!g2200) & (!g2189) & (g2187) & (g2188) & (!g2076) & (g2077)) + ((!g2200) & (!g2189) & (g2187) & (g2188) & (g2076) & (g2077)) + ((!g2200) & (g2189) & (!g2187) & (!g2188) & (g2076) & (!g2077)) + ((!g2200) & (g2189) & (!g2187) & (g2188) & (g2076) & (!g2077)) + ((!g2200) & (g2189) & (!g2187) & (g2188) & (g2076) & (g2077)) + ((!g2200) & (g2189) & (g2187) & (!g2188) & (!g2076) & (g2077)) + ((!g2200) & (g2189) & (g2187) & (!g2188) & (g2076) & (!g2077)) + ((!g2200) & (g2189) & (g2187) & (g2188) & (!g2076) & (g2077)) + ((!g2200) & (g2189) & (g2187) & (g2188) & (g2076) & (!g2077)) + ((!g2200) & (g2189) & (g2187) & (g2188) & (g2076) & (g2077)) + ((g2200) & (!g2189) & (!g2187) & (!g2188) & (!g2076) & (!g2077)) + ((g2200) & (!g2189) & (!g2187) & (g2188) & (!g2076) & (!g2077)) + ((g2200) & (!g2189) & (!g2187) & (g2188) & (g2076) & (g2077)) + ((g2200) & (!g2189) & (g2187) & (!g2188) & (!g2076) & (!g2077)) + ((g2200) & (!g2189) & (g2187) & (!g2188) & (!g2076) & (g2077)) + ((g2200) & (!g2189) & (g2187) & (g2188) & (!g2076) & (!g2077)) + ((g2200) & (!g2189) & (g2187) & (g2188) & (!g2076) & (g2077)) + ((g2200) & (!g2189) & (g2187) & (g2188) & (g2076) & (g2077)) + ((g2200) & (g2189) & (!g2187) & (!g2188) & (!g2076) & (!g2077)) + ((g2200) & (g2189) & (!g2187) & (!g2188) & (g2076) & (!g2077)) + ((g2200) & (g2189) & (!g2187) & (g2188) & (!g2076) & (!g2077)) + ((g2200) & (g2189) & (!g2187) & (g2188) & (g2076) & (!g2077)) + ((g2200) & (g2189) & (!g2187) & (g2188) & (g2076) & (g2077)) + ((g2200) & (g2189) & (g2187) & (!g2188) & (!g2076) & (!g2077)) + ((g2200) & (g2189) & (g2187) & (!g2188) & (!g2076) & (g2077)) + ((g2200) & (g2189) & (g2187) & (!g2188) & (g2076) & (!g2077)) + ((g2200) & (g2189) & (g2187) & (g2188) & (!g2076) & (!g2077)) + ((g2200) & (g2189) & (g2187) & (g2188) & (!g2076) & (g2077)) + ((g2200) & (g2189) & (g2187) & (g2188) & (g2076) & (!g2077)) + ((g2200) & (g2189) & (g2187) & (g2188) & (g2076) & (g2077)));
	assign g2493 = (((!g2399) & (!g2400) & (!sk[70]) & (!g2489) & (g2491) & (!g2492)) + ((!g2399) & (!g2400) & (!sk[70]) & (!g2489) & (g2491) & (g2492)) + ((!g2399) & (!g2400) & (!sk[70]) & (g2489) & (!g2491) & (!g2492)) + ((!g2399) & (!g2400) & (!sk[70]) & (g2489) & (!g2491) & (g2492)) + ((!g2399) & (!g2400) & (!sk[70]) & (g2489) & (g2491) & (!g2492)) + ((!g2399) & (!g2400) & (!sk[70]) & (g2489) & (g2491) & (g2492)) + ((!g2399) & (!g2400) & (sk[70]) & (!g2489) & (g2491) & (!g2492)) + ((!g2399) & (!g2400) & (sk[70]) & (!g2489) & (g2491) & (g2492)) + ((!g2399) & (!g2400) & (sk[70]) & (g2489) & (g2491) & (!g2492)) + ((!g2399) & (!g2400) & (sk[70]) & (g2489) & (g2491) & (g2492)) + ((!g2399) & (g2400) & (!sk[70]) & (!g2489) & (!g2491) & (!g2492)) + ((!g2399) & (g2400) & (!sk[70]) & (!g2489) & (!g2491) & (g2492)) + ((!g2399) & (g2400) & (!sk[70]) & (!g2489) & (g2491) & (!g2492)) + ((!g2399) & (g2400) & (!sk[70]) & (!g2489) & (g2491) & (g2492)) + ((!g2399) & (g2400) & (!sk[70]) & (g2489) & (!g2491) & (!g2492)) + ((!g2399) & (g2400) & (!sk[70]) & (g2489) & (!g2491) & (g2492)) + ((!g2399) & (g2400) & (!sk[70]) & (g2489) & (g2491) & (!g2492)) + ((!g2399) & (g2400) & (!sk[70]) & (g2489) & (g2491) & (g2492)) + ((!g2399) & (g2400) & (sk[70]) & (g2489) & (!g2491) & (!g2492)) + ((!g2399) & (g2400) & (sk[70]) & (g2489) & (!g2491) & (g2492)) + ((!g2399) & (g2400) & (sk[70]) & (g2489) & (g2491) & (!g2492)) + ((!g2399) & (g2400) & (sk[70]) & (g2489) & (g2491) & (g2492)) + ((g2399) & (!g2400) & (!sk[70]) & (!g2489) & (g2491) & (!g2492)) + ((g2399) & (!g2400) & (!sk[70]) & (!g2489) & (g2491) & (g2492)) + ((g2399) & (!g2400) & (!sk[70]) & (g2489) & (!g2491) & (!g2492)) + ((g2399) & (!g2400) & (!sk[70]) & (g2489) & (!g2491) & (g2492)) + ((g2399) & (!g2400) & (!sk[70]) & (g2489) & (g2491) & (!g2492)) + ((g2399) & (!g2400) & (!sk[70]) & (g2489) & (g2491) & (g2492)) + ((g2399) & (!g2400) & (sk[70]) & (!g2489) & (!g2491) & (g2492)) + ((g2399) & (!g2400) & (sk[70]) & (!g2489) & (g2491) & (g2492)) + ((g2399) & (!g2400) & (sk[70]) & (g2489) & (!g2491) & (g2492)) + ((g2399) & (!g2400) & (sk[70]) & (g2489) & (g2491) & (g2492)) + ((g2399) & (g2400) & (!sk[70]) & (!g2489) & (!g2491) & (!g2492)) + ((g2399) & (g2400) & (!sk[70]) & (!g2489) & (!g2491) & (g2492)) + ((g2399) & (g2400) & (!sk[70]) & (!g2489) & (g2491) & (!g2492)) + ((g2399) & (g2400) & (!sk[70]) & (!g2489) & (g2491) & (g2492)) + ((g2399) & (g2400) & (!sk[70]) & (g2489) & (!g2491) & (!g2492)) + ((g2399) & (g2400) & (!sk[70]) & (g2489) & (!g2491) & (g2492)) + ((g2399) & (g2400) & (!sk[70]) & (g2489) & (g2491) & (!g2492)) + ((g2399) & (g2400) & (!sk[70]) & (g2489) & (g2491) & (g2492)));
	assign g2494 = (((!g2482) & (!g2119) & (!g2124) & (!g2264) & (!g3588) & (!g2493)) + ((!g2482) & (!g2119) & (!g2124) & (!g2264) & (g3588) & (!g2493)) + ((!g2482) & (!g2119) & (!g2124) & (g2264) & (!g3588) & (!g2493)) + ((!g2482) & (!g2119) & (!g2124) & (g2264) & (!g3588) & (g2493)) + ((!g2482) & (!g2119) & (g2124) & (!g2264) & (!g3588) & (!g2493)) + ((!g2482) & (!g2119) & (g2124) & (!g2264) & (!g3588) & (g2493)) + ((!g2482) & (!g2119) & (g2124) & (!g2264) & (g3588) & (!g2493)) + ((!g2482) & (!g2119) & (g2124) & (!g2264) & (g3588) & (g2493)) + ((!g2482) & (!g2119) & (g2124) & (g2264) & (!g3588) & (!g2493)) + ((!g2482) & (!g2119) & (g2124) & (g2264) & (!g3588) & (g2493)) + ((!g2482) & (!g2119) & (g2124) & (g2264) & (g3588) & (!g2493)) + ((!g2482) & (!g2119) & (g2124) & (g2264) & (g3588) & (g2493)) + ((!g2482) & (g2119) & (!g2124) & (!g2264) & (!g3588) & (!g2493)) + ((!g2482) & (g2119) & (!g2124) & (!g2264) & (g3588) & (!g2493)) + ((!g2482) & (g2119) & (!g2124) & (g2264) & (!g3588) & (!g2493)) + ((!g2482) & (g2119) & (!g2124) & (g2264) & (!g3588) & (g2493)) + ((g2482) & (!g2119) & (!g2124) & (!g2264) & (!g3588) & (!g2493)) + ((g2482) & (!g2119) & (!g2124) & (!g2264) & (g3588) & (!g2493)) + ((g2482) & (!g2119) & (!g2124) & (g2264) & (!g3588) & (!g2493)) + ((g2482) & (!g2119) & (!g2124) & (g2264) & (!g3588) & (g2493)) + ((g2482) & (g2119) & (!g2124) & (!g2264) & (!g3588) & (!g2493)) + ((g2482) & (g2119) & (!g2124) & (!g2264) & (g3588) & (!g2493)) + ((g2482) & (g2119) & (!g2124) & (g2264) & (!g3588) & (!g2493)) + ((g2482) & (g2119) & (!g2124) & (g2264) & (!g3588) & (g2493)) + ((g2482) & (g2119) & (g2124) & (g2264) & (!g3588) & (!g2493)) + ((g2482) & (g2119) & (g2124) & (g2264) & (!g3588) & (g2493)) + ((g2482) & (g2119) & (g2124) & (g2264) & (g3588) & (!g2493)) + ((g2482) & (g2119) & (g2124) & (g2264) & (g3588) & (g2493)));
	assign g2495 = (((!g75) & (!g2119) & (!g2280) & (!g2480) & (!g2481) & (!g2494)) + ((!g75) & (!g2119) & (!g2280) & (!g2480) & (g2481) & (!g2494)) + ((!g75) & (!g2119) & (!g2280) & (g2480) & (!g2481) & (!g2494)) + ((!g75) & (!g2119) & (!g2280) & (g2480) & (g2481) & (!g2494)) + ((!g75) & (g2119) & (!g2280) & (!g2480) & (!g2481) & (!g2494)) + ((!g75) & (g2119) & (!g2280) & (!g2480) & (g2481) & (!g2494)) + ((!g75) & (g2119) & (!g2280) & (g2480) & (!g2481) & (!g2494)) + ((!g75) & (g2119) & (!g2280) & (g2480) & (g2481) & (!g2494)) + ((!g75) & (g2119) & (g2280) & (!g2480) & (!g2481) & (!g2494)) + ((!g75) & (g2119) & (g2280) & (!g2480) & (!g2481) & (g2494)) + ((!g75) & (g2119) & (g2280) & (!g2480) & (g2481) & (!g2494)) + ((!g75) & (g2119) & (g2280) & (!g2480) & (g2481) & (g2494)) + ((!g75) & (g2119) & (g2280) & (g2480) & (!g2481) & (!g2494)) + ((!g75) & (g2119) & (g2280) & (g2480) & (!g2481) & (g2494)) + ((!g75) & (g2119) & (g2280) & (g2480) & (g2481) & (!g2494)) + ((!g75) & (g2119) & (g2280) & (g2480) & (g2481) & (g2494)) + ((g75) & (!g2119) & (!g2280) & (!g2480) & (g2481) & (!g2494)) + ((g75) & (!g2119) & (!g2280) & (!g2480) & (g2481) & (g2494)) + ((g75) & (!g2119) & (!g2280) & (g2480) & (!g2481) & (!g2494)) + ((g75) & (!g2119) & (!g2280) & (g2480) & (!g2481) & (g2494)) + ((g75) & (!g2119) & (!g2280) & (g2480) & (g2481) & (!g2494)) + ((g75) & (!g2119) & (!g2280) & (g2480) & (g2481) & (g2494)) + ((g75) & (!g2119) & (g2280) & (!g2480) & (g2481) & (!g2494)) + ((g75) & (!g2119) & (g2280) & (!g2480) & (g2481) & (g2494)) + ((g75) & (!g2119) & (g2280) & (g2480) & (!g2481) & (!g2494)) + ((g75) & (!g2119) & (g2280) & (g2480) & (!g2481) & (g2494)) + ((g75) & (!g2119) & (g2280) & (g2480) & (g2481) & (!g2494)) + ((g75) & (!g2119) & (g2280) & (g2480) & (g2481) & (g2494)) + ((g75) & (g2119) & (!g2280) & (!g2480) & (g2481) & (!g2494)) + ((g75) & (g2119) & (!g2280) & (!g2480) & (g2481) & (g2494)) + ((g75) & (g2119) & (!g2280) & (g2480) & (!g2481) & (!g2494)) + ((g75) & (g2119) & (!g2280) & (g2480) & (!g2481) & (g2494)) + ((g75) & (g2119) & (!g2280) & (g2480) & (g2481) & (!g2494)) + ((g75) & (g2119) & (!g2280) & (g2480) & (g2481) & (g2494)) + ((g75) & (g2119) & (g2280) & (!g2480) & (g2481) & (!g2494)) + ((g75) & (g2119) & (g2280) & (!g2480) & (g2481) & (g2494)) + ((g75) & (g2119) & (g2280) & (g2480) & (!g2481) & (!g2494)) + ((g75) & (g2119) & (g2280) & (g2480) & (!g2481) & (g2494)) + ((g75) & (g2119) & (g2280) & (g2480) & (g2481) & (!g2494)) + ((g75) & (g2119) & (g2280) & (g2480) & (g2481) & (g2494)));
	assign g2496 = (((!g630) & (!g587) & (!sk[73]) & (!g2409) & (g724)) + ((!g630) & (!g587) & (!sk[73]) & (g2409) & (!g724)) + ((!g630) & (!g587) & (!sk[73]) & (g2409) & (g724)) + ((!g630) & (g587) & (!sk[73]) & (!g2409) & (!g724)) + ((!g630) & (g587) & (!sk[73]) & (!g2409) & (g724)) + ((!g630) & (g587) & (!sk[73]) & (g2409) & (!g724)) + ((!g630) & (g587) & (!sk[73]) & (g2409) & (g724)) + ((g630) & (!g587) & (!sk[73]) & (!g2409) & (g724)) + ((g630) & (!g587) & (!sk[73]) & (g2409) & (!g724)) + ((g630) & (!g587) & (!sk[73]) & (g2409) & (g724)) + ((g630) & (g587) & (!sk[73]) & (!g2409) & (!g724)) + ((g630) & (g587) & (!sk[73]) & (!g2409) & (g724)) + ((g630) & (g587) & (!sk[73]) & (g2409) & (!g724)) + ((g630) & (g587) & (!sk[73]) & (g2409) & (g724)) + ((g630) & (g587) & (sk[73]) & (g2409) & (g724)));
	assign g2497 = (((!sk[74]) & (g771) & (!g2496)) + ((!sk[74]) & (g771) & (g2496)) + ((sk[74]) & (!g771) & (g2496)) + ((sk[74]) & (g771) & (!g2496)));
	assign g2498 = (((!sk[75]) & (!g1772) & (!g2033) & (g2034)) + ((!sk[75]) & (!g1772) & (g2033) & (!g2034)) + ((!sk[75]) & (!g1772) & (g2033) & (g2034)) + ((!sk[75]) & (g1772) & (!g2033) & (g2034)) + ((!sk[75]) & (g1772) & (g2033) & (!g2034)) + ((!sk[75]) & (g1772) & (g2033) & (g2034)) + ((sk[75]) & (g1772) & (!g2033) & (g2034)));
	assign g5037 = (((!g2921) & (!g3080) & (!sk[76]) & (g2499)) + ((!g2921) & (!g3080) & (sk[76]) & (g2499)) + ((!g2921) & (g3080) & (!sk[76]) & (!g2499)) + ((!g2921) & (g3080) & (!sk[76]) & (g2499)) + ((!g2921) & (g3080) & (sk[76]) & (g2499)) + ((g2921) & (!g3080) & (!sk[76]) & (g2499)) + ((g2921) & (g3080) & (!sk[76]) & (!g2499)) + ((g2921) & (g3080) & (!sk[76]) & (g2499)) + ((g2921) & (g3080) & (sk[76]) & (!g2499)) + ((g2921) & (g3080) & (sk[76]) & (g2499)));
	assign g2500 = (((!g91) & (!g630) & (!sk[77]) & (!g586) & (g2433) & (!g724)) + ((!g91) & (!g630) & (!sk[77]) & (!g586) & (g2433) & (g724)) + ((!g91) & (!g630) & (!sk[77]) & (g586) & (!g2433) & (!g724)) + ((!g91) & (!g630) & (!sk[77]) & (g586) & (!g2433) & (g724)) + ((!g91) & (!g630) & (!sk[77]) & (g586) & (g2433) & (!g724)) + ((!g91) & (!g630) & (!sk[77]) & (g586) & (g2433) & (g724)) + ((!g91) & (g630) & (!sk[77]) & (!g586) & (!g2433) & (!g724)) + ((!g91) & (g630) & (!sk[77]) & (!g586) & (!g2433) & (g724)) + ((!g91) & (g630) & (!sk[77]) & (!g586) & (g2433) & (!g724)) + ((!g91) & (g630) & (!sk[77]) & (!g586) & (g2433) & (g724)) + ((!g91) & (g630) & (!sk[77]) & (g586) & (!g2433) & (!g724)) + ((!g91) & (g630) & (!sk[77]) & (g586) & (!g2433) & (g724)) + ((!g91) & (g630) & (!sk[77]) & (g586) & (g2433) & (!g724)) + ((!g91) & (g630) & (!sk[77]) & (g586) & (g2433) & (g724)) + ((!g91) & (g630) & (sk[77]) & (!g586) & (g2433) & (g724)) + ((!g91) & (g630) & (sk[77]) & (g586) & (g2433) & (!g724)) + ((g91) & (!g630) & (!sk[77]) & (!g586) & (g2433) & (!g724)) + ((g91) & (!g630) & (!sk[77]) & (!g586) & (g2433) & (g724)) + ((g91) & (!g630) & (!sk[77]) & (g586) & (!g2433) & (!g724)) + ((g91) & (!g630) & (!sk[77]) & (g586) & (!g2433) & (g724)) + ((g91) & (!g630) & (!sk[77]) & (g586) & (g2433) & (!g724)) + ((g91) & (!g630) & (!sk[77]) & (g586) & (g2433) & (g724)) + ((g91) & (!g630) & (sk[77]) & (!g586) & (g2433) & (g724)) + ((g91) & (!g630) & (sk[77]) & (g586) & (g2433) & (!g724)) + ((g91) & (g630) & (!sk[77]) & (!g586) & (!g2433) & (!g724)) + ((g91) & (g630) & (!sk[77]) & (!g586) & (!g2433) & (g724)) + ((g91) & (g630) & (!sk[77]) & (!g586) & (g2433) & (!g724)) + ((g91) & (g630) & (!sk[77]) & (!g586) & (g2433) & (g724)) + ((g91) & (g630) & (!sk[77]) & (g586) & (!g2433) & (!g724)) + ((g91) & (g630) & (!sk[77]) & (g586) & (!g2433) & (g724)) + ((g91) & (g630) & (!sk[77]) & (g586) & (g2433) & (!g724)) + ((g91) & (g630) & (!sk[77]) & (g586) & (g2433) & (g724)) + ((g91) & (g630) & (sk[77]) & (!g586) & (!g2433) & (g724)) + ((g91) & (g630) & (sk[77]) & (!g586) & (g2433) & (g724)) + ((g91) & (g630) & (sk[77]) & (g586) & (!g2433) & (!g724)) + ((g91) & (g630) & (sk[77]) & (g586) & (g2433) & (!g724)));
	assign g2501 = (((g586) & (!sk[78]) & (!g724)) + ((g586) & (!sk[78]) & (g724)) + ((g586) & (sk[78]) & (g724)));
	assign g2502 = (((!g2500) & (sk[79]) & (!g2501)) + ((g2500) & (!sk[79]) & (!g2501)) + ((g2500) & (!sk[79]) & (g2501)));
	assign g2503 = (((!g677) & (!g2033) & (!g2034) & (!g771) & (g2499) & (!g2502)) + ((!g677) & (!g2033) & (!g2034) & (!g771) & (g2499) & (g2502)) + ((!g677) & (!g2033) & (!g2034) & (g771) & (g2499) & (!g2502)) + ((!g677) & (!g2033) & (!g2034) & (g771) & (g2499) & (g2502)) + ((!g677) & (g2033) & (!g2034) & (!g771) & (!g2499) & (!g2502)) + ((!g677) & (g2033) & (!g2034) & (!g771) & (g2499) & (!g2502)) + ((!g677) & (g2033) & (!g2034) & (g771) & (!g2499) & (g2502)) + ((!g677) & (g2033) & (!g2034) & (g771) & (g2499) & (g2502)) + ((g677) & (!g2033) & (!g2034) & (!g771) & (g2499) & (!g2502)) + ((g677) & (!g2033) & (!g2034) & (!g771) & (g2499) & (g2502)) + ((g677) & (!g2033) & (!g2034) & (g771) & (g2499) & (!g2502)) + ((g677) & (!g2033) & (!g2034) & (g771) & (g2499) & (g2502)) + ((g677) & (g2033) & (!g2034) & (!g771) & (!g2499) & (g2502)) + ((g677) & (g2033) & (!g2034) & (!g771) & (g2499) & (g2502)) + ((g677) & (g2033) & (!g2034) & (g771) & (!g2499) & (!g2502)) + ((g677) & (g2033) & (!g2034) & (g771) & (g2499) & (!g2502)));
	assign g2504 = (((g2329) & (!g2029) & (g2408) & (!g2497) & (!g2498) & (g2503)) + ((g2329) & (!g2029) & (g2408) & (!g2497) & (g2498) & (!g2503)) + ((g2329) & (!g2029) & (g2408) & (!g2497) & (g2498) & (g2503)) + ((g2329) & (!g2029) & (g2408) & (g2497) & (!g2498) & (g2503)) + ((g2329) & (!g2029) & (g2408) & (g2497) & (g2498) & (!g2503)) + ((g2329) & (!g2029) & (g2408) & (g2497) & (g2498) & (g2503)) + ((g2329) & (g2029) & (g2408) & (g2497) & (!g2498) & (!g2503)) + ((g2329) & (g2029) & (g2408) & (g2497) & (!g2498) & (g2503)) + ((g2329) & (g2029) & (g2408) & (g2497) & (g2498) & (!g2503)) + ((g2329) & (g2029) & (g2408) & (g2497) & (g2498) & (g2503)));
	assign g2505 = (((g2131) & (g2132) & (!dmem_dat_ix30x) & (!g2128) & (g2129) & (dmem_dat_ix14x)) + ((g2131) & (g2132) & (dmem_dat_ix30x) & (!g2128) & (!g2129) & (!dmem_dat_ix14x)) + ((g2131) & (g2132) & (dmem_dat_ix30x) & (!g2128) & (!g2129) & (dmem_dat_ix14x)) + ((g2131) & (g2132) & (dmem_dat_ix30x) & (!g2128) & (g2129) & (dmem_dat_ix14x)));
	assign g2506 = (((!g2363) & (!g2131) & (!g2132) & (dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((!g2363) & (!g2131) & (!g2132) & (dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((!g2363) & (!g2131) & (g2132) & (!dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((!g2363) & (!g2131) & (g2132) & (!dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((!g2363) & (!g2131) & (g2132) & (dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((!g2363) & (!g2131) & (g2132) & (dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((!g2363) & (g2131) & (!g2132) & (!dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((!g2363) & (g2131) & (!g2132) & (!dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((!g2363) & (g2131) & (!g2132) & (dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((!g2363) & (g2131) & (!g2132) & (dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((!g2363) & (g2131) & (!g2132) & (dmem_dat_ix14x) & (sk[83]) & (!g2338)) + ((!g2363) & (g2131) & (!g2132) & (dmem_dat_ix14x) & (sk[83]) & (g2338)) + ((!g2363) & (g2131) & (g2132) & (!dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((!g2363) & (g2131) & (g2132) & (!dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((!g2363) & (g2131) & (g2132) & (dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((!g2363) & (g2131) & (g2132) & (dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((g2363) & (!g2131) & (!g2132) & (!dmem_dat_ix14x) & (sk[83]) & (g2338)) + ((g2363) & (!g2131) & (!g2132) & (dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((g2363) & (!g2131) & (!g2132) & (dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((g2363) & (!g2131) & (!g2132) & (dmem_dat_ix14x) & (sk[83]) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (!dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((g2363) & (!g2131) & (g2132) & (!dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (!dmem_dat_ix14x) & (sk[83]) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((g2363) & (!g2131) & (g2132) & (dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((g2363) & (!g2131) & (g2132) & (dmem_dat_ix14x) & (sk[83]) & (g2338)) + ((g2363) & (g2131) & (!g2132) & (!dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((g2363) & (g2131) & (!g2132) & (!dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((g2363) & (g2131) & (!g2132) & (dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((g2363) & (g2131) & (!g2132) & (dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((g2363) & (g2131) & (!g2132) & (dmem_dat_ix14x) & (sk[83]) & (!g2338)) + ((g2363) & (g2131) & (!g2132) & (dmem_dat_ix14x) & (sk[83]) & (g2338)) + ((g2363) & (g2131) & (g2132) & (!dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((g2363) & (g2131) & (g2132) & (!dmem_dat_ix14x) & (!sk[83]) & (g2338)) + ((g2363) & (g2131) & (g2132) & (dmem_dat_ix14x) & (!sk[83]) & (!g2338)) + ((g2363) & (g2131) & (g2132) & (dmem_dat_ix14x) & (!sk[83]) & (g2338)));
	assign g2508 = (((!g2119) & (!g2120) & (!sk[84]) & (!g2482) & (g2483) & (!g2507)) + ((!g2119) & (!g2120) & (!sk[84]) & (!g2482) & (g2483) & (g2507)) + ((!g2119) & (!g2120) & (!sk[84]) & (g2482) & (!g2483) & (!g2507)) + ((!g2119) & (!g2120) & (!sk[84]) & (g2482) & (!g2483) & (g2507)) + ((!g2119) & (!g2120) & (!sk[84]) & (g2482) & (g2483) & (!g2507)) + ((!g2119) & (!g2120) & (!sk[84]) & (g2482) & (g2483) & (g2507)) + ((!g2119) & (!g2120) & (sk[84]) & (!g2482) & (!g2483) & (g2507)) + ((!g2119) & (!g2120) & (sk[84]) & (!g2482) & (g2483) & (g2507)) + ((!g2119) & (!g2120) & (sk[84]) & (g2482) & (!g2483) & (g2507)) + ((!g2119) & (!g2120) & (sk[84]) & (g2482) & (g2483) & (!g2507)) + ((!g2119) & (g2120) & (!sk[84]) & (!g2482) & (!g2483) & (!g2507)) + ((!g2119) & (g2120) & (!sk[84]) & (!g2482) & (!g2483) & (g2507)) + ((!g2119) & (g2120) & (!sk[84]) & (!g2482) & (g2483) & (!g2507)) + ((!g2119) & (g2120) & (!sk[84]) & (!g2482) & (g2483) & (g2507)) + ((!g2119) & (g2120) & (!sk[84]) & (g2482) & (!g2483) & (!g2507)) + ((!g2119) & (g2120) & (!sk[84]) & (g2482) & (!g2483) & (g2507)) + ((!g2119) & (g2120) & (!sk[84]) & (g2482) & (g2483) & (!g2507)) + ((!g2119) & (g2120) & (!sk[84]) & (g2482) & (g2483) & (g2507)) + ((!g2119) & (g2120) & (sk[84]) & (!g2482) & (!g2483) & (!g2507)) + ((!g2119) & (g2120) & (sk[84]) & (!g2482) & (g2483) & (!g2507)) + ((!g2119) & (g2120) & (sk[84]) & (g2482) & (!g2483) & (!g2507)) + ((!g2119) & (g2120) & (sk[84]) & (g2482) & (g2483) & (g2507)) + ((g2119) & (!g2120) & (!sk[84]) & (!g2482) & (g2483) & (!g2507)) + ((g2119) & (!g2120) & (!sk[84]) & (!g2482) & (g2483) & (g2507)) + ((g2119) & (!g2120) & (!sk[84]) & (g2482) & (!g2483) & (!g2507)) + ((g2119) & (!g2120) & (!sk[84]) & (g2482) & (!g2483) & (g2507)) + ((g2119) & (!g2120) & (!sk[84]) & (g2482) & (g2483) & (!g2507)) + ((g2119) & (!g2120) & (!sk[84]) & (g2482) & (g2483) & (g2507)) + ((g2119) & (!g2120) & (sk[84]) & (!g2482) & (!g2483) & (g2507)) + ((g2119) & (!g2120) & (sk[84]) & (!g2482) & (g2483) & (!g2507)) + ((g2119) & (!g2120) & (sk[84]) & (g2482) & (!g2483) & (!g2507)) + ((g2119) & (!g2120) & (sk[84]) & (g2482) & (g2483) & (!g2507)) + ((g2119) & (g2120) & (!sk[84]) & (!g2482) & (!g2483) & (!g2507)) + ((g2119) & (g2120) & (!sk[84]) & (!g2482) & (!g2483) & (g2507)) + ((g2119) & (g2120) & (!sk[84]) & (!g2482) & (g2483) & (!g2507)) + ((g2119) & (g2120) & (!sk[84]) & (!g2482) & (g2483) & (g2507)) + ((g2119) & (g2120) & (!sk[84]) & (g2482) & (!g2483) & (!g2507)) + ((g2119) & (g2120) & (!sk[84]) & (g2482) & (!g2483) & (g2507)) + ((g2119) & (g2120) & (!sk[84]) & (g2482) & (g2483) & (!g2507)) + ((g2119) & (g2120) & (!sk[84]) & (g2482) & (g2483) & (g2507)) + ((g2119) & (g2120) & (sk[84]) & (!g2482) & (!g2483) & (!g2507)) + ((g2119) & (g2120) & (sk[84]) & (!g2482) & (g2483) & (g2507)) + ((g2119) & (g2120) & (sk[84]) & (g2482) & (!g2483) & (g2507)) + ((g2119) & (g2120) & (sk[84]) & (g2482) & (g2483) & (g2507)));
	assign g2509 = (((!g2461) & (!g2462) & (!g2464) & (!g2465) & (!g2486) & (!g2487)) + ((!g2461) & (!g2462) & (!g2464) & (!g2465) & (!g2486) & (g2487)) + ((!g2461) & (!g2462) & (!g2464) & (!g2465) & (g2486) & (!g2487)) + ((!g2461) & (!g2462) & (!g2464) & (g2465) & (!g2486) & (!g2487)) + ((!g2461) & (!g2462) & (!g2464) & (g2465) & (!g2486) & (g2487)) + ((!g2461) & (!g2462) & (!g2464) & (g2465) & (g2486) & (!g2487)) + ((!g2461) & (!g2462) & (g2464) & (!g2465) & (!g2486) & (!g2487)) + ((!g2461) & (!g2462) & (g2464) & (!g2465) & (!g2486) & (g2487)) + ((!g2461) & (!g2462) & (g2464) & (!g2465) & (g2486) & (!g2487)) + ((!g2461) & (!g2462) & (g2464) & (g2465) & (!g2486) & (!g2487)) + ((!g2461) & (g2462) & (!g2464) & (!g2465) & (!g2486) & (!g2487)) + ((!g2461) & (g2462) & (!g2464) & (!g2465) & (!g2486) & (g2487)) + ((!g2461) & (g2462) & (!g2464) & (!g2465) & (g2486) & (!g2487)) + ((!g2461) & (g2462) & (!g2464) & (g2465) & (!g2486) & (!g2487)) + ((!g2461) & (g2462) & (g2464) & (!g2465) & (!g2486) & (!g2487)) + ((!g2461) & (g2462) & (g2464) & (g2465) & (!g2486) & (!g2487)) + ((g2461) & (!g2462) & (!g2464) & (!g2465) & (!g2486) & (!g2487)) + ((g2461) & (!g2462) & (!g2464) & (!g2465) & (!g2486) & (g2487)) + ((g2461) & (!g2462) & (!g2464) & (!g2465) & (g2486) & (!g2487)) + ((g2461) & (!g2462) & (!g2464) & (g2465) & (!g2486) & (!g2487)) + ((g2461) & (!g2462) & (g2464) & (!g2465) & (!g2486) & (!g2487)) + ((g2461) & (!g2462) & (g2464) & (g2465) & (!g2486) & (!g2487)) + ((g2461) & (g2462) & (!g2464) & (!g2465) & (!g2486) & (!g2487)) + ((g2461) & (g2462) & (!g2464) & (!g2465) & (!g2486) & (g2487)) + ((g2461) & (g2462) & (!g2464) & (!g2465) & (g2486) & (!g2487)) + ((g2461) & (g2462) & (!g2464) & (g2465) & (!g2486) & (!g2487)) + ((g2461) & (g2462) & (g2464) & (!g2465) & (!g2486) & (!g2487)) + ((g2461) & (g2462) & (g2464) & (g2465) & (!g2486) & (!g2487)));
	assign g2510 = (((g2119) & (!sk[86]) & (!g2482)) + ((g2119) & (!sk[86]) & (g2482)) + ((g2119) & (sk[86]) & (!g2482)));
	assign g2511 = (((!sk[87]) & (g2120) & (!g2507)) + ((!sk[87]) & (g2120) & (g2507)) + ((sk[87]) & (!g2120) & (!g2507)) + ((sk[87]) & (g2120) & (g2507)));
	assign g2512 = (((!g2509) & (!g2510) & (!sk[88]) & (g2511)) + ((!g2509) & (!g2510) & (sk[88]) & (!g2511)) + ((!g2509) & (g2510) & (!sk[88]) & (!g2511)) + ((!g2509) & (g2510) & (!sk[88]) & (g2511)) + ((!g2509) & (g2510) & (sk[88]) & (g2511)) + ((g2509) & (!g2510) & (!sk[88]) & (g2511)) + ((g2509) & (!g2510) & (sk[88]) & (g2511)) + ((g2509) & (g2510) & (!sk[88]) & (!g2511)) + ((g2509) & (g2510) & (!sk[88]) & (g2511)) + ((g2509) & (g2510) & (sk[88]) & (!g2511)));
	assign g2513 = (((!sk[89]) & (g2120) & (!g2507)) + ((!sk[89]) & (g2120) & (g2507)) + ((sk[89]) & (g2120) & (g2507)));
	assign g2514 = (((!g2120) & (!g2119) & (!g2118) & (g2111) & (g2071) & (g2074)) + ((!g2120) & (!g2119) & (g2118) & (!g2111) & (!g2071) & (g2074)) + ((!g2120) & (!g2119) & (g2118) & (g2111) & (!g2071) & (g2074)) + ((!g2120) & (!g2119) & (g2118) & (g2111) & (g2071) & (g2074)) + ((!g2120) & (g2119) & (!g2118) & (!g2111) & (g2071) & (!g2074)) + ((!g2120) & (g2119) & (!g2118) & (g2111) & (g2071) & (!g2074)) + ((!g2120) & (g2119) & (!g2118) & (g2111) & (g2071) & (g2074)) + ((!g2120) & (g2119) & (g2118) & (!g2111) & (!g2071) & (g2074)) + ((!g2120) & (g2119) & (g2118) & (!g2111) & (g2071) & (!g2074)) + ((!g2120) & (g2119) & (g2118) & (g2111) & (!g2071) & (g2074)) + ((!g2120) & (g2119) & (g2118) & (g2111) & (g2071) & (!g2074)) + ((!g2120) & (g2119) & (g2118) & (g2111) & (g2071) & (g2074)) + ((g2120) & (!g2119) & (!g2118) & (!g2111) & (!g2071) & (!g2074)) + ((g2120) & (!g2119) & (!g2118) & (g2111) & (!g2071) & (!g2074)) + ((g2120) & (!g2119) & (!g2118) & (g2111) & (g2071) & (g2074)) + ((g2120) & (!g2119) & (g2118) & (!g2111) & (!g2071) & (!g2074)) + ((g2120) & (!g2119) & (g2118) & (!g2111) & (!g2071) & (g2074)) + ((g2120) & (!g2119) & (g2118) & (g2111) & (!g2071) & (!g2074)) + ((g2120) & (!g2119) & (g2118) & (g2111) & (!g2071) & (g2074)) + ((g2120) & (!g2119) & (g2118) & (g2111) & (g2071) & (g2074)) + ((g2120) & (g2119) & (!g2118) & (!g2111) & (!g2071) & (!g2074)) + ((g2120) & (g2119) & (!g2118) & (!g2111) & (g2071) & (!g2074)) + ((g2120) & (g2119) & (!g2118) & (g2111) & (!g2071) & (!g2074)) + ((g2120) & (g2119) & (!g2118) & (g2111) & (g2071) & (!g2074)) + ((g2120) & (g2119) & (!g2118) & (g2111) & (g2071) & (g2074)) + ((g2120) & (g2119) & (g2118) & (!g2111) & (!g2071) & (!g2074)) + ((g2120) & (g2119) & (g2118) & (!g2111) & (!g2071) & (g2074)) + ((g2120) & (g2119) & (g2118) & (!g2111) & (g2071) & (!g2074)) + ((g2120) & (g2119) & (g2118) & (g2111) & (!g2071) & (!g2074)) + ((g2120) & (g2119) & (g2118) & (g2111) & (!g2071) & (g2074)) + ((g2120) & (g2119) & (g2118) & (g2111) & (g2071) & (!g2074)) + ((g2120) & (g2119) & (g2118) & (g2111) & (g2071) & (g2074)));
	assign g2515 = (((!g2514) & (!g2320) & (!g2426) & (g2211) & (g2076) & (g2077)) + ((!g2514) & (!g2320) & (g2426) & (!g2211) & (!g2076) & (g2077)) + ((!g2514) & (!g2320) & (g2426) & (g2211) & (!g2076) & (g2077)) + ((!g2514) & (!g2320) & (g2426) & (g2211) & (g2076) & (g2077)) + ((!g2514) & (g2320) & (!g2426) & (!g2211) & (g2076) & (!g2077)) + ((!g2514) & (g2320) & (!g2426) & (g2211) & (g2076) & (!g2077)) + ((!g2514) & (g2320) & (!g2426) & (g2211) & (g2076) & (g2077)) + ((!g2514) & (g2320) & (g2426) & (!g2211) & (!g2076) & (g2077)) + ((!g2514) & (g2320) & (g2426) & (!g2211) & (g2076) & (!g2077)) + ((!g2514) & (g2320) & (g2426) & (g2211) & (!g2076) & (g2077)) + ((!g2514) & (g2320) & (g2426) & (g2211) & (g2076) & (!g2077)) + ((!g2514) & (g2320) & (g2426) & (g2211) & (g2076) & (g2077)) + ((g2514) & (!g2320) & (!g2426) & (!g2211) & (!g2076) & (!g2077)) + ((g2514) & (!g2320) & (!g2426) & (g2211) & (!g2076) & (!g2077)) + ((g2514) & (!g2320) & (!g2426) & (g2211) & (g2076) & (g2077)) + ((g2514) & (!g2320) & (g2426) & (!g2211) & (!g2076) & (!g2077)) + ((g2514) & (!g2320) & (g2426) & (!g2211) & (!g2076) & (g2077)) + ((g2514) & (!g2320) & (g2426) & (g2211) & (!g2076) & (!g2077)) + ((g2514) & (!g2320) & (g2426) & (g2211) & (!g2076) & (g2077)) + ((g2514) & (!g2320) & (g2426) & (g2211) & (g2076) & (g2077)) + ((g2514) & (g2320) & (!g2426) & (!g2211) & (!g2076) & (!g2077)) + ((g2514) & (g2320) & (!g2426) & (!g2211) & (g2076) & (!g2077)) + ((g2514) & (g2320) & (!g2426) & (g2211) & (!g2076) & (!g2077)) + ((g2514) & (g2320) & (!g2426) & (g2211) & (g2076) & (!g2077)) + ((g2514) & (g2320) & (!g2426) & (g2211) & (g2076) & (g2077)) + ((g2514) & (g2320) & (g2426) & (!g2211) & (!g2076) & (!g2077)) + ((g2514) & (g2320) & (g2426) & (!g2211) & (!g2076) & (g2077)) + ((g2514) & (g2320) & (g2426) & (!g2211) & (g2076) & (!g2077)) + ((g2514) & (g2320) & (g2426) & (g2211) & (!g2076) & (!g2077)) + ((g2514) & (g2320) & (g2426) & (g2211) & (!g2076) & (g2077)) + ((g2514) & (g2320) & (g2426) & (g2211) & (g2076) & (!g2077)) + ((g2514) & (g2320) & (g2426) & (g2211) & (g2076) & (g2077)));
	assign g2516 = (((!sk[92]) & (!g2076) & (!g2077) & (!g2192) & (g2218)) + ((!sk[92]) & (!g2076) & (!g2077) & (g2192) & (!g2218)) + ((!sk[92]) & (!g2076) & (!g2077) & (g2192) & (g2218)) + ((!sk[92]) & (!g2076) & (g2077) & (!g2192) & (!g2218)) + ((!sk[92]) & (!g2076) & (g2077) & (!g2192) & (g2218)) + ((!sk[92]) & (!g2076) & (g2077) & (g2192) & (!g2218)) + ((!sk[92]) & (!g2076) & (g2077) & (g2192) & (g2218)) + ((!sk[92]) & (g2076) & (!g2077) & (!g2192) & (g2218)) + ((!sk[92]) & (g2076) & (!g2077) & (g2192) & (!g2218)) + ((!sk[92]) & (g2076) & (!g2077) & (g2192) & (g2218)) + ((!sk[92]) & (g2076) & (g2077) & (!g2192) & (!g2218)) + ((!sk[92]) & (g2076) & (g2077) & (!g2192) & (g2218)) + ((!sk[92]) & (g2076) & (g2077) & (g2192) & (!g2218)) + ((!sk[92]) & (g2076) & (g2077) & (g2192) & (g2218)) + ((sk[92]) & (!g2076) & (!g2077) & (!g2192) & (g2218)) + ((sk[92]) & (!g2076) & (!g2077) & (g2192) & (g2218)) + ((sk[92]) & (!g2076) & (g2077) & (g2192) & (!g2218)) + ((sk[92]) & (!g2076) & (g2077) & (g2192) & (g2218)) + ((sk[92]) & (g2076) & (!g2077) & (g2192) & (!g2218)) + ((sk[92]) & (g2076) & (!g2077) & (g2192) & (g2218)) + ((sk[92]) & (g2076) & (g2077) & (g2192) & (!g2218)) + ((sk[92]) & (g2076) & (g2077) & (g2192) & (g2218)));
	assign g2517 = (((!g2223) & (!g2217) & (!g2215) & (g2216) & (g2076) & (g2077)) + ((!g2223) & (!g2217) & (g2215) & (!g2216) & (!g2076) & (g2077)) + ((!g2223) & (!g2217) & (g2215) & (g2216) & (!g2076) & (g2077)) + ((!g2223) & (!g2217) & (g2215) & (g2216) & (g2076) & (g2077)) + ((!g2223) & (g2217) & (!g2215) & (!g2216) & (g2076) & (!g2077)) + ((!g2223) & (g2217) & (!g2215) & (g2216) & (g2076) & (!g2077)) + ((!g2223) & (g2217) & (!g2215) & (g2216) & (g2076) & (g2077)) + ((!g2223) & (g2217) & (g2215) & (!g2216) & (!g2076) & (g2077)) + ((!g2223) & (g2217) & (g2215) & (!g2216) & (g2076) & (!g2077)) + ((!g2223) & (g2217) & (g2215) & (g2216) & (!g2076) & (g2077)) + ((!g2223) & (g2217) & (g2215) & (g2216) & (g2076) & (!g2077)) + ((!g2223) & (g2217) & (g2215) & (g2216) & (g2076) & (g2077)) + ((g2223) & (!g2217) & (!g2215) & (!g2216) & (!g2076) & (!g2077)) + ((g2223) & (!g2217) & (!g2215) & (g2216) & (!g2076) & (!g2077)) + ((g2223) & (!g2217) & (!g2215) & (g2216) & (g2076) & (g2077)) + ((g2223) & (!g2217) & (g2215) & (!g2216) & (!g2076) & (!g2077)) + ((g2223) & (!g2217) & (g2215) & (!g2216) & (!g2076) & (g2077)) + ((g2223) & (!g2217) & (g2215) & (g2216) & (!g2076) & (!g2077)) + ((g2223) & (!g2217) & (g2215) & (g2216) & (!g2076) & (g2077)) + ((g2223) & (!g2217) & (g2215) & (g2216) & (g2076) & (g2077)) + ((g2223) & (g2217) & (!g2215) & (!g2216) & (!g2076) & (!g2077)) + ((g2223) & (g2217) & (!g2215) & (!g2216) & (g2076) & (!g2077)) + ((g2223) & (g2217) & (!g2215) & (g2216) & (!g2076) & (!g2077)) + ((g2223) & (g2217) & (!g2215) & (g2216) & (g2076) & (!g2077)) + ((g2223) & (g2217) & (!g2215) & (g2216) & (g2076) & (g2077)) + ((g2223) & (g2217) & (g2215) & (!g2216) & (!g2076) & (!g2077)) + ((g2223) & (g2217) & (g2215) & (!g2216) & (!g2076) & (g2077)) + ((g2223) & (g2217) & (g2215) & (!g2216) & (g2076) & (!g2077)) + ((g2223) & (g2217) & (g2215) & (g2216) & (!g2076) & (!g2077)) + ((g2223) & (g2217) & (g2215) & (g2216) & (!g2076) & (g2077)) + ((g2223) & (g2217) & (g2215) & (g2216) & (g2076) & (!g2077)) + ((g2223) & (g2217) & (g2215) & (g2216) & (g2076) & (g2077)));
	assign g2518 = (((!g2073) & (!g2080) & (!g2125) & (g2515) & (!g2516) & (!g2517)) + ((!g2073) & (!g2080) & (!g2125) & (g2515) & (!g2516) & (g2517)) + ((!g2073) & (!g2080) & (!g2125) & (g2515) & (g2516) & (!g2517)) + ((!g2073) & (!g2080) & (!g2125) & (g2515) & (g2516) & (g2517)) + ((!g2073) & (!g2080) & (g2125) & (!g2515) & (!g2516) & (g2517)) + ((!g2073) & (!g2080) & (g2125) & (!g2515) & (g2516) & (g2517)) + ((!g2073) & (!g2080) & (g2125) & (g2515) & (!g2516) & (g2517)) + ((!g2073) & (!g2080) & (g2125) & (g2515) & (g2516) & (g2517)) + ((!g2073) & (g2080) & (!g2125) & (g2515) & (!g2516) & (!g2517)) + ((!g2073) & (g2080) & (!g2125) & (g2515) & (!g2516) & (g2517)) + ((!g2073) & (g2080) & (!g2125) & (g2515) & (g2516) & (!g2517)) + ((!g2073) & (g2080) & (!g2125) & (g2515) & (g2516) & (g2517)) + ((!g2073) & (g2080) & (g2125) & (!g2515) & (!g2516) & (g2517)) + ((!g2073) & (g2080) & (g2125) & (!g2515) & (g2516) & (g2517)) + ((!g2073) & (g2080) & (g2125) & (g2515) & (!g2516) & (g2517)) + ((!g2073) & (g2080) & (g2125) & (g2515) & (g2516) & (g2517)) + ((g2073) & (!g2080) & (g2125) & (!g2515) & (g2516) & (!g2517)) + ((g2073) & (!g2080) & (g2125) & (!g2515) & (g2516) & (g2517)) + ((g2073) & (!g2080) & (g2125) & (g2515) & (g2516) & (!g2517)) + ((g2073) & (!g2080) & (g2125) & (g2515) & (g2516) & (g2517)) + ((g2073) & (g2080) & (!g2125) & (g2515) & (!g2516) & (!g2517)) + ((g2073) & (g2080) & (!g2125) & (g2515) & (!g2516) & (g2517)) + ((g2073) & (g2080) & (!g2125) & (g2515) & (g2516) & (!g2517)) + ((g2073) & (g2080) & (!g2125) & (g2515) & (g2516) & (g2517)) + ((g2073) & (g2080) & (g2125) & (!g2515) & (g2516) & (!g2517)) + ((g2073) & (g2080) & (g2125) & (!g2515) & (g2516) & (g2517)) + ((g2073) & (g2080) & (g2125) & (g2515) & (g2516) & (!g2517)) + ((g2073) & (g2080) & (g2125) & (g2515) & (g2516) & (g2517)));
	assign g2519 = (((!g2507) & (!g2120) & (!g2124) & (!g2264) & (!g3575) & (!g2518)) + ((!g2507) & (!g2120) & (!g2124) & (!g2264) & (g3575) & (!g2518)) + ((!g2507) & (!g2120) & (!g2124) & (g2264) & (!g3575) & (!g2518)) + ((!g2507) & (!g2120) & (!g2124) & (g2264) & (!g3575) & (g2518)) + ((!g2507) & (!g2120) & (g2124) & (!g2264) & (!g3575) & (!g2518)) + ((!g2507) & (!g2120) & (g2124) & (!g2264) & (!g3575) & (g2518)) + ((!g2507) & (!g2120) & (g2124) & (!g2264) & (g3575) & (!g2518)) + ((!g2507) & (!g2120) & (g2124) & (!g2264) & (g3575) & (g2518)) + ((!g2507) & (!g2120) & (g2124) & (g2264) & (!g3575) & (!g2518)) + ((!g2507) & (!g2120) & (g2124) & (g2264) & (!g3575) & (g2518)) + ((!g2507) & (!g2120) & (g2124) & (g2264) & (g3575) & (!g2518)) + ((!g2507) & (!g2120) & (g2124) & (g2264) & (g3575) & (g2518)) + ((!g2507) & (g2120) & (!g2124) & (!g2264) & (!g3575) & (!g2518)) + ((!g2507) & (g2120) & (!g2124) & (!g2264) & (g3575) & (!g2518)) + ((!g2507) & (g2120) & (!g2124) & (g2264) & (!g3575) & (!g2518)) + ((!g2507) & (g2120) & (!g2124) & (g2264) & (!g3575) & (g2518)) + ((g2507) & (!g2120) & (!g2124) & (!g2264) & (!g3575) & (!g2518)) + ((g2507) & (!g2120) & (!g2124) & (!g2264) & (g3575) & (!g2518)) + ((g2507) & (!g2120) & (!g2124) & (g2264) & (!g3575) & (!g2518)) + ((g2507) & (!g2120) & (!g2124) & (g2264) & (!g3575) & (g2518)) + ((g2507) & (g2120) & (!g2124) & (!g2264) & (!g3575) & (!g2518)) + ((g2507) & (g2120) & (!g2124) & (!g2264) & (g3575) & (!g2518)) + ((g2507) & (g2120) & (!g2124) & (g2264) & (!g3575) & (!g2518)) + ((g2507) & (g2120) & (!g2124) & (g2264) & (!g3575) & (g2518)) + ((g2507) & (g2120) & (g2124) & (g2264) & (!g3575) & (!g2518)) + ((g2507) & (g2120) & (g2124) & (g2264) & (!g3575) & (g2518)) + ((g2507) & (g2120) & (g2124) & (g2264) & (g3575) & (!g2518)) + ((g2507) & (g2120) & (g2124) & (g2264) & (g3575) & (g2518)));
	assign g2520 = (((!g75) & (!g2120) & (!g2280) & (!g2505) & (!g2506) & (!g2519)) + ((!g75) & (!g2120) & (!g2280) & (!g2505) & (g2506) & (!g2519)) + ((!g75) & (!g2120) & (!g2280) & (g2505) & (!g2506) & (!g2519)) + ((!g75) & (!g2120) & (!g2280) & (g2505) & (g2506) & (!g2519)) + ((!g75) & (g2120) & (!g2280) & (!g2505) & (!g2506) & (!g2519)) + ((!g75) & (g2120) & (!g2280) & (!g2505) & (g2506) & (!g2519)) + ((!g75) & (g2120) & (!g2280) & (g2505) & (!g2506) & (!g2519)) + ((!g75) & (g2120) & (!g2280) & (g2505) & (g2506) & (!g2519)) + ((!g75) & (g2120) & (g2280) & (!g2505) & (!g2506) & (!g2519)) + ((!g75) & (g2120) & (g2280) & (!g2505) & (!g2506) & (g2519)) + ((!g75) & (g2120) & (g2280) & (!g2505) & (g2506) & (!g2519)) + ((!g75) & (g2120) & (g2280) & (!g2505) & (g2506) & (g2519)) + ((!g75) & (g2120) & (g2280) & (g2505) & (!g2506) & (!g2519)) + ((!g75) & (g2120) & (g2280) & (g2505) & (!g2506) & (g2519)) + ((!g75) & (g2120) & (g2280) & (g2505) & (g2506) & (!g2519)) + ((!g75) & (g2120) & (g2280) & (g2505) & (g2506) & (g2519)) + ((g75) & (!g2120) & (!g2280) & (!g2505) & (g2506) & (!g2519)) + ((g75) & (!g2120) & (!g2280) & (!g2505) & (g2506) & (g2519)) + ((g75) & (!g2120) & (!g2280) & (g2505) & (!g2506) & (!g2519)) + ((g75) & (!g2120) & (!g2280) & (g2505) & (!g2506) & (g2519)) + ((g75) & (!g2120) & (!g2280) & (g2505) & (g2506) & (!g2519)) + ((g75) & (!g2120) & (!g2280) & (g2505) & (g2506) & (g2519)) + ((g75) & (!g2120) & (g2280) & (!g2505) & (g2506) & (!g2519)) + ((g75) & (!g2120) & (g2280) & (!g2505) & (g2506) & (g2519)) + ((g75) & (!g2120) & (g2280) & (g2505) & (!g2506) & (!g2519)) + ((g75) & (!g2120) & (g2280) & (g2505) & (!g2506) & (g2519)) + ((g75) & (!g2120) & (g2280) & (g2505) & (g2506) & (!g2519)) + ((g75) & (!g2120) & (g2280) & (g2505) & (g2506) & (g2519)) + ((g75) & (g2120) & (!g2280) & (!g2505) & (g2506) & (!g2519)) + ((g75) & (g2120) & (!g2280) & (!g2505) & (g2506) & (g2519)) + ((g75) & (g2120) & (!g2280) & (g2505) & (!g2506) & (!g2519)) + ((g75) & (g2120) & (!g2280) & (g2505) & (!g2506) & (g2519)) + ((g75) & (g2120) & (!g2280) & (g2505) & (g2506) & (!g2519)) + ((g75) & (g2120) & (!g2280) & (g2505) & (g2506) & (g2519)) + ((g75) & (g2120) & (g2280) & (!g2505) & (g2506) & (!g2519)) + ((g75) & (g2120) & (g2280) & (!g2505) & (g2506) & (g2519)) + ((g75) & (g2120) & (g2280) & (g2505) & (!g2506) & (!g2519)) + ((g75) & (g2120) & (g2280) & (g2505) & (!g2506) & (g2519)) + ((g75) & (g2120) & (g2280) & (g2505) & (g2506) & (!g2519)) + ((g75) & (g2120) & (g2280) & (g2505) & (g2506) & (g2519)));
	assign g2521 = (((!sk[97]) & (!g771) & (!g2496) & (g818)) + ((!sk[97]) & (!g771) & (g2496) & (!g818)) + ((!sk[97]) & (!g771) & (g2496) & (g818)) + ((!sk[97]) & (g771) & (!g2496) & (g818)) + ((!sk[97]) & (g771) & (g2496) & (!g818)) + ((!sk[97]) & (g771) & (g2496) & (g818)) + ((sk[97]) & (!g771) & (!g2496) & (g818)) + ((sk[97]) & (!g771) & (g2496) & (g818)) + ((sk[97]) & (g771) & (!g2496) & (g818)) + ((sk[97]) & (g771) & (g2496) & (!g818)));
	assign g2522 = (((!g1785) & (!sk[98]) & (!g2033) & (g2034)) + ((!g1785) & (!sk[98]) & (g2033) & (!g2034)) + ((!g1785) & (!sk[98]) & (g2033) & (g2034)) + ((g1785) & (!sk[98]) & (!g2033) & (g2034)) + ((g1785) & (!sk[98]) & (g2033) & (!g2034)) + ((g1785) & (!sk[98]) & (g2033) & (g2034)) + ((g1785) & (sk[98]) & (!g2033) & (g2034)));
	assign g5038 = (((!g2921) & (!sk[99]) & (!g3226) & (g2523)) + ((!g2921) & (!sk[99]) & (g3226) & (!g2523)) + ((!g2921) & (!sk[99]) & (g3226) & (g2523)) + ((!g2921) & (sk[99]) & (!g3226) & (g2523)) + ((!g2921) & (sk[99]) & (g3226) & (g2523)) + ((g2921) & (!sk[99]) & (!g3226) & (g2523)) + ((g2921) & (!sk[99]) & (g3226) & (!g2523)) + ((g2921) & (!sk[99]) & (g3226) & (g2523)) + ((g2921) & (sk[99]) & (g3226) & (!g2523)) + ((g2921) & (sk[99]) & (g3226) & (g2523)));
	assign g2524 = (((!g677) & (!g726) & (!g771) & (!g2502) & (sk[100]) & (g818)) + ((!g677) & (!g726) & (!g771) & (g2502) & (!sk[100]) & (!g818)) + ((!g677) & (!g726) & (!g771) & (g2502) & (!sk[100]) & (g818)) + ((!g677) & (!g726) & (!g771) & (g2502) & (sk[100]) & (g818)) + ((!g677) & (!g726) & (g771) & (!g2502) & (!sk[100]) & (!g818)) + ((!g677) & (!g726) & (g771) & (!g2502) & (!sk[100]) & (g818)) + ((!g677) & (!g726) & (g771) & (!g2502) & (sk[100]) & (!g818)) + ((!g677) & (!g726) & (g771) & (g2502) & (!sk[100]) & (!g818)) + ((!g677) & (!g726) & (g771) & (g2502) & (!sk[100]) & (g818)) + ((!g677) & (!g726) & (g771) & (g2502) & (sk[100]) & (g818)) + ((!g677) & (g726) & (!g771) & (!g2502) & (!sk[100]) & (!g818)) + ((!g677) & (g726) & (!g771) & (!g2502) & (!sk[100]) & (g818)) + ((!g677) & (g726) & (!g771) & (!g2502) & (sk[100]) & (!g818)) + ((!g677) & (g726) & (!g771) & (g2502) & (!sk[100]) & (!g818)) + ((!g677) & (g726) & (!g771) & (g2502) & (!sk[100]) & (g818)) + ((!g677) & (g726) & (!g771) & (g2502) & (sk[100]) & (!g818)) + ((!g677) & (g726) & (g771) & (!g2502) & (!sk[100]) & (!g818)) + ((!g677) & (g726) & (g771) & (!g2502) & (!sk[100]) & (g818)) + ((!g677) & (g726) & (g771) & (!g2502) & (sk[100]) & (g818)) + ((!g677) & (g726) & (g771) & (g2502) & (!sk[100]) & (!g818)) + ((!g677) & (g726) & (g771) & (g2502) & (!sk[100]) & (g818)) + ((!g677) & (g726) & (g771) & (g2502) & (sk[100]) & (!g818)) + ((g677) & (!g726) & (!g771) & (!g2502) & (sk[100]) & (!g818)) + ((g677) & (!g726) & (!g771) & (g2502) & (!sk[100]) & (!g818)) + ((g677) & (!g726) & (!g771) & (g2502) & (!sk[100]) & (g818)) + ((g677) & (!g726) & (!g771) & (g2502) & (sk[100]) & (g818)) + ((g677) & (!g726) & (g771) & (!g2502) & (!sk[100]) & (!g818)) + ((g677) & (!g726) & (g771) & (!g2502) & (!sk[100]) & (g818)) + ((g677) & (!g726) & (g771) & (!g2502) & (sk[100]) & (!g818)) + ((g677) & (!g726) & (g771) & (g2502) & (!sk[100]) & (!g818)) + ((g677) & (!g726) & (g771) & (g2502) & (!sk[100]) & (g818)) + ((g677) & (!g726) & (g771) & (g2502) & (sk[100]) & (!g818)) + ((g677) & (g726) & (!g771) & (!g2502) & (!sk[100]) & (!g818)) + ((g677) & (g726) & (!g771) & (!g2502) & (!sk[100]) & (g818)) + ((g677) & (g726) & (!g771) & (!g2502) & (sk[100]) & (g818)) + ((g677) & (g726) & (!g771) & (g2502) & (!sk[100]) & (!g818)) + ((g677) & (g726) & (!g771) & (g2502) & (!sk[100]) & (g818)) + ((g677) & (g726) & (!g771) & (g2502) & (sk[100]) & (!g818)) + ((g677) & (g726) & (g771) & (!g2502) & (!sk[100]) & (!g818)) + ((g677) & (g726) & (g771) & (!g2502) & (!sk[100]) & (g818)) + ((g677) & (g726) & (g771) & (!g2502) & (sk[100]) & (g818)) + ((g677) & (g726) & (g771) & (g2502) & (!sk[100]) & (!g818)) + ((g677) & (g726) & (g771) & (g2502) & (!sk[100]) & (g818)) + ((g677) & (g726) & (g771) & (g2502) & (sk[100]) & (g818)));
	assign g2525 = (((!g2033) & (!sk[101]) & (!g2034) & (!g2523) & (g2524)) + ((!g2033) & (!sk[101]) & (!g2034) & (g2523) & (!g2524)) + ((!g2033) & (!sk[101]) & (!g2034) & (g2523) & (g2524)) + ((!g2033) & (!sk[101]) & (g2034) & (!g2523) & (!g2524)) + ((!g2033) & (!sk[101]) & (g2034) & (!g2523) & (g2524)) + ((!g2033) & (!sk[101]) & (g2034) & (g2523) & (!g2524)) + ((!g2033) & (!sk[101]) & (g2034) & (g2523) & (g2524)) + ((!g2033) & (sk[101]) & (!g2034) & (g2523) & (!g2524)) + ((!g2033) & (sk[101]) & (!g2034) & (g2523) & (g2524)) + ((g2033) & (!sk[101]) & (!g2034) & (!g2523) & (g2524)) + ((g2033) & (!sk[101]) & (!g2034) & (g2523) & (!g2524)) + ((g2033) & (!sk[101]) & (!g2034) & (g2523) & (g2524)) + ((g2033) & (!sk[101]) & (g2034) & (!g2523) & (!g2524)) + ((g2033) & (!sk[101]) & (g2034) & (!g2523) & (g2524)) + ((g2033) & (!sk[101]) & (g2034) & (g2523) & (!g2524)) + ((g2033) & (!sk[101]) & (g2034) & (g2523) & (g2524)) + ((g2033) & (sk[101]) & (!g2034) & (!g2523) & (g2524)) + ((g2033) & (sk[101]) & (!g2034) & (g2523) & (g2524)));
	assign g2526 = (((g2329) & (!g2029) & (g2408) & (!g2521) & (!g2522) & (g2525)) + ((g2329) & (!g2029) & (g2408) & (!g2521) & (g2522) & (!g2525)) + ((g2329) & (!g2029) & (g2408) & (!g2521) & (g2522) & (g2525)) + ((g2329) & (!g2029) & (g2408) & (g2521) & (!g2522) & (g2525)) + ((g2329) & (!g2029) & (g2408) & (g2521) & (g2522) & (!g2525)) + ((g2329) & (!g2029) & (g2408) & (g2521) & (g2522) & (g2525)) + ((g2329) & (g2029) & (g2408) & (g2521) & (!g2522) & (!g2525)) + ((g2329) & (g2029) & (g2408) & (g2521) & (!g2522) & (g2525)) + ((g2329) & (g2029) & (g2408) & (g2521) & (g2522) & (!g2525)) + ((g2329) & (g2029) & (g2408) & (g2521) & (g2522) & (g2525)));
	assign g2527 = (((!dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[103]) & (!g2128) & (g2129)) + ((!dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[103]) & (g2128) & (!g2129)) + ((!dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[103]) & (g2128) & (g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[103]) & (!g2128) & (!g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[103]) & (!g2128) & (g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[103]) & (g2128) & (!g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[103]) & (g2128) & (g2129)) + ((!dmem_dat_ix31x) & (dmem_dat_ix15x) & (sk[103]) & (!g2128) & (g2129)) + ((dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[103]) & (!g2128) & (g2129)) + ((dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[103]) & (g2128) & (!g2129)) + ((dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[103]) & (g2128) & (g2129)) + ((dmem_dat_ix31x) & (!dmem_dat_ix15x) & (sk[103]) & (!g2128) & (!g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[103]) & (!g2128) & (!g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[103]) & (!g2128) & (g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[103]) & (g2128) & (!g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[103]) & (g2128) & (g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix15x) & (sk[103]) & (!g2128) & (!g2129)) + ((dmem_dat_ix31x) & (dmem_dat_ix15x) & (sk[103]) & (!g2128) & (g2129)));
	assign g2528 = (((!g2363) & (g2131) & (!g2132) & (dmem_dat_ix15x) & (!g2338) & (!g2527)) + ((!g2363) & (g2131) & (!g2132) & (dmem_dat_ix15x) & (!g2338) & (g2527)) + ((!g2363) & (g2131) & (!g2132) & (dmem_dat_ix15x) & (g2338) & (!g2527)) + ((!g2363) & (g2131) & (!g2132) & (dmem_dat_ix15x) & (g2338) & (g2527)) + ((!g2363) & (g2131) & (g2132) & (!dmem_dat_ix15x) & (!g2338) & (g2527)) + ((!g2363) & (g2131) & (g2132) & (!dmem_dat_ix15x) & (g2338) & (g2527)) + ((!g2363) & (g2131) & (g2132) & (dmem_dat_ix15x) & (!g2338) & (g2527)) + ((!g2363) & (g2131) & (g2132) & (dmem_dat_ix15x) & (g2338) & (g2527)) + ((g2363) & (!g2131) & (!g2132) & (!dmem_dat_ix15x) & (g2338) & (!g2527)) + ((g2363) & (!g2131) & (!g2132) & (!dmem_dat_ix15x) & (g2338) & (g2527)) + ((g2363) & (!g2131) & (!g2132) & (dmem_dat_ix15x) & (g2338) & (!g2527)) + ((g2363) & (!g2131) & (!g2132) & (dmem_dat_ix15x) & (g2338) & (g2527)) + ((g2363) & (!g2131) & (g2132) & (!dmem_dat_ix15x) & (g2338) & (!g2527)) + ((g2363) & (!g2131) & (g2132) & (!dmem_dat_ix15x) & (g2338) & (g2527)) + ((g2363) & (!g2131) & (g2132) & (dmem_dat_ix15x) & (g2338) & (!g2527)) + ((g2363) & (!g2131) & (g2132) & (dmem_dat_ix15x) & (g2338) & (g2527)) + ((g2363) & (g2131) & (!g2132) & (dmem_dat_ix15x) & (!g2338) & (!g2527)) + ((g2363) & (g2131) & (!g2132) & (dmem_dat_ix15x) & (!g2338) & (g2527)) + ((g2363) & (g2131) & (!g2132) & (dmem_dat_ix15x) & (g2338) & (!g2527)) + ((g2363) & (g2131) & (!g2132) & (dmem_dat_ix15x) & (g2338) & (g2527)) + ((g2363) & (g2131) & (g2132) & (!dmem_dat_ix15x) & (!g2338) & (g2527)) + ((g2363) & (g2131) & (g2132) & (!dmem_dat_ix15x) & (g2338) & (g2527)) + ((g2363) & (g2131) & (g2132) & (dmem_dat_ix15x) & (!g2338) & (g2527)) + ((g2363) & (g2131) & (g2132) & (dmem_dat_ix15x) & (g2338) & (g2527)));
	assign g2530 = (((!g2119) & (!g2120) & (!g2482) & (!g2483) & (!g2507) & (!g3119)) + ((!g2119) & (!g2120) & (!g2482) & (!g2483) & (g2507) & (!g3119)) + ((!g2119) & (!g2120) & (!g2482) & (g2483) & (!g2507) & (!g3119)) + ((!g2119) & (!g2120) & (!g2482) & (g2483) & (g2507) & (!g3119)) + ((!g2119) & (!g2120) & (g2482) & (!g2483) & (!g2507) & (!g3119)) + ((!g2119) & (!g2120) & (g2482) & (!g2483) & (g2507) & (!g3119)) + ((!g2119) & (!g2120) & (g2482) & (g2483) & (!g2507) & (!g3119)) + ((!g2119) & (!g2120) & (g2482) & (g2483) & (g2507) & (g3119)) + ((!g2119) & (g2120) & (!g2482) & (!g2483) & (!g2507) & (!g3119)) + ((!g2119) & (g2120) & (!g2482) & (!g2483) & (g2507) & (g3119)) + ((!g2119) & (g2120) & (!g2482) & (g2483) & (!g2507) & (!g3119)) + ((!g2119) & (g2120) & (!g2482) & (g2483) & (g2507) & (g3119)) + ((!g2119) & (g2120) & (g2482) & (!g2483) & (!g2507) & (!g3119)) + ((!g2119) & (g2120) & (g2482) & (!g2483) & (g2507) & (g3119)) + ((!g2119) & (g2120) & (g2482) & (g2483) & (!g2507) & (g3119)) + ((!g2119) & (g2120) & (g2482) & (g2483) & (g2507) & (g3119)) + ((g2119) & (!g2120) & (!g2482) & (!g2483) & (!g2507) & (!g3119)) + ((g2119) & (!g2120) & (!g2482) & (!g2483) & (g2507) & (!g3119)) + ((g2119) & (!g2120) & (!g2482) & (g2483) & (!g2507) & (!g3119)) + ((g2119) & (!g2120) & (!g2482) & (g2483) & (g2507) & (g3119)) + ((g2119) & (!g2120) & (g2482) & (!g2483) & (!g2507) & (!g3119)) + ((g2119) & (!g2120) & (g2482) & (!g2483) & (g2507) & (g3119)) + ((g2119) & (!g2120) & (g2482) & (g2483) & (!g2507) & (!g3119)) + ((g2119) & (!g2120) & (g2482) & (g2483) & (g2507) & (g3119)) + ((g2119) & (g2120) & (!g2482) & (!g2483) & (!g2507) & (!g3119)) + ((g2119) & (g2120) & (!g2482) & (!g2483) & (g2507) & (g3119)) + ((g2119) & (g2120) & (!g2482) & (g2483) & (!g2507) & (g3119)) + ((g2119) & (g2120) & (!g2482) & (g2483) & (g2507) & (g3119)) + ((g2119) & (g2120) & (g2482) & (!g2483) & (!g2507) & (g3119)) + ((g2119) & (g2120) & (g2482) & (!g2483) & (g2507) & (g3119)) + ((g2119) & (g2120) & (g2482) & (g2483) & (!g2507) & (g3119)) + ((g2119) & (g2120) & (g2482) & (g2483) & (g2507) & (g3119)));
	assign g2531 = (((!g2484) & (!g2485) & (!sk[106]) & (!g2508) & (g2530)) + ((!g2484) & (!g2485) & (!sk[106]) & (g2508) & (!g2530)) + ((!g2484) & (!g2485) & (!sk[106]) & (g2508) & (g2530)) + ((!g2484) & (!g2485) & (sk[106]) & (!g2508) & (g2530)) + ((!g2484) & (!g2485) & (sk[106]) & (g2508) & (g2530)) + ((!g2484) & (g2485) & (!sk[106]) & (!g2508) & (!g2530)) + ((!g2484) & (g2485) & (!sk[106]) & (!g2508) & (g2530)) + ((!g2484) & (g2485) & (!sk[106]) & (g2508) & (!g2530)) + ((!g2484) & (g2485) & (!sk[106]) & (g2508) & (g2530)) + ((!g2484) & (g2485) & (sk[106]) & (!g2508) & (g2530)) + ((!g2484) & (g2485) & (sk[106]) & (g2508) & (g2530)) + ((g2484) & (!g2485) & (!sk[106]) & (!g2508) & (g2530)) + ((g2484) & (!g2485) & (!sk[106]) & (g2508) & (!g2530)) + ((g2484) & (!g2485) & (!sk[106]) & (g2508) & (g2530)) + ((g2484) & (!g2485) & (sk[106]) & (!g2508) & (g2530)) + ((g2484) & (!g2485) & (sk[106]) & (g2508) & (g2530)) + ((g2484) & (g2485) & (!sk[106]) & (!g2508) & (!g2530)) + ((g2484) & (g2485) & (!sk[106]) & (!g2508) & (g2530)) + ((g2484) & (g2485) & (!sk[106]) & (g2508) & (!g2530)) + ((g2484) & (g2485) & (!sk[106]) & (g2508) & (g2530)) + ((g2484) & (g2485) & (sk[106]) & (!g2508) & (g2530)) + ((g2484) & (g2485) & (sk[106]) & (g2508) & (!g2530)));
	assign g2532 = (((!g2509) & (!sk[107]) & (!g2510) & (g2511)) + ((!g2509) & (!sk[107]) & (g2510) & (!g2511)) + ((!g2509) & (!sk[107]) & (g2510) & (g2511)) + ((!g2509) & (sk[107]) & (!g2510) & (g2511)) + ((!g2509) & (sk[107]) & (g2510) & (!g2511)) + ((!g2509) & (sk[107]) & (g2510) & (g2511)) + ((g2509) & (!sk[107]) & (!g2510) & (g2511)) + ((g2509) & (!sk[107]) & (g2510) & (!g2511)) + ((g2509) & (!sk[107]) & (g2510) & (g2511)) + ((g2509) & (sk[107]) & (g2510) & (g2511)));
	assign g2533 = (((g2120) & (!sk[108]) & (!g2507)) + ((g2120) & (!sk[108]) & (g2507)) + ((g2120) & (sk[108]) & (!g2507)));
	assign g2534 = (((!sk[109]) & (g2121) & (!g2529)) + ((!sk[109]) & (g2121) & (g2529)) + ((sk[109]) & (!g2121) & (!g2529)) + ((sk[109]) & (g2121) & (g2529)));
	assign g2535 = (((!sk[110]) & (!g2532) & (!g2533) & (g2534)) + ((!sk[110]) & (!g2532) & (g2533) & (!g2534)) + ((!sk[110]) & (!g2532) & (g2533) & (g2534)) + ((!sk[110]) & (g2532) & (!g2533) & (g2534)) + ((!sk[110]) & (g2532) & (g2533) & (!g2534)) + ((!sk[110]) & (g2532) & (g2533) & (g2534)) + ((sk[110]) & (!g2532) & (!g2533) & (g2534)) + ((sk[110]) & (!g2532) & (g2533) & (!g2534)) + ((sk[110]) & (g2532) & (!g2533) & (!g2534)) + ((sk[110]) & (g2532) & (g2533) & (g2534)));
	assign g2536 = (((!g2121) & (!g2120) & (!g2119) & (g2118) & (g2071) & (g2074)) + ((!g2121) & (!g2120) & (g2119) & (!g2118) & (!g2071) & (g2074)) + ((!g2121) & (!g2120) & (g2119) & (g2118) & (!g2071) & (g2074)) + ((!g2121) & (!g2120) & (g2119) & (g2118) & (g2071) & (g2074)) + ((!g2121) & (g2120) & (!g2119) & (!g2118) & (g2071) & (!g2074)) + ((!g2121) & (g2120) & (!g2119) & (g2118) & (g2071) & (!g2074)) + ((!g2121) & (g2120) & (!g2119) & (g2118) & (g2071) & (g2074)) + ((!g2121) & (g2120) & (g2119) & (!g2118) & (!g2071) & (g2074)) + ((!g2121) & (g2120) & (g2119) & (!g2118) & (g2071) & (!g2074)) + ((!g2121) & (g2120) & (g2119) & (g2118) & (!g2071) & (g2074)) + ((!g2121) & (g2120) & (g2119) & (g2118) & (g2071) & (!g2074)) + ((!g2121) & (g2120) & (g2119) & (g2118) & (g2071) & (g2074)) + ((g2121) & (!g2120) & (!g2119) & (!g2118) & (!g2071) & (!g2074)) + ((g2121) & (!g2120) & (!g2119) & (g2118) & (!g2071) & (!g2074)) + ((g2121) & (!g2120) & (!g2119) & (g2118) & (g2071) & (g2074)) + ((g2121) & (!g2120) & (g2119) & (!g2118) & (!g2071) & (!g2074)) + ((g2121) & (!g2120) & (g2119) & (!g2118) & (!g2071) & (g2074)) + ((g2121) & (!g2120) & (g2119) & (g2118) & (!g2071) & (!g2074)) + ((g2121) & (!g2120) & (g2119) & (g2118) & (!g2071) & (g2074)) + ((g2121) & (!g2120) & (g2119) & (g2118) & (g2071) & (g2074)) + ((g2121) & (g2120) & (!g2119) & (!g2118) & (!g2071) & (!g2074)) + ((g2121) & (g2120) & (!g2119) & (!g2118) & (g2071) & (!g2074)) + ((g2121) & (g2120) & (!g2119) & (g2118) & (!g2071) & (!g2074)) + ((g2121) & (g2120) & (!g2119) & (g2118) & (g2071) & (!g2074)) + ((g2121) & (g2120) & (!g2119) & (g2118) & (g2071) & (g2074)) + ((g2121) & (g2120) & (g2119) & (!g2118) & (!g2071) & (!g2074)) + ((g2121) & (g2120) & (g2119) & (!g2118) & (!g2071) & (g2074)) + ((g2121) & (g2120) & (g2119) & (!g2118) & (g2071) & (!g2074)) + ((g2121) & (g2120) & (g2119) & (g2118) & (!g2071) & (!g2074)) + ((g2121) & (g2120) & (g2119) & (g2118) & (!g2071) & (g2074)) + ((g2121) & (g2120) & (g2119) & (g2118) & (g2071) & (!g2074)) + ((g2121) & (g2120) & (g2119) & (g2118) & (g2071) & (g2074)));
	assign g2537 = (((!g2536) & (!g2350) & (!g2449) & (g2236) & (g2076) & (g2077)) + ((!g2536) & (!g2350) & (g2449) & (!g2236) & (!g2076) & (g2077)) + ((!g2536) & (!g2350) & (g2449) & (g2236) & (!g2076) & (g2077)) + ((!g2536) & (!g2350) & (g2449) & (g2236) & (g2076) & (g2077)) + ((!g2536) & (g2350) & (!g2449) & (!g2236) & (g2076) & (!g2077)) + ((!g2536) & (g2350) & (!g2449) & (g2236) & (g2076) & (!g2077)) + ((!g2536) & (g2350) & (!g2449) & (g2236) & (g2076) & (g2077)) + ((!g2536) & (g2350) & (g2449) & (!g2236) & (!g2076) & (g2077)) + ((!g2536) & (g2350) & (g2449) & (!g2236) & (g2076) & (!g2077)) + ((!g2536) & (g2350) & (g2449) & (g2236) & (!g2076) & (g2077)) + ((!g2536) & (g2350) & (g2449) & (g2236) & (g2076) & (!g2077)) + ((!g2536) & (g2350) & (g2449) & (g2236) & (g2076) & (g2077)) + ((g2536) & (!g2350) & (!g2449) & (!g2236) & (!g2076) & (!g2077)) + ((g2536) & (!g2350) & (!g2449) & (g2236) & (!g2076) & (!g2077)) + ((g2536) & (!g2350) & (!g2449) & (g2236) & (g2076) & (g2077)) + ((g2536) & (!g2350) & (g2449) & (!g2236) & (!g2076) & (!g2077)) + ((g2536) & (!g2350) & (g2449) & (!g2236) & (!g2076) & (g2077)) + ((g2536) & (!g2350) & (g2449) & (g2236) & (!g2076) & (!g2077)) + ((g2536) & (!g2350) & (g2449) & (g2236) & (!g2076) & (g2077)) + ((g2536) & (!g2350) & (g2449) & (g2236) & (g2076) & (g2077)) + ((g2536) & (g2350) & (!g2449) & (!g2236) & (!g2076) & (!g2077)) + ((g2536) & (g2350) & (!g2449) & (!g2236) & (g2076) & (!g2077)) + ((g2536) & (g2350) & (!g2449) & (g2236) & (!g2076) & (!g2077)) + ((g2536) & (g2350) & (!g2449) & (g2236) & (g2076) & (!g2077)) + ((g2536) & (g2350) & (!g2449) & (g2236) & (g2076) & (g2077)) + ((g2536) & (g2350) & (g2449) & (!g2236) & (!g2076) & (!g2077)) + ((g2536) & (g2350) & (g2449) & (!g2236) & (!g2076) & (g2077)) + ((g2536) & (g2350) & (g2449) & (!g2236) & (g2076) & (!g2077)) + ((g2536) & (g2350) & (g2449) & (g2236) & (!g2076) & (!g2077)) + ((g2536) & (g2350) & (g2449) & (g2236) & (!g2076) & (g2077)) + ((g2536) & (g2350) & (g2449) & (g2236) & (g2076) & (!g2077)) + ((g2536) & (g2350) & (g2449) & (g2236) & (g2076) & (g2077)));
	assign g2538 = (((!g2076) & (!g2077) & (!sk[113]) & (!g2192) & (g2245)) + ((!g2076) & (!g2077) & (!sk[113]) & (g2192) & (!g2245)) + ((!g2076) & (!g2077) & (!sk[113]) & (g2192) & (g2245)) + ((!g2076) & (!g2077) & (sk[113]) & (!g2192) & (g2245)) + ((!g2076) & (!g2077) & (sk[113]) & (g2192) & (g2245)) + ((!g2076) & (g2077) & (!sk[113]) & (!g2192) & (!g2245)) + ((!g2076) & (g2077) & (!sk[113]) & (!g2192) & (g2245)) + ((!g2076) & (g2077) & (!sk[113]) & (g2192) & (!g2245)) + ((!g2076) & (g2077) & (!sk[113]) & (g2192) & (g2245)) + ((!g2076) & (g2077) & (sk[113]) & (g2192) & (!g2245)) + ((!g2076) & (g2077) & (sk[113]) & (g2192) & (g2245)) + ((g2076) & (!g2077) & (!sk[113]) & (!g2192) & (g2245)) + ((g2076) & (!g2077) & (!sk[113]) & (g2192) & (!g2245)) + ((g2076) & (!g2077) & (!sk[113]) & (g2192) & (g2245)) + ((g2076) & (!g2077) & (sk[113]) & (g2192) & (!g2245)) + ((g2076) & (!g2077) & (sk[113]) & (g2192) & (g2245)) + ((g2076) & (g2077) & (!sk[113]) & (!g2192) & (!g2245)) + ((g2076) & (g2077) & (!sk[113]) & (!g2192) & (g2245)) + ((g2076) & (g2077) & (!sk[113]) & (g2192) & (!g2245)) + ((g2076) & (g2077) & (!sk[113]) & (g2192) & (g2245)) + ((g2076) & (g2077) & (sk[113]) & (g2192) & (!g2245)) + ((g2076) & (g2077) & (sk[113]) & (g2192) & (g2245)));
	assign g2539 = (((!g2250) & (!g2244) & (!g2242) & (g2243) & (g2076) & (g2077)) + ((!g2250) & (!g2244) & (g2242) & (!g2243) & (!g2076) & (g2077)) + ((!g2250) & (!g2244) & (g2242) & (g2243) & (!g2076) & (g2077)) + ((!g2250) & (!g2244) & (g2242) & (g2243) & (g2076) & (g2077)) + ((!g2250) & (g2244) & (!g2242) & (!g2243) & (g2076) & (!g2077)) + ((!g2250) & (g2244) & (!g2242) & (g2243) & (g2076) & (!g2077)) + ((!g2250) & (g2244) & (!g2242) & (g2243) & (g2076) & (g2077)) + ((!g2250) & (g2244) & (g2242) & (!g2243) & (!g2076) & (g2077)) + ((!g2250) & (g2244) & (g2242) & (!g2243) & (g2076) & (!g2077)) + ((!g2250) & (g2244) & (g2242) & (g2243) & (!g2076) & (g2077)) + ((!g2250) & (g2244) & (g2242) & (g2243) & (g2076) & (!g2077)) + ((!g2250) & (g2244) & (g2242) & (g2243) & (g2076) & (g2077)) + ((g2250) & (!g2244) & (!g2242) & (!g2243) & (!g2076) & (!g2077)) + ((g2250) & (!g2244) & (!g2242) & (g2243) & (!g2076) & (!g2077)) + ((g2250) & (!g2244) & (!g2242) & (g2243) & (g2076) & (g2077)) + ((g2250) & (!g2244) & (g2242) & (!g2243) & (!g2076) & (!g2077)) + ((g2250) & (!g2244) & (g2242) & (!g2243) & (!g2076) & (g2077)) + ((g2250) & (!g2244) & (g2242) & (g2243) & (!g2076) & (!g2077)) + ((g2250) & (!g2244) & (g2242) & (g2243) & (!g2076) & (g2077)) + ((g2250) & (!g2244) & (g2242) & (g2243) & (g2076) & (g2077)) + ((g2250) & (g2244) & (!g2242) & (!g2243) & (!g2076) & (!g2077)) + ((g2250) & (g2244) & (!g2242) & (!g2243) & (g2076) & (!g2077)) + ((g2250) & (g2244) & (!g2242) & (g2243) & (!g2076) & (!g2077)) + ((g2250) & (g2244) & (!g2242) & (g2243) & (g2076) & (!g2077)) + ((g2250) & (g2244) & (!g2242) & (g2243) & (g2076) & (g2077)) + ((g2250) & (g2244) & (g2242) & (!g2243) & (!g2076) & (!g2077)) + ((g2250) & (g2244) & (g2242) & (!g2243) & (!g2076) & (g2077)) + ((g2250) & (g2244) & (g2242) & (!g2243) & (g2076) & (!g2077)) + ((g2250) & (g2244) & (g2242) & (g2243) & (!g2076) & (!g2077)) + ((g2250) & (g2244) & (g2242) & (g2243) & (!g2076) & (g2077)) + ((g2250) & (g2244) & (g2242) & (g2243) & (g2076) & (!g2077)) + ((g2250) & (g2244) & (g2242) & (g2243) & (g2076) & (g2077)));
	assign g2540 = (((!g2073) & (!g2080) & (!g2125) & (g2537) & (!g2538) & (!g2539)) + ((!g2073) & (!g2080) & (!g2125) & (g2537) & (!g2538) & (g2539)) + ((!g2073) & (!g2080) & (!g2125) & (g2537) & (g2538) & (!g2539)) + ((!g2073) & (!g2080) & (!g2125) & (g2537) & (g2538) & (g2539)) + ((!g2073) & (!g2080) & (g2125) & (!g2537) & (!g2538) & (g2539)) + ((!g2073) & (!g2080) & (g2125) & (!g2537) & (g2538) & (g2539)) + ((!g2073) & (!g2080) & (g2125) & (g2537) & (!g2538) & (g2539)) + ((!g2073) & (!g2080) & (g2125) & (g2537) & (g2538) & (g2539)) + ((!g2073) & (g2080) & (!g2125) & (g2537) & (!g2538) & (!g2539)) + ((!g2073) & (g2080) & (!g2125) & (g2537) & (!g2538) & (g2539)) + ((!g2073) & (g2080) & (!g2125) & (g2537) & (g2538) & (!g2539)) + ((!g2073) & (g2080) & (!g2125) & (g2537) & (g2538) & (g2539)) + ((!g2073) & (g2080) & (g2125) & (!g2537) & (!g2538) & (g2539)) + ((!g2073) & (g2080) & (g2125) & (!g2537) & (g2538) & (g2539)) + ((!g2073) & (g2080) & (g2125) & (g2537) & (!g2538) & (g2539)) + ((!g2073) & (g2080) & (g2125) & (g2537) & (g2538) & (g2539)) + ((g2073) & (!g2080) & (g2125) & (!g2537) & (g2538) & (!g2539)) + ((g2073) & (!g2080) & (g2125) & (!g2537) & (g2538) & (g2539)) + ((g2073) & (!g2080) & (g2125) & (g2537) & (g2538) & (!g2539)) + ((g2073) & (!g2080) & (g2125) & (g2537) & (g2538) & (g2539)) + ((g2073) & (g2080) & (!g2125) & (g2537) & (!g2538) & (!g2539)) + ((g2073) & (g2080) & (!g2125) & (g2537) & (!g2538) & (g2539)) + ((g2073) & (g2080) & (!g2125) & (g2537) & (g2538) & (!g2539)) + ((g2073) & (g2080) & (!g2125) & (g2537) & (g2538) & (g2539)) + ((g2073) & (g2080) & (g2125) & (!g2537) & (g2538) & (!g2539)) + ((g2073) & (g2080) & (g2125) & (!g2537) & (g2538) & (g2539)) + ((g2073) & (g2080) & (g2125) & (g2537) & (g2538) & (!g2539)) + ((g2073) & (g2080) & (g2125) & (g2537) & (g2538) & (g2539)));
	assign g2541 = (((!g2529) & (!g2121) & (!g2124) & (!g2264) & (!g3562) & (!g2540)) + ((!g2529) & (!g2121) & (!g2124) & (!g2264) & (g3562) & (!g2540)) + ((!g2529) & (!g2121) & (!g2124) & (g2264) & (!g3562) & (!g2540)) + ((!g2529) & (!g2121) & (!g2124) & (g2264) & (!g3562) & (g2540)) + ((!g2529) & (!g2121) & (g2124) & (!g2264) & (!g3562) & (!g2540)) + ((!g2529) & (!g2121) & (g2124) & (!g2264) & (!g3562) & (g2540)) + ((!g2529) & (!g2121) & (g2124) & (!g2264) & (g3562) & (!g2540)) + ((!g2529) & (!g2121) & (g2124) & (!g2264) & (g3562) & (g2540)) + ((!g2529) & (!g2121) & (g2124) & (g2264) & (!g3562) & (!g2540)) + ((!g2529) & (!g2121) & (g2124) & (g2264) & (!g3562) & (g2540)) + ((!g2529) & (!g2121) & (g2124) & (g2264) & (g3562) & (!g2540)) + ((!g2529) & (!g2121) & (g2124) & (g2264) & (g3562) & (g2540)) + ((!g2529) & (g2121) & (!g2124) & (!g2264) & (!g3562) & (!g2540)) + ((!g2529) & (g2121) & (!g2124) & (!g2264) & (g3562) & (!g2540)) + ((!g2529) & (g2121) & (!g2124) & (g2264) & (!g3562) & (!g2540)) + ((!g2529) & (g2121) & (!g2124) & (g2264) & (!g3562) & (g2540)) + ((g2529) & (!g2121) & (!g2124) & (!g2264) & (!g3562) & (!g2540)) + ((g2529) & (!g2121) & (!g2124) & (!g2264) & (g3562) & (!g2540)) + ((g2529) & (!g2121) & (!g2124) & (g2264) & (!g3562) & (!g2540)) + ((g2529) & (!g2121) & (!g2124) & (g2264) & (!g3562) & (g2540)) + ((g2529) & (g2121) & (!g2124) & (!g2264) & (!g3562) & (!g2540)) + ((g2529) & (g2121) & (!g2124) & (!g2264) & (g3562) & (!g2540)) + ((g2529) & (g2121) & (!g2124) & (g2264) & (!g3562) & (!g2540)) + ((g2529) & (g2121) & (!g2124) & (g2264) & (!g3562) & (g2540)) + ((g2529) & (g2121) & (g2124) & (g2264) & (!g3562) & (!g2540)) + ((g2529) & (g2121) & (g2124) & (g2264) & (!g3562) & (g2540)) + ((g2529) & (g2121) & (g2124) & (g2264) & (g3562) & (!g2540)) + ((g2529) & (g2121) & (g2124) & (g2264) & (g3562) & (g2540)));
	assign g2542 = (((!sk[117]) & (!g75) & (!g2121) & (!g2280) & (g2528) & (!g2541)) + ((!sk[117]) & (!g75) & (!g2121) & (!g2280) & (g2528) & (g2541)) + ((!sk[117]) & (!g75) & (!g2121) & (g2280) & (!g2528) & (!g2541)) + ((!sk[117]) & (!g75) & (!g2121) & (g2280) & (!g2528) & (g2541)) + ((!sk[117]) & (!g75) & (!g2121) & (g2280) & (g2528) & (!g2541)) + ((!sk[117]) & (!g75) & (!g2121) & (g2280) & (g2528) & (g2541)) + ((!sk[117]) & (!g75) & (g2121) & (!g2280) & (!g2528) & (!g2541)) + ((!sk[117]) & (!g75) & (g2121) & (!g2280) & (!g2528) & (g2541)) + ((!sk[117]) & (!g75) & (g2121) & (!g2280) & (g2528) & (!g2541)) + ((!sk[117]) & (!g75) & (g2121) & (!g2280) & (g2528) & (g2541)) + ((!sk[117]) & (!g75) & (g2121) & (g2280) & (!g2528) & (!g2541)) + ((!sk[117]) & (!g75) & (g2121) & (g2280) & (!g2528) & (g2541)) + ((!sk[117]) & (!g75) & (g2121) & (g2280) & (g2528) & (!g2541)) + ((!sk[117]) & (!g75) & (g2121) & (g2280) & (g2528) & (g2541)) + ((!sk[117]) & (g75) & (!g2121) & (!g2280) & (g2528) & (!g2541)) + ((!sk[117]) & (g75) & (!g2121) & (!g2280) & (g2528) & (g2541)) + ((!sk[117]) & (g75) & (!g2121) & (g2280) & (!g2528) & (!g2541)) + ((!sk[117]) & (g75) & (!g2121) & (g2280) & (!g2528) & (g2541)) + ((!sk[117]) & (g75) & (!g2121) & (g2280) & (g2528) & (!g2541)) + ((!sk[117]) & (g75) & (!g2121) & (g2280) & (g2528) & (g2541)) + ((!sk[117]) & (g75) & (g2121) & (!g2280) & (!g2528) & (!g2541)) + ((!sk[117]) & (g75) & (g2121) & (!g2280) & (!g2528) & (g2541)) + ((!sk[117]) & (g75) & (g2121) & (!g2280) & (g2528) & (!g2541)) + ((!sk[117]) & (g75) & (g2121) & (!g2280) & (g2528) & (g2541)) + ((!sk[117]) & (g75) & (g2121) & (g2280) & (!g2528) & (!g2541)) + ((!sk[117]) & (g75) & (g2121) & (g2280) & (!g2528) & (g2541)) + ((!sk[117]) & (g75) & (g2121) & (g2280) & (g2528) & (!g2541)) + ((!sk[117]) & (g75) & (g2121) & (g2280) & (g2528) & (g2541)) + ((sk[117]) & (!g75) & (!g2121) & (!g2280) & (!g2528) & (!g2541)) + ((sk[117]) & (!g75) & (!g2121) & (!g2280) & (g2528) & (!g2541)) + ((sk[117]) & (!g75) & (g2121) & (!g2280) & (!g2528) & (!g2541)) + ((sk[117]) & (!g75) & (g2121) & (!g2280) & (g2528) & (!g2541)) + ((sk[117]) & (!g75) & (g2121) & (g2280) & (!g2528) & (!g2541)) + ((sk[117]) & (!g75) & (g2121) & (g2280) & (!g2528) & (g2541)) + ((sk[117]) & (!g75) & (g2121) & (g2280) & (g2528) & (!g2541)) + ((sk[117]) & (!g75) & (g2121) & (g2280) & (g2528) & (g2541)) + ((sk[117]) & (g75) & (!g2121) & (!g2280) & (g2528) & (!g2541)) + ((sk[117]) & (g75) & (!g2121) & (!g2280) & (g2528) & (g2541)) + ((sk[117]) & (g75) & (!g2121) & (g2280) & (g2528) & (!g2541)) + ((sk[117]) & (g75) & (!g2121) & (g2280) & (g2528) & (g2541)) + ((sk[117]) & (g75) & (g2121) & (!g2280) & (g2528) & (!g2541)) + ((sk[117]) & (g75) & (g2121) & (!g2280) & (g2528) & (g2541)) + ((sk[117]) & (g75) & (g2121) & (g2280) & (g2528) & (!g2541)) + ((sk[117]) & (g75) & (g2121) & (g2280) & (g2528) & (g2541)));
	assign g2543 = (((!g771) & (!sk[118]) & (!g2496) & (!g818) & (g865)) + ((!g771) & (!sk[118]) & (!g2496) & (g818) & (!g865)) + ((!g771) & (!sk[118]) & (!g2496) & (g818) & (g865)) + ((!g771) & (!sk[118]) & (g2496) & (!g818) & (!g865)) + ((!g771) & (!sk[118]) & (g2496) & (!g818) & (g865)) + ((!g771) & (!sk[118]) & (g2496) & (g818) & (!g865)) + ((!g771) & (!sk[118]) & (g2496) & (g818) & (g865)) + ((!g771) & (sk[118]) & (!g2496) & (!g818) & (g865)) + ((!g771) & (sk[118]) & (!g2496) & (g818) & (g865)) + ((!g771) & (sk[118]) & (g2496) & (!g818) & (g865)) + ((!g771) & (sk[118]) & (g2496) & (g818) & (g865)) + ((g771) & (!sk[118]) & (!g2496) & (!g818) & (g865)) + ((g771) & (!sk[118]) & (!g2496) & (g818) & (!g865)) + ((g771) & (!sk[118]) & (!g2496) & (g818) & (g865)) + ((g771) & (!sk[118]) & (g2496) & (!g818) & (!g865)) + ((g771) & (!sk[118]) & (g2496) & (!g818) & (g865)) + ((g771) & (!sk[118]) & (g2496) & (g818) & (!g865)) + ((g771) & (!sk[118]) & (g2496) & (g818) & (g865)) + ((g771) & (sk[118]) & (!g2496) & (!g818) & (g865)) + ((g771) & (sk[118]) & (!g2496) & (g818) & (g865)) + ((g771) & (sk[118]) & (g2496) & (!g818) & (g865)) + ((g771) & (sk[118]) & (g2496) & (g818) & (!g865)));
	assign g5039 = (((!sk[119]) & (!g2921) & (!g3083) & (g2544)) + ((!sk[119]) & (!g2921) & (g3083) & (!g2544)) + ((!sk[119]) & (!g2921) & (g3083) & (g2544)) + ((!sk[119]) & (g2921) & (!g3083) & (g2544)) + ((!sk[119]) & (g2921) & (g3083) & (!g2544)) + ((!sk[119]) & (g2921) & (g3083) & (g2544)) + ((sk[119]) & (!g2921) & (!g3083) & (g2544)) + ((sk[119]) & (!g2921) & (g3083) & (g2544)) + ((sk[119]) & (g2921) & (g3083) & (!g2544)) + ((sk[119]) & (g2921) & (g3083) & (g2544)));
	assign g2545 = (((!g677) & (!g726) & (!g771) & (!g2500) & (!g2501) & (!g818)) + ((!g677) & (!g726) & (!g771) & (!g2500) & (!g2501) & (g818)) + ((!g677) & (!g726) & (!g771) & (!g2500) & (g2501) & (!g818)) + ((!g677) & (!g726) & (!g771) & (!g2500) & (g2501) & (g818)) + ((!g677) & (!g726) & (!g771) & (g2500) & (!g2501) & (!g818)) + ((!g677) & (!g726) & (!g771) & (g2500) & (!g2501) & (g818)) + ((!g677) & (!g726) & (!g771) & (g2500) & (g2501) & (!g818)) + ((!g677) & (!g726) & (!g771) & (g2500) & (g2501) & (g818)) + ((!g677) & (!g726) & (g771) & (!g2500) & (!g2501) & (!g818)) + ((!g677) & (!g726) & (g771) & (!g2500) & (!g2501) & (g818)) + ((!g677) & (!g726) & (g771) & (!g2500) & (g2501) & (!g818)) + ((!g677) & (!g726) & (g771) & (g2500) & (!g2501) & (!g818)) + ((!g677) & (!g726) & (g771) & (g2500) & (g2501) & (!g818)) + ((!g677) & (g726) & (!g771) & (!g2500) & (!g2501) & (!g818)) + ((!g677) & (g726) & (!g771) & (!g2500) & (g2501) & (!g818)) + ((!g677) & (g726) & (!g771) & (g2500) & (!g2501) & (!g818)) + ((!g677) & (g726) & (!g771) & (g2500) & (g2501) & (!g818)) + ((!g677) & (g726) & (g771) & (!g2500) & (!g2501) & (!g818)) + ((g677) & (!g726) & (!g771) & (!g2500) & (!g2501) & (!g818)) + ((g677) & (!g726) & (!g771) & (!g2500) & (!g2501) & (g818)) + ((g677) & (!g726) & (!g771) & (!g2500) & (g2501) & (!g818)) + ((g677) & (!g726) & (!g771) & (g2500) & (!g2501) & (!g818)) + ((g677) & (!g726) & (!g771) & (g2500) & (g2501) & (!g818)) + ((g677) & (!g726) & (g771) & (!g2500) & (!g2501) & (!g818)) + ((g677) & (!g726) & (g771) & (!g2500) & (g2501) & (!g818)) + ((g677) & (!g726) & (g771) & (g2500) & (!g2501) & (!g818)) + ((g677) & (!g726) & (g771) & (g2500) & (g2501) & (!g818)) + ((g677) & (g726) & (!g771) & (!g2500) & (!g2501) & (!g818)));
	assign g2546 = (((!g773) & (!sk[121]) & (!g865) & (g2545)) + ((!g773) & (!sk[121]) & (g865) & (!g2545)) + ((!g773) & (!sk[121]) & (g865) & (g2545)) + ((!g773) & (sk[121]) & (!g865) & (!g2545)) + ((!g773) & (sk[121]) & (g865) & (g2545)) + ((g773) & (!sk[121]) & (!g865) & (g2545)) + ((g773) & (!sk[121]) & (g865) & (!g2545)) + ((g773) & (!sk[121]) & (g865) & (g2545)) + ((g773) & (sk[121]) & (!g865) & (g2545)) + ((g773) & (sk[121]) & (g865) & (!g2545)));
	assign g2547 = (((!g1798) & (!g2033) & (!sk[122]) & (!g2034) & (g2544) & (!g2546)) + ((!g1798) & (!g2033) & (!sk[122]) & (!g2034) & (g2544) & (g2546)) + ((!g1798) & (!g2033) & (!sk[122]) & (g2034) & (!g2544) & (!g2546)) + ((!g1798) & (!g2033) & (!sk[122]) & (g2034) & (!g2544) & (g2546)) + ((!g1798) & (!g2033) & (!sk[122]) & (g2034) & (g2544) & (!g2546)) + ((!g1798) & (!g2033) & (!sk[122]) & (g2034) & (g2544) & (g2546)) + ((!g1798) & (!g2033) & (sk[122]) & (!g2034) & (g2544) & (!g2546)) + ((!g1798) & (!g2033) & (sk[122]) & (!g2034) & (g2544) & (g2546)) + ((!g1798) & (g2033) & (!sk[122]) & (!g2034) & (!g2544) & (!g2546)) + ((!g1798) & (g2033) & (!sk[122]) & (!g2034) & (!g2544) & (g2546)) + ((!g1798) & (g2033) & (!sk[122]) & (!g2034) & (g2544) & (!g2546)) + ((!g1798) & (g2033) & (!sk[122]) & (!g2034) & (g2544) & (g2546)) + ((!g1798) & (g2033) & (!sk[122]) & (g2034) & (!g2544) & (!g2546)) + ((!g1798) & (g2033) & (!sk[122]) & (g2034) & (!g2544) & (g2546)) + ((!g1798) & (g2033) & (!sk[122]) & (g2034) & (g2544) & (!g2546)) + ((!g1798) & (g2033) & (!sk[122]) & (g2034) & (g2544) & (g2546)) + ((!g1798) & (g2033) & (sk[122]) & (!g2034) & (!g2544) & (g2546)) + ((!g1798) & (g2033) & (sk[122]) & (!g2034) & (g2544) & (g2546)) + ((g1798) & (!g2033) & (!sk[122]) & (!g2034) & (g2544) & (!g2546)) + ((g1798) & (!g2033) & (!sk[122]) & (!g2034) & (g2544) & (g2546)) + ((g1798) & (!g2033) & (!sk[122]) & (g2034) & (!g2544) & (!g2546)) + ((g1798) & (!g2033) & (!sk[122]) & (g2034) & (!g2544) & (g2546)) + ((g1798) & (!g2033) & (!sk[122]) & (g2034) & (g2544) & (!g2546)) + ((g1798) & (!g2033) & (!sk[122]) & (g2034) & (g2544) & (g2546)) + ((g1798) & (!g2033) & (sk[122]) & (!g2034) & (g2544) & (!g2546)) + ((g1798) & (!g2033) & (sk[122]) & (!g2034) & (g2544) & (g2546)) + ((g1798) & (!g2033) & (sk[122]) & (g2034) & (!g2544) & (!g2546)) + ((g1798) & (!g2033) & (sk[122]) & (g2034) & (!g2544) & (g2546)) + ((g1798) & (!g2033) & (sk[122]) & (g2034) & (g2544) & (!g2546)) + ((g1798) & (!g2033) & (sk[122]) & (g2034) & (g2544) & (g2546)) + ((g1798) & (g2033) & (!sk[122]) & (!g2034) & (!g2544) & (!g2546)) + ((g1798) & (g2033) & (!sk[122]) & (!g2034) & (!g2544) & (g2546)) + ((g1798) & (g2033) & (!sk[122]) & (!g2034) & (g2544) & (!g2546)) + ((g1798) & (g2033) & (!sk[122]) & (!g2034) & (g2544) & (g2546)) + ((g1798) & (g2033) & (!sk[122]) & (g2034) & (!g2544) & (!g2546)) + ((g1798) & (g2033) & (!sk[122]) & (g2034) & (!g2544) & (g2546)) + ((g1798) & (g2033) & (!sk[122]) & (g2034) & (g2544) & (!g2546)) + ((g1798) & (g2033) & (!sk[122]) & (g2034) & (g2544) & (g2546)) + ((g1798) & (g2033) & (sk[122]) & (!g2034) & (!g2544) & (g2546)) + ((g1798) & (g2033) & (sk[122]) & (!g2034) & (g2544) & (g2546)));
	assign g2548 = (((!g2329) & (!g2029) & (!g2408) & (!sk[123]) & (g2543) & (!g2547)) + ((!g2329) & (!g2029) & (!g2408) & (!sk[123]) & (g2543) & (g2547)) + ((!g2329) & (!g2029) & (g2408) & (!sk[123]) & (!g2543) & (!g2547)) + ((!g2329) & (!g2029) & (g2408) & (!sk[123]) & (!g2543) & (g2547)) + ((!g2329) & (!g2029) & (g2408) & (!sk[123]) & (g2543) & (!g2547)) + ((!g2329) & (!g2029) & (g2408) & (!sk[123]) & (g2543) & (g2547)) + ((!g2329) & (g2029) & (!g2408) & (!sk[123]) & (!g2543) & (!g2547)) + ((!g2329) & (g2029) & (!g2408) & (!sk[123]) & (!g2543) & (g2547)) + ((!g2329) & (g2029) & (!g2408) & (!sk[123]) & (g2543) & (!g2547)) + ((!g2329) & (g2029) & (!g2408) & (!sk[123]) & (g2543) & (g2547)) + ((!g2329) & (g2029) & (g2408) & (!sk[123]) & (!g2543) & (!g2547)) + ((!g2329) & (g2029) & (g2408) & (!sk[123]) & (!g2543) & (g2547)) + ((!g2329) & (g2029) & (g2408) & (!sk[123]) & (g2543) & (!g2547)) + ((!g2329) & (g2029) & (g2408) & (!sk[123]) & (g2543) & (g2547)) + ((g2329) & (!g2029) & (!g2408) & (!sk[123]) & (g2543) & (!g2547)) + ((g2329) & (!g2029) & (!g2408) & (!sk[123]) & (g2543) & (g2547)) + ((g2329) & (!g2029) & (g2408) & (!sk[123]) & (!g2543) & (!g2547)) + ((g2329) & (!g2029) & (g2408) & (!sk[123]) & (!g2543) & (g2547)) + ((g2329) & (!g2029) & (g2408) & (!sk[123]) & (g2543) & (!g2547)) + ((g2329) & (!g2029) & (g2408) & (!sk[123]) & (g2543) & (g2547)) + ((g2329) & (!g2029) & (g2408) & (sk[123]) & (!g2543) & (g2547)) + ((g2329) & (!g2029) & (g2408) & (sk[123]) & (g2543) & (g2547)) + ((g2329) & (g2029) & (!g2408) & (!sk[123]) & (!g2543) & (!g2547)) + ((g2329) & (g2029) & (!g2408) & (!sk[123]) & (!g2543) & (g2547)) + ((g2329) & (g2029) & (!g2408) & (!sk[123]) & (g2543) & (!g2547)) + ((g2329) & (g2029) & (!g2408) & (!sk[123]) & (g2543) & (g2547)) + ((g2329) & (g2029) & (g2408) & (!sk[123]) & (!g2543) & (!g2547)) + ((g2329) & (g2029) & (g2408) & (!sk[123]) & (!g2543) & (g2547)) + ((g2329) & (g2029) & (g2408) & (!sk[123]) & (g2543) & (!g2547)) + ((g2329) & (g2029) & (g2408) & (!sk[123]) & (g2543) & (g2547)) + ((g2329) & (g2029) & (g2408) & (sk[123]) & (g2543) & (!g2547)) + ((g2329) & (g2029) & (g2408) & (sk[123]) & (g2543) & (g2547)));
	assign g2549 = (((g78) & (g79) & (g80) & (!g81) & (!g82) & (!g83)));
	assign g2550 = (((!g2363) & (g2131) & (g2549) & (g2132) & (!g2338) & (g2527)) + ((!g2363) & (g2131) & (g2549) & (g2132) & (g2338) & (g2527)) + ((g2363) & (!g2131) & (!g2549) & (!g2132) & (g2338) & (!g2527)) + ((g2363) & (!g2131) & (!g2549) & (!g2132) & (g2338) & (g2527)) + ((g2363) & (!g2131) & (!g2549) & (g2132) & (g2338) & (!g2527)) + ((g2363) & (!g2131) & (!g2549) & (g2132) & (g2338) & (g2527)) + ((g2363) & (!g2131) & (g2549) & (!g2132) & (g2338) & (!g2527)) + ((g2363) & (!g2131) & (g2549) & (!g2132) & (g2338) & (g2527)) + ((g2363) & (!g2131) & (g2549) & (g2132) & (g2338) & (!g2527)) + ((g2363) & (!g2131) & (g2549) & (g2132) & (g2338) & (g2527)) + ((g2363) & (g2131) & (g2549) & (g2132) & (!g2338) & (g2527)) + ((g2363) & (g2131) & (g2549) & (g2132) & (g2338) & (g2527)));
	assign g2552 = (((!g2111) & (!g2439) & (!g2441) & (!g2442) & (!g3137) & (g3138)) + ((!g2111) & (!g2439) & (!g2441) & (g2442) & (!g3137) & (g3138)) + ((!g2111) & (!g2439) & (g2441) & (!g2442) & (!g3137) & (g3138)) + ((!g2111) & (!g2439) & (g2441) & (g2442) & (!g3137) & (g3138)) + ((!g2111) & (g2439) & (!g2441) & (!g2442) & (!g3137) & (g3138)) + ((!g2111) & (g2439) & (!g2441) & (g2442) & (!g3137) & (g3138)) + ((!g2111) & (g2439) & (!g2441) & (g2442) & (g3137) & (g3138)) + ((!g2111) & (g2439) & (g2441) & (!g2442) & (!g3137) & (g3138)) + ((!g2111) & (g2439) & (g2441) & (!g2442) & (g3137) & (g3138)) + ((!g2111) & (g2439) & (g2441) & (g2442) & (!g3137) & (g3138)) + ((!g2111) & (g2439) & (g2441) & (g2442) & (g3137) & (g3138)) + ((g2111) & (!g2439) & (!g2441) & (!g2442) & (!g3137) & (g3138)) + ((g2111) & (!g2439) & (!g2441) & (g2442) & (!g3137) & (g3138)) + ((g2111) & (!g2439) & (!g2441) & (g2442) & (g3137) & (g3138)) + ((g2111) & (!g2439) & (g2441) & (!g2442) & (!g3137) & (g3138)) + ((g2111) & (!g2439) & (g2441) & (!g2442) & (g3137) & (g3138)) + ((g2111) & (!g2439) & (g2441) & (g2442) & (!g3137) & (g3138)) + ((g2111) & (!g2439) & (g2441) & (g2442) & (g3137) & (g3138)) + ((g2111) & (g2439) & (!g2441) & (!g2442) & (!g3137) & (g3138)) + ((g2111) & (g2439) & (!g2441) & (!g2442) & (g3137) & (g3138)) + ((g2111) & (g2439) & (!g2441) & (g2442) & (!g3137) & (g3138)) + ((g2111) & (g2439) & (!g2441) & (g2442) & (g3137) & (g3138)) + ((g2111) & (g2439) & (g2441) & (!g2442) & (!g3137) & (g3138)) + ((g2111) & (g2439) & (g2441) & (!g2442) & (g3137) & (g3138)) + ((g2111) & (g2439) & (g2441) & (g2442) & (!g3137) & (g3138)) + ((g2111) & (g2439) & (g2441) & (g2442) & (g3137) & (g3138)));
	assign g2553 = (((g2121) & (!sk[127]) & (!g2529)) + ((g2121) & (!sk[127]) & (g2529)) + ((g2121) & (sk[127]) & (g2529)));
	assign g2554 = (((!g2083) & (!g2551) & (!g2552) & (!sk[0]) & (g2553)) + ((!g2083) & (!g2551) & (!g2552) & (sk[0]) & (g2553)) + ((!g2083) & (!g2551) & (g2552) & (!sk[0]) & (!g2553)) + ((!g2083) & (!g2551) & (g2552) & (!sk[0]) & (g2553)) + ((!g2083) & (!g2551) & (g2552) & (sk[0]) & (!g2553)) + ((!g2083) & (!g2551) & (g2552) & (sk[0]) & (g2553)) + ((!g2083) & (g2551) & (!g2552) & (!sk[0]) & (!g2553)) + ((!g2083) & (g2551) & (!g2552) & (!sk[0]) & (g2553)) + ((!g2083) & (g2551) & (!g2552) & (sk[0]) & (!g2553)) + ((!g2083) & (g2551) & (g2552) & (!sk[0]) & (!g2553)) + ((!g2083) & (g2551) & (g2552) & (!sk[0]) & (g2553)) + ((g2083) & (!g2551) & (!g2552) & (!sk[0]) & (g2553)) + ((g2083) & (!g2551) & (!g2552) & (sk[0]) & (!g2553)) + ((g2083) & (!g2551) & (g2552) & (!sk[0]) & (!g2553)) + ((g2083) & (!g2551) & (g2552) & (!sk[0]) & (g2553)) + ((g2083) & (g2551) & (!g2552) & (!sk[0]) & (!g2553)) + ((g2083) & (g2551) & (!g2552) & (!sk[0]) & (g2553)) + ((g2083) & (g2551) & (!g2552) & (sk[0]) & (g2553)) + ((g2083) & (g2551) & (g2552) & (!sk[0]) & (!g2553)) + ((g2083) & (g2551) & (g2552) & (!sk[0]) & (g2553)) + ((g2083) & (g2551) & (g2552) & (sk[0]) & (!g2553)) + ((g2083) & (g2551) & (g2552) & (sk[0]) & (g2553)));
	assign g2555 = (((!g2484) & (!g2485) & (!g2508) & (!sk[1]) & (g2530)) + ((!g2484) & (!g2485) & (g2508) & (!sk[1]) & (!g2530)) + ((!g2484) & (!g2485) & (g2508) & (!sk[1]) & (g2530)) + ((!g2484) & (g2485) & (!g2508) & (!sk[1]) & (!g2530)) + ((!g2484) & (g2485) & (!g2508) & (!sk[1]) & (g2530)) + ((!g2484) & (g2485) & (g2508) & (!sk[1]) & (!g2530)) + ((!g2484) & (g2485) & (g2508) & (!sk[1]) & (g2530)) + ((g2484) & (!g2485) & (!g2508) & (!sk[1]) & (g2530)) + ((g2484) & (!g2485) & (g2508) & (!sk[1]) & (!g2530)) + ((g2484) & (!g2485) & (g2508) & (!sk[1]) & (g2530)) + ((g2484) & (g2485) & (!g2508) & (!sk[1]) & (!g2530)) + ((g2484) & (g2485) & (!g2508) & (!sk[1]) & (g2530)) + ((g2484) & (g2485) & (g2508) & (!sk[1]) & (!g2530)) + ((g2484) & (g2485) & (g2508) & (!sk[1]) & (g2530)) + ((g2484) & (g2485) & (g2508) & (sk[1]) & (g2530)));
	assign g2556 = (((!sk[2]) & (g2121) & (!g2529)) + ((!sk[2]) & (g2121) & (g2529)) + ((sk[2]) & (g2121) & (!g2529)));
	assign g2557 = (((!sk[3]) & (g2551) & (!g2083)) + ((!sk[3]) & (g2551) & (g2083)) + ((sk[3]) & (!g2551) & (!g2083)) + ((sk[3]) & (g2551) & (g2083)));
	assign g2558 = (((!g2532) & (!g2533) & (!sk[4]) & (!g2534) & (g2556) & (!g2557)) + ((!g2532) & (!g2533) & (!sk[4]) & (!g2534) & (g2556) & (g2557)) + ((!g2532) & (!g2533) & (!sk[4]) & (g2534) & (!g2556) & (!g2557)) + ((!g2532) & (!g2533) & (!sk[4]) & (g2534) & (!g2556) & (g2557)) + ((!g2532) & (!g2533) & (!sk[4]) & (g2534) & (g2556) & (!g2557)) + ((!g2532) & (!g2533) & (!sk[4]) & (g2534) & (g2556) & (g2557)) + ((!g2532) & (!g2533) & (sk[4]) & (!g2534) & (!g2556) & (g2557)) + ((!g2532) & (!g2533) & (sk[4]) & (!g2534) & (g2556) & (!g2557)) + ((!g2532) & (!g2533) & (sk[4]) & (g2534) & (!g2556) & (g2557)) + ((!g2532) & (!g2533) & (sk[4]) & (g2534) & (g2556) & (!g2557)) + ((!g2532) & (g2533) & (!sk[4]) & (!g2534) & (!g2556) & (!g2557)) + ((!g2532) & (g2533) & (!sk[4]) & (!g2534) & (!g2556) & (g2557)) + ((!g2532) & (g2533) & (!sk[4]) & (!g2534) & (g2556) & (!g2557)) + ((!g2532) & (g2533) & (!sk[4]) & (!g2534) & (g2556) & (g2557)) + ((!g2532) & (g2533) & (!sk[4]) & (g2534) & (!g2556) & (!g2557)) + ((!g2532) & (g2533) & (!sk[4]) & (g2534) & (!g2556) & (g2557)) + ((!g2532) & (g2533) & (!sk[4]) & (g2534) & (g2556) & (!g2557)) + ((!g2532) & (g2533) & (!sk[4]) & (g2534) & (g2556) & (g2557)) + ((!g2532) & (g2533) & (sk[4]) & (!g2534) & (!g2556) & (g2557)) + ((!g2532) & (g2533) & (sk[4]) & (!g2534) & (g2556) & (!g2557)) + ((!g2532) & (g2533) & (sk[4]) & (g2534) & (!g2556) & (!g2557)) + ((!g2532) & (g2533) & (sk[4]) & (g2534) & (g2556) & (g2557)) + ((g2532) & (!g2533) & (!sk[4]) & (!g2534) & (g2556) & (!g2557)) + ((g2532) & (!g2533) & (!sk[4]) & (!g2534) & (g2556) & (g2557)) + ((g2532) & (!g2533) & (!sk[4]) & (g2534) & (!g2556) & (!g2557)) + ((g2532) & (!g2533) & (!sk[4]) & (g2534) & (!g2556) & (g2557)) + ((g2532) & (!g2533) & (!sk[4]) & (g2534) & (g2556) & (!g2557)) + ((g2532) & (!g2533) & (!sk[4]) & (g2534) & (g2556) & (g2557)) + ((g2532) & (!g2533) & (sk[4]) & (!g2534) & (!g2556) & (g2557)) + ((g2532) & (!g2533) & (sk[4]) & (!g2534) & (g2556) & (!g2557)) + ((g2532) & (!g2533) & (sk[4]) & (g2534) & (!g2556) & (!g2557)) + ((g2532) & (!g2533) & (sk[4]) & (g2534) & (g2556) & (g2557)) + ((g2532) & (g2533) & (!sk[4]) & (!g2534) & (!g2556) & (!g2557)) + ((g2532) & (g2533) & (!sk[4]) & (!g2534) & (!g2556) & (g2557)) + ((g2532) & (g2533) & (!sk[4]) & (!g2534) & (g2556) & (!g2557)) + ((g2532) & (g2533) & (!sk[4]) & (!g2534) & (g2556) & (g2557)) + ((g2532) & (g2533) & (!sk[4]) & (g2534) & (!g2556) & (!g2557)) + ((g2532) & (g2533) & (!sk[4]) & (g2534) & (!g2556) & (g2557)) + ((g2532) & (g2533) & (!sk[4]) & (g2534) & (g2556) & (!g2557)) + ((g2532) & (g2533) & (!sk[4]) & (g2534) & (g2556) & (g2557)) + ((g2532) & (g2533) & (sk[4]) & (!g2534) & (!g2556) & (!g2557)) + ((g2532) & (g2533) & (sk[4]) & (!g2534) & (g2556) & (g2557)) + ((g2532) & (g2533) & (sk[4]) & (g2534) & (!g2556) & (!g2557)) + ((g2532) & (g2533) & (sk[4]) & (g2534) & (g2556) & (g2557)));
	assign g2559 = (((!g2083) & (!g2121) & (!g2120) & (g2119) & (g2071) & (g2074)) + ((!g2083) & (!g2121) & (g2120) & (!g2119) & (!g2071) & (g2074)) + ((!g2083) & (!g2121) & (g2120) & (g2119) & (!g2071) & (g2074)) + ((!g2083) & (!g2121) & (g2120) & (g2119) & (g2071) & (g2074)) + ((!g2083) & (g2121) & (!g2120) & (!g2119) & (g2071) & (!g2074)) + ((!g2083) & (g2121) & (!g2120) & (g2119) & (g2071) & (!g2074)) + ((!g2083) & (g2121) & (!g2120) & (g2119) & (g2071) & (g2074)) + ((!g2083) & (g2121) & (g2120) & (!g2119) & (!g2071) & (g2074)) + ((!g2083) & (g2121) & (g2120) & (!g2119) & (g2071) & (!g2074)) + ((!g2083) & (g2121) & (g2120) & (g2119) & (!g2071) & (g2074)) + ((!g2083) & (g2121) & (g2120) & (g2119) & (g2071) & (!g2074)) + ((!g2083) & (g2121) & (g2120) & (g2119) & (g2071) & (g2074)) + ((g2083) & (!g2121) & (!g2120) & (!g2119) & (!g2071) & (!g2074)) + ((g2083) & (!g2121) & (!g2120) & (g2119) & (!g2071) & (!g2074)) + ((g2083) & (!g2121) & (!g2120) & (g2119) & (g2071) & (g2074)) + ((g2083) & (!g2121) & (g2120) & (!g2119) & (!g2071) & (!g2074)) + ((g2083) & (!g2121) & (g2120) & (!g2119) & (!g2071) & (g2074)) + ((g2083) & (!g2121) & (g2120) & (g2119) & (!g2071) & (!g2074)) + ((g2083) & (!g2121) & (g2120) & (g2119) & (!g2071) & (g2074)) + ((g2083) & (!g2121) & (g2120) & (g2119) & (g2071) & (g2074)) + ((g2083) & (g2121) & (!g2120) & (!g2119) & (!g2071) & (!g2074)) + ((g2083) & (g2121) & (!g2120) & (!g2119) & (g2071) & (!g2074)) + ((g2083) & (g2121) & (!g2120) & (g2119) & (!g2071) & (!g2074)) + ((g2083) & (g2121) & (!g2120) & (g2119) & (g2071) & (!g2074)) + ((g2083) & (g2121) & (!g2120) & (g2119) & (g2071) & (g2074)) + ((g2083) & (g2121) & (g2120) & (!g2119) & (!g2071) & (!g2074)) + ((g2083) & (g2121) & (g2120) & (!g2119) & (!g2071) & (g2074)) + ((g2083) & (g2121) & (g2120) & (!g2119) & (g2071) & (!g2074)) + ((g2083) & (g2121) & (g2120) & (g2119) & (!g2071) & (!g2074)) + ((g2083) & (g2121) & (g2120) & (g2119) & (!g2071) & (g2074)) + ((g2083) & (g2121) & (g2120) & (g2119) & (g2071) & (!g2074)) + ((g2083) & (g2121) & (g2120) & (g2119) & (g2071) & (g2074)));
	assign g2560 = (((!g2559) & (!g2372) & (!g2467) & (g2272) & (g2076) & (g2077)) + ((!g2559) & (!g2372) & (g2467) & (!g2272) & (!g2076) & (g2077)) + ((!g2559) & (!g2372) & (g2467) & (g2272) & (!g2076) & (g2077)) + ((!g2559) & (!g2372) & (g2467) & (g2272) & (g2076) & (g2077)) + ((!g2559) & (g2372) & (!g2467) & (!g2272) & (g2076) & (!g2077)) + ((!g2559) & (g2372) & (!g2467) & (g2272) & (g2076) & (!g2077)) + ((!g2559) & (g2372) & (!g2467) & (g2272) & (g2076) & (g2077)) + ((!g2559) & (g2372) & (g2467) & (!g2272) & (!g2076) & (g2077)) + ((!g2559) & (g2372) & (g2467) & (!g2272) & (g2076) & (!g2077)) + ((!g2559) & (g2372) & (g2467) & (g2272) & (!g2076) & (g2077)) + ((!g2559) & (g2372) & (g2467) & (g2272) & (g2076) & (!g2077)) + ((!g2559) & (g2372) & (g2467) & (g2272) & (g2076) & (g2077)) + ((g2559) & (!g2372) & (!g2467) & (!g2272) & (!g2076) & (!g2077)) + ((g2559) & (!g2372) & (!g2467) & (g2272) & (!g2076) & (!g2077)) + ((g2559) & (!g2372) & (!g2467) & (g2272) & (g2076) & (g2077)) + ((g2559) & (!g2372) & (g2467) & (!g2272) & (!g2076) & (!g2077)) + ((g2559) & (!g2372) & (g2467) & (!g2272) & (!g2076) & (g2077)) + ((g2559) & (!g2372) & (g2467) & (g2272) & (!g2076) & (!g2077)) + ((g2559) & (!g2372) & (g2467) & (g2272) & (!g2076) & (g2077)) + ((g2559) & (!g2372) & (g2467) & (g2272) & (g2076) & (g2077)) + ((g2559) & (g2372) & (!g2467) & (!g2272) & (!g2076) & (!g2077)) + ((g2559) & (g2372) & (!g2467) & (!g2272) & (g2076) & (!g2077)) + ((g2559) & (g2372) & (!g2467) & (g2272) & (!g2076) & (!g2077)) + ((g2559) & (g2372) & (!g2467) & (g2272) & (g2076) & (!g2077)) + ((g2559) & (g2372) & (!g2467) & (g2272) & (g2076) & (g2077)) + ((g2559) & (g2372) & (g2467) & (!g2272) & (!g2076) & (!g2077)) + ((g2559) & (g2372) & (g2467) & (!g2272) & (!g2076) & (g2077)) + ((g2559) & (g2372) & (g2467) & (!g2272) & (g2076) & (!g2077)) + ((g2559) & (g2372) & (g2467) & (g2272) & (!g2076) & (!g2077)) + ((g2559) & (g2372) & (g2467) & (g2272) & (!g2076) & (g2077)) + ((g2559) & (g2372) & (g2467) & (g2272) & (g2076) & (!g2077)) + ((g2559) & (g2372) & (g2467) & (g2272) & (g2076) & (g2077)));
	assign g2561 = (((!g2560) & (!g2078) & (!g2103) & (g2191) & (g2073) & (g2125)) + ((!g2560) & (!g2078) & (g2103) & (!g2191) & (!g2073) & (g2125)) + ((!g2560) & (!g2078) & (g2103) & (g2191) & (!g2073) & (g2125)) + ((!g2560) & (!g2078) & (g2103) & (g2191) & (g2073) & (g2125)) + ((!g2560) & (g2078) & (!g2103) & (!g2191) & (g2073) & (!g2125)) + ((!g2560) & (g2078) & (!g2103) & (g2191) & (g2073) & (!g2125)) + ((!g2560) & (g2078) & (!g2103) & (g2191) & (g2073) & (g2125)) + ((!g2560) & (g2078) & (g2103) & (!g2191) & (!g2073) & (g2125)) + ((!g2560) & (g2078) & (g2103) & (!g2191) & (g2073) & (!g2125)) + ((!g2560) & (g2078) & (g2103) & (g2191) & (!g2073) & (g2125)) + ((!g2560) & (g2078) & (g2103) & (g2191) & (g2073) & (!g2125)) + ((!g2560) & (g2078) & (g2103) & (g2191) & (g2073) & (g2125)) + ((g2560) & (!g2078) & (!g2103) & (!g2191) & (!g2073) & (!g2125)) + ((g2560) & (!g2078) & (!g2103) & (g2191) & (!g2073) & (!g2125)) + ((g2560) & (!g2078) & (!g2103) & (g2191) & (g2073) & (g2125)) + ((g2560) & (!g2078) & (g2103) & (!g2191) & (!g2073) & (!g2125)) + ((g2560) & (!g2078) & (g2103) & (!g2191) & (!g2073) & (g2125)) + ((g2560) & (!g2078) & (g2103) & (g2191) & (!g2073) & (!g2125)) + ((g2560) & (!g2078) & (g2103) & (g2191) & (!g2073) & (g2125)) + ((g2560) & (!g2078) & (g2103) & (g2191) & (g2073) & (g2125)) + ((g2560) & (g2078) & (!g2103) & (!g2191) & (!g2073) & (!g2125)) + ((g2560) & (g2078) & (!g2103) & (!g2191) & (g2073) & (!g2125)) + ((g2560) & (g2078) & (!g2103) & (g2191) & (!g2073) & (!g2125)) + ((g2560) & (g2078) & (!g2103) & (g2191) & (g2073) & (!g2125)) + ((g2560) & (g2078) & (!g2103) & (g2191) & (g2073) & (g2125)) + ((g2560) & (g2078) & (g2103) & (!g2191) & (!g2073) & (!g2125)) + ((g2560) & (g2078) & (g2103) & (!g2191) & (!g2073) & (g2125)) + ((g2560) & (g2078) & (g2103) & (!g2191) & (g2073) & (!g2125)) + ((g2560) & (g2078) & (g2103) & (g2191) & (!g2073) & (!g2125)) + ((g2560) & (g2078) & (g2103) & (g2191) & (!g2073) & (g2125)) + ((g2560) & (g2078) & (g2103) & (g2191) & (g2073) & (!g2125)) + ((g2560) & (g2078) & (g2103) & (g2191) & (g2073) & (g2125)));
	assign g2562 = (((!g2083) & (!g2551) & (!g2124) & (!g2264) & (!g3550) & (g2561)) + ((!g2083) & (!g2551) & (!g2124) & (!g2264) & (g3550) & (g2561)) + ((!g2083) & (!g2551) & (!g2124) & (g2264) & (g3550) & (!g2561)) + ((!g2083) & (!g2551) & (!g2124) & (g2264) & (g3550) & (g2561)) + ((!g2083) & (g2551) & (!g2124) & (!g2264) & (!g3550) & (g2561)) + ((!g2083) & (g2551) & (!g2124) & (!g2264) & (g3550) & (g2561)) + ((!g2083) & (g2551) & (!g2124) & (g2264) & (g3550) & (!g2561)) + ((!g2083) & (g2551) & (!g2124) & (g2264) & (g3550) & (g2561)) + ((!g2083) & (g2551) & (g2124) & (!g2264) & (!g3550) & (!g2561)) + ((!g2083) & (g2551) & (g2124) & (!g2264) & (!g3550) & (g2561)) + ((!g2083) & (g2551) & (g2124) & (!g2264) & (g3550) & (!g2561)) + ((!g2083) & (g2551) & (g2124) & (!g2264) & (g3550) & (g2561)) + ((!g2083) & (g2551) & (g2124) & (g2264) & (!g3550) & (!g2561)) + ((!g2083) & (g2551) & (g2124) & (g2264) & (!g3550) & (g2561)) + ((!g2083) & (g2551) & (g2124) & (g2264) & (g3550) & (!g2561)) + ((!g2083) & (g2551) & (g2124) & (g2264) & (g3550) & (g2561)) + ((g2083) & (!g2551) & (!g2124) & (!g2264) & (!g3550) & (g2561)) + ((g2083) & (!g2551) & (!g2124) & (!g2264) & (g3550) & (g2561)) + ((g2083) & (!g2551) & (!g2124) & (g2264) & (g3550) & (!g2561)) + ((g2083) & (!g2551) & (!g2124) & (g2264) & (g3550) & (g2561)) + ((g2083) & (!g2551) & (g2124) & (!g2264) & (!g3550) & (!g2561)) + ((g2083) & (!g2551) & (g2124) & (!g2264) & (!g3550) & (g2561)) + ((g2083) & (!g2551) & (g2124) & (!g2264) & (g3550) & (!g2561)) + ((g2083) & (!g2551) & (g2124) & (!g2264) & (g3550) & (g2561)) + ((g2083) & (!g2551) & (g2124) & (g2264) & (!g3550) & (!g2561)) + ((g2083) & (!g2551) & (g2124) & (g2264) & (!g3550) & (g2561)) + ((g2083) & (!g2551) & (g2124) & (g2264) & (g3550) & (!g2561)) + ((g2083) & (!g2551) & (g2124) & (g2264) & (g3550) & (g2561)) + ((g2083) & (g2551) & (!g2124) & (!g2264) & (!g3550) & (g2561)) + ((g2083) & (g2551) & (!g2124) & (!g2264) & (g3550) & (g2561)) + ((g2083) & (g2551) & (!g2124) & (g2264) & (g3550) & (!g2561)) + ((g2083) & (g2551) & (!g2124) & (g2264) & (g3550) & (g2561)) + ((g2083) & (g2551) & (g2124) & (!g2264) & (!g3550) & (!g2561)) + ((g2083) & (g2551) & (g2124) & (!g2264) & (!g3550) & (g2561)) + ((g2083) & (g2551) & (g2124) & (!g2264) & (g3550) & (!g2561)) + ((g2083) & (g2551) & (g2124) & (!g2264) & (g3550) & (g2561)));
	assign g2563 = (((!g771) & (!sk[9]) & (!g2496) & (!g818) & (g865)) + ((!g771) & (!sk[9]) & (!g2496) & (g818) & (!g865)) + ((!g771) & (!sk[9]) & (!g2496) & (g818) & (g865)) + ((!g771) & (!sk[9]) & (g2496) & (!g818) & (!g865)) + ((!g771) & (!sk[9]) & (g2496) & (!g818) & (g865)) + ((!g771) & (!sk[9]) & (g2496) & (g818) & (!g865)) + ((!g771) & (!sk[9]) & (g2496) & (g818) & (g865)) + ((g771) & (!sk[9]) & (!g2496) & (!g818) & (g865)) + ((g771) & (!sk[9]) & (!g2496) & (g818) & (!g865)) + ((g771) & (!sk[9]) & (!g2496) & (g818) & (g865)) + ((g771) & (!sk[9]) & (g2496) & (!g818) & (!g865)) + ((g771) & (!sk[9]) & (g2496) & (!g818) & (g865)) + ((g771) & (!sk[9]) & (g2496) & (g818) & (!g865)) + ((g771) & (!sk[9]) & (g2496) & (g818) & (g865)) + ((g771) & (sk[9]) & (g2496) & (g818) & (g865)));
	assign g2564 = (((!sk[10]) & (g912) & (!g2563)) + ((!sk[10]) & (g912) & (g2563)) + ((sk[10]) & (!g912) & (g2563)) + ((sk[10]) & (g912) & (!g2563)));
	assign g2565 = (((!sk[11]) & (!g1810) & (!g2033) & (g2034)) + ((!sk[11]) & (!g1810) & (g2033) & (!g2034)) + ((!sk[11]) & (!g1810) & (g2033) & (g2034)) + ((!sk[11]) & (g1810) & (!g2033) & (g2034)) + ((!sk[11]) & (g1810) & (g2033) & (!g2034)) + ((!sk[11]) & (g1810) & (g2033) & (g2034)) + ((sk[11]) & (g1810) & (!g2033) & (g2034)));
	assign g5040 = (((!sk[12]) & (!g2921) & (!g3087) & (g2566)) + ((!sk[12]) & (!g2921) & (g3087) & (!g2566)) + ((!sk[12]) & (!g2921) & (g3087) & (g2566)) + ((!sk[12]) & (g2921) & (!g3087) & (g2566)) + ((!sk[12]) & (g2921) & (g3087) & (!g2566)) + ((!sk[12]) & (g2921) & (g3087) & (g2566)) + ((sk[12]) & (!g2921) & (!g3087) & (g2566)) + ((sk[12]) & (!g2921) & (g3087) & (g2566)) + ((sk[12]) & (g2921) & (g3087) & (!g2566)) + ((sk[12]) & (g2921) & (g3087) & (g2566)));
	assign g2567 = (((!sk[13]) & (!g773) & (!g865) & (g2545)) + ((!sk[13]) & (!g773) & (g865) & (!g2545)) + ((!sk[13]) & (!g773) & (g865) & (g2545)) + ((!sk[13]) & (g773) & (!g865) & (g2545)) + ((!sk[13]) & (g773) & (g865) & (!g2545)) + ((!sk[13]) & (g773) & (g865) & (g2545)) + ((sk[13]) & (!g773) & (g865) & (!g2545)) + ((sk[13]) & (g773) & (!g865) & (!g2545)) + ((sk[13]) & (g773) & (g865) & (!g2545)) + ((sk[13]) & (g773) & (g865) & (g2545)));
	assign g2568 = (((!g820) & (!g2033) & (!g2034) & (!g912) & (g2566) & (!g2567)) + ((!g820) & (!g2033) & (!g2034) & (!g912) & (g2566) & (g2567)) + ((!g820) & (!g2033) & (!g2034) & (g912) & (g2566) & (!g2567)) + ((!g820) & (!g2033) & (!g2034) & (g912) & (g2566) & (g2567)) + ((!g820) & (g2033) & (!g2034) & (!g912) & (!g2566) & (g2567)) + ((!g820) & (g2033) & (!g2034) & (!g912) & (g2566) & (g2567)) + ((!g820) & (g2033) & (!g2034) & (g912) & (!g2566) & (!g2567)) + ((!g820) & (g2033) & (!g2034) & (g912) & (g2566) & (!g2567)) + ((g820) & (!g2033) & (!g2034) & (!g912) & (g2566) & (!g2567)) + ((g820) & (!g2033) & (!g2034) & (!g912) & (g2566) & (g2567)) + ((g820) & (!g2033) & (!g2034) & (g912) & (g2566) & (!g2567)) + ((g820) & (!g2033) & (!g2034) & (g912) & (g2566) & (g2567)) + ((g820) & (g2033) & (!g2034) & (!g912) & (!g2566) & (!g2567)) + ((g820) & (g2033) & (!g2034) & (!g912) & (g2566) & (!g2567)) + ((g820) & (g2033) & (!g2034) & (g912) & (!g2566) & (g2567)) + ((g820) & (g2033) & (!g2034) & (g912) & (g2566) & (g2567)));
	assign g2569 = (((g2329) & (!g2029) & (g2408) & (!g2564) & (!g2565) & (g2568)) + ((g2329) & (!g2029) & (g2408) & (!g2564) & (g2565) & (!g2568)) + ((g2329) & (!g2029) & (g2408) & (!g2564) & (g2565) & (g2568)) + ((g2329) & (!g2029) & (g2408) & (g2564) & (!g2565) & (g2568)) + ((g2329) & (!g2029) & (g2408) & (g2564) & (g2565) & (!g2568)) + ((g2329) & (!g2029) & (g2408) & (g2564) & (g2565) & (g2568)) + ((g2329) & (g2029) & (g2408) & (g2564) & (!g2565) & (!g2568)) + ((g2329) & (g2029) & (g2408) & (g2564) & (!g2565) & (g2568)) + ((g2329) & (g2029) & (g2408) & (g2564) & (g2565) & (!g2568)) + ((g2329) & (g2029) & (g2408) & (g2564) & (g2565) & (g2568)));
	assign g2571 = (((!g2083) & (!g2084) & (!g2551) & (!g2552) & (!g2553) & (g2570)) + ((!g2083) & (!g2084) & (!g2551) & (!g2552) & (g2553) & (g2570)) + ((!g2083) & (!g2084) & (!g2551) & (g2552) & (!g2553) & (g2570)) + ((!g2083) & (!g2084) & (!g2551) & (g2552) & (g2553) & (g2570)) + ((!g2083) & (!g2084) & (g2551) & (!g2552) & (!g2553) & (g2570)) + ((!g2083) & (!g2084) & (g2551) & (!g2552) & (g2553) & (!g2570)) + ((!g2083) & (!g2084) & (g2551) & (g2552) & (!g2553) & (!g2570)) + ((!g2083) & (!g2084) & (g2551) & (g2552) & (g2553) & (!g2570)) + ((!g2083) & (g2084) & (!g2551) & (!g2552) & (!g2553) & (!g2570)) + ((!g2083) & (g2084) & (!g2551) & (!g2552) & (g2553) & (!g2570)) + ((!g2083) & (g2084) & (!g2551) & (g2552) & (!g2553) & (!g2570)) + ((!g2083) & (g2084) & (!g2551) & (g2552) & (g2553) & (!g2570)) + ((!g2083) & (g2084) & (g2551) & (!g2552) & (!g2553) & (!g2570)) + ((!g2083) & (g2084) & (g2551) & (!g2552) & (g2553) & (g2570)) + ((!g2083) & (g2084) & (g2551) & (g2552) & (!g2553) & (g2570)) + ((!g2083) & (g2084) & (g2551) & (g2552) & (g2553) & (g2570)) + ((g2083) & (!g2084) & (!g2551) & (!g2552) & (!g2553) & (g2570)) + ((g2083) & (!g2084) & (!g2551) & (!g2552) & (g2553) & (!g2570)) + ((g2083) & (!g2084) & (!g2551) & (g2552) & (!g2553) & (!g2570)) + ((g2083) & (!g2084) & (!g2551) & (g2552) & (g2553) & (!g2570)) + ((g2083) & (!g2084) & (g2551) & (!g2552) & (!g2553) & (!g2570)) + ((g2083) & (!g2084) & (g2551) & (!g2552) & (g2553) & (!g2570)) + ((g2083) & (!g2084) & (g2551) & (g2552) & (!g2553) & (!g2570)) + ((g2083) & (!g2084) & (g2551) & (g2552) & (g2553) & (!g2570)) + ((g2083) & (g2084) & (!g2551) & (!g2552) & (!g2553) & (!g2570)) + ((g2083) & (g2084) & (!g2551) & (!g2552) & (g2553) & (g2570)) + ((g2083) & (g2084) & (!g2551) & (g2552) & (!g2553) & (g2570)) + ((g2083) & (g2084) & (!g2551) & (g2552) & (g2553) & (g2570)) + ((g2083) & (g2084) & (g2551) & (!g2552) & (!g2553) & (g2570)) + ((g2083) & (g2084) & (g2551) & (!g2552) & (g2553) & (g2570)) + ((g2083) & (g2084) & (g2551) & (g2552) & (!g2553) & (g2570)) + ((g2083) & (g2084) & (g2551) & (g2552) & (g2553) & (g2570)));
	assign g2572 = (((!sk[17]) & (g2556) & (!g2557)) + ((!sk[17]) & (g2556) & (g2557)) + ((sk[17]) & (!g2556) & (g2557)) + ((sk[17]) & (g2556) & (!g2557)));
	assign g2573 = (((!g2509) & (!g2510) & (!g2511) & (g2533) & (g2534) & (g2572)) + ((!g2509) & (!g2510) & (g2511) & (!g2533) & (g2534) & (g2572)) + ((!g2509) & (!g2510) & (g2511) & (g2533) & (!g2534) & (g2572)) + ((!g2509) & (!g2510) & (g2511) & (g2533) & (g2534) & (g2572)) + ((!g2509) & (g2510) & (!g2511) & (!g2533) & (g2534) & (g2572)) + ((!g2509) & (g2510) & (!g2511) & (g2533) & (!g2534) & (g2572)) + ((!g2509) & (g2510) & (!g2511) & (g2533) & (g2534) & (g2572)) + ((!g2509) & (g2510) & (g2511) & (!g2533) & (g2534) & (g2572)) + ((!g2509) & (g2510) & (g2511) & (g2533) & (!g2534) & (g2572)) + ((!g2509) & (g2510) & (g2511) & (g2533) & (g2534) & (g2572)) + ((g2509) & (!g2510) & (!g2511) & (g2533) & (g2534) & (g2572)) + ((g2509) & (!g2510) & (g2511) & (g2533) & (g2534) & (g2572)) + ((g2509) & (g2510) & (!g2511) & (g2533) & (g2534) & (g2572)) + ((g2509) & (g2510) & (g2511) & (!g2533) & (g2534) & (g2572)) + ((g2509) & (g2510) & (g2511) & (g2533) & (!g2534) & (g2572)) + ((g2509) & (g2510) & (g2511) & (g2533) & (g2534) & (g2572)));
	assign g2574 = (((g2556) & (!sk[19]) & (!g2557)) + ((g2556) & (!sk[19]) & (g2557)) + ((g2556) & (sk[19]) & (g2557)));
	assign g2575 = (((!sk[20]) & (g2573) & (!g2574)) + ((!sk[20]) & (g2573) & (g2574)) + ((sk[20]) & (!g2573) & (!g2574)));
	assign g2576 = (((!g2551) & (sk[21]) & (g2083)) + ((g2551) & (!sk[21]) & (!g2083)) + ((g2551) & (!sk[21]) & (g2083)));
	assign g2577 = (((!g2570) & (sk[22]) & (!g2084)) + ((g2570) & (!sk[22]) & (!g2084)) + ((g2570) & (!sk[22]) & (g2084)) + ((g2570) & (sk[22]) & (g2084)));
	assign g2578 = (((!g2575) & (!g2576) & (!sk[23]) & (g2577)) + ((!g2575) & (!g2576) & (sk[23]) & (!g2577)) + ((!g2575) & (g2576) & (!sk[23]) & (!g2577)) + ((!g2575) & (g2576) & (!sk[23]) & (g2577)) + ((!g2575) & (g2576) & (sk[23]) & (g2577)) + ((g2575) & (!g2576) & (!sk[23]) & (g2577)) + ((g2575) & (!g2576) & (sk[23]) & (g2577)) + ((g2575) & (g2576) & (!sk[23]) & (!g2577)) + ((g2575) & (g2576) & (!sk[23]) & (g2577)) + ((g2575) & (g2576) & (sk[23]) & (!g2577)));
	assign g2579 = (((!sk[24]) & (g2084) & (!g2570)) + ((!sk[24]) & (g2084) & (g2570)) + ((sk[24]) & (g2084) & (g2570)));
	assign g2580 = (((!g2084) & (!g2083) & (!g2121) & (g2120) & (g2071) & (g2074)) + ((!g2084) & (!g2083) & (g2121) & (!g2120) & (!g2071) & (g2074)) + ((!g2084) & (!g2083) & (g2121) & (g2120) & (!g2071) & (g2074)) + ((!g2084) & (!g2083) & (g2121) & (g2120) & (g2071) & (g2074)) + ((!g2084) & (g2083) & (!g2121) & (!g2120) & (g2071) & (!g2074)) + ((!g2084) & (g2083) & (!g2121) & (g2120) & (g2071) & (!g2074)) + ((!g2084) & (g2083) & (!g2121) & (g2120) & (g2071) & (g2074)) + ((!g2084) & (g2083) & (g2121) & (!g2120) & (!g2071) & (g2074)) + ((!g2084) & (g2083) & (g2121) & (!g2120) & (g2071) & (!g2074)) + ((!g2084) & (g2083) & (g2121) & (g2120) & (!g2071) & (g2074)) + ((!g2084) & (g2083) & (g2121) & (g2120) & (g2071) & (!g2074)) + ((!g2084) & (g2083) & (g2121) & (g2120) & (g2071) & (g2074)) + ((g2084) & (!g2083) & (!g2121) & (!g2120) & (!g2071) & (!g2074)) + ((g2084) & (!g2083) & (!g2121) & (g2120) & (!g2071) & (!g2074)) + ((g2084) & (!g2083) & (!g2121) & (g2120) & (g2071) & (g2074)) + ((g2084) & (!g2083) & (g2121) & (!g2120) & (!g2071) & (!g2074)) + ((g2084) & (!g2083) & (g2121) & (!g2120) & (!g2071) & (g2074)) + ((g2084) & (!g2083) & (g2121) & (g2120) & (!g2071) & (!g2074)) + ((g2084) & (!g2083) & (g2121) & (g2120) & (!g2071) & (g2074)) + ((g2084) & (!g2083) & (g2121) & (g2120) & (g2071) & (g2074)) + ((g2084) & (g2083) & (!g2121) & (!g2120) & (!g2071) & (!g2074)) + ((g2084) & (g2083) & (!g2121) & (!g2120) & (g2071) & (!g2074)) + ((g2084) & (g2083) & (!g2121) & (g2120) & (!g2071) & (!g2074)) + ((g2084) & (g2083) & (!g2121) & (g2120) & (g2071) & (!g2074)) + ((g2084) & (g2083) & (!g2121) & (g2120) & (g2071) & (g2074)) + ((g2084) & (g2083) & (g2121) & (!g2120) & (!g2071) & (!g2074)) + ((g2084) & (g2083) & (g2121) & (!g2120) & (!g2071) & (g2074)) + ((g2084) & (g2083) & (g2121) & (!g2120) & (g2071) & (!g2074)) + ((g2084) & (g2083) & (g2121) & (g2120) & (!g2071) & (!g2074)) + ((g2084) & (g2083) & (g2121) & (g2120) & (!g2071) & (g2074)) + ((g2084) & (g2083) & (g2121) & (g2120) & (g2071) & (!g2074)) + ((g2084) & (g2083) & (g2121) & (g2120) & (g2071) & (g2074)));
	assign g2581 = (((!g2580) & (!g2402) & (!g2490) & (g2296) & (g2076) & (g2077)) + ((!g2580) & (!g2402) & (g2490) & (!g2296) & (!g2076) & (g2077)) + ((!g2580) & (!g2402) & (g2490) & (g2296) & (!g2076) & (g2077)) + ((!g2580) & (!g2402) & (g2490) & (g2296) & (g2076) & (g2077)) + ((!g2580) & (g2402) & (!g2490) & (!g2296) & (g2076) & (!g2077)) + ((!g2580) & (g2402) & (!g2490) & (g2296) & (g2076) & (!g2077)) + ((!g2580) & (g2402) & (!g2490) & (g2296) & (g2076) & (g2077)) + ((!g2580) & (g2402) & (g2490) & (!g2296) & (!g2076) & (g2077)) + ((!g2580) & (g2402) & (g2490) & (!g2296) & (g2076) & (!g2077)) + ((!g2580) & (g2402) & (g2490) & (g2296) & (!g2076) & (g2077)) + ((!g2580) & (g2402) & (g2490) & (g2296) & (g2076) & (!g2077)) + ((!g2580) & (g2402) & (g2490) & (g2296) & (g2076) & (g2077)) + ((g2580) & (!g2402) & (!g2490) & (!g2296) & (!g2076) & (!g2077)) + ((g2580) & (!g2402) & (!g2490) & (g2296) & (!g2076) & (!g2077)) + ((g2580) & (!g2402) & (!g2490) & (g2296) & (g2076) & (g2077)) + ((g2580) & (!g2402) & (g2490) & (!g2296) & (!g2076) & (!g2077)) + ((g2580) & (!g2402) & (g2490) & (!g2296) & (!g2076) & (g2077)) + ((g2580) & (!g2402) & (g2490) & (g2296) & (!g2076) & (!g2077)) + ((g2580) & (!g2402) & (g2490) & (g2296) & (!g2076) & (g2077)) + ((g2580) & (!g2402) & (g2490) & (g2296) & (g2076) & (g2077)) + ((g2580) & (g2402) & (!g2490) & (!g2296) & (!g2076) & (!g2077)) + ((g2580) & (g2402) & (!g2490) & (!g2296) & (g2076) & (!g2077)) + ((g2580) & (g2402) & (!g2490) & (g2296) & (!g2076) & (!g2077)) + ((g2580) & (g2402) & (!g2490) & (g2296) & (g2076) & (!g2077)) + ((g2580) & (g2402) & (!g2490) & (g2296) & (g2076) & (g2077)) + ((g2580) & (g2402) & (g2490) & (!g2296) & (!g2076) & (!g2077)) + ((g2580) & (g2402) & (g2490) & (!g2296) & (!g2076) & (g2077)) + ((g2580) & (g2402) & (g2490) & (!g2296) & (g2076) & (!g2077)) + ((g2580) & (g2402) & (g2490) & (g2296) & (!g2076) & (!g2077)) + ((g2580) & (g2402) & (g2490) & (g2296) & (!g2076) & (g2077)) + ((g2580) & (g2402) & (g2490) & (g2296) & (g2076) & (!g2077)) + ((g2580) & (g2402) & (g2490) & (g2296) & (g2076) & (g2077)));
	assign g2582 = (((!g2581) & (!g2184) & (!g2194) & (g2191) & (g2073) & (g2125)) + ((!g2581) & (!g2184) & (g2194) & (!g2191) & (!g2073) & (g2125)) + ((!g2581) & (!g2184) & (g2194) & (g2191) & (!g2073) & (g2125)) + ((!g2581) & (!g2184) & (g2194) & (g2191) & (g2073) & (g2125)) + ((!g2581) & (g2184) & (!g2194) & (!g2191) & (g2073) & (!g2125)) + ((!g2581) & (g2184) & (!g2194) & (g2191) & (g2073) & (!g2125)) + ((!g2581) & (g2184) & (!g2194) & (g2191) & (g2073) & (g2125)) + ((!g2581) & (g2184) & (g2194) & (!g2191) & (!g2073) & (g2125)) + ((!g2581) & (g2184) & (g2194) & (!g2191) & (g2073) & (!g2125)) + ((!g2581) & (g2184) & (g2194) & (g2191) & (!g2073) & (g2125)) + ((!g2581) & (g2184) & (g2194) & (g2191) & (g2073) & (!g2125)) + ((!g2581) & (g2184) & (g2194) & (g2191) & (g2073) & (g2125)) + ((g2581) & (!g2184) & (!g2194) & (!g2191) & (!g2073) & (!g2125)) + ((g2581) & (!g2184) & (!g2194) & (g2191) & (!g2073) & (!g2125)) + ((g2581) & (!g2184) & (!g2194) & (g2191) & (g2073) & (g2125)) + ((g2581) & (!g2184) & (g2194) & (!g2191) & (!g2073) & (!g2125)) + ((g2581) & (!g2184) & (g2194) & (!g2191) & (!g2073) & (g2125)) + ((g2581) & (!g2184) & (g2194) & (g2191) & (!g2073) & (!g2125)) + ((g2581) & (!g2184) & (g2194) & (g2191) & (!g2073) & (g2125)) + ((g2581) & (!g2184) & (g2194) & (g2191) & (g2073) & (g2125)) + ((g2581) & (g2184) & (!g2194) & (!g2191) & (!g2073) & (!g2125)) + ((g2581) & (g2184) & (!g2194) & (!g2191) & (g2073) & (!g2125)) + ((g2581) & (g2184) & (!g2194) & (g2191) & (!g2073) & (!g2125)) + ((g2581) & (g2184) & (!g2194) & (g2191) & (g2073) & (!g2125)) + ((g2581) & (g2184) & (!g2194) & (g2191) & (g2073) & (g2125)) + ((g2581) & (g2184) & (g2194) & (!g2191) & (!g2073) & (!g2125)) + ((g2581) & (g2184) & (g2194) & (!g2191) & (!g2073) & (g2125)) + ((g2581) & (g2184) & (g2194) & (!g2191) & (g2073) & (!g2125)) + ((g2581) & (g2184) & (g2194) & (g2191) & (!g2073) & (!g2125)) + ((g2581) & (g2184) & (g2194) & (g2191) & (!g2073) & (g2125)) + ((g2581) & (g2184) & (g2194) & (g2191) & (g2073) & (!g2125)) + ((g2581) & (g2184) & (g2194) & (g2191) & (g2073) & (g2125)));
	assign g2583 = (((!g2084) & (!g2570) & (!g2124) & (!g2264) & (!g3526) & (g2582)) + ((!g2084) & (!g2570) & (!g2124) & (!g2264) & (g3526) & (g2582)) + ((!g2084) & (!g2570) & (!g2124) & (g2264) & (g3526) & (!g2582)) + ((!g2084) & (!g2570) & (!g2124) & (g2264) & (g3526) & (g2582)) + ((!g2084) & (g2570) & (!g2124) & (!g2264) & (!g3526) & (g2582)) + ((!g2084) & (g2570) & (!g2124) & (!g2264) & (g3526) & (g2582)) + ((!g2084) & (g2570) & (!g2124) & (g2264) & (g3526) & (!g2582)) + ((!g2084) & (g2570) & (!g2124) & (g2264) & (g3526) & (g2582)) + ((!g2084) & (g2570) & (g2124) & (!g2264) & (!g3526) & (!g2582)) + ((!g2084) & (g2570) & (g2124) & (!g2264) & (!g3526) & (g2582)) + ((!g2084) & (g2570) & (g2124) & (!g2264) & (g3526) & (!g2582)) + ((!g2084) & (g2570) & (g2124) & (!g2264) & (g3526) & (g2582)) + ((!g2084) & (g2570) & (g2124) & (g2264) & (!g3526) & (!g2582)) + ((!g2084) & (g2570) & (g2124) & (g2264) & (!g3526) & (g2582)) + ((!g2084) & (g2570) & (g2124) & (g2264) & (g3526) & (!g2582)) + ((!g2084) & (g2570) & (g2124) & (g2264) & (g3526) & (g2582)) + ((g2084) & (!g2570) & (!g2124) & (!g2264) & (!g3526) & (g2582)) + ((g2084) & (!g2570) & (!g2124) & (!g2264) & (g3526) & (g2582)) + ((g2084) & (!g2570) & (!g2124) & (g2264) & (g3526) & (!g2582)) + ((g2084) & (!g2570) & (!g2124) & (g2264) & (g3526) & (g2582)) + ((g2084) & (!g2570) & (g2124) & (!g2264) & (!g3526) & (!g2582)) + ((g2084) & (!g2570) & (g2124) & (!g2264) & (!g3526) & (g2582)) + ((g2084) & (!g2570) & (g2124) & (!g2264) & (g3526) & (!g2582)) + ((g2084) & (!g2570) & (g2124) & (!g2264) & (g3526) & (g2582)) + ((g2084) & (!g2570) & (g2124) & (g2264) & (!g3526) & (!g2582)) + ((g2084) & (!g2570) & (g2124) & (g2264) & (!g3526) & (g2582)) + ((g2084) & (!g2570) & (g2124) & (g2264) & (g3526) & (!g2582)) + ((g2084) & (!g2570) & (g2124) & (g2264) & (g3526) & (g2582)) + ((g2084) & (g2570) & (!g2124) & (!g2264) & (!g3526) & (g2582)) + ((g2084) & (g2570) & (!g2124) & (!g2264) & (g3526) & (g2582)) + ((g2084) & (g2570) & (!g2124) & (g2264) & (g3526) & (!g2582)) + ((g2084) & (g2570) & (!g2124) & (g2264) & (g3526) & (g2582)) + ((g2084) & (g2570) & (g2124) & (!g2264) & (!g3526) & (!g2582)) + ((g2084) & (g2570) & (g2124) & (!g2264) & (!g3526) & (g2582)) + ((g2084) & (g2570) & (g2124) & (!g2264) & (g3526) & (!g2582)) + ((g2084) & (g2570) & (g2124) & (!g2264) & (g3526) & (g2582)));
	assign g2584 = (((!g912) & (!sk[29]) & (!g2563) & (g960)) + ((!g912) & (!sk[29]) & (g2563) & (!g960)) + ((!g912) & (!sk[29]) & (g2563) & (g960)) + ((!g912) & (sk[29]) & (!g2563) & (g960)) + ((!g912) & (sk[29]) & (g2563) & (g960)) + ((g912) & (!sk[29]) & (!g2563) & (g960)) + ((g912) & (!sk[29]) & (g2563) & (!g960)) + ((g912) & (!sk[29]) & (g2563) & (g960)) + ((g912) & (sk[29]) & (!g2563) & (g960)) + ((g912) & (sk[29]) & (g2563) & (!g960)));
	assign g2585 = (((!sk[30]) & (g2033) & (!g2034)) + ((!sk[30]) & (g2033) & (g2034)) + ((sk[30]) & (g2033) & (!g2034)));
	assign g2586 = (((!g867) & (!g820) & (!g912) & (!g2567) & (g960) & (g2585)) + ((!g867) & (!g820) & (!g912) & (g2567) & (g960) & (g2585)) + ((!g867) & (!g820) & (g912) & (!g2567) & (g960) & (g2585)) + ((!g867) & (!g820) & (g912) & (g2567) & (!g960) & (g2585)) + ((!g867) & (g820) & (!g912) & (!g2567) & (g960) & (g2585)) + ((!g867) & (g820) & (!g912) & (g2567) & (!g960) & (g2585)) + ((!g867) & (g820) & (g912) & (!g2567) & (!g960) & (g2585)) + ((!g867) & (g820) & (g912) & (g2567) & (!g960) & (g2585)) + ((g867) & (!g820) & (!g912) & (!g2567) & (!g960) & (g2585)) + ((g867) & (!g820) & (!g912) & (g2567) & (!g960) & (g2585)) + ((g867) & (!g820) & (g912) & (!g2567) & (!g960) & (g2585)) + ((g867) & (!g820) & (g912) & (g2567) & (g960) & (g2585)) + ((g867) & (g820) & (!g912) & (!g2567) & (!g960) & (g2585)) + ((g867) & (g820) & (!g912) & (g2567) & (g960) & (g2585)) + ((g867) & (g820) & (g912) & (!g2567) & (g960) & (g2585)) + ((g867) & (g820) & (g912) & (g2567) & (g960) & (g2585)));
	assign g5041 = (((!g2921) & (!sk[32]) & (!g3213) & (g2587)) + ((!g2921) & (!sk[32]) & (g3213) & (!g2587)) + ((!g2921) & (!sk[32]) & (g3213) & (g2587)) + ((!g2921) & (sk[32]) & (!g3213) & (g2587)) + ((!g2921) & (sk[32]) & (g3213) & (g2587)) + ((g2921) & (!sk[32]) & (!g3213) & (g2587)) + ((g2921) & (!sk[32]) & (g3213) & (!g2587)) + ((g2921) & (!sk[32]) & (g3213) & (g2587)) + ((g2921) & (sk[32]) & (g3213) & (!g2587)) + ((g2921) & (sk[32]) & (g3213) & (g2587)));
	assign g2588 = (((!g1824) & (!g2033) & (!sk[33]) & (!g2034) & (g2587)) + ((!g1824) & (!g2033) & (!sk[33]) & (g2034) & (!g2587)) + ((!g1824) & (!g2033) & (!sk[33]) & (g2034) & (g2587)) + ((!g1824) & (!g2033) & (sk[33]) & (!g2034) & (g2587)) + ((!g1824) & (g2033) & (!sk[33]) & (!g2034) & (!g2587)) + ((!g1824) & (g2033) & (!sk[33]) & (!g2034) & (g2587)) + ((!g1824) & (g2033) & (!sk[33]) & (g2034) & (!g2587)) + ((!g1824) & (g2033) & (!sk[33]) & (g2034) & (g2587)) + ((g1824) & (!g2033) & (!sk[33]) & (!g2034) & (g2587)) + ((g1824) & (!g2033) & (!sk[33]) & (g2034) & (!g2587)) + ((g1824) & (!g2033) & (!sk[33]) & (g2034) & (g2587)) + ((g1824) & (!g2033) & (sk[33]) & (!g2034) & (g2587)) + ((g1824) & (!g2033) & (sk[33]) & (g2034) & (!g2587)) + ((g1824) & (!g2033) & (sk[33]) & (g2034) & (g2587)) + ((g1824) & (g2033) & (!sk[33]) & (!g2034) & (!g2587)) + ((g1824) & (g2033) & (!sk[33]) & (!g2034) & (g2587)) + ((g1824) & (g2033) & (!sk[33]) & (g2034) & (!g2587)) + ((g1824) & (g2033) & (!sk[33]) & (g2034) & (g2587)));
	assign g2589 = (((g2329) & (!g2029) & (g2408) & (!g2584) & (!g2586) & (g2588)) + ((g2329) & (!g2029) & (g2408) & (!g2584) & (g2586) & (!g2588)) + ((g2329) & (!g2029) & (g2408) & (!g2584) & (g2586) & (g2588)) + ((g2329) & (!g2029) & (g2408) & (g2584) & (!g2586) & (g2588)) + ((g2329) & (!g2029) & (g2408) & (g2584) & (g2586) & (!g2588)) + ((g2329) & (!g2029) & (g2408) & (g2584) & (g2586) & (g2588)) + ((g2329) & (g2029) & (g2408) & (g2584) & (!g2586) & (!g2588)) + ((g2329) & (g2029) & (g2408) & (g2584) & (!g2586) & (g2588)) + ((g2329) & (g2029) & (g2408) & (g2584) & (g2586) & (!g2588)) + ((g2329) & (g2029) & (g2408) & (g2584) & (g2586) & (g2588)));
	assign g2591 = (((!g2083) & (!g2084) & (g2551) & (!g2552) & (g2553) & (g2570)) + ((!g2083) & (!g2084) & (g2551) & (g2552) & (!g2553) & (g2570)) + ((!g2083) & (!g2084) & (g2551) & (g2552) & (g2553) & (g2570)) + ((!g2083) & (g2084) & (!g2551) & (!g2552) & (!g2553) & (g2570)) + ((!g2083) & (g2084) & (!g2551) & (!g2552) & (g2553) & (g2570)) + ((!g2083) & (g2084) & (!g2551) & (g2552) & (!g2553) & (g2570)) + ((!g2083) & (g2084) & (!g2551) & (g2552) & (g2553) & (g2570)) + ((!g2083) & (g2084) & (g2551) & (!g2552) & (!g2553) & (g2570)) + ((!g2083) & (g2084) & (g2551) & (!g2552) & (g2553) & (!g2570)) + ((!g2083) & (g2084) & (g2551) & (!g2552) & (g2553) & (g2570)) + ((!g2083) & (g2084) & (g2551) & (g2552) & (!g2553) & (!g2570)) + ((!g2083) & (g2084) & (g2551) & (g2552) & (!g2553) & (g2570)) + ((!g2083) & (g2084) & (g2551) & (g2552) & (g2553) & (!g2570)) + ((!g2083) & (g2084) & (g2551) & (g2552) & (g2553) & (g2570)) + ((g2083) & (!g2084) & (!g2551) & (!g2552) & (g2553) & (g2570)) + ((g2083) & (!g2084) & (!g2551) & (g2552) & (!g2553) & (g2570)) + ((g2083) & (!g2084) & (!g2551) & (g2552) & (g2553) & (g2570)) + ((g2083) & (!g2084) & (g2551) & (!g2552) & (!g2553) & (g2570)) + ((g2083) & (!g2084) & (g2551) & (!g2552) & (g2553) & (g2570)) + ((g2083) & (!g2084) & (g2551) & (g2552) & (!g2553) & (g2570)) + ((g2083) & (!g2084) & (g2551) & (g2552) & (g2553) & (g2570)) + ((g2083) & (g2084) & (!g2551) & (!g2552) & (!g2553) & (g2570)) + ((g2083) & (g2084) & (!g2551) & (!g2552) & (g2553) & (!g2570)) + ((g2083) & (g2084) & (!g2551) & (!g2552) & (g2553) & (g2570)) + ((g2083) & (g2084) & (!g2551) & (g2552) & (!g2553) & (!g2570)) + ((g2083) & (g2084) & (!g2551) & (g2552) & (!g2553) & (g2570)) + ((g2083) & (g2084) & (!g2551) & (g2552) & (g2553) & (!g2570)) + ((g2083) & (g2084) & (!g2551) & (g2552) & (g2553) & (g2570)) + ((g2083) & (g2084) & (g2551) & (!g2552) & (!g2553) & (!g2570)) + ((g2083) & (g2084) & (g2551) & (!g2552) & (!g2553) & (g2570)) + ((g2083) & (g2084) & (g2551) & (!g2552) & (g2553) & (!g2570)) + ((g2083) & (g2084) & (g2551) & (!g2552) & (g2553) & (g2570)) + ((g2083) & (g2084) & (g2551) & (g2552) & (!g2553) & (!g2570)) + ((g2083) & (g2084) & (g2551) & (g2552) & (!g2553) & (g2570)) + ((g2083) & (g2084) & (g2551) & (g2552) & (g2553) & (!g2570)) + ((g2083) & (g2084) & (g2551) & (g2552) & (g2553) & (g2570)));
	assign g2592 = (((!g2570) & (sk[36]) & (g2084)) + ((g2570) & (!sk[36]) & (!g2084)) + ((g2570) & (!sk[36]) & (g2084)));
	assign g2593 = (((!g2590) & (sk[37]) & (!g2085)) + ((g2590) & (!sk[37]) & (!g2085)) + ((g2590) & (!sk[37]) & (g2085)) + ((g2590) & (sk[37]) & (g2085)));
	assign g2594 = (((!g2575) & (!g2576) & (!sk[38]) & (!g2577) & (g2592) & (!g2593)) + ((!g2575) & (!g2576) & (!sk[38]) & (!g2577) & (g2592) & (g2593)) + ((!g2575) & (!g2576) & (!sk[38]) & (g2577) & (!g2592) & (!g2593)) + ((!g2575) & (!g2576) & (!sk[38]) & (g2577) & (!g2592) & (g2593)) + ((!g2575) & (!g2576) & (!sk[38]) & (g2577) & (g2592) & (!g2593)) + ((!g2575) & (!g2576) & (!sk[38]) & (g2577) & (g2592) & (g2593)) + ((!g2575) & (!g2576) & (sk[38]) & (!g2577) & (!g2592) & (g2593)) + ((!g2575) & (!g2576) & (sk[38]) & (!g2577) & (g2592) & (!g2593)) + ((!g2575) & (!g2576) & (sk[38]) & (g2577) & (!g2592) & (!g2593)) + ((!g2575) & (!g2576) & (sk[38]) & (g2577) & (g2592) & (g2593)) + ((!g2575) & (g2576) & (!sk[38]) & (!g2577) & (!g2592) & (!g2593)) + ((!g2575) & (g2576) & (!sk[38]) & (!g2577) & (!g2592) & (g2593)) + ((!g2575) & (g2576) & (!sk[38]) & (!g2577) & (g2592) & (!g2593)) + ((!g2575) & (g2576) & (!sk[38]) & (!g2577) & (g2592) & (g2593)) + ((!g2575) & (g2576) & (!sk[38]) & (g2577) & (!g2592) & (!g2593)) + ((!g2575) & (g2576) & (!sk[38]) & (g2577) & (!g2592) & (g2593)) + ((!g2575) & (g2576) & (!sk[38]) & (g2577) & (g2592) & (!g2593)) + ((!g2575) & (g2576) & (!sk[38]) & (g2577) & (g2592) & (g2593)) + ((!g2575) & (g2576) & (sk[38]) & (!g2577) & (!g2592) & (!g2593)) + ((!g2575) & (g2576) & (sk[38]) & (!g2577) & (g2592) & (g2593)) + ((!g2575) & (g2576) & (sk[38]) & (g2577) & (!g2592) & (!g2593)) + ((!g2575) & (g2576) & (sk[38]) & (g2577) & (g2592) & (g2593)) + ((g2575) & (!g2576) & (!sk[38]) & (!g2577) & (g2592) & (!g2593)) + ((g2575) & (!g2576) & (!sk[38]) & (!g2577) & (g2592) & (g2593)) + ((g2575) & (!g2576) & (!sk[38]) & (g2577) & (!g2592) & (!g2593)) + ((g2575) & (!g2576) & (!sk[38]) & (g2577) & (!g2592) & (g2593)) + ((g2575) & (!g2576) & (!sk[38]) & (g2577) & (g2592) & (!g2593)) + ((g2575) & (!g2576) & (!sk[38]) & (g2577) & (g2592) & (g2593)) + ((g2575) & (!g2576) & (sk[38]) & (!g2577) & (!g2592) & (g2593)) + ((g2575) & (!g2576) & (sk[38]) & (!g2577) & (g2592) & (!g2593)) + ((g2575) & (!g2576) & (sk[38]) & (g2577) & (!g2592) & (g2593)) + ((g2575) & (!g2576) & (sk[38]) & (g2577) & (g2592) & (!g2593)) + ((g2575) & (g2576) & (!sk[38]) & (!g2577) & (!g2592) & (!g2593)) + ((g2575) & (g2576) & (!sk[38]) & (!g2577) & (!g2592) & (g2593)) + ((g2575) & (g2576) & (!sk[38]) & (!g2577) & (g2592) & (!g2593)) + ((g2575) & (g2576) & (!sk[38]) & (!g2577) & (g2592) & (g2593)) + ((g2575) & (g2576) & (!sk[38]) & (g2577) & (!g2592) & (!g2593)) + ((g2575) & (g2576) & (!sk[38]) & (g2577) & (!g2592) & (g2593)) + ((g2575) & (g2576) & (!sk[38]) & (g2577) & (g2592) & (!g2593)) + ((g2575) & (g2576) & (!sk[38]) & (g2577) & (g2592) & (g2593)) + ((g2575) & (g2576) & (sk[38]) & (!g2577) & (!g2592) & (g2593)) + ((g2575) & (g2576) & (sk[38]) & (!g2577) & (g2592) & (!g2593)) + ((g2575) & (g2576) & (sk[38]) & (g2577) & (!g2592) & (!g2593)) + ((g2575) & (g2576) & (sk[38]) & (g2577) & (g2592) & (g2593)));
	assign g2595 = (((!g2085) & (!g2084) & (!g2083) & (g2121) & (g2071) & (g2074)) + ((!g2085) & (!g2084) & (g2083) & (!g2121) & (!g2071) & (g2074)) + ((!g2085) & (!g2084) & (g2083) & (g2121) & (!g2071) & (g2074)) + ((!g2085) & (!g2084) & (g2083) & (g2121) & (g2071) & (g2074)) + ((!g2085) & (g2084) & (!g2083) & (!g2121) & (g2071) & (!g2074)) + ((!g2085) & (g2084) & (!g2083) & (g2121) & (g2071) & (!g2074)) + ((!g2085) & (g2084) & (!g2083) & (g2121) & (g2071) & (g2074)) + ((!g2085) & (g2084) & (g2083) & (!g2121) & (!g2071) & (g2074)) + ((!g2085) & (g2084) & (g2083) & (!g2121) & (g2071) & (!g2074)) + ((!g2085) & (g2084) & (g2083) & (g2121) & (!g2071) & (g2074)) + ((!g2085) & (g2084) & (g2083) & (g2121) & (g2071) & (!g2074)) + ((!g2085) & (g2084) & (g2083) & (g2121) & (g2071) & (g2074)) + ((g2085) & (!g2084) & (!g2083) & (!g2121) & (!g2071) & (!g2074)) + ((g2085) & (!g2084) & (!g2083) & (g2121) & (!g2071) & (!g2074)) + ((g2085) & (!g2084) & (!g2083) & (g2121) & (g2071) & (g2074)) + ((g2085) & (!g2084) & (g2083) & (!g2121) & (!g2071) & (!g2074)) + ((g2085) & (!g2084) & (g2083) & (!g2121) & (!g2071) & (g2074)) + ((g2085) & (!g2084) & (g2083) & (g2121) & (!g2071) & (!g2074)) + ((g2085) & (!g2084) & (g2083) & (g2121) & (!g2071) & (g2074)) + ((g2085) & (!g2084) & (g2083) & (g2121) & (g2071) & (g2074)) + ((g2085) & (g2084) & (!g2083) & (!g2121) & (!g2071) & (!g2074)) + ((g2085) & (g2084) & (!g2083) & (!g2121) & (g2071) & (!g2074)) + ((g2085) & (g2084) & (!g2083) & (g2121) & (!g2071) & (!g2074)) + ((g2085) & (g2084) & (!g2083) & (g2121) & (g2071) & (!g2074)) + ((g2085) & (g2084) & (!g2083) & (g2121) & (g2071) & (g2074)) + ((g2085) & (g2084) & (g2083) & (!g2121) & (!g2071) & (!g2074)) + ((g2085) & (g2084) & (g2083) & (!g2121) & (!g2071) & (g2074)) + ((g2085) & (g2084) & (g2083) & (!g2121) & (g2071) & (!g2074)) + ((g2085) & (g2084) & (g2083) & (g2121) & (!g2071) & (!g2074)) + ((g2085) & (g2084) & (g2083) & (g2121) & (!g2071) & (g2074)) + ((g2085) & (g2084) & (g2083) & (g2121) & (g2071) & (!g2074)) + ((g2085) & (g2084) & (g2083) & (g2121) & (g2071) & (g2074)));
	assign g2596 = (((!g2595) & (!g2426) & (!g2514) & (g2320) & (g2076) & (g2077)) + ((!g2595) & (!g2426) & (g2514) & (!g2320) & (!g2076) & (g2077)) + ((!g2595) & (!g2426) & (g2514) & (g2320) & (!g2076) & (g2077)) + ((!g2595) & (!g2426) & (g2514) & (g2320) & (g2076) & (g2077)) + ((!g2595) & (g2426) & (!g2514) & (!g2320) & (g2076) & (!g2077)) + ((!g2595) & (g2426) & (!g2514) & (g2320) & (g2076) & (!g2077)) + ((!g2595) & (g2426) & (!g2514) & (g2320) & (g2076) & (g2077)) + ((!g2595) & (g2426) & (g2514) & (!g2320) & (!g2076) & (g2077)) + ((!g2595) & (g2426) & (g2514) & (!g2320) & (g2076) & (!g2077)) + ((!g2595) & (g2426) & (g2514) & (g2320) & (!g2076) & (g2077)) + ((!g2595) & (g2426) & (g2514) & (g2320) & (g2076) & (!g2077)) + ((!g2595) & (g2426) & (g2514) & (g2320) & (g2076) & (g2077)) + ((g2595) & (!g2426) & (!g2514) & (!g2320) & (!g2076) & (!g2077)) + ((g2595) & (!g2426) & (!g2514) & (g2320) & (!g2076) & (!g2077)) + ((g2595) & (!g2426) & (!g2514) & (g2320) & (g2076) & (g2077)) + ((g2595) & (!g2426) & (g2514) & (!g2320) & (!g2076) & (!g2077)) + ((g2595) & (!g2426) & (g2514) & (!g2320) & (!g2076) & (g2077)) + ((g2595) & (!g2426) & (g2514) & (g2320) & (!g2076) & (!g2077)) + ((g2595) & (!g2426) & (g2514) & (g2320) & (!g2076) & (g2077)) + ((g2595) & (!g2426) & (g2514) & (g2320) & (g2076) & (g2077)) + ((g2595) & (g2426) & (!g2514) & (!g2320) & (!g2076) & (!g2077)) + ((g2595) & (g2426) & (!g2514) & (!g2320) & (g2076) & (!g2077)) + ((g2595) & (g2426) & (!g2514) & (g2320) & (!g2076) & (!g2077)) + ((g2595) & (g2426) & (!g2514) & (g2320) & (g2076) & (!g2077)) + ((g2595) & (g2426) & (!g2514) & (g2320) & (g2076) & (g2077)) + ((g2595) & (g2426) & (g2514) & (!g2320) & (!g2076) & (!g2077)) + ((g2595) & (g2426) & (g2514) & (!g2320) & (!g2076) & (g2077)) + ((g2595) & (g2426) & (g2514) & (!g2320) & (g2076) & (!g2077)) + ((g2595) & (g2426) & (g2514) & (g2320) & (!g2076) & (!g2077)) + ((g2595) & (g2426) & (g2514) & (g2320) & (!g2076) & (g2077)) + ((g2595) & (g2426) & (g2514) & (g2320) & (g2076) & (!g2077)) + ((g2595) & (g2426) & (g2514) & (g2320) & (g2076) & (g2077)));
	assign g2597 = (((!g2596) & (!g2212) & (!g2219) & (g2191) & (g2073) & (g2125)) + ((!g2596) & (!g2212) & (g2219) & (!g2191) & (!g2073) & (g2125)) + ((!g2596) & (!g2212) & (g2219) & (g2191) & (!g2073) & (g2125)) + ((!g2596) & (!g2212) & (g2219) & (g2191) & (g2073) & (g2125)) + ((!g2596) & (g2212) & (!g2219) & (!g2191) & (g2073) & (!g2125)) + ((!g2596) & (g2212) & (!g2219) & (g2191) & (g2073) & (!g2125)) + ((!g2596) & (g2212) & (!g2219) & (g2191) & (g2073) & (g2125)) + ((!g2596) & (g2212) & (g2219) & (!g2191) & (!g2073) & (g2125)) + ((!g2596) & (g2212) & (g2219) & (!g2191) & (g2073) & (!g2125)) + ((!g2596) & (g2212) & (g2219) & (g2191) & (!g2073) & (g2125)) + ((!g2596) & (g2212) & (g2219) & (g2191) & (g2073) & (!g2125)) + ((!g2596) & (g2212) & (g2219) & (g2191) & (g2073) & (g2125)) + ((g2596) & (!g2212) & (!g2219) & (!g2191) & (!g2073) & (!g2125)) + ((g2596) & (!g2212) & (!g2219) & (g2191) & (!g2073) & (!g2125)) + ((g2596) & (!g2212) & (!g2219) & (g2191) & (g2073) & (g2125)) + ((g2596) & (!g2212) & (g2219) & (!g2191) & (!g2073) & (!g2125)) + ((g2596) & (!g2212) & (g2219) & (!g2191) & (!g2073) & (g2125)) + ((g2596) & (!g2212) & (g2219) & (g2191) & (!g2073) & (!g2125)) + ((g2596) & (!g2212) & (g2219) & (g2191) & (!g2073) & (g2125)) + ((g2596) & (!g2212) & (g2219) & (g2191) & (g2073) & (g2125)) + ((g2596) & (g2212) & (!g2219) & (!g2191) & (!g2073) & (!g2125)) + ((g2596) & (g2212) & (!g2219) & (!g2191) & (g2073) & (!g2125)) + ((g2596) & (g2212) & (!g2219) & (g2191) & (!g2073) & (!g2125)) + ((g2596) & (g2212) & (!g2219) & (g2191) & (g2073) & (!g2125)) + ((g2596) & (g2212) & (!g2219) & (g2191) & (g2073) & (g2125)) + ((g2596) & (g2212) & (g2219) & (!g2191) & (!g2073) & (!g2125)) + ((g2596) & (g2212) & (g2219) & (!g2191) & (!g2073) & (g2125)) + ((g2596) & (g2212) & (g2219) & (!g2191) & (g2073) & (!g2125)) + ((g2596) & (g2212) & (g2219) & (g2191) & (!g2073) & (!g2125)) + ((g2596) & (g2212) & (g2219) & (g2191) & (!g2073) & (g2125)) + ((g2596) & (g2212) & (g2219) & (g2191) & (g2073) & (!g2125)) + ((g2596) & (g2212) & (g2219) & (g2191) & (g2073) & (g2125)));
	assign g2598 = (((!g2085) & (!g2590) & (!g2124) & (!g2264) & (!g3502) & (g2597)) + ((!g2085) & (!g2590) & (!g2124) & (!g2264) & (g3502) & (g2597)) + ((!g2085) & (!g2590) & (!g2124) & (g2264) & (g3502) & (!g2597)) + ((!g2085) & (!g2590) & (!g2124) & (g2264) & (g3502) & (g2597)) + ((!g2085) & (g2590) & (!g2124) & (!g2264) & (!g3502) & (g2597)) + ((!g2085) & (g2590) & (!g2124) & (!g2264) & (g3502) & (g2597)) + ((!g2085) & (g2590) & (!g2124) & (g2264) & (g3502) & (!g2597)) + ((!g2085) & (g2590) & (!g2124) & (g2264) & (g3502) & (g2597)) + ((!g2085) & (g2590) & (g2124) & (!g2264) & (!g3502) & (!g2597)) + ((!g2085) & (g2590) & (g2124) & (!g2264) & (!g3502) & (g2597)) + ((!g2085) & (g2590) & (g2124) & (!g2264) & (g3502) & (!g2597)) + ((!g2085) & (g2590) & (g2124) & (!g2264) & (g3502) & (g2597)) + ((!g2085) & (g2590) & (g2124) & (g2264) & (!g3502) & (!g2597)) + ((!g2085) & (g2590) & (g2124) & (g2264) & (!g3502) & (g2597)) + ((!g2085) & (g2590) & (g2124) & (g2264) & (g3502) & (!g2597)) + ((!g2085) & (g2590) & (g2124) & (g2264) & (g3502) & (g2597)) + ((g2085) & (!g2590) & (!g2124) & (!g2264) & (!g3502) & (g2597)) + ((g2085) & (!g2590) & (!g2124) & (!g2264) & (g3502) & (g2597)) + ((g2085) & (!g2590) & (!g2124) & (g2264) & (g3502) & (!g2597)) + ((g2085) & (!g2590) & (!g2124) & (g2264) & (g3502) & (g2597)) + ((g2085) & (!g2590) & (g2124) & (!g2264) & (!g3502) & (!g2597)) + ((g2085) & (!g2590) & (g2124) & (!g2264) & (!g3502) & (g2597)) + ((g2085) & (!g2590) & (g2124) & (!g2264) & (g3502) & (!g2597)) + ((g2085) & (!g2590) & (g2124) & (!g2264) & (g3502) & (g2597)) + ((g2085) & (!g2590) & (g2124) & (g2264) & (!g3502) & (!g2597)) + ((g2085) & (!g2590) & (g2124) & (g2264) & (!g3502) & (g2597)) + ((g2085) & (!g2590) & (g2124) & (g2264) & (g3502) & (!g2597)) + ((g2085) & (!g2590) & (g2124) & (g2264) & (g3502) & (g2597)) + ((g2085) & (g2590) & (!g2124) & (!g2264) & (!g3502) & (g2597)) + ((g2085) & (g2590) & (!g2124) & (!g2264) & (g3502) & (g2597)) + ((g2085) & (g2590) & (!g2124) & (g2264) & (g3502) & (!g2597)) + ((g2085) & (g2590) & (!g2124) & (g2264) & (g3502) & (g2597)) + ((g2085) & (g2590) & (g2124) & (!g2264) & (!g3502) & (!g2597)) + ((g2085) & (g2590) & (g2124) & (!g2264) & (!g3502) & (g2597)) + ((g2085) & (g2590) & (g2124) & (!g2264) & (g3502) & (!g2597)) + ((g2085) & (g2590) & (g2124) & (!g2264) & (g3502) & (g2597)));
	assign g2599 = (((!g912) & (!g2563) & (!g960) & (!sk[43]) & (g1005)) + ((!g912) & (!g2563) & (!g960) & (sk[43]) & (g1005)) + ((!g912) & (!g2563) & (g960) & (!sk[43]) & (!g1005)) + ((!g912) & (!g2563) & (g960) & (!sk[43]) & (g1005)) + ((!g912) & (!g2563) & (g960) & (sk[43]) & (g1005)) + ((!g912) & (g2563) & (!g960) & (!sk[43]) & (!g1005)) + ((!g912) & (g2563) & (!g960) & (!sk[43]) & (g1005)) + ((!g912) & (g2563) & (!g960) & (sk[43]) & (g1005)) + ((!g912) & (g2563) & (g960) & (!sk[43]) & (!g1005)) + ((!g912) & (g2563) & (g960) & (!sk[43]) & (g1005)) + ((!g912) & (g2563) & (g960) & (sk[43]) & (g1005)) + ((g912) & (!g2563) & (!g960) & (!sk[43]) & (g1005)) + ((g912) & (!g2563) & (!g960) & (sk[43]) & (g1005)) + ((g912) & (!g2563) & (g960) & (!sk[43]) & (!g1005)) + ((g912) & (!g2563) & (g960) & (!sk[43]) & (g1005)) + ((g912) & (!g2563) & (g960) & (sk[43]) & (g1005)) + ((g912) & (g2563) & (!g960) & (!sk[43]) & (!g1005)) + ((g912) & (g2563) & (!g960) & (!sk[43]) & (g1005)) + ((g912) & (g2563) & (!g960) & (sk[43]) & (g1005)) + ((g912) & (g2563) & (g960) & (!sk[43]) & (!g1005)) + ((g912) & (g2563) & (g960) & (!sk[43]) & (g1005)) + ((g912) & (g2563) & (g960) & (sk[43]) & (!g1005)));
	assign g2600 = (((!g867) & (sk[44]) & (g960)) + ((g867) & (!sk[44]) & (!g960)) + ((g867) & (!sk[44]) & (g960)) + ((g867) & (sk[44]) & (!g960)));
	assign g2601 = (((!g820) & (!g773) & (g865) & (!g2545) & (g912) & (g2600)) + ((!g820) & (g773) & (!g865) & (!g2545) & (g912) & (g2600)) + ((!g820) & (g773) & (g865) & (!g2545) & (g912) & (g2600)) + ((!g820) & (g773) & (g865) & (g2545) & (g912) & (g2600)) + ((g820) & (!g773) & (!g865) & (!g2545) & (g912) & (g2600)) + ((g820) & (!g773) & (!g865) & (g2545) & (g912) & (g2600)) + ((g820) & (!g773) & (g865) & (!g2545) & (!g912) & (g2600)) + ((g820) & (!g773) & (g865) & (!g2545) & (g912) & (g2600)) + ((g820) & (!g773) & (g865) & (g2545) & (g912) & (g2600)) + ((g820) & (g773) & (!g865) & (!g2545) & (!g912) & (g2600)) + ((g820) & (g773) & (!g865) & (!g2545) & (g912) & (g2600)) + ((g820) & (g773) & (!g865) & (g2545) & (g912) & (g2600)) + ((g820) & (g773) & (g865) & (!g2545) & (!g912) & (g2600)) + ((g820) & (g773) & (g865) & (!g2545) & (g912) & (g2600)) + ((g820) & (g773) & (g865) & (g2545) & (!g912) & (g2600)) + ((g820) & (g773) & (g865) & (g2545) & (g912) & (g2600)));
	assign g2602 = (((g867) & (!sk[46]) & (!g960)) + ((g867) & (!sk[46]) & (g960)) + ((g867) & (sk[46]) & (g960)));
	assign g2603 = (((!g2601) & (sk[47]) & (!g2602)) + ((g2601) & (!sk[47]) & (!g2602)) + ((g2601) & (!sk[47]) & (g2602)));
	assign g2604 = (((!sk[48]) & (!g165) & (!g2585) & (!g1005) & (g2603)) + ((!sk[48]) & (!g165) & (!g2585) & (g1005) & (!g2603)) + ((!sk[48]) & (!g165) & (!g2585) & (g1005) & (g2603)) + ((!sk[48]) & (!g165) & (g2585) & (!g1005) & (!g2603)) + ((!sk[48]) & (!g165) & (g2585) & (!g1005) & (g2603)) + ((!sk[48]) & (!g165) & (g2585) & (g1005) & (!g2603)) + ((!sk[48]) & (!g165) & (g2585) & (g1005) & (g2603)) + ((!sk[48]) & (g165) & (!g2585) & (!g1005) & (g2603)) + ((!sk[48]) & (g165) & (!g2585) & (g1005) & (!g2603)) + ((!sk[48]) & (g165) & (!g2585) & (g1005) & (g2603)) + ((!sk[48]) & (g165) & (g2585) & (!g1005) & (!g2603)) + ((!sk[48]) & (g165) & (g2585) & (!g1005) & (g2603)) + ((!sk[48]) & (g165) & (g2585) & (g1005) & (!g2603)) + ((!sk[48]) & (g165) & (g2585) & (g1005) & (g2603)) + ((sk[48]) & (!g165) & (g2585) & (!g1005) & (!g2603)) + ((sk[48]) & (!g165) & (g2585) & (g1005) & (g2603)) + ((sk[48]) & (g165) & (g2585) & (!g1005) & (g2603)) + ((sk[48]) & (g165) & (g2585) & (g1005) & (!g2603)));
	assign g5042 = (((!g2921) & (!g3200) & (!sk[49]) & (g2605)) + ((!g2921) & (!g3200) & (sk[49]) & (g2605)) + ((!g2921) & (g3200) & (!sk[49]) & (!g2605)) + ((!g2921) & (g3200) & (!sk[49]) & (g2605)) + ((!g2921) & (g3200) & (sk[49]) & (g2605)) + ((g2921) & (!g3200) & (!sk[49]) & (g2605)) + ((g2921) & (g3200) & (!sk[49]) & (!g2605)) + ((g2921) & (g3200) & (!sk[49]) & (g2605)) + ((g2921) & (g3200) & (sk[49]) & (!g2605)) + ((g2921) & (g3200) & (sk[49]) & (g2605)));
	assign g2606 = (((!g1837) & (!g2033) & (!g2034) & (!sk[50]) & (g2605)) + ((!g1837) & (!g2033) & (!g2034) & (sk[50]) & (g2605)) + ((!g1837) & (!g2033) & (g2034) & (!sk[50]) & (!g2605)) + ((!g1837) & (!g2033) & (g2034) & (!sk[50]) & (g2605)) + ((!g1837) & (g2033) & (!g2034) & (!sk[50]) & (!g2605)) + ((!g1837) & (g2033) & (!g2034) & (!sk[50]) & (g2605)) + ((!g1837) & (g2033) & (g2034) & (!sk[50]) & (!g2605)) + ((!g1837) & (g2033) & (g2034) & (!sk[50]) & (g2605)) + ((g1837) & (!g2033) & (!g2034) & (!sk[50]) & (g2605)) + ((g1837) & (!g2033) & (!g2034) & (sk[50]) & (g2605)) + ((g1837) & (!g2033) & (g2034) & (!sk[50]) & (!g2605)) + ((g1837) & (!g2033) & (g2034) & (!sk[50]) & (g2605)) + ((g1837) & (!g2033) & (g2034) & (sk[50]) & (!g2605)) + ((g1837) & (!g2033) & (g2034) & (sk[50]) & (g2605)) + ((g1837) & (g2033) & (!g2034) & (!sk[50]) & (!g2605)) + ((g1837) & (g2033) & (!g2034) & (!sk[50]) & (g2605)) + ((g1837) & (g2033) & (g2034) & (!sk[50]) & (!g2605)) + ((g1837) & (g2033) & (g2034) & (!sk[50]) & (g2605)));
	assign g2607 = (((g2329) & (!g2029) & (g2408) & (!g2599) & (!g2604) & (g2606)) + ((g2329) & (!g2029) & (g2408) & (!g2599) & (g2604) & (!g2606)) + ((g2329) & (!g2029) & (g2408) & (!g2599) & (g2604) & (g2606)) + ((g2329) & (!g2029) & (g2408) & (g2599) & (!g2604) & (g2606)) + ((g2329) & (!g2029) & (g2408) & (g2599) & (g2604) & (!g2606)) + ((g2329) & (!g2029) & (g2408) & (g2599) & (g2604) & (g2606)) + ((g2329) & (g2029) & (g2408) & (g2599) & (!g2604) & (!g2606)) + ((g2329) & (g2029) & (g2408) & (g2599) & (!g2604) & (g2606)) + ((g2329) & (g2029) & (g2408) & (g2599) & (g2604) & (!g2606)) + ((g2329) & (g2029) & (g2408) & (g2599) & (g2604) & (g2606)));
	assign g2609 = (((!g2086) & (!g2608) & (!sk[52]) & (!g2085) & (g2590) & (!g2591)) + ((!g2086) & (!g2608) & (!sk[52]) & (!g2085) & (g2590) & (g2591)) + ((!g2086) & (!g2608) & (!sk[52]) & (g2085) & (!g2590) & (!g2591)) + ((!g2086) & (!g2608) & (!sk[52]) & (g2085) & (!g2590) & (g2591)) + ((!g2086) & (!g2608) & (!sk[52]) & (g2085) & (g2590) & (!g2591)) + ((!g2086) & (!g2608) & (!sk[52]) & (g2085) & (g2590) & (g2591)) + ((!g2086) & (!g2608) & (sk[52]) & (!g2085) & (g2590) & (g2591)) + ((!g2086) & (!g2608) & (sk[52]) & (g2085) & (!g2590) & (g2591)) + ((!g2086) & (!g2608) & (sk[52]) & (g2085) & (g2590) & (!g2591)) + ((!g2086) & (!g2608) & (sk[52]) & (g2085) & (g2590) & (g2591)) + ((!g2086) & (g2608) & (!sk[52]) & (!g2085) & (!g2590) & (!g2591)) + ((!g2086) & (g2608) & (!sk[52]) & (!g2085) & (!g2590) & (g2591)) + ((!g2086) & (g2608) & (!sk[52]) & (!g2085) & (g2590) & (!g2591)) + ((!g2086) & (g2608) & (!sk[52]) & (!g2085) & (g2590) & (g2591)) + ((!g2086) & (g2608) & (!sk[52]) & (g2085) & (!g2590) & (!g2591)) + ((!g2086) & (g2608) & (!sk[52]) & (g2085) & (!g2590) & (g2591)) + ((!g2086) & (g2608) & (!sk[52]) & (g2085) & (g2590) & (!g2591)) + ((!g2086) & (g2608) & (!sk[52]) & (g2085) & (g2590) & (g2591)) + ((!g2086) & (g2608) & (sk[52]) & (!g2085) & (!g2590) & (!g2591)) + ((!g2086) & (g2608) & (sk[52]) & (!g2085) & (!g2590) & (g2591)) + ((!g2086) & (g2608) & (sk[52]) & (!g2085) & (g2590) & (!g2591)) + ((!g2086) & (g2608) & (sk[52]) & (g2085) & (!g2590) & (!g2591)) + ((g2086) & (!g2608) & (!sk[52]) & (!g2085) & (g2590) & (!g2591)) + ((g2086) & (!g2608) & (!sk[52]) & (!g2085) & (g2590) & (g2591)) + ((g2086) & (!g2608) & (!sk[52]) & (g2085) & (!g2590) & (!g2591)) + ((g2086) & (!g2608) & (!sk[52]) & (g2085) & (!g2590) & (g2591)) + ((g2086) & (!g2608) & (!sk[52]) & (g2085) & (g2590) & (!g2591)) + ((g2086) & (!g2608) & (!sk[52]) & (g2085) & (g2590) & (g2591)) + ((g2086) & (!g2608) & (sk[52]) & (!g2085) & (!g2590) & (!g2591)) + ((g2086) & (!g2608) & (sk[52]) & (!g2085) & (!g2590) & (g2591)) + ((g2086) & (!g2608) & (sk[52]) & (!g2085) & (g2590) & (!g2591)) + ((g2086) & (!g2608) & (sk[52]) & (g2085) & (!g2590) & (!g2591)) + ((g2086) & (g2608) & (!sk[52]) & (!g2085) & (!g2590) & (!g2591)) + ((g2086) & (g2608) & (!sk[52]) & (!g2085) & (!g2590) & (g2591)) + ((g2086) & (g2608) & (!sk[52]) & (!g2085) & (g2590) & (!g2591)) + ((g2086) & (g2608) & (!sk[52]) & (!g2085) & (g2590) & (g2591)) + ((g2086) & (g2608) & (!sk[52]) & (g2085) & (!g2590) & (!g2591)) + ((g2086) & (g2608) & (!sk[52]) & (g2085) & (!g2590) & (g2591)) + ((g2086) & (g2608) & (!sk[52]) & (g2085) & (g2590) & (!g2591)) + ((g2086) & (g2608) & (!sk[52]) & (g2085) & (g2590) & (g2591)) + ((g2086) & (g2608) & (sk[52]) & (!g2085) & (g2590) & (g2591)) + ((g2086) & (g2608) & (sk[52]) & (g2085) & (!g2590) & (g2591)) + ((g2086) & (g2608) & (sk[52]) & (g2085) & (g2590) & (!g2591)) + ((g2086) & (g2608) & (sk[52]) & (g2085) & (g2590) & (g2591)));
	assign g2610 = (((g2554) & (g2555) & (g2571) & (!g2085) & (!g2590) & (g2591)) + ((g2554) & (g2555) & (g2571) & (!g2085) & (g2590) & (!g2591)) + ((g2554) & (g2555) & (g2571) & (g2085) & (!g2590) & (!g2591)) + ((g2554) & (g2555) & (g2571) & (g2085) & (g2590) & (g2591)));
	assign g2611 = (((!g2573) & (!g2574) & (!g2576) & (!g2577) & (!g2592) & (!g2593)) + ((!g2573) & (!g2574) & (!g2576) & (!g2577) & (!g2592) & (g2593)) + ((!g2573) & (!g2574) & (!g2576) & (!g2577) & (g2592) & (!g2593)) + ((!g2573) & (!g2574) & (!g2576) & (g2577) & (!g2592) & (!g2593)) + ((!g2573) & (!g2574) & (!g2576) & (g2577) & (!g2592) & (g2593)) + ((!g2573) & (!g2574) & (!g2576) & (g2577) & (g2592) & (!g2593)) + ((!g2573) & (!g2574) & (g2576) & (!g2577) & (!g2592) & (!g2593)) + ((!g2573) & (!g2574) & (g2576) & (!g2577) & (!g2592) & (g2593)) + ((!g2573) & (!g2574) & (g2576) & (!g2577) & (g2592) & (!g2593)) + ((!g2573) & (!g2574) & (g2576) & (g2577) & (!g2592) & (!g2593)) + ((!g2573) & (g2574) & (!g2576) & (!g2577) & (!g2592) & (!g2593)) + ((!g2573) & (g2574) & (!g2576) & (!g2577) & (!g2592) & (g2593)) + ((!g2573) & (g2574) & (!g2576) & (!g2577) & (g2592) & (!g2593)) + ((!g2573) & (g2574) & (!g2576) & (g2577) & (!g2592) & (!g2593)) + ((!g2573) & (g2574) & (g2576) & (!g2577) & (!g2592) & (!g2593)) + ((!g2573) & (g2574) & (g2576) & (g2577) & (!g2592) & (!g2593)) + ((g2573) & (!g2574) & (!g2576) & (!g2577) & (!g2592) & (!g2593)) + ((g2573) & (!g2574) & (!g2576) & (!g2577) & (!g2592) & (g2593)) + ((g2573) & (!g2574) & (!g2576) & (!g2577) & (g2592) & (!g2593)) + ((g2573) & (!g2574) & (!g2576) & (g2577) & (!g2592) & (!g2593)) + ((g2573) & (!g2574) & (g2576) & (!g2577) & (!g2592) & (!g2593)) + ((g2573) & (!g2574) & (g2576) & (g2577) & (!g2592) & (!g2593)) + ((g2573) & (g2574) & (!g2576) & (!g2577) & (!g2592) & (!g2593)) + ((g2573) & (g2574) & (!g2576) & (!g2577) & (!g2592) & (g2593)) + ((g2573) & (g2574) & (!g2576) & (!g2577) & (g2592) & (!g2593)) + ((g2573) & (g2574) & (!g2576) & (g2577) & (!g2592) & (!g2593)) + ((g2573) & (g2574) & (g2576) & (!g2577) & (!g2592) & (!g2593)) + ((g2573) & (g2574) & (g2576) & (g2577) & (!g2592) & (!g2593)));
	assign g2612 = (((!g2590) & (sk[55]) & (g2085)) + ((g2590) & (!sk[55]) & (!g2085)) + ((g2590) & (!sk[55]) & (g2085)));
	assign g2613 = (((!g2608) & (sk[56]) & (!g2086)) + ((g2608) & (!sk[56]) & (!g2086)) + ((g2608) & (!sk[56]) & (g2086)) + ((g2608) & (sk[56]) & (g2086)));
	assign g2614 = (((!g2611) & (!sk[57]) & (!g2612) & (g2613)) + ((!g2611) & (!sk[57]) & (g2612) & (!g2613)) + ((!g2611) & (!sk[57]) & (g2612) & (g2613)) + ((!g2611) & (sk[57]) & (!g2612) & (!g2613)) + ((!g2611) & (sk[57]) & (g2612) & (g2613)) + ((g2611) & (!sk[57]) & (!g2612) & (g2613)) + ((g2611) & (!sk[57]) & (g2612) & (!g2613)) + ((g2611) & (!sk[57]) & (g2612) & (g2613)) + ((g2611) & (sk[57]) & (!g2612) & (g2613)) + ((g2611) & (sk[57]) & (g2612) & (!g2613)));
	assign g2615 = (((!g2086) & (!g2085) & (!g2084) & (g2083) & (g2071) & (g2074)) + ((!g2086) & (!g2085) & (g2084) & (!g2083) & (!g2071) & (g2074)) + ((!g2086) & (!g2085) & (g2084) & (g2083) & (!g2071) & (g2074)) + ((!g2086) & (!g2085) & (g2084) & (g2083) & (g2071) & (g2074)) + ((!g2086) & (g2085) & (!g2084) & (!g2083) & (g2071) & (!g2074)) + ((!g2086) & (g2085) & (!g2084) & (g2083) & (g2071) & (!g2074)) + ((!g2086) & (g2085) & (!g2084) & (g2083) & (g2071) & (g2074)) + ((!g2086) & (g2085) & (g2084) & (!g2083) & (!g2071) & (g2074)) + ((!g2086) & (g2085) & (g2084) & (!g2083) & (g2071) & (!g2074)) + ((!g2086) & (g2085) & (g2084) & (g2083) & (!g2071) & (g2074)) + ((!g2086) & (g2085) & (g2084) & (g2083) & (g2071) & (!g2074)) + ((!g2086) & (g2085) & (g2084) & (g2083) & (g2071) & (g2074)) + ((g2086) & (!g2085) & (!g2084) & (!g2083) & (!g2071) & (!g2074)) + ((g2086) & (!g2085) & (!g2084) & (g2083) & (!g2071) & (!g2074)) + ((g2086) & (!g2085) & (!g2084) & (g2083) & (g2071) & (g2074)) + ((g2086) & (!g2085) & (g2084) & (!g2083) & (!g2071) & (!g2074)) + ((g2086) & (!g2085) & (g2084) & (!g2083) & (!g2071) & (g2074)) + ((g2086) & (!g2085) & (g2084) & (g2083) & (!g2071) & (!g2074)) + ((g2086) & (!g2085) & (g2084) & (g2083) & (!g2071) & (g2074)) + ((g2086) & (!g2085) & (g2084) & (g2083) & (g2071) & (g2074)) + ((g2086) & (g2085) & (!g2084) & (!g2083) & (!g2071) & (!g2074)) + ((g2086) & (g2085) & (!g2084) & (!g2083) & (g2071) & (!g2074)) + ((g2086) & (g2085) & (!g2084) & (g2083) & (!g2071) & (!g2074)) + ((g2086) & (g2085) & (!g2084) & (g2083) & (g2071) & (!g2074)) + ((g2086) & (g2085) & (!g2084) & (g2083) & (g2071) & (g2074)) + ((g2086) & (g2085) & (g2084) & (!g2083) & (!g2071) & (!g2074)) + ((g2086) & (g2085) & (g2084) & (!g2083) & (!g2071) & (g2074)) + ((g2086) & (g2085) & (g2084) & (!g2083) & (g2071) & (!g2074)) + ((g2086) & (g2085) & (g2084) & (g2083) & (!g2071) & (!g2074)) + ((g2086) & (g2085) & (g2084) & (g2083) & (!g2071) & (g2074)) + ((g2086) & (g2085) & (g2084) & (g2083) & (g2071) & (!g2074)) + ((g2086) & (g2085) & (g2084) & (g2083) & (g2071) & (g2074)));
	assign g2616 = (((!g2615) & (!g2449) & (!g2536) & (g2350) & (g2076) & (g2077)) + ((!g2615) & (!g2449) & (g2536) & (!g2350) & (!g2076) & (g2077)) + ((!g2615) & (!g2449) & (g2536) & (g2350) & (!g2076) & (g2077)) + ((!g2615) & (!g2449) & (g2536) & (g2350) & (g2076) & (g2077)) + ((!g2615) & (g2449) & (!g2536) & (!g2350) & (g2076) & (!g2077)) + ((!g2615) & (g2449) & (!g2536) & (g2350) & (g2076) & (!g2077)) + ((!g2615) & (g2449) & (!g2536) & (g2350) & (g2076) & (g2077)) + ((!g2615) & (g2449) & (g2536) & (!g2350) & (!g2076) & (g2077)) + ((!g2615) & (g2449) & (g2536) & (!g2350) & (g2076) & (!g2077)) + ((!g2615) & (g2449) & (g2536) & (g2350) & (!g2076) & (g2077)) + ((!g2615) & (g2449) & (g2536) & (g2350) & (g2076) & (!g2077)) + ((!g2615) & (g2449) & (g2536) & (g2350) & (g2076) & (g2077)) + ((g2615) & (!g2449) & (!g2536) & (!g2350) & (!g2076) & (!g2077)) + ((g2615) & (!g2449) & (!g2536) & (g2350) & (!g2076) & (!g2077)) + ((g2615) & (!g2449) & (!g2536) & (g2350) & (g2076) & (g2077)) + ((g2615) & (!g2449) & (g2536) & (!g2350) & (!g2076) & (!g2077)) + ((g2615) & (!g2449) & (g2536) & (!g2350) & (!g2076) & (g2077)) + ((g2615) & (!g2449) & (g2536) & (g2350) & (!g2076) & (!g2077)) + ((g2615) & (!g2449) & (g2536) & (g2350) & (!g2076) & (g2077)) + ((g2615) & (!g2449) & (g2536) & (g2350) & (g2076) & (g2077)) + ((g2615) & (g2449) & (!g2536) & (!g2350) & (!g2076) & (!g2077)) + ((g2615) & (g2449) & (!g2536) & (!g2350) & (g2076) & (!g2077)) + ((g2615) & (g2449) & (!g2536) & (g2350) & (!g2076) & (!g2077)) + ((g2615) & (g2449) & (!g2536) & (g2350) & (g2076) & (!g2077)) + ((g2615) & (g2449) & (!g2536) & (g2350) & (g2076) & (g2077)) + ((g2615) & (g2449) & (g2536) & (!g2350) & (!g2076) & (!g2077)) + ((g2615) & (g2449) & (g2536) & (!g2350) & (!g2076) & (g2077)) + ((g2615) & (g2449) & (g2536) & (!g2350) & (g2076) & (!g2077)) + ((g2615) & (g2449) & (g2536) & (g2350) & (!g2076) & (!g2077)) + ((g2615) & (g2449) & (g2536) & (g2350) & (!g2076) & (g2077)) + ((g2615) & (g2449) & (g2536) & (g2350) & (g2076) & (!g2077)) + ((g2615) & (g2449) & (g2536) & (g2350) & (g2076) & (g2077)));
	assign g2617 = (((!g2616) & (!g2237) & (!g2246) & (g2191) & (g2073) & (g2125)) + ((!g2616) & (!g2237) & (g2246) & (!g2191) & (!g2073) & (g2125)) + ((!g2616) & (!g2237) & (g2246) & (g2191) & (!g2073) & (g2125)) + ((!g2616) & (!g2237) & (g2246) & (g2191) & (g2073) & (g2125)) + ((!g2616) & (g2237) & (!g2246) & (!g2191) & (g2073) & (!g2125)) + ((!g2616) & (g2237) & (!g2246) & (g2191) & (g2073) & (!g2125)) + ((!g2616) & (g2237) & (!g2246) & (g2191) & (g2073) & (g2125)) + ((!g2616) & (g2237) & (g2246) & (!g2191) & (!g2073) & (g2125)) + ((!g2616) & (g2237) & (g2246) & (!g2191) & (g2073) & (!g2125)) + ((!g2616) & (g2237) & (g2246) & (g2191) & (!g2073) & (g2125)) + ((!g2616) & (g2237) & (g2246) & (g2191) & (g2073) & (!g2125)) + ((!g2616) & (g2237) & (g2246) & (g2191) & (g2073) & (g2125)) + ((g2616) & (!g2237) & (!g2246) & (!g2191) & (!g2073) & (!g2125)) + ((g2616) & (!g2237) & (!g2246) & (g2191) & (!g2073) & (!g2125)) + ((g2616) & (!g2237) & (!g2246) & (g2191) & (g2073) & (g2125)) + ((g2616) & (!g2237) & (g2246) & (!g2191) & (!g2073) & (!g2125)) + ((g2616) & (!g2237) & (g2246) & (!g2191) & (!g2073) & (g2125)) + ((g2616) & (!g2237) & (g2246) & (g2191) & (!g2073) & (!g2125)) + ((g2616) & (!g2237) & (g2246) & (g2191) & (!g2073) & (g2125)) + ((g2616) & (!g2237) & (g2246) & (g2191) & (g2073) & (g2125)) + ((g2616) & (g2237) & (!g2246) & (!g2191) & (!g2073) & (!g2125)) + ((g2616) & (g2237) & (!g2246) & (!g2191) & (g2073) & (!g2125)) + ((g2616) & (g2237) & (!g2246) & (g2191) & (!g2073) & (!g2125)) + ((g2616) & (g2237) & (!g2246) & (g2191) & (g2073) & (!g2125)) + ((g2616) & (g2237) & (!g2246) & (g2191) & (g2073) & (g2125)) + ((g2616) & (g2237) & (g2246) & (!g2191) & (!g2073) & (!g2125)) + ((g2616) & (g2237) & (g2246) & (!g2191) & (!g2073) & (g2125)) + ((g2616) & (g2237) & (g2246) & (!g2191) & (g2073) & (!g2125)) + ((g2616) & (g2237) & (g2246) & (g2191) & (!g2073) & (!g2125)) + ((g2616) & (g2237) & (g2246) & (g2191) & (!g2073) & (g2125)) + ((g2616) & (g2237) & (g2246) & (g2191) & (g2073) & (!g2125)) + ((g2616) & (g2237) & (g2246) & (g2191) & (g2073) & (g2125)));
	assign g2618 = (((!g2086) & (!g2608) & (!g2124) & (!g2264) & (!g3479) & (g2617)) + ((!g2086) & (!g2608) & (!g2124) & (!g2264) & (g3479) & (g2617)) + ((!g2086) & (!g2608) & (!g2124) & (g2264) & (g3479) & (!g2617)) + ((!g2086) & (!g2608) & (!g2124) & (g2264) & (g3479) & (g2617)) + ((!g2086) & (g2608) & (!g2124) & (!g2264) & (!g3479) & (g2617)) + ((!g2086) & (g2608) & (!g2124) & (!g2264) & (g3479) & (g2617)) + ((!g2086) & (g2608) & (!g2124) & (g2264) & (g3479) & (!g2617)) + ((!g2086) & (g2608) & (!g2124) & (g2264) & (g3479) & (g2617)) + ((!g2086) & (g2608) & (g2124) & (!g2264) & (!g3479) & (!g2617)) + ((!g2086) & (g2608) & (g2124) & (!g2264) & (!g3479) & (g2617)) + ((!g2086) & (g2608) & (g2124) & (!g2264) & (g3479) & (!g2617)) + ((!g2086) & (g2608) & (g2124) & (!g2264) & (g3479) & (g2617)) + ((!g2086) & (g2608) & (g2124) & (g2264) & (!g3479) & (!g2617)) + ((!g2086) & (g2608) & (g2124) & (g2264) & (!g3479) & (g2617)) + ((!g2086) & (g2608) & (g2124) & (g2264) & (g3479) & (!g2617)) + ((!g2086) & (g2608) & (g2124) & (g2264) & (g3479) & (g2617)) + ((g2086) & (!g2608) & (!g2124) & (!g2264) & (!g3479) & (g2617)) + ((g2086) & (!g2608) & (!g2124) & (!g2264) & (g3479) & (g2617)) + ((g2086) & (!g2608) & (!g2124) & (g2264) & (g3479) & (!g2617)) + ((g2086) & (!g2608) & (!g2124) & (g2264) & (g3479) & (g2617)) + ((g2086) & (!g2608) & (g2124) & (!g2264) & (!g3479) & (!g2617)) + ((g2086) & (!g2608) & (g2124) & (!g2264) & (!g3479) & (g2617)) + ((g2086) & (!g2608) & (g2124) & (!g2264) & (g3479) & (!g2617)) + ((g2086) & (!g2608) & (g2124) & (!g2264) & (g3479) & (g2617)) + ((g2086) & (!g2608) & (g2124) & (g2264) & (!g3479) & (!g2617)) + ((g2086) & (!g2608) & (g2124) & (g2264) & (!g3479) & (g2617)) + ((g2086) & (!g2608) & (g2124) & (g2264) & (g3479) & (!g2617)) + ((g2086) & (!g2608) & (g2124) & (g2264) & (g3479) & (g2617)) + ((g2086) & (g2608) & (!g2124) & (!g2264) & (!g3479) & (g2617)) + ((g2086) & (g2608) & (!g2124) & (!g2264) & (g3479) & (g2617)) + ((g2086) & (g2608) & (!g2124) & (g2264) & (g3479) & (!g2617)) + ((g2086) & (g2608) & (!g2124) & (g2264) & (g3479) & (g2617)) + ((g2086) & (g2608) & (g2124) & (!g2264) & (!g3479) & (!g2617)) + ((g2086) & (g2608) & (g2124) & (!g2264) & (!g3479) & (g2617)) + ((g2086) & (g2608) & (g2124) & (!g2264) & (g3479) & (!g2617)) + ((g2086) & (g2608) & (g2124) & (!g2264) & (g3479) & (g2617)));
	assign g2619 = (((!g912) & (!sk[62]) & (!g2563) & (!g960) & (g1005)) + ((!g912) & (!sk[62]) & (!g2563) & (g960) & (!g1005)) + ((!g912) & (!sk[62]) & (!g2563) & (g960) & (g1005)) + ((!g912) & (!sk[62]) & (g2563) & (!g960) & (!g1005)) + ((!g912) & (!sk[62]) & (g2563) & (!g960) & (g1005)) + ((!g912) & (!sk[62]) & (g2563) & (g960) & (!g1005)) + ((!g912) & (!sk[62]) & (g2563) & (g960) & (g1005)) + ((g912) & (!sk[62]) & (!g2563) & (!g960) & (g1005)) + ((g912) & (!sk[62]) & (!g2563) & (g960) & (!g1005)) + ((g912) & (!sk[62]) & (!g2563) & (g960) & (g1005)) + ((g912) & (!sk[62]) & (g2563) & (!g960) & (!g1005)) + ((g912) & (!sk[62]) & (g2563) & (!g960) & (g1005)) + ((g912) & (!sk[62]) & (g2563) & (g960) & (!g1005)) + ((g912) & (!sk[62]) & (g2563) & (g960) & (g1005)) + ((g912) & (sk[62]) & (g2563) & (g960) & (g1005)));
	assign g2620 = (((!g1050) & (sk[63]) & (g2619)) + ((g1050) & (!sk[63]) & (!g2619)) + ((g1050) & (!sk[63]) & (g2619)) + ((g1050) & (sk[63]) & (!g2619)));
	assign g2621 = (((!g165) & (!sk[64]) & (!g166) & (!g1005) & (g2603) & (!g1050)) + ((!g165) & (!sk[64]) & (!g166) & (!g1005) & (g2603) & (g1050)) + ((!g165) & (!sk[64]) & (!g166) & (g1005) & (!g2603) & (!g1050)) + ((!g165) & (!sk[64]) & (!g166) & (g1005) & (!g2603) & (g1050)) + ((!g165) & (!sk[64]) & (!g166) & (g1005) & (g2603) & (!g1050)) + ((!g165) & (!sk[64]) & (!g166) & (g1005) & (g2603) & (g1050)) + ((!g165) & (!sk[64]) & (g166) & (!g1005) & (!g2603) & (!g1050)) + ((!g165) & (!sk[64]) & (g166) & (!g1005) & (!g2603) & (g1050)) + ((!g165) & (!sk[64]) & (g166) & (!g1005) & (g2603) & (!g1050)) + ((!g165) & (!sk[64]) & (g166) & (!g1005) & (g2603) & (g1050)) + ((!g165) & (!sk[64]) & (g166) & (g1005) & (!g2603) & (!g1050)) + ((!g165) & (!sk[64]) & (g166) & (g1005) & (!g2603) & (g1050)) + ((!g165) & (!sk[64]) & (g166) & (g1005) & (g2603) & (!g1050)) + ((!g165) & (!sk[64]) & (g166) & (g1005) & (g2603) & (g1050)) + ((!g165) & (sk[64]) & (!g166) & (!g1005) & (!g2603) & (g1050)) + ((!g165) & (sk[64]) & (!g166) & (!g1005) & (g2603) & (g1050)) + ((!g165) & (sk[64]) & (!g166) & (g1005) & (!g2603) & (!g1050)) + ((!g165) & (sk[64]) & (!g166) & (g1005) & (g2603) & (g1050)) + ((!g165) & (sk[64]) & (g166) & (!g1005) & (!g2603) & (!g1050)) + ((!g165) & (sk[64]) & (g166) & (!g1005) & (g2603) & (!g1050)) + ((!g165) & (sk[64]) & (g166) & (g1005) & (!g2603) & (g1050)) + ((!g165) & (sk[64]) & (g166) & (g1005) & (g2603) & (!g1050)) + ((g165) & (!sk[64]) & (!g166) & (!g1005) & (g2603) & (!g1050)) + ((g165) & (!sk[64]) & (!g166) & (!g1005) & (g2603) & (g1050)) + ((g165) & (!sk[64]) & (!g166) & (g1005) & (!g2603) & (!g1050)) + ((g165) & (!sk[64]) & (!g166) & (g1005) & (!g2603) & (g1050)) + ((g165) & (!sk[64]) & (!g166) & (g1005) & (g2603) & (!g1050)) + ((g165) & (!sk[64]) & (!g166) & (g1005) & (g2603) & (g1050)) + ((g165) & (!sk[64]) & (g166) & (!g1005) & (!g2603) & (!g1050)) + ((g165) & (!sk[64]) & (g166) & (!g1005) & (!g2603) & (g1050)) + ((g165) & (!sk[64]) & (g166) & (!g1005) & (g2603) & (!g1050)) + ((g165) & (!sk[64]) & (g166) & (!g1005) & (g2603) & (g1050)) + ((g165) & (!sk[64]) & (g166) & (g1005) & (!g2603) & (!g1050)) + ((g165) & (!sk[64]) & (g166) & (g1005) & (!g2603) & (g1050)) + ((g165) & (!sk[64]) & (g166) & (g1005) & (g2603) & (!g1050)) + ((g165) & (!sk[64]) & (g166) & (g1005) & (g2603) & (g1050)) + ((g165) & (sk[64]) & (!g166) & (!g1005) & (!g2603) & (!g1050)) + ((g165) & (sk[64]) & (!g166) & (!g1005) & (g2603) & (g1050)) + ((g165) & (sk[64]) & (!g166) & (g1005) & (!g2603) & (!g1050)) + ((g165) & (sk[64]) & (!g166) & (g1005) & (g2603) & (!g1050)) + ((g165) & (sk[64]) & (g166) & (!g1005) & (!g2603) & (g1050)) + ((g165) & (sk[64]) & (g166) & (!g1005) & (g2603) & (!g1050)) + ((g165) & (sk[64]) & (g166) & (g1005) & (!g2603) & (g1050)) + ((g165) & (sk[64]) & (g166) & (g1005) & (g2603) & (g1050)));
	assign g5043 = (((!sk[65]) & (!g2921) & (!g3091) & (g2622)) + ((!sk[65]) & (!g2921) & (g3091) & (!g2622)) + ((!sk[65]) & (!g2921) & (g3091) & (g2622)) + ((!sk[65]) & (g2921) & (!g3091) & (g2622)) + ((!sk[65]) & (g2921) & (g3091) & (!g2622)) + ((!sk[65]) & (g2921) & (g3091) & (g2622)) + ((sk[65]) & (!g2921) & (!g3091) & (g2622)) + ((sk[65]) & (!g2921) & (g3091) & (g2622)) + ((sk[65]) & (g2921) & (g3091) & (!g2622)) + ((sk[65]) & (g2921) & (g3091) & (g2622)));
	assign g2623 = (((!g1850) & (!g2033) & (!g2034) & (!sk[66]) & (g2621) & (!g2622)) + ((!g1850) & (!g2033) & (!g2034) & (!sk[66]) & (g2621) & (g2622)) + ((!g1850) & (!g2033) & (!g2034) & (sk[66]) & (!g2621) & (g2622)) + ((!g1850) & (!g2033) & (!g2034) & (sk[66]) & (g2621) & (g2622)) + ((!g1850) & (!g2033) & (g2034) & (!sk[66]) & (!g2621) & (!g2622)) + ((!g1850) & (!g2033) & (g2034) & (!sk[66]) & (!g2621) & (g2622)) + ((!g1850) & (!g2033) & (g2034) & (!sk[66]) & (g2621) & (!g2622)) + ((!g1850) & (!g2033) & (g2034) & (!sk[66]) & (g2621) & (g2622)) + ((!g1850) & (g2033) & (!g2034) & (!sk[66]) & (!g2621) & (!g2622)) + ((!g1850) & (g2033) & (!g2034) & (!sk[66]) & (!g2621) & (g2622)) + ((!g1850) & (g2033) & (!g2034) & (!sk[66]) & (g2621) & (!g2622)) + ((!g1850) & (g2033) & (!g2034) & (!sk[66]) & (g2621) & (g2622)) + ((!g1850) & (g2033) & (!g2034) & (sk[66]) & (g2621) & (!g2622)) + ((!g1850) & (g2033) & (!g2034) & (sk[66]) & (g2621) & (g2622)) + ((!g1850) & (g2033) & (g2034) & (!sk[66]) & (!g2621) & (!g2622)) + ((!g1850) & (g2033) & (g2034) & (!sk[66]) & (!g2621) & (g2622)) + ((!g1850) & (g2033) & (g2034) & (!sk[66]) & (g2621) & (!g2622)) + ((!g1850) & (g2033) & (g2034) & (!sk[66]) & (g2621) & (g2622)) + ((g1850) & (!g2033) & (!g2034) & (!sk[66]) & (g2621) & (!g2622)) + ((g1850) & (!g2033) & (!g2034) & (!sk[66]) & (g2621) & (g2622)) + ((g1850) & (!g2033) & (!g2034) & (sk[66]) & (!g2621) & (g2622)) + ((g1850) & (!g2033) & (!g2034) & (sk[66]) & (g2621) & (g2622)) + ((g1850) & (!g2033) & (g2034) & (!sk[66]) & (!g2621) & (!g2622)) + ((g1850) & (!g2033) & (g2034) & (!sk[66]) & (!g2621) & (g2622)) + ((g1850) & (!g2033) & (g2034) & (!sk[66]) & (g2621) & (!g2622)) + ((g1850) & (!g2033) & (g2034) & (!sk[66]) & (g2621) & (g2622)) + ((g1850) & (!g2033) & (g2034) & (sk[66]) & (!g2621) & (!g2622)) + ((g1850) & (!g2033) & (g2034) & (sk[66]) & (!g2621) & (g2622)) + ((g1850) & (!g2033) & (g2034) & (sk[66]) & (g2621) & (!g2622)) + ((g1850) & (!g2033) & (g2034) & (sk[66]) & (g2621) & (g2622)) + ((g1850) & (g2033) & (!g2034) & (!sk[66]) & (!g2621) & (!g2622)) + ((g1850) & (g2033) & (!g2034) & (!sk[66]) & (!g2621) & (g2622)) + ((g1850) & (g2033) & (!g2034) & (!sk[66]) & (g2621) & (!g2622)) + ((g1850) & (g2033) & (!g2034) & (!sk[66]) & (g2621) & (g2622)) + ((g1850) & (g2033) & (!g2034) & (sk[66]) & (g2621) & (!g2622)) + ((g1850) & (g2033) & (!g2034) & (sk[66]) & (g2621) & (g2622)) + ((g1850) & (g2033) & (g2034) & (!sk[66]) & (!g2621) & (!g2622)) + ((g1850) & (g2033) & (g2034) & (!sk[66]) & (!g2621) & (g2622)) + ((g1850) & (g2033) & (g2034) & (!sk[66]) & (g2621) & (!g2622)) + ((g1850) & (g2033) & (g2034) & (!sk[66]) & (g2621) & (g2622)));
	assign g2624 = (((!sk[67]) & (!g2329) & (!g2029) & (!g2408) & (g2620) & (!g2623)) + ((!sk[67]) & (!g2329) & (!g2029) & (!g2408) & (g2620) & (g2623)) + ((!sk[67]) & (!g2329) & (!g2029) & (g2408) & (g2620) & (!g2623)) + ((!sk[67]) & (!g2329) & (!g2029) & (g2408) & (g2620) & (g2623)) + ((!sk[67]) & (!g2329) & (g2029) & (!g2408) & (!g2620) & (!g2623)) + ((!sk[67]) & (!g2329) & (g2029) & (!g2408) & (!g2620) & (g2623)) + ((!sk[67]) & (!g2329) & (g2029) & (!g2408) & (g2620) & (!g2623)) + ((!sk[67]) & (!g2329) & (g2029) & (!g2408) & (g2620) & (g2623)) + ((!sk[67]) & (!g2329) & (g2029) & (g2408) & (!g2620) & (!g2623)) + ((!sk[67]) & (!g2329) & (g2029) & (g2408) & (!g2620) & (g2623)) + ((!sk[67]) & (!g2329) & (g2029) & (g2408) & (g2620) & (!g2623)) + ((!sk[67]) & (!g2329) & (g2029) & (g2408) & (g2620) & (g2623)) + ((!sk[67]) & (g2329) & (!g2029) & (!g2408) & (g2620) & (!g2623)) + ((!sk[67]) & (g2329) & (!g2029) & (!g2408) & (g2620) & (g2623)) + ((!sk[67]) & (g2329) & (!g2029) & (g2408) & (g2620) & (!g2623)) + ((!sk[67]) & (g2329) & (!g2029) & (g2408) & (g2620) & (g2623)) + ((!sk[67]) & (g2329) & (g2029) & (!g2408) & (!g2620) & (!g2623)) + ((!sk[67]) & (g2329) & (g2029) & (!g2408) & (!g2620) & (g2623)) + ((!sk[67]) & (g2329) & (g2029) & (!g2408) & (g2620) & (!g2623)) + ((!sk[67]) & (g2329) & (g2029) & (!g2408) & (g2620) & (g2623)) + ((!sk[67]) & (g2329) & (g2029) & (g2408) & (!g2620) & (!g2623)) + ((!sk[67]) & (g2329) & (g2029) & (g2408) & (!g2620) & (g2623)) + ((!sk[67]) & (g2329) & (g2029) & (g2408) & (g2620) & (!g2623)) + ((!sk[67]) & (g2329) & (g2029) & (g2408) & (g2620) & (g2623)) + ((sk[67]) & (g2329) & (!g2029) & (g2408) & (!g2620) & (g2623)) + ((sk[67]) & (g2329) & (!g2029) & (g2408) & (g2620) & (g2623)) + ((sk[67]) & (g2329) & (g2029) & (g2408) & (g2620) & (!g2623)) + ((sk[67]) & (g2329) & (g2029) & (g2408) & (g2620) & (g2623)));
	assign g2626 = (((!g2086) & (!g2608) & (!g2085) & (!g2590) & (!g2591) & (!g3127)) + ((!g2086) & (!g2608) & (!g2085) & (!g2590) & (g2591) & (!g3127)) + ((!g2086) & (!g2608) & (!g2085) & (g2590) & (!g2591) & (!g3127)) + ((!g2086) & (!g2608) & (!g2085) & (g2590) & (g2591) & (!g3127)) + ((!g2086) & (!g2608) & (g2085) & (!g2590) & (!g2591) & (!g3127)) + ((!g2086) & (!g2608) & (g2085) & (!g2590) & (g2591) & (!g3127)) + ((!g2086) & (!g2608) & (g2085) & (g2590) & (!g2591) & (!g3127)) + ((!g2086) & (!g2608) & (g2085) & (g2590) & (g2591) & (!g3127)) + ((!g2086) & (g2608) & (!g2085) & (!g2590) & (!g2591) & (!g3127)) + ((!g2086) & (g2608) & (!g2085) & (!g2590) & (g2591) & (!g3127)) + ((!g2086) & (g2608) & (!g2085) & (g2590) & (!g2591) & (!g3127)) + ((!g2086) & (g2608) & (!g2085) & (g2590) & (g2591) & (g3127)) + ((!g2086) & (g2608) & (g2085) & (!g2590) & (!g2591) & (!g3127)) + ((!g2086) & (g2608) & (g2085) & (!g2590) & (g2591) & (g3127)) + ((!g2086) & (g2608) & (g2085) & (g2590) & (!g2591) & (g3127)) + ((!g2086) & (g2608) & (g2085) & (g2590) & (g2591) & (g3127)) + ((g2086) & (!g2608) & (!g2085) & (!g2590) & (!g2591) & (!g3127)) + ((g2086) & (!g2608) & (!g2085) & (!g2590) & (g2591) & (!g3127)) + ((g2086) & (!g2608) & (!g2085) & (g2590) & (!g2591) & (!g3127)) + ((g2086) & (!g2608) & (!g2085) & (g2590) & (g2591) & (g3127)) + ((g2086) & (!g2608) & (g2085) & (!g2590) & (!g2591) & (!g3127)) + ((g2086) & (!g2608) & (g2085) & (!g2590) & (g2591) & (g3127)) + ((g2086) & (!g2608) & (g2085) & (g2590) & (!g2591) & (g3127)) + ((g2086) & (!g2608) & (g2085) & (g2590) & (g2591) & (g3127)) + ((g2086) & (g2608) & (!g2085) & (!g2590) & (!g2591) & (g3127)) + ((g2086) & (g2608) & (!g2085) & (!g2590) & (g2591) & (g3127)) + ((g2086) & (g2608) & (!g2085) & (g2590) & (!g2591) & (g3127)) + ((g2086) & (g2608) & (!g2085) & (g2590) & (g2591) & (g3127)) + ((g2086) & (g2608) & (g2085) & (!g2590) & (!g2591) & (g3127)) + ((g2086) & (g2608) & (g2085) & (!g2590) & (g2591) & (g3127)) + ((g2086) & (g2608) & (g2085) & (g2590) & (!g2591) & (g3127)) + ((g2086) & (g2608) & (g2085) & (g2590) & (g2591) & (g3127)));
	assign g2627 = (((!g2611) & (!sk[69]) & (g2612) & (!g2613)) + ((!g2611) & (!sk[69]) & (g2612) & (g2613)) + ((!g2611) & (sk[69]) & (!g2612) & (g2613)) + ((!g2611) & (sk[69]) & (g2612) & (!g2613)) + ((!g2611) & (sk[69]) & (g2612) & (g2613)) + ((g2611) & (!sk[69]) & (g2612) & (!g2613)) + ((g2611) & (!sk[69]) & (g2612) & (g2613)) + ((g2611) & (sk[69]) & (g2612) & (g2613)));
	assign g2628 = (((!sk[70]) & (!g2608) & (g2086)) + ((!sk[70]) & (g2608) & (g2086)) + ((sk[70]) & (!g2608) & (g2086)));
	assign g2629 = (((!sk[71]) & (!g2625) & (g2093)) + ((!sk[71]) & (g2625) & (g2093)) + ((sk[71]) & (!g2625) & (!g2093)) + ((sk[71]) & (g2625) & (g2093)));
	assign g2630 = (((!g2627) & (!g2628) & (sk[72]) & (g2629)) + ((!g2627) & (g2628) & (!sk[72]) & (!g2629)) + ((!g2627) & (g2628) & (!sk[72]) & (g2629)) + ((!g2627) & (g2628) & (sk[72]) & (!g2629)) + ((g2627) & (!g2628) & (sk[72]) & (!g2629)) + ((g2627) & (g2628) & (!sk[72]) & (!g2629)) + ((g2627) & (g2628) & (!sk[72]) & (g2629)) + ((g2627) & (g2628) & (sk[72]) & (g2629)));
	assign g2631 = (((!sk[73]) & (!g2093) & (g2625)) + ((!sk[73]) & (g2093) & (g2625)) + ((sk[73]) & (g2093) & (g2625)));
	assign g2632 = (((!g2093) & (!g2086) & (!g2085) & (g2084) & (g2071) & (g2074)) + ((!g2093) & (!g2086) & (g2085) & (!g2084) & (!g2071) & (g2074)) + ((!g2093) & (!g2086) & (g2085) & (g2084) & (!g2071) & (g2074)) + ((!g2093) & (!g2086) & (g2085) & (g2084) & (g2071) & (g2074)) + ((!g2093) & (g2086) & (!g2085) & (!g2084) & (g2071) & (!g2074)) + ((!g2093) & (g2086) & (!g2085) & (g2084) & (g2071) & (!g2074)) + ((!g2093) & (g2086) & (!g2085) & (g2084) & (g2071) & (g2074)) + ((!g2093) & (g2086) & (g2085) & (!g2084) & (!g2071) & (g2074)) + ((!g2093) & (g2086) & (g2085) & (!g2084) & (g2071) & (!g2074)) + ((!g2093) & (g2086) & (g2085) & (g2084) & (!g2071) & (g2074)) + ((!g2093) & (g2086) & (g2085) & (g2084) & (g2071) & (!g2074)) + ((!g2093) & (g2086) & (g2085) & (g2084) & (g2071) & (g2074)) + ((g2093) & (!g2086) & (!g2085) & (!g2084) & (!g2071) & (!g2074)) + ((g2093) & (!g2086) & (!g2085) & (g2084) & (!g2071) & (!g2074)) + ((g2093) & (!g2086) & (!g2085) & (g2084) & (g2071) & (g2074)) + ((g2093) & (!g2086) & (g2085) & (!g2084) & (!g2071) & (!g2074)) + ((g2093) & (!g2086) & (g2085) & (!g2084) & (!g2071) & (g2074)) + ((g2093) & (!g2086) & (g2085) & (g2084) & (!g2071) & (!g2074)) + ((g2093) & (!g2086) & (g2085) & (g2084) & (!g2071) & (g2074)) + ((g2093) & (!g2086) & (g2085) & (g2084) & (g2071) & (g2074)) + ((g2093) & (g2086) & (!g2085) & (!g2084) & (!g2071) & (!g2074)) + ((g2093) & (g2086) & (!g2085) & (!g2084) & (g2071) & (!g2074)) + ((g2093) & (g2086) & (!g2085) & (g2084) & (!g2071) & (!g2074)) + ((g2093) & (g2086) & (!g2085) & (g2084) & (g2071) & (!g2074)) + ((g2093) & (g2086) & (!g2085) & (g2084) & (g2071) & (g2074)) + ((g2093) & (g2086) & (g2085) & (!g2084) & (!g2071) & (!g2074)) + ((g2093) & (g2086) & (g2085) & (!g2084) & (!g2071) & (g2074)) + ((g2093) & (g2086) & (g2085) & (!g2084) & (g2071) & (!g2074)) + ((g2093) & (g2086) & (g2085) & (g2084) & (!g2071) & (!g2074)) + ((g2093) & (g2086) & (g2085) & (g2084) & (!g2071) & (g2074)) + ((g2093) & (g2086) & (g2085) & (g2084) & (g2071) & (!g2074)) + ((g2093) & (g2086) & (g2085) & (g2084) & (g2071) & (g2074)));
	assign g2633 = (((!g2632) & (!g2467) & (!g2559) & (g2372) & (g2076) & (g2077)) + ((!g2632) & (!g2467) & (g2559) & (!g2372) & (!g2076) & (g2077)) + ((!g2632) & (!g2467) & (g2559) & (g2372) & (!g2076) & (g2077)) + ((!g2632) & (!g2467) & (g2559) & (g2372) & (g2076) & (g2077)) + ((!g2632) & (g2467) & (!g2559) & (!g2372) & (g2076) & (!g2077)) + ((!g2632) & (g2467) & (!g2559) & (g2372) & (g2076) & (!g2077)) + ((!g2632) & (g2467) & (!g2559) & (g2372) & (g2076) & (g2077)) + ((!g2632) & (g2467) & (g2559) & (!g2372) & (!g2076) & (g2077)) + ((!g2632) & (g2467) & (g2559) & (!g2372) & (g2076) & (!g2077)) + ((!g2632) & (g2467) & (g2559) & (g2372) & (!g2076) & (g2077)) + ((!g2632) & (g2467) & (g2559) & (g2372) & (g2076) & (!g2077)) + ((!g2632) & (g2467) & (g2559) & (g2372) & (g2076) & (g2077)) + ((g2632) & (!g2467) & (!g2559) & (!g2372) & (!g2076) & (!g2077)) + ((g2632) & (!g2467) & (!g2559) & (g2372) & (!g2076) & (!g2077)) + ((g2632) & (!g2467) & (!g2559) & (g2372) & (g2076) & (g2077)) + ((g2632) & (!g2467) & (g2559) & (!g2372) & (!g2076) & (!g2077)) + ((g2632) & (!g2467) & (g2559) & (!g2372) & (!g2076) & (g2077)) + ((g2632) & (!g2467) & (g2559) & (g2372) & (!g2076) & (!g2077)) + ((g2632) & (!g2467) & (g2559) & (g2372) & (!g2076) & (g2077)) + ((g2632) & (!g2467) & (g2559) & (g2372) & (g2076) & (g2077)) + ((g2632) & (g2467) & (!g2559) & (!g2372) & (!g2076) & (!g2077)) + ((g2632) & (g2467) & (!g2559) & (!g2372) & (g2076) & (!g2077)) + ((g2632) & (g2467) & (!g2559) & (g2372) & (!g2076) & (!g2077)) + ((g2632) & (g2467) & (!g2559) & (g2372) & (g2076) & (!g2077)) + ((g2632) & (g2467) & (!g2559) & (g2372) & (g2076) & (g2077)) + ((g2632) & (g2467) & (g2559) & (!g2372) & (!g2076) & (!g2077)) + ((g2632) & (g2467) & (g2559) & (!g2372) & (!g2076) & (g2077)) + ((g2632) & (g2467) & (g2559) & (!g2372) & (g2076) & (!g2077)) + ((g2632) & (g2467) & (g2559) & (g2372) & (!g2076) & (!g2077)) + ((g2632) & (g2467) & (g2559) & (g2372) & (!g2076) & (g2077)) + ((g2632) & (g2467) & (g2559) & (g2372) & (g2076) & (!g2077)) + ((g2632) & (g2467) & (g2559) & (g2372) & (g2076) & (g2077)));
	assign g2634 = (((!g2633) & (!g2273) & (!g2274) & (g2191) & (g2073) & (g2125)) + ((!g2633) & (!g2273) & (g2274) & (!g2191) & (!g2073) & (g2125)) + ((!g2633) & (!g2273) & (g2274) & (g2191) & (!g2073) & (g2125)) + ((!g2633) & (!g2273) & (g2274) & (g2191) & (g2073) & (g2125)) + ((!g2633) & (g2273) & (!g2274) & (!g2191) & (g2073) & (!g2125)) + ((!g2633) & (g2273) & (!g2274) & (g2191) & (g2073) & (!g2125)) + ((!g2633) & (g2273) & (!g2274) & (g2191) & (g2073) & (g2125)) + ((!g2633) & (g2273) & (g2274) & (!g2191) & (!g2073) & (g2125)) + ((!g2633) & (g2273) & (g2274) & (!g2191) & (g2073) & (!g2125)) + ((!g2633) & (g2273) & (g2274) & (g2191) & (!g2073) & (g2125)) + ((!g2633) & (g2273) & (g2274) & (g2191) & (g2073) & (!g2125)) + ((!g2633) & (g2273) & (g2274) & (g2191) & (g2073) & (g2125)) + ((g2633) & (!g2273) & (!g2274) & (!g2191) & (!g2073) & (!g2125)) + ((g2633) & (!g2273) & (!g2274) & (g2191) & (!g2073) & (!g2125)) + ((g2633) & (!g2273) & (!g2274) & (g2191) & (g2073) & (g2125)) + ((g2633) & (!g2273) & (g2274) & (!g2191) & (!g2073) & (!g2125)) + ((g2633) & (!g2273) & (g2274) & (!g2191) & (!g2073) & (g2125)) + ((g2633) & (!g2273) & (g2274) & (g2191) & (!g2073) & (!g2125)) + ((g2633) & (!g2273) & (g2274) & (g2191) & (!g2073) & (g2125)) + ((g2633) & (!g2273) & (g2274) & (g2191) & (g2073) & (g2125)) + ((g2633) & (g2273) & (!g2274) & (!g2191) & (!g2073) & (!g2125)) + ((g2633) & (g2273) & (!g2274) & (!g2191) & (g2073) & (!g2125)) + ((g2633) & (g2273) & (!g2274) & (g2191) & (!g2073) & (!g2125)) + ((g2633) & (g2273) & (!g2274) & (g2191) & (g2073) & (!g2125)) + ((g2633) & (g2273) & (!g2274) & (g2191) & (g2073) & (g2125)) + ((g2633) & (g2273) & (g2274) & (!g2191) & (!g2073) & (!g2125)) + ((g2633) & (g2273) & (g2274) & (!g2191) & (!g2073) & (g2125)) + ((g2633) & (g2273) & (g2274) & (!g2191) & (g2073) & (!g2125)) + ((g2633) & (g2273) & (g2274) & (g2191) & (!g2073) & (!g2125)) + ((g2633) & (g2273) & (g2274) & (g2191) & (!g2073) & (g2125)) + ((g2633) & (g2273) & (g2274) & (g2191) & (g2073) & (!g2125)) + ((g2633) & (g2273) & (g2274) & (g2191) & (g2073) & (g2125)));
	assign g2635 = (((!g2093) & (!g2625) & (!g2124) & (!g2264) & (!g3455) & (g2634)) + ((!g2093) & (!g2625) & (!g2124) & (!g2264) & (g3455) & (g2634)) + ((!g2093) & (!g2625) & (!g2124) & (g2264) & (g3455) & (!g2634)) + ((!g2093) & (!g2625) & (!g2124) & (g2264) & (g3455) & (g2634)) + ((!g2093) & (g2625) & (!g2124) & (!g2264) & (!g3455) & (g2634)) + ((!g2093) & (g2625) & (!g2124) & (!g2264) & (g3455) & (g2634)) + ((!g2093) & (g2625) & (!g2124) & (g2264) & (g3455) & (!g2634)) + ((!g2093) & (g2625) & (!g2124) & (g2264) & (g3455) & (g2634)) + ((!g2093) & (g2625) & (g2124) & (!g2264) & (!g3455) & (!g2634)) + ((!g2093) & (g2625) & (g2124) & (!g2264) & (!g3455) & (g2634)) + ((!g2093) & (g2625) & (g2124) & (!g2264) & (g3455) & (!g2634)) + ((!g2093) & (g2625) & (g2124) & (!g2264) & (g3455) & (g2634)) + ((!g2093) & (g2625) & (g2124) & (g2264) & (!g3455) & (!g2634)) + ((!g2093) & (g2625) & (g2124) & (g2264) & (!g3455) & (g2634)) + ((!g2093) & (g2625) & (g2124) & (g2264) & (g3455) & (!g2634)) + ((!g2093) & (g2625) & (g2124) & (g2264) & (g3455) & (g2634)) + ((g2093) & (!g2625) & (!g2124) & (!g2264) & (!g3455) & (g2634)) + ((g2093) & (!g2625) & (!g2124) & (!g2264) & (g3455) & (g2634)) + ((g2093) & (!g2625) & (!g2124) & (g2264) & (g3455) & (!g2634)) + ((g2093) & (!g2625) & (!g2124) & (g2264) & (g3455) & (g2634)) + ((g2093) & (!g2625) & (g2124) & (!g2264) & (!g3455) & (!g2634)) + ((g2093) & (!g2625) & (g2124) & (!g2264) & (!g3455) & (g2634)) + ((g2093) & (!g2625) & (g2124) & (!g2264) & (g3455) & (!g2634)) + ((g2093) & (!g2625) & (g2124) & (!g2264) & (g3455) & (g2634)) + ((g2093) & (!g2625) & (g2124) & (g2264) & (!g3455) & (!g2634)) + ((g2093) & (!g2625) & (g2124) & (g2264) & (!g3455) & (g2634)) + ((g2093) & (!g2625) & (g2124) & (g2264) & (g3455) & (!g2634)) + ((g2093) & (!g2625) & (g2124) & (g2264) & (g3455) & (g2634)) + ((g2093) & (g2625) & (!g2124) & (!g2264) & (!g3455) & (g2634)) + ((g2093) & (g2625) & (!g2124) & (!g2264) & (g3455) & (g2634)) + ((g2093) & (g2625) & (!g2124) & (g2264) & (g3455) & (!g2634)) + ((g2093) & (g2625) & (!g2124) & (g2264) & (g3455) & (g2634)) + ((g2093) & (g2625) & (g2124) & (!g2264) & (!g3455) & (!g2634)) + ((g2093) & (g2625) & (g2124) & (!g2264) & (!g3455) & (g2634)) + ((g2093) & (g2625) & (g2124) & (!g2264) & (g3455) & (!g2634)) + ((g2093) & (g2625) & (g2124) & (!g2264) & (g3455) & (g2634)));
	assign g2636 = (((!g1050) & (!g2619) & (sk[78]) & (g1095)) + ((!g1050) & (g2619) & (!sk[78]) & (!g1095)) + ((!g1050) & (g2619) & (!sk[78]) & (g1095)) + ((!g1050) & (g2619) & (sk[78]) & (g1095)) + ((g1050) & (!g2619) & (sk[78]) & (g1095)) + ((g1050) & (g2619) & (!sk[78]) & (!g1095)) + ((g1050) & (g2619) & (!sk[78]) & (g1095)) + ((g1050) & (g2619) & (sk[78]) & (!g1095)));
	assign g2637 = (((!g165) & (!g166) & (!g1005) & (!g2601) & (!g2602) & (!g1050)) + ((!g165) & (!g166) & (!g1005) & (!g2601) & (!g2602) & (g1050)) + ((!g165) & (!g166) & (!g1005) & (!g2601) & (g2602) & (!g1050)) + ((!g165) & (!g166) & (!g1005) & (!g2601) & (g2602) & (g1050)) + ((!g165) & (!g166) & (!g1005) & (g2601) & (!g2602) & (!g1050)) + ((!g165) & (!g166) & (!g1005) & (g2601) & (!g2602) & (g1050)) + ((!g165) & (!g166) & (!g1005) & (g2601) & (g2602) & (!g1050)) + ((!g165) & (!g166) & (!g1005) & (g2601) & (g2602) & (g1050)) + ((!g165) & (!g166) & (g1005) & (!g2601) & (!g2602) & (!g1050)) + ((!g165) & (!g166) & (g1005) & (!g2601) & (!g2602) & (g1050)) + ((!g165) & (!g166) & (g1005) & (!g2601) & (g2602) & (!g1050)) + ((!g165) & (!g166) & (g1005) & (g2601) & (!g2602) & (!g1050)) + ((!g165) & (!g166) & (g1005) & (g2601) & (g2602) & (!g1050)) + ((!g165) & (g166) & (!g1005) & (!g2601) & (!g2602) & (!g1050)) + ((!g165) & (g166) & (!g1005) & (!g2601) & (g2602) & (!g1050)) + ((!g165) & (g166) & (!g1005) & (g2601) & (!g2602) & (!g1050)) + ((!g165) & (g166) & (!g1005) & (g2601) & (g2602) & (!g1050)) + ((!g165) & (g166) & (g1005) & (!g2601) & (!g2602) & (!g1050)) + ((g165) & (!g166) & (!g1005) & (!g2601) & (!g2602) & (!g1050)) + ((g165) & (!g166) & (!g1005) & (!g2601) & (!g2602) & (g1050)) + ((g165) & (!g166) & (!g1005) & (!g2601) & (g2602) & (!g1050)) + ((g165) & (!g166) & (!g1005) & (g2601) & (!g2602) & (!g1050)) + ((g165) & (!g166) & (!g1005) & (g2601) & (g2602) & (!g1050)) + ((g165) & (!g166) & (g1005) & (!g2601) & (!g2602) & (!g1050)) + ((g165) & (!g166) & (g1005) & (!g2601) & (g2602) & (!g1050)) + ((g165) & (!g166) & (g1005) & (g2601) & (!g2602) & (!g1050)) + ((g165) & (!g166) & (g1005) & (g2601) & (g2602) & (!g1050)) + ((g165) & (g166) & (!g1005) & (!g2601) & (!g2602) & (!g1050)));
	assign g2638 = (((!g148) & (!g1095) & (sk[80]) & (!g2637)) + ((!g148) & (g1095) & (!sk[80]) & (!g2637)) + ((!g148) & (g1095) & (!sk[80]) & (g2637)) + ((!g148) & (g1095) & (sk[80]) & (g2637)) + ((g148) & (!g1095) & (sk[80]) & (g2637)) + ((g148) & (g1095) & (!sk[80]) & (!g2637)) + ((g148) & (g1095) & (!sk[80]) & (g2637)) + ((g148) & (g1095) & (sk[80]) & (!g2637)));
	assign g5044 = (((!sk[81]) & (!g2921) & (g3093) & (!g2639)) + ((!sk[81]) & (!g2921) & (g3093) & (g2639)) + ((!sk[81]) & (g2921) & (g3093) & (!g2639)) + ((!sk[81]) & (g2921) & (g3093) & (g2639)) + ((sk[81]) & (!g2921) & (!g3093) & (g2639)) + ((sk[81]) & (!g2921) & (g3093) & (g2639)) + ((sk[81]) & (g2921) & (g3093) & (!g2639)) + ((sk[81]) & (g2921) & (g3093) & (g2639)));
	assign g2640 = (((!g1863) & (!g2033) & (!sk[82]) & (!g2034) & (g2638) & (!g2639)) + ((!g1863) & (!g2033) & (!sk[82]) & (!g2034) & (g2638) & (g2639)) + ((!g1863) & (!g2033) & (!sk[82]) & (g2034) & (g2638) & (!g2639)) + ((!g1863) & (!g2033) & (!sk[82]) & (g2034) & (g2638) & (g2639)) + ((!g1863) & (!g2033) & (sk[82]) & (!g2034) & (!g2638) & (g2639)) + ((!g1863) & (!g2033) & (sk[82]) & (!g2034) & (g2638) & (g2639)) + ((!g1863) & (g2033) & (!sk[82]) & (!g2034) & (!g2638) & (!g2639)) + ((!g1863) & (g2033) & (!sk[82]) & (!g2034) & (!g2638) & (g2639)) + ((!g1863) & (g2033) & (!sk[82]) & (!g2034) & (g2638) & (!g2639)) + ((!g1863) & (g2033) & (!sk[82]) & (!g2034) & (g2638) & (g2639)) + ((!g1863) & (g2033) & (!sk[82]) & (g2034) & (!g2638) & (!g2639)) + ((!g1863) & (g2033) & (!sk[82]) & (g2034) & (!g2638) & (g2639)) + ((!g1863) & (g2033) & (!sk[82]) & (g2034) & (g2638) & (!g2639)) + ((!g1863) & (g2033) & (!sk[82]) & (g2034) & (g2638) & (g2639)) + ((!g1863) & (g2033) & (sk[82]) & (!g2034) & (g2638) & (!g2639)) + ((!g1863) & (g2033) & (sk[82]) & (!g2034) & (g2638) & (g2639)) + ((g1863) & (!g2033) & (!sk[82]) & (!g2034) & (g2638) & (!g2639)) + ((g1863) & (!g2033) & (!sk[82]) & (!g2034) & (g2638) & (g2639)) + ((g1863) & (!g2033) & (!sk[82]) & (g2034) & (g2638) & (!g2639)) + ((g1863) & (!g2033) & (!sk[82]) & (g2034) & (g2638) & (g2639)) + ((g1863) & (!g2033) & (sk[82]) & (!g2034) & (!g2638) & (g2639)) + ((g1863) & (!g2033) & (sk[82]) & (!g2034) & (g2638) & (g2639)) + ((g1863) & (!g2033) & (sk[82]) & (g2034) & (!g2638) & (!g2639)) + ((g1863) & (!g2033) & (sk[82]) & (g2034) & (!g2638) & (g2639)) + ((g1863) & (!g2033) & (sk[82]) & (g2034) & (g2638) & (!g2639)) + ((g1863) & (!g2033) & (sk[82]) & (g2034) & (g2638) & (g2639)) + ((g1863) & (g2033) & (!sk[82]) & (!g2034) & (!g2638) & (!g2639)) + ((g1863) & (g2033) & (!sk[82]) & (!g2034) & (!g2638) & (g2639)) + ((g1863) & (g2033) & (!sk[82]) & (!g2034) & (g2638) & (!g2639)) + ((g1863) & (g2033) & (!sk[82]) & (!g2034) & (g2638) & (g2639)) + ((g1863) & (g2033) & (!sk[82]) & (g2034) & (!g2638) & (!g2639)) + ((g1863) & (g2033) & (!sk[82]) & (g2034) & (!g2638) & (g2639)) + ((g1863) & (g2033) & (!sk[82]) & (g2034) & (g2638) & (!g2639)) + ((g1863) & (g2033) & (!sk[82]) & (g2034) & (g2638) & (g2639)) + ((g1863) & (g2033) & (sk[82]) & (!g2034) & (g2638) & (!g2639)) + ((g1863) & (g2033) & (sk[82]) & (!g2034) & (g2638) & (g2639)));
	assign g2641 = (((!g2329) & (!g2029) & (!g2408) & (g2636) & (!sk[83]) & (!g2640)) + ((!g2329) & (!g2029) & (!g2408) & (g2636) & (!sk[83]) & (g2640)) + ((!g2329) & (!g2029) & (g2408) & (g2636) & (!sk[83]) & (!g2640)) + ((!g2329) & (!g2029) & (g2408) & (g2636) & (!sk[83]) & (g2640)) + ((!g2329) & (g2029) & (!g2408) & (!g2636) & (!sk[83]) & (!g2640)) + ((!g2329) & (g2029) & (!g2408) & (!g2636) & (!sk[83]) & (g2640)) + ((!g2329) & (g2029) & (!g2408) & (g2636) & (!sk[83]) & (!g2640)) + ((!g2329) & (g2029) & (!g2408) & (g2636) & (!sk[83]) & (g2640)) + ((!g2329) & (g2029) & (g2408) & (!g2636) & (!sk[83]) & (!g2640)) + ((!g2329) & (g2029) & (g2408) & (!g2636) & (!sk[83]) & (g2640)) + ((!g2329) & (g2029) & (g2408) & (g2636) & (!sk[83]) & (!g2640)) + ((!g2329) & (g2029) & (g2408) & (g2636) & (!sk[83]) & (g2640)) + ((g2329) & (!g2029) & (!g2408) & (g2636) & (!sk[83]) & (!g2640)) + ((g2329) & (!g2029) & (!g2408) & (g2636) & (!sk[83]) & (g2640)) + ((g2329) & (!g2029) & (g2408) & (!g2636) & (sk[83]) & (g2640)) + ((g2329) & (!g2029) & (g2408) & (g2636) & (!sk[83]) & (!g2640)) + ((g2329) & (!g2029) & (g2408) & (g2636) & (!sk[83]) & (g2640)) + ((g2329) & (!g2029) & (g2408) & (g2636) & (sk[83]) & (g2640)) + ((g2329) & (g2029) & (!g2408) & (!g2636) & (!sk[83]) & (!g2640)) + ((g2329) & (g2029) & (!g2408) & (!g2636) & (!sk[83]) & (g2640)) + ((g2329) & (g2029) & (!g2408) & (g2636) & (!sk[83]) & (!g2640)) + ((g2329) & (g2029) & (!g2408) & (g2636) & (!sk[83]) & (g2640)) + ((g2329) & (g2029) & (g2408) & (!g2636) & (!sk[83]) & (!g2640)) + ((g2329) & (g2029) & (g2408) & (!g2636) & (!sk[83]) & (g2640)) + ((g2329) & (g2029) & (g2408) & (g2636) & (!sk[83]) & (!g2640)) + ((g2329) & (g2029) & (g2408) & (g2636) & (!sk[83]) & (g2640)) + ((g2329) & (g2029) & (g2408) & (g2636) & (sk[83]) & (!g2640)) + ((g2329) & (g2029) & (g2408) & (g2636) & (sk[83]) & (g2640)));
	assign g2643 = (((!sk[84]) & (!g2093) & (g2625)) + ((!sk[84]) & (g2093) & (g2625)) + ((sk[84]) & (!g2093) & (g2625)) + ((sk[84]) & (g2093) & (!g2625)));
	assign g2644 = (((!g2085) & (!g2086) & (g2590) & (g2591) & (g2608) & (g2643)) + ((!g2085) & (g2086) & (!g2590) & (!g2591) & (g2608) & (g2643)) + ((!g2085) & (g2086) & (!g2590) & (g2591) & (g2608) & (g2643)) + ((!g2085) & (g2086) & (g2590) & (!g2591) & (g2608) & (g2643)) + ((!g2085) & (g2086) & (g2590) & (g2591) & (!g2608) & (g2643)) + ((!g2085) & (g2086) & (g2590) & (g2591) & (g2608) & (g2643)) + ((g2085) & (!g2086) & (!g2590) & (g2591) & (g2608) & (g2643)) + ((g2085) & (!g2086) & (g2590) & (!g2591) & (g2608) & (g2643)) + ((g2085) & (!g2086) & (g2590) & (g2591) & (g2608) & (g2643)) + ((g2085) & (g2086) & (!g2590) & (!g2591) & (g2608) & (g2643)) + ((g2085) & (g2086) & (!g2590) & (g2591) & (!g2608) & (g2643)) + ((g2085) & (g2086) & (!g2590) & (g2591) & (g2608) & (g2643)) + ((g2085) & (g2086) & (g2590) & (!g2591) & (!g2608) & (g2643)) + ((g2085) & (g2086) & (g2590) & (!g2591) & (g2608) & (g2643)) + ((g2085) & (g2086) & (g2590) & (g2591) & (!g2608) & (g2643)) + ((g2085) & (g2086) & (g2590) & (g2591) & (g2608) & (g2643)));
	assign g2645 = (((!g2644) & (!sk[86]) & (!g2631) & (g2094) & (!g2642)) + ((!g2644) & (!sk[86]) & (!g2631) & (g2094) & (g2642)) + ((!g2644) & (!sk[86]) & (g2631) & (!g2094) & (g2642)) + ((!g2644) & (!sk[86]) & (g2631) & (g2094) & (!g2642)) + ((!g2644) & (!sk[86]) & (g2631) & (g2094) & (g2642)) + ((!g2644) & (sk[86]) & (!g2631) & (!g2094) & (g2642)) + ((!g2644) & (sk[86]) & (!g2631) & (g2094) & (!g2642)) + ((!g2644) & (sk[86]) & (g2631) & (!g2094) & (!g2642)) + ((!g2644) & (sk[86]) & (g2631) & (g2094) & (g2642)) + ((g2644) & (!sk[86]) & (!g2631) & (!g2094) & (g2642)) + ((g2644) & (!sk[86]) & (!g2631) & (g2094) & (!g2642)) + ((g2644) & (!sk[86]) & (!g2631) & (g2094) & (g2642)) + ((g2644) & (!sk[86]) & (g2631) & (!g2094) & (g2642)) + ((g2644) & (!sk[86]) & (g2631) & (g2094) & (!g2642)) + ((g2644) & (!sk[86]) & (g2631) & (g2094) & (g2642)) + ((g2644) & (sk[86]) & (!g2631) & (!g2094) & (!g2642)) + ((g2644) & (sk[86]) & (!g2631) & (g2094) & (g2642)) + ((g2644) & (sk[86]) & (g2631) & (!g2094) & (!g2642)) + ((g2644) & (sk[86]) & (g2631) & (g2094) & (g2642)));
	assign g2646 = (((!g2609) & (!sk[87]) & (!g2610) & (g2626) & (!g2645)) + ((!g2609) & (!sk[87]) & (!g2610) & (g2626) & (g2645)) + ((!g2609) & (!sk[87]) & (g2610) & (!g2626) & (g2645)) + ((!g2609) & (!sk[87]) & (g2610) & (g2626) & (!g2645)) + ((!g2609) & (!sk[87]) & (g2610) & (g2626) & (g2645)) + ((!g2609) & (sk[87]) & (!g2610) & (!g2626) & (g2645)) + ((!g2609) & (sk[87]) & (!g2610) & (g2626) & (g2645)) + ((!g2609) & (sk[87]) & (g2610) & (!g2626) & (g2645)) + ((!g2609) & (sk[87]) & (g2610) & (g2626) & (g2645)) + ((g2609) & (!sk[87]) & (!g2610) & (!g2626) & (g2645)) + ((g2609) & (!sk[87]) & (!g2610) & (g2626) & (!g2645)) + ((g2609) & (!sk[87]) & (!g2610) & (g2626) & (g2645)) + ((g2609) & (!sk[87]) & (g2610) & (!g2626) & (g2645)) + ((g2609) & (!sk[87]) & (g2610) & (g2626) & (!g2645)) + ((g2609) & (!sk[87]) & (g2610) & (g2626) & (g2645)) + ((g2609) & (sk[87]) & (!g2610) & (!g2626) & (g2645)) + ((g2609) & (sk[87]) & (!g2610) & (g2626) & (g2645)) + ((g2609) & (sk[87]) & (g2610) & (!g2626) & (g2645)) + ((g2609) & (sk[87]) & (g2610) & (g2626) & (!g2645)));
	assign g2647 = (((!sk[88]) & (!g2625) & (g2093)) + ((!sk[88]) & (g2625) & (g2093)) + ((sk[88]) & (!g2625) & (g2093)));
	assign g2648 = (((!sk[89]) & (!g2642) & (g2094)) + ((!sk[89]) & (g2642) & (g2094)) + ((sk[89]) & (!g2642) & (!g2094)) + ((sk[89]) & (g2642) & (g2094)));
	assign g2649 = (((!g2627) & (!g2628) & (!g2629) & (!g2647) & (sk[90]) & (g2648)) + ((!g2627) & (!g2628) & (!g2629) & (g2647) & (!sk[90]) & (!g2648)) + ((!g2627) & (!g2628) & (!g2629) & (g2647) & (!sk[90]) & (g2648)) + ((!g2627) & (!g2628) & (!g2629) & (g2647) & (sk[90]) & (!g2648)) + ((!g2627) & (!g2628) & (g2629) & (!g2647) & (sk[90]) & (g2648)) + ((!g2627) & (!g2628) & (g2629) & (g2647) & (!sk[90]) & (!g2648)) + ((!g2627) & (!g2628) & (g2629) & (g2647) & (!sk[90]) & (g2648)) + ((!g2627) & (!g2628) & (g2629) & (g2647) & (sk[90]) & (!g2648)) + ((!g2627) & (g2628) & (!g2629) & (!g2647) & (!sk[90]) & (!g2648)) + ((!g2627) & (g2628) & (!g2629) & (!g2647) & (!sk[90]) & (g2648)) + ((!g2627) & (g2628) & (!g2629) & (!g2647) & (sk[90]) & (g2648)) + ((!g2627) & (g2628) & (!g2629) & (g2647) & (!sk[90]) & (!g2648)) + ((!g2627) & (g2628) & (!g2629) & (g2647) & (!sk[90]) & (g2648)) + ((!g2627) & (g2628) & (!g2629) & (g2647) & (sk[90]) & (!g2648)) + ((!g2627) & (g2628) & (g2629) & (!g2647) & (!sk[90]) & (!g2648)) + ((!g2627) & (g2628) & (g2629) & (!g2647) & (!sk[90]) & (g2648)) + ((!g2627) & (g2628) & (g2629) & (!g2647) & (sk[90]) & (!g2648)) + ((!g2627) & (g2628) & (g2629) & (g2647) & (!sk[90]) & (!g2648)) + ((!g2627) & (g2628) & (g2629) & (g2647) & (!sk[90]) & (g2648)) + ((!g2627) & (g2628) & (g2629) & (g2647) & (sk[90]) & (g2648)) + ((g2627) & (!g2628) & (!g2629) & (!g2647) & (sk[90]) & (g2648)) + ((g2627) & (!g2628) & (!g2629) & (g2647) & (!sk[90]) & (!g2648)) + ((g2627) & (!g2628) & (!g2629) & (g2647) & (!sk[90]) & (g2648)) + ((g2627) & (!g2628) & (!g2629) & (g2647) & (sk[90]) & (!g2648)) + ((g2627) & (!g2628) & (g2629) & (!g2647) & (sk[90]) & (!g2648)) + ((g2627) & (!g2628) & (g2629) & (g2647) & (!sk[90]) & (!g2648)) + ((g2627) & (!g2628) & (g2629) & (g2647) & (!sk[90]) & (g2648)) + ((g2627) & (!g2628) & (g2629) & (g2647) & (sk[90]) & (g2648)) + ((g2627) & (g2628) & (!g2629) & (!g2647) & (!sk[90]) & (!g2648)) + ((g2627) & (g2628) & (!g2629) & (!g2647) & (!sk[90]) & (g2648)) + ((g2627) & (g2628) & (!g2629) & (!g2647) & (sk[90]) & (!g2648)) + ((g2627) & (g2628) & (!g2629) & (g2647) & (!sk[90]) & (!g2648)) + ((g2627) & (g2628) & (!g2629) & (g2647) & (!sk[90]) & (g2648)) + ((g2627) & (g2628) & (!g2629) & (g2647) & (sk[90]) & (g2648)) + ((g2627) & (g2628) & (g2629) & (!g2647) & (!sk[90]) & (!g2648)) + ((g2627) & (g2628) & (g2629) & (!g2647) & (!sk[90]) & (g2648)) + ((g2627) & (g2628) & (g2629) & (!g2647) & (sk[90]) & (!g2648)) + ((g2627) & (g2628) & (g2629) & (g2647) & (!sk[90]) & (!g2648)) + ((g2627) & (g2628) & (g2629) & (g2647) & (!sk[90]) & (g2648)) + ((g2627) & (g2628) & (g2629) & (g2647) & (sk[90]) & (g2648)));
	assign g2650 = (((!g2094) & (!g2093) & (!g2086) & (g2085) & (g2071) & (g2074)) + ((!g2094) & (!g2093) & (g2086) & (!g2085) & (!g2071) & (g2074)) + ((!g2094) & (!g2093) & (g2086) & (g2085) & (!g2071) & (g2074)) + ((!g2094) & (!g2093) & (g2086) & (g2085) & (g2071) & (g2074)) + ((!g2094) & (g2093) & (!g2086) & (!g2085) & (g2071) & (!g2074)) + ((!g2094) & (g2093) & (!g2086) & (g2085) & (g2071) & (!g2074)) + ((!g2094) & (g2093) & (!g2086) & (g2085) & (g2071) & (g2074)) + ((!g2094) & (g2093) & (g2086) & (!g2085) & (!g2071) & (g2074)) + ((!g2094) & (g2093) & (g2086) & (!g2085) & (g2071) & (!g2074)) + ((!g2094) & (g2093) & (g2086) & (g2085) & (!g2071) & (g2074)) + ((!g2094) & (g2093) & (g2086) & (g2085) & (g2071) & (!g2074)) + ((!g2094) & (g2093) & (g2086) & (g2085) & (g2071) & (g2074)) + ((g2094) & (!g2093) & (!g2086) & (!g2085) & (!g2071) & (!g2074)) + ((g2094) & (!g2093) & (!g2086) & (g2085) & (!g2071) & (!g2074)) + ((g2094) & (!g2093) & (!g2086) & (g2085) & (g2071) & (g2074)) + ((g2094) & (!g2093) & (g2086) & (!g2085) & (!g2071) & (!g2074)) + ((g2094) & (!g2093) & (g2086) & (!g2085) & (!g2071) & (g2074)) + ((g2094) & (!g2093) & (g2086) & (g2085) & (!g2071) & (!g2074)) + ((g2094) & (!g2093) & (g2086) & (g2085) & (!g2071) & (g2074)) + ((g2094) & (!g2093) & (g2086) & (g2085) & (g2071) & (g2074)) + ((g2094) & (g2093) & (!g2086) & (!g2085) & (!g2071) & (!g2074)) + ((g2094) & (g2093) & (!g2086) & (!g2085) & (g2071) & (!g2074)) + ((g2094) & (g2093) & (!g2086) & (g2085) & (!g2071) & (!g2074)) + ((g2094) & (g2093) & (!g2086) & (g2085) & (g2071) & (!g2074)) + ((g2094) & (g2093) & (!g2086) & (g2085) & (g2071) & (g2074)) + ((g2094) & (g2093) & (g2086) & (!g2085) & (!g2071) & (!g2074)) + ((g2094) & (g2093) & (g2086) & (!g2085) & (!g2071) & (g2074)) + ((g2094) & (g2093) & (g2086) & (!g2085) & (g2071) & (!g2074)) + ((g2094) & (g2093) & (g2086) & (g2085) & (!g2071) & (!g2074)) + ((g2094) & (g2093) & (g2086) & (g2085) & (!g2071) & (g2074)) + ((g2094) & (g2093) & (g2086) & (g2085) & (g2071) & (!g2074)) + ((g2094) & (g2093) & (g2086) & (g2085) & (g2071) & (g2074)));
	assign g2651 = (((!g2650) & (!g2490) & (!g2580) & (g2402) & (g2076) & (g2077)) + ((!g2650) & (!g2490) & (g2580) & (!g2402) & (!g2076) & (g2077)) + ((!g2650) & (!g2490) & (g2580) & (g2402) & (!g2076) & (g2077)) + ((!g2650) & (!g2490) & (g2580) & (g2402) & (g2076) & (g2077)) + ((!g2650) & (g2490) & (!g2580) & (!g2402) & (g2076) & (!g2077)) + ((!g2650) & (g2490) & (!g2580) & (g2402) & (g2076) & (!g2077)) + ((!g2650) & (g2490) & (!g2580) & (g2402) & (g2076) & (g2077)) + ((!g2650) & (g2490) & (g2580) & (!g2402) & (!g2076) & (g2077)) + ((!g2650) & (g2490) & (g2580) & (!g2402) & (g2076) & (!g2077)) + ((!g2650) & (g2490) & (g2580) & (g2402) & (!g2076) & (g2077)) + ((!g2650) & (g2490) & (g2580) & (g2402) & (g2076) & (!g2077)) + ((!g2650) & (g2490) & (g2580) & (g2402) & (g2076) & (g2077)) + ((g2650) & (!g2490) & (!g2580) & (!g2402) & (!g2076) & (!g2077)) + ((g2650) & (!g2490) & (!g2580) & (g2402) & (!g2076) & (!g2077)) + ((g2650) & (!g2490) & (!g2580) & (g2402) & (g2076) & (g2077)) + ((g2650) & (!g2490) & (g2580) & (!g2402) & (!g2076) & (!g2077)) + ((g2650) & (!g2490) & (g2580) & (!g2402) & (!g2076) & (g2077)) + ((g2650) & (!g2490) & (g2580) & (g2402) & (!g2076) & (!g2077)) + ((g2650) & (!g2490) & (g2580) & (g2402) & (!g2076) & (g2077)) + ((g2650) & (!g2490) & (g2580) & (g2402) & (g2076) & (g2077)) + ((g2650) & (g2490) & (!g2580) & (!g2402) & (!g2076) & (!g2077)) + ((g2650) & (g2490) & (!g2580) & (!g2402) & (g2076) & (!g2077)) + ((g2650) & (g2490) & (!g2580) & (g2402) & (!g2076) & (!g2077)) + ((g2650) & (g2490) & (!g2580) & (g2402) & (g2076) & (!g2077)) + ((g2650) & (g2490) & (!g2580) & (g2402) & (g2076) & (g2077)) + ((g2650) & (g2490) & (g2580) & (!g2402) & (!g2076) & (!g2077)) + ((g2650) & (g2490) & (g2580) & (!g2402) & (!g2076) & (g2077)) + ((g2650) & (g2490) & (g2580) & (!g2402) & (g2076) & (!g2077)) + ((g2650) & (g2490) & (g2580) & (g2402) & (!g2076) & (!g2077)) + ((g2650) & (g2490) & (g2580) & (g2402) & (!g2076) & (g2077)) + ((g2650) & (g2490) & (g2580) & (g2402) & (g2076) & (!g2077)) + ((g2650) & (g2490) & (g2580) & (g2402) & (g2076) & (g2077)));
	assign g2652 = (((!g2651) & (!g2297) & (!g2299) & (g2191) & (g2073) & (g2125)) + ((!g2651) & (!g2297) & (g2299) & (!g2191) & (!g2073) & (g2125)) + ((!g2651) & (!g2297) & (g2299) & (g2191) & (!g2073) & (g2125)) + ((!g2651) & (!g2297) & (g2299) & (g2191) & (g2073) & (g2125)) + ((!g2651) & (g2297) & (!g2299) & (!g2191) & (g2073) & (!g2125)) + ((!g2651) & (g2297) & (!g2299) & (g2191) & (g2073) & (!g2125)) + ((!g2651) & (g2297) & (!g2299) & (g2191) & (g2073) & (g2125)) + ((!g2651) & (g2297) & (g2299) & (!g2191) & (!g2073) & (g2125)) + ((!g2651) & (g2297) & (g2299) & (!g2191) & (g2073) & (!g2125)) + ((!g2651) & (g2297) & (g2299) & (g2191) & (!g2073) & (g2125)) + ((!g2651) & (g2297) & (g2299) & (g2191) & (g2073) & (!g2125)) + ((!g2651) & (g2297) & (g2299) & (g2191) & (g2073) & (g2125)) + ((g2651) & (!g2297) & (!g2299) & (!g2191) & (!g2073) & (!g2125)) + ((g2651) & (!g2297) & (!g2299) & (g2191) & (!g2073) & (!g2125)) + ((g2651) & (!g2297) & (!g2299) & (g2191) & (g2073) & (g2125)) + ((g2651) & (!g2297) & (g2299) & (!g2191) & (!g2073) & (!g2125)) + ((g2651) & (!g2297) & (g2299) & (!g2191) & (!g2073) & (g2125)) + ((g2651) & (!g2297) & (g2299) & (g2191) & (!g2073) & (!g2125)) + ((g2651) & (!g2297) & (g2299) & (g2191) & (!g2073) & (g2125)) + ((g2651) & (!g2297) & (g2299) & (g2191) & (g2073) & (g2125)) + ((g2651) & (g2297) & (!g2299) & (!g2191) & (!g2073) & (!g2125)) + ((g2651) & (g2297) & (!g2299) & (!g2191) & (g2073) & (!g2125)) + ((g2651) & (g2297) & (!g2299) & (g2191) & (!g2073) & (!g2125)) + ((g2651) & (g2297) & (!g2299) & (g2191) & (g2073) & (!g2125)) + ((g2651) & (g2297) & (!g2299) & (g2191) & (g2073) & (g2125)) + ((g2651) & (g2297) & (g2299) & (!g2191) & (!g2073) & (!g2125)) + ((g2651) & (g2297) & (g2299) & (!g2191) & (!g2073) & (g2125)) + ((g2651) & (g2297) & (g2299) & (!g2191) & (g2073) & (!g2125)) + ((g2651) & (g2297) & (g2299) & (g2191) & (!g2073) & (!g2125)) + ((g2651) & (g2297) & (g2299) & (g2191) & (!g2073) & (g2125)) + ((g2651) & (g2297) & (g2299) & (g2191) & (g2073) & (!g2125)) + ((g2651) & (g2297) & (g2299) & (g2191) & (g2073) & (g2125)));
	assign g2653 = (((!g2094) & (!g2642) & (!g2124) & (!g2264) & (!g3431) & (g2652)) + ((!g2094) & (!g2642) & (!g2124) & (!g2264) & (g3431) & (g2652)) + ((!g2094) & (!g2642) & (!g2124) & (g2264) & (g3431) & (!g2652)) + ((!g2094) & (!g2642) & (!g2124) & (g2264) & (g3431) & (g2652)) + ((!g2094) & (g2642) & (!g2124) & (!g2264) & (!g3431) & (g2652)) + ((!g2094) & (g2642) & (!g2124) & (!g2264) & (g3431) & (g2652)) + ((!g2094) & (g2642) & (!g2124) & (g2264) & (g3431) & (!g2652)) + ((!g2094) & (g2642) & (!g2124) & (g2264) & (g3431) & (g2652)) + ((!g2094) & (g2642) & (g2124) & (!g2264) & (!g3431) & (!g2652)) + ((!g2094) & (g2642) & (g2124) & (!g2264) & (!g3431) & (g2652)) + ((!g2094) & (g2642) & (g2124) & (!g2264) & (g3431) & (!g2652)) + ((!g2094) & (g2642) & (g2124) & (!g2264) & (g3431) & (g2652)) + ((!g2094) & (g2642) & (g2124) & (g2264) & (!g3431) & (!g2652)) + ((!g2094) & (g2642) & (g2124) & (g2264) & (!g3431) & (g2652)) + ((!g2094) & (g2642) & (g2124) & (g2264) & (g3431) & (!g2652)) + ((!g2094) & (g2642) & (g2124) & (g2264) & (g3431) & (g2652)) + ((g2094) & (!g2642) & (!g2124) & (!g2264) & (!g3431) & (g2652)) + ((g2094) & (!g2642) & (!g2124) & (!g2264) & (g3431) & (g2652)) + ((g2094) & (!g2642) & (!g2124) & (g2264) & (g3431) & (!g2652)) + ((g2094) & (!g2642) & (!g2124) & (g2264) & (g3431) & (g2652)) + ((g2094) & (!g2642) & (g2124) & (!g2264) & (!g3431) & (!g2652)) + ((g2094) & (!g2642) & (g2124) & (!g2264) & (!g3431) & (g2652)) + ((g2094) & (!g2642) & (g2124) & (!g2264) & (g3431) & (!g2652)) + ((g2094) & (!g2642) & (g2124) & (!g2264) & (g3431) & (g2652)) + ((g2094) & (!g2642) & (g2124) & (g2264) & (!g3431) & (!g2652)) + ((g2094) & (!g2642) & (g2124) & (g2264) & (!g3431) & (g2652)) + ((g2094) & (!g2642) & (g2124) & (g2264) & (g3431) & (!g2652)) + ((g2094) & (!g2642) & (g2124) & (g2264) & (g3431) & (g2652)) + ((g2094) & (g2642) & (!g2124) & (!g2264) & (!g3431) & (g2652)) + ((g2094) & (g2642) & (!g2124) & (!g2264) & (g3431) & (g2652)) + ((g2094) & (g2642) & (!g2124) & (g2264) & (g3431) & (!g2652)) + ((g2094) & (g2642) & (!g2124) & (g2264) & (g3431) & (g2652)) + ((g2094) & (g2642) & (g2124) & (!g2264) & (!g3431) & (!g2652)) + ((g2094) & (g2642) & (g2124) & (!g2264) & (!g3431) & (g2652)) + ((g2094) & (g2642) & (g2124) & (!g2264) & (g3431) & (!g2652)) + ((g2094) & (g2642) & (g2124) & (!g2264) & (g3431) & (g2652)));
	assign g2654 = (((!g1050) & (!g2619) & (!g1095) & (sk[95]) & (g1140)) + ((!g1050) & (!g2619) & (g1095) & (!sk[95]) & (!g1140)) + ((!g1050) & (!g2619) & (g1095) & (!sk[95]) & (g1140)) + ((!g1050) & (!g2619) & (g1095) & (sk[95]) & (g1140)) + ((!g1050) & (g2619) & (!g1095) & (!sk[95]) & (g1140)) + ((!g1050) & (g2619) & (!g1095) & (sk[95]) & (g1140)) + ((!g1050) & (g2619) & (g1095) & (!sk[95]) & (!g1140)) + ((!g1050) & (g2619) & (g1095) & (!sk[95]) & (g1140)) + ((!g1050) & (g2619) & (g1095) & (sk[95]) & (g1140)) + ((g1050) & (!g2619) & (!g1095) & (!sk[95]) & (g1140)) + ((g1050) & (!g2619) & (!g1095) & (sk[95]) & (g1140)) + ((g1050) & (!g2619) & (g1095) & (!sk[95]) & (!g1140)) + ((g1050) & (!g2619) & (g1095) & (!sk[95]) & (g1140)) + ((g1050) & (!g2619) & (g1095) & (sk[95]) & (g1140)) + ((g1050) & (g2619) & (!g1095) & (!sk[95]) & (g1140)) + ((g1050) & (g2619) & (!g1095) & (sk[95]) & (g1140)) + ((g1050) & (g2619) & (g1095) & (!sk[95]) & (!g1140)) + ((g1050) & (g2619) & (g1095) & (!sk[95]) & (g1140)) + ((g1050) & (g2619) & (g1095) & (sk[95]) & (!g1140)));
	assign g2655 = (((!g148) & (!sk[96]) & (g1095) & (!g2637)) + ((!g148) & (!sk[96]) & (g1095) & (g2637)) + ((!g148) & (sk[96]) & (g1095) & (!g2637)) + ((g148) & (!sk[96]) & (g1095) & (!g2637)) + ((g148) & (!sk[96]) & (g1095) & (g2637)) + ((g148) & (sk[96]) & (!g1095) & (!g2637)) + ((g148) & (sk[96]) & (g1095) & (!g2637)) + ((g148) & (sk[96]) & (g1095) & (g2637)));
	assign g2656 = (((!g147) & (!g2585) & (g1140) & (!sk[97]) & (!g2655)) + ((!g147) & (!g2585) & (g1140) & (!sk[97]) & (g2655)) + ((!g147) & (g2585) & (!g1140) & (!sk[97]) & (g2655)) + ((!g147) & (g2585) & (!g1140) & (sk[97]) & (g2655)) + ((!g147) & (g2585) & (g1140) & (!sk[97]) & (!g2655)) + ((!g147) & (g2585) & (g1140) & (!sk[97]) & (g2655)) + ((!g147) & (g2585) & (g1140) & (sk[97]) & (!g2655)) + ((g147) & (!g2585) & (!g1140) & (!sk[97]) & (g2655)) + ((g147) & (!g2585) & (g1140) & (!sk[97]) & (!g2655)) + ((g147) & (!g2585) & (g1140) & (!sk[97]) & (g2655)) + ((g147) & (g2585) & (!g1140) & (!sk[97]) & (g2655)) + ((g147) & (g2585) & (!g1140) & (sk[97]) & (!g2655)) + ((g147) & (g2585) & (g1140) & (!sk[97]) & (!g2655)) + ((g147) & (g2585) & (g1140) & (!sk[97]) & (g2655)) + ((g147) & (g2585) & (g1140) & (sk[97]) & (g2655)));
	assign g5045 = (((!g2921) & (!sk[98]) & (g3187) & (!g2657)) + ((!g2921) & (!sk[98]) & (g3187) & (g2657)) + ((!g2921) & (sk[98]) & (!g3187) & (g2657)) + ((!g2921) & (sk[98]) & (g3187) & (g2657)) + ((g2921) & (!sk[98]) & (g3187) & (!g2657)) + ((g2921) & (!sk[98]) & (g3187) & (g2657)) + ((g2921) & (sk[98]) & (g3187) & (!g2657)) + ((g2921) & (sk[98]) & (g3187) & (g2657)));
	assign g2658 = (((!g1876) & (!sk[99]) & (!g2033) & (g2034) & (!g2657)) + ((!g1876) & (!sk[99]) & (!g2033) & (g2034) & (g2657)) + ((!g1876) & (!sk[99]) & (g2033) & (!g2034) & (g2657)) + ((!g1876) & (!sk[99]) & (g2033) & (g2034) & (!g2657)) + ((!g1876) & (!sk[99]) & (g2033) & (g2034) & (g2657)) + ((!g1876) & (sk[99]) & (!g2033) & (!g2034) & (g2657)) + ((g1876) & (!sk[99]) & (!g2033) & (!g2034) & (g2657)) + ((g1876) & (!sk[99]) & (!g2033) & (g2034) & (!g2657)) + ((g1876) & (!sk[99]) & (!g2033) & (g2034) & (g2657)) + ((g1876) & (!sk[99]) & (g2033) & (!g2034) & (g2657)) + ((g1876) & (!sk[99]) & (g2033) & (g2034) & (!g2657)) + ((g1876) & (!sk[99]) & (g2033) & (g2034) & (g2657)) + ((g1876) & (sk[99]) & (!g2033) & (!g2034) & (g2657)) + ((g1876) & (sk[99]) & (!g2033) & (g2034) & (!g2657)) + ((g1876) & (sk[99]) & (!g2033) & (g2034) & (g2657)));
	assign g2659 = (((g2329) & (!g2029) & (g2408) & (!g2654) & (!g2656) & (g2658)) + ((g2329) & (!g2029) & (g2408) & (!g2654) & (g2656) & (!g2658)) + ((g2329) & (!g2029) & (g2408) & (!g2654) & (g2656) & (g2658)) + ((g2329) & (!g2029) & (g2408) & (g2654) & (!g2656) & (g2658)) + ((g2329) & (!g2029) & (g2408) & (g2654) & (g2656) & (!g2658)) + ((g2329) & (!g2029) & (g2408) & (g2654) & (g2656) & (g2658)) + ((g2329) & (g2029) & (g2408) & (g2654) & (!g2656) & (!g2658)) + ((g2329) & (g2029) & (g2408) & (g2654) & (!g2656) & (g2658)) + ((g2329) & (g2029) & (g2408) & (g2654) & (g2656) & (!g2658)) + ((g2329) & (g2029) & (g2408) & (g2654) & (g2656) & (g2658)));
	assign g2661 = (((!g2094) & (!g2095) & (!g2642) & (g2660) & (!g2644) & (!g2631)) + ((!g2094) & (!g2095) & (!g2642) & (g2660) & (!g2644) & (g2631)) + ((!g2094) & (!g2095) & (!g2642) & (g2660) & (g2644) & (!g2631)) + ((!g2094) & (!g2095) & (!g2642) & (g2660) & (g2644) & (g2631)) + ((!g2094) & (!g2095) & (g2642) & (!g2660) & (!g2644) & (g2631)) + ((!g2094) & (!g2095) & (g2642) & (!g2660) & (g2644) & (!g2631)) + ((!g2094) & (!g2095) & (g2642) & (!g2660) & (g2644) & (g2631)) + ((!g2094) & (!g2095) & (g2642) & (g2660) & (!g2644) & (!g2631)) + ((!g2094) & (g2095) & (!g2642) & (!g2660) & (!g2644) & (!g2631)) + ((!g2094) & (g2095) & (!g2642) & (!g2660) & (!g2644) & (g2631)) + ((!g2094) & (g2095) & (!g2642) & (!g2660) & (g2644) & (!g2631)) + ((!g2094) & (g2095) & (!g2642) & (!g2660) & (g2644) & (g2631)) + ((!g2094) & (g2095) & (g2642) & (!g2660) & (!g2644) & (!g2631)) + ((!g2094) & (g2095) & (g2642) & (g2660) & (!g2644) & (g2631)) + ((!g2094) & (g2095) & (g2642) & (g2660) & (g2644) & (!g2631)) + ((!g2094) & (g2095) & (g2642) & (g2660) & (g2644) & (g2631)) + ((g2094) & (!g2095) & (!g2642) & (!g2660) & (!g2644) & (g2631)) + ((g2094) & (!g2095) & (!g2642) & (!g2660) & (g2644) & (!g2631)) + ((g2094) & (!g2095) & (!g2642) & (!g2660) & (g2644) & (g2631)) + ((g2094) & (!g2095) & (!g2642) & (g2660) & (!g2644) & (!g2631)) + ((g2094) & (!g2095) & (g2642) & (!g2660) & (!g2644) & (!g2631)) + ((g2094) & (!g2095) & (g2642) & (!g2660) & (!g2644) & (g2631)) + ((g2094) & (!g2095) & (g2642) & (!g2660) & (g2644) & (!g2631)) + ((g2094) & (!g2095) & (g2642) & (!g2660) & (g2644) & (g2631)) + ((g2094) & (g2095) & (!g2642) & (!g2660) & (!g2644) & (!g2631)) + ((g2094) & (g2095) & (!g2642) & (g2660) & (!g2644) & (g2631)) + ((g2094) & (g2095) & (!g2642) & (g2660) & (g2644) & (!g2631)) + ((g2094) & (g2095) & (!g2642) & (g2660) & (g2644) & (g2631)) + ((g2094) & (g2095) & (g2642) & (g2660) & (!g2644) & (!g2631)) + ((g2094) & (g2095) & (g2642) & (g2660) & (!g2644) & (g2631)) + ((g2094) & (g2095) & (g2642) & (g2660) & (g2644) & (!g2631)) + ((g2094) & (g2095) & (g2642) & (g2660) & (g2644) & (g2631)));
	assign g2662 = (((g2609) & (g2610) & (g2626) & (!g2644) & (!g2631) & (!g3126)) + ((g2609) & (g2610) & (g2626) & (!g2644) & (g2631) & (g3126)) + ((g2609) & (g2610) & (g2626) & (g2644) & (!g2631) & (g3126)) + ((g2609) & (g2610) & (g2626) & (g2644) & (g2631) & (g3126)));
	assign g2663 = (((!g2647) & (!sk[103]) & (g2648)) + ((!g2647) & (sk[103]) & (g2648)) + ((g2647) & (!sk[103]) & (g2648)) + ((g2647) & (sk[103]) & (!g2648)));
	assign g2664 = (((!g2611) & (!g2612) & (!g2613) & (g2628) & (g2629) & (g2663)) + ((!g2611) & (!g2612) & (g2613) & (!g2628) & (g2629) & (g2663)) + ((!g2611) & (!g2612) & (g2613) & (g2628) & (!g2629) & (g2663)) + ((!g2611) & (!g2612) & (g2613) & (g2628) & (g2629) & (g2663)) + ((!g2611) & (g2612) & (!g2613) & (!g2628) & (g2629) & (g2663)) + ((!g2611) & (g2612) & (!g2613) & (g2628) & (!g2629) & (g2663)) + ((!g2611) & (g2612) & (!g2613) & (g2628) & (g2629) & (g2663)) + ((!g2611) & (g2612) & (g2613) & (!g2628) & (g2629) & (g2663)) + ((!g2611) & (g2612) & (g2613) & (g2628) & (!g2629) & (g2663)) + ((!g2611) & (g2612) & (g2613) & (g2628) & (g2629) & (g2663)) + ((g2611) & (!g2612) & (!g2613) & (g2628) & (g2629) & (g2663)) + ((g2611) & (!g2612) & (g2613) & (g2628) & (g2629) & (g2663)) + ((g2611) & (g2612) & (!g2613) & (g2628) & (g2629) & (g2663)) + ((g2611) & (g2612) & (g2613) & (!g2628) & (g2629) & (g2663)) + ((g2611) & (g2612) & (g2613) & (g2628) & (!g2629) & (g2663)) + ((g2611) & (g2612) & (g2613) & (g2628) & (g2629) & (g2663)));
	assign g2665 = (((!g2647) & (!sk[105]) & (g2648)) + ((g2647) & (!sk[105]) & (g2648)) + ((g2647) & (sk[105]) & (g2648)));
	assign g2666 = (((!sk[106]) & (!g2642) & (g2094)) + ((!sk[106]) & (g2642) & (g2094)) + ((sk[106]) & (!g2642) & (g2094)));
	assign g2667 = (((!g2660) & (!sk[107]) & (g2095)) + ((!g2660) & (sk[107]) & (!g2095)) + ((g2660) & (!sk[107]) & (g2095)) + ((g2660) & (sk[107]) & (g2095)));
	assign g2668 = (((!g2664) & (!sk[108]) & (!g2665) & (g2666) & (!g2667)) + ((!g2664) & (!sk[108]) & (!g2665) & (g2666) & (g2667)) + ((!g2664) & (!sk[108]) & (g2665) & (!g2666) & (g2667)) + ((!g2664) & (!sk[108]) & (g2665) & (g2666) & (!g2667)) + ((!g2664) & (!sk[108]) & (g2665) & (g2666) & (g2667)) + ((!g2664) & (sk[108]) & (!g2665) & (!g2666) & (g2667)) + ((!g2664) & (sk[108]) & (!g2665) & (g2666) & (!g2667)) + ((!g2664) & (sk[108]) & (g2665) & (!g2666) & (!g2667)) + ((!g2664) & (sk[108]) & (g2665) & (g2666) & (g2667)) + ((g2664) & (!sk[108]) & (!g2665) & (!g2666) & (g2667)) + ((g2664) & (!sk[108]) & (!g2665) & (g2666) & (!g2667)) + ((g2664) & (!sk[108]) & (!g2665) & (g2666) & (g2667)) + ((g2664) & (!sk[108]) & (g2665) & (!g2666) & (g2667)) + ((g2664) & (!sk[108]) & (g2665) & (g2666) & (!g2667)) + ((g2664) & (!sk[108]) & (g2665) & (g2666) & (g2667)) + ((g2664) & (sk[108]) & (!g2665) & (!g2666) & (!g2667)) + ((g2664) & (sk[108]) & (!g2665) & (g2666) & (g2667)) + ((g2664) & (sk[108]) & (g2665) & (!g2666) & (!g2667)) + ((g2664) & (sk[108]) & (g2665) & (g2666) & (g2667)));
	assign g2669 = (((!g2095) & (!g2094) & (!g2093) & (g2086) & (g2071) & (g2074)) + ((!g2095) & (!g2094) & (g2093) & (!g2086) & (!g2071) & (g2074)) + ((!g2095) & (!g2094) & (g2093) & (g2086) & (!g2071) & (g2074)) + ((!g2095) & (!g2094) & (g2093) & (g2086) & (g2071) & (g2074)) + ((!g2095) & (g2094) & (!g2093) & (!g2086) & (g2071) & (!g2074)) + ((!g2095) & (g2094) & (!g2093) & (g2086) & (g2071) & (!g2074)) + ((!g2095) & (g2094) & (!g2093) & (g2086) & (g2071) & (g2074)) + ((!g2095) & (g2094) & (g2093) & (!g2086) & (!g2071) & (g2074)) + ((!g2095) & (g2094) & (g2093) & (!g2086) & (g2071) & (!g2074)) + ((!g2095) & (g2094) & (g2093) & (g2086) & (!g2071) & (g2074)) + ((!g2095) & (g2094) & (g2093) & (g2086) & (g2071) & (!g2074)) + ((!g2095) & (g2094) & (g2093) & (g2086) & (g2071) & (g2074)) + ((g2095) & (!g2094) & (!g2093) & (!g2086) & (!g2071) & (!g2074)) + ((g2095) & (!g2094) & (!g2093) & (g2086) & (!g2071) & (!g2074)) + ((g2095) & (!g2094) & (!g2093) & (g2086) & (g2071) & (g2074)) + ((g2095) & (!g2094) & (g2093) & (!g2086) & (!g2071) & (!g2074)) + ((g2095) & (!g2094) & (g2093) & (!g2086) & (!g2071) & (g2074)) + ((g2095) & (!g2094) & (g2093) & (g2086) & (!g2071) & (!g2074)) + ((g2095) & (!g2094) & (g2093) & (g2086) & (!g2071) & (g2074)) + ((g2095) & (!g2094) & (g2093) & (g2086) & (g2071) & (g2074)) + ((g2095) & (g2094) & (!g2093) & (!g2086) & (!g2071) & (!g2074)) + ((g2095) & (g2094) & (!g2093) & (!g2086) & (g2071) & (!g2074)) + ((g2095) & (g2094) & (!g2093) & (g2086) & (!g2071) & (!g2074)) + ((g2095) & (g2094) & (!g2093) & (g2086) & (g2071) & (!g2074)) + ((g2095) & (g2094) & (!g2093) & (g2086) & (g2071) & (g2074)) + ((g2095) & (g2094) & (g2093) & (!g2086) & (!g2071) & (!g2074)) + ((g2095) & (g2094) & (g2093) & (!g2086) & (!g2071) & (g2074)) + ((g2095) & (g2094) & (g2093) & (!g2086) & (g2071) & (!g2074)) + ((g2095) & (g2094) & (g2093) & (g2086) & (!g2071) & (!g2074)) + ((g2095) & (g2094) & (g2093) & (g2086) & (!g2071) & (g2074)) + ((g2095) & (g2094) & (g2093) & (g2086) & (g2071) & (!g2074)) + ((g2095) & (g2094) & (g2093) & (g2086) & (g2071) & (g2074)));
	assign g2670 = (((!g2669) & (!g2514) & (!g2595) & (g2426) & (g2076) & (g2077)) + ((!g2669) & (!g2514) & (g2595) & (!g2426) & (!g2076) & (g2077)) + ((!g2669) & (!g2514) & (g2595) & (g2426) & (!g2076) & (g2077)) + ((!g2669) & (!g2514) & (g2595) & (g2426) & (g2076) & (g2077)) + ((!g2669) & (g2514) & (!g2595) & (!g2426) & (g2076) & (!g2077)) + ((!g2669) & (g2514) & (!g2595) & (g2426) & (g2076) & (!g2077)) + ((!g2669) & (g2514) & (!g2595) & (g2426) & (g2076) & (g2077)) + ((!g2669) & (g2514) & (g2595) & (!g2426) & (!g2076) & (g2077)) + ((!g2669) & (g2514) & (g2595) & (!g2426) & (g2076) & (!g2077)) + ((!g2669) & (g2514) & (g2595) & (g2426) & (!g2076) & (g2077)) + ((!g2669) & (g2514) & (g2595) & (g2426) & (g2076) & (!g2077)) + ((!g2669) & (g2514) & (g2595) & (g2426) & (g2076) & (g2077)) + ((g2669) & (!g2514) & (!g2595) & (!g2426) & (!g2076) & (!g2077)) + ((g2669) & (!g2514) & (!g2595) & (g2426) & (!g2076) & (!g2077)) + ((g2669) & (!g2514) & (!g2595) & (g2426) & (g2076) & (g2077)) + ((g2669) & (!g2514) & (g2595) & (!g2426) & (!g2076) & (!g2077)) + ((g2669) & (!g2514) & (g2595) & (!g2426) & (!g2076) & (g2077)) + ((g2669) & (!g2514) & (g2595) & (g2426) & (!g2076) & (!g2077)) + ((g2669) & (!g2514) & (g2595) & (g2426) & (!g2076) & (g2077)) + ((g2669) & (!g2514) & (g2595) & (g2426) & (g2076) & (g2077)) + ((g2669) & (g2514) & (!g2595) & (!g2426) & (!g2076) & (!g2077)) + ((g2669) & (g2514) & (!g2595) & (!g2426) & (g2076) & (!g2077)) + ((g2669) & (g2514) & (!g2595) & (g2426) & (!g2076) & (!g2077)) + ((g2669) & (g2514) & (!g2595) & (g2426) & (g2076) & (!g2077)) + ((g2669) & (g2514) & (!g2595) & (g2426) & (g2076) & (g2077)) + ((g2669) & (g2514) & (g2595) & (!g2426) & (!g2076) & (!g2077)) + ((g2669) & (g2514) & (g2595) & (!g2426) & (!g2076) & (g2077)) + ((g2669) & (g2514) & (g2595) & (!g2426) & (g2076) & (!g2077)) + ((g2669) & (g2514) & (g2595) & (g2426) & (!g2076) & (!g2077)) + ((g2669) & (g2514) & (g2595) & (g2426) & (!g2076) & (g2077)) + ((g2669) & (g2514) & (g2595) & (g2426) & (g2076) & (!g2077)) + ((g2669) & (g2514) & (g2595) & (g2426) & (g2076) & (g2077)));
	assign g2671 = (((!g2670) & (!g2321) & (!g2323) & (g2191) & (g2073) & (g2125)) + ((!g2670) & (!g2321) & (g2323) & (!g2191) & (!g2073) & (g2125)) + ((!g2670) & (!g2321) & (g2323) & (g2191) & (!g2073) & (g2125)) + ((!g2670) & (!g2321) & (g2323) & (g2191) & (g2073) & (g2125)) + ((!g2670) & (g2321) & (!g2323) & (!g2191) & (g2073) & (!g2125)) + ((!g2670) & (g2321) & (!g2323) & (g2191) & (g2073) & (!g2125)) + ((!g2670) & (g2321) & (!g2323) & (g2191) & (g2073) & (g2125)) + ((!g2670) & (g2321) & (g2323) & (!g2191) & (!g2073) & (g2125)) + ((!g2670) & (g2321) & (g2323) & (!g2191) & (g2073) & (!g2125)) + ((!g2670) & (g2321) & (g2323) & (g2191) & (!g2073) & (g2125)) + ((!g2670) & (g2321) & (g2323) & (g2191) & (g2073) & (!g2125)) + ((!g2670) & (g2321) & (g2323) & (g2191) & (g2073) & (g2125)) + ((g2670) & (!g2321) & (!g2323) & (!g2191) & (!g2073) & (!g2125)) + ((g2670) & (!g2321) & (!g2323) & (g2191) & (!g2073) & (!g2125)) + ((g2670) & (!g2321) & (!g2323) & (g2191) & (g2073) & (g2125)) + ((g2670) & (!g2321) & (g2323) & (!g2191) & (!g2073) & (!g2125)) + ((g2670) & (!g2321) & (g2323) & (!g2191) & (!g2073) & (g2125)) + ((g2670) & (!g2321) & (g2323) & (g2191) & (!g2073) & (!g2125)) + ((g2670) & (!g2321) & (g2323) & (g2191) & (!g2073) & (g2125)) + ((g2670) & (!g2321) & (g2323) & (g2191) & (g2073) & (g2125)) + ((g2670) & (g2321) & (!g2323) & (!g2191) & (!g2073) & (!g2125)) + ((g2670) & (g2321) & (!g2323) & (!g2191) & (g2073) & (!g2125)) + ((g2670) & (g2321) & (!g2323) & (g2191) & (!g2073) & (!g2125)) + ((g2670) & (g2321) & (!g2323) & (g2191) & (g2073) & (!g2125)) + ((g2670) & (g2321) & (!g2323) & (g2191) & (g2073) & (g2125)) + ((g2670) & (g2321) & (g2323) & (!g2191) & (!g2073) & (!g2125)) + ((g2670) & (g2321) & (g2323) & (!g2191) & (!g2073) & (g2125)) + ((g2670) & (g2321) & (g2323) & (!g2191) & (g2073) & (!g2125)) + ((g2670) & (g2321) & (g2323) & (g2191) & (!g2073) & (!g2125)) + ((g2670) & (g2321) & (g2323) & (g2191) & (!g2073) & (g2125)) + ((g2670) & (g2321) & (g2323) & (g2191) & (g2073) & (!g2125)) + ((g2670) & (g2321) & (g2323) & (g2191) & (g2073) & (g2125)));
	assign g2672 = (((!g2095) & (!g2660) & (!g2124) & (!g2264) & (!g3408) & (g2671)) + ((!g2095) & (!g2660) & (!g2124) & (!g2264) & (g3408) & (g2671)) + ((!g2095) & (!g2660) & (!g2124) & (g2264) & (g3408) & (!g2671)) + ((!g2095) & (!g2660) & (!g2124) & (g2264) & (g3408) & (g2671)) + ((!g2095) & (g2660) & (!g2124) & (!g2264) & (!g3408) & (g2671)) + ((!g2095) & (g2660) & (!g2124) & (!g2264) & (g3408) & (g2671)) + ((!g2095) & (g2660) & (!g2124) & (g2264) & (g3408) & (!g2671)) + ((!g2095) & (g2660) & (!g2124) & (g2264) & (g3408) & (g2671)) + ((!g2095) & (g2660) & (g2124) & (!g2264) & (!g3408) & (!g2671)) + ((!g2095) & (g2660) & (g2124) & (!g2264) & (!g3408) & (g2671)) + ((!g2095) & (g2660) & (g2124) & (!g2264) & (g3408) & (!g2671)) + ((!g2095) & (g2660) & (g2124) & (!g2264) & (g3408) & (g2671)) + ((!g2095) & (g2660) & (g2124) & (g2264) & (!g3408) & (!g2671)) + ((!g2095) & (g2660) & (g2124) & (g2264) & (!g3408) & (g2671)) + ((!g2095) & (g2660) & (g2124) & (g2264) & (g3408) & (!g2671)) + ((!g2095) & (g2660) & (g2124) & (g2264) & (g3408) & (g2671)) + ((g2095) & (!g2660) & (!g2124) & (!g2264) & (!g3408) & (g2671)) + ((g2095) & (!g2660) & (!g2124) & (!g2264) & (g3408) & (g2671)) + ((g2095) & (!g2660) & (!g2124) & (g2264) & (g3408) & (!g2671)) + ((g2095) & (!g2660) & (!g2124) & (g2264) & (g3408) & (g2671)) + ((g2095) & (!g2660) & (g2124) & (!g2264) & (!g3408) & (!g2671)) + ((g2095) & (!g2660) & (g2124) & (!g2264) & (!g3408) & (g2671)) + ((g2095) & (!g2660) & (g2124) & (!g2264) & (g3408) & (!g2671)) + ((g2095) & (!g2660) & (g2124) & (!g2264) & (g3408) & (g2671)) + ((g2095) & (!g2660) & (g2124) & (g2264) & (!g3408) & (!g2671)) + ((g2095) & (!g2660) & (g2124) & (g2264) & (!g3408) & (g2671)) + ((g2095) & (!g2660) & (g2124) & (g2264) & (g3408) & (!g2671)) + ((g2095) & (!g2660) & (g2124) & (g2264) & (g3408) & (g2671)) + ((g2095) & (g2660) & (!g2124) & (!g2264) & (!g3408) & (g2671)) + ((g2095) & (g2660) & (!g2124) & (!g2264) & (g3408) & (g2671)) + ((g2095) & (g2660) & (!g2124) & (g2264) & (g3408) & (!g2671)) + ((g2095) & (g2660) & (!g2124) & (g2264) & (g3408) & (g2671)) + ((g2095) & (g2660) & (g2124) & (!g2264) & (!g3408) & (!g2671)) + ((g2095) & (g2660) & (g2124) & (!g2264) & (!g3408) & (g2671)) + ((g2095) & (g2660) & (g2124) & (!g2264) & (g3408) & (!g2671)) + ((g2095) & (g2660) & (g2124) & (!g2264) & (g3408) & (g2671)));
	assign g2673 = (((!sk[113]) & (!g1050) & (!g2619) & (g1095) & (!g1140)) + ((!sk[113]) & (!g1050) & (!g2619) & (g1095) & (g1140)) + ((!sk[113]) & (!g1050) & (g2619) & (!g1095) & (g1140)) + ((!sk[113]) & (!g1050) & (g2619) & (g1095) & (!g1140)) + ((!sk[113]) & (!g1050) & (g2619) & (g1095) & (g1140)) + ((!sk[113]) & (g1050) & (!g2619) & (!g1095) & (g1140)) + ((!sk[113]) & (g1050) & (!g2619) & (g1095) & (!g1140)) + ((!sk[113]) & (g1050) & (!g2619) & (g1095) & (g1140)) + ((!sk[113]) & (g1050) & (g2619) & (!g1095) & (g1140)) + ((!sk[113]) & (g1050) & (g2619) & (g1095) & (!g1140)) + ((!sk[113]) & (g1050) & (g2619) & (g1095) & (g1140)) + ((sk[113]) & (g1050) & (g2619) & (g1095) & (g1140)));
	assign g2674 = (((!sk[114]) & (!g1185) & (g2673)) + ((!sk[114]) & (g1185) & (g2673)) + ((sk[114]) & (!g1185) & (g2673)) + ((sk[114]) & (g1185) & (!g2673)));
	assign g2675 = (((!g147) & (!sk[115]) & (g1140) & (!g2655)) + ((!g147) & (!sk[115]) & (g1140) & (g2655)) + ((!g147) & (sk[115]) & (g1140) & (g2655)) + ((g147) & (!sk[115]) & (g1140) & (!g2655)) + ((g147) & (!sk[115]) & (g1140) & (g2655)) + ((g147) & (sk[115]) & (!g1140) & (g2655)) + ((g147) & (sk[115]) & (g1140) & (!g2655)) + ((g147) & (sk[115]) & (g1140) & (g2655)));
	assign g2676 = (((!sk[116]) & (!g142) & (!g2585) & (g1185) & (!g2675)) + ((!sk[116]) & (!g142) & (!g2585) & (g1185) & (g2675)) + ((!sk[116]) & (!g142) & (g2585) & (!g1185) & (g2675)) + ((!sk[116]) & (!g142) & (g2585) & (g1185) & (!g2675)) + ((!sk[116]) & (!g142) & (g2585) & (g1185) & (g2675)) + ((!sk[116]) & (g142) & (!g2585) & (!g1185) & (g2675)) + ((!sk[116]) & (g142) & (!g2585) & (g1185) & (!g2675)) + ((!sk[116]) & (g142) & (!g2585) & (g1185) & (g2675)) + ((!sk[116]) & (g142) & (g2585) & (!g1185) & (g2675)) + ((!sk[116]) & (g142) & (g2585) & (g1185) & (!g2675)) + ((!sk[116]) & (g142) & (g2585) & (g1185) & (g2675)) + ((sk[116]) & (!g142) & (g2585) & (!g1185) & (g2675)) + ((sk[116]) & (!g142) & (g2585) & (g1185) & (!g2675)) + ((sk[116]) & (g142) & (g2585) & (!g1185) & (!g2675)) + ((sk[116]) & (g142) & (g2585) & (g1185) & (g2675)));
	assign g5046 = (((!g2921) & (!g3098) & (sk[117]) & (g2677)) + ((!g2921) & (g3098) & (!sk[117]) & (!g2677)) + ((!g2921) & (g3098) & (!sk[117]) & (g2677)) + ((!g2921) & (g3098) & (sk[117]) & (g2677)) + ((g2921) & (g3098) & (!sk[117]) & (!g2677)) + ((g2921) & (g3098) & (!sk[117]) & (g2677)) + ((g2921) & (g3098) & (sk[117]) & (!g2677)) + ((g2921) & (g3098) & (sk[117]) & (g2677)));
	assign g2678 = (((!g1889) & (!sk[118]) & (!g2033) & (g2034) & (!g2677)) + ((!g1889) & (!sk[118]) & (!g2033) & (g2034) & (g2677)) + ((!g1889) & (!sk[118]) & (g2033) & (!g2034) & (g2677)) + ((!g1889) & (!sk[118]) & (g2033) & (g2034) & (!g2677)) + ((!g1889) & (!sk[118]) & (g2033) & (g2034) & (g2677)) + ((!g1889) & (sk[118]) & (!g2033) & (!g2034) & (g2677)) + ((g1889) & (!sk[118]) & (!g2033) & (!g2034) & (g2677)) + ((g1889) & (!sk[118]) & (!g2033) & (g2034) & (!g2677)) + ((g1889) & (!sk[118]) & (!g2033) & (g2034) & (g2677)) + ((g1889) & (!sk[118]) & (g2033) & (!g2034) & (g2677)) + ((g1889) & (!sk[118]) & (g2033) & (g2034) & (!g2677)) + ((g1889) & (!sk[118]) & (g2033) & (g2034) & (g2677)) + ((g1889) & (sk[118]) & (!g2033) & (!g2034) & (g2677)) + ((g1889) & (sk[118]) & (!g2033) & (g2034) & (!g2677)) + ((g1889) & (sk[118]) & (!g2033) & (g2034) & (g2677)));
	assign g2679 = (((g2329) & (!g2029) & (g2408) & (!g2674) & (!g2676) & (g2678)) + ((g2329) & (!g2029) & (g2408) & (!g2674) & (g2676) & (!g2678)) + ((g2329) & (!g2029) & (g2408) & (!g2674) & (g2676) & (g2678)) + ((g2329) & (!g2029) & (g2408) & (g2674) & (!g2676) & (g2678)) + ((g2329) & (!g2029) & (g2408) & (g2674) & (g2676) & (!g2678)) + ((g2329) & (!g2029) & (g2408) & (g2674) & (g2676) & (g2678)) + ((g2329) & (g2029) & (g2408) & (g2674) & (!g2676) & (!g2678)) + ((g2329) & (g2029) & (g2408) & (g2674) & (!g2676) & (g2678)) + ((g2329) & (g2029) & (g2408) & (g2674) & (g2676) & (!g2678)) + ((g2329) & (g2029) & (g2408) & (g2674) & (g2676) & (g2678)));
	assign g2681 = (((!g2094) & (!g2095) & (g2642) & (!g2644) & (g2631) & (g2660)) + ((!g2094) & (!g2095) & (g2642) & (g2644) & (!g2631) & (g2660)) + ((!g2094) & (!g2095) & (g2642) & (g2644) & (g2631) & (g2660)) + ((!g2094) & (g2095) & (!g2642) & (!g2644) & (!g2631) & (g2660)) + ((!g2094) & (g2095) & (!g2642) & (!g2644) & (g2631) & (g2660)) + ((!g2094) & (g2095) & (!g2642) & (g2644) & (!g2631) & (g2660)) + ((!g2094) & (g2095) & (!g2642) & (g2644) & (g2631) & (g2660)) + ((!g2094) & (g2095) & (g2642) & (!g2644) & (!g2631) & (g2660)) + ((!g2094) & (g2095) & (g2642) & (!g2644) & (g2631) & (!g2660)) + ((!g2094) & (g2095) & (g2642) & (!g2644) & (g2631) & (g2660)) + ((!g2094) & (g2095) & (g2642) & (g2644) & (!g2631) & (!g2660)) + ((!g2094) & (g2095) & (g2642) & (g2644) & (!g2631) & (g2660)) + ((!g2094) & (g2095) & (g2642) & (g2644) & (g2631) & (!g2660)) + ((!g2094) & (g2095) & (g2642) & (g2644) & (g2631) & (g2660)) + ((g2094) & (!g2095) & (!g2642) & (!g2644) & (g2631) & (g2660)) + ((g2094) & (!g2095) & (!g2642) & (g2644) & (!g2631) & (g2660)) + ((g2094) & (!g2095) & (!g2642) & (g2644) & (g2631) & (g2660)) + ((g2094) & (!g2095) & (g2642) & (!g2644) & (!g2631) & (g2660)) + ((g2094) & (!g2095) & (g2642) & (!g2644) & (g2631) & (g2660)) + ((g2094) & (!g2095) & (g2642) & (g2644) & (!g2631) & (g2660)) + ((g2094) & (!g2095) & (g2642) & (g2644) & (g2631) & (g2660)) + ((g2094) & (g2095) & (!g2642) & (!g2644) & (!g2631) & (g2660)) + ((g2094) & (g2095) & (!g2642) & (!g2644) & (g2631) & (!g2660)) + ((g2094) & (g2095) & (!g2642) & (!g2644) & (g2631) & (g2660)) + ((g2094) & (g2095) & (!g2642) & (g2644) & (!g2631) & (!g2660)) + ((g2094) & (g2095) & (!g2642) & (g2644) & (!g2631) & (g2660)) + ((g2094) & (g2095) & (!g2642) & (g2644) & (g2631) & (!g2660)) + ((g2094) & (g2095) & (!g2642) & (g2644) & (g2631) & (g2660)) + ((g2094) & (g2095) & (g2642) & (!g2644) & (!g2631) & (!g2660)) + ((g2094) & (g2095) & (g2642) & (!g2644) & (!g2631) & (g2660)) + ((g2094) & (g2095) & (g2642) & (!g2644) & (g2631) & (!g2660)) + ((g2094) & (g2095) & (g2642) & (!g2644) & (g2631) & (g2660)) + ((g2094) & (g2095) & (g2642) & (g2644) & (!g2631) & (!g2660)) + ((g2094) & (g2095) & (g2642) & (g2644) & (!g2631) & (g2660)) + ((g2094) & (g2095) & (g2642) & (g2644) & (g2631) & (!g2660)) + ((g2094) & (g2095) & (g2642) & (g2644) & (g2631) & (g2660)));
	assign g2682 = (((!g2096) & (!sk[121]) & (g2680) & (!g2681)) + ((!g2096) & (!sk[121]) & (g2680) & (g2681)) + ((!g2096) & (sk[121]) & (!g2680) & (g2681)) + ((!g2096) & (sk[121]) & (g2680) & (!g2681)) + ((g2096) & (!sk[121]) & (g2680) & (!g2681)) + ((g2096) & (!sk[121]) & (g2680) & (g2681)) + ((g2096) & (sk[121]) & (!g2680) & (!g2681)) + ((g2096) & (sk[121]) & (g2680) & (g2681)));
	assign g2683 = (((!sk[122]) & (!g2661) & (g2662) & (!g2682)) + ((!sk[122]) & (!g2661) & (g2662) & (g2682)) + ((!sk[122]) & (g2661) & (g2662) & (!g2682)) + ((!sk[122]) & (g2661) & (g2662) & (g2682)) + ((sk[122]) & (!g2661) & (!g2662) & (g2682)) + ((sk[122]) & (!g2661) & (g2662) & (g2682)) + ((sk[122]) & (g2661) & (!g2662) & (g2682)) + ((sk[122]) & (g2661) & (g2662) & (!g2682)));
	assign g2684 = (((!sk[123]) & (!g2660) & (g2095)) + ((!sk[123]) & (g2660) & (g2095)) + ((sk[123]) & (!g2660) & (g2095)));
	assign g2685 = (((!sk[124]) & (!g2680) & (g2096)) + ((!sk[124]) & (g2680) & (g2096)) + ((sk[124]) & (!g2680) & (!g2096)) + ((sk[124]) & (g2680) & (g2096)));
	assign g2686 = (((!g2664) & (!g2665) & (!g2666) & (!g2667) & (!g2684) & (g2685)) + ((!g2664) & (!g2665) & (!g2666) & (!g2667) & (g2684) & (!g2685)) + ((!g2664) & (!g2665) & (!g2666) & (g2667) & (!g2684) & (g2685)) + ((!g2664) & (!g2665) & (!g2666) & (g2667) & (g2684) & (!g2685)) + ((!g2664) & (!g2665) & (g2666) & (!g2667) & (!g2684) & (g2685)) + ((!g2664) & (!g2665) & (g2666) & (!g2667) & (g2684) & (!g2685)) + ((!g2664) & (!g2665) & (g2666) & (g2667) & (!g2684) & (!g2685)) + ((!g2664) & (!g2665) & (g2666) & (g2667) & (g2684) & (g2685)) + ((!g2664) & (g2665) & (!g2666) & (!g2667) & (!g2684) & (g2685)) + ((!g2664) & (g2665) & (!g2666) & (!g2667) & (g2684) & (!g2685)) + ((!g2664) & (g2665) & (!g2666) & (g2667) & (!g2684) & (!g2685)) + ((!g2664) & (g2665) & (!g2666) & (g2667) & (g2684) & (g2685)) + ((!g2664) & (g2665) & (g2666) & (!g2667) & (!g2684) & (!g2685)) + ((!g2664) & (g2665) & (g2666) & (!g2667) & (g2684) & (g2685)) + ((!g2664) & (g2665) & (g2666) & (g2667) & (!g2684) & (!g2685)) + ((!g2664) & (g2665) & (g2666) & (g2667) & (g2684) & (g2685)) + ((g2664) & (!g2665) & (!g2666) & (!g2667) & (!g2684) & (g2685)) + ((g2664) & (!g2665) & (!g2666) & (!g2667) & (g2684) & (!g2685)) + ((g2664) & (!g2665) & (!g2666) & (g2667) & (!g2684) & (!g2685)) + ((g2664) & (!g2665) & (!g2666) & (g2667) & (g2684) & (g2685)) + ((g2664) & (!g2665) & (g2666) & (!g2667) & (!g2684) & (!g2685)) + ((g2664) & (!g2665) & (g2666) & (!g2667) & (g2684) & (g2685)) + ((g2664) & (!g2665) & (g2666) & (g2667) & (!g2684) & (!g2685)) + ((g2664) & (!g2665) & (g2666) & (g2667) & (g2684) & (g2685)) + ((g2664) & (g2665) & (!g2666) & (!g2667) & (!g2684) & (g2685)) + ((g2664) & (g2665) & (!g2666) & (!g2667) & (g2684) & (!g2685)) + ((g2664) & (g2665) & (!g2666) & (g2667) & (!g2684) & (!g2685)) + ((g2664) & (g2665) & (!g2666) & (g2667) & (g2684) & (g2685)) + ((g2664) & (g2665) & (g2666) & (!g2667) & (!g2684) & (!g2685)) + ((g2664) & (g2665) & (g2666) & (!g2667) & (g2684) & (g2685)) + ((g2664) & (g2665) & (g2666) & (g2667) & (!g2684) & (!g2685)) + ((g2664) & (g2665) & (g2666) & (g2667) & (g2684) & (g2685)));
	assign g2687 = (((!g2096) & (!g2095) & (!g2094) & (g2093) & (g2071) & (g2074)) + ((!g2096) & (!g2095) & (g2094) & (!g2093) & (!g2071) & (g2074)) + ((!g2096) & (!g2095) & (g2094) & (g2093) & (!g2071) & (g2074)) + ((!g2096) & (!g2095) & (g2094) & (g2093) & (g2071) & (g2074)) + ((!g2096) & (g2095) & (!g2094) & (!g2093) & (g2071) & (!g2074)) + ((!g2096) & (g2095) & (!g2094) & (g2093) & (g2071) & (!g2074)) + ((!g2096) & (g2095) & (!g2094) & (g2093) & (g2071) & (g2074)) + ((!g2096) & (g2095) & (g2094) & (!g2093) & (!g2071) & (g2074)) + ((!g2096) & (g2095) & (g2094) & (!g2093) & (g2071) & (!g2074)) + ((!g2096) & (g2095) & (g2094) & (g2093) & (!g2071) & (g2074)) + ((!g2096) & (g2095) & (g2094) & (g2093) & (g2071) & (!g2074)) + ((!g2096) & (g2095) & (g2094) & (g2093) & (g2071) & (g2074)) + ((g2096) & (!g2095) & (!g2094) & (!g2093) & (!g2071) & (!g2074)) + ((g2096) & (!g2095) & (!g2094) & (g2093) & (!g2071) & (!g2074)) + ((g2096) & (!g2095) & (!g2094) & (g2093) & (g2071) & (g2074)) + ((g2096) & (!g2095) & (g2094) & (!g2093) & (!g2071) & (!g2074)) + ((g2096) & (!g2095) & (g2094) & (!g2093) & (!g2071) & (g2074)) + ((g2096) & (!g2095) & (g2094) & (g2093) & (!g2071) & (!g2074)) + ((g2096) & (!g2095) & (g2094) & (g2093) & (!g2071) & (g2074)) + ((g2096) & (!g2095) & (g2094) & (g2093) & (g2071) & (g2074)) + ((g2096) & (g2095) & (!g2094) & (!g2093) & (!g2071) & (!g2074)) + ((g2096) & (g2095) & (!g2094) & (!g2093) & (g2071) & (!g2074)) + ((g2096) & (g2095) & (!g2094) & (g2093) & (!g2071) & (!g2074)) + ((g2096) & (g2095) & (!g2094) & (g2093) & (g2071) & (!g2074)) + ((g2096) & (g2095) & (!g2094) & (g2093) & (g2071) & (g2074)) + ((g2096) & (g2095) & (g2094) & (!g2093) & (!g2071) & (!g2074)) + ((g2096) & (g2095) & (g2094) & (!g2093) & (!g2071) & (g2074)) + ((g2096) & (g2095) & (g2094) & (!g2093) & (g2071) & (!g2074)) + ((g2096) & (g2095) & (g2094) & (g2093) & (!g2071) & (!g2074)) + ((g2096) & (g2095) & (g2094) & (g2093) & (!g2071) & (g2074)) + ((g2096) & (g2095) & (g2094) & (g2093) & (g2071) & (!g2074)) + ((g2096) & (g2095) & (g2094) & (g2093) & (g2071) & (g2074)));
	assign g2688 = (((!g2687) & (!g2536) & (!g2615) & (g2449) & (g2076) & (g2077)) + ((!g2687) & (!g2536) & (g2615) & (!g2449) & (!g2076) & (g2077)) + ((!g2687) & (!g2536) & (g2615) & (g2449) & (!g2076) & (g2077)) + ((!g2687) & (!g2536) & (g2615) & (g2449) & (g2076) & (g2077)) + ((!g2687) & (g2536) & (!g2615) & (!g2449) & (g2076) & (!g2077)) + ((!g2687) & (g2536) & (!g2615) & (g2449) & (g2076) & (!g2077)) + ((!g2687) & (g2536) & (!g2615) & (g2449) & (g2076) & (g2077)) + ((!g2687) & (g2536) & (g2615) & (!g2449) & (!g2076) & (g2077)) + ((!g2687) & (g2536) & (g2615) & (!g2449) & (g2076) & (!g2077)) + ((!g2687) & (g2536) & (g2615) & (g2449) & (!g2076) & (g2077)) + ((!g2687) & (g2536) & (g2615) & (g2449) & (g2076) & (!g2077)) + ((!g2687) & (g2536) & (g2615) & (g2449) & (g2076) & (g2077)) + ((g2687) & (!g2536) & (!g2615) & (!g2449) & (!g2076) & (!g2077)) + ((g2687) & (!g2536) & (!g2615) & (g2449) & (!g2076) & (!g2077)) + ((g2687) & (!g2536) & (!g2615) & (g2449) & (g2076) & (g2077)) + ((g2687) & (!g2536) & (g2615) & (!g2449) & (!g2076) & (!g2077)) + ((g2687) & (!g2536) & (g2615) & (!g2449) & (!g2076) & (g2077)) + ((g2687) & (!g2536) & (g2615) & (g2449) & (!g2076) & (!g2077)) + ((g2687) & (!g2536) & (g2615) & (g2449) & (!g2076) & (g2077)) + ((g2687) & (!g2536) & (g2615) & (g2449) & (g2076) & (g2077)) + ((g2687) & (g2536) & (!g2615) & (!g2449) & (!g2076) & (!g2077)) + ((g2687) & (g2536) & (!g2615) & (!g2449) & (g2076) & (!g2077)) + ((g2687) & (g2536) & (!g2615) & (g2449) & (!g2076) & (!g2077)) + ((g2687) & (g2536) & (!g2615) & (g2449) & (g2076) & (!g2077)) + ((g2687) & (g2536) & (!g2615) & (g2449) & (g2076) & (g2077)) + ((g2687) & (g2536) & (g2615) & (!g2449) & (!g2076) & (!g2077)) + ((g2687) & (g2536) & (g2615) & (!g2449) & (!g2076) & (g2077)) + ((g2687) & (g2536) & (g2615) & (!g2449) & (g2076) & (!g2077)) + ((g2687) & (g2536) & (g2615) & (g2449) & (!g2076) & (!g2077)) + ((g2687) & (g2536) & (g2615) & (g2449) & (!g2076) & (g2077)) + ((g2687) & (g2536) & (g2615) & (g2449) & (g2076) & (!g2077)) + ((g2687) & (g2536) & (g2615) & (g2449) & (g2076) & (g2077)));
	assign g2689 = (((!g2688) & (!g2351) & (!g2353) & (g2191) & (g2073) & (g2125)) + ((!g2688) & (!g2351) & (g2353) & (!g2191) & (!g2073) & (g2125)) + ((!g2688) & (!g2351) & (g2353) & (g2191) & (!g2073) & (g2125)) + ((!g2688) & (!g2351) & (g2353) & (g2191) & (g2073) & (g2125)) + ((!g2688) & (g2351) & (!g2353) & (!g2191) & (g2073) & (!g2125)) + ((!g2688) & (g2351) & (!g2353) & (g2191) & (g2073) & (!g2125)) + ((!g2688) & (g2351) & (!g2353) & (g2191) & (g2073) & (g2125)) + ((!g2688) & (g2351) & (g2353) & (!g2191) & (!g2073) & (g2125)) + ((!g2688) & (g2351) & (g2353) & (!g2191) & (g2073) & (!g2125)) + ((!g2688) & (g2351) & (g2353) & (g2191) & (!g2073) & (g2125)) + ((!g2688) & (g2351) & (g2353) & (g2191) & (g2073) & (!g2125)) + ((!g2688) & (g2351) & (g2353) & (g2191) & (g2073) & (g2125)) + ((g2688) & (!g2351) & (!g2353) & (!g2191) & (!g2073) & (!g2125)) + ((g2688) & (!g2351) & (!g2353) & (g2191) & (!g2073) & (!g2125)) + ((g2688) & (!g2351) & (!g2353) & (g2191) & (g2073) & (g2125)) + ((g2688) & (!g2351) & (g2353) & (!g2191) & (!g2073) & (!g2125)) + ((g2688) & (!g2351) & (g2353) & (!g2191) & (!g2073) & (g2125)) + ((g2688) & (!g2351) & (g2353) & (g2191) & (!g2073) & (!g2125)) + ((g2688) & (!g2351) & (g2353) & (g2191) & (!g2073) & (g2125)) + ((g2688) & (!g2351) & (g2353) & (g2191) & (g2073) & (g2125)) + ((g2688) & (g2351) & (!g2353) & (!g2191) & (!g2073) & (!g2125)) + ((g2688) & (g2351) & (!g2353) & (!g2191) & (g2073) & (!g2125)) + ((g2688) & (g2351) & (!g2353) & (g2191) & (!g2073) & (!g2125)) + ((g2688) & (g2351) & (!g2353) & (g2191) & (g2073) & (!g2125)) + ((g2688) & (g2351) & (!g2353) & (g2191) & (g2073) & (g2125)) + ((g2688) & (g2351) & (g2353) & (!g2191) & (!g2073) & (!g2125)) + ((g2688) & (g2351) & (g2353) & (!g2191) & (!g2073) & (g2125)) + ((g2688) & (g2351) & (g2353) & (!g2191) & (g2073) & (!g2125)) + ((g2688) & (g2351) & (g2353) & (g2191) & (!g2073) & (!g2125)) + ((g2688) & (g2351) & (g2353) & (g2191) & (!g2073) & (g2125)) + ((g2688) & (g2351) & (g2353) & (g2191) & (g2073) & (!g2125)) + ((g2688) & (g2351) & (g2353) & (g2191) & (g2073) & (g2125)));
	assign g2690 = (((!g2096) & (!g2680) & (!g2124) & (!g2264) & (!g3384) & (g2689)) + ((!g2096) & (!g2680) & (!g2124) & (!g2264) & (g3384) & (g2689)) + ((!g2096) & (!g2680) & (!g2124) & (g2264) & (g3384) & (!g2689)) + ((!g2096) & (!g2680) & (!g2124) & (g2264) & (g3384) & (g2689)) + ((!g2096) & (g2680) & (!g2124) & (!g2264) & (!g3384) & (g2689)) + ((!g2096) & (g2680) & (!g2124) & (!g2264) & (g3384) & (g2689)) + ((!g2096) & (g2680) & (!g2124) & (g2264) & (g3384) & (!g2689)) + ((!g2096) & (g2680) & (!g2124) & (g2264) & (g3384) & (g2689)) + ((!g2096) & (g2680) & (g2124) & (!g2264) & (!g3384) & (!g2689)) + ((!g2096) & (g2680) & (g2124) & (!g2264) & (!g3384) & (g2689)) + ((!g2096) & (g2680) & (g2124) & (!g2264) & (g3384) & (!g2689)) + ((!g2096) & (g2680) & (g2124) & (!g2264) & (g3384) & (g2689)) + ((!g2096) & (g2680) & (g2124) & (g2264) & (!g3384) & (!g2689)) + ((!g2096) & (g2680) & (g2124) & (g2264) & (!g3384) & (g2689)) + ((!g2096) & (g2680) & (g2124) & (g2264) & (g3384) & (!g2689)) + ((!g2096) & (g2680) & (g2124) & (g2264) & (g3384) & (g2689)) + ((g2096) & (!g2680) & (!g2124) & (!g2264) & (!g3384) & (g2689)) + ((g2096) & (!g2680) & (!g2124) & (!g2264) & (g3384) & (g2689)) + ((g2096) & (!g2680) & (!g2124) & (g2264) & (g3384) & (!g2689)) + ((g2096) & (!g2680) & (!g2124) & (g2264) & (g3384) & (g2689)) + ((g2096) & (!g2680) & (g2124) & (!g2264) & (!g3384) & (!g2689)) + ((g2096) & (!g2680) & (g2124) & (!g2264) & (!g3384) & (g2689)) + ((g2096) & (!g2680) & (g2124) & (!g2264) & (g3384) & (!g2689)) + ((g2096) & (!g2680) & (g2124) & (!g2264) & (g3384) & (g2689)) + ((g2096) & (!g2680) & (g2124) & (g2264) & (!g3384) & (!g2689)) + ((g2096) & (!g2680) & (g2124) & (g2264) & (!g3384) & (g2689)) + ((g2096) & (!g2680) & (g2124) & (g2264) & (g3384) & (!g2689)) + ((g2096) & (!g2680) & (g2124) & (g2264) & (g3384) & (g2689)) + ((g2096) & (g2680) & (!g2124) & (!g2264) & (!g3384) & (g2689)) + ((g2096) & (g2680) & (!g2124) & (!g2264) & (g3384) & (g2689)) + ((g2096) & (g2680) & (!g2124) & (g2264) & (g3384) & (!g2689)) + ((g2096) & (g2680) & (!g2124) & (g2264) & (g3384) & (g2689)) + ((g2096) & (g2680) & (g2124) & (!g2264) & (!g3384) & (!g2689)) + ((g2096) & (g2680) & (g2124) & (!g2264) & (!g3384) & (g2689)) + ((g2096) & (g2680) & (g2124) & (!g2264) & (g3384) & (!g2689)) + ((g2096) & (g2680) & (g2124) & (!g2264) & (g3384) & (g2689)));
	assign g2691 = (((!g1185) & (!sk[2]) & (g2673) & (!g1230)) + ((!g1185) & (!sk[2]) & (g2673) & (g1230)) + ((!g1185) & (sk[2]) & (!g2673) & (g1230)) + ((!g1185) & (sk[2]) & (g2673) & (g1230)) + ((g1185) & (!sk[2]) & (g2673) & (!g1230)) + ((g1185) & (!sk[2]) & (g2673) & (g1230)) + ((g1185) & (sk[2]) & (!g2673) & (g1230)) + ((g1185) & (sk[2]) & (g2673) & (!g1230)));
	assign g2692 = (((!g142) & (!sk[3]) & (g1185)) + ((!g142) & (sk[3]) & (g1185)) + ((g142) & (!sk[3]) & (g1185)) + ((g142) & (sk[3]) & (!g1185)));
	assign g2693 = (((!g147) & (!g148) & (g1095) & (!g2637) & (g1140) & (g2692)) + ((!g147) & (g148) & (!g1095) & (!g2637) & (g1140) & (g2692)) + ((!g147) & (g148) & (g1095) & (!g2637) & (g1140) & (g2692)) + ((!g147) & (g148) & (g1095) & (g2637) & (g1140) & (g2692)) + ((g147) & (!g148) & (!g1095) & (!g2637) & (g1140) & (g2692)) + ((g147) & (!g148) & (!g1095) & (g2637) & (g1140) & (g2692)) + ((g147) & (!g148) & (g1095) & (!g2637) & (!g1140) & (g2692)) + ((g147) & (!g148) & (g1095) & (!g2637) & (g1140) & (g2692)) + ((g147) & (!g148) & (g1095) & (g2637) & (g1140) & (g2692)) + ((g147) & (g148) & (!g1095) & (!g2637) & (!g1140) & (g2692)) + ((g147) & (g148) & (!g1095) & (!g2637) & (g1140) & (g2692)) + ((g147) & (g148) & (!g1095) & (g2637) & (g1140) & (g2692)) + ((g147) & (g148) & (g1095) & (!g2637) & (!g1140) & (g2692)) + ((g147) & (g148) & (g1095) & (!g2637) & (g1140) & (g2692)) + ((g147) & (g148) & (g1095) & (g2637) & (!g1140) & (g2692)) + ((g147) & (g148) & (g1095) & (g2637) & (g1140) & (g2692)));
	assign g2694 = (((!g142) & (!sk[5]) & (g1185)) + ((g142) & (!sk[5]) & (g1185)) + ((g142) & (sk[5]) & (g1185)));
	assign g2695 = (((!g678) & (!g2585) & (!g1230) & (!sk[6]) & (g2693) & (!g2694)) + ((!g678) & (!g2585) & (!g1230) & (!sk[6]) & (g2693) & (g2694)) + ((!g678) & (!g2585) & (g1230) & (!sk[6]) & (g2693) & (!g2694)) + ((!g678) & (!g2585) & (g1230) & (!sk[6]) & (g2693) & (g2694)) + ((!g678) & (g2585) & (!g1230) & (!sk[6]) & (!g2693) & (!g2694)) + ((!g678) & (g2585) & (!g1230) & (!sk[6]) & (!g2693) & (g2694)) + ((!g678) & (g2585) & (!g1230) & (!sk[6]) & (g2693) & (!g2694)) + ((!g678) & (g2585) & (!g1230) & (!sk[6]) & (g2693) & (g2694)) + ((!g678) & (g2585) & (!g1230) & (sk[6]) & (!g2693) & (g2694)) + ((!g678) & (g2585) & (!g1230) & (sk[6]) & (g2693) & (!g2694)) + ((!g678) & (g2585) & (!g1230) & (sk[6]) & (g2693) & (g2694)) + ((!g678) & (g2585) & (g1230) & (!sk[6]) & (!g2693) & (!g2694)) + ((!g678) & (g2585) & (g1230) & (!sk[6]) & (!g2693) & (g2694)) + ((!g678) & (g2585) & (g1230) & (!sk[6]) & (g2693) & (!g2694)) + ((!g678) & (g2585) & (g1230) & (!sk[6]) & (g2693) & (g2694)) + ((!g678) & (g2585) & (g1230) & (sk[6]) & (!g2693) & (!g2694)) + ((g678) & (!g2585) & (!g1230) & (!sk[6]) & (g2693) & (!g2694)) + ((g678) & (!g2585) & (!g1230) & (!sk[6]) & (g2693) & (g2694)) + ((g678) & (!g2585) & (g1230) & (!sk[6]) & (g2693) & (!g2694)) + ((g678) & (!g2585) & (g1230) & (!sk[6]) & (g2693) & (g2694)) + ((g678) & (g2585) & (!g1230) & (!sk[6]) & (!g2693) & (!g2694)) + ((g678) & (g2585) & (!g1230) & (!sk[6]) & (!g2693) & (g2694)) + ((g678) & (g2585) & (!g1230) & (!sk[6]) & (g2693) & (!g2694)) + ((g678) & (g2585) & (!g1230) & (!sk[6]) & (g2693) & (g2694)) + ((g678) & (g2585) & (!g1230) & (sk[6]) & (!g2693) & (!g2694)) + ((g678) & (g2585) & (g1230) & (!sk[6]) & (!g2693) & (!g2694)) + ((g678) & (g2585) & (g1230) & (!sk[6]) & (!g2693) & (g2694)) + ((g678) & (g2585) & (g1230) & (!sk[6]) & (g2693) & (!g2694)) + ((g678) & (g2585) & (g1230) & (!sk[6]) & (g2693) & (g2694)) + ((g678) & (g2585) & (g1230) & (sk[6]) & (!g2693) & (g2694)) + ((g678) & (g2585) & (g1230) & (sk[6]) & (g2693) & (!g2694)) + ((g678) & (g2585) & (g1230) & (sk[6]) & (g2693) & (g2694)));
	assign g5047 = (((!g2921) & (!g3174) & (sk[7]) & (g2696)) + ((!g2921) & (g3174) & (!sk[7]) & (!g2696)) + ((!g2921) & (g3174) & (!sk[7]) & (g2696)) + ((!g2921) & (g3174) & (sk[7]) & (g2696)) + ((g2921) & (g3174) & (!sk[7]) & (!g2696)) + ((g2921) & (g3174) & (!sk[7]) & (g2696)) + ((g2921) & (g3174) & (sk[7]) & (!g2696)) + ((g2921) & (g3174) & (sk[7]) & (g2696)));
	assign g2697 = (((!g1902) & (!g2033) & (!sk[8]) & (g2034) & (!g2696)) + ((!g1902) & (!g2033) & (!sk[8]) & (g2034) & (g2696)) + ((!g1902) & (!g2033) & (sk[8]) & (!g2034) & (g2696)) + ((!g1902) & (g2033) & (!sk[8]) & (!g2034) & (g2696)) + ((!g1902) & (g2033) & (!sk[8]) & (g2034) & (!g2696)) + ((!g1902) & (g2033) & (!sk[8]) & (g2034) & (g2696)) + ((g1902) & (!g2033) & (!sk[8]) & (!g2034) & (g2696)) + ((g1902) & (!g2033) & (!sk[8]) & (g2034) & (!g2696)) + ((g1902) & (!g2033) & (!sk[8]) & (g2034) & (g2696)) + ((g1902) & (!g2033) & (sk[8]) & (!g2034) & (g2696)) + ((g1902) & (!g2033) & (sk[8]) & (g2034) & (!g2696)) + ((g1902) & (!g2033) & (sk[8]) & (g2034) & (g2696)) + ((g1902) & (g2033) & (!sk[8]) & (!g2034) & (g2696)) + ((g1902) & (g2033) & (!sk[8]) & (g2034) & (!g2696)) + ((g1902) & (g2033) & (!sk[8]) & (g2034) & (g2696)));
	assign g2698 = (((g2329) & (!g2029) & (g2408) & (!g2691) & (!g2695) & (g2697)) + ((g2329) & (!g2029) & (g2408) & (!g2691) & (g2695) & (!g2697)) + ((g2329) & (!g2029) & (g2408) & (!g2691) & (g2695) & (g2697)) + ((g2329) & (!g2029) & (g2408) & (g2691) & (!g2695) & (g2697)) + ((g2329) & (!g2029) & (g2408) & (g2691) & (g2695) & (!g2697)) + ((g2329) & (!g2029) & (g2408) & (g2691) & (g2695) & (g2697)) + ((g2329) & (g2029) & (g2408) & (g2691) & (!g2695) & (!g2697)) + ((g2329) & (g2029) & (g2408) & (g2691) & (!g2695) & (g2697)) + ((g2329) & (g2029) & (g2408) & (g2691) & (g2695) & (!g2697)) + ((g2329) & (g2029) & (g2408) & (g2691) & (g2695) & (g2697)));
	assign g2700 = (((!g2088) & (!g2096) & (!g2680) & (!sk[10]) & (g2681) & (!g2699)) + ((!g2088) & (!g2096) & (!g2680) & (!sk[10]) & (g2681) & (g2699)) + ((!g2088) & (!g2096) & (!g2680) & (sk[10]) & (!g2681) & (g2699)) + ((!g2088) & (!g2096) & (!g2680) & (sk[10]) & (g2681) & (g2699)) + ((!g2088) & (!g2096) & (g2680) & (!sk[10]) & (g2681) & (!g2699)) + ((!g2088) & (!g2096) & (g2680) & (!sk[10]) & (g2681) & (g2699)) + ((!g2088) & (!g2096) & (g2680) & (sk[10]) & (!g2681) & (g2699)) + ((!g2088) & (!g2096) & (g2680) & (sk[10]) & (g2681) & (!g2699)) + ((!g2088) & (g2096) & (!g2680) & (!sk[10]) & (!g2681) & (!g2699)) + ((!g2088) & (g2096) & (!g2680) & (!sk[10]) & (!g2681) & (g2699)) + ((!g2088) & (g2096) & (!g2680) & (!sk[10]) & (g2681) & (!g2699)) + ((!g2088) & (g2096) & (!g2680) & (!sk[10]) & (g2681) & (g2699)) + ((!g2088) & (g2096) & (!g2680) & (sk[10]) & (!g2681) & (g2699)) + ((!g2088) & (g2096) & (!g2680) & (sk[10]) & (g2681) & (!g2699)) + ((!g2088) & (g2096) & (g2680) & (!sk[10]) & (!g2681) & (!g2699)) + ((!g2088) & (g2096) & (g2680) & (!sk[10]) & (!g2681) & (g2699)) + ((!g2088) & (g2096) & (g2680) & (!sk[10]) & (g2681) & (!g2699)) + ((!g2088) & (g2096) & (g2680) & (!sk[10]) & (g2681) & (g2699)) + ((!g2088) & (g2096) & (g2680) & (sk[10]) & (!g2681) & (!g2699)) + ((!g2088) & (g2096) & (g2680) & (sk[10]) & (g2681) & (!g2699)) + ((g2088) & (!g2096) & (!g2680) & (!sk[10]) & (g2681) & (!g2699)) + ((g2088) & (!g2096) & (!g2680) & (!sk[10]) & (g2681) & (g2699)) + ((g2088) & (!g2096) & (!g2680) & (sk[10]) & (!g2681) & (!g2699)) + ((g2088) & (!g2096) & (!g2680) & (sk[10]) & (g2681) & (!g2699)) + ((g2088) & (!g2096) & (g2680) & (!sk[10]) & (g2681) & (!g2699)) + ((g2088) & (!g2096) & (g2680) & (!sk[10]) & (g2681) & (g2699)) + ((g2088) & (!g2096) & (g2680) & (sk[10]) & (!g2681) & (!g2699)) + ((g2088) & (!g2096) & (g2680) & (sk[10]) & (g2681) & (g2699)) + ((g2088) & (g2096) & (!g2680) & (!sk[10]) & (!g2681) & (!g2699)) + ((g2088) & (g2096) & (!g2680) & (!sk[10]) & (!g2681) & (g2699)) + ((g2088) & (g2096) & (!g2680) & (!sk[10]) & (g2681) & (!g2699)) + ((g2088) & (g2096) & (!g2680) & (!sk[10]) & (g2681) & (g2699)) + ((g2088) & (g2096) & (!g2680) & (sk[10]) & (!g2681) & (!g2699)) + ((g2088) & (g2096) & (!g2680) & (sk[10]) & (g2681) & (g2699)) + ((g2088) & (g2096) & (g2680) & (!sk[10]) & (!g2681) & (!g2699)) + ((g2088) & (g2096) & (g2680) & (!sk[10]) & (!g2681) & (g2699)) + ((g2088) & (g2096) & (g2680) & (!sk[10]) & (g2681) & (!g2699)) + ((g2088) & (g2096) & (g2680) & (!sk[10]) & (g2681) & (g2699)) + ((g2088) & (g2096) & (g2680) & (sk[10]) & (!g2681) & (g2699)) + ((g2088) & (g2096) & (g2680) & (sk[10]) & (g2681) & (g2699)));
	assign g2701 = (((!g2661) & (!g2662) & (!g2682) & (sk[11]) & (g2700)) + ((!g2661) & (!g2662) & (g2682) & (!sk[11]) & (!g2700)) + ((!g2661) & (!g2662) & (g2682) & (!sk[11]) & (g2700)) + ((!g2661) & (!g2662) & (g2682) & (sk[11]) & (g2700)) + ((!g2661) & (g2662) & (!g2682) & (!sk[11]) & (g2700)) + ((!g2661) & (g2662) & (!g2682) & (sk[11]) & (g2700)) + ((!g2661) & (g2662) & (g2682) & (!sk[11]) & (!g2700)) + ((!g2661) & (g2662) & (g2682) & (!sk[11]) & (g2700)) + ((!g2661) & (g2662) & (g2682) & (sk[11]) & (g2700)) + ((g2661) & (!g2662) & (!g2682) & (!sk[11]) & (g2700)) + ((g2661) & (!g2662) & (!g2682) & (sk[11]) & (g2700)) + ((g2661) & (!g2662) & (g2682) & (!sk[11]) & (!g2700)) + ((g2661) & (!g2662) & (g2682) & (!sk[11]) & (g2700)) + ((g2661) & (!g2662) & (g2682) & (sk[11]) & (g2700)) + ((g2661) & (g2662) & (!g2682) & (!sk[11]) & (g2700)) + ((g2661) & (g2662) & (!g2682) & (sk[11]) & (g2700)) + ((g2661) & (g2662) & (g2682) & (!sk[11]) & (!g2700)) + ((g2661) & (g2662) & (g2682) & (!sk[11]) & (g2700)) + ((g2661) & (g2662) & (g2682) & (sk[11]) & (!g2700)));
	assign g2702 = (((!g2664) & (!g2665) & (!g2666) & (!g2667) & (!g2684) & (!g2685)) + ((!g2664) & (!g2665) & (!g2666) & (!g2667) & (!g2684) & (g2685)) + ((!g2664) & (!g2665) & (!g2666) & (!g2667) & (g2684) & (!g2685)) + ((!g2664) & (!g2665) & (!g2666) & (g2667) & (!g2684) & (!g2685)) + ((!g2664) & (!g2665) & (!g2666) & (g2667) & (!g2684) & (g2685)) + ((!g2664) & (!g2665) & (!g2666) & (g2667) & (g2684) & (!g2685)) + ((!g2664) & (!g2665) & (g2666) & (!g2667) & (!g2684) & (!g2685)) + ((!g2664) & (!g2665) & (g2666) & (!g2667) & (!g2684) & (g2685)) + ((!g2664) & (!g2665) & (g2666) & (!g2667) & (g2684) & (!g2685)) + ((!g2664) & (!g2665) & (g2666) & (g2667) & (!g2684) & (!g2685)) + ((!g2664) & (g2665) & (!g2666) & (!g2667) & (!g2684) & (!g2685)) + ((!g2664) & (g2665) & (!g2666) & (!g2667) & (!g2684) & (g2685)) + ((!g2664) & (g2665) & (!g2666) & (!g2667) & (g2684) & (!g2685)) + ((!g2664) & (g2665) & (!g2666) & (g2667) & (!g2684) & (!g2685)) + ((!g2664) & (g2665) & (g2666) & (!g2667) & (!g2684) & (!g2685)) + ((!g2664) & (g2665) & (g2666) & (g2667) & (!g2684) & (!g2685)) + ((g2664) & (!g2665) & (!g2666) & (!g2667) & (!g2684) & (!g2685)) + ((g2664) & (!g2665) & (!g2666) & (!g2667) & (!g2684) & (g2685)) + ((g2664) & (!g2665) & (!g2666) & (!g2667) & (g2684) & (!g2685)) + ((g2664) & (!g2665) & (!g2666) & (g2667) & (!g2684) & (!g2685)) + ((g2664) & (!g2665) & (g2666) & (!g2667) & (!g2684) & (!g2685)) + ((g2664) & (!g2665) & (g2666) & (g2667) & (!g2684) & (!g2685)) + ((g2664) & (g2665) & (!g2666) & (!g2667) & (!g2684) & (!g2685)) + ((g2664) & (g2665) & (!g2666) & (!g2667) & (!g2684) & (g2685)) + ((g2664) & (g2665) & (!g2666) & (!g2667) & (g2684) & (!g2685)) + ((g2664) & (g2665) & (!g2666) & (g2667) & (!g2684) & (!g2685)) + ((g2664) & (g2665) & (g2666) & (!g2667) & (!g2684) & (!g2685)) + ((g2664) & (g2665) & (g2666) & (g2667) & (!g2684) & (!g2685)));
	assign g2703 = (((!g2680) & (!sk[13]) & (g2096)) + ((!g2680) & (sk[13]) & (g2096)) + ((g2680) & (!sk[13]) & (g2096)));
	assign g2704 = (((!sk[14]) & (!g2699) & (g2088)) + ((!sk[14]) & (g2699) & (g2088)) + ((sk[14]) & (!g2699) & (!g2088)) + ((sk[14]) & (g2699) & (g2088)));
	assign g2705 = (((!sk[15]) & (!g2702) & (g2703) & (!g2704)) + ((!sk[15]) & (!g2702) & (g2703) & (g2704)) + ((!sk[15]) & (g2702) & (g2703) & (!g2704)) + ((!sk[15]) & (g2702) & (g2703) & (g2704)) + ((sk[15]) & (!g2702) & (!g2703) & (!g2704)) + ((sk[15]) & (!g2702) & (g2703) & (g2704)) + ((sk[15]) & (g2702) & (!g2703) & (g2704)) + ((sk[15]) & (g2702) & (g2703) & (!g2704)));
	assign g2706 = (((!g2088) & (!g2096) & (!g2095) & (g2094) & (g2071) & (g2074)) + ((!g2088) & (!g2096) & (g2095) & (!g2094) & (!g2071) & (g2074)) + ((!g2088) & (!g2096) & (g2095) & (g2094) & (!g2071) & (g2074)) + ((!g2088) & (!g2096) & (g2095) & (g2094) & (g2071) & (g2074)) + ((!g2088) & (g2096) & (!g2095) & (!g2094) & (g2071) & (!g2074)) + ((!g2088) & (g2096) & (!g2095) & (g2094) & (g2071) & (!g2074)) + ((!g2088) & (g2096) & (!g2095) & (g2094) & (g2071) & (g2074)) + ((!g2088) & (g2096) & (g2095) & (!g2094) & (!g2071) & (g2074)) + ((!g2088) & (g2096) & (g2095) & (!g2094) & (g2071) & (!g2074)) + ((!g2088) & (g2096) & (g2095) & (g2094) & (!g2071) & (g2074)) + ((!g2088) & (g2096) & (g2095) & (g2094) & (g2071) & (!g2074)) + ((!g2088) & (g2096) & (g2095) & (g2094) & (g2071) & (g2074)) + ((g2088) & (!g2096) & (!g2095) & (!g2094) & (!g2071) & (!g2074)) + ((g2088) & (!g2096) & (!g2095) & (g2094) & (!g2071) & (!g2074)) + ((g2088) & (!g2096) & (!g2095) & (g2094) & (g2071) & (g2074)) + ((g2088) & (!g2096) & (g2095) & (!g2094) & (!g2071) & (!g2074)) + ((g2088) & (!g2096) & (g2095) & (!g2094) & (!g2071) & (g2074)) + ((g2088) & (!g2096) & (g2095) & (g2094) & (!g2071) & (!g2074)) + ((g2088) & (!g2096) & (g2095) & (g2094) & (!g2071) & (g2074)) + ((g2088) & (!g2096) & (g2095) & (g2094) & (g2071) & (g2074)) + ((g2088) & (g2096) & (!g2095) & (!g2094) & (!g2071) & (!g2074)) + ((g2088) & (g2096) & (!g2095) & (!g2094) & (g2071) & (!g2074)) + ((g2088) & (g2096) & (!g2095) & (g2094) & (!g2071) & (!g2074)) + ((g2088) & (g2096) & (!g2095) & (g2094) & (g2071) & (!g2074)) + ((g2088) & (g2096) & (!g2095) & (g2094) & (g2071) & (g2074)) + ((g2088) & (g2096) & (g2095) & (!g2094) & (!g2071) & (!g2074)) + ((g2088) & (g2096) & (g2095) & (!g2094) & (!g2071) & (g2074)) + ((g2088) & (g2096) & (g2095) & (!g2094) & (g2071) & (!g2074)) + ((g2088) & (g2096) & (g2095) & (g2094) & (!g2071) & (!g2074)) + ((g2088) & (g2096) & (g2095) & (g2094) & (!g2071) & (g2074)) + ((g2088) & (g2096) & (g2095) & (g2094) & (g2071) & (!g2074)) + ((g2088) & (g2096) & (g2095) & (g2094) & (g2071) & (g2074)));
	assign g2707 = (((!g2706) & (!g2559) & (!g2632) & (g2467) & (g2076) & (g2077)) + ((!g2706) & (!g2559) & (g2632) & (!g2467) & (!g2076) & (g2077)) + ((!g2706) & (!g2559) & (g2632) & (g2467) & (!g2076) & (g2077)) + ((!g2706) & (!g2559) & (g2632) & (g2467) & (g2076) & (g2077)) + ((!g2706) & (g2559) & (!g2632) & (!g2467) & (g2076) & (!g2077)) + ((!g2706) & (g2559) & (!g2632) & (g2467) & (g2076) & (!g2077)) + ((!g2706) & (g2559) & (!g2632) & (g2467) & (g2076) & (g2077)) + ((!g2706) & (g2559) & (g2632) & (!g2467) & (!g2076) & (g2077)) + ((!g2706) & (g2559) & (g2632) & (!g2467) & (g2076) & (!g2077)) + ((!g2706) & (g2559) & (g2632) & (g2467) & (!g2076) & (g2077)) + ((!g2706) & (g2559) & (g2632) & (g2467) & (g2076) & (!g2077)) + ((!g2706) & (g2559) & (g2632) & (g2467) & (g2076) & (g2077)) + ((g2706) & (!g2559) & (!g2632) & (!g2467) & (!g2076) & (!g2077)) + ((g2706) & (!g2559) & (!g2632) & (g2467) & (!g2076) & (!g2077)) + ((g2706) & (!g2559) & (!g2632) & (g2467) & (g2076) & (g2077)) + ((g2706) & (!g2559) & (g2632) & (!g2467) & (!g2076) & (!g2077)) + ((g2706) & (!g2559) & (g2632) & (!g2467) & (!g2076) & (g2077)) + ((g2706) & (!g2559) & (g2632) & (g2467) & (!g2076) & (!g2077)) + ((g2706) & (!g2559) & (g2632) & (g2467) & (!g2076) & (g2077)) + ((g2706) & (!g2559) & (g2632) & (g2467) & (g2076) & (g2077)) + ((g2706) & (g2559) & (!g2632) & (!g2467) & (!g2076) & (!g2077)) + ((g2706) & (g2559) & (!g2632) & (!g2467) & (g2076) & (!g2077)) + ((g2706) & (g2559) & (!g2632) & (g2467) & (!g2076) & (!g2077)) + ((g2706) & (g2559) & (!g2632) & (g2467) & (g2076) & (!g2077)) + ((g2706) & (g2559) & (!g2632) & (g2467) & (g2076) & (g2077)) + ((g2706) & (g2559) & (g2632) & (!g2467) & (!g2076) & (!g2077)) + ((g2706) & (g2559) & (g2632) & (!g2467) & (!g2076) & (g2077)) + ((g2706) & (g2559) & (g2632) & (!g2467) & (g2076) & (!g2077)) + ((g2706) & (g2559) & (g2632) & (g2467) & (!g2076) & (!g2077)) + ((g2706) & (g2559) & (g2632) & (g2467) & (!g2076) & (g2077)) + ((g2706) & (g2559) & (g2632) & (g2467) & (g2076) & (!g2077)) + ((g2706) & (g2559) & (g2632) & (g2467) & (g2076) & (g2077)));
	assign g2708 = (((!g2707) & (!g2373) & (!g2374) & (g2191) & (g2073) & (g2125)) + ((!g2707) & (!g2373) & (g2374) & (!g2191) & (!g2073) & (g2125)) + ((!g2707) & (!g2373) & (g2374) & (g2191) & (!g2073) & (g2125)) + ((!g2707) & (!g2373) & (g2374) & (g2191) & (g2073) & (g2125)) + ((!g2707) & (g2373) & (!g2374) & (!g2191) & (g2073) & (!g2125)) + ((!g2707) & (g2373) & (!g2374) & (g2191) & (g2073) & (!g2125)) + ((!g2707) & (g2373) & (!g2374) & (g2191) & (g2073) & (g2125)) + ((!g2707) & (g2373) & (g2374) & (!g2191) & (!g2073) & (g2125)) + ((!g2707) & (g2373) & (g2374) & (!g2191) & (g2073) & (!g2125)) + ((!g2707) & (g2373) & (g2374) & (g2191) & (!g2073) & (g2125)) + ((!g2707) & (g2373) & (g2374) & (g2191) & (g2073) & (!g2125)) + ((!g2707) & (g2373) & (g2374) & (g2191) & (g2073) & (g2125)) + ((g2707) & (!g2373) & (!g2374) & (!g2191) & (!g2073) & (!g2125)) + ((g2707) & (!g2373) & (!g2374) & (g2191) & (!g2073) & (!g2125)) + ((g2707) & (!g2373) & (!g2374) & (g2191) & (g2073) & (g2125)) + ((g2707) & (!g2373) & (g2374) & (!g2191) & (!g2073) & (!g2125)) + ((g2707) & (!g2373) & (g2374) & (!g2191) & (!g2073) & (g2125)) + ((g2707) & (!g2373) & (g2374) & (g2191) & (!g2073) & (!g2125)) + ((g2707) & (!g2373) & (g2374) & (g2191) & (!g2073) & (g2125)) + ((g2707) & (!g2373) & (g2374) & (g2191) & (g2073) & (g2125)) + ((g2707) & (g2373) & (!g2374) & (!g2191) & (!g2073) & (!g2125)) + ((g2707) & (g2373) & (!g2374) & (!g2191) & (g2073) & (!g2125)) + ((g2707) & (g2373) & (!g2374) & (g2191) & (!g2073) & (!g2125)) + ((g2707) & (g2373) & (!g2374) & (g2191) & (g2073) & (!g2125)) + ((g2707) & (g2373) & (!g2374) & (g2191) & (g2073) & (g2125)) + ((g2707) & (g2373) & (g2374) & (!g2191) & (!g2073) & (!g2125)) + ((g2707) & (g2373) & (g2374) & (!g2191) & (!g2073) & (g2125)) + ((g2707) & (g2373) & (g2374) & (!g2191) & (g2073) & (!g2125)) + ((g2707) & (g2373) & (g2374) & (g2191) & (!g2073) & (!g2125)) + ((g2707) & (g2373) & (g2374) & (g2191) & (!g2073) & (g2125)) + ((g2707) & (g2373) & (g2374) & (g2191) & (g2073) & (!g2125)) + ((g2707) & (g2373) & (g2374) & (g2191) & (g2073) & (g2125)));
	assign g2709 = (((!g2088) & (!g2699) & (!g2124) & (!g2264) & (!g3360) & (g2708)) + ((!g2088) & (!g2699) & (!g2124) & (!g2264) & (g3360) & (g2708)) + ((!g2088) & (!g2699) & (!g2124) & (g2264) & (g3360) & (!g2708)) + ((!g2088) & (!g2699) & (!g2124) & (g2264) & (g3360) & (g2708)) + ((!g2088) & (g2699) & (!g2124) & (!g2264) & (!g3360) & (g2708)) + ((!g2088) & (g2699) & (!g2124) & (!g2264) & (g3360) & (g2708)) + ((!g2088) & (g2699) & (!g2124) & (g2264) & (g3360) & (!g2708)) + ((!g2088) & (g2699) & (!g2124) & (g2264) & (g3360) & (g2708)) + ((!g2088) & (g2699) & (g2124) & (!g2264) & (!g3360) & (!g2708)) + ((!g2088) & (g2699) & (g2124) & (!g2264) & (!g3360) & (g2708)) + ((!g2088) & (g2699) & (g2124) & (!g2264) & (g3360) & (!g2708)) + ((!g2088) & (g2699) & (g2124) & (!g2264) & (g3360) & (g2708)) + ((!g2088) & (g2699) & (g2124) & (g2264) & (!g3360) & (!g2708)) + ((!g2088) & (g2699) & (g2124) & (g2264) & (!g3360) & (g2708)) + ((!g2088) & (g2699) & (g2124) & (g2264) & (g3360) & (!g2708)) + ((!g2088) & (g2699) & (g2124) & (g2264) & (g3360) & (g2708)) + ((g2088) & (!g2699) & (!g2124) & (!g2264) & (!g3360) & (g2708)) + ((g2088) & (!g2699) & (!g2124) & (!g2264) & (g3360) & (g2708)) + ((g2088) & (!g2699) & (!g2124) & (g2264) & (g3360) & (!g2708)) + ((g2088) & (!g2699) & (!g2124) & (g2264) & (g3360) & (g2708)) + ((g2088) & (!g2699) & (g2124) & (!g2264) & (!g3360) & (!g2708)) + ((g2088) & (!g2699) & (g2124) & (!g2264) & (!g3360) & (g2708)) + ((g2088) & (!g2699) & (g2124) & (!g2264) & (g3360) & (!g2708)) + ((g2088) & (!g2699) & (g2124) & (!g2264) & (g3360) & (g2708)) + ((g2088) & (!g2699) & (g2124) & (g2264) & (!g3360) & (!g2708)) + ((g2088) & (!g2699) & (g2124) & (g2264) & (!g3360) & (g2708)) + ((g2088) & (!g2699) & (g2124) & (g2264) & (g3360) & (!g2708)) + ((g2088) & (!g2699) & (g2124) & (g2264) & (g3360) & (g2708)) + ((g2088) & (g2699) & (!g2124) & (!g2264) & (!g3360) & (g2708)) + ((g2088) & (g2699) & (!g2124) & (!g2264) & (g3360) & (g2708)) + ((g2088) & (g2699) & (!g2124) & (g2264) & (g3360) & (!g2708)) + ((g2088) & (g2699) & (!g2124) & (g2264) & (g3360) & (g2708)) + ((g2088) & (g2699) & (g2124) & (!g2264) & (!g3360) & (!g2708)) + ((g2088) & (g2699) & (g2124) & (!g2264) & (!g3360) & (g2708)) + ((g2088) & (g2699) & (g2124) & (!g2264) & (g3360) & (!g2708)) + ((g2088) & (g2699) & (g2124) & (!g2264) & (g3360) & (g2708)));
	assign g2710 = (((!g1185) & (!g2673) & (!sk[20]) & (g1230) & (!g1275)) + ((!g1185) & (!g2673) & (!sk[20]) & (g1230) & (g1275)) + ((!g1185) & (!g2673) & (sk[20]) & (!g1230) & (g1275)) + ((!g1185) & (!g2673) & (sk[20]) & (g1230) & (g1275)) + ((!g1185) & (g2673) & (!sk[20]) & (!g1230) & (g1275)) + ((!g1185) & (g2673) & (!sk[20]) & (g1230) & (!g1275)) + ((!g1185) & (g2673) & (!sk[20]) & (g1230) & (g1275)) + ((!g1185) & (g2673) & (sk[20]) & (!g1230) & (g1275)) + ((!g1185) & (g2673) & (sk[20]) & (g1230) & (g1275)) + ((g1185) & (!g2673) & (!sk[20]) & (!g1230) & (g1275)) + ((g1185) & (!g2673) & (!sk[20]) & (g1230) & (!g1275)) + ((g1185) & (!g2673) & (!sk[20]) & (g1230) & (g1275)) + ((g1185) & (!g2673) & (sk[20]) & (!g1230) & (g1275)) + ((g1185) & (!g2673) & (sk[20]) & (g1230) & (g1275)) + ((g1185) & (g2673) & (!sk[20]) & (!g1230) & (g1275)) + ((g1185) & (g2673) & (!sk[20]) & (g1230) & (!g1275)) + ((g1185) & (g2673) & (!sk[20]) & (g1230) & (g1275)) + ((g1185) & (g2673) & (sk[20]) & (!g1230) & (g1275)) + ((g1185) & (g2673) & (sk[20]) & (g1230) & (!g1275)));
	assign g2711 = (((!g109) & (!g678) & (!g1230) & (!g2693) & (!g2694) & (g1275)) + ((!g109) & (!g678) & (!g1230) & (!g2693) & (g2694) & (g1275)) + ((!g109) & (!g678) & (!g1230) & (g2693) & (!g2694) & (g1275)) + ((!g109) & (!g678) & (!g1230) & (g2693) & (g2694) & (g1275)) + ((!g109) & (!g678) & (g1230) & (!g2693) & (!g2694) & (g1275)) + ((!g109) & (!g678) & (g1230) & (!g2693) & (g2694) & (!g1275)) + ((!g109) & (!g678) & (g1230) & (g2693) & (!g2694) & (!g1275)) + ((!g109) & (!g678) & (g1230) & (g2693) & (g2694) & (!g1275)) + ((!g109) & (g678) & (!g1230) & (!g2693) & (!g2694) & (g1275)) + ((!g109) & (g678) & (!g1230) & (!g2693) & (g2694) & (!g1275)) + ((!g109) & (g678) & (!g1230) & (g2693) & (!g2694) & (!g1275)) + ((!g109) & (g678) & (!g1230) & (g2693) & (g2694) & (!g1275)) + ((!g109) & (g678) & (g1230) & (!g2693) & (!g2694) & (!g1275)) + ((!g109) & (g678) & (g1230) & (!g2693) & (g2694) & (!g1275)) + ((!g109) & (g678) & (g1230) & (g2693) & (!g2694) & (!g1275)) + ((!g109) & (g678) & (g1230) & (g2693) & (g2694) & (!g1275)) + ((g109) & (!g678) & (!g1230) & (!g2693) & (!g2694) & (!g1275)) + ((g109) & (!g678) & (!g1230) & (!g2693) & (g2694) & (!g1275)) + ((g109) & (!g678) & (!g1230) & (g2693) & (!g2694) & (!g1275)) + ((g109) & (!g678) & (!g1230) & (g2693) & (g2694) & (!g1275)) + ((g109) & (!g678) & (g1230) & (!g2693) & (!g2694) & (!g1275)) + ((g109) & (!g678) & (g1230) & (!g2693) & (g2694) & (g1275)) + ((g109) & (!g678) & (g1230) & (g2693) & (!g2694) & (g1275)) + ((g109) & (!g678) & (g1230) & (g2693) & (g2694) & (g1275)) + ((g109) & (g678) & (!g1230) & (!g2693) & (!g2694) & (!g1275)) + ((g109) & (g678) & (!g1230) & (!g2693) & (g2694) & (g1275)) + ((g109) & (g678) & (!g1230) & (g2693) & (!g2694) & (g1275)) + ((g109) & (g678) & (!g1230) & (g2693) & (g2694) & (g1275)) + ((g109) & (g678) & (g1230) & (!g2693) & (!g2694) & (g1275)) + ((g109) & (g678) & (g1230) & (!g2693) & (g2694) & (g1275)) + ((g109) & (g678) & (g1230) & (g2693) & (!g2694) & (g1275)) + ((g109) & (g678) & (g1230) & (g2693) & (g2694) & (g1275)));
	assign g5048 = (((!g2921) & (!sk[22]) & (g3101) & (!g2712)) + ((!g2921) & (!sk[22]) & (g3101) & (g2712)) + ((!g2921) & (sk[22]) & (!g3101) & (g2712)) + ((!g2921) & (sk[22]) & (g3101) & (g2712)) + ((g2921) & (!sk[22]) & (g3101) & (!g2712)) + ((g2921) & (!sk[22]) & (g3101) & (g2712)) + ((g2921) & (sk[22]) & (g3101) & (!g2712)) + ((g2921) & (sk[22]) & (g3101) & (g2712)));
	assign g2713 = (((!g1915) & (!sk[23]) & (!g2033) & (!g2034) & (g2711) & (!g2712)) + ((!g1915) & (!sk[23]) & (!g2033) & (!g2034) & (g2711) & (g2712)) + ((!g1915) & (!sk[23]) & (!g2033) & (g2034) & (g2711) & (!g2712)) + ((!g1915) & (!sk[23]) & (!g2033) & (g2034) & (g2711) & (g2712)) + ((!g1915) & (!sk[23]) & (g2033) & (!g2034) & (!g2711) & (!g2712)) + ((!g1915) & (!sk[23]) & (g2033) & (!g2034) & (!g2711) & (g2712)) + ((!g1915) & (!sk[23]) & (g2033) & (!g2034) & (g2711) & (!g2712)) + ((!g1915) & (!sk[23]) & (g2033) & (!g2034) & (g2711) & (g2712)) + ((!g1915) & (!sk[23]) & (g2033) & (g2034) & (!g2711) & (!g2712)) + ((!g1915) & (!sk[23]) & (g2033) & (g2034) & (!g2711) & (g2712)) + ((!g1915) & (!sk[23]) & (g2033) & (g2034) & (g2711) & (!g2712)) + ((!g1915) & (!sk[23]) & (g2033) & (g2034) & (g2711) & (g2712)) + ((!g1915) & (sk[23]) & (!g2033) & (!g2034) & (!g2711) & (g2712)) + ((!g1915) & (sk[23]) & (!g2033) & (!g2034) & (g2711) & (g2712)) + ((!g1915) & (sk[23]) & (g2033) & (!g2034) & (g2711) & (!g2712)) + ((!g1915) & (sk[23]) & (g2033) & (!g2034) & (g2711) & (g2712)) + ((g1915) & (!sk[23]) & (!g2033) & (!g2034) & (g2711) & (!g2712)) + ((g1915) & (!sk[23]) & (!g2033) & (!g2034) & (g2711) & (g2712)) + ((g1915) & (!sk[23]) & (!g2033) & (g2034) & (g2711) & (!g2712)) + ((g1915) & (!sk[23]) & (!g2033) & (g2034) & (g2711) & (g2712)) + ((g1915) & (!sk[23]) & (g2033) & (!g2034) & (!g2711) & (!g2712)) + ((g1915) & (!sk[23]) & (g2033) & (!g2034) & (!g2711) & (g2712)) + ((g1915) & (!sk[23]) & (g2033) & (!g2034) & (g2711) & (!g2712)) + ((g1915) & (!sk[23]) & (g2033) & (!g2034) & (g2711) & (g2712)) + ((g1915) & (!sk[23]) & (g2033) & (g2034) & (!g2711) & (!g2712)) + ((g1915) & (!sk[23]) & (g2033) & (g2034) & (!g2711) & (g2712)) + ((g1915) & (!sk[23]) & (g2033) & (g2034) & (g2711) & (!g2712)) + ((g1915) & (!sk[23]) & (g2033) & (g2034) & (g2711) & (g2712)) + ((g1915) & (sk[23]) & (!g2033) & (!g2034) & (!g2711) & (g2712)) + ((g1915) & (sk[23]) & (!g2033) & (!g2034) & (g2711) & (g2712)) + ((g1915) & (sk[23]) & (!g2033) & (g2034) & (!g2711) & (!g2712)) + ((g1915) & (sk[23]) & (!g2033) & (g2034) & (!g2711) & (g2712)) + ((g1915) & (sk[23]) & (!g2033) & (g2034) & (g2711) & (!g2712)) + ((g1915) & (sk[23]) & (!g2033) & (g2034) & (g2711) & (g2712)) + ((g1915) & (sk[23]) & (g2033) & (!g2034) & (g2711) & (!g2712)) + ((g1915) & (sk[23]) & (g2033) & (!g2034) & (g2711) & (g2712)));
	assign g2714 = (((!g2329) & (!g2029) & (!g2408) & (g2710) & (!sk[24]) & (!g2713)) + ((!g2329) & (!g2029) & (!g2408) & (g2710) & (!sk[24]) & (g2713)) + ((!g2329) & (!g2029) & (g2408) & (g2710) & (!sk[24]) & (!g2713)) + ((!g2329) & (!g2029) & (g2408) & (g2710) & (!sk[24]) & (g2713)) + ((!g2329) & (g2029) & (!g2408) & (!g2710) & (!sk[24]) & (!g2713)) + ((!g2329) & (g2029) & (!g2408) & (!g2710) & (!sk[24]) & (g2713)) + ((!g2329) & (g2029) & (!g2408) & (g2710) & (!sk[24]) & (!g2713)) + ((!g2329) & (g2029) & (!g2408) & (g2710) & (!sk[24]) & (g2713)) + ((!g2329) & (g2029) & (g2408) & (!g2710) & (!sk[24]) & (!g2713)) + ((!g2329) & (g2029) & (g2408) & (!g2710) & (!sk[24]) & (g2713)) + ((!g2329) & (g2029) & (g2408) & (g2710) & (!sk[24]) & (!g2713)) + ((!g2329) & (g2029) & (g2408) & (g2710) & (!sk[24]) & (g2713)) + ((g2329) & (!g2029) & (!g2408) & (g2710) & (!sk[24]) & (!g2713)) + ((g2329) & (!g2029) & (!g2408) & (g2710) & (!sk[24]) & (g2713)) + ((g2329) & (!g2029) & (g2408) & (!g2710) & (sk[24]) & (g2713)) + ((g2329) & (!g2029) & (g2408) & (g2710) & (!sk[24]) & (!g2713)) + ((g2329) & (!g2029) & (g2408) & (g2710) & (!sk[24]) & (g2713)) + ((g2329) & (!g2029) & (g2408) & (g2710) & (sk[24]) & (g2713)) + ((g2329) & (g2029) & (!g2408) & (!g2710) & (!sk[24]) & (!g2713)) + ((g2329) & (g2029) & (!g2408) & (!g2710) & (!sk[24]) & (g2713)) + ((g2329) & (g2029) & (!g2408) & (g2710) & (!sk[24]) & (!g2713)) + ((g2329) & (g2029) & (!g2408) & (g2710) & (!sk[24]) & (g2713)) + ((g2329) & (g2029) & (g2408) & (!g2710) & (!sk[24]) & (!g2713)) + ((g2329) & (g2029) & (g2408) & (!g2710) & (!sk[24]) & (g2713)) + ((g2329) & (g2029) & (g2408) & (g2710) & (!sk[24]) & (!g2713)) + ((g2329) & (g2029) & (g2408) & (g2710) & (!sk[24]) & (g2713)) + ((g2329) & (g2029) & (g2408) & (g2710) & (sk[24]) & (!g2713)) + ((g2329) & (g2029) & (g2408) & (g2710) & (sk[24]) & (g2713)));
	assign g2716 = (((!g2089) & (!sk[25]) & (g2715)) + ((!g2089) & (sk[25]) & (g2715)) + ((g2089) & (!sk[25]) & (g2715)) + ((g2089) & (sk[25]) & (!g2715)));
	assign g2717 = (((!g2088) & (!g2096) & (!g2680) & (!g2681) & (!g2699) & (g2716)) + ((!g2088) & (!g2096) & (!g2680) & (!g2681) & (g2699) & (g2716)) + ((!g2088) & (!g2096) & (!g2680) & (g2681) & (!g2699) & (g2716)) + ((!g2088) & (!g2096) & (!g2680) & (g2681) & (g2699) & (g2716)) + ((!g2088) & (!g2096) & (g2680) & (!g2681) & (!g2699) & (g2716)) + ((!g2088) & (!g2096) & (g2680) & (!g2681) & (g2699) & (g2716)) + ((!g2088) & (!g2096) & (g2680) & (g2681) & (!g2699) & (g2716)) + ((!g2088) & (!g2096) & (g2680) & (g2681) & (g2699) & (!g2716)) + ((!g2088) & (g2096) & (!g2680) & (!g2681) & (!g2699) & (g2716)) + ((!g2088) & (g2096) & (!g2680) & (!g2681) & (g2699) & (g2716)) + ((!g2088) & (g2096) & (!g2680) & (g2681) & (!g2699) & (g2716)) + ((!g2088) & (g2096) & (!g2680) & (g2681) & (g2699) & (!g2716)) + ((!g2088) & (g2096) & (g2680) & (!g2681) & (!g2699) & (g2716)) + ((!g2088) & (g2096) & (g2680) & (!g2681) & (g2699) & (!g2716)) + ((!g2088) & (g2096) & (g2680) & (g2681) & (!g2699) & (g2716)) + ((!g2088) & (g2096) & (g2680) & (g2681) & (g2699) & (!g2716)) + ((g2088) & (!g2096) & (!g2680) & (!g2681) & (!g2699) & (g2716)) + ((g2088) & (!g2096) & (!g2680) & (!g2681) & (g2699) & (!g2716)) + ((g2088) & (!g2096) & (!g2680) & (g2681) & (!g2699) & (g2716)) + ((g2088) & (!g2096) & (!g2680) & (g2681) & (g2699) & (!g2716)) + ((g2088) & (!g2096) & (g2680) & (!g2681) & (!g2699) & (g2716)) + ((g2088) & (!g2096) & (g2680) & (!g2681) & (g2699) & (!g2716)) + ((g2088) & (!g2096) & (g2680) & (g2681) & (!g2699) & (!g2716)) + ((g2088) & (!g2096) & (g2680) & (g2681) & (g2699) & (!g2716)) + ((g2088) & (g2096) & (!g2680) & (!g2681) & (!g2699) & (g2716)) + ((g2088) & (g2096) & (!g2680) & (!g2681) & (g2699) & (!g2716)) + ((g2088) & (g2096) & (!g2680) & (g2681) & (!g2699) & (!g2716)) + ((g2088) & (g2096) & (!g2680) & (g2681) & (g2699) & (!g2716)) + ((g2088) & (g2096) & (g2680) & (!g2681) & (!g2699) & (!g2716)) + ((g2088) & (g2096) & (g2680) & (!g2681) & (g2699) & (!g2716)) + ((g2088) & (g2096) & (g2680) & (g2681) & (!g2699) & (!g2716)) + ((g2088) & (g2096) & (g2680) & (g2681) & (g2699) & (!g2716)));
	assign g2718 = (((!g2661) & (!sk[27]) & (!g2662) & (!g2682) & (g2700) & (!g2717)) + ((!g2661) & (!sk[27]) & (!g2662) & (!g2682) & (g2700) & (g2717)) + ((!g2661) & (!sk[27]) & (!g2662) & (g2682) & (g2700) & (!g2717)) + ((!g2661) & (!sk[27]) & (!g2662) & (g2682) & (g2700) & (g2717)) + ((!g2661) & (!sk[27]) & (g2662) & (!g2682) & (!g2700) & (!g2717)) + ((!g2661) & (!sk[27]) & (g2662) & (!g2682) & (!g2700) & (g2717)) + ((!g2661) & (!sk[27]) & (g2662) & (!g2682) & (g2700) & (!g2717)) + ((!g2661) & (!sk[27]) & (g2662) & (!g2682) & (g2700) & (g2717)) + ((!g2661) & (!sk[27]) & (g2662) & (g2682) & (!g2700) & (!g2717)) + ((!g2661) & (!sk[27]) & (g2662) & (g2682) & (!g2700) & (g2717)) + ((!g2661) & (!sk[27]) & (g2662) & (g2682) & (g2700) & (!g2717)) + ((!g2661) & (!sk[27]) & (g2662) & (g2682) & (g2700) & (g2717)) + ((!g2661) & (sk[27]) & (!g2662) & (!g2682) & (!g2700) & (g2717)) + ((!g2661) & (sk[27]) & (!g2662) & (!g2682) & (g2700) & (g2717)) + ((!g2661) & (sk[27]) & (!g2662) & (g2682) & (!g2700) & (g2717)) + ((!g2661) & (sk[27]) & (!g2662) & (g2682) & (g2700) & (g2717)) + ((!g2661) & (sk[27]) & (g2662) & (!g2682) & (!g2700) & (g2717)) + ((!g2661) & (sk[27]) & (g2662) & (!g2682) & (g2700) & (g2717)) + ((!g2661) & (sk[27]) & (g2662) & (g2682) & (!g2700) & (g2717)) + ((!g2661) & (sk[27]) & (g2662) & (g2682) & (g2700) & (g2717)) + ((g2661) & (!sk[27]) & (!g2662) & (!g2682) & (g2700) & (!g2717)) + ((g2661) & (!sk[27]) & (!g2662) & (!g2682) & (g2700) & (g2717)) + ((g2661) & (!sk[27]) & (!g2662) & (g2682) & (g2700) & (!g2717)) + ((g2661) & (!sk[27]) & (!g2662) & (g2682) & (g2700) & (g2717)) + ((g2661) & (!sk[27]) & (g2662) & (!g2682) & (!g2700) & (!g2717)) + ((g2661) & (!sk[27]) & (g2662) & (!g2682) & (!g2700) & (g2717)) + ((g2661) & (!sk[27]) & (g2662) & (!g2682) & (g2700) & (!g2717)) + ((g2661) & (!sk[27]) & (g2662) & (!g2682) & (g2700) & (g2717)) + ((g2661) & (!sk[27]) & (g2662) & (g2682) & (!g2700) & (!g2717)) + ((g2661) & (!sk[27]) & (g2662) & (g2682) & (!g2700) & (g2717)) + ((g2661) & (!sk[27]) & (g2662) & (g2682) & (g2700) & (!g2717)) + ((g2661) & (!sk[27]) & (g2662) & (g2682) & (g2700) & (g2717)) + ((g2661) & (sk[27]) & (!g2662) & (!g2682) & (!g2700) & (g2717)) + ((g2661) & (sk[27]) & (!g2662) & (!g2682) & (g2700) & (g2717)) + ((g2661) & (sk[27]) & (!g2662) & (g2682) & (!g2700) & (g2717)) + ((g2661) & (sk[27]) & (!g2662) & (g2682) & (g2700) & (g2717)) + ((g2661) & (sk[27]) & (g2662) & (!g2682) & (!g2700) & (g2717)) + ((g2661) & (sk[27]) & (g2662) & (!g2682) & (g2700) & (g2717)) + ((g2661) & (sk[27]) & (g2662) & (g2682) & (!g2700) & (g2717)) + ((g2661) & (sk[27]) & (g2662) & (g2682) & (g2700) & (!g2717)));
	assign g2719 = (((!sk[28]) & (g2702) & (!g2703) & (!g2704)) + ((!sk[28]) & (g2702) & (!g2703) & (g2704)) + ((!sk[28]) & (g2702) & (g2703) & (!g2704)) + ((!sk[28]) & (g2702) & (g2703) & (g2704)) + ((sk[28]) & (!g2702) & (!g2703) & (g2704)) + ((sk[28]) & (!g2702) & (g2703) & (!g2704)) + ((sk[28]) & (!g2702) & (g2703) & (g2704)) + ((sk[28]) & (g2702) & (g2703) & (g2704)));
	assign g2720 = (((!g2699) & (!sk[29]) & (g2088)) + ((!g2699) & (sk[29]) & (g2088)) + ((g2699) & (!sk[29]) & (g2088)));
	assign g2721 = (((!sk[30]) & (!g2715) & (g2089)) + ((!sk[30]) & (g2715) & (g2089)) + ((sk[30]) & (!g2715) & (!g2089)) + ((sk[30]) & (g2715) & (g2089)));
	assign g2722 = (((!g2719) & (!g2720) & (sk[31]) & (g2721)) + ((!g2719) & (g2720) & (sk[31]) & (!g2721)) + ((g2719) & (!g2720) & (!sk[31]) & (!g2721)) + ((g2719) & (!g2720) & (!sk[31]) & (g2721)) + ((g2719) & (!g2720) & (sk[31]) & (!g2721)) + ((g2719) & (g2720) & (!sk[31]) & (!g2721)) + ((g2719) & (g2720) & (!sk[31]) & (g2721)) + ((g2719) & (g2720) & (sk[31]) & (g2721)));
	assign g2723 = (((!g2089) & (!g2088) & (!g2096) & (g2095) & (g2071) & (g2074)) + ((!g2089) & (!g2088) & (g2096) & (!g2095) & (!g2071) & (g2074)) + ((!g2089) & (!g2088) & (g2096) & (g2095) & (!g2071) & (g2074)) + ((!g2089) & (!g2088) & (g2096) & (g2095) & (g2071) & (g2074)) + ((!g2089) & (g2088) & (!g2096) & (!g2095) & (g2071) & (!g2074)) + ((!g2089) & (g2088) & (!g2096) & (g2095) & (g2071) & (!g2074)) + ((!g2089) & (g2088) & (!g2096) & (g2095) & (g2071) & (g2074)) + ((!g2089) & (g2088) & (g2096) & (!g2095) & (!g2071) & (g2074)) + ((!g2089) & (g2088) & (g2096) & (!g2095) & (g2071) & (!g2074)) + ((!g2089) & (g2088) & (g2096) & (g2095) & (!g2071) & (g2074)) + ((!g2089) & (g2088) & (g2096) & (g2095) & (g2071) & (!g2074)) + ((!g2089) & (g2088) & (g2096) & (g2095) & (g2071) & (g2074)) + ((g2089) & (!g2088) & (!g2096) & (!g2095) & (!g2071) & (!g2074)) + ((g2089) & (!g2088) & (!g2096) & (g2095) & (!g2071) & (!g2074)) + ((g2089) & (!g2088) & (!g2096) & (g2095) & (g2071) & (g2074)) + ((g2089) & (!g2088) & (g2096) & (!g2095) & (!g2071) & (!g2074)) + ((g2089) & (!g2088) & (g2096) & (!g2095) & (!g2071) & (g2074)) + ((g2089) & (!g2088) & (g2096) & (g2095) & (!g2071) & (!g2074)) + ((g2089) & (!g2088) & (g2096) & (g2095) & (!g2071) & (g2074)) + ((g2089) & (!g2088) & (g2096) & (g2095) & (g2071) & (g2074)) + ((g2089) & (g2088) & (!g2096) & (!g2095) & (!g2071) & (!g2074)) + ((g2089) & (g2088) & (!g2096) & (!g2095) & (g2071) & (!g2074)) + ((g2089) & (g2088) & (!g2096) & (g2095) & (!g2071) & (!g2074)) + ((g2089) & (g2088) & (!g2096) & (g2095) & (g2071) & (!g2074)) + ((g2089) & (g2088) & (!g2096) & (g2095) & (g2071) & (g2074)) + ((g2089) & (g2088) & (g2096) & (!g2095) & (!g2071) & (!g2074)) + ((g2089) & (g2088) & (g2096) & (!g2095) & (!g2071) & (g2074)) + ((g2089) & (g2088) & (g2096) & (!g2095) & (g2071) & (!g2074)) + ((g2089) & (g2088) & (g2096) & (g2095) & (!g2071) & (!g2074)) + ((g2089) & (g2088) & (g2096) & (g2095) & (!g2071) & (g2074)) + ((g2089) & (g2088) & (g2096) & (g2095) & (g2071) & (!g2074)) + ((g2089) & (g2088) & (g2096) & (g2095) & (g2071) & (g2074)));
	assign g2724 = (((!g2723) & (!g2580) & (!g2650) & (g2490) & (g2076) & (g2077)) + ((!g2723) & (!g2580) & (g2650) & (!g2490) & (!g2076) & (g2077)) + ((!g2723) & (!g2580) & (g2650) & (g2490) & (!g2076) & (g2077)) + ((!g2723) & (!g2580) & (g2650) & (g2490) & (g2076) & (g2077)) + ((!g2723) & (g2580) & (!g2650) & (!g2490) & (g2076) & (!g2077)) + ((!g2723) & (g2580) & (!g2650) & (g2490) & (g2076) & (!g2077)) + ((!g2723) & (g2580) & (!g2650) & (g2490) & (g2076) & (g2077)) + ((!g2723) & (g2580) & (g2650) & (!g2490) & (!g2076) & (g2077)) + ((!g2723) & (g2580) & (g2650) & (!g2490) & (g2076) & (!g2077)) + ((!g2723) & (g2580) & (g2650) & (g2490) & (!g2076) & (g2077)) + ((!g2723) & (g2580) & (g2650) & (g2490) & (g2076) & (!g2077)) + ((!g2723) & (g2580) & (g2650) & (g2490) & (g2076) & (g2077)) + ((g2723) & (!g2580) & (!g2650) & (!g2490) & (!g2076) & (!g2077)) + ((g2723) & (!g2580) & (!g2650) & (g2490) & (!g2076) & (!g2077)) + ((g2723) & (!g2580) & (!g2650) & (g2490) & (g2076) & (g2077)) + ((g2723) & (!g2580) & (g2650) & (!g2490) & (!g2076) & (!g2077)) + ((g2723) & (!g2580) & (g2650) & (!g2490) & (!g2076) & (g2077)) + ((g2723) & (!g2580) & (g2650) & (g2490) & (!g2076) & (!g2077)) + ((g2723) & (!g2580) & (g2650) & (g2490) & (!g2076) & (g2077)) + ((g2723) & (!g2580) & (g2650) & (g2490) & (g2076) & (g2077)) + ((g2723) & (g2580) & (!g2650) & (!g2490) & (!g2076) & (!g2077)) + ((g2723) & (g2580) & (!g2650) & (!g2490) & (g2076) & (!g2077)) + ((g2723) & (g2580) & (!g2650) & (g2490) & (!g2076) & (!g2077)) + ((g2723) & (g2580) & (!g2650) & (g2490) & (g2076) & (!g2077)) + ((g2723) & (g2580) & (!g2650) & (g2490) & (g2076) & (g2077)) + ((g2723) & (g2580) & (g2650) & (!g2490) & (!g2076) & (!g2077)) + ((g2723) & (g2580) & (g2650) & (!g2490) & (!g2076) & (g2077)) + ((g2723) & (g2580) & (g2650) & (!g2490) & (g2076) & (!g2077)) + ((g2723) & (g2580) & (g2650) & (g2490) & (!g2076) & (!g2077)) + ((g2723) & (g2580) & (g2650) & (g2490) & (!g2076) & (g2077)) + ((g2723) & (g2580) & (g2650) & (g2490) & (g2076) & (!g2077)) + ((g2723) & (g2580) & (g2650) & (g2490) & (g2076) & (g2077)));
	assign g2725 = (((!g2724) & (!g2403) & (!g2401) & (g2191) & (g2073) & (g2125)) + ((!g2724) & (!g2403) & (g2401) & (!g2191) & (!g2073) & (g2125)) + ((!g2724) & (!g2403) & (g2401) & (g2191) & (!g2073) & (g2125)) + ((!g2724) & (!g2403) & (g2401) & (g2191) & (g2073) & (g2125)) + ((!g2724) & (g2403) & (!g2401) & (!g2191) & (g2073) & (!g2125)) + ((!g2724) & (g2403) & (!g2401) & (g2191) & (g2073) & (!g2125)) + ((!g2724) & (g2403) & (!g2401) & (g2191) & (g2073) & (g2125)) + ((!g2724) & (g2403) & (g2401) & (!g2191) & (!g2073) & (g2125)) + ((!g2724) & (g2403) & (g2401) & (!g2191) & (g2073) & (!g2125)) + ((!g2724) & (g2403) & (g2401) & (g2191) & (!g2073) & (g2125)) + ((!g2724) & (g2403) & (g2401) & (g2191) & (g2073) & (!g2125)) + ((!g2724) & (g2403) & (g2401) & (g2191) & (g2073) & (g2125)) + ((g2724) & (!g2403) & (!g2401) & (!g2191) & (!g2073) & (!g2125)) + ((g2724) & (!g2403) & (!g2401) & (g2191) & (!g2073) & (!g2125)) + ((g2724) & (!g2403) & (!g2401) & (g2191) & (g2073) & (g2125)) + ((g2724) & (!g2403) & (g2401) & (!g2191) & (!g2073) & (!g2125)) + ((g2724) & (!g2403) & (g2401) & (!g2191) & (!g2073) & (g2125)) + ((g2724) & (!g2403) & (g2401) & (g2191) & (!g2073) & (!g2125)) + ((g2724) & (!g2403) & (g2401) & (g2191) & (!g2073) & (g2125)) + ((g2724) & (!g2403) & (g2401) & (g2191) & (g2073) & (g2125)) + ((g2724) & (g2403) & (!g2401) & (!g2191) & (!g2073) & (!g2125)) + ((g2724) & (g2403) & (!g2401) & (!g2191) & (g2073) & (!g2125)) + ((g2724) & (g2403) & (!g2401) & (g2191) & (!g2073) & (!g2125)) + ((g2724) & (g2403) & (!g2401) & (g2191) & (g2073) & (!g2125)) + ((g2724) & (g2403) & (!g2401) & (g2191) & (g2073) & (g2125)) + ((g2724) & (g2403) & (g2401) & (!g2191) & (!g2073) & (!g2125)) + ((g2724) & (g2403) & (g2401) & (!g2191) & (!g2073) & (g2125)) + ((g2724) & (g2403) & (g2401) & (!g2191) & (g2073) & (!g2125)) + ((g2724) & (g2403) & (g2401) & (g2191) & (!g2073) & (!g2125)) + ((g2724) & (g2403) & (g2401) & (g2191) & (!g2073) & (g2125)) + ((g2724) & (g2403) & (g2401) & (g2191) & (g2073) & (!g2125)) + ((g2724) & (g2403) & (g2401) & (g2191) & (g2073) & (g2125)));
	assign g2726 = (((!g2089) & (!g2715) & (!g2124) & (!g2264) & (!g3336) & (g2725)) + ((!g2089) & (!g2715) & (!g2124) & (!g2264) & (g3336) & (g2725)) + ((!g2089) & (!g2715) & (!g2124) & (g2264) & (g3336) & (!g2725)) + ((!g2089) & (!g2715) & (!g2124) & (g2264) & (g3336) & (g2725)) + ((!g2089) & (g2715) & (!g2124) & (!g2264) & (!g3336) & (g2725)) + ((!g2089) & (g2715) & (!g2124) & (!g2264) & (g3336) & (g2725)) + ((!g2089) & (g2715) & (!g2124) & (g2264) & (g3336) & (!g2725)) + ((!g2089) & (g2715) & (!g2124) & (g2264) & (g3336) & (g2725)) + ((!g2089) & (g2715) & (g2124) & (!g2264) & (!g3336) & (!g2725)) + ((!g2089) & (g2715) & (g2124) & (!g2264) & (!g3336) & (g2725)) + ((!g2089) & (g2715) & (g2124) & (!g2264) & (g3336) & (!g2725)) + ((!g2089) & (g2715) & (g2124) & (!g2264) & (g3336) & (g2725)) + ((!g2089) & (g2715) & (g2124) & (g2264) & (!g3336) & (!g2725)) + ((!g2089) & (g2715) & (g2124) & (g2264) & (!g3336) & (g2725)) + ((!g2089) & (g2715) & (g2124) & (g2264) & (g3336) & (!g2725)) + ((!g2089) & (g2715) & (g2124) & (g2264) & (g3336) & (g2725)) + ((g2089) & (!g2715) & (!g2124) & (!g2264) & (!g3336) & (g2725)) + ((g2089) & (!g2715) & (!g2124) & (!g2264) & (g3336) & (g2725)) + ((g2089) & (!g2715) & (!g2124) & (g2264) & (g3336) & (!g2725)) + ((g2089) & (!g2715) & (!g2124) & (g2264) & (g3336) & (g2725)) + ((g2089) & (!g2715) & (g2124) & (!g2264) & (!g3336) & (!g2725)) + ((g2089) & (!g2715) & (g2124) & (!g2264) & (!g3336) & (g2725)) + ((g2089) & (!g2715) & (g2124) & (!g2264) & (g3336) & (!g2725)) + ((g2089) & (!g2715) & (g2124) & (!g2264) & (g3336) & (g2725)) + ((g2089) & (!g2715) & (g2124) & (g2264) & (!g3336) & (!g2725)) + ((g2089) & (!g2715) & (g2124) & (g2264) & (!g3336) & (g2725)) + ((g2089) & (!g2715) & (g2124) & (g2264) & (g3336) & (!g2725)) + ((g2089) & (!g2715) & (g2124) & (g2264) & (g3336) & (g2725)) + ((g2089) & (g2715) & (!g2124) & (!g2264) & (!g3336) & (g2725)) + ((g2089) & (g2715) & (!g2124) & (!g2264) & (g3336) & (g2725)) + ((g2089) & (g2715) & (!g2124) & (g2264) & (g3336) & (!g2725)) + ((g2089) & (g2715) & (!g2124) & (g2264) & (g3336) & (g2725)) + ((g2089) & (g2715) & (g2124) & (!g2264) & (!g3336) & (!g2725)) + ((g2089) & (g2715) & (g2124) & (!g2264) & (!g3336) & (g2725)) + ((g2089) & (g2715) & (g2124) & (!g2264) & (g3336) & (!g2725)) + ((g2089) & (g2715) & (g2124) & (!g2264) & (g3336) & (g2725)));
	assign g2727 = (((!g1185) & (!sk[36]) & (!g2673) & (!g1230) & (g1275)) + ((!g1185) & (!sk[36]) & (!g2673) & (g1230) & (!g1275)) + ((!g1185) & (!sk[36]) & (!g2673) & (g1230) & (g1275)) + ((!g1185) & (!sk[36]) & (g2673) & (!g1230) & (g1275)) + ((!g1185) & (!sk[36]) & (g2673) & (g1230) & (!g1275)) + ((!g1185) & (!sk[36]) & (g2673) & (g1230) & (g1275)) + ((g1185) & (!sk[36]) & (!g2673) & (!g1230) & (g1275)) + ((g1185) & (!sk[36]) & (!g2673) & (g1230) & (!g1275)) + ((g1185) & (!sk[36]) & (!g2673) & (g1230) & (g1275)) + ((g1185) & (!sk[36]) & (g2673) & (!g1230) & (g1275)) + ((g1185) & (!sk[36]) & (g2673) & (g1230) & (!g1275)) + ((g1185) & (!sk[36]) & (g2673) & (g1230) & (g1275)) + ((g1185) & (sk[36]) & (g2673) & (g1230) & (g1275)));
	assign g2728 = (((!g1320) & (!sk[37]) & (g2727)) + ((!g1320) & (sk[37]) & (g2727)) + ((g1320) & (!sk[37]) & (g2727)) + ((g1320) & (sk[37]) & (!g2727)));
	assign g2729 = (((!g109) & (!g678) & (!g1230) & (!g2693) & (!g2694) & (!g1275)) + ((!g109) & (!g678) & (!g1230) & (!g2693) & (!g2694) & (g1275)) + ((!g109) & (!g678) & (!g1230) & (!g2693) & (g2694) & (!g1275)) + ((!g109) & (!g678) & (!g1230) & (!g2693) & (g2694) & (g1275)) + ((!g109) & (!g678) & (!g1230) & (g2693) & (!g2694) & (!g1275)) + ((!g109) & (!g678) & (!g1230) & (g2693) & (!g2694) & (g1275)) + ((!g109) & (!g678) & (!g1230) & (g2693) & (g2694) & (!g1275)) + ((!g109) & (!g678) & (!g1230) & (g2693) & (g2694) & (g1275)) + ((!g109) & (!g678) & (g1230) & (!g2693) & (!g2694) & (!g1275)) + ((!g109) & (!g678) & (g1230) & (!g2693) & (!g2694) & (g1275)) + ((!g109) & (!g678) & (g1230) & (!g2693) & (g2694) & (!g1275)) + ((!g109) & (!g678) & (g1230) & (g2693) & (!g2694) & (!g1275)) + ((!g109) & (!g678) & (g1230) & (g2693) & (g2694) & (!g1275)) + ((!g109) & (g678) & (!g1230) & (!g2693) & (!g2694) & (!g1275)) + ((!g109) & (g678) & (!g1230) & (!g2693) & (!g2694) & (g1275)) + ((!g109) & (g678) & (!g1230) & (!g2693) & (g2694) & (!g1275)) + ((!g109) & (g678) & (!g1230) & (g2693) & (!g2694) & (!g1275)) + ((!g109) & (g678) & (!g1230) & (g2693) & (g2694) & (!g1275)) + ((!g109) & (g678) & (g1230) & (!g2693) & (!g2694) & (!g1275)) + ((!g109) & (g678) & (g1230) & (!g2693) & (g2694) & (!g1275)) + ((!g109) & (g678) & (g1230) & (g2693) & (!g2694) & (!g1275)) + ((!g109) & (g678) & (g1230) & (g2693) & (g2694) & (!g1275)) + ((g109) & (!g678) & (!g1230) & (!g2693) & (!g2694) & (!g1275)) + ((g109) & (!g678) & (!g1230) & (!g2693) & (g2694) & (!g1275)) + ((g109) & (!g678) & (!g1230) & (g2693) & (!g2694) & (!g1275)) + ((g109) & (!g678) & (!g1230) & (g2693) & (g2694) & (!g1275)) + ((g109) & (!g678) & (g1230) & (!g2693) & (!g2694) & (!g1275)) + ((g109) & (g678) & (!g1230) & (!g2693) & (!g2694) & (!g1275)));
	assign g2730 = (((!sk[39]) & (g108) & (!g1320) & (!g2729)) + ((!sk[39]) & (g108) & (!g1320) & (g2729)) + ((!sk[39]) & (g108) & (g1320) & (!g2729)) + ((!sk[39]) & (g108) & (g1320) & (g2729)) + ((sk[39]) & (!g108) & (!g1320) & (!g2729)) + ((sk[39]) & (!g108) & (g1320) & (g2729)) + ((sk[39]) & (g108) & (!g1320) & (g2729)) + ((sk[39]) & (g108) & (g1320) & (!g2729)));
	assign g5049 = (((!g2921) & (!g3103) & (sk[40]) & (g2731)) + ((!g2921) & (g3103) & (sk[40]) & (g2731)) + ((g2921) & (!g3103) & (!sk[40]) & (!g2731)) + ((g2921) & (!g3103) & (!sk[40]) & (g2731)) + ((g2921) & (g3103) & (!sk[40]) & (!g2731)) + ((g2921) & (g3103) & (!sk[40]) & (g2731)) + ((g2921) & (g3103) & (sk[40]) & (!g2731)) + ((g2921) & (g3103) & (sk[40]) & (g2731)));
	assign g2732 = (((!g1929) & (!g2033) & (!g2034) & (!sk[41]) & (g2730) & (!g2731)) + ((!g1929) & (!g2033) & (!g2034) & (!sk[41]) & (g2730) & (g2731)) + ((!g1929) & (!g2033) & (!g2034) & (sk[41]) & (!g2730) & (g2731)) + ((!g1929) & (!g2033) & (!g2034) & (sk[41]) & (g2730) & (g2731)) + ((!g1929) & (!g2033) & (g2034) & (!sk[41]) & (!g2730) & (!g2731)) + ((!g1929) & (!g2033) & (g2034) & (!sk[41]) & (!g2730) & (g2731)) + ((!g1929) & (!g2033) & (g2034) & (!sk[41]) & (g2730) & (!g2731)) + ((!g1929) & (!g2033) & (g2034) & (!sk[41]) & (g2730) & (g2731)) + ((!g1929) & (g2033) & (!g2034) & (!sk[41]) & (g2730) & (!g2731)) + ((!g1929) & (g2033) & (!g2034) & (!sk[41]) & (g2730) & (g2731)) + ((!g1929) & (g2033) & (!g2034) & (sk[41]) & (g2730) & (!g2731)) + ((!g1929) & (g2033) & (!g2034) & (sk[41]) & (g2730) & (g2731)) + ((!g1929) & (g2033) & (g2034) & (!sk[41]) & (!g2730) & (!g2731)) + ((!g1929) & (g2033) & (g2034) & (!sk[41]) & (!g2730) & (g2731)) + ((!g1929) & (g2033) & (g2034) & (!sk[41]) & (g2730) & (!g2731)) + ((!g1929) & (g2033) & (g2034) & (!sk[41]) & (g2730) & (g2731)) + ((g1929) & (!g2033) & (!g2034) & (!sk[41]) & (g2730) & (!g2731)) + ((g1929) & (!g2033) & (!g2034) & (!sk[41]) & (g2730) & (g2731)) + ((g1929) & (!g2033) & (!g2034) & (sk[41]) & (!g2730) & (g2731)) + ((g1929) & (!g2033) & (!g2034) & (sk[41]) & (g2730) & (g2731)) + ((g1929) & (!g2033) & (g2034) & (!sk[41]) & (!g2730) & (!g2731)) + ((g1929) & (!g2033) & (g2034) & (!sk[41]) & (!g2730) & (g2731)) + ((g1929) & (!g2033) & (g2034) & (!sk[41]) & (g2730) & (!g2731)) + ((g1929) & (!g2033) & (g2034) & (!sk[41]) & (g2730) & (g2731)) + ((g1929) & (!g2033) & (g2034) & (sk[41]) & (!g2730) & (!g2731)) + ((g1929) & (!g2033) & (g2034) & (sk[41]) & (!g2730) & (g2731)) + ((g1929) & (!g2033) & (g2034) & (sk[41]) & (g2730) & (!g2731)) + ((g1929) & (!g2033) & (g2034) & (sk[41]) & (g2730) & (g2731)) + ((g1929) & (g2033) & (!g2034) & (!sk[41]) & (g2730) & (!g2731)) + ((g1929) & (g2033) & (!g2034) & (!sk[41]) & (g2730) & (g2731)) + ((g1929) & (g2033) & (!g2034) & (sk[41]) & (g2730) & (!g2731)) + ((g1929) & (g2033) & (!g2034) & (sk[41]) & (g2730) & (g2731)) + ((g1929) & (g2033) & (g2034) & (!sk[41]) & (!g2730) & (!g2731)) + ((g1929) & (g2033) & (g2034) & (!sk[41]) & (!g2730) & (g2731)) + ((g1929) & (g2033) & (g2034) & (!sk[41]) & (g2730) & (!g2731)) + ((g1929) & (g2033) & (g2034) & (!sk[41]) & (g2730) & (g2731)));
	assign g2733 = (((!g2329) & (!g2029) & (!sk[42]) & (!g2408) & (g2728) & (!g2732)) + ((!g2329) & (!g2029) & (!sk[42]) & (!g2408) & (g2728) & (g2732)) + ((!g2329) & (!g2029) & (!sk[42]) & (g2408) & (!g2728) & (!g2732)) + ((!g2329) & (!g2029) & (!sk[42]) & (g2408) & (!g2728) & (g2732)) + ((!g2329) & (!g2029) & (!sk[42]) & (g2408) & (g2728) & (!g2732)) + ((!g2329) & (!g2029) & (!sk[42]) & (g2408) & (g2728) & (g2732)) + ((!g2329) & (g2029) & (!sk[42]) & (!g2408) & (g2728) & (!g2732)) + ((!g2329) & (g2029) & (!sk[42]) & (!g2408) & (g2728) & (g2732)) + ((!g2329) & (g2029) & (!sk[42]) & (g2408) & (!g2728) & (!g2732)) + ((!g2329) & (g2029) & (!sk[42]) & (g2408) & (!g2728) & (g2732)) + ((!g2329) & (g2029) & (!sk[42]) & (g2408) & (g2728) & (!g2732)) + ((!g2329) & (g2029) & (!sk[42]) & (g2408) & (g2728) & (g2732)) + ((g2329) & (!g2029) & (!sk[42]) & (!g2408) & (g2728) & (!g2732)) + ((g2329) & (!g2029) & (!sk[42]) & (!g2408) & (g2728) & (g2732)) + ((g2329) & (!g2029) & (!sk[42]) & (g2408) & (!g2728) & (!g2732)) + ((g2329) & (!g2029) & (!sk[42]) & (g2408) & (!g2728) & (g2732)) + ((g2329) & (!g2029) & (!sk[42]) & (g2408) & (g2728) & (!g2732)) + ((g2329) & (!g2029) & (!sk[42]) & (g2408) & (g2728) & (g2732)) + ((g2329) & (!g2029) & (sk[42]) & (g2408) & (!g2728) & (g2732)) + ((g2329) & (!g2029) & (sk[42]) & (g2408) & (g2728) & (g2732)) + ((g2329) & (g2029) & (!sk[42]) & (!g2408) & (g2728) & (!g2732)) + ((g2329) & (g2029) & (!sk[42]) & (!g2408) & (g2728) & (g2732)) + ((g2329) & (g2029) & (!sk[42]) & (g2408) & (!g2728) & (!g2732)) + ((g2329) & (g2029) & (!sk[42]) & (g2408) & (!g2728) & (g2732)) + ((g2329) & (g2029) & (!sk[42]) & (g2408) & (g2728) & (!g2732)) + ((g2329) & (g2029) & (!sk[42]) & (g2408) & (g2728) & (g2732)) + ((g2329) & (g2029) & (sk[42]) & (g2408) & (g2728) & (!g2732)) + ((g2329) & (g2029) & (sk[42]) & (g2408) & (g2728) & (g2732)));
	assign g2735 = (((!g2088) & (!g2096) & (g2680) & (g2681) & (g2699) & (g2716)) + ((!g2088) & (g2096) & (!g2680) & (g2681) & (g2699) & (g2716)) + ((!g2088) & (g2096) & (g2680) & (!g2681) & (g2699) & (g2716)) + ((!g2088) & (g2096) & (g2680) & (g2681) & (g2699) & (g2716)) + ((g2088) & (!g2096) & (!g2680) & (!g2681) & (g2699) & (g2716)) + ((g2088) & (!g2096) & (!g2680) & (g2681) & (g2699) & (g2716)) + ((g2088) & (!g2096) & (g2680) & (!g2681) & (g2699) & (g2716)) + ((g2088) & (!g2096) & (g2680) & (g2681) & (!g2699) & (g2716)) + ((g2088) & (!g2096) & (g2680) & (g2681) & (g2699) & (g2716)) + ((g2088) & (g2096) & (!g2680) & (!g2681) & (g2699) & (g2716)) + ((g2088) & (g2096) & (!g2680) & (g2681) & (!g2699) & (g2716)) + ((g2088) & (g2096) & (!g2680) & (g2681) & (g2699) & (g2716)) + ((g2088) & (g2096) & (g2680) & (!g2681) & (!g2699) & (g2716)) + ((g2088) & (g2096) & (g2680) & (!g2681) & (g2699) & (g2716)) + ((g2088) & (g2096) & (g2680) & (g2681) & (!g2699) & (g2716)) + ((g2088) & (g2096) & (g2680) & (g2681) & (g2699) & (g2716)));
	assign g2736 = (((!sk[44]) & (!g2089) & (g2715)) + ((!sk[44]) & (g2089) & (g2715)) + ((sk[44]) & (g2089) & (g2715)));
	assign g2737 = (((!g2090) & (!g2734) & (!g2735) & (!sk[45]) & (g2736)) + ((!g2090) & (!g2734) & (!g2735) & (sk[45]) & (g2736)) + ((!g2090) & (!g2734) & (g2735) & (!sk[45]) & (!g2736)) + ((!g2090) & (!g2734) & (g2735) & (!sk[45]) & (g2736)) + ((!g2090) & (!g2734) & (g2735) & (sk[45]) & (!g2736)) + ((!g2090) & (!g2734) & (g2735) & (sk[45]) & (g2736)) + ((!g2090) & (g2734) & (!g2735) & (!sk[45]) & (g2736)) + ((!g2090) & (g2734) & (!g2735) & (sk[45]) & (!g2736)) + ((!g2090) & (g2734) & (g2735) & (!sk[45]) & (!g2736)) + ((!g2090) & (g2734) & (g2735) & (!sk[45]) & (g2736)) + ((g2090) & (!g2734) & (!g2735) & (!sk[45]) & (g2736)) + ((g2090) & (!g2734) & (!g2735) & (sk[45]) & (!g2736)) + ((g2090) & (!g2734) & (g2735) & (!sk[45]) & (!g2736)) + ((g2090) & (!g2734) & (g2735) & (!sk[45]) & (g2736)) + ((g2090) & (g2734) & (!g2735) & (!sk[45]) & (g2736)) + ((g2090) & (g2734) & (!g2735) & (sk[45]) & (g2736)) + ((g2090) & (g2734) & (g2735) & (!sk[45]) & (!g2736)) + ((g2090) & (g2734) & (g2735) & (!sk[45]) & (g2736)) + ((g2090) & (g2734) & (g2735) & (sk[45]) & (!g2736)) + ((g2090) & (g2734) & (g2735) & (sk[45]) & (g2736)));
	assign g2738 = (((!g2661) & (!g2662) & (!g2682) & (!sk[46]) & (g2700) & (!g2717)) + ((!g2661) & (!g2662) & (!g2682) & (!sk[46]) & (g2700) & (g2717)) + ((!g2661) & (!g2662) & (g2682) & (!sk[46]) & (!g2700) & (!g2717)) + ((!g2661) & (!g2662) & (g2682) & (!sk[46]) & (!g2700) & (g2717)) + ((!g2661) & (!g2662) & (g2682) & (!sk[46]) & (g2700) & (!g2717)) + ((!g2661) & (!g2662) & (g2682) & (!sk[46]) & (g2700) & (g2717)) + ((!g2661) & (g2662) & (!g2682) & (!sk[46]) & (g2700) & (!g2717)) + ((!g2661) & (g2662) & (!g2682) & (!sk[46]) & (g2700) & (g2717)) + ((!g2661) & (g2662) & (g2682) & (!sk[46]) & (!g2700) & (!g2717)) + ((!g2661) & (g2662) & (g2682) & (!sk[46]) & (!g2700) & (g2717)) + ((!g2661) & (g2662) & (g2682) & (!sk[46]) & (g2700) & (!g2717)) + ((!g2661) & (g2662) & (g2682) & (!sk[46]) & (g2700) & (g2717)) + ((g2661) & (!g2662) & (!g2682) & (!sk[46]) & (!g2700) & (!g2717)) + ((g2661) & (!g2662) & (!g2682) & (!sk[46]) & (!g2700) & (g2717)) + ((g2661) & (!g2662) & (!g2682) & (!sk[46]) & (g2700) & (!g2717)) + ((g2661) & (!g2662) & (!g2682) & (!sk[46]) & (g2700) & (g2717)) + ((g2661) & (!g2662) & (g2682) & (!sk[46]) & (!g2700) & (!g2717)) + ((g2661) & (!g2662) & (g2682) & (!sk[46]) & (!g2700) & (g2717)) + ((g2661) & (!g2662) & (g2682) & (!sk[46]) & (g2700) & (!g2717)) + ((g2661) & (!g2662) & (g2682) & (!sk[46]) & (g2700) & (g2717)) + ((g2661) & (g2662) & (!g2682) & (!sk[46]) & (!g2700) & (!g2717)) + ((g2661) & (g2662) & (!g2682) & (!sk[46]) & (!g2700) & (g2717)) + ((g2661) & (g2662) & (!g2682) & (!sk[46]) & (g2700) & (!g2717)) + ((g2661) & (g2662) & (!g2682) & (!sk[46]) & (g2700) & (g2717)) + ((g2661) & (g2662) & (g2682) & (!sk[46]) & (!g2700) & (!g2717)) + ((g2661) & (g2662) & (g2682) & (!sk[46]) & (!g2700) & (g2717)) + ((g2661) & (g2662) & (g2682) & (!sk[46]) & (g2700) & (!g2717)) + ((g2661) & (g2662) & (g2682) & (!sk[46]) & (g2700) & (g2717)) + ((g2661) & (g2662) & (g2682) & (sk[46]) & (g2700) & (g2717)));
	assign g2739 = (((!g2715) & (!sk[47]) & (g2089)) + ((!g2715) & (sk[47]) & (g2089)) + ((g2715) & (!sk[47]) & (g2089)));
	assign g2740 = (((!g2734) & (!sk[48]) & (g2090)) + ((!g2734) & (sk[48]) & (!g2090)) + ((g2734) & (!sk[48]) & (g2090)) + ((g2734) & (sk[48]) & (g2090)));
	assign g2741 = (((!g2719) & (!g2720) & (!g2721) & (!g2739) & (sk[49]) & (g2740)) + ((!g2719) & (!g2720) & (!g2721) & (g2739) & (!sk[49]) & (!g2740)) + ((!g2719) & (!g2720) & (!g2721) & (g2739) & (!sk[49]) & (g2740)) + ((!g2719) & (!g2720) & (!g2721) & (g2739) & (sk[49]) & (!g2740)) + ((!g2719) & (!g2720) & (g2721) & (!g2739) & (!sk[49]) & (!g2740)) + ((!g2719) & (!g2720) & (g2721) & (!g2739) & (!sk[49]) & (g2740)) + ((!g2719) & (!g2720) & (g2721) & (!g2739) & (sk[49]) & (g2740)) + ((!g2719) & (!g2720) & (g2721) & (g2739) & (!sk[49]) & (!g2740)) + ((!g2719) & (!g2720) & (g2721) & (g2739) & (!sk[49]) & (g2740)) + ((!g2719) & (!g2720) & (g2721) & (g2739) & (sk[49]) & (!g2740)) + ((!g2719) & (g2720) & (!g2721) & (!g2739) & (sk[49]) & (g2740)) + ((!g2719) & (g2720) & (!g2721) & (g2739) & (!sk[49]) & (!g2740)) + ((!g2719) & (g2720) & (!g2721) & (g2739) & (!sk[49]) & (g2740)) + ((!g2719) & (g2720) & (!g2721) & (g2739) & (sk[49]) & (!g2740)) + ((!g2719) & (g2720) & (g2721) & (!g2739) & (!sk[49]) & (!g2740)) + ((!g2719) & (g2720) & (g2721) & (!g2739) & (!sk[49]) & (g2740)) + ((!g2719) & (g2720) & (g2721) & (!g2739) & (sk[49]) & (!g2740)) + ((!g2719) & (g2720) & (g2721) & (g2739) & (!sk[49]) & (!g2740)) + ((!g2719) & (g2720) & (g2721) & (g2739) & (!sk[49]) & (g2740)) + ((!g2719) & (g2720) & (g2721) & (g2739) & (sk[49]) & (g2740)) + ((g2719) & (!g2720) & (!g2721) & (!g2739) & (!sk[49]) & (!g2740)) + ((g2719) & (!g2720) & (!g2721) & (!g2739) & (!sk[49]) & (g2740)) + ((g2719) & (!g2720) & (!g2721) & (!g2739) & (sk[49]) & (g2740)) + ((g2719) & (!g2720) & (!g2721) & (g2739) & (!sk[49]) & (!g2740)) + ((g2719) & (!g2720) & (!g2721) & (g2739) & (!sk[49]) & (g2740)) + ((g2719) & (!g2720) & (!g2721) & (g2739) & (sk[49]) & (!g2740)) + ((g2719) & (!g2720) & (g2721) & (!g2739) & (!sk[49]) & (!g2740)) + ((g2719) & (!g2720) & (g2721) & (!g2739) & (!sk[49]) & (g2740)) + ((g2719) & (!g2720) & (g2721) & (!g2739) & (sk[49]) & (!g2740)) + ((g2719) & (!g2720) & (g2721) & (g2739) & (!sk[49]) & (!g2740)) + ((g2719) & (!g2720) & (g2721) & (g2739) & (!sk[49]) & (g2740)) + ((g2719) & (!g2720) & (g2721) & (g2739) & (sk[49]) & (g2740)) + ((g2719) & (g2720) & (!g2721) & (!g2739) & (!sk[49]) & (!g2740)) + ((g2719) & (g2720) & (!g2721) & (!g2739) & (!sk[49]) & (g2740)) + ((g2719) & (g2720) & (!g2721) & (!g2739) & (sk[49]) & (!g2740)) + ((g2719) & (g2720) & (!g2721) & (g2739) & (!sk[49]) & (!g2740)) + ((g2719) & (g2720) & (!g2721) & (g2739) & (!sk[49]) & (g2740)) + ((g2719) & (g2720) & (!g2721) & (g2739) & (sk[49]) & (g2740)) + ((g2719) & (g2720) & (g2721) & (!g2739) & (!sk[49]) & (!g2740)) + ((g2719) & (g2720) & (g2721) & (!g2739) & (!sk[49]) & (g2740)) + ((g2719) & (g2720) & (g2721) & (!g2739) & (sk[49]) & (!g2740)) + ((g2719) & (g2720) & (g2721) & (g2739) & (!sk[49]) & (!g2740)) + ((g2719) & (g2720) & (g2721) & (g2739) & (!sk[49]) & (g2740)) + ((g2719) & (g2720) & (g2721) & (g2739) & (sk[49]) & (g2740)));
	assign g2742 = (((!g2090) & (!g2089) & (!g2088) & (g2096) & (g2071) & (g2074)) + ((!g2090) & (!g2089) & (g2088) & (!g2096) & (!g2071) & (g2074)) + ((!g2090) & (!g2089) & (g2088) & (g2096) & (!g2071) & (g2074)) + ((!g2090) & (!g2089) & (g2088) & (g2096) & (g2071) & (g2074)) + ((!g2090) & (g2089) & (!g2088) & (!g2096) & (g2071) & (!g2074)) + ((!g2090) & (g2089) & (!g2088) & (g2096) & (g2071) & (!g2074)) + ((!g2090) & (g2089) & (!g2088) & (g2096) & (g2071) & (g2074)) + ((!g2090) & (g2089) & (g2088) & (!g2096) & (!g2071) & (g2074)) + ((!g2090) & (g2089) & (g2088) & (!g2096) & (g2071) & (!g2074)) + ((!g2090) & (g2089) & (g2088) & (g2096) & (!g2071) & (g2074)) + ((!g2090) & (g2089) & (g2088) & (g2096) & (g2071) & (!g2074)) + ((!g2090) & (g2089) & (g2088) & (g2096) & (g2071) & (g2074)) + ((g2090) & (!g2089) & (!g2088) & (!g2096) & (!g2071) & (!g2074)) + ((g2090) & (!g2089) & (!g2088) & (g2096) & (!g2071) & (!g2074)) + ((g2090) & (!g2089) & (!g2088) & (g2096) & (g2071) & (g2074)) + ((g2090) & (!g2089) & (g2088) & (!g2096) & (!g2071) & (!g2074)) + ((g2090) & (!g2089) & (g2088) & (!g2096) & (!g2071) & (g2074)) + ((g2090) & (!g2089) & (g2088) & (g2096) & (!g2071) & (!g2074)) + ((g2090) & (!g2089) & (g2088) & (g2096) & (!g2071) & (g2074)) + ((g2090) & (!g2089) & (g2088) & (g2096) & (g2071) & (g2074)) + ((g2090) & (g2089) & (!g2088) & (!g2096) & (!g2071) & (!g2074)) + ((g2090) & (g2089) & (!g2088) & (!g2096) & (g2071) & (!g2074)) + ((g2090) & (g2089) & (!g2088) & (g2096) & (!g2071) & (!g2074)) + ((g2090) & (g2089) & (!g2088) & (g2096) & (g2071) & (!g2074)) + ((g2090) & (g2089) & (!g2088) & (g2096) & (g2071) & (g2074)) + ((g2090) & (g2089) & (g2088) & (!g2096) & (!g2071) & (!g2074)) + ((g2090) & (g2089) & (g2088) & (!g2096) & (!g2071) & (g2074)) + ((g2090) & (g2089) & (g2088) & (!g2096) & (g2071) & (!g2074)) + ((g2090) & (g2089) & (g2088) & (g2096) & (!g2071) & (!g2074)) + ((g2090) & (g2089) & (g2088) & (g2096) & (!g2071) & (g2074)) + ((g2090) & (g2089) & (g2088) & (g2096) & (g2071) & (!g2074)) + ((g2090) & (g2089) & (g2088) & (g2096) & (g2071) & (g2074)));
	assign g2743 = (((!g2742) & (!g2595) & (!g2669) & (g2514) & (g2076) & (g2077)) + ((!g2742) & (!g2595) & (g2669) & (!g2514) & (!g2076) & (g2077)) + ((!g2742) & (!g2595) & (g2669) & (g2514) & (!g2076) & (g2077)) + ((!g2742) & (!g2595) & (g2669) & (g2514) & (g2076) & (g2077)) + ((!g2742) & (g2595) & (!g2669) & (!g2514) & (g2076) & (!g2077)) + ((!g2742) & (g2595) & (!g2669) & (g2514) & (g2076) & (!g2077)) + ((!g2742) & (g2595) & (!g2669) & (g2514) & (g2076) & (g2077)) + ((!g2742) & (g2595) & (g2669) & (!g2514) & (!g2076) & (g2077)) + ((!g2742) & (g2595) & (g2669) & (!g2514) & (g2076) & (!g2077)) + ((!g2742) & (g2595) & (g2669) & (g2514) & (!g2076) & (g2077)) + ((!g2742) & (g2595) & (g2669) & (g2514) & (g2076) & (!g2077)) + ((!g2742) & (g2595) & (g2669) & (g2514) & (g2076) & (g2077)) + ((g2742) & (!g2595) & (!g2669) & (!g2514) & (!g2076) & (!g2077)) + ((g2742) & (!g2595) & (!g2669) & (g2514) & (!g2076) & (!g2077)) + ((g2742) & (!g2595) & (!g2669) & (g2514) & (g2076) & (g2077)) + ((g2742) & (!g2595) & (g2669) & (!g2514) & (!g2076) & (!g2077)) + ((g2742) & (!g2595) & (g2669) & (!g2514) & (!g2076) & (g2077)) + ((g2742) & (!g2595) & (g2669) & (g2514) & (!g2076) & (!g2077)) + ((g2742) & (!g2595) & (g2669) & (g2514) & (!g2076) & (g2077)) + ((g2742) & (!g2595) & (g2669) & (g2514) & (g2076) & (g2077)) + ((g2742) & (g2595) & (!g2669) & (!g2514) & (!g2076) & (!g2077)) + ((g2742) & (g2595) & (!g2669) & (!g2514) & (g2076) & (!g2077)) + ((g2742) & (g2595) & (!g2669) & (g2514) & (!g2076) & (!g2077)) + ((g2742) & (g2595) & (!g2669) & (g2514) & (g2076) & (!g2077)) + ((g2742) & (g2595) & (!g2669) & (g2514) & (g2076) & (g2077)) + ((g2742) & (g2595) & (g2669) & (!g2514) & (!g2076) & (!g2077)) + ((g2742) & (g2595) & (g2669) & (!g2514) & (!g2076) & (g2077)) + ((g2742) & (g2595) & (g2669) & (!g2514) & (g2076) & (!g2077)) + ((g2742) & (g2595) & (g2669) & (g2514) & (!g2076) & (!g2077)) + ((g2742) & (g2595) & (g2669) & (g2514) & (!g2076) & (g2077)) + ((g2742) & (g2595) & (g2669) & (g2514) & (g2076) & (!g2077)) + ((g2742) & (g2595) & (g2669) & (g2514) & (g2076) & (g2077)));
	assign g2744 = (((!g2743) & (!g2427) & (!g2425) & (g2191) & (g2073) & (g2125)) + ((!g2743) & (!g2427) & (g2425) & (!g2191) & (!g2073) & (g2125)) + ((!g2743) & (!g2427) & (g2425) & (g2191) & (!g2073) & (g2125)) + ((!g2743) & (!g2427) & (g2425) & (g2191) & (g2073) & (g2125)) + ((!g2743) & (g2427) & (!g2425) & (!g2191) & (g2073) & (!g2125)) + ((!g2743) & (g2427) & (!g2425) & (g2191) & (g2073) & (!g2125)) + ((!g2743) & (g2427) & (!g2425) & (g2191) & (g2073) & (g2125)) + ((!g2743) & (g2427) & (g2425) & (!g2191) & (!g2073) & (g2125)) + ((!g2743) & (g2427) & (g2425) & (!g2191) & (g2073) & (!g2125)) + ((!g2743) & (g2427) & (g2425) & (g2191) & (!g2073) & (g2125)) + ((!g2743) & (g2427) & (g2425) & (g2191) & (g2073) & (!g2125)) + ((!g2743) & (g2427) & (g2425) & (g2191) & (g2073) & (g2125)) + ((g2743) & (!g2427) & (!g2425) & (!g2191) & (!g2073) & (!g2125)) + ((g2743) & (!g2427) & (!g2425) & (g2191) & (!g2073) & (!g2125)) + ((g2743) & (!g2427) & (!g2425) & (g2191) & (g2073) & (g2125)) + ((g2743) & (!g2427) & (g2425) & (!g2191) & (!g2073) & (!g2125)) + ((g2743) & (!g2427) & (g2425) & (!g2191) & (!g2073) & (g2125)) + ((g2743) & (!g2427) & (g2425) & (g2191) & (!g2073) & (!g2125)) + ((g2743) & (!g2427) & (g2425) & (g2191) & (!g2073) & (g2125)) + ((g2743) & (!g2427) & (g2425) & (g2191) & (g2073) & (g2125)) + ((g2743) & (g2427) & (!g2425) & (!g2191) & (!g2073) & (!g2125)) + ((g2743) & (g2427) & (!g2425) & (!g2191) & (g2073) & (!g2125)) + ((g2743) & (g2427) & (!g2425) & (g2191) & (!g2073) & (!g2125)) + ((g2743) & (g2427) & (!g2425) & (g2191) & (g2073) & (!g2125)) + ((g2743) & (g2427) & (!g2425) & (g2191) & (g2073) & (g2125)) + ((g2743) & (g2427) & (g2425) & (!g2191) & (!g2073) & (!g2125)) + ((g2743) & (g2427) & (g2425) & (!g2191) & (!g2073) & (g2125)) + ((g2743) & (g2427) & (g2425) & (!g2191) & (g2073) & (!g2125)) + ((g2743) & (g2427) & (g2425) & (g2191) & (!g2073) & (!g2125)) + ((g2743) & (g2427) & (g2425) & (g2191) & (!g2073) & (g2125)) + ((g2743) & (g2427) & (g2425) & (g2191) & (g2073) & (!g2125)) + ((g2743) & (g2427) & (g2425) & (g2191) & (g2073) & (g2125)));
	assign g2745 = (((!g2090) & (!g2734) & (!g2124) & (!g2264) & (!g3313) & (g2744)) + ((!g2090) & (!g2734) & (!g2124) & (!g2264) & (g3313) & (g2744)) + ((!g2090) & (!g2734) & (!g2124) & (g2264) & (g3313) & (!g2744)) + ((!g2090) & (!g2734) & (!g2124) & (g2264) & (g3313) & (g2744)) + ((!g2090) & (g2734) & (!g2124) & (!g2264) & (!g3313) & (g2744)) + ((!g2090) & (g2734) & (!g2124) & (!g2264) & (g3313) & (g2744)) + ((!g2090) & (g2734) & (!g2124) & (g2264) & (g3313) & (!g2744)) + ((!g2090) & (g2734) & (!g2124) & (g2264) & (g3313) & (g2744)) + ((!g2090) & (g2734) & (g2124) & (!g2264) & (!g3313) & (!g2744)) + ((!g2090) & (g2734) & (g2124) & (!g2264) & (!g3313) & (g2744)) + ((!g2090) & (g2734) & (g2124) & (!g2264) & (g3313) & (!g2744)) + ((!g2090) & (g2734) & (g2124) & (!g2264) & (g3313) & (g2744)) + ((!g2090) & (g2734) & (g2124) & (g2264) & (!g3313) & (!g2744)) + ((!g2090) & (g2734) & (g2124) & (g2264) & (!g3313) & (g2744)) + ((!g2090) & (g2734) & (g2124) & (g2264) & (g3313) & (!g2744)) + ((!g2090) & (g2734) & (g2124) & (g2264) & (g3313) & (g2744)) + ((g2090) & (!g2734) & (!g2124) & (!g2264) & (!g3313) & (g2744)) + ((g2090) & (!g2734) & (!g2124) & (!g2264) & (g3313) & (g2744)) + ((g2090) & (!g2734) & (!g2124) & (g2264) & (g3313) & (!g2744)) + ((g2090) & (!g2734) & (!g2124) & (g2264) & (g3313) & (g2744)) + ((g2090) & (!g2734) & (g2124) & (!g2264) & (!g3313) & (!g2744)) + ((g2090) & (!g2734) & (g2124) & (!g2264) & (!g3313) & (g2744)) + ((g2090) & (!g2734) & (g2124) & (!g2264) & (g3313) & (!g2744)) + ((g2090) & (!g2734) & (g2124) & (!g2264) & (g3313) & (g2744)) + ((g2090) & (!g2734) & (g2124) & (g2264) & (!g3313) & (!g2744)) + ((g2090) & (!g2734) & (g2124) & (g2264) & (!g3313) & (g2744)) + ((g2090) & (!g2734) & (g2124) & (g2264) & (g3313) & (!g2744)) + ((g2090) & (!g2734) & (g2124) & (g2264) & (g3313) & (g2744)) + ((g2090) & (g2734) & (!g2124) & (!g2264) & (!g3313) & (g2744)) + ((g2090) & (g2734) & (!g2124) & (!g2264) & (g3313) & (g2744)) + ((g2090) & (g2734) & (!g2124) & (g2264) & (g3313) & (!g2744)) + ((g2090) & (g2734) & (!g2124) & (g2264) & (g3313) & (g2744)) + ((g2090) & (g2734) & (g2124) & (!g2264) & (!g3313) & (!g2744)) + ((g2090) & (g2734) & (g2124) & (!g2264) & (!g3313) & (g2744)) + ((g2090) & (g2734) & (g2124) & (!g2264) & (g3313) & (!g2744)) + ((g2090) & (g2734) & (g2124) & (!g2264) & (g3313) & (g2744)));
	assign g2746 = (((!g1320) & (!sk[54]) & (g2727) & (!g1365)) + ((!g1320) & (!sk[54]) & (g2727) & (g1365)) + ((!g1320) & (sk[54]) & (!g2727) & (g1365)) + ((!g1320) & (sk[54]) & (g2727) & (g1365)) + ((g1320) & (!sk[54]) & (!g2727) & (!g1365)) + ((g1320) & (!sk[54]) & (!g2727) & (g1365)) + ((g1320) & (!sk[54]) & (g2727) & (!g1365)) + ((g1320) & (!sk[54]) & (g2727) & (g1365)) + ((g1320) & (sk[54]) & (!g2727) & (g1365)) + ((g1320) & (sk[54]) & (g2727) & (!g1365)));
	assign g2747 = (((!g108) & (!g110) & (g2585) & (!g1320) & (!g2729) & (g1365)) + ((!g108) & (!g110) & (g2585) & (!g1320) & (g2729) & (g1365)) + ((!g108) & (!g110) & (g2585) & (g1320) & (!g2729) & (!g1365)) + ((!g108) & (!g110) & (g2585) & (g1320) & (g2729) & (g1365)) + ((!g108) & (g110) & (g2585) & (!g1320) & (!g2729) & (!g1365)) + ((!g108) & (g110) & (g2585) & (!g1320) & (g2729) & (!g1365)) + ((!g108) & (g110) & (g2585) & (g1320) & (!g2729) & (g1365)) + ((!g108) & (g110) & (g2585) & (g1320) & (g2729) & (!g1365)) + ((g108) & (!g110) & (g2585) & (!g1320) & (!g2729) & (!g1365)) + ((g108) & (!g110) & (g2585) & (!g1320) & (g2729) & (g1365)) + ((g108) & (!g110) & (g2585) & (g1320) & (!g2729) & (!g1365)) + ((g108) & (!g110) & (g2585) & (g1320) & (g2729) & (!g1365)) + ((g108) & (g110) & (g2585) & (!g1320) & (!g2729) & (g1365)) + ((g108) & (g110) & (g2585) & (!g1320) & (g2729) & (!g1365)) + ((g108) & (g110) & (g2585) & (g1320) & (!g2729) & (g1365)) + ((g108) & (g110) & (g2585) & (g1320) & (g2729) & (g1365)));
	assign g5050 = (((!g2921) & (!sk[56]) & (g3161) & (!g2748)) + ((!g2921) & (!sk[56]) & (g3161) & (g2748)) + ((!g2921) & (sk[56]) & (!g3161) & (g2748)) + ((!g2921) & (sk[56]) & (g3161) & (g2748)) + ((g2921) & (!sk[56]) & (!g3161) & (!g2748)) + ((g2921) & (!sk[56]) & (!g3161) & (g2748)) + ((g2921) & (!sk[56]) & (g3161) & (!g2748)) + ((g2921) & (!sk[56]) & (g3161) & (g2748)) + ((g2921) & (sk[56]) & (g3161) & (!g2748)) + ((g2921) & (sk[56]) & (g3161) & (g2748)));
	assign g2749 = (((!sk[57]) & (!g1942) & (!g2033) & (!g2034) & (g2748)) + ((!sk[57]) & (!g1942) & (!g2033) & (g2034) & (g2748)) + ((!sk[57]) & (!g1942) & (g2033) & (!g2034) & (!g2748)) + ((!sk[57]) & (!g1942) & (g2033) & (!g2034) & (g2748)) + ((!sk[57]) & (!g1942) & (g2033) & (g2034) & (!g2748)) + ((!sk[57]) & (!g1942) & (g2033) & (g2034) & (g2748)) + ((!sk[57]) & (g1942) & (!g2033) & (!g2034) & (!g2748)) + ((!sk[57]) & (g1942) & (!g2033) & (!g2034) & (g2748)) + ((!sk[57]) & (g1942) & (!g2033) & (g2034) & (!g2748)) + ((!sk[57]) & (g1942) & (!g2033) & (g2034) & (g2748)) + ((!sk[57]) & (g1942) & (g2033) & (!g2034) & (!g2748)) + ((!sk[57]) & (g1942) & (g2033) & (!g2034) & (g2748)) + ((!sk[57]) & (g1942) & (g2033) & (g2034) & (!g2748)) + ((!sk[57]) & (g1942) & (g2033) & (g2034) & (g2748)) + ((sk[57]) & (!g1942) & (!g2033) & (!g2034) & (g2748)) + ((sk[57]) & (g1942) & (!g2033) & (!g2034) & (g2748)) + ((sk[57]) & (g1942) & (!g2033) & (g2034) & (!g2748)) + ((sk[57]) & (g1942) & (!g2033) & (g2034) & (g2748)));
	assign g2750 = (((g2329) & (!g2029) & (g2408) & (!g2746) & (!g2747) & (g2749)) + ((g2329) & (!g2029) & (g2408) & (!g2746) & (g2747) & (!g2749)) + ((g2329) & (!g2029) & (g2408) & (!g2746) & (g2747) & (g2749)) + ((g2329) & (!g2029) & (g2408) & (g2746) & (!g2747) & (g2749)) + ((g2329) & (!g2029) & (g2408) & (g2746) & (g2747) & (!g2749)) + ((g2329) & (!g2029) & (g2408) & (g2746) & (g2747) & (g2749)) + ((g2329) & (g2029) & (g2408) & (g2746) & (!g2747) & (!g2749)) + ((g2329) & (g2029) & (g2408) & (g2746) & (!g2747) & (g2749)) + ((g2329) & (g2029) & (g2408) & (g2746) & (g2747) & (!g2749)) + ((g2329) & (g2029) & (g2408) & (g2746) & (g2747) & (g2749)));
	assign g2752 = (((!g2090) & (!g2091) & (!g2734) & (!g2735) & (!g2736) & (g2751)) + ((!g2090) & (!g2091) & (!g2734) & (!g2735) & (g2736) & (g2751)) + ((!g2090) & (!g2091) & (!g2734) & (g2735) & (!g2736) & (g2751)) + ((!g2090) & (!g2091) & (!g2734) & (g2735) & (g2736) & (g2751)) + ((!g2090) & (!g2091) & (g2734) & (!g2735) & (!g2736) & (g2751)) + ((!g2090) & (!g2091) & (g2734) & (!g2735) & (g2736) & (!g2751)) + ((!g2090) & (!g2091) & (g2734) & (g2735) & (!g2736) & (!g2751)) + ((!g2090) & (!g2091) & (g2734) & (g2735) & (g2736) & (!g2751)) + ((!g2090) & (g2091) & (!g2734) & (!g2735) & (!g2736) & (!g2751)) + ((!g2090) & (g2091) & (!g2734) & (!g2735) & (g2736) & (!g2751)) + ((!g2090) & (g2091) & (!g2734) & (g2735) & (!g2736) & (!g2751)) + ((!g2090) & (g2091) & (!g2734) & (g2735) & (g2736) & (!g2751)) + ((!g2090) & (g2091) & (g2734) & (!g2735) & (!g2736) & (!g2751)) + ((!g2090) & (g2091) & (g2734) & (!g2735) & (g2736) & (g2751)) + ((!g2090) & (g2091) & (g2734) & (g2735) & (!g2736) & (g2751)) + ((!g2090) & (g2091) & (g2734) & (g2735) & (g2736) & (g2751)) + ((g2090) & (!g2091) & (!g2734) & (!g2735) & (!g2736) & (g2751)) + ((g2090) & (!g2091) & (!g2734) & (!g2735) & (g2736) & (!g2751)) + ((g2090) & (!g2091) & (!g2734) & (g2735) & (!g2736) & (!g2751)) + ((g2090) & (!g2091) & (!g2734) & (g2735) & (g2736) & (!g2751)) + ((g2090) & (!g2091) & (g2734) & (!g2735) & (!g2736) & (!g2751)) + ((g2090) & (!g2091) & (g2734) & (!g2735) & (g2736) & (!g2751)) + ((g2090) & (!g2091) & (g2734) & (g2735) & (!g2736) & (!g2751)) + ((g2090) & (!g2091) & (g2734) & (g2735) & (g2736) & (!g2751)) + ((g2090) & (g2091) & (!g2734) & (!g2735) & (!g2736) & (!g2751)) + ((g2090) & (g2091) & (!g2734) & (!g2735) & (g2736) & (g2751)) + ((g2090) & (g2091) & (!g2734) & (g2735) & (!g2736) & (g2751)) + ((g2090) & (g2091) & (!g2734) & (g2735) & (g2736) & (g2751)) + ((g2090) & (g2091) & (g2734) & (!g2735) & (!g2736) & (g2751)) + ((g2090) & (g2091) & (g2734) & (!g2735) & (g2736) & (g2751)) + ((g2090) & (g2091) & (g2734) & (g2735) & (!g2736) & (g2751)) + ((g2090) & (g2091) & (g2734) & (g2735) & (g2736) & (g2751)));
	assign g2753 = (((!g2739) & (!sk[60]) & (g2740)) + ((!g2739) & (sk[60]) & (g2740)) + ((g2739) & (!sk[60]) & (g2740)) + ((g2739) & (sk[60]) & (!g2740)));
	assign g2754 = (((!g2702) & (!g2703) & (!g2704) & (g2720) & (g2721) & (g2753)) + ((!g2702) & (!g2703) & (g2704) & (!g2720) & (g2721) & (g2753)) + ((!g2702) & (!g2703) & (g2704) & (g2720) & (!g2721) & (g2753)) + ((!g2702) & (!g2703) & (g2704) & (g2720) & (g2721) & (g2753)) + ((!g2702) & (g2703) & (!g2704) & (!g2720) & (g2721) & (g2753)) + ((!g2702) & (g2703) & (!g2704) & (g2720) & (!g2721) & (g2753)) + ((!g2702) & (g2703) & (!g2704) & (g2720) & (g2721) & (g2753)) + ((!g2702) & (g2703) & (g2704) & (!g2720) & (g2721) & (g2753)) + ((!g2702) & (g2703) & (g2704) & (g2720) & (!g2721) & (g2753)) + ((!g2702) & (g2703) & (g2704) & (g2720) & (g2721) & (g2753)) + ((g2702) & (!g2703) & (!g2704) & (g2720) & (g2721) & (g2753)) + ((g2702) & (!g2703) & (g2704) & (g2720) & (g2721) & (g2753)) + ((g2702) & (g2703) & (!g2704) & (g2720) & (g2721) & (g2753)) + ((g2702) & (g2703) & (g2704) & (!g2720) & (g2721) & (g2753)) + ((g2702) & (g2703) & (g2704) & (g2720) & (!g2721) & (g2753)) + ((g2702) & (g2703) & (g2704) & (g2720) & (g2721) & (g2753)));
	assign g2755 = (((!sk[62]) & (!g2739) & (g2740)) + ((!sk[62]) & (g2739) & (g2740)) + ((sk[62]) & (g2739) & (g2740)));
	assign g2756 = (((!g2734) & (!sk[63]) & (g2090)) + ((!g2734) & (sk[63]) & (g2090)) + ((g2734) & (!sk[63]) & (g2090)));
	assign g2757 = (((!g2751) & (!sk[64]) & (g2091)) + ((!g2751) & (sk[64]) & (!g2091)) + ((g2751) & (!sk[64]) & (g2091)) + ((g2751) & (sk[64]) & (g2091)));
	assign g2758 = (((!g2754) & (!sk[65]) & (!g2755) & (!g2756) & (g2757)) + ((!g2754) & (!sk[65]) & (!g2755) & (g2756) & (g2757)) + ((!g2754) & (!sk[65]) & (g2755) & (!g2756) & (!g2757)) + ((!g2754) & (!sk[65]) & (g2755) & (!g2756) & (g2757)) + ((!g2754) & (!sk[65]) & (g2755) & (g2756) & (!g2757)) + ((!g2754) & (!sk[65]) & (g2755) & (g2756) & (g2757)) + ((!g2754) & (sk[65]) & (!g2755) & (!g2756) & (g2757)) + ((!g2754) & (sk[65]) & (!g2755) & (g2756) & (!g2757)) + ((!g2754) & (sk[65]) & (g2755) & (!g2756) & (!g2757)) + ((!g2754) & (sk[65]) & (g2755) & (g2756) & (g2757)) + ((g2754) & (!sk[65]) & (!g2755) & (!g2756) & (!g2757)) + ((g2754) & (!sk[65]) & (!g2755) & (!g2756) & (g2757)) + ((g2754) & (!sk[65]) & (!g2755) & (g2756) & (!g2757)) + ((g2754) & (!sk[65]) & (!g2755) & (g2756) & (g2757)) + ((g2754) & (!sk[65]) & (g2755) & (!g2756) & (!g2757)) + ((g2754) & (!sk[65]) & (g2755) & (!g2756) & (g2757)) + ((g2754) & (!sk[65]) & (g2755) & (g2756) & (!g2757)) + ((g2754) & (!sk[65]) & (g2755) & (g2756) & (g2757)) + ((g2754) & (sk[65]) & (!g2755) & (!g2756) & (!g2757)) + ((g2754) & (sk[65]) & (!g2755) & (g2756) & (g2757)) + ((g2754) & (sk[65]) & (g2755) & (!g2756) & (!g2757)) + ((g2754) & (sk[65]) & (g2755) & (g2756) & (g2757)));
	assign g2759 = (((!g2091) & (!sk[66]) & (g2751)) + ((g2091) & (!sk[66]) & (g2751)) + ((g2091) & (sk[66]) & (g2751)));
	assign g2760 = (((!g2091) & (!g2090) & (!g2089) & (g2088) & (g2071) & (g2074)) + ((!g2091) & (!g2090) & (g2089) & (!g2088) & (!g2071) & (g2074)) + ((!g2091) & (!g2090) & (g2089) & (g2088) & (!g2071) & (g2074)) + ((!g2091) & (!g2090) & (g2089) & (g2088) & (g2071) & (g2074)) + ((!g2091) & (g2090) & (!g2089) & (!g2088) & (g2071) & (!g2074)) + ((!g2091) & (g2090) & (!g2089) & (g2088) & (g2071) & (!g2074)) + ((!g2091) & (g2090) & (!g2089) & (g2088) & (g2071) & (g2074)) + ((!g2091) & (g2090) & (g2089) & (!g2088) & (!g2071) & (g2074)) + ((!g2091) & (g2090) & (g2089) & (!g2088) & (g2071) & (!g2074)) + ((!g2091) & (g2090) & (g2089) & (g2088) & (!g2071) & (g2074)) + ((!g2091) & (g2090) & (g2089) & (g2088) & (g2071) & (!g2074)) + ((!g2091) & (g2090) & (g2089) & (g2088) & (g2071) & (g2074)) + ((g2091) & (!g2090) & (!g2089) & (!g2088) & (!g2071) & (!g2074)) + ((g2091) & (!g2090) & (!g2089) & (g2088) & (!g2071) & (!g2074)) + ((g2091) & (!g2090) & (!g2089) & (g2088) & (g2071) & (g2074)) + ((g2091) & (!g2090) & (g2089) & (!g2088) & (!g2071) & (!g2074)) + ((g2091) & (!g2090) & (g2089) & (!g2088) & (!g2071) & (g2074)) + ((g2091) & (!g2090) & (g2089) & (g2088) & (!g2071) & (!g2074)) + ((g2091) & (!g2090) & (g2089) & (g2088) & (!g2071) & (g2074)) + ((g2091) & (!g2090) & (g2089) & (g2088) & (g2071) & (g2074)) + ((g2091) & (g2090) & (!g2089) & (!g2088) & (!g2071) & (!g2074)) + ((g2091) & (g2090) & (!g2089) & (!g2088) & (g2071) & (!g2074)) + ((g2091) & (g2090) & (!g2089) & (g2088) & (!g2071) & (!g2074)) + ((g2091) & (g2090) & (!g2089) & (g2088) & (g2071) & (!g2074)) + ((g2091) & (g2090) & (!g2089) & (g2088) & (g2071) & (g2074)) + ((g2091) & (g2090) & (g2089) & (!g2088) & (!g2071) & (!g2074)) + ((g2091) & (g2090) & (g2089) & (!g2088) & (!g2071) & (g2074)) + ((g2091) & (g2090) & (g2089) & (!g2088) & (g2071) & (!g2074)) + ((g2091) & (g2090) & (g2089) & (g2088) & (!g2071) & (!g2074)) + ((g2091) & (g2090) & (g2089) & (g2088) & (!g2071) & (g2074)) + ((g2091) & (g2090) & (g2089) & (g2088) & (g2071) & (!g2074)) + ((g2091) & (g2090) & (g2089) & (g2088) & (g2071) & (g2074)));
	assign g2761 = (((!g2760) & (!g2615) & (!g2687) & (g2536) & (g2076) & (g2077)) + ((!g2760) & (!g2615) & (g2687) & (!g2536) & (!g2076) & (g2077)) + ((!g2760) & (!g2615) & (g2687) & (g2536) & (!g2076) & (g2077)) + ((!g2760) & (!g2615) & (g2687) & (g2536) & (g2076) & (g2077)) + ((!g2760) & (g2615) & (!g2687) & (!g2536) & (g2076) & (!g2077)) + ((!g2760) & (g2615) & (!g2687) & (g2536) & (g2076) & (!g2077)) + ((!g2760) & (g2615) & (!g2687) & (g2536) & (g2076) & (g2077)) + ((!g2760) & (g2615) & (g2687) & (!g2536) & (!g2076) & (g2077)) + ((!g2760) & (g2615) & (g2687) & (!g2536) & (g2076) & (!g2077)) + ((!g2760) & (g2615) & (g2687) & (g2536) & (!g2076) & (g2077)) + ((!g2760) & (g2615) & (g2687) & (g2536) & (g2076) & (!g2077)) + ((!g2760) & (g2615) & (g2687) & (g2536) & (g2076) & (g2077)) + ((g2760) & (!g2615) & (!g2687) & (!g2536) & (!g2076) & (!g2077)) + ((g2760) & (!g2615) & (!g2687) & (g2536) & (!g2076) & (!g2077)) + ((g2760) & (!g2615) & (!g2687) & (g2536) & (g2076) & (g2077)) + ((g2760) & (!g2615) & (g2687) & (!g2536) & (!g2076) & (!g2077)) + ((g2760) & (!g2615) & (g2687) & (!g2536) & (!g2076) & (g2077)) + ((g2760) & (!g2615) & (g2687) & (g2536) & (!g2076) & (!g2077)) + ((g2760) & (!g2615) & (g2687) & (g2536) & (!g2076) & (g2077)) + ((g2760) & (!g2615) & (g2687) & (g2536) & (g2076) & (g2077)) + ((g2760) & (g2615) & (!g2687) & (!g2536) & (!g2076) & (!g2077)) + ((g2760) & (g2615) & (!g2687) & (!g2536) & (g2076) & (!g2077)) + ((g2760) & (g2615) & (!g2687) & (g2536) & (!g2076) & (!g2077)) + ((g2760) & (g2615) & (!g2687) & (g2536) & (g2076) & (!g2077)) + ((g2760) & (g2615) & (!g2687) & (g2536) & (g2076) & (g2077)) + ((g2760) & (g2615) & (g2687) & (!g2536) & (!g2076) & (!g2077)) + ((g2760) & (g2615) & (g2687) & (!g2536) & (!g2076) & (g2077)) + ((g2760) & (g2615) & (g2687) & (!g2536) & (g2076) & (!g2077)) + ((g2760) & (g2615) & (g2687) & (g2536) & (!g2076) & (!g2077)) + ((g2760) & (g2615) & (g2687) & (g2536) & (!g2076) & (g2077)) + ((g2760) & (g2615) & (g2687) & (g2536) & (g2076) & (!g2077)) + ((g2760) & (g2615) & (g2687) & (g2536) & (g2076) & (g2077)));
	assign g2762 = (((!g2761) & (!g2450) & (!g2448) & (g2191) & (g2073) & (g2125)) + ((!g2761) & (!g2450) & (g2448) & (!g2191) & (!g2073) & (g2125)) + ((!g2761) & (!g2450) & (g2448) & (g2191) & (!g2073) & (g2125)) + ((!g2761) & (!g2450) & (g2448) & (g2191) & (g2073) & (g2125)) + ((!g2761) & (g2450) & (!g2448) & (!g2191) & (g2073) & (!g2125)) + ((!g2761) & (g2450) & (!g2448) & (g2191) & (g2073) & (!g2125)) + ((!g2761) & (g2450) & (!g2448) & (g2191) & (g2073) & (g2125)) + ((!g2761) & (g2450) & (g2448) & (!g2191) & (!g2073) & (g2125)) + ((!g2761) & (g2450) & (g2448) & (!g2191) & (g2073) & (!g2125)) + ((!g2761) & (g2450) & (g2448) & (g2191) & (!g2073) & (g2125)) + ((!g2761) & (g2450) & (g2448) & (g2191) & (g2073) & (!g2125)) + ((!g2761) & (g2450) & (g2448) & (g2191) & (g2073) & (g2125)) + ((g2761) & (!g2450) & (!g2448) & (!g2191) & (!g2073) & (!g2125)) + ((g2761) & (!g2450) & (!g2448) & (g2191) & (!g2073) & (!g2125)) + ((g2761) & (!g2450) & (!g2448) & (g2191) & (g2073) & (g2125)) + ((g2761) & (!g2450) & (g2448) & (!g2191) & (!g2073) & (!g2125)) + ((g2761) & (!g2450) & (g2448) & (!g2191) & (!g2073) & (g2125)) + ((g2761) & (!g2450) & (g2448) & (g2191) & (!g2073) & (!g2125)) + ((g2761) & (!g2450) & (g2448) & (g2191) & (!g2073) & (g2125)) + ((g2761) & (!g2450) & (g2448) & (g2191) & (g2073) & (g2125)) + ((g2761) & (g2450) & (!g2448) & (!g2191) & (!g2073) & (!g2125)) + ((g2761) & (g2450) & (!g2448) & (!g2191) & (g2073) & (!g2125)) + ((g2761) & (g2450) & (!g2448) & (g2191) & (!g2073) & (!g2125)) + ((g2761) & (g2450) & (!g2448) & (g2191) & (g2073) & (!g2125)) + ((g2761) & (g2450) & (!g2448) & (g2191) & (g2073) & (g2125)) + ((g2761) & (g2450) & (g2448) & (!g2191) & (!g2073) & (!g2125)) + ((g2761) & (g2450) & (g2448) & (!g2191) & (!g2073) & (g2125)) + ((g2761) & (g2450) & (g2448) & (!g2191) & (g2073) & (!g2125)) + ((g2761) & (g2450) & (g2448) & (g2191) & (!g2073) & (!g2125)) + ((g2761) & (g2450) & (g2448) & (g2191) & (!g2073) & (g2125)) + ((g2761) & (g2450) & (g2448) & (g2191) & (g2073) & (!g2125)) + ((g2761) & (g2450) & (g2448) & (g2191) & (g2073) & (g2125)));
	assign g2763 = (((!g2091) & (!g2751) & (!g2124) & (!g2264) & (!g3289) & (g2762)) + ((!g2091) & (!g2751) & (!g2124) & (!g2264) & (g3289) & (g2762)) + ((!g2091) & (!g2751) & (!g2124) & (g2264) & (g3289) & (!g2762)) + ((!g2091) & (!g2751) & (!g2124) & (g2264) & (g3289) & (g2762)) + ((!g2091) & (g2751) & (!g2124) & (!g2264) & (!g3289) & (g2762)) + ((!g2091) & (g2751) & (!g2124) & (!g2264) & (g3289) & (g2762)) + ((!g2091) & (g2751) & (!g2124) & (g2264) & (g3289) & (!g2762)) + ((!g2091) & (g2751) & (!g2124) & (g2264) & (g3289) & (g2762)) + ((!g2091) & (g2751) & (g2124) & (!g2264) & (!g3289) & (!g2762)) + ((!g2091) & (g2751) & (g2124) & (!g2264) & (!g3289) & (g2762)) + ((!g2091) & (g2751) & (g2124) & (!g2264) & (g3289) & (!g2762)) + ((!g2091) & (g2751) & (g2124) & (!g2264) & (g3289) & (g2762)) + ((!g2091) & (g2751) & (g2124) & (g2264) & (!g3289) & (!g2762)) + ((!g2091) & (g2751) & (g2124) & (g2264) & (!g3289) & (g2762)) + ((!g2091) & (g2751) & (g2124) & (g2264) & (g3289) & (!g2762)) + ((!g2091) & (g2751) & (g2124) & (g2264) & (g3289) & (g2762)) + ((g2091) & (!g2751) & (!g2124) & (!g2264) & (!g3289) & (g2762)) + ((g2091) & (!g2751) & (!g2124) & (!g2264) & (g3289) & (g2762)) + ((g2091) & (!g2751) & (!g2124) & (g2264) & (g3289) & (!g2762)) + ((g2091) & (!g2751) & (!g2124) & (g2264) & (g3289) & (g2762)) + ((g2091) & (!g2751) & (g2124) & (!g2264) & (!g3289) & (!g2762)) + ((g2091) & (!g2751) & (g2124) & (!g2264) & (!g3289) & (g2762)) + ((g2091) & (!g2751) & (g2124) & (!g2264) & (g3289) & (!g2762)) + ((g2091) & (!g2751) & (g2124) & (!g2264) & (g3289) & (g2762)) + ((g2091) & (!g2751) & (g2124) & (g2264) & (!g3289) & (!g2762)) + ((g2091) & (!g2751) & (g2124) & (g2264) & (!g3289) & (g2762)) + ((g2091) & (!g2751) & (g2124) & (g2264) & (g3289) & (!g2762)) + ((g2091) & (!g2751) & (g2124) & (g2264) & (g3289) & (g2762)) + ((g2091) & (g2751) & (!g2124) & (!g2264) & (!g3289) & (g2762)) + ((g2091) & (g2751) & (!g2124) & (!g2264) & (g3289) & (g2762)) + ((g2091) & (g2751) & (!g2124) & (g2264) & (g3289) & (!g2762)) + ((g2091) & (g2751) & (!g2124) & (g2264) & (g3289) & (g2762)) + ((g2091) & (g2751) & (g2124) & (!g2264) & (!g3289) & (!g2762)) + ((g2091) & (g2751) & (g2124) & (!g2264) & (!g3289) & (g2762)) + ((g2091) & (g2751) & (g2124) & (!g2264) & (g3289) & (!g2762)) + ((g2091) & (g2751) & (g2124) & (!g2264) & (g3289) & (g2762)));
	assign g2764 = (((!g1320) & (!sk[71]) & (!g2727) & (!g1365) & (g1410)) + ((!g1320) & (!sk[71]) & (!g2727) & (g1365) & (g1410)) + ((!g1320) & (!sk[71]) & (g2727) & (!g1365) & (!g1410)) + ((!g1320) & (!sk[71]) & (g2727) & (!g1365) & (g1410)) + ((!g1320) & (!sk[71]) & (g2727) & (g1365) & (!g1410)) + ((!g1320) & (!sk[71]) & (g2727) & (g1365) & (g1410)) + ((!g1320) & (sk[71]) & (!g2727) & (!g1365) & (g1410)) + ((!g1320) & (sk[71]) & (!g2727) & (g1365) & (g1410)) + ((!g1320) & (sk[71]) & (g2727) & (!g1365) & (g1410)) + ((!g1320) & (sk[71]) & (g2727) & (g1365) & (g1410)) + ((g1320) & (!sk[71]) & (!g2727) & (!g1365) & (!g1410)) + ((g1320) & (!sk[71]) & (!g2727) & (!g1365) & (g1410)) + ((g1320) & (!sk[71]) & (!g2727) & (g1365) & (!g1410)) + ((g1320) & (!sk[71]) & (!g2727) & (g1365) & (g1410)) + ((g1320) & (!sk[71]) & (g2727) & (!g1365) & (!g1410)) + ((g1320) & (!sk[71]) & (g2727) & (!g1365) & (g1410)) + ((g1320) & (!sk[71]) & (g2727) & (g1365) & (!g1410)) + ((g1320) & (!sk[71]) & (g2727) & (g1365) & (g1410)) + ((g1320) & (sk[71]) & (!g2727) & (!g1365) & (g1410)) + ((g1320) & (sk[71]) & (!g2727) & (g1365) & (g1410)) + ((g1320) & (sk[71]) & (g2727) & (!g1365) & (g1410)) + ((g1320) & (sk[71]) & (g2727) & (g1365) & (!g1410)));
	assign g2765 = (((!g108) & (!g110) & (!sk[72]) & (!g1320) & (g2729) & (!g1365)) + ((!g108) & (!g110) & (!sk[72]) & (!g1320) & (g2729) & (g1365)) + ((!g108) & (!g110) & (!sk[72]) & (g1320) & (!g2729) & (!g1365)) + ((!g108) & (!g110) & (!sk[72]) & (g1320) & (!g2729) & (g1365)) + ((!g108) & (!g110) & (!sk[72]) & (g1320) & (g2729) & (!g1365)) + ((!g108) & (!g110) & (!sk[72]) & (g1320) & (g2729) & (g1365)) + ((!g108) & (!g110) & (sk[72]) & (g1320) & (!g2729) & (g1365)) + ((!g108) & (g110) & (!sk[72]) & (!g1320) & (g2729) & (!g1365)) + ((!g108) & (g110) & (!sk[72]) & (!g1320) & (g2729) & (g1365)) + ((!g108) & (g110) & (!sk[72]) & (g1320) & (!g2729) & (!g1365)) + ((!g108) & (g110) & (!sk[72]) & (g1320) & (!g2729) & (g1365)) + ((!g108) & (g110) & (!sk[72]) & (g1320) & (g2729) & (!g1365)) + ((!g108) & (g110) & (!sk[72]) & (g1320) & (g2729) & (g1365)) + ((!g108) & (g110) & (sk[72]) & (!g1320) & (!g2729) & (g1365)) + ((!g108) & (g110) & (sk[72]) & (!g1320) & (g2729) & (g1365)) + ((!g108) & (g110) & (sk[72]) & (g1320) & (!g2729) & (!g1365)) + ((!g108) & (g110) & (sk[72]) & (g1320) & (!g2729) & (g1365)) + ((!g108) & (g110) & (sk[72]) & (g1320) & (g2729) & (g1365)) + ((g108) & (!g110) & (!sk[72]) & (!g1320) & (!g2729) & (!g1365)) + ((g108) & (!g110) & (!sk[72]) & (!g1320) & (!g2729) & (g1365)) + ((g108) & (!g110) & (!sk[72]) & (!g1320) & (g2729) & (!g1365)) + ((g108) & (!g110) & (!sk[72]) & (!g1320) & (g2729) & (g1365)) + ((g108) & (!g110) & (!sk[72]) & (g1320) & (!g2729) & (!g1365)) + ((g108) & (!g110) & (!sk[72]) & (g1320) & (!g2729) & (g1365)) + ((g108) & (!g110) & (!sk[72]) & (g1320) & (g2729) & (!g1365)) + ((g108) & (!g110) & (!sk[72]) & (g1320) & (g2729) & (g1365)) + ((g108) & (!g110) & (sk[72]) & (!g1320) & (!g2729) & (g1365)) + ((g108) & (!g110) & (sk[72]) & (g1320) & (!g2729) & (g1365)) + ((g108) & (!g110) & (sk[72]) & (g1320) & (g2729) & (g1365)) + ((g108) & (g110) & (!sk[72]) & (!g1320) & (!g2729) & (!g1365)) + ((g108) & (g110) & (!sk[72]) & (!g1320) & (!g2729) & (g1365)) + ((g108) & (g110) & (!sk[72]) & (!g1320) & (g2729) & (!g1365)) + ((g108) & (g110) & (!sk[72]) & (!g1320) & (g2729) & (g1365)) + ((g108) & (g110) & (!sk[72]) & (g1320) & (!g2729) & (!g1365)) + ((g108) & (g110) & (!sk[72]) & (g1320) & (!g2729) & (g1365)) + ((g108) & (g110) & (!sk[72]) & (g1320) & (g2729) & (!g1365)) + ((g108) & (g110) & (!sk[72]) & (g1320) & (g2729) & (g1365)) + ((g108) & (g110) & (sk[72]) & (!g1320) & (!g2729) & (!g1365)) + ((g108) & (g110) & (sk[72]) & (!g1320) & (!g2729) & (g1365)) + ((g108) & (g110) & (sk[72]) & (!g1320) & (g2729) & (g1365)) + ((g108) & (g110) & (sk[72]) & (g1320) & (!g2729) & (!g1365)) + ((g108) & (g110) & (sk[72]) & (g1320) & (!g2729) & (g1365)) + ((g108) & (g110) & (sk[72]) & (g1320) & (g2729) & (!g1365)) + ((g108) & (g110) & (sk[72]) & (g1320) & (g2729) & (g1365)));
	assign g2766 = (((!sk[73]) & (!g107) & (!g2585) & (!g1410) & (g2765)) + ((!sk[73]) & (!g107) & (!g2585) & (g1410) & (g2765)) + ((!sk[73]) & (!g107) & (g2585) & (!g1410) & (!g2765)) + ((!sk[73]) & (!g107) & (g2585) & (!g1410) & (g2765)) + ((!sk[73]) & (!g107) & (g2585) & (g1410) & (!g2765)) + ((!sk[73]) & (!g107) & (g2585) & (g1410) & (g2765)) + ((!sk[73]) & (g107) & (!g2585) & (!g1410) & (!g2765)) + ((!sk[73]) & (g107) & (!g2585) & (!g1410) & (g2765)) + ((!sk[73]) & (g107) & (!g2585) & (g1410) & (!g2765)) + ((!sk[73]) & (g107) & (!g2585) & (g1410) & (g2765)) + ((!sk[73]) & (g107) & (g2585) & (!g1410) & (!g2765)) + ((!sk[73]) & (g107) & (g2585) & (!g1410) & (g2765)) + ((!sk[73]) & (g107) & (g2585) & (g1410) & (!g2765)) + ((!sk[73]) & (g107) & (g2585) & (g1410) & (g2765)) + ((sk[73]) & (!g107) & (g2585) & (!g1410) & (g2765)) + ((sk[73]) & (!g107) & (g2585) & (g1410) & (!g2765)) + ((sk[73]) & (g107) & (g2585) & (!g1410) & (!g2765)) + ((sk[73]) & (g107) & (g2585) & (g1410) & (g2765)));
	assign g5051 = (((!g2921) & (!sk[74]) & (g3148) & (!g2767)) + ((!g2921) & (!sk[74]) & (g3148) & (g2767)) + ((!g2921) & (sk[74]) & (!g3148) & (g2767)) + ((!g2921) & (sk[74]) & (g3148) & (g2767)) + ((g2921) & (!sk[74]) & (!g3148) & (!g2767)) + ((g2921) & (!sk[74]) & (!g3148) & (g2767)) + ((g2921) & (!sk[74]) & (g3148) & (!g2767)) + ((g2921) & (!sk[74]) & (g3148) & (g2767)) + ((g2921) & (sk[74]) & (g3148) & (!g2767)) + ((g2921) & (sk[74]) & (g3148) & (g2767)));
	assign g2768 = (((!g1955) & (!g2033) & (!g2034) & (!sk[75]) & (g2767)) + ((!g1955) & (!g2033) & (!g2034) & (sk[75]) & (g2767)) + ((!g1955) & (!g2033) & (g2034) & (!sk[75]) & (g2767)) + ((!g1955) & (g2033) & (!g2034) & (!sk[75]) & (!g2767)) + ((!g1955) & (g2033) & (!g2034) & (!sk[75]) & (g2767)) + ((!g1955) & (g2033) & (g2034) & (!sk[75]) & (!g2767)) + ((!g1955) & (g2033) & (g2034) & (!sk[75]) & (g2767)) + ((g1955) & (!g2033) & (!g2034) & (!sk[75]) & (!g2767)) + ((g1955) & (!g2033) & (!g2034) & (!sk[75]) & (g2767)) + ((g1955) & (!g2033) & (!g2034) & (sk[75]) & (g2767)) + ((g1955) & (!g2033) & (g2034) & (!sk[75]) & (!g2767)) + ((g1955) & (!g2033) & (g2034) & (!sk[75]) & (g2767)) + ((g1955) & (!g2033) & (g2034) & (sk[75]) & (!g2767)) + ((g1955) & (!g2033) & (g2034) & (sk[75]) & (g2767)) + ((g1955) & (g2033) & (!g2034) & (!sk[75]) & (!g2767)) + ((g1955) & (g2033) & (!g2034) & (!sk[75]) & (g2767)) + ((g1955) & (g2033) & (g2034) & (!sk[75]) & (!g2767)) + ((g1955) & (g2033) & (g2034) & (!sk[75]) & (g2767)));
	assign g2769 = (((g2329) & (!g2029) & (g2408) & (!g2764) & (!g2766) & (g2768)) + ((g2329) & (!g2029) & (g2408) & (!g2764) & (g2766) & (!g2768)) + ((g2329) & (!g2029) & (g2408) & (!g2764) & (g2766) & (g2768)) + ((g2329) & (!g2029) & (g2408) & (g2764) & (!g2766) & (g2768)) + ((g2329) & (!g2029) & (g2408) & (g2764) & (g2766) & (!g2768)) + ((g2329) & (!g2029) & (g2408) & (g2764) & (g2766) & (g2768)) + ((g2329) & (g2029) & (g2408) & (g2764) & (!g2766) & (!g2768)) + ((g2329) & (g2029) & (g2408) & (g2764) & (!g2766) & (g2768)) + ((g2329) & (g2029) & (g2408) & (g2764) & (g2766) & (!g2768)) + ((g2329) & (g2029) & (g2408) & (g2764) & (g2766) & (g2768)));
	assign g2770 = (((!g2080) & (!sk[77]) & (!g2081) & (!g2124) & (g2125) & (!g2181)) + ((!g2080) & (!sk[77]) & (!g2081) & (!g2124) & (g2125) & (g2181)) + ((!g2080) & (!sk[77]) & (!g2081) & (g2124) & (!g2125) & (!g2181)) + ((!g2080) & (!sk[77]) & (!g2081) & (g2124) & (!g2125) & (g2181)) + ((!g2080) & (!sk[77]) & (!g2081) & (g2124) & (g2125) & (!g2181)) + ((!g2080) & (!sk[77]) & (!g2081) & (g2124) & (g2125) & (g2181)) + ((!g2080) & (!sk[77]) & (g2081) & (!g2124) & (g2125) & (!g2181)) + ((!g2080) & (!sk[77]) & (g2081) & (!g2124) & (g2125) & (g2181)) + ((!g2080) & (!sk[77]) & (g2081) & (g2124) & (!g2125) & (!g2181)) + ((!g2080) & (!sk[77]) & (g2081) & (g2124) & (!g2125) & (g2181)) + ((!g2080) & (!sk[77]) & (g2081) & (g2124) & (g2125) & (!g2181)) + ((!g2080) & (!sk[77]) & (g2081) & (g2124) & (g2125) & (g2181)) + ((!g2080) & (sk[77]) & (!g2081) & (!g2124) & (!g2125) & (!g2181)) + ((!g2080) & (sk[77]) & (!g2081) & (!g2124) & (!g2125) & (g2181)) + ((!g2080) & (sk[77]) & (!g2081) & (g2124) & (g2125) & (!g2181)) + ((!g2080) & (sk[77]) & (!g2081) & (g2124) & (g2125) & (g2181)) + ((!g2080) & (sk[77]) & (g2081) & (!g2124) & (!g2125) & (g2181)) + ((!g2080) & (sk[77]) & (g2081) & (g2124) & (g2125) & (!g2181)) + ((!g2080) & (sk[77]) & (g2081) & (g2124) & (g2125) & (g2181)) + ((g2080) & (!sk[77]) & (!g2081) & (!g2124) & (!g2125) & (!g2181)) + ((g2080) & (!sk[77]) & (!g2081) & (!g2124) & (!g2125) & (g2181)) + ((g2080) & (!sk[77]) & (!g2081) & (!g2124) & (g2125) & (!g2181)) + ((g2080) & (!sk[77]) & (!g2081) & (!g2124) & (g2125) & (g2181)) + ((g2080) & (!sk[77]) & (!g2081) & (g2124) & (!g2125) & (!g2181)) + ((g2080) & (!sk[77]) & (!g2081) & (g2124) & (!g2125) & (g2181)) + ((g2080) & (!sk[77]) & (!g2081) & (g2124) & (g2125) & (!g2181)) + ((g2080) & (!sk[77]) & (!g2081) & (g2124) & (g2125) & (g2181)) + ((g2080) & (!sk[77]) & (g2081) & (!g2124) & (!g2125) & (!g2181)) + ((g2080) & (!sk[77]) & (g2081) & (!g2124) & (!g2125) & (g2181)) + ((g2080) & (!sk[77]) & (g2081) & (!g2124) & (g2125) & (!g2181)) + ((g2080) & (!sk[77]) & (g2081) & (!g2124) & (g2125) & (g2181)) + ((g2080) & (!sk[77]) & (g2081) & (g2124) & (!g2125) & (!g2181)) + ((g2080) & (!sk[77]) & (g2081) & (g2124) & (!g2125) & (g2181)) + ((g2080) & (!sk[77]) & (g2081) & (g2124) & (g2125) & (!g2181)) + ((g2080) & (!sk[77]) & (g2081) & (g2124) & (g2125) & (g2181)) + ((g2080) & (sk[77]) & (!g2081) & (g2124) & (!g2125) & (!g2181)) + ((g2080) & (sk[77]) & (!g2081) & (g2124) & (!g2125) & (g2181)) + ((g2080) & (sk[77]) & (!g2081) & (g2124) & (g2125) & (!g2181)) + ((g2080) & (sk[77]) & (!g2081) & (g2124) & (g2125) & (g2181)) + ((g2080) & (sk[77]) & (g2081) & (g2124) & (!g2125) & (!g2181)) + ((g2080) & (sk[77]) & (g2081) & (g2124) & (!g2125) & (g2181)) + ((g2080) & (sk[77]) & (g2081) & (g2124) & (g2125) & (!g2181)) + ((g2080) & (sk[77]) & (g2081) & (g2124) & (g2125) & (g2181)));
	assign g2772 = (((!g2090) & (!g2091) & (g2734) & (!g2735) & (g2736) & (g2751)) + ((!g2090) & (!g2091) & (g2734) & (g2735) & (!g2736) & (g2751)) + ((!g2090) & (!g2091) & (g2734) & (g2735) & (g2736) & (g2751)) + ((!g2090) & (g2091) & (!g2734) & (!g2735) & (!g2736) & (g2751)) + ((!g2090) & (g2091) & (!g2734) & (!g2735) & (g2736) & (g2751)) + ((!g2090) & (g2091) & (!g2734) & (g2735) & (!g2736) & (g2751)) + ((!g2090) & (g2091) & (!g2734) & (g2735) & (g2736) & (g2751)) + ((!g2090) & (g2091) & (g2734) & (!g2735) & (!g2736) & (g2751)) + ((!g2090) & (g2091) & (g2734) & (!g2735) & (g2736) & (!g2751)) + ((!g2090) & (g2091) & (g2734) & (!g2735) & (g2736) & (g2751)) + ((!g2090) & (g2091) & (g2734) & (g2735) & (!g2736) & (!g2751)) + ((!g2090) & (g2091) & (g2734) & (g2735) & (!g2736) & (g2751)) + ((!g2090) & (g2091) & (g2734) & (g2735) & (g2736) & (!g2751)) + ((!g2090) & (g2091) & (g2734) & (g2735) & (g2736) & (g2751)) + ((g2090) & (!g2091) & (!g2734) & (!g2735) & (g2736) & (g2751)) + ((g2090) & (!g2091) & (!g2734) & (g2735) & (!g2736) & (g2751)) + ((g2090) & (!g2091) & (!g2734) & (g2735) & (g2736) & (g2751)) + ((g2090) & (!g2091) & (g2734) & (!g2735) & (!g2736) & (g2751)) + ((g2090) & (!g2091) & (g2734) & (!g2735) & (g2736) & (g2751)) + ((g2090) & (!g2091) & (g2734) & (g2735) & (!g2736) & (g2751)) + ((g2090) & (!g2091) & (g2734) & (g2735) & (g2736) & (g2751)) + ((g2090) & (g2091) & (!g2734) & (!g2735) & (!g2736) & (g2751)) + ((g2090) & (g2091) & (!g2734) & (!g2735) & (g2736) & (!g2751)) + ((g2090) & (g2091) & (!g2734) & (!g2735) & (g2736) & (g2751)) + ((g2090) & (g2091) & (!g2734) & (g2735) & (!g2736) & (!g2751)) + ((g2090) & (g2091) & (!g2734) & (g2735) & (!g2736) & (g2751)) + ((g2090) & (g2091) & (!g2734) & (g2735) & (g2736) & (!g2751)) + ((g2090) & (g2091) & (!g2734) & (g2735) & (g2736) & (g2751)) + ((g2090) & (g2091) & (g2734) & (!g2735) & (!g2736) & (!g2751)) + ((g2090) & (g2091) & (g2734) & (!g2735) & (!g2736) & (g2751)) + ((g2090) & (g2091) & (g2734) & (!g2735) & (g2736) & (!g2751)) + ((g2090) & (g2091) & (g2734) & (!g2735) & (g2736) & (g2751)) + ((g2090) & (g2091) & (g2734) & (g2735) & (!g2736) & (!g2751)) + ((g2090) & (g2091) & (g2734) & (g2735) & (!g2736) & (g2751)) + ((g2090) & (g2091) & (g2734) & (g2735) & (g2736) & (!g2751)) + ((g2090) & (g2091) & (g2734) & (g2735) & (g2736) & (g2751)));
	assign g2773 = (((!sk[79]) & (!g2098) & (g2771)) + ((!sk[79]) & (g2098) & (g2771)) + ((sk[79]) & (!g2098) & (g2771)) + ((sk[79]) & (g2098) & (!g2771)));
	assign g2774 = (((!sk[80]) & (!g2737) & (!g2738) & (!g2752) & (g2772) & (!g2773)) + ((!sk[80]) & (!g2737) & (!g2738) & (!g2752) & (g2772) & (g2773)) + ((!sk[80]) & (!g2737) & (!g2738) & (g2752) & (!g2772) & (!g2773)) + ((!sk[80]) & (!g2737) & (!g2738) & (g2752) & (!g2772) & (g2773)) + ((!sk[80]) & (!g2737) & (!g2738) & (g2752) & (g2772) & (!g2773)) + ((!sk[80]) & (!g2737) & (!g2738) & (g2752) & (g2772) & (g2773)) + ((!sk[80]) & (!g2737) & (g2738) & (!g2752) & (g2772) & (!g2773)) + ((!sk[80]) & (!g2737) & (g2738) & (!g2752) & (g2772) & (g2773)) + ((!sk[80]) & (!g2737) & (g2738) & (g2752) & (!g2772) & (!g2773)) + ((!sk[80]) & (!g2737) & (g2738) & (g2752) & (!g2772) & (g2773)) + ((!sk[80]) & (!g2737) & (g2738) & (g2752) & (g2772) & (!g2773)) + ((!sk[80]) & (!g2737) & (g2738) & (g2752) & (g2772) & (g2773)) + ((!sk[80]) & (g2737) & (!g2738) & (!g2752) & (!g2772) & (!g2773)) + ((!sk[80]) & (g2737) & (!g2738) & (!g2752) & (!g2772) & (g2773)) + ((!sk[80]) & (g2737) & (!g2738) & (!g2752) & (g2772) & (!g2773)) + ((!sk[80]) & (g2737) & (!g2738) & (!g2752) & (g2772) & (g2773)) + ((!sk[80]) & (g2737) & (!g2738) & (g2752) & (!g2772) & (!g2773)) + ((!sk[80]) & (g2737) & (!g2738) & (g2752) & (!g2772) & (g2773)) + ((!sk[80]) & (g2737) & (!g2738) & (g2752) & (g2772) & (!g2773)) + ((!sk[80]) & (g2737) & (!g2738) & (g2752) & (g2772) & (g2773)) + ((!sk[80]) & (g2737) & (g2738) & (!g2752) & (!g2772) & (!g2773)) + ((!sk[80]) & (g2737) & (g2738) & (!g2752) & (!g2772) & (g2773)) + ((!sk[80]) & (g2737) & (g2738) & (!g2752) & (g2772) & (!g2773)) + ((!sk[80]) & (g2737) & (g2738) & (!g2752) & (g2772) & (g2773)) + ((!sk[80]) & (g2737) & (g2738) & (g2752) & (!g2772) & (!g2773)) + ((!sk[80]) & (g2737) & (g2738) & (g2752) & (!g2772) & (g2773)) + ((!sk[80]) & (g2737) & (g2738) & (g2752) & (g2772) & (!g2773)) + ((!sk[80]) & (g2737) & (g2738) & (g2752) & (g2772) & (g2773)) + ((sk[80]) & (!g2737) & (!g2738) & (!g2752) & (!g2772) & (g2773)) + ((sk[80]) & (!g2737) & (!g2738) & (!g2752) & (g2772) & (!g2773)) + ((sk[80]) & (!g2737) & (!g2738) & (g2752) & (!g2772) & (g2773)) + ((sk[80]) & (!g2737) & (!g2738) & (g2752) & (g2772) & (!g2773)) + ((sk[80]) & (!g2737) & (g2738) & (!g2752) & (!g2772) & (g2773)) + ((sk[80]) & (!g2737) & (g2738) & (!g2752) & (g2772) & (!g2773)) + ((sk[80]) & (!g2737) & (g2738) & (g2752) & (!g2772) & (g2773)) + ((sk[80]) & (!g2737) & (g2738) & (g2752) & (g2772) & (!g2773)) + ((sk[80]) & (g2737) & (!g2738) & (!g2752) & (!g2772) & (g2773)) + ((sk[80]) & (g2737) & (!g2738) & (!g2752) & (g2772) & (!g2773)) + ((sk[80]) & (g2737) & (!g2738) & (g2752) & (!g2772) & (g2773)) + ((sk[80]) & (g2737) & (!g2738) & (g2752) & (g2772) & (!g2773)) + ((sk[80]) & (g2737) & (g2738) & (!g2752) & (!g2772) & (g2773)) + ((sk[80]) & (g2737) & (g2738) & (!g2752) & (g2772) & (!g2773)) + ((sk[80]) & (g2737) & (g2738) & (g2752) & (!g2772) & (!g2773)) + ((sk[80]) & (g2737) & (g2738) & (g2752) & (g2772) & (g2773)));
	assign g2775 = (((!sk[81]) & (!g2751) & (g2091)) + ((!sk[81]) & (g2751) & (g2091)) + ((sk[81]) & (!g2751) & (g2091)));
	assign g2776 = (((!sk[82]) & (!g2771) & (g2098)) + ((!sk[82]) & (g2771) & (g2098)) + ((sk[82]) & (!g2771) & (!g2098)) + ((sk[82]) & (g2771) & (g2098)));
	assign g2777 = (((!g2754) & (!g2755) & (!g2756) & (!g2757) & (!g2775) & (g2776)) + ((!g2754) & (!g2755) & (!g2756) & (!g2757) & (g2775) & (!g2776)) + ((!g2754) & (!g2755) & (!g2756) & (g2757) & (!g2775) & (g2776)) + ((!g2754) & (!g2755) & (!g2756) & (g2757) & (g2775) & (!g2776)) + ((!g2754) & (!g2755) & (g2756) & (!g2757) & (!g2775) & (g2776)) + ((!g2754) & (!g2755) & (g2756) & (!g2757) & (g2775) & (!g2776)) + ((!g2754) & (!g2755) & (g2756) & (g2757) & (!g2775) & (!g2776)) + ((!g2754) & (!g2755) & (g2756) & (g2757) & (g2775) & (g2776)) + ((!g2754) & (g2755) & (!g2756) & (!g2757) & (!g2775) & (g2776)) + ((!g2754) & (g2755) & (!g2756) & (!g2757) & (g2775) & (!g2776)) + ((!g2754) & (g2755) & (!g2756) & (g2757) & (!g2775) & (!g2776)) + ((!g2754) & (g2755) & (!g2756) & (g2757) & (g2775) & (g2776)) + ((!g2754) & (g2755) & (g2756) & (!g2757) & (!g2775) & (!g2776)) + ((!g2754) & (g2755) & (g2756) & (!g2757) & (g2775) & (g2776)) + ((!g2754) & (g2755) & (g2756) & (g2757) & (!g2775) & (!g2776)) + ((!g2754) & (g2755) & (g2756) & (g2757) & (g2775) & (g2776)) + ((g2754) & (!g2755) & (!g2756) & (!g2757) & (!g2775) & (g2776)) + ((g2754) & (!g2755) & (!g2756) & (!g2757) & (g2775) & (!g2776)) + ((g2754) & (!g2755) & (!g2756) & (g2757) & (!g2775) & (!g2776)) + ((g2754) & (!g2755) & (!g2756) & (g2757) & (g2775) & (g2776)) + ((g2754) & (!g2755) & (g2756) & (!g2757) & (!g2775) & (!g2776)) + ((g2754) & (!g2755) & (g2756) & (!g2757) & (g2775) & (g2776)) + ((g2754) & (!g2755) & (g2756) & (g2757) & (!g2775) & (!g2776)) + ((g2754) & (!g2755) & (g2756) & (g2757) & (g2775) & (g2776)) + ((g2754) & (g2755) & (!g2756) & (!g2757) & (!g2775) & (g2776)) + ((g2754) & (g2755) & (!g2756) & (!g2757) & (g2775) & (!g2776)) + ((g2754) & (g2755) & (!g2756) & (g2757) & (!g2775) & (!g2776)) + ((g2754) & (g2755) & (!g2756) & (g2757) & (g2775) & (g2776)) + ((g2754) & (g2755) & (g2756) & (!g2757) & (!g2775) & (!g2776)) + ((g2754) & (g2755) & (g2756) & (!g2757) & (g2775) & (g2776)) + ((g2754) & (g2755) & (g2756) & (g2757) & (!g2775) & (!g2776)) + ((g2754) & (g2755) & (g2756) & (g2757) & (g2775) & (g2776)));
	assign g2778 = (((!g2706) & (!g2091) & (!g2090) & (g2089) & (g2196) & (g2197)) + ((!g2706) & (!g2091) & (g2090) & (!g2089) & (!g2196) & (g2197)) + ((!g2706) & (!g2091) & (g2090) & (g2089) & (!g2196) & (g2197)) + ((!g2706) & (!g2091) & (g2090) & (g2089) & (g2196) & (g2197)) + ((!g2706) & (g2091) & (!g2090) & (!g2089) & (g2196) & (!g2197)) + ((!g2706) & (g2091) & (!g2090) & (g2089) & (g2196) & (!g2197)) + ((!g2706) & (g2091) & (!g2090) & (g2089) & (g2196) & (g2197)) + ((!g2706) & (g2091) & (g2090) & (!g2089) & (!g2196) & (g2197)) + ((!g2706) & (g2091) & (g2090) & (!g2089) & (g2196) & (!g2197)) + ((!g2706) & (g2091) & (g2090) & (g2089) & (!g2196) & (g2197)) + ((!g2706) & (g2091) & (g2090) & (g2089) & (g2196) & (!g2197)) + ((!g2706) & (g2091) & (g2090) & (g2089) & (g2196) & (g2197)) + ((g2706) & (!g2091) & (!g2090) & (!g2089) & (!g2196) & (!g2197)) + ((g2706) & (!g2091) & (!g2090) & (g2089) & (!g2196) & (!g2197)) + ((g2706) & (!g2091) & (!g2090) & (g2089) & (g2196) & (g2197)) + ((g2706) & (!g2091) & (g2090) & (!g2089) & (!g2196) & (!g2197)) + ((g2706) & (!g2091) & (g2090) & (!g2089) & (!g2196) & (g2197)) + ((g2706) & (!g2091) & (g2090) & (g2089) & (!g2196) & (!g2197)) + ((g2706) & (!g2091) & (g2090) & (g2089) & (!g2196) & (g2197)) + ((g2706) & (!g2091) & (g2090) & (g2089) & (g2196) & (g2197)) + ((g2706) & (g2091) & (!g2090) & (!g2089) & (!g2196) & (!g2197)) + ((g2706) & (g2091) & (!g2090) & (!g2089) & (g2196) & (!g2197)) + ((g2706) & (g2091) & (!g2090) & (g2089) & (!g2196) & (!g2197)) + ((g2706) & (g2091) & (!g2090) & (g2089) & (g2196) & (!g2197)) + ((g2706) & (g2091) & (!g2090) & (g2089) & (g2196) & (g2197)) + ((g2706) & (g2091) & (g2090) & (!g2089) & (!g2196) & (!g2197)) + ((g2706) & (g2091) & (g2090) & (!g2089) & (!g2196) & (g2197)) + ((g2706) & (g2091) & (g2090) & (!g2089) & (g2196) & (!g2197)) + ((g2706) & (g2091) & (g2090) & (g2089) & (!g2196) & (!g2197)) + ((g2706) & (g2091) & (g2090) & (g2089) & (!g2196) & (g2197)) + ((g2706) & (g2091) & (g2090) & (g2089) & (g2196) & (!g2197)) + ((g2706) & (g2091) & (g2090) & (g2089) & (g2196) & (g2197)));
	assign g2779 = (((!g2468) & (!g2778) & (!g2632) & (g2559) & (g2201) & (g2202)) + ((!g2468) & (!g2778) & (g2632) & (!g2559) & (!g2201) & (g2202)) + ((!g2468) & (!g2778) & (g2632) & (g2559) & (!g2201) & (g2202)) + ((!g2468) & (!g2778) & (g2632) & (g2559) & (g2201) & (g2202)) + ((!g2468) & (g2778) & (!g2632) & (!g2559) & (g2201) & (!g2202)) + ((!g2468) & (g2778) & (!g2632) & (g2559) & (g2201) & (!g2202)) + ((!g2468) & (g2778) & (!g2632) & (g2559) & (g2201) & (g2202)) + ((!g2468) & (g2778) & (g2632) & (!g2559) & (!g2201) & (g2202)) + ((!g2468) & (g2778) & (g2632) & (!g2559) & (g2201) & (!g2202)) + ((!g2468) & (g2778) & (g2632) & (g2559) & (!g2201) & (g2202)) + ((!g2468) & (g2778) & (g2632) & (g2559) & (g2201) & (!g2202)) + ((!g2468) & (g2778) & (g2632) & (g2559) & (g2201) & (g2202)) + ((g2468) & (!g2778) & (!g2632) & (!g2559) & (!g2201) & (!g2202)) + ((g2468) & (!g2778) & (!g2632) & (g2559) & (!g2201) & (!g2202)) + ((g2468) & (!g2778) & (!g2632) & (g2559) & (g2201) & (g2202)) + ((g2468) & (!g2778) & (g2632) & (!g2559) & (!g2201) & (!g2202)) + ((g2468) & (!g2778) & (g2632) & (!g2559) & (!g2201) & (g2202)) + ((g2468) & (!g2778) & (g2632) & (g2559) & (!g2201) & (!g2202)) + ((g2468) & (!g2778) & (g2632) & (g2559) & (!g2201) & (g2202)) + ((g2468) & (!g2778) & (g2632) & (g2559) & (g2201) & (g2202)) + ((g2468) & (g2778) & (!g2632) & (!g2559) & (!g2201) & (!g2202)) + ((g2468) & (g2778) & (!g2632) & (!g2559) & (g2201) & (!g2202)) + ((g2468) & (g2778) & (!g2632) & (g2559) & (!g2201) & (!g2202)) + ((g2468) & (g2778) & (!g2632) & (g2559) & (g2201) & (!g2202)) + ((g2468) & (g2778) & (!g2632) & (g2559) & (g2201) & (g2202)) + ((g2468) & (g2778) & (g2632) & (!g2559) & (!g2201) & (!g2202)) + ((g2468) & (g2778) & (g2632) & (!g2559) & (!g2201) & (g2202)) + ((g2468) & (g2778) & (g2632) & (!g2559) & (g2201) & (!g2202)) + ((g2468) & (g2778) & (g2632) & (g2559) & (!g2201) & (!g2202)) + ((g2468) & (g2778) & (g2632) & (g2559) & (!g2201) & (g2202)) + ((g2468) & (g2778) & (g2632) & (g2559) & (g2201) & (!g2202)) + ((g2468) & (g2778) & (g2632) & (g2559) & (g2201) & (g2202)));
	assign g2780 = (((!g2073) & (!sk[86]) & (g2080) & (!g2125)) + ((!g2073) & (!sk[86]) & (g2080) & (g2125)) + ((!g2073) & (sk[86]) & (!g2080) & (!g2125)) + ((g2073) & (!sk[86]) & (!g2080) & (!g2125)) + ((g2073) & (!sk[86]) & (!g2080) & (g2125)) + ((g2073) & (!sk[86]) & (g2080) & (!g2125)) + ((g2073) & (!sk[86]) & (g2080) & (g2125)) + ((g2073) & (sk[86]) & (!g2080) & (!g2125)) + ((g2073) & (sk[86]) & (!g2080) & (g2125)));
	assign g2781 = (((!g3265) & (!g2779) & (!g2469) & (g2192) & (g2780) & (g2190)) + ((!g3265) & (!g2779) & (g2469) & (!g2192) & (!g2780) & (g2190)) + ((!g3265) & (!g2779) & (g2469) & (g2192) & (!g2780) & (g2190)) + ((!g3265) & (!g2779) & (g2469) & (g2192) & (g2780) & (g2190)) + ((!g3265) & (g2779) & (!g2469) & (!g2192) & (g2780) & (!g2190)) + ((!g3265) & (g2779) & (!g2469) & (g2192) & (g2780) & (!g2190)) + ((!g3265) & (g2779) & (!g2469) & (g2192) & (g2780) & (g2190)) + ((!g3265) & (g2779) & (g2469) & (!g2192) & (!g2780) & (g2190)) + ((!g3265) & (g2779) & (g2469) & (!g2192) & (g2780) & (!g2190)) + ((!g3265) & (g2779) & (g2469) & (g2192) & (!g2780) & (g2190)) + ((!g3265) & (g2779) & (g2469) & (g2192) & (g2780) & (!g2190)) + ((!g3265) & (g2779) & (g2469) & (g2192) & (g2780) & (g2190)) + ((g3265) & (!g2779) & (!g2469) & (!g2192) & (!g2780) & (!g2190)) + ((g3265) & (!g2779) & (!g2469) & (g2192) & (!g2780) & (!g2190)) + ((g3265) & (!g2779) & (!g2469) & (g2192) & (g2780) & (g2190)) + ((g3265) & (!g2779) & (g2469) & (!g2192) & (!g2780) & (!g2190)) + ((g3265) & (!g2779) & (g2469) & (!g2192) & (!g2780) & (g2190)) + ((g3265) & (!g2779) & (g2469) & (g2192) & (!g2780) & (!g2190)) + ((g3265) & (!g2779) & (g2469) & (g2192) & (!g2780) & (g2190)) + ((g3265) & (!g2779) & (g2469) & (g2192) & (g2780) & (g2190)) + ((g3265) & (g2779) & (!g2469) & (!g2192) & (!g2780) & (!g2190)) + ((g3265) & (g2779) & (!g2469) & (!g2192) & (g2780) & (!g2190)) + ((g3265) & (g2779) & (!g2469) & (g2192) & (!g2780) & (!g2190)) + ((g3265) & (g2779) & (!g2469) & (g2192) & (g2780) & (!g2190)) + ((g3265) & (g2779) & (!g2469) & (g2192) & (g2780) & (g2190)) + ((g3265) & (g2779) & (g2469) & (!g2192) & (!g2780) & (!g2190)) + ((g3265) & (g2779) & (g2469) & (!g2192) & (!g2780) & (g2190)) + ((g3265) & (g2779) & (g2469) & (!g2192) & (g2780) & (!g2190)) + ((g3265) & (g2779) & (g2469) & (g2192) & (!g2780) & (!g2190)) + ((g3265) & (g2779) & (g2469) & (g2192) & (!g2780) & (g2190)) + ((g3265) & (g2779) & (g2469) & (g2192) & (g2780) & (!g2190)) + ((g3265) & (g2779) & (g2469) & (g2192) & (g2780) & (g2190)));
	assign g2782 = (((!g2081) & (!g2124) & (!g2770) & (!g2771) & (!g2781) & (!g2098)) + ((!g2081) & (!g2124) & (!g2770) & (!g2771) & (!g2781) & (g2098)) + ((!g2081) & (!g2124) & (!g2770) & (g2771) & (!g2781) & (!g2098)) + ((!g2081) & (!g2124) & (!g2770) & (g2771) & (!g2781) & (g2098)) + ((!g2081) & (!g2124) & (g2770) & (!g2771) & (!g2781) & (!g2098)) + ((!g2081) & (!g2124) & (g2770) & (!g2771) & (g2781) & (!g2098)) + ((!g2081) & (!g2124) & (g2770) & (g2771) & (!g2781) & (!g2098)) + ((!g2081) & (!g2124) & (g2770) & (g2771) & (g2781) & (!g2098)) + ((!g2081) & (g2124) & (!g2770) & (!g2771) & (!g2781) & (!g2098)) + ((!g2081) & (g2124) & (!g2770) & (!g2771) & (g2781) & (!g2098)) + ((!g2081) & (g2124) & (g2770) & (!g2771) & (!g2781) & (!g2098)) + ((!g2081) & (g2124) & (g2770) & (!g2771) & (g2781) & (!g2098)) + ((!g2081) & (g2124) & (g2770) & (g2771) & (!g2781) & (!g2098)) + ((!g2081) & (g2124) & (g2770) & (g2771) & (g2781) & (!g2098)) + ((g2081) & (!g2124) & (!g2770) & (!g2771) & (!g2781) & (!g2098)) + ((g2081) & (!g2124) & (!g2770) & (!g2771) & (!g2781) & (g2098)) + ((g2081) & (!g2124) & (!g2770) & (g2771) & (!g2781) & (!g2098)) + ((g2081) & (!g2124) & (!g2770) & (g2771) & (!g2781) & (g2098)) + ((g2081) & (!g2124) & (g2770) & (!g2771) & (!g2781) & (!g2098)) + ((g2081) & (!g2124) & (g2770) & (!g2771) & (g2781) & (!g2098)) + ((g2081) & (!g2124) & (g2770) & (g2771) & (!g2781) & (!g2098)) + ((g2081) & (!g2124) & (g2770) & (g2771) & (g2781) & (!g2098)) + ((g2081) & (g2124) & (!g2770) & (!g2771) & (!g2781) & (!g2098)) + ((g2081) & (g2124) & (!g2770) & (!g2771) & (g2781) & (!g2098)) + ((g2081) & (g2124) & (!g2770) & (g2771) & (!g2781) & (g2098)) + ((g2081) & (g2124) & (!g2770) & (g2771) & (g2781) & (g2098)) + ((g2081) & (g2124) & (g2770) & (!g2771) & (!g2781) & (!g2098)) + ((g2081) & (g2124) & (g2770) & (!g2771) & (g2781) & (!g2098)) + ((g2081) & (g2124) & (g2770) & (g2771) & (!g2781) & (!g2098)) + ((g2081) & (g2124) & (g2770) & (g2771) & (g2781) & (!g2098)));
	assign g2783 = (((!g2363) & (!sk[89]) & (g2338)) + ((g2363) & (!sk[89]) & (g2338)) + ((g2363) & (sk[89]) & (g2338)));
	assign g2784 = (((!g2549) & (!dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[90]) & (g2128) & (!g2129)) + ((!g2549) & (!dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[90]) & (g2128) & (g2129)) + ((!g2549) & (!dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (!g2128) & (!g2129)) + ((!g2549) & (!dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (!g2128) & (g2129)) + ((!g2549) & (!dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (g2128) & (!g2129)) + ((!g2549) & (!dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (g2128) & (g2129)) + ((!g2549) & (dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[90]) & (g2128) & (!g2129)) + ((!g2549) & (dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[90]) & (g2128) & (g2129)) + ((!g2549) & (dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (!g2128) & (!g2129)) + ((!g2549) & (dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (!g2128) & (g2129)) + ((!g2549) & (dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (g2128) & (!g2129)) + ((!g2549) & (dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (g2128) & (g2129)) + ((g2549) & (!dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[90]) & (!g2128) & (!g2129)) + ((g2549) & (!dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[90]) & (!g2128) & (g2129)) + ((g2549) & (!dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[90]) & (g2128) & (!g2129)) + ((g2549) & (!dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[90]) & (g2128) & (g2129)) + ((g2549) & (!dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (!g2128) & (!g2129)) + ((g2549) & (!dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (!g2128) & (g2129)) + ((g2549) & (!dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (g2128) & (!g2129)) + ((g2549) & (!dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (g2128) & (g2129)) + ((g2549) & (!dmem_dat_ix31x) & (dmem_dat_ix15x) & (sk[90]) & (!g2128) & (g2129)) + ((g2549) & (dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[90]) & (!g2128) & (!g2129)) + ((g2549) & (dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[90]) & (!g2128) & (g2129)) + ((g2549) & (dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[90]) & (g2128) & (!g2129)) + ((g2549) & (dmem_dat_ix31x) & (!dmem_dat_ix15x) & (!sk[90]) & (g2128) & (g2129)) + ((g2549) & (dmem_dat_ix31x) & (!dmem_dat_ix15x) & (sk[90]) & (!g2128) & (!g2129)) + ((g2549) & (dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (!g2128) & (!g2129)) + ((g2549) & (dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (!g2128) & (g2129)) + ((g2549) & (dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (g2128) & (!g2129)) + ((g2549) & (dmem_dat_ix31x) & (dmem_dat_ix15x) & (!sk[90]) & (g2128) & (g2129)) + ((g2549) & (dmem_dat_ix31x) & (dmem_dat_ix15x) & (sk[90]) & (!g2128) & (!g2129)) + ((g2549) & (dmem_dat_ix31x) & (dmem_dat_ix15x) & (sk[90]) & (!g2128) & (g2129)));
	assign g2785 = (((!sk[91]) & (!g75) & (g2131)) + ((!sk[91]) & (g75) & (g2131)) + ((sk[91]) & (g75) & (g2131)));
	assign g2786 = (((!g75) & (!sk[92]) & (g2127)) + ((g75) & (!sk[92]) & (g2127)) + ((g75) & (sk[92]) & (!g2127)));
	assign g2787 = (((!g2782) & (!dmem_dat_ix28x) & (!g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2782) & (!dmem_dat_ix28x) & (!g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2782) & (!dmem_dat_ix28x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((!g2782) & (!dmem_dat_ix28x) & (g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2782) & (!dmem_dat_ix28x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((!g2782) & (!dmem_dat_ix28x) & (g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2782) & (!dmem_dat_ix28x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((!g2782) & (!dmem_dat_ix28x) & (g2783) & (g2784) & (g2785) & (g2786)) + ((!g2782) & (dmem_dat_ix28x) & (!g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2782) & (dmem_dat_ix28x) & (!g2783) & (!g2784) & (g2785) & (!g2786)) + ((!g2782) & (dmem_dat_ix28x) & (!g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2782) & (dmem_dat_ix28x) & (!g2783) & (g2784) & (g2785) & (!g2786)) + ((!g2782) & (dmem_dat_ix28x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((!g2782) & (dmem_dat_ix28x) & (g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2782) & (dmem_dat_ix28x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((!g2782) & (dmem_dat_ix28x) & (g2783) & (!g2784) & (g2785) & (!g2786)) + ((!g2782) & (dmem_dat_ix28x) & (g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2782) & (dmem_dat_ix28x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((!g2782) & (dmem_dat_ix28x) & (g2783) & (g2784) & (g2785) & (!g2786)) + ((!g2782) & (dmem_dat_ix28x) & (g2783) & (g2784) & (g2785) & (g2786)) + ((g2782) & (!dmem_dat_ix28x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((g2782) & (!dmem_dat_ix28x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((g2782) & (!dmem_dat_ix28x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((g2782) & (!dmem_dat_ix28x) & (g2783) & (g2784) & (g2785) & (g2786)) + ((g2782) & (dmem_dat_ix28x) & (!g2783) & (!g2784) & (g2785) & (!g2786)) + ((g2782) & (dmem_dat_ix28x) & (!g2783) & (g2784) & (g2785) & (!g2786)) + ((g2782) & (dmem_dat_ix28x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((g2782) & (dmem_dat_ix28x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((g2782) & (dmem_dat_ix28x) & (g2783) & (!g2784) & (g2785) & (!g2786)) + ((g2782) & (dmem_dat_ix28x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((g2782) & (dmem_dat_ix28x) & (g2783) & (g2784) & (g2785) & (!g2786)) + ((g2782) & (dmem_dat_ix28x) & (g2783) & (g2784) & (g2785) & (g2786)));
	assign g2788 = (((!g1320) & (!g2727) & (!sk[94]) & (!g1365) & (g1410)) + ((!g1320) & (!g2727) & (!sk[94]) & (g1365) & (g1410)) + ((!g1320) & (g2727) & (!sk[94]) & (!g1365) & (!g1410)) + ((!g1320) & (g2727) & (!sk[94]) & (!g1365) & (g1410)) + ((!g1320) & (g2727) & (!sk[94]) & (g1365) & (!g1410)) + ((!g1320) & (g2727) & (!sk[94]) & (g1365) & (g1410)) + ((g1320) & (!g2727) & (!sk[94]) & (!g1365) & (!g1410)) + ((g1320) & (!g2727) & (!sk[94]) & (!g1365) & (g1410)) + ((g1320) & (!g2727) & (!sk[94]) & (g1365) & (!g1410)) + ((g1320) & (!g2727) & (!sk[94]) & (g1365) & (g1410)) + ((g1320) & (g2727) & (!sk[94]) & (!g1365) & (!g1410)) + ((g1320) & (g2727) & (!sk[94]) & (!g1365) & (g1410)) + ((g1320) & (g2727) & (!sk[94]) & (g1365) & (!g1410)) + ((g1320) & (g2727) & (!sk[94]) & (g1365) & (g1410)) + ((g1320) & (g2727) & (sk[94]) & (g1365) & (g1410)));
	assign g2789 = (((!g1455) & (!sk[95]) & (g2788)) + ((!g1455) & (sk[95]) & (g2788)) + ((g1455) & (!sk[95]) & (g2788)) + ((g1455) & (sk[95]) & (!g2788)));
	assign g2790 = (((!sk[96]) & (!g107) & (!g1410) & (!g2765) & (g1455)) + ((!sk[96]) & (!g107) & (!g1410) & (g2765) & (g1455)) + ((!sk[96]) & (!g107) & (g1410) & (!g2765) & (!g1455)) + ((!sk[96]) & (!g107) & (g1410) & (!g2765) & (g1455)) + ((!sk[96]) & (!g107) & (g1410) & (g2765) & (!g1455)) + ((!sk[96]) & (!g107) & (g1410) & (g2765) & (g1455)) + ((!sk[96]) & (g107) & (!g1410) & (!g2765) & (!g1455)) + ((!sk[96]) & (g107) & (!g1410) & (!g2765) & (g1455)) + ((!sk[96]) & (g107) & (!g1410) & (g2765) & (!g1455)) + ((!sk[96]) & (g107) & (!g1410) & (g2765) & (g1455)) + ((!sk[96]) & (g107) & (g1410) & (!g2765) & (!g1455)) + ((!sk[96]) & (g107) & (g1410) & (!g2765) & (g1455)) + ((!sk[96]) & (g107) & (g1410) & (g2765) & (!g1455)) + ((!sk[96]) & (g107) & (g1410) & (g2765) & (g1455)) + ((sk[96]) & (!g107) & (!g1410) & (!g2765) & (g1455)) + ((sk[96]) & (!g107) & (!g1410) & (g2765) & (g1455)) + ((sk[96]) & (!g107) & (g1410) & (!g2765) & (g1455)) + ((sk[96]) & (!g107) & (g1410) & (g2765) & (!g1455)) + ((sk[96]) & (g107) & (!g1410) & (!g2765) & (!g1455)) + ((sk[96]) & (g107) & (!g1410) & (g2765) & (g1455)) + ((sk[96]) & (g107) & (g1410) & (!g2765) & (g1455)) + ((sk[96]) & (g107) & (g1410) & (g2765) & (g1455)));
	assign g5052 = (((!g2921) & (!g3107) & (sk[97]) & (g2791)) + ((!g2921) & (g3107) & (!sk[97]) & (!g2791)) + ((!g2921) & (g3107) & (!sk[97]) & (g2791)) + ((!g2921) & (g3107) & (sk[97]) & (g2791)) + ((g2921) & (!g3107) & (!sk[97]) & (!g2791)) + ((g2921) & (!g3107) & (!sk[97]) & (g2791)) + ((g2921) & (g3107) & (!sk[97]) & (!g2791)) + ((g2921) & (g3107) & (!sk[97]) & (g2791)) + ((g2921) & (g3107) & (sk[97]) & (!g2791)) + ((g2921) & (g3107) & (sk[97]) & (g2791)));
	assign g2792 = (((!sk[98]) & (!g1968) & (!g2033) & (!g2034) & (g2790) & (!g2791)) + ((!sk[98]) & (!g1968) & (!g2033) & (!g2034) & (g2790) & (g2791)) + ((!sk[98]) & (!g1968) & (!g2033) & (g2034) & (!g2790) & (!g2791)) + ((!sk[98]) & (!g1968) & (!g2033) & (g2034) & (!g2790) & (g2791)) + ((!sk[98]) & (!g1968) & (!g2033) & (g2034) & (g2790) & (!g2791)) + ((!sk[98]) & (!g1968) & (!g2033) & (g2034) & (g2790) & (g2791)) + ((!sk[98]) & (!g1968) & (g2033) & (!g2034) & (g2790) & (!g2791)) + ((!sk[98]) & (!g1968) & (g2033) & (!g2034) & (g2790) & (g2791)) + ((!sk[98]) & (!g1968) & (g2033) & (g2034) & (!g2790) & (!g2791)) + ((!sk[98]) & (!g1968) & (g2033) & (g2034) & (!g2790) & (g2791)) + ((!sk[98]) & (!g1968) & (g2033) & (g2034) & (g2790) & (!g2791)) + ((!sk[98]) & (!g1968) & (g2033) & (g2034) & (g2790) & (g2791)) + ((!sk[98]) & (g1968) & (!g2033) & (!g2034) & (!g2790) & (!g2791)) + ((!sk[98]) & (g1968) & (!g2033) & (!g2034) & (!g2790) & (g2791)) + ((!sk[98]) & (g1968) & (!g2033) & (!g2034) & (g2790) & (!g2791)) + ((!sk[98]) & (g1968) & (!g2033) & (!g2034) & (g2790) & (g2791)) + ((!sk[98]) & (g1968) & (!g2033) & (g2034) & (!g2790) & (!g2791)) + ((!sk[98]) & (g1968) & (!g2033) & (g2034) & (!g2790) & (g2791)) + ((!sk[98]) & (g1968) & (!g2033) & (g2034) & (g2790) & (!g2791)) + ((!sk[98]) & (g1968) & (!g2033) & (g2034) & (g2790) & (g2791)) + ((!sk[98]) & (g1968) & (g2033) & (!g2034) & (!g2790) & (!g2791)) + ((!sk[98]) & (g1968) & (g2033) & (!g2034) & (!g2790) & (g2791)) + ((!sk[98]) & (g1968) & (g2033) & (!g2034) & (g2790) & (!g2791)) + ((!sk[98]) & (g1968) & (g2033) & (!g2034) & (g2790) & (g2791)) + ((!sk[98]) & (g1968) & (g2033) & (g2034) & (!g2790) & (!g2791)) + ((!sk[98]) & (g1968) & (g2033) & (g2034) & (!g2790) & (g2791)) + ((!sk[98]) & (g1968) & (g2033) & (g2034) & (g2790) & (!g2791)) + ((!sk[98]) & (g1968) & (g2033) & (g2034) & (g2790) & (g2791)) + ((sk[98]) & (!g1968) & (!g2033) & (!g2034) & (!g2790) & (g2791)) + ((sk[98]) & (!g1968) & (!g2033) & (!g2034) & (g2790) & (g2791)) + ((sk[98]) & (!g1968) & (g2033) & (!g2034) & (g2790) & (!g2791)) + ((sk[98]) & (!g1968) & (g2033) & (!g2034) & (g2790) & (g2791)) + ((sk[98]) & (g1968) & (!g2033) & (!g2034) & (!g2790) & (g2791)) + ((sk[98]) & (g1968) & (!g2033) & (!g2034) & (g2790) & (g2791)) + ((sk[98]) & (g1968) & (!g2033) & (g2034) & (!g2790) & (!g2791)) + ((sk[98]) & (g1968) & (!g2033) & (g2034) & (!g2790) & (g2791)) + ((sk[98]) & (g1968) & (!g2033) & (g2034) & (g2790) & (!g2791)) + ((sk[98]) & (g1968) & (!g2033) & (g2034) & (g2790) & (g2791)) + ((sk[98]) & (g1968) & (g2033) & (!g2034) & (g2790) & (!g2791)) + ((sk[98]) & (g1968) & (g2033) & (!g2034) & (g2790) & (g2791)));
	assign g2793 = (((!g2329) & (!g2029) & (!g2408) & (g2789) & (!sk[99]) & (!g2792)) + ((!g2329) & (!g2029) & (!g2408) & (g2789) & (!sk[99]) & (g2792)) + ((!g2329) & (!g2029) & (g2408) & (!g2789) & (!sk[99]) & (!g2792)) + ((!g2329) & (!g2029) & (g2408) & (!g2789) & (!sk[99]) & (g2792)) + ((!g2329) & (!g2029) & (g2408) & (g2789) & (!sk[99]) & (!g2792)) + ((!g2329) & (!g2029) & (g2408) & (g2789) & (!sk[99]) & (g2792)) + ((!g2329) & (g2029) & (!g2408) & (g2789) & (!sk[99]) & (!g2792)) + ((!g2329) & (g2029) & (!g2408) & (g2789) & (!sk[99]) & (g2792)) + ((!g2329) & (g2029) & (g2408) & (!g2789) & (!sk[99]) & (!g2792)) + ((!g2329) & (g2029) & (g2408) & (!g2789) & (!sk[99]) & (g2792)) + ((!g2329) & (g2029) & (g2408) & (g2789) & (!sk[99]) & (!g2792)) + ((!g2329) & (g2029) & (g2408) & (g2789) & (!sk[99]) & (g2792)) + ((g2329) & (!g2029) & (!g2408) & (!g2789) & (!sk[99]) & (!g2792)) + ((g2329) & (!g2029) & (!g2408) & (!g2789) & (!sk[99]) & (g2792)) + ((g2329) & (!g2029) & (!g2408) & (g2789) & (!sk[99]) & (!g2792)) + ((g2329) & (!g2029) & (!g2408) & (g2789) & (!sk[99]) & (g2792)) + ((g2329) & (!g2029) & (g2408) & (!g2789) & (!sk[99]) & (!g2792)) + ((g2329) & (!g2029) & (g2408) & (!g2789) & (!sk[99]) & (g2792)) + ((g2329) & (!g2029) & (g2408) & (!g2789) & (sk[99]) & (g2792)) + ((g2329) & (!g2029) & (g2408) & (g2789) & (!sk[99]) & (!g2792)) + ((g2329) & (!g2029) & (g2408) & (g2789) & (!sk[99]) & (g2792)) + ((g2329) & (!g2029) & (g2408) & (g2789) & (sk[99]) & (g2792)) + ((g2329) & (g2029) & (!g2408) & (!g2789) & (!sk[99]) & (!g2792)) + ((g2329) & (g2029) & (!g2408) & (!g2789) & (!sk[99]) & (g2792)) + ((g2329) & (g2029) & (!g2408) & (g2789) & (!sk[99]) & (!g2792)) + ((g2329) & (g2029) & (!g2408) & (g2789) & (!sk[99]) & (g2792)) + ((g2329) & (g2029) & (g2408) & (!g2789) & (!sk[99]) & (!g2792)) + ((g2329) & (g2029) & (g2408) & (!g2789) & (!sk[99]) & (g2792)) + ((g2329) & (g2029) & (g2408) & (g2789) & (!sk[99]) & (!g2792)) + ((g2329) & (g2029) & (g2408) & (g2789) & (!sk[99]) & (g2792)) + ((g2329) & (g2029) & (g2408) & (g2789) & (sk[99]) & (!g2792)) + ((g2329) & (g2029) & (g2408) & (g2789) & (sk[99]) & (g2792)));
	assign g2795 = (((!sk[100]) & (!g2098) & (!g2099) & (!g2771) & (g2772) & (!g2794)) + ((!sk[100]) & (!g2098) & (!g2099) & (!g2771) & (g2772) & (g2794)) + ((!sk[100]) & (!g2098) & (!g2099) & (g2771) & (!g2772) & (!g2794)) + ((!sk[100]) & (!g2098) & (!g2099) & (g2771) & (!g2772) & (g2794)) + ((!sk[100]) & (!g2098) & (!g2099) & (g2771) & (g2772) & (!g2794)) + ((!sk[100]) & (!g2098) & (!g2099) & (g2771) & (g2772) & (g2794)) + ((!sk[100]) & (!g2098) & (g2099) & (!g2771) & (g2772) & (!g2794)) + ((!sk[100]) & (!g2098) & (g2099) & (!g2771) & (g2772) & (g2794)) + ((!sk[100]) & (!g2098) & (g2099) & (g2771) & (!g2772) & (!g2794)) + ((!sk[100]) & (!g2098) & (g2099) & (g2771) & (!g2772) & (g2794)) + ((!sk[100]) & (!g2098) & (g2099) & (g2771) & (g2772) & (!g2794)) + ((!sk[100]) & (!g2098) & (g2099) & (g2771) & (g2772) & (g2794)) + ((!sk[100]) & (g2098) & (!g2099) & (!g2771) & (!g2772) & (!g2794)) + ((!sk[100]) & (g2098) & (!g2099) & (!g2771) & (!g2772) & (g2794)) + ((!sk[100]) & (g2098) & (!g2099) & (!g2771) & (g2772) & (!g2794)) + ((!sk[100]) & (g2098) & (!g2099) & (!g2771) & (g2772) & (g2794)) + ((!sk[100]) & (g2098) & (!g2099) & (g2771) & (!g2772) & (!g2794)) + ((!sk[100]) & (g2098) & (!g2099) & (g2771) & (!g2772) & (g2794)) + ((!sk[100]) & (g2098) & (!g2099) & (g2771) & (g2772) & (!g2794)) + ((!sk[100]) & (g2098) & (!g2099) & (g2771) & (g2772) & (g2794)) + ((!sk[100]) & (g2098) & (g2099) & (!g2771) & (!g2772) & (!g2794)) + ((!sk[100]) & (g2098) & (g2099) & (!g2771) & (!g2772) & (g2794)) + ((!sk[100]) & (g2098) & (g2099) & (!g2771) & (g2772) & (!g2794)) + ((!sk[100]) & (g2098) & (g2099) & (!g2771) & (g2772) & (g2794)) + ((!sk[100]) & (g2098) & (g2099) & (g2771) & (!g2772) & (!g2794)) + ((!sk[100]) & (g2098) & (g2099) & (g2771) & (!g2772) & (g2794)) + ((!sk[100]) & (g2098) & (g2099) & (g2771) & (g2772) & (!g2794)) + ((!sk[100]) & (g2098) & (g2099) & (g2771) & (g2772) & (g2794)) + ((sk[100]) & (!g2098) & (!g2099) & (!g2771) & (!g2772) & (g2794)) + ((sk[100]) & (!g2098) & (!g2099) & (!g2771) & (g2772) & (g2794)) + ((sk[100]) & (!g2098) & (!g2099) & (g2771) & (!g2772) & (g2794)) + ((sk[100]) & (!g2098) & (!g2099) & (g2771) & (g2772) & (!g2794)) + ((sk[100]) & (!g2098) & (g2099) & (!g2771) & (!g2772) & (!g2794)) + ((sk[100]) & (!g2098) & (g2099) & (!g2771) & (g2772) & (!g2794)) + ((sk[100]) & (!g2098) & (g2099) & (g2771) & (!g2772) & (!g2794)) + ((sk[100]) & (!g2098) & (g2099) & (g2771) & (g2772) & (g2794)) + ((sk[100]) & (g2098) & (!g2099) & (!g2771) & (!g2772) & (g2794)) + ((sk[100]) & (g2098) & (!g2099) & (!g2771) & (g2772) & (!g2794)) + ((sk[100]) & (g2098) & (!g2099) & (g2771) & (!g2772) & (!g2794)) + ((sk[100]) & (g2098) & (!g2099) & (g2771) & (g2772) & (!g2794)) + ((sk[100]) & (g2098) & (g2099) & (!g2771) & (!g2772) & (!g2794)) + ((sk[100]) & (g2098) & (g2099) & (!g2771) & (g2772) & (g2794)) + ((sk[100]) & (g2098) & (g2099) & (g2771) & (!g2772) & (g2794)) + ((sk[100]) & (g2098) & (g2099) & (g2771) & (g2772) & (g2794)));
	assign g2796 = (((!g2737) & (!sk[101]) & (!g2738) & (!g2752) & (g2772) & (!g2773)) + ((!g2737) & (!sk[101]) & (!g2738) & (!g2752) & (g2772) & (g2773)) + ((!g2737) & (!sk[101]) & (!g2738) & (g2752) & (!g2772) & (!g2773)) + ((!g2737) & (!sk[101]) & (!g2738) & (g2752) & (!g2772) & (g2773)) + ((!g2737) & (!sk[101]) & (!g2738) & (g2752) & (g2772) & (!g2773)) + ((!g2737) & (!sk[101]) & (!g2738) & (g2752) & (g2772) & (g2773)) + ((!g2737) & (!sk[101]) & (g2738) & (!g2752) & (g2772) & (!g2773)) + ((!g2737) & (!sk[101]) & (g2738) & (!g2752) & (g2772) & (g2773)) + ((!g2737) & (!sk[101]) & (g2738) & (g2752) & (!g2772) & (!g2773)) + ((!g2737) & (!sk[101]) & (g2738) & (g2752) & (!g2772) & (g2773)) + ((!g2737) & (!sk[101]) & (g2738) & (g2752) & (g2772) & (!g2773)) + ((!g2737) & (!sk[101]) & (g2738) & (g2752) & (g2772) & (g2773)) + ((g2737) & (!sk[101]) & (!g2738) & (!g2752) & (!g2772) & (!g2773)) + ((g2737) & (!sk[101]) & (!g2738) & (!g2752) & (!g2772) & (g2773)) + ((g2737) & (!sk[101]) & (!g2738) & (!g2752) & (g2772) & (!g2773)) + ((g2737) & (!sk[101]) & (!g2738) & (!g2752) & (g2772) & (g2773)) + ((g2737) & (!sk[101]) & (!g2738) & (g2752) & (!g2772) & (!g2773)) + ((g2737) & (!sk[101]) & (!g2738) & (g2752) & (!g2772) & (g2773)) + ((g2737) & (!sk[101]) & (!g2738) & (g2752) & (g2772) & (!g2773)) + ((g2737) & (!sk[101]) & (!g2738) & (g2752) & (g2772) & (g2773)) + ((g2737) & (!sk[101]) & (g2738) & (!g2752) & (!g2772) & (!g2773)) + ((g2737) & (!sk[101]) & (g2738) & (!g2752) & (!g2772) & (g2773)) + ((g2737) & (!sk[101]) & (g2738) & (!g2752) & (g2772) & (!g2773)) + ((g2737) & (!sk[101]) & (g2738) & (!g2752) & (g2772) & (g2773)) + ((g2737) & (!sk[101]) & (g2738) & (g2752) & (!g2772) & (!g2773)) + ((g2737) & (!sk[101]) & (g2738) & (g2752) & (!g2772) & (g2773)) + ((g2737) & (!sk[101]) & (g2738) & (g2752) & (g2772) & (!g2773)) + ((g2737) & (!sk[101]) & (g2738) & (g2752) & (g2772) & (g2773)) + ((g2737) & (sk[101]) & (g2738) & (g2752) & (!g2772) & (g2773)) + ((g2737) & (sk[101]) & (g2738) & (g2752) & (g2772) & (!g2773)));
	assign g2797 = (((!g2754) & (!g2755) & (!g2756) & (!g2757) & (!g2775) & (!g2776)) + ((!g2754) & (!g2755) & (!g2756) & (!g2757) & (!g2775) & (g2776)) + ((!g2754) & (!g2755) & (!g2756) & (!g2757) & (g2775) & (!g2776)) + ((!g2754) & (!g2755) & (!g2756) & (g2757) & (!g2775) & (!g2776)) + ((!g2754) & (!g2755) & (!g2756) & (g2757) & (!g2775) & (g2776)) + ((!g2754) & (!g2755) & (!g2756) & (g2757) & (g2775) & (!g2776)) + ((!g2754) & (!g2755) & (g2756) & (!g2757) & (!g2775) & (!g2776)) + ((!g2754) & (!g2755) & (g2756) & (!g2757) & (!g2775) & (g2776)) + ((!g2754) & (!g2755) & (g2756) & (!g2757) & (g2775) & (!g2776)) + ((!g2754) & (!g2755) & (g2756) & (g2757) & (!g2775) & (!g2776)) + ((!g2754) & (g2755) & (!g2756) & (!g2757) & (!g2775) & (!g2776)) + ((!g2754) & (g2755) & (!g2756) & (!g2757) & (!g2775) & (g2776)) + ((!g2754) & (g2755) & (!g2756) & (!g2757) & (g2775) & (!g2776)) + ((!g2754) & (g2755) & (!g2756) & (g2757) & (!g2775) & (!g2776)) + ((!g2754) & (g2755) & (g2756) & (!g2757) & (!g2775) & (!g2776)) + ((!g2754) & (g2755) & (g2756) & (g2757) & (!g2775) & (!g2776)) + ((g2754) & (!g2755) & (!g2756) & (!g2757) & (!g2775) & (!g2776)) + ((g2754) & (!g2755) & (!g2756) & (!g2757) & (!g2775) & (g2776)) + ((g2754) & (!g2755) & (!g2756) & (!g2757) & (g2775) & (!g2776)) + ((g2754) & (!g2755) & (!g2756) & (g2757) & (!g2775) & (!g2776)) + ((g2754) & (!g2755) & (g2756) & (!g2757) & (!g2775) & (!g2776)) + ((g2754) & (!g2755) & (g2756) & (g2757) & (!g2775) & (!g2776)) + ((g2754) & (g2755) & (!g2756) & (!g2757) & (!g2775) & (!g2776)) + ((g2754) & (g2755) & (!g2756) & (!g2757) & (!g2775) & (g2776)) + ((g2754) & (g2755) & (!g2756) & (!g2757) & (g2775) & (!g2776)) + ((g2754) & (g2755) & (!g2756) & (g2757) & (!g2775) & (!g2776)) + ((g2754) & (g2755) & (g2756) & (!g2757) & (!g2775) & (!g2776)) + ((g2754) & (g2755) & (g2756) & (g2757) & (!g2775) & (!g2776)));
	assign g2798 = (((!sk[103]) & (!g2771) & (g2098)) + ((!sk[103]) & (g2771) & (g2098)) + ((sk[103]) & (!g2771) & (g2098)));
	assign g2799 = (((!g2794) & (!sk[104]) & (g2099)) + ((!g2794) & (sk[104]) & (!g2099)) + ((g2794) & (!sk[104]) & (g2099)) + ((g2794) & (sk[104]) & (g2099)));
	assign g2800 = (((!g2795) & (!g2081) & (g2125) & (!g2796) & (!g2797) & (g3116)) + ((!g2795) & (!g2081) & (g2125) & (!g2796) & (g2797) & (!g3116)) + ((!g2795) & (!g2081) & (g2125) & (g2796) & (!g2797) & (g3116)) + ((!g2795) & (!g2081) & (g2125) & (g2796) & (g2797) & (!g3116)) + ((!g2795) & (g2081) & (!g2125) & (g2796) & (!g2797) & (!g3116)) + ((!g2795) & (g2081) & (!g2125) & (g2796) & (!g2797) & (g3116)) + ((!g2795) & (g2081) & (!g2125) & (g2796) & (g2797) & (!g3116)) + ((!g2795) & (g2081) & (!g2125) & (g2796) & (g2797) & (g3116)) + ((!g2795) & (g2081) & (g2125) & (!g2796) & (!g2797) & (g3116)) + ((!g2795) & (g2081) & (g2125) & (!g2796) & (g2797) & (g3116)) + ((!g2795) & (g2081) & (g2125) & (g2796) & (!g2797) & (g3116)) + ((!g2795) & (g2081) & (g2125) & (g2796) & (g2797) & (g3116)) + ((g2795) & (!g2081) & (!g2125) & (!g2796) & (!g2797) & (!g3116)) + ((g2795) & (!g2081) & (!g2125) & (!g2796) & (!g2797) & (g3116)) + ((g2795) & (!g2081) & (!g2125) & (!g2796) & (g2797) & (!g3116)) + ((g2795) & (!g2081) & (!g2125) & (!g2796) & (g2797) & (g3116)) + ((g2795) & (!g2081) & (!g2125) & (g2796) & (!g2797) & (!g3116)) + ((g2795) & (!g2081) & (!g2125) & (g2796) & (!g2797) & (g3116)) + ((g2795) & (!g2081) & (!g2125) & (g2796) & (g2797) & (!g3116)) + ((g2795) & (!g2081) & (!g2125) & (g2796) & (g2797) & (g3116)) + ((g2795) & (!g2081) & (g2125) & (!g2796) & (!g2797) & (g3116)) + ((g2795) & (!g2081) & (g2125) & (!g2796) & (g2797) & (!g3116)) + ((g2795) & (!g2081) & (g2125) & (g2796) & (!g2797) & (g3116)) + ((g2795) & (!g2081) & (g2125) & (g2796) & (g2797) & (!g3116)) + ((g2795) & (g2081) & (!g2125) & (!g2796) & (!g2797) & (!g3116)) + ((g2795) & (g2081) & (!g2125) & (!g2796) & (!g2797) & (g3116)) + ((g2795) & (g2081) & (!g2125) & (!g2796) & (g2797) & (!g3116)) + ((g2795) & (g2081) & (!g2125) & (!g2796) & (g2797) & (g3116)) + ((g2795) & (g2081) & (g2125) & (!g2796) & (!g2797) & (g3116)) + ((g2795) & (g2081) & (g2125) & (!g2796) & (g2797) & (g3116)) + ((g2795) & (g2081) & (g2125) & (g2796) & (!g2797) & (g3116)) + ((g2795) & (g2081) & (g2125) & (g2796) & (g2797) & (g3116)));
	assign g2801 = (((!g2723) & (!g2098) & (!g2091) & (g2090) & (g2196) & (g2197)) + ((!g2723) & (!g2098) & (g2091) & (!g2090) & (!g2196) & (g2197)) + ((!g2723) & (!g2098) & (g2091) & (g2090) & (!g2196) & (g2197)) + ((!g2723) & (!g2098) & (g2091) & (g2090) & (g2196) & (g2197)) + ((!g2723) & (g2098) & (!g2091) & (!g2090) & (g2196) & (!g2197)) + ((!g2723) & (g2098) & (!g2091) & (g2090) & (g2196) & (!g2197)) + ((!g2723) & (g2098) & (!g2091) & (g2090) & (g2196) & (g2197)) + ((!g2723) & (g2098) & (g2091) & (!g2090) & (!g2196) & (g2197)) + ((!g2723) & (g2098) & (g2091) & (!g2090) & (g2196) & (!g2197)) + ((!g2723) & (g2098) & (g2091) & (g2090) & (!g2196) & (g2197)) + ((!g2723) & (g2098) & (g2091) & (g2090) & (g2196) & (!g2197)) + ((!g2723) & (g2098) & (g2091) & (g2090) & (g2196) & (g2197)) + ((g2723) & (!g2098) & (!g2091) & (!g2090) & (!g2196) & (!g2197)) + ((g2723) & (!g2098) & (!g2091) & (g2090) & (!g2196) & (!g2197)) + ((g2723) & (!g2098) & (!g2091) & (g2090) & (g2196) & (g2197)) + ((g2723) & (!g2098) & (g2091) & (!g2090) & (!g2196) & (!g2197)) + ((g2723) & (!g2098) & (g2091) & (!g2090) & (!g2196) & (g2197)) + ((g2723) & (!g2098) & (g2091) & (g2090) & (!g2196) & (!g2197)) + ((g2723) & (!g2098) & (g2091) & (g2090) & (!g2196) & (g2197)) + ((g2723) & (!g2098) & (g2091) & (g2090) & (g2196) & (g2197)) + ((g2723) & (g2098) & (!g2091) & (!g2090) & (!g2196) & (!g2197)) + ((g2723) & (g2098) & (!g2091) & (!g2090) & (g2196) & (!g2197)) + ((g2723) & (g2098) & (!g2091) & (g2090) & (!g2196) & (!g2197)) + ((g2723) & (g2098) & (!g2091) & (g2090) & (g2196) & (!g2197)) + ((g2723) & (g2098) & (!g2091) & (g2090) & (g2196) & (g2197)) + ((g2723) & (g2098) & (g2091) & (!g2090) & (!g2196) & (!g2197)) + ((g2723) & (g2098) & (g2091) & (!g2090) & (!g2196) & (g2197)) + ((g2723) & (g2098) & (g2091) & (!g2090) & (g2196) & (!g2197)) + ((g2723) & (g2098) & (g2091) & (g2090) & (!g2196) & (!g2197)) + ((g2723) & (g2098) & (g2091) & (g2090) & (!g2196) & (g2197)) + ((g2723) & (g2098) & (g2091) & (g2090) & (g2196) & (!g2197)) + ((g2723) & (g2098) & (g2091) & (g2090) & (g2196) & (g2197)));
	assign g2802 = (((!g2491) & (!g2801) & (!g2650) & (g2580) & (g2201) & (g2202)) + ((!g2491) & (!g2801) & (g2650) & (!g2580) & (!g2201) & (g2202)) + ((!g2491) & (!g2801) & (g2650) & (g2580) & (!g2201) & (g2202)) + ((!g2491) & (!g2801) & (g2650) & (g2580) & (g2201) & (g2202)) + ((!g2491) & (g2801) & (!g2650) & (!g2580) & (g2201) & (!g2202)) + ((!g2491) & (g2801) & (!g2650) & (g2580) & (g2201) & (!g2202)) + ((!g2491) & (g2801) & (!g2650) & (g2580) & (g2201) & (g2202)) + ((!g2491) & (g2801) & (g2650) & (!g2580) & (!g2201) & (g2202)) + ((!g2491) & (g2801) & (g2650) & (!g2580) & (g2201) & (!g2202)) + ((!g2491) & (g2801) & (g2650) & (g2580) & (!g2201) & (g2202)) + ((!g2491) & (g2801) & (g2650) & (g2580) & (g2201) & (!g2202)) + ((!g2491) & (g2801) & (g2650) & (g2580) & (g2201) & (g2202)) + ((g2491) & (!g2801) & (!g2650) & (!g2580) & (!g2201) & (!g2202)) + ((g2491) & (!g2801) & (!g2650) & (g2580) & (!g2201) & (!g2202)) + ((g2491) & (!g2801) & (!g2650) & (g2580) & (g2201) & (g2202)) + ((g2491) & (!g2801) & (g2650) & (!g2580) & (!g2201) & (!g2202)) + ((g2491) & (!g2801) & (g2650) & (!g2580) & (!g2201) & (g2202)) + ((g2491) & (!g2801) & (g2650) & (g2580) & (!g2201) & (!g2202)) + ((g2491) & (!g2801) & (g2650) & (g2580) & (!g2201) & (g2202)) + ((g2491) & (!g2801) & (g2650) & (g2580) & (g2201) & (g2202)) + ((g2491) & (g2801) & (!g2650) & (!g2580) & (!g2201) & (!g2202)) + ((g2491) & (g2801) & (!g2650) & (!g2580) & (g2201) & (!g2202)) + ((g2491) & (g2801) & (!g2650) & (g2580) & (!g2201) & (!g2202)) + ((g2491) & (g2801) & (!g2650) & (g2580) & (g2201) & (!g2202)) + ((g2491) & (g2801) & (!g2650) & (g2580) & (g2201) & (g2202)) + ((g2491) & (g2801) & (g2650) & (!g2580) & (!g2201) & (!g2202)) + ((g2491) & (g2801) & (g2650) & (!g2580) & (!g2201) & (g2202)) + ((g2491) & (g2801) & (g2650) & (!g2580) & (g2201) & (!g2202)) + ((g2491) & (g2801) & (g2650) & (g2580) & (!g2201) & (!g2202)) + ((g2491) & (g2801) & (g2650) & (g2580) & (!g2201) & (g2202)) + ((g2491) & (g2801) & (g2650) & (g2580) & (g2201) & (!g2202)) + ((g2491) & (g2801) & (g2650) & (g2580) & (g2201) & (g2202)));
	assign g2803 = (((!g2800) & (!g2802) & (!g2489) & (g2192) & (g2780) & (g2190)) + ((!g2800) & (!g2802) & (g2489) & (!g2192) & (!g2780) & (g2190)) + ((!g2800) & (!g2802) & (g2489) & (g2192) & (!g2780) & (g2190)) + ((!g2800) & (!g2802) & (g2489) & (g2192) & (g2780) & (g2190)) + ((!g2800) & (g2802) & (!g2489) & (!g2192) & (g2780) & (!g2190)) + ((!g2800) & (g2802) & (!g2489) & (g2192) & (g2780) & (!g2190)) + ((!g2800) & (g2802) & (!g2489) & (g2192) & (g2780) & (g2190)) + ((!g2800) & (g2802) & (g2489) & (!g2192) & (!g2780) & (g2190)) + ((!g2800) & (g2802) & (g2489) & (!g2192) & (g2780) & (!g2190)) + ((!g2800) & (g2802) & (g2489) & (g2192) & (!g2780) & (g2190)) + ((!g2800) & (g2802) & (g2489) & (g2192) & (g2780) & (!g2190)) + ((!g2800) & (g2802) & (g2489) & (g2192) & (g2780) & (g2190)) + ((g2800) & (!g2802) & (!g2489) & (!g2192) & (!g2780) & (!g2190)) + ((g2800) & (!g2802) & (!g2489) & (g2192) & (!g2780) & (!g2190)) + ((g2800) & (!g2802) & (!g2489) & (g2192) & (g2780) & (g2190)) + ((g2800) & (!g2802) & (g2489) & (!g2192) & (!g2780) & (!g2190)) + ((g2800) & (!g2802) & (g2489) & (!g2192) & (!g2780) & (g2190)) + ((g2800) & (!g2802) & (g2489) & (g2192) & (!g2780) & (!g2190)) + ((g2800) & (!g2802) & (g2489) & (g2192) & (!g2780) & (g2190)) + ((g2800) & (!g2802) & (g2489) & (g2192) & (g2780) & (g2190)) + ((g2800) & (g2802) & (!g2489) & (!g2192) & (!g2780) & (!g2190)) + ((g2800) & (g2802) & (!g2489) & (!g2192) & (g2780) & (!g2190)) + ((g2800) & (g2802) & (!g2489) & (g2192) & (!g2780) & (!g2190)) + ((g2800) & (g2802) & (!g2489) & (g2192) & (g2780) & (!g2190)) + ((g2800) & (g2802) & (!g2489) & (g2192) & (g2780) & (g2190)) + ((g2800) & (g2802) & (g2489) & (!g2192) & (!g2780) & (!g2190)) + ((g2800) & (g2802) & (g2489) & (!g2192) & (!g2780) & (g2190)) + ((g2800) & (g2802) & (g2489) & (!g2192) & (g2780) & (!g2190)) + ((g2800) & (g2802) & (g2489) & (g2192) & (!g2780) & (!g2190)) + ((g2800) & (g2802) & (g2489) & (g2192) & (!g2780) & (g2190)) + ((g2800) & (g2802) & (g2489) & (g2192) & (g2780) & (!g2190)) + ((g2800) & (g2802) & (g2489) & (g2192) & (g2780) & (g2190)));
	assign g2804 = (((!g2081) & (!g2124) & (!g2770) & (!g2794) & (!g2803) & (!g2099)) + ((!g2081) & (!g2124) & (!g2770) & (!g2794) & (!g2803) & (g2099)) + ((!g2081) & (!g2124) & (!g2770) & (g2794) & (!g2803) & (!g2099)) + ((!g2081) & (!g2124) & (!g2770) & (g2794) & (!g2803) & (g2099)) + ((!g2081) & (!g2124) & (g2770) & (!g2794) & (!g2803) & (!g2099)) + ((!g2081) & (!g2124) & (g2770) & (!g2794) & (g2803) & (!g2099)) + ((!g2081) & (!g2124) & (g2770) & (g2794) & (!g2803) & (!g2099)) + ((!g2081) & (!g2124) & (g2770) & (g2794) & (g2803) & (!g2099)) + ((!g2081) & (g2124) & (!g2770) & (!g2794) & (!g2803) & (!g2099)) + ((!g2081) & (g2124) & (!g2770) & (!g2794) & (g2803) & (!g2099)) + ((!g2081) & (g2124) & (g2770) & (!g2794) & (!g2803) & (!g2099)) + ((!g2081) & (g2124) & (g2770) & (!g2794) & (g2803) & (!g2099)) + ((!g2081) & (g2124) & (g2770) & (g2794) & (!g2803) & (!g2099)) + ((!g2081) & (g2124) & (g2770) & (g2794) & (g2803) & (!g2099)) + ((g2081) & (!g2124) & (!g2770) & (!g2794) & (!g2803) & (!g2099)) + ((g2081) & (!g2124) & (!g2770) & (!g2794) & (!g2803) & (g2099)) + ((g2081) & (!g2124) & (!g2770) & (g2794) & (!g2803) & (!g2099)) + ((g2081) & (!g2124) & (!g2770) & (g2794) & (!g2803) & (g2099)) + ((g2081) & (!g2124) & (g2770) & (!g2794) & (!g2803) & (!g2099)) + ((g2081) & (!g2124) & (g2770) & (!g2794) & (g2803) & (!g2099)) + ((g2081) & (!g2124) & (g2770) & (g2794) & (!g2803) & (!g2099)) + ((g2081) & (!g2124) & (g2770) & (g2794) & (g2803) & (!g2099)) + ((g2081) & (g2124) & (!g2770) & (!g2794) & (!g2803) & (!g2099)) + ((g2081) & (g2124) & (!g2770) & (!g2794) & (g2803) & (!g2099)) + ((g2081) & (g2124) & (!g2770) & (g2794) & (!g2803) & (g2099)) + ((g2081) & (g2124) & (!g2770) & (g2794) & (g2803) & (g2099)) + ((g2081) & (g2124) & (g2770) & (!g2794) & (!g2803) & (!g2099)) + ((g2081) & (g2124) & (g2770) & (!g2794) & (g2803) & (!g2099)) + ((g2081) & (g2124) & (g2770) & (g2794) & (!g2803) & (!g2099)) + ((g2081) & (g2124) & (g2770) & (g2794) & (g2803) & (!g2099)));
	assign g2805 = (((!g2804) & (!dmem_dat_ix29x) & (!g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2804) & (!dmem_dat_ix29x) & (!g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2804) & (!dmem_dat_ix29x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((!g2804) & (!dmem_dat_ix29x) & (g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2804) & (!dmem_dat_ix29x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((!g2804) & (!dmem_dat_ix29x) & (g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2804) & (!dmem_dat_ix29x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((!g2804) & (!dmem_dat_ix29x) & (g2783) & (g2784) & (g2785) & (g2786)) + ((!g2804) & (dmem_dat_ix29x) & (!g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2804) & (dmem_dat_ix29x) & (!g2783) & (!g2784) & (g2785) & (!g2786)) + ((!g2804) & (dmem_dat_ix29x) & (!g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2804) & (dmem_dat_ix29x) & (!g2783) & (g2784) & (g2785) & (!g2786)) + ((!g2804) & (dmem_dat_ix29x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((!g2804) & (dmem_dat_ix29x) & (g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2804) & (dmem_dat_ix29x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((!g2804) & (dmem_dat_ix29x) & (g2783) & (!g2784) & (g2785) & (!g2786)) + ((!g2804) & (dmem_dat_ix29x) & (g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2804) & (dmem_dat_ix29x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((!g2804) & (dmem_dat_ix29x) & (g2783) & (g2784) & (g2785) & (!g2786)) + ((!g2804) & (dmem_dat_ix29x) & (g2783) & (g2784) & (g2785) & (g2786)) + ((g2804) & (!dmem_dat_ix29x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((g2804) & (!dmem_dat_ix29x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((g2804) & (!dmem_dat_ix29x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((g2804) & (!dmem_dat_ix29x) & (g2783) & (g2784) & (g2785) & (g2786)) + ((g2804) & (dmem_dat_ix29x) & (!g2783) & (!g2784) & (g2785) & (!g2786)) + ((g2804) & (dmem_dat_ix29x) & (!g2783) & (g2784) & (g2785) & (!g2786)) + ((g2804) & (dmem_dat_ix29x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((g2804) & (dmem_dat_ix29x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((g2804) & (dmem_dat_ix29x) & (g2783) & (!g2784) & (g2785) & (!g2786)) + ((g2804) & (dmem_dat_ix29x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((g2804) & (dmem_dat_ix29x) & (g2783) & (g2784) & (g2785) & (!g2786)) + ((g2804) & (dmem_dat_ix29x) & (g2783) & (g2784) & (g2785) & (g2786)));
	assign g2806 = (((!g1455) & (!g2788) & (sk[111]) & (g1500)) + ((!g1455) & (g2788) & (!sk[111]) & (!g1500)) + ((!g1455) & (g2788) & (!sk[111]) & (g1500)) + ((!g1455) & (g2788) & (sk[111]) & (g1500)) + ((g1455) & (!g2788) & (!sk[111]) & (!g1500)) + ((g1455) & (!g2788) & (!sk[111]) & (g1500)) + ((g1455) & (!g2788) & (sk[111]) & (g1500)) + ((g1455) & (g2788) & (!sk[111]) & (!g1500)) + ((g1455) & (g2788) & (!sk[111]) & (g1500)) + ((g1455) & (g2788) & (sk[111]) & (!g1500)));
	assign g2807 = (((!g107) & (!g1410) & (!g2765) & (!g1455) & (sk[112]) & (g1500)) + ((!g107) & (!g1410) & (!g2765) & (g1455) & (!sk[112]) & (!g1500)) + ((!g107) & (!g1410) & (!g2765) & (g1455) & (!sk[112]) & (g1500)) + ((!g107) & (!g1410) & (!g2765) & (g1455) & (sk[112]) & (g1500)) + ((!g107) & (!g1410) & (g2765) & (!g1455) & (!sk[112]) & (!g1500)) + ((!g107) & (!g1410) & (g2765) & (!g1455) & (!sk[112]) & (g1500)) + ((!g107) & (!g1410) & (g2765) & (!g1455) & (sk[112]) & (g1500)) + ((!g107) & (!g1410) & (g2765) & (g1455) & (!sk[112]) & (!g1500)) + ((!g107) & (!g1410) & (g2765) & (g1455) & (!sk[112]) & (g1500)) + ((!g107) & (!g1410) & (g2765) & (g1455) & (sk[112]) & (g1500)) + ((!g107) & (g1410) & (!g2765) & (!g1455) & (sk[112]) & (g1500)) + ((!g107) & (g1410) & (!g2765) & (g1455) & (!sk[112]) & (!g1500)) + ((!g107) & (g1410) & (!g2765) & (g1455) & (!sk[112]) & (g1500)) + ((!g107) & (g1410) & (!g2765) & (g1455) & (sk[112]) & (g1500)) + ((!g107) & (g1410) & (g2765) & (!g1455) & (!sk[112]) & (!g1500)) + ((!g107) & (g1410) & (g2765) & (!g1455) & (!sk[112]) & (g1500)) + ((!g107) & (g1410) & (g2765) & (!g1455) & (sk[112]) & (g1500)) + ((!g107) & (g1410) & (g2765) & (g1455) & (!sk[112]) & (!g1500)) + ((!g107) & (g1410) & (g2765) & (g1455) & (!sk[112]) & (g1500)) + ((!g107) & (g1410) & (g2765) & (g1455) & (sk[112]) & (!g1500)) + ((g107) & (!g1410) & (!g2765) & (!g1455) & (!sk[112]) & (!g1500)) + ((g107) & (!g1410) & (!g2765) & (!g1455) & (!sk[112]) & (g1500)) + ((g107) & (!g1410) & (!g2765) & (!g1455) & (sk[112]) & (!g1500)) + ((g107) & (!g1410) & (!g2765) & (g1455) & (!sk[112]) & (!g1500)) + ((g107) & (!g1410) & (!g2765) & (g1455) & (!sk[112]) & (g1500)) + ((g107) & (!g1410) & (!g2765) & (g1455) & (sk[112]) & (g1500)) + ((g107) & (!g1410) & (g2765) & (!g1455) & (!sk[112]) & (!g1500)) + ((g107) & (!g1410) & (g2765) & (!g1455) & (!sk[112]) & (g1500)) + ((g107) & (!g1410) & (g2765) & (!g1455) & (sk[112]) & (g1500)) + ((g107) & (!g1410) & (g2765) & (g1455) & (!sk[112]) & (!g1500)) + ((g107) & (!g1410) & (g2765) & (g1455) & (!sk[112]) & (g1500)) + ((g107) & (!g1410) & (g2765) & (g1455) & (sk[112]) & (g1500)) + ((g107) & (g1410) & (!g2765) & (!g1455) & (!sk[112]) & (!g1500)) + ((g107) & (g1410) & (!g2765) & (!g1455) & (!sk[112]) & (g1500)) + ((g107) & (g1410) & (!g2765) & (!g1455) & (sk[112]) & (g1500)) + ((g107) & (g1410) & (!g2765) & (g1455) & (!sk[112]) & (!g1500)) + ((g107) & (g1410) & (!g2765) & (g1455) & (!sk[112]) & (g1500)) + ((g107) & (g1410) & (!g2765) & (g1455) & (sk[112]) & (g1500)) + ((g107) & (g1410) & (g2765) & (!g1455) & (!sk[112]) & (!g1500)) + ((g107) & (g1410) & (g2765) & (!g1455) & (!sk[112]) & (g1500)) + ((g107) & (g1410) & (g2765) & (!g1455) & (sk[112]) & (g1500)) + ((g107) & (g1410) & (g2765) & (g1455) & (!sk[112]) & (!g1500)) + ((g107) & (g1410) & (g2765) & (g1455) & (!sk[112]) & (g1500)) + ((g107) & (g1410) & (g2765) & (g1455) & (sk[112]) & (g1500)));
	assign g5053 = (((!g2921) & (!g3109) & (sk[113]) & (g2808)) + ((!g2921) & (g3109) & (!sk[113]) & (!g2808)) + ((!g2921) & (g3109) & (!sk[113]) & (g2808)) + ((!g2921) & (g3109) & (sk[113]) & (g2808)) + ((g2921) & (!g3109) & (!sk[113]) & (!g2808)) + ((g2921) & (!g3109) & (!sk[113]) & (g2808)) + ((g2921) & (g3109) & (!sk[113]) & (!g2808)) + ((g2921) & (g3109) & (!sk[113]) & (g2808)) + ((g2921) & (g3109) & (sk[113]) & (!g2808)) + ((g2921) & (g3109) & (sk[113]) & (g2808)));
	assign g2809 = (((!sk[114]) & (!g1981) & (!g2033) & (!g2034) & (g2807) & (!g2808)) + ((!sk[114]) & (!g1981) & (!g2033) & (!g2034) & (g2807) & (g2808)) + ((!sk[114]) & (!g1981) & (!g2033) & (g2034) & (!g2807) & (!g2808)) + ((!sk[114]) & (!g1981) & (!g2033) & (g2034) & (!g2807) & (g2808)) + ((!sk[114]) & (!g1981) & (!g2033) & (g2034) & (g2807) & (!g2808)) + ((!sk[114]) & (!g1981) & (!g2033) & (g2034) & (g2807) & (g2808)) + ((!sk[114]) & (!g1981) & (g2033) & (!g2034) & (g2807) & (!g2808)) + ((!sk[114]) & (!g1981) & (g2033) & (!g2034) & (g2807) & (g2808)) + ((!sk[114]) & (!g1981) & (g2033) & (g2034) & (!g2807) & (!g2808)) + ((!sk[114]) & (!g1981) & (g2033) & (g2034) & (!g2807) & (g2808)) + ((!sk[114]) & (!g1981) & (g2033) & (g2034) & (g2807) & (!g2808)) + ((!sk[114]) & (!g1981) & (g2033) & (g2034) & (g2807) & (g2808)) + ((!sk[114]) & (g1981) & (!g2033) & (!g2034) & (!g2807) & (!g2808)) + ((!sk[114]) & (g1981) & (!g2033) & (!g2034) & (!g2807) & (g2808)) + ((!sk[114]) & (g1981) & (!g2033) & (!g2034) & (g2807) & (!g2808)) + ((!sk[114]) & (g1981) & (!g2033) & (!g2034) & (g2807) & (g2808)) + ((!sk[114]) & (g1981) & (!g2033) & (g2034) & (!g2807) & (!g2808)) + ((!sk[114]) & (g1981) & (!g2033) & (g2034) & (!g2807) & (g2808)) + ((!sk[114]) & (g1981) & (!g2033) & (g2034) & (g2807) & (!g2808)) + ((!sk[114]) & (g1981) & (!g2033) & (g2034) & (g2807) & (g2808)) + ((!sk[114]) & (g1981) & (g2033) & (!g2034) & (!g2807) & (!g2808)) + ((!sk[114]) & (g1981) & (g2033) & (!g2034) & (!g2807) & (g2808)) + ((!sk[114]) & (g1981) & (g2033) & (!g2034) & (g2807) & (!g2808)) + ((!sk[114]) & (g1981) & (g2033) & (!g2034) & (g2807) & (g2808)) + ((!sk[114]) & (g1981) & (g2033) & (g2034) & (!g2807) & (!g2808)) + ((!sk[114]) & (g1981) & (g2033) & (g2034) & (!g2807) & (g2808)) + ((!sk[114]) & (g1981) & (g2033) & (g2034) & (g2807) & (!g2808)) + ((!sk[114]) & (g1981) & (g2033) & (g2034) & (g2807) & (g2808)) + ((sk[114]) & (!g1981) & (!g2033) & (!g2034) & (!g2807) & (g2808)) + ((sk[114]) & (!g1981) & (!g2033) & (!g2034) & (g2807) & (g2808)) + ((sk[114]) & (!g1981) & (g2033) & (!g2034) & (g2807) & (!g2808)) + ((sk[114]) & (!g1981) & (g2033) & (!g2034) & (g2807) & (g2808)) + ((sk[114]) & (g1981) & (!g2033) & (!g2034) & (!g2807) & (g2808)) + ((sk[114]) & (g1981) & (!g2033) & (!g2034) & (g2807) & (g2808)) + ((sk[114]) & (g1981) & (!g2033) & (g2034) & (!g2807) & (!g2808)) + ((sk[114]) & (g1981) & (!g2033) & (g2034) & (!g2807) & (g2808)) + ((sk[114]) & (g1981) & (!g2033) & (g2034) & (g2807) & (!g2808)) + ((sk[114]) & (g1981) & (!g2033) & (g2034) & (g2807) & (g2808)) + ((sk[114]) & (g1981) & (g2033) & (!g2034) & (g2807) & (!g2808)) + ((sk[114]) & (g1981) & (g2033) & (!g2034) & (g2807) & (g2808)));
	assign g2810 = (((!sk[115]) & (!g2329) & (!g2029) & (!g2408) & (g2806) & (!g2809)) + ((!sk[115]) & (!g2329) & (!g2029) & (!g2408) & (g2806) & (g2809)) + ((!sk[115]) & (!g2329) & (!g2029) & (g2408) & (!g2806) & (!g2809)) + ((!sk[115]) & (!g2329) & (!g2029) & (g2408) & (!g2806) & (g2809)) + ((!sk[115]) & (!g2329) & (!g2029) & (g2408) & (g2806) & (!g2809)) + ((!sk[115]) & (!g2329) & (!g2029) & (g2408) & (g2806) & (g2809)) + ((!sk[115]) & (!g2329) & (g2029) & (!g2408) & (g2806) & (!g2809)) + ((!sk[115]) & (!g2329) & (g2029) & (!g2408) & (g2806) & (g2809)) + ((!sk[115]) & (!g2329) & (g2029) & (g2408) & (!g2806) & (!g2809)) + ((!sk[115]) & (!g2329) & (g2029) & (g2408) & (!g2806) & (g2809)) + ((!sk[115]) & (!g2329) & (g2029) & (g2408) & (g2806) & (!g2809)) + ((!sk[115]) & (!g2329) & (g2029) & (g2408) & (g2806) & (g2809)) + ((!sk[115]) & (g2329) & (!g2029) & (!g2408) & (!g2806) & (!g2809)) + ((!sk[115]) & (g2329) & (!g2029) & (!g2408) & (!g2806) & (g2809)) + ((!sk[115]) & (g2329) & (!g2029) & (!g2408) & (g2806) & (!g2809)) + ((!sk[115]) & (g2329) & (!g2029) & (!g2408) & (g2806) & (g2809)) + ((!sk[115]) & (g2329) & (!g2029) & (g2408) & (!g2806) & (!g2809)) + ((!sk[115]) & (g2329) & (!g2029) & (g2408) & (!g2806) & (g2809)) + ((!sk[115]) & (g2329) & (!g2029) & (g2408) & (g2806) & (!g2809)) + ((!sk[115]) & (g2329) & (!g2029) & (g2408) & (g2806) & (g2809)) + ((!sk[115]) & (g2329) & (g2029) & (!g2408) & (!g2806) & (!g2809)) + ((!sk[115]) & (g2329) & (g2029) & (!g2408) & (!g2806) & (g2809)) + ((!sk[115]) & (g2329) & (g2029) & (!g2408) & (g2806) & (!g2809)) + ((!sk[115]) & (g2329) & (g2029) & (!g2408) & (g2806) & (g2809)) + ((!sk[115]) & (g2329) & (g2029) & (g2408) & (!g2806) & (!g2809)) + ((!sk[115]) & (g2329) & (g2029) & (g2408) & (!g2806) & (g2809)) + ((!sk[115]) & (g2329) & (g2029) & (g2408) & (g2806) & (!g2809)) + ((!sk[115]) & (g2329) & (g2029) & (g2408) & (g2806) & (g2809)) + ((sk[115]) & (g2329) & (!g2029) & (g2408) & (!g2806) & (g2809)) + ((sk[115]) & (g2329) & (!g2029) & (g2408) & (g2806) & (g2809)) + ((sk[115]) & (g2329) & (g2029) & (g2408) & (g2806) & (!g2809)) + ((sk[115]) & (g2329) & (g2029) & (g2408) & (g2806) & (g2809)));
	assign g2812 = (((!g2100) & (!sk[116]) & (g2811)) + ((!g2100) & (sk[116]) & (g2811)) + ((g2100) & (!sk[116]) & (g2811)) + ((g2100) & (sk[116]) & (!g2811)));
	assign g2813 = (((!g2098) & (!g2099) & (!g2771) & (!g2772) & (!g2794) & (g2812)) + ((!g2098) & (!g2099) & (!g2771) & (!g2772) & (g2794) & (g2812)) + ((!g2098) & (!g2099) & (!g2771) & (g2772) & (!g2794) & (g2812)) + ((!g2098) & (!g2099) & (!g2771) & (g2772) & (g2794) & (g2812)) + ((!g2098) & (!g2099) & (g2771) & (!g2772) & (!g2794) & (g2812)) + ((!g2098) & (!g2099) & (g2771) & (!g2772) & (g2794) & (g2812)) + ((!g2098) & (!g2099) & (g2771) & (g2772) & (!g2794) & (g2812)) + ((!g2098) & (!g2099) & (g2771) & (g2772) & (g2794) & (!g2812)) + ((!g2098) & (g2099) & (!g2771) & (!g2772) & (!g2794) & (g2812)) + ((!g2098) & (g2099) & (!g2771) & (!g2772) & (g2794) & (!g2812)) + ((!g2098) & (g2099) & (!g2771) & (g2772) & (!g2794) & (g2812)) + ((!g2098) & (g2099) & (!g2771) & (g2772) & (g2794) & (!g2812)) + ((!g2098) & (g2099) & (g2771) & (!g2772) & (!g2794) & (g2812)) + ((!g2098) & (g2099) & (g2771) & (!g2772) & (g2794) & (!g2812)) + ((!g2098) & (g2099) & (g2771) & (g2772) & (!g2794) & (!g2812)) + ((!g2098) & (g2099) & (g2771) & (g2772) & (g2794) & (!g2812)) + ((g2098) & (!g2099) & (!g2771) & (!g2772) & (!g2794) & (g2812)) + ((g2098) & (!g2099) & (!g2771) & (!g2772) & (g2794) & (g2812)) + ((g2098) & (!g2099) & (!g2771) & (g2772) & (!g2794) & (g2812)) + ((g2098) & (!g2099) & (!g2771) & (g2772) & (g2794) & (!g2812)) + ((g2098) & (!g2099) & (g2771) & (!g2772) & (!g2794) & (g2812)) + ((g2098) & (!g2099) & (g2771) & (!g2772) & (g2794) & (!g2812)) + ((g2098) & (!g2099) & (g2771) & (g2772) & (!g2794) & (g2812)) + ((g2098) & (!g2099) & (g2771) & (g2772) & (g2794) & (!g2812)) + ((g2098) & (g2099) & (!g2771) & (!g2772) & (!g2794) & (g2812)) + ((g2098) & (g2099) & (!g2771) & (!g2772) & (g2794) & (!g2812)) + ((g2098) & (g2099) & (!g2771) & (g2772) & (!g2794) & (!g2812)) + ((g2098) & (g2099) & (!g2771) & (g2772) & (g2794) & (!g2812)) + ((g2098) & (g2099) & (g2771) & (!g2772) & (!g2794) & (!g2812)) + ((g2098) & (g2099) & (g2771) & (!g2772) & (g2794) & (!g2812)) + ((g2098) & (g2099) & (g2771) & (g2772) & (!g2794) & (!g2812)) + ((g2098) & (g2099) & (g2771) & (g2772) & (g2794) & (!g2812)));
	assign g2814 = (((!g2794) & (!sk[118]) & (g2099)) + ((!g2794) & (sk[118]) & (g2099)) + ((g2794) & (!sk[118]) & (g2099)));
	assign g2815 = (((!sk[119]) & (!g2811) & (g2100)) + ((!sk[119]) & (g2811) & (g2100)) + ((sk[119]) & (!g2811) & (!g2100)) + ((sk[119]) & (g2811) & (g2100)));
	assign g2816 = (((!g2813) & (!g2125) & (!g2797) & (g2795) & (!g3131) & (g3132)) + ((!g2813) & (!g2125) & (!g2797) & (g2795) & (g3131) & (g3132)) + ((!g2813) & (!g2125) & (g2797) & (g2795) & (!g3131) & (g3132)) + ((!g2813) & (!g2125) & (g2797) & (g2795) & (g3131) & (g3132)) + ((!g2813) & (g2125) & (!g2797) & (!g2795) & (!g3131) & (!g3132)) + ((!g2813) & (g2125) & (!g2797) & (!g2795) & (g3131) & (!g3132)) + ((!g2813) & (g2125) & (!g2797) & (g2795) & (!g3131) & (!g3132)) + ((!g2813) & (g2125) & (!g2797) & (g2795) & (g3131) & (!g3132)) + ((!g2813) & (g2125) & (g2797) & (!g2795) & (g3131) & (!g3132)) + ((!g2813) & (g2125) & (g2797) & (!g2795) & (g3131) & (g3132)) + ((!g2813) & (g2125) & (g2797) & (g2795) & (g3131) & (!g3132)) + ((!g2813) & (g2125) & (g2797) & (g2795) & (g3131) & (g3132)) + ((g2813) & (!g2125) & (!g2797) & (!g2795) & (!g3131) & (!g3132)) + ((g2813) & (!g2125) & (!g2797) & (!g2795) & (!g3131) & (g3132)) + ((g2813) & (!g2125) & (!g2797) & (!g2795) & (g3131) & (!g3132)) + ((g2813) & (!g2125) & (!g2797) & (!g2795) & (g3131) & (g3132)) + ((g2813) & (!g2125) & (!g2797) & (g2795) & (!g3131) & (!g3132)) + ((g2813) & (!g2125) & (!g2797) & (g2795) & (g3131) & (!g3132)) + ((g2813) & (!g2125) & (g2797) & (!g2795) & (!g3131) & (!g3132)) + ((g2813) & (!g2125) & (g2797) & (!g2795) & (!g3131) & (g3132)) + ((g2813) & (!g2125) & (g2797) & (!g2795) & (g3131) & (!g3132)) + ((g2813) & (!g2125) & (g2797) & (!g2795) & (g3131) & (g3132)) + ((g2813) & (!g2125) & (g2797) & (g2795) & (!g3131) & (!g3132)) + ((g2813) & (!g2125) & (g2797) & (g2795) & (g3131) & (!g3132)) + ((g2813) & (g2125) & (!g2797) & (!g2795) & (!g3131) & (!g3132)) + ((g2813) & (g2125) & (!g2797) & (!g2795) & (g3131) & (!g3132)) + ((g2813) & (g2125) & (!g2797) & (g2795) & (!g3131) & (!g3132)) + ((g2813) & (g2125) & (!g2797) & (g2795) & (g3131) & (!g3132)) + ((g2813) & (g2125) & (g2797) & (!g2795) & (g3131) & (!g3132)) + ((g2813) & (g2125) & (g2797) & (!g2795) & (g3131) & (g3132)) + ((g2813) & (g2125) & (g2797) & (g2795) & (g3131) & (!g3132)) + ((g2813) & (g2125) & (g2797) & (g2795) & (g3131) & (g3132)));
	assign g2817 = (((!g2742) & (!g2099) & (!g2098) & (g2091) & (g2196) & (g2197)) + ((!g2742) & (!g2099) & (g2098) & (!g2091) & (!g2196) & (g2197)) + ((!g2742) & (!g2099) & (g2098) & (g2091) & (!g2196) & (g2197)) + ((!g2742) & (!g2099) & (g2098) & (g2091) & (g2196) & (g2197)) + ((!g2742) & (g2099) & (!g2098) & (!g2091) & (g2196) & (!g2197)) + ((!g2742) & (g2099) & (!g2098) & (g2091) & (g2196) & (!g2197)) + ((!g2742) & (g2099) & (!g2098) & (g2091) & (g2196) & (g2197)) + ((!g2742) & (g2099) & (g2098) & (!g2091) & (!g2196) & (g2197)) + ((!g2742) & (g2099) & (g2098) & (!g2091) & (g2196) & (!g2197)) + ((!g2742) & (g2099) & (g2098) & (g2091) & (!g2196) & (g2197)) + ((!g2742) & (g2099) & (g2098) & (g2091) & (g2196) & (!g2197)) + ((!g2742) & (g2099) & (g2098) & (g2091) & (g2196) & (g2197)) + ((g2742) & (!g2099) & (!g2098) & (!g2091) & (!g2196) & (!g2197)) + ((g2742) & (!g2099) & (!g2098) & (g2091) & (!g2196) & (!g2197)) + ((g2742) & (!g2099) & (!g2098) & (g2091) & (g2196) & (g2197)) + ((g2742) & (!g2099) & (g2098) & (!g2091) & (!g2196) & (!g2197)) + ((g2742) & (!g2099) & (g2098) & (!g2091) & (!g2196) & (g2197)) + ((g2742) & (!g2099) & (g2098) & (g2091) & (!g2196) & (!g2197)) + ((g2742) & (!g2099) & (g2098) & (g2091) & (!g2196) & (g2197)) + ((g2742) & (!g2099) & (g2098) & (g2091) & (g2196) & (g2197)) + ((g2742) & (g2099) & (!g2098) & (!g2091) & (!g2196) & (!g2197)) + ((g2742) & (g2099) & (!g2098) & (!g2091) & (g2196) & (!g2197)) + ((g2742) & (g2099) & (!g2098) & (g2091) & (!g2196) & (!g2197)) + ((g2742) & (g2099) & (!g2098) & (g2091) & (g2196) & (!g2197)) + ((g2742) & (g2099) & (!g2098) & (g2091) & (g2196) & (g2197)) + ((g2742) & (g2099) & (g2098) & (!g2091) & (!g2196) & (!g2197)) + ((g2742) & (g2099) & (g2098) & (!g2091) & (!g2196) & (g2197)) + ((g2742) & (g2099) & (g2098) & (!g2091) & (g2196) & (!g2197)) + ((g2742) & (g2099) & (g2098) & (g2091) & (!g2196) & (!g2197)) + ((g2742) & (g2099) & (g2098) & (g2091) & (!g2196) & (g2197)) + ((g2742) & (g2099) & (g2098) & (g2091) & (g2196) & (!g2197)) + ((g2742) & (g2099) & (g2098) & (g2091) & (g2196) & (g2197)));
	assign g2818 = (((!g2515) & (!g2817) & (!g2669) & (g2595) & (g2201) & (g2202)) + ((!g2515) & (!g2817) & (g2669) & (!g2595) & (!g2201) & (g2202)) + ((!g2515) & (!g2817) & (g2669) & (g2595) & (!g2201) & (g2202)) + ((!g2515) & (!g2817) & (g2669) & (g2595) & (g2201) & (g2202)) + ((!g2515) & (g2817) & (!g2669) & (!g2595) & (g2201) & (!g2202)) + ((!g2515) & (g2817) & (!g2669) & (g2595) & (g2201) & (!g2202)) + ((!g2515) & (g2817) & (!g2669) & (g2595) & (g2201) & (g2202)) + ((!g2515) & (g2817) & (g2669) & (!g2595) & (!g2201) & (g2202)) + ((!g2515) & (g2817) & (g2669) & (!g2595) & (g2201) & (!g2202)) + ((!g2515) & (g2817) & (g2669) & (g2595) & (!g2201) & (g2202)) + ((!g2515) & (g2817) & (g2669) & (g2595) & (g2201) & (!g2202)) + ((!g2515) & (g2817) & (g2669) & (g2595) & (g2201) & (g2202)) + ((g2515) & (!g2817) & (!g2669) & (!g2595) & (!g2201) & (!g2202)) + ((g2515) & (!g2817) & (!g2669) & (g2595) & (!g2201) & (!g2202)) + ((g2515) & (!g2817) & (!g2669) & (g2595) & (g2201) & (g2202)) + ((g2515) & (!g2817) & (g2669) & (!g2595) & (!g2201) & (!g2202)) + ((g2515) & (!g2817) & (g2669) & (!g2595) & (!g2201) & (g2202)) + ((g2515) & (!g2817) & (g2669) & (g2595) & (!g2201) & (!g2202)) + ((g2515) & (!g2817) & (g2669) & (g2595) & (!g2201) & (g2202)) + ((g2515) & (!g2817) & (g2669) & (g2595) & (g2201) & (g2202)) + ((g2515) & (g2817) & (!g2669) & (!g2595) & (!g2201) & (!g2202)) + ((g2515) & (g2817) & (!g2669) & (!g2595) & (g2201) & (!g2202)) + ((g2515) & (g2817) & (!g2669) & (g2595) & (!g2201) & (!g2202)) + ((g2515) & (g2817) & (!g2669) & (g2595) & (g2201) & (!g2202)) + ((g2515) & (g2817) & (!g2669) & (g2595) & (g2201) & (g2202)) + ((g2515) & (g2817) & (g2669) & (!g2595) & (!g2201) & (!g2202)) + ((g2515) & (g2817) & (g2669) & (!g2595) & (!g2201) & (g2202)) + ((g2515) & (g2817) & (g2669) & (!g2595) & (g2201) & (!g2202)) + ((g2515) & (g2817) & (g2669) & (g2595) & (!g2201) & (!g2202)) + ((g2515) & (g2817) & (g2669) & (g2595) & (!g2201) & (g2202)) + ((g2515) & (g2817) & (g2669) & (g2595) & (g2201) & (!g2202)) + ((g2515) & (g2817) & (g2669) & (g2595) & (g2201) & (g2202)));
	assign g2819 = (((!g2816) & (!g2818) & (!g2516) & (g2192) & (g2780) & (g2190)) + ((!g2816) & (!g2818) & (g2516) & (!g2192) & (!g2780) & (g2190)) + ((!g2816) & (!g2818) & (g2516) & (g2192) & (!g2780) & (g2190)) + ((!g2816) & (!g2818) & (g2516) & (g2192) & (g2780) & (g2190)) + ((!g2816) & (g2818) & (!g2516) & (!g2192) & (g2780) & (!g2190)) + ((!g2816) & (g2818) & (!g2516) & (g2192) & (g2780) & (!g2190)) + ((!g2816) & (g2818) & (!g2516) & (g2192) & (g2780) & (g2190)) + ((!g2816) & (g2818) & (g2516) & (!g2192) & (!g2780) & (g2190)) + ((!g2816) & (g2818) & (g2516) & (!g2192) & (g2780) & (!g2190)) + ((!g2816) & (g2818) & (g2516) & (g2192) & (!g2780) & (g2190)) + ((!g2816) & (g2818) & (g2516) & (g2192) & (g2780) & (!g2190)) + ((!g2816) & (g2818) & (g2516) & (g2192) & (g2780) & (g2190)) + ((g2816) & (!g2818) & (!g2516) & (!g2192) & (!g2780) & (!g2190)) + ((g2816) & (!g2818) & (!g2516) & (g2192) & (!g2780) & (!g2190)) + ((g2816) & (!g2818) & (!g2516) & (g2192) & (g2780) & (g2190)) + ((g2816) & (!g2818) & (g2516) & (!g2192) & (!g2780) & (!g2190)) + ((g2816) & (!g2818) & (g2516) & (!g2192) & (!g2780) & (g2190)) + ((g2816) & (!g2818) & (g2516) & (g2192) & (!g2780) & (!g2190)) + ((g2816) & (!g2818) & (g2516) & (g2192) & (!g2780) & (g2190)) + ((g2816) & (!g2818) & (g2516) & (g2192) & (g2780) & (g2190)) + ((g2816) & (g2818) & (!g2516) & (!g2192) & (!g2780) & (!g2190)) + ((g2816) & (g2818) & (!g2516) & (!g2192) & (g2780) & (!g2190)) + ((g2816) & (g2818) & (!g2516) & (g2192) & (!g2780) & (!g2190)) + ((g2816) & (g2818) & (!g2516) & (g2192) & (g2780) & (!g2190)) + ((g2816) & (g2818) & (!g2516) & (g2192) & (g2780) & (g2190)) + ((g2816) & (g2818) & (g2516) & (!g2192) & (!g2780) & (!g2190)) + ((g2816) & (g2818) & (g2516) & (!g2192) & (!g2780) & (g2190)) + ((g2816) & (g2818) & (g2516) & (!g2192) & (g2780) & (!g2190)) + ((g2816) & (g2818) & (g2516) & (g2192) & (!g2780) & (!g2190)) + ((g2816) & (g2818) & (g2516) & (g2192) & (!g2780) & (g2190)) + ((g2816) & (g2818) & (g2516) & (g2192) & (g2780) & (!g2190)) + ((g2816) & (g2818) & (g2516) & (g2192) & (g2780) & (g2190)));
	assign g2820 = (((!g2081) & (!g2124) & (!g2770) & (!g2811) & (!g2819) & (!g2100)) + ((!g2081) & (!g2124) & (!g2770) & (!g2811) & (!g2819) & (g2100)) + ((!g2081) & (!g2124) & (!g2770) & (g2811) & (!g2819) & (!g2100)) + ((!g2081) & (!g2124) & (!g2770) & (g2811) & (!g2819) & (g2100)) + ((!g2081) & (!g2124) & (g2770) & (!g2811) & (!g2819) & (!g2100)) + ((!g2081) & (!g2124) & (g2770) & (!g2811) & (g2819) & (!g2100)) + ((!g2081) & (!g2124) & (g2770) & (g2811) & (!g2819) & (!g2100)) + ((!g2081) & (!g2124) & (g2770) & (g2811) & (g2819) & (!g2100)) + ((!g2081) & (g2124) & (!g2770) & (!g2811) & (!g2819) & (!g2100)) + ((!g2081) & (g2124) & (!g2770) & (!g2811) & (g2819) & (!g2100)) + ((!g2081) & (g2124) & (g2770) & (!g2811) & (!g2819) & (!g2100)) + ((!g2081) & (g2124) & (g2770) & (!g2811) & (g2819) & (!g2100)) + ((!g2081) & (g2124) & (g2770) & (g2811) & (!g2819) & (!g2100)) + ((!g2081) & (g2124) & (g2770) & (g2811) & (g2819) & (!g2100)) + ((g2081) & (!g2124) & (!g2770) & (!g2811) & (!g2819) & (!g2100)) + ((g2081) & (!g2124) & (!g2770) & (!g2811) & (!g2819) & (g2100)) + ((g2081) & (!g2124) & (!g2770) & (g2811) & (!g2819) & (!g2100)) + ((g2081) & (!g2124) & (!g2770) & (g2811) & (!g2819) & (g2100)) + ((g2081) & (!g2124) & (g2770) & (!g2811) & (!g2819) & (!g2100)) + ((g2081) & (!g2124) & (g2770) & (!g2811) & (g2819) & (!g2100)) + ((g2081) & (!g2124) & (g2770) & (g2811) & (!g2819) & (!g2100)) + ((g2081) & (!g2124) & (g2770) & (g2811) & (g2819) & (!g2100)) + ((g2081) & (g2124) & (!g2770) & (!g2811) & (!g2819) & (!g2100)) + ((g2081) & (g2124) & (!g2770) & (!g2811) & (g2819) & (!g2100)) + ((g2081) & (g2124) & (!g2770) & (g2811) & (!g2819) & (g2100)) + ((g2081) & (g2124) & (!g2770) & (g2811) & (g2819) & (g2100)) + ((g2081) & (g2124) & (g2770) & (!g2811) & (!g2819) & (!g2100)) + ((g2081) & (g2124) & (g2770) & (!g2811) & (g2819) & (!g2100)) + ((g2081) & (g2124) & (g2770) & (g2811) & (!g2819) & (!g2100)) + ((g2081) & (g2124) & (g2770) & (g2811) & (g2819) & (!g2100)));
	assign g2821 = (((!g2820) & (!dmem_dat_ix30x) & (!g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2820) & (!dmem_dat_ix30x) & (!g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2820) & (!dmem_dat_ix30x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((!g2820) & (!dmem_dat_ix30x) & (g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2820) & (!dmem_dat_ix30x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((!g2820) & (!dmem_dat_ix30x) & (g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2820) & (!dmem_dat_ix30x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((!g2820) & (!dmem_dat_ix30x) & (g2783) & (g2784) & (g2785) & (g2786)) + ((!g2820) & (dmem_dat_ix30x) & (!g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2820) & (dmem_dat_ix30x) & (!g2783) & (!g2784) & (g2785) & (!g2786)) + ((!g2820) & (dmem_dat_ix30x) & (!g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2820) & (dmem_dat_ix30x) & (!g2783) & (g2784) & (g2785) & (!g2786)) + ((!g2820) & (dmem_dat_ix30x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((!g2820) & (dmem_dat_ix30x) & (g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2820) & (dmem_dat_ix30x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((!g2820) & (dmem_dat_ix30x) & (g2783) & (!g2784) & (g2785) & (!g2786)) + ((!g2820) & (dmem_dat_ix30x) & (g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2820) & (dmem_dat_ix30x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((!g2820) & (dmem_dat_ix30x) & (g2783) & (g2784) & (g2785) & (!g2786)) + ((!g2820) & (dmem_dat_ix30x) & (g2783) & (g2784) & (g2785) & (g2786)) + ((g2820) & (!dmem_dat_ix30x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((g2820) & (!dmem_dat_ix30x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((g2820) & (!dmem_dat_ix30x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((g2820) & (!dmem_dat_ix30x) & (g2783) & (g2784) & (g2785) & (g2786)) + ((g2820) & (dmem_dat_ix30x) & (!g2783) & (!g2784) & (g2785) & (!g2786)) + ((g2820) & (dmem_dat_ix30x) & (!g2783) & (g2784) & (g2785) & (!g2786)) + ((g2820) & (dmem_dat_ix30x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((g2820) & (dmem_dat_ix30x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((g2820) & (dmem_dat_ix30x) & (g2783) & (!g2784) & (g2785) & (!g2786)) + ((g2820) & (dmem_dat_ix30x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((g2820) & (dmem_dat_ix30x) & (g2783) & (g2784) & (g2785) & (!g2786)) + ((g2820) & (dmem_dat_ix30x) & (g2783) & (g2784) & (g2785) & (g2786)));
	assign g2822 = (((!sk[126]) & (!g1455) & (!g2788) & (!g1500) & (g1544)) + ((!sk[126]) & (!g1455) & (!g2788) & (g1500) & (g1544)) + ((!sk[126]) & (!g1455) & (g2788) & (!g1500) & (!g1544)) + ((!sk[126]) & (!g1455) & (g2788) & (!g1500) & (g1544)) + ((!sk[126]) & (!g1455) & (g2788) & (g1500) & (!g1544)) + ((!sk[126]) & (!g1455) & (g2788) & (g1500) & (g1544)) + ((!sk[126]) & (g1455) & (!g2788) & (!g1500) & (!g1544)) + ((!sk[126]) & (g1455) & (!g2788) & (!g1500) & (g1544)) + ((!sk[126]) & (g1455) & (!g2788) & (g1500) & (!g1544)) + ((!sk[126]) & (g1455) & (!g2788) & (g1500) & (g1544)) + ((!sk[126]) & (g1455) & (g2788) & (!g1500) & (!g1544)) + ((!sk[126]) & (g1455) & (g2788) & (!g1500) & (g1544)) + ((!sk[126]) & (g1455) & (g2788) & (g1500) & (!g1544)) + ((!sk[126]) & (g1455) & (g2788) & (g1500) & (g1544)) + ((sk[126]) & (!g1455) & (!g2788) & (!g1500) & (g1544)) + ((sk[126]) & (!g1455) & (!g2788) & (g1500) & (g1544)) + ((sk[126]) & (!g1455) & (g2788) & (!g1500) & (g1544)) + ((sk[126]) & (!g1455) & (g2788) & (g1500) & (g1544)) + ((sk[126]) & (g1455) & (!g2788) & (!g1500) & (g1544)) + ((sk[126]) & (g1455) & (!g2788) & (g1500) & (g1544)) + ((sk[126]) & (g1455) & (g2788) & (!g1500) & (g1544)) + ((sk[126]) & (g1455) & (g2788) & (g1500) & (!g1544)));
	assign g2823 = (((!g107) & (!g1410) & (!g2765) & (g1455) & (!sk[127]) & (!g1500)) + ((!g107) & (!g1410) & (!g2765) & (g1455) & (!sk[127]) & (g1500)) + ((!g107) & (!g1410) & (g2765) & (!g1455) & (!sk[127]) & (!g1500)) + ((!g107) & (!g1410) & (g2765) & (!g1455) & (!sk[127]) & (g1500)) + ((!g107) & (!g1410) & (g2765) & (g1455) & (!sk[127]) & (!g1500)) + ((!g107) & (!g1410) & (g2765) & (g1455) & (!sk[127]) & (g1500)) + ((!g107) & (g1410) & (!g2765) & (g1455) & (!sk[127]) & (!g1500)) + ((!g107) & (g1410) & (!g2765) & (g1455) & (!sk[127]) & (g1500)) + ((!g107) & (g1410) & (g2765) & (!g1455) & (!sk[127]) & (!g1500)) + ((!g107) & (g1410) & (g2765) & (!g1455) & (!sk[127]) & (g1500)) + ((!g107) & (g1410) & (g2765) & (g1455) & (!sk[127]) & (!g1500)) + ((!g107) & (g1410) & (g2765) & (g1455) & (!sk[127]) & (g1500)) + ((!g107) & (g1410) & (g2765) & (g1455) & (sk[127]) & (g1500)) + ((g107) & (!g1410) & (!g2765) & (!g1455) & (!sk[127]) & (!g1500)) + ((g107) & (!g1410) & (!g2765) & (!g1455) & (!sk[127]) & (g1500)) + ((g107) & (!g1410) & (!g2765) & (!g1455) & (sk[127]) & (g1500)) + ((g107) & (!g1410) & (!g2765) & (g1455) & (!sk[127]) & (!g1500)) + ((g107) & (!g1410) & (!g2765) & (g1455) & (!sk[127]) & (g1500)) + ((g107) & (!g1410) & (!g2765) & (g1455) & (sk[127]) & (!g1500)) + ((g107) & (!g1410) & (!g2765) & (g1455) & (sk[127]) & (g1500)) + ((g107) & (!g1410) & (g2765) & (!g1455) & (!sk[127]) & (!g1500)) + ((g107) & (!g1410) & (g2765) & (!g1455) & (!sk[127]) & (g1500)) + ((g107) & (!g1410) & (g2765) & (!g1455) & (sk[127]) & (!g1500)) + ((g107) & (!g1410) & (g2765) & (!g1455) & (sk[127]) & (g1500)) + ((g107) & (!g1410) & (g2765) & (g1455) & (!sk[127]) & (!g1500)) + ((g107) & (!g1410) & (g2765) & (g1455) & (!sk[127]) & (g1500)) + ((g107) & (!g1410) & (g2765) & (g1455) & (sk[127]) & (!g1500)) + ((g107) & (!g1410) & (g2765) & (g1455) & (sk[127]) & (g1500)) + ((g107) & (g1410) & (!g2765) & (!g1455) & (!sk[127]) & (!g1500)) + ((g107) & (g1410) & (!g2765) & (!g1455) & (!sk[127]) & (g1500)) + ((g107) & (g1410) & (!g2765) & (!g1455) & (sk[127]) & (!g1500)) + ((g107) & (g1410) & (!g2765) & (!g1455) & (sk[127]) & (g1500)) + ((g107) & (g1410) & (!g2765) & (g1455) & (!sk[127]) & (!g1500)) + ((g107) & (g1410) & (!g2765) & (g1455) & (!sk[127]) & (g1500)) + ((g107) & (g1410) & (!g2765) & (g1455) & (sk[127]) & (!g1500)) + ((g107) & (g1410) & (!g2765) & (g1455) & (sk[127]) & (g1500)) + ((g107) & (g1410) & (g2765) & (!g1455) & (!sk[127]) & (!g1500)) + ((g107) & (g1410) & (g2765) & (!g1455) & (!sk[127]) & (g1500)) + ((g107) & (g1410) & (g2765) & (!g1455) & (sk[127]) & (!g1500)) + ((g107) & (g1410) & (g2765) & (!g1455) & (sk[127]) & (g1500)) + ((g107) & (g1410) & (g2765) & (g1455) & (!sk[127]) & (!g1500)) + ((g107) & (g1410) & (g2765) & (g1455) & (!sk[127]) & (g1500)) + ((g107) & (g1410) & (g2765) & (g1455) & (sk[127]) & (!g1500)) + ((g107) & (g1410) & (g2765) & (g1455) & (sk[127]) & (g1500)));
	assign g5054 = (((!g2921) & (!sk[0]) & (g3111) & (!g2824)) + ((!g2921) & (!sk[0]) & (g3111) & (g2824)) + ((!g2921) & (sk[0]) & (!g3111) & (g2824)) + ((!g2921) & (sk[0]) & (g3111) & (g2824)) + ((g2921) & (!sk[0]) & (!g3111) & (!g2824)) + ((g2921) & (!sk[0]) & (!g3111) & (g2824)) + ((g2921) & (!sk[0]) & (g3111) & (!g2824)) + ((g2921) & (!sk[0]) & (g3111) & (g2824)) + ((g2921) & (sk[0]) & (g3111) & (!g2824)) + ((g2921) & (sk[0]) & (g3111) & (g2824)));
	assign g2825 = (((!g2329) & (!g2029) & (!g2408) & (g2822) & (!sk[1]) & (!g3252)) + ((!g2329) & (!g2029) & (!g2408) & (g2822) & (!sk[1]) & (g3252)) + ((!g2329) & (!g2029) & (g2408) & (!g2822) & (!sk[1]) & (!g3252)) + ((!g2329) & (!g2029) & (g2408) & (!g2822) & (!sk[1]) & (g3252)) + ((!g2329) & (!g2029) & (g2408) & (g2822) & (!sk[1]) & (!g3252)) + ((!g2329) & (!g2029) & (g2408) & (g2822) & (!sk[1]) & (g3252)) + ((!g2329) & (g2029) & (!g2408) & (g2822) & (!sk[1]) & (!g3252)) + ((!g2329) & (g2029) & (!g2408) & (g2822) & (!sk[1]) & (g3252)) + ((!g2329) & (g2029) & (g2408) & (!g2822) & (!sk[1]) & (!g3252)) + ((!g2329) & (g2029) & (g2408) & (!g2822) & (!sk[1]) & (g3252)) + ((!g2329) & (g2029) & (g2408) & (g2822) & (!sk[1]) & (!g3252)) + ((!g2329) & (g2029) & (g2408) & (g2822) & (!sk[1]) & (g3252)) + ((g2329) & (!g2029) & (!g2408) & (!g2822) & (!sk[1]) & (!g3252)) + ((g2329) & (!g2029) & (!g2408) & (!g2822) & (!sk[1]) & (g3252)) + ((g2329) & (!g2029) & (!g2408) & (g2822) & (!sk[1]) & (!g3252)) + ((g2329) & (!g2029) & (!g2408) & (g2822) & (!sk[1]) & (g3252)) + ((g2329) & (!g2029) & (g2408) & (!g2822) & (!sk[1]) & (!g3252)) + ((g2329) & (!g2029) & (g2408) & (!g2822) & (!sk[1]) & (g3252)) + ((g2329) & (!g2029) & (g2408) & (!g2822) & (sk[1]) & (g3252)) + ((g2329) & (!g2029) & (g2408) & (g2822) & (!sk[1]) & (!g3252)) + ((g2329) & (!g2029) & (g2408) & (g2822) & (!sk[1]) & (g3252)) + ((g2329) & (!g2029) & (g2408) & (g2822) & (sk[1]) & (g3252)) + ((g2329) & (g2029) & (!g2408) & (!g2822) & (!sk[1]) & (!g3252)) + ((g2329) & (g2029) & (!g2408) & (!g2822) & (!sk[1]) & (g3252)) + ((g2329) & (g2029) & (!g2408) & (g2822) & (!sk[1]) & (!g3252)) + ((g2329) & (g2029) & (!g2408) & (g2822) & (!sk[1]) & (g3252)) + ((g2329) & (g2029) & (g2408) & (!g2822) & (!sk[1]) & (!g3252)) + ((g2329) & (g2029) & (g2408) & (!g2822) & (!sk[1]) & (g3252)) + ((g2329) & (g2029) & (g2408) & (g2822) & (!sk[1]) & (!g3252)) + ((g2329) & (g2029) & (g2408) & (g2822) & (!sk[1]) & (g3252)) + ((g2329) & (g2029) & (g2408) & (g2822) & (sk[1]) & (!g3252)) + ((g2329) & (g2029) & (g2408) & (g2822) & (sk[1]) & (g3252)));
	assign g2826 = (((!g1455) & (!g2788) & (!sk[2]) & (!g1500) & (g1544) & (!g1547)) + ((!g1455) & (!g2788) & (!sk[2]) & (!g1500) & (g1544) & (g1547)) + ((!g1455) & (!g2788) & (!sk[2]) & (g1500) & (!g1544) & (!g1547)) + ((!g1455) & (!g2788) & (!sk[2]) & (g1500) & (!g1544) & (g1547)) + ((!g1455) & (!g2788) & (!sk[2]) & (g1500) & (g1544) & (!g1547)) + ((!g1455) & (!g2788) & (!sk[2]) & (g1500) & (g1544) & (g1547)) + ((!g1455) & (!g2788) & (sk[2]) & (!g1500) & (!g1544) & (g1547)) + ((!g1455) & (!g2788) & (sk[2]) & (!g1500) & (g1544) & (g1547)) + ((!g1455) & (!g2788) & (sk[2]) & (g1500) & (!g1544) & (g1547)) + ((!g1455) & (!g2788) & (sk[2]) & (g1500) & (g1544) & (g1547)) + ((!g1455) & (g2788) & (!sk[2]) & (!g1500) & (g1544) & (!g1547)) + ((!g1455) & (g2788) & (!sk[2]) & (!g1500) & (g1544) & (g1547)) + ((!g1455) & (g2788) & (!sk[2]) & (g1500) & (!g1544) & (!g1547)) + ((!g1455) & (g2788) & (!sk[2]) & (g1500) & (!g1544) & (g1547)) + ((!g1455) & (g2788) & (!sk[2]) & (g1500) & (g1544) & (!g1547)) + ((!g1455) & (g2788) & (!sk[2]) & (g1500) & (g1544) & (g1547)) + ((!g1455) & (g2788) & (sk[2]) & (!g1500) & (!g1544) & (g1547)) + ((!g1455) & (g2788) & (sk[2]) & (!g1500) & (g1544) & (g1547)) + ((!g1455) & (g2788) & (sk[2]) & (g1500) & (!g1544) & (g1547)) + ((!g1455) & (g2788) & (sk[2]) & (g1500) & (g1544) & (g1547)) + ((g1455) & (!g2788) & (!sk[2]) & (!g1500) & (!g1544) & (!g1547)) + ((g1455) & (!g2788) & (!sk[2]) & (!g1500) & (!g1544) & (g1547)) + ((g1455) & (!g2788) & (!sk[2]) & (!g1500) & (g1544) & (!g1547)) + ((g1455) & (!g2788) & (!sk[2]) & (!g1500) & (g1544) & (g1547)) + ((g1455) & (!g2788) & (!sk[2]) & (g1500) & (!g1544) & (!g1547)) + ((g1455) & (!g2788) & (!sk[2]) & (g1500) & (!g1544) & (g1547)) + ((g1455) & (!g2788) & (!sk[2]) & (g1500) & (g1544) & (!g1547)) + ((g1455) & (!g2788) & (!sk[2]) & (g1500) & (g1544) & (g1547)) + ((g1455) & (!g2788) & (sk[2]) & (!g1500) & (!g1544) & (g1547)) + ((g1455) & (!g2788) & (sk[2]) & (!g1500) & (g1544) & (g1547)) + ((g1455) & (!g2788) & (sk[2]) & (g1500) & (!g1544) & (g1547)) + ((g1455) & (!g2788) & (sk[2]) & (g1500) & (g1544) & (g1547)) + ((g1455) & (g2788) & (!sk[2]) & (!g1500) & (!g1544) & (!g1547)) + ((g1455) & (g2788) & (!sk[2]) & (!g1500) & (!g1544) & (g1547)) + ((g1455) & (g2788) & (!sk[2]) & (!g1500) & (g1544) & (!g1547)) + ((g1455) & (g2788) & (!sk[2]) & (!g1500) & (g1544) & (g1547)) + ((g1455) & (g2788) & (!sk[2]) & (g1500) & (!g1544) & (!g1547)) + ((g1455) & (g2788) & (!sk[2]) & (g1500) & (!g1544) & (g1547)) + ((g1455) & (g2788) & (!sk[2]) & (g1500) & (g1544) & (!g1547)) + ((g1455) & (g2788) & (!sk[2]) & (g1500) & (g1544) & (g1547)) + ((g1455) & (g2788) & (sk[2]) & (!g1500) & (!g1544) & (g1547)) + ((g1455) & (g2788) & (sk[2]) & (!g1500) & (g1544) & (g1547)) + ((g1455) & (g2788) & (sk[2]) & (g1500) & (!g1544) & (g1547)) + ((g1455) & (g2788) & (sk[2]) & (g1500) & (g1544) & (!g1547)));
	assign g5055 = (((!g2921) & (!g3112) & (sk[3]) & (g2827)) + ((!g2921) & (g3112) & (!sk[3]) & (!g2827)) + ((!g2921) & (g3112) & (!sk[3]) & (g2827)) + ((!g2921) & (g3112) & (sk[3]) & (g2827)) + ((g2921) & (!g3112) & (!sk[3]) & (!g2827)) + ((g2921) & (!g3112) & (!sk[3]) & (g2827)) + ((g2921) & (g3112) & (!sk[3]) & (!g2827)) + ((g2921) & (g3112) & (!sk[3]) & (g2827)) + ((g2921) & (g3112) & (sk[3]) & (!g2827)) + ((g2921) & (g3112) & (sk[3]) & (g2827)));
	assign g2828 = (((!g2007) & (!sk[4]) & (!g2033) & (!g2034) & (g2827)) + ((!g2007) & (!sk[4]) & (!g2033) & (g2034) & (g2827)) + ((!g2007) & (!sk[4]) & (g2033) & (!g2034) & (!g2827)) + ((!g2007) & (!sk[4]) & (g2033) & (!g2034) & (g2827)) + ((!g2007) & (!sk[4]) & (g2033) & (g2034) & (!g2827)) + ((!g2007) & (!sk[4]) & (g2033) & (g2034) & (g2827)) + ((!g2007) & (sk[4]) & (!g2033) & (!g2034) & (g2827)) + ((g2007) & (!sk[4]) & (!g2033) & (!g2034) & (!g2827)) + ((g2007) & (!sk[4]) & (!g2033) & (!g2034) & (g2827)) + ((g2007) & (!sk[4]) & (!g2033) & (g2034) & (!g2827)) + ((g2007) & (!sk[4]) & (!g2033) & (g2034) & (g2827)) + ((g2007) & (!sk[4]) & (g2033) & (!g2034) & (!g2827)) + ((g2007) & (!sk[4]) & (g2033) & (!g2034) & (g2827)) + ((g2007) & (!sk[4]) & (g2033) & (g2034) & (!g2827)) + ((g2007) & (!sk[4]) & (g2033) & (g2034) & (g2827)) + ((g2007) & (sk[4]) & (!g2033) & (!g2034) & (g2827)) + ((g2007) & (sk[4]) & (!g2033) & (g2034) & (!g2827)) + ((g2007) & (sk[4]) & (!g2033) & (g2034) & (g2827)));
	assign g2829 = (((!g107) & (!g2585) & (!g1544) & (!g2823) & (!g1547) & (!g2828)) + ((!g107) & (!g2585) & (!g1544) & (!g2823) & (g1547) & (!g2828)) + ((!g107) & (!g2585) & (!g1544) & (g2823) & (!g1547) & (!g2828)) + ((!g107) & (!g2585) & (!g1544) & (g2823) & (g1547) & (!g2828)) + ((!g107) & (!g2585) & (g1544) & (!g2823) & (!g1547) & (!g2828)) + ((!g107) & (!g2585) & (g1544) & (!g2823) & (g1547) & (!g2828)) + ((!g107) & (!g2585) & (g1544) & (g2823) & (!g1547) & (!g2828)) + ((!g107) & (!g2585) & (g1544) & (g2823) & (g1547) & (!g2828)) + ((!g107) & (g2585) & (!g1544) & (!g2823) & (!g1547) & (!g2828)) + ((!g107) & (g2585) & (!g1544) & (g2823) & (!g1547) & (!g2828)) + ((!g107) & (g2585) & (g1544) & (!g2823) & (!g1547) & (!g2828)) + ((!g107) & (g2585) & (g1544) & (g2823) & (g1547) & (!g2828)) + ((g107) & (!g2585) & (!g1544) & (!g2823) & (!g1547) & (!g2828)) + ((g107) & (!g2585) & (!g1544) & (!g2823) & (g1547) & (!g2828)) + ((g107) & (!g2585) & (!g1544) & (g2823) & (!g1547) & (!g2828)) + ((g107) & (!g2585) & (!g1544) & (g2823) & (g1547) & (!g2828)) + ((g107) & (!g2585) & (g1544) & (!g2823) & (!g1547) & (!g2828)) + ((g107) & (!g2585) & (g1544) & (!g2823) & (g1547) & (!g2828)) + ((g107) & (!g2585) & (g1544) & (g2823) & (!g1547) & (!g2828)) + ((g107) & (!g2585) & (g1544) & (g2823) & (g1547) & (!g2828)) + ((g107) & (g2585) & (!g1544) & (!g2823) & (g1547) & (!g2828)) + ((g107) & (g2585) & (!g1544) & (g2823) & (!g1547) & (!g2828)) + ((g107) & (g2585) & (g1544) & (!g2823) & (!g1547) & (!g2828)) + ((g107) & (g2585) & (g1544) & (g2823) & (!g1547) & (!g2828)));
	assign g2830 = (((!g2329) & (!sk[6]) & (!g2029) & (!g2408) & (g2826) & (!g2829)) + ((!g2329) & (!sk[6]) & (!g2029) & (!g2408) & (g2826) & (g2829)) + ((!g2329) & (!sk[6]) & (!g2029) & (g2408) & (!g2826) & (!g2829)) + ((!g2329) & (!sk[6]) & (!g2029) & (g2408) & (!g2826) & (g2829)) + ((!g2329) & (!sk[6]) & (!g2029) & (g2408) & (g2826) & (!g2829)) + ((!g2329) & (!sk[6]) & (!g2029) & (g2408) & (g2826) & (g2829)) + ((!g2329) & (!sk[6]) & (g2029) & (!g2408) & (g2826) & (!g2829)) + ((!g2329) & (!sk[6]) & (g2029) & (!g2408) & (g2826) & (g2829)) + ((!g2329) & (!sk[6]) & (g2029) & (g2408) & (!g2826) & (!g2829)) + ((!g2329) & (!sk[6]) & (g2029) & (g2408) & (!g2826) & (g2829)) + ((!g2329) & (!sk[6]) & (g2029) & (g2408) & (g2826) & (!g2829)) + ((!g2329) & (!sk[6]) & (g2029) & (g2408) & (g2826) & (g2829)) + ((g2329) & (!sk[6]) & (!g2029) & (!g2408) & (!g2826) & (!g2829)) + ((g2329) & (!sk[6]) & (!g2029) & (!g2408) & (!g2826) & (g2829)) + ((g2329) & (!sk[6]) & (!g2029) & (!g2408) & (g2826) & (!g2829)) + ((g2329) & (!sk[6]) & (!g2029) & (!g2408) & (g2826) & (g2829)) + ((g2329) & (!sk[6]) & (!g2029) & (g2408) & (!g2826) & (!g2829)) + ((g2329) & (!sk[6]) & (!g2029) & (g2408) & (!g2826) & (g2829)) + ((g2329) & (!sk[6]) & (!g2029) & (g2408) & (g2826) & (!g2829)) + ((g2329) & (!sk[6]) & (!g2029) & (g2408) & (g2826) & (g2829)) + ((g2329) & (!sk[6]) & (g2029) & (!g2408) & (!g2826) & (!g2829)) + ((g2329) & (!sk[6]) & (g2029) & (!g2408) & (!g2826) & (g2829)) + ((g2329) & (!sk[6]) & (g2029) & (!g2408) & (g2826) & (!g2829)) + ((g2329) & (!sk[6]) & (g2029) & (!g2408) & (g2826) & (g2829)) + ((g2329) & (!sk[6]) & (g2029) & (g2408) & (!g2826) & (!g2829)) + ((g2329) & (!sk[6]) & (g2029) & (g2408) & (!g2826) & (g2829)) + ((g2329) & (!sk[6]) & (g2029) & (g2408) & (g2826) & (!g2829)) + ((g2329) & (!sk[6]) & (g2029) & (g2408) & (g2826) & (g2829)) + ((g2329) & (sk[6]) & (!g2029) & (g2408) & (!g2826) & (!g2829)) + ((g2329) & (sk[6]) & (!g2029) & (g2408) & (g2826) & (!g2829)) + ((g2329) & (sk[6]) & (g2029) & (g2408) & (g2826) & (!g2829)) + ((g2329) & (sk[6]) & (g2029) & (g2408) & (g2826) & (g2829)));
	assign g2832 = (((!g2098) & (!g2099) & (!g2771) & (g2772) & (!sk[7]) & (!g2794)) + ((!g2098) & (!g2099) & (!g2771) & (g2772) & (!sk[7]) & (g2794)) + ((!g2098) & (!g2099) & (g2771) & (!g2772) & (!sk[7]) & (!g2794)) + ((!g2098) & (!g2099) & (g2771) & (!g2772) & (!sk[7]) & (g2794)) + ((!g2098) & (!g2099) & (g2771) & (g2772) & (!sk[7]) & (!g2794)) + ((!g2098) & (!g2099) & (g2771) & (g2772) & (!sk[7]) & (g2794)) + ((!g2098) & (!g2099) & (g2771) & (g2772) & (sk[7]) & (g2794)) + ((!g2098) & (g2099) & (!g2771) & (!g2772) & (sk[7]) & (g2794)) + ((!g2098) & (g2099) & (!g2771) & (g2772) & (!sk[7]) & (!g2794)) + ((!g2098) & (g2099) & (!g2771) & (g2772) & (!sk[7]) & (g2794)) + ((!g2098) & (g2099) & (!g2771) & (g2772) & (sk[7]) & (g2794)) + ((!g2098) & (g2099) & (g2771) & (!g2772) & (!sk[7]) & (!g2794)) + ((!g2098) & (g2099) & (g2771) & (!g2772) & (!sk[7]) & (g2794)) + ((!g2098) & (g2099) & (g2771) & (!g2772) & (sk[7]) & (g2794)) + ((!g2098) & (g2099) & (g2771) & (g2772) & (!sk[7]) & (!g2794)) + ((!g2098) & (g2099) & (g2771) & (g2772) & (!sk[7]) & (g2794)) + ((!g2098) & (g2099) & (g2771) & (g2772) & (sk[7]) & (!g2794)) + ((!g2098) & (g2099) & (g2771) & (g2772) & (sk[7]) & (g2794)) + ((g2098) & (!g2099) & (!g2771) & (!g2772) & (!sk[7]) & (!g2794)) + ((g2098) & (!g2099) & (!g2771) & (!g2772) & (!sk[7]) & (g2794)) + ((g2098) & (!g2099) & (!g2771) & (g2772) & (!sk[7]) & (!g2794)) + ((g2098) & (!g2099) & (!g2771) & (g2772) & (!sk[7]) & (g2794)) + ((g2098) & (!g2099) & (!g2771) & (g2772) & (sk[7]) & (g2794)) + ((g2098) & (!g2099) & (g2771) & (!g2772) & (!sk[7]) & (!g2794)) + ((g2098) & (!g2099) & (g2771) & (!g2772) & (!sk[7]) & (g2794)) + ((g2098) & (!g2099) & (g2771) & (!g2772) & (sk[7]) & (g2794)) + ((g2098) & (!g2099) & (g2771) & (g2772) & (!sk[7]) & (!g2794)) + ((g2098) & (!g2099) & (g2771) & (g2772) & (!sk[7]) & (g2794)) + ((g2098) & (!g2099) & (g2771) & (g2772) & (sk[7]) & (g2794)) + ((g2098) & (g2099) & (!g2771) & (!g2772) & (!sk[7]) & (!g2794)) + ((g2098) & (g2099) & (!g2771) & (!g2772) & (!sk[7]) & (g2794)) + ((g2098) & (g2099) & (!g2771) & (!g2772) & (sk[7]) & (g2794)) + ((g2098) & (g2099) & (!g2771) & (g2772) & (!sk[7]) & (!g2794)) + ((g2098) & (g2099) & (!g2771) & (g2772) & (!sk[7]) & (g2794)) + ((g2098) & (g2099) & (!g2771) & (g2772) & (sk[7]) & (!g2794)) + ((g2098) & (g2099) & (!g2771) & (g2772) & (sk[7]) & (g2794)) + ((g2098) & (g2099) & (g2771) & (!g2772) & (!sk[7]) & (!g2794)) + ((g2098) & (g2099) & (g2771) & (!g2772) & (!sk[7]) & (g2794)) + ((g2098) & (g2099) & (g2771) & (!g2772) & (sk[7]) & (!g2794)) + ((g2098) & (g2099) & (g2771) & (!g2772) & (sk[7]) & (g2794)) + ((g2098) & (g2099) & (g2771) & (g2772) & (!sk[7]) & (!g2794)) + ((g2098) & (g2099) & (g2771) & (g2772) & (!sk[7]) & (g2794)) + ((g2098) & (g2099) & (g2771) & (g2772) & (sk[7]) & (!g2794)) + ((g2098) & (g2099) & (g2771) & (g2772) & (sk[7]) & (g2794)));
	assign g2833 = (((!g2101) & (!sk[8]) & (g2831)) + ((!g2101) & (sk[8]) & (g2831)) + ((g2101) & (!sk[8]) & (g2831)) + ((g2101) & (sk[8]) & (!g2831)));
	assign g2834 = (((!g2100) & (!g2795) & (!g2796) & (!g2811) & (!g2832) & (g2833)) + ((!g2100) & (!g2795) & (!g2796) & (!g2811) & (g2832) & (g2833)) + ((!g2100) & (!g2795) & (!g2796) & (g2811) & (!g2832) & (g2833)) + ((!g2100) & (!g2795) & (!g2796) & (g2811) & (g2832) & (!g2833)) + ((!g2100) & (!g2795) & (g2796) & (!g2811) & (!g2832) & (g2833)) + ((!g2100) & (!g2795) & (g2796) & (!g2811) & (g2832) & (g2833)) + ((!g2100) & (!g2795) & (g2796) & (g2811) & (!g2832) & (g2833)) + ((!g2100) & (!g2795) & (g2796) & (g2811) & (g2832) & (!g2833)) + ((!g2100) & (g2795) & (!g2796) & (!g2811) & (!g2832) & (g2833)) + ((!g2100) & (g2795) & (!g2796) & (!g2811) & (g2832) & (g2833)) + ((!g2100) & (g2795) & (!g2796) & (g2811) & (!g2832) & (g2833)) + ((!g2100) & (g2795) & (!g2796) & (g2811) & (g2832) & (!g2833)) + ((!g2100) & (g2795) & (g2796) & (!g2811) & (!g2832) & (g2833)) + ((!g2100) & (g2795) & (g2796) & (!g2811) & (g2832) & (!g2833)) + ((!g2100) & (g2795) & (g2796) & (g2811) & (!g2832) & (!g2833)) + ((!g2100) & (g2795) & (g2796) & (g2811) & (g2832) & (!g2833)) + ((g2100) & (!g2795) & (!g2796) & (!g2811) & (!g2832) & (g2833)) + ((g2100) & (!g2795) & (!g2796) & (!g2811) & (g2832) & (!g2833)) + ((g2100) & (!g2795) & (!g2796) & (g2811) & (!g2832) & (!g2833)) + ((g2100) & (!g2795) & (!g2796) & (g2811) & (g2832) & (!g2833)) + ((g2100) & (!g2795) & (g2796) & (!g2811) & (!g2832) & (g2833)) + ((g2100) & (!g2795) & (g2796) & (!g2811) & (g2832) & (!g2833)) + ((g2100) & (!g2795) & (g2796) & (g2811) & (!g2832) & (!g2833)) + ((g2100) & (!g2795) & (g2796) & (g2811) & (g2832) & (!g2833)) + ((g2100) & (g2795) & (!g2796) & (!g2811) & (!g2832) & (g2833)) + ((g2100) & (g2795) & (!g2796) & (!g2811) & (g2832) & (!g2833)) + ((g2100) & (g2795) & (!g2796) & (g2811) & (!g2832) & (!g2833)) + ((g2100) & (g2795) & (!g2796) & (g2811) & (g2832) & (!g2833)) + ((g2100) & (g2795) & (g2796) & (!g2811) & (!g2832) & (!g2833)) + ((g2100) & (g2795) & (g2796) & (!g2811) & (g2832) & (!g2833)) + ((g2100) & (g2795) & (g2796) & (g2811) & (!g2832) & (!g2833)) + ((g2100) & (g2795) & (g2796) & (g2811) & (g2832) & (g2833)));
	assign g2835 = (((!g2831) & (!g2101) & (!sk[10]) & (!g2811) & (g2100)) + ((!g2831) & (!g2101) & (!sk[10]) & (g2811) & (g2100)) + ((!g2831) & (!g2101) & (sk[10]) & (!g2811) & (!g2100)) + ((!g2831) & (!g2101) & (sk[10]) & (g2811) & (!g2100)) + ((!g2831) & (!g2101) & (sk[10]) & (g2811) & (g2100)) + ((!g2831) & (g2101) & (!sk[10]) & (!g2811) & (!g2100)) + ((!g2831) & (g2101) & (!sk[10]) & (!g2811) & (g2100)) + ((!g2831) & (g2101) & (!sk[10]) & (g2811) & (!g2100)) + ((!g2831) & (g2101) & (!sk[10]) & (g2811) & (g2100)) + ((!g2831) & (g2101) & (sk[10]) & (!g2811) & (g2100)) + ((g2831) & (!g2101) & (!sk[10]) & (!g2811) & (!g2100)) + ((g2831) & (!g2101) & (!sk[10]) & (!g2811) & (g2100)) + ((g2831) & (!g2101) & (!sk[10]) & (g2811) & (!g2100)) + ((g2831) & (!g2101) & (!sk[10]) & (g2811) & (g2100)) + ((g2831) & (!g2101) & (sk[10]) & (!g2811) & (g2100)) + ((g2831) & (g2101) & (!sk[10]) & (!g2811) & (!g2100)) + ((g2831) & (g2101) & (!sk[10]) & (!g2811) & (g2100)) + ((g2831) & (g2101) & (!sk[10]) & (g2811) & (!g2100)) + ((g2831) & (g2101) & (!sk[10]) & (g2811) & (g2100)) + ((g2831) & (g2101) & (sk[10]) & (!g2811) & (!g2100)) + ((g2831) & (g2101) & (sk[10]) & (g2811) & (!g2100)) + ((g2831) & (g2101) & (sk[10]) & (g2811) & (g2100)));
	assign g2836 = (((!g2797) & (!g2798) & (!g2799) & (!g2814) & (!g2815) & (g2835)) + ((!g2797) & (!g2798) & (!g2799) & (!g2814) & (g2815) & (g2835)) + ((!g2797) & (!g2798) & (!g2799) & (g2814) & (!g2815) & (g2835)) + ((!g2797) & (!g2798) & (!g2799) & (g2814) & (g2815) & (!g2835)) + ((!g2797) & (!g2798) & (g2799) & (!g2814) & (!g2815) & (g2835)) + ((!g2797) & (!g2798) & (g2799) & (!g2814) & (g2815) & (!g2835)) + ((!g2797) & (!g2798) & (g2799) & (g2814) & (!g2815) & (!g2835)) + ((!g2797) & (!g2798) & (g2799) & (g2814) & (g2815) & (!g2835)) + ((!g2797) & (g2798) & (!g2799) & (!g2814) & (!g2815) & (g2835)) + ((!g2797) & (g2798) & (!g2799) & (!g2814) & (g2815) & (!g2835)) + ((!g2797) & (g2798) & (!g2799) & (g2814) & (!g2815) & (!g2835)) + ((!g2797) & (g2798) & (!g2799) & (g2814) & (g2815) & (!g2835)) + ((!g2797) & (g2798) & (g2799) & (!g2814) & (!g2815) & (g2835)) + ((!g2797) & (g2798) & (g2799) & (!g2814) & (g2815) & (!g2835)) + ((!g2797) & (g2798) & (g2799) & (g2814) & (!g2815) & (!g2835)) + ((!g2797) & (g2798) & (g2799) & (g2814) & (g2815) & (!g2835)) + ((g2797) & (!g2798) & (!g2799) & (!g2814) & (!g2815) & (g2835)) + ((g2797) & (!g2798) & (!g2799) & (!g2814) & (g2815) & (g2835)) + ((g2797) & (!g2798) & (!g2799) & (g2814) & (!g2815) & (g2835)) + ((g2797) & (!g2798) & (!g2799) & (g2814) & (g2815) & (!g2835)) + ((g2797) & (!g2798) & (g2799) & (!g2814) & (!g2815) & (g2835)) + ((g2797) & (!g2798) & (g2799) & (!g2814) & (g2815) & (g2835)) + ((g2797) & (!g2798) & (g2799) & (g2814) & (!g2815) & (g2835)) + ((g2797) & (!g2798) & (g2799) & (g2814) & (g2815) & (!g2835)) + ((g2797) & (g2798) & (!g2799) & (!g2814) & (!g2815) & (g2835)) + ((g2797) & (g2798) & (!g2799) & (!g2814) & (g2815) & (g2835)) + ((g2797) & (g2798) & (!g2799) & (g2814) & (!g2815) & (g2835)) + ((g2797) & (g2798) & (!g2799) & (g2814) & (g2815) & (!g2835)) + ((g2797) & (g2798) & (g2799) & (!g2814) & (!g2815) & (g2835)) + ((g2797) & (g2798) & (g2799) & (!g2814) & (g2815) & (!g2835)) + ((g2797) & (g2798) & (g2799) & (g2814) & (!g2815) & (!g2835)) + ((g2797) & (g2798) & (g2799) & (g2814) & (g2815) & (!g2835)));
	assign g2837 = (((!sk[12]) & (!g2101) & (g2831)) + ((!sk[12]) & (g2101) & (g2831)) + ((sk[12]) & (g2101) & (g2831)));
	assign g2838 = (((!g2760) & (!g2100) & (!g2099) & (g2098) & (g2196) & (g2197)) + ((!g2760) & (!g2100) & (g2099) & (!g2098) & (!g2196) & (g2197)) + ((!g2760) & (!g2100) & (g2099) & (g2098) & (!g2196) & (g2197)) + ((!g2760) & (!g2100) & (g2099) & (g2098) & (g2196) & (g2197)) + ((!g2760) & (g2100) & (!g2099) & (!g2098) & (g2196) & (!g2197)) + ((!g2760) & (g2100) & (!g2099) & (g2098) & (g2196) & (!g2197)) + ((!g2760) & (g2100) & (!g2099) & (g2098) & (g2196) & (g2197)) + ((!g2760) & (g2100) & (g2099) & (!g2098) & (!g2196) & (g2197)) + ((!g2760) & (g2100) & (g2099) & (!g2098) & (g2196) & (!g2197)) + ((!g2760) & (g2100) & (g2099) & (g2098) & (!g2196) & (g2197)) + ((!g2760) & (g2100) & (g2099) & (g2098) & (g2196) & (!g2197)) + ((!g2760) & (g2100) & (g2099) & (g2098) & (g2196) & (g2197)) + ((g2760) & (!g2100) & (!g2099) & (!g2098) & (!g2196) & (!g2197)) + ((g2760) & (!g2100) & (!g2099) & (g2098) & (!g2196) & (!g2197)) + ((g2760) & (!g2100) & (!g2099) & (g2098) & (g2196) & (g2197)) + ((g2760) & (!g2100) & (g2099) & (!g2098) & (!g2196) & (!g2197)) + ((g2760) & (!g2100) & (g2099) & (!g2098) & (!g2196) & (g2197)) + ((g2760) & (!g2100) & (g2099) & (g2098) & (!g2196) & (!g2197)) + ((g2760) & (!g2100) & (g2099) & (g2098) & (!g2196) & (g2197)) + ((g2760) & (!g2100) & (g2099) & (g2098) & (g2196) & (g2197)) + ((g2760) & (g2100) & (!g2099) & (!g2098) & (!g2196) & (!g2197)) + ((g2760) & (g2100) & (!g2099) & (!g2098) & (g2196) & (!g2197)) + ((g2760) & (g2100) & (!g2099) & (g2098) & (!g2196) & (!g2197)) + ((g2760) & (g2100) & (!g2099) & (g2098) & (g2196) & (!g2197)) + ((g2760) & (g2100) & (!g2099) & (g2098) & (g2196) & (g2197)) + ((g2760) & (g2100) & (g2099) & (!g2098) & (!g2196) & (!g2197)) + ((g2760) & (g2100) & (g2099) & (!g2098) & (!g2196) & (g2197)) + ((g2760) & (g2100) & (g2099) & (!g2098) & (g2196) & (!g2197)) + ((g2760) & (g2100) & (g2099) & (g2098) & (!g2196) & (!g2197)) + ((g2760) & (g2100) & (g2099) & (g2098) & (!g2196) & (g2197)) + ((g2760) & (g2100) & (g2099) & (g2098) & (g2196) & (!g2197)) + ((g2760) & (g2100) & (g2099) & (g2098) & (g2196) & (g2197)));
	assign g2839 = (((!g2537) & (!g2838) & (!g2687) & (g2615) & (g2201) & (g2202)) + ((!g2537) & (!g2838) & (g2687) & (!g2615) & (!g2201) & (g2202)) + ((!g2537) & (!g2838) & (g2687) & (g2615) & (!g2201) & (g2202)) + ((!g2537) & (!g2838) & (g2687) & (g2615) & (g2201) & (g2202)) + ((!g2537) & (g2838) & (!g2687) & (!g2615) & (g2201) & (!g2202)) + ((!g2537) & (g2838) & (!g2687) & (g2615) & (g2201) & (!g2202)) + ((!g2537) & (g2838) & (!g2687) & (g2615) & (g2201) & (g2202)) + ((!g2537) & (g2838) & (g2687) & (!g2615) & (!g2201) & (g2202)) + ((!g2537) & (g2838) & (g2687) & (!g2615) & (g2201) & (!g2202)) + ((!g2537) & (g2838) & (g2687) & (g2615) & (!g2201) & (g2202)) + ((!g2537) & (g2838) & (g2687) & (g2615) & (g2201) & (!g2202)) + ((!g2537) & (g2838) & (g2687) & (g2615) & (g2201) & (g2202)) + ((g2537) & (!g2838) & (!g2687) & (!g2615) & (!g2201) & (!g2202)) + ((g2537) & (!g2838) & (!g2687) & (g2615) & (!g2201) & (!g2202)) + ((g2537) & (!g2838) & (!g2687) & (g2615) & (g2201) & (g2202)) + ((g2537) & (!g2838) & (g2687) & (!g2615) & (!g2201) & (!g2202)) + ((g2537) & (!g2838) & (g2687) & (!g2615) & (!g2201) & (g2202)) + ((g2537) & (!g2838) & (g2687) & (g2615) & (!g2201) & (!g2202)) + ((g2537) & (!g2838) & (g2687) & (g2615) & (!g2201) & (g2202)) + ((g2537) & (!g2838) & (g2687) & (g2615) & (g2201) & (g2202)) + ((g2537) & (g2838) & (!g2687) & (!g2615) & (!g2201) & (!g2202)) + ((g2537) & (g2838) & (!g2687) & (!g2615) & (g2201) & (!g2202)) + ((g2537) & (g2838) & (!g2687) & (g2615) & (!g2201) & (!g2202)) + ((g2537) & (g2838) & (!g2687) & (g2615) & (g2201) & (!g2202)) + ((g2537) & (g2838) & (!g2687) & (g2615) & (g2201) & (g2202)) + ((g2537) & (g2838) & (g2687) & (!g2615) & (!g2201) & (!g2202)) + ((g2537) & (g2838) & (g2687) & (!g2615) & (!g2201) & (g2202)) + ((g2537) & (g2838) & (g2687) & (!g2615) & (g2201) & (!g2202)) + ((g2537) & (g2838) & (g2687) & (g2615) & (!g2201) & (!g2202)) + ((g2537) & (g2838) & (g2687) & (g2615) & (!g2201) & (g2202)) + ((g2537) & (g2838) & (g2687) & (g2615) & (g2201) & (!g2202)) + ((g2537) & (g2838) & (g2687) & (g2615) & (g2201) & (g2202)));
	assign g2840 = (((!g2081) & (!g2124) & (!g2770) & (!g2831) & (!g3140) & (!g2101)) + ((!g2081) & (!g2124) & (!g2770) & (!g2831) & (!g3140) & (g2101)) + ((!g2081) & (!g2124) & (!g2770) & (g2831) & (!g3140) & (!g2101)) + ((!g2081) & (!g2124) & (!g2770) & (g2831) & (!g3140) & (g2101)) + ((!g2081) & (!g2124) & (g2770) & (!g2831) & (!g3140) & (!g2101)) + ((!g2081) & (!g2124) & (g2770) & (!g2831) & (g3140) & (!g2101)) + ((!g2081) & (!g2124) & (g2770) & (g2831) & (!g3140) & (!g2101)) + ((!g2081) & (!g2124) & (g2770) & (g2831) & (g3140) & (!g2101)) + ((!g2081) & (g2124) & (!g2770) & (!g2831) & (!g3140) & (!g2101)) + ((!g2081) & (g2124) & (!g2770) & (!g2831) & (g3140) & (!g2101)) + ((!g2081) & (g2124) & (g2770) & (!g2831) & (!g3140) & (!g2101)) + ((!g2081) & (g2124) & (g2770) & (!g2831) & (g3140) & (!g2101)) + ((!g2081) & (g2124) & (g2770) & (g2831) & (!g3140) & (!g2101)) + ((!g2081) & (g2124) & (g2770) & (g2831) & (g3140) & (!g2101)) + ((g2081) & (!g2124) & (!g2770) & (!g2831) & (!g3140) & (!g2101)) + ((g2081) & (!g2124) & (!g2770) & (!g2831) & (!g3140) & (g2101)) + ((g2081) & (!g2124) & (!g2770) & (g2831) & (!g3140) & (!g2101)) + ((g2081) & (!g2124) & (!g2770) & (g2831) & (!g3140) & (g2101)) + ((g2081) & (!g2124) & (g2770) & (!g2831) & (!g3140) & (!g2101)) + ((g2081) & (!g2124) & (g2770) & (!g2831) & (g3140) & (!g2101)) + ((g2081) & (!g2124) & (g2770) & (g2831) & (!g3140) & (!g2101)) + ((g2081) & (!g2124) & (g2770) & (g2831) & (g3140) & (!g2101)) + ((g2081) & (g2124) & (!g2770) & (!g2831) & (!g3140) & (!g2101)) + ((g2081) & (g2124) & (!g2770) & (!g2831) & (g3140) & (!g2101)) + ((g2081) & (g2124) & (!g2770) & (g2831) & (!g3140) & (g2101)) + ((g2081) & (g2124) & (!g2770) & (g2831) & (g3140) & (g2101)) + ((g2081) & (g2124) & (g2770) & (!g2831) & (!g3140) & (!g2101)) + ((g2081) & (g2124) & (g2770) & (!g2831) & (g3140) & (!g2101)) + ((g2081) & (g2124) & (g2770) & (g2831) & (!g3140) & (!g2101)) + ((g2081) & (g2124) & (g2770) & (g2831) & (g3140) & (!g2101)));
	assign g2841 = (((!g2840) & (!dmem_dat_ix31x) & (!g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2840) & (!dmem_dat_ix31x) & (!g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2840) & (!dmem_dat_ix31x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((!g2840) & (!dmem_dat_ix31x) & (g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2840) & (!dmem_dat_ix31x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((!g2840) & (!dmem_dat_ix31x) & (g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2840) & (!dmem_dat_ix31x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((!g2840) & (!dmem_dat_ix31x) & (g2783) & (g2784) & (g2785) & (g2786)) + ((!g2840) & (dmem_dat_ix31x) & (!g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2840) & (dmem_dat_ix31x) & (!g2783) & (!g2784) & (g2785) & (!g2786)) + ((!g2840) & (dmem_dat_ix31x) & (!g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2840) & (dmem_dat_ix31x) & (!g2783) & (g2784) & (g2785) & (!g2786)) + ((!g2840) & (dmem_dat_ix31x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((!g2840) & (dmem_dat_ix31x) & (g2783) & (!g2784) & (!g2785) & (!g2786)) + ((!g2840) & (dmem_dat_ix31x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((!g2840) & (dmem_dat_ix31x) & (g2783) & (!g2784) & (g2785) & (!g2786)) + ((!g2840) & (dmem_dat_ix31x) & (g2783) & (g2784) & (!g2785) & (!g2786)) + ((!g2840) & (dmem_dat_ix31x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((!g2840) & (dmem_dat_ix31x) & (g2783) & (g2784) & (g2785) & (!g2786)) + ((!g2840) & (dmem_dat_ix31x) & (g2783) & (g2784) & (g2785) & (g2786)) + ((g2840) & (!dmem_dat_ix31x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((g2840) & (!dmem_dat_ix31x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((g2840) & (!dmem_dat_ix31x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((g2840) & (!dmem_dat_ix31x) & (g2783) & (g2784) & (g2785) & (g2786)) + ((g2840) & (dmem_dat_ix31x) & (!g2783) & (!g2784) & (g2785) & (!g2786)) + ((g2840) & (dmem_dat_ix31x) & (!g2783) & (g2784) & (g2785) & (!g2786)) + ((g2840) & (dmem_dat_ix31x) & (!g2783) & (g2784) & (g2785) & (g2786)) + ((g2840) & (dmem_dat_ix31x) & (g2783) & (!g2784) & (!g2785) & (g2786)) + ((g2840) & (dmem_dat_ix31x) & (g2783) & (!g2784) & (g2785) & (!g2786)) + ((g2840) & (dmem_dat_ix31x) & (g2783) & (g2784) & (!g2785) & (g2786)) + ((g2840) & (dmem_dat_ix31x) & (g2783) & (g2784) & (g2785) & (!g2786)) + ((g2840) & (dmem_dat_ix31x) & (g2783) & (g2784) & (g2785) & (g2786)));
	assign g2842 = (((!sk[17]) & (!g74) & (!dmem_ack_i) & (!g75) & (g128)) + ((!sk[17]) & (!g74) & (!dmem_ack_i) & (g75) & (g128)) + ((!sk[17]) & (!g74) & (dmem_ack_i) & (!g75) & (!g128)) + ((!sk[17]) & (!g74) & (dmem_ack_i) & (!g75) & (g128)) + ((!sk[17]) & (!g74) & (dmem_ack_i) & (g75) & (!g128)) + ((!sk[17]) & (!g74) & (dmem_ack_i) & (g75) & (g128)) + ((!sk[17]) & (g74) & (!dmem_ack_i) & (!g75) & (!g128)) + ((!sk[17]) & (g74) & (!dmem_ack_i) & (!g75) & (g128)) + ((!sk[17]) & (g74) & (!dmem_ack_i) & (g75) & (!g128)) + ((!sk[17]) & (g74) & (!dmem_ack_i) & (g75) & (g128)) + ((!sk[17]) & (g74) & (dmem_ack_i) & (!g75) & (!g128)) + ((!sk[17]) & (g74) & (dmem_ack_i) & (!g75) & (g128)) + ((!sk[17]) & (g74) & (dmem_ack_i) & (g75) & (!g128)) + ((!sk[17]) & (g74) & (dmem_ack_i) & (g75) & (g128)) + ((sk[17]) & (!g74) & (!dmem_ack_i) & (!g75) & (!g128)) + ((sk[17]) & (!g74) & (!dmem_ack_i) & (g75) & (!g128)) + ((sk[17]) & (!g74) & (dmem_ack_i) & (!g75) & (!g128)) + ((sk[17]) & (!g74) & (dmem_ack_i) & (g75) & (!g128)) + ((sk[17]) & (!g74) & (dmem_ack_i) & (g75) & (g128)) + ((sk[17]) & (g74) & (!dmem_ack_i) & (!g75) & (!g128)) + ((sk[17]) & (g74) & (!dmem_ack_i) & (!g75) & (g128)) + ((sk[17]) & (g74) & (!dmem_ack_i) & (g75) & (!g128)) + ((sk[17]) & (g74) & (!dmem_ack_i) & (g75) & (g128)) + ((sk[17]) & (g74) & (dmem_ack_i) & (!g75) & (!g128)) + ((sk[17]) & (g74) & (dmem_ack_i) & (!g75) & (g128)) + ((sk[17]) & (g74) & (dmem_ack_i) & (g75) & (!g128)) + ((sk[17]) & (g74) & (dmem_ack_i) & (g75) & (g128)));
	assign g2843 = (((!g2022) & (!g76) & (!g77) & (g104) & (!sk[18]) & (!g122)) + ((!g2022) & (!g76) & (!g77) & (g104) & (!sk[18]) & (g122)) + ((!g2022) & (!g76) & (g77) & (!g104) & (!sk[18]) & (!g122)) + ((!g2022) & (!g76) & (g77) & (!g104) & (!sk[18]) & (g122)) + ((!g2022) & (!g76) & (g77) & (g104) & (!sk[18]) & (!g122)) + ((!g2022) & (!g76) & (g77) & (g104) & (!sk[18]) & (g122)) + ((!g2022) & (g76) & (!g77) & (g104) & (!sk[18]) & (!g122)) + ((!g2022) & (g76) & (!g77) & (g104) & (!sk[18]) & (g122)) + ((!g2022) & (g76) & (g77) & (!g104) & (!sk[18]) & (!g122)) + ((!g2022) & (g76) & (g77) & (!g104) & (!sk[18]) & (g122)) + ((!g2022) & (g76) & (g77) & (g104) & (!sk[18]) & (!g122)) + ((!g2022) & (g76) & (g77) & (g104) & (!sk[18]) & (g122)) + ((g2022) & (!g76) & (!g77) & (!g104) & (!sk[18]) & (!g122)) + ((g2022) & (!g76) & (!g77) & (!g104) & (!sk[18]) & (g122)) + ((g2022) & (!g76) & (!g77) & (!g104) & (sk[18]) & (!g122)) + ((g2022) & (!g76) & (!g77) & (!g104) & (sk[18]) & (g122)) + ((g2022) & (!g76) & (!g77) & (g104) & (!sk[18]) & (!g122)) + ((g2022) & (!g76) & (!g77) & (g104) & (!sk[18]) & (g122)) + ((g2022) & (!g76) & (!g77) & (g104) & (sk[18]) & (!g122)) + ((g2022) & (!g76) & (g77) & (!g104) & (!sk[18]) & (!g122)) + ((g2022) & (!g76) & (g77) & (!g104) & (!sk[18]) & (g122)) + ((g2022) & (!g76) & (g77) & (g104) & (!sk[18]) & (!g122)) + ((g2022) & (!g76) & (g77) & (g104) & (!sk[18]) & (g122)) + ((g2022) & (g76) & (!g77) & (!g104) & (!sk[18]) & (!g122)) + ((g2022) & (g76) & (!g77) & (!g104) & (!sk[18]) & (g122)) + ((g2022) & (g76) & (!g77) & (g104) & (!sk[18]) & (!g122)) + ((g2022) & (g76) & (!g77) & (g104) & (!sk[18]) & (g122)) + ((g2022) & (g76) & (g77) & (!g104) & (!sk[18]) & (!g122)) + ((g2022) & (g76) & (g77) & (!g104) & (!sk[18]) & (g122)) + ((g2022) & (g76) & (g77) & (g104) & (!sk[18]) & (!g122)) + ((g2022) & (g76) & (g77) & (g104) & (!sk[18]) & (g122)));
	assign g2844 = (((!g74) & (!dmem_ack_i) & (!g75) & (!nmi_i) & (g2023) & (!g2843)) + ((!g74) & (!dmem_ack_i) & (!g75) & (!nmi_i) & (g2023) & (g2843)) + ((!g74) & (!dmem_ack_i) & (!g75) & (nmi_i) & (!g2023) & (!g2843)) + ((!g74) & (!dmem_ack_i) & (!g75) & (nmi_i) & (!g2023) & (g2843)) + ((!g74) & (!dmem_ack_i) & (!g75) & (nmi_i) & (g2023) & (!g2843)) + ((!g74) & (!dmem_ack_i) & (!g75) & (nmi_i) & (g2023) & (g2843)) + ((!g74) & (!dmem_ack_i) & (g75) & (!nmi_i) & (g2023) & (!g2843)) + ((!g74) & (!dmem_ack_i) & (g75) & (!nmi_i) & (g2023) & (g2843)) + ((!g74) & (!dmem_ack_i) & (g75) & (nmi_i) & (!g2023) & (!g2843)) + ((!g74) & (!dmem_ack_i) & (g75) & (nmi_i) & (!g2023) & (g2843)) + ((!g74) & (!dmem_ack_i) & (g75) & (nmi_i) & (g2023) & (!g2843)) + ((!g74) & (!dmem_ack_i) & (g75) & (nmi_i) & (g2023) & (g2843)) + ((!g74) & (dmem_ack_i) & (!g75) & (!nmi_i) & (g2023) & (!g2843)) + ((!g74) & (dmem_ack_i) & (!g75) & (!nmi_i) & (g2023) & (g2843)) + ((!g74) & (dmem_ack_i) & (!g75) & (nmi_i) & (!g2023) & (!g2843)) + ((!g74) & (dmem_ack_i) & (!g75) & (nmi_i) & (!g2023) & (g2843)) + ((!g74) & (dmem_ack_i) & (!g75) & (nmi_i) & (g2023) & (!g2843)) + ((!g74) & (dmem_ack_i) & (!g75) & (nmi_i) & (g2023) & (g2843)) + ((!g74) & (dmem_ack_i) & (g75) & (!nmi_i) & (g2023) & (!g2843)) + ((!g74) & (dmem_ack_i) & (g75) & (nmi_i) & (!g2023) & (!g2843)) + ((!g74) & (dmem_ack_i) & (g75) & (nmi_i) & (g2023) & (!g2843)) + ((g74) & (!dmem_ack_i) & (!g75) & (!nmi_i) & (g2023) & (!g2843)) + ((g74) & (!dmem_ack_i) & (!g75) & (nmi_i) & (!g2023) & (!g2843)) + ((g74) & (!dmem_ack_i) & (!g75) & (nmi_i) & (g2023) & (!g2843)) + ((g74) & (!dmem_ack_i) & (g75) & (!nmi_i) & (g2023) & (!g2843)) + ((g74) & (!dmem_ack_i) & (g75) & (nmi_i) & (!g2023) & (!g2843)) + ((g74) & (!dmem_ack_i) & (g75) & (nmi_i) & (g2023) & (!g2843)) + ((g74) & (dmem_ack_i) & (!g75) & (!nmi_i) & (g2023) & (!g2843)) + ((g74) & (dmem_ack_i) & (!g75) & (nmi_i) & (!g2023) & (!g2843)) + ((g74) & (dmem_ack_i) & (!g75) & (nmi_i) & (g2023) & (!g2843)) + ((g74) & (dmem_ack_i) & (g75) & (!nmi_i) & (g2023) & (!g2843)) + ((g74) & (dmem_ack_i) & (g75) & (nmi_i) & (!g2023) & (!g2843)) + ((g74) & (dmem_ack_i) & (g75) & (nmi_i) & (g2023) & (!g2843)));
	assign g2845 = (((!sk[20]) & (!g80) & (g82) & (!g83)) + ((!sk[20]) & (!g80) & (g82) & (g83)) + ((!sk[20]) & (g80) & (!g82) & (!g83)) + ((!sk[20]) & (g80) & (!g82) & (g83)) + ((!sk[20]) & (g80) & (g82) & (!g83)) + ((!sk[20]) & (g80) & (g82) & (g83)) + ((sk[20]) & (g80) & (g82) & (g83)));
	assign g2846 = (((!sk[21]) & (!g2845) & (g107)) + ((!sk[21]) & (g2845) & (g107)) + ((sk[21]) & (g2845) & (!g107)));
	assign g2847 = (((!sk[22]) & (!g108) & (g109) & (!g2846)) + ((!sk[22]) & (!g108) & (g109) & (g2846)) + ((!sk[22]) & (g108) & (!g109) & (!g2846)) + ((!sk[22]) & (g108) & (!g109) & (g2846)) + ((!sk[22]) & (g108) & (g109) & (!g2846)) + ((!sk[22]) & (g108) & (g109) & (g2846)) + ((sk[22]) & (!g108) & (g109) & (g2846)));
	assign g2848 = (((!g2090) & (!g2091) & (!g2098) & (!g2734) & (!g2751) & (!g2771)) + ((!g2090) & (!g2091) & (g2098) & (!g2734) & (!g2751) & (g2771)) + ((!g2090) & (g2091) & (!g2098) & (!g2734) & (g2751) & (!g2771)) + ((!g2090) & (g2091) & (g2098) & (!g2734) & (g2751) & (g2771)) + ((g2090) & (!g2091) & (!g2098) & (g2734) & (!g2751) & (!g2771)) + ((g2090) & (!g2091) & (g2098) & (g2734) & (!g2751) & (g2771)) + ((g2090) & (g2091) & (!g2098) & (g2734) & (g2751) & (!g2771)) + ((g2090) & (g2091) & (g2098) & (g2734) & (g2751) & (g2771)));
	assign g2849 = (((!g2088) & (!sk[24]) & (!g2089) & (!g2699) & (g2715) & (!g2848)) + ((!g2088) & (!sk[24]) & (!g2089) & (!g2699) & (g2715) & (g2848)) + ((!g2088) & (!sk[24]) & (!g2089) & (g2699) & (!g2715) & (!g2848)) + ((!g2088) & (!sk[24]) & (!g2089) & (g2699) & (!g2715) & (g2848)) + ((!g2088) & (!sk[24]) & (!g2089) & (g2699) & (g2715) & (!g2848)) + ((!g2088) & (!sk[24]) & (!g2089) & (g2699) & (g2715) & (g2848)) + ((!g2088) & (!sk[24]) & (g2089) & (!g2699) & (g2715) & (!g2848)) + ((!g2088) & (!sk[24]) & (g2089) & (!g2699) & (g2715) & (g2848)) + ((!g2088) & (!sk[24]) & (g2089) & (g2699) & (!g2715) & (!g2848)) + ((!g2088) & (!sk[24]) & (g2089) & (g2699) & (!g2715) & (g2848)) + ((!g2088) & (!sk[24]) & (g2089) & (g2699) & (g2715) & (!g2848)) + ((!g2088) & (!sk[24]) & (g2089) & (g2699) & (g2715) & (g2848)) + ((!g2088) & (sk[24]) & (!g2089) & (!g2699) & (!g2715) & (g2848)) + ((!g2088) & (sk[24]) & (g2089) & (!g2699) & (g2715) & (g2848)) + ((g2088) & (!sk[24]) & (!g2089) & (!g2699) & (!g2715) & (!g2848)) + ((g2088) & (!sk[24]) & (!g2089) & (!g2699) & (!g2715) & (g2848)) + ((g2088) & (!sk[24]) & (!g2089) & (!g2699) & (g2715) & (!g2848)) + ((g2088) & (!sk[24]) & (!g2089) & (!g2699) & (g2715) & (g2848)) + ((g2088) & (!sk[24]) & (!g2089) & (g2699) & (!g2715) & (!g2848)) + ((g2088) & (!sk[24]) & (!g2089) & (g2699) & (!g2715) & (g2848)) + ((g2088) & (!sk[24]) & (!g2089) & (g2699) & (g2715) & (!g2848)) + ((g2088) & (!sk[24]) & (!g2089) & (g2699) & (g2715) & (g2848)) + ((g2088) & (!sk[24]) & (g2089) & (!g2699) & (!g2715) & (!g2848)) + ((g2088) & (!sk[24]) & (g2089) & (!g2699) & (!g2715) & (g2848)) + ((g2088) & (!sk[24]) & (g2089) & (!g2699) & (g2715) & (!g2848)) + ((g2088) & (!sk[24]) & (g2089) & (!g2699) & (g2715) & (g2848)) + ((g2088) & (!sk[24]) & (g2089) & (g2699) & (!g2715) & (!g2848)) + ((g2088) & (!sk[24]) & (g2089) & (g2699) & (!g2715) & (g2848)) + ((g2088) & (!sk[24]) & (g2089) & (g2699) & (g2715) & (!g2848)) + ((g2088) & (!sk[24]) & (g2089) & (g2699) & (g2715) & (g2848)) + ((g2088) & (sk[24]) & (!g2089) & (g2699) & (!g2715) & (g2848)) + ((g2088) & (sk[24]) & (g2089) & (g2699) & (g2715) & (g2848)));
	assign g2850 = (((!g2095) & (!sk[25]) & (!g2096) & (!g2660) & (g2680) & (!g2849)) + ((!g2095) & (!sk[25]) & (!g2096) & (!g2660) & (g2680) & (g2849)) + ((!g2095) & (!sk[25]) & (!g2096) & (g2660) & (!g2680) & (!g2849)) + ((!g2095) & (!sk[25]) & (!g2096) & (g2660) & (!g2680) & (g2849)) + ((!g2095) & (!sk[25]) & (!g2096) & (g2660) & (g2680) & (!g2849)) + ((!g2095) & (!sk[25]) & (!g2096) & (g2660) & (g2680) & (g2849)) + ((!g2095) & (!sk[25]) & (g2096) & (!g2660) & (g2680) & (!g2849)) + ((!g2095) & (!sk[25]) & (g2096) & (!g2660) & (g2680) & (g2849)) + ((!g2095) & (!sk[25]) & (g2096) & (g2660) & (!g2680) & (!g2849)) + ((!g2095) & (!sk[25]) & (g2096) & (g2660) & (!g2680) & (g2849)) + ((!g2095) & (!sk[25]) & (g2096) & (g2660) & (g2680) & (!g2849)) + ((!g2095) & (!sk[25]) & (g2096) & (g2660) & (g2680) & (g2849)) + ((!g2095) & (sk[25]) & (!g2096) & (!g2660) & (!g2680) & (g2849)) + ((!g2095) & (sk[25]) & (g2096) & (!g2660) & (g2680) & (g2849)) + ((g2095) & (!sk[25]) & (!g2096) & (!g2660) & (!g2680) & (!g2849)) + ((g2095) & (!sk[25]) & (!g2096) & (!g2660) & (!g2680) & (g2849)) + ((g2095) & (!sk[25]) & (!g2096) & (!g2660) & (g2680) & (!g2849)) + ((g2095) & (!sk[25]) & (!g2096) & (!g2660) & (g2680) & (g2849)) + ((g2095) & (!sk[25]) & (!g2096) & (g2660) & (!g2680) & (!g2849)) + ((g2095) & (!sk[25]) & (!g2096) & (g2660) & (!g2680) & (g2849)) + ((g2095) & (!sk[25]) & (!g2096) & (g2660) & (g2680) & (!g2849)) + ((g2095) & (!sk[25]) & (!g2096) & (g2660) & (g2680) & (g2849)) + ((g2095) & (!sk[25]) & (g2096) & (!g2660) & (!g2680) & (!g2849)) + ((g2095) & (!sk[25]) & (g2096) & (!g2660) & (!g2680) & (g2849)) + ((g2095) & (!sk[25]) & (g2096) & (!g2660) & (g2680) & (!g2849)) + ((g2095) & (!sk[25]) & (g2096) & (!g2660) & (g2680) & (g2849)) + ((g2095) & (!sk[25]) & (g2096) & (g2660) & (!g2680) & (!g2849)) + ((g2095) & (!sk[25]) & (g2096) & (g2660) & (!g2680) & (g2849)) + ((g2095) & (!sk[25]) & (g2096) & (g2660) & (g2680) & (!g2849)) + ((g2095) & (!sk[25]) & (g2096) & (g2660) & (g2680) & (g2849)) + ((g2095) & (sk[25]) & (!g2096) & (g2660) & (!g2680) & (g2849)) + ((g2095) & (sk[25]) & (g2096) & (g2660) & (g2680) & (g2849)));
	assign g2851 = (((!g2110) & (!g2111) & (!g2418) & (!sk[26]) & (g2439)) + ((!g2110) & (!g2111) & (!g2418) & (sk[26]) & (!g2439)) + ((!g2110) & (!g2111) & (g2418) & (!sk[26]) & (g2439)) + ((!g2110) & (g2111) & (!g2418) & (!sk[26]) & (!g2439)) + ((!g2110) & (g2111) & (!g2418) & (!sk[26]) & (g2439)) + ((!g2110) & (g2111) & (!g2418) & (sk[26]) & (g2439)) + ((!g2110) & (g2111) & (g2418) & (!sk[26]) & (!g2439)) + ((!g2110) & (g2111) & (g2418) & (!sk[26]) & (g2439)) + ((g2110) & (!g2111) & (!g2418) & (!sk[26]) & (!g2439)) + ((g2110) & (!g2111) & (!g2418) & (!sk[26]) & (g2439)) + ((g2110) & (!g2111) & (g2418) & (!sk[26]) & (!g2439)) + ((g2110) & (!g2111) & (g2418) & (!sk[26]) & (g2439)) + ((g2110) & (!g2111) & (g2418) & (sk[26]) & (!g2439)) + ((g2110) & (g2111) & (!g2418) & (!sk[26]) & (!g2439)) + ((g2110) & (g2111) & (!g2418) & (!sk[26]) & (g2439)) + ((g2110) & (g2111) & (g2418) & (!sk[26]) & (!g2439)) + ((g2110) & (g2111) & (g2418) & (!sk[26]) & (g2439)) + ((g2110) & (g2111) & (g2418) & (sk[26]) & (g2439)));
	assign g2852 = (((!sk[27]) & (!g2109) & (g2391) & (!g2851)) + ((!sk[27]) & (!g2109) & (g2391) & (g2851)) + ((!sk[27]) & (g2109) & (!g2391) & (!g2851)) + ((!sk[27]) & (g2109) & (!g2391) & (g2851)) + ((!sk[27]) & (g2109) & (g2391) & (!g2851)) + ((!sk[27]) & (g2109) & (g2391) & (g2851)) + ((sk[27]) & (!g2109) & (!g2391) & (g2851)) + ((sk[27]) & (g2109) & (g2391) & (g2851)));
	assign g2853 = (((!g2108) & (!g2116) & (!g2340) & (!g2365) & (sk[28]) & (g2852)) + ((!g2108) & (!g2116) & (!g2340) & (g2365) & (!sk[28]) & (!g2852)) + ((!g2108) & (!g2116) & (!g2340) & (g2365) & (!sk[28]) & (g2852)) + ((!g2108) & (!g2116) & (g2340) & (!g2365) & (!sk[28]) & (!g2852)) + ((!g2108) & (!g2116) & (g2340) & (!g2365) & (!sk[28]) & (g2852)) + ((!g2108) & (!g2116) & (g2340) & (g2365) & (!sk[28]) & (!g2852)) + ((!g2108) & (!g2116) & (g2340) & (g2365) & (!sk[28]) & (g2852)) + ((!g2108) & (g2116) & (!g2340) & (g2365) & (!sk[28]) & (!g2852)) + ((!g2108) & (g2116) & (!g2340) & (g2365) & (!sk[28]) & (g2852)) + ((!g2108) & (g2116) & (g2340) & (!g2365) & (!sk[28]) & (!g2852)) + ((!g2108) & (g2116) & (g2340) & (!g2365) & (!sk[28]) & (g2852)) + ((!g2108) & (g2116) & (g2340) & (!g2365) & (sk[28]) & (g2852)) + ((!g2108) & (g2116) & (g2340) & (g2365) & (!sk[28]) & (!g2852)) + ((!g2108) & (g2116) & (g2340) & (g2365) & (!sk[28]) & (g2852)) + ((g2108) & (!g2116) & (!g2340) & (!g2365) & (!sk[28]) & (!g2852)) + ((g2108) & (!g2116) & (!g2340) & (!g2365) & (!sk[28]) & (g2852)) + ((g2108) & (!g2116) & (!g2340) & (g2365) & (!sk[28]) & (!g2852)) + ((g2108) & (!g2116) & (!g2340) & (g2365) & (!sk[28]) & (g2852)) + ((g2108) & (!g2116) & (!g2340) & (g2365) & (sk[28]) & (g2852)) + ((g2108) & (!g2116) & (g2340) & (!g2365) & (!sk[28]) & (!g2852)) + ((g2108) & (!g2116) & (g2340) & (!g2365) & (!sk[28]) & (g2852)) + ((g2108) & (!g2116) & (g2340) & (g2365) & (!sk[28]) & (!g2852)) + ((g2108) & (!g2116) & (g2340) & (g2365) & (!sk[28]) & (g2852)) + ((g2108) & (g2116) & (!g2340) & (!g2365) & (!sk[28]) & (!g2852)) + ((g2108) & (g2116) & (!g2340) & (!g2365) & (!sk[28]) & (g2852)) + ((g2108) & (g2116) & (!g2340) & (g2365) & (!sk[28]) & (!g2852)) + ((g2108) & (g2116) & (!g2340) & (g2365) & (!sk[28]) & (g2852)) + ((g2108) & (g2116) & (g2340) & (!g2365) & (!sk[28]) & (!g2852)) + ((g2108) & (g2116) & (g2340) & (!g2365) & (!sk[28]) & (g2852)) + ((g2108) & (g2116) & (g2340) & (g2365) & (!sk[28]) & (!g2852)) + ((g2108) & (g2116) & (g2340) & (g2365) & (!sk[28]) & (g2852)) + ((g2108) & (g2116) & (g2340) & (g2365) & (sk[28]) & (g2852)));
	assign g2854 = (((!g2086) & (!g2093) & (!g2094) & (!g2608) & (!g2625) & (!g2642)) + ((!g2086) & (!g2093) & (g2094) & (!g2608) & (!g2625) & (g2642)) + ((!g2086) & (g2093) & (!g2094) & (!g2608) & (g2625) & (!g2642)) + ((!g2086) & (g2093) & (g2094) & (!g2608) & (g2625) & (g2642)) + ((g2086) & (!g2093) & (!g2094) & (g2608) & (!g2625) & (!g2642)) + ((g2086) & (!g2093) & (g2094) & (g2608) & (!g2625) & (g2642)) + ((g2086) & (g2093) & (!g2094) & (g2608) & (g2625) & (!g2642)) + ((g2086) & (g2093) & (g2094) & (g2608) & (g2625) & (g2642)));
	assign g2855 = (((!sk[30]) & (!g2084) & (!g2085) & (!g2570) & (g2590) & (!g2854)) + ((!sk[30]) & (!g2084) & (!g2085) & (!g2570) & (g2590) & (g2854)) + ((!sk[30]) & (!g2084) & (!g2085) & (g2570) & (!g2590) & (!g2854)) + ((!sk[30]) & (!g2084) & (!g2085) & (g2570) & (!g2590) & (g2854)) + ((!sk[30]) & (!g2084) & (!g2085) & (g2570) & (g2590) & (!g2854)) + ((!sk[30]) & (!g2084) & (!g2085) & (g2570) & (g2590) & (g2854)) + ((!sk[30]) & (!g2084) & (g2085) & (!g2570) & (g2590) & (!g2854)) + ((!sk[30]) & (!g2084) & (g2085) & (!g2570) & (g2590) & (g2854)) + ((!sk[30]) & (!g2084) & (g2085) & (g2570) & (!g2590) & (!g2854)) + ((!sk[30]) & (!g2084) & (g2085) & (g2570) & (!g2590) & (g2854)) + ((!sk[30]) & (!g2084) & (g2085) & (g2570) & (g2590) & (!g2854)) + ((!sk[30]) & (!g2084) & (g2085) & (g2570) & (g2590) & (g2854)) + ((!sk[30]) & (g2084) & (!g2085) & (!g2570) & (!g2590) & (!g2854)) + ((!sk[30]) & (g2084) & (!g2085) & (!g2570) & (!g2590) & (g2854)) + ((!sk[30]) & (g2084) & (!g2085) & (!g2570) & (g2590) & (!g2854)) + ((!sk[30]) & (g2084) & (!g2085) & (!g2570) & (g2590) & (g2854)) + ((!sk[30]) & (g2084) & (!g2085) & (g2570) & (!g2590) & (!g2854)) + ((!sk[30]) & (g2084) & (!g2085) & (g2570) & (!g2590) & (g2854)) + ((!sk[30]) & (g2084) & (!g2085) & (g2570) & (g2590) & (!g2854)) + ((!sk[30]) & (g2084) & (!g2085) & (g2570) & (g2590) & (g2854)) + ((!sk[30]) & (g2084) & (g2085) & (!g2570) & (!g2590) & (!g2854)) + ((!sk[30]) & (g2084) & (g2085) & (!g2570) & (!g2590) & (g2854)) + ((!sk[30]) & (g2084) & (g2085) & (!g2570) & (g2590) & (!g2854)) + ((!sk[30]) & (g2084) & (g2085) & (!g2570) & (g2590) & (g2854)) + ((!sk[30]) & (g2084) & (g2085) & (g2570) & (!g2590) & (!g2854)) + ((!sk[30]) & (g2084) & (g2085) & (g2570) & (!g2590) & (g2854)) + ((!sk[30]) & (g2084) & (g2085) & (g2570) & (g2590) & (!g2854)) + ((!sk[30]) & (g2084) & (g2085) & (g2570) & (g2590) & (g2854)) + ((sk[30]) & (!g2084) & (!g2085) & (!g2570) & (!g2590) & (g2854)) + ((sk[30]) & (!g2084) & (g2085) & (!g2570) & (g2590) & (g2854)) + ((sk[30]) & (g2084) & (!g2085) & (g2570) & (!g2590) & (g2854)) + ((sk[30]) & (g2084) & (g2085) & (g2570) & (g2590) & (g2854)));
	assign g2856 = (((!sk[31]) & (!g2083) & (!g2121) & (!g2529) & (g2551) & (!g2855)) + ((!sk[31]) & (!g2083) & (!g2121) & (!g2529) & (g2551) & (g2855)) + ((!sk[31]) & (!g2083) & (!g2121) & (g2529) & (!g2551) & (!g2855)) + ((!sk[31]) & (!g2083) & (!g2121) & (g2529) & (!g2551) & (g2855)) + ((!sk[31]) & (!g2083) & (!g2121) & (g2529) & (g2551) & (!g2855)) + ((!sk[31]) & (!g2083) & (!g2121) & (g2529) & (g2551) & (g2855)) + ((!sk[31]) & (!g2083) & (g2121) & (!g2529) & (g2551) & (!g2855)) + ((!sk[31]) & (!g2083) & (g2121) & (!g2529) & (g2551) & (g2855)) + ((!sk[31]) & (!g2083) & (g2121) & (g2529) & (!g2551) & (!g2855)) + ((!sk[31]) & (!g2083) & (g2121) & (g2529) & (!g2551) & (g2855)) + ((!sk[31]) & (!g2083) & (g2121) & (g2529) & (g2551) & (!g2855)) + ((!sk[31]) & (!g2083) & (g2121) & (g2529) & (g2551) & (g2855)) + ((!sk[31]) & (g2083) & (!g2121) & (!g2529) & (!g2551) & (!g2855)) + ((!sk[31]) & (g2083) & (!g2121) & (!g2529) & (!g2551) & (g2855)) + ((!sk[31]) & (g2083) & (!g2121) & (!g2529) & (g2551) & (!g2855)) + ((!sk[31]) & (g2083) & (!g2121) & (!g2529) & (g2551) & (g2855)) + ((!sk[31]) & (g2083) & (!g2121) & (g2529) & (!g2551) & (!g2855)) + ((!sk[31]) & (g2083) & (!g2121) & (g2529) & (!g2551) & (g2855)) + ((!sk[31]) & (g2083) & (!g2121) & (g2529) & (g2551) & (!g2855)) + ((!sk[31]) & (g2083) & (!g2121) & (g2529) & (g2551) & (g2855)) + ((!sk[31]) & (g2083) & (g2121) & (!g2529) & (!g2551) & (!g2855)) + ((!sk[31]) & (g2083) & (g2121) & (!g2529) & (!g2551) & (g2855)) + ((!sk[31]) & (g2083) & (g2121) & (!g2529) & (g2551) & (!g2855)) + ((!sk[31]) & (g2083) & (g2121) & (!g2529) & (g2551) & (g2855)) + ((!sk[31]) & (g2083) & (g2121) & (g2529) & (!g2551) & (!g2855)) + ((!sk[31]) & (g2083) & (g2121) & (g2529) & (!g2551) & (g2855)) + ((!sk[31]) & (g2083) & (g2121) & (g2529) & (g2551) & (!g2855)) + ((!sk[31]) & (g2083) & (g2121) & (g2529) & (g2551) & (g2855)) + ((sk[31]) & (!g2083) & (!g2121) & (!g2529) & (!g2551) & (g2855)) + ((sk[31]) & (!g2083) & (g2121) & (g2529) & (!g2551) & (g2855)) + ((sk[31]) & (g2083) & (!g2121) & (!g2529) & (g2551) & (g2855)) + ((sk[31]) & (g2083) & (g2121) & (g2529) & (g2551) & (g2855)));
	assign g2857 = (((!g2100) & (!g2101) & (!g2811) & (!sk[32]) & (g2831)) + ((!g2100) & (!g2101) & (!g2811) & (sk[32]) & (!g2831)) + ((!g2100) & (!g2101) & (g2811) & (!sk[32]) & (g2831)) + ((!g2100) & (g2101) & (!g2811) & (!sk[32]) & (!g2831)) + ((!g2100) & (g2101) & (!g2811) & (!sk[32]) & (g2831)) + ((!g2100) & (g2101) & (!g2811) & (sk[32]) & (g2831)) + ((!g2100) & (g2101) & (g2811) & (!sk[32]) & (!g2831)) + ((!g2100) & (g2101) & (g2811) & (!sk[32]) & (g2831)) + ((g2100) & (!g2101) & (!g2811) & (!sk[32]) & (!g2831)) + ((g2100) & (!g2101) & (!g2811) & (!sk[32]) & (g2831)) + ((g2100) & (!g2101) & (g2811) & (!sk[32]) & (!g2831)) + ((g2100) & (!g2101) & (g2811) & (!sk[32]) & (g2831)) + ((g2100) & (!g2101) & (g2811) & (sk[32]) & (!g2831)) + ((g2100) & (g2101) & (!g2811) & (!sk[32]) & (!g2831)) + ((g2100) & (g2101) & (!g2811) & (!sk[32]) & (g2831)) + ((g2100) & (g2101) & (g2811) & (!sk[32]) & (!g2831)) + ((g2100) & (g2101) & (g2811) & (!sk[32]) & (g2831)) + ((g2100) & (g2101) & (g2811) & (sk[32]) & (g2831)));
	assign g2858 = (((!g2119) & (!g2120) & (!sk[33]) & (!g2482) & (g2507)) + ((!g2119) & (!g2120) & (!sk[33]) & (g2482) & (g2507)) + ((!g2119) & (!g2120) & (sk[33]) & (!g2482) & (!g2507)) + ((!g2119) & (g2120) & (!sk[33]) & (!g2482) & (!g2507)) + ((!g2119) & (g2120) & (!sk[33]) & (!g2482) & (g2507)) + ((!g2119) & (g2120) & (!sk[33]) & (g2482) & (!g2507)) + ((!g2119) & (g2120) & (!sk[33]) & (g2482) & (g2507)) + ((!g2119) & (g2120) & (sk[33]) & (!g2482) & (g2507)) + ((g2119) & (!g2120) & (!sk[33]) & (!g2482) & (!g2507)) + ((g2119) & (!g2120) & (!sk[33]) & (!g2482) & (g2507)) + ((g2119) & (!g2120) & (!sk[33]) & (g2482) & (!g2507)) + ((g2119) & (!g2120) & (!sk[33]) & (g2482) & (g2507)) + ((g2119) & (!g2120) & (sk[33]) & (g2482) & (!g2507)) + ((g2119) & (g2120) & (!sk[33]) & (!g2482) & (!g2507)) + ((g2119) & (g2120) & (!sk[33]) & (!g2482) & (g2507)) + ((g2119) & (g2120) & (!sk[33]) & (g2482) & (!g2507)) + ((g2119) & (g2120) & (!sk[33]) & (g2482) & (g2507)) + ((g2119) & (g2120) & (sk[33]) & (g2482) & (g2507)));
	assign g2859 = (((!sk[34]) & (!g2118) & (g2457) & (!g2858)) + ((!sk[34]) & (!g2118) & (g2457) & (g2858)) + ((!sk[34]) & (g2118) & (!g2457) & (!g2858)) + ((!sk[34]) & (g2118) & (!g2457) & (g2858)) + ((!sk[34]) & (g2118) & (g2457) & (!g2858)) + ((!sk[34]) & (g2118) & (g2457) & (g2858)) + ((sk[34]) & (!g2118) & (!g2457) & (g2858)) + ((sk[34]) & (g2118) & (g2457) & (g2858)));
	assign g2860 = (((!g2073) & (!sk[35]) & (!g2113) & (!g2114) & (g2289)) + ((!g2073) & (!sk[35]) & (!g2113) & (g2114) & (g2289)) + ((!g2073) & (!sk[35]) & (g2113) & (!g2114) & (!g2289)) + ((!g2073) & (!sk[35]) & (g2113) & (!g2114) & (g2289)) + ((!g2073) & (!sk[35]) & (g2113) & (g2114) & (!g2289)) + ((!g2073) & (!sk[35]) & (g2113) & (g2114) & (g2289)) + ((!g2073) & (sk[35]) & (!g2113) & (!g2114) & (!g2289)) + ((!g2073) & (sk[35]) & (!g2113) & (g2114) & (g2289)) + ((g2073) & (!sk[35]) & (!g2113) & (!g2114) & (!g2289)) + ((g2073) & (!sk[35]) & (!g2113) & (!g2114) & (g2289)) + ((g2073) & (!sk[35]) & (!g2113) & (g2114) & (!g2289)) + ((g2073) & (!sk[35]) & (!g2113) & (g2114) & (g2289)) + ((g2073) & (!sk[35]) & (g2113) & (!g2114) & (!g2289)) + ((g2073) & (!sk[35]) & (g2113) & (!g2114) & (g2289)) + ((g2073) & (!sk[35]) & (g2113) & (g2114) & (!g2289)) + ((g2073) & (!sk[35]) & (g2113) & (g2114) & (g2289)) + ((g2073) & (sk[35]) & (g2113) & (!g2114) & (!g2289)) + ((g2073) & (sk[35]) & (g2113) & (g2114) & (g2289)));
	assign g2861 = (((!g2074) & (!g2076) & (!g2077) & (!g2105) & (!g2104) & (!g2106)) + ((!g2074) & (!g2076) & (g2077) & (g2105) & (!g2104) & (!g2106)) + ((!g2074) & (g2076) & (!g2077) & (!g2105) & (!g2104) & (g2106)) + ((!g2074) & (g2076) & (g2077) & (g2105) & (!g2104) & (g2106)) + ((g2074) & (!g2076) & (!g2077) & (!g2105) & (g2104) & (!g2106)) + ((g2074) & (!g2076) & (g2077) & (g2105) & (g2104) & (!g2106)) + ((g2074) & (g2076) & (!g2077) & (!g2105) & (g2104) & (g2106)) + ((g2074) & (g2076) & (g2077) & (g2105) & (g2104) & (g2106)));
	assign g2862 = (((!g2071) & (!sk[37]) & (!g2070) & (!g2859) & (g2860) & (!g2861)) + ((!g2071) & (!sk[37]) & (!g2070) & (!g2859) & (g2860) & (g2861)) + ((!g2071) & (!sk[37]) & (!g2070) & (g2859) & (!g2860) & (!g2861)) + ((!g2071) & (!sk[37]) & (!g2070) & (g2859) & (!g2860) & (g2861)) + ((!g2071) & (!sk[37]) & (!g2070) & (g2859) & (g2860) & (!g2861)) + ((!g2071) & (!sk[37]) & (!g2070) & (g2859) & (g2860) & (g2861)) + ((!g2071) & (!sk[37]) & (g2070) & (!g2859) & (g2860) & (!g2861)) + ((!g2071) & (!sk[37]) & (g2070) & (!g2859) & (g2860) & (g2861)) + ((!g2071) & (!sk[37]) & (g2070) & (g2859) & (!g2860) & (!g2861)) + ((!g2071) & (!sk[37]) & (g2070) & (g2859) & (!g2860) & (g2861)) + ((!g2071) & (!sk[37]) & (g2070) & (g2859) & (g2860) & (!g2861)) + ((!g2071) & (!sk[37]) & (g2070) & (g2859) & (g2860) & (g2861)) + ((!g2071) & (sk[37]) & (!g2070) & (g2859) & (g2860) & (g2861)) + ((g2071) & (!sk[37]) & (!g2070) & (!g2859) & (!g2860) & (!g2861)) + ((g2071) & (!sk[37]) & (!g2070) & (!g2859) & (!g2860) & (g2861)) + ((g2071) & (!sk[37]) & (!g2070) & (!g2859) & (g2860) & (!g2861)) + ((g2071) & (!sk[37]) & (!g2070) & (!g2859) & (g2860) & (g2861)) + ((g2071) & (!sk[37]) & (!g2070) & (g2859) & (!g2860) & (!g2861)) + ((g2071) & (!sk[37]) & (!g2070) & (g2859) & (!g2860) & (g2861)) + ((g2071) & (!sk[37]) & (!g2070) & (g2859) & (g2860) & (!g2861)) + ((g2071) & (!sk[37]) & (!g2070) & (g2859) & (g2860) & (g2861)) + ((g2071) & (!sk[37]) & (g2070) & (!g2859) & (!g2860) & (!g2861)) + ((g2071) & (!sk[37]) & (g2070) & (!g2859) & (!g2860) & (g2861)) + ((g2071) & (!sk[37]) & (g2070) & (!g2859) & (g2860) & (!g2861)) + ((g2071) & (!sk[37]) & (g2070) & (!g2859) & (g2860) & (g2861)) + ((g2071) & (!sk[37]) & (g2070) & (g2859) & (!g2860) & (!g2861)) + ((g2071) & (!sk[37]) & (g2070) & (g2859) & (!g2860) & (g2861)) + ((g2071) & (!sk[37]) & (g2070) & (g2859) & (g2860) & (!g2861)) + ((g2071) & (!sk[37]) & (g2070) & (g2859) & (g2860) & (g2861)) + ((g2071) & (sk[37]) & (g2070) & (g2859) & (g2860) & (g2861)));
	assign g2863 = (((!g2099) & (!g2794) & (!g2856) & (g2857) & (!sk[38]) & (!g2862)) + ((!g2099) & (!g2794) & (!g2856) & (g2857) & (!sk[38]) & (g2862)) + ((!g2099) & (!g2794) & (g2856) & (!g2857) & (!sk[38]) & (!g2862)) + ((!g2099) & (!g2794) & (g2856) & (!g2857) & (!sk[38]) & (g2862)) + ((!g2099) & (!g2794) & (g2856) & (g2857) & (!sk[38]) & (!g2862)) + ((!g2099) & (!g2794) & (g2856) & (g2857) & (!sk[38]) & (g2862)) + ((!g2099) & (!g2794) & (g2856) & (g2857) & (sk[38]) & (g2862)) + ((!g2099) & (g2794) & (!g2856) & (g2857) & (!sk[38]) & (!g2862)) + ((!g2099) & (g2794) & (!g2856) & (g2857) & (!sk[38]) & (g2862)) + ((!g2099) & (g2794) & (g2856) & (!g2857) & (!sk[38]) & (!g2862)) + ((!g2099) & (g2794) & (g2856) & (!g2857) & (!sk[38]) & (g2862)) + ((!g2099) & (g2794) & (g2856) & (g2857) & (!sk[38]) & (!g2862)) + ((!g2099) & (g2794) & (g2856) & (g2857) & (!sk[38]) & (g2862)) + ((g2099) & (!g2794) & (!g2856) & (!g2857) & (!sk[38]) & (!g2862)) + ((g2099) & (!g2794) & (!g2856) & (!g2857) & (!sk[38]) & (g2862)) + ((g2099) & (!g2794) & (!g2856) & (g2857) & (!sk[38]) & (!g2862)) + ((g2099) & (!g2794) & (!g2856) & (g2857) & (!sk[38]) & (g2862)) + ((g2099) & (!g2794) & (g2856) & (!g2857) & (!sk[38]) & (!g2862)) + ((g2099) & (!g2794) & (g2856) & (!g2857) & (!sk[38]) & (g2862)) + ((g2099) & (!g2794) & (g2856) & (g2857) & (!sk[38]) & (!g2862)) + ((g2099) & (!g2794) & (g2856) & (g2857) & (!sk[38]) & (g2862)) + ((g2099) & (g2794) & (!g2856) & (!g2857) & (!sk[38]) & (!g2862)) + ((g2099) & (g2794) & (!g2856) & (!g2857) & (!sk[38]) & (g2862)) + ((g2099) & (g2794) & (!g2856) & (g2857) & (!sk[38]) & (!g2862)) + ((g2099) & (g2794) & (!g2856) & (g2857) & (!sk[38]) & (g2862)) + ((g2099) & (g2794) & (g2856) & (!g2857) & (!sk[38]) & (!g2862)) + ((g2099) & (g2794) & (g2856) & (!g2857) & (!sk[38]) & (g2862)) + ((g2099) & (g2794) & (g2856) & (g2857) & (!sk[38]) & (!g2862)) + ((g2099) & (g2794) & (g2856) & (g2857) & (!sk[38]) & (g2862)) + ((g2099) & (g2794) & (g2856) & (g2857) & (sk[38]) & (g2862)));
	assign g2864 = (((!sk[39]) & (!g2115) & (!g2312) & (!g2850) & (g2853) & (!g2863)) + ((!sk[39]) & (!g2115) & (!g2312) & (!g2850) & (g2853) & (g2863)) + ((!sk[39]) & (!g2115) & (!g2312) & (g2850) & (!g2853) & (!g2863)) + ((!sk[39]) & (!g2115) & (!g2312) & (g2850) & (!g2853) & (g2863)) + ((!sk[39]) & (!g2115) & (!g2312) & (g2850) & (g2853) & (!g2863)) + ((!sk[39]) & (!g2115) & (!g2312) & (g2850) & (g2853) & (g2863)) + ((!sk[39]) & (!g2115) & (g2312) & (!g2850) & (g2853) & (!g2863)) + ((!sk[39]) & (!g2115) & (g2312) & (!g2850) & (g2853) & (g2863)) + ((!sk[39]) & (!g2115) & (g2312) & (g2850) & (!g2853) & (!g2863)) + ((!sk[39]) & (!g2115) & (g2312) & (g2850) & (!g2853) & (g2863)) + ((!sk[39]) & (!g2115) & (g2312) & (g2850) & (g2853) & (!g2863)) + ((!sk[39]) & (!g2115) & (g2312) & (g2850) & (g2853) & (g2863)) + ((!sk[39]) & (g2115) & (!g2312) & (!g2850) & (!g2853) & (!g2863)) + ((!sk[39]) & (g2115) & (!g2312) & (!g2850) & (!g2853) & (g2863)) + ((!sk[39]) & (g2115) & (!g2312) & (!g2850) & (g2853) & (!g2863)) + ((!sk[39]) & (g2115) & (!g2312) & (!g2850) & (g2853) & (g2863)) + ((!sk[39]) & (g2115) & (!g2312) & (g2850) & (!g2853) & (!g2863)) + ((!sk[39]) & (g2115) & (!g2312) & (g2850) & (!g2853) & (g2863)) + ((!sk[39]) & (g2115) & (!g2312) & (g2850) & (g2853) & (!g2863)) + ((!sk[39]) & (g2115) & (!g2312) & (g2850) & (g2853) & (g2863)) + ((!sk[39]) & (g2115) & (g2312) & (!g2850) & (!g2853) & (!g2863)) + ((!sk[39]) & (g2115) & (g2312) & (!g2850) & (!g2853) & (g2863)) + ((!sk[39]) & (g2115) & (g2312) & (!g2850) & (g2853) & (!g2863)) + ((!sk[39]) & (g2115) & (g2312) & (!g2850) & (g2853) & (g2863)) + ((!sk[39]) & (g2115) & (g2312) & (g2850) & (!g2853) & (!g2863)) + ((!sk[39]) & (g2115) & (g2312) & (g2850) & (!g2853) & (g2863)) + ((!sk[39]) & (g2115) & (g2312) & (g2850) & (g2853) & (!g2863)) + ((!sk[39]) & (g2115) & (g2312) & (g2850) & (g2853) & (g2863)) + ((sk[39]) & (!g2115) & (!g2312) & (g2850) & (g2853) & (g2863)) + ((sk[39]) & (g2115) & (g2312) & (g2850) & (g2853) & (g2863)));
	assign g2865 = (((!g110) & (!g106) & (!g678) & (!sk[40]) & (g2847) & (!g2864)) + ((!g110) & (!g106) & (!g678) & (!sk[40]) & (g2847) & (g2864)) + ((!g110) & (!g106) & (g678) & (!sk[40]) & (!g2847) & (!g2864)) + ((!g110) & (!g106) & (g678) & (!sk[40]) & (!g2847) & (g2864)) + ((!g110) & (!g106) & (g678) & (!sk[40]) & (g2847) & (!g2864)) + ((!g110) & (!g106) & (g678) & (!sk[40]) & (g2847) & (g2864)) + ((!g110) & (g106) & (!g678) & (!sk[40]) & (g2847) & (!g2864)) + ((!g110) & (g106) & (!g678) & (!sk[40]) & (g2847) & (g2864)) + ((!g110) & (g106) & (g678) & (!sk[40]) & (!g2847) & (!g2864)) + ((!g110) & (g106) & (g678) & (!sk[40]) & (!g2847) & (g2864)) + ((!g110) & (g106) & (g678) & (!sk[40]) & (g2847) & (!g2864)) + ((!g110) & (g106) & (g678) & (!sk[40]) & (g2847) & (g2864)) + ((g110) & (!g106) & (!g678) & (!sk[40]) & (!g2847) & (!g2864)) + ((g110) & (!g106) & (!g678) & (!sk[40]) & (!g2847) & (g2864)) + ((g110) & (!g106) & (!g678) & (!sk[40]) & (g2847) & (!g2864)) + ((g110) & (!g106) & (!g678) & (!sk[40]) & (g2847) & (g2864)) + ((g110) & (!g106) & (g678) & (!sk[40]) & (!g2847) & (!g2864)) + ((g110) & (!g106) & (g678) & (!sk[40]) & (!g2847) & (g2864)) + ((g110) & (!g106) & (g678) & (!sk[40]) & (g2847) & (!g2864)) + ((g110) & (!g106) & (g678) & (!sk[40]) & (g2847) & (g2864)) + ((g110) & (g106) & (!g678) & (!sk[40]) & (!g2847) & (!g2864)) + ((g110) & (g106) & (!g678) & (!sk[40]) & (!g2847) & (g2864)) + ((g110) & (g106) & (!g678) & (!sk[40]) & (g2847) & (!g2864)) + ((g110) & (g106) & (!g678) & (!sk[40]) & (g2847) & (g2864)) + ((g110) & (g106) & (!g678) & (sk[40]) & (g2847) & (!g2864)) + ((g110) & (g106) & (g678) & (!sk[40]) & (!g2847) & (!g2864)) + ((g110) & (g106) & (g678) & (!sk[40]) & (!g2847) & (g2864)) + ((g110) & (g106) & (g678) & (!sk[40]) & (g2847) & (!g2864)) + ((g110) & (g106) & (g678) & (!sk[40]) & (g2847) & (g2864)) + ((g110) & (g106) & (g678) & (sk[40]) & (g2847) & (!g2864)) + ((g110) & (g106) & (g678) & (sk[40]) & (g2847) & (g2864)));
	assign g2866 = (((!g108) & (g109) & (!sk[41]) & (!g2846)) + ((!g108) & (g109) & (!sk[41]) & (g2846)) + ((g108) & (!g109) & (!sk[41]) & (!g2846)) + ((g108) & (!g109) & (!sk[41]) & (g2846)) + ((g108) & (!g109) & (sk[41]) & (g2846)) + ((g108) & (g109) & (!sk[41]) & (!g2846)) + ((g108) & (g109) & (!sk[41]) & (g2846)));
	assign g2867 = (((!g110) & (!sk[42]) & (g106) & (!g2866)) + ((!g110) & (!sk[42]) & (g106) & (g2866)) + ((g110) & (!sk[42]) & (!g106) & (!g2866)) + ((g110) & (!sk[42]) & (!g106) & (g2866)) + ((g110) & (!sk[42]) & (g106) & (!g2866)) + ((g110) & (!sk[42]) & (g106) & (g2866)) + ((g110) & (sk[42]) & (g106) & (g2866)));
	assign g2868 = (((!g2074) & (!g2071) & (!sk[43]) & (!g2070) & (g2104)) + ((!g2074) & (!g2071) & (!sk[43]) & (g2070) & (g2104)) + ((!g2074) & (g2071) & (!sk[43]) & (!g2070) & (!g2104)) + ((!g2074) & (g2071) & (!sk[43]) & (!g2070) & (g2104)) + ((!g2074) & (g2071) & (!sk[43]) & (g2070) & (!g2104)) + ((!g2074) & (g2071) & (!sk[43]) & (g2070) & (g2104)) + ((!g2074) & (g2071) & (sk[43]) & (!g2070) & (!g2104)) + ((g2074) & (!g2071) & (!sk[43]) & (!g2070) & (!g2104)) + ((g2074) & (!g2071) & (!sk[43]) & (!g2070) & (g2104)) + ((g2074) & (!g2071) & (!sk[43]) & (g2070) & (!g2104)) + ((g2074) & (!g2071) & (!sk[43]) & (g2070) & (g2104)) + ((g2074) & (!g2071) & (sk[43]) & (!g2070) & (!g2104)) + ((g2074) & (!g2071) & (sk[43]) & (g2070) & (!g2104)) + ((g2074) & (g2071) & (!sk[43]) & (!g2070) & (!g2104)) + ((g2074) & (g2071) & (!sk[43]) & (!g2070) & (g2104)) + ((g2074) & (g2071) & (!sk[43]) & (g2070) & (!g2104)) + ((g2074) & (g2071) & (!sk[43]) & (g2070) & (g2104)) + ((g2074) & (g2071) & (sk[43]) & (!g2070) & (!g2104)) + ((g2074) & (g2071) & (sk[43]) & (!g2070) & (g2104)) + ((g2074) & (g2071) & (sk[43]) & (g2070) & (!g2104)));
	assign g2869 = (((!g2076) & (!sk[44]) & (!g2077) & (!g2105) & (g2106) & (!g2868)) + ((!g2076) & (!sk[44]) & (!g2077) & (!g2105) & (g2106) & (g2868)) + ((!g2076) & (!sk[44]) & (!g2077) & (g2105) & (!g2106) & (!g2868)) + ((!g2076) & (!sk[44]) & (!g2077) & (g2105) & (!g2106) & (g2868)) + ((!g2076) & (!sk[44]) & (!g2077) & (g2105) & (g2106) & (!g2868)) + ((!g2076) & (!sk[44]) & (!g2077) & (g2105) & (g2106) & (g2868)) + ((!g2076) & (!sk[44]) & (g2077) & (!g2105) & (g2106) & (!g2868)) + ((!g2076) & (!sk[44]) & (g2077) & (!g2105) & (g2106) & (g2868)) + ((!g2076) & (!sk[44]) & (g2077) & (g2105) & (!g2106) & (!g2868)) + ((!g2076) & (!sk[44]) & (g2077) & (g2105) & (!g2106) & (g2868)) + ((!g2076) & (!sk[44]) & (g2077) & (g2105) & (g2106) & (!g2868)) + ((!g2076) & (!sk[44]) & (g2077) & (g2105) & (g2106) & (g2868)) + ((!g2076) & (sk[44]) & (!g2077) & (!g2105) & (!g2106) & (g2868)) + ((!g2076) & (sk[44]) & (g2077) & (!g2105) & (!g2106) & (!g2868)) + ((!g2076) & (sk[44]) & (g2077) & (!g2105) & (!g2106) & (g2868)) + ((!g2076) & (sk[44]) & (g2077) & (g2105) & (!g2106) & (g2868)) + ((g2076) & (!sk[44]) & (!g2077) & (!g2105) & (!g2106) & (!g2868)) + ((g2076) & (!sk[44]) & (!g2077) & (!g2105) & (!g2106) & (g2868)) + ((g2076) & (!sk[44]) & (!g2077) & (!g2105) & (g2106) & (!g2868)) + ((g2076) & (!sk[44]) & (!g2077) & (!g2105) & (g2106) & (g2868)) + ((g2076) & (!sk[44]) & (!g2077) & (g2105) & (!g2106) & (!g2868)) + ((g2076) & (!sk[44]) & (!g2077) & (g2105) & (!g2106) & (g2868)) + ((g2076) & (!sk[44]) & (!g2077) & (g2105) & (g2106) & (!g2868)) + ((g2076) & (!sk[44]) & (!g2077) & (g2105) & (g2106) & (g2868)) + ((g2076) & (!sk[44]) & (g2077) & (!g2105) & (!g2106) & (!g2868)) + ((g2076) & (!sk[44]) & (g2077) & (!g2105) & (!g2106) & (g2868)) + ((g2076) & (!sk[44]) & (g2077) & (!g2105) & (g2106) & (!g2868)) + ((g2076) & (!sk[44]) & (g2077) & (!g2105) & (g2106) & (g2868)) + ((g2076) & (!sk[44]) & (g2077) & (g2105) & (!g2106) & (!g2868)) + ((g2076) & (!sk[44]) & (g2077) & (g2105) & (!g2106) & (g2868)) + ((g2076) & (!sk[44]) & (g2077) & (g2105) & (g2106) & (!g2868)) + ((g2076) & (!sk[44]) & (g2077) & (g2105) & (g2106) & (g2868)) + ((g2076) & (sk[44]) & (!g2077) & (!g2105) & (!g2106) & (!g2868)) + ((g2076) & (sk[44]) & (!g2077) & (!g2105) & (!g2106) & (g2868)) + ((g2076) & (sk[44]) & (!g2077) & (!g2105) & (g2106) & (g2868)) + ((g2076) & (sk[44]) & (!g2077) & (g2105) & (!g2106) & (!g2868)) + ((g2076) & (sk[44]) & (!g2077) & (g2105) & (!g2106) & (g2868)) + ((g2076) & (sk[44]) & (g2077) & (!g2105) & (!g2106) & (!g2868)) + ((g2076) & (sk[44]) & (g2077) & (!g2105) & (!g2106) & (g2868)) + ((g2076) & (sk[44]) & (g2077) & (!g2105) & (g2106) & (!g2868)) + ((g2076) & (sk[44]) & (g2077) & (!g2105) & (g2106) & (g2868)) + ((g2076) & (sk[44]) & (g2077) & (g2105) & (!g2106) & (!g2868)) + ((g2076) & (sk[44]) & (g2077) & (g2105) & (!g2106) & (g2868)) + ((g2076) & (sk[44]) & (g2077) & (g2105) & (g2106) & (g2868)));
	assign g2870 = (((!g2073) & (!sk[45]) & (!g2113) & (!g2114) & (g2289) & (!g2869)) + ((!g2073) & (!sk[45]) & (!g2113) & (!g2114) & (g2289) & (g2869)) + ((!g2073) & (!sk[45]) & (!g2113) & (g2114) & (!g2289) & (!g2869)) + ((!g2073) & (!sk[45]) & (!g2113) & (g2114) & (!g2289) & (g2869)) + ((!g2073) & (!sk[45]) & (!g2113) & (g2114) & (g2289) & (!g2869)) + ((!g2073) & (!sk[45]) & (!g2113) & (g2114) & (g2289) & (g2869)) + ((!g2073) & (!sk[45]) & (g2113) & (!g2114) & (g2289) & (!g2869)) + ((!g2073) & (!sk[45]) & (g2113) & (!g2114) & (g2289) & (g2869)) + ((!g2073) & (!sk[45]) & (g2113) & (g2114) & (!g2289) & (!g2869)) + ((!g2073) & (!sk[45]) & (g2113) & (g2114) & (!g2289) & (g2869)) + ((!g2073) & (!sk[45]) & (g2113) & (g2114) & (g2289) & (!g2869)) + ((!g2073) & (!sk[45]) & (g2113) & (g2114) & (g2289) & (g2869)) + ((!g2073) & (sk[45]) & (!g2113) & (!g2114) & (!g2289) & (g2869)) + ((!g2073) & (sk[45]) & (!g2113) & (!g2114) & (g2289) & (!g2869)) + ((!g2073) & (sk[45]) & (!g2113) & (!g2114) & (g2289) & (g2869)) + ((!g2073) & (sk[45]) & (!g2113) & (g2114) & (g2289) & (g2869)) + ((!g2073) & (sk[45]) & (g2113) & (!g2114) & (g2289) & (!g2869)) + ((!g2073) & (sk[45]) & (g2113) & (!g2114) & (g2289) & (g2869)) + ((g2073) & (!sk[45]) & (!g2113) & (!g2114) & (!g2289) & (!g2869)) + ((g2073) & (!sk[45]) & (!g2113) & (!g2114) & (!g2289) & (g2869)) + ((g2073) & (!sk[45]) & (!g2113) & (!g2114) & (g2289) & (!g2869)) + ((g2073) & (!sk[45]) & (!g2113) & (!g2114) & (g2289) & (g2869)) + ((g2073) & (!sk[45]) & (!g2113) & (g2114) & (!g2289) & (!g2869)) + ((g2073) & (!sk[45]) & (!g2113) & (g2114) & (!g2289) & (g2869)) + ((g2073) & (!sk[45]) & (!g2113) & (g2114) & (g2289) & (!g2869)) + ((g2073) & (!sk[45]) & (!g2113) & (g2114) & (g2289) & (g2869)) + ((g2073) & (!sk[45]) & (g2113) & (!g2114) & (!g2289) & (!g2869)) + ((g2073) & (!sk[45]) & (g2113) & (!g2114) & (!g2289) & (g2869)) + ((g2073) & (!sk[45]) & (g2113) & (!g2114) & (g2289) & (!g2869)) + ((g2073) & (!sk[45]) & (g2113) & (!g2114) & (g2289) & (g2869)) + ((g2073) & (!sk[45]) & (g2113) & (g2114) & (!g2289) & (!g2869)) + ((g2073) & (!sk[45]) & (g2113) & (g2114) & (!g2289) & (g2869)) + ((g2073) & (!sk[45]) & (g2113) & (g2114) & (g2289) & (!g2869)) + ((g2073) & (!sk[45]) & (g2113) & (g2114) & (g2289) & (g2869)) + ((g2073) & (sk[45]) & (!g2113) & (!g2114) & (!g2289) & (!g2869)) + ((g2073) & (sk[45]) & (!g2113) & (!g2114) & (!g2289) & (g2869)) + ((g2073) & (sk[45]) & (!g2113) & (!g2114) & (g2289) & (!g2869)) + ((g2073) & (sk[45]) & (!g2113) & (!g2114) & (g2289) & (g2869)) + ((g2073) & (sk[45]) & (!g2113) & (g2114) & (g2289) & (!g2869)) + ((g2073) & (sk[45]) & (!g2113) & (g2114) & (g2289) & (g2869)) + ((g2073) & (sk[45]) & (g2113) & (!g2114) & (!g2289) & (g2869)) + ((g2073) & (sk[45]) & (g2113) & (!g2114) & (g2289) & (!g2869)) + ((g2073) & (sk[45]) & (g2113) & (!g2114) & (g2289) & (g2869)) + ((g2073) & (sk[45]) & (g2113) & (g2114) & (g2289) & (g2869)));
	assign g2871 = (((!g2109) & (!g2110) & (!g2111) & (!g2391) & (!g2418) & (g2439)) + ((!g2109) & (!g2110) & (!g2111) & (!g2391) & (g2418) & (!g2439)) + ((!g2109) & (!g2110) & (!g2111) & (!g2391) & (g2418) & (g2439)) + ((!g2109) & (!g2110) & (!g2111) & (g2391) & (!g2418) & (!g2439)) + ((!g2109) & (!g2110) & (!g2111) & (g2391) & (!g2418) & (g2439)) + ((!g2109) & (!g2110) & (!g2111) & (g2391) & (g2418) & (!g2439)) + ((!g2109) & (!g2110) & (!g2111) & (g2391) & (g2418) & (g2439)) + ((!g2109) & (!g2110) & (g2111) & (!g2391) & (g2418) & (g2439)) + ((!g2109) & (!g2110) & (g2111) & (g2391) & (!g2418) & (g2439)) + ((!g2109) & (!g2110) & (g2111) & (g2391) & (g2418) & (g2439)) + ((!g2109) & (g2110) & (!g2111) & (!g2391) & (!g2418) & (g2439)) + ((!g2109) & (g2110) & (!g2111) & (!g2391) & (g2418) & (g2439)) + ((!g2109) & (g2110) & (!g2111) & (g2391) & (!g2418) & (g2439)) + ((!g2109) & (g2110) & (!g2111) & (g2391) & (g2418) & (!g2439)) + ((!g2109) & (g2110) & (!g2111) & (g2391) & (g2418) & (g2439)) + ((!g2109) & (g2110) & (g2111) & (g2391) & (g2418) & (g2439)) + ((g2109) & (!g2110) & (!g2111) & (!g2391) & (!g2418) & (g2439)) + ((g2109) & (!g2110) & (!g2111) & (!g2391) & (g2418) & (!g2439)) + ((g2109) & (!g2110) & (!g2111) & (!g2391) & (g2418) & (g2439)) + ((g2109) & (!g2110) & (!g2111) & (g2391) & (!g2418) & (g2439)) + ((g2109) & (!g2110) & (!g2111) & (g2391) & (g2418) & (!g2439)) + ((g2109) & (!g2110) & (!g2111) & (g2391) & (g2418) & (g2439)) + ((g2109) & (!g2110) & (g2111) & (!g2391) & (g2418) & (g2439)) + ((g2109) & (!g2110) & (g2111) & (g2391) & (g2418) & (g2439)) + ((g2109) & (g2110) & (!g2111) & (!g2391) & (!g2418) & (g2439)) + ((g2109) & (g2110) & (!g2111) & (!g2391) & (g2418) & (g2439)) + ((g2109) & (g2110) & (!g2111) & (g2391) & (!g2418) & (g2439)) + ((g2109) & (g2110) & (!g2111) & (g2391) & (g2418) & (g2439)));
	assign g2872 = (((!g2108) & (!g2116) & (!g2340) & (!g2365) & (!g2852) & (!g2871)) + ((!g2108) & (!g2116) & (!g2340) & (!g2365) & (g2852) & (!g2871)) + ((!g2108) & (!g2116) & (!g2340) & (g2365) & (!g2852) & (!g2871)) + ((!g2108) & (!g2116) & (g2340) & (!g2365) & (!g2852) & (!g2871)) + ((!g2108) & (!g2116) & (g2340) & (g2365) & (!g2852) & (!g2871)) + ((!g2108) & (g2116) & (!g2340) & (!g2365) & (!g2852) & (!g2871)) + ((!g2108) & (g2116) & (!g2340) & (!g2365) & (g2852) & (!g2871)) + ((!g2108) & (g2116) & (!g2340) & (g2365) & (!g2852) & (!g2871)) + ((!g2108) & (g2116) & (g2340) & (!g2365) & (!g2852) & (!g2871)) + ((!g2108) & (g2116) & (g2340) & (!g2365) & (g2852) & (!g2871)) + ((!g2108) & (g2116) & (g2340) & (g2365) & (!g2852) & (!g2871)) + ((g2108) & (!g2116) & (!g2340) & (!g2365) & (!g2852) & (!g2871)) + ((g2108) & (!g2116) & (!g2340) & (!g2365) & (g2852) & (!g2871)) + ((g2108) & (!g2116) & (!g2340) & (g2365) & (!g2852) & (!g2871)) + ((g2108) & (!g2116) & (!g2340) & (g2365) & (g2852) & (!g2871)) + ((g2108) & (!g2116) & (g2340) & (!g2365) & (!g2852) & (!g2871)) + ((g2108) & (!g2116) & (g2340) & (!g2365) & (g2852) & (!g2871)) + ((g2108) & (!g2116) & (g2340) & (g2365) & (!g2852) & (!g2871)) + ((g2108) & (g2116) & (!g2340) & (!g2365) & (!g2852) & (!g2871)) + ((g2108) & (g2116) & (!g2340) & (!g2365) & (g2852) & (!g2871)) + ((g2108) & (g2116) & (!g2340) & (g2365) & (!g2852) & (!g2871)) + ((g2108) & (g2116) & (!g2340) & (g2365) & (g2852) & (!g2871)) + ((g2108) & (g2116) & (g2340) & (!g2365) & (!g2852) & (!g2871)) + ((g2108) & (g2116) & (g2340) & (!g2365) & (g2852) & (!g2871)) + ((g2108) & (g2116) & (g2340) & (g2365) & (!g2852) & (!g2871)) + ((g2108) & (g2116) & (g2340) & (g2365) & (g2852) & (!g2871)));
	assign g2873 = (((!g2115) & (!g2312) & (!g2853) & (!sk[48]) & (g2870) & (!g2872)) + ((!g2115) & (!g2312) & (!g2853) & (!sk[48]) & (g2870) & (g2872)) + ((!g2115) & (!g2312) & (!g2853) & (sk[48]) & (!g2870) & (g2872)) + ((!g2115) & (!g2312) & (!g2853) & (sk[48]) & (g2870) & (g2872)) + ((!g2115) & (!g2312) & (g2853) & (!sk[48]) & (!g2870) & (!g2872)) + ((!g2115) & (!g2312) & (g2853) & (!sk[48]) & (!g2870) & (g2872)) + ((!g2115) & (!g2312) & (g2853) & (!sk[48]) & (g2870) & (!g2872)) + ((!g2115) & (!g2312) & (g2853) & (!sk[48]) & (g2870) & (g2872)) + ((!g2115) & (!g2312) & (g2853) & (sk[48]) & (!g2870) & (g2872)) + ((!g2115) & (g2312) & (!g2853) & (!sk[48]) & (g2870) & (!g2872)) + ((!g2115) & (g2312) & (!g2853) & (!sk[48]) & (g2870) & (g2872)) + ((!g2115) & (g2312) & (!g2853) & (sk[48]) & (!g2870) & (g2872)) + ((!g2115) & (g2312) & (!g2853) & (sk[48]) & (g2870) & (g2872)) + ((!g2115) & (g2312) & (g2853) & (!sk[48]) & (!g2870) & (!g2872)) + ((!g2115) & (g2312) & (g2853) & (!sk[48]) & (!g2870) & (g2872)) + ((!g2115) & (g2312) & (g2853) & (!sk[48]) & (g2870) & (!g2872)) + ((!g2115) & (g2312) & (g2853) & (!sk[48]) & (g2870) & (g2872)) + ((g2115) & (!g2312) & (!g2853) & (!sk[48]) & (!g2870) & (!g2872)) + ((g2115) & (!g2312) & (!g2853) & (!sk[48]) & (!g2870) & (g2872)) + ((g2115) & (!g2312) & (!g2853) & (!sk[48]) & (g2870) & (!g2872)) + ((g2115) & (!g2312) & (!g2853) & (!sk[48]) & (g2870) & (g2872)) + ((g2115) & (!g2312) & (!g2853) & (sk[48]) & (!g2870) & (g2872)) + ((g2115) & (!g2312) & (!g2853) & (sk[48]) & (g2870) & (g2872)) + ((g2115) & (!g2312) & (g2853) & (!sk[48]) & (!g2870) & (!g2872)) + ((g2115) & (!g2312) & (g2853) & (!sk[48]) & (!g2870) & (g2872)) + ((g2115) & (!g2312) & (g2853) & (!sk[48]) & (g2870) & (!g2872)) + ((g2115) & (!g2312) & (g2853) & (!sk[48]) & (g2870) & (g2872)) + ((g2115) & (!g2312) & (g2853) & (sk[48]) & (!g2870) & (g2872)) + ((g2115) & (!g2312) & (g2853) & (sk[48]) & (g2870) & (g2872)) + ((g2115) & (g2312) & (!g2853) & (!sk[48]) & (!g2870) & (!g2872)) + ((g2115) & (g2312) & (!g2853) & (!sk[48]) & (!g2870) & (g2872)) + ((g2115) & (g2312) & (!g2853) & (!sk[48]) & (g2870) & (!g2872)) + ((g2115) & (g2312) & (!g2853) & (!sk[48]) & (g2870) & (g2872)) + ((g2115) & (g2312) & (!g2853) & (sk[48]) & (!g2870) & (g2872)) + ((g2115) & (g2312) & (!g2853) & (sk[48]) & (g2870) & (g2872)) + ((g2115) & (g2312) & (g2853) & (!sk[48]) & (!g2870) & (!g2872)) + ((g2115) & (g2312) & (g2853) & (!sk[48]) & (!g2870) & (g2872)) + ((g2115) & (g2312) & (g2853) & (!sk[48]) & (g2870) & (!g2872)) + ((g2115) & (g2312) & (g2853) & (!sk[48]) & (g2870) & (g2872)) + ((g2115) & (g2312) & (g2853) & (sk[48]) & (!g2870) & (g2872)));
	assign g2874 = (((!g2119) & (!sk[49]) & (!g2120) & (!g2482) & (g2507)) + ((!g2119) & (!sk[49]) & (!g2120) & (g2482) & (g2507)) + ((!g2119) & (!sk[49]) & (g2120) & (!g2482) & (!g2507)) + ((!g2119) & (!sk[49]) & (g2120) & (!g2482) & (g2507)) + ((!g2119) & (!sk[49]) & (g2120) & (g2482) & (!g2507)) + ((!g2119) & (!sk[49]) & (g2120) & (g2482) & (g2507)) + ((!g2119) & (sk[49]) & (!g2120) & (!g2482) & (g2507)) + ((!g2119) & (sk[49]) & (!g2120) & (g2482) & (!g2507)) + ((!g2119) & (sk[49]) & (!g2120) & (g2482) & (g2507)) + ((!g2119) & (sk[49]) & (g2120) & (g2482) & (g2507)) + ((g2119) & (!sk[49]) & (!g2120) & (!g2482) & (!g2507)) + ((g2119) & (!sk[49]) & (!g2120) & (!g2482) & (g2507)) + ((g2119) & (!sk[49]) & (!g2120) & (g2482) & (!g2507)) + ((g2119) & (!sk[49]) & (!g2120) & (g2482) & (g2507)) + ((g2119) & (!sk[49]) & (g2120) & (!g2482) & (!g2507)) + ((g2119) & (!sk[49]) & (g2120) & (!g2482) & (g2507)) + ((g2119) & (!sk[49]) & (g2120) & (g2482) & (!g2507)) + ((g2119) & (!sk[49]) & (g2120) & (g2482) & (g2507)) + ((g2119) & (sk[49]) & (!g2120) & (!g2482) & (g2507)) + ((g2119) & (sk[49]) & (!g2120) & (g2482) & (g2507)));
	assign g2875 = (((!g2118) & (!sk[50]) & (!g2457) & (!g2858) & (g2873) & (!g2874)) + ((!g2118) & (!sk[50]) & (!g2457) & (!g2858) & (g2873) & (g2874)) + ((!g2118) & (!sk[50]) & (!g2457) & (g2858) & (!g2873) & (!g2874)) + ((!g2118) & (!sk[50]) & (!g2457) & (g2858) & (!g2873) & (g2874)) + ((!g2118) & (!sk[50]) & (!g2457) & (g2858) & (g2873) & (!g2874)) + ((!g2118) & (!sk[50]) & (!g2457) & (g2858) & (g2873) & (g2874)) + ((!g2118) & (!sk[50]) & (g2457) & (!g2858) & (g2873) & (!g2874)) + ((!g2118) & (!sk[50]) & (g2457) & (!g2858) & (g2873) & (g2874)) + ((!g2118) & (!sk[50]) & (g2457) & (g2858) & (!g2873) & (!g2874)) + ((!g2118) & (!sk[50]) & (g2457) & (g2858) & (!g2873) & (g2874)) + ((!g2118) & (!sk[50]) & (g2457) & (g2858) & (g2873) & (!g2874)) + ((!g2118) & (!sk[50]) & (g2457) & (g2858) & (g2873) & (g2874)) + ((!g2118) & (sk[50]) & (!g2457) & (!g2858) & (!g2873) & (!g2874)) + ((!g2118) & (sk[50]) & (!g2457) & (!g2858) & (g2873) & (!g2874)) + ((!g2118) & (sk[50]) & (!g2457) & (g2858) & (g2873) & (!g2874)) + ((!g2118) & (sk[50]) & (g2457) & (!g2858) & (!g2873) & (!g2874)) + ((!g2118) & (sk[50]) & (g2457) & (!g2858) & (g2873) & (!g2874)) + ((g2118) & (!sk[50]) & (!g2457) & (!g2858) & (!g2873) & (!g2874)) + ((g2118) & (!sk[50]) & (!g2457) & (!g2858) & (!g2873) & (g2874)) + ((g2118) & (!sk[50]) & (!g2457) & (!g2858) & (g2873) & (!g2874)) + ((g2118) & (!sk[50]) & (!g2457) & (!g2858) & (g2873) & (g2874)) + ((g2118) & (!sk[50]) & (!g2457) & (g2858) & (!g2873) & (!g2874)) + ((g2118) & (!sk[50]) & (!g2457) & (g2858) & (!g2873) & (g2874)) + ((g2118) & (!sk[50]) & (!g2457) & (g2858) & (g2873) & (!g2874)) + ((g2118) & (!sk[50]) & (!g2457) & (g2858) & (g2873) & (g2874)) + ((g2118) & (!sk[50]) & (g2457) & (!g2858) & (!g2873) & (!g2874)) + ((g2118) & (!sk[50]) & (g2457) & (!g2858) & (!g2873) & (g2874)) + ((g2118) & (!sk[50]) & (g2457) & (!g2858) & (g2873) & (!g2874)) + ((g2118) & (!sk[50]) & (g2457) & (!g2858) & (g2873) & (g2874)) + ((g2118) & (!sk[50]) & (g2457) & (g2858) & (!g2873) & (!g2874)) + ((g2118) & (!sk[50]) & (g2457) & (g2858) & (!g2873) & (g2874)) + ((g2118) & (!sk[50]) & (g2457) & (g2858) & (g2873) & (!g2874)) + ((g2118) & (!sk[50]) & (g2457) & (g2858) & (g2873) & (g2874)) + ((g2118) & (sk[50]) & (!g2457) & (!g2858) & (!g2873) & (!g2874)) + ((g2118) & (sk[50]) & (!g2457) & (!g2858) & (g2873) & (!g2874)) + ((g2118) & (sk[50]) & (!g2457) & (g2858) & (!g2873) & (!g2874)) + ((g2118) & (sk[50]) & (!g2457) & (g2858) & (g2873) & (!g2874)) + ((g2118) & (sk[50]) & (g2457) & (!g2858) & (!g2873) & (!g2874)) + ((g2118) & (sk[50]) & (g2457) & (!g2858) & (g2873) & (!g2874)) + ((g2118) & (sk[50]) & (g2457) & (g2858) & (g2873) & (!g2874)));
	assign g2876 = (((!g2086) & (!g2093) & (!g2094) & (!g2608) & (!g2625) & (g2642)) + ((!g2086) & (!g2093) & (!g2094) & (!g2608) & (g2625) & (!g2642)) + ((!g2086) & (!g2093) & (!g2094) & (!g2608) & (g2625) & (g2642)) + ((!g2086) & (!g2093) & (!g2094) & (g2608) & (!g2625) & (!g2642)) + ((!g2086) & (!g2093) & (!g2094) & (g2608) & (!g2625) & (g2642)) + ((!g2086) & (!g2093) & (!g2094) & (g2608) & (g2625) & (!g2642)) + ((!g2086) & (!g2093) & (!g2094) & (g2608) & (g2625) & (g2642)) + ((!g2086) & (!g2093) & (g2094) & (!g2608) & (g2625) & (g2642)) + ((!g2086) & (!g2093) & (g2094) & (g2608) & (!g2625) & (g2642)) + ((!g2086) & (!g2093) & (g2094) & (g2608) & (g2625) & (g2642)) + ((!g2086) & (g2093) & (!g2094) & (!g2608) & (!g2625) & (g2642)) + ((!g2086) & (g2093) & (!g2094) & (!g2608) & (g2625) & (g2642)) + ((!g2086) & (g2093) & (!g2094) & (g2608) & (!g2625) & (g2642)) + ((!g2086) & (g2093) & (!g2094) & (g2608) & (g2625) & (!g2642)) + ((!g2086) & (g2093) & (!g2094) & (g2608) & (g2625) & (g2642)) + ((!g2086) & (g2093) & (g2094) & (g2608) & (g2625) & (g2642)) + ((g2086) & (!g2093) & (!g2094) & (!g2608) & (!g2625) & (g2642)) + ((g2086) & (!g2093) & (!g2094) & (!g2608) & (g2625) & (!g2642)) + ((g2086) & (!g2093) & (!g2094) & (!g2608) & (g2625) & (g2642)) + ((g2086) & (!g2093) & (!g2094) & (g2608) & (!g2625) & (g2642)) + ((g2086) & (!g2093) & (!g2094) & (g2608) & (g2625) & (!g2642)) + ((g2086) & (!g2093) & (!g2094) & (g2608) & (g2625) & (g2642)) + ((g2086) & (!g2093) & (g2094) & (!g2608) & (g2625) & (g2642)) + ((g2086) & (!g2093) & (g2094) & (g2608) & (g2625) & (g2642)) + ((g2086) & (g2093) & (!g2094) & (!g2608) & (!g2625) & (g2642)) + ((g2086) & (g2093) & (!g2094) & (!g2608) & (g2625) & (g2642)) + ((g2086) & (g2093) & (!g2094) & (g2608) & (!g2625) & (g2642)) + ((g2086) & (g2093) & (!g2094) & (g2608) & (g2625) & (g2642)));
	assign g2877 = (((!g2084) & (!g2085) & (!g2570) & (!g2590) & (!g2854) & (!g2876)) + ((!g2084) & (!g2085) & (!g2570) & (!g2590) & (g2854) & (!g2876)) + ((!g2084) & (!g2085) & (!g2570) & (g2590) & (!g2854) & (!g2876)) + ((!g2084) & (!g2085) & (g2570) & (!g2590) & (!g2854) & (!g2876)) + ((!g2084) & (!g2085) & (g2570) & (g2590) & (!g2854) & (!g2876)) + ((!g2084) & (g2085) & (!g2570) & (!g2590) & (!g2854) & (!g2876)) + ((!g2084) & (g2085) & (!g2570) & (!g2590) & (g2854) & (!g2876)) + ((!g2084) & (g2085) & (!g2570) & (g2590) & (!g2854) & (!g2876)) + ((!g2084) & (g2085) & (!g2570) & (g2590) & (g2854) & (!g2876)) + ((!g2084) & (g2085) & (g2570) & (!g2590) & (!g2854) & (!g2876)) + ((!g2084) & (g2085) & (g2570) & (!g2590) & (g2854) & (!g2876)) + ((!g2084) & (g2085) & (g2570) & (g2590) & (!g2854) & (!g2876)) + ((g2084) & (!g2085) & (!g2570) & (!g2590) & (!g2854) & (!g2876)) + ((g2084) & (!g2085) & (!g2570) & (!g2590) & (g2854) & (!g2876)) + ((g2084) & (!g2085) & (!g2570) & (g2590) & (!g2854) & (!g2876)) + ((g2084) & (!g2085) & (g2570) & (!g2590) & (!g2854) & (!g2876)) + ((g2084) & (!g2085) & (g2570) & (!g2590) & (g2854) & (!g2876)) + ((g2084) & (!g2085) & (g2570) & (g2590) & (!g2854) & (!g2876)) + ((g2084) & (g2085) & (!g2570) & (!g2590) & (!g2854) & (!g2876)) + ((g2084) & (g2085) & (!g2570) & (!g2590) & (g2854) & (!g2876)) + ((g2084) & (g2085) & (!g2570) & (g2590) & (!g2854) & (!g2876)) + ((g2084) & (g2085) & (!g2570) & (g2590) & (g2854) & (!g2876)) + ((g2084) & (g2085) & (g2570) & (!g2590) & (!g2854) & (!g2876)) + ((g2084) & (g2085) & (g2570) & (!g2590) & (g2854) & (!g2876)) + ((g2084) & (g2085) & (g2570) & (g2590) & (!g2854) & (!g2876)) + ((g2084) & (g2085) & (g2570) & (g2590) & (g2854) & (!g2876)));
	assign g2878 = (((!g2083) & (!g2121) & (!g2529) & (!sk[53]) & (g2551) & (!g2855)) + ((!g2083) & (!g2121) & (!g2529) & (!sk[53]) & (g2551) & (g2855)) + ((!g2083) & (!g2121) & (!g2529) & (sk[53]) & (g2551) & (g2855)) + ((!g2083) & (!g2121) & (g2529) & (!sk[53]) & (!g2551) & (!g2855)) + ((!g2083) & (!g2121) & (g2529) & (!sk[53]) & (!g2551) & (g2855)) + ((!g2083) & (!g2121) & (g2529) & (!sk[53]) & (g2551) & (!g2855)) + ((!g2083) & (!g2121) & (g2529) & (!sk[53]) & (g2551) & (g2855)) + ((!g2083) & (!g2121) & (g2529) & (sk[53]) & (!g2551) & (g2855)) + ((!g2083) & (!g2121) & (g2529) & (sk[53]) & (g2551) & (g2855)) + ((!g2083) & (g2121) & (!g2529) & (!sk[53]) & (g2551) & (!g2855)) + ((!g2083) & (g2121) & (!g2529) & (!sk[53]) & (g2551) & (g2855)) + ((!g2083) & (g2121) & (!g2529) & (sk[53]) & (g2551) & (g2855)) + ((!g2083) & (g2121) & (g2529) & (!sk[53]) & (!g2551) & (!g2855)) + ((!g2083) & (g2121) & (g2529) & (!sk[53]) & (!g2551) & (g2855)) + ((!g2083) & (g2121) & (g2529) & (!sk[53]) & (g2551) & (!g2855)) + ((!g2083) & (g2121) & (g2529) & (!sk[53]) & (g2551) & (g2855)) + ((!g2083) & (g2121) & (g2529) & (sk[53]) & (g2551) & (g2855)) + ((g2083) & (!g2121) & (!g2529) & (!sk[53]) & (!g2551) & (!g2855)) + ((g2083) & (!g2121) & (!g2529) & (!sk[53]) & (!g2551) & (g2855)) + ((g2083) & (!g2121) & (!g2529) & (!sk[53]) & (g2551) & (!g2855)) + ((g2083) & (!g2121) & (!g2529) & (!sk[53]) & (g2551) & (g2855)) + ((g2083) & (!g2121) & (g2529) & (!sk[53]) & (!g2551) & (!g2855)) + ((g2083) & (!g2121) & (g2529) & (!sk[53]) & (!g2551) & (g2855)) + ((g2083) & (!g2121) & (g2529) & (!sk[53]) & (g2551) & (!g2855)) + ((g2083) & (!g2121) & (g2529) & (!sk[53]) & (g2551) & (g2855)) + ((g2083) & (!g2121) & (g2529) & (sk[53]) & (g2551) & (g2855)) + ((g2083) & (g2121) & (!g2529) & (!sk[53]) & (!g2551) & (!g2855)) + ((g2083) & (g2121) & (!g2529) & (!sk[53]) & (!g2551) & (g2855)) + ((g2083) & (g2121) & (!g2529) & (!sk[53]) & (g2551) & (!g2855)) + ((g2083) & (g2121) & (!g2529) & (!sk[53]) & (g2551) & (g2855)) + ((g2083) & (g2121) & (g2529) & (!sk[53]) & (!g2551) & (!g2855)) + ((g2083) & (g2121) & (g2529) & (!sk[53]) & (!g2551) & (g2855)) + ((g2083) & (g2121) & (g2529) & (!sk[53]) & (g2551) & (!g2855)) + ((g2083) & (g2121) & (g2529) & (!sk[53]) & (g2551) & (g2855)));
	assign g2879 = (((!g2856) & (!g2875) & (!g2877) & (!sk[54]) & (g2878)) + ((!g2856) & (!g2875) & (g2877) & (!sk[54]) & (g2878)) + ((!g2856) & (!g2875) & (g2877) & (sk[54]) & (!g2878)) + ((!g2856) & (g2875) & (!g2877) & (!sk[54]) & (!g2878)) + ((!g2856) & (g2875) & (!g2877) & (!sk[54]) & (g2878)) + ((!g2856) & (g2875) & (g2877) & (!sk[54]) & (!g2878)) + ((!g2856) & (g2875) & (g2877) & (!sk[54]) & (g2878)) + ((!g2856) & (g2875) & (g2877) & (sk[54]) & (!g2878)) + ((g2856) & (!g2875) & (!g2877) & (!sk[54]) & (!g2878)) + ((g2856) & (!g2875) & (!g2877) & (!sk[54]) & (g2878)) + ((g2856) & (!g2875) & (g2877) & (!sk[54]) & (!g2878)) + ((g2856) & (!g2875) & (g2877) & (!sk[54]) & (g2878)) + ((g2856) & (g2875) & (!g2877) & (!sk[54]) & (!g2878)) + ((g2856) & (g2875) & (!g2877) & (!sk[54]) & (g2878)) + ((g2856) & (g2875) & (g2877) & (!sk[54]) & (!g2878)) + ((g2856) & (g2875) & (g2877) & (!sk[54]) & (g2878)) + ((g2856) & (g2875) & (g2877) & (sk[54]) & (!g2878)));
	assign g2880 = (((!g2090) & (!g2091) & (!g2098) & (!g2734) & (!g2751) & (g2771)) + ((!g2090) & (!g2091) & (!g2098) & (!g2734) & (g2751) & (!g2771)) + ((!g2090) & (!g2091) & (!g2098) & (!g2734) & (g2751) & (g2771)) + ((!g2090) & (!g2091) & (!g2098) & (g2734) & (!g2751) & (!g2771)) + ((!g2090) & (!g2091) & (!g2098) & (g2734) & (!g2751) & (g2771)) + ((!g2090) & (!g2091) & (!g2098) & (g2734) & (g2751) & (!g2771)) + ((!g2090) & (!g2091) & (!g2098) & (g2734) & (g2751) & (g2771)) + ((!g2090) & (!g2091) & (g2098) & (!g2734) & (g2751) & (g2771)) + ((!g2090) & (!g2091) & (g2098) & (g2734) & (!g2751) & (g2771)) + ((!g2090) & (!g2091) & (g2098) & (g2734) & (g2751) & (g2771)) + ((!g2090) & (g2091) & (!g2098) & (!g2734) & (!g2751) & (g2771)) + ((!g2090) & (g2091) & (!g2098) & (!g2734) & (g2751) & (g2771)) + ((!g2090) & (g2091) & (!g2098) & (g2734) & (!g2751) & (g2771)) + ((!g2090) & (g2091) & (!g2098) & (g2734) & (g2751) & (!g2771)) + ((!g2090) & (g2091) & (!g2098) & (g2734) & (g2751) & (g2771)) + ((!g2090) & (g2091) & (g2098) & (g2734) & (g2751) & (g2771)) + ((g2090) & (!g2091) & (!g2098) & (!g2734) & (!g2751) & (g2771)) + ((g2090) & (!g2091) & (!g2098) & (!g2734) & (g2751) & (!g2771)) + ((g2090) & (!g2091) & (!g2098) & (!g2734) & (g2751) & (g2771)) + ((g2090) & (!g2091) & (!g2098) & (g2734) & (!g2751) & (g2771)) + ((g2090) & (!g2091) & (!g2098) & (g2734) & (g2751) & (!g2771)) + ((g2090) & (!g2091) & (!g2098) & (g2734) & (g2751) & (g2771)) + ((g2090) & (!g2091) & (g2098) & (!g2734) & (g2751) & (g2771)) + ((g2090) & (!g2091) & (g2098) & (g2734) & (g2751) & (g2771)) + ((g2090) & (g2091) & (!g2098) & (!g2734) & (!g2751) & (g2771)) + ((g2090) & (g2091) & (!g2098) & (!g2734) & (g2751) & (g2771)) + ((g2090) & (g2091) & (!g2098) & (g2734) & (!g2751) & (g2771)) + ((g2090) & (g2091) & (!g2098) & (g2734) & (g2751) & (g2771)));
	assign g2881 = (((!g2088) & (!g2089) & (!g2699) & (!g2715) & (!g2848) & (!g2880)) + ((!g2088) & (!g2089) & (!g2699) & (!g2715) & (g2848) & (!g2880)) + ((!g2088) & (!g2089) & (!g2699) & (g2715) & (!g2848) & (!g2880)) + ((!g2088) & (!g2089) & (g2699) & (!g2715) & (!g2848) & (!g2880)) + ((!g2088) & (!g2089) & (g2699) & (g2715) & (!g2848) & (!g2880)) + ((!g2088) & (g2089) & (!g2699) & (!g2715) & (!g2848) & (!g2880)) + ((!g2088) & (g2089) & (!g2699) & (!g2715) & (g2848) & (!g2880)) + ((!g2088) & (g2089) & (!g2699) & (g2715) & (!g2848) & (!g2880)) + ((!g2088) & (g2089) & (!g2699) & (g2715) & (g2848) & (!g2880)) + ((!g2088) & (g2089) & (g2699) & (!g2715) & (!g2848) & (!g2880)) + ((!g2088) & (g2089) & (g2699) & (!g2715) & (g2848) & (!g2880)) + ((!g2088) & (g2089) & (g2699) & (g2715) & (!g2848) & (!g2880)) + ((g2088) & (!g2089) & (!g2699) & (!g2715) & (!g2848) & (!g2880)) + ((g2088) & (!g2089) & (!g2699) & (!g2715) & (g2848) & (!g2880)) + ((g2088) & (!g2089) & (!g2699) & (g2715) & (!g2848) & (!g2880)) + ((g2088) & (!g2089) & (g2699) & (!g2715) & (!g2848) & (!g2880)) + ((g2088) & (!g2089) & (g2699) & (!g2715) & (g2848) & (!g2880)) + ((g2088) & (!g2089) & (g2699) & (g2715) & (!g2848) & (!g2880)) + ((g2088) & (g2089) & (!g2699) & (!g2715) & (!g2848) & (!g2880)) + ((g2088) & (g2089) & (!g2699) & (!g2715) & (g2848) & (!g2880)) + ((g2088) & (g2089) & (!g2699) & (g2715) & (!g2848) & (!g2880)) + ((g2088) & (g2089) & (!g2699) & (g2715) & (g2848) & (!g2880)) + ((g2088) & (g2089) & (g2699) & (!g2715) & (!g2848) & (!g2880)) + ((g2088) & (g2089) & (g2699) & (!g2715) & (g2848) & (!g2880)) + ((g2088) & (g2089) & (g2699) & (g2715) & (!g2848) & (!g2880)) + ((g2088) & (g2089) & (g2699) & (g2715) & (g2848) & (!g2880)));
	assign g2882 = (((!g2095) & (!g2096) & (!g2660) & (g2680) & (!sk[57]) & (!g2849)) + ((!g2095) & (!g2096) & (!g2660) & (g2680) & (!sk[57]) & (g2849)) + ((!g2095) & (!g2096) & (!g2660) & (g2680) & (sk[57]) & (g2849)) + ((!g2095) & (!g2096) & (g2660) & (!g2680) & (!sk[57]) & (!g2849)) + ((!g2095) & (!g2096) & (g2660) & (!g2680) & (!sk[57]) & (g2849)) + ((!g2095) & (!g2096) & (g2660) & (!g2680) & (sk[57]) & (g2849)) + ((!g2095) & (!g2096) & (g2660) & (g2680) & (!sk[57]) & (!g2849)) + ((!g2095) & (!g2096) & (g2660) & (g2680) & (!sk[57]) & (g2849)) + ((!g2095) & (!g2096) & (g2660) & (g2680) & (sk[57]) & (g2849)) + ((!g2095) & (g2096) & (!g2660) & (g2680) & (!sk[57]) & (!g2849)) + ((!g2095) & (g2096) & (!g2660) & (g2680) & (!sk[57]) & (g2849)) + ((!g2095) & (g2096) & (g2660) & (!g2680) & (!sk[57]) & (!g2849)) + ((!g2095) & (g2096) & (g2660) & (!g2680) & (!sk[57]) & (g2849)) + ((!g2095) & (g2096) & (g2660) & (g2680) & (!sk[57]) & (!g2849)) + ((!g2095) & (g2096) & (g2660) & (g2680) & (!sk[57]) & (g2849)) + ((!g2095) & (g2096) & (g2660) & (g2680) & (sk[57]) & (g2849)) + ((g2095) & (!g2096) & (!g2660) & (!g2680) & (!sk[57]) & (!g2849)) + ((g2095) & (!g2096) & (!g2660) & (!g2680) & (!sk[57]) & (g2849)) + ((g2095) & (!g2096) & (!g2660) & (g2680) & (!sk[57]) & (!g2849)) + ((g2095) & (!g2096) & (!g2660) & (g2680) & (!sk[57]) & (g2849)) + ((g2095) & (!g2096) & (!g2660) & (g2680) & (sk[57]) & (g2849)) + ((g2095) & (!g2096) & (g2660) & (!g2680) & (!sk[57]) & (!g2849)) + ((g2095) & (!g2096) & (g2660) & (!g2680) & (!sk[57]) & (g2849)) + ((g2095) & (!g2096) & (g2660) & (g2680) & (!sk[57]) & (!g2849)) + ((g2095) & (!g2096) & (g2660) & (g2680) & (!sk[57]) & (g2849)) + ((g2095) & (!g2096) & (g2660) & (g2680) & (sk[57]) & (g2849)) + ((g2095) & (g2096) & (!g2660) & (!g2680) & (!sk[57]) & (!g2849)) + ((g2095) & (g2096) & (!g2660) & (!g2680) & (!sk[57]) & (g2849)) + ((g2095) & (g2096) & (!g2660) & (g2680) & (!sk[57]) & (!g2849)) + ((g2095) & (g2096) & (!g2660) & (g2680) & (!sk[57]) & (g2849)) + ((g2095) & (g2096) & (g2660) & (!g2680) & (!sk[57]) & (!g2849)) + ((g2095) & (g2096) & (g2660) & (!g2680) & (!sk[57]) & (g2849)) + ((g2095) & (g2096) & (g2660) & (g2680) & (!sk[57]) & (!g2849)) + ((g2095) & (g2096) & (g2660) & (g2680) & (!sk[57]) & (g2849)));
	assign g2883 = (((!g2850) & (!g2879) & (!sk[58]) & (!g2881) & (g2882)) + ((!g2850) & (!g2879) & (!sk[58]) & (g2881) & (g2882)) + ((!g2850) & (!g2879) & (sk[58]) & (g2881) & (!g2882)) + ((!g2850) & (g2879) & (!sk[58]) & (!g2881) & (!g2882)) + ((!g2850) & (g2879) & (!sk[58]) & (!g2881) & (g2882)) + ((!g2850) & (g2879) & (!sk[58]) & (g2881) & (!g2882)) + ((!g2850) & (g2879) & (!sk[58]) & (g2881) & (g2882)) + ((!g2850) & (g2879) & (sk[58]) & (g2881) & (!g2882)) + ((g2850) & (!g2879) & (!sk[58]) & (!g2881) & (!g2882)) + ((g2850) & (!g2879) & (!sk[58]) & (!g2881) & (g2882)) + ((g2850) & (!g2879) & (!sk[58]) & (g2881) & (!g2882)) + ((g2850) & (!g2879) & (!sk[58]) & (g2881) & (g2882)) + ((g2850) & (g2879) & (!sk[58]) & (!g2881) & (!g2882)) + ((g2850) & (g2879) & (!sk[58]) & (!g2881) & (g2882)) + ((g2850) & (g2879) & (!sk[58]) & (g2881) & (!g2882)) + ((g2850) & (g2879) & (!sk[58]) & (g2881) & (g2882)) + ((g2850) & (g2879) & (sk[58]) & (g2881) & (!g2882)));
	assign g2884 = (((!g2100) & (!g2101) & (!g2811) & (!sk[59]) & (g2831)) + ((!g2100) & (!g2101) & (!g2811) & (sk[59]) & (g2831)) + ((!g2100) & (!g2101) & (g2811) & (!sk[59]) & (g2831)) + ((!g2100) & (!g2101) & (g2811) & (sk[59]) & (!g2831)) + ((!g2100) & (!g2101) & (g2811) & (sk[59]) & (g2831)) + ((!g2100) & (g2101) & (!g2811) & (!sk[59]) & (!g2831)) + ((!g2100) & (g2101) & (!g2811) & (!sk[59]) & (g2831)) + ((!g2100) & (g2101) & (g2811) & (!sk[59]) & (!g2831)) + ((!g2100) & (g2101) & (g2811) & (!sk[59]) & (g2831)) + ((!g2100) & (g2101) & (g2811) & (sk[59]) & (g2831)) + ((g2100) & (!g2101) & (!g2811) & (!sk[59]) & (!g2831)) + ((g2100) & (!g2101) & (!g2811) & (!sk[59]) & (g2831)) + ((g2100) & (!g2101) & (!g2811) & (sk[59]) & (g2831)) + ((g2100) & (!g2101) & (g2811) & (!sk[59]) & (!g2831)) + ((g2100) & (!g2101) & (g2811) & (!sk[59]) & (g2831)) + ((g2100) & (!g2101) & (g2811) & (sk[59]) & (g2831)) + ((g2100) & (g2101) & (!g2811) & (!sk[59]) & (!g2831)) + ((g2100) & (g2101) & (!g2811) & (!sk[59]) & (g2831)) + ((g2100) & (g2101) & (g2811) & (!sk[59]) & (!g2831)) + ((g2100) & (g2101) & (g2811) & (!sk[59]) & (g2831)));
	assign g2885 = (((!g2099) & (!g2794) & (!g2857) & (!g2883) & (sk[60]) & (!g2884)) + ((!g2099) & (!g2794) & (!g2857) & (g2883) & (!sk[60]) & (!g2884)) + ((!g2099) & (!g2794) & (!g2857) & (g2883) & (!sk[60]) & (g2884)) + ((!g2099) & (!g2794) & (!g2857) & (g2883) & (sk[60]) & (!g2884)) + ((!g2099) & (!g2794) & (g2857) & (!g2883) & (!sk[60]) & (!g2884)) + ((!g2099) & (!g2794) & (g2857) & (!g2883) & (!sk[60]) & (g2884)) + ((!g2099) & (!g2794) & (g2857) & (g2883) & (!sk[60]) & (!g2884)) + ((!g2099) & (!g2794) & (g2857) & (g2883) & (!sk[60]) & (g2884)) + ((!g2099) & (!g2794) & (g2857) & (g2883) & (sk[60]) & (!g2884)) + ((!g2099) & (g2794) & (!g2857) & (!g2883) & (sk[60]) & (!g2884)) + ((!g2099) & (g2794) & (!g2857) & (g2883) & (!sk[60]) & (!g2884)) + ((!g2099) & (g2794) & (!g2857) & (g2883) & (!sk[60]) & (g2884)) + ((!g2099) & (g2794) & (!g2857) & (g2883) & (sk[60]) & (!g2884)) + ((!g2099) & (g2794) & (g2857) & (!g2883) & (!sk[60]) & (!g2884)) + ((!g2099) & (g2794) & (g2857) & (!g2883) & (!sk[60]) & (g2884)) + ((!g2099) & (g2794) & (g2857) & (g2883) & (!sk[60]) & (!g2884)) + ((!g2099) & (g2794) & (g2857) & (g2883) & (!sk[60]) & (g2884)) + ((g2099) & (!g2794) & (!g2857) & (!g2883) & (!sk[60]) & (!g2884)) + ((g2099) & (!g2794) & (!g2857) & (!g2883) & (!sk[60]) & (g2884)) + ((g2099) & (!g2794) & (!g2857) & (!g2883) & (sk[60]) & (!g2884)) + ((g2099) & (!g2794) & (!g2857) & (g2883) & (!sk[60]) & (!g2884)) + ((g2099) & (!g2794) & (!g2857) & (g2883) & (!sk[60]) & (g2884)) + ((g2099) & (!g2794) & (!g2857) & (g2883) & (sk[60]) & (!g2884)) + ((g2099) & (!g2794) & (g2857) & (!g2883) & (!sk[60]) & (!g2884)) + ((g2099) & (!g2794) & (g2857) & (!g2883) & (!sk[60]) & (g2884)) + ((g2099) & (!g2794) & (g2857) & (!g2883) & (sk[60]) & (!g2884)) + ((g2099) & (!g2794) & (g2857) & (g2883) & (!sk[60]) & (!g2884)) + ((g2099) & (!g2794) & (g2857) & (g2883) & (!sk[60]) & (g2884)) + ((g2099) & (!g2794) & (g2857) & (g2883) & (sk[60]) & (!g2884)) + ((g2099) & (g2794) & (!g2857) & (!g2883) & (!sk[60]) & (!g2884)) + ((g2099) & (g2794) & (!g2857) & (!g2883) & (!sk[60]) & (g2884)) + ((g2099) & (g2794) & (!g2857) & (!g2883) & (sk[60]) & (!g2884)) + ((g2099) & (g2794) & (!g2857) & (g2883) & (!sk[60]) & (!g2884)) + ((g2099) & (g2794) & (!g2857) & (g2883) & (!sk[60]) & (g2884)) + ((g2099) & (g2794) & (!g2857) & (g2883) & (sk[60]) & (!g2884)) + ((g2099) & (g2794) & (g2857) & (!g2883) & (!sk[60]) & (!g2884)) + ((g2099) & (g2794) & (g2857) & (!g2883) & (!sk[60]) & (g2884)) + ((g2099) & (g2794) & (g2857) & (g2883) & (!sk[60]) & (!g2884)) + ((g2099) & (g2794) & (g2857) & (g2883) & (!sk[60]) & (g2884)) + ((g2099) & (g2794) & (g2857) & (g2883) & (sk[60]) & (!g2884)));
	assign g2886 = (((!g110) & (!sk[61]) & (g106) & (!g2866)) + ((!g110) & (!sk[61]) & (g106) & (g2866)) + ((!g110) & (sk[61]) & (g106) & (g2866)) + ((g110) & (!sk[61]) & (!g106) & (!g2866)) + ((g110) & (!sk[61]) & (!g106) & (g2866)) + ((g110) & (!sk[61]) & (g106) & (!g2866)) + ((g110) & (!sk[61]) & (g106) & (g2866)));
	assign g2887 = (((!g2074) & (!g2071) & (!g2070) & (!sk[62]) & (g2104)) + ((!g2074) & (!g2071) & (!g2070) & (sk[62]) & (g2104)) + ((!g2074) & (!g2071) & (g2070) & (!sk[62]) & (g2104)) + ((!g2074) & (!g2071) & (g2070) & (sk[62]) & (!g2104)) + ((!g2074) & (!g2071) & (g2070) & (sk[62]) & (g2104)) + ((!g2074) & (g2071) & (!g2070) & (!sk[62]) & (!g2104)) + ((!g2074) & (g2071) & (!g2070) & (!sk[62]) & (g2104)) + ((!g2074) & (g2071) & (!g2070) & (sk[62]) & (g2104)) + ((!g2074) & (g2071) & (g2070) & (!sk[62]) & (!g2104)) + ((!g2074) & (g2071) & (g2070) & (!sk[62]) & (g2104)) + ((!g2074) & (g2071) & (g2070) & (sk[62]) & (g2104)) + ((g2074) & (!g2071) & (!g2070) & (!sk[62]) & (!g2104)) + ((g2074) & (!g2071) & (!g2070) & (!sk[62]) & (g2104)) + ((g2074) & (!g2071) & (g2070) & (!sk[62]) & (!g2104)) + ((g2074) & (!g2071) & (g2070) & (!sk[62]) & (g2104)) + ((g2074) & (!g2071) & (g2070) & (sk[62]) & (g2104)) + ((g2074) & (g2071) & (!g2070) & (!sk[62]) & (!g2104)) + ((g2074) & (g2071) & (!g2070) & (!sk[62]) & (g2104)) + ((g2074) & (g2071) & (g2070) & (!sk[62]) & (!g2104)) + ((g2074) & (g2071) & (g2070) & (!sk[62]) & (g2104)));
	assign g2888 = (((!g2076) & (!g2077) & (!sk[63]) & (!g2105) & (g2106) & (!g2887)) + ((!g2076) & (!g2077) & (!sk[63]) & (!g2105) & (g2106) & (g2887)) + ((!g2076) & (!g2077) & (!sk[63]) & (g2105) & (!g2106) & (!g2887)) + ((!g2076) & (!g2077) & (!sk[63]) & (g2105) & (!g2106) & (g2887)) + ((!g2076) & (!g2077) & (!sk[63]) & (g2105) & (g2106) & (!g2887)) + ((!g2076) & (!g2077) & (!sk[63]) & (g2105) & (g2106) & (g2887)) + ((!g2076) & (!g2077) & (sk[63]) & (!g2105) & (!g2106) & (g2887)) + ((!g2076) & (!g2077) & (sk[63]) & (!g2105) & (g2106) & (!g2887)) + ((!g2076) & (!g2077) & (sk[63]) & (!g2105) & (g2106) & (g2887)) + ((!g2076) & (!g2077) & (sk[63]) & (g2105) & (!g2106) & (!g2887)) + ((!g2076) & (!g2077) & (sk[63]) & (g2105) & (!g2106) & (g2887)) + ((!g2076) & (!g2077) & (sk[63]) & (g2105) & (g2106) & (!g2887)) + ((!g2076) & (!g2077) & (sk[63]) & (g2105) & (g2106) & (g2887)) + ((!g2076) & (g2077) & (!sk[63]) & (!g2105) & (g2106) & (!g2887)) + ((!g2076) & (g2077) & (!sk[63]) & (!g2105) & (g2106) & (g2887)) + ((!g2076) & (g2077) & (!sk[63]) & (g2105) & (!g2106) & (!g2887)) + ((!g2076) & (g2077) & (!sk[63]) & (g2105) & (!g2106) & (g2887)) + ((!g2076) & (g2077) & (!sk[63]) & (g2105) & (g2106) & (!g2887)) + ((!g2076) & (g2077) & (!sk[63]) & (g2105) & (g2106) & (g2887)) + ((!g2076) & (g2077) & (sk[63]) & (!g2105) & (g2106) & (!g2887)) + ((!g2076) & (g2077) & (sk[63]) & (!g2105) & (g2106) & (g2887)) + ((!g2076) & (g2077) & (sk[63]) & (g2105) & (!g2106) & (g2887)) + ((!g2076) & (g2077) & (sk[63]) & (g2105) & (g2106) & (!g2887)) + ((!g2076) & (g2077) & (sk[63]) & (g2105) & (g2106) & (g2887)) + ((g2076) & (!g2077) & (!sk[63]) & (!g2105) & (!g2106) & (!g2887)) + ((g2076) & (!g2077) & (!sk[63]) & (!g2105) & (!g2106) & (g2887)) + ((g2076) & (!g2077) & (!sk[63]) & (!g2105) & (g2106) & (!g2887)) + ((g2076) & (!g2077) & (!sk[63]) & (!g2105) & (g2106) & (g2887)) + ((g2076) & (!g2077) & (!sk[63]) & (g2105) & (!g2106) & (!g2887)) + ((g2076) & (!g2077) & (!sk[63]) & (g2105) & (!g2106) & (g2887)) + ((g2076) & (!g2077) & (!sk[63]) & (g2105) & (g2106) & (!g2887)) + ((g2076) & (!g2077) & (!sk[63]) & (g2105) & (g2106) & (g2887)) + ((g2076) & (!g2077) & (sk[63]) & (!g2105) & (g2106) & (g2887)) + ((g2076) & (!g2077) & (sk[63]) & (g2105) & (g2106) & (!g2887)) + ((g2076) & (!g2077) & (sk[63]) & (g2105) & (g2106) & (g2887)) + ((g2076) & (g2077) & (!sk[63]) & (!g2105) & (!g2106) & (!g2887)) + ((g2076) & (g2077) & (!sk[63]) & (!g2105) & (!g2106) & (g2887)) + ((g2076) & (g2077) & (!sk[63]) & (!g2105) & (g2106) & (!g2887)) + ((g2076) & (g2077) & (!sk[63]) & (!g2105) & (g2106) & (g2887)) + ((g2076) & (g2077) & (!sk[63]) & (g2105) & (!g2106) & (!g2887)) + ((g2076) & (g2077) & (!sk[63]) & (g2105) & (!g2106) & (g2887)) + ((g2076) & (g2077) & (!sk[63]) & (g2105) & (g2106) & (!g2887)) + ((g2076) & (g2077) & (!sk[63]) & (g2105) & (g2106) & (g2887)) + ((g2076) & (g2077) & (sk[63]) & (g2105) & (g2106) & (g2887)));
	assign g2889 = (((!g2073) & (!g2113) & (!sk[64]) & (!g2114) & (g2289) & (!g2888)) + ((!g2073) & (!g2113) & (!sk[64]) & (!g2114) & (g2289) & (g2888)) + ((!g2073) & (!g2113) & (!sk[64]) & (g2114) & (!g2289) & (!g2888)) + ((!g2073) & (!g2113) & (!sk[64]) & (g2114) & (!g2289) & (g2888)) + ((!g2073) & (!g2113) & (!sk[64]) & (g2114) & (g2289) & (!g2888)) + ((!g2073) & (!g2113) & (!sk[64]) & (g2114) & (g2289) & (g2888)) + ((!g2073) & (!g2113) & (sk[64]) & (!g2114) & (!g2289) & (g2888)) + ((!g2073) & (!g2113) & (sk[64]) & (g2114) & (!g2289) & (!g2888)) + ((!g2073) & (!g2113) & (sk[64]) & (g2114) & (!g2289) & (g2888)) + ((!g2073) & (!g2113) & (sk[64]) & (g2114) & (g2289) & (g2888)) + ((!g2073) & (g2113) & (!sk[64]) & (!g2114) & (g2289) & (!g2888)) + ((!g2073) & (g2113) & (!sk[64]) & (!g2114) & (g2289) & (g2888)) + ((!g2073) & (g2113) & (!sk[64]) & (g2114) & (!g2289) & (!g2888)) + ((!g2073) & (g2113) & (!sk[64]) & (g2114) & (!g2289) & (g2888)) + ((!g2073) & (g2113) & (!sk[64]) & (g2114) & (g2289) & (!g2888)) + ((!g2073) & (g2113) & (!sk[64]) & (g2114) & (g2289) & (g2888)) + ((!g2073) & (g2113) & (sk[64]) & (!g2114) & (!g2289) & (!g2888)) + ((!g2073) & (g2113) & (sk[64]) & (!g2114) & (!g2289) & (g2888)) + ((!g2073) & (g2113) & (sk[64]) & (g2114) & (!g2289) & (!g2888)) + ((!g2073) & (g2113) & (sk[64]) & (g2114) & (!g2289) & (g2888)) + ((!g2073) & (g2113) & (sk[64]) & (g2114) & (g2289) & (!g2888)) + ((!g2073) & (g2113) & (sk[64]) & (g2114) & (g2289) & (g2888)) + ((g2073) & (!g2113) & (!sk[64]) & (!g2114) & (!g2289) & (!g2888)) + ((g2073) & (!g2113) & (!sk[64]) & (!g2114) & (!g2289) & (g2888)) + ((g2073) & (!g2113) & (!sk[64]) & (!g2114) & (g2289) & (!g2888)) + ((g2073) & (!g2113) & (!sk[64]) & (!g2114) & (g2289) & (g2888)) + ((g2073) & (!g2113) & (!sk[64]) & (g2114) & (!g2289) & (!g2888)) + ((g2073) & (!g2113) & (!sk[64]) & (g2114) & (!g2289) & (g2888)) + ((g2073) & (!g2113) & (!sk[64]) & (g2114) & (g2289) & (!g2888)) + ((g2073) & (!g2113) & (!sk[64]) & (g2114) & (g2289) & (g2888)) + ((g2073) & (!g2113) & (sk[64]) & (g2114) & (!g2289) & (!g2888)) + ((g2073) & (!g2113) & (sk[64]) & (g2114) & (!g2289) & (g2888)) + ((g2073) & (g2113) & (!sk[64]) & (!g2114) & (!g2289) & (!g2888)) + ((g2073) & (g2113) & (!sk[64]) & (!g2114) & (!g2289) & (g2888)) + ((g2073) & (g2113) & (!sk[64]) & (!g2114) & (g2289) & (!g2888)) + ((g2073) & (g2113) & (!sk[64]) & (!g2114) & (g2289) & (g2888)) + ((g2073) & (g2113) & (!sk[64]) & (g2114) & (!g2289) & (!g2888)) + ((g2073) & (g2113) & (!sk[64]) & (g2114) & (!g2289) & (g2888)) + ((g2073) & (g2113) & (!sk[64]) & (g2114) & (g2289) & (!g2888)) + ((g2073) & (g2113) & (!sk[64]) & (g2114) & (g2289) & (g2888)) + ((g2073) & (g2113) & (sk[64]) & (!g2114) & (!g2289) & (g2888)) + ((g2073) & (g2113) & (sk[64]) & (g2114) & (!g2289) & (!g2888)) + ((g2073) & (g2113) & (sk[64]) & (g2114) & (!g2289) & (g2888)) + ((g2073) & (g2113) & (sk[64]) & (g2114) & (g2289) & (g2888)));
	assign g2890 = (((!g2115) & (!g2116) & (!g2312) & (!g2340) & (sk[65]) & (g2889)) + ((!g2115) & (!g2116) & (!g2312) & (g2340) & (!sk[65]) & (!g2889)) + ((!g2115) & (!g2116) & (!g2312) & (g2340) & (!sk[65]) & (g2889)) + ((!g2115) & (!g2116) & (g2312) & (!g2340) & (!sk[65]) & (!g2889)) + ((!g2115) & (!g2116) & (g2312) & (!g2340) & (!sk[65]) & (g2889)) + ((!g2115) & (!g2116) & (g2312) & (g2340) & (!sk[65]) & (!g2889)) + ((!g2115) & (!g2116) & (g2312) & (g2340) & (!sk[65]) & (g2889)) + ((!g2115) & (g2116) & (!g2312) & (!g2340) & (sk[65]) & (!g2889)) + ((!g2115) & (g2116) & (!g2312) & (!g2340) & (sk[65]) & (g2889)) + ((!g2115) & (g2116) & (!g2312) & (g2340) & (!sk[65]) & (!g2889)) + ((!g2115) & (g2116) & (!g2312) & (g2340) & (!sk[65]) & (g2889)) + ((!g2115) & (g2116) & (!g2312) & (g2340) & (sk[65]) & (g2889)) + ((!g2115) & (g2116) & (g2312) & (!g2340) & (!sk[65]) & (!g2889)) + ((!g2115) & (g2116) & (g2312) & (!g2340) & (!sk[65]) & (g2889)) + ((!g2115) & (g2116) & (g2312) & (!g2340) & (sk[65]) & (!g2889)) + ((!g2115) & (g2116) & (g2312) & (!g2340) & (sk[65]) & (g2889)) + ((!g2115) & (g2116) & (g2312) & (g2340) & (!sk[65]) & (!g2889)) + ((!g2115) & (g2116) & (g2312) & (g2340) & (!sk[65]) & (g2889)) + ((g2115) & (!g2116) & (!g2312) & (!g2340) & (!sk[65]) & (!g2889)) + ((g2115) & (!g2116) & (!g2312) & (!g2340) & (!sk[65]) & (g2889)) + ((g2115) & (!g2116) & (!g2312) & (!g2340) & (sk[65]) & (!g2889)) + ((g2115) & (!g2116) & (!g2312) & (!g2340) & (sk[65]) & (g2889)) + ((g2115) & (!g2116) & (!g2312) & (g2340) & (!sk[65]) & (!g2889)) + ((g2115) & (!g2116) & (!g2312) & (g2340) & (!sk[65]) & (g2889)) + ((g2115) & (!g2116) & (g2312) & (!g2340) & (!sk[65]) & (!g2889)) + ((g2115) & (!g2116) & (g2312) & (!g2340) & (!sk[65]) & (g2889)) + ((g2115) & (!g2116) & (g2312) & (!g2340) & (sk[65]) & (g2889)) + ((g2115) & (!g2116) & (g2312) & (g2340) & (!sk[65]) & (!g2889)) + ((g2115) & (!g2116) & (g2312) & (g2340) & (!sk[65]) & (g2889)) + ((g2115) & (g2116) & (!g2312) & (!g2340) & (!sk[65]) & (!g2889)) + ((g2115) & (g2116) & (!g2312) & (!g2340) & (!sk[65]) & (g2889)) + ((g2115) & (g2116) & (!g2312) & (!g2340) & (sk[65]) & (!g2889)) + ((g2115) & (g2116) & (!g2312) & (!g2340) & (sk[65]) & (g2889)) + ((g2115) & (g2116) & (!g2312) & (g2340) & (!sk[65]) & (!g2889)) + ((g2115) & (g2116) & (!g2312) & (g2340) & (!sk[65]) & (g2889)) + ((g2115) & (g2116) & (!g2312) & (g2340) & (sk[65]) & (!g2889)) + ((g2115) & (g2116) & (!g2312) & (g2340) & (sk[65]) & (g2889)) + ((g2115) & (g2116) & (g2312) & (!g2340) & (!sk[65]) & (!g2889)) + ((g2115) & (g2116) & (g2312) & (!g2340) & (!sk[65]) & (g2889)) + ((g2115) & (g2116) & (g2312) & (!g2340) & (sk[65]) & (!g2889)) + ((g2115) & (g2116) & (g2312) & (!g2340) & (sk[65]) & (g2889)) + ((g2115) & (g2116) & (g2312) & (g2340) & (!sk[65]) & (!g2889)) + ((g2115) & (g2116) & (g2312) & (g2340) & (!sk[65]) & (g2889)) + ((g2115) & (g2116) & (g2312) & (g2340) & (sk[65]) & (g2889)));
	assign g2891 = (((!g2118) & (!g2119) & (g2120) & (!g2457) & (!g2482) & (!g2507)) + ((!g2118) & (!g2119) & (g2120) & (!g2457) & (g2482) & (!g2507)) + ((!g2118) & (!g2119) & (g2120) & (g2457) & (!g2482) & (!g2507)) + ((!g2118) & (!g2119) & (g2120) & (g2457) & (g2482) & (!g2507)) + ((!g2118) & (g2119) & (!g2120) & (!g2457) & (!g2482) & (!g2507)) + ((!g2118) & (g2119) & (!g2120) & (g2457) & (!g2482) & (!g2507)) + ((!g2118) & (g2119) & (g2120) & (!g2457) & (!g2482) & (!g2507)) + ((!g2118) & (g2119) & (g2120) & (!g2457) & (!g2482) & (g2507)) + ((!g2118) & (g2119) & (g2120) & (!g2457) & (g2482) & (!g2507)) + ((!g2118) & (g2119) & (g2120) & (g2457) & (!g2482) & (!g2507)) + ((!g2118) & (g2119) & (g2120) & (g2457) & (!g2482) & (g2507)) + ((!g2118) & (g2119) & (g2120) & (g2457) & (g2482) & (!g2507)) + ((g2118) & (!g2119) & (!g2120) & (!g2457) & (!g2482) & (!g2507)) + ((g2118) & (!g2119) & (g2120) & (!g2457) & (!g2482) & (!g2507)) + ((g2118) & (!g2119) & (g2120) & (!g2457) & (!g2482) & (g2507)) + ((g2118) & (!g2119) & (g2120) & (!g2457) & (g2482) & (!g2507)) + ((g2118) & (!g2119) & (g2120) & (g2457) & (!g2482) & (!g2507)) + ((g2118) & (!g2119) & (g2120) & (g2457) & (g2482) & (!g2507)) + ((g2118) & (g2119) & (!g2120) & (!g2457) & (!g2482) & (!g2507)) + ((g2118) & (g2119) & (!g2120) & (!g2457) & (g2482) & (!g2507)) + ((g2118) & (g2119) & (!g2120) & (g2457) & (!g2482) & (!g2507)) + ((g2118) & (g2119) & (g2120) & (!g2457) & (!g2482) & (!g2507)) + ((g2118) & (g2119) & (g2120) & (!g2457) & (!g2482) & (g2507)) + ((g2118) & (g2119) & (g2120) & (!g2457) & (g2482) & (!g2507)) + ((g2118) & (g2119) & (g2120) & (!g2457) & (g2482) & (g2507)) + ((g2118) & (g2119) & (g2120) & (g2457) & (!g2482) & (!g2507)) + ((g2118) & (g2119) & (g2120) & (g2457) & (!g2482) & (g2507)) + ((g2118) & (g2119) & (g2120) & (g2457) & (g2482) & (!g2507)));
	assign g2892 = (((!g2109) & (!g2391) & (!g2859) & (!g2851) & (sk[67]) & (!g2891)) + ((!g2109) & (!g2391) & (!g2859) & (g2851) & (!sk[67]) & (!g2891)) + ((!g2109) & (!g2391) & (!g2859) & (g2851) & (!sk[67]) & (g2891)) + ((!g2109) & (!g2391) & (!g2859) & (g2851) & (sk[67]) & (!g2891)) + ((!g2109) & (!g2391) & (g2859) & (!g2851) & (!sk[67]) & (!g2891)) + ((!g2109) & (!g2391) & (g2859) & (!g2851) & (!sk[67]) & (g2891)) + ((!g2109) & (!g2391) & (g2859) & (!g2851) & (sk[67]) & (!g2891)) + ((!g2109) & (!g2391) & (g2859) & (g2851) & (!sk[67]) & (!g2891)) + ((!g2109) & (!g2391) & (g2859) & (g2851) & (!sk[67]) & (g2891)) + ((!g2109) & (!g2391) & (g2859) & (g2851) & (sk[67]) & (!g2891)) + ((!g2109) & (g2391) & (!g2859) & (!g2851) & (sk[67]) & (!g2891)) + ((!g2109) & (g2391) & (!g2859) & (g2851) & (!sk[67]) & (!g2891)) + ((!g2109) & (g2391) & (!g2859) & (g2851) & (!sk[67]) & (g2891)) + ((!g2109) & (g2391) & (!g2859) & (g2851) & (sk[67]) & (!g2891)) + ((!g2109) & (g2391) & (g2859) & (!g2851) & (!sk[67]) & (!g2891)) + ((!g2109) & (g2391) & (g2859) & (!g2851) & (!sk[67]) & (g2891)) + ((!g2109) & (g2391) & (g2859) & (!g2851) & (sk[67]) & (!g2891)) + ((!g2109) & (g2391) & (g2859) & (g2851) & (!sk[67]) & (!g2891)) + ((!g2109) & (g2391) & (g2859) & (g2851) & (!sk[67]) & (g2891)) + ((!g2109) & (g2391) & (g2859) & (g2851) & (sk[67]) & (!g2891)) + ((g2109) & (!g2391) & (!g2859) & (!g2851) & (!sk[67]) & (!g2891)) + ((g2109) & (!g2391) & (!g2859) & (!g2851) & (!sk[67]) & (g2891)) + ((g2109) & (!g2391) & (!g2859) & (!g2851) & (sk[67]) & (!g2891)) + ((g2109) & (!g2391) & (!g2859) & (g2851) & (!sk[67]) & (!g2891)) + ((g2109) & (!g2391) & (!g2859) & (g2851) & (!sk[67]) & (g2891)) + ((g2109) & (!g2391) & (!g2859) & (g2851) & (sk[67]) & (!g2891)) + ((g2109) & (!g2391) & (g2859) & (!g2851) & (!sk[67]) & (!g2891)) + ((g2109) & (!g2391) & (g2859) & (!g2851) & (!sk[67]) & (g2891)) + ((g2109) & (!g2391) & (g2859) & (!g2851) & (sk[67]) & (!g2891)) + ((g2109) & (!g2391) & (g2859) & (g2851) & (!sk[67]) & (!g2891)) + ((g2109) & (!g2391) & (g2859) & (g2851) & (!sk[67]) & (g2891)) + ((g2109) & (g2391) & (!g2859) & (!g2851) & (!sk[67]) & (!g2891)) + ((g2109) & (g2391) & (!g2859) & (!g2851) & (!sk[67]) & (g2891)) + ((g2109) & (g2391) & (!g2859) & (!g2851) & (sk[67]) & (!g2891)) + ((g2109) & (g2391) & (!g2859) & (g2851) & (!sk[67]) & (!g2891)) + ((g2109) & (g2391) & (!g2859) & (g2851) & (!sk[67]) & (g2891)) + ((g2109) & (g2391) & (!g2859) & (g2851) & (sk[67]) & (!g2891)) + ((g2109) & (g2391) & (g2859) & (!g2851) & (!sk[67]) & (!g2891)) + ((g2109) & (g2391) & (g2859) & (!g2851) & (!sk[67]) & (g2891)) + ((g2109) & (g2391) & (g2859) & (!g2851) & (sk[67]) & (!g2891)) + ((g2109) & (g2391) & (g2859) & (g2851) & (!sk[67]) & (!g2891)) + ((g2109) & (g2391) & (g2859) & (g2851) & (!sk[67]) & (g2891)) + ((g2109) & (g2391) & (g2859) & (g2851) & (sk[67]) & (!g2891)));
	assign g2893 = (((!g2110) & (!g2111) & (!g2418) & (!g2439) & (!g2859) & (g2892)) + ((!g2110) & (!g2111) & (!g2418) & (!g2439) & (g2859) & (g2892)) + ((!g2110) & (!g2111) & (!g2418) & (g2439) & (!g2859) & (g2892)) + ((!g2110) & (!g2111) & (!g2418) & (g2439) & (g2859) & (g2892)) + ((!g2110) & (!g2111) & (g2418) & (!g2439) & (!g2859) & (g2892)) + ((!g2110) & (!g2111) & (g2418) & (!g2439) & (g2859) & (g2892)) + ((!g2110) & (!g2111) & (g2418) & (g2439) & (!g2859) & (g2892)) + ((!g2110) & (!g2111) & (g2418) & (g2439) & (g2859) & (g2892)) + ((!g2110) & (g2111) & (!g2418) & (!g2439) & (!g2859) & (g2892)) + ((!g2110) & (g2111) & (!g2418) & (g2439) & (!g2859) & (g2892)) + ((!g2110) & (g2111) & (!g2418) & (g2439) & (g2859) & (g2892)) + ((!g2110) & (g2111) & (g2418) & (!g2439) & (!g2859) & (g2892)) + ((!g2110) & (g2111) & (g2418) & (g2439) & (!g2859) & (g2892)) + ((!g2110) & (g2111) & (g2418) & (g2439) & (g2859) & (g2892)) + ((g2110) & (!g2111) & (!g2418) & (!g2439) & (!g2859) & (g2892)) + ((g2110) & (!g2111) & (!g2418) & (g2439) & (!g2859) & (g2892)) + ((g2110) & (!g2111) & (!g2418) & (g2439) & (g2859) & (g2892)) + ((g2110) & (!g2111) & (g2418) & (!g2439) & (!g2859) & (g2892)) + ((g2110) & (!g2111) & (g2418) & (!g2439) & (g2859) & (g2892)) + ((g2110) & (!g2111) & (g2418) & (g2439) & (!g2859) & (g2892)) + ((g2110) & (!g2111) & (g2418) & (g2439) & (g2859) & (g2892)) + ((g2110) & (g2111) & (!g2418) & (!g2439) & (!g2859) & (g2892)) + ((g2110) & (g2111) & (!g2418) & (g2439) & (!g2859) & (g2892)) + ((g2110) & (g2111) & (g2418) & (!g2439) & (!g2859) & (g2892)) + ((g2110) & (g2111) & (g2418) & (g2439) & (!g2859) & (g2892)) + ((g2110) & (g2111) & (g2418) & (g2439) & (g2859) & (g2892)));
	assign g2894 = (((!g2108) & (!g2365) & (!g2859) & (!g2852) & (!g2890) & (g2893)) + ((!g2108) & (!g2365) & (!g2859) & (!g2852) & (g2890) & (g2893)) + ((!g2108) & (!g2365) & (!g2859) & (g2852) & (!g2890) & (g2893)) + ((!g2108) & (!g2365) & (!g2859) & (g2852) & (g2890) & (g2893)) + ((!g2108) & (!g2365) & (g2859) & (!g2852) & (!g2890) & (g2893)) + ((!g2108) & (!g2365) & (g2859) & (!g2852) & (g2890) & (g2893)) + ((!g2108) & (!g2365) & (g2859) & (g2852) & (!g2890) & (g2893)) + ((!g2108) & (g2365) & (!g2859) & (!g2852) & (!g2890) & (g2893)) + ((!g2108) & (g2365) & (!g2859) & (!g2852) & (g2890) & (g2893)) + ((!g2108) & (g2365) & (!g2859) & (g2852) & (!g2890) & (g2893)) + ((!g2108) & (g2365) & (!g2859) & (g2852) & (g2890) & (g2893)) + ((!g2108) & (g2365) & (g2859) & (!g2852) & (!g2890) & (g2893)) + ((!g2108) & (g2365) & (g2859) & (!g2852) & (g2890) & (g2893)) + ((!g2108) & (g2365) & (g2859) & (g2852) & (!g2890) & (g2893)) + ((!g2108) & (g2365) & (g2859) & (g2852) & (g2890) & (g2893)) + ((g2108) & (!g2365) & (!g2859) & (!g2852) & (!g2890) & (g2893)) + ((g2108) & (!g2365) & (!g2859) & (!g2852) & (g2890) & (g2893)) + ((g2108) & (!g2365) & (!g2859) & (g2852) & (!g2890) & (g2893)) + ((g2108) & (!g2365) & (!g2859) & (g2852) & (g2890) & (g2893)) + ((g2108) & (!g2365) & (g2859) & (!g2852) & (!g2890) & (g2893)) + ((g2108) & (!g2365) & (g2859) & (!g2852) & (g2890) & (g2893)) + ((g2108) & (g2365) & (!g2859) & (!g2852) & (!g2890) & (g2893)) + ((g2108) & (g2365) & (!g2859) & (!g2852) & (g2890) & (g2893)) + ((g2108) & (g2365) & (!g2859) & (g2852) & (!g2890) & (g2893)) + ((g2108) & (g2365) & (!g2859) & (g2852) & (g2890) & (g2893)) + ((g2108) & (g2365) & (g2859) & (!g2852) & (!g2890) & (g2893)) + ((g2108) & (g2365) & (g2859) & (!g2852) & (g2890) & (g2893)) + ((g2108) & (g2365) & (g2859) & (g2852) & (!g2890) & (g2893)));
	assign g2895 = (((!g2086) & (!g2093) & (g2094) & (!g2608) & (!g2625) & (!g2642)) + ((!g2086) & (!g2093) & (g2094) & (!g2608) & (g2625) & (!g2642)) + ((!g2086) & (!g2093) & (g2094) & (g2608) & (!g2625) & (!g2642)) + ((!g2086) & (!g2093) & (g2094) & (g2608) & (g2625) & (!g2642)) + ((!g2086) & (g2093) & (!g2094) & (!g2608) & (!g2625) & (!g2642)) + ((!g2086) & (g2093) & (!g2094) & (g2608) & (!g2625) & (!g2642)) + ((!g2086) & (g2093) & (g2094) & (!g2608) & (!g2625) & (!g2642)) + ((!g2086) & (g2093) & (g2094) & (!g2608) & (!g2625) & (g2642)) + ((!g2086) & (g2093) & (g2094) & (!g2608) & (g2625) & (!g2642)) + ((!g2086) & (g2093) & (g2094) & (g2608) & (!g2625) & (!g2642)) + ((!g2086) & (g2093) & (g2094) & (g2608) & (!g2625) & (g2642)) + ((!g2086) & (g2093) & (g2094) & (g2608) & (g2625) & (!g2642)) + ((g2086) & (!g2093) & (!g2094) & (!g2608) & (!g2625) & (!g2642)) + ((g2086) & (!g2093) & (g2094) & (!g2608) & (!g2625) & (!g2642)) + ((g2086) & (!g2093) & (g2094) & (!g2608) & (!g2625) & (g2642)) + ((g2086) & (!g2093) & (g2094) & (!g2608) & (g2625) & (!g2642)) + ((g2086) & (!g2093) & (g2094) & (g2608) & (!g2625) & (!g2642)) + ((g2086) & (!g2093) & (g2094) & (g2608) & (g2625) & (!g2642)) + ((g2086) & (g2093) & (!g2094) & (!g2608) & (!g2625) & (!g2642)) + ((g2086) & (g2093) & (!g2094) & (!g2608) & (g2625) & (!g2642)) + ((g2086) & (g2093) & (!g2094) & (g2608) & (!g2625) & (!g2642)) + ((g2086) & (g2093) & (g2094) & (!g2608) & (!g2625) & (!g2642)) + ((g2086) & (g2093) & (g2094) & (!g2608) & (!g2625) & (g2642)) + ((g2086) & (g2093) & (g2094) & (!g2608) & (g2625) & (!g2642)) + ((g2086) & (g2093) & (g2094) & (!g2608) & (g2625) & (g2642)) + ((g2086) & (g2093) & (g2094) & (g2608) & (!g2625) & (!g2642)) + ((g2086) & (g2093) & (g2094) & (g2608) & (!g2625) & (g2642)) + ((g2086) & (g2093) & (g2094) & (g2608) & (g2625) & (!g2642)));
	assign g2896 = (((!g2084) & (!g2085) & (!g2570) & (!g2590) & (!g2854) & (!g2895)) + ((!g2084) & (!g2085) & (!g2570) & (!g2590) & (g2854) & (!g2895)) + ((!g2084) & (!g2085) & (!g2570) & (g2590) & (!g2854) & (!g2895)) + ((!g2084) & (!g2085) & (!g2570) & (g2590) & (g2854) & (!g2895)) + ((!g2084) & (!g2085) & (g2570) & (!g2590) & (!g2854) & (!g2895)) + ((!g2084) & (!g2085) & (g2570) & (!g2590) & (g2854) & (!g2895)) + ((!g2084) & (!g2085) & (g2570) & (g2590) & (!g2854) & (!g2895)) + ((!g2084) & (!g2085) & (g2570) & (g2590) & (g2854) & (!g2895)) + ((!g2084) & (g2085) & (!g2570) & (!g2590) & (!g2854) & (!g2895)) + ((!g2084) & (g2085) & (!g2570) & (g2590) & (!g2854) & (!g2895)) + ((!g2084) & (g2085) & (!g2570) & (g2590) & (g2854) & (!g2895)) + ((!g2084) & (g2085) & (g2570) & (!g2590) & (!g2854) & (!g2895)) + ((!g2084) & (g2085) & (g2570) & (g2590) & (!g2854) & (!g2895)) + ((!g2084) & (g2085) & (g2570) & (g2590) & (g2854) & (!g2895)) + ((g2084) & (!g2085) & (!g2570) & (!g2590) & (!g2854) & (!g2895)) + ((g2084) & (!g2085) & (!g2570) & (g2590) & (!g2854) & (!g2895)) + ((g2084) & (!g2085) & (!g2570) & (g2590) & (g2854) & (!g2895)) + ((g2084) & (!g2085) & (g2570) & (!g2590) & (!g2854) & (!g2895)) + ((g2084) & (!g2085) & (g2570) & (!g2590) & (g2854) & (!g2895)) + ((g2084) & (!g2085) & (g2570) & (g2590) & (!g2854) & (!g2895)) + ((g2084) & (!g2085) & (g2570) & (g2590) & (g2854) & (!g2895)) + ((g2084) & (g2085) & (!g2570) & (!g2590) & (!g2854) & (!g2895)) + ((g2084) & (g2085) & (!g2570) & (g2590) & (!g2854) & (!g2895)) + ((g2084) & (g2085) & (g2570) & (!g2590) & (!g2854) & (!g2895)) + ((g2084) & (g2085) & (g2570) & (g2590) & (!g2854) & (!g2895)) + ((g2084) & (g2085) & (g2570) & (g2590) & (g2854) & (!g2895)));
	assign g2897 = (((!g2083) & (!sk[72]) & (!g2121) & (!g2529) & (g2551) & (!g2855)) + ((!g2083) & (!sk[72]) & (!g2121) & (!g2529) & (g2551) & (g2855)) + ((!g2083) & (!sk[72]) & (!g2121) & (g2529) & (!g2551) & (!g2855)) + ((!g2083) & (!sk[72]) & (!g2121) & (g2529) & (!g2551) & (g2855)) + ((!g2083) & (!sk[72]) & (!g2121) & (g2529) & (g2551) & (!g2855)) + ((!g2083) & (!sk[72]) & (!g2121) & (g2529) & (g2551) & (g2855)) + ((!g2083) & (!sk[72]) & (g2121) & (!g2529) & (g2551) & (!g2855)) + ((!g2083) & (!sk[72]) & (g2121) & (!g2529) & (g2551) & (g2855)) + ((!g2083) & (!sk[72]) & (g2121) & (g2529) & (!g2551) & (!g2855)) + ((!g2083) & (!sk[72]) & (g2121) & (g2529) & (!g2551) & (g2855)) + ((!g2083) & (!sk[72]) & (g2121) & (g2529) & (g2551) & (!g2855)) + ((!g2083) & (!sk[72]) & (g2121) & (g2529) & (g2551) & (g2855)) + ((!g2083) & (sk[72]) & (g2121) & (!g2529) & (!g2551) & (g2855)) + ((g2083) & (!sk[72]) & (!g2121) & (!g2529) & (!g2551) & (!g2855)) + ((g2083) & (!sk[72]) & (!g2121) & (!g2529) & (!g2551) & (g2855)) + ((g2083) & (!sk[72]) & (!g2121) & (!g2529) & (g2551) & (!g2855)) + ((g2083) & (!sk[72]) & (!g2121) & (!g2529) & (g2551) & (g2855)) + ((g2083) & (!sk[72]) & (!g2121) & (g2529) & (!g2551) & (!g2855)) + ((g2083) & (!sk[72]) & (!g2121) & (g2529) & (!g2551) & (g2855)) + ((g2083) & (!sk[72]) & (!g2121) & (g2529) & (g2551) & (!g2855)) + ((g2083) & (!sk[72]) & (!g2121) & (g2529) & (g2551) & (g2855)) + ((g2083) & (!sk[72]) & (g2121) & (!g2529) & (!g2551) & (!g2855)) + ((g2083) & (!sk[72]) & (g2121) & (!g2529) & (!g2551) & (g2855)) + ((g2083) & (!sk[72]) & (g2121) & (!g2529) & (g2551) & (!g2855)) + ((g2083) & (!sk[72]) & (g2121) & (!g2529) & (g2551) & (g2855)) + ((g2083) & (!sk[72]) & (g2121) & (g2529) & (!g2551) & (!g2855)) + ((g2083) & (!sk[72]) & (g2121) & (g2529) & (!g2551) & (g2855)) + ((g2083) & (!sk[72]) & (g2121) & (g2529) & (g2551) & (!g2855)) + ((g2083) & (!sk[72]) & (g2121) & (g2529) & (g2551) & (g2855)) + ((g2083) & (sk[72]) & (!g2121) & (!g2529) & (!g2551) & (g2855)) + ((g2083) & (sk[72]) & (!g2121) & (g2529) & (!g2551) & (g2855)) + ((g2083) & (sk[72]) & (g2121) & (!g2529) & (!g2551) & (g2855)) + ((g2083) & (sk[72]) & (g2121) & (!g2529) & (g2551) & (g2855)) + ((g2083) & (sk[72]) & (g2121) & (g2529) & (!g2551) & (g2855)));
	assign g2898 = (((!g2856) & (!g2894) & (!g2896) & (!sk[73]) & (g2897)) + ((!g2856) & (!g2894) & (g2896) & (!sk[73]) & (g2897)) + ((!g2856) & (!g2894) & (g2896) & (sk[73]) & (!g2897)) + ((!g2856) & (g2894) & (!g2896) & (!sk[73]) & (!g2897)) + ((!g2856) & (g2894) & (!g2896) & (!sk[73]) & (g2897)) + ((!g2856) & (g2894) & (g2896) & (!sk[73]) & (!g2897)) + ((!g2856) & (g2894) & (g2896) & (!sk[73]) & (g2897)) + ((!g2856) & (g2894) & (g2896) & (sk[73]) & (!g2897)) + ((g2856) & (!g2894) & (!g2896) & (!sk[73]) & (!g2897)) + ((g2856) & (!g2894) & (!g2896) & (!sk[73]) & (g2897)) + ((g2856) & (!g2894) & (g2896) & (!sk[73]) & (!g2897)) + ((g2856) & (!g2894) & (g2896) & (!sk[73]) & (g2897)) + ((g2856) & (g2894) & (!g2896) & (!sk[73]) & (!g2897)) + ((g2856) & (g2894) & (!g2896) & (!sk[73]) & (g2897)) + ((g2856) & (g2894) & (g2896) & (!sk[73]) & (!g2897)) + ((g2856) & (g2894) & (g2896) & (!sk[73]) & (g2897)) + ((g2856) & (g2894) & (g2896) & (sk[73]) & (!g2897)));
	assign g2899 = (((!g2090) & (!g2091) & (g2098) & (!g2734) & (!g2751) & (!g2771)) + ((!g2090) & (!g2091) & (g2098) & (!g2734) & (g2751) & (!g2771)) + ((!g2090) & (!g2091) & (g2098) & (g2734) & (!g2751) & (!g2771)) + ((!g2090) & (!g2091) & (g2098) & (g2734) & (g2751) & (!g2771)) + ((!g2090) & (g2091) & (!g2098) & (!g2734) & (!g2751) & (!g2771)) + ((!g2090) & (g2091) & (!g2098) & (g2734) & (!g2751) & (!g2771)) + ((!g2090) & (g2091) & (g2098) & (!g2734) & (!g2751) & (!g2771)) + ((!g2090) & (g2091) & (g2098) & (!g2734) & (!g2751) & (g2771)) + ((!g2090) & (g2091) & (g2098) & (!g2734) & (g2751) & (!g2771)) + ((!g2090) & (g2091) & (g2098) & (g2734) & (!g2751) & (!g2771)) + ((!g2090) & (g2091) & (g2098) & (g2734) & (!g2751) & (g2771)) + ((!g2090) & (g2091) & (g2098) & (g2734) & (g2751) & (!g2771)) + ((g2090) & (!g2091) & (!g2098) & (!g2734) & (!g2751) & (!g2771)) + ((g2090) & (!g2091) & (g2098) & (!g2734) & (!g2751) & (!g2771)) + ((g2090) & (!g2091) & (g2098) & (!g2734) & (!g2751) & (g2771)) + ((g2090) & (!g2091) & (g2098) & (!g2734) & (g2751) & (!g2771)) + ((g2090) & (!g2091) & (g2098) & (g2734) & (!g2751) & (!g2771)) + ((g2090) & (!g2091) & (g2098) & (g2734) & (g2751) & (!g2771)) + ((g2090) & (g2091) & (!g2098) & (!g2734) & (!g2751) & (!g2771)) + ((g2090) & (g2091) & (!g2098) & (!g2734) & (g2751) & (!g2771)) + ((g2090) & (g2091) & (!g2098) & (g2734) & (!g2751) & (!g2771)) + ((g2090) & (g2091) & (g2098) & (!g2734) & (!g2751) & (!g2771)) + ((g2090) & (g2091) & (g2098) & (!g2734) & (!g2751) & (g2771)) + ((g2090) & (g2091) & (g2098) & (!g2734) & (g2751) & (!g2771)) + ((g2090) & (g2091) & (g2098) & (!g2734) & (g2751) & (g2771)) + ((g2090) & (g2091) & (g2098) & (g2734) & (!g2751) & (!g2771)) + ((g2090) & (g2091) & (g2098) & (g2734) & (!g2751) & (g2771)) + ((g2090) & (g2091) & (g2098) & (g2734) & (g2751) & (!g2771)));
	assign g2900 = (((!g2088) & (!g2089) & (!g2699) & (!g2715) & (!g2848) & (!g2899)) + ((!g2088) & (!g2089) & (!g2699) & (!g2715) & (g2848) & (!g2899)) + ((!g2088) & (!g2089) & (!g2699) & (g2715) & (!g2848) & (!g2899)) + ((!g2088) & (!g2089) & (!g2699) & (g2715) & (g2848) & (!g2899)) + ((!g2088) & (!g2089) & (g2699) & (!g2715) & (!g2848) & (!g2899)) + ((!g2088) & (!g2089) & (g2699) & (!g2715) & (g2848) & (!g2899)) + ((!g2088) & (!g2089) & (g2699) & (g2715) & (!g2848) & (!g2899)) + ((!g2088) & (!g2089) & (g2699) & (g2715) & (g2848) & (!g2899)) + ((!g2088) & (g2089) & (!g2699) & (!g2715) & (!g2848) & (!g2899)) + ((!g2088) & (g2089) & (!g2699) & (g2715) & (!g2848) & (!g2899)) + ((!g2088) & (g2089) & (!g2699) & (g2715) & (g2848) & (!g2899)) + ((!g2088) & (g2089) & (g2699) & (!g2715) & (!g2848) & (!g2899)) + ((!g2088) & (g2089) & (g2699) & (g2715) & (!g2848) & (!g2899)) + ((!g2088) & (g2089) & (g2699) & (g2715) & (g2848) & (!g2899)) + ((g2088) & (!g2089) & (!g2699) & (!g2715) & (!g2848) & (!g2899)) + ((g2088) & (!g2089) & (!g2699) & (g2715) & (!g2848) & (!g2899)) + ((g2088) & (!g2089) & (!g2699) & (g2715) & (g2848) & (!g2899)) + ((g2088) & (!g2089) & (g2699) & (!g2715) & (!g2848) & (!g2899)) + ((g2088) & (!g2089) & (g2699) & (!g2715) & (g2848) & (!g2899)) + ((g2088) & (!g2089) & (g2699) & (g2715) & (!g2848) & (!g2899)) + ((g2088) & (!g2089) & (g2699) & (g2715) & (g2848) & (!g2899)) + ((g2088) & (g2089) & (!g2699) & (!g2715) & (!g2848) & (!g2899)) + ((g2088) & (g2089) & (!g2699) & (g2715) & (!g2848) & (!g2899)) + ((g2088) & (g2089) & (g2699) & (!g2715) & (!g2848) & (!g2899)) + ((g2088) & (g2089) & (g2699) & (g2715) & (!g2848) & (!g2899)) + ((g2088) & (g2089) & (g2699) & (g2715) & (g2848) & (!g2899)));
	assign g2901 = (((!g2095) & (!g2096) & (!g2660) & (g2680) & (!sk[76]) & (!g2849)) + ((!g2095) & (!g2096) & (!g2660) & (g2680) & (!sk[76]) & (g2849)) + ((!g2095) & (!g2096) & (g2660) & (!g2680) & (!sk[76]) & (!g2849)) + ((!g2095) & (!g2096) & (g2660) & (!g2680) & (!sk[76]) & (g2849)) + ((!g2095) & (!g2096) & (g2660) & (g2680) & (!sk[76]) & (!g2849)) + ((!g2095) & (!g2096) & (g2660) & (g2680) & (!sk[76]) & (g2849)) + ((!g2095) & (g2096) & (!g2660) & (!g2680) & (sk[76]) & (g2849)) + ((!g2095) & (g2096) & (!g2660) & (g2680) & (!sk[76]) & (!g2849)) + ((!g2095) & (g2096) & (!g2660) & (g2680) & (!sk[76]) & (g2849)) + ((!g2095) & (g2096) & (g2660) & (!g2680) & (!sk[76]) & (!g2849)) + ((!g2095) & (g2096) & (g2660) & (!g2680) & (!sk[76]) & (g2849)) + ((!g2095) & (g2096) & (g2660) & (!g2680) & (sk[76]) & (g2849)) + ((!g2095) & (g2096) & (g2660) & (g2680) & (!sk[76]) & (!g2849)) + ((!g2095) & (g2096) & (g2660) & (g2680) & (!sk[76]) & (g2849)) + ((g2095) & (!g2096) & (!g2660) & (!g2680) & (!sk[76]) & (!g2849)) + ((g2095) & (!g2096) & (!g2660) & (!g2680) & (!sk[76]) & (g2849)) + ((g2095) & (!g2096) & (!g2660) & (!g2680) & (sk[76]) & (g2849)) + ((g2095) & (!g2096) & (!g2660) & (g2680) & (!sk[76]) & (!g2849)) + ((g2095) & (!g2096) & (!g2660) & (g2680) & (!sk[76]) & (g2849)) + ((g2095) & (!g2096) & (g2660) & (!g2680) & (!sk[76]) & (!g2849)) + ((g2095) & (!g2096) & (g2660) & (!g2680) & (!sk[76]) & (g2849)) + ((g2095) & (!g2096) & (g2660) & (g2680) & (!sk[76]) & (!g2849)) + ((g2095) & (!g2096) & (g2660) & (g2680) & (!sk[76]) & (g2849)) + ((g2095) & (g2096) & (!g2660) & (!g2680) & (!sk[76]) & (!g2849)) + ((g2095) & (g2096) & (!g2660) & (!g2680) & (!sk[76]) & (g2849)) + ((g2095) & (g2096) & (!g2660) & (!g2680) & (sk[76]) & (g2849)) + ((g2095) & (g2096) & (!g2660) & (g2680) & (!sk[76]) & (!g2849)) + ((g2095) & (g2096) & (!g2660) & (g2680) & (!sk[76]) & (g2849)) + ((g2095) & (g2096) & (!g2660) & (g2680) & (sk[76]) & (g2849)) + ((g2095) & (g2096) & (g2660) & (!g2680) & (!sk[76]) & (!g2849)) + ((g2095) & (g2096) & (g2660) & (!g2680) & (!sk[76]) & (g2849)) + ((g2095) & (g2096) & (g2660) & (!g2680) & (sk[76]) & (g2849)) + ((g2095) & (g2096) & (g2660) & (g2680) & (!sk[76]) & (!g2849)) + ((g2095) & (g2096) & (g2660) & (g2680) & (!sk[76]) & (g2849)));
	assign g2902 = (((!g2850) & (!sk[77]) & (!g2898) & (!g2900) & (g2901)) + ((!g2850) & (!sk[77]) & (!g2898) & (g2900) & (g2901)) + ((!g2850) & (!sk[77]) & (g2898) & (!g2900) & (!g2901)) + ((!g2850) & (!sk[77]) & (g2898) & (!g2900) & (g2901)) + ((!g2850) & (!sk[77]) & (g2898) & (g2900) & (!g2901)) + ((!g2850) & (!sk[77]) & (g2898) & (g2900) & (g2901)) + ((!g2850) & (sk[77]) & (!g2898) & (g2900) & (!g2901)) + ((!g2850) & (sk[77]) & (g2898) & (g2900) & (!g2901)) + ((g2850) & (!sk[77]) & (!g2898) & (!g2900) & (!g2901)) + ((g2850) & (!sk[77]) & (!g2898) & (!g2900) & (g2901)) + ((g2850) & (!sk[77]) & (!g2898) & (g2900) & (!g2901)) + ((g2850) & (!sk[77]) & (!g2898) & (g2900) & (g2901)) + ((g2850) & (!sk[77]) & (g2898) & (!g2900) & (!g2901)) + ((g2850) & (!sk[77]) & (g2898) & (!g2900) & (g2901)) + ((g2850) & (!sk[77]) & (g2898) & (g2900) & (!g2901)) + ((g2850) & (!sk[77]) & (g2898) & (g2900) & (g2901)) + ((g2850) & (sk[77]) & (g2898) & (g2900) & (!g2901)));
	assign g2903 = (((!g2100) & (!g2101) & (!sk[78]) & (!g2811) & (g2831)) + ((!g2100) & (!g2101) & (!sk[78]) & (g2811) & (g2831)) + ((!g2100) & (g2101) & (!sk[78]) & (!g2811) & (!g2831)) + ((!g2100) & (g2101) & (!sk[78]) & (!g2811) & (g2831)) + ((!g2100) & (g2101) & (!sk[78]) & (g2811) & (!g2831)) + ((!g2100) & (g2101) & (!sk[78]) & (g2811) & (g2831)) + ((!g2100) & (g2101) & (sk[78]) & (!g2811) & (!g2831)) + ((!g2100) & (g2101) & (sk[78]) & (g2811) & (!g2831)) + ((g2100) & (!g2101) & (!sk[78]) & (!g2811) & (!g2831)) + ((g2100) & (!g2101) & (!sk[78]) & (!g2811) & (g2831)) + ((g2100) & (!g2101) & (!sk[78]) & (g2811) & (!g2831)) + ((g2100) & (!g2101) & (!sk[78]) & (g2811) & (g2831)) + ((g2100) & (!g2101) & (sk[78]) & (!g2811) & (!g2831)) + ((g2100) & (g2101) & (!sk[78]) & (!g2811) & (!g2831)) + ((g2100) & (g2101) & (!sk[78]) & (!g2811) & (g2831)) + ((g2100) & (g2101) & (!sk[78]) & (g2811) & (!g2831)) + ((g2100) & (g2101) & (!sk[78]) & (g2811) & (g2831)) + ((g2100) & (g2101) & (sk[78]) & (!g2811) & (!g2831)) + ((g2100) & (g2101) & (sk[78]) & (!g2811) & (g2831)) + ((g2100) & (g2101) & (sk[78]) & (g2811) & (!g2831)));
	assign g2904 = (((!g2099) & (!sk[79]) & (!g2794) & (!g2857) & (g2902) & (!g2903)) + ((!g2099) & (!sk[79]) & (!g2794) & (!g2857) & (g2902) & (g2903)) + ((!g2099) & (!sk[79]) & (!g2794) & (g2857) & (!g2902) & (!g2903)) + ((!g2099) & (!sk[79]) & (!g2794) & (g2857) & (!g2902) & (g2903)) + ((!g2099) & (!sk[79]) & (!g2794) & (g2857) & (g2902) & (!g2903)) + ((!g2099) & (!sk[79]) & (!g2794) & (g2857) & (g2902) & (g2903)) + ((!g2099) & (!sk[79]) & (g2794) & (!g2857) & (g2902) & (!g2903)) + ((!g2099) & (!sk[79]) & (g2794) & (!g2857) & (g2902) & (g2903)) + ((!g2099) & (!sk[79]) & (g2794) & (g2857) & (!g2902) & (!g2903)) + ((!g2099) & (!sk[79]) & (g2794) & (g2857) & (!g2902) & (g2903)) + ((!g2099) & (!sk[79]) & (g2794) & (g2857) & (g2902) & (!g2903)) + ((!g2099) & (!sk[79]) & (g2794) & (g2857) & (g2902) & (g2903)) + ((!g2099) & (sk[79]) & (!g2794) & (!g2857) & (!g2902) & (!g2903)) + ((!g2099) & (sk[79]) & (!g2794) & (!g2857) & (g2902) & (!g2903)) + ((!g2099) & (sk[79]) & (!g2794) & (g2857) & (g2902) & (!g2903)) + ((!g2099) & (sk[79]) & (g2794) & (!g2857) & (!g2902) & (!g2903)) + ((!g2099) & (sk[79]) & (g2794) & (!g2857) & (g2902) & (!g2903)) + ((!g2099) & (sk[79]) & (g2794) & (g2857) & (!g2902) & (!g2903)) + ((!g2099) & (sk[79]) & (g2794) & (g2857) & (g2902) & (!g2903)) + ((g2099) & (!sk[79]) & (!g2794) & (!g2857) & (!g2902) & (!g2903)) + ((g2099) & (!sk[79]) & (!g2794) & (!g2857) & (!g2902) & (g2903)) + ((g2099) & (!sk[79]) & (!g2794) & (!g2857) & (g2902) & (!g2903)) + ((g2099) & (!sk[79]) & (!g2794) & (!g2857) & (g2902) & (g2903)) + ((g2099) & (!sk[79]) & (!g2794) & (g2857) & (!g2902) & (!g2903)) + ((g2099) & (!sk[79]) & (!g2794) & (g2857) & (!g2902) & (g2903)) + ((g2099) & (!sk[79]) & (!g2794) & (g2857) & (g2902) & (!g2903)) + ((g2099) & (!sk[79]) & (!g2794) & (g2857) & (g2902) & (g2903)) + ((g2099) & (!sk[79]) & (g2794) & (!g2857) & (!g2902) & (!g2903)) + ((g2099) & (!sk[79]) & (g2794) & (!g2857) & (!g2902) & (g2903)) + ((g2099) & (!sk[79]) & (g2794) & (!g2857) & (g2902) & (!g2903)) + ((g2099) & (!sk[79]) & (g2794) & (!g2857) & (g2902) & (g2903)) + ((g2099) & (!sk[79]) & (g2794) & (g2857) & (!g2902) & (!g2903)) + ((g2099) & (!sk[79]) & (g2794) & (g2857) & (!g2902) & (g2903)) + ((g2099) & (!sk[79]) & (g2794) & (g2857) & (g2902) & (!g2903)) + ((g2099) & (!sk[79]) & (g2794) & (g2857) & (g2902) & (g2903)) + ((g2099) & (sk[79]) & (!g2794) & (!g2857) & (!g2902) & (!g2903)) + ((g2099) & (sk[79]) & (!g2794) & (!g2857) & (g2902) & (!g2903)) + ((g2099) & (sk[79]) & (g2794) & (!g2857) & (!g2902) & (!g2903)) + ((g2099) & (sk[79]) & (g2794) & (!g2857) & (g2902) & (!g2903)) + ((g2099) & (sk[79]) & (g2794) & (g2857) & (g2902) & (!g2903)));
	assign g2905 = (((!sk[80]) & (!g110) & (g106) & (!g2847)) + ((!sk[80]) & (!g110) & (g106) & (g2847)) + ((!sk[80]) & (g110) & (!g106) & (!g2847)) + ((!sk[80]) & (g110) & (!g106) & (g2847)) + ((!sk[80]) & (g110) & (g106) & (!g2847)) + ((!sk[80]) & (g110) & (g106) & (g2847)) + ((sk[80]) & (!g110) & (g106) & (g2847)));
	assign g2906 = (((!g108) & (!g109) & (!g110) & (!sk[81]) & (g678) & (!g2846)) + ((!g108) & (!g109) & (!g110) & (!sk[81]) & (g678) & (g2846)) + ((!g108) & (!g109) & (!g110) & (sk[81]) & (g678) & (g2846)) + ((!g108) & (!g109) & (g110) & (!sk[81]) & (!g678) & (!g2846)) + ((!g108) & (!g109) & (g110) & (!sk[81]) & (!g678) & (g2846)) + ((!g108) & (!g109) & (g110) & (!sk[81]) & (g678) & (!g2846)) + ((!g108) & (!g109) & (g110) & (!sk[81]) & (g678) & (g2846)) + ((!g108) & (g109) & (!g110) & (!sk[81]) & (g678) & (!g2846)) + ((!g108) & (g109) & (!g110) & (!sk[81]) & (g678) & (g2846)) + ((!g108) & (g109) & (g110) & (!sk[81]) & (!g678) & (!g2846)) + ((!g108) & (g109) & (g110) & (!sk[81]) & (!g678) & (g2846)) + ((!g108) & (g109) & (g110) & (!sk[81]) & (g678) & (!g2846)) + ((!g108) & (g109) & (g110) & (!sk[81]) & (g678) & (g2846)) + ((g108) & (!g109) & (!g110) & (!sk[81]) & (!g678) & (!g2846)) + ((g108) & (!g109) & (!g110) & (!sk[81]) & (!g678) & (g2846)) + ((g108) & (!g109) & (!g110) & (!sk[81]) & (g678) & (!g2846)) + ((g108) & (!g109) & (!g110) & (!sk[81]) & (g678) & (g2846)) + ((g108) & (!g109) & (g110) & (!sk[81]) & (!g678) & (!g2846)) + ((g108) & (!g109) & (g110) & (!sk[81]) & (!g678) & (g2846)) + ((g108) & (!g109) & (g110) & (!sk[81]) & (g678) & (!g2846)) + ((g108) & (!g109) & (g110) & (!sk[81]) & (g678) & (g2846)) + ((g108) & (g109) & (!g110) & (!sk[81]) & (!g678) & (!g2846)) + ((g108) & (g109) & (!g110) & (!sk[81]) & (!g678) & (g2846)) + ((g108) & (g109) & (!g110) & (!sk[81]) & (g678) & (!g2846)) + ((g108) & (g109) & (!g110) & (!sk[81]) & (g678) & (g2846)) + ((g108) & (g109) & (g110) & (!sk[81]) & (!g678) & (!g2846)) + ((g108) & (g109) & (g110) & (!sk[81]) & (!g678) & (g2846)) + ((g108) & (g109) & (g110) & (!sk[81]) & (g678) & (!g2846)) + ((g108) & (g109) & (g110) & (!sk[81]) & (g678) & (g2846)));
	assign g2907 = (((!g108) & (!g109) & (!g110) & (g678) & (!sk[82]) & (!g2846)) + ((!g108) & (!g109) & (!g110) & (g678) & (!sk[82]) & (g2846)) + ((!g108) & (!g109) & (!g110) & (g678) & (sk[82]) & (g2846)) + ((!g108) & (!g109) & (g110) & (!g678) & (!sk[82]) & (!g2846)) + ((!g108) & (!g109) & (g110) & (!g678) & (!sk[82]) & (g2846)) + ((!g108) & (!g109) & (g110) & (g678) & (!sk[82]) & (!g2846)) + ((!g108) & (!g109) & (g110) & (g678) & (!sk[82]) & (g2846)) + ((!g108) & (g109) & (!g110) & (!g678) & (sk[82]) & (g2846)) + ((!g108) & (g109) & (!g110) & (g678) & (!sk[82]) & (!g2846)) + ((!g108) & (g109) & (!g110) & (g678) & (!sk[82]) & (g2846)) + ((!g108) & (g109) & (g110) & (!g678) & (!sk[82]) & (!g2846)) + ((!g108) & (g109) & (g110) & (!g678) & (!sk[82]) & (g2846)) + ((!g108) & (g109) & (g110) & (!g678) & (sk[82]) & (g2846)) + ((!g108) & (g109) & (g110) & (g678) & (!sk[82]) & (!g2846)) + ((!g108) & (g109) & (g110) & (g678) & (!sk[82]) & (g2846)) + ((g108) & (!g109) & (!g110) & (!g678) & (!sk[82]) & (!g2846)) + ((g108) & (!g109) & (!g110) & (!g678) & (!sk[82]) & (g2846)) + ((g108) & (!g109) & (!g110) & (!g678) & (sk[82]) & (g2846)) + ((g108) & (!g109) & (!g110) & (g678) & (!sk[82]) & (!g2846)) + ((g108) & (!g109) & (!g110) & (g678) & (!sk[82]) & (g2846)) + ((g108) & (!g109) & (g110) & (!g678) & (!sk[82]) & (!g2846)) + ((g108) & (!g109) & (g110) & (!g678) & (!sk[82]) & (g2846)) + ((g108) & (!g109) & (g110) & (!g678) & (sk[82]) & (g2846)) + ((g108) & (!g109) & (g110) & (g678) & (!sk[82]) & (!g2846)) + ((g108) & (!g109) & (g110) & (g678) & (!sk[82]) & (g2846)) + ((g108) & (g109) & (!g110) & (!g678) & (!sk[82]) & (!g2846)) + ((g108) & (g109) & (!g110) & (!g678) & (!sk[82]) & (g2846)) + ((g108) & (g109) & (!g110) & (g678) & (!sk[82]) & (!g2846)) + ((g108) & (g109) & (!g110) & (g678) & (!sk[82]) & (g2846)) + ((g108) & (g109) & (g110) & (!g678) & (!sk[82]) & (!g2846)) + ((g108) & (g109) & (g110) & (!g678) & (!sk[82]) & (g2846)) + ((g108) & (g109) & (g110) & (g678) & (!sk[82]) & (!g2846)) + ((g108) & (g109) & (g110) & (g678) & (!sk[82]) & (g2846)));
	assign g2908 = (((!g106) & (!g2864) & (!g2906) & (!sk[83]) & (g2907)) + ((!g106) & (!g2864) & (g2906) & (!sk[83]) & (g2907)) + ((!g106) & (g2864) & (!g2906) & (!sk[83]) & (!g2907)) + ((!g106) & (g2864) & (!g2906) & (!sk[83]) & (g2907)) + ((!g106) & (g2864) & (!g2906) & (sk[83]) & (!g2907)) + ((!g106) & (g2864) & (!g2906) & (sk[83]) & (g2907)) + ((!g106) & (g2864) & (g2906) & (!sk[83]) & (!g2907)) + ((!g106) & (g2864) & (g2906) & (!sk[83]) & (g2907)) + ((!g106) & (g2864) & (g2906) & (sk[83]) & (!g2907)) + ((!g106) & (g2864) & (g2906) & (sk[83]) & (g2907)) + ((g106) & (!g2864) & (!g2906) & (!sk[83]) & (!g2907)) + ((g106) & (!g2864) & (!g2906) & (!sk[83]) & (g2907)) + ((g106) & (!g2864) & (g2906) & (!sk[83]) & (!g2907)) + ((g106) & (!g2864) & (g2906) & (!sk[83]) & (g2907)) + ((g106) & (!g2864) & (g2906) & (sk[83]) & (!g2907)) + ((g106) & (!g2864) & (g2906) & (sk[83]) & (g2907)) + ((g106) & (g2864) & (!g2906) & (!sk[83]) & (!g2907)) + ((g106) & (g2864) & (!g2906) & (!sk[83]) & (g2907)) + ((g106) & (g2864) & (!g2906) & (sk[83]) & (!g2907)) + ((g106) & (g2864) & (g2906) & (!sk[83]) & (!g2907)) + ((g106) & (g2864) & (g2906) & (!sk[83]) & (g2907)) + ((g106) & (g2864) & (g2906) & (sk[83]) & (!g2907)));
	assign g2909 = (((!g2885) & (!g2886) & (!g2904) & (!g2905) & (sk[84]) & (!g2908)) + ((!g2885) & (!g2886) & (!g2904) & (g2905) & (!sk[84]) & (!g2908)) + ((!g2885) & (!g2886) & (!g2904) & (g2905) & (!sk[84]) & (g2908)) + ((!g2885) & (!g2886) & (g2904) & (!g2905) & (!sk[84]) & (!g2908)) + ((!g2885) & (!g2886) & (g2904) & (!g2905) & (!sk[84]) & (g2908)) + ((!g2885) & (!g2886) & (g2904) & (!g2905) & (sk[84]) & (!g2908)) + ((!g2885) & (!g2886) & (g2904) & (g2905) & (!sk[84]) & (!g2908)) + ((!g2885) & (!g2886) & (g2904) & (g2905) & (!sk[84]) & (g2908)) + ((!g2885) & (!g2886) & (g2904) & (g2905) & (sk[84]) & (!g2908)) + ((!g2885) & (g2886) & (!g2904) & (g2905) & (!sk[84]) & (!g2908)) + ((!g2885) & (g2886) & (!g2904) & (g2905) & (!sk[84]) & (g2908)) + ((!g2885) & (g2886) & (g2904) & (!g2905) & (!sk[84]) & (!g2908)) + ((!g2885) & (g2886) & (g2904) & (!g2905) & (!sk[84]) & (g2908)) + ((!g2885) & (g2886) & (g2904) & (g2905) & (!sk[84]) & (!g2908)) + ((!g2885) & (g2886) & (g2904) & (g2905) & (!sk[84]) & (g2908)) + ((g2885) & (!g2886) & (!g2904) & (!g2905) & (!sk[84]) & (!g2908)) + ((g2885) & (!g2886) & (!g2904) & (!g2905) & (!sk[84]) & (g2908)) + ((g2885) & (!g2886) & (!g2904) & (!g2905) & (sk[84]) & (!g2908)) + ((g2885) & (!g2886) & (!g2904) & (g2905) & (!sk[84]) & (!g2908)) + ((g2885) & (!g2886) & (!g2904) & (g2905) & (!sk[84]) & (g2908)) + ((g2885) & (!g2886) & (g2904) & (!g2905) & (!sk[84]) & (!g2908)) + ((g2885) & (!g2886) & (g2904) & (!g2905) & (!sk[84]) & (g2908)) + ((g2885) & (!g2886) & (g2904) & (!g2905) & (sk[84]) & (!g2908)) + ((g2885) & (!g2886) & (g2904) & (g2905) & (!sk[84]) & (!g2908)) + ((g2885) & (!g2886) & (g2904) & (g2905) & (!sk[84]) & (g2908)) + ((g2885) & (!g2886) & (g2904) & (g2905) & (sk[84]) & (!g2908)) + ((g2885) & (g2886) & (!g2904) & (!g2905) & (!sk[84]) & (!g2908)) + ((g2885) & (g2886) & (!g2904) & (!g2905) & (!sk[84]) & (g2908)) + ((g2885) & (g2886) & (!g2904) & (!g2905) & (sk[84]) & (!g2908)) + ((g2885) & (g2886) & (!g2904) & (g2905) & (!sk[84]) & (!g2908)) + ((g2885) & (g2886) & (!g2904) & (g2905) & (!sk[84]) & (g2908)) + ((g2885) & (g2886) & (g2904) & (!g2905) & (!sk[84]) & (!g2908)) + ((g2885) & (g2886) & (g2904) & (!g2905) & (!sk[84]) & (g2908)) + ((g2885) & (g2886) & (g2904) & (!g2905) & (sk[84]) & (!g2908)) + ((g2885) & (g2886) & (g2904) & (g2905) & (!sk[84]) & (!g2908)) + ((g2885) & (g2886) & (g2904) & (g2905) & (!sk[84]) & (g2908)) + ((g2885) & (g2886) & (g2904) & (g2905) & (sk[84]) & (!g2908)));
	assign g2910 = (((!g2101) & (!g2831) & (!g2836) & (!g2865) & (!g2867) & (g2909)) + ((!g2101) & (!g2831) & (!g2836) & (!g2865) & (g2867) & (g2909)) + ((!g2101) & (!g2831) & (g2836) & (!g2865) & (!g2867) & (g2909)) + ((!g2101) & (!g2831) & (g2836) & (g2865) & (!g2867) & (g2909)) + ((!g2101) & (g2831) & (!g2836) & (!g2865) & (!g2867) & (g2909)) + ((!g2101) & (g2831) & (!g2836) & (!g2865) & (g2867) & (g2909)) + ((!g2101) & (g2831) & (g2836) & (!g2865) & (!g2867) & (g2909)) + ((!g2101) & (g2831) & (g2836) & (!g2865) & (g2867) & (g2909)) + ((g2101) & (!g2831) & (!g2836) & (!g2865) & (!g2867) & (g2909)) + ((g2101) & (!g2831) & (!g2836) & (g2865) & (!g2867) & (g2909)) + ((g2101) & (!g2831) & (g2836) & (!g2865) & (!g2867) & (g2909)) + ((g2101) & (!g2831) & (g2836) & (g2865) & (!g2867) & (g2909)) + ((g2101) & (g2831) & (!g2836) & (!g2865) & (!g2867) & (g2909)) + ((g2101) & (g2831) & (!g2836) & (!g2865) & (g2867) & (g2909)) + ((g2101) & (g2831) & (g2836) & (!g2865) & (!g2867) & (g2909)) + ((g2101) & (g2831) & (g2836) & (g2865) & (!g2867) & (g2909)));
	assign g2911 = (((!sk[86]) & (!g2081) & (g2124) & (!g2190)) + ((!sk[86]) & (!g2081) & (g2124) & (g2190)) + ((!sk[86]) & (g2081) & (!g2124) & (!g2190)) + ((!sk[86]) & (g2081) & (!g2124) & (g2190)) + ((!sk[86]) & (g2081) & (g2124) & (!g2190)) + ((!sk[86]) & (g2081) & (g2124) & (g2190)) + ((sk[86]) & (!g2081) & (g2124) & (g2190)));
	assign g2912 = (((!g2040) & (!g106) & (!sk[87]) & (!g2030) & (g2049) & (!g2054)) + ((!g2040) & (!g106) & (!sk[87]) & (!g2030) & (g2049) & (g2054)) + ((!g2040) & (!g106) & (!sk[87]) & (g2030) & (!g2049) & (!g2054)) + ((!g2040) & (!g106) & (!sk[87]) & (g2030) & (!g2049) & (g2054)) + ((!g2040) & (!g106) & (!sk[87]) & (g2030) & (g2049) & (!g2054)) + ((!g2040) & (!g106) & (!sk[87]) & (g2030) & (g2049) & (g2054)) + ((!g2040) & (!g106) & (sk[87]) & (!g2030) & (!g2049) & (!g2054)) + ((!g2040) & (!g106) & (sk[87]) & (!g2030) & (!g2049) & (g2054)) + ((!g2040) & (!g106) & (sk[87]) & (!g2030) & (g2049) & (!g2054)) + ((!g2040) & (!g106) & (sk[87]) & (!g2030) & (g2049) & (g2054)) + ((!g2040) & (g106) & (!sk[87]) & (!g2030) & (g2049) & (!g2054)) + ((!g2040) & (g106) & (!sk[87]) & (!g2030) & (g2049) & (g2054)) + ((!g2040) & (g106) & (!sk[87]) & (g2030) & (!g2049) & (!g2054)) + ((!g2040) & (g106) & (!sk[87]) & (g2030) & (!g2049) & (g2054)) + ((!g2040) & (g106) & (!sk[87]) & (g2030) & (g2049) & (!g2054)) + ((!g2040) & (g106) & (!sk[87]) & (g2030) & (g2049) & (g2054)) + ((g2040) & (!g106) & (!sk[87]) & (!g2030) & (!g2049) & (!g2054)) + ((g2040) & (!g106) & (!sk[87]) & (!g2030) & (!g2049) & (g2054)) + ((g2040) & (!g106) & (!sk[87]) & (!g2030) & (g2049) & (!g2054)) + ((g2040) & (!g106) & (!sk[87]) & (!g2030) & (g2049) & (g2054)) + ((g2040) & (!g106) & (!sk[87]) & (g2030) & (!g2049) & (!g2054)) + ((g2040) & (!g106) & (!sk[87]) & (g2030) & (!g2049) & (g2054)) + ((g2040) & (!g106) & (!sk[87]) & (g2030) & (g2049) & (!g2054)) + ((g2040) & (!g106) & (!sk[87]) & (g2030) & (g2049) & (g2054)) + ((g2040) & (!g106) & (sk[87]) & (!g2030) & (!g2049) & (!g2054)) + ((g2040) & (!g106) & (sk[87]) & (!g2030) & (!g2049) & (g2054)) + ((g2040) & (!g106) & (sk[87]) & (!g2030) & (g2049) & (!g2054)) + ((g2040) & (!g106) & (sk[87]) & (g2030) & (!g2049) & (!g2054)) + ((g2040) & (!g106) & (sk[87]) & (g2030) & (!g2049) & (g2054)) + ((g2040) & (!g106) & (sk[87]) & (g2030) & (g2049) & (!g2054)) + ((g2040) & (g106) & (!sk[87]) & (!g2030) & (!g2049) & (!g2054)) + ((g2040) & (g106) & (!sk[87]) & (!g2030) & (!g2049) & (g2054)) + ((g2040) & (g106) & (!sk[87]) & (!g2030) & (g2049) & (!g2054)) + ((g2040) & (g106) & (!sk[87]) & (!g2030) & (g2049) & (g2054)) + ((g2040) & (g106) & (!sk[87]) & (g2030) & (!g2049) & (!g2054)) + ((g2040) & (g106) & (!sk[87]) & (g2030) & (!g2049) & (g2054)) + ((g2040) & (g106) & (!sk[87]) & (g2030) & (g2049) & (!g2054)) + ((g2040) & (g106) & (!sk[87]) & (g2030) & (g2049) & (g2054)) + ((g2040) & (g106) & (sk[87]) & (!g2030) & (!g2049) & (!g2054)) + ((g2040) & (g106) & (sk[87]) & (!g2030) & (!g2049) & (g2054)) + ((g2040) & (g106) & (sk[87]) & (!g2030) & (g2049) & (!g2054)) + ((g2040) & (g106) & (sk[87]) & (g2030) & (!g2049) & (!g2054)) + ((g2040) & (g106) & (sk[87]) & (g2030) & (!g2049) & (g2054)) + ((g2040) & (g106) & (sk[87]) & (g2030) & (g2049) & (!g2054)));
	assign g2913 = (((!g2040) & (g2049) & (!sk[88]) & (!g2054)) + ((!g2040) & (g2049) & (!sk[88]) & (g2054)) + ((g2040) & (!g2049) & (!sk[88]) & (!g2054)) + ((g2040) & (!g2049) & (!sk[88]) & (g2054)) + ((g2040) & (g2049) & (!sk[88]) & (!g2054)) + ((g2040) & (g2049) & (!sk[88]) & (g2054)) + ((g2040) & (g2049) & (sk[88]) & (g2054)));
	assign g5056 = (((!g2924) & (!sk[89]) & (g3114) & (!g2914)) + ((!g2924) & (!sk[89]) & (g3114) & (g2914)) + ((!g2924) & (sk[89]) & (!g3114) & (g2914)) + ((!g2924) & (sk[89]) & (g3114) & (g2914)) + ((g2924) & (!sk[89]) & (!g3114) & (!g2914)) + ((g2924) & (!sk[89]) & (!g3114) & (g2914)) + ((g2924) & (!sk[89]) & (g3114) & (!g2914)) + ((g2924) & (!sk[89]) & (g3114) & (g2914)) + ((g2924) & (sk[89]) & (g3114) & (!g2914)) + ((g2924) & (sk[89]) & (g3114) & (g2914)));
	assign g2915 = (((!g2030) & (!g1720) & (!sk[90]) & (!g2913) & (g2914)) + ((!g2030) & (!g1720) & (!sk[90]) & (g2913) & (g2914)) + ((!g2030) & (g1720) & (!sk[90]) & (!g2913) & (!g2914)) + ((!g2030) & (g1720) & (!sk[90]) & (!g2913) & (g2914)) + ((!g2030) & (g1720) & (!sk[90]) & (g2913) & (!g2914)) + ((!g2030) & (g1720) & (!sk[90]) & (g2913) & (g2914)) + ((!g2030) & (g1720) & (sk[90]) & (g2913) & (!g2914)) + ((!g2030) & (g1720) & (sk[90]) & (g2913) & (g2914)) + ((g2030) & (!g1720) & (!sk[90]) & (!g2913) & (!g2914)) + ((g2030) & (!g1720) & (!sk[90]) & (!g2913) & (g2914)) + ((g2030) & (!g1720) & (!sk[90]) & (g2913) & (!g2914)) + ((g2030) & (!g1720) & (!sk[90]) & (g2913) & (g2914)) + ((g2030) & (!g1720) & (sk[90]) & (!g2913) & (g2914)) + ((g2030) & (!g1720) & (sk[90]) & (g2913) & (g2914)) + ((g2030) & (g1720) & (!sk[90]) & (!g2913) & (!g2914)) + ((g2030) & (g1720) & (!sk[90]) & (!g2913) & (g2914)) + ((g2030) & (g1720) & (!sk[90]) & (g2913) & (!g2914)) + ((g2030) & (g1720) & (!sk[90]) & (g2913) & (g2914)) + ((g2030) & (g1720) & (sk[90]) & (!g2913) & (g2914)) + ((g2030) & (g1720) & (sk[90]) & (g2913) & (!g2914)) + ((g2030) & (g1720) & (sk[90]) & (g2913) & (g2914)));
	assign g2916 = (((!g106) & (!g2026) & (!g2910) & (!g2911) & (!g2912) & (!g2915)) + ((!g106) & (!g2026) & (!g2910) & (!g2911) & (g2912) & (!g2915)) + ((!g106) & (!g2026) & (!g2910) & (g2911) & (!g2912) & (!g2915)) + ((!g106) & (!g2026) & (g2910) & (!g2911) & (!g2912) & (!g2915)) + ((!g106) & (!g2026) & (g2910) & (!g2911) & (g2912) & (!g2915)) + ((!g106) & (!g2026) & (g2910) & (g2911) & (!g2912) & (!g2915)) + ((!g106) & (!g2026) & (g2910) & (g2911) & (g2912) & (!g2915)) + ((!g106) & (g2026) & (!g2910) & (!g2911) & (!g2912) & (!g2915)) + ((!g106) & (g2026) & (!g2910) & (g2911) & (!g2912) & (!g2915)) + ((!g106) & (g2026) & (g2910) & (!g2911) & (!g2912) & (!g2915)) + ((!g106) & (g2026) & (g2910) & (g2911) & (!g2912) & (!g2915)) + ((!g106) & (g2026) & (g2910) & (g2911) & (g2912) & (!g2915)) + ((g106) & (!g2026) & (g2910) & (!g2911) & (!g2912) & (!g2915)) + ((g106) & (!g2026) & (g2910) & (!g2911) & (g2912) & (!g2915)) + ((g106) & (!g2026) & (g2910) & (g2911) & (!g2912) & (!g2915)) + ((g106) & (!g2026) & (g2910) & (g2911) & (g2912) & (!g2915)) + ((g106) & (g2026) & (g2910) & (!g2911) & (!g2912) & (!g2915)) + ((g106) & (g2026) & (g2910) & (g2911) & (!g2912) & (!g2915)) + ((g106) & (g2026) & (g2910) & (g2911) & (g2912) & (!g2915)));
	assign g2917 = (((!nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (g2843) & (!g2916)) + ((!nmi_i) & (!g2023) & (!intr_i) & (g2330) & (g2843) & (!g2916)) + ((!nmi_i) & (!g2023) & (intr_i) & (g2330) & (g2843) & (!g2916)));
	assign g2918 = (((!g76) & (!g1620) & (g2028) & (g2036) & (!g2356) & (g2843)) + ((!g76) & (g1620) & (!g2028) & (!g2036) & (g2356) & (g2843)) + ((!g76) & (g1620) & (!g2028) & (g2036) & (g2356) & (g2843)) + ((!g76) & (g1620) & (g2028) & (!g2036) & (g2356) & (g2843)) + ((!g76) & (g1620) & (g2028) & (g2036) & (!g2356) & (g2843)) + ((!g76) & (g1620) & (g2028) & (g2036) & (g2356) & (g2843)) + ((g76) & (!g1620) & (!g2028) & (!g2036) & (!g2356) & (!g2843)) + ((g76) & (!g1620) & (!g2028) & (!g2036) & (!g2356) & (g2843)) + ((g76) & (!g1620) & (!g2028) & (!g2036) & (g2356) & (!g2843)) + ((g76) & (!g1620) & (!g2028) & (!g2036) & (g2356) & (g2843)) + ((g76) & (!g1620) & (!g2028) & (g2036) & (!g2356) & (!g2843)) + ((g76) & (!g1620) & (!g2028) & (g2036) & (!g2356) & (g2843)) + ((g76) & (!g1620) & (!g2028) & (g2036) & (g2356) & (!g2843)) + ((g76) & (!g1620) & (!g2028) & (g2036) & (g2356) & (g2843)) + ((g76) & (!g1620) & (g2028) & (!g2036) & (!g2356) & (!g2843)) + ((g76) & (!g1620) & (g2028) & (!g2036) & (!g2356) & (g2843)) + ((g76) & (!g1620) & (g2028) & (!g2036) & (g2356) & (!g2843)) + ((g76) & (!g1620) & (g2028) & (!g2036) & (g2356) & (g2843)) + ((g76) & (!g1620) & (g2028) & (g2036) & (!g2356) & (!g2843)) + ((g76) & (!g1620) & (g2028) & (g2036) & (!g2356) & (g2843)) + ((g76) & (!g1620) & (g2028) & (g2036) & (g2356) & (!g2843)) + ((g76) & (!g1620) & (g2028) & (g2036) & (g2356) & (g2843)) + ((g76) & (g1620) & (!g2028) & (!g2036) & (!g2356) & (!g2843)) + ((g76) & (g1620) & (!g2028) & (!g2036) & (!g2356) & (g2843)) + ((g76) & (g1620) & (!g2028) & (!g2036) & (g2356) & (!g2843)) + ((g76) & (g1620) & (!g2028) & (!g2036) & (g2356) & (g2843)) + ((g76) & (g1620) & (!g2028) & (g2036) & (!g2356) & (!g2843)) + ((g76) & (g1620) & (!g2028) & (g2036) & (!g2356) & (g2843)) + ((g76) & (g1620) & (!g2028) & (g2036) & (g2356) & (!g2843)) + ((g76) & (g1620) & (!g2028) & (g2036) & (g2356) & (g2843)) + ((g76) & (g1620) & (g2028) & (!g2036) & (!g2356) & (!g2843)) + ((g76) & (g1620) & (g2028) & (!g2036) & (!g2356) & (g2843)) + ((g76) & (g1620) & (g2028) & (!g2036) & (g2356) & (!g2843)) + ((g76) & (g1620) & (g2028) & (!g2036) & (g2356) & (g2843)) + ((g76) & (g1620) & (g2028) & (g2036) & (!g2356) & (!g2843)) + ((g76) & (g1620) & (g2028) & (g2036) & (!g2356) & (g2843)) + ((g76) & (g1620) & (g2028) & (g2036) & (g2356) & (!g2843)) + ((g76) & (g1620) & (g2028) & (g2036) & (g2356) & (g2843)));
	assign g2919 = (((!nmi_i) & (!g2023) & (!intr_i) & (!g2039) & (!g2056) & (g2843)) + ((!nmi_i) & (!g2023) & (!intr_i) & (!g2039) & (g2056) & (g2843)) + ((!nmi_i) & (!g2023) & (!intr_i) & (g2039) & (!g2056) & (g2843)) + ((!nmi_i) & (!g2023) & (!intr_i) & (g2039) & (g2056) & (g2843)) + ((!nmi_i) & (!g2023) & (intr_i) & (!g2039) & (!g2056) & (g2843)));
	assign g2920 = (((!g2050) & (!g2051) & (!sk[95]) & (!g2052) & (g2053) & (!g2049)) + ((!g2050) & (!g2051) & (!sk[95]) & (!g2052) & (g2053) & (g2049)) + ((!g2050) & (!g2051) & (!sk[95]) & (g2052) & (!g2053) & (!g2049)) + ((!g2050) & (!g2051) & (!sk[95]) & (g2052) & (!g2053) & (g2049)) + ((!g2050) & (!g2051) & (!sk[95]) & (g2052) & (g2053) & (!g2049)) + ((!g2050) & (!g2051) & (!sk[95]) & (g2052) & (g2053) & (g2049)) + ((!g2050) & (g2051) & (!sk[95]) & (!g2052) & (g2053) & (!g2049)) + ((!g2050) & (g2051) & (!sk[95]) & (!g2052) & (g2053) & (g2049)) + ((!g2050) & (g2051) & (!sk[95]) & (g2052) & (!g2053) & (!g2049)) + ((!g2050) & (g2051) & (!sk[95]) & (g2052) & (!g2053) & (g2049)) + ((!g2050) & (g2051) & (!sk[95]) & (g2052) & (g2053) & (!g2049)) + ((!g2050) & (g2051) & (!sk[95]) & (g2052) & (g2053) & (g2049)) + ((g2050) & (!g2051) & (!sk[95]) & (!g2052) & (!g2053) & (!g2049)) + ((g2050) & (!g2051) & (!sk[95]) & (!g2052) & (!g2053) & (g2049)) + ((g2050) & (!g2051) & (!sk[95]) & (!g2052) & (g2053) & (!g2049)) + ((g2050) & (!g2051) & (!sk[95]) & (!g2052) & (g2053) & (g2049)) + ((g2050) & (!g2051) & (!sk[95]) & (g2052) & (!g2053) & (!g2049)) + ((g2050) & (!g2051) & (!sk[95]) & (g2052) & (!g2053) & (g2049)) + ((g2050) & (!g2051) & (!sk[95]) & (g2052) & (g2053) & (!g2049)) + ((g2050) & (!g2051) & (!sk[95]) & (g2052) & (g2053) & (g2049)) + ((g2050) & (g2051) & (!sk[95]) & (!g2052) & (!g2053) & (!g2049)) + ((g2050) & (g2051) & (!sk[95]) & (!g2052) & (!g2053) & (g2049)) + ((g2050) & (g2051) & (!sk[95]) & (!g2052) & (g2053) & (!g2049)) + ((g2050) & (g2051) & (!sk[95]) & (!g2052) & (g2053) & (g2049)) + ((g2050) & (g2051) & (!sk[95]) & (g2052) & (!g2053) & (!g2049)) + ((g2050) & (g2051) & (!sk[95]) & (g2052) & (!g2053) & (g2049)) + ((g2050) & (g2051) & (!sk[95]) & (g2052) & (g2053) & (!g2049)) + ((g2050) & (g2051) & (!sk[95]) & (g2052) & (g2053) & (g2049)) + ((g2050) & (g2051) & (sk[95]) & (g2052) & (!g2053) & (g2049)));
	assign g2921 = (((!sk[96]) & (!g2059) & (!g2040) & (!g2028) & (g2919) & (!g2920)) + ((!sk[96]) & (!g2059) & (!g2040) & (!g2028) & (g2919) & (g2920)) + ((!sk[96]) & (!g2059) & (!g2040) & (g2028) & (!g2919) & (!g2920)) + ((!sk[96]) & (!g2059) & (!g2040) & (g2028) & (!g2919) & (g2920)) + ((!sk[96]) & (!g2059) & (!g2040) & (g2028) & (g2919) & (!g2920)) + ((!sk[96]) & (!g2059) & (!g2040) & (g2028) & (g2919) & (g2920)) + ((!sk[96]) & (!g2059) & (g2040) & (!g2028) & (g2919) & (!g2920)) + ((!sk[96]) & (!g2059) & (g2040) & (!g2028) & (g2919) & (g2920)) + ((!sk[96]) & (!g2059) & (g2040) & (g2028) & (!g2919) & (!g2920)) + ((!sk[96]) & (!g2059) & (g2040) & (g2028) & (!g2919) & (g2920)) + ((!sk[96]) & (!g2059) & (g2040) & (g2028) & (g2919) & (!g2920)) + ((!sk[96]) & (!g2059) & (g2040) & (g2028) & (g2919) & (g2920)) + ((!sk[96]) & (g2059) & (!g2040) & (!g2028) & (!g2919) & (!g2920)) + ((!sk[96]) & (g2059) & (!g2040) & (!g2028) & (!g2919) & (g2920)) + ((!sk[96]) & (g2059) & (!g2040) & (!g2028) & (g2919) & (!g2920)) + ((!sk[96]) & (g2059) & (!g2040) & (!g2028) & (g2919) & (g2920)) + ((!sk[96]) & (g2059) & (!g2040) & (g2028) & (!g2919) & (!g2920)) + ((!sk[96]) & (g2059) & (!g2040) & (g2028) & (!g2919) & (g2920)) + ((!sk[96]) & (g2059) & (!g2040) & (g2028) & (g2919) & (!g2920)) + ((!sk[96]) & (g2059) & (!g2040) & (g2028) & (g2919) & (g2920)) + ((!sk[96]) & (g2059) & (g2040) & (!g2028) & (!g2919) & (!g2920)) + ((!sk[96]) & (g2059) & (g2040) & (!g2028) & (!g2919) & (g2920)) + ((!sk[96]) & (g2059) & (g2040) & (!g2028) & (g2919) & (!g2920)) + ((!sk[96]) & (g2059) & (g2040) & (!g2028) & (g2919) & (g2920)) + ((!sk[96]) & (g2059) & (g2040) & (g2028) & (!g2919) & (!g2920)) + ((!sk[96]) & (g2059) & (g2040) & (g2028) & (!g2919) & (g2920)) + ((!sk[96]) & (g2059) & (g2040) & (g2028) & (g2919) & (!g2920)) + ((!sk[96]) & (g2059) & (g2040) & (g2028) & (g2919) & (g2920)) + ((sk[96]) & (g2059) & (!g2040) & (!g2028) & (!g2919) & (!g2920)) + ((sk[96]) & (g2059) & (!g2040) & (!g2028) & (!g2919) & (g2920)) + ((sk[96]) & (g2059) & (!g2040) & (g2028) & (!g2919) & (!g2920)) + ((sk[96]) & (g2059) & (!g2040) & (g2028) & (!g2919) & (g2920)) + ((sk[96]) & (g2059) & (g2040) & (!g2028) & (!g2919) & (!g2920)) + ((sk[96]) & (g2059) & (g2040) & (!g2028) & (!g2919) & (g2920)) + ((sk[96]) & (g2059) & (g2040) & (!g2028) & (g2919) & (g2920)) + ((sk[96]) & (g2059) & (g2040) & (g2028) & (!g2919) & (!g2920)) + ((sk[96]) & (g2059) & (g2040) & (g2028) & (!g2919) & (g2920)));
	assign g2922 = (((!g1632) & (!nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (!g2843)) + ((!g1632) & (!nmi_i) & (!g2023) & (intr_i) & (!g2330) & (!g2843)) + ((!g1632) & (!nmi_i) & (!g2023) & (intr_i) & (!g2330) & (g2843)) + ((!g1632) & (!nmi_i) & (g2023) & (!intr_i) & (!g2330) & (!g2843)) + ((!g1632) & (!nmi_i) & (g2023) & (!intr_i) & (!g2330) & (g2843)) + ((!g1632) & (!nmi_i) & (g2023) & (intr_i) & (!g2330) & (!g2843)) + ((!g1632) & (!nmi_i) & (g2023) & (intr_i) & (!g2330) & (g2843)) + ((!g1632) & (nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (!g2843)) + ((!g1632) & (nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (g2843)) + ((!g1632) & (nmi_i) & (!g2023) & (intr_i) & (!g2330) & (!g2843)) + ((!g1632) & (nmi_i) & (!g2023) & (intr_i) & (!g2330) & (g2843)) + ((!g1632) & (nmi_i) & (g2023) & (!intr_i) & (!g2330) & (!g2843)) + ((!g1632) & (nmi_i) & (g2023) & (!intr_i) & (!g2330) & (g2843)) + ((!g1632) & (nmi_i) & (g2023) & (intr_i) & (!g2330) & (!g2843)) + ((!g1632) & (nmi_i) & (g2023) & (intr_i) & (!g2330) & (g2843)) + ((g1632) & (!nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (!g2843)) + ((g1632) & (!nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (g2843)) + ((g1632) & (!nmi_i) & (!g2023) & (!intr_i) & (g2330) & (g2843)) + ((g1632) & (!nmi_i) & (!g2023) & (intr_i) & (!g2330) & (!g2843)) + ((g1632) & (!nmi_i) & (!g2023) & (intr_i) & (!g2330) & (g2843)) + ((g1632) & (!nmi_i) & (!g2023) & (intr_i) & (g2330) & (g2843)) + ((g1632) & (!nmi_i) & (g2023) & (!intr_i) & (!g2330) & (!g2843)) + ((g1632) & (!nmi_i) & (g2023) & (!intr_i) & (!g2330) & (g2843)) + ((g1632) & (!nmi_i) & (g2023) & (intr_i) & (!g2330) & (!g2843)) + ((g1632) & (!nmi_i) & (g2023) & (intr_i) & (!g2330) & (g2843)) + ((g1632) & (nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (!g2843)) + ((g1632) & (nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (g2843)) + ((g1632) & (nmi_i) & (!g2023) & (intr_i) & (!g2330) & (!g2843)) + ((g1632) & (nmi_i) & (!g2023) & (intr_i) & (!g2330) & (g2843)) + ((g1632) & (nmi_i) & (g2023) & (!intr_i) & (!g2330) & (!g2843)) + ((g1632) & (nmi_i) & (g2023) & (!intr_i) & (!g2330) & (g2843)) + ((g1632) & (nmi_i) & (g2023) & (intr_i) & (!g2330) & (!g2843)) + ((g1632) & (nmi_i) & (g2023) & (intr_i) & (!g2330) & (g2843)));
	assign g2923 = (((!sk[98]) & (!g2050) & (!g2051) & (!g2052) & (g2053) & (!g2049)) + ((!sk[98]) & (!g2050) & (!g2051) & (!g2052) & (g2053) & (g2049)) + ((!sk[98]) & (!g2050) & (!g2051) & (g2052) & (!g2053) & (!g2049)) + ((!sk[98]) & (!g2050) & (!g2051) & (g2052) & (!g2053) & (g2049)) + ((!sk[98]) & (!g2050) & (!g2051) & (g2052) & (g2053) & (!g2049)) + ((!sk[98]) & (!g2050) & (!g2051) & (g2052) & (g2053) & (g2049)) + ((!sk[98]) & (!g2050) & (g2051) & (!g2052) & (g2053) & (!g2049)) + ((!sk[98]) & (!g2050) & (g2051) & (!g2052) & (g2053) & (g2049)) + ((!sk[98]) & (!g2050) & (g2051) & (g2052) & (!g2053) & (!g2049)) + ((!sk[98]) & (!g2050) & (g2051) & (g2052) & (!g2053) & (g2049)) + ((!sk[98]) & (!g2050) & (g2051) & (g2052) & (g2053) & (!g2049)) + ((!sk[98]) & (!g2050) & (g2051) & (g2052) & (g2053) & (g2049)) + ((!sk[98]) & (g2050) & (!g2051) & (!g2052) & (!g2053) & (!g2049)) + ((!sk[98]) & (g2050) & (!g2051) & (!g2052) & (!g2053) & (g2049)) + ((!sk[98]) & (g2050) & (!g2051) & (!g2052) & (g2053) & (!g2049)) + ((!sk[98]) & (g2050) & (!g2051) & (!g2052) & (g2053) & (g2049)) + ((!sk[98]) & (g2050) & (!g2051) & (g2052) & (!g2053) & (!g2049)) + ((!sk[98]) & (g2050) & (!g2051) & (g2052) & (!g2053) & (g2049)) + ((!sk[98]) & (g2050) & (!g2051) & (g2052) & (g2053) & (!g2049)) + ((!sk[98]) & (g2050) & (!g2051) & (g2052) & (g2053) & (g2049)) + ((!sk[98]) & (g2050) & (g2051) & (!g2052) & (!g2053) & (!g2049)) + ((!sk[98]) & (g2050) & (g2051) & (!g2052) & (!g2053) & (g2049)) + ((!sk[98]) & (g2050) & (g2051) & (!g2052) & (g2053) & (!g2049)) + ((!sk[98]) & (g2050) & (g2051) & (!g2052) & (g2053) & (g2049)) + ((!sk[98]) & (g2050) & (g2051) & (g2052) & (!g2053) & (!g2049)) + ((!sk[98]) & (g2050) & (g2051) & (g2052) & (!g2053) & (g2049)) + ((!sk[98]) & (g2050) & (g2051) & (g2052) & (g2053) & (!g2049)) + ((!sk[98]) & (g2050) & (g2051) & (g2052) & (g2053) & (g2049)) + ((sk[98]) & (g2050) & (g2051) & (!g2052) & (g2053) & (g2049)));
	assign g2924 = (((!g2059) & (!g2040) & (!sk[99]) & (!g2028) & (g2919) & (!g2923)) + ((!g2059) & (!g2040) & (!sk[99]) & (!g2028) & (g2919) & (g2923)) + ((!g2059) & (!g2040) & (!sk[99]) & (g2028) & (!g2919) & (!g2923)) + ((!g2059) & (!g2040) & (!sk[99]) & (g2028) & (!g2919) & (g2923)) + ((!g2059) & (!g2040) & (!sk[99]) & (g2028) & (g2919) & (!g2923)) + ((!g2059) & (!g2040) & (!sk[99]) & (g2028) & (g2919) & (g2923)) + ((!g2059) & (g2040) & (!sk[99]) & (!g2028) & (g2919) & (!g2923)) + ((!g2059) & (g2040) & (!sk[99]) & (!g2028) & (g2919) & (g2923)) + ((!g2059) & (g2040) & (!sk[99]) & (g2028) & (!g2919) & (!g2923)) + ((!g2059) & (g2040) & (!sk[99]) & (g2028) & (!g2919) & (g2923)) + ((!g2059) & (g2040) & (!sk[99]) & (g2028) & (g2919) & (!g2923)) + ((!g2059) & (g2040) & (!sk[99]) & (g2028) & (g2919) & (g2923)) + ((g2059) & (!g2040) & (!sk[99]) & (!g2028) & (!g2919) & (!g2923)) + ((g2059) & (!g2040) & (!sk[99]) & (!g2028) & (!g2919) & (g2923)) + ((g2059) & (!g2040) & (!sk[99]) & (!g2028) & (g2919) & (!g2923)) + ((g2059) & (!g2040) & (!sk[99]) & (!g2028) & (g2919) & (g2923)) + ((g2059) & (!g2040) & (!sk[99]) & (g2028) & (!g2919) & (!g2923)) + ((g2059) & (!g2040) & (!sk[99]) & (g2028) & (!g2919) & (g2923)) + ((g2059) & (!g2040) & (!sk[99]) & (g2028) & (g2919) & (!g2923)) + ((g2059) & (!g2040) & (!sk[99]) & (g2028) & (g2919) & (g2923)) + ((g2059) & (!g2040) & (sk[99]) & (!g2028) & (!g2919) & (!g2923)) + ((g2059) & (!g2040) & (sk[99]) & (!g2028) & (!g2919) & (g2923)) + ((g2059) & (!g2040) & (sk[99]) & (g2028) & (!g2919) & (!g2923)) + ((g2059) & (!g2040) & (sk[99]) & (g2028) & (!g2919) & (g2923)) + ((g2059) & (g2040) & (!sk[99]) & (!g2028) & (!g2919) & (!g2923)) + ((g2059) & (g2040) & (!sk[99]) & (!g2028) & (!g2919) & (g2923)) + ((g2059) & (g2040) & (!sk[99]) & (!g2028) & (g2919) & (!g2923)) + ((g2059) & (g2040) & (!sk[99]) & (!g2028) & (g2919) & (g2923)) + ((g2059) & (g2040) & (!sk[99]) & (g2028) & (!g2919) & (!g2923)) + ((g2059) & (g2040) & (!sk[99]) & (g2028) & (!g2919) & (g2923)) + ((g2059) & (g2040) & (!sk[99]) & (g2028) & (g2919) & (!g2923)) + ((g2059) & (g2040) & (!sk[99]) & (g2028) & (g2919) & (g2923)) + ((g2059) & (g2040) & (sk[99]) & (!g2028) & (!g2919) & (!g2923)) + ((g2059) & (g2040) & (sk[99]) & (!g2028) & (!g2919) & (g2923)) + ((g2059) & (g2040) & (sk[99]) & (!g2028) & (g2919) & (g2923)) + ((g2059) & (g2040) & (sk[99]) & (g2028) & (!g2919) & (!g2923)) + ((g2059) & (g2040) & (sk[99]) & (g2028) & (!g2919) & (g2923)));
	assign g2925 = (((!nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (sk[100]) & (g2843)) + ((!nmi_i) & (!g2023) & (!intr_i) & (g2330) & (!sk[100]) & (!g2843)) + ((!nmi_i) & (!g2023) & (!intr_i) & (g2330) & (!sk[100]) & (g2843)) + ((!nmi_i) & (!g2023) & (intr_i) & (!g2330) & (!sk[100]) & (!g2843)) + ((!nmi_i) & (!g2023) & (intr_i) & (!g2330) & (!sk[100]) & (g2843)) + ((!nmi_i) & (!g2023) & (intr_i) & (g2330) & (!sk[100]) & (!g2843)) + ((!nmi_i) & (!g2023) & (intr_i) & (g2330) & (!sk[100]) & (g2843)) + ((!nmi_i) & (g2023) & (!intr_i) & (g2330) & (!sk[100]) & (!g2843)) + ((!nmi_i) & (g2023) & (!intr_i) & (g2330) & (!sk[100]) & (g2843)) + ((!nmi_i) & (g2023) & (intr_i) & (!g2330) & (!sk[100]) & (!g2843)) + ((!nmi_i) & (g2023) & (intr_i) & (!g2330) & (!sk[100]) & (g2843)) + ((!nmi_i) & (g2023) & (intr_i) & (g2330) & (!sk[100]) & (!g2843)) + ((!nmi_i) & (g2023) & (intr_i) & (g2330) & (!sk[100]) & (g2843)) + ((nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (!sk[100]) & (!g2843)) + ((nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (!sk[100]) & (g2843)) + ((nmi_i) & (!g2023) & (!intr_i) & (g2330) & (!sk[100]) & (!g2843)) + ((nmi_i) & (!g2023) & (!intr_i) & (g2330) & (!sk[100]) & (g2843)) + ((nmi_i) & (!g2023) & (intr_i) & (!g2330) & (!sk[100]) & (!g2843)) + ((nmi_i) & (!g2023) & (intr_i) & (!g2330) & (!sk[100]) & (g2843)) + ((nmi_i) & (!g2023) & (intr_i) & (g2330) & (!sk[100]) & (!g2843)) + ((nmi_i) & (!g2023) & (intr_i) & (g2330) & (!sk[100]) & (g2843)) + ((nmi_i) & (g2023) & (!intr_i) & (!g2330) & (!sk[100]) & (!g2843)) + ((nmi_i) & (g2023) & (!intr_i) & (!g2330) & (!sk[100]) & (g2843)) + ((nmi_i) & (g2023) & (!intr_i) & (g2330) & (!sk[100]) & (!g2843)) + ((nmi_i) & (g2023) & (!intr_i) & (g2330) & (!sk[100]) & (g2843)) + ((nmi_i) & (g2023) & (intr_i) & (!g2330) & (!sk[100]) & (!g2843)) + ((nmi_i) & (g2023) & (intr_i) & (!g2330) & (!sk[100]) & (g2843)) + ((nmi_i) & (g2023) & (intr_i) & (g2330) & (!sk[100]) & (!g2843)) + ((nmi_i) & (g2023) & (intr_i) & (g2330) & (!sk[100]) & (g2843)));
	assign g2926 = (((!g77) & (!g1604) & (g2028) & (g2061) & (!g2356) & (g2843)) + ((!g77) & (g1604) & (!g2028) & (!g2061) & (g2356) & (g2843)) + ((!g77) & (g1604) & (!g2028) & (g2061) & (g2356) & (g2843)) + ((!g77) & (g1604) & (g2028) & (!g2061) & (g2356) & (g2843)) + ((!g77) & (g1604) & (g2028) & (g2061) & (!g2356) & (g2843)) + ((!g77) & (g1604) & (g2028) & (g2061) & (g2356) & (g2843)) + ((g77) & (!g1604) & (!g2028) & (!g2061) & (!g2356) & (!g2843)) + ((g77) & (!g1604) & (!g2028) & (!g2061) & (!g2356) & (g2843)) + ((g77) & (!g1604) & (!g2028) & (!g2061) & (g2356) & (!g2843)) + ((g77) & (!g1604) & (!g2028) & (!g2061) & (g2356) & (g2843)) + ((g77) & (!g1604) & (!g2028) & (g2061) & (!g2356) & (!g2843)) + ((g77) & (!g1604) & (!g2028) & (g2061) & (!g2356) & (g2843)) + ((g77) & (!g1604) & (!g2028) & (g2061) & (g2356) & (!g2843)) + ((g77) & (!g1604) & (!g2028) & (g2061) & (g2356) & (g2843)) + ((g77) & (!g1604) & (g2028) & (!g2061) & (!g2356) & (!g2843)) + ((g77) & (!g1604) & (g2028) & (!g2061) & (!g2356) & (g2843)) + ((g77) & (!g1604) & (g2028) & (!g2061) & (g2356) & (!g2843)) + ((g77) & (!g1604) & (g2028) & (!g2061) & (g2356) & (g2843)) + ((g77) & (!g1604) & (g2028) & (g2061) & (!g2356) & (!g2843)) + ((g77) & (!g1604) & (g2028) & (g2061) & (!g2356) & (g2843)) + ((g77) & (!g1604) & (g2028) & (g2061) & (g2356) & (!g2843)) + ((g77) & (!g1604) & (g2028) & (g2061) & (g2356) & (g2843)) + ((g77) & (g1604) & (!g2028) & (!g2061) & (!g2356) & (!g2843)) + ((g77) & (g1604) & (!g2028) & (!g2061) & (!g2356) & (g2843)) + ((g77) & (g1604) & (!g2028) & (!g2061) & (g2356) & (!g2843)) + ((g77) & (g1604) & (!g2028) & (!g2061) & (g2356) & (g2843)) + ((g77) & (g1604) & (!g2028) & (g2061) & (!g2356) & (!g2843)) + ((g77) & (g1604) & (!g2028) & (g2061) & (!g2356) & (g2843)) + ((g77) & (g1604) & (!g2028) & (g2061) & (g2356) & (!g2843)) + ((g77) & (g1604) & (!g2028) & (g2061) & (g2356) & (g2843)) + ((g77) & (g1604) & (g2028) & (!g2061) & (!g2356) & (!g2843)) + ((g77) & (g1604) & (g2028) & (!g2061) & (!g2356) & (g2843)) + ((g77) & (g1604) & (g2028) & (!g2061) & (g2356) & (!g2843)) + ((g77) & (g1604) & (g2028) & (!g2061) & (g2356) & (g2843)) + ((g77) & (g1604) & (g2028) & (g2061) & (!g2356) & (!g2843)) + ((g77) & (g1604) & (g2028) & (g2061) & (!g2356) & (g2843)) + ((g77) & (g1604) & (g2028) & (g2061) & (g2356) & (!g2843)) + ((g77) & (g1604) & (g2028) & (g2061) & (g2356) & (g2843)));
	assign g2927 = (((!g1632) & (!g2028) & (!g141) & (!g2067) & (!g2356) & (!g2843)) + ((!g1632) & (!g2028) & (!g141) & (!g2067) & (!g2356) & (g2843)) + ((!g1632) & (!g2028) & (!g141) & (!g2067) & (g2356) & (!g2843)) + ((!g1632) & (!g2028) & (!g141) & (g2067) & (!g2356) & (!g2843)) + ((!g1632) & (!g2028) & (!g141) & (g2067) & (!g2356) & (g2843)) + ((!g1632) & (!g2028) & (!g141) & (g2067) & (g2356) & (!g2843)) + ((!g1632) & (g2028) & (!g141) & (!g2067) & (!g2356) & (!g2843)) + ((!g1632) & (g2028) & (!g141) & (!g2067) & (g2356) & (!g2843)) + ((!g1632) & (g2028) & (!g141) & (g2067) & (!g2356) & (!g2843)) + ((!g1632) & (g2028) & (!g141) & (g2067) & (!g2356) & (g2843)) + ((!g1632) & (g2028) & (!g141) & (g2067) & (g2356) & (!g2843)) + ((!g1632) & (g2028) & (g141) & (g2067) & (!g2356) & (g2843)) + ((g1632) & (!g2028) & (!g141) & (!g2067) & (!g2356) & (!g2843)) + ((g1632) & (!g2028) & (!g141) & (!g2067) & (!g2356) & (g2843)) + ((g1632) & (!g2028) & (!g141) & (!g2067) & (g2356) & (!g2843)) + ((g1632) & (!g2028) & (!g141) & (!g2067) & (g2356) & (g2843)) + ((g1632) & (!g2028) & (!g141) & (g2067) & (!g2356) & (!g2843)) + ((g1632) & (!g2028) & (!g141) & (g2067) & (!g2356) & (g2843)) + ((g1632) & (!g2028) & (!g141) & (g2067) & (g2356) & (!g2843)) + ((g1632) & (!g2028) & (!g141) & (g2067) & (g2356) & (g2843)) + ((g1632) & (!g2028) & (g141) & (!g2067) & (g2356) & (g2843)) + ((g1632) & (!g2028) & (g141) & (g2067) & (g2356) & (g2843)) + ((g1632) & (g2028) & (!g141) & (!g2067) & (!g2356) & (!g2843)) + ((g1632) & (g2028) & (!g141) & (!g2067) & (g2356) & (!g2843)) + ((g1632) & (g2028) & (!g141) & (!g2067) & (g2356) & (g2843)) + ((g1632) & (g2028) & (!g141) & (g2067) & (!g2356) & (!g2843)) + ((g1632) & (g2028) & (!g141) & (g2067) & (!g2356) & (g2843)) + ((g1632) & (g2028) & (!g141) & (g2067) & (g2356) & (!g2843)) + ((g1632) & (g2028) & (!g141) & (g2067) & (g2356) & (g2843)) + ((g1632) & (g2028) & (g141) & (!g2067) & (g2356) & (g2843)) + ((g1632) & (g2028) & (g141) & (g2067) & (!g2356) & (g2843)) + ((g1632) & (g2028) & (g141) & (g2067) & (g2356) & (g2843)));
	assign g2928 = (((g78) & (!g79) & (g80) & (!g81) & (g82) & (g83)));
	assign g2929 = (((!sk[104]) & (!g2024) & (!g77) & (!g142) & (g167) & (!g187)) + ((!sk[104]) & (!g2024) & (!g77) & (!g142) & (g167) & (g187)) + ((!sk[104]) & (!g2024) & (!g77) & (g142) & (!g167) & (!g187)) + ((!sk[104]) & (!g2024) & (!g77) & (g142) & (!g167) & (g187)) + ((!sk[104]) & (!g2024) & (!g77) & (g142) & (g167) & (!g187)) + ((!sk[104]) & (!g2024) & (!g77) & (g142) & (g167) & (g187)) + ((!sk[104]) & (!g2024) & (g77) & (!g142) & (g167) & (!g187)) + ((!sk[104]) & (!g2024) & (g77) & (!g142) & (g167) & (g187)) + ((!sk[104]) & (!g2024) & (g77) & (g142) & (!g167) & (!g187)) + ((!sk[104]) & (!g2024) & (g77) & (g142) & (!g167) & (g187)) + ((!sk[104]) & (!g2024) & (g77) & (g142) & (g167) & (!g187)) + ((!sk[104]) & (!g2024) & (g77) & (g142) & (g167) & (g187)) + ((!sk[104]) & (g2024) & (!g77) & (!g142) & (!g167) & (!g187)) + ((!sk[104]) & (g2024) & (!g77) & (!g142) & (!g167) & (g187)) + ((!sk[104]) & (g2024) & (!g77) & (!g142) & (g167) & (!g187)) + ((!sk[104]) & (g2024) & (!g77) & (!g142) & (g167) & (g187)) + ((!sk[104]) & (g2024) & (!g77) & (g142) & (!g167) & (!g187)) + ((!sk[104]) & (g2024) & (!g77) & (g142) & (!g167) & (g187)) + ((!sk[104]) & (g2024) & (!g77) & (g142) & (g167) & (!g187)) + ((!sk[104]) & (g2024) & (!g77) & (g142) & (g167) & (g187)) + ((!sk[104]) & (g2024) & (g77) & (!g142) & (!g167) & (!g187)) + ((!sk[104]) & (g2024) & (g77) & (!g142) & (!g167) & (g187)) + ((!sk[104]) & (g2024) & (g77) & (!g142) & (g167) & (!g187)) + ((!sk[104]) & (g2024) & (g77) & (!g142) & (g167) & (g187)) + ((!sk[104]) & (g2024) & (g77) & (g142) & (!g167) & (!g187)) + ((!sk[104]) & (g2024) & (g77) & (g142) & (!g167) & (g187)) + ((!sk[104]) & (g2024) & (g77) & (g142) & (g167) & (!g187)) + ((!sk[104]) & (g2024) & (g77) & (g142) & (g167) & (g187)) + ((sk[104]) & (!g2024) & (!g77) & (!g142) & (!g167) & (g187)) + ((sk[104]) & (!g2024) & (!g77) & (!g142) & (g167) & (g187)) + ((sk[104]) & (!g2024) & (!g77) & (g142) & (g167) & (!g187)) + ((sk[104]) & (!g2024) & (!g77) & (g142) & (g167) & (g187)) + ((sk[104]) & (!g2024) & (g77) & (!g142) & (!g167) & (g187)) + ((sk[104]) & (!g2024) & (g77) & (!g142) & (g167) & (g187)) + ((sk[104]) & (!g2024) & (g77) & (g142) & (g167) & (!g187)) + ((sk[104]) & (!g2024) & (g77) & (g142) & (g167) & (g187)) + ((sk[104]) & (g2024) & (g77) & (!g142) & (!g167) & (!g187)) + ((sk[104]) & (g2024) & (g77) & (!g142) & (!g167) & (g187)) + ((sk[104]) & (g2024) & (g77) & (!g142) & (g167) & (!g187)) + ((sk[104]) & (g2024) & (g77) & (!g142) & (g167) & (g187)) + ((sk[104]) & (g2024) & (g77) & (g142) & (!g167) & (!g187)) + ((sk[104]) & (g2024) & (g77) & (g142) & (!g167) & (g187)) + ((sk[104]) & (g2024) & (g77) & (g142) & (g167) & (!g187)) + ((sk[104]) & (g2024) & (g77) & (g142) & (g167) & (g187)));
	assign g2930 = (((!g80) & (!sk[105]) & (!g81) & (!g82) & (g83)) + ((!g80) & (!sk[105]) & (!g81) & (g82) & (g83)) + ((!g80) & (!sk[105]) & (g81) & (!g82) & (!g83)) + ((!g80) & (!sk[105]) & (g81) & (!g82) & (g83)) + ((!g80) & (!sk[105]) & (g81) & (g82) & (!g83)) + ((!g80) & (!sk[105]) & (g81) & (g82) & (g83)) + ((g80) & (!sk[105]) & (!g81) & (!g82) & (!g83)) + ((g80) & (!sk[105]) & (!g81) & (!g82) & (g83)) + ((g80) & (!sk[105]) & (!g81) & (g82) & (!g83)) + ((g80) & (!sk[105]) & (!g81) & (g82) & (g83)) + ((g80) & (!sk[105]) & (g81) & (!g82) & (!g83)) + ((g80) & (!sk[105]) & (g81) & (!g82) & (g83)) + ((g80) & (!sk[105]) & (g81) & (g82) & (!g83)) + ((g80) & (!sk[105]) & (g81) & (g82) & (g83)) + ((g80) & (sk[105]) & (!g81) & (g82) & (g83)));
	assign g2931 = (((g78) & (g79) & (g80) & (!g81) & (!g82) & (g83)));
	assign g2932 = (((!g87) & (!sk[107]) & (!g88) & (!g89) & (g102) & (!g3139)) + ((!g87) & (!sk[107]) & (!g88) & (!g89) & (g102) & (g3139)) + ((!g87) & (!sk[107]) & (!g88) & (g89) & (!g102) & (!g3139)) + ((!g87) & (!sk[107]) & (!g88) & (g89) & (!g102) & (g3139)) + ((!g87) & (!sk[107]) & (!g88) & (g89) & (g102) & (!g3139)) + ((!g87) & (!sk[107]) & (!g88) & (g89) & (g102) & (g3139)) + ((!g87) & (!sk[107]) & (g88) & (!g89) & (g102) & (!g3139)) + ((!g87) & (!sk[107]) & (g88) & (!g89) & (g102) & (g3139)) + ((!g87) & (!sk[107]) & (g88) & (g89) & (!g102) & (!g3139)) + ((!g87) & (!sk[107]) & (g88) & (g89) & (!g102) & (g3139)) + ((!g87) & (!sk[107]) & (g88) & (g89) & (g102) & (!g3139)) + ((!g87) & (!sk[107]) & (g88) & (g89) & (g102) & (g3139)) + ((!g87) & (sk[107]) & (!g88) & (!g89) & (!g102) & (g3139)) + ((!g87) & (sk[107]) & (!g88) & (!g89) & (g102) & (g3139)) + ((!g87) & (sk[107]) & (!g88) & (g89) & (!g102) & (g3139)) + ((!g87) & (sk[107]) & (!g88) & (g89) & (g102) & (g3139)) + ((!g87) & (sk[107]) & (g88) & (!g89) & (!g102) & (g3139)) + ((!g87) & (sk[107]) & (g88) & (g89) & (!g102) & (g3139)) + ((!g87) & (sk[107]) & (g88) & (g89) & (g102) & (g3139)) + ((g87) & (!sk[107]) & (!g88) & (!g89) & (!g102) & (!g3139)) + ((g87) & (!sk[107]) & (!g88) & (!g89) & (!g102) & (g3139)) + ((g87) & (!sk[107]) & (!g88) & (!g89) & (g102) & (!g3139)) + ((g87) & (!sk[107]) & (!g88) & (!g89) & (g102) & (g3139)) + ((g87) & (!sk[107]) & (!g88) & (g89) & (!g102) & (!g3139)) + ((g87) & (!sk[107]) & (!g88) & (g89) & (!g102) & (g3139)) + ((g87) & (!sk[107]) & (!g88) & (g89) & (g102) & (!g3139)) + ((g87) & (!sk[107]) & (!g88) & (g89) & (g102) & (g3139)) + ((g87) & (!sk[107]) & (g88) & (!g89) & (!g102) & (!g3139)) + ((g87) & (!sk[107]) & (g88) & (!g89) & (!g102) & (g3139)) + ((g87) & (!sk[107]) & (g88) & (!g89) & (g102) & (!g3139)) + ((g87) & (!sk[107]) & (g88) & (!g89) & (g102) & (g3139)) + ((g87) & (!sk[107]) & (g88) & (g89) & (!g102) & (!g3139)) + ((g87) & (!sk[107]) & (g88) & (g89) & (!g102) & (g3139)) + ((g87) & (!sk[107]) & (g88) & (g89) & (g102) & (!g3139)) + ((g87) & (!sk[107]) & (g88) & (g89) & (g102) & (g3139)) + ((g87) & (sk[107]) & (!g88) & (!g89) & (!g102) & (g3139)) + ((g87) & (sk[107]) & (!g88) & (!g89) & (g102) & (g3139)) + ((g87) & (sk[107]) & (!g88) & (g89) & (!g102) & (g3139)) + ((g87) & (sk[107]) & (g88) & (!g89) & (!g102) & (g3139)) + ((g87) & (sk[107]) & (g88) & (!g89) & (g102) & (g3139)) + ((g87) & (sk[107]) & (g88) & (g89) & (!g102) & (g3139)) + ((g87) & (sk[107]) & (g88) & (g89) & (g102) & (g3139)));
	assign g2933 = (((!g85) & (!g86) & (!g88) & (g91) & (!sk[108]) & (!g92)) + ((!g85) & (!g86) & (!g88) & (g91) & (!sk[108]) & (g92)) + ((!g85) & (!g86) & (g88) & (!g91) & (!sk[108]) & (!g92)) + ((!g85) & (!g86) & (g88) & (!g91) & (!sk[108]) & (g92)) + ((!g85) & (!g86) & (g88) & (g91) & (!sk[108]) & (!g92)) + ((!g85) & (!g86) & (g88) & (g91) & (!sk[108]) & (g92)) + ((!g85) & (!g86) & (g88) & (g91) & (sk[108]) & (g92)) + ((!g85) & (g86) & (!g88) & (g91) & (!sk[108]) & (!g92)) + ((!g85) & (g86) & (!g88) & (g91) & (!sk[108]) & (g92)) + ((!g85) & (g86) & (g88) & (!g91) & (!sk[108]) & (!g92)) + ((!g85) & (g86) & (g88) & (!g91) & (!sk[108]) & (g92)) + ((!g85) & (g86) & (g88) & (g91) & (!sk[108]) & (!g92)) + ((!g85) & (g86) & (g88) & (g91) & (!sk[108]) & (g92)) + ((g85) & (!g86) & (!g88) & (!g91) & (!sk[108]) & (!g92)) + ((g85) & (!g86) & (!g88) & (!g91) & (!sk[108]) & (g92)) + ((g85) & (!g86) & (!g88) & (g91) & (!sk[108]) & (!g92)) + ((g85) & (!g86) & (!g88) & (g91) & (!sk[108]) & (g92)) + ((g85) & (!g86) & (g88) & (!g91) & (!sk[108]) & (!g92)) + ((g85) & (!g86) & (g88) & (!g91) & (!sk[108]) & (g92)) + ((g85) & (!g86) & (g88) & (g91) & (!sk[108]) & (!g92)) + ((g85) & (!g86) & (g88) & (g91) & (!sk[108]) & (g92)) + ((g85) & (g86) & (!g88) & (!g91) & (!sk[108]) & (!g92)) + ((g85) & (g86) & (!g88) & (!g91) & (!sk[108]) & (g92)) + ((g85) & (g86) & (!g88) & (g91) & (!sk[108]) & (!g92)) + ((g85) & (g86) & (!g88) & (g91) & (!sk[108]) & (g92)) + ((g85) & (g86) & (g88) & (!g91) & (!sk[108]) & (!g92)) + ((g85) & (g86) & (g88) & (!g91) & (!sk[108]) & (g92)) + ((g85) & (g86) & (g88) & (g91) & (!sk[108]) & (!g92)) + ((g85) & (g86) & (g88) & (g91) & (!sk[108]) & (g92)));
	assign g2934 = (((!g87) & (!g89) & (!sk[109]) & (!g90) & (g2933)) + ((!g87) & (!g89) & (!sk[109]) & (g90) & (g2933)) + ((!g87) & (g89) & (!sk[109]) & (!g90) & (!g2933)) + ((!g87) & (g89) & (!sk[109]) & (!g90) & (g2933)) + ((!g87) & (g89) & (!sk[109]) & (g90) & (!g2933)) + ((!g87) & (g89) & (!sk[109]) & (g90) & (g2933)) + ((!g87) & (g89) & (sk[109]) & (g90) & (g2933)) + ((g87) & (!g89) & (!sk[109]) & (!g90) & (!g2933)) + ((g87) & (!g89) & (!sk[109]) & (!g90) & (g2933)) + ((g87) & (!g89) & (!sk[109]) & (g90) & (!g2933)) + ((g87) & (!g89) & (!sk[109]) & (g90) & (g2933)) + ((g87) & (!g89) & (sk[109]) & (!g90) & (g2933)) + ((g87) & (g89) & (!sk[109]) & (!g90) & (!g2933)) + ((g87) & (g89) & (!sk[109]) & (!g90) & (g2933)) + ((g87) & (g89) & (!sk[109]) & (g90) & (!g2933)) + ((g87) & (g89) & (!sk[109]) & (g90) & (g2933)));
	assign g2935 = (((!g2931) & (!sk[110]) & (!g84) & (!g99) & (g2932) & (!g2934)) + ((!g2931) & (!sk[110]) & (!g84) & (!g99) & (g2932) & (g2934)) + ((!g2931) & (!sk[110]) & (!g84) & (g99) & (!g2932) & (!g2934)) + ((!g2931) & (!sk[110]) & (!g84) & (g99) & (!g2932) & (g2934)) + ((!g2931) & (!sk[110]) & (!g84) & (g99) & (g2932) & (!g2934)) + ((!g2931) & (!sk[110]) & (!g84) & (g99) & (g2932) & (g2934)) + ((!g2931) & (!sk[110]) & (g84) & (!g99) & (g2932) & (!g2934)) + ((!g2931) & (!sk[110]) & (g84) & (!g99) & (g2932) & (g2934)) + ((!g2931) & (!sk[110]) & (g84) & (g99) & (!g2932) & (!g2934)) + ((!g2931) & (!sk[110]) & (g84) & (g99) & (!g2932) & (g2934)) + ((!g2931) & (!sk[110]) & (g84) & (g99) & (g2932) & (!g2934)) + ((!g2931) & (!sk[110]) & (g84) & (g99) & (g2932) & (g2934)) + ((!g2931) & (sk[110]) & (!g84) & (!g99) & (!g2932) & (!g2934)) + ((!g2931) & (sk[110]) & (!g84) & (!g99) & (!g2932) & (g2934)) + ((!g2931) & (sk[110]) & (!g84) & (!g99) & (g2932) & (!g2934)) + ((!g2931) & (sk[110]) & (!g84) & (!g99) & (g2932) & (g2934)) + ((!g2931) & (sk[110]) & (g84) & (!g99) & (g2932) & (!g2934)) + ((g2931) & (!sk[110]) & (!g84) & (!g99) & (!g2932) & (!g2934)) + ((g2931) & (!sk[110]) & (!g84) & (!g99) & (!g2932) & (g2934)) + ((g2931) & (!sk[110]) & (!g84) & (!g99) & (g2932) & (!g2934)) + ((g2931) & (!sk[110]) & (!g84) & (!g99) & (g2932) & (g2934)) + ((g2931) & (!sk[110]) & (!g84) & (g99) & (!g2932) & (!g2934)) + ((g2931) & (!sk[110]) & (!g84) & (g99) & (!g2932) & (g2934)) + ((g2931) & (!sk[110]) & (!g84) & (g99) & (g2932) & (!g2934)) + ((g2931) & (!sk[110]) & (!g84) & (g99) & (g2932) & (g2934)) + ((g2931) & (!sk[110]) & (g84) & (!g99) & (!g2932) & (!g2934)) + ((g2931) & (!sk[110]) & (g84) & (!g99) & (!g2932) & (g2934)) + ((g2931) & (!sk[110]) & (g84) & (!g99) & (g2932) & (!g2934)) + ((g2931) & (!sk[110]) & (g84) & (!g99) & (g2932) & (g2934)) + ((g2931) & (!sk[110]) & (g84) & (g99) & (!g2932) & (!g2934)) + ((g2931) & (!sk[110]) & (g84) & (g99) & (!g2932) & (g2934)) + ((g2931) & (!sk[110]) & (g84) & (g99) & (g2932) & (!g2934)) + ((g2931) & (!sk[110]) & (g84) & (g99) & (g2932) & (g2934)));
	assign g2936 = (((!g118) & (!g86) & (!g119) & (!sk[111]) & (g2935)) + ((!g118) & (!g86) & (!g119) & (sk[111]) & (g2935)) + ((!g118) & (!g86) & (g119) & (!sk[111]) & (g2935)) + ((!g118) & (g86) & (!g119) & (!sk[111]) & (!g2935)) + ((!g118) & (g86) & (!g119) & (!sk[111]) & (g2935)) + ((!g118) & (g86) & (!g119) & (sk[111]) & (g2935)) + ((!g118) & (g86) & (g119) & (!sk[111]) & (!g2935)) + ((!g118) & (g86) & (g119) & (!sk[111]) & (g2935)) + ((g118) & (!g86) & (!g119) & (!sk[111]) & (!g2935)) + ((g118) & (!g86) & (!g119) & (!sk[111]) & (g2935)) + ((g118) & (!g86) & (g119) & (!sk[111]) & (!g2935)) + ((g118) & (!g86) & (g119) & (!sk[111]) & (g2935)) + ((g118) & (g86) & (!g119) & (!sk[111]) & (!g2935)) + ((g118) & (g86) & (!g119) & (!sk[111]) & (g2935)) + ((g118) & (g86) & (!g119) & (sk[111]) & (g2935)) + ((g118) & (g86) & (g119) & (!sk[111]) & (!g2935)) + ((g118) & (g86) & (g119) & (!sk[111]) & (g2935)));
	assign g2937 = (((!sk[112]) & (!g118) & (!g85) & (!g86) & (g2936)) + ((!sk[112]) & (!g118) & (!g85) & (g86) & (g2936)) + ((!sk[112]) & (!g118) & (g85) & (!g86) & (!g2936)) + ((!sk[112]) & (!g118) & (g85) & (!g86) & (g2936)) + ((!sk[112]) & (!g118) & (g85) & (g86) & (!g2936)) + ((!sk[112]) & (!g118) & (g85) & (g86) & (g2936)) + ((!sk[112]) & (g118) & (!g85) & (!g86) & (!g2936)) + ((!sk[112]) & (g118) & (!g85) & (!g86) & (g2936)) + ((!sk[112]) & (g118) & (!g85) & (g86) & (!g2936)) + ((!sk[112]) & (g118) & (!g85) & (g86) & (g2936)) + ((!sk[112]) & (g118) & (g85) & (!g86) & (!g2936)) + ((!sk[112]) & (g118) & (g85) & (!g86) & (g2936)) + ((!sk[112]) & (g118) & (g85) & (g86) & (!g2936)) + ((!sk[112]) & (g118) & (g85) & (g86) & (g2936)) + ((sk[112]) & (!g118) & (!g85) & (!g86) & (g2936)) + ((sk[112]) & (!g118) & (!g85) & (g86) & (g2936)) + ((sk[112]) & (!g118) & (g85) & (!g86) & (g2936)) + ((sk[112]) & (!g118) & (g85) & (g86) & (g2936)) + ((sk[112]) & (g118) & (!g85) & (!g86) & (g2936)) + ((sk[112]) & (g118) & (g85) & (!g86) & (g2936)) + ((sk[112]) & (g118) & (g85) & (g86) & (g2936)));
	assign g2938 = (((!g78) & (!sk[113]) & (!g79) & (!g81) & (g2845) & (!g2937)) + ((!g78) & (!sk[113]) & (!g79) & (!g81) & (g2845) & (g2937)) + ((!g78) & (!sk[113]) & (!g79) & (g81) & (!g2845) & (!g2937)) + ((!g78) & (!sk[113]) & (!g79) & (g81) & (!g2845) & (g2937)) + ((!g78) & (!sk[113]) & (!g79) & (g81) & (g2845) & (!g2937)) + ((!g78) & (!sk[113]) & (!g79) & (g81) & (g2845) & (g2937)) + ((!g78) & (!sk[113]) & (g79) & (!g81) & (g2845) & (!g2937)) + ((!g78) & (!sk[113]) & (g79) & (!g81) & (g2845) & (g2937)) + ((!g78) & (!sk[113]) & (g79) & (g81) & (!g2845) & (!g2937)) + ((!g78) & (!sk[113]) & (g79) & (g81) & (!g2845) & (g2937)) + ((!g78) & (!sk[113]) & (g79) & (g81) & (g2845) & (!g2937)) + ((!g78) & (!sk[113]) & (g79) & (g81) & (g2845) & (g2937)) + ((!g78) & (sk[113]) & (!g79) & (!g81) & (!g2845) & (g2937)) + ((!g78) & (sk[113]) & (!g79) & (!g81) & (g2845) & (g2937)) + ((!g78) & (sk[113]) & (!g79) & (g81) & (!g2845) & (g2937)) + ((!g78) & (sk[113]) & (g79) & (!g81) & (!g2845) & (g2937)) + ((!g78) & (sk[113]) & (g79) & (!g81) & (g2845) & (g2937)) + ((!g78) & (sk[113]) & (g79) & (g81) & (!g2845) & (g2937)) + ((!g78) & (sk[113]) & (g79) & (g81) & (g2845) & (g2937)) + ((g78) & (!sk[113]) & (!g79) & (!g81) & (!g2845) & (!g2937)) + ((g78) & (!sk[113]) & (!g79) & (!g81) & (!g2845) & (g2937)) + ((g78) & (!sk[113]) & (!g79) & (!g81) & (g2845) & (!g2937)) + ((g78) & (!sk[113]) & (!g79) & (!g81) & (g2845) & (g2937)) + ((g78) & (!sk[113]) & (!g79) & (g81) & (!g2845) & (!g2937)) + ((g78) & (!sk[113]) & (!g79) & (g81) & (!g2845) & (g2937)) + ((g78) & (!sk[113]) & (!g79) & (g81) & (g2845) & (!g2937)) + ((g78) & (!sk[113]) & (!g79) & (g81) & (g2845) & (g2937)) + ((g78) & (!sk[113]) & (g79) & (!g81) & (!g2845) & (!g2937)) + ((g78) & (!sk[113]) & (g79) & (!g81) & (!g2845) & (g2937)) + ((g78) & (!sk[113]) & (g79) & (!g81) & (g2845) & (!g2937)) + ((g78) & (!sk[113]) & (g79) & (!g81) & (g2845) & (g2937)) + ((g78) & (!sk[113]) & (g79) & (g81) & (!g2845) & (!g2937)) + ((g78) & (!sk[113]) & (g79) & (g81) & (!g2845) & (g2937)) + ((g78) & (!sk[113]) & (g79) & (g81) & (g2845) & (!g2937)) + ((g78) & (!sk[113]) & (g79) & (g81) & (g2845) & (g2937)) + ((g78) & (sk[113]) & (!g79) & (!g81) & (!g2845) & (g2937)) + ((g78) & (sk[113]) & (!g79) & (!g81) & (g2845) & (g2937)) + ((g78) & (sk[113]) & (!g79) & (g81) & (!g2845) & (g2937)) + ((g78) & (sk[113]) & (!g79) & (g81) & (g2845) & (g2937)) + ((g78) & (sk[113]) & (g79) & (!g81) & (!g2845) & (g2937)) + ((g78) & (sk[113]) & (g79) & (g81) & (!g2845) & (g2937)) + ((g78) & (sk[113]) & (g79) & (g81) & (g2845) & (g2937)));
	assign g2939 = (((!g78) & (!g79) & (!g135) & (!g82) & (!g83) & (g2938)) + ((!g78) & (!g79) & (!g135) & (!g82) & (g83) & (g2938)) + ((!g78) & (!g79) & (!g135) & (g82) & (!g83) & (g2938)) + ((!g78) & (!g79) & (!g135) & (g82) & (g83) & (g2938)) + ((!g78) & (!g79) & (g135) & (!g82) & (!g83) & (g2938)) + ((!g78) & (!g79) & (g135) & (g82) & (!g83) & (g2938)) + ((!g78) & (!g79) & (g135) & (g82) & (g83) & (g2938)) + ((!g78) & (g79) & (!g135) & (!g82) & (!g83) & (g2938)) + ((!g78) & (g79) & (!g135) & (!g82) & (g83) & (g2938)) + ((!g78) & (g79) & (!g135) & (g82) & (!g83) & (g2938)) + ((!g78) & (g79) & (!g135) & (g82) & (g83) & (g2938)) + ((!g78) & (g79) & (g135) & (g82) & (!g83) & (g2938)) + ((!g78) & (g79) & (g135) & (g82) & (g83) & (g2938)) + ((g78) & (!g79) & (!g135) & (!g82) & (!g83) & (g2938)) + ((g78) & (!g79) & (!g135) & (!g82) & (g83) & (g2938)) + ((g78) & (!g79) & (!g135) & (g82) & (!g83) & (g2938)) + ((g78) & (!g79) & (!g135) & (g82) & (g83) & (g2938)) + ((g78) & (!g79) & (g135) & (g82) & (!g83) & (g2938)) + ((g78) & (!g79) & (g135) & (g82) & (g83) & (g2938)) + ((g78) & (g79) & (!g135) & (!g82) & (!g83) & (g2938)) + ((g78) & (g79) & (!g135) & (!g82) & (g83) & (g2938)) + ((g78) & (g79) & (!g135) & (g82) & (!g83) & (g2938)) + ((g78) & (g79) & (!g135) & (g82) & (g83) & (g2938)) + ((g78) & (g79) & (g135) & (!g82) & (g83) & (g2938)) + ((g78) & (g79) & (g135) & (g82) & (!g83) & (g2938)) + ((g78) & (g79) & (g135) & (g82) & (g83) & (g2938)));
	assign g2940 = (((!g78) & (!g79) & (!g2930) & (!sk[115]) & (g2939)) + ((!g78) & (!g79) & (!g2930) & (sk[115]) & (g2939)) + ((!g78) & (!g79) & (g2930) & (!sk[115]) & (g2939)) + ((!g78) & (!g79) & (g2930) & (sk[115]) & (g2939)) + ((!g78) & (g79) & (!g2930) & (!sk[115]) & (!g2939)) + ((!g78) & (g79) & (!g2930) & (!sk[115]) & (g2939)) + ((!g78) & (g79) & (!g2930) & (sk[115]) & (g2939)) + ((!g78) & (g79) & (g2930) & (!sk[115]) & (!g2939)) + ((!g78) & (g79) & (g2930) & (!sk[115]) & (g2939)) + ((g78) & (!g79) & (!g2930) & (!sk[115]) & (!g2939)) + ((g78) & (!g79) & (!g2930) & (!sk[115]) & (g2939)) + ((g78) & (!g79) & (!g2930) & (sk[115]) & (g2939)) + ((g78) & (!g79) & (g2930) & (!sk[115]) & (!g2939)) + ((g78) & (!g79) & (g2930) & (!sk[115]) & (g2939)) + ((g78) & (!g79) & (g2930) & (sk[115]) & (g2939)) + ((g78) & (g79) & (!g2930) & (!sk[115]) & (!g2939)) + ((g78) & (g79) & (!g2930) & (!sk[115]) & (g2939)) + ((g78) & (g79) & (!g2930) & (sk[115]) & (g2939)) + ((g78) & (g79) & (g2930) & (!sk[115]) & (!g2939)) + ((g78) & (g79) & (g2930) & (!sk[115]) & (g2939)) + ((g78) & (g79) & (g2930) & (sk[115]) & (g2939)));
	assign g2941 = (((!g2928) & (!g2024) & (sk[116]) & (g2935)) + ((!g2928) & (g2024) & (!sk[116]) & (!g2935)) + ((!g2928) & (g2024) & (!sk[116]) & (g2935)) + ((g2928) & (!g2024) & (!sk[116]) & (!g2935)) + ((g2928) & (!g2024) & (!sk[116]) & (g2935)) + ((g2928) & (g2024) & (!sk[116]) & (!g2935)) + ((g2928) & (g2024) & (!sk[116]) & (g2935)));
	assign g2942 = (((!g79) & (!g80) & (!g81) & (g133) & (!sk[117]) & (!g2941)) + ((!g79) & (!g80) & (!g81) & (g133) & (!sk[117]) & (g2941)) + ((!g79) & (!g80) & (g81) & (!g133) & (!sk[117]) & (!g2941)) + ((!g79) & (!g80) & (g81) & (!g133) & (!sk[117]) & (g2941)) + ((!g79) & (!g80) & (g81) & (g133) & (!sk[117]) & (!g2941)) + ((!g79) & (!g80) & (g81) & (g133) & (!sk[117]) & (g2941)) + ((!g79) & (g80) & (!g81) & (g133) & (!sk[117]) & (!g2941)) + ((!g79) & (g80) & (!g81) & (g133) & (!sk[117]) & (g2941)) + ((!g79) & (g80) & (g81) & (!g133) & (!sk[117]) & (!g2941)) + ((!g79) & (g80) & (g81) & (!g133) & (!sk[117]) & (g2941)) + ((!g79) & (g80) & (g81) & (g133) & (!sk[117]) & (!g2941)) + ((!g79) & (g80) & (g81) & (g133) & (!sk[117]) & (g2941)) + ((g79) & (!g80) & (!g81) & (!g133) & (!sk[117]) & (!g2941)) + ((g79) & (!g80) & (!g81) & (!g133) & (!sk[117]) & (g2941)) + ((g79) & (!g80) & (!g81) & (g133) & (!sk[117]) & (!g2941)) + ((g79) & (!g80) & (!g81) & (g133) & (!sk[117]) & (g2941)) + ((g79) & (!g80) & (!g81) & (g133) & (sk[117]) & (g2941)) + ((g79) & (!g80) & (g81) & (!g133) & (!sk[117]) & (!g2941)) + ((g79) & (!g80) & (g81) & (!g133) & (!sk[117]) & (g2941)) + ((g79) & (!g80) & (g81) & (g133) & (!sk[117]) & (!g2941)) + ((g79) & (!g80) & (g81) & (g133) & (!sk[117]) & (g2941)) + ((g79) & (g80) & (!g81) & (!g133) & (!sk[117]) & (!g2941)) + ((g79) & (g80) & (!g81) & (!g133) & (!sk[117]) & (g2941)) + ((g79) & (g80) & (!g81) & (g133) & (!sk[117]) & (!g2941)) + ((g79) & (g80) & (!g81) & (g133) & (!sk[117]) & (g2941)) + ((g79) & (g80) & (g81) & (!g133) & (!sk[117]) & (!g2941)) + ((g79) & (g80) & (g81) & (!g133) & (!sk[117]) & (g2941)) + ((g79) & (g80) & (g81) & (g133) & (!sk[117]) & (!g2941)) + ((g79) & (g80) & (g81) & (g133) & (!sk[117]) & (g2941)));
	assign g2943 = (((!sk[118]) & (!g79) & (g80) & (!g81)) + ((!sk[118]) & (!g79) & (g80) & (g81)) + ((!sk[118]) & (g79) & (!g80) & (!g81)) + ((!sk[118]) & (g79) & (!g80) & (g81)) + ((!sk[118]) & (g79) & (g80) & (!g81)) + ((!sk[118]) & (g79) & (g80) & (g81)) + ((sk[118]) & (g79) & (g80) & (!g81)));
	assign g2944 = (((!sk[119]) & (!g2363) & (g2938)) + ((!sk[119]) & (g2363) & (g2938)) + ((sk[119]) & (!g2363) & (g2938)));
	assign g2945 = (((g84) & (!g87) & (g89) & (g90) & (g2932) & (g2933)) + ((g84) & (g87) & (!g89) & (!g90) & (g2932) & (g2933)));
	assign g2946 = (((!sk[121]) & (!g2363) & (g2938) & (!g2945)) + ((!sk[121]) & (!g2363) & (g2938) & (g2945)) + ((!sk[121]) & (g2363) & (!g2938) & (!g2945)) + ((!sk[121]) & (g2363) & (!g2938) & (g2945)) + ((!sk[121]) & (g2363) & (g2938) & (!g2945)) + ((!sk[121]) & (g2363) & (g2938) & (g2945)) + ((sk[121]) & (!g2363) & (!g2938) & (!g2945)) + ((sk[121]) & (!g2363) & (g2938) & (!g2945)) + ((sk[121]) & (g2363) & (!g2938) & (!g2945)));
	assign g2947 = (((!g78) & (!g2943) & (!g82) & (!g83) & (!g2944) & (g2946)) + ((!g78) & (!g2943) & (!g82) & (!g83) & (g2944) & (g2946)) + ((!g78) & (!g2943) & (!g82) & (g83) & (!g2944) & (g2946)) + ((!g78) & (!g2943) & (!g82) & (g83) & (g2944) & (g2946)) + ((!g78) & (!g2943) & (g82) & (!g83) & (!g2944) & (g2946)) + ((!g78) & (!g2943) & (g82) & (!g83) & (g2944) & (g2946)) + ((!g78) & (!g2943) & (g82) & (g83) & (!g2944) & (g2946)) + ((!g78) & (!g2943) & (g82) & (g83) & (g2944) & (g2946)) + ((!g78) & (g2943) & (!g82) & (!g83) & (!g2944) & (g2946)) + ((!g78) & (g2943) & (!g82) & (g83) & (!g2944) & (g2946)) + ((!g78) & (g2943) & (g82) & (!g83) & (!g2944) & (g2946)) + ((!g78) & (g2943) & (g82) & (!g83) & (g2944) & (g2946)) + ((!g78) & (g2943) & (g82) & (g83) & (!g2944) & (g2946)) + ((!g78) & (g2943) & (g82) & (g83) & (g2944) & (g2946)) + ((g78) & (!g2943) & (!g82) & (!g83) & (!g2944) & (g2946)) + ((g78) & (!g2943) & (!g82) & (!g83) & (g2944) & (g2946)) + ((g78) & (!g2943) & (!g82) & (g83) & (!g2944) & (g2946)) + ((g78) & (!g2943) & (!g82) & (g83) & (g2944) & (g2946)) + ((g78) & (!g2943) & (g82) & (!g83) & (!g2944) & (g2946)) + ((g78) & (!g2943) & (g82) & (!g83) & (g2944) & (g2946)) + ((g78) & (!g2943) & (g82) & (g83) & (!g2944) & (g2946)) + ((g78) & (!g2943) & (g82) & (g83) & (g2944) & (g2946)) + ((g78) & (g2943) & (!g82) & (!g83) & (!g2944) & (g2946)) + ((g78) & (g2943) & (!g82) & (g83) & (!g2944) & (g2946)) + ((g78) & (g2943) & (!g82) & (g83) & (g2944) & (g2946)) + ((g78) & (g2943) & (g82) & (!g83) & (!g2944) & (g2946)) + ((g78) & (g2943) & (g82) & (!g83) & (g2944) & (g2946)) + ((g78) & (g2943) & (g82) & (g83) & (!g2944) & (g2946)) + ((g78) & (g2943) & (g82) & (g83) & (g2944) & (g2946)));
	assign g2948 = (((!g79) & (!g135) & (!g82) & (!g83) & (!g2938) & (g2947)) + ((!g79) & (!g135) & (!g82) & (!g83) & (g2938) & (g2947)) + ((!g79) & (!g135) & (!g82) & (g83) & (!g2938) & (g2947)) + ((!g79) & (!g135) & (!g82) & (g83) & (g2938) & (g2947)) + ((!g79) & (!g135) & (g82) & (!g83) & (!g2938) & (g2947)) + ((!g79) & (!g135) & (g82) & (!g83) & (g2938) & (g2947)) + ((!g79) & (!g135) & (g82) & (g83) & (!g2938) & (g2947)) + ((!g79) & (!g135) & (g82) & (g83) & (g2938) & (g2947)) + ((!g79) & (g135) & (!g82) & (!g83) & (!g2938) & (g2947)) + ((!g79) & (g135) & (!g82) & (!g83) & (g2938) & (g2947)) + ((!g79) & (g135) & (!g82) & (g83) & (!g2938) & (g2947)) + ((!g79) & (g135) & (g82) & (!g83) & (!g2938) & (g2947)) + ((!g79) & (g135) & (g82) & (!g83) & (g2938) & (g2947)) + ((!g79) & (g135) & (g82) & (g83) & (!g2938) & (g2947)) + ((!g79) & (g135) & (g82) & (g83) & (g2938) & (g2947)) + ((g79) & (!g135) & (!g82) & (!g83) & (!g2938) & (g2947)) + ((g79) & (!g135) & (!g82) & (!g83) & (g2938) & (g2947)) + ((g79) & (!g135) & (!g82) & (g83) & (!g2938) & (g2947)) + ((g79) & (!g135) & (!g82) & (g83) & (g2938) & (g2947)) + ((g79) & (!g135) & (g82) & (!g83) & (!g2938) & (g2947)) + ((g79) & (!g135) & (g82) & (!g83) & (g2938) & (g2947)) + ((g79) & (!g135) & (g82) & (g83) & (!g2938) & (g2947)) + ((g79) & (!g135) & (g82) & (g83) & (g2938) & (g2947)) + ((g79) & (g135) & (!g82) & (!g83) & (!g2938) & (g2947)) + ((g79) & (g135) & (!g82) & (!g83) & (g2938) & (g2947)) + ((g79) & (g135) & (!g82) & (g83) & (!g2938) & (g2947)) + ((g79) & (g135) & (!g82) & (g83) & (g2938) & (g2947)) + ((g79) & (g135) & (g82) & (!g83) & (!g2938) & (g2947)) + ((g79) & (g135) & (g82) & (!g83) & (g2938) & (g2947)) + ((g79) & (g135) & (g82) & (g83) & (!g2938) & (g2947)) + ((g79) & (g135) & (g82) & (g83) & (g2938) & (g2947)));
	assign g2949 = (((!g2942) & (!sk[124]) & (g2948)) + ((!g2942) & (sk[124]) & (g2948)) + ((g2942) & (!sk[124]) & (g2948)));
	assign g2950 = (((!sk[125]) & (!g2940) & (g2949)) + ((!sk[125]) & (g2940) & (g2949)) + ((sk[125]) & (!g2940) & (g2949)));
	assign g2951 = (((!g2928) & (!sk[126]) & (g2920)) + ((g2928) & (!sk[126]) & (g2920)) + ((g2928) & (sk[126]) & (!g2920)));
	assign g2952 = (((!g2928) & (!g2024) & (!g2950) & (!sk[127]) & (g2951)) + ((!g2928) & (!g2024) & (g2950) & (!sk[127]) & (g2951)) + ((!g2928) & (!g2024) & (g2950) & (sk[127]) & (!g2951)) + ((!g2928) & (g2024) & (!g2950) & (!sk[127]) & (!g2951)) + ((!g2928) & (g2024) & (!g2950) & (!sk[127]) & (g2951)) + ((!g2928) & (g2024) & (!g2950) & (sk[127]) & (!g2951)) + ((!g2928) & (g2024) & (g2950) & (!sk[127]) & (!g2951)) + ((!g2928) & (g2024) & (g2950) & (!sk[127]) & (g2951)) + ((!g2928) & (g2024) & (g2950) & (sk[127]) & (!g2951)) + ((g2928) & (!g2024) & (!g2950) & (!sk[127]) & (!g2951)) + ((g2928) & (!g2024) & (!g2950) & (!sk[127]) & (g2951)) + ((g2928) & (!g2024) & (!g2950) & (sk[127]) & (!g2951)) + ((g2928) & (!g2024) & (g2950) & (!sk[127]) & (!g2951)) + ((g2928) & (!g2024) & (g2950) & (!sk[127]) & (g2951)) + ((g2928) & (!g2024) & (g2950) & (sk[127]) & (!g2951)) + ((g2928) & (g2024) & (!g2950) & (!sk[127]) & (!g2951)) + ((g2928) & (g2024) & (!g2950) & (!sk[127]) & (g2951)) + ((g2928) & (g2024) & (!g2950) & (sk[127]) & (!g2951)) + ((g2928) & (g2024) & (g2950) & (!sk[127]) & (!g2951)) + ((g2928) & (g2024) & (g2950) & (!sk[127]) & (g2951)) + ((g2928) & (g2024) & (g2950) & (sk[127]) & (!g2951)));
	assign g2953 = (((!g2928) & (!sk[0]) & (!g2060) & (!g2929) & (g2952)) + ((!g2928) & (!sk[0]) & (!g2060) & (g2929) & (g2952)) + ((!g2928) & (!sk[0]) & (g2060) & (!g2929) & (!g2952)) + ((!g2928) & (!sk[0]) & (g2060) & (!g2929) & (g2952)) + ((!g2928) & (!sk[0]) & (g2060) & (g2929) & (!g2952)) + ((!g2928) & (!sk[0]) & (g2060) & (g2929) & (g2952)) + ((!g2928) & (sk[0]) & (!g2060) & (g2929) & (g2952)) + ((!g2928) & (sk[0]) & (g2060) & (g2929) & (g2952)) + ((g2928) & (!sk[0]) & (!g2060) & (!g2929) & (!g2952)) + ((g2928) & (!sk[0]) & (!g2060) & (!g2929) & (g2952)) + ((g2928) & (!sk[0]) & (!g2060) & (g2929) & (!g2952)) + ((g2928) & (!sk[0]) & (!g2060) & (g2929) & (g2952)) + ((g2928) & (!sk[0]) & (g2060) & (!g2929) & (!g2952)) + ((g2928) & (!sk[0]) & (g2060) & (!g2929) & (g2952)) + ((g2928) & (!sk[0]) & (g2060) & (g2929) & (!g2952)) + ((g2928) & (!sk[0]) & (g2060) & (g2929) & (g2952)) + ((g2928) & (sk[0]) & (g2060) & (!g2929) & (g2952)) + ((g2928) & (sk[0]) & (g2060) & (g2929) & (g2952)));
	assign g2954 = (((!g2928) & (!g2024) & (sk[1]) & (g2950)) + ((!g2928) & (g2024) & (!sk[1]) & (!g2950)) + ((!g2928) & (g2024) & (!sk[1]) & (g2950)) + ((g2928) & (!g2024) & (!sk[1]) & (!g2950)) + ((g2928) & (!g2024) & (!sk[1]) & (g2950)) + ((g2928) & (g2024) & (!sk[1]) & (!g2950)) + ((g2928) & (g2024) & (!sk[1]) & (g2950)));
	assign g2955 = (((!g78) & (!sk[2]) & (!g79) & (!g2930) & (g2937)) + ((!g78) & (!sk[2]) & (!g79) & (g2930) & (g2937)) + ((!g78) & (!sk[2]) & (g79) & (!g2930) & (!g2937)) + ((!g78) & (!sk[2]) & (g79) & (!g2930) & (g2937)) + ((!g78) & (!sk[2]) & (g79) & (g2930) & (!g2937)) + ((!g78) & (!sk[2]) & (g79) & (g2930) & (g2937)) + ((g78) & (!sk[2]) & (!g79) & (!g2930) & (!g2937)) + ((g78) & (!sk[2]) & (!g79) & (!g2930) & (g2937)) + ((g78) & (!sk[2]) & (!g79) & (g2930) & (!g2937)) + ((g78) & (!sk[2]) & (!g79) & (g2930) & (g2937)) + ((g78) & (!sk[2]) & (g79) & (!g2930) & (!g2937)) + ((g78) & (!sk[2]) & (g79) & (!g2930) & (g2937)) + ((g78) & (!sk[2]) & (g79) & (g2930) & (!g2937)) + ((g78) & (!sk[2]) & (g79) & (g2930) & (g2937)) + ((g78) & (sk[2]) & (g79) & (g2930) & (g2937)));
	assign g2956 = (((!g118) & (!g85) & (!sk[3]) & (!g86) & (g2936)) + ((!g118) & (!g85) & (!sk[3]) & (g86) & (g2936)) + ((!g118) & (g85) & (!sk[3]) & (!g86) & (!g2936)) + ((!g118) & (g85) & (!sk[3]) & (!g86) & (g2936)) + ((!g118) & (g85) & (!sk[3]) & (g86) & (!g2936)) + ((!g118) & (g85) & (!sk[3]) & (g86) & (g2936)) + ((g118) & (!g85) & (!sk[3]) & (!g86) & (!g2936)) + ((g118) & (!g85) & (!sk[3]) & (!g86) & (g2936)) + ((g118) & (!g85) & (!sk[3]) & (g86) & (!g2936)) + ((g118) & (!g85) & (!sk[3]) & (g86) & (g2936)) + ((g118) & (!g85) & (sk[3]) & (g86) & (g2936)) + ((g118) & (g85) & (!sk[3]) & (!g86) & (!g2936)) + ((g118) & (g85) & (!sk[3]) & (!g86) & (g2936)) + ((g118) & (g85) & (!sk[3]) & (g86) & (!g2936)) + ((g118) & (g85) & (!sk[3]) & (g86) & (g2936)));
	assign g2957 = (((!g119) & (!sk[4]) & (g2935)) + ((!g119) & (sk[4]) & (g2935)) + ((g119) & (!sk[4]) & (g2935)));
	assign g2958 = (((!g78) & (!g79) & (!g2930) & (!sk[5]) & (g2939)) + ((!g78) & (!g79) & (g2930) & (!sk[5]) & (g2939)) + ((!g78) & (g79) & (!g2930) & (!sk[5]) & (!g2939)) + ((!g78) & (g79) & (!g2930) & (!sk[5]) & (g2939)) + ((!g78) & (g79) & (g2930) & (!sk[5]) & (!g2939)) + ((!g78) & (g79) & (g2930) & (!sk[5]) & (g2939)) + ((!g78) & (g79) & (g2930) & (sk[5]) & (g2939)) + ((g78) & (!g79) & (!g2930) & (!sk[5]) & (!g2939)) + ((g78) & (!g79) & (!g2930) & (!sk[5]) & (g2939)) + ((g78) & (!g79) & (g2930) & (!sk[5]) & (!g2939)) + ((g78) & (!g79) & (g2930) & (!sk[5]) & (g2939)) + ((g78) & (g79) & (!g2930) & (!sk[5]) & (!g2939)) + ((g78) & (g79) & (!g2930) & (!sk[5]) & (g2939)) + ((g78) & (g79) & (g2930) & (!sk[5]) & (!g2939)) + ((g78) & (g79) & (g2930) & (!sk[5]) & (g2939)));
	assign g2959 = (((!sk[6]) & (!g118) & (!g86) & (!g2957) & (g2958)) + ((!sk[6]) & (!g118) & (!g86) & (g2957) & (g2958)) + ((!sk[6]) & (!g118) & (g86) & (!g2957) & (!g2958)) + ((!sk[6]) & (!g118) & (g86) & (!g2957) & (g2958)) + ((!sk[6]) & (!g118) & (g86) & (g2957) & (!g2958)) + ((!sk[6]) & (!g118) & (g86) & (g2957) & (g2958)) + ((!sk[6]) & (g118) & (!g86) & (!g2957) & (!g2958)) + ((!sk[6]) & (g118) & (!g86) & (!g2957) & (g2958)) + ((!sk[6]) & (g118) & (!g86) & (g2957) & (!g2958)) + ((!sk[6]) & (g118) & (!g86) & (g2957) & (g2958)) + ((!sk[6]) & (g118) & (g86) & (!g2957) & (!g2958)) + ((!sk[6]) & (g118) & (g86) & (!g2957) & (g2958)) + ((!sk[6]) & (g118) & (g86) & (g2957) & (!g2958)) + ((!sk[6]) & (g118) & (g86) & (g2957) & (g2958)) + ((sk[6]) & (!g118) & (!g86) & (!g2957) & (!g2958)) + ((sk[6]) & (!g118) & (!g86) & (g2957) & (!g2958)) + ((sk[6]) & (!g118) & (g86) & (!g2957) & (!g2958)) + ((sk[6]) & (!g118) & (g86) & (g2957) & (!g2958)) + ((sk[6]) & (g118) & (!g86) & (!g2957) & (!g2958)) + ((sk[6]) & (g118) & (g86) & (!g2957) & (!g2958)) + ((sk[6]) & (g118) & (g86) & (g2957) & (!g2958)));
	assign g2960 = (((!g78) & (g79) & (g80) & (!g81) & (g82) & (!g83)));
	assign g2961 = (((!g2941) & (!sk[8]) & (g2960)) + ((g2941) & (!sk[8]) & (g2960)) + ((g2941) & (sk[8]) & (g2960)));
	assign g2962 = (((!g2931) & (!sk[9]) & (!g2956) & (!g2959) & (g2961)) + ((!g2931) & (!sk[9]) & (!g2956) & (g2959) & (g2961)) + ((!g2931) & (!sk[9]) & (g2956) & (!g2959) & (!g2961)) + ((!g2931) & (!sk[9]) & (g2956) & (!g2959) & (g2961)) + ((!g2931) & (!sk[9]) & (g2956) & (g2959) & (!g2961)) + ((!g2931) & (!sk[9]) & (g2956) & (g2959) & (g2961)) + ((!g2931) & (sk[9]) & (!g2956) & (g2959) & (!g2961)) + ((g2931) & (!sk[9]) & (!g2956) & (!g2959) & (!g2961)) + ((g2931) & (!sk[9]) & (!g2956) & (!g2959) & (g2961)) + ((g2931) & (!sk[9]) & (!g2956) & (g2959) & (!g2961)) + ((g2931) & (!sk[9]) & (!g2956) & (g2959) & (g2961)) + ((g2931) & (!sk[9]) & (g2956) & (!g2959) & (!g2961)) + ((g2931) & (!sk[9]) & (g2956) & (!g2959) & (g2961)) + ((g2931) & (!sk[9]) & (g2956) & (g2959) & (!g2961)) + ((g2931) & (!sk[9]) & (g2956) & (g2959) & (g2961)));
	assign g2963 = (((!g99) & (!g2955) & (sk[10]) & (g2962)) + ((!g99) & (g2955) & (!sk[10]) & (!g2962)) + ((!g99) & (g2955) & (!sk[10]) & (g2962)) + ((g99) & (!g2955) & (!sk[10]) & (!g2962)) + ((g99) & (!g2955) & (!sk[10]) & (g2962)) + ((g99) & (g2955) & (!sk[10]) & (!g2962)) + ((g99) & (g2955) & (!sk[10]) & (g2962)));
	assign g2964 = (((!g89) & (!sk[11]) & (!g1604) & (!g2954) & (g2963)) + ((!g89) & (!sk[11]) & (!g1604) & (g2954) & (g2963)) + ((!g89) & (!sk[11]) & (g1604) & (!g2954) & (!g2963)) + ((!g89) & (!sk[11]) & (g1604) & (!g2954) & (g2963)) + ((!g89) & (!sk[11]) & (g1604) & (g2954) & (!g2963)) + ((!g89) & (!sk[11]) & (g1604) & (g2954) & (g2963)) + ((!g89) & (sk[11]) & (g1604) & (g2954) & (g2963)) + ((g89) & (!sk[11]) & (!g1604) & (!g2954) & (!g2963)) + ((g89) & (!sk[11]) & (!g1604) & (!g2954) & (g2963)) + ((g89) & (!sk[11]) & (!g1604) & (g2954) & (!g2963)) + ((g89) & (!sk[11]) & (!g1604) & (g2954) & (g2963)) + ((g89) & (!sk[11]) & (g1604) & (!g2954) & (!g2963)) + ((g89) & (!sk[11]) & (g1604) & (!g2954) & (g2963)) + ((g89) & (!sk[11]) & (g1604) & (g2954) & (!g2963)) + ((g89) & (!sk[11]) & (g1604) & (g2954) & (g2963)) + ((g89) & (sk[11]) & (!g1604) & (g2954) & (!g2963)) + ((g89) & (sk[11]) & (g1604) & (g2954) & (!g2963)) + ((g89) & (sk[11]) & (g1604) & (g2954) & (g2963)));
	assign g2965 = (((!g1656) & (!g318) & (!sk[12]) & (!g2954) & (g2963)) + ((!g1656) & (!g318) & (!sk[12]) & (g2954) & (g2963)) + ((!g1656) & (g318) & (!sk[12]) & (!g2954) & (!g2963)) + ((!g1656) & (g318) & (!sk[12]) & (!g2954) & (g2963)) + ((!g1656) & (g318) & (!sk[12]) & (g2954) & (!g2963)) + ((!g1656) & (g318) & (!sk[12]) & (g2954) & (g2963)) + ((!g1656) & (g318) & (sk[12]) & (g2954) & (!g2963)) + ((g1656) & (!g318) & (!sk[12]) & (!g2954) & (!g2963)) + ((g1656) & (!g318) & (!sk[12]) & (!g2954) & (g2963)) + ((g1656) & (!g318) & (!sk[12]) & (g2954) & (!g2963)) + ((g1656) & (!g318) & (!sk[12]) & (g2954) & (g2963)) + ((g1656) & (!g318) & (sk[12]) & (g2954) & (g2963)) + ((g1656) & (g318) & (!sk[12]) & (!g2954) & (!g2963)) + ((g1656) & (g318) & (!sk[12]) & (!g2954) & (g2963)) + ((g1656) & (g318) & (!sk[12]) & (g2954) & (!g2963)) + ((g1656) & (g318) & (!sk[12]) & (g2954) & (g2963)) + ((g1656) & (g318) & (sk[12]) & (g2954) & (!g2963)) + ((g1656) & (g318) & (sk[12]) & (g2954) & (g2963)));
	assign g2966 = (((!g88) & (!sk[13]) & (!g1620) & (!g2954) & (g2963)) + ((!g88) & (!sk[13]) & (!g1620) & (g2954) & (g2963)) + ((!g88) & (!sk[13]) & (g1620) & (!g2954) & (!g2963)) + ((!g88) & (!sk[13]) & (g1620) & (!g2954) & (g2963)) + ((!g88) & (!sk[13]) & (g1620) & (g2954) & (!g2963)) + ((!g88) & (!sk[13]) & (g1620) & (g2954) & (g2963)) + ((!g88) & (sk[13]) & (g1620) & (g2954) & (g2963)) + ((g88) & (!sk[13]) & (!g1620) & (!g2954) & (!g2963)) + ((g88) & (!sk[13]) & (!g1620) & (!g2954) & (g2963)) + ((g88) & (!sk[13]) & (!g1620) & (g2954) & (!g2963)) + ((g88) & (!sk[13]) & (!g1620) & (g2954) & (g2963)) + ((g88) & (!sk[13]) & (g1620) & (!g2954) & (!g2963)) + ((g88) & (!sk[13]) & (g1620) & (!g2954) & (g2963)) + ((g88) & (!sk[13]) & (g1620) & (g2954) & (!g2963)) + ((g88) & (!sk[13]) & (g1620) & (g2954) & (g2963)) + ((g88) & (sk[13]) & (!g1620) & (g2954) & (!g2963)) + ((g88) & (sk[13]) & (g1620) & (g2954) & (!g2963)) + ((g88) & (sk[13]) & (g1620) & (g2954) & (g2963)));
	assign g2967 = (((!g90) & (!sk[14]) & (!g1644) & (!g2954) & (g2963)) + ((!g90) & (!sk[14]) & (!g1644) & (g2954) & (g2963)) + ((!g90) & (!sk[14]) & (g1644) & (!g2954) & (!g2963)) + ((!g90) & (!sk[14]) & (g1644) & (!g2954) & (g2963)) + ((!g90) & (!sk[14]) & (g1644) & (g2954) & (!g2963)) + ((!g90) & (!sk[14]) & (g1644) & (g2954) & (g2963)) + ((!g90) & (sk[14]) & (g1644) & (g2954) & (g2963)) + ((g90) & (!sk[14]) & (!g1644) & (!g2954) & (!g2963)) + ((g90) & (!sk[14]) & (!g1644) & (!g2954) & (g2963)) + ((g90) & (!sk[14]) & (!g1644) & (g2954) & (!g2963)) + ((g90) & (!sk[14]) & (!g1644) & (g2954) & (g2963)) + ((g90) & (!sk[14]) & (g1644) & (!g2954) & (!g2963)) + ((g90) & (!sk[14]) & (g1644) & (!g2954) & (g2963)) + ((g90) & (!sk[14]) & (g1644) & (g2954) & (!g2963)) + ((g90) & (!sk[14]) & (g1644) & (g2954) & (g2963)) + ((g90) & (sk[14]) & (!g1644) & (g2954) & (!g2963)) + ((g90) & (sk[14]) & (g1644) & (g2954) & (!g2963)) + ((g90) & (sk[14]) & (g1644) & (g2954) & (g2963)));
	assign g2968 = (((!g87) & (!g1632) & (!g2954) & (!sk[15]) & (g2963)) + ((!g87) & (!g1632) & (g2954) & (!sk[15]) & (g2963)) + ((!g87) & (g1632) & (!g2954) & (!sk[15]) & (!g2963)) + ((!g87) & (g1632) & (!g2954) & (!sk[15]) & (g2963)) + ((!g87) & (g1632) & (g2954) & (!sk[15]) & (!g2963)) + ((!g87) & (g1632) & (g2954) & (!sk[15]) & (g2963)) + ((!g87) & (g1632) & (g2954) & (sk[15]) & (g2963)) + ((g87) & (!g1632) & (!g2954) & (!sk[15]) & (!g2963)) + ((g87) & (!g1632) & (!g2954) & (!sk[15]) & (g2963)) + ((g87) & (!g1632) & (g2954) & (!sk[15]) & (!g2963)) + ((g87) & (!g1632) & (g2954) & (!sk[15]) & (g2963)) + ((g87) & (!g1632) & (g2954) & (sk[15]) & (!g2963)) + ((g87) & (g1632) & (!g2954) & (!sk[15]) & (!g2963)) + ((g87) & (g1632) & (!g2954) & (!sk[15]) & (g2963)) + ((g87) & (g1632) & (g2954) & (!sk[15]) & (!g2963)) + ((g87) & (g1632) & (g2954) & (!sk[15]) & (g2963)) + ((g87) & (g1632) & (g2954) & (sk[15]) & (!g2963)) + ((g87) & (g1632) & (g2954) & (sk[15]) & (g2963)));
	assign g5057 = (((!sk[16]) & (!g2924) & (g3115) & (!g2969)) + ((!sk[16]) & (!g2924) & (g3115) & (g2969)) + ((!sk[16]) & (g2924) & (!g3115) & (!g2969)) + ((!sk[16]) & (g2924) & (!g3115) & (g2969)) + ((!sk[16]) & (g2924) & (g3115) & (!g2969)) + ((!sk[16]) & (g2924) & (g3115) & (g2969)) + ((sk[16]) & (!g2924) & (!g3115) & (g2969)) + ((sk[16]) & (!g2924) & (g3115) & (g2969)) + ((sk[16]) & (g2924) & (g3115) & (!g2969)) + ((sk[16]) & (g2924) & (g3115) & (g2969)));
	assign g2970 = (((!g2795) & (!g2796) & (!sk[17]) & (!g2813) & (g3120) & (!g3121)) + ((!g2795) & (!g2796) & (!sk[17]) & (!g2813) & (g3120) & (g3121)) + ((!g2795) & (!g2796) & (!sk[17]) & (g2813) & (!g3120) & (!g3121)) + ((!g2795) & (!g2796) & (!sk[17]) & (g2813) & (!g3120) & (g3121)) + ((!g2795) & (!g2796) & (!sk[17]) & (g2813) & (g3120) & (!g3121)) + ((!g2795) & (!g2796) & (!sk[17]) & (g2813) & (g3120) & (g3121)) + ((!g2795) & (!g2796) & (sk[17]) & (!g2813) & (!g3120) & (g3121)) + ((!g2795) & (!g2796) & (sk[17]) & (!g2813) & (g3120) & (g3121)) + ((!g2795) & (!g2796) & (sk[17]) & (g2813) & (!g3120) & (g3121)) + ((!g2795) & (!g2796) & (sk[17]) & (g2813) & (g3120) & (g3121)) + ((!g2795) & (g2796) & (!sk[17]) & (!g2813) & (g3120) & (!g3121)) + ((!g2795) & (g2796) & (!sk[17]) & (!g2813) & (g3120) & (g3121)) + ((!g2795) & (g2796) & (!sk[17]) & (g2813) & (!g3120) & (!g3121)) + ((!g2795) & (g2796) & (!sk[17]) & (g2813) & (!g3120) & (g3121)) + ((!g2795) & (g2796) & (!sk[17]) & (g2813) & (g3120) & (!g3121)) + ((!g2795) & (g2796) & (!sk[17]) & (g2813) & (g3120) & (g3121)) + ((!g2795) & (g2796) & (sk[17]) & (!g2813) & (!g3120) & (g3121)) + ((!g2795) & (g2796) & (sk[17]) & (!g2813) & (g3120) & (g3121)) + ((!g2795) & (g2796) & (sk[17]) & (g2813) & (!g3120) & (g3121)) + ((!g2795) & (g2796) & (sk[17]) & (g2813) & (g3120) & (g3121)) + ((g2795) & (!g2796) & (!sk[17]) & (!g2813) & (!g3120) & (!g3121)) + ((g2795) & (!g2796) & (!sk[17]) & (!g2813) & (!g3120) & (g3121)) + ((g2795) & (!g2796) & (!sk[17]) & (!g2813) & (g3120) & (!g3121)) + ((g2795) & (!g2796) & (!sk[17]) & (!g2813) & (g3120) & (g3121)) + ((g2795) & (!g2796) & (!sk[17]) & (g2813) & (!g3120) & (!g3121)) + ((g2795) & (!g2796) & (!sk[17]) & (g2813) & (!g3120) & (g3121)) + ((g2795) & (!g2796) & (!sk[17]) & (g2813) & (g3120) & (!g3121)) + ((g2795) & (!g2796) & (!sk[17]) & (g2813) & (g3120) & (g3121)) + ((g2795) & (!g2796) & (sk[17]) & (!g2813) & (!g3120) & (g3121)) + ((g2795) & (!g2796) & (sk[17]) & (!g2813) & (g3120) & (g3121)) + ((g2795) & (!g2796) & (sk[17]) & (g2813) & (!g3120) & (g3121)) + ((g2795) & (!g2796) & (sk[17]) & (g2813) & (g3120) & (g3121)) + ((g2795) & (g2796) & (!sk[17]) & (!g2813) & (!g3120) & (!g3121)) + ((g2795) & (g2796) & (!sk[17]) & (!g2813) & (!g3120) & (g3121)) + ((g2795) & (g2796) & (!sk[17]) & (!g2813) & (g3120) & (!g3121)) + ((g2795) & (g2796) & (!sk[17]) & (!g2813) & (g3120) & (g3121)) + ((g2795) & (g2796) & (!sk[17]) & (g2813) & (!g3120) & (!g3121)) + ((g2795) & (g2796) & (!sk[17]) & (g2813) & (!g3120) & (g3121)) + ((g2795) & (g2796) & (!sk[17]) & (g2813) & (g3120) & (!g3121)) + ((g2795) & (g2796) & (!sk[17]) & (g2813) & (g3120) & (g3121)) + ((g2795) & (g2796) & (sk[17]) & (!g2813) & (!g3120) & (g3121)) + ((g2795) & (g2796) & (sk[17]) & (!g2813) & (g3120) & (g3121)) + ((g2795) & (g2796) & (sk[17]) & (g2813) & (!g3120) & (!g3121)) + ((g2795) & (g2796) & (sk[17]) & (g2813) & (!g3120) & (g3121)));
	assign g2971 = (((!g2080) & (!g2079) & (!sk[18]) & (!g2124) & (g2125) & (!g2970)) + ((!g2080) & (!g2079) & (!sk[18]) & (!g2124) & (g2125) & (g2970)) + ((!g2080) & (!g2079) & (!sk[18]) & (g2124) & (!g2125) & (!g2970)) + ((!g2080) & (!g2079) & (!sk[18]) & (g2124) & (!g2125) & (g2970)) + ((!g2080) & (!g2079) & (!sk[18]) & (g2124) & (g2125) & (!g2970)) + ((!g2080) & (!g2079) & (!sk[18]) & (g2124) & (g2125) & (g2970)) + ((!g2080) & (g2079) & (!sk[18]) & (!g2124) & (g2125) & (!g2970)) + ((!g2080) & (g2079) & (!sk[18]) & (!g2124) & (g2125) & (g2970)) + ((!g2080) & (g2079) & (!sk[18]) & (g2124) & (!g2125) & (!g2970)) + ((!g2080) & (g2079) & (!sk[18]) & (g2124) & (!g2125) & (g2970)) + ((!g2080) & (g2079) & (!sk[18]) & (g2124) & (g2125) & (!g2970)) + ((!g2080) & (g2079) & (!sk[18]) & (g2124) & (g2125) & (g2970)) + ((!g2080) & (g2079) & (sk[18]) & (!g2124) & (!g2125) & (!g2970)) + ((!g2080) & (g2079) & (sk[18]) & (!g2124) & (!g2125) & (g2970)) + ((!g2080) & (g2079) & (sk[18]) & (!g2124) & (g2125) & (!g2970)) + ((!g2080) & (g2079) & (sk[18]) & (!g2124) & (g2125) & (g2970)) + ((!g2080) & (g2079) & (sk[18]) & (g2124) & (!g2125) & (!g2970)) + ((!g2080) & (g2079) & (sk[18]) & (g2124) & (!g2125) & (g2970)) + ((!g2080) & (g2079) & (sk[18]) & (g2124) & (g2125) & (!g2970)) + ((!g2080) & (g2079) & (sk[18]) & (g2124) & (g2125) & (g2970)) + ((g2080) & (!g2079) & (!sk[18]) & (!g2124) & (!g2125) & (!g2970)) + ((g2080) & (!g2079) & (!sk[18]) & (!g2124) & (!g2125) & (g2970)) + ((g2080) & (!g2079) & (!sk[18]) & (!g2124) & (g2125) & (!g2970)) + ((g2080) & (!g2079) & (!sk[18]) & (!g2124) & (g2125) & (g2970)) + ((g2080) & (!g2079) & (!sk[18]) & (g2124) & (!g2125) & (!g2970)) + ((g2080) & (!g2079) & (!sk[18]) & (g2124) & (!g2125) & (g2970)) + ((g2080) & (!g2079) & (!sk[18]) & (g2124) & (g2125) & (!g2970)) + ((g2080) & (!g2079) & (!sk[18]) & (g2124) & (g2125) & (g2970)) + ((g2080) & (!g2079) & (sk[18]) & (!g2124) & (!g2125) & (g2970)) + ((g2080) & (g2079) & (!sk[18]) & (!g2124) & (!g2125) & (!g2970)) + ((g2080) & (g2079) & (!sk[18]) & (!g2124) & (!g2125) & (g2970)) + ((g2080) & (g2079) & (!sk[18]) & (!g2124) & (g2125) & (!g2970)) + ((g2080) & (g2079) & (!sk[18]) & (!g2124) & (g2125) & (g2970)) + ((g2080) & (g2079) & (!sk[18]) & (g2124) & (!g2125) & (!g2970)) + ((g2080) & (g2079) & (!sk[18]) & (g2124) & (!g2125) & (g2970)) + ((g2080) & (g2079) & (!sk[18]) & (g2124) & (g2125) & (!g2970)) + ((g2080) & (g2079) & (!sk[18]) & (g2124) & (g2125) & (g2970)) + ((g2080) & (g2079) & (sk[18]) & (!g2124) & (!g2125) & (g2970)) + ((g2080) & (g2079) & (sk[18]) & (!g2124) & (g2125) & (!g2970)) + ((g2080) & (g2079) & (sk[18]) & (!g2124) & (g2125) & (g2970)) + ((g2080) & (g2079) & (sk[18]) & (g2124) & (!g2125) & (!g2970)) + ((g2080) & (g2079) & (sk[18]) & (g2124) & (!g2125) & (g2970)) + ((g2080) & (g2079) & (sk[18]) & (g2124) & (g2125) & (!g2970)) + ((g2080) & (g2079) & (sk[18]) & (g2124) & (g2125) & (g2970)));
	assign g2972 = (((!g2030) & (!g2913) & (!g2969) & (!g2079) & (g2970) & (g3122)) + ((!g2030) & (!g2913) & (!g2969) & (g2079) & (!g2970) & (!g3122)) + ((!g2030) & (!g2913) & (!g2969) & (g2079) & (g2970) & (!g3122)) + ((!g2030) & (!g2913) & (!g2969) & (g2079) & (g2970) & (g3122)) + ((!g2030) & (!g2913) & (g2969) & (!g2079) & (g2970) & (g3122)) + ((!g2030) & (!g2913) & (g2969) & (g2079) & (!g2970) & (!g3122)) + ((!g2030) & (!g2913) & (g2969) & (g2079) & (g2970) & (!g3122)) + ((!g2030) & (!g2913) & (g2969) & (g2079) & (g2970) & (g3122)) + ((!g2030) & (g2913) & (!g2969) & (!g2079) & (!g2970) & (g3122)) + ((!g2030) & (g2913) & (!g2969) & (!g2079) & (g2970) & (g3122)) + ((!g2030) & (g2913) & (!g2969) & (g2079) & (!g2970) & (g3122)) + ((!g2030) & (g2913) & (!g2969) & (g2079) & (g2970) & (g3122)) + ((!g2030) & (g2913) & (g2969) & (!g2079) & (!g2970) & (g3122)) + ((!g2030) & (g2913) & (g2969) & (!g2079) & (g2970) & (g3122)) + ((!g2030) & (g2913) & (g2969) & (g2079) & (!g2970) & (g3122)) + ((!g2030) & (g2913) & (g2969) & (g2079) & (g2970) & (g3122)) + ((g2030) & (!g2913) & (g2969) & (!g2079) & (!g2970) & (!g3122)) + ((g2030) & (!g2913) & (g2969) & (!g2079) & (!g2970) & (g3122)) + ((g2030) & (!g2913) & (g2969) & (!g2079) & (g2970) & (!g3122)) + ((g2030) & (!g2913) & (g2969) & (!g2079) & (g2970) & (g3122)) + ((g2030) & (!g2913) & (g2969) & (g2079) & (!g2970) & (!g3122)) + ((g2030) & (!g2913) & (g2969) & (g2079) & (!g2970) & (g3122)) + ((g2030) & (!g2913) & (g2969) & (g2079) & (g2970) & (!g3122)) + ((g2030) & (!g2913) & (g2969) & (g2079) & (g2970) & (g3122)) + ((g2030) & (g2913) & (g2969) & (!g2079) & (!g2970) & (!g3122)) + ((g2030) & (g2913) & (g2969) & (!g2079) & (!g2970) & (g3122)) + ((g2030) & (g2913) & (g2969) & (!g2079) & (g2970) & (!g3122)) + ((g2030) & (g2913) & (g2969) & (!g2079) & (g2970) & (g3122)) + ((g2030) & (g2913) & (g2969) & (g2079) & (!g2970) & (!g3122)) + ((g2030) & (g2913) & (g2969) & (g2079) & (!g2970) & (g3122)) + ((g2030) & (g2913) & (g2969) & (g2079) & (g2970) & (!g3122)) + ((g2030) & (g2913) & (g2969) & (g2079) & (g2970) & (g3122)));
	assign g2973 = (((!nmi_i) & (!g2023) & (!intr_i) & (!g2330) & (g2843) & (g2972)) + ((!nmi_i) & (!g2023) & (!intr_i) & (g2330) & (g2843) & (g2972)) + ((!nmi_i) & (!g2023) & (intr_i) & (g2330) & (g2843) & (g2972)));
	assign g2974 = (((g84) & (!g87) & (!g88) & (!g89) & (g102) & (!g3139)) + ((g84) & (!g87) & (!g88) & (!g89) & (g102) & (g3139)) + ((g84) & (!g87) & (!g88) & (g89) & (g102) & (!g3139)) + ((g84) & (!g87) & (!g88) & (g89) & (g102) & (g3139)) + ((g84) & (!g87) & (g88) & (!g89) & (g102) & (g3139)) + ((g84) & (!g87) & (g88) & (g89) & (g102) & (!g3139)) + ((g84) & (!g87) & (g88) & (g89) & (g102) & (g3139)));
	assign g2975 = (((!sk[22]) & (!g2931) & (g99) & (!g2974)) + ((!sk[22]) & (!g2931) & (g99) & (g2974)) + ((!sk[22]) & (g2931) & (!g99) & (!g2974)) + ((!sk[22]) & (g2931) & (!g99) & (g2974)) + ((!sk[22]) & (g2931) & (g99) & (!g2974)) + ((!sk[22]) & (g2931) & (g99) & (g2974)) + ((sk[22]) & (!g2931) & (!g99) & (g2974)) + ((sk[22]) & (!g2931) & (g99) & (!g2974)) + ((sk[22]) & (!g2931) & (g99) & (g2974)) + ((sk[22]) & (g2931) & (!g99) & (!g2974)) + ((sk[22]) & (g2931) & (!g99) & (g2974)) + ((sk[22]) & (g2931) & (g99) & (!g2974)) + ((sk[22]) & (g2931) & (g99) & (g2974)));
	assign g2976 = (((!sk[23]) & (!g84) & (!g95) & (!g100) & (g101) & (!g2959)) + ((!sk[23]) & (!g84) & (!g95) & (!g100) & (g101) & (g2959)) + ((!sk[23]) & (!g84) & (!g95) & (g100) & (!g101) & (!g2959)) + ((!sk[23]) & (!g84) & (!g95) & (g100) & (!g101) & (g2959)) + ((!sk[23]) & (!g84) & (!g95) & (g100) & (g101) & (!g2959)) + ((!sk[23]) & (!g84) & (!g95) & (g100) & (g101) & (g2959)) + ((!sk[23]) & (!g84) & (g95) & (!g100) & (g101) & (!g2959)) + ((!sk[23]) & (!g84) & (g95) & (!g100) & (g101) & (g2959)) + ((!sk[23]) & (!g84) & (g95) & (g100) & (!g101) & (!g2959)) + ((!sk[23]) & (!g84) & (g95) & (g100) & (!g101) & (g2959)) + ((!sk[23]) & (!g84) & (g95) & (g100) & (g101) & (!g2959)) + ((!sk[23]) & (!g84) & (g95) & (g100) & (g101) & (g2959)) + ((!sk[23]) & (g84) & (!g95) & (!g100) & (!g101) & (!g2959)) + ((!sk[23]) & (g84) & (!g95) & (!g100) & (!g101) & (g2959)) + ((!sk[23]) & (g84) & (!g95) & (!g100) & (g101) & (!g2959)) + ((!sk[23]) & (g84) & (!g95) & (!g100) & (g101) & (g2959)) + ((!sk[23]) & (g84) & (!g95) & (g100) & (!g101) & (!g2959)) + ((!sk[23]) & (g84) & (!g95) & (g100) & (!g101) & (g2959)) + ((!sk[23]) & (g84) & (!g95) & (g100) & (g101) & (!g2959)) + ((!sk[23]) & (g84) & (!g95) & (g100) & (g101) & (g2959)) + ((!sk[23]) & (g84) & (g95) & (!g100) & (!g101) & (!g2959)) + ((!sk[23]) & (g84) & (g95) & (!g100) & (!g101) & (g2959)) + ((!sk[23]) & (g84) & (g95) & (!g100) & (g101) & (!g2959)) + ((!sk[23]) & (g84) & (g95) & (!g100) & (g101) & (g2959)) + ((!sk[23]) & (g84) & (g95) & (g100) & (!g101) & (!g2959)) + ((!sk[23]) & (g84) & (g95) & (g100) & (!g101) & (g2959)) + ((!sk[23]) & (g84) & (g95) & (g100) & (g101) & (!g2959)) + ((!sk[23]) & (g84) & (g95) & (g100) & (g101) & (g2959)) + ((sk[23]) & (!g84) & (!g95) & (!g100) & (!g101) & (!g2959)) + ((sk[23]) & (!g84) & (!g95) & (!g100) & (!g101) & (g2959)) + ((sk[23]) & (!g84) & (!g95) & (!g100) & (g101) & (!g2959)) + ((sk[23]) & (!g84) & (!g95) & (!g100) & (g101) & (g2959)) + ((sk[23]) & (!g84) & (!g95) & (g100) & (!g101) & (!g2959)) + ((sk[23]) & (!g84) & (!g95) & (g100) & (g101) & (!g2959)) + ((sk[23]) & (!g84) & (!g95) & (g100) & (g101) & (g2959)) + ((sk[23]) & (!g84) & (g95) & (!g100) & (!g101) & (!g2959)) + ((sk[23]) & (!g84) & (g95) & (!g100) & (!g101) & (g2959)) + ((sk[23]) & (!g84) & (g95) & (!g100) & (g101) & (!g2959)) + ((sk[23]) & (!g84) & (g95) & (!g100) & (g101) & (g2959)) + ((sk[23]) & (!g84) & (g95) & (g100) & (!g101) & (!g2959)) + ((sk[23]) & (!g84) & (g95) & (g100) & (g101) & (!g2959)) + ((sk[23]) & (!g84) & (g95) & (g100) & (g101) & (g2959)) + ((sk[23]) & (g84) & (!g95) & (!g100) & (!g101) & (!g2959)) + ((sk[23]) & (g84) & (!g95) & (!g100) & (!g101) & (g2959)) + ((sk[23]) & (g84) & (!g95) & (!g100) & (g101) & (!g2959)) + ((sk[23]) & (g84) & (!g95) & (!g100) & (g101) & (g2959)) + ((sk[23]) & (g84) & (!g95) & (g100) & (!g101) & (!g2959)) + ((sk[23]) & (g84) & (!g95) & (g100) & (g101) & (!g2959)) + ((sk[23]) & (g84) & (!g95) & (g100) & (g101) & (g2959)) + ((sk[23]) & (g84) & (g95) & (!g100) & (!g101) & (!g2959)) + ((sk[23]) & (g84) & (g95) & (!g100) & (!g101) & (g2959)) + ((sk[23]) & (g84) & (g95) & (!g100) & (g101) & (!g2959)) + ((sk[23]) & (g84) & (g95) & (!g100) & (g101) & (g2959)) + ((sk[23]) & (g84) & (g95) & (g100) & (!g101) & (!g2959)) + ((sk[23]) & (g84) & (g95) & (g100) & (!g101) & (g2959)) + ((sk[23]) & (g84) & (g95) & (g100) & (g101) & (!g2959)) + ((sk[23]) & (g84) & (g95) & (g100) & (g101) & (g2959)));
	assign g2977 = (((!sk[24]) & (!g2928) & (g2024) & (!g2935)) + ((!sk[24]) & (!g2928) & (g2024) & (g2935)) + ((!sk[24]) & (g2928) & (!g2024) & (!g2935)) + ((!sk[24]) & (g2928) & (!g2024) & (g2935)) + ((!sk[24]) & (g2928) & (g2024) & (!g2935)) + ((!sk[24]) & (g2928) & (g2024) & (g2935)) + ((sk[24]) & (!g2928) & (g2024) & (g2935)) + ((sk[24]) & (g2928) & (!g2024) & (g2935)) + ((sk[24]) & (g2928) & (g2024) & (g2935)));
	assign g2978 = (((!sk[25]) & (!g2928) & (g2942)) + ((!sk[25]) & (g2928) & (g2942)) + ((sk[25]) & (!g2928) & (!g2942)));
	assign g2979 = (((!g911) & (!g2564) & (!g89) & (g2566) & (g2977) & (!g2978)) + ((!g911) & (!g2564) & (g89) & (!g2566) & (!g2977) & (!g2978)) + ((!g911) & (!g2564) & (g89) & (g2566) & (!g2977) & (!g2978)) + ((!g911) & (!g2564) & (g89) & (g2566) & (g2977) & (!g2978)) + ((!g911) & (g2564) & (!g89) & (!g2566) & (g2977) & (g2978)) + ((!g911) & (g2564) & (!g89) & (g2566) & (g2977) & (!g2978)) + ((!g911) & (g2564) & (!g89) & (g2566) & (g2977) & (g2978)) + ((!g911) & (g2564) & (g89) & (!g2566) & (!g2977) & (!g2978)) + ((!g911) & (g2564) & (g89) & (!g2566) & (g2977) & (g2978)) + ((!g911) & (g2564) & (g89) & (g2566) & (!g2977) & (!g2978)) + ((!g911) & (g2564) & (g89) & (g2566) & (g2977) & (!g2978)) + ((!g911) & (g2564) & (g89) & (g2566) & (g2977) & (g2978)) + ((g911) & (!g2564) & (!g89) & (!g2566) & (!g2977) & (g2978)) + ((g911) & (!g2564) & (!g89) & (g2566) & (!g2977) & (g2978)) + ((g911) & (!g2564) & (!g89) & (g2566) & (g2977) & (!g2978)) + ((g911) & (!g2564) & (g89) & (!g2566) & (!g2977) & (!g2978)) + ((g911) & (!g2564) & (g89) & (!g2566) & (!g2977) & (g2978)) + ((g911) & (!g2564) & (g89) & (g2566) & (!g2977) & (!g2978)) + ((g911) & (!g2564) & (g89) & (g2566) & (!g2977) & (g2978)) + ((g911) & (!g2564) & (g89) & (g2566) & (g2977) & (!g2978)) + ((g911) & (g2564) & (!g89) & (!g2566) & (!g2977) & (g2978)) + ((g911) & (g2564) & (!g89) & (!g2566) & (g2977) & (g2978)) + ((g911) & (g2564) & (!g89) & (g2566) & (!g2977) & (g2978)) + ((g911) & (g2564) & (!g89) & (g2566) & (g2977) & (!g2978)) + ((g911) & (g2564) & (!g89) & (g2566) & (g2977) & (g2978)) + ((g911) & (g2564) & (g89) & (!g2566) & (!g2977) & (!g2978)) + ((g911) & (g2564) & (g89) & (!g2566) & (!g2977) & (g2978)) + ((g911) & (g2564) & (g89) & (!g2566) & (g2977) & (g2978)) + ((g911) & (g2564) & (g89) & (g2566) & (!g2977) & (!g2978)) + ((g911) & (g2564) & (g89) & (g2566) & (!g2977) & (g2978)) + ((g911) & (g2564) & (g89) & (g2566) & (g2977) & (!g2978)) + ((g911) & (g2564) & (g89) & (g2566) & (g2977) & (g2978)));
	assign g2980 = (((!g2940) & (!sk[27]) & (g2948)) + ((!g2940) & (sk[27]) & (g2948)) + ((g2940) & (!sk[27]) & (g2948)));
	assign g2981 = (((!g2928) & (!g2024) & (!g2935) & (!g2942) & (!g2951) & (!g2980)) + ((!g2928) & (!g2024) & (!g2935) & (!g2942) & (g2951) & (!g2980)) + ((!g2928) & (!g2024) & (g2935) & (!g2942) & (!g2951) & (!g2980)) + ((!g2928) & (!g2024) & (g2935) & (!g2942) & (g2951) & (!g2980)) + ((!g2928) & (!g2024) & (g2935) & (!g2942) & (g2951) & (g2980)) + ((!g2928) & (g2024) & (!g2935) & (!g2942) & (!g2951) & (!g2980)) + ((!g2928) & (g2024) & (!g2935) & (!g2942) & (g2951) & (!g2980)) + ((g2928) & (!g2024) & (!g2935) & (!g2942) & (!g2951) & (!g2980)) + ((g2928) & (!g2024) & (!g2935) & (!g2942) & (g2951) & (!g2980)) + ((g2928) & (!g2024) & (g2935) & (!g2942) & (g2951) & (!g2980)) + ((g2928) & (!g2024) & (g2935) & (!g2942) & (g2951) & (g2980)) + ((g2928) & (g2024) & (!g2935) & (!g2942) & (!g2951) & (!g2980)) + ((g2928) & (g2024) & (!g2935) & (!g2942) & (g2951) & (!g2980)));
	assign g2982 = (((!g2979) & (!sk[29]) & (g2981)) + ((g2979) & (!sk[29]) & (g2981)) + ((g2979) & (sk[29]) & (!g2981)));
	assign g2983 = (((!g959) & (!g2584) & (!g88) & (g2587) & (g2977) & (!g2978)) + ((!g959) & (!g2584) & (g88) & (!g2587) & (!g2977) & (!g2978)) + ((!g959) & (!g2584) & (g88) & (g2587) & (!g2977) & (!g2978)) + ((!g959) & (!g2584) & (g88) & (g2587) & (g2977) & (!g2978)) + ((!g959) & (g2584) & (!g88) & (!g2587) & (g2977) & (g2978)) + ((!g959) & (g2584) & (!g88) & (g2587) & (g2977) & (!g2978)) + ((!g959) & (g2584) & (!g88) & (g2587) & (g2977) & (g2978)) + ((!g959) & (g2584) & (g88) & (!g2587) & (!g2977) & (!g2978)) + ((!g959) & (g2584) & (g88) & (!g2587) & (g2977) & (g2978)) + ((!g959) & (g2584) & (g88) & (g2587) & (!g2977) & (!g2978)) + ((!g959) & (g2584) & (g88) & (g2587) & (g2977) & (!g2978)) + ((!g959) & (g2584) & (g88) & (g2587) & (g2977) & (g2978)) + ((g959) & (!g2584) & (!g88) & (!g2587) & (!g2977) & (g2978)) + ((g959) & (!g2584) & (!g88) & (g2587) & (!g2977) & (g2978)) + ((g959) & (!g2584) & (!g88) & (g2587) & (g2977) & (!g2978)) + ((g959) & (!g2584) & (g88) & (!g2587) & (!g2977) & (!g2978)) + ((g959) & (!g2584) & (g88) & (!g2587) & (!g2977) & (g2978)) + ((g959) & (!g2584) & (g88) & (g2587) & (!g2977) & (!g2978)) + ((g959) & (!g2584) & (g88) & (g2587) & (!g2977) & (g2978)) + ((g959) & (!g2584) & (g88) & (g2587) & (g2977) & (!g2978)) + ((g959) & (g2584) & (!g88) & (!g2587) & (!g2977) & (g2978)) + ((g959) & (g2584) & (!g88) & (!g2587) & (g2977) & (g2978)) + ((g959) & (g2584) & (!g88) & (g2587) & (!g2977) & (g2978)) + ((g959) & (g2584) & (!g88) & (g2587) & (g2977) & (!g2978)) + ((g959) & (g2584) & (!g88) & (g2587) & (g2977) & (g2978)) + ((g959) & (g2584) & (g88) & (!g2587) & (!g2977) & (!g2978)) + ((g959) & (g2584) & (g88) & (!g2587) & (!g2977) & (g2978)) + ((g959) & (g2584) & (g88) & (!g2587) & (g2977) & (g2978)) + ((g959) & (g2584) & (g88) & (g2587) & (!g2977) & (!g2978)) + ((g959) & (g2584) & (g88) & (g2587) & (!g2977) & (g2978)) + ((g959) & (g2584) & (g88) & (g2587) & (g2977) & (!g2978)) + ((g959) & (g2584) & (g88) & (g2587) & (g2977) & (g2978)));
	assign g2984 = (((!sk[31]) & (!g2981) & (g2983)) + ((!sk[31]) & (g2981) & (g2983)) + ((sk[31]) & (!g2981) & (g2983)));
	assign g2985 = (((!g1004) & (!g2599) & (!g87) & (g2605) & (g2977) & (!g2978)) + ((!g1004) & (!g2599) & (g87) & (!g2605) & (!g2977) & (!g2978)) + ((!g1004) & (!g2599) & (g87) & (g2605) & (!g2977) & (!g2978)) + ((!g1004) & (!g2599) & (g87) & (g2605) & (g2977) & (!g2978)) + ((!g1004) & (g2599) & (!g87) & (!g2605) & (g2977) & (g2978)) + ((!g1004) & (g2599) & (!g87) & (g2605) & (g2977) & (!g2978)) + ((!g1004) & (g2599) & (!g87) & (g2605) & (g2977) & (g2978)) + ((!g1004) & (g2599) & (g87) & (!g2605) & (!g2977) & (!g2978)) + ((!g1004) & (g2599) & (g87) & (!g2605) & (g2977) & (g2978)) + ((!g1004) & (g2599) & (g87) & (g2605) & (!g2977) & (!g2978)) + ((!g1004) & (g2599) & (g87) & (g2605) & (g2977) & (!g2978)) + ((!g1004) & (g2599) & (g87) & (g2605) & (g2977) & (g2978)) + ((g1004) & (!g2599) & (!g87) & (!g2605) & (!g2977) & (g2978)) + ((g1004) & (!g2599) & (!g87) & (g2605) & (!g2977) & (g2978)) + ((g1004) & (!g2599) & (!g87) & (g2605) & (g2977) & (!g2978)) + ((g1004) & (!g2599) & (g87) & (!g2605) & (!g2977) & (!g2978)) + ((g1004) & (!g2599) & (g87) & (!g2605) & (!g2977) & (g2978)) + ((g1004) & (!g2599) & (g87) & (g2605) & (!g2977) & (!g2978)) + ((g1004) & (!g2599) & (g87) & (g2605) & (!g2977) & (g2978)) + ((g1004) & (!g2599) & (g87) & (g2605) & (g2977) & (!g2978)) + ((g1004) & (g2599) & (!g87) & (!g2605) & (!g2977) & (g2978)) + ((g1004) & (g2599) & (!g87) & (!g2605) & (g2977) & (g2978)) + ((g1004) & (g2599) & (!g87) & (g2605) & (!g2977) & (g2978)) + ((g1004) & (g2599) & (!g87) & (g2605) & (g2977) & (!g2978)) + ((g1004) & (g2599) & (!g87) & (g2605) & (g2977) & (g2978)) + ((g1004) & (g2599) & (g87) & (!g2605) & (!g2977) & (!g2978)) + ((g1004) & (g2599) & (g87) & (!g2605) & (!g2977) & (g2978)) + ((g1004) & (g2599) & (g87) & (!g2605) & (g2977) & (g2978)) + ((g1004) & (g2599) & (g87) & (g2605) & (!g2977) & (!g2978)) + ((g1004) & (g2599) & (g87) & (g2605) & (!g2977) & (g2978)) + ((g1004) & (g2599) & (g87) & (g2605) & (g2977) & (!g2978)) + ((g1004) & (g2599) & (g87) & (g2605) & (g2977) & (g2978)));
	assign g2986 = (((!g2981) & (!sk[33]) & (g2985)) + ((!g2981) & (sk[33]) & (g2985)) + ((g2981) & (!sk[33]) & (g2985)));
	assign g2987 = (((!g1049) & (!g2620) & (!g90) & (g2622) & (g2977) & (!g2978)) + ((!g1049) & (!g2620) & (g90) & (!g2622) & (!g2977) & (!g2978)) + ((!g1049) & (!g2620) & (g90) & (g2622) & (!g2977) & (!g2978)) + ((!g1049) & (!g2620) & (g90) & (g2622) & (g2977) & (!g2978)) + ((!g1049) & (g2620) & (!g90) & (!g2622) & (g2977) & (g2978)) + ((!g1049) & (g2620) & (!g90) & (g2622) & (g2977) & (!g2978)) + ((!g1049) & (g2620) & (!g90) & (g2622) & (g2977) & (g2978)) + ((!g1049) & (g2620) & (g90) & (!g2622) & (!g2977) & (!g2978)) + ((!g1049) & (g2620) & (g90) & (!g2622) & (g2977) & (g2978)) + ((!g1049) & (g2620) & (g90) & (g2622) & (!g2977) & (!g2978)) + ((!g1049) & (g2620) & (g90) & (g2622) & (g2977) & (!g2978)) + ((!g1049) & (g2620) & (g90) & (g2622) & (g2977) & (g2978)) + ((g1049) & (!g2620) & (!g90) & (!g2622) & (!g2977) & (g2978)) + ((g1049) & (!g2620) & (!g90) & (g2622) & (!g2977) & (g2978)) + ((g1049) & (!g2620) & (!g90) & (g2622) & (g2977) & (!g2978)) + ((g1049) & (!g2620) & (g90) & (!g2622) & (!g2977) & (!g2978)) + ((g1049) & (!g2620) & (g90) & (!g2622) & (!g2977) & (g2978)) + ((g1049) & (!g2620) & (g90) & (g2622) & (!g2977) & (!g2978)) + ((g1049) & (!g2620) & (g90) & (g2622) & (!g2977) & (g2978)) + ((g1049) & (!g2620) & (g90) & (g2622) & (g2977) & (!g2978)) + ((g1049) & (g2620) & (!g90) & (!g2622) & (!g2977) & (g2978)) + ((g1049) & (g2620) & (!g90) & (!g2622) & (g2977) & (g2978)) + ((g1049) & (g2620) & (!g90) & (g2622) & (!g2977) & (g2978)) + ((g1049) & (g2620) & (!g90) & (g2622) & (g2977) & (!g2978)) + ((g1049) & (g2620) & (!g90) & (g2622) & (g2977) & (g2978)) + ((g1049) & (g2620) & (g90) & (!g2622) & (!g2977) & (!g2978)) + ((g1049) & (g2620) & (g90) & (!g2622) & (!g2977) & (g2978)) + ((g1049) & (g2620) & (g90) & (!g2622) & (g2977) & (g2978)) + ((g1049) & (g2620) & (g90) & (g2622) & (!g2977) & (!g2978)) + ((g1049) & (g2620) & (g90) & (g2622) & (!g2977) & (g2978)) + ((g1049) & (g2620) & (g90) & (g2622) & (g2977) & (!g2978)) + ((g1049) & (g2620) & (g90) & (g2622) & (g2977) & (g2978)));
	assign g2988 = (((!sk[35]) & (!g2981) & (g2987)) + ((!sk[35]) & (g2981) & (g2987)) + ((sk[35]) & (!g2981) & (g2987)));
	assign g2989 = (((!g1274) & (!g2710) & (!g92) & (g2712) & (g2977) & (!g2978)) + ((!g1274) & (!g2710) & (g92) & (!g2712) & (!g2977) & (!g2978)) + ((!g1274) & (!g2710) & (g92) & (g2712) & (!g2977) & (!g2978)) + ((!g1274) & (!g2710) & (g92) & (g2712) & (g2977) & (!g2978)) + ((!g1274) & (g2710) & (!g92) & (!g2712) & (g2977) & (g2978)) + ((!g1274) & (g2710) & (!g92) & (g2712) & (g2977) & (!g2978)) + ((!g1274) & (g2710) & (!g92) & (g2712) & (g2977) & (g2978)) + ((!g1274) & (g2710) & (g92) & (!g2712) & (!g2977) & (!g2978)) + ((!g1274) & (g2710) & (g92) & (!g2712) & (g2977) & (g2978)) + ((!g1274) & (g2710) & (g92) & (g2712) & (!g2977) & (!g2978)) + ((!g1274) & (g2710) & (g92) & (g2712) & (g2977) & (!g2978)) + ((!g1274) & (g2710) & (g92) & (g2712) & (g2977) & (g2978)) + ((g1274) & (!g2710) & (!g92) & (!g2712) & (!g2977) & (g2978)) + ((g1274) & (!g2710) & (!g92) & (g2712) & (!g2977) & (g2978)) + ((g1274) & (!g2710) & (!g92) & (g2712) & (g2977) & (!g2978)) + ((g1274) & (!g2710) & (g92) & (!g2712) & (!g2977) & (!g2978)) + ((g1274) & (!g2710) & (g92) & (!g2712) & (!g2977) & (g2978)) + ((g1274) & (!g2710) & (g92) & (g2712) & (!g2977) & (!g2978)) + ((g1274) & (!g2710) & (g92) & (g2712) & (!g2977) & (g2978)) + ((g1274) & (!g2710) & (g92) & (g2712) & (g2977) & (!g2978)) + ((g1274) & (g2710) & (!g92) & (!g2712) & (!g2977) & (g2978)) + ((g1274) & (g2710) & (!g92) & (!g2712) & (g2977) & (g2978)) + ((g1274) & (g2710) & (!g92) & (g2712) & (!g2977) & (g2978)) + ((g1274) & (g2710) & (!g92) & (g2712) & (g2977) & (!g2978)) + ((g1274) & (g2710) & (!g92) & (g2712) & (g2977) & (g2978)) + ((g1274) & (g2710) & (g92) & (!g2712) & (!g2977) & (!g2978)) + ((g1274) & (g2710) & (g92) & (!g2712) & (!g2977) & (g2978)) + ((g1274) & (g2710) & (g92) & (!g2712) & (g2977) & (g2978)) + ((g1274) & (g2710) & (g92) & (g2712) & (!g2977) & (!g2978)) + ((g1274) & (g2710) & (g92) & (g2712) & (!g2977) & (g2978)) + ((g1274) & (g2710) & (g92) & (g2712) & (g2977) & (!g2978)) + ((g1274) & (g2710) & (g92) & (g2712) & (g2977) & (g2978)));
	assign g2990 = (((!sk[37]) & (!g2981) & (g2989)) + ((!sk[37]) & (g2981) & (g2989)) + ((sk[37]) & (!g2981) & (g2989)));
	assign g2991 = (((!g1319) & (!g2728) & (!g91) & (g2731) & (g2977) & (!g2978)) + ((!g1319) & (!g2728) & (g91) & (!g2731) & (!g2977) & (!g2978)) + ((!g1319) & (!g2728) & (g91) & (g2731) & (!g2977) & (!g2978)) + ((!g1319) & (!g2728) & (g91) & (g2731) & (g2977) & (!g2978)) + ((!g1319) & (g2728) & (!g91) & (!g2731) & (g2977) & (g2978)) + ((!g1319) & (g2728) & (!g91) & (g2731) & (g2977) & (!g2978)) + ((!g1319) & (g2728) & (!g91) & (g2731) & (g2977) & (g2978)) + ((!g1319) & (g2728) & (g91) & (!g2731) & (!g2977) & (!g2978)) + ((!g1319) & (g2728) & (g91) & (!g2731) & (g2977) & (g2978)) + ((!g1319) & (g2728) & (g91) & (g2731) & (!g2977) & (!g2978)) + ((!g1319) & (g2728) & (g91) & (g2731) & (g2977) & (!g2978)) + ((!g1319) & (g2728) & (g91) & (g2731) & (g2977) & (g2978)) + ((g1319) & (!g2728) & (!g91) & (!g2731) & (!g2977) & (g2978)) + ((g1319) & (!g2728) & (!g91) & (g2731) & (!g2977) & (g2978)) + ((g1319) & (!g2728) & (!g91) & (g2731) & (g2977) & (!g2978)) + ((g1319) & (!g2728) & (g91) & (!g2731) & (!g2977) & (!g2978)) + ((g1319) & (!g2728) & (g91) & (!g2731) & (!g2977) & (g2978)) + ((g1319) & (!g2728) & (g91) & (g2731) & (!g2977) & (!g2978)) + ((g1319) & (!g2728) & (g91) & (g2731) & (!g2977) & (g2978)) + ((g1319) & (!g2728) & (g91) & (g2731) & (g2977) & (!g2978)) + ((g1319) & (g2728) & (!g91) & (!g2731) & (!g2977) & (g2978)) + ((g1319) & (g2728) & (!g91) & (!g2731) & (g2977) & (g2978)) + ((g1319) & (g2728) & (!g91) & (g2731) & (!g2977) & (g2978)) + ((g1319) & (g2728) & (!g91) & (g2731) & (g2977) & (!g2978)) + ((g1319) & (g2728) & (!g91) & (g2731) & (g2977) & (g2978)) + ((g1319) & (g2728) & (g91) & (!g2731) & (!g2977) & (!g2978)) + ((g1319) & (g2728) & (g91) & (!g2731) & (!g2977) & (g2978)) + ((g1319) & (g2728) & (g91) & (!g2731) & (g2977) & (g2978)) + ((g1319) & (g2728) & (g91) & (g2731) & (!g2977) & (!g2978)) + ((g1319) & (g2728) & (g91) & (g2731) & (!g2977) & (g2978)) + ((g1319) & (g2728) & (g91) & (g2731) & (g2977) & (!g2978)) + ((g1319) & (g2728) & (g91) & (g2731) & (g2977) & (g2978)));
	assign g2992 = (((!g2981) & (!sk[39]) & (g2991)) + ((!g2981) & (sk[39]) & (g2991)) + ((g2981) & (!sk[39]) & (g2991)));
	assign g2993 = (((!g1364) & (!g2746) & (!g586) & (g2748) & (g2977) & (!g2978)) + ((!g1364) & (!g2746) & (g586) & (!g2748) & (!g2977) & (!g2978)) + ((!g1364) & (!g2746) & (g586) & (g2748) & (!g2977) & (!g2978)) + ((!g1364) & (!g2746) & (g586) & (g2748) & (g2977) & (!g2978)) + ((!g1364) & (g2746) & (!g586) & (!g2748) & (g2977) & (g2978)) + ((!g1364) & (g2746) & (!g586) & (g2748) & (g2977) & (!g2978)) + ((!g1364) & (g2746) & (!g586) & (g2748) & (g2977) & (g2978)) + ((!g1364) & (g2746) & (g586) & (!g2748) & (!g2977) & (!g2978)) + ((!g1364) & (g2746) & (g586) & (!g2748) & (g2977) & (g2978)) + ((!g1364) & (g2746) & (g586) & (g2748) & (!g2977) & (!g2978)) + ((!g1364) & (g2746) & (g586) & (g2748) & (g2977) & (!g2978)) + ((!g1364) & (g2746) & (g586) & (g2748) & (g2977) & (g2978)) + ((g1364) & (!g2746) & (!g586) & (!g2748) & (!g2977) & (g2978)) + ((g1364) & (!g2746) & (!g586) & (g2748) & (!g2977) & (g2978)) + ((g1364) & (!g2746) & (!g586) & (g2748) & (g2977) & (!g2978)) + ((g1364) & (!g2746) & (g586) & (!g2748) & (!g2977) & (!g2978)) + ((g1364) & (!g2746) & (g586) & (!g2748) & (!g2977) & (g2978)) + ((g1364) & (!g2746) & (g586) & (g2748) & (!g2977) & (!g2978)) + ((g1364) & (!g2746) & (g586) & (g2748) & (!g2977) & (g2978)) + ((g1364) & (!g2746) & (g586) & (g2748) & (g2977) & (!g2978)) + ((g1364) & (g2746) & (!g586) & (!g2748) & (!g2977) & (g2978)) + ((g1364) & (g2746) & (!g586) & (!g2748) & (g2977) & (g2978)) + ((g1364) & (g2746) & (!g586) & (g2748) & (!g2977) & (g2978)) + ((g1364) & (g2746) & (!g586) & (g2748) & (g2977) & (!g2978)) + ((g1364) & (g2746) & (!g586) & (g2748) & (g2977) & (g2978)) + ((g1364) & (g2746) & (g586) & (!g2748) & (!g2977) & (!g2978)) + ((g1364) & (g2746) & (g586) & (!g2748) & (!g2977) & (g2978)) + ((g1364) & (g2746) & (g586) & (!g2748) & (g2977) & (g2978)) + ((g1364) & (g2746) & (g586) & (g2748) & (!g2977) & (!g2978)) + ((g1364) & (g2746) & (g586) & (g2748) & (!g2977) & (g2978)) + ((g1364) & (g2746) & (g586) & (g2748) & (g2977) & (!g2978)) + ((g1364) & (g2746) & (g586) & (g2748) & (g2977) & (g2978)));
	assign g2994 = (((!sk[41]) & (!g2981) & (g2993)) + ((!sk[41]) & (g2981) & (g2993)) + ((sk[41]) & (!g2981) & (g2993)));
	assign g2995 = (((!g1409) & (!g2764) & (!g677) & (g2767) & (g2977) & (!g2978)) + ((!g1409) & (!g2764) & (g677) & (!g2767) & (!g2977) & (!g2978)) + ((!g1409) & (!g2764) & (g677) & (g2767) & (!g2977) & (!g2978)) + ((!g1409) & (!g2764) & (g677) & (g2767) & (g2977) & (!g2978)) + ((!g1409) & (g2764) & (!g677) & (!g2767) & (g2977) & (g2978)) + ((!g1409) & (g2764) & (!g677) & (g2767) & (g2977) & (!g2978)) + ((!g1409) & (g2764) & (!g677) & (g2767) & (g2977) & (g2978)) + ((!g1409) & (g2764) & (g677) & (!g2767) & (!g2977) & (!g2978)) + ((!g1409) & (g2764) & (g677) & (!g2767) & (g2977) & (g2978)) + ((!g1409) & (g2764) & (g677) & (g2767) & (!g2977) & (!g2978)) + ((!g1409) & (g2764) & (g677) & (g2767) & (g2977) & (!g2978)) + ((!g1409) & (g2764) & (g677) & (g2767) & (g2977) & (g2978)) + ((g1409) & (!g2764) & (!g677) & (!g2767) & (!g2977) & (g2978)) + ((g1409) & (!g2764) & (!g677) & (g2767) & (!g2977) & (g2978)) + ((g1409) & (!g2764) & (!g677) & (g2767) & (g2977) & (!g2978)) + ((g1409) & (!g2764) & (g677) & (!g2767) & (!g2977) & (!g2978)) + ((g1409) & (!g2764) & (g677) & (!g2767) & (!g2977) & (g2978)) + ((g1409) & (!g2764) & (g677) & (g2767) & (!g2977) & (!g2978)) + ((g1409) & (!g2764) & (g677) & (g2767) & (!g2977) & (g2978)) + ((g1409) & (!g2764) & (g677) & (g2767) & (g2977) & (!g2978)) + ((g1409) & (g2764) & (!g677) & (!g2767) & (!g2977) & (g2978)) + ((g1409) & (g2764) & (!g677) & (!g2767) & (g2977) & (g2978)) + ((g1409) & (g2764) & (!g677) & (g2767) & (!g2977) & (g2978)) + ((g1409) & (g2764) & (!g677) & (g2767) & (g2977) & (!g2978)) + ((g1409) & (g2764) & (!g677) & (g2767) & (g2977) & (g2978)) + ((g1409) & (g2764) & (g677) & (!g2767) & (!g2977) & (!g2978)) + ((g1409) & (g2764) & (g677) & (!g2767) & (!g2977) & (g2978)) + ((g1409) & (g2764) & (g677) & (!g2767) & (g2977) & (g2978)) + ((g1409) & (g2764) & (g677) & (g2767) & (!g2977) & (!g2978)) + ((g1409) & (g2764) & (g677) & (g2767) & (!g2977) & (g2978)) + ((g1409) & (g2764) & (g677) & (g2767) & (g2977) & (!g2978)) + ((g1409) & (g2764) & (g677) & (g2767) & (g2977) & (g2978)));
	assign g2996 = (((!g2981) & (!sk[43]) & (g2995)) + ((!g2981) & (sk[43]) & (g2995)) + ((g2981) & (!sk[43]) & (g2995)));
	assign g2997 = (((!g1094) & (!g2636) & (!g318) & (g2639) & (g2977) & (!g2978)) + ((!g1094) & (!g2636) & (g318) & (!g2639) & (!g2977) & (!g2978)) + ((!g1094) & (!g2636) & (g318) & (g2639) & (!g2977) & (!g2978)) + ((!g1094) & (!g2636) & (g318) & (g2639) & (g2977) & (!g2978)) + ((!g1094) & (g2636) & (!g318) & (!g2639) & (g2977) & (g2978)) + ((!g1094) & (g2636) & (!g318) & (g2639) & (g2977) & (!g2978)) + ((!g1094) & (g2636) & (!g318) & (g2639) & (g2977) & (g2978)) + ((!g1094) & (g2636) & (g318) & (!g2639) & (!g2977) & (!g2978)) + ((!g1094) & (g2636) & (g318) & (!g2639) & (g2977) & (g2978)) + ((!g1094) & (g2636) & (g318) & (g2639) & (!g2977) & (!g2978)) + ((!g1094) & (g2636) & (g318) & (g2639) & (g2977) & (!g2978)) + ((!g1094) & (g2636) & (g318) & (g2639) & (g2977) & (g2978)) + ((g1094) & (!g2636) & (!g318) & (!g2639) & (!g2977) & (g2978)) + ((g1094) & (!g2636) & (!g318) & (g2639) & (!g2977) & (g2978)) + ((g1094) & (!g2636) & (!g318) & (g2639) & (g2977) & (!g2978)) + ((g1094) & (!g2636) & (g318) & (!g2639) & (!g2977) & (!g2978)) + ((g1094) & (!g2636) & (g318) & (!g2639) & (!g2977) & (g2978)) + ((g1094) & (!g2636) & (g318) & (g2639) & (!g2977) & (!g2978)) + ((g1094) & (!g2636) & (g318) & (g2639) & (!g2977) & (g2978)) + ((g1094) & (!g2636) & (g318) & (g2639) & (g2977) & (!g2978)) + ((g1094) & (g2636) & (!g318) & (!g2639) & (!g2977) & (g2978)) + ((g1094) & (g2636) & (!g318) & (!g2639) & (g2977) & (g2978)) + ((g1094) & (g2636) & (!g318) & (g2639) & (!g2977) & (g2978)) + ((g1094) & (g2636) & (!g318) & (g2639) & (g2977) & (!g2978)) + ((g1094) & (g2636) & (!g318) & (g2639) & (g2977) & (g2978)) + ((g1094) & (g2636) & (g318) & (!g2639) & (!g2977) & (!g2978)) + ((g1094) & (g2636) & (g318) & (!g2639) & (!g2977) & (g2978)) + ((g1094) & (g2636) & (g318) & (!g2639) & (g2977) & (g2978)) + ((g1094) & (g2636) & (g318) & (g2639) & (!g2977) & (!g2978)) + ((g1094) & (g2636) & (g318) & (g2639) & (!g2977) & (g2978)) + ((g1094) & (g2636) & (g318) & (g2639) & (g2977) & (!g2978)) + ((g1094) & (g2636) & (g318) & (g2639) & (g2977) & (g2978)));
	assign g2998 = (((!sk[45]) & (!g2981) & (g2997)) + ((!sk[45]) & (g2981) & (g2997)) + ((sk[45]) & (!g2981) & (g2997)));
	assign g2999 = (((!g1139) & (!g2654) & (!g364) & (g2657) & (g2977) & (!g2978)) + ((!g1139) & (!g2654) & (g364) & (!g2657) & (!g2977) & (!g2978)) + ((!g1139) & (!g2654) & (g364) & (g2657) & (!g2977) & (!g2978)) + ((!g1139) & (!g2654) & (g364) & (g2657) & (g2977) & (!g2978)) + ((!g1139) & (g2654) & (!g364) & (!g2657) & (g2977) & (g2978)) + ((!g1139) & (g2654) & (!g364) & (g2657) & (g2977) & (!g2978)) + ((!g1139) & (g2654) & (!g364) & (g2657) & (g2977) & (g2978)) + ((!g1139) & (g2654) & (g364) & (!g2657) & (!g2977) & (!g2978)) + ((!g1139) & (g2654) & (g364) & (!g2657) & (g2977) & (g2978)) + ((!g1139) & (g2654) & (g364) & (g2657) & (!g2977) & (!g2978)) + ((!g1139) & (g2654) & (g364) & (g2657) & (g2977) & (!g2978)) + ((!g1139) & (g2654) & (g364) & (g2657) & (g2977) & (g2978)) + ((g1139) & (!g2654) & (!g364) & (!g2657) & (!g2977) & (g2978)) + ((g1139) & (!g2654) & (!g364) & (g2657) & (!g2977) & (g2978)) + ((g1139) & (!g2654) & (!g364) & (g2657) & (g2977) & (!g2978)) + ((g1139) & (!g2654) & (g364) & (!g2657) & (!g2977) & (!g2978)) + ((g1139) & (!g2654) & (g364) & (!g2657) & (!g2977) & (g2978)) + ((g1139) & (!g2654) & (g364) & (g2657) & (!g2977) & (!g2978)) + ((g1139) & (!g2654) & (g364) & (g2657) & (!g2977) & (g2978)) + ((g1139) & (!g2654) & (g364) & (g2657) & (g2977) & (!g2978)) + ((g1139) & (g2654) & (!g364) & (!g2657) & (!g2977) & (g2978)) + ((g1139) & (g2654) & (!g364) & (!g2657) & (g2977) & (g2978)) + ((g1139) & (g2654) & (!g364) & (g2657) & (!g2977) & (g2978)) + ((g1139) & (g2654) & (!g364) & (g2657) & (g2977) & (!g2978)) + ((g1139) & (g2654) & (!g364) & (g2657) & (g2977) & (g2978)) + ((g1139) & (g2654) & (g364) & (!g2657) & (!g2977) & (!g2978)) + ((g1139) & (g2654) & (g364) & (!g2657) & (!g2977) & (g2978)) + ((g1139) & (g2654) & (g364) & (!g2657) & (g2977) & (g2978)) + ((g1139) & (g2654) & (g364) & (g2657) & (!g2977) & (!g2978)) + ((g1139) & (g2654) & (g364) & (g2657) & (!g2977) & (g2978)) + ((g1139) & (g2654) & (g364) & (g2657) & (g2977) & (!g2978)) + ((g1139) & (g2654) & (g364) & (g2657) & (g2977) & (g2978)));
	assign g3000 = (((!g2981) & (!sk[47]) & (g2999)) + ((!g2981) & (sk[47]) & (g2999)) + ((g2981) & (!sk[47]) & (g2999)));
	assign g3001 = (((!g1184) & (!g2674) & (!g86) & (g2677) & (g2977) & (!g2978)) + ((!g1184) & (!g2674) & (g86) & (!g2677) & (!g2977) & (!g2978)) + ((!g1184) & (!g2674) & (g86) & (g2677) & (!g2977) & (!g2978)) + ((!g1184) & (!g2674) & (g86) & (g2677) & (g2977) & (!g2978)) + ((!g1184) & (g2674) & (!g86) & (!g2677) & (g2977) & (g2978)) + ((!g1184) & (g2674) & (!g86) & (g2677) & (g2977) & (!g2978)) + ((!g1184) & (g2674) & (!g86) & (g2677) & (g2977) & (g2978)) + ((!g1184) & (g2674) & (g86) & (!g2677) & (!g2977) & (!g2978)) + ((!g1184) & (g2674) & (g86) & (!g2677) & (g2977) & (g2978)) + ((!g1184) & (g2674) & (g86) & (g2677) & (!g2977) & (!g2978)) + ((!g1184) & (g2674) & (g86) & (g2677) & (g2977) & (!g2978)) + ((!g1184) & (g2674) & (g86) & (g2677) & (g2977) & (g2978)) + ((g1184) & (!g2674) & (!g86) & (!g2677) & (!g2977) & (g2978)) + ((g1184) & (!g2674) & (!g86) & (g2677) & (!g2977) & (g2978)) + ((g1184) & (!g2674) & (!g86) & (g2677) & (g2977) & (!g2978)) + ((g1184) & (!g2674) & (g86) & (!g2677) & (!g2977) & (!g2978)) + ((g1184) & (!g2674) & (g86) & (!g2677) & (!g2977) & (g2978)) + ((g1184) & (!g2674) & (g86) & (g2677) & (!g2977) & (!g2978)) + ((g1184) & (!g2674) & (g86) & (g2677) & (!g2977) & (g2978)) + ((g1184) & (!g2674) & (g86) & (g2677) & (g2977) & (!g2978)) + ((g1184) & (g2674) & (!g86) & (!g2677) & (!g2977) & (g2978)) + ((g1184) & (g2674) & (!g86) & (!g2677) & (g2977) & (g2978)) + ((g1184) & (g2674) & (!g86) & (g2677) & (!g2977) & (g2978)) + ((g1184) & (g2674) & (!g86) & (g2677) & (g2977) & (!g2978)) + ((g1184) & (g2674) & (!g86) & (g2677) & (g2977) & (g2978)) + ((g1184) & (g2674) & (g86) & (!g2677) & (!g2977) & (!g2978)) + ((g1184) & (g2674) & (g86) & (!g2677) & (!g2977) & (g2978)) + ((g1184) & (g2674) & (g86) & (!g2677) & (g2977) & (g2978)) + ((g1184) & (g2674) & (g86) & (g2677) & (!g2977) & (!g2978)) + ((g1184) & (g2674) & (g86) & (g2677) & (!g2977) & (g2978)) + ((g1184) & (g2674) & (g86) & (g2677) & (g2977) & (!g2978)) + ((g1184) & (g2674) & (g86) & (g2677) & (g2977) & (g2978)));
	assign g3002 = (((!sk[49]) & (!g2981) & (g3001)) + ((!sk[49]) & (g2981) & (g3001)) + ((sk[49]) & (!g2981) & (g3001)));
	assign g3003 = (((!g1229) & (!g2691) & (!g85) & (g2696) & (g2977) & (!g2978)) + ((!g1229) & (!g2691) & (g85) & (!g2696) & (!g2977) & (!g2978)) + ((!g1229) & (!g2691) & (g85) & (g2696) & (!g2977) & (!g2978)) + ((!g1229) & (!g2691) & (g85) & (g2696) & (g2977) & (!g2978)) + ((!g1229) & (g2691) & (!g85) & (!g2696) & (g2977) & (g2978)) + ((!g1229) & (g2691) & (!g85) & (g2696) & (g2977) & (!g2978)) + ((!g1229) & (g2691) & (!g85) & (g2696) & (g2977) & (g2978)) + ((!g1229) & (g2691) & (g85) & (!g2696) & (!g2977) & (!g2978)) + ((!g1229) & (g2691) & (g85) & (!g2696) & (g2977) & (g2978)) + ((!g1229) & (g2691) & (g85) & (g2696) & (!g2977) & (!g2978)) + ((!g1229) & (g2691) & (g85) & (g2696) & (g2977) & (!g2978)) + ((!g1229) & (g2691) & (g85) & (g2696) & (g2977) & (g2978)) + ((g1229) & (!g2691) & (!g85) & (!g2696) & (!g2977) & (g2978)) + ((g1229) & (!g2691) & (!g85) & (g2696) & (!g2977) & (g2978)) + ((g1229) & (!g2691) & (!g85) & (g2696) & (g2977) & (!g2978)) + ((g1229) & (!g2691) & (g85) & (!g2696) & (!g2977) & (!g2978)) + ((g1229) & (!g2691) & (g85) & (!g2696) & (!g2977) & (g2978)) + ((g1229) & (!g2691) & (g85) & (g2696) & (!g2977) & (!g2978)) + ((g1229) & (!g2691) & (g85) & (g2696) & (!g2977) & (g2978)) + ((g1229) & (!g2691) & (g85) & (g2696) & (g2977) & (!g2978)) + ((g1229) & (g2691) & (!g85) & (!g2696) & (!g2977) & (g2978)) + ((g1229) & (g2691) & (!g85) & (!g2696) & (g2977) & (g2978)) + ((g1229) & (g2691) & (!g85) & (g2696) & (!g2977) & (g2978)) + ((g1229) & (g2691) & (!g85) & (g2696) & (g2977) & (!g2978)) + ((g1229) & (g2691) & (!g85) & (g2696) & (g2977) & (g2978)) + ((g1229) & (g2691) & (g85) & (!g2696) & (!g2977) & (!g2978)) + ((g1229) & (g2691) & (g85) & (!g2696) & (!g2977) & (g2978)) + ((g1229) & (g2691) & (g85) & (!g2696) & (g2977) & (g2978)) + ((g1229) & (g2691) & (g85) & (g2696) & (!g2977) & (!g2978)) + ((g1229) & (g2691) & (g85) & (g2696) & (!g2977) & (g2978)) + ((g1229) & (g2691) & (g85) & (g2696) & (g2977) & (!g2978)) + ((g1229) & (g2691) & (g85) & (g2696) & (g2977) & (g2978)));
	assign g3004 = (((!sk[51]) & (!g2981) & (g3003)) + ((!sk[51]) & (g2981) & (g3003)) + ((sk[51]) & (!g2981) & (g3003)));
	assign g3005 = (((!g1454) & (!g2789) & (!g726) & (g2791) & (g2977) & (!g2978)) + ((!g1454) & (!g2789) & (g726) & (!g2791) & (!g2977) & (!g2978)) + ((!g1454) & (!g2789) & (g726) & (g2791) & (!g2977) & (!g2978)) + ((!g1454) & (!g2789) & (g726) & (g2791) & (g2977) & (!g2978)) + ((!g1454) & (g2789) & (!g726) & (!g2791) & (g2977) & (g2978)) + ((!g1454) & (g2789) & (!g726) & (g2791) & (g2977) & (!g2978)) + ((!g1454) & (g2789) & (!g726) & (g2791) & (g2977) & (g2978)) + ((!g1454) & (g2789) & (g726) & (!g2791) & (!g2977) & (!g2978)) + ((!g1454) & (g2789) & (g726) & (!g2791) & (g2977) & (g2978)) + ((!g1454) & (g2789) & (g726) & (g2791) & (!g2977) & (!g2978)) + ((!g1454) & (g2789) & (g726) & (g2791) & (g2977) & (!g2978)) + ((!g1454) & (g2789) & (g726) & (g2791) & (g2977) & (g2978)) + ((g1454) & (!g2789) & (!g726) & (!g2791) & (!g2977) & (g2978)) + ((g1454) & (!g2789) & (!g726) & (g2791) & (!g2977) & (g2978)) + ((g1454) & (!g2789) & (!g726) & (g2791) & (g2977) & (!g2978)) + ((g1454) & (!g2789) & (g726) & (!g2791) & (!g2977) & (!g2978)) + ((g1454) & (!g2789) & (g726) & (!g2791) & (!g2977) & (g2978)) + ((g1454) & (!g2789) & (g726) & (g2791) & (!g2977) & (!g2978)) + ((g1454) & (!g2789) & (g726) & (g2791) & (!g2977) & (g2978)) + ((g1454) & (!g2789) & (g726) & (g2791) & (g2977) & (!g2978)) + ((g1454) & (g2789) & (!g726) & (!g2791) & (!g2977) & (g2978)) + ((g1454) & (g2789) & (!g726) & (!g2791) & (g2977) & (g2978)) + ((g1454) & (g2789) & (!g726) & (g2791) & (!g2977) & (g2978)) + ((g1454) & (g2789) & (!g726) & (g2791) & (g2977) & (!g2978)) + ((g1454) & (g2789) & (!g726) & (g2791) & (g2977) & (g2978)) + ((g1454) & (g2789) & (g726) & (!g2791) & (!g2977) & (!g2978)) + ((g1454) & (g2789) & (g726) & (!g2791) & (!g2977) & (g2978)) + ((g1454) & (g2789) & (g726) & (!g2791) & (g2977) & (g2978)) + ((g1454) & (g2789) & (g726) & (g2791) & (!g2977) & (!g2978)) + ((g1454) & (g2789) & (g726) & (g2791) & (!g2977) & (g2978)) + ((g1454) & (g2789) & (g726) & (g2791) & (g2977) & (!g2978)) + ((g1454) & (g2789) & (g726) & (g2791) & (g2977) & (g2978)));
	assign g3006 = (((!sk[53]) & (!g2981) & (g3005)) + ((!sk[53]) & (g2981) & (g3005)) + ((sk[53]) & (!g2981) & (g3005)));
	assign g3007 = (((!g1499) & (!g2806) & (!g773) & (g2808) & (g2977) & (!g2978)) + ((!g1499) & (!g2806) & (g773) & (!g2808) & (!g2977) & (!g2978)) + ((!g1499) & (!g2806) & (g773) & (g2808) & (!g2977) & (!g2978)) + ((!g1499) & (!g2806) & (g773) & (g2808) & (g2977) & (!g2978)) + ((!g1499) & (g2806) & (!g773) & (!g2808) & (g2977) & (g2978)) + ((!g1499) & (g2806) & (!g773) & (g2808) & (g2977) & (!g2978)) + ((!g1499) & (g2806) & (!g773) & (g2808) & (g2977) & (g2978)) + ((!g1499) & (g2806) & (g773) & (!g2808) & (!g2977) & (!g2978)) + ((!g1499) & (g2806) & (g773) & (!g2808) & (g2977) & (g2978)) + ((!g1499) & (g2806) & (g773) & (g2808) & (!g2977) & (!g2978)) + ((!g1499) & (g2806) & (g773) & (g2808) & (g2977) & (!g2978)) + ((!g1499) & (g2806) & (g773) & (g2808) & (g2977) & (g2978)) + ((g1499) & (!g2806) & (!g773) & (!g2808) & (!g2977) & (g2978)) + ((g1499) & (!g2806) & (!g773) & (g2808) & (!g2977) & (g2978)) + ((g1499) & (!g2806) & (!g773) & (g2808) & (g2977) & (!g2978)) + ((g1499) & (!g2806) & (g773) & (!g2808) & (!g2977) & (!g2978)) + ((g1499) & (!g2806) & (g773) & (!g2808) & (!g2977) & (g2978)) + ((g1499) & (!g2806) & (g773) & (g2808) & (!g2977) & (!g2978)) + ((g1499) & (!g2806) & (g773) & (g2808) & (!g2977) & (g2978)) + ((g1499) & (!g2806) & (g773) & (g2808) & (g2977) & (!g2978)) + ((g1499) & (g2806) & (!g773) & (!g2808) & (!g2977) & (g2978)) + ((g1499) & (g2806) & (!g773) & (!g2808) & (g2977) & (g2978)) + ((g1499) & (g2806) & (!g773) & (g2808) & (!g2977) & (g2978)) + ((g1499) & (g2806) & (!g773) & (g2808) & (g2977) & (!g2978)) + ((g1499) & (g2806) & (!g773) & (g2808) & (g2977) & (g2978)) + ((g1499) & (g2806) & (g773) & (!g2808) & (!g2977) & (!g2978)) + ((g1499) & (g2806) & (g773) & (!g2808) & (!g2977) & (g2978)) + ((g1499) & (g2806) & (g773) & (!g2808) & (g2977) & (g2978)) + ((g1499) & (g2806) & (g773) & (g2808) & (!g2977) & (!g2978)) + ((g1499) & (g2806) & (g773) & (g2808) & (!g2977) & (g2978)) + ((g1499) & (g2806) & (g773) & (g2808) & (g2977) & (!g2978)) + ((g1499) & (g2806) & (g773) & (g2808) & (g2977) & (g2978)));
	assign g3008 = (((!g2981) & (!sk[55]) & (g3007)) + ((!g2981) & (sk[55]) & (g3007)) + ((g2981) & (!sk[55]) & (g3007)));
	assign g3009 = (((!g1543) & (!g2822) & (!g820) & (g2824) & (g2977) & (!g2978)) + ((!g1543) & (!g2822) & (g820) & (!g2824) & (!g2977) & (!g2978)) + ((!g1543) & (!g2822) & (g820) & (g2824) & (!g2977) & (!g2978)) + ((!g1543) & (!g2822) & (g820) & (g2824) & (g2977) & (!g2978)) + ((!g1543) & (g2822) & (!g820) & (!g2824) & (g2977) & (g2978)) + ((!g1543) & (g2822) & (!g820) & (g2824) & (g2977) & (!g2978)) + ((!g1543) & (g2822) & (!g820) & (g2824) & (g2977) & (g2978)) + ((!g1543) & (g2822) & (g820) & (!g2824) & (!g2977) & (!g2978)) + ((!g1543) & (g2822) & (g820) & (!g2824) & (g2977) & (g2978)) + ((!g1543) & (g2822) & (g820) & (g2824) & (!g2977) & (!g2978)) + ((!g1543) & (g2822) & (g820) & (g2824) & (g2977) & (!g2978)) + ((!g1543) & (g2822) & (g820) & (g2824) & (g2977) & (g2978)) + ((g1543) & (!g2822) & (!g820) & (!g2824) & (!g2977) & (g2978)) + ((g1543) & (!g2822) & (!g820) & (g2824) & (!g2977) & (g2978)) + ((g1543) & (!g2822) & (!g820) & (g2824) & (g2977) & (!g2978)) + ((g1543) & (!g2822) & (g820) & (!g2824) & (!g2977) & (!g2978)) + ((g1543) & (!g2822) & (g820) & (!g2824) & (!g2977) & (g2978)) + ((g1543) & (!g2822) & (g820) & (g2824) & (!g2977) & (!g2978)) + ((g1543) & (!g2822) & (g820) & (g2824) & (!g2977) & (g2978)) + ((g1543) & (!g2822) & (g820) & (g2824) & (g2977) & (!g2978)) + ((g1543) & (g2822) & (!g820) & (!g2824) & (!g2977) & (g2978)) + ((g1543) & (g2822) & (!g820) & (!g2824) & (g2977) & (g2978)) + ((g1543) & (g2822) & (!g820) & (g2824) & (!g2977) & (g2978)) + ((g1543) & (g2822) & (!g820) & (g2824) & (g2977) & (!g2978)) + ((g1543) & (g2822) & (!g820) & (g2824) & (g2977) & (g2978)) + ((g1543) & (g2822) & (g820) & (!g2824) & (!g2977) & (!g2978)) + ((g1543) & (g2822) & (g820) & (!g2824) & (!g2977) & (g2978)) + ((g1543) & (g2822) & (g820) & (!g2824) & (g2977) & (g2978)) + ((g1543) & (g2822) & (g820) & (g2824) & (!g2977) & (!g2978)) + ((g1543) & (g2822) & (g820) & (g2824) & (!g2977) & (g2978)) + ((g1543) & (g2822) & (g820) & (g2824) & (g2977) & (!g2978)) + ((g1543) & (g2822) & (g820) & (g2824) & (g2977) & (g2978)));
	assign g3010 = (((!g2981) & (!sk[57]) & (g3009)) + ((!g2981) & (sk[57]) & (g3009)) + ((g2981) & (!sk[57]) & (g3009)));
	assign g3011 = (((!g1589) & (!g2826) & (!g867) & (g2827) & (g2977) & (!g2978)) + ((!g1589) & (!g2826) & (g867) & (!g2827) & (!g2977) & (!g2978)) + ((!g1589) & (!g2826) & (g867) & (g2827) & (!g2977) & (!g2978)) + ((!g1589) & (!g2826) & (g867) & (g2827) & (g2977) & (!g2978)) + ((!g1589) & (g2826) & (!g867) & (!g2827) & (g2977) & (g2978)) + ((!g1589) & (g2826) & (!g867) & (g2827) & (g2977) & (!g2978)) + ((!g1589) & (g2826) & (!g867) & (g2827) & (g2977) & (g2978)) + ((!g1589) & (g2826) & (g867) & (!g2827) & (!g2977) & (!g2978)) + ((!g1589) & (g2826) & (g867) & (!g2827) & (g2977) & (g2978)) + ((!g1589) & (g2826) & (g867) & (g2827) & (!g2977) & (!g2978)) + ((!g1589) & (g2826) & (g867) & (g2827) & (g2977) & (!g2978)) + ((!g1589) & (g2826) & (g867) & (g2827) & (g2977) & (g2978)) + ((g1589) & (!g2826) & (!g867) & (!g2827) & (!g2977) & (g2978)) + ((g1589) & (!g2826) & (!g867) & (g2827) & (!g2977) & (g2978)) + ((g1589) & (!g2826) & (!g867) & (g2827) & (g2977) & (!g2978)) + ((g1589) & (!g2826) & (g867) & (!g2827) & (!g2977) & (!g2978)) + ((g1589) & (!g2826) & (g867) & (!g2827) & (!g2977) & (g2978)) + ((g1589) & (!g2826) & (g867) & (g2827) & (!g2977) & (!g2978)) + ((g1589) & (!g2826) & (g867) & (g2827) & (!g2977) & (g2978)) + ((g1589) & (!g2826) & (g867) & (g2827) & (g2977) & (!g2978)) + ((g1589) & (g2826) & (!g867) & (!g2827) & (!g2977) & (g2978)) + ((g1589) & (g2826) & (!g867) & (!g2827) & (g2977) & (g2978)) + ((g1589) & (g2826) & (!g867) & (g2827) & (!g2977) & (g2978)) + ((g1589) & (g2826) & (!g867) & (g2827) & (g2977) & (!g2978)) + ((g1589) & (g2826) & (!g867) & (g2827) & (g2977) & (g2978)) + ((g1589) & (g2826) & (g867) & (!g2827) & (!g2977) & (!g2978)) + ((g1589) & (g2826) & (g867) & (!g2827) & (!g2977) & (g2978)) + ((g1589) & (g2826) & (g867) & (!g2827) & (g2977) & (g2978)) + ((g1589) & (g2826) & (g867) & (g2827) & (!g2977) & (!g2978)) + ((g1589) & (g2826) & (g867) & (g2827) & (!g2977) & (g2978)) + ((g1589) & (g2826) & (g867) & (g2827) & (g2977) & (!g2978)) + ((g1589) & (g2826) & (g867) & (g2827) & (g2977) & (g2978)));
	assign g3012 = (((!sk[59]) & (!g2981) & (g3011)) + ((!sk[59]) & (g2981) & (g3011)) + ((sk[59]) & (!g2981) & (g3011)));
	assign g3013 = (((!sk[60]) & (!g2024) & (!g76) & (!g142) & (g209) & (!g229)) + ((!sk[60]) & (!g2024) & (!g76) & (!g142) & (g209) & (g229)) + ((!sk[60]) & (!g2024) & (!g76) & (g142) & (!g209) & (!g229)) + ((!sk[60]) & (!g2024) & (!g76) & (g142) & (!g209) & (g229)) + ((!sk[60]) & (!g2024) & (!g76) & (g142) & (g209) & (!g229)) + ((!sk[60]) & (!g2024) & (!g76) & (g142) & (g209) & (g229)) + ((!sk[60]) & (!g2024) & (g76) & (!g142) & (g209) & (!g229)) + ((!sk[60]) & (!g2024) & (g76) & (!g142) & (g209) & (g229)) + ((!sk[60]) & (!g2024) & (g76) & (g142) & (!g209) & (!g229)) + ((!sk[60]) & (!g2024) & (g76) & (g142) & (!g209) & (g229)) + ((!sk[60]) & (!g2024) & (g76) & (g142) & (g209) & (!g229)) + ((!sk[60]) & (!g2024) & (g76) & (g142) & (g209) & (g229)) + ((!sk[60]) & (g2024) & (!g76) & (!g142) & (!g209) & (!g229)) + ((!sk[60]) & (g2024) & (!g76) & (!g142) & (!g209) & (g229)) + ((!sk[60]) & (g2024) & (!g76) & (!g142) & (g209) & (!g229)) + ((!sk[60]) & (g2024) & (!g76) & (!g142) & (g209) & (g229)) + ((!sk[60]) & (g2024) & (!g76) & (g142) & (!g209) & (!g229)) + ((!sk[60]) & (g2024) & (!g76) & (g142) & (!g209) & (g229)) + ((!sk[60]) & (g2024) & (!g76) & (g142) & (g209) & (!g229)) + ((!sk[60]) & (g2024) & (!g76) & (g142) & (g209) & (g229)) + ((!sk[60]) & (g2024) & (g76) & (!g142) & (!g209) & (!g229)) + ((!sk[60]) & (g2024) & (g76) & (!g142) & (!g209) & (g229)) + ((!sk[60]) & (g2024) & (g76) & (!g142) & (g209) & (!g229)) + ((!sk[60]) & (g2024) & (g76) & (!g142) & (g209) & (g229)) + ((!sk[60]) & (g2024) & (g76) & (g142) & (!g209) & (!g229)) + ((!sk[60]) & (g2024) & (g76) & (g142) & (!g209) & (g229)) + ((!sk[60]) & (g2024) & (g76) & (g142) & (g209) & (!g229)) + ((!sk[60]) & (g2024) & (g76) & (g142) & (g209) & (g229)) + ((sk[60]) & (!g2024) & (!g76) & (!g142) & (!g209) & (g229)) + ((sk[60]) & (!g2024) & (!g76) & (!g142) & (g209) & (g229)) + ((sk[60]) & (!g2024) & (!g76) & (g142) & (g209) & (!g229)) + ((sk[60]) & (!g2024) & (!g76) & (g142) & (g209) & (g229)) + ((sk[60]) & (!g2024) & (g76) & (!g142) & (!g209) & (g229)) + ((sk[60]) & (!g2024) & (g76) & (!g142) & (g209) & (g229)) + ((sk[60]) & (!g2024) & (g76) & (g142) & (g209) & (!g229)) + ((sk[60]) & (!g2024) & (g76) & (g142) & (g209) & (g229)) + ((sk[60]) & (g2024) & (g76) & (!g142) & (!g209) & (!g229)) + ((sk[60]) & (g2024) & (g76) & (!g142) & (!g209) & (g229)) + ((sk[60]) & (g2024) & (g76) & (!g142) & (g209) & (!g229)) + ((sk[60]) & (g2024) & (g76) & (!g142) & (g209) & (g229)) + ((sk[60]) & (g2024) & (g76) & (g142) & (!g209) & (!g229)) + ((sk[60]) & (g2024) & (g76) & (g142) & (!g209) & (g229)) + ((sk[60]) & (g2024) & (g76) & (g142) & (g209) & (!g229)) + ((sk[60]) & (g2024) & (g76) & (g142) & (g209) & (g229)));
	assign g3014 = (((!g2928) & (!sk[61]) & (!g2035) & (!g2952) & (g3013)) + ((!g2928) & (!sk[61]) & (!g2035) & (g2952) & (g3013)) + ((!g2928) & (!sk[61]) & (g2035) & (!g2952) & (!g3013)) + ((!g2928) & (!sk[61]) & (g2035) & (!g2952) & (g3013)) + ((!g2928) & (!sk[61]) & (g2035) & (g2952) & (!g3013)) + ((!g2928) & (!sk[61]) & (g2035) & (g2952) & (g3013)) + ((!g2928) & (sk[61]) & (!g2035) & (g2952) & (g3013)) + ((!g2928) & (sk[61]) & (g2035) & (g2952) & (g3013)) + ((g2928) & (!sk[61]) & (!g2035) & (!g2952) & (!g3013)) + ((g2928) & (!sk[61]) & (!g2035) & (!g2952) & (g3013)) + ((g2928) & (!sk[61]) & (!g2035) & (g2952) & (!g3013)) + ((g2928) & (!sk[61]) & (!g2035) & (g2952) & (g3013)) + ((g2928) & (!sk[61]) & (g2035) & (!g2952) & (!g3013)) + ((g2928) & (!sk[61]) & (g2035) & (!g2952) & (g3013)) + ((g2928) & (!sk[61]) & (g2035) & (g2952) & (!g3013)) + ((g2928) & (!sk[61]) & (g2035) & (g2952) & (g3013)) + ((g2928) & (sk[61]) & (g2035) & (g2952) & (!g3013)) + ((g2928) & (sk[61]) & (g2035) & (g2952) & (g3013)));
	assign g3015 = (((!sk[62]) & (!g142) & (g252) & (!g272)) + ((!sk[62]) & (!g142) & (g252) & (g272)) + ((!sk[62]) & (g142) & (!g252) & (!g272)) + ((!sk[62]) & (g142) & (!g252) & (g272)) + ((!sk[62]) & (g142) & (g252) & (!g272)) + ((!sk[62]) & (g142) & (g252) & (g272)) + ((sk[62]) & (!g142) & (!g252) & (g272)) + ((sk[62]) & (!g142) & (g252) & (g272)) + ((sk[62]) & (g142) & (g252) & (!g272)) + ((sk[62]) & (g142) & (g252) & (g272)));
	assign g3016 = (((!g2928) & (!sk[63]) & (g2024) & (!g2950)) + ((!g2928) & (!sk[63]) & (g2024) & (g2950)) + ((!g2928) & (sk[63]) & (!g2024) & (!g2950)) + ((!g2928) & (sk[63]) & (g2024) & (!g2950)) + ((!g2928) & (sk[63]) & (g2024) & (g2950)) + ((g2928) & (!sk[63]) & (!g2024) & (!g2950)) + ((g2928) & (!sk[63]) & (!g2024) & (g2950)) + ((g2928) & (!sk[63]) & (g2024) & (!g2950)) + ((g2928) & (!sk[63]) & (g2024) & (g2950)));
	assign g3017 = (((!sk[64]) & (!g2920) & (g2923)) + ((!sk[64]) & (g2920) & (g2923)) + ((sk[64]) & (!g2920) & (!g2923)));
	assign g3018 = (((!g2049) & (!g2054) & (sk[65]) & (!g2923)) + ((!g2049) & (g2054) & (!sk[65]) & (!g2923)) + ((!g2049) & (g2054) & (!sk[65]) & (g2923)) + ((!g2049) & (g2054) & (sk[65]) & (!g2923)) + ((g2049) & (!g2054) & (!sk[65]) & (!g2923)) + ((g2049) & (!g2054) & (!sk[65]) & (g2923)) + ((g2049) & (!g2054) & (sk[65]) & (!g2923)) + ((g2049) & (g2054) & (!sk[65]) & (!g2923)) + ((g2049) & (g2054) & (!sk[65]) & (g2923)));
	assign g3019 = (((!g2038) & (!sk[66]) & (!g2330) & (!g2066) & (g3017) & (!g3018)) + ((!g2038) & (!sk[66]) & (!g2330) & (!g2066) & (g3017) & (g3018)) + ((!g2038) & (!sk[66]) & (!g2330) & (g2066) & (!g3017) & (!g3018)) + ((!g2038) & (!sk[66]) & (!g2330) & (g2066) & (!g3017) & (g3018)) + ((!g2038) & (!sk[66]) & (!g2330) & (g2066) & (g3017) & (!g3018)) + ((!g2038) & (!sk[66]) & (!g2330) & (g2066) & (g3017) & (g3018)) + ((!g2038) & (!sk[66]) & (g2330) & (!g2066) & (g3017) & (!g3018)) + ((!g2038) & (!sk[66]) & (g2330) & (!g2066) & (g3017) & (g3018)) + ((!g2038) & (!sk[66]) & (g2330) & (g2066) & (!g3017) & (!g3018)) + ((!g2038) & (!sk[66]) & (g2330) & (g2066) & (!g3017) & (g3018)) + ((!g2038) & (!sk[66]) & (g2330) & (g2066) & (g3017) & (!g3018)) + ((!g2038) & (!sk[66]) & (g2330) & (g2066) & (g3017) & (g3018)) + ((!g2038) & (sk[66]) & (!g2330) & (!g2066) & (g3017) & (!g3018)) + ((!g2038) & (sk[66]) & (!g2330) & (g2066) & (!g3017) & (g3018)) + ((!g2038) & (sk[66]) & (!g2330) & (g2066) & (g3017) & (!g3018)) + ((!g2038) & (sk[66]) & (g2330) & (g2066) & (!g3017) & (g3018)) + ((g2038) & (!sk[66]) & (!g2330) & (!g2066) & (!g3017) & (!g3018)) + ((g2038) & (!sk[66]) & (!g2330) & (!g2066) & (!g3017) & (g3018)) + ((g2038) & (!sk[66]) & (!g2330) & (!g2066) & (g3017) & (!g3018)) + ((g2038) & (!sk[66]) & (!g2330) & (!g2066) & (g3017) & (g3018)) + ((g2038) & (!sk[66]) & (!g2330) & (g2066) & (!g3017) & (!g3018)) + ((g2038) & (!sk[66]) & (!g2330) & (g2066) & (!g3017) & (g3018)) + ((g2038) & (!sk[66]) & (!g2330) & (g2066) & (g3017) & (!g3018)) + ((g2038) & (!sk[66]) & (!g2330) & (g2066) & (g3017) & (g3018)) + ((g2038) & (!sk[66]) & (g2330) & (!g2066) & (!g3017) & (!g3018)) + ((g2038) & (!sk[66]) & (g2330) & (!g2066) & (!g3017) & (g3018)) + ((g2038) & (!sk[66]) & (g2330) & (!g2066) & (g3017) & (!g3018)) + ((g2038) & (!sk[66]) & (g2330) & (!g2066) & (g3017) & (g3018)) + ((g2038) & (!sk[66]) & (g2330) & (g2066) & (!g3017) & (!g3018)) + ((g2038) & (!sk[66]) & (g2330) & (g2066) & (!g3017) & (g3018)) + ((g2038) & (!sk[66]) & (g2330) & (g2066) & (g3017) & (!g3018)) + ((g2038) & (!sk[66]) & (g2330) & (g2066) & (g3017) & (g3018)) + ((g2038) & (sk[66]) & (!g2330) & (!g2066) & (!g3017) & (!g3018)) + ((g2038) & (sk[66]) & (!g2330) & (!g2066) & (g3017) & (!g3018)) + ((g2038) & (sk[66]) & (!g2330) & (g2066) & (!g3017) & (!g3018)) + ((g2038) & (sk[66]) & (!g2330) & (g2066) & (!g3017) & (g3018)) + ((g2038) & (sk[66]) & (!g2330) & (g2066) & (g3017) & (!g3018)) + ((g2038) & (sk[66]) & (g2330) & (!g2066) & (!g3017) & (!g3018)) + ((g2038) & (sk[66]) & (g2330) & (g2066) & (!g3017) & (!g3018)) + ((g2038) & (sk[66]) & (g2330) & (g2066) & (!g3017) & (g3018)));
	assign g3020 = (((!g3015) & (!g141) & (!g2977) & (!sk[67]) & (g3016) & (!g3019)) + ((!g3015) & (!g141) & (!g2977) & (!sk[67]) & (g3016) & (g3019)) + ((!g3015) & (!g141) & (g2977) & (!sk[67]) & (!g3016) & (!g3019)) + ((!g3015) & (!g141) & (g2977) & (!sk[67]) & (!g3016) & (g3019)) + ((!g3015) & (!g141) & (g2977) & (!sk[67]) & (g3016) & (!g3019)) + ((!g3015) & (!g141) & (g2977) & (!sk[67]) & (g3016) & (g3019)) + ((!g3015) & (!g141) & (g2977) & (sk[67]) & (!g3016) & (g3019)) + ((!g3015) & (!g141) & (g2977) & (sk[67]) & (g3016) & (!g3019)) + ((!g3015) & (!g141) & (g2977) & (sk[67]) & (g3016) & (g3019)) + ((!g3015) & (g141) & (!g2977) & (!sk[67]) & (g3016) & (!g3019)) + ((!g3015) & (g141) & (!g2977) & (!sk[67]) & (g3016) & (g3019)) + ((!g3015) & (g141) & (g2977) & (!sk[67]) & (!g3016) & (!g3019)) + ((!g3015) & (g141) & (g2977) & (!sk[67]) & (!g3016) & (g3019)) + ((!g3015) & (g141) & (g2977) & (!sk[67]) & (g3016) & (!g3019)) + ((!g3015) & (g141) & (g2977) & (!sk[67]) & (g3016) & (g3019)) + ((!g3015) & (g141) & (g2977) & (sk[67]) & (!g3016) & (g3019)) + ((g3015) & (!g141) & (!g2977) & (!sk[67]) & (!g3016) & (!g3019)) + ((g3015) & (!g141) & (!g2977) & (!sk[67]) & (!g3016) & (g3019)) + ((g3015) & (!g141) & (!g2977) & (!sk[67]) & (g3016) & (!g3019)) + ((g3015) & (!g141) & (!g2977) & (!sk[67]) & (g3016) & (g3019)) + ((g3015) & (!g141) & (!g2977) & (sk[67]) & (!g3016) & (!g3019)) + ((g3015) & (!g141) & (!g2977) & (sk[67]) & (!g3016) & (g3019)) + ((g3015) & (!g141) & (g2977) & (!sk[67]) & (!g3016) & (!g3019)) + ((g3015) & (!g141) & (g2977) & (!sk[67]) & (!g3016) & (g3019)) + ((g3015) & (!g141) & (g2977) & (!sk[67]) & (g3016) & (!g3019)) + ((g3015) & (!g141) & (g2977) & (!sk[67]) & (g3016) & (g3019)) + ((g3015) & (!g141) & (g2977) & (sk[67]) & (!g3016) & (g3019)) + ((g3015) & (!g141) & (g2977) & (sk[67]) & (g3016) & (!g3019)) + ((g3015) & (!g141) & (g2977) & (sk[67]) & (g3016) & (g3019)) + ((g3015) & (g141) & (!g2977) & (!sk[67]) & (!g3016) & (!g3019)) + ((g3015) & (g141) & (!g2977) & (!sk[67]) & (!g3016) & (g3019)) + ((g3015) & (g141) & (!g2977) & (!sk[67]) & (g3016) & (!g3019)) + ((g3015) & (g141) & (!g2977) & (!sk[67]) & (g3016) & (g3019)) + ((g3015) & (g141) & (!g2977) & (sk[67]) & (!g3016) & (!g3019)) + ((g3015) & (g141) & (!g2977) & (sk[67]) & (!g3016) & (g3019)) + ((g3015) & (g141) & (g2977) & (!sk[67]) & (!g3016) & (!g3019)) + ((g3015) & (g141) & (g2977) & (!sk[67]) & (!g3016) & (g3019)) + ((g3015) & (g141) & (g2977) & (!sk[67]) & (g3016) & (!g3019)) + ((g3015) & (g141) & (g2977) & (!sk[67]) & (g3016) & (g3019)) + ((g3015) & (g141) & (g2977) & (sk[67]) & (!g3016) & (g3019)));
	assign g3021 = (((!g2024) & (!g142) & (!g296) & (!sk[68]) & (g316) & (!g2230)) + ((!g2024) & (!g142) & (!g296) & (!sk[68]) & (g316) & (g2230)) + ((!g2024) & (!g142) & (!g296) & (sk[68]) & (g316) & (!g2230)) + ((!g2024) & (!g142) & (!g296) & (sk[68]) & (g316) & (g2230)) + ((!g2024) & (!g142) & (g296) & (!sk[68]) & (!g316) & (!g2230)) + ((!g2024) & (!g142) & (g296) & (!sk[68]) & (!g316) & (g2230)) + ((!g2024) & (!g142) & (g296) & (!sk[68]) & (g316) & (!g2230)) + ((!g2024) & (!g142) & (g296) & (!sk[68]) & (g316) & (g2230)) + ((!g2024) & (!g142) & (g296) & (sk[68]) & (g316) & (!g2230)) + ((!g2024) & (!g142) & (g296) & (sk[68]) & (g316) & (g2230)) + ((!g2024) & (g142) & (!g296) & (!sk[68]) & (g316) & (!g2230)) + ((!g2024) & (g142) & (!g296) & (!sk[68]) & (g316) & (g2230)) + ((!g2024) & (g142) & (g296) & (!sk[68]) & (!g316) & (!g2230)) + ((!g2024) & (g142) & (g296) & (!sk[68]) & (!g316) & (g2230)) + ((!g2024) & (g142) & (g296) & (!sk[68]) & (g316) & (!g2230)) + ((!g2024) & (g142) & (g296) & (!sk[68]) & (g316) & (g2230)) + ((!g2024) & (g142) & (g296) & (sk[68]) & (!g316) & (!g2230)) + ((!g2024) & (g142) & (g296) & (sk[68]) & (!g316) & (g2230)) + ((!g2024) & (g142) & (g296) & (sk[68]) & (g316) & (!g2230)) + ((!g2024) & (g142) & (g296) & (sk[68]) & (g316) & (g2230)) + ((g2024) & (!g142) & (!g296) & (!sk[68]) & (!g316) & (!g2230)) + ((g2024) & (!g142) & (!g296) & (!sk[68]) & (!g316) & (g2230)) + ((g2024) & (!g142) & (!g296) & (!sk[68]) & (g316) & (!g2230)) + ((g2024) & (!g142) & (!g296) & (!sk[68]) & (g316) & (g2230)) + ((g2024) & (!g142) & (!g296) & (sk[68]) & (!g316) & (g2230)) + ((g2024) & (!g142) & (!g296) & (sk[68]) & (g316) & (g2230)) + ((g2024) & (!g142) & (g296) & (!sk[68]) & (!g316) & (!g2230)) + ((g2024) & (!g142) & (g296) & (!sk[68]) & (!g316) & (g2230)) + ((g2024) & (!g142) & (g296) & (!sk[68]) & (g316) & (!g2230)) + ((g2024) & (!g142) & (g296) & (!sk[68]) & (g316) & (g2230)) + ((g2024) & (!g142) & (g296) & (sk[68]) & (!g316) & (g2230)) + ((g2024) & (!g142) & (g296) & (sk[68]) & (g316) & (g2230)) + ((g2024) & (g142) & (!g296) & (!sk[68]) & (!g316) & (!g2230)) + ((g2024) & (g142) & (!g296) & (!sk[68]) & (!g316) & (g2230)) + ((g2024) & (g142) & (!g296) & (!sk[68]) & (g316) & (!g2230)) + ((g2024) & (g142) & (!g296) & (!sk[68]) & (g316) & (g2230)) + ((g2024) & (g142) & (!g296) & (sk[68]) & (!g316) & (g2230)) + ((g2024) & (g142) & (!g296) & (sk[68]) & (g316) & (g2230)) + ((g2024) & (g142) & (g296) & (!sk[68]) & (!g316) & (!g2230)) + ((g2024) & (g142) & (g296) & (!sk[68]) & (!g316) & (g2230)) + ((g2024) & (g142) & (g296) & (!sk[68]) & (g316) & (!g2230)) + ((g2024) & (g142) & (g296) & (!sk[68]) & (g316) & (g2230)) + ((g2024) & (g142) & (g296) & (sk[68]) & (!g316) & (g2230)) + ((g2024) & (g142) & (g296) & (sk[68]) & (g316) & (g2230)));
	assign g3022 = (((!g2928) & (!sk[69]) & (!g2231) & (!g2952) & (g3021)) + ((!g2928) & (!sk[69]) & (!g2231) & (g2952) & (g3021)) + ((!g2928) & (!sk[69]) & (g2231) & (!g2952) & (!g3021)) + ((!g2928) & (!sk[69]) & (g2231) & (!g2952) & (g3021)) + ((!g2928) & (!sk[69]) & (g2231) & (g2952) & (!g3021)) + ((!g2928) & (!sk[69]) & (g2231) & (g2952) & (g3021)) + ((!g2928) & (sk[69]) & (!g2231) & (g2952) & (g3021)) + ((!g2928) & (sk[69]) & (g2231) & (g2952) & (g3021)) + ((g2928) & (!sk[69]) & (!g2231) & (!g2952) & (!g3021)) + ((g2928) & (!sk[69]) & (!g2231) & (!g2952) & (g3021)) + ((g2928) & (!sk[69]) & (!g2231) & (g2952) & (!g3021)) + ((g2928) & (!sk[69]) & (!g2231) & (g2952) & (g3021)) + ((g2928) & (!sk[69]) & (g2231) & (!g2952) & (!g3021)) + ((g2928) & (!sk[69]) & (g2231) & (!g2952) & (g3021)) + ((g2928) & (!sk[69]) & (g2231) & (g2952) & (!g3021)) + ((g2928) & (!sk[69]) & (g2231) & (g2952) & (g3021)) + ((g2928) & (sk[69]) & (g2231) & (g2952) & (!g3021)) + ((g2928) & (sk[69]) & (g2231) & (g2952) & (g3021)));
	assign g3023 = (((!sk[70]) & (!g2024) & (!g142) & (!g518) & (g538) & (!g2355)) + ((!sk[70]) & (!g2024) & (!g142) & (!g518) & (g538) & (g2355)) + ((!sk[70]) & (!g2024) & (!g142) & (g518) & (!g538) & (!g2355)) + ((!sk[70]) & (!g2024) & (!g142) & (g518) & (!g538) & (g2355)) + ((!sk[70]) & (!g2024) & (!g142) & (g518) & (g538) & (!g2355)) + ((!sk[70]) & (!g2024) & (!g142) & (g518) & (g538) & (g2355)) + ((!sk[70]) & (!g2024) & (g142) & (!g518) & (g538) & (!g2355)) + ((!sk[70]) & (!g2024) & (g142) & (!g518) & (g538) & (g2355)) + ((!sk[70]) & (!g2024) & (g142) & (g518) & (!g538) & (!g2355)) + ((!sk[70]) & (!g2024) & (g142) & (g518) & (!g538) & (g2355)) + ((!sk[70]) & (!g2024) & (g142) & (g518) & (g538) & (!g2355)) + ((!sk[70]) & (!g2024) & (g142) & (g518) & (g538) & (g2355)) + ((!sk[70]) & (g2024) & (!g142) & (!g518) & (!g538) & (!g2355)) + ((!sk[70]) & (g2024) & (!g142) & (!g518) & (!g538) & (g2355)) + ((!sk[70]) & (g2024) & (!g142) & (!g518) & (g538) & (!g2355)) + ((!sk[70]) & (g2024) & (!g142) & (!g518) & (g538) & (g2355)) + ((!sk[70]) & (g2024) & (!g142) & (g518) & (!g538) & (!g2355)) + ((!sk[70]) & (g2024) & (!g142) & (g518) & (!g538) & (g2355)) + ((!sk[70]) & (g2024) & (!g142) & (g518) & (g538) & (!g2355)) + ((!sk[70]) & (g2024) & (!g142) & (g518) & (g538) & (g2355)) + ((!sk[70]) & (g2024) & (g142) & (!g518) & (!g538) & (!g2355)) + ((!sk[70]) & (g2024) & (g142) & (!g518) & (!g538) & (g2355)) + ((!sk[70]) & (g2024) & (g142) & (!g518) & (g538) & (!g2355)) + ((!sk[70]) & (g2024) & (g142) & (!g518) & (g538) & (g2355)) + ((!sk[70]) & (g2024) & (g142) & (g518) & (!g538) & (!g2355)) + ((!sk[70]) & (g2024) & (g142) & (g518) & (!g538) & (g2355)) + ((!sk[70]) & (g2024) & (g142) & (g518) & (g538) & (!g2355)) + ((!sk[70]) & (g2024) & (g142) & (g518) & (g538) & (g2355)) + ((sk[70]) & (!g2024) & (!g142) & (!g518) & (g538) & (!g2355)) + ((sk[70]) & (!g2024) & (!g142) & (!g518) & (g538) & (g2355)) + ((sk[70]) & (!g2024) & (!g142) & (g518) & (g538) & (!g2355)) + ((sk[70]) & (!g2024) & (!g142) & (g518) & (g538) & (g2355)) + ((sk[70]) & (!g2024) & (g142) & (g518) & (!g538) & (!g2355)) + ((sk[70]) & (!g2024) & (g142) & (g518) & (!g538) & (g2355)) + ((sk[70]) & (!g2024) & (g142) & (g518) & (g538) & (!g2355)) + ((sk[70]) & (!g2024) & (g142) & (g518) & (g538) & (g2355)) + ((sk[70]) & (g2024) & (!g142) & (!g518) & (!g538) & (g2355)) + ((sk[70]) & (g2024) & (!g142) & (!g518) & (g538) & (g2355)) + ((sk[70]) & (g2024) & (!g142) & (g518) & (!g538) & (g2355)) + ((sk[70]) & (g2024) & (!g142) & (g518) & (g538) & (g2355)) + ((sk[70]) & (g2024) & (g142) & (!g518) & (!g538) & (g2355)) + ((sk[70]) & (g2024) & (g142) & (!g518) & (g538) & (g2355)) + ((sk[70]) & (g2024) & (g142) & (g518) & (!g538) & (g2355)) + ((sk[70]) & (g2024) & (g142) & (g518) & (g538) & (g2355)));
	assign g3024 = (((!g2928) & (!g2357) & (!sk[71]) & (!g2952) & (g3023)) + ((!g2928) & (!g2357) & (!sk[71]) & (g2952) & (g3023)) + ((!g2928) & (!g2357) & (sk[71]) & (g2952) & (g3023)) + ((!g2928) & (g2357) & (!sk[71]) & (!g2952) & (!g3023)) + ((!g2928) & (g2357) & (!sk[71]) & (!g2952) & (g3023)) + ((!g2928) & (g2357) & (!sk[71]) & (g2952) & (!g3023)) + ((!g2928) & (g2357) & (!sk[71]) & (g2952) & (g3023)) + ((!g2928) & (g2357) & (sk[71]) & (g2952) & (g3023)) + ((g2928) & (!g2357) & (!sk[71]) & (!g2952) & (!g3023)) + ((g2928) & (!g2357) & (!sk[71]) & (!g2952) & (g3023)) + ((g2928) & (!g2357) & (!sk[71]) & (g2952) & (!g3023)) + ((g2928) & (!g2357) & (!sk[71]) & (g2952) & (g3023)) + ((g2928) & (g2357) & (!sk[71]) & (!g2952) & (!g3023)) + ((g2928) & (g2357) & (!sk[71]) & (!g2952) & (g3023)) + ((g2928) & (g2357) & (!sk[71]) & (g2952) & (!g3023)) + ((g2928) & (g2357) & (!sk[71]) & (g2952) & (g3023)) + ((g2928) & (g2357) & (sk[71]) & (g2952) & (!g3023)) + ((g2928) & (g2357) & (sk[71]) & (g2952) & (g3023)));
	assign g3025 = (((!g2977) & (!g3016) & (!g2916) & (!g3017) & (!g2380) & (g3124)) + ((!g2977) & (!g3016) & (!g2916) & (!g3017) & (g2380) & (g3124)) + ((!g2977) & (!g3016) & (!g2916) & (g3017) & (!g2380) & (g3124)) + ((!g2977) & (!g3016) & (!g2916) & (g3017) & (g2380) & (g3124)) + ((!g2977) & (!g3016) & (g2916) & (!g3017) & (!g2380) & (g3124)) + ((!g2977) & (!g3016) & (g2916) & (!g3017) & (g2380) & (g3124)) + ((!g2977) & (!g3016) & (g2916) & (g3017) & (!g2380) & (g3124)) + ((!g2977) & (!g3016) & (g2916) & (g3017) & (g2380) & (g3124)) + ((g2977) & (!g3016) & (!g2916) & (!g3017) & (!g2380) & (g3124)) + ((g2977) & (!g3016) & (!g2916) & (!g3017) & (g2380) & (g3124)) + ((g2977) & (!g3016) & (!g2916) & (g3017) & (!g2380) & (g3124)) + ((g2977) & (!g3016) & (!g2916) & (g3017) & (g2380) & (g3124)) + ((g2977) & (!g3016) & (g2916) & (!g3017) & (!g2380) & (g3124)) + ((g2977) & (!g3016) & (g2916) & (!g3017) & (g2380) & (g3124)) + ((g2977) & (g3016) & (!g2916) & (!g3017) & (g2380) & (!g3124)) + ((g2977) & (g3016) & (!g2916) & (!g3017) & (g2380) & (g3124)) + ((g2977) & (g3016) & (!g2916) & (g3017) & (g2380) & (!g3124)) + ((g2977) & (g3016) & (!g2916) & (g3017) & (g2380) & (g3124)) + ((g2977) & (g3016) & (g2916) & (!g3017) & (g2380) & (!g3124)) + ((g2977) & (g3016) & (g2916) & (!g3017) & (g2380) & (g3124)) + ((g2977) & (g3016) & (g2916) & (g3017) & (g2380) & (!g3124)) + ((g2977) & (g3016) & (g2916) & (g3017) & (g2380) & (g3124)));
	assign g3026 = (((!sk[73]) & (!g142) & (g608) & (!g628)) + ((!sk[73]) & (!g142) & (g608) & (g628)) + ((!sk[73]) & (g142) & (!g608) & (!g628)) + ((!sk[73]) & (g142) & (!g608) & (g628)) + ((!sk[73]) & (g142) & (g608) & (!g628)) + ((!sk[73]) & (g142) & (g608) & (g628)) + ((sk[73]) & (!g142) & (!g608) & (g628)) + ((sk[73]) & (!g142) & (g608) & (g628)) + ((sk[73]) & (g142) & (g608) & (!g628)) + ((sk[73]) & (g142) & (g608) & (g628)));
	assign g3027 = (((!g2413) & (!g3017) & (!g3018) & (!sk[74]) & (g2969)) + ((!g2413) & (!g3017) & (!g3018) & (sk[74]) & (g2969)) + ((!g2413) & (!g3017) & (g3018) & (!sk[74]) & (g2969)) + ((!g2413) & (g3017) & (!g3018) & (!sk[74]) & (!g2969)) + ((!g2413) & (g3017) & (!g3018) & (!sk[74]) & (g2969)) + ((!g2413) & (g3017) & (g3018) & (!sk[74]) & (!g2969)) + ((!g2413) & (g3017) & (g3018) & (!sk[74]) & (g2969)) + ((g2413) & (!g3017) & (!g3018) & (!sk[74]) & (!g2969)) + ((g2413) & (!g3017) & (!g3018) & (!sk[74]) & (g2969)) + ((g2413) & (!g3017) & (!g3018) & (sk[74]) & (g2969)) + ((g2413) & (!g3017) & (g3018) & (!sk[74]) & (!g2969)) + ((g2413) & (!g3017) & (g3018) & (!sk[74]) & (g2969)) + ((g2413) & (!g3017) & (g3018) & (sk[74]) & (!g2969)) + ((g2413) & (!g3017) & (g3018) & (sk[74]) & (g2969)) + ((g2413) & (g3017) & (!g3018) & (!sk[74]) & (!g2969)) + ((g2413) & (g3017) & (!g3018) & (!sk[74]) & (g2969)) + ((g2413) & (g3017) & (g3018) & (!sk[74]) & (!g2969)) + ((g2413) & (g3017) & (g3018) & (!sk[74]) & (g2969)));
	assign g3028 = (((!g3026) & (!sk[75]) & (!g2410) & (!g2977) & (g3016) & (!g3027)) + ((!g3026) & (!sk[75]) & (!g2410) & (!g2977) & (g3016) & (g3027)) + ((!g3026) & (!sk[75]) & (!g2410) & (g2977) & (!g3016) & (!g3027)) + ((!g3026) & (!sk[75]) & (!g2410) & (g2977) & (!g3016) & (g3027)) + ((!g3026) & (!sk[75]) & (!g2410) & (g2977) & (g3016) & (!g3027)) + ((!g3026) & (!sk[75]) & (!g2410) & (g2977) & (g3016) & (g3027)) + ((!g3026) & (!sk[75]) & (g2410) & (!g2977) & (g3016) & (!g3027)) + ((!g3026) & (!sk[75]) & (g2410) & (!g2977) & (g3016) & (g3027)) + ((!g3026) & (!sk[75]) & (g2410) & (g2977) & (!g3016) & (!g3027)) + ((!g3026) & (!sk[75]) & (g2410) & (g2977) & (!g3016) & (g3027)) + ((!g3026) & (!sk[75]) & (g2410) & (g2977) & (g3016) & (!g3027)) + ((!g3026) & (!sk[75]) & (g2410) & (g2977) & (g3016) & (g3027)) + ((!g3026) & (sk[75]) & (!g2410) & (g2977) & (!g3016) & (g3027)) + ((!g3026) & (sk[75]) & (g2410) & (g2977) & (!g3016) & (g3027)) + ((!g3026) & (sk[75]) & (g2410) & (g2977) & (g3016) & (!g3027)) + ((!g3026) & (sk[75]) & (g2410) & (g2977) & (g3016) & (g3027)) + ((g3026) & (!sk[75]) & (!g2410) & (!g2977) & (!g3016) & (!g3027)) + ((g3026) & (!sk[75]) & (!g2410) & (!g2977) & (!g3016) & (g3027)) + ((g3026) & (!sk[75]) & (!g2410) & (!g2977) & (g3016) & (!g3027)) + ((g3026) & (!sk[75]) & (!g2410) & (!g2977) & (g3016) & (g3027)) + ((g3026) & (!sk[75]) & (!g2410) & (g2977) & (!g3016) & (!g3027)) + ((g3026) & (!sk[75]) & (!g2410) & (g2977) & (!g3016) & (g3027)) + ((g3026) & (!sk[75]) & (!g2410) & (g2977) & (g3016) & (!g3027)) + ((g3026) & (!sk[75]) & (!g2410) & (g2977) & (g3016) & (g3027)) + ((g3026) & (!sk[75]) & (g2410) & (!g2977) & (!g3016) & (!g3027)) + ((g3026) & (!sk[75]) & (g2410) & (!g2977) & (!g3016) & (g3027)) + ((g3026) & (!sk[75]) & (g2410) & (!g2977) & (g3016) & (!g3027)) + ((g3026) & (!sk[75]) & (g2410) & (!g2977) & (g3016) & (g3027)) + ((g3026) & (!sk[75]) & (g2410) & (g2977) & (!g3016) & (!g3027)) + ((g3026) & (!sk[75]) & (g2410) & (g2977) & (!g3016) & (g3027)) + ((g3026) & (!sk[75]) & (g2410) & (g2977) & (g3016) & (!g3027)) + ((g3026) & (!sk[75]) & (g2410) & (g2977) & (g3016) & (g3027)) + ((g3026) & (sk[75]) & (!g2410) & (!g2977) & (!g3016) & (!g3027)) + ((g3026) & (sk[75]) & (!g2410) & (!g2977) & (!g3016) & (g3027)) + ((g3026) & (sk[75]) & (!g2410) & (g2977) & (!g3016) & (g3027)) + ((g3026) & (sk[75]) & (g2410) & (!g2977) & (!g3016) & (!g3027)) + ((g3026) & (sk[75]) & (g2410) & (!g2977) & (!g3016) & (g3027)) + ((g3026) & (sk[75]) & (g2410) & (g2977) & (!g3016) & (g3027)) + ((g3026) & (sk[75]) & (g2410) & (g2977) & (g3016) & (!g3027)) + ((g3026) & (sk[75]) & (g2410) & (g2977) & (g3016) & (g3027)));
	assign g3029 = (((!g2977) & (!g3016) & (!g3017) & (!g3018) & (!g2972) & (g3028)) + ((!g2977) & (!g3016) & (!g3017) & (!g3018) & (g2972) & (g3028)) + ((!g2977) & (!g3016) & (!g3017) & (g3018) & (!g2972) & (g3028)) + ((!g2977) & (!g3016) & (!g3017) & (g3018) & (g2972) & (g3028)) + ((!g2977) & (!g3016) & (g3017) & (!g3018) & (!g2972) & (g3028)) + ((!g2977) & (!g3016) & (g3017) & (!g3018) & (g2972) & (g3028)) + ((!g2977) & (!g3016) & (g3017) & (g3018) & (!g2972) & (g3028)) + ((!g2977) & (!g3016) & (g3017) & (g3018) & (g2972) & (g3028)) + ((!g2977) & (g3016) & (!g3017) & (!g3018) & (!g2972) & (g3028)) + ((!g2977) & (g3016) & (!g3017) & (!g3018) & (g2972) & (g3028)) + ((!g2977) & (g3016) & (!g3017) & (g3018) & (!g2972) & (g3028)) + ((!g2977) & (g3016) & (!g3017) & (g3018) & (g2972) & (g3028)) + ((!g2977) & (g3016) & (g3017) & (!g3018) & (!g2972) & (g3028)) + ((!g2977) & (g3016) & (g3017) & (!g3018) & (g2972) & (g3028)) + ((!g2977) & (g3016) & (g3017) & (g3018) & (!g2972) & (g3028)) + ((!g2977) & (g3016) & (g3017) & (g3018) & (g2972) & (g3028)) + ((g2977) & (!g3016) & (!g3017) & (!g3018) & (!g2972) & (g3028)) + ((g2977) & (!g3016) & (!g3017) & (!g3018) & (g2972) & (g3028)) + ((g2977) & (!g3016) & (!g3017) & (g3018) & (!g2972) & (g3028)) + ((g2977) & (!g3016) & (!g3017) & (g3018) & (g2972) & (g3028)) + ((g2977) & (!g3016) & (g3017) & (!g3018) & (!g2972) & (g3028)) + ((g2977) & (!g3016) & (g3017) & (!g3018) & (g2972) & (!g3028)) + ((g2977) & (!g3016) & (g3017) & (!g3018) & (g2972) & (g3028)) + ((g2977) & (!g3016) & (g3017) & (g3018) & (!g2972) & (g3028)) + ((g2977) & (!g3016) & (g3017) & (g3018) & (g2972) & (g3028)) + ((g2977) & (g3016) & (!g3017) & (!g3018) & (!g2972) & (g3028)) + ((g2977) & (g3016) & (!g3017) & (!g3018) & (g2972) & (g3028)) + ((g2977) & (g3016) & (!g3017) & (g3018) & (!g2972) & (g3028)) + ((g2977) & (g3016) & (!g3017) & (g3018) & (g2972) & (g3028)) + ((g2977) & (g3016) & (g3017) & (!g3018) & (!g2972) & (g3028)) + ((g2977) & (g3016) & (g3017) & (!g3018) & (g2972) & (g3028)) + ((g2977) & (g3016) & (g3017) & (g3018) & (!g2972) & (g3028)) + ((g2977) & (g3016) & (g3017) & (g3018) & (g2972) & (g3028)));
	assign g3030 = (((!g2928) & (!g2024) & (g672) & (!g2432) & (!g2436) & (g2952)) + ((!g2928) & (!g2024) & (g672) & (!g2432) & (g2436) & (g2952)) + ((!g2928) & (!g2024) & (g672) & (g2432) & (!g2436) & (g2952)) + ((!g2928) & (!g2024) & (g672) & (g2432) & (g2436) & (g2952)) + ((!g2928) & (g2024) & (!g672) & (!g2432) & (g2436) & (g2952)) + ((!g2928) & (g2024) & (!g672) & (g2432) & (g2436) & (g2952)) + ((!g2928) & (g2024) & (g672) & (!g2432) & (g2436) & (g2952)) + ((!g2928) & (g2024) & (g672) & (g2432) & (g2436) & (g2952)) + ((g2928) & (!g2024) & (!g672) & (g2432) & (!g2436) & (g2952)) + ((g2928) & (!g2024) & (!g672) & (g2432) & (g2436) & (g2952)) + ((g2928) & (!g2024) & (g672) & (g2432) & (!g2436) & (g2952)) + ((g2928) & (!g2024) & (g672) & (g2432) & (g2436) & (g2952)) + ((g2928) & (g2024) & (!g672) & (g2432) & (!g2436) & (g2952)) + ((g2928) & (g2024) & (!g672) & (g2432) & (g2436) & (g2952)) + ((g2928) & (g2024) & (g672) & (g2432) & (!g2436) & (g2952)) + ((g2928) & (g2024) & (g672) & (g2432) & (g2436) & (g2952)));
	assign g3031 = (((!g2024) & (!g142) & (!g341) & (g361) & (!sk[78]) & (!g2257)) + ((!g2024) & (!g142) & (!g341) & (g361) & (!sk[78]) & (g2257)) + ((!g2024) & (!g142) & (!g341) & (g361) & (sk[78]) & (!g2257)) + ((!g2024) & (!g142) & (!g341) & (g361) & (sk[78]) & (g2257)) + ((!g2024) & (!g142) & (g341) & (!g361) & (!sk[78]) & (!g2257)) + ((!g2024) & (!g142) & (g341) & (!g361) & (!sk[78]) & (g2257)) + ((!g2024) & (!g142) & (g341) & (g361) & (!sk[78]) & (!g2257)) + ((!g2024) & (!g142) & (g341) & (g361) & (!sk[78]) & (g2257)) + ((!g2024) & (!g142) & (g341) & (g361) & (sk[78]) & (!g2257)) + ((!g2024) & (!g142) & (g341) & (g361) & (sk[78]) & (g2257)) + ((!g2024) & (g142) & (!g341) & (g361) & (!sk[78]) & (!g2257)) + ((!g2024) & (g142) & (!g341) & (g361) & (!sk[78]) & (g2257)) + ((!g2024) & (g142) & (g341) & (!g361) & (!sk[78]) & (!g2257)) + ((!g2024) & (g142) & (g341) & (!g361) & (!sk[78]) & (g2257)) + ((!g2024) & (g142) & (g341) & (!g361) & (sk[78]) & (!g2257)) + ((!g2024) & (g142) & (g341) & (!g361) & (sk[78]) & (g2257)) + ((!g2024) & (g142) & (g341) & (g361) & (!sk[78]) & (!g2257)) + ((!g2024) & (g142) & (g341) & (g361) & (!sk[78]) & (g2257)) + ((!g2024) & (g142) & (g341) & (g361) & (sk[78]) & (!g2257)) + ((!g2024) & (g142) & (g341) & (g361) & (sk[78]) & (g2257)) + ((g2024) & (!g142) & (!g341) & (!g361) & (!sk[78]) & (!g2257)) + ((g2024) & (!g142) & (!g341) & (!g361) & (!sk[78]) & (g2257)) + ((g2024) & (!g142) & (!g341) & (!g361) & (sk[78]) & (g2257)) + ((g2024) & (!g142) & (!g341) & (g361) & (!sk[78]) & (!g2257)) + ((g2024) & (!g142) & (!g341) & (g361) & (!sk[78]) & (g2257)) + ((g2024) & (!g142) & (!g341) & (g361) & (sk[78]) & (g2257)) + ((g2024) & (!g142) & (g341) & (!g361) & (!sk[78]) & (!g2257)) + ((g2024) & (!g142) & (g341) & (!g361) & (!sk[78]) & (g2257)) + ((g2024) & (!g142) & (g341) & (!g361) & (sk[78]) & (g2257)) + ((g2024) & (!g142) & (g341) & (g361) & (!sk[78]) & (!g2257)) + ((g2024) & (!g142) & (g341) & (g361) & (!sk[78]) & (g2257)) + ((g2024) & (!g142) & (g341) & (g361) & (sk[78]) & (g2257)) + ((g2024) & (g142) & (!g341) & (!g361) & (!sk[78]) & (!g2257)) + ((g2024) & (g142) & (!g341) & (!g361) & (!sk[78]) & (g2257)) + ((g2024) & (g142) & (!g341) & (!g361) & (sk[78]) & (g2257)) + ((g2024) & (g142) & (!g341) & (g361) & (!sk[78]) & (!g2257)) + ((g2024) & (g142) & (!g341) & (g361) & (!sk[78]) & (g2257)) + ((g2024) & (g142) & (!g341) & (g361) & (sk[78]) & (g2257)) + ((g2024) & (g142) & (g341) & (!g361) & (!sk[78]) & (!g2257)) + ((g2024) & (g142) & (g341) & (!g361) & (!sk[78]) & (g2257)) + ((g2024) & (g142) & (g341) & (!g361) & (sk[78]) & (g2257)) + ((g2024) & (g142) & (g341) & (g361) & (!sk[78]) & (!g2257)) + ((g2024) & (g142) & (g341) & (g361) & (!sk[78]) & (g2257)) + ((g2024) & (g142) & (g341) & (g361) & (sk[78]) & (g2257)));
	assign g3032 = (((!sk[79]) & (!g2928) & (!g2258) & (!g2952) & (g3031)) + ((!sk[79]) & (!g2928) & (!g2258) & (g2952) & (g3031)) + ((!sk[79]) & (!g2928) & (g2258) & (!g2952) & (!g3031)) + ((!sk[79]) & (!g2928) & (g2258) & (!g2952) & (g3031)) + ((!sk[79]) & (!g2928) & (g2258) & (g2952) & (!g3031)) + ((!sk[79]) & (!g2928) & (g2258) & (g2952) & (g3031)) + ((!sk[79]) & (g2928) & (!g2258) & (!g2952) & (!g3031)) + ((!sk[79]) & (g2928) & (!g2258) & (!g2952) & (g3031)) + ((!sk[79]) & (g2928) & (!g2258) & (g2952) & (!g3031)) + ((!sk[79]) & (g2928) & (!g2258) & (g2952) & (g3031)) + ((!sk[79]) & (g2928) & (g2258) & (!g2952) & (!g3031)) + ((!sk[79]) & (g2928) & (g2258) & (!g2952) & (g3031)) + ((!sk[79]) & (g2928) & (g2258) & (g2952) & (!g3031)) + ((!sk[79]) & (g2928) & (g2258) & (g2952) & (g3031)) + ((sk[79]) & (!g2928) & (!g2258) & (g2952) & (g3031)) + ((sk[79]) & (!g2928) & (g2258) & (g2952) & (g3031)) + ((sk[79]) & (g2928) & (g2258) & (g2952) & (!g3031)) + ((sk[79]) & (g2928) & (g2258) & (g2952) & (g3031)));
	assign g3033 = (((!sk[80]) & (!g2024) & (!g142) & (!g386) & (g406) & (!g2283)) + ((!sk[80]) & (!g2024) & (!g142) & (!g386) & (g406) & (g2283)) + ((!sk[80]) & (!g2024) & (!g142) & (g386) & (!g406) & (!g2283)) + ((!sk[80]) & (!g2024) & (!g142) & (g386) & (!g406) & (g2283)) + ((!sk[80]) & (!g2024) & (!g142) & (g386) & (g406) & (!g2283)) + ((!sk[80]) & (!g2024) & (!g142) & (g386) & (g406) & (g2283)) + ((!sk[80]) & (!g2024) & (g142) & (!g386) & (g406) & (!g2283)) + ((!sk[80]) & (!g2024) & (g142) & (!g386) & (g406) & (g2283)) + ((!sk[80]) & (!g2024) & (g142) & (g386) & (!g406) & (!g2283)) + ((!sk[80]) & (!g2024) & (g142) & (g386) & (!g406) & (g2283)) + ((!sk[80]) & (!g2024) & (g142) & (g386) & (g406) & (!g2283)) + ((!sk[80]) & (!g2024) & (g142) & (g386) & (g406) & (g2283)) + ((!sk[80]) & (g2024) & (!g142) & (!g386) & (!g406) & (!g2283)) + ((!sk[80]) & (g2024) & (!g142) & (!g386) & (!g406) & (g2283)) + ((!sk[80]) & (g2024) & (!g142) & (!g386) & (g406) & (!g2283)) + ((!sk[80]) & (g2024) & (!g142) & (!g386) & (g406) & (g2283)) + ((!sk[80]) & (g2024) & (!g142) & (g386) & (!g406) & (!g2283)) + ((!sk[80]) & (g2024) & (!g142) & (g386) & (!g406) & (g2283)) + ((!sk[80]) & (g2024) & (!g142) & (g386) & (g406) & (!g2283)) + ((!sk[80]) & (g2024) & (!g142) & (g386) & (g406) & (g2283)) + ((!sk[80]) & (g2024) & (g142) & (!g386) & (!g406) & (!g2283)) + ((!sk[80]) & (g2024) & (g142) & (!g386) & (!g406) & (g2283)) + ((!sk[80]) & (g2024) & (g142) & (!g386) & (g406) & (!g2283)) + ((!sk[80]) & (g2024) & (g142) & (!g386) & (g406) & (g2283)) + ((!sk[80]) & (g2024) & (g142) & (g386) & (!g406) & (!g2283)) + ((!sk[80]) & (g2024) & (g142) & (g386) & (!g406) & (g2283)) + ((!sk[80]) & (g2024) & (g142) & (g386) & (g406) & (!g2283)) + ((!sk[80]) & (g2024) & (g142) & (g386) & (g406) & (g2283)) + ((sk[80]) & (!g2024) & (!g142) & (!g386) & (g406) & (!g2283)) + ((sk[80]) & (!g2024) & (!g142) & (!g386) & (g406) & (g2283)) + ((sk[80]) & (!g2024) & (!g142) & (g386) & (g406) & (!g2283)) + ((sk[80]) & (!g2024) & (!g142) & (g386) & (g406) & (g2283)) + ((sk[80]) & (!g2024) & (g142) & (g386) & (!g406) & (!g2283)) + ((sk[80]) & (!g2024) & (g142) & (g386) & (!g406) & (g2283)) + ((sk[80]) & (!g2024) & (g142) & (g386) & (g406) & (!g2283)) + ((sk[80]) & (!g2024) & (g142) & (g386) & (g406) & (g2283)) + ((sk[80]) & (g2024) & (!g142) & (!g386) & (!g406) & (g2283)) + ((sk[80]) & (g2024) & (!g142) & (!g386) & (g406) & (g2283)) + ((sk[80]) & (g2024) & (!g142) & (g386) & (!g406) & (g2283)) + ((sk[80]) & (g2024) & (!g142) & (g386) & (g406) & (g2283)) + ((sk[80]) & (g2024) & (g142) & (!g386) & (!g406) & (g2283)) + ((sk[80]) & (g2024) & (g142) & (!g386) & (g406) & (g2283)) + ((sk[80]) & (g2024) & (g142) & (g386) & (!g406) & (g2283)) + ((sk[80]) & (g2024) & (g142) & (g386) & (g406) & (g2283)));
	assign g3034 = (((!g2928) & (!g2284) & (!sk[81]) & (!g2952) & (g3033)) + ((!g2928) & (!g2284) & (!sk[81]) & (g2952) & (g3033)) + ((!g2928) & (!g2284) & (sk[81]) & (g2952) & (g3033)) + ((!g2928) & (g2284) & (!sk[81]) & (!g2952) & (!g3033)) + ((!g2928) & (g2284) & (!sk[81]) & (!g2952) & (g3033)) + ((!g2928) & (g2284) & (!sk[81]) & (g2952) & (!g3033)) + ((!g2928) & (g2284) & (!sk[81]) & (g2952) & (g3033)) + ((!g2928) & (g2284) & (sk[81]) & (g2952) & (g3033)) + ((g2928) & (!g2284) & (!sk[81]) & (!g2952) & (!g3033)) + ((g2928) & (!g2284) & (!sk[81]) & (!g2952) & (g3033)) + ((g2928) & (!g2284) & (!sk[81]) & (g2952) & (!g3033)) + ((g2928) & (!g2284) & (!sk[81]) & (g2952) & (g3033)) + ((g2928) & (g2284) & (!sk[81]) & (!g2952) & (!g3033)) + ((g2928) & (g2284) & (!sk[81]) & (!g2952) & (g3033)) + ((g2928) & (g2284) & (!sk[81]) & (g2952) & (!g3033)) + ((g2928) & (g2284) & (!sk[81]) & (g2952) & (g3033)) + ((g2928) & (g2284) & (sk[81]) & (g2952) & (!g3033)) + ((g2928) & (g2284) & (sk[81]) & (g2952) & (g3033)));
	assign g3035 = (((!g2024) & (!g142) & (!g430) & (!sk[82]) & (g450) & (!g2305)) + ((!g2024) & (!g142) & (!g430) & (!sk[82]) & (g450) & (g2305)) + ((!g2024) & (!g142) & (!g430) & (sk[82]) & (g450) & (!g2305)) + ((!g2024) & (!g142) & (!g430) & (sk[82]) & (g450) & (g2305)) + ((!g2024) & (!g142) & (g430) & (!sk[82]) & (!g450) & (!g2305)) + ((!g2024) & (!g142) & (g430) & (!sk[82]) & (!g450) & (g2305)) + ((!g2024) & (!g142) & (g430) & (!sk[82]) & (g450) & (!g2305)) + ((!g2024) & (!g142) & (g430) & (!sk[82]) & (g450) & (g2305)) + ((!g2024) & (!g142) & (g430) & (sk[82]) & (g450) & (!g2305)) + ((!g2024) & (!g142) & (g430) & (sk[82]) & (g450) & (g2305)) + ((!g2024) & (g142) & (!g430) & (!sk[82]) & (g450) & (!g2305)) + ((!g2024) & (g142) & (!g430) & (!sk[82]) & (g450) & (g2305)) + ((!g2024) & (g142) & (g430) & (!sk[82]) & (!g450) & (!g2305)) + ((!g2024) & (g142) & (g430) & (!sk[82]) & (!g450) & (g2305)) + ((!g2024) & (g142) & (g430) & (!sk[82]) & (g450) & (!g2305)) + ((!g2024) & (g142) & (g430) & (!sk[82]) & (g450) & (g2305)) + ((!g2024) & (g142) & (g430) & (sk[82]) & (!g450) & (!g2305)) + ((!g2024) & (g142) & (g430) & (sk[82]) & (!g450) & (g2305)) + ((!g2024) & (g142) & (g430) & (sk[82]) & (g450) & (!g2305)) + ((!g2024) & (g142) & (g430) & (sk[82]) & (g450) & (g2305)) + ((g2024) & (!g142) & (!g430) & (!sk[82]) & (!g450) & (!g2305)) + ((g2024) & (!g142) & (!g430) & (!sk[82]) & (!g450) & (g2305)) + ((g2024) & (!g142) & (!g430) & (!sk[82]) & (g450) & (!g2305)) + ((g2024) & (!g142) & (!g430) & (!sk[82]) & (g450) & (g2305)) + ((g2024) & (!g142) & (!g430) & (sk[82]) & (!g450) & (g2305)) + ((g2024) & (!g142) & (!g430) & (sk[82]) & (g450) & (g2305)) + ((g2024) & (!g142) & (g430) & (!sk[82]) & (!g450) & (!g2305)) + ((g2024) & (!g142) & (g430) & (!sk[82]) & (!g450) & (g2305)) + ((g2024) & (!g142) & (g430) & (!sk[82]) & (g450) & (!g2305)) + ((g2024) & (!g142) & (g430) & (!sk[82]) & (g450) & (g2305)) + ((g2024) & (!g142) & (g430) & (sk[82]) & (!g450) & (g2305)) + ((g2024) & (!g142) & (g430) & (sk[82]) & (g450) & (g2305)) + ((g2024) & (g142) & (!g430) & (!sk[82]) & (!g450) & (!g2305)) + ((g2024) & (g142) & (!g430) & (!sk[82]) & (!g450) & (g2305)) + ((g2024) & (g142) & (!g430) & (!sk[82]) & (g450) & (!g2305)) + ((g2024) & (g142) & (!g430) & (!sk[82]) & (g450) & (g2305)) + ((g2024) & (g142) & (!g430) & (sk[82]) & (!g450) & (g2305)) + ((g2024) & (g142) & (!g430) & (sk[82]) & (g450) & (g2305)) + ((g2024) & (g142) & (g430) & (!sk[82]) & (!g450) & (!g2305)) + ((g2024) & (g142) & (g430) & (!sk[82]) & (!g450) & (g2305)) + ((g2024) & (g142) & (g430) & (!sk[82]) & (g450) & (!g2305)) + ((g2024) & (g142) & (g430) & (!sk[82]) & (g450) & (g2305)) + ((g2024) & (g142) & (g430) & (sk[82]) & (!g450) & (g2305)) + ((g2024) & (g142) & (g430) & (sk[82]) & (g450) & (g2305)));
	assign g3036 = (((!g2928) & (!g2306) & (!g2952) & (!sk[83]) & (g3035)) + ((!g2928) & (!g2306) & (g2952) & (!sk[83]) & (g3035)) + ((!g2928) & (!g2306) & (g2952) & (sk[83]) & (g3035)) + ((!g2928) & (g2306) & (!g2952) & (!sk[83]) & (!g3035)) + ((!g2928) & (g2306) & (!g2952) & (!sk[83]) & (g3035)) + ((!g2928) & (g2306) & (g2952) & (!sk[83]) & (!g3035)) + ((!g2928) & (g2306) & (g2952) & (!sk[83]) & (g3035)) + ((!g2928) & (g2306) & (g2952) & (sk[83]) & (g3035)) + ((g2928) & (!g2306) & (!g2952) & (!sk[83]) & (!g3035)) + ((g2928) & (!g2306) & (!g2952) & (!sk[83]) & (g3035)) + ((g2928) & (!g2306) & (g2952) & (!sk[83]) & (!g3035)) + ((g2928) & (!g2306) & (g2952) & (!sk[83]) & (g3035)) + ((g2928) & (g2306) & (!g2952) & (!sk[83]) & (!g3035)) + ((g2928) & (g2306) & (!g2952) & (!sk[83]) & (g3035)) + ((g2928) & (g2306) & (g2952) & (!sk[83]) & (!g3035)) + ((g2928) & (g2306) & (g2952) & (!sk[83]) & (g3035)) + ((g2928) & (g2306) & (g2952) & (sk[83]) & (!g3035)) + ((g2928) & (g2306) & (g2952) & (sk[83]) & (g3035)));
	assign g3037 = (((!g2024) & (!g142) & (!g474) & (g494) & (!sk[84]) & (!g2332)) + ((!g2024) & (!g142) & (!g474) & (g494) & (!sk[84]) & (g2332)) + ((!g2024) & (!g142) & (!g474) & (g494) & (sk[84]) & (!g2332)) + ((!g2024) & (!g142) & (!g474) & (g494) & (sk[84]) & (g2332)) + ((!g2024) & (!g142) & (g474) & (!g494) & (!sk[84]) & (!g2332)) + ((!g2024) & (!g142) & (g474) & (!g494) & (!sk[84]) & (g2332)) + ((!g2024) & (!g142) & (g474) & (g494) & (!sk[84]) & (!g2332)) + ((!g2024) & (!g142) & (g474) & (g494) & (!sk[84]) & (g2332)) + ((!g2024) & (!g142) & (g474) & (g494) & (sk[84]) & (!g2332)) + ((!g2024) & (!g142) & (g474) & (g494) & (sk[84]) & (g2332)) + ((!g2024) & (g142) & (!g474) & (g494) & (!sk[84]) & (!g2332)) + ((!g2024) & (g142) & (!g474) & (g494) & (!sk[84]) & (g2332)) + ((!g2024) & (g142) & (g474) & (!g494) & (!sk[84]) & (!g2332)) + ((!g2024) & (g142) & (g474) & (!g494) & (!sk[84]) & (g2332)) + ((!g2024) & (g142) & (g474) & (!g494) & (sk[84]) & (!g2332)) + ((!g2024) & (g142) & (g474) & (!g494) & (sk[84]) & (g2332)) + ((!g2024) & (g142) & (g474) & (g494) & (!sk[84]) & (!g2332)) + ((!g2024) & (g142) & (g474) & (g494) & (!sk[84]) & (g2332)) + ((!g2024) & (g142) & (g474) & (g494) & (sk[84]) & (!g2332)) + ((!g2024) & (g142) & (g474) & (g494) & (sk[84]) & (g2332)) + ((g2024) & (!g142) & (!g474) & (!g494) & (!sk[84]) & (!g2332)) + ((g2024) & (!g142) & (!g474) & (!g494) & (!sk[84]) & (g2332)) + ((g2024) & (!g142) & (!g474) & (!g494) & (sk[84]) & (g2332)) + ((g2024) & (!g142) & (!g474) & (g494) & (!sk[84]) & (!g2332)) + ((g2024) & (!g142) & (!g474) & (g494) & (!sk[84]) & (g2332)) + ((g2024) & (!g142) & (!g474) & (g494) & (sk[84]) & (g2332)) + ((g2024) & (!g142) & (g474) & (!g494) & (!sk[84]) & (!g2332)) + ((g2024) & (!g142) & (g474) & (!g494) & (!sk[84]) & (g2332)) + ((g2024) & (!g142) & (g474) & (!g494) & (sk[84]) & (g2332)) + ((g2024) & (!g142) & (g474) & (g494) & (!sk[84]) & (!g2332)) + ((g2024) & (!g142) & (g474) & (g494) & (!sk[84]) & (g2332)) + ((g2024) & (!g142) & (g474) & (g494) & (sk[84]) & (g2332)) + ((g2024) & (g142) & (!g474) & (!g494) & (!sk[84]) & (!g2332)) + ((g2024) & (g142) & (!g474) & (!g494) & (!sk[84]) & (g2332)) + ((g2024) & (g142) & (!g474) & (!g494) & (sk[84]) & (g2332)) + ((g2024) & (g142) & (!g474) & (g494) & (!sk[84]) & (!g2332)) + ((g2024) & (g142) & (!g474) & (g494) & (!sk[84]) & (g2332)) + ((g2024) & (g142) & (!g474) & (g494) & (sk[84]) & (g2332)) + ((g2024) & (g142) & (g474) & (!g494) & (!sk[84]) & (!g2332)) + ((g2024) & (g142) & (g474) & (!g494) & (!sk[84]) & (g2332)) + ((g2024) & (g142) & (g474) & (!g494) & (sk[84]) & (g2332)) + ((g2024) & (g142) & (g474) & (g494) & (!sk[84]) & (!g2332)) + ((g2024) & (g142) & (g474) & (g494) & (!sk[84]) & (g2332)) + ((g2024) & (g142) & (g474) & (g494) & (sk[84]) & (g2332)));
	assign g3038 = (((!sk[85]) & (!g2928) & (!g2333) & (!g2952) & (g3037)) + ((!sk[85]) & (!g2928) & (!g2333) & (g2952) & (g3037)) + ((!sk[85]) & (!g2928) & (g2333) & (!g2952) & (!g3037)) + ((!sk[85]) & (!g2928) & (g2333) & (!g2952) & (g3037)) + ((!sk[85]) & (!g2928) & (g2333) & (g2952) & (!g3037)) + ((!sk[85]) & (!g2928) & (g2333) & (g2952) & (g3037)) + ((!sk[85]) & (g2928) & (!g2333) & (!g2952) & (!g3037)) + ((!sk[85]) & (g2928) & (!g2333) & (!g2952) & (g3037)) + ((!sk[85]) & (g2928) & (!g2333) & (g2952) & (!g3037)) + ((!sk[85]) & (g2928) & (!g2333) & (g2952) & (g3037)) + ((!sk[85]) & (g2928) & (g2333) & (!g2952) & (!g3037)) + ((!sk[85]) & (g2928) & (g2333) & (!g2952) & (g3037)) + ((!sk[85]) & (g2928) & (g2333) & (g2952) & (!g3037)) + ((!sk[85]) & (g2928) & (g2333) & (g2952) & (g3037)) + ((sk[85]) & (!g2928) & (!g2333) & (g2952) & (g3037)) + ((sk[85]) & (!g2928) & (g2333) & (g2952) & (g3037)) + ((sk[85]) & (g2928) & (g2333) & (g2952) & (!g3037)) + ((sk[85]) & (g2928) & (g2333) & (g2952) & (g3037)));
	assign g3039 = (((!g2928) & (!g2024) & (g723) & (!g2474) & (!g2476) & (g2952)) + ((!g2928) & (!g2024) & (g723) & (!g2474) & (g2476) & (g2952)) + ((!g2928) & (!g2024) & (g723) & (g2474) & (!g2476) & (g2952)) + ((!g2928) & (!g2024) & (g723) & (g2474) & (g2476) & (g2952)) + ((!g2928) & (g2024) & (!g723) & (g2474) & (!g2476) & (g2952)) + ((!g2928) & (g2024) & (!g723) & (g2474) & (g2476) & (g2952)) + ((!g2928) & (g2024) & (g723) & (g2474) & (!g2476) & (g2952)) + ((!g2928) & (g2024) & (g723) & (g2474) & (g2476) & (g2952)) + ((g2928) & (!g2024) & (!g723) & (!g2474) & (g2476) & (g2952)) + ((g2928) & (!g2024) & (!g723) & (g2474) & (g2476) & (g2952)) + ((g2928) & (!g2024) & (g723) & (!g2474) & (g2476) & (g2952)) + ((g2928) & (!g2024) & (g723) & (g2474) & (g2476) & (g2952)) + ((g2928) & (g2024) & (!g723) & (!g2474) & (g2476) & (g2952)) + ((g2928) & (g2024) & (!g723) & (g2474) & (g2476) & (g2952)) + ((g2928) & (g2024) & (g723) & (!g2474) & (g2476) & (g2952)) + ((g2928) & (g2024) & (g723) & (g2474) & (g2476) & (g2952)));
	assign g3040 = (((!g2928) & (!g2024) & (g770) & (!g2497) & (!g2499) & (g2952)) + ((!g2928) & (!g2024) & (g770) & (!g2497) & (g2499) & (g2952)) + ((!g2928) & (!g2024) & (g770) & (g2497) & (!g2499) & (g2952)) + ((!g2928) & (!g2024) & (g770) & (g2497) & (g2499) & (g2952)) + ((!g2928) & (g2024) & (!g770) & (g2497) & (!g2499) & (g2952)) + ((!g2928) & (g2024) & (!g770) & (g2497) & (g2499) & (g2952)) + ((!g2928) & (g2024) & (g770) & (g2497) & (!g2499) & (g2952)) + ((!g2928) & (g2024) & (g770) & (g2497) & (g2499) & (g2952)) + ((g2928) & (!g2024) & (!g770) & (!g2497) & (g2499) & (g2952)) + ((g2928) & (!g2024) & (!g770) & (g2497) & (g2499) & (g2952)) + ((g2928) & (!g2024) & (g770) & (!g2497) & (g2499) & (g2952)) + ((g2928) & (!g2024) & (g770) & (g2497) & (g2499) & (g2952)) + ((g2928) & (g2024) & (!g770) & (!g2497) & (g2499) & (g2952)) + ((g2928) & (g2024) & (!g770) & (g2497) & (g2499) & (g2952)) + ((g2928) & (g2024) & (g770) & (!g2497) & (g2499) & (g2952)) + ((g2928) & (g2024) & (g770) & (g2497) & (g2499) & (g2952)));
	assign g3041 = (((!g2928) & (!g2024) & (g817) & (!g2521) & (!g2523) & (g2952)) + ((!g2928) & (!g2024) & (g817) & (!g2521) & (g2523) & (g2952)) + ((!g2928) & (!g2024) & (g817) & (g2521) & (!g2523) & (g2952)) + ((!g2928) & (!g2024) & (g817) & (g2521) & (g2523) & (g2952)) + ((!g2928) & (g2024) & (!g817) & (g2521) & (!g2523) & (g2952)) + ((!g2928) & (g2024) & (!g817) & (g2521) & (g2523) & (g2952)) + ((!g2928) & (g2024) & (g817) & (g2521) & (!g2523) & (g2952)) + ((!g2928) & (g2024) & (g817) & (g2521) & (g2523) & (g2952)) + ((g2928) & (!g2024) & (!g817) & (!g2521) & (g2523) & (g2952)) + ((g2928) & (!g2024) & (!g817) & (g2521) & (g2523) & (g2952)) + ((g2928) & (!g2024) & (g817) & (!g2521) & (g2523) & (g2952)) + ((g2928) & (!g2024) & (g817) & (g2521) & (g2523) & (g2952)) + ((g2928) & (g2024) & (!g817) & (!g2521) & (g2523) & (g2952)) + ((g2928) & (g2024) & (!g817) & (g2521) & (g2523) & (g2952)) + ((g2928) & (g2024) & (g817) & (!g2521) & (g2523) & (g2952)) + ((g2928) & (g2024) & (g817) & (g2521) & (g2523) & (g2952)));
	assign g3042 = (((!g2928) & (!g2024) & (g864) & (!g2543) & (!g2544) & (g2952)) + ((!g2928) & (!g2024) & (g864) & (!g2543) & (g2544) & (g2952)) + ((!g2928) & (!g2024) & (g864) & (g2543) & (!g2544) & (g2952)) + ((!g2928) & (!g2024) & (g864) & (g2543) & (g2544) & (g2952)) + ((!g2928) & (g2024) & (!g864) & (g2543) & (!g2544) & (g2952)) + ((!g2928) & (g2024) & (!g864) & (g2543) & (g2544) & (g2952)) + ((!g2928) & (g2024) & (g864) & (g2543) & (!g2544) & (g2952)) + ((!g2928) & (g2024) & (g864) & (g2543) & (g2544) & (g2952)) + ((g2928) & (!g2024) & (!g864) & (!g2543) & (g2544) & (g2952)) + ((g2928) & (!g2024) & (!g864) & (g2543) & (g2544) & (g2952)) + ((g2928) & (!g2024) & (g864) & (!g2543) & (g2544) & (g2952)) + ((g2928) & (!g2024) & (g864) & (g2543) & (g2544) & (g2952)) + ((g2928) & (g2024) & (!g864) & (!g2543) & (g2544) & (g2952)) + ((g2928) & (g2024) & (!g864) & (g2543) & (g2544) & (g2952)) + ((g2928) & (g2024) & (g864) & (!g2543) & (g2544) & (g2952)) + ((g2928) & (g2024) & (g864) & (g2543) & (g2544) & (g2952)));
	assign g3043 = (((!g84) & (!sk[90]) & (!g87) & (!g88) & (g102)) + ((!g84) & (!sk[90]) & (!g87) & (g88) & (g102)) + ((!g84) & (!sk[90]) & (g87) & (!g88) & (!g102)) + ((!g84) & (!sk[90]) & (g87) & (!g88) & (g102)) + ((!g84) & (!sk[90]) & (g87) & (g88) & (!g102)) + ((!g84) & (!sk[90]) & (g87) & (g88) & (g102)) + ((g84) & (!sk[90]) & (!g87) & (!g88) & (!g102)) + ((g84) & (!sk[90]) & (!g87) & (!g88) & (g102)) + ((g84) & (!sk[90]) & (!g87) & (g88) & (!g102)) + ((g84) & (!sk[90]) & (!g87) & (g88) & (g102)) + ((g84) & (!sk[90]) & (g87) & (!g88) & (!g102)) + ((g84) & (!sk[90]) & (g87) & (!g88) & (g102)) + ((g84) & (!sk[90]) & (g87) & (g88) & (!g102)) + ((g84) & (!sk[90]) & (g87) & (g88) & (g102)) + ((g84) & (sk[90]) & (g87) & (!g88) & (g102)));
	assign g3044 = (((!sk[91]) & (!g106) & (!g2937) & (!g2958) & (g2961) & (!g3043)) + ((!sk[91]) & (!g106) & (!g2937) & (!g2958) & (g2961) & (g3043)) + ((!sk[91]) & (!g106) & (!g2937) & (g2958) & (!g2961) & (!g3043)) + ((!sk[91]) & (!g106) & (!g2937) & (g2958) & (!g2961) & (g3043)) + ((!sk[91]) & (!g106) & (!g2937) & (g2958) & (g2961) & (!g3043)) + ((!sk[91]) & (!g106) & (!g2937) & (g2958) & (g2961) & (g3043)) + ((!sk[91]) & (!g106) & (g2937) & (!g2958) & (g2961) & (!g3043)) + ((!sk[91]) & (!g106) & (g2937) & (!g2958) & (g2961) & (g3043)) + ((!sk[91]) & (!g106) & (g2937) & (g2958) & (!g2961) & (!g3043)) + ((!sk[91]) & (!g106) & (g2937) & (g2958) & (!g2961) & (g3043)) + ((!sk[91]) & (!g106) & (g2937) & (g2958) & (g2961) & (!g3043)) + ((!sk[91]) & (!g106) & (g2937) & (g2958) & (g2961) & (g3043)) + ((!sk[91]) & (g106) & (!g2937) & (!g2958) & (!g2961) & (!g3043)) + ((!sk[91]) & (g106) & (!g2937) & (!g2958) & (!g2961) & (g3043)) + ((!sk[91]) & (g106) & (!g2937) & (!g2958) & (g2961) & (!g3043)) + ((!sk[91]) & (g106) & (!g2937) & (!g2958) & (g2961) & (g3043)) + ((!sk[91]) & (g106) & (!g2937) & (g2958) & (!g2961) & (!g3043)) + ((!sk[91]) & (g106) & (!g2937) & (g2958) & (!g2961) & (g3043)) + ((!sk[91]) & (g106) & (!g2937) & (g2958) & (g2961) & (!g3043)) + ((!sk[91]) & (g106) & (!g2937) & (g2958) & (g2961) & (g3043)) + ((!sk[91]) & (g106) & (g2937) & (!g2958) & (!g2961) & (!g3043)) + ((!sk[91]) & (g106) & (g2937) & (!g2958) & (!g2961) & (g3043)) + ((!sk[91]) & (g106) & (g2937) & (!g2958) & (g2961) & (!g3043)) + ((!sk[91]) & (g106) & (g2937) & (!g2958) & (g2961) & (g3043)) + ((!sk[91]) & (g106) & (g2937) & (g2958) & (!g2961) & (!g3043)) + ((!sk[91]) & (g106) & (g2937) & (g2958) & (!g2961) & (g3043)) + ((!sk[91]) & (g106) & (g2937) & (g2958) & (g2961) & (!g3043)) + ((!sk[91]) & (g106) & (g2937) & (g2958) & (g2961) & (g3043)) + ((sk[91]) & (!g106) & (!g2937) & (!g2958) & (!g2961) & (g3043)) + ((sk[91]) & (!g106) & (!g2937) & (!g2958) & (g2961) & (!g3043)) + ((sk[91]) & (!g106) & (!g2937) & (!g2958) & (g2961) & (g3043)) + ((sk[91]) & (!g106) & (!g2937) & (g2958) & (!g2961) & (!g3043)) + ((sk[91]) & (!g106) & (!g2937) & (g2958) & (!g2961) & (g3043)) + ((sk[91]) & (!g106) & (!g2937) & (g2958) & (g2961) & (!g3043)) + ((sk[91]) & (!g106) & (!g2937) & (g2958) & (g2961) & (g3043)) + ((sk[91]) & (!g106) & (g2937) & (!g2958) & (!g2961) & (g3043)) + ((sk[91]) & (!g106) & (g2937) & (!g2958) & (g2961) & (!g3043)) + ((sk[91]) & (!g106) & (g2937) & (!g2958) & (g2961) & (g3043)) + ((sk[91]) & (!g106) & (g2937) & (g2958) & (!g2961) & (!g3043)) + ((sk[91]) & (!g106) & (g2937) & (g2958) & (!g2961) & (g3043)) + ((sk[91]) & (!g106) & (g2937) & (g2958) & (g2961) & (!g3043)) + ((sk[91]) & (!g106) & (g2937) & (g2958) & (g2961) & (g3043)) + ((sk[91]) & (g106) & (!g2937) & (!g2958) & (!g2961) & (g3043)) + ((sk[91]) & (g106) & (!g2937) & (!g2958) & (g2961) & (!g3043)) + ((sk[91]) & (g106) & (!g2937) & (!g2958) & (g2961) & (g3043)) + ((sk[91]) & (g106) & (!g2937) & (g2958) & (!g2961) & (!g3043)) + ((sk[91]) & (g106) & (!g2937) & (g2958) & (!g2961) & (g3043)) + ((sk[91]) & (g106) & (!g2937) & (g2958) & (g2961) & (!g3043)) + ((sk[91]) & (g106) & (!g2937) & (g2958) & (g2961) & (g3043)) + ((sk[91]) & (g106) & (g2937) & (!g2958) & (!g2961) & (!g3043)) + ((sk[91]) & (g106) & (g2937) & (!g2958) & (!g2961) & (g3043)) + ((sk[91]) & (g106) & (g2937) & (!g2958) & (g2961) & (!g3043)) + ((sk[91]) & (g106) & (g2937) & (!g2958) & (g2961) & (g3043)) + ((sk[91]) & (g106) & (g2937) & (g2958) & (!g2961) & (!g3043)) + ((sk[91]) & (g106) & (g2937) & (g2958) & (!g2961) & (g3043)) + ((sk[91]) & (g106) & (g2937) & (g2958) & (g2961) & (!g3043)) + ((sk[91]) & (g106) & (g2937) & (g2958) & (g2961) & (g3043)));
	assign g3045 = (((!g113) & (!sk[92]) & (g3139)) + ((g113) & (!sk[92]) & (g3139)) + ((g113) & (sk[92]) & (g3139)));
	assign g3046 = (((!g118) & (!sk[93]) & (!g96) & (!g94) & (g2956) & (!g2957)) + ((!g118) & (!sk[93]) & (!g96) & (!g94) & (g2956) & (g2957)) + ((!g118) & (!sk[93]) & (!g96) & (g94) & (!g2956) & (!g2957)) + ((!g118) & (!sk[93]) & (!g96) & (g94) & (!g2956) & (g2957)) + ((!g118) & (!sk[93]) & (!g96) & (g94) & (g2956) & (!g2957)) + ((!g118) & (!sk[93]) & (!g96) & (g94) & (g2956) & (g2957)) + ((!g118) & (!sk[93]) & (g96) & (!g94) & (g2956) & (!g2957)) + ((!g118) & (!sk[93]) & (g96) & (!g94) & (g2956) & (g2957)) + ((!g118) & (!sk[93]) & (g96) & (g94) & (!g2956) & (!g2957)) + ((!g118) & (!sk[93]) & (g96) & (g94) & (!g2956) & (g2957)) + ((!g118) & (!sk[93]) & (g96) & (g94) & (g2956) & (!g2957)) + ((!g118) & (!sk[93]) & (g96) & (g94) & (g2956) & (g2957)) + ((!g118) & (sk[93]) & (!g96) & (!g94) & (!g2956) & (!g2957)) + ((!g118) & (sk[93]) & (!g96) & (!g94) & (!g2956) & (g2957)) + ((!g118) & (sk[93]) & (g96) & (!g94) & (!g2956) & (!g2957)) + ((!g118) & (sk[93]) & (g96) & (!g94) & (!g2956) & (g2957)) + ((g118) & (!sk[93]) & (!g96) & (!g94) & (!g2956) & (!g2957)) + ((g118) & (!sk[93]) & (!g96) & (!g94) & (!g2956) & (g2957)) + ((g118) & (!sk[93]) & (!g96) & (!g94) & (g2956) & (!g2957)) + ((g118) & (!sk[93]) & (!g96) & (!g94) & (g2956) & (g2957)) + ((g118) & (!sk[93]) & (!g96) & (g94) & (!g2956) & (!g2957)) + ((g118) & (!sk[93]) & (!g96) & (g94) & (!g2956) & (g2957)) + ((g118) & (!sk[93]) & (!g96) & (g94) & (g2956) & (!g2957)) + ((g118) & (!sk[93]) & (!g96) & (g94) & (g2956) & (g2957)) + ((g118) & (!sk[93]) & (g96) & (!g94) & (!g2956) & (!g2957)) + ((g118) & (!sk[93]) & (g96) & (!g94) & (!g2956) & (g2957)) + ((g118) & (!sk[93]) & (g96) & (!g94) & (g2956) & (!g2957)) + ((g118) & (!sk[93]) & (g96) & (!g94) & (g2956) & (g2957)) + ((g118) & (!sk[93]) & (g96) & (g94) & (!g2956) & (!g2957)) + ((g118) & (!sk[93]) & (g96) & (g94) & (!g2956) & (g2957)) + ((g118) & (!sk[93]) & (g96) & (g94) & (g2956) & (!g2957)) + ((g118) & (!sk[93]) & (g96) & (g94) & (g2956) & (g2957)) + ((g118) & (sk[93]) & (!g96) & (!g94) & (!g2956) & (!g2957)) + ((g118) & (sk[93]) & (!g96) & (!g94) & (!g2956) & (g2957)) + ((g118) & (sk[93]) & (g96) & (!g94) & (!g2956) & (!g2957)));
	assign g3047 = (((!g106) & (!g100) & (!g2937) & (!g3045) & (sk[94]) & (!g3046)) + ((!g106) & (!g100) & (!g2937) & (!g3045) & (sk[94]) & (g3046)) + ((!g106) & (!g100) & (!g2937) & (g3045) & (!sk[94]) & (!g3046)) + ((!g106) & (!g100) & (!g2937) & (g3045) & (!sk[94]) & (g3046)) + ((!g106) & (!g100) & (!g2937) & (g3045) & (sk[94]) & (!g3046)) + ((!g106) & (!g100) & (!g2937) & (g3045) & (sk[94]) & (g3046)) + ((!g106) & (!g100) & (g2937) & (!g3045) & (!sk[94]) & (!g3046)) + ((!g106) & (!g100) & (g2937) & (!g3045) & (!sk[94]) & (g3046)) + ((!g106) & (!g100) & (g2937) & (!g3045) & (sk[94]) & (!g3046)) + ((!g106) & (!g100) & (g2937) & (!g3045) & (sk[94]) & (g3046)) + ((!g106) & (!g100) & (g2937) & (g3045) & (!sk[94]) & (!g3046)) + ((!g106) & (!g100) & (g2937) & (g3045) & (!sk[94]) & (g3046)) + ((!g106) & (!g100) & (g2937) & (g3045) & (sk[94]) & (!g3046)) + ((!g106) & (!g100) & (g2937) & (g3045) & (sk[94]) & (g3046)) + ((!g106) & (g100) & (!g2937) & (!g3045) & (sk[94]) & (!g3046)) + ((!g106) & (g100) & (!g2937) & (g3045) & (!sk[94]) & (!g3046)) + ((!g106) & (g100) & (!g2937) & (g3045) & (!sk[94]) & (g3046)) + ((!g106) & (g100) & (!g2937) & (g3045) & (sk[94]) & (!g3046)) + ((!g106) & (g100) & (!g2937) & (g3045) & (sk[94]) & (g3046)) + ((!g106) & (g100) & (g2937) & (!g3045) & (!sk[94]) & (!g3046)) + ((!g106) & (g100) & (g2937) & (!g3045) & (!sk[94]) & (g3046)) + ((!g106) & (g100) & (g2937) & (!g3045) & (sk[94]) & (!g3046)) + ((!g106) & (g100) & (g2937) & (g3045) & (!sk[94]) & (!g3046)) + ((!g106) & (g100) & (g2937) & (g3045) & (!sk[94]) & (g3046)) + ((!g106) & (g100) & (g2937) & (g3045) & (sk[94]) & (!g3046)) + ((!g106) & (g100) & (g2937) & (g3045) & (sk[94]) & (g3046)) + ((g106) & (!g100) & (!g2937) & (!g3045) & (!sk[94]) & (!g3046)) + ((g106) & (!g100) & (!g2937) & (!g3045) & (!sk[94]) & (g3046)) + ((g106) & (!g100) & (!g2937) & (!g3045) & (sk[94]) & (!g3046)) + ((g106) & (!g100) & (!g2937) & (!g3045) & (sk[94]) & (g3046)) + ((g106) & (!g100) & (!g2937) & (g3045) & (!sk[94]) & (!g3046)) + ((g106) & (!g100) & (!g2937) & (g3045) & (!sk[94]) & (g3046)) + ((g106) & (!g100) & (!g2937) & (g3045) & (sk[94]) & (!g3046)) + ((g106) & (!g100) & (!g2937) & (g3045) & (sk[94]) & (g3046)) + ((g106) & (!g100) & (g2937) & (!g3045) & (!sk[94]) & (!g3046)) + ((g106) & (!g100) & (g2937) & (!g3045) & (!sk[94]) & (g3046)) + ((g106) & (!g100) & (g2937) & (!g3045) & (sk[94]) & (!g3046)) + ((g106) & (!g100) & (g2937) & (!g3045) & (sk[94]) & (g3046)) + ((g106) & (!g100) & (g2937) & (g3045) & (!sk[94]) & (!g3046)) + ((g106) & (!g100) & (g2937) & (g3045) & (!sk[94]) & (g3046)) + ((g106) & (!g100) & (g2937) & (g3045) & (sk[94]) & (!g3046)) + ((g106) & (!g100) & (g2937) & (g3045) & (sk[94]) & (g3046)) + ((g106) & (g100) & (!g2937) & (!g3045) & (!sk[94]) & (!g3046)) + ((g106) & (g100) & (!g2937) & (!g3045) & (!sk[94]) & (g3046)) + ((g106) & (g100) & (!g2937) & (!g3045) & (sk[94]) & (!g3046)) + ((g106) & (g100) & (!g2937) & (g3045) & (!sk[94]) & (!g3046)) + ((g106) & (g100) & (!g2937) & (g3045) & (!sk[94]) & (g3046)) + ((g106) & (g100) & (!g2937) & (g3045) & (sk[94]) & (!g3046)) + ((g106) & (g100) & (!g2937) & (g3045) & (sk[94]) & (g3046)) + ((g106) & (g100) & (g2937) & (!g3045) & (!sk[94]) & (!g3046)) + ((g106) & (g100) & (g2937) & (!g3045) & (!sk[94]) & (g3046)) + ((g106) & (g100) & (g2937) & (!g3045) & (sk[94]) & (!g3046)) + ((g106) & (g100) & (g2937) & (!g3045) & (sk[94]) & (g3046)) + ((g106) & (g100) & (g2937) & (g3045) & (!sk[94]) & (!g3046)) + ((g106) & (g100) & (g2937) & (g3045) & (!sk[94]) & (g3046)) + ((g106) & (g100) & (g2937) & (g3045) & (sk[94]) & (!g3046)) + ((g106) & (g100) & (g2937) & (g3045) & (sk[94]) & (g3046)));
	assign g3048 = (((!sk[95]) & (!g2024) & (g104) & (!g3045)) + ((!sk[95]) & (!g2024) & (g104) & (g3045)) + ((!sk[95]) & (g2024) & (!g104) & (!g3045)) + ((!sk[95]) & (g2024) & (!g104) & (g3045)) + ((!sk[95]) & (g2024) & (g104) & (!g3045)) + ((!sk[95]) & (g2024) & (g104) & (g3045)) + ((sk[95]) & (!g2024) & (g104) & (!g3045)));
	assign g3049 = (((!g2928) & (!g2920) & (g2949) & (g2962) & (!g3018) & (g3048)) + ((!g2928) & (!g2920) & (g2949) & (g2962) & (g3018) & (g3048)) + ((!g2928) & (g2920) & (g2949) & (g2962) & (!g3018) & (g3048)) + ((!g2928) & (g2920) & (g2949) & (g2962) & (g3018) & (g3048)) + ((g2928) & (!g2920) & (g2949) & (g2962) & (g3018) & (g3048)));
	assign g3050 = (((!sk[97]) & (!g2024) & (g3049)) + ((!sk[97]) & (g2024) & (g3049)) + ((sk[97]) & (!g2024) & (!g3049)));
	assign g3051 = (((!g109) & (!sk[98]) & (g3050)) + ((g109) & (!sk[98]) & (g3050)) + ((g109) & (sk[98]) & (g3050)));
	assign g3052 = (((!g2024) & (!sk[99]) & (g678) & (!g3049)) + ((!g2024) & (!sk[99]) & (g678) & (g3049)) + ((!g2024) & (sk[99]) & (g678) & (!g3049)) + ((g2024) & (!sk[99]) & (!g678) & (!g3049)) + ((g2024) & (!sk[99]) & (!g678) & (g3049)) + ((g2024) & (!sk[99]) & (g678) & (!g3049)) + ((g2024) & (!sk[99]) & (g678) & (g3049)) + ((g2024) & (sk[99]) & (!g678) & (!g3049)) + ((g2024) & (sk[99]) & (!g678) & (g3049)) + ((g2024) & (sk[99]) & (g678) & (!g3049)) + ((g2024) & (sk[99]) & (g678) & (g3049)));
	assign g3053 = (((!g108) & (!sk[100]) & (g3050)) + ((g108) & (!sk[100]) & (g3050)) + ((g108) & (sk[100]) & (g3050)));
	assign g3054 = (((!sk[101]) & (!g107) & (g3050)) + ((!sk[101]) & (g107) & (g3050)) + ((sk[101]) & (g107) & (g3050)));
	assign g3055 = (((!sk[102]) & (!g110) & (g2024) & (!g3049)) + ((!sk[102]) & (!g110) & (g2024) & (g3049)) + ((!sk[102]) & (g110) & (!g2024) & (!g3049)) + ((!sk[102]) & (g110) & (!g2024) & (g3049)) + ((!sk[102]) & (g110) & (g2024) & (!g3049)) + ((!sk[102]) & (g110) & (g2024) & (g3049)) + ((sk[102]) & (!g110) & (g2024) & (!g3049)) + ((sk[102]) & (!g110) & (g2024) & (g3049)) + ((sk[102]) & (g110) & (!g2024) & (!g3049)) + ((sk[102]) & (g110) & (g2024) & (!g3049)) + ((sk[102]) & (g110) & (g2024) & (g3049)));
	assign g3056 = (((!g1644) & (!g2028) & (g2230) & (!g2233) & (!g2356) & (!g2843)) + ((!g1644) & (!g2028) & (g2230) & (!g2233) & (!g2356) & (g2843)) + ((!g1644) & (!g2028) & (g2230) & (!g2233) & (g2356) & (!g2843)) + ((!g1644) & (!g2028) & (g2230) & (g2233) & (!g2356) & (!g2843)) + ((!g1644) & (!g2028) & (g2230) & (g2233) & (!g2356) & (g2843)) + ((!g1644) & (!g2028) & (g2230) & (g2233) & (g2356) & (!g2843)) + ((!g1644) & (g2028) & (!g2230) & (g2233) & (!g2356) & (g2843)) + ((!g1644) & (g2028) & (g2230) & (!g2233) & (!g2356) & (!g2843)) + ((!g1644) & (g2028) & (g2230) & (!g2233) & (g2356) & (!g2843)) + ((!g1644) & (g2028) & (g2230) & (g2233) & (!g2356) & (!g2843)) + ((!g1644) & (g2028) & (g2230) & (g2233) & (!g2356) & (g2843)) + ((!g1644) & (g2028) & (g2230) & (g2233) & (g2356) & (!g2843)) + ((g1644) & (!g2028) & (!g2230) & (!g2233) & (g2356) & (g2843)) + ((g1644) & (!g2028) & (!g2230) & (g2233) & (g2356) & (g2843)) + ((g1644) & (!g2028) & (g2230) & (!g2233) & (!g2356) & (!g2843)) + ((g1644) & (!g2028) & (g2230) & (!g2233) & (!g2356) & (g2843)) + ((g1644) & (!g2028) & (g2230) & (!g2233) & (g2356) & (!g2843)) + ((g1644) & (!g2028) & (g2230) & (!g2233) & (g2356) & (g2843)) + ((g1644) & (!g2028) & (g2230) & (g2233) & (!g2356) & (!g2843)) + ((g1644) & (!g2028) & (g2230) & (g2233) & (!g2356) & (g2843)) + ((g1644) & (!g2028) & (g2230) & (g2233) & (g2356) & (!g2843)) + ((g1644) & (!g2028) & (g2230) & (g2233) & (g2356) & (g2843)) + ((g1644) & (g2028) & (!g2230) & (!g2233) & (g2356) & (g2843)) + ((g1644) & (g2028) & (!g2230) & (g2233) & (!g2356) & (g2843)) + ((g1644) & (g2028) & (!g2230) & (g2233) & (g2356) & (g2843)) + ((g1644) & (g2028) & (g2230) & (!g2233) & (!g2356) & (!g2843)) + ((g1644) & (g2028) & (g2230) & (!g2233) & (g2356) & (!g2843)) + ((g1644) & (g2028) & (g2230) & (!g2233) & (g2356) & (g2843)) + ((g1644) & (g2028) & (g2230) & (g2233) & (!g2356) & (!g2843)) + ((g1644) & (g2028) & (g2230) & (g2233) & (!g2356) & (g2843)) + ((g1644) & (g2028) & (g2230) & (g2233) & (g2356) & (!g2843)) + ((g1644) & (g2028) & (g2230) & (g2233) & (g2356) & (g2843)));
	assign g3057 = (((!g1656) & (!g2028) & (g2257) & (!g2261) & (!g2356) & (!g2843)) + ((!g1656) & (!g2028) & (g2257) & (!g2261) & (!g2356) & (g2843)) + ((!g1656) & (!g2028) & (g2257) & (!g2261) & (g2356) & (!g2843)) + ((!g1656) & (!g2028) & (g2257) & (g2261) & (!g2356) & (!g2843)) + ((!g1656) & (!g2028) & (g2257) & (g2261) & (!g2356) & (g2843)) + ((!g1656) & (!g2028) & (g2257) & (g2261) & (g2356) & (!g2843)) + ((!g1656) & (g2028) & (!g2257) & (g2261) & (!g2356) & (g2843)) + ((!g1656) & (g2028) & (g2257) & (!g2261) & (!g2356) & (!g2843)) + ((!g1656) & (g2028) & (g2257) & (!g2261) & (g2356) & (!g2843)) + ((!g1656) & (g2028) & (g2257) & (g2261) & (!g2356) & (!g2843)) + ((!g1656) & (g2028) & (g2257) & (g2261) & (!g2356) & (g2843)) + ((!g1656) & (g2028) & (g2257) & (g2261) & (g2356) & (!g2843)) + ((g1656) & (!g2028) & (!g2257) & (!g2261) & (g2356) & (g2843)) + ((g1656) & (!g2028) & (!g2257) & (g2261) & (g2356) & (g2843)) + ((g1656) & (!g2028) & (g2257) & (!g2261) & (!g2356) & (!g2843)) + ((g1656) & (!g2028) & (g2257) & (!g2261) & (!g2356) & (g2843)) + ((g1656) & (!g2028) & (g2257) & (!g2261) & (g2356) & (!g2843)) + ((g1656) & (!g2028) & (g2257) & (!g2261) & (g2356) & (g2843)) + ((g1656) & (!g2028) & (g2257) & (g2261) & (!g2356) & (!g2843)) + ((g1656) & (!g2028) & (g2257) & (g2261) & (!g2356) & (g2843)) + ((g1656) & (!g2028) & (g2257) & (g2261) & (g2356) & (!g2843)) + ((g1656) & (!g2028) & (g2257) & (g2261) & (g2356) & (g2843)) + ((g1656) & (g2028) & (!g2257) & (!g2261) & (g2356) & (g2843)) + ((g1656) & (g2028) & (!g2257) & (g2261) & (!g2356) & (g2843)) + ((g1656) & (g2028) & (!g2257) & (g2261) & (g2356) & (g2843)) + ((g1656) & (g2028) & (g2257) & (!g2261) & (!g2356) & (!g2843)) + ((g1656) & (g2028) & (g2257) & (!g2261) & (g2356) & (!g2843)) + ((g1656) & (g2028) & (g2257) & (!g2261) & (g2356) & (g2843)) + ((g1656) & (g2028) & (g2257) & (g2261) & (!g2356) & (!g2843)) + ((g1656) & (g2028) & (g2257) & (g2261) & (!g2356) & (g2843)) + ((g1656) & (g2028) & (g2257) & (g2261) & (g2356) & (!g2843)) + ((g1656) & (g2028) & (g2257) & (g2261) & (g2356) & (g2843)));
	assign g3058 = (((!g1668) & (!g2028) & (g2283) & (!g2286) & (!g2356) & (!g2843)) + ((!g1668) & (!g2028) & (g2283) & (!g2286) & (!g2356) & (g2843)) + ((!g1668) & (!g2028) & (g2283) & (!g2286) & (g2356) & (!g2843)) + ((!g1668) & (!g2028) & (g2283) & (g2286) & (!g2356) & (!g2843)) + ((!g1668) & (!g2028) & (g2283) & (g2286) & (!g2356) & (g2843)) + ((!g1668) & (!g2028) & (g2283) & (g2286) & (g2356) & (!g2843)) + ((!g1668) & (g2028) & (!g2283) & (g2286) & (!g2356) & (g2843)) + ((!g1668) & (g2028) & (g2283) & (!g2286) & (!g2356) & (!g2843)) + ((!g1668) & (g2028) & (g2283) & (!g2286) & (g2356) & (!g2843)) + ((!g1668) & (g2028) & (g2283) & (g2286) & (!g2356) & (!g2843)) + ((!g1668) & (g2028) & (g2283) & (g2286) & (!g2356) & (g2843)) + ((!g1668) & (g2028) & (g2283) & (g2286) & (g2356) & (!g2843)) + ((g1668) & (!g2028) & (!g2283) & (!g2286) & (g2356) & (g2843)) + ((g1668) & (!g2028) & (!g2283) & (g2286) & (g2356) & (g2843)) + ((g1668) & (!g2028) & (g2283) & (!g2286) & (!g2356) & (!g2843)) + ((g1668) & (!g2028) & (g2283) & (!g2286) & (!g2356) & (g2843)) + ((g1668) & (!g2028) & (g2283) & (!g2286) & (g2356) & (!g2843)) + ((g1668) & (!g2028) & (g2283) & (!g2286) & (g2356) & (g2843)) + ((g1668) & (!g2028) & (g2283) & (g2286) & (!g2356) & (!g2843)) + ((g1668) & (!g2028) & (g2283) & (g2286) & (!g2356) & (g2843)) + ((g1668) & (!g2028) & (g2283) & (g2286) & (g2356) & (!g2843)) + ((g1668) & (!g2028) & (g2283) & (g2286) & (g2356) & (g2843)) + ((g1668) & (g2028) & (!g2283) & (!g2286) & (g2356) & (g2843)) + ((g1668) & (g2028) & (!g2283) & (g2286) & (!g2356) & (g2843)) + ((g1668) & (g2028) & (!g2283) & (g2286) & (g2356) & (g2843)) + ((g1668) & (g2028) & (g2283) & (!g2286) & (!g2356) & (!g2843)) + ((g1668) & (g2028) & (g2283) & (!g2286) & (g2356) & (!g2843)) + ((g1668) & (g2028) & (g2283) & (!g2286) & (g2356) & (g2843)) + ((g1668) & (g2028) & (g2283) & (g2286) & (!g2356) & (!g2843)) + ((g1668) & (g2028) & (g2283) & (g2286) & (!g2356) & (g2843)) + ((g1668) & (g2028) & (g2283) & (g2286) & (g2356) & (!g2843)) + ((g1668) & (g2028) & (g2283) & (g2286) & (g2356) & (g2843)));
	assign g3059 = (((!g1668) & (!g364) & (!g2954) & (!sk[106]) & (g2963)) + ((!g1668) & (!g364) & (g2954) & (!sk[106]) & (g2963)) + ((!g1668) & (g364) & (!g2954) & (!sk[106]) & (!g2963)) + ((!g1668) & (g364) & (!g2954) & (!sk[106]) & (g2963)) + ((!g1668) & (g364) & (g2954) & (!sk[106]) & (!g2963)) + ((!g1668) & (g364) & (g2954) & (!sk[106]) & (g2963)) + ((!g1668) & (g364) & (g2954) & (sk[106]) & (!g2963)) + ((g1668) & (!g364) & (!g2954) & (!sk[106]) & (!g2963)) + ((g1668) & (!g364) & (!g2954) & (!sk[106]) & (g2963)) + ((g1668) & (!g364) & (g2954) & (!sk[106]) & (!g2963)) + ((g1668) & (!g364) & (g2954) & (!sk[106]) & (g2963)) + ((g1668) & (!g364) & (g2954) & (sk[106]) & (g2963)) + ((g1668) & (g364) & (!g2954) & (!sk[106]) & (!g2963)) + ((g1668) & (g364) & (!g2954) & (!sk[106]) & (g2963)) + ((g1668) & (g364) & (g2954) & (!sk[106]) & (!g2963)) + ((g1668) & (g364) & (g2954) & (!sk[106]) & (g2963)) + ((g1668) & (g364) & (g2954) & (sk[106]) & (!g2963)) + ((g1668) & (g364) & (g2954) & (sk[106]) & (g2963)));
	assign g3060 = (((!g1680) & (!g2028) & (g2305) & (!g2309) & (!g2356) & (!g2843)) + ((!g1680) & (!g2028) & (g2305) & (!g2309) & (!g2356) & (g2843)) + ((!g1680) & (!g2028) & (g2305) & (!g2309) & (g2356) & (!g2843)) + ((!g1680) & (!g2028) & (g2305) & (g2309) & (!g2356) & (!g2843)) + ((!g1680) & (!g2028) & (g2305) & (g2309) & (!g2356) & (g2843)) + ((!g1680) & (!g2028) & (g2305) & (g2309) & (g2356) & (!g2843)) + ((!g1680) & (g2028) & (!g2305) & (g2309) & (!g2356) & (g2843)) + ((!g1680) & (g2028) & (g2305) & (!g2309) & (!g2356) & (!g2843)) + ((!g1680) & (g2028) & (g2305) & (!g2309) & (g2356) & (!g2843)) + ((!g1680) & (g2028) & (g2305) & (g2309) & (!g2356) & (!g2843)) + ((!g1680) & (g2028) & (g2305) & (g2309) & (!g2356) & (g2843)) + ((!g1680) & (g2028) & (g2305) & (g2309) & (g2356) & (!g2843)) + ((g1680) & (!g2028) & (!g2305) & (!g2309) & (g2356) & (g2843)) + ((g1680) & (!g2028) & (!g2305) & (g2309) & (g2356) & (g2843)) + ((g1680) & (!g2028) & (g2305) & (!g2309) & (!g2356) & (!g2843)) + ((g1680) & (!g2028) & (g2305) & (!g2309) & (!g2356) & (g2843)) + ((g1680) & (!g2028) & (g2305) & (!g2309) & (g2356) & (!g2843)) + ((g1680) & (!g2028) & (g2305) & (!g2309) & (g2356) & (g2843)) + ((g1680) & (!g2028) & (g2305) & (g2309) & (!g2356) & (!g2843)) + ((g1680) & (!g2028) & (g2305) & (g2309) & (!g2356) & (g2843)) + ((g1680) & (!g2028) & (g2305) & (g2309) & (g2356) & (!g2843)) + ((g1680) & (!g2028) & (g2305) & (g2309) & (g2356) & (g2843)) + ((g1680) & (g2028) & (!g2305) & (!g2309) & (g2356) & (g2843)) + ((g1680) & (g2028) & (!g2305) & (g2309) & (!g2356) & (g2843)) + ((g1680) & (g2028) & (!g2305) & (g2309) & (g2356) & (g2843)) + ((g1680) & (g2028) & (g2305) & (!g2309) & (!g2356) & (!g2843)) + ((g1680) & (g2028) & (g2305) & (!g2309) & (g2356) & (!g2843)) + ((g1680) & (g2028) & (g2305) & (!g2309) & (g2356) & (g2843)) + ((g1680) & (g2028) & (g2305) & (g2309) & (!g2356) & (!g2843)) + ((g1680) & (g2028) & (g2305) & (g2309) & (!g2356) & (g2843)) + ((g1680) & (g2028) & (g2305) & (g2309) & (g2356) & (!g2843)) + ((g1680) & (g2028) & (g2305) & (g2309) & (g2356) & (g2843)));
	assign g3061 = (((!g78) & (!g79) & (!g81) & (g2845) & (!sk[108]) & (!g2937)) + ((!g78) & (!g79) & (!g81) & (g2845) & (!sk[108]) & (g2937)) + ((!g78) & (!g79) & (g81) & (!g2845) & (!sk[108]) & (!g2937)) + ((!g78) & (!g79) & (g81) & (!g2845) & (!sk[108]) & (g2937)) + ((!g78) & (!g79) & (g81) & (g2845) & (!sk[108]) & (!g2937)) + ((!g78) & (!g79) & (g81) & (g2845) & (!sk[108]) & (g2937)) + ((!g78) & (!g79) & (g81) & (g2845) & (sk[108]) & (g2937)) + ((!g78) & (g79) & (!g81) & (g2845) & (!sk[108]) & (!g2937)) + ((!g78) & (g79) & (!g81) & (g2845) & (!sk[108]) & (g2937)) + ((!g78) & (g79) & (g81) & (!g2845) & (!sk[108]) & (!g2937)) + ((!g78) & (g79) & (g81) & (!g2845) & (!sk[108]) & (g2937)) + ((!g78) & (g79) & (g81) & (g2845) & (!sk[108]) & (!g2937)) + ((!g78) & (g79) & (g81) & (g2845) & (!sk[108]) & (g2937)) + ((g78) & (!g79) & (!g81) & (!g2845) & (!sk[108]) & (!g2937)) + ((g78) & (!g79) & (!g81) & (!g2845) & (!sk[108]) & (g2937)) + ((g78) & (!g79) & (!g81) & (g2845) & (!sk[108]) & (!g2937)) + ((g78) & (!g79) & (!g81) & (g2845) & (!sk[108]) & (g2937)) + ((g78) & (!g79) & (g81) & (!g2845) & (!sk[108]) & (!g2937)) + ((g78) & (!g79) & (g81) & (!g2845) & (!sk[108]) & (g2937)) + ((g78) & (!g79) & (g81) & (g2845) & (!sk[108]) & (!g2937)) + ((g78) & (!g79) & (g81) & (g2845) & (!sk[108]) & (g2937)) + ((g78) & (g79) & (!g81) & (!g2845) & (!sk[108]) & (!g2937)) + ((g78) & (g79) & (!g81) & (!g2845) & (!sk[108]) & (g2937)) + ((g78) & (g79) & (!g81) & (g2845) & (!sk[108]) & (!g2937)) + ((g78) & (g79) & (!g81) & (g2845) & (!sk[108]) & (g2937)) + ((g78) & (g79) & (g81) & (!g2845) & (!sk[108]) & (!g2937)) + ((g78) & (g79) & (g81) & (!g2845) & (!sk[108]) & (g2937)) + ((g78) & (g79) & (g81) & (g2845) & (!sk[108]) & (!g2937)) + ((g78) & (g79) & (g81) & (g2845) & (!sk[108]) & (g2937)));
	assign g3062 = (((!g2974) & (!g3043) & (sk[109]) & (!g3061)) + ((!g2974) & (g3043) & (!sk[109]) & (!g3061)) + ((!g2974) & (g3043) & (!sk[109]) & (g3061)) + ((g2974) & (!g3043) & (!sk[109]) & (!g3061)) + ((g2974) & (!g3043) & (!sk[109]) & (g3061)) + ((g2974) & (g3043) & (!sk[109]) & (!g3061)) + ((g2974) & (g3043) & (!sk[109]) & (g3061)));
	assign g3063 = (((!g118) & (!g85) & (!g86) & (g84) & (g93) & (!g2957)) + ((!g118) & (!g85) & (!g86) & (g84) & (g93) & (g2957)) + ((!g118) & (g85) & (!g86) & (g84) & (g93) & (!g2957)) + ((!g118) & (g85) & (!g86) & (g84) & (g93) & (g2957)) + ((g118) & (!g85) & (!g86) & (!g84) & (!g93) & (g2957)) + ((g118) & (!g85) & (!g86) & (!g84) & (g93) & (g2957)) + ((g118) & (!g85) & (!g86) & (g84) & (!g93) & (g2957)) + ((g118) & (!g85) & (!g86) & (g84) & (g93) & (!g2957)) + ((g118) & (!g85) & (!g86) & (g84) & (g93) & (g2957)) + ((g118) & (g85) & (!g86) & (g84) & (g93) & (!g2957)) + ((g118) & (g85) & (!g86) & (g84) & (g93) & (g2957)));
	assign g3064 = (((!g2954) & (!sk[111]) & (g3046) & (!g3063)) + ((!g2954) & (!sk[111]) & (g3046) & (g3063)) + ((g2954) & (!sk[111]) & (!g3046) & (!g3063)) + ((g2954) & (!sk[111]) & (!g3046) & (g3063)) + ((g2954) & (!sk[111]) & (g3046) & (!g3063)) + ((g2954) & (!sk[111]) & (g3046) & (g3063)) + ((g2954) & (sk[111]) & (g3046) & (!g3063)));
	assign g3065 = (((!g86) & (!g1680) & (!g3062) & (!sk[112]) & (g3064)) + ((!g86) & (!g1680) & (g3062) & (!sk[112]) & (g3064)) + ((!g86) & (g1680) & (!g3062) & (!sk[112]) & (!g3064)) + ((!g86) & (g1680) & (!g3062) & (!sk[112]) & (g3064)) + ((!g86) & (g1680) & (!g3062) & (sk[112]) & (g3064)) + ((!g86) & (g1680) & (g3062) & (!sk[112]) & (!g3064)) + ((!g86) & (g1680) & (g3062) & (!sk[112]) & (g3064)) + ((g86) & (!g1680) & (!g3062) & (!sk[112]) & (!g3064)) + ((g86) & (!g1680) & (!g3062) & (!sk[112]) & (g3064)) + ((g86) & (!g1680) & (g3062) & (!sk[112]) & (!g3064)) + ((g86) & (!g1680) & (g3062) & (!sk[112]) & (g3064)) + ((g86) & (!g1680) & (g3062) & (sk[112]) & (g3064)) + ((g86) & (g1680) & (!g3062) & (!sk[112]) & (!g3064)) + ((g86) & (g1680) & (!g3062) & (!sk[112]) & (g3064)) + ((g86) & (g1680) & (!g3062) & (sk[112]) & (g3064)) + ((g86) & (g1680) & (g3062) & (!sk[112]) & (!g3064)) + ((g86) & (g1680) & (g3062) & (!sk[112]) & (g3064)) + ((g86) & (g1680) & (g3062) & (sk[112]) & (g3064)));
	assign g3066 = (((!g1692) & (!g2028) & (g2332) & (!g2335) & (!g2356) & (!g2843)) + ((!g1692) & (!g2028) & (g2332) & (!g2335) & (!g2356) & (g2843)) + ((!g1692) & (!g2028) & (g2332) & (!g2335) & (g2356) & (!g2843)) + ((!g1692) & (!g2028) & (g2332) & (g2335) & (!g2356) & (!g2843)) + ((!g1692) & (!g2028) & (g2332) & (g2335) & (!g2356) & (g2843)) + ((!g1692) & (!g2028) & (g2332) & (g2335) & (g2356) & (!g2843)) + ((!g1692) & (g2028) & (!g2332) & (g2335) & (!g2356) & (g2843)) + ((!g1692) & (g2028) & (g2332) & (!g2335) & (!g2356) & (!g2843)) + ((!g1692) & (g2028) & (g2332) & (!g2335) & (g2356) & (!g2843)) + ((!g1692) & (g2028) & (g2332) & (g2335) & (!g2356) & (!g2843)) + ((!g1692) & (g2028) & (g2332) & (g2335) & (!g2356) & (g2843)) + ((!g1692) & (g2028) & (g2332) & (g2335) & (g2356) & (!g2843)) + ((g1692) & (!g2028) & (!g2332) & (!g2335) & (g2356) & (g2843)) + ((g1692) & (!g2028) & (!g2332) & (g2335) & (g2356) & (g2843)) + ((g1692) & (!g2028) & (g2332) & (!g2335) & (!g2356) & (!g2843)) + ((g1692) & (!g2028) & (g2332) & (!g2335) & (!g2356) & (g2843)) + ((g1692) & (!g2028) & (g2332) & (!g2335) & (g2356) & (!g2843)) + ((g1692) & (!g2028) & (g2332) & (!g2335) & (g2356) & (g2843)) + ((g1692) & (!g2028) & (g2332) & (g2335) & (!g2356) & (!g2843)) + ((g1692) & (!g2028) & (g2332) & (g2335) & (!g2356) & (g2843)) + ((g1692) & (!g2028) & (g2332) & (g2335) & (g2356) & (!g2843)) + ((g1692) & (!g2028) & (g2332) & (g2335) & (g2356) & (g2843)) + ((g1692) & (g2028) & (!g2332) & (!g2335) & (g2356) & (g2843)) + ((g1692) & (g2028) & (!g2332) & (g2335) & (!g2356) & (g2843)) + ((g1692) & (g2028) & (!g2332) & (g2335) & (g2356) & (g2843)) + ((g1692) & (g2028) & (g2332) & (!g2335) & (!g2356) & (!g2843)) + ((g1692) & (g2028) & (g2332) & (!g2335) & (g2356) & (!g2843)) + ((g1692) & (g2028) & (g2332) & (!g2335) & (g2356) & (g2843)) + ((g1692) & (g2028) & (g2332) & (g2335) & (!g2356) & (!g2843)) + ((g1692) & (g2028) & (g2332) & (g2335) & (!g2356) & (g2843)) + ((g1692) & (g2028) & (g2332) & (g2335) & (g2356) & (!g2843)) + ((g1692) & (g2028) & (g2332) & (g2335) & (g2356) & (g2843)));
	assign g3067 = (((!g85) & (!g1692) & (!g3062) & (!sk[114]) & (g3064)) + ((!g85) & (!g1692) & (g3062) & (!sk[114]) & (g3064)) + ((!g85) & (g1692) & (!g3062) & (!sk[114]) & (!g3064)) + ((!g85) & (g1692) & (!g3062) & (!sk[114]) & (g3064)) + ((!g85) & (g1692) & (!g3062) & (sk[114]) & (g3064)) + ((!g85) & (g1692) & (g3062) & (!sk[114]) & (!g3064)) + ((!g85) & (g1692) & (g3062) & (!sk[114]) & (g3064)) + ((g85) & (!g1692) & (!g3062) & (!sk[114]) & (!g3064)) + ((g85) & (!g1692) & (!g3062) & (!sk[114]) & (g3064)) + ((g85) & (!g1692) & (g3062) & (!sk[114]) & (!g3064)) + ((g85) & (!g1692) & (g3062) & (!sk[114]) & (g3064)) + ((g85) & (!g1692) & (g3062) & (sk[114]) & (g3064)) + ((g85) & (g1692) & (!g3062) & (!sk[114]) & (!g3064)) + ((g85) & (g1692) & (!g3062) & (!sk[114]) & (g3064)) + ((g85) & (g1692) & (!g3062) & (sk[114]) & (g3064)) + ((g85) & (g1692) & (g3062) & (!sk[114]) & (!g3064)) + ((g85) & (g1692) & (g3062) & (!sk[114]) & (g3064)) + ((g85) & (g1692) & (g3062) & (sk[114]) & (g3064)));
	assign g3068 = (((!g1705) & (!g2028) & (g2355) & (!g2356) & (!g2360) & (!g2843)) + ((!g1705) & (!g2028) & (g2355) & (!g2356) & (!g2360) & (g2843)) + ((!g1705) & (!g2028) & (g2355) & (!g2356) & (g2360) & (!g2843)) + ((!g1705) & (!g2028) & (g2355) & (!g2356) & (g2360) & (g2843)) + ((!g1705) & (!g2028) & (g2355) & (g2356) & (!g2360) & (!g2843)) + ((!g1705) & (!g2028) & (g2355) & (g2356) & (g2360) & (!g2843)) + ((!g1705) & (g2028) & (!g2355) & (!g2356) & (g2360) & (g2843)) + ((!g1705) & (g2028) & (g2355) & (!g2356) & (!g2360) & (!g2843)) + ((!g1705) & (g2028) & (g2355) & (!g2356) & (g2360) & (!g2843)) + ((!g1705) & (g2028) & (g2355) & (!g2356) & (g2360) & (g2843)) + ((!g1705) & (g2028) & (g2355) & (g2356) & (!g2360) & (!g2843)) + ((!g1705) & (g2028) & (g2355) & (g2356) & (g2360) & (!g2843)) + ((g1705) & (!g2028) & (!g2355) & (g2356) & (!g2360) & (g2843)) + ((g1705) & (!g2028) & (!g2355) & (g2356) & (g2360) & (g2843)) + ((g1705) & (!g2028) & (g2355) & (!g2356) & (!g2360) & (!g2843)) + ((g1705) & (!g2028) & (g2355) & (!g2356) & (!g2360) & (g2843)) + ((g1705) & (!g2028) & (g2355) & (!g2356) & (g2360) & (!g2843)) + ((g1705) & (!g2028) & (g2355) & (!g2356) & (g2360) & (g2843)) + ((g1705) & (!g2028) & (g2355) & (g2356) & (!g2360) & (!g2843)) + ((g1705) & (!g2028) & (g2355) & (g2356) & (!g2360) & (g2843)) + ((g1705) & (!g2028) & (g2355) & (g2356) & (g2360) & (!g2843)) + ((g1705) & (!g2028) & (g2355) & (g2356) & (g2360) & (g2843)) + ((g1705) & (g2028) & (!g2355) & (!g2356) & (g2360) & (g2843)) + ((g1705) & (g2028) & (!g2355) & (g2356) & (!g2360) & (g2843)) + ((g1705) & (g2028) & (!g2355) & (g2356) & (g2360) & (g2843)) + ((g1705) & (g2028) & (g2355) & (!g2356) & (!g2360) & (!g2843)) + ((g1705) & (g2028) & (g2355) & (!g2356) & (g2360) & (!g2843)) + ((g1705) & (g2028) & (g2355) & (!g2356) & (g2360) & (g2843)) + ((g1705) & (g2028) & (g2355) & (g2356) & (!g2360) & (!g2843)) + ((g1705) & (g2028) & (g2355) & (g2356) & (!g2360) & (g2843)) + ((g1705) & (g2028) & (g2355) & (g2356) & (g2360) & (!g2843)) + ((g1705) & (g2028) & (g2355) & (g2356) & (g2360) & (g2843)));
	assign g3069 = (((!g92) & (!sk[116]) & (!g1705) & (!g3062) & (g3064)) + ((!g92) & (!sk[116]) & (!g1705) & (g3062) & (g3064)) + ((!g92) & (!sk[116]) & (g1705) & (!g3062) & (!g3064)) + ((!g92) & (!sk[116]) & (g1705) & (!g3062) & (g3064)) + ((!g92) & (!sk[116]) & (g1705) & (g3062) & (!g3064)) + ((!g92) & (!sk[116]) & (g1705) & (g3062) & (g3064)) + ((!g92) & (sk[116]) & (g1705) & (!g3062) & (g3064)) + ((g92) & (!sk[116]) & (!g1705) & (!g3062) & (!g3064)) + ((g92) & (!sk[116]) & (!g1705) & (!g3062) & (g3064)) + ((g92) & (!sk[116]) & (!g1705) & (g3062) & (!g3064)) + ((g92) & (!sk[116]) & (!g1705) & (g3062) & (g3064)) + ((g92) & (!sk[116]) & (g1705) & (!g3062) & (!g3064)) + ((g92) & (!sk[116]) & (g1705) & (!g3062) & (g3064)) + ((g92) & (!sk[116]) & (g1705) & (g3062) & (!g3064)) + ((g92) & (!sk[116]) & (g1705) & (g3062) & (g3064)) + ((g92) & (sk[116]) & (!g1705) & (g3062) & (g3064)) + ((g92) & (sk[116]) & (g1705) & (!g3062) & (g3064)) + ((g92) & (sk[116]) & (g1705) & (g3062) & (g3064)));
	assign g3070 = (((!g1720) & (!g2028) & (!g2356) & (g2380) & (!g2387) & (!g2843)) + ((!g1720) & (!g2028) & (!g2356) & (g2380) & (!g2387) & (g2843)) + ((!g1720) & (!g2028) & (!g2356) & (g2380) & (g2387) & (!g2843)) + ((!g1720) & (!g2028) & (!g2356) & (g2380) & (g2387) & (g2843)) + ((!g1720) & (!g2028) & (g2356) & (g2380) & (!g2387) & (!g2843)) + ((!g1720) & (!g2028) & (g2356) & (g2380) & (g2387) & (!g2843)) + ((!g1720) & (g2028) & (!g2356) & (!g2380) & (!g2387) & (g2843)) + ((!g1720) & (g2028) & (!g2356) & (g2380) & (!g2387) & (!g2843)) + ((!g1720) & (g2028) & (!g2356) & (g2380) & (!g2387) & (g2843)) + ((!g1720) & (g2028) & (!g2356) & (g2380) & (g2387) & (!g2843)) + ((!g1720) & (g2028) & (g2356) & (g2380) & (!g2387) & (!g2843)) + ((!g1720) & (g2028) & (g2356) & (g2380) & (g2387) & (!g2843)) + ((g1720) & (!g2028) & (!g2356) & (g2380) & (!g2387) & (!g2843)) + ((g1720) & (!g2028) & (!g2356) & (g2380) & (!g2387) & (g2843)) + ((g1720) & (!g2028) & (!g2356) & (g2380) & (g2387) & (!g2843)) + ((g1720) & (!g2028) & (!g2356) & (g2380) & (g2387) & (g2843)) + ((g1720) & (!g2028) & (g2356) & (!g2380) & (!g2387) & (g2843)) + ((g1720) & (!g2028) & (g2356) & (!g2380) & (g2387) & (g2843)) + ((g1720) & (!g2028) & (g2356) & (g2380) & (!g2387) & (!g2843)) + ((g1720) & (!g2028) & (g2356) & (g2380) & (!g2387) & (g2843)) + ((g1720) & (!g2028) & (g2356) & (g2380) & (g2387) & (!g2843)) + ((g1720) & (!g2028) & (g2356) & (g2380) & (g2387) & (g2843)) + ((g1720) & (g2028) & (!g2356) & (!g2380) & (!g2387) & (g2843)) + ((g1720) & (g2028) & (!g2356) & (g2380) & (!g2387) & (!g2843)) + ((g1720) & (g2028) & (!g2356) & (g2380) & (!g2387) & (g2843)) + ((g1720) & (g2028) & (!g2356) & (g2380) & (g2387) & (!g2843)) + ((g1720) & (g2028) & (g2356) & (!g2380) & (!g2387) & (g2843)) + ((g1720) & (g2028) & (g2356) & (!g2380) & (g2387) & (g2843)) + ((g1720) & (g2028) & (g2356) & (g2380) & (!g2387) & (!g2843)) + ((g1720) & (g2028) & (g2356) & (g2380) & (!g2387) & (g2843)) + ((g1720) & (g2028) & (g2356) & (g2380) & (g2387) & (!g2843)) + ((g1720) & (g2028) & (g2356) & (g2380) & (g2387) & (g2843)));
	assign g3071 = (((!g91) & (!sk[118]) & (!g1720) & (!g3062) & (g3064)) + ((!g91) & (!sk[118]) & (!g1720) & (g3062) & (g3064)) + ((!g91) & (!sk[118]) & (g1720) & (!g3062) & (!g3064)) + ((!g91) & (!sk[118]) & (g1720) & (!g3062) & (g3064)) + ((!g91) & (!sk[118]) & (g1720) & (g3062) & (!g3064)) + ((!g91) & (!sk[118]) & (g1720) & (g3062) & (g3064)) + ((!g91) & (sk[118]) & (g1720) & (!g3062) & (g3064)) + ((g91) & (!sk[118]) & (!g1720) & (!g3062) & (!g3064)) + ((g91) & (!sk[118]) & (!g1720) & (!g3062) & (g3064)) + ((g91) & (!sk[118]) & (!g1720) & (g3062) & (!g3064)) + ((g91) & (!sk[118]) & (!g1720) & (g3062) & (g3064)) + ((g91) & (!sk[118]) & (g1720) & (!g3062) & (!g3064)) + ((g91) & (!sk[118]) & (g1720) & (!g3062) & (g3064)) + ((g91) & (!sk[118]) & (g1720) & (g3062) & (!g3064)) + ((g91) & (!sk[118]) & (g1720) & (g3062) & (g3064)) + ((g91) & (sk[118]) & (!g1720) & (g3062) & (g3064)) + ((g91) & (sk[118]) & (g1720) & (!g3062) & (g3064)) + ((g91) & (sk[118]) & (g1720) & (g3062) & (g3064)));
	assign g3072 = (((!g2412) & (!sk[119]) & (g2414)) + ((!g2412) & (sk[119]) & (!g2414)) + ((g2412) & (!sk[119]) & (g2414)));
	assign g3073 = (((!g1733) & (!g2028) & (!g2356) & (g2410) & (!g3072) & (!g2843)) + ((!g1733) & (!g2028) & (!g2356) & (g2410) & (!g3072) & (g2843)) + ((!g1733) & (!g2028) & (!g2356) & (g2410) & (g3072) & (!g2843)) + ((!g1733) & (!g2028) & (!g2356) & (g2410) & (g3072) & (g2843)) + ((!g1733) & (!g2028) & (g2356) & (g2410) & (!g3072) & (!g2843)) + ((!g1733) & (!g2028) & (g2356) & (g2410) & (g3072) & (!g2843)) + ((!g1733) & (g2028) & (!g2356) & (!g2410) & (!g3072) & (g2843)) + ((!g1733) & (g2028) & (!g2356) & (g2410) & (!g3072) & (!g2843)) + ((!g1733) & (g2028) & (!g2356) & (g2410) & (!g3072) & (g2843)) + ((!g1733) & (g2028) & (!g2356) & (g2410) & (g3072) & (!g2843)) + ((!g1733) & (g2028) & (g2356) & (g2410) & (!g3072) & (!g2843)) + ((!g1733) & (g2028) & (g2356) & (g2410) & (g3072) & (!g2843)) + ((g1733) & (!g2028) & (!g2356) & (g2410) & (!g3072) & (!g2843)) + ((g1733) & (!g2028) & (!g2356) & (g2410) & (!g3072) & (g2843)) + ((g1733) & (!g2028) & (!g2356) & (g2410) & (g3072) & (!g2843)) + ((g1733) & (!g2028) & (!g2356) & (g2410) & (g3072) & (g2843)) + ((g1733) & (!g2028) & (g2356) & (!g2410) & (!g3072) & (g2843)) + ((g1733) & (!g2028) & (g2356) & (!g2410) & (g3072) & (g2843)) + ((g1733) & (!g2028) & (g2356) & (g2410) & (!g3072) & (!g2843)) + ((g1733) & (!g2028) & (g2356) & (g2410) & (!g3072) & (g2843)) + ((g1733) & (!g2028) & (g2356) & (g2410) & (g3072) & (!g2843)) + ((g1733) & (!g2028) & (g2356) & (g2410) & (g3072) & (g2843)) + ((g1733) & (g2028) & (!g2356) & (!g2410) & (!g3072) & (g2843)) + ((g1733) & (g2028) & (!g2356) & (g2410) & (!g3072) & (!g2843)) + ((g1733) & (g2028) & (!g2356) & (g2410) & (!g3072) & (g2843)) + ((g1733) & (g2028) & (!g2356) & (g2410) & (g3072) & (!g2843)) + ((g1733) & (g2028) & (g2356) & (!g2410) & (!g3072) & (g2843)) + ((g1733) & (g2028) & (g2356) & (!g2410) & (g3072) & (g2843)) + ((g1733) & (g2028) & (g2356) & (g2410) & (!g3072) & (!g2843)) + ((g1733) & (g2028) & (g2356) & (g2410) & (!g3072) & (g2843)) + ((g1733) & (g2028) & (g2356) & (g2410) & (g3072) & (!g2843)) + ((g1733) & (g2028) & (g2356) & (g2410) & (g3072) & (g2843)));
	assign g3074 = (((!g1733) & (!g586) & (!sk[121]) & (!g3062) & (g3064)) + ((!g1733) & (!g586) & (!sk[121]) & (g3062) & (g3064)) + ((!g1733) & (g586) & (!sk[121]) & (!g3062) & (!g3064)) + ((!g1733) & (g586) & (!sk[121]) & (!g3062) & (g3064)) + ((!g1733) & (g586) & (!sk[121]) & (g3062) & (!g3064)) + ((!g1733) & (g586) & (!sk[121]) & (g3062) & (g3064)) + ((!g1733) & (g586) & (sk[121]) & (g3062) & (g3064)) + ((g1733) & (!g586) & (!sk[121]) & (!g3062) & (!g3064)) + ((g1733) & (!g586) & (!sk[121]) & (!g3062) & (g3064)) + ((g1733) & (!g586) & (!sk[121]) & (g3062) & (!g3064)) + ((g1733) & (!g586) & (!sk[121]) & (g3062) & (g3064)) + ((g1733) & (!g586) & (sk[121]) & (!g3062) & (g3064)) + ((g1733) & (g586) & (!sk[121]) & (!g3062) & (!g3064)) + ((g1733) & (g586) & (!sk[121]) & (!g3062) & (g3064)) + ((g1733) & (g586) & (!sk[121]) & (g3062) & (!g3064)) + ((g1733) & (g586) & (!sk[121]) & (g3062) & (g3064)) + ((g1733) & (g586) & (sk[121]) & (!g3062) & (g3064)) + ((g1733) & (g586) & (sk[121]) & (g3062) & (g3064)));
	assign g3075 = (((!g1746) & (!g2028) & (!g2356) & (!g2435) & (g2436) & (!g2843)) + ((!g1746) & (!g2028) & (!g2356) & (!g2435) & (g2436) & (g2843)) + ((!g1746) & (!g2028) & (!g2356) & (g2435) & (g2436) & (!g2843)) + ((!g1746) & (!g2028) & (!g2356) & (g2435) & (g2436) & (g2843)) + ((!g1746) & (!g2028) & (g2356) & (!g2435) & (g2436) & (!g2843)) + ((!g1746) & (!g2028) & (g2356) & (g2435) & (g2436) & (!g2843)) + ((!g1746) & (g2028) & (!g2356) & (!g2435) & (g2436) & (!g2843)) + ((!g1746) & (g2028) & (!g2356) & (g2435) & (!g2436) & (g2843)) + ((!g1746) & (g2028) & (!g2356) & (g2435) & (g2436) & (!g2843)) + ((!g1746) & (g2028) & (!g2356) & (g2435) & (g2436) & (g2843)) + ((!g1746) & (g2028) & (g2356) & (!g2435) & (g2436) & (!g2843)) + ((!g1746) & (g2028) & (g2356) & (g2435) & (g2436) & (!g2843)) + ((g1746) & (!g2028) & (!g2356) & (!g2435) & (g2436) & (!g2843)) + ((g1746) & (!g2028) & (!g2356) & (!g2435) & (g2436) & (g2843)) + ((g1746) & (!g2028) & (!g2356) & (g2435) & (g2436) & (!g2843)) + ((g1746) & (!g2028) & (!g2356) & (g2435) & (g2436) & (g2843)) + ((g1746) & (!g2028) & (g2356) & (!g2435) & (!g2436) & (g2843)) + ((g1746) & (!g2028) & (g2356) & (!g2435) & (g2436) & (!g2843)) + ((g1746) & (!g2028) & (g2356) & (!g2435) & (g2436) & (g2843)) + ((g1746) & (!g2028) & (g2356) & (g2435) & (!g2436) & (g2843)) + ((g1746) & (!g2028) & (g2356) & (g2435) & (g2436) & (!g2843)) + ((g1746) & (!g2028) & (g2356) & (g2435) & (g2436) & (g2843)) + ((g1746) & (g2028) & (!g2356) & (!g2435) & (g2436) & (!g2843)) + ((g1746) & (g2028) & (!g2356) & (g2435) & (!g2436) & (g2843)) + ((g1746) & (g2028) & (!g2356) & (g2435) & (g2436) & (!g2843)) + ((g1746) & (g2028) & (!g2356) & (g2435) & (g2436) & (g2843)) + ((g1746) & (g2028) & (g2356) & (!g2435) & (!g2436) & (g2843)) + ((g1746) & (g2028) & (g2356) & (!g2435) & (g2436) & (!g2843)) + ((g1746) & (g2028) & (g2356) & (!g2435) & (g2436) & (g2843)) + ((g1746) & (g2028) & (g2356) & (g2435) & (!g2436) & (g2843)) + ((g1746) & (g2028) & (g2356) & (g2435) & (g2436) & (!g2843)) + ((g1746) & (g2028) & (g2356) & (g2435) & (g2436) & (g2843)));
	assign g3076 = (((!g677) & (!g1746) & (!sk[123]) & (!g3062) & (g3064)) + ((!g677) & (!g1746) & (!sk[123]) & (g3062) & (g3064)) + ((!g677) & (g1746) & (!sk[123]) & (!g3062) & (!g3064)) + ((!g677) & (g1746) & (!sk[123]) & (!g3062) & (g3064)) + ((!g677) & (g1746) & (!sk[123]) & (g3062) & (!g3064)) + ((!g677) & (g1746) & (!sk[123]) & (g3062) & (g3064)) + ((!g677) & (g1746) & (sk[123]) & (!g3062) & (g3064)) + ((g677) & (!g1746) & (!sk[123]) & (!g3062) & (!g3064)) + ((g677) & (!g1746) & (!sk[123]) & (!g3062) & (g3064)) + ((g677) & (!g1746) & (!sk[123]) & (g3062) & (!g3064)) + ((g677) & (!g1746) & (!sk[123]) & (g3062) & (g3064)) + ((g677) & (!g1746) & (sk[123]) & (g3062) & (g3064)) + ((g677) & (g1746) & (!sk[123]) & (!g3062) & (!g3064)) + ((g677) & (g1746) & (!sk[123]) & (!g3062) & (g3064)) + ((g677) & (g1746) & (!sk[123]) & (g3062) & (!g3064)) + ((g677) & (g1746) & (!sk[123]) & (g3062) & (g3064)) + ((g677) & (g1746) & (sk[123]) & (!g3062) & (g3064)) + ((g677) & (g1746) & (sk[123]) & (g3062) & (g3064)));
	assign g3077 = (((!g726) & (!g1759) & (!g3062) & (!sk[124]) & (g3064)) + ((!g726) & (!g1759) & (g3062) & (!sk[124]) & (g3064)) + ((!g726) & (g1759) & (!g3062) & (!sk[124]) & (!g3064)) + ((!g726) & (g1759) & (!g3062) & (!sk[124]) & (g3064)) + ((!g726) & (g1759) & (!g3062) & (sk[124]) & (g3064)) + ((!g726) & (g1759) & (g3062) & (!sk[124]) & (!g3064)) + ((!g726) & (g1759) & (g3062) & (!sk[124]) & (g3064)) + ((g726) & (!g1759) & (!g3062) & (!sk[124]) & (!g3064)) + ((g726) & (!g1759) & (!g3062) & (!sk[124]) & (g3064)) + ((g726) & (!g1759) & (g3062) & (!sk[124]) & (!g3064)) + ((g726) & (!g1759) & (g3062) & (!sk[124]) & (g3064)) + ((g726) & (!g1759) & (g3062) & (sk[124]) & (g3064)) + ((g726) & (g1759) & (!g3062) & (!sk[124]) & (!g3064)) + ((g726) & (g1759) & (!g3062) & (!sk[124]) & (g3064)) + ((g726) & (g1759) & (!g3062) & (sk[124]) & (g3064)) + ((g726) & (g1759) & (g3062) & (!sk[124]) & (!g3064)) + ((g726) & (g1759) & (g3062) & (!sk[124]) & (g3064)) + ((g726) & (g1759) & (g3062) & (sk[124]) & (g3064)));
	assign g3078 = (((!sk[125]) & (!g773) & (!g1772) & (!g3062) & (g3064)) + ((!sk[125]) & (!g773) & (!g1772) & (g3062) & (g3064)) + ((!sk[125]) & (!g773) & (g1772) & (!g3062) & (!g3064)) + ((!sk[125]) & (!g773) & (g1772) & (!g3062) & (g3064)) + ((!sk[125]) & (!g773) & (g1772) & (g3062) & (!g3064)) + ((!sk[125]) & (!g773) & (g1772) & (g3062) & (g3064)) + ((!sk[125]) & (g773) & (!g1772) & (!g3062) & (!g3064)) + ((!sk[125]) & (g773) & (!g1772) & (!g3062) & (g3064)) + ((!sk[125]) & (g773) & (!g1772) & (g3062) & (!g3064)) + ((!sk[125]) & (g773) & (!g1772) & (g3062) & (g3064)) + ((!sk[125]) & (g773) & (g1772) & (!g3062) & (!g3064)) + ((!sk[125]) & (g773) & (g1772) & (!g3062) & (g3064)) + ((!sk[125]) & (g773) & (g1772) & (g3062) & (!g3064)) + ((!sk[125]) & (g773) & (g1772) & (g3062) & (g3064)) + ((sk[125]) & (!g773) & (g1772) & (!g3062) & (g3064)) + ((sk[125]) & (g773) & (!g1772) & (g3062) & (g3064)) + ((sk[125]) & (g773) & (g1772) & (!g3062) & (g3064)) + ((sk[125]) & (g773) & (g1772) & (g3062) & (g3064)));
	assign g3079 = (((!sk[126]) & (!g2498) & (g2503)) + ((!sk[126]) & (g2498) & (g2503)) + ((sk[126]) & (!g2498) & (!g2503)));
	assign g3080 = (((!g1772) & (!g2028) & (!g2356) & (g2497) & (!g3079) & (!g2843)) + ((!g1772) & (!g2028) & (!g2356) & (g2497) & (!g3079) & (g2843)) + ((!g1772) & (!g2028) & (!g2356) & (g2497) & (g3079) & (!g2843)) + ((!g1772) & (!g2028) & (!g2356) & (g2497) & (g3079) & (g2843)) + ((!g1772) & (!g2028) & (g2356) & (g2497) & (!g3079) & (!g2843)) + ((!g1772) & (!g2028) & (g2356) & (g2497) & (g3079) & (!g2843)) + ((!g1772) & (g2028) & (!g2356) & (!g2497) & (!g3079) & (g2843)) + ((!g1772) & (g2028) & (!g2356) & (g2497) & (!g3079) & (!g2843)) + ((!g1772) & (g2028) & (!g2356) & (g2497) & (!g3079) & (g2843)) + ((!g1772) & (g2028) & (!g2356) & (g2497) & (g3079) & (!g2843)) + ((!g1772) & (g2028) & (g2356) & (g2497) & (!g3079) & (!g2843)) + ((!g1772) & (g2028) & (g2356) & (g2497) & (g3079) & (!g2843)) + ((g1772) & (!g2028) & (!g2356) & (g2497) & (!g3079) & (!g2843)) + ((g1772) & (!g2028) & (!g2356) & (g2497) & (!g3079) & (g2843)) + ((g1772) & (!g2028) & (!g2356) & (g2497) & (g3079) & (!g2843)) + ((g1772) & (!g2028) & (!g2356) & (g2497) & (g3079) & (g2843)) + ((g1772) & (!g2028) & (g2356) & (!g2497) & (!g3079) & (g2843)) + ((g1772) & (!g2028) & (g2356) & (!g2497) & (g3079) & (g2843)) + ((g1772) & (!g2028) & (g2356) & (g2497) & (!g3079) & (!g2843)) + ((g1772) & (!g2028) & (g2356) & (g2497) & (!g3079) & (g2843)) + ((g1772) & (!g2028) & (g2356) & (g2497) & (g3079) & (!g2843)) + ((g1772) & (!g2028) & (g2356) & (g2497) & (g3079) & (g2843)) + ((g1772) & (g2028) & (!g2356) & (!g2497) & (!g3079) & (g2843)) + ((g1772) & (g2028) & (!g2356) & (g2497) & (!g3079) & (!g2843)) + ((g1772) & (g2028) & (!g2356) & (g2497) & (!g3079) & (g2843)) + ((g1772) & (g2028) & (!g2356) & (g2497) & (g3079) & (!g2843)) + ((g1772) & (g2028) & (g2356) & (!g2497) & (!g3079) & (g2843)) + ((g1772) & (g2028) & (g2356) & (!g2497) & (g3079) & (g2843)) + ((g1772) & (g2028) & (g2356) & (g2497) & (!g3079) & (!g2843)) + ((g1772) & (g2028) & (g2356) & (g2497) & (!g3079) & (g2843)) + ((g1772) & (g2028) & (g2356) & (g2497) & (g3079) & (!g2843)) + ((g1772) & (g2028) & (g2356) & (g2497) & (g3079) & (g2843)));
	assign g3081 = (((!g820) & (!sk[0]) & (!g1785) & (!g3062) & (g3064)) + ((!g820) & (!sk[0]) & (!g1785) & (g3062) & (g3064)) + ((!g820) & (!sk[0]) & (g1785) & (!g3062) & (!g3064)) + ((!g820) & (!sk[0]) & (g1785) & (!g3062) & (g3064)) + ((!g820) & (!sk[0]) & (g1785) & (g3062) & (!g3064)) + ((!g820) & (!sk[0]) & (g1785) & (g3062) & (g3064)) + ((!g820) & (sk[0]) & (g1785) & (!g3062) & (g3064)) + ((g820) & (!sk[0]) & (!g1785) & (!g3062) & (!g3064)) + ((g820) & (!sk[0]) & (!g1785) & (!g3062) & (g3064)) + ((g820) & (!sk[0]) & (!g1785) & (g3062) & (!g3064)) + ((g820) & (!sk[0]) & (!g1785) & (g3062) & (g3064)) + ((g820) & (!sk[0]) & (g1785) & (!g3062) & (!g3064)) + ((g820) & (!sk[0]) & (g1785) & (!g3062) & (g3064)) + ((g820) & (!sk[0]) & (g1785) & (g3062) & (!g3064)) + ((g820) & (!sk[0]) & (g1785) & (g3062) & (g3064)) + ((g820) & (sk[0]) & (!g1785) & (g3062) & (g3064)) + ((g820) & (sk[0]) & (g1785) & (!g3062) & (g3064)) + ((g820) & (sk[0]) & (g1785) & (g3062) & (g3064)));
	assign g3082 = (((!g867) & (!g1798) & (!g3062) & (!sk[1]) & (g3064)) + ((!g867) & (!g1798) & (g3062) & (!sk[1]) & (g3064)) + ((!g867) & (g1798) & (!g3062) & (!sk[1]) & (!g3064)) + ((!g867) & (g1798) & (!g3062) & (!sk[1]) & (g3064)) + ((!g867) & (g1798) & (!g3062) & (sk[1]) & (g3064)) + ((!g867) & (g1798) & (g3062) & (!sk[1]) & (!g3064)) + ((!g867) & (g1798) & (g3062) & (!sk[1]) & (g3064)) + ((g867) & (!g1798) & (!g3062) & (!sk[1]) & (!g3064)) + ((g867) & (!g1798) & (!g3062) & (!sk[1]) & (g3064)) + ((g867) & (!g1798) & (g3062) & (!sk[1]) & (!g3064)) + ((g867) & (!g1798) & (g3062) & (!sk[1]) & (g3064)) + ((g867) & (!g1798) & (g3062) & (sk[1]) & (g3064)) + ((g867) & (g1798) & (!g3062) & (!sk[1]) & (!g3064)) + ((g867) & (g1798) & (!g3062) & (!sk[1]) & (g3064)) + ((g867) & (g1798) & (!g3062) & (sk[1]) & (g3064)) + ((g867) & (g1798) & (g3062) & (!sk[1]) & (!g3064)) + ((g867) & (g1798) & (g3062) & (!sk[1]) & (g3064)) + ((g867) & (g1798) & (g3062) & (sk[1]) & (g3064)));
	assign g3083 = (((!g1798) & (!g2028) & (!g2356) & (g2543) & (!g2547) & (!g2843)) + ((!g1798) & (!g2028) & (!g2356) & (g2543) & (!g2547) & (g2843)) + ((!g1798) & (!g2028) & (!g2356) & (g2543) & (g2547) & (!g2843)) + ((!g1798) & (!g2028) & (!g2356) & (g2543) & (g2547) & (g2843)) + ((!g1798) & (!g2028) & (g2356) & (g2543) & (!g2547) & (!g2843)) + ((!g1798) & (!g2028) & (g2356) & (g2543) & (g2547) & (!g2843)) + ((!g1798) & (g2028) & (!g2356) & (!g2543) & (g2547) & (g2843)) + ((!g1798) & (g2028) & (!g2356) & (g2543) & (!g2547) & (!g2843)) + ((!g1798) & (g2028) & (!g2356) & (g2543) & (g2547) & (!g2843)) + ((!g1798) & (g2028) & (!g2356) & (g2543) & (g2547) & (g2843)) + ((!g1798) & (g2028) & (g2356) & (g2543) & (!g2547) & (!g2843)) + ((!g1798) & (g2028) & (g2356) & (g2543) & (g2547) & (!g2843)) + ((g1798) & (!g2028) & (!g2356) & (g2543) & (!g2547) & (!g2843)) + ((g1798) & (!g2028) & (!g2356) & (g2543) & (!g2547) & (g2843)) + ((g1798) & (!g2028) & (!g2356) & (g2543) & (g2547) & (!g2843)) + ((g1798) & (!g2028) & (!g2356) & (g2543) & (g2547) & (g2843)) + ((g1798) & (!g2028) & (g2356) & (!g2543) & (!g2547) & (g2843)) + ((g1798) & (!g2028) & (g2356) & (!g2543) & (g2547) & (g2843)) + ((g1798) & (!g2028) & (g2356) & (g2543) & (!g2547) & (!g2843)) + ((g1798) & (!g2028) & (g2356) & (g2543) & (!g2547) & (g2843)) + ((g1798) & (!g2028) & (g2356) & (g2543) & (g2547) & (!g2843)) + ((g1798) & (!g2028) & (g2356) & (g2543) & (g2547) & (g2843)) + ((g1798) & (g2028) & (!g2356) & (!g2543) & (g2547) & (g2843)) + ((g1798) & (g2028) & (!g2356) & (g2543) & (!g2547) & (!g2843)) + ((g1798) & (g2028) & (!g2356) & (g2543) & (g2547) & (!g2843)) + ((g1798) & (g2028) & (!g2356) & (g2543) & (g2547) & (g2843)) + ((g1798) & (g2028) & (g2356) & (!g2543) & (!g2547) & (g2843)) + ((g1798) & (g2028) & (g2356) & (!g2543) & (g2547) & (g2843)) + ((g1798) & (g2028) & (g2356) & (g2543) & (!g2547) & (!g2843)) + ((g1798) & (g2028) & (g2356) & (g2543) & (!g2547) & (g2843)) + ((g1798) & (g2028) & (g2356) & (g2543) & (g2547) & (!g2843)) + ((g1798) & (g2028) & (g2356) & (g2543) & (g2547) & (g2843)));
	assign g3084 = (((!sk[3]) & (!g2931) & (!g867) & (!g2955) & (g2958)) + ((!sk[3]) & (!g2931) & (!g867) & (g2955) & (g2958)) + ((!sk[3]) & (!g2931) & (g867) & (!g2955) & (!g2958)) + ((!sk[3]) & (!g2931) & (g867) & (!g2955) & (g2958)) + ((!sk[3]) & (!g2931) & (g867) & (g2955) & (!g2958)) + ((!sk[3]) & (!g2931) & (g867) & (g2955) & (g2958)) + ((!sk[3]) & (g2931) & (!g867) & (!g2955) & (!g2958)) + ((!sk[3]) & (g2931) & (!g867) & (!g2955) & (g2958)) + ((!sk[3]) & (g2931) & (!g867) & (g2955) & (!g2958)) + ((!sk[3]) & (g2931) & (!g867) & (g2955) & (g2958)) + ((!sk[3]) & (g2931) & (g867) & (!g2955) & (!g2958)) + ((!sk[3]) & (g2931) & (g867) & (!g2955) & (g2958)) + ((!sk[3]) & (g2931) & (g867) & (g2955) & (!g2958)) + ((!sk[3]) & (g2931) & (g867) & (g2955) & (g2958)) + ((sk[3]) & (!g2931) & (g867) & (!g2955) & (g2958)) + ((sk[3]) & (!g2931) & (g867) & (g2955) & (!g2958)) + ((sk[3]) & (!g2931) & (g867) & (g2955) & (g2958)) + ((sk[3]) & (g2931) & (g867) & (!g2955) & (!g2958)) + ((sk[3]) & (g2931) & (g867) & (!g2955) & (g2958)) + ((sk[3]) & (g2931) & (g867) & (g2955) & (!g2958)) + ((sk[3]) & (g2931) & (g867) & (g2955) & (g2958)));
	assign g3085 = (((!g1810) & (!g3062) & (sk[4]) & (g3084)) + ((!g1810) & (g3062) & (!sk[4]) & (!g3084)) + ((!g1810) & (g3062) & (!sk[4]) & (g3084)) + ((!g1810) & (g3062) & (sk[4]) & (g3084)) + ((g1810) & (!g3062) & (!sk[4]) & (!g3084)) + ((g1810) & (!g3062) & (!sk[4]) & (g3084)) + ((g1810) & (!g3062) & (sk[4]) & (!g3084)) + ((g1810) & (!g3062) & (sk[4]) & (g3084)) + ((g1810) & (g3062) & (!sk[4]) & (!g3084)) + ((g1810) & (g3062) & (!sk[4]) & (g3084)) + ((g1810) & (g3062) & (sk[4]) & (g3084)));
	assign g3086 = (((!g2565) & (!sk[5]) & (g2568)) + ((!g2565) & (sk[5]) & (!g2568)) + ((g2565) & (!sk[5]) & (g2568)));
	assign g3087 = (((!g1810) & (!g2028) & (!g2356) & (g2564) & (!g3086) & (!g2843)) + ((!g1810) & (!g2028) & (!g2356) & (g2564) & (!g3086) & (g2843)) + ((!g1810) & (!g2028) & (!g2356) & (g2564) & (g3086) & (!g2843)) + ((!g1810) & (!g2028) & (!g2356) & (g2564) & (g3086) & (g2843)) + ((!g1810) & (!g2028) & (g2356) & (g2564) & (!g3086) & (!g2843)) + ((!g1810) & (!g2028) & (g2356) & (g2564) & (g3086) & (!g2843)) + ((!g1810) & (g2028) & (!g2356) & (!g2564) & (!g3086) & (g2843)) + ((!g1810) & (g2028) & (!g2356) & (g2564) & (!g3086) & (!g2843)) + ((!g1810) & (g2028) & (!g2356) & (g2564) & (!g3086) & (g2843)) + ((!g1810) & (g2028) & (!g2356) & (g2564) & (g3086) & (!g2843)) + ((!g1810) & (g2028) & (g2356) & (g2564) & (!g3086) & (!g2843)) + ((!g1810) & (g2028) & (g2356) & (g2564) & (g3086) & (!g2843)) + ((g1810) & (!g2028) & (!g2356) & (g2564) & (!g3086) & (!g2843)) + ((g1810) & (!g2028) & (!g2356) & (g2564) & (!g3086) & (g2843)) + ((g1810) & (!g2028) & (!g2356) & (g2564) & (g3086) & (!g2843)) + ((g1810) & (!g2028) & (!g2356) & (g2564) & (g3086) & (g2843)) + ((g1810) & (!g2028) & (g2356) & (!g2564) & (!g3086) & (g2843)) + ((g1810) & (!g2028) & (g2356) & (!g2564) & (g3086) & (g2843)) + ((g1810) & (!g2028) & (g2356) & (g2564) & (!g3086) & (!g2843)) + ((g1810) & (!g2028) & (g2356) & (g2564) & (!g3086) & (g2843)) + ((g1810) & (!g2028) & (g2356) & (g2564) & (g3086) & (!g2843)) + ((g1810) & (!g2028) & (g2356) & (g2564) & (g3086) & (g2843)) + ((g1810) & (g2028) & (!g2356) & (!g2564) & (!g3086) & (g2843)) + ((g1810) & (g2028) & (!g2356) & (g2564) & (!g3086) & (!g2843)) + ((g1810) & (g2028) & (!g2356) & (g2564) & (!g3086) & (g2843)) + ((g1810) & (g2028) & (!g2356) & (g2564) & (g3086) & (!g2843)) + ((g1810) & (g2028) & (g2356) & (!g2564) & (!g3086) & (g2843)) + ((g1810) & (g2028) & (g2356) & (!g2564) & (g3086) & (g2843)) + ((g1810) & (g2028) & (g2356) & (g2564) & (!g3086) & (!g2843)) + ((g1810) & (g2028) & (g2356) & (g2564) & (!g3086) & (g2843)) + ((g1810) & (g2028) & (g2356) & (g2564) & (g3086) & (!g2843)) + ((g1810) & (g2028) & (g2356) & (g2564) & (g3086) & (g2843)));
	assign g3088 = (((!g1824) & (!sk[7]) & (g3062) & (!g3084)) + ((!g1824) & (!sk[7]) & (g3062) & (g3084)) + ((!g1824) & (sk[7]) & (!g3062) & (g3084)) + ((!g1824) & (sk[7]) & (g3062) & (g3084)) + ((g1824) & (!sk[7]) & (!g3062) & (!g3084)) + ((g1824) & (!sk[7]) & (!g3062) & (g3084)) + ((g1824) & (!sk[7]) & (g3062) & (!g3084)) + ((g1824) & (!sk[7]) & (g3062) & (g3084)) + ((g1824) & (sk[7]) & (!g3062) & (!g3084)) + ((g1824) & (sk[7]) & (!g3062) & (g3084)) + ((g1824) & (sk[7]) & (g3062) & (g3084)));
	assign g3089 = (((!sk[8]) & (!g1837) & (g3062) & (!g3084)) + ((!sk[8]) & (!g1837) & (g3062) & (g3084)) + ((!sk[8]) & (g1837) & (!g3062) & (!g3084)) + ((!sk[8]) & (g1837) & (!g3062) & (g3084)) + ((!sk[8]) & (g1837) & (g3062) & (!g3084)) + ((!sk[8]) & (g1837) & (g3062) & (g3084)) + ((sk[8]) & (!g1837) & (!g3062) & (g3084)) + ((sk[8]) & (!g1837) & (g3062) & (g3084)) + ((sk[8]) & (g1837) & (!g3062) & (!g3084)) + ((sk[8]) & (g1837) & (!g3062) & (g3084)) + ((sk[8]) & (g1837) & (g3062) & (g3084)));
	assign g3090 = (((!sk[9]) & (!g1850) & (g3062) & (!g3084)) + ((!sk[9]) & (!g1850) & (g3062) & (g3084)) + ((!sk[9]) & (g1850) & (!g3062) & (!g3084)) + ((!sk[9]) & (g1850) & (!g3062) & (g3084)) + ((!sk[9]) & (g1850) & (g3062) & (!g3084)) + ((!sk[9]) & (g1850) & (g3062) & (g3084)) + ((sk[9]) & (!g1850) & (!g3062) & (g3084)) + ((sk[9]) & (!g1850) & (g3062) & (g3084)) + ((sk[9]) & (g1850) & (!g3062) & (!g3084)) + ((sk[9]) & (g1850) & (!g3062) & (g3084)) + ((sk[9]) & (g1850) & (g3062) & (g3084)));
	assign g3091 = (((!g1850) & (!g2028) & (!g2356) & (g2620) & (!g2623) & (!g2843)) + ((!g1850) & (!g2028) & (!g2356) & (g2620) & (!g2623) & (g2843)) + ((!g1850) & (!g2028) & (!g2356) & (g2620) & (g2623) & (!g2843)) + ((!g1850) & (!g2028) & (!g2356) & (g2620) & (g2623) & (g2843)) + ((!g1850) & (!g2028) & (g2356) & (g2620) & (!g2623) & (!g2843)) + ((!g1850) & (!g2028) & (g2356) & (g2620) & (g2623) & (!g2843)) + ((!g1850) & (g2028) & (!g2356) & (!g2620) & (g2623) & (g2843)) + ((!g1850) & (g2028) & (!g2356) & (g2620) & (!g2623) & (!g2843)) + ((!g1850) & (g2028) & (!g2356) & (g2620) & (g2623) & (!g2843)) + ((!g1850) & (g2028) & (!g2356) & (g2620) & (g2623) & (g2843)) + ((!g1850) & (g2028) & (g2356) & (g2620) & (!g2623) & (!g2843)) + ((!g1850) & (g2028) & (g2356) & (g2620) & (g2623) & (!g2843)) + ((g1850) & (!g2028) & (!g2356) & (g2620) & (!g2623) & (!g2843)) + ((g1850) & (!g2028) & (!g2356) & (g2620) & (!g2623) & (g2843)) + ((g1850) & (!g2028) & (!g2356) & (g2620) & (g2623) & (!g2843)) + ((g1850) & (!g2028) & (!g2356) & (g2620) & (g2623) & (g2843)) + ((g1850) & (!g2028) & (g2356) & (!g2620) & (!g2623) & (g2843)) + ((g1850) & (!g2028) & (g2356) & (!g2620) & (g2623) & (g2843)) + ((g1850) & (!g2028) & (g2356) & (g2620) & (!g2623) & (!g2843)) + ((g1850) & (!g2028) & (g2356) & (g2620) & (!g2623) & (g2843)) + ((g1850) & (!g2028) & (g2356) & (g2620) & (g2623) & (!g2843)) + ((g1850) & (!g2028) & (g2356) & (g2620) & (g2623) & (g2843)) + ((g1850) & (g2028) & (!g2356) & (!g2620) & (g2623) & (g2843)) + ((g1850) & (g2028) & (!g2356) & (g2620) & (!g2623) & (!g2843)) + ((g1850) & (g2028) & (!g2356) & (g2620) & (g2623) & (!g2843)) + ((g1850) & (g2028) & (!g2356) & (g2620) & (g2623) & (g2843)) + ((g1850) & (g2028) & (g2356) & (!g2620) & (!g2623) & (g2843)) + ((g1850) & (g2028) & (g2356) & (!g2620) & (g2623) & (g2843)) + ((g1850) & (g2028) & (g2356) & (g2620) & (!g2623) & (!g2843)) + ((g1850) & (g2028) & (g2356) & (g2620) & (!g2623) & (g2843)) + ((g1850) & (g2028) & (g2356) & (g2620) & (g2623) & (!g2843)) + ((g1850) & (g2028) & (g2356) & (g2620) & (g2623) & (g2843)));
	assign g3092 = (((!g1863) & (!g3062) & (sk[11]) & (g3084)) + ((!g1863) & (g3062) & (!sk[11]) & (!g3084)) + ((!g1863) & (g3062) & (!sk[11]) & (g3084)) + ((!g1863) & (g3062) & (sk[11]) & (g3084)) + ((g1863) & (!g3062) & (!sk[11]) & (!g3084)) + ((g1863) & (!g3062) & (!sk[11]) & (g3084)) + ((g1863) & (!g3062) & (sk[11]) & (!g3084)) + ((g1863) & (!g3062) & (sk[11]) & (g3084)) + ((g1863) & (g3062) & (!sk[11]) & (!g3084)) + ((g1863) & (g3062) & (!sk[11]) & (g3084)) + ((g1863) & (g3062) & (sk[11]) & (g3084)));
	assign g3093 = (((!g1863) & (!g2028) & (!g2356) & (g2636) & (!g2640) & (!g2843)) + ((!g1863) & (!g2028) & (!g2356) & (g2636) & (!g2640) & (g2843)) + ((!g1863) & (!g2028) & (!g2356) & (g2636) & (g2640) & (!g2843)) + ((!g1863) & (!g2028) & (!g2356) & (g2636) & (g2640) & (g2843)) + ((!g1863) & (!g2028) & (g2356) & (g2636) & (!g2640) & (!g2843)) + ((!g1863) & (!g2028) & (g2356) & (g2636) & (g2640) & (!g2843)) + ((!g1863) & (g2028) & (!g2356) & (!g2636) & (g2640) & (g2843)) + ((!g1863) & (g2028) & (!g2356) & (g2636) & (!g2640) & (!g2843)) + ((!g1863) & (g2028) & (!g2356) & (g2636) & (g2640) & (!g2843)) + ((!g1863) & (g2028) & (!g2356) & (g2636) & (g2640) & (g2843)) + ((!g1863) & (g2028) & (g2356) & (g2636) & (!g2640) & (!g2843)) + ((!g1863) & (g2028) & (g2356) & (g2636) & (g2640) & (!g2843)) + ((g1863) & (!g2028) & (!g2356) & (g2636) & (!g2640) & (!g2843)) + ((g1863) & (!g2028) & (!g2356) & (g2636) & (!g2640) & (g2843)) + ((g1863) & (!g2028) & (!g2356) & (g2636) & (g2640) & (!g2843)) + ((g1863) & (!g2028) & (!g2356) & (g2636) & (g2640) & (g2843)) + ((g1863) & (!g2028) & (g2356) & (!g2636) & (!g2640) & (g2843)) + ((g1863) & (!g2028) & (g2356) & (!g2636) & (g2640) & (g2843)) + ((g1863) & (!g2028) & (g2356) & (g2636) & (!g2640) & (!g2843)) + ((g1863) & (!g2028) & (g2356) & (g2636) & (!g2640) & (g2843)) + ((g1863) & (!g2028) & (g2356) & (g2636) & (g2640) & (!g2843)) + ((g1863) & (!g2028) & (g2356) & (g2636) & (g2640) & (g2843)) + ((g1863) & (g2028) & (!g2356) & (!g2636) & (g2640) & (g2843)) + ((g1863) & (g2028) & (!g2356) & (g2636) & (!g2640) & (!g2843)) + ((g1863) & (g2028) & (!g2356) & (g2636) & (g2640) & (!g2843)) + ((g1863) & (g2028) & (!g2356) & (g2636) & (g2640) & (g2843)) + ((g1863) & (g2028) & (g2356) & (!g2636) & (!g2640) & (g2843)) + ((g1863) & (g2028) & (g2356) & (!g2636) & (g2640) & (g2843)) + ((g1863) & (g2028) & (g2356) & (g2636) & (!g2640) & (!g2843)) + ((g1863) & (g2028) & (g2356) & (g2636) & (!g2640) & (g2843)) + ((g1863) & (g2028) & (g2356) & (g2636) & (g2640) & (!g2843)) + ((g1863) & (g2028) & (g2356) & (g2636) & (g2640) & (g2843)));
	assign g3094 = (((!sk[13]) & (!g1876) & (g3062) & (!g3084)) + ((!sk[13]) & (!g1876) & (g3062) & (g3084)) + ((!sk[13]) & (g1876) & (!g3062) & (!g3084)) + ((!sk[13]) & (g1876) & (!g3062) & (g3084)) + ((!sk[13]) & (g1876) & (g3062) & (!g3084)) + ((!sk[13]) & (g1876) & (g3062) & (g3084)) + ((sk[13]) & (!g1876) & (!g3062) & (g3084)) + ((sk[13]) & (!g1876) & (g3062) & (g3084)) + ((sk[13]) & (g1876) & (!g3062) & (!g3084)) + ((sk[13]) & (g1876) & (!g3062) & (g3084)) + ((sk[13]) & (g1876) & (g3062) & (g3084)));
	assign g3095 = (((!sk[14]) & (!g1889) & (g3062) & (!g3084)) + ((!sk[14]) & (!g1889) & (g3062) & (g3084)) + ((!sk[14]) & (g1889) & (!g3062) & (!g3084)) + ((!sk[14]) & (g1889) & (!g3062) & (g3084)) + ((!sk[14]) & (g1889) & (g3062) & (!g3084)) + ((!sk[14]) & (g1889) & (g3062) & (g3084)) + ((sk[14]) & (!g1889) & (!g3062) & (g3084)) + ((sk[14]) & (!g1889) & (g3062) & (g3084)) + ((sk[14]) & (g1889) & (!g3062) & (!g3084)) + ((sk[14]) & (g1889) & (!g3062) & (g3084)) + ((sk[14]) & (g1889) & (g3062) & (g3084)));
	assign g3096 = (((!g142) & (!sk[15]) & (g1185) & (!g2675)) + ((!g142) & (!sk[15]) & (g1185) & (g2675)) + ((!g142) & (sk[15]) & (!g1185) & (g2675)) + ((!g142) & (sk[15]) & (g1185) & (!g2675)) + ((g142) & (!sk[15]) & (!g1185) & (!g2675)) + ((g142) & (!sk[15]) & (!g1185) & (g2675)) + ((g142) & (!sk[15]) & (g1185) & (!g2675)) + ((g142) & (!sk[15]) & (g1185) & (g2675)) + ((g142) & (sk[15]) & (!g1185) & (!g2675)) + ((g142) & (sk[15]) & (g1185) & (g2675)));
	assign g3097 = (((!g1889) & (!sk[16]) & (!g2033) & (!g2034) & (g3096) & (!g2677)) + ((!g1889) & (!sk[16]) & (!g2033) & (!g2034) & (g3096) & (g2677)) + ((!g1889) & (!sk[16]) & (!g2033) & (g2034) & (!g3096) & (!g2677)) + ((!g1889) & (!sk[16]) & (!g2033) & (g2034) & (!g3096) & (g2677)) + ((!g1889) & (!sk[16]) & (!g2033) & (g2034) & (g3096) & (!g2677)) + ((!g1889) & (!sk[16]) & (!g2033) & (g2034) & (g3096) & (g2677)) + ((!g1889) & (!sk[16]) & (g2033) & (!g2034) & (g3096) & (!g2677)) + ((!g1889) & (!sk[16]) & (g2033) & (!g2034) & (g3096) & (g2677)) + ((!g1889) & (!sk[16]) & (g2033) & (g2034) & (!g3096) & (!g2677)) + ((!g1889) & (!sk[16]) & (g2033) & (g2034) & (!g3096) & (g2677)) + ((!g1889) & (!sk[16]) & (g2033) & (g2034) & (g3096) & (!g2677)) + ((!g1889) & (!sk[16]) & (g2033) & (g2034) & (g3096) & (g2677)) + ((!g1889) & (sk[16]) & (!g2033) & (!g2034) & (!g3096) & (g2677)) + ((!g1889) & (sk[16]) & (!g2033) & (!g2034) & (g3096) & (g2677)) + ((!g1889) & (sk[16]) & (g2033) & (!g2034) & (g3096) & (!g2677)) + ((!g1889) & (sk[16]) & (g2033) & (!g2034) & (g3096) & (g2677)) + ((g1889) & (!sk[16]) & (!g2033) & (!g2034) & (!g3096) & (!g2677)) + ((g1889) & (!sk[16]) & (!g2033) & (!g2034) & (!g3096) & (g2677)) + ((g1889) & (!sk[16]) & (!g2033) & (!g2034) & (g3096) & (!g2677)) + ((g1889) & (!sk[16]) & (!g2033) & (!g2034) & (g3096) & (g2677)) + ((g1889) & (!sk[16]) & (!g2033) & (g2034) & (!g3096) & (!g2677)) + ((g1889) & (!sk[16]) & (!g2033) & (g2034) & (!g3096) & (g2677)) + ((g1889) & (!sk[16]) & (!g2033) & (g2034) & (g3096) & (!g2677)) + ((g1889) & (!sk[16]) & (!g2033) & (g2034) & (g3096) & (g2677)) + ((g1889) & (!sk[16]) & (g2033) & (!g2034) & (!g3096) & (!g2677)) + ((g1889) & (!sk[16]) & (g2033) & (!g2034) & (!g3096) & (g2677)) + ((g1889) & (!sk[16]) & (g2033) & (!g2034) & (g3096) & (!g2677)) + ((g1889) & (!sk[16]) & (g2033) & (!g2034) & (g3096) & (g2677)) + ((g1889) & (!sk[16]) & (g2033) & (g2034) & (!g3096) & (!g2677)) + ((g1889) & (!sk[16]) & (g2033) & (g2034) & (!g3096) & (g2677)) + ((g1889) & (!sk[16]) & (g2033) & (g2034) & (g3096) & (!g2677)) + ((g1889) & (!sk[16]) & (g2033) & (g2034) & (g3096) & (g2677)) + ((g1889) & (sk[16]) & (!g2033) & (!g2034) & (!g3096) & (g2677)) + ((g1889) & (sk[16]) & (!g2033) & (!g2034) & (g3096) & (g2677)) + ((g1889) & (sk[16]) & (!g2033) & (g2034) & (!g3096) & (!g2677)) + ((g1889) & (sk[16]) & (!g2033) & (g2034) & (!g3096) & (g2677)) + ((g1889) & (sk[16]) & (!g2033) & (g2034) & (g3096) & (!g2677)) + ((g1889) & (sk[16]) & (!g2033) & (g2034) & (g3096) & (g2677)) + ((g1889) & (sk[16]) & (g2033) & (!g2034) & (g3096) & (!g2677)) + ((g1889) & (sk[16]) & (g2033) & (!g2034) & (g3096) & (g2677)));
	assign g3098 = (((!g1889) & (!g2028) & (!g2356) & (g2674) & (!g3097) & (!g2843)) + ((!g1889) & (!g2028) & (!g2356) & (g2674) & (!g3097) & (g2843)) + ((!g1889) & (!g2028) & (!g2356) & (g2674) & (g3097) & (!g2843)) + ((!g1889) & (!g2028) & (!g2356) & (g2674) & (g3097) & (g2843)) + ((!g1889) & (!g2028) & (g2356) & (g2674) & (!g3097) & (!g2843)) + ((!g1889) & (!g2028) & (g2356) & (g2674) & (g3097) & (!g2843)) + ((!g1889) & (g2028) & (!g2356) & (!g2674) & (g3097) & (g2843)) + ((!g1889) & (g2028) & (!g2356) & (g2674) & (!g3097) & (!g2843)) + ((!g1889) & (g2028) & (!g2356) & (g2674) & (g3097) & (!g2843)) + ((!g1889) & (g2028) & (!g2356) & (g2674) & (g3097) & (g2843)) + ((!g1889) & (g2028) & (g2356) & (g2674) & (!g3097) & (!g2843)) + ((!g1889) & (g2028) & (g2356) & (g2674) & (g3097) & (!g2843)) + ((g1889) & (!g2028) & (!g2356) & (g2674) & (!g3097) & (!g2843)) + ((g1889) & (!g2028) & (!g2356) & (g2674) & (!g3097) & (g2843)) + ((g1889) & (!g2028) & (!g2356) & (g2674) & (g3097) & (!g2843)) + ((g1889) & (!g2028) & (!g2356) & (g2674) & (g3097) & (g2843)) + ((g1889) & (!g2028) & (g2356) & (!g2674) & (!g3097) & (g2843)) + ((g1889) & (!g2028) & (g2356) & (!g2674) & (g3097) & (g2843)) + ((g1889) & (!g2028) & (g2356) & (g2674) & (!g3097) & (!g2843)) + ((g1889) & (!g2028) & (g2356) & (g2674) & (!g3097) & (g2843)) + ((g1889) & (!g2028) & (g2356) & (g2674) & (g3097) & (!g2843)) + ((g1889) & (!g2028) & (g2356) & (g2674) & (g3097) & (g2843)) + ((g1889) & (g2028) & (!g2356) & (!g2674) & (g3097) & (g2843)) + ((g1889) & (g2028) & (!g2356) & (g2674) & (!g3097) & (!g2843)) + ((g1889) & (g2028) & (!g2356) & (g2674) & (g3097) & (!g2843)) + ((g1889) & (g2028) & (!g2356) & (g2674) & (g3097) & (g2843)) + ((g1889) & (g2028) & (g2356) & (!g2674) & (!g3097) & (g2843)) + ((g1889) & (g2028) & (g2356) & (!g2674) & (g3097) & (g2843)) + ((g1889) & (g2028) & (g2356) & (g2674) & (!g3097) & (!g2843)) + ((g1889) & (g2028) & (g2356) & (g2674) & (!g3097) & (g2843)) + ((g1889) & (g2028) & (g2356) & (g2674) & (g3097) & (!g2843)) + ((g1889) & (g2028) & (g2356) & (g2674) & (g3097) & (g2843)));
	assign g3099 = (((!g1902) & (!sk[18]) & (g3062) & (!g3084)) + ((!g1902) & (!sk[18]) & (g3062) & (g3084)) + ((!g1902) & (sk[18]) & (!g3062) & (g3084)) + ((!g1902) & (sk[18]) & (g3062) & (g3084)) + ((g1902) & (!sk[18]) & (!g3062) & (!g3084)) + ((g1902) & (!sk[18]) & (!g3062) & (g3084)) + ((g1902) & (!sk[18]) & (g3062) & (!g3084)) + ((g1902) & (!sk[18]) & (g3062) & (g3084)) + ((g1902) & (sk[18]) & (!g3062) & (!g3084)) + ((g1902) & (sk[18]) & (!g3062) & (g3084)) + ((g1902) & (sk[18]) & (g3062) & (g3084)));
	assign g3100 = (((!sk[19]) & (!g1915) & (g3062) & (!g3084)) + ((!sk[19]) & (!g1915) & (g3062) & (g3084)) + ((!sk[19]) & (g1915) & (!g3062) & (!g3084)) + ((!sk[19]) & (g1915) & (!g3062) & (g3084)) + ((!sk[19]) & (g1915) & (g3062) & (!g3084)) + ((!sk[19]) & (g1915) & (g3062) & (g3084)) + ((sk[19]) & (!g1915) & (!g3062) & (g3084)) + ((sk[19]) & (!g1915) & (g3062) & (g3084)) + ((sk[19]) & (g1915) & (!g3062) & (!g3084)) + ((sk[19]) & (g1915) & (!g3062) & (g3084)) + ((sk[19]) & (g1915) & (g3062) & (g3084)));
	assign g3101 = (((!g1915) & (!g2028) & (!g2356) & (g2710) & (!g2713) & (!g2843)) + ((!g1915) & (!g2028) & (!g2356) & (g2710) & (!g2713) & (g2843)) + ((!g1915) & (!g2028) & (!g2356) & (g2710) & (g2713) & (!g2843)) + ((!g1915) & (!g2028) & (!g2356) & (g2710) & (g2713) & (g2843)) + ((!g1915) & (!g2028) & (g2356) & (g2710) & (!g2713) & (!g2843)) + ((!g1915) & (!g2028) & (g2356) & (g2710) & (g2713) & (!g2843)) + ((!g1915) & (g2028) & (!g2356) & (!g2710) & (g2713) & (g2843)) + ((!g1915) & (g2028) & (!g2356) & (g2710) & (!g2713) & (!g2843)) + ((!g1915) & (g2028) & (!g2356) & (g2710) & (g2713) & (!g2843)) + ((!g1915) & (g2028) & (!g2356) & (g2710) & (g2713) & (g2843)) + ((!g1915) & (g2028) & (g2356) & (g2710) & (!g2713) & (!g2843)) + ((!g1915) & (g2028) & (g2356) & (g2710) & (g2713) & (!g2843)) + ((g1915) & (!g2028) & (!g2356) & (g2710) & (!g2713) & (!g2843)) + ((g1915) & (!g2028) & (!g2356) & (g2710) & (!g2713) & (g2843)) + ((g1915) & (!g2028) & (!g2356) & (g2710) & (g2713) & (!g2843)) + ((g1915) & (!g2028) & (!g2356) & (g2710) & (g2713) & (g2843)) + ((g1915) & (!g2028) & (g2356) & (!g2710) & (!g2713) & (g2843)) + ((g1915) & (!g2028) & (g2356) & (!g2710) & (g2713) & (g2843)) + ((g1915) & (!g2028) & (g2356) & (g2710) & (!g2713) & (!g2843)) + ((g1915) & (!g2028) & (g2356) & (g2710) & (!g2713) & (g2843)) + ((g1915) & (!g2028) & (g2356) & (g2710) & (g2713) & (!g2843)) + ((g1915) & (!g2028) & (g2356) & (g2710) & (g2713) & (g2843)) + ((g1915) & (g2028) & (!g2356) & (!g2710) & (g2713) & (g2843)) + ((g1915) & (g2028) & (!g2356) & (g2710) & (!g2713) & (!g2843)) + ((g1915) & (g2028) & (!g2356) & (g2710) & (g2713) & (!g2843)) + ((g1915) & (g2028) & (!g2356) & (g2710) & (g2713) & (g2843)) + ((g1915) & (g2028) & (g2356) & (!g2710) & (!g2713) & (g2843)) + ((g1915) & (g2028) & (g2356) & (!g2710) & (g2713) & (g2843)) + ((g1915) & (g2028) & (g2356) & (g2710) & (!g2713) & (!g2843)) + ((g1915) & (g2028) & (g2356) & (g2710) & (!g2713) & (g2843)) + ((g1915) & (g2028) & (g2356) & (g2710) & (g2713) & (!g2843)) + ((g1915) & (g2028) & (g2356) & (g2710) & (g2713) & (g2843)));
	assign g3102 = (((!g1929) & (!sk[21]) & (g3062) & (!g3084)) + ((!g1929) & (!sk[21]) & (g3062) & (g3084)) + ((!g1929) & (sk[21]) & (!g3062) & (g3084)) + ((!g1929) & (sk[21]) & (g3062) & (g3084)) + ((g1929) & (!sk[21]) & (!g3062) & (!g3084)) + ((g1929) & (!sk[21]) & (!g3062) & (g3084)) + ((g1929) & (!sk[21]) & (g3062) & (!g3084)) + ((g1929) & (!sk[21]) & (g3062) & (g3084)) + ((g1929) & (sk[21]) & (!g3062) & (!g3084)) + ((g1929) & (sk[21]) & (!g3062) & (g3084)) + ((g1929) & (sk[21]) & (g3062) & (g3084)));
	assign g3103 = (((!g1929) & (!g2028) & (!g2356) & (g2728) & (!g2732) & (!g2843)) + ((!g1929) & (!g2028) & (!g2356) & (g2728) & (!g2732) & (g2843)) + ((!g1929) & (!g2028) & (!g2356) & (g2728) & (g2732) & (!g2843)) + ((!g1929) & (!g2028) & (!g2356) & (g2728) & (g2732) & (g2843)) + ((!g1929) & (!g2028) & (g2356) & (g2728) & (!g2732) & (!g2843)) + ((!g1929) & (!g2028) & (g2356) & (g2728) & (g2732) & (!g2843)) + ((!g1929) & (g2028) & (!g2356) & (!g2728) & (g2732) & (g2843)) + ((!g1929) & (g2028) & (!g2356) & (g2728) & (!g2732) & (!g2843)) + ((!g1929) & (g2028) & (!g2356) & (g2728) & (g2732) & (!g2843)) + ((!g1929) & (g2028) & (!g2356) & (g2728) & (g2732) & (g2843)) + ((!g1929) & (g2028) & (g2356) & (g2728) & (!g2732) & (!g2843)) + ((!g1929) & (g2028) & (g2356) & (g2728) & (g2732) & (!g2843)) + ((g1929) & (!g2028) & (!g2356) & (g2728) & (!g2732) & (!g2843)) + ((g1929) & (!g2028) & (!g2356) & (g2728) & (!g2732) & (g2843)) + ((g1929) & (!g2028) & (!g2356) & (g2728) & (g2732) & (!g2843)) + ((g1929) & (!g2028) & (!g2356) & (g2728) & (g2732) & (g2843)) + ((g1929) & (!g2028) & (g2356) & (!g2728) & (!g2732) & (g2843)) + ((g1929) & (!g2028) & (g2356) & (!g2728) & (g2732) & (g2843)) + ((g1929) & (!g2028) & (g2356) & (g2728) & (!g2732) & (!g2843)) + ((g1929) & (!g2028) & (g2356) & (g2728) & (!g2732) & (g2843)) + ((g1929) & (!g2028) & (g2356) & (g2728) & (g2732) & (!g2843)) + ((g1929) & (!g2028) & (g2356) & (g2728) & (g2732) & (g2843)) + ((g1929) & (g2028) & (!g2356) & (!g2728) & (g2732) & (g2843)) + ((g1929) & (g2028) & (!g2356) & (g2728) & (!g2732) & (!g2843)) + ((g1929) & (g2028) & (!g2356) & (g2728) & (g2732) & (!g2843)) + ((g1929) & (g2028) & (!g2356) & (g2728) & (g2732) & (g2843)) + ((g1929) & (g2028) & (g2356) & (!g2728) & (!g2732) & (g2843)) + ((g1929) & (g2028) & (g2356) & (!g2728) & (g2732) & (g2843)) + ((g1929) & (g2028) & (g2356) & (g2728) & (!g2732) & (!g2843)) + ((g1929) & (g2028) & (g2356) & (g2728) & (!g2732) & (g2843)) + ((g1929) & (g2028) & (g2356) & (g2728) & (g2732) & (!g2843)) + ((g1929) & (g2028) & (g2356) & (g2728) & (g2732) & (g2843)));
	assign g3104 = (((!g1942) & (!sk[23]) & (g3062) & (!g3084)) + ((!g1942) & (!sk[23]) & (g3062) & (g3084)) + ((!g1942) & (sk[23]) & (!g3062) & (g3084)) + ((!g1942) & (sk[23]) & (g3062) & (g3084)) + ((g1942) & (!sk[23]) & (!g3062) & (!g3084)) + ((g1942) & (!sk[23]) & (!g3062) & (g3084)) + ((g1942) & (!sk[23]) & (g3062) & (!g3084)) + ((g1942) & (!sk[23]) & (g3062) & (g3084)) + ((g1942) & (sk[23]) & (!g3062) & (!g3084)) + ((g1942) & (sk[23]) & (!g3062) & (g3084)) + ((g1942) & (sk[23]) & (g3062) & (g3084)));
	assign g3105 = (((!g1955) & (!g3062) & (sk[24]) & (g3084)) + ((!g1955) & (g3062) & (!sk[24]) & (!g3084)) + ((!g1955) & (g3062) & (!sk[24]) & (g3084)) + ((!g1955) & (g3062) & (sk[24]) & (g3084)) + ((g1955) & (!g3062) & (!sk[24]) & (!g3084)) + ((g1955) & (!g3062) & (!sk[24]) & (g3084)) + ((g1955) & (!g3062) & (sk[24]) & (!g3084)) + ((g1955) & (!g3062) & (sk[24]) & (g3084)) + ((g1955) & (g3062) & (!sk[24]) & (!g3084)) + ((g1955) & (g3062) & (!sk[24]) & (g3084)) + ((g1955) & (g3062) & (sk[24]) & (g3084)));
	assign g3106 = (((!g1968) & (!g3062) & (sk[25]) & (g3084)) + ((!g1968) & (g3062) & (!sk[25]) & (!g3084)) + ((!g1968) & (g3062) & (!sk[25]) & (g3084)) + ((!g1968) & (g3062) & (sk[25]) & (g3084)) + ((g1968) & (!g3062) & (!sk[25]) & (!g3084)) + ((g1968) & (!g3062) & (!sk[25]) & (g3084)) + ((g1968) & (!g3062) & (sk[25]) & (!g3084)) + ((g1968) & (!g3062) & (sk[25]) & (g3084)) + ((g1968) & (g3062) & (!sk[25]) & (!g3084)) + ((g1968) & (g3062) & (!sk[25]) & (g3084)) + ((g1968) & (g3062) & (sk[25]) & (g3084)));
	assign g3107 = (((!g1968) & (!g2028) & (!g2356) & (g2789) & (!g2792) & (!g2843)) + ((!g1968) & (!g2028) & (!g2356) & (g2789) & (!g2792) & (g2843)) + ((!g1968) & (!g2028) & (!g2356) & (g2789) & (g2792) & (!g2843)) + ((!g1968) & (!g2028) & (!g2356) & (g2789) & (g2792) & (g2843)) + ((!g1968) & (!g2028) & (g2356) & (g2789) & (!g2792) & (!g2843)) + ((!g1968) & (!g2028) & (g2356) & (g2789) & (g2792) & (!g2843)) + ((!g1968) & (g2028) & (!g2356) & (!g2789) & (g2792) & (g2843)) + ((!g1968) & (g2028) & (!g2356) & (g2789) & (!g2792) & (!g2843)) + ((!g1968) & (g2028) & (!g2356) & (g2789) & (g2792) & (!g2843)) + ((!g1968) & (g2028) & (!g2356) & (g2789) & (g2792) & (g2843)) + ((!g1968) & (g2028) & (g2356) & (g2789) & (!g2792) & (!g2843)) + ((!g1968) & (g2028) & (g2356) & (g2789) & (g2792) & (!g2843)) + ((g1968) & (!g2028) & (!g2356) & (g2789) & (!g2792) & (!g2843)) + ((g1968) & (!g2028) & (!g2356) & (g2789) & (!g2792) & (g2843)) + ((g1968) & (!g2028) & (!g2356) & (g2789) & (g2792) & (!g2843)) + ((g1968) & (!g2028) & (!g2356) & (g2789) & (g2792) & (g2843)) + ((g1968) & (!g2028) & (g2356) & (!g2789) & (!g2792) & (g2843)) + ((g1968) & (!g2028) & (g2356) & (!g2789) & (g2792) & (g2843)) + ((g1968) & (!g2028) & (g2356) & (g2789) & (!g2792) & (!g2843)) + ((g1968) & (!g2028) & (g2356) & (g2789) & (!g2792) & (g2843)) + ((g1968) & (!g2028) & (g2356) & (g2789) & (g2792) & (!g2843)) + ((g1968) & (!g2028) & (g2356) & (g2789) & (g2792) & (g2843)) + ((g1968) & (g2028) & (!g2356) & (!g2789) & (g2792) & (g2843)) + ((g1968) & (g2028) & (!g2356) & (g2789) & (!g2792) & (!g2843)) + ((g1968) & (g2028) & (!g2356) & (g2789) & (g2792) & (!g2843)) + ((g1968) & (g2028) & (!g2356) & (g2789) & (g2792) & (g2843)) + ((g1968) & (g2028) & (g2356) & (!g2789) & (!g2792) & (g2843)) + ((g1968) & (g2028) & (g2356) & (!g2789) & (g2792) & (g2843)) + ((g1968) & (g2028) & (g2356) & (g2789) & (!g2792) & (!g2843)) + ((g1968) & (g2028) & (g2356) & (g2789) & (!g2792) & (g2843)) + ((g1968) & (g2028) & (g2356) & (g2789) & (g2792) & (!g2843)) + ((g1968) & (g2028) & (g2356) & (g2789) & (g2792) & (g2843)));
	assign g3108 = (((!g1981) & (!g3062) & (sk[27]) & (g3084)) + ((!g1981) & (g3062) & (!sk[27]) & (!g3084)) + ((!g1981) & (g3062) & (!sk[27]) & (g3084)) + ((!g1981) & (g3062) & (sk[27]) & (g3084)) + ((g1981) & (!g3062) & (!sk[27]) & (!g3084)) + ((g1981) & (!g3062) & (!sk[27]) & (g3084)) + ((g1981) & (!g3062) & (sk[27]) & (!g3084)) + ((g1981) & (!g3062) & (sk[27]) & (g3084)) + ((g1981) & (g3062) & (!sk[27]) & (!g3084)) + ((g1981) & (g3062) & (!sk[27]) & (g3084)) + ((g1981) & (g3062) & (sk[27]) & (g3084)));
	assign g3109 = (((!g1981) & (!g2028) & (!g2356) & (g2806) & (!g2809) & (!g2843)) + ((!g1981) & (!g2028) & (!g2356) & (g2806) & (!g2809) & (g2843)) + ((!g1981) & (!g2028) & (!g2356) & (g2806) & (g2809) & (!g2843)) + ((!g1981) & (!g2028) & (!g2356) & (g2806) & (g2809) & (g2843)) + ((!g1981) & (!g2028) & (g2356) & (g2806) & (!g2809) & (!g2843)) + ((!g1981) & (!g2028) & (g2356) & (g2806) & (g2809) & (!g2843)) + ((!g1981) & (g2028) & (!g2356) & (!g2806) & (g2809) & (g2843)) + ((!g1981) & (g2028) & (!g2356) & (g2806) & (!g2809) & (!g2843)) + ((!g1981) & (g2028) & (!g2356) & (g2806) & (g2809) & (!g2843)) + ((!g1981) & (g2028) & (!g2356) & (g2806) & (g2809) & (g2843)) + ((!g1981) & (g2028) & (g2356) & (g2806) & (!g2809) & (!g2843)) + ((!g1981) & (g2028) & (g2356) & (g2806) & (g2809) & (!g2843)) + ((g1981) & (!g2028) & (!g2356) & (g2806) & (!g2809) & (!g2843)) + ((g1981) & (!g2028) & (!g2356) & (g2806) & (!g2809) & (g2843)) + ((g1981) & (!g2028) & (!g2356) & (g2806) & (g2809) & (!g2843)) + ((g1981) & (!g2028) & (!g2356) & (g2806) & (g2809) & (g2843)) + ((g1981) & (!g2028) & (g2356) & (!g2806) & (!g2809) & (g2843)) + ((g1981) & (!g2028) & (g2356) & (!g2806) & (g2809) & (g2843)) + ((g1981) & (!g2028) & (g2356) & (g2806) & (!g2809) & (!g2843)) + ((g1981) & (!g2028) & (g2356) & (g2806) & (!g2809) & (g2843)) + ((g1981) & (!g2028) & (g2356) & (g2806) & (g2809) & (!g2843)) + ((g1981) & (!g2028) & (g2356) & (g2806) & (g2809) & (g2843)) + ((g1981) & (g2028) & (!g2356) & (!g2806) & (g2809) & (g2843)) + ((g1981) & (g2028) & (!g2356) & (g2806) & (!g2809) & (!g2843)) + ((g1981) & (g2028) & (!g2356) & (g2806) & (g2809) & (!g2843)) + ((g1981) & (g2028) & (!g2356) & (g2806) & (g2809) & (g2843)) + ((g1981) & (g2028) & (g2356) & (!g2806) & (!g2809) & (g2843)) + ((g1981) & (g2028) & (g2356) & (!g2806) & (g2809) & (g2843)) + ((g1981) & (g2028) & (g2356) & (g2806) & (!g2809) & (!g2843)) + ((g1981) & (g2028) & (g2356) & (g2806) & (!g2809) & (g2843)) + ((g1981) & (g2028) & (g2356) & (g2806) & (g2809) & (!g2843)) + ((g1981) & (g2028) & (g2356) & (g2806) & (g2809) & (g2843)));
	assign g3110 = (((!g1994) & (!sk[29]) & (g3062) & (!g3084)) + ((!g1994) & (!sk[29]) & (g3062) & (g3084)) + ((!g1994) & (sk[29]) & (!g3062) & (g3084)) + ((!g1994) & (sk[29]) & (g3062) & (g3084)) + ((g1994) & (!sk[29]) & (!g3062) & (!g3084)) + ((g1994) & (!sk[29]) & (!g3062) & (g3084)) + ((g1994) & (!sk[29]) & (g3062) & (!g3084)) + ((g1994) & (!sk[29]) & (g3062) & (g3084)) + ((g1994) & (sk[29]) & (!g3062) & (!g3084)) + ((g1994) & (sk[29]) & (!g3062) & (g3084)) + ((g1994) & (sk[29]) & (g3062) & (g3084)));
	assign g3111 = (((!g1994) & (!g2028) & (!g2356) & (g2822) & (!g3252) & (!g2843)) + ((!g1994) & (!g2028) & (!g2356) & (g2822) & (!g3252) & (g2843)) + ((!g1994) & (!g2028) & (!g2356) & (g2822) & (g3252) & (!g2843)) + ((!g1994) & (!g2028) & (!g2356) & (g2822) & (g3252) & (g2843)) + ((!g1994) & (!g2028) & (g2356) & (g2822) & (!g3252) & (!g2843)) + ((!g1994) & (!g2028) & (g2356) & (g2822) & (g3252) & (!g2843)) + ((!g1994) & (g2028) & (!g2356) & (!g2822) & (g3252) & (g2843)) + ((!g1994) & (g2028) & (!g2356) & (g2822) & (!g3252) & (!g2843)) + ((!g1994) & (g2028) & (!g2356) & (g2822) & (g3252) & (!g2843)) + ((!g1994) & (g2028) & (!g2356) & (g2822) & (g3252) & (g2843)) + ((!g1994) & (g2028) & (g2356) & (g2822) & (!g3252) & (!g2843)) + ((!g1994) & (g2028) & (g2356) & (g2822) & (g3252) & (!g2843)) + ((g1994) & (!g2028) & (!g2356) & (g2822) & (!g3252) & (!g2843)) + ((g1994) & (!g2028) & (!g2356) & (g2822) & (!g3252) & (g2843)) + ((g1994) & (!g2028) & (!g2356) & (g2822) & (g3252) & (!g2843)) + ((g1994) & (!g2028) & (!g2356) & (g2822) & (g3252) & (g2843)) + ((g1994) & (!g2028) & (g2356) & (!g2822) & (!g3252) & (g2843)) + ((g1994) & (!g2028) & (g2356) & (!g2822) & (g3252) & (g2843)) + ((g1994) & (!g2028) & (g2356) & (g2822) & (!g3252) & (!g2843)) + ((g1994) & (!g2028) & (g2356) & (g2822) & (!g3252) & (g2843)) + ((g1994) & (!g2028) & (g2356) & (g2822) & (g3252) & (!g2843)) + ((g1994) & (!g2028) & (g2356) & (g2822) & (g3252) & (g2843)) + ((g1994) & (g2028) & (!g2356) & (!g2822) & (g3252) & (g2843)) + ((g1994) & (g2028) & (!g2356) & (g2822) & (!g3252) & (!g2843)) + ((g1994) & (g2028) & (!g2356) & (g2822) & (g3252) & (!g2843)) + ((g1994) & (g2028) & (!g2356) & (g2822) & (g3252) & (g2843)) + ((g1994) & (g2028) & (g2356) & (!g2822) & (!g3252) & (g2843)) + ((g1994) & (g2028) & (g2356) & (!g2822) & (g3252) & (g2843)) + ((g1994) & (g2028) & (g2356) & (g2822) & (!g3252) & (!g2843)) + ((g1994) & (g2028) & (g2356) & (g2822) & (!g3252) & (g2843)) + ((g1994) & (g2028) & (g2356) & (g2822) & (g3252) & (!g2843)) + ((g1994) & (g2028) & (g2356) & (g2822) & (g3252) & (g2843)));
	assign g3112 = (((!g2007) & (!g2028) & (!g2356) & (g2826) & (!g2829) & (!g2843)) + ((!g2007) & (!g2028) & (!g2356) & (g2826) & (!g2829) & (g2843)) + ((!g2007) & (!g2028) & (!g2356) & (g2826) & (g2829) & (!g2843)) + ((!g2007) & (!g2028) & (!g2356) & (g2826) & (g2829) & (g2843)) + ((!g2007) & (!g2028) & (g2356) & (g2826) & (!g2829) & (!g2843)) + ((!g2007) & (!g2028) & (g2356) & (g2826) & (g2829) & (!g2843)) + ((!g2007) & (g2028) & (!g2356) & (!g2826) & (!g2829) & (g2843)) + ((!g2007) & (g2028) & (!g2356) & (g2826) & (!g2829) & (!g2843)) + ((!g2007) & (g2028) & (!g2356) & (g2826) & (!g2829) & (g2843)) + ((!g2007) & (g2028) & (!g2356) & (g2826) & (g2829) & (!g2843)) + ((!g2007) & (g2028) & (g2356) & (g2826) & (!g2829) & (!g2843)) + ((!g2007) & (g2028) & (g2356) & (g2826) & (g2829) & (!g2843)) + ((g2007) & (!g2028) & (!g2356) & (g2826) & (!g2829) & (!g2843)) + ((g2007) & (!g2028) & (!g2356) & (g2826) & (!g2829) & (g2843)) + ((g2007) & (!g2028) & (!g2356) & (g2826) & (g2829) & (!g2843)) + ((g2007) & (!g2028) & (!g2356) & (g2826) & (g2829) & (g2843)) + ((g2007) & (!g2028) & (g2356) & (!g2826) & (!g2829) & (g2843)) + ((g2007) & (!g2028) & (g2356) & (!g2826) & (g2829) & (g2843)) + ((g2007) & (!g2028) & (g2356) & (g2826) & (!g2829) & (!g2843)) + ((g2007) & (!g2028) & (g2356) & (g2826) & (!g2829) & (g2843)) + ((g2007) & (!g2028) & (g2356) & (g2826) & (g2829) & (!g2843)) + ((g2007) & (!g2028) & (g2356) & (g2826) & (g2829) & (g2843)) + ((g2007) & (g2028) & (!g2356) & (!g2826) & (!g2829) & (g2843)) + ((g2007) & (g2028) & (!g2356) & (g2826) & (!g2829) & (!g2843)) + ((g2007) & (g2028) & (!g2356) & (g2826) & (!g2829) & (g2843)) + ((g2007) & (g2028) & (!g2356) & (g2826) & (g2829) & (!g2843)) + ((g2007) & (g2028) & (g2356) & (!g2826) & (!g2829) & (g2843)) + ((g2007) & (g2028) & (g2356) & (!g2826) & (g2829) & (g2843)) + ((g2007) & (g2028) & (g2356) & (g2826) & (!g2829) & (!g2843)) + ((g2007) & (g2028) & (g2356) & (g2826) & (!g2829) & (g2843)) + ((g2007) & (g2028) & (g2356) & (g2826) & (g2829) & (!g2843)) + ((g2007) & (g2028) & (g2356) & (g2826) & (g2829) & (g2843)));
	assign g3113 = (((!g2007) & (!g3062) & (sk[32]) & (g3084)) + ((!g2007) & (g3062) & (!sk[32]) & (!g3084)) + ((!g2007) & (g3062) & (!sk[32]) & (g3084)) + ((!g2007) & (g3062) & (sk[32]) & (g3084)) + ((g2007) & (!g3062) & (!sk[32]) & (!g3084)) + ((g2007) & (!g3062) & (!sk[32]) & (g3084)) + ((g2007) & (!g3062) & (sk[32]) & (!g3084)) + ((g2007) & (!g3062) & (sk[32]) & (g3084)) + ((g2007) & (g3062) & (!sk[32]) & (!g3084)) + ((g2007) & (g3062) & (!sk[32]) & (g3084)) + ((g2007) & (g3062) & (sk[32]) & (g3084)));
	assign g3114 = (((!sk[33]) & (!g1720) & (g2919) & (!g2916)) + ((!sk[33]) & (!g1720) & (g2919) & (g2916)) + ((!sk[33]) & (g1720) & (!g2919) & (!g2916)) + ((!sk[33]) & (g1720) & (!g2919) & (g2916)) + ((!sk[33]) & (g1720) & (g2919) & (!g2916)) + ((!sk[33]) & (g1720) & (g2919) & (g2916)) + ((sk[33]) & (!g1720) & (!g2919) & (!g2916)) + ((sk[33]) & (g1720) & (!g2919) & (!g2916)) + ((sk[33]) & (g1720) & (g2919) & (!g2916)) + ((sk[33]) & (g1720) & (g2919) & (g2916)));
	assign g3115 = (((!g2030) & (!g1733) & (!g2913) & (!g2919) & (!g2969) & (g2971)) + ((!g2030) & (!g1733) & (!g2913) & (!g2919) & (g2969) & (g2971)) + ((!g2030) & (g1733) & (!g2913) & (!g2919) & (!g2969) & (g2971)) + ((!g2030) & (g1733) & (!g2913) & (!g2919) & (g2969) & (g2971)) + ((!g2030) & (g1733) & (!g2913) & (g2919) & (!g2969) & (!g2971)) + ((!g2030) & (g1733) & (!g2913) & (g2919) & (!g2969) & (g2971)) + ((!g2030) & (g1733) & (!g2913) & (g2919) & (g2969) & (!g2971)) + ((!g2030) & (g1733) & (!g2913) & (g2919) & (g2969) & (g2971)) + ((!g2030) & (g1733) & (g2913) & (!g2919) & (!g2969) & (!g2971)) + ((!g2030) & (g1733) & (g2913) & (!g2919) & (!g2969) & (g2971)) + ((!g2030) & (g1733) & (g2913) & (!g2919) & (g2969) & (!g2971)) + ((!g2030) & (g1733) & (g2913) & (!g2919) & (g2969) & (g2971)) + ((!g2030) & (g1733) & (g2913) & (g2919) & (!g2969) & (!g2971)) + ((!g2030) & (g1733) & (g2913) & (g2919) & (!g2969) & (g2971)) + ((!g2030) & (g1733) & (g2913) & (g2919) & (g2969) & (!g2971)) + ((!g2030) & (g1733) & (g2913) & (g2919) & (g2969) & (g2971)) + ((g2030) & (!g1733) & (!g2913) & (!g2919) & (g2969) & (!g2971)) + ((g2030) & (!g1733) & (!g2913) & (!g2919) & (g2969) & (g2971)) + ((g2030) & (!g1733) & (g2913) & (!g2919) & (g2969) & (!g2971)) + ((g2030) & (!g1733) & (g2913) & (!g2919) & (g2969) & (g2971)) + ((g2030) & (g1733) & (!g2913) & (!g2919) & (g2969) & (!g2971)) + ((g2030) & (g1733) & (!g2913) & (!g2919) & (g2969) & (g2971)) + ((g2030) & (g1733) & (!g2913) & (g2919) & (!g2969) & (!g2971)) + ((g2030) & (g1733) & (!g2913) & (g2919) & (!g2969) & (g2971)) + ((g2030) & (g1733) & (!g2913) & (g2919) & (g2969) & (!g2971)) + ((g2030) & (g1733) & (!g2913) & (g2919) & (g2969) & (g2971)) + ((g2030) & (g1733) & (g2913) & (!g2919) & (g2969) & (!g2971)) + ((g2030) & (g1733) & (g2913) & (!g2919) & (g2969) & (g2971)) + ((g2030) & (g1733) & (g2913) & (g2919) & (!g2969) & (!g2971)) + ((g2030) & (g1733) & (g2913) & (g2919) & (!g2969) & (g2971)) + ((g2030) & (g1733) & (g2913) & (g2919) & (g2969) & (!g2971)) + ((g2030) & (g1733) & (g2913) & (g2919) & (g2969) & (g2971)));
	assign g3116 = (((!g2081) & (!g2798) & (!g2799) & (!sk[35]) & (g2099) & (!g2794)) + ((!g2081) & (!g2798) & (!g2799) & (!sk[35]) & (g2099) & (g2794)) + ((!g2081) & (!g2798) & (!g2799) & (sk[35]) & (!g2099) & (!g2794)) + ((!g2081) & (!g2798) & (!g2799) & (sk[35]) & (!g2099) & (g2794)) + ((!g2081) & (!g2798) & (!g2799) & (sk[35]) & (g2099) & (!g2794)) + ((!g2081) & (!g2798) & (!g2799) & (sk[35]) & (g2099) & (g2794)) + ((!g2081) & (!g2798) & (g2799) & (!sk[35]) & (!g2099) & (!g2794)) + ((!g2081) & (!g2798) & (g2799) & (!sk[35]) & (!g2099) & (g2794)) + ((!g2081) & (!g2798) & (g2799) & (!sk[35]) & (g2099) & (!g2794)) + ((!g2081) & (!g2798) & (g2799) & (!sk[35]) & (g2099) & (g2794)) + ((!g2081) & (g2798) & (!g2799) & (!sk[35]) & (g2099) & (!g2794)) + ((!g2081) & (g2798) & (!g2799) & (!sk[35]) & (g2099) & (g2794)) + ((!g2081) & (g2798) & (g2799) & (!sk[35]) & (!g2099) & (!g2794)) + ((!g2081) & (g2798) & (g2799) & (!sk[35]) & (!g2099) & (g2794)) + ((!g2081) & (g2798) & (g2799) & (!sk[35]) & (g2099) & (!g2794)) + ((!g2081) & (g2798) & (g2799) & (!sk[35]) & (g2099) & (g2794)) + ((!g2081) & (g2798) & (g2799) & (sk[35]) & (!g2099) & (!g2794)) + ((!g2081) & (g2798) & (g2799) & (sk[35]) & (!g2099) & (g2794)) + ((!g2081) & (g2798) & (g2799) & (sk[35]) & (g2099) & (!g2794)) + ((!g2081) & (g2798) & (g2799) & (sk[35]) & (g2099) & (g2794)) + ((g2081) & (!g2798) & (!g2799) & (!sk[35]) & (!g2099) & (!g2794)) + ((g2081) & (!g2798) & (!g2799) & (!sk[35]) & (!g2099) & (g2794)) + ((g2081) & (!g2798) & (!g2799) & (!sk[35]) & (g2099) & (!g2794)) + ((g2081) & (!g2798) & (!g2799) & (!sk[35]) & (g2099) & (g2794)) + ((g2081) & (!g2798) & (!g2799) & (sk[35]) & (g2099) & (g2794)) + ((g2081) & (!g2798) & (g2799) & (!sk[35]) & (!g2099) & (!g2794)) + ((g2081) & (!g2798) & (g2799) & (!sk[35]) & (!g2099) & (g2794)) + ((g2081) & (!g2798) & (g2799) & (!sk[35]) & (g2099) & (!g2794)) + ((g2081) & (!g2798) & (g2799) & (!sk[35]) & (g2099) & (g2794)) + ((g2081) & (!g2798) & (g2799) & (sk[35]) & (g2099) & (g2794)) + ((g2081) & (g2798) & (!g2799) & (!sk[35]) & (!g2099) & (!g2794)) + ((g2081) & (g2798) & (!g2799) & (!sk[35]) & (!g2099) & (g2794)) + ((g2081) & (g2798) & (!g2799) & (!sk[35]) & (g2099) & (!g2794)) + ((g2081) & (g2798) & (!g2799) & (!sk[35]) & (g2099) & (g2794)) + ((g2081) & (g2798) & (!g2799) & (sk[35]) & (g2099) & (g2794)) + ((g2081) & (g2798) & (g2799) & (!sk[35]) & (!g2099) & (!g2794)) + ((g2081) & (g2798) & (g2799) & (!sk[35]) & (!g2099) & (g2794)) + ((g2081) & (g2798) & (g2799) & (!sk[35]) & (g2099) & (!g2794)) + ((g2081) & (g2798) & (g2799) & (!sk[35]) & (g2099) & (g2794)) + ((g2081) & (g2798) & (g2799) & (sk[35]) & (g2099) & (g2794)));
	assign g3117 = (((!g87) & (g88) & (!sk[36]) & (!g89)) + ((!g87) & (g88) & (!sk[36]) & (g89)) + ((!g87) & (g88) & (sk[36]) & (!g89)) + ((g87) & (!g88) & (!sk[36]) & (!g89)) + ((g87) & (!g88) & (!sk[36]) & (g89)) + ((g87) & (!g88) & (sk[36]) & (g89)) + ((g87) & (g88) & (!sk[36]) & (!g89)) + ((g87) & (g88) & (!sk[36]) & (g89)) + ((g87) & (g88) & (sk[36]) & (!g89)) + ((g87) & (g88) & (sk[36]) & (g89)));
	assign g3118 = (((!g126) & (g1500) & (!sk[37]) & (!g1454)) + ((!g126) & (g1500) & (!sk[37]) & (g1454)) + ((!g126) & (g1500) & (sk[37]) & (!g1454)) + ((!g126) & (g1500) & (sk[37]) & (g1454)) + ((g126) & (!g1500) & (!sk[37]) & (!g1454)) + ((g126) & (!g1500) & (!sk[37]) & (g1454)) + ((g126) & (!g1500) & (sk[37]) & (!g1454)) + ((g126) & (g1500) & (!sk[37]) & (!g1454)) + ((g126) & (g1500) & (!sk[37]) & (g1454)) + ((g126) & (g1500) & (sk[37]) & (!g1454)));
	assign g3119 = (((!g2121) & (!sk[38]) & (g2529)) + ((!g2121) & (sk[38]) & (!g2529)) + ((g2121) & (!sk[38]) & (g2529)) + ((g2121) & (sk[38]) & (g2529)));
	assign g3120 = (((!g2081) & (!g2101) & (!g2831) & (!g2100) & (!g2811) & (!g2832)) + ((!g2081) & (!g2101) & (!g2831) & (!g2100) & (!g2811) & (g2832)) + ((!g2081) & (!g2101) & (!g2831) & (!g2100) & (g2811) & (!g2832)) + ((!g2081) & (!g2101) & (!g2831) & (!g2100) & (g2811) & (g2832)) + ((!g2081) & (!g2101) & (!g2831) & (g2100) & (!g2811) & (!g2832)) + ((!g2081) & (!g2101) & (!g2831) & (g2100) & (!g2811) & (g2832)) + ((!g2081) & (!g2101) & (!g2831) & (g2100) & (g2811) & (!g2832)) + ((!g2081) & (!g2101) & (!g2831) & (g2100) & (g2811) & (g2832)) + ((!g2081) & (!g2101) & (g2831) & (!g2100) & (!g2811) & (!g2832)) + ((!g2081) & (!g2101) & (g2831) & (!g2100) & (!g2811) & (g2832)) + ((!g2081) & (!g2101) & (g2831) & (!g2100) & (g2811) & (!g2832)) + ((!g2081) & (!g2101) & (g2831) & (g2100) & (!g2811) & (!g2832)) + ((!g2081) & (g2101) & (!g2831) & (!g2100) & (!g2811) & (!g2832)) + ((!g2081) & (g2101) & (!g2831) & (!g2100) & (!g2811) & (g2832)) + ((!g2081) & (g2101) & (!g2831) & (!g2100) & (g2811) & (!g2832)) + ((!g2081) & (g2101) & (!g2831) & (g2100) & (!g2811) & (!g2832)) + ((g2081) & (!g2101) & (!g2831) & (!g2100) & (!g2811) & (!g2832)) + ((g2081) & (!g2101) & (!g2831) & (!g2100) & (!g2811) & (g2832)) + ((g2081) & (!g2101) & (!g2831) & (!g2100) & (g2811) & (!g2832)) + ((g2081) & (!g2101) & (!g2831) & (g2100) & (!g2811) & (!g2832)) + ((g2081) & (g2101) & (g2831) & (!g2100) & (g2811) & (g2832)) + ((g2081) & (g2101) & (g2831) & (g2100) & (!g2811) & (g2832)) + ((g2081) & (g2101) & (g2831) & (g2100) & (g2811) & (!g2832)) + ((g2081) & (g2101) & (g2831) & (g2100) & (g2811) & (g2832)));
	assign g3121 = (((!g2101) & (!sk[40]) & (!g2831) & (!g2100) & (g2811) & (!g2832)) + ((!g2101) & (!sk[40]) & (!g2831) & (!g2100) & (g2811) & (g2832)) + ((!g2101) & (!sk[40]) & (!g2831) & (g2100) & (!g2811) & (!g2832)) + ((!g2101) & (!sk[40]) & (!g2831) & (g2100) & (!g2811) & (g2832)) + ((!g2101) & (!sk[40]) & (!g2831) & (g2100) & (g2811) & (!g2832)) + ((!g2101) & (!sk[40]) & (!g2831) & (g2100) & (g2811) & (g2832)) + ((!g2101) & (!sk[40]) & (g2831) & (!g2100) & (g2811) & (!g2832)) + ((!g2101) & (!sk[40]) & (g2831) & (!g2100) & (g2811) & (g2832)) + ((!g2101) & (!sk[40]) & (g2831) & (g2100) & (!g2811) & (!g2832)) + ((!g2101) & (!sk[40]) & (g2831) & (g2100) & (!g2811) & (g2832)) + ((!g2101) & (!sk[40]) & (g2831) & (g2100) & (g2811) & (!g2832)) + ((!g2101) & (!sk[40]) & (g2831) & (g2100) & (g2811) & (g2832)) + ((!g2101) & (sk[40]) & (g2831) & (!g2100) & (g2811) & (g2832)) + ((!g2101) & (sk[40]) & (g2831) & (g2100) & (!g2811) & (g2832)) + ((!g2101) & (sk[40]) & (g2831) & (g2100) & (g2811) & (!g2832)) + ((!g2101) & (sk[40]) & (g2831) & (g2100) & (g2811) & (g2832)) + ((g2101) & (!sk[40]) & (!g2831) & (!g2100) & (!g2811) & (!g2832)) + ((g2101) & (!sk[40]) & (!g2831) & (!g2100) & (!g2811) & (g2832)) + ((g2101) & (!sk[40]) & (!g2831) & (!g2100) & (g2811) & (!g2832)) + ((g2101) & (!sk[40]) & (!g2831) & (!g2100) & (g2811) & (g2832)) + ((g2101) & (!sk[40]) & (!g2831) & (g2100) & (!g2811) & (!g2832)) + ((g2101) & (!sk[40]) & (!g2831) & (g2100) & (!g2811) & (g2832)) + ((g2101) & (!sk[40]) & (!g2831) & (g2100) & (g2811) & (!g2832)) + ((g2101) & (!sk[40]) & (!g2831) & (g2100) & (g2811) & (g2832)) + ((g2101) & (!sk[40]) & (g2831) & (!g2100) & (!g2811) & (!g2832)) + ((g2101) & (!sk[40]) & (g2831) & (!g2100) & (!g2811) & (g2832)) + ((g2101) & (!sk[40]) & (g2831) & (!g2100) & (g2811) & (!g2832)) + ((g2101) & (!sk[40]) & (g2831) & (!g2100) & (g2811) & (g2832)) + ((g2101) & (!sk[40]) & (g2831) & (g2100) & (!g2811) & (!g2832)) + ((g2101) & (!sk[40]) & (g2831) & (g2100) & (!g2811) & (g2832)) + ((g2101) & (!sk[40]) & (g2831) & (g2100) & (g2811) & (!g2832)) + ((g2101) & (!sk[40]) & (g2831) & (g2100) & (g2811) & (g2832)) + ((g2101) & (sk[40]) & (!g2831) & (!g2100) & (g2811) & (g2832)) + ((g2101) & (sk[40]) & (!g2831) & (g2100) & (!g2811) & (g2832)) + ((g2101) & (sk[40]) & (!g2831) & (g2100) & (g2811) & (!g2832)) + ((g2101) & (sk[40]) & (!g2831) & (g2100) & (g2811) & (g2832)) + ((g2101) & (sk[40]) & (g2831) & (!g2100) & (!g2811) & (!g2832)) + ((g2101) & (sk[40]) & (g2831) & (!g2100) & (!g2811) & (g2832)) + ((g2101) & (sk[40]) & (g2831) & (!g2100) & (g2811) & (!g2832)) + ((g2101) & (sk[40]) & (g2831) & (!g2100) & (g2811) & (g2832)) + ((g2101) & (sk[40]) & (g2831) & (g2100) & (!g2811) & (!g2832)) + ((g2101) & (sk[40]) & (g2831) & (g2100) & (!g2811) & (g2832)) + ((g2101) & (sk[40]) & (g2831) & (g2100) & (g2811) & (!g2832)) + ((g2101) & (sk[40]) & (g2831) & (g2100) & (g2811) & (g2832)));
	assign g3122 = (((!sk[41]) & (!g1733) & (!g2913) & (!g2080) & (g2124) & (!g2125)) + ((!sk[41]) & (!g1733) & (!g2913) & (!g2080) & (g2124) & (g2125)) + ((!sk[41]) & (!g1733) & (!g2913) & (g2080) & (!g2124) & (!g2125)) + ((!sk[41]) & (!g1733) & (!g2913) & (g2080) & (!g2124) & (g2125)) + ((!sk[41]) & (!g1733) & (!g2913) & (g2080) & (g2124) & (!g2125)) + ((!sk[41]) & (!g1733) & (!g2913) & (g2080) & (g2124) & (g2125)) + ((!sk[41]) & (!g1733) & (g2913) & (!g2080) & (g2124) & (!g2125)) + ((!sk[41]) & (!g1733) & (g2913) & (!g2080) & (g2124) & (g2125)) + ((!sk[41]) & (!g1733) & (g2913) & (g2080) & (!g2124) & (!g2125)) + ((!sk[41]) & (!g1733) & (g2913) & (g2080) & (!g2124) & (g2125)) + ((!sk[41]) & (!g1733) & (g2913) & (g2080) & (g2124) & (!g2125)) + ((!sk[41]) & (!g1733) & (g2913) & (g2080) & (g2124) & (g2125)) + ((!sk[41]) & (g1733) & (!g2913) & (!g2080) & (!g2124) & (!g2125)) + ((!sk[41]) & (g1733) & (!g2913) & (!g2080) & (!g2124) & (g2125)) + ((!sk[41]) & (g1733) & (!g2913) & (!g2080) & (g2124) & (!g2125)) + ((!sk[41]) & (g1733) & (!g2913) & (!g2080) & (g2124) & (g2125)) + ((!sk[41]) & (g1733) & (!g2913) & (g2080) & (!g2124) & (!g2125)) + ((!sk[41]) & (g1733) & (!g2913) & (g2080) & (!g2124) & (g2125)) + ((!sk[41]) & (g1733) & (!g2913) & (g2080) & (g2124) & (!g2125)) + ((!sk[41]) & (g1733) & (!g2913) & (g2080) & (g2124) & (g2125)) + ((!sk[41]) & (g1733) & (g2913) & (!g2080) & (!g2124) & (!g2125)) + ((!sk[41]) & (g1733) & (g2913) & (!g2080) & (!g2124) & (g2125)) + ((!sk[41]) & (g1733) & (g2913) & (!g2080) & (g2124) & (!g2125)) + ((!sk[41]) & (g1733) & (g2913) & (!g2080) & (g2124) & (g2125)) + ((!sk[41]) & (g1733) & (g2913) & (g2080) & (!g2124) & (!g2125)) + ((!sk[41]) & (g1733) & (g2913) & (g2080) & (!g2124) & (g2125)) + ((!sk[41]) & (g1733) & (g2913) & (g2080) & (g2124) & (!g2125)) + ((!sk[41]) & (g1733) & (g2913) & (g2080) & (g2124) & (g2125)) + ((sk[41]) & (!g1733) & (!g2913) & (g2080) & (!g2124) & (!g2125)) + ((sk[41]) & (g1733) & (!g2913) & (g2080) & (!g2124) & (!g2125)) + ((sk[41]) & (g1733) & (g2913) & (!g2080) & (!g2124) & (!g2125)) + ((sk[41]) & (g1733) & (g2913) & (!g2080) & (!g2124) & (g2125)) + ((sk[41]) & (g1733) & (g2913) & (!g2080) & (g2124) & (!g2125)) + ((sk[41]) & (g1733) & (g2913) & (!g2080) & (g2124) & (g2125)) + ((sk[41]) & (g1733) & (g2913) & (g2080) & (!g2124) & (!g2125)) + ((sk[41]) & (g1733) & (g2913) & (g2080) & (!g2124) & (g2125)) + ((sk[41]) & (g1733) & (g2913) & (g2080) & (g2124) & (!g2125)) + ((sk[41]) & (g1733) & (g2913) & (g2080) & (g2124) & (g2125)));
	assign g3123 = (((!g2383) & (!g2914) & (!sk[42]) & (!g3017) & (g3018)) + ((!g2383) & (!g2914) & (!sk[42]) & (g3017) & (g3018)) + ((!g2383) & (!g2914) & (sk[42]) & (g3017) & (!g3018)) + ((!g2383) & (g2914) & (!sk[42]) & (!g3017) & (!g3018)) + ((!g2383) & (g2914) & (!sk[42]) & (!g3017) & (g3018)) + ((!g2383) & (g2914) & (!sk[42]) & (g3017) & (!g3018)) + ((!g2383) & (g2914) & (!sk[42]) & (g3017) & (g3018)) + ((!g2383) & (g2914) & (sk[42]) & (!g3017) & (!g3018)) + ((!g2383) & (g2914) & (sk[42]) & (g3017) & (!g3018)) + ((g2383) & (!g2914) & (!sk[42]) & (!g3017) & (!g3018)) + ((g2383) & (!g2914) & (!sk[42]) & (!g3017) & (g3018)) + ((g2383) & (!g2914) & (!sk[42]) & (g3017) & (!g3018)) + ((g2383) & (!g2914) & (!sk[42]) & (g3017) & (g3018)) + ((g2383) & (!g2914) & (sk[42]) & (!g3017) & (g3018)) + ((g2383) & (!g2914) & (sk[42]) & (g3017) & (!g3018)) + ((g2383) & (g2914) & (!sk[42]) & (!g3017) & (!g3018)) + ((g2383) & (g2914) & (!sk[42]) & (!g3017) & (g3018)) + ((g2383) & (g2914) & (!sk[42]) & (g3017) & (!g3018)) + ((g2383) & (g2914) & (!sk[42]) & (g3017) & (g3018)) + ((g2383) & (g2914) & (sk[42]) & (!g3017) & (!g3018)) + ((g2383) & (g2914) & (sk[42]) & (!g3017) & (g3018)) + ((g2383) & (g2914) & (sk[42]) & (g3017) & (!g3018)));
	assign g3124 = (((!g2977) & (!g142) & (!sk[43]) & (!g563) & (g583) & (!g3123)) + ((!g2977) & (!g142) & (!sk[43]) & (!g563) & (g583) & (g3123)) + ((!g2977) & (!g142) & (!sk[43]) & (g563) & (!g583) & (!g3123)) + ((!g2977) & (!g142) & (!sk[43]) & (g563) & (!g583) & (g3123)) + ((!g2977) & (!g142) & (!sk[43]) & (g563) & (g583) & (!g3123)) + ((!g2977) & (!g142) & (!sk[43]) & (g563) & (g583) & (g3123)) + ((!g2977) & (!g142) & (sk[43]) & (!g563) & (g583) & (!g3123)) + ((!g2977) & (!g142) & (sk[43]) & (!g563) & (g583) & (g3123)) + ((!g2977) & (!g142) & (sk[43]) & (g563) & (g583) & (!g3123)) + ((!g2977) & (!g142) & (sk[43]) & (g563) & (g583) & (g3123)) + ((!g2977) & (g142) & (!sk[43]) & (!g563) & (g583) & (!g3123)) + ((!g2977) & (g142) & (!sk[43]) & (!g563) & (g583) & (g3123)) + ((!g2977) & (g142) & (!sk[43]) & (g563) & (!g583) & (!g3123)) + ((!g2977) & (g142) & (!sk[43]) & (g563) & (!g583) & (g3123)) + ((!g2977) & (g142) & (!sk[43]) & (g563) & (g583) & (!g3123)) + ((!g2977) & (g142) & (!sk[43]) & (g563) & (g583) & (g3123)) + ((!g2977) & (g142) & (sk[43]) & (g563) & (!g583) & (!g3123)) + ((!g2977) & (g142) & (sk[43]) & (g563) & (!g583) & (g3123)) + ((!g2977) & (g142) & (sk[43]) & (g563) & (g583) & (!g3123)) + ((!g2977) & (g142) & (sk[43]) & (g563) & (g583) & (g3123)) + ((g2977) & (!g142) & (!sk[43]) & (!g563) & (!g583) & (!g3123)) + ((g2977) & (!g142) & (!sk[43]) & (!g563) & (!g583) & (g3123)) + ((g2977) & (!g142) & (!sk[43]) & (!g563) & (g583) & (!g3123)) + ((g2977) & (!g142) & (!sk[43]) & (!g563) & (g583) & (g3123)) + ((g2977) & (!g142) & (!sk[43]) & (g563) & (!g583) & (!g3123)) + ((g2977) & (!g142) & (!sk[43]) & (g563) & (!g583) & (g3123)) + ((g2977) & (!g142) & (!sk[43]) & (g563) & (g583) & (!g3123)) + ((g2977) & (!g142) & (!sk[43]) & (g563) & (g583) & (g3123)) + ((g2977) & (!g142) & (sk[43]) & (!g563) & (!g583) & (g3123)) + ((g2977) & (!g142) & (sk[43]) & (!g563) & (g583) & (g3123)) + ((g2977) & (!g142) & (sk[43]) & (g563) & (!g583) & (g3123)) + ((g2977) & (!g142) & (sk[43]) & (g563) & (g583) & (g3123)) + ((g2977) & (g142) & (!sk[43]) & (!g563) & (!g583) & (!g3123)) + ((g2977) & (g142) & (!sk[43]) & (!g563) & (!g583) & (g3123)) + ((g2977) & (g142) & (!sk[43]) & (!g563) & (g583) & (!g3123)) + ((g2977) & (g142) & (!sk[43]) & (!g563) & (g583) & (g3123)) + ((g2977) & (g142) & (!sk[43]) & (g563) & (!g583) & (!g3123)) + ((g2977) & (g142) & (!sk[43]) & (g563) & (!g583) & (g3123)) + ((g2977) & (g142) & (!sk[43]) & (g563) & (g583) & (!g3123)) + ((g2977) & (g142) & (!sk[43]) & (g563) & (g583) & (g3123)) + ((g2977) & (g142) & (sk[43]) & (!g563) & (!g583) & (g3123)) + ((g2977) & (g142) & (sk[43]) & (!g563) & (g583) & (g3123)) + ((g2977) & (g142) & (sk[43]) & (g563) & (!g583) & (g3123)) + ((g2977) & (g142) & (sk[43]) & (g563) & (g583) & (g3123)));
	assign g3125 = (((!g2071) & (!g2070) & (!g2074) & (!g2104) & (!g2105) & (g2077)) + ((!g2071) & (!g2070) & (!g2074) & (g2104) & (!g2105) & (g2077)) + ((!g2071) & (!g2070) & (g2074) & (!g2104) & (!g2105) & (!g2077)) + ((!g2071) & (!g2070) & (g2074) & (!g2104) & (!g2105) & (g2077)) + ((!g2071) & (!g2070) & (g2074) & (!g2104) & (g2105) & (g2077)) + ((!g2071) & (!g2070) & (g2074) & (g2104) & (!g2105) & (g2077)) + ((!g2071) & (g2070) & (!g2074) & (!g2104) & (!g2105) & (g2077)) + ((!g2071) & (g2070) & (!g2074) & (g2104) & (!g2105) & (g2077)) + ((!g2071) & (g2070) & (g2074) & (!g2104) & (!g2105) & (!g2077)) + ((!g2071) & (g2070) & (g2074) & (!g2104) & (!g2105) & (g2077)) + ((!g2071) & (g2070) & (g2074) & (!g2104) & (g2105) & (g2077)) + ((!g2071) & (g2070) & (g2074) & (g2104) & (!g2105) & (g2077)) + ((g2071) & (!g2070) & (!g2074) & (!g2104) & (!g2105) & (!g2077)) + ((g2071) & (!g2070) & (!g2074) & (!g2104) & (!g2105) & (g2077)) + ((g2071) & (!g2070) & (!g2074) & (!g2104) & (g2105) & (g2077)) + ((g2071) & (!g2070) & (!g2074) & (g2104) & (!g2105) & (g2077)) + ((g2071) & (!g2070) & (g2074) & (!g2104) & (!g2105) & (!g2077)) + ((g2071) & (!g2070) & (g2074) & (!g2104) & (!g2105) & (g2077)) + ((g2071) & (!g2070) & (g2074) & (!g2104) & (g2105) & (g2077)) + ((g2071) & (!g2070) & (g2074) & (g2104) & (!g2105) & (!g2077)) + ((g2071) & (!g2070) & (g2074) & (g2104) & (!g2105) & (g2077)) + ((g2071) & (!g2070) & (g2074) & (g2104) & (g2105) & (g2077)) + ((g2071) & (g2070) & (!g2074) & (!g2104) & (!g2105) & (g2077)) + ((g2071) & (g2070) & (!g2074) & (g2104) & (!g2105) & (g2077)) + ((g2071) & (g2070) & (g2074) & (!g2104) & (!g2105) & (!g2077)) + ((g2071) & (g2070) & (g2074) & (!g2104) & (!g2105) & (g2077)) + ((g2071) & (g2070) & (g2074) & (!g2104) & (g2105) & (g2077)) + ((g2071) & (g2070) & (g2074) & (g2104) & (!g2105) & (g2077)));
	assign g3126 = (((!sk[45]) & (!g2094) & (g2642)) + ((!sk[45]) & (g2094) & (g2642)) + ((sk[45]) & (!g2094) & (!g2642)) + ((sk[45]) & (g2094) & (g2642)));
	assign g3127 = (((!sk[46]) & (!g2093) & (g2625)) + ((!sk[46]) & (g2093) & (g2625)) + ((sk[46]) & (!g2093) & (!g2625)) + ((sk[46]) & (g2093) & (g2625)));
	assign g3128 = (((!g2839) & (!g2538) & (!g2192) & (!g2780) & (!g2190) & (g2837)) + ((!g2839) & (!g2538) & (g2192) & (!g2780) & (!g2190) & (g2837)) + ((!g2839) & (!g2538) & (g2192) & (g2780) & (g2190) & (!g2837)) + ((!g2839) & (!g2538) & (g2192) & (g2780) & (g2190) & (g2837)) + ((!g2839) & (g2538) & (!g2192) & (!g2780) & (!g2190) & (g2837)) + ((!g2839) & (g2538) & (!g2192) & (!g2780) & (g2190) & (!g2837)) + ((!g2839) & (g2538) & (!g2192) & (!g2780) & (g2190) & (g2837)) + ((!g2839) & (g2538) & (g2192) & (!g2780) & (!g2190) & (g2837)) + ((!g2839) & (g2538) & (g2192) & (!g2780) & (g2190) & (!g2837)) + ((!g2839) & (g2538) & (g2192) & (!g2780) & (g2190) & (g2837)) + ((!g2839) & (g2538) & (g2192) & (g2780) & (g2190) & (!g2837)) + ((!g2839) & (g2538) & (g2192) & (g2780) & (g2190) & (g2837)) + ((g2839) & (!g2538) & (!g2192) & (!g2780) & (!g2190) & (g2837)) + ((g2839) & (!g2538) & (!g2192) & (g2780) & (!g2190) & (!g2837)) + ((g2839) & (!g2538) & (!g2192) & (g2780) & (!g2190) & (g2837)) + ((g2839) & (!g2538) & (g2192) & (!g2780) & (!g2190) & (g2837)) + ((g2839) & (!g2538) & (g2192) & (g2780) & (!g2190) & (!g2837)) + ((g2839) & (!g2538) & (g2192) & (g2780) & (!g2190) & (g2837)) + ((g2839) & (!g2538) & (g2192) & (g2780) & (g2190) & (!g2837)) + ((g2839) & (!g2538) & (g2192) & (g2780) & (g2190) & (g2837)) + ((g2839) & (g2538) & (!g2192) & (!g2780) & (!g2190) & (g2837)) + ((g2839) & (g2538) & (!g2192) & (!g2780) & (g2190) & (!g2837)) + ((g2839) & (g2538) & (!g2192) & (!g2780) & (g2190) & (g2837)) + ((g2839) & (g2538) & (!g2192) & (g2780) & (!g2190) & (!g2837)) + ((g2839) & (g2538) & (!g2192) & (g2780) & (!g2190) & (g2837)) + ((g2839) & (g2538) & (g2192) & (!g2780) & (!g2190) & (g2837)) + ((g2839) & (g2538) & (g2192) & (!g2780) & (g2190) & (!g2837)) + ((g2839) & (g2538) & (g2192) & (!g2780) & (g2190) & (g2837)) + ((g2839) & (g2538) & (g2192) & (g2780) & (!g2190) & (!g2837)) + ((g2839) & (g2538) & (g2192) & (g2780) & (!g2190) & (g2837)) + ((g2839) & (g2538) & (g2192) & (g2780) & (g2190) & (!g2837)) + ((g2839) & (g2538) & (g2192) & (g2780) & (g2190) & (g2837)));
	assign g3129 = (((!g2081) & (!g2125) & (!g2100) & (!g2811) & (!g2832) & (!g2833)) + ((!g2081) & (!g2125) & (!g2100) & (!g2811) & (g2832) & (!g2833)) + ((!g2081) & (!g2125) & (!g2100) & (g2811) & (!g2832) & (!g2833)) + ((!g2081) & (!g2125) & (!g2100) & (g2811) & (g2832) & (g2833)) + ((!g2081) & (!g2125) & (g2100) & (!g2811) & (!g2832) & (!g2833)) + ((!g2081) & (!g2125) & (g2100) & (!g2811) & (g2832) & (g2833)) + ((!g2081) & (!g2125) & (g2100) & (g2811) & (!g2832) & (g2833)) + ((!g2081) & (!g2125) & (g2100) & (g2811) & (g2832) & (g2833)) + ((g2081) & (g2125) & (!g2100) & (!g2811) & (!g2832) & (!g2833)) + ((g2081) & (g2125) & (!g2100) & (!g2811) & (!g2832) & (g2833)) + ((g2081) & (g2125) & (!g2100) & (!g2811) & (g2832) & (!g2833)) + ((g2081) & (g2125) & (!g2100) & (!g2811) & (g2832) & (g2833)) + ((g2081) & (g2125) & (!g2100) & (g2811) & (!g2832) & (!g2833)) + ((g2081) & (g2125) & (!g2100) & (g2811) & (!g2832) & (g2833)) + ((g2081) & (g2125) & (!g2100) & (g2811) & (g2832) & (!g2833)) + ((g2081) & (g2125) & (!g2100) & (g2811) & (g2832) & (g2833)) + ((g2081) & (g2125) & (g2100) & (!g2811) & (!g2832) & (!g2833)) + ((g2081) & (g2125) & (g2100) & (!g2811) & (!g2832) & (g2833)) + ((g2081) & (g2125) & (g2100) & (!g2811) & (g2832) & (!g2833)) + ((g2081) & (g2125) & (g2100) & (!g2811) & (g2832) & (g2833)) + ((g2081) & (g2125) & (g2100) & (g2811) & (!g2832) & (!g2833)) + ((g2081) & (g2125) & (g2100) & (g2811) & (!g2832) & (g2833)) + ((g2081) & (g2125) & (g2100) & (g2811) & (g2832) & (!g2833)) + ((g2081) & (g2125) & (g2100) & (g2811) & (g2832) & (g2833)));
	assign g3130 = (((!g2798) & (!g2799) & (!g2814) & (!sk[49]) & (g2815)) + ((!g2798) & (!g2799) & (!g2814) & (sk[49]) & (g2815)) + ((!g2798) & (!g2799) & (g2814) & (!sk[49]) & (g2815)) + ((!g2798) & (!g2799) & (g2814) & (sk[49]) & (!g2815)) + ((!g2798) & (g2799) & (!g2814) & (!sk[49]) & (!g2815)) + ((!g2798) & (g2799) & (!g2814) & (!sk[49]) & (g2815)) + ((!g2798) & (g2799) & (!g2814) & (sk[49]) & (!g2815)) + ((!g2798) & (g2799) & (g2814) & (!sk[49]) & (!g2815)) + ((!g2798) & (g2799) & (g2814) & (!sk[49]) & (g2815)) + ((!g2798) & (g2799) & (g2814) & (sk[49]) & (g2815)) + ((g2798) & (!g2799) & (!g2814) & (!sk[49]) & (!g2815)) + ((g2798) & (!g2799) & (!g2814) & (!sk[49]) & (g2815)) + ((g2798) & (!g2799) & (!g2814) & (sk[49]) & (!g2815)) + ((g2798) & (!g2799) & (g2814) & (!sk[49]) & (!g2815)) + ((g2798) & (!g2799) & (g2814) & (!sk[49]) & (g2815)) + ((g2798) & (!g2799) & (g2814) & (sk[49]) & (g2815)) + ((g2798) & (g2799) & (!g2814) & (!sk[49]) & (!g2815)) + ((g2798) & (g2799) & (!g2814) & (!sk[49]) & (g2815)) + ((g2798) & (g2799) & (!g2814) & (sk[49]) & (!g2815)) + ((g2798) & (g2799) & (g2814) & (!sk[49]) & (!g2815)) + ((g2798) & (g2799) & (g2814) & (!sk[49]) & (g2815)) + ((g2798) & (g2799) & (g2814) & (sk[49]) & (g2815)));
	assign g3131 = (((!g2081) & (!g2798) & (!g2799) & (!g2100) & (!g2811) & (g3130)) + ((!g2081) & (!g2798) & (!g2799) & (!g2100) & (g2811) & (g3130)) + ((!g2081) & (!g2798) & (!g2799) & (g2100) & (!g2811) & (g3130)) + ((!g2081) & (!g2798) & (!g2799) & (g2100) & (g2811) & (g3130)) + ((!g2081) & (!g2798) & (g2799) & (!g2100) & (!g2811) & (!g3130)) + ((!g2081) & (!g2798) & (g2799) & (!g2100) & (g2811) & (!g3130)) + ((!g2081) & (!g2798) & (g2799) & (g2100) & (!g2811) & (!g3130)) + ((!g2081) & (!g2798) & (g2799) & (g2100) & (g2811) & (!g3130)) + ((!g2081) & (g2798) & (!g2799) & (!g2100) & (!g2811) & (!g3130)) + ((!g2081) & (g2798) & (!g2799) & (!g2100) & (g2811) & (!g3130)) + ((!g2081) & (g2798) & (!g2799) & (g2100) & (!g2811) & (!g3130)) + ((!g2081) & (g2798) & (!g2799) & (g2100) & (g2811) & (!g3130)) + ((!g2081) & (g2798) & (g2799) & (!g2100) & (!g2811) & (g3130)) + ((!g2081) & (g2798) & (g2799) & (!g2100) & (g2811) & (g3130)) + ((!g2081) & (g2798) & (g2799) & (g2100) & (!g2811) & (g3130)) + ((!g2081) & (g2798) & (g2799) & (g2100) & (g2811) & (g3130)) + ((g2081) & (!g2798) & (!g2799) & (g2100) & (g2811) & (!g3130)) + ((g2081) & (!g2798) & (!g2799) & (g2100) & (g2811) & (g3130)) + ((g2081) & (!g2798) & (g2799) & (g2100) & (g2811) & (!g3130)) + ((g2081) & (!g2798) & (g2799) & (g2100) & (g2811) & (g3130)) + ((g2081) & (g2798) & (!g2799) & (g2100) & (g2811) & (!g3130)) + ((g2081) & (g2798) & (!g2799) & (g2100) & (g2811) & (g3130)) + ((g2081) & (g2798) & (g2799) & (g2100) & (g2811) & (!g3130)) + ((g2081) & (g2798) & (g2799) & (g2100) & (g2811) & (g3130)));
	assign g3132 = (((!g2081) & (!g2125) & (!g2796) & (!sk[51]) & (g3130) & (!g3131)) + ((!g2081) & (!g2125) & (!g2796) & (!sk[51]) & (g3130) & (g3131)) + ((!g2081) & (!g2125) & (g2796) & (!sk[51]) & (!g3130) & (!g3131)) + ((!g2081) & (!g2125) & (g2796) & (!sk[51]) & (!g3130) & (g3131)) + ((!g2081) & (!g2125) & (g2796) & (!sk[51]) & (g3130) & (!g3131)) + ((!g2081) & (!g2125) & (g2796) & (!sk[51]) & (g3130) & (g3131)) + ((!g2081) & (g2125) & (!g2796) & (!sk[51]) & (g3130) & (!g3131)) + ((!g2081) & (g2125) & (!g2796) & (!sk[51]) & (g3130) & (g3131)) + ((!g2081) & (g2125) & (!g2796) & (sk[51]) & (!g3130) & (!g3131)) + ((!g2081) & (g2125) & (!g2796) & (sk[51]) & (!g3130) & (g3131)) + ((!g2081) & (g2125) & (g2796) & (!sk[51]) & (!g3130) & (!g3131)) + ((!g2081) & (g2125) & (g2796) & (!sk[51]) & (!g3130) & (g3131)) + ((!g2081) & (g2125) & (g2796) & (!sk[51]) & (g3130) & (!g3131)) + ((!g2081) & (g2125) & (g2796) & (!sk[51]) & (g3130) & (g3131)) + ((!g2081) & (g2125) & (g2796) & (sk[51]) & (!g3130) & (!g3131)) + ((!g2081) & (g2125) & (g2796) & (sk[51]) & (!g3130) & (g3131)) + ((g2081) & (!g2125) & (!g2796) & (!sk[51]) & (!g3130) & (!g3131)) + ((g2081) & (!g2125) & (!g2796) & (!sk[51]) & (!g3130) & (g3131)) + ((g2081) & (!g2125) & (!g2796) & (!sk[51]) & (g3130) & (!g3131)) + ((g2081) & (!g2125) & (!g2796) & (!sk[51]) & (g3130) & (g3131)) + ((g2081) & (!g2125) & (g2796) & (!sk[51]) & (!g3130) & (!g3131)) + ((g2081) & (!g2125) & (g2796) & (!sk[51]) & (!g3130) & (g3131)) + ((g2081) & (!g2125) & (g2796) & (!sk[51]) & (g3130) & (!g3131)) + ((g2081) & (!g2125) & (g2796) & (!sk[51]) & (g3130) & (g3131)) + ((g2081) & (!g2125) & (g2796) & (sk[51]) & (!g3130) & (!g3131)) + ((g2081) & (!g2125) & (g2796) & (sk[51]) & (!g3130) & (g3131)) + ((g2081) & (!g2125) & (g2796) & (sk[51]) & (g3130) & (!g3131)) + ((g2081) & (!g2125) & (g2796) & (sk[51]) & (g3130) & (g3131)) + ((g2081) & (g2125) & (!g2796) & (!sk[51]) & (!g3130) & (!g3131)) + ((g2081) & (g2125) & (!g2796) & (!sk[51]) & (!g3130) & (g3131)) + ((g2081) & (g2125) & (!g2796) & (!sk[51]) & (g3130) & (!g3131)) + ((g2081) & (g2125) & (!g2796) & (!sk[51]) & (g3130) & (g3131)) + ((g2081) & (g2125) & (!g2796) & (sk[51]) & (!g3130) & (!g3131)) + ((g2081) & (g2125) & (!g2796) & (sk[51]) & (g3130) & (!g3131)) + ((g2081) & (g2125) & (g2796) & (!sk[51]) & (!g3130) & (!g3131)) + ((g2081) & (g2125) & (g2796) & (!sk[51]) & (!g3130) & (g3131)) + ((g2081) & (g2125) & (g2796) & (!sk[51]) & (g3130) & (!g3131)) + ((g2081) & (g2125) & (g2796) & (!sk[51]) & (g3130) & (g3131)) + ((g2081) & (g2125) & (g2796) & (sk[51]) & (!g3130) & (!g3131)) + ((g2081) & (g2125) & (g2796) & (sk[51]) & (g3130) & (!g3131)));
	assign g3133 = (((!g817) & (!g770) & (!g774) & (!g821) & (!g864) & (!g868)) + ((!g817) & (!g770) & (!g774) & (!g821) & (g864) & (g868)) + ((!g817) & (g770) & (!g774) & (!g821) & (!g864) & (!g868)) + ((!g817) & (g770) & (!g774) & (!g821) & (g864) & (g868)) + ((!g817) & (g770) & (g774) & (!g821) & (!g864) & (!g868)) + ((!g817) & (g770) & (g774) & (!g821) & (g864) & (g868)) + ((g817) & (!g770) & (!g774) & (!g821) & (!g864) & (!g868)) + ((g817) & (!g770) & (!g774) & (!g821) & (g864) & (g868)) + ((g817) & (!g770) & (!g774) & (g821) & (!g864) & (!g868)) + ((g817) & (!g770) & (!g774) & (g821) & (g864) & (g868)) + ((g817) & (!g770) & (g774) & (!g821) & (!g864) & (!g868)) + ((g817) & (!g770) & (g774) & (!g821) & (g864) & (g868)) + ((g817) & (g770) & (!g774) & (!g821) & (!g864) & (!g868)) + ((g817) & (g770) & (!g774) & (!g821) & (g864) & (g868)) + ((g817) & (g770) & (!g774) & (g821) & (!g864) & (!g868)) + ((g817) & (g770) & (!g774) & (g821) & (g864) & (g868)) + ((g817) & (g770) & (g774) & (!g821) & (!g864) & (!g868)) + ((g817) & (g770) & (g774) & (!g821) & (g864) & (g868)) + ((g817) & (g770) & (g774) & (g821) & (!g864) & (!g868)) + ((g817) & (g770) & (g774) & (g821) & (g864) & (g868)));
	assign g3134 = (((!g817) & (!g770) & (!g774) & (!g821) & (!g723) & (!g727)) + ((!g817) & (!g770) & (!g774) & (!g821) & (!g723) & (g727)) + ((!g817) & (!g770) & (!g774) & (!g821) & (g723) & (g727)) + ((!g817) & (!g770) & (!g774) & (g821) & (!g723) & (!g727)) + ((!g817) & (!g770) & (!g774) & (g821) & (!g723) & (g727)) + ((!g817) & (!g770) & (!g774) & (g821) & (g723) & (g727)) + ((!g817) & (!g770) & (g774) & (!g821) & (!g723) & (!g727)) + ((!g817) & (!g770) & (g774) & (!g821) & (!g723) & (g727)) + ((!g817) & (!g770) & (g774) & (!g821) & (g723) & (g727)) + ((!g817) & (!g770) & (g774) & (g821) & (!g723) & (!g727)) + ((!g817) & (!g770) & (g774) & (g821) & (!g723) & (g727)) + ((!g817) & (!g770) & (g774) & (g821) & (g723) & (g727)) + ((!g817) & (g770) & (g774) & (!g821) & (!g723) & (!g727)) + ((!g817) & (g770) & (g774) & (!g821) & (!g723) & (g727)) + ((!g817) & (g770) & (g774) & (!g821) & (g723) & (g727)) + ((!g817) & (g770) & (g774) & (g821) & (!g723) & (!g727)) + ((!g817) & (g770) & (g774) & (g821) & (!g723) & (g727)) + ((!g817) & (g770) & (g774) & (g821) & (g723) & (g727)) + ((g817) & (!g770) & (!g774) & (g821) & (!g723) & (!g727)) + ((g817) & (!g770) & (!g774) & (g821) & (!g723) & (g727)) + ((g817) & (!g770) & (!g774) & (g821) & (g723) & (g727)) + ((g817) & (!g770) & (g774) & (g821) & (!g723) & (!g727)) + ((g817) & (!g770) & (g774) & (g821) & (!g723) & (g727)) + ((g817) & (!g770) & (g774) & (g821) & (g723) & (g727)) + ((g817) & (g770) & (g774) & (g821) & (!g723) & (!g727)) + ((g817) & (g770) & (g774) & (g821) & (!g723) & (g727)) + ((g817) & (g770) & (g774) & (g821) & (g723) & (g727)));
	assign g3135 = (((!g723) & (!sk[54]) & (!g727) & (!g3133) & (g3134)) + ((!g723) & (!sk[54]) & (!g727) & (g3133) & (g3134)) + ((!g723) & (!sk[54]) & (g727) & (!g3133) & (!g3134)) + ((!g723) & (!sk[54]) & (g727) & (!g3133) & (g3134)) + ((!g723) & (!sk[54]) & (g727) & (g3133) & (!g3134)) + ((!g723) & (!sk[54]) & (g727) & (g3133) & (g3134)) + ((!g723) & (sk[54]) & (!g727) & (g3133) & (!g3134)) + ((!g723) & (sk[54]) & (!g727) & (g3133) & (g3134)) + ((!g723) & (sk[54]) & (g727) & (g3133) & (!g3134)) + ((g723) & (!sk[54]) & (!g727) & (!g3133) & (!g3134)) + ((g723) & (!sk[54]) & (!g727) & (!g3133) & (g3134)) + ((g723) & (!sk[54]) & (!g727) & (g3133) & (!g3134)) + ((g723) & (!sk[54]) & (!g727) & (g3133) & (g3134)) + ((g723) & (!sk[54]) & (g727) & (!g3133) & (!g3134)) + ((g723) & (!sk[54]) & (g727) & (!g3133) & (g3134)) + ((g723) & (!sk[54]) & (g727) & (g3133) & (!g3134)) + ((g723) & (!sk[54]) & (g727) & (g3133) & (g3134)) + ((g723) & (sk[54]) & (!g727) & (g3133) & (!g3134)) + ((g723) & (sk[54]) & (!g727) & (g3133) & (g3134)) + ((g723) & (sk[54]) & (g727) & (g3133) & (!g3134)) + ((g723) & (sk[54]) & (g727) & (g3133) & (g3134)));
	assign g3136 = (((!g2119) & (!g2120) & (g2482) & (g2507) & (!g2121) & (g2529)) + ((!g2119) & (!g2120) & (g2482) & (g2507) & (g2121) & (!g2529)) + ((!g2119) & (g2120) & (!g2482) & (g2507) & (!g2121) & (g2529)) + ((!g2119) & (g2120) & (!g2482) & (g2507) & (g2121) & (!g2529)) + ((!g2119) & (g2120) & (g2482) & (!g2507) & (!g2121) & (g2529)) + ((!g2119) & (g2120) & (g2482) & (!g2507) & (g2121) & (!g2529)) + ((!g2119) & (g2120) & (g2482) & (g2507) & (!g2121) & (g2529)) + ((!g2119) & (g2120) & (g2482) & (g2507) & (g2121) & (!g2529)) + ((g2119) & (!g2120) & (!g2482) & (g2507) & (!g2121) & (g2529)) + ((g2119) & (!g2120) & (!g2482) & (g2507) & (g2121) & (!g2529)) + ((g2119) & (!g2120) & (g2482) & (g2507) & (!g2121) & (g2529)) + ((g2119) & (!g2120) & (g2482) & (g2507) & (g2121) & (!g2529)) + ((g2119) & (g2120) & (!g2482) & (!g2507) & (!g2121) & (g2529)) + ((g2119) & (g2120) & (!g2482) & (!g2507) & (g2121) & (!g2529)) + ((g2119) & (g2120) & (!g2482) & (g2507) & (!g2121) & (g2529)) + ((g2119) & (g2120) & (!g2482) & (g2507) & (g2121) & (!g2529)) + ((g2119) & (g2120) & (g2482) & (!g2507) & (!g2121) & (g2529)) + ((g2119) & (g2120) & (g2482) & (!g2507) & (g2121) & (!g2529)) + ((g2119) & (g2120) & (g2482) & (g2507) & (!g2121) & (g2529)) + ((g2119) & (g2120) & (g2482) & (g2507) & (g2121) & (!g2529)));
	assign g3137 = (((!g2119) & (!g2120) & (!g2482) & (!g2507) & (!g2118) & (!g2457)) + ((!g2119) & (!g2120) & (!g2482) & (!g2507) & (!g2118) & (g2457)) + ((!g2119) & (!g2120) & (!g2482) & (!g2507) & (g2118) & (!g2457)) + ((!g2119) & (!g2120) & (!g2482) & (g2507) & (!g2118) & (!g2457)) + ((!g2119) & (!g2120) & (!g2482) & (g2507) & (!g2118) & (g2457)) + ((!g2119) & (!g2120) & (!g2482) & (g2507) & (g2118) & (!g2457)) + ((!g2119) & (!g2120) & (g2482) & (!g2507) & (!g2118) & (!g2457)) + ((!g2119) & (!g2120) & (g2482) & (!g2507) & (!g2118) & (g2457)) + ((!g2119) & (!g2120) & (g2482) & (!g2507) & (g2118) & (!g2457)) + ((!g2119) & (!g2120) & (g2482) & (g2507) & (!g2118) & (!g2457)) + ((!g2119) & (!g2120) & (g2482) & (g2507) & (!g2118) & (g2457)) + ((!g2119) & (!g2120) & (g2482) & (g2507) & (g2118) & (!g2457)) + ((!g2119) & (g2120) & (!g2482) & (!g2507) & (!g2118) & (!g2457)) + ((!g2119) & (g2120) & (!g2482) & (!g2507) & (!g2118) & (g2457)) + ((!g2119) & (g2120) & (!g2482) & (!g2507) & (g2118) & (!g2457)) + ((!g2119) & (g2120) & (g2482) & (!g2507) & (!g2118) & (!g2457)) + ((!g2119) & (g2120) & (g2482) & (!g2507) & (!g2118) & (g2457)) + ((!g2119) & (g2120) & (g2482) & (!g2507) & (g2118) & (!g2457)) + ((g2119) & (!g2120) & (!g2482) & (!g2507) & (!g2118) & (!g2457)) + ((g2119) & (!g2120) & (!g2482) & (!g2507) & (!g2118) & (g2457)) + ((g2119) & (!g2120) & (!g2482) & (!g2507) & (g2118) & (!g2457)) + ((g2119) & (!g2120) & (!g2482) & (g2507) & (!g2118) & (!g2457)) + ((g2119) & (!g2120) & (!g2482) & (g2507) & (!g2118) & (g2457)) + ((g2119) & (!g2120) & (!g2482) & (g2507) & (g2118) & (!g2457)) + ((g2119) & (g2120) & (!g2482) & (!g2507) & (!g2118) & (!g2457)) + ((g2119) & (g2120) & (!g2482) & (!g2507) & (!g2118) & (g2457)) + ((g2119) & (g2120) & (!g2482) & (!g2507) & (g2118) & (!g2457)));
	assign g3138 = (((!g2118) & (!g2457) & (!g3136) & (!sk[57]) & (g3137)) + ((!g2118) & (!g2457) & (g3136) & (!sk[57]) & (g3137)) + ((!g2118) & (!g2457) & (g3136) & (sk[57]) & (!g3137)) + ((!g2118) & (g2457) & (!g3136) & (!sk[57]) & (!g3137)) + ((!g2118) & (g2457) & (!g3136) & (!sk[57]) & (g3137)) + ((!g2118) & (g2457) & (g3136) & (!sk[57]) & (!g3137)) + ((!g2118) & (g2457) & (g3136) & (!sk[57]) & (g3137)) + ((!g2118) & (g2457) & (g3136) & (sk[57]) & (!g3137)) + ((!g2118) & (g2457) & (g3136) & (sk[57]) & (g3137)) + ((g2118) & (!g2457) & (!g3136) & (!sk[57]) & (!g3137)) + ((g2118) & (!g2457) & (!g3136) & (!sk[57]) & (g3137)) + ((g2118) & (!g2457) & (g3136) & (!sk[57]) & (!g3137)) + ((g2118) & (!g2457) & (g3136) & (!sk[57]) & (g3137)) + ((g2118) & (!g2457) & (g3136) & (sk[57]) & (!g3137)) + ((g2118) & (!g2457) & (g3136) & (sk[57]) & (g3137)) + ((g2118) & (g2457) & (!g3136) & (!sk[57]) & (!g3137)) + ((g2118) & (g2457) & (!g3136) & (!sk[57]) & (g3137)) + ((g2118) & (g2457) & (g3136) & (!sk[57]) & (!g3137)) + ((g2118) & (g2457) & (g3136) & (!sk[57]) & (g3137)) + ((g2118) & (g2457) & (g3136) & (sk[57]) & (!g3137)) + ((g2118) & (g2457) & (g3136) & (sk[57]) & (g3137)));
	assign g3139 = (((!g3117) & (!g102) & (!sk[58]) & (!g93) & (g86) & (!g85)) + ((!g3117) & (!g102) & (!sk[58]) & (!g93) & (g86) & (g85)) + ((!g3117) & (!g102) & (!sk[58]) & (g93) & (!g86) & (!g85)) + ((!g3117) & (!g102) & (!sk[58]) & (g93) & (!g86) & (g85)) + ((!g3117) & (!g102) & (!sk[58]) & (g93) & (g86) & (!g85)) + ((!g3117) & (!g102) & (!sk[58]) & (g93) & (g86) & (g85)) + ((!g3117) & (!g102) & (sk[58]) & (!g93) & (!g86) & (!g85)) + ((!g3117) & (!g102) & (sk[58]) & (!g93) & (!g86) & (g85)) + ((!g3117) & (!g102) & (sk[58]) & (!g93) & (g86) & (!g85)) + ((!g3117) & (!g102) & (sk[58]) & (!g93) & (g86) & (g85)) + ((!g3117) & (!g102) & (sk[58]) & (g93) & (g86) & (g85)) + ((!g3117) & (g102) & (!sk[58]) & (!g93) & (g86) & (!g85)) + ((!g3117) & (g102) & (!sk[58]) & (!g93) & (g86) & (g85)) + ((!g3117) & (g102) & (!sk[58]) & (g93) & (!g86) & (!g85)) + ((!g3117) & (g102) & (!sk[58]) & (g93) & (!g86) & (g85)) + ((!g3117) & (g102) & (!sk[58]) & (g93) & (g86) & (!g85)) + ((!g3117) & (g102) & (!sk[58]) & (g93) & (g86) & (g85)) + ((g3117) & (!g102) & (!sk[58]) & (!g93) & (!g86) & (!g85)) + ((g3117) & (!g102) & (!sk[58]) & (!g93) & (!g86) & (g85)) + ((g3117) & (!g102) & (!sk[58]) & (!g93) & (g86) & (!g85)) + ((g3117) & (!g102) & (!sk[58]) & (!g93) & (g86) & (g85)) + ((g3117) & (!g102) & (!sk[58]) & (g93) & (!g86) & (!g85)) + ((g3117) & (!g102) & (!sk[58]) & (g93) & (!g86) & (g85)) + ((g3117) & (!g102) & (!sk[58]) & (g93) & (g86) & (!g85)) + ((g3117) & (!g102) & (!sk[58]) & (g93) & (g86) & (g85)) + ((g3117) & (!g102) & (sk[58]) & (!g93) & (!g86) & (!g85)) + ((g3117) & (!g102) & (sk[58]) & (!g93) & (!g86) & (g85)) + ((g3117) & (!g102) & (sk[58]) & (!g93) & (g86) & (!g85)) + ((g3117) & (!g102) & (sk[58]) & (!g93) & (g86) & (g85)) + ((g3117) & (!g102) & (sk[58]) & (g93) & (g86) & (g85)) + ((g3117) & (g102) & (!sk[58]) & (!g93) & (!g86) & (!g85)) + ((g3117) & (g102) & (!sk[58]) & (!g93) & (!g86) & (g85)) + ((g3117) & (g102) & (!sk[58]) & (!g93) & (g86) & (!g85)) + ((g3117) & (g102) & (!sk[58]) & (!g93) & (g86) & (g85)) + ((g3117) & (g102) & (!sk[58]) & (g93) & (!g86) & (!g85)) + ((g3117) & (g102) & (!sk[58]) & (g93) & (!g86) & (g85)) + ((g3117) & (g102) & (!sk[58]) & (g93) & (g86) & (!g85)) + ((g3117) & (g102) & (!sk[58]) & (g93) & (g86) & (g85)) + ((g3117) & (g102) & (sk[58]) & (!g93) & (!g86) & (!g85)) + ((g3117) & (g102) & (sk[58]) & (!g93) & (!g86) & (g85)) + ((g3117) & (g102) & (sk[58]) & (!g93) & (g86) & (!g85)) + ((g3117) & (g102) & (sk[58]) & (!g93) & (g86) & (g85)) + ((g3117) & (g102) & (sk[58]) & (g93) & (g86) & (g85)));
	assign g3140 = (((!g2081) & (!g2080) & (!g3141) & (!g2125) & (!g2836) & (!g2834)) + ((!g2081) & (!g2080) & (!g3141) & (!g2125) & (!g2836) & (g2834)) + ((!g2081) & (!g2080) & (!g3141) & (!g2125) & (g2836) & (!g2834)) + ((!g2081) & (!g2080) & (!g3141) & (!g2125) & (g2836) & (g2834)) + ((!g2081) & (!g2080) & (!g3141) & (g2125) & (!g2836) & (!g2834)) + ((!g2081) & (!g2080) & (!g3141) & (g2125) & (!g2836) & (g2834)) + ((!g2081) & (!g2080) & (!g3141) & (g2125) & (g2836) & (!g2834)) + ((!g2081) & (!g2080) & (!g3141) & (g2125) & (g2836) & (g2834)) + ((!g2081) & (g2080) & (!g3141) & (!g2125) & (!g2836) & (!g2834)) + ((!g2081) & (g2080) & (!g3141) & (!g2125) & (!g2836) & (g2834)) + ((!g2081) & (g2080) & (!g3141) & (!g2125) & (g2836) & (!g2834)) + ((!g2081) & (g2080) & (!g3141) & (!g2125) & (g2836) & (g2834)) + ((!g2081) & (g2080) & (!g3141) & (g2125) & (g2836) & (!g2834)) + ((!g2081) & (g2080) & (!g3141) & (g2125) & (g2836) & (g2834)) + ((g2081) & (!g2080) & (!g3141) & (!g2125) & (!g2836) & (!g2834)) + ((g2081) & (!g2080) & (!g3141) & (!g2125) & (!g2836) & (g2834)) + ((g2081) & (!g2080) & (!g3141) & (!g2125) & (g2836) & (!g2834)) + ((g2081) & (!g2080) & (!g3141) & (!g2125) & (g2836) & (g2834)) + ((g2081) & (!g2080) & (!g3141) & (g2125) & (!g2836) & (!g2834)) + ((g2081) & (!g2080) & (!g3141) & (g2125) & (!g2836) & (g2834)) + ((g2081) & (!g2080) & (!g3141) & (g2125) & (g2836) & (!g2834)) + ((g2081) & (!g2080) & (!g3141) & (g2125) & (g2836) & (g2834)) + ((g2081) & (g2080) & (!g3141) & (!g2125) & (!g2836) & (g2834)) + ((g2081) & (g2080) & (!g3141) & (!g2125) & (g2836) & (g2834)) + ((g2081) & (g2080) & (!g3141) & (g2125) & (!g2836) & (!g2834)) + ((g2081) & (g2080) & (!g3141) & (g2125) & (!g2836) & (g2834)) + ((g2081) & (g2080) & (!g3141) & (g2125) & (g2836) & (!g2834)) + ((g2081) & (g2080) & (!g3141) & (g2125) & (g2836) & (g2834)));
	assign g3141 = (((!g2080) & (!g3129) & (!g3128) & (!sk[60]) & (g2125)) + ((!g2080) & (!g3129) & (!g3128) & (sk[60]) & (!g2125)) + ((!g2080) & (!g3129) & (!g3128) & (sk[60]) & (g2125)) + ((!g2080) & (!g3129) & (g3128) & (!sk[60]) & (g2125)) + ((!g2080) & (g3129) & (!g3128) & (!sk[60]) & (!g2125)) + ((!g2080) & (g3129) & (!g3128) & (!sk[60]) & (g2125)) + ((!g2080) & (g3129) & (!g3128) & (sk[60]) & (!g2125)) + ((!g2080) & (g3129) & (!g3128) & (sk[60]) & (g2125)) + ((!g2080) & (g3129) & (g3128) & (!sk[60]) & (!g2125)) + ((!g2080) & (g3129) & (g3128) & (!sk[60]) & (g2125)) + ((g2080) & (!g3129) & (!g3128) & (!sk[60]) & (!g2125)) + ((g2080) & (!g3129) & (!g3128) & (!sk[60]) & (g2125)) + ((g2080) & (!g3129) & (g3128) & (!sk[60]) & (!g2125)) + ((g2080) & (!g3129) & (g3128) & (!sk[60]) & (g2125)) + ((g2080) & (g3129) & (!g3128) & (!sk[60]) & (!g2125)) + ((g2080) & (g3129) & (!g3128) & (!sk[60]) & (g2125)) + ((g2080) & (g3129) & (!g3128) & (sk[60]) & (!g2125)) + ((g2080) & (g3129) & (!g3128) & (sk[60]) & (g2125)) + ((g2080) & (g3129) & (g3128) & (!sk[60]) & (!g2125)) + ((g2080) & (g3129) & (g3128) & (!sk[60]) & (g2125)) + ((g2080) & (g3129) & (g3128) & (sk[60]) & (!g2125)));
	assign g3142 = (((!g2591) & (!g2590) & (!g2085) & (g2571) & (g2555) & (g2554)) + ((!g2591) & (!g2590) & (g2085) & (!g2571) & (!g2555) & (!g2554)) + ((!g2591) & (!g2590) & (g2085) & (!g2571) & (!g2555) & (g2554)) + ((!g2591) & (!g2590) & (g2085) & (!g2571) & (g2555) & (!g2554)) + ((!g2591) & (!g2590) & (g2085) & (!g2571) & (g2555) & (g2554)) + ((!g2591) & (!g2590) & (g2085) & (g2571) & (!g2555) & (!g2554)) + ((!g2591) & (!g2590) & (g2085) & (g2571) & (!g2555) & (g2554)) + ((!g2591) & (!g2590) & (g2085) & (g2571) & (g2555) & (!g2554)) + ((!g2591) & (g2590) & (!g2085) & (!g2571) & (!g2555) & (!g2554)) + ((!g2591) & (g2590) & (!g2085) & (!g2571) & (!g2555) & (g2554)) + ((!g2591) & (g2590) & (!g2085) & (!g2571) & (g2555) & (!g2554)) + ((!g2591) & (g2590) & (!g2085) & (!g2571) & (g2555) & (g2554)) + ((!g2591) & (g2590) & (!g2085) & (g2571) & (!g2555) & (!g2554)) + ((!g2591) & (g2590) & (!g2085) & (g2571) & (!g2555) & (g2554)) + ((!g2591) & (g2590) & (!g2085) & (g2571) & (g2555) & (!g2554)) + ((!g2591) & (g2590) & (g2085) & (g2571) & (g2555) & (g2554)) + ((g2591) & (!g2590) & (!g2085) & (!g2571) & (!g2555) & (!g2554)) + ((g2591) & (!g2590) & (!g2085) & (!g2571) & (!g2555) & (g2554)) + ((g2591) & (!g2590) & (!g2085) & (!g2571) & (g2555) & (!g2554)) + ((g2591) & (!g2590) & (!g2085) & (!g2571) & (g2555) & (g2554)) + ((g2591) & (!g2590) & (!g2085) & (g2571) & (!g2555) & (!g2554)) + ((g2591) & (!g2590) & (!g2085) & (g2571) & (!g2555) & (g2554)) + ((g2591) & (!g2590) & (!g2085) & (g2571) & (g2555) & (!g2554)) + ((g2591) & (!g2590) & (g2085) & (g2571) & (g2555) & (g2554)) + ((g2591) & (g2590) & (!g2085) & (g2571) & (g2555) & (g2554)) + ((g2591) & (g2590) & (g2085) & (!g2571) & (!g2555) & (!g2554)) + ((g2591) & (g2590) & (g2085) & (!g2571) & (!g2555) & (g2554)) + ((g2591) & (g2590) & (g2085) & (!g2571) & (g2555) & (!g2554)) + ((g2591) & (g2590) & (g2085) & (!g2571) & (g2555) & (g2554)) + ((g2591) & (g2590) & (g2085) & (g2571) & (!g2555) & (!g2554)) + ((g2591) & (g2590) & (g2085) & (g2571) & (!g2555) & (g2554)) + ((g2591) & (g2590) & (g2085) & (g2571) & (g2555) & (!g2554)));
	assign g3143 = (((!g2077) & (!g2105) & (!g2104) & (!g2074) & (!g2241) & (!g2186)) + ((!g2077) & (!g2105) & (!g2104) & (!g2074) & (g2241) & (g2186)) + ((!g2077) & (!g2105) & (!g2104) & (g2074) & (g2241) & (!g2186)) + ((!g2077) & (!g2105) & (!g2104) & (g2074) & (g2241) & (g2186)) + ((!g2077) & (!g2105) & (g2104) & (!g2074) & (!g2241) & (!g2186)) + ((!g2077) & (!g2105) & (g2104) & (!g2074) & (!g2241) & (g2186)) + ((!g2077) & (!g2105) & (g2104) & (g2074) & (!g2241) & (!g2186)) + ((!g2077) & (!g2105) & (g2104) & (g2074) & (g2241) & (g2186)) + ((!g2077) & (g2105) & (!g2104) & (!g2074) & (!g2241) & (!g2186)) + ((!g2077) & (g2105) & (!g2104) & (!g2074) & (!g2241) & (g2186)) + ((!g2077) & (g2105) & (!g2104) & (g2074) & (!g2241) & (!g2186)) + ((!g2077) & (g2105) & (!g2104) & (g2074) & (!g2241) & (g2186)) + ((!g2077) & (g2105) & (g2104) & (!g2074) & (!g2241) & (!g2186)) + ((!g2077) & (g2105) & (g2104) & (!g2074) & (!g2241) & (g2186)) + ((!g2077) & (g2105) & (g2104) & (g2074) & (!g2241) & (!g2186)) + ((!g2077) & (g2105) & (g2104) & (g2074) & (!g2241) & (g2186)) + ((g2077) & (!g2105) & (!g2104) & (!g2074) & (g2241) & (!g2186)) + ((g2077) & (!g2105) & (!g2104) & (!g2074) & (g2241) & (g2186)) + ((g2077) & (!g2105) & (!g2104) & (g2074) & (g2241) & (!g2186)) + ((g2077) & (!g2105) & (!g2104) & (g2074) & (g2241) & (g2186)) + ((g2077) & (!g2105) & (g2104) & (!g2074) & (g2241) & (!g2186)) + ((g2077) & (!g2105) & (g2104) & (!g2074) & (g2241) & (g2186)) + ((g2077) & (!g2105) & (g2104) & (g2074) & (g2241) & (!g2186)) + ((g2077) & (!g2105) & (g2104) & (g2074) & (g2241) & (g2186)) + ((g2077) & (g2105) & (!g2104) & (!g2074) & (!g2241) & (!g2186)) + ((g2077) & (g2105) & (!g2104) & (!g2074) & (g2241) & (g2186)) + ((g2077) & (g2105) & (!g2104) & (g2074) & (g2241) & (!g2186)) + ((g2077) & (g2105) & (!g2104) & (g2074) & (g2241) & (g2186)) + ((g2077) & (g2105) & (g2104) & (!g2074) & (!g2241) & (!g2186)) + ((g2077) & (g2105) & (g2104) & (!g2074) & (!g2241) & (g2186)) + ((g2077) & (g2105) & (g2104) & (g2074) & (!g2241) & (!g2186)) + ((g2077) & (g2105) & (g2104) & (g2074) & (g2241) & (g2186)));
	assign g3144 = (((!g2077) & (!g2105) & (!g2104) & (!g2074) & (!g2070) & (g2071)) + ((!g2077) & (!g2105) & (!g2104) & (g2074) & (!g2070) & (!g2071)) + ((!g2077) & (!g2105) & (!g2104) & (g2074) & (!g2070) & (g2071)) + ((!g2077) & (!g2105) & (!g2104) & (g2074) & (g2070) & (!g2071)) + ((!g2077) & (!g2105) & (!g2104) & (g2074) & (g2070) & (g2071)) + ((!g2077) & (!g2105) & (g2104) & (g2074) & (!g2070) & (g2071)) + ((!g2077) & (g2105) & (!g2104) & (!g2074) & (!g2070) & (!g2071)) + ((!g2077) & (g2105) & (!g2104) & (!g2074) & (g2070) & (!g2071)) + ((!g2077) & (g2105) & (!g2104) & (!g2074) & (g2070) & (g2071)) + ((!g2077) & (g2105) & (g2104) & (!g2074) & (!g2070) & (!g2071)) + ((!g2077) & (g2105) & (g2104) & (!g2074) & (!g2070) & (g2071)) + ((!g2077) & (g2105) & (g2104) & (!g2074) & (g2070) & (!g2071)) + ((!g2077) & (g2105) & (g2104) & (!g2074) & (g2070) & (g2071)) + ((!g2077) & (g2105) & (g2104) & (g2074) & (!g2070) & (!g2071)) + ((!g2077) & (g2105) & (g2104) & (g2074) & (g2070) & (!g2071)) + ((!g2077) & (g2105) & (g2104) & (g2074) & (g2070) & (g2071)) + ((g2077) & (!g2105) & (!g2104) & (!g2074) & (!g2070) & (!g2071)) + ((g2077) & (!g2105) & (!g2104) & (!g2074) & (g2070) & (!g2071)) + ((g2077) & (!g2105) & (!g2104) & (!g2074) & (g2070) & (g2071)) + ((g2077) & (!g2105) & (g2104) & (!g2074) & (!g2070) & (!g2071)) + ((g2077) & (!g2105) & (g2104) & (!g2074) & (!g2070) & (g2071)) + ((g2077) & (!g2105) & (g2104) & (!g2074) & (g2070) & (!g2071)) + ((g2077) & (!g2105) & (g2104) & (!g2074) & (g2070) & (g2071)) + ((g2077) & (!g2105) & (g2104) & (g2074) & (!g2070) & (!g2071)) + ((g2077) & (!g2105) & (g2104) & (g2074) & (g2070) & (!g2071)) + ((g2077) & (!g2105) & (g2104) & (g2074) & (g2070) & (g2071)) + ((g2077) & (g2105) & (!g2104) & (!g2074) & (!g2070) & (g2071)) + ((g2077) & (g2105) & (!g2104) & (g2074) & (!g2070) & (!g2071)) + ((g2077) & (g2105) & (!g2104) & (g2074) & (!g2070) & (g2071)) + ((g2077) & (g2105) & (!g2104) & (g2074) & (g2070) & (!g2071)) + ((g2077) & (g2105) & (!g2104) & (g2074) & (g2070) & (g2071)) + ((g2077) & (g2105) & (g2104) & (g2074) & (!g2070) & (g2071)));
	assign g3145 = (((!g2104) & (!g2070) & (!g2071) & (!sk[64]) & (g2074) & (!g2125)) + ((!g2104) & (!g2070) & (!g2071) & (!sk[64]) & (g2074) & (g2125)) + ((!g2104) & (!g2070) & (!g2071) & (sk[64]) & (g2074) & (!g2125)) + ((!g2104) & (!g2070) & (!g2071) & (sk[64]) & (g2074) & (g2125)) + ((!g2104) & (!g2070) & (g2071) & (!sk[64]) & (!g2074) & (!g2125)) + ((!g2104) & (!g2070) & (g2071) & (!sk[64]) & (!g2074) & (g2125)) + ((!g2104) & (!g2070) & (g2071) & (!sk[64]) & (g2074) & (!g2125)) + ((!g2104) & (!g2070) & (g2071) & (!sk[64]) & (g2074) & (g2125)) + ((!g2104) & (!g2070) & (g2071) & (sk[64]) & (!g2074) & (g2125)) + ((!g2104) & (!g2070) & (g2071) & (sk[64]) & (g2074) & (!g2125)) + ((!g2104) & (g2070) & (!g2071) & (!sk[64]) & (g2074) & (!g2125)) + ((!g2104) & (g2070) & (!g2071) & (!sk[64]) & (g2074) & (g2125)) + ((!g2104) & (g2070) & (!g2071) & (sk[64]) & (g2074) & (!g2125)) + ((!g2104) & (g2070) & (!g2071) & (sk[64]) & (g2074) & (g2125)) + ((!g2104) & (g2070) & (g2071) & (!sk[64]) & (!g2074) & (!g2125)) + ((!g2104) & (g2070) & (g2071) & (!sk[64]) & (!g2074) & (g2125)) + ((!g2104) & (g2070) & (g2071) & (!sk[64]) & (g2074) & (!g2125)) + ((!g2104) & (g2070) & (g2071) & (!sk[64]) & (g2074) & (g2125)) + ((!g2104) & (g2070) & (g2071) & (sk[64]) & (!g2074) & (!g2125)) + ((!g2104) & (g2070) & (g2071) & (sk[64]) & (g2074) & (g2125)) + ((g2104) & (!g2070) & (!g2071) & (!sk[64]) & (!g2074) & (!g2125)) + ((g2104) & (!g2070) & (!g2071) & (!sk[64]) & (!g2074) & (g2125)) + ((g2104) & (!g2070) & (!g2071) & (!sk[64]) & (g2074) & (!g2125)) + ((g2104) & (!g2070) & (!g2071) & (!sk[64]) & (g2074) & (g2125)) + ((g2104) & (!g2070) & (!g2071) & (sk[64]) & (!g2074) & (!g2125)) + ((g2104) & (!g2070) & (!g2071) & (sk[64]) & (!g2074) & (g2125)) + ((g2104) & (!g2070) & (g2071) & (!sk[64]) & (!g2074) & (!g2125)) + ((g2104) & (!g2070) & (g2071) & (!sk[64]) & (!g2074) & (g2125)) + ((g2104) & (!g2070) & (g2071) & (!sk[64]) & (g2074) & (!g2125)) + ((g2104) & (!g2070) & (g2071) & (!sk[64]) & (g2074) & (g2125)) + ((g2104) & (!g2070) & (g2071) & (sk[64]) & (!g2074) & (!g2125)) + ((g2104) & (!g2070) & (g2071) & (sk[64]) & (g2074) & (g2125)) + ((g2104) & (g2070) & (!g2071) & (!sk[64]) & (!g2074) & (!g2125)) + ((g2104) & (g2070) & (!g2071) & (!sk[64]) & (!g2074) & (g2125)) + ((g2104) & (g2070) & (!g2071) & (!sk[64]) & (g2074) & (!g2125)) + ((g2104) & (g2070) & (!g2071) & (!sk[64]) & (g2074) & (g2125)) + ((g2104) & (g2070) & (!g2071) & (sk[64]) & (!g2074) & (!g2125)) + ((g2104) & (g2070) & (!g2071) & (sk[64]) & (!g2074) & (g2125)) + ((g2104) & (g2070) & (g2071) & (!sk[64]) & (!g2074) & (!g2125)) + ((g2104) & (g2070) & (g2071) & (!sk[64]) & (!g2074) & (g2125)) + ((g2104) & (g2070) & (g2071) & (!sk[64]) & (g2074) & (!g2125)) + ((g2104) & (g2070) & (g2071) & (!sk[64]) & (g2074) & (g2125)) + ((g2104) & (g2070) & (g2071) & (sk[64]) & (!g2074) & (g2125)) + ((g2104) & (g2070) & (g2071) & (sk[64]) & (g2074) & (!g2125)));
	assign g3146 = (((!g2079) & (!g2104) & (!g2070) & (!g2071) & (g2074) & (!g2125)) + ((!g2079) & (!g2104) & (!g2070) & (g2071) & (g2074) & (!g2125)) + ((!g2079) & (!g2104) & (g2070) & (!g2071) & (g2074) & (!g2125)) + ((!g2079) & (!g2104) & (g2070) & (g2071) & (!g2074) & (!g2125)) + ((!g2079) & (g2104) & (!g2070) & (!g2071) & (!g2074) & (!g2125)) + ((!g2079) & (g2104) & (!g2070) & (!g2071) & (g2074) & (g2125)) + ((!g2079) & (g2104) & (!g2070) & (g2071) & (!g2074) & (!g2125)) + ((!g2079) & (g2104) & (!g2070) & (g2071) & (g2074) & (g2125)) + ((!g2079) & (g2104) & (g2070) & (!g2071) & (!g2074) & (!g2125)) + ((!g2079) & (g2104) & (g2070) & (!g2071) & (g2074) & (g2125)) + ((!g2079) & (g2104) & (g2070) & (g2071) & (g2074) & (!g2125)) + ((!g2079) & (g2104) & (g2070) & (g2071) & (g2074) & (g2125)) + ((g2079) & (!g2104) & (!g2070) & (!g2071) & (g2074) & (!g2125)) + ((g2079) & (!g2104) & (!g2070) & (g2071) & (!g2074) & (!g2125)) + ((g2079) & (!g2104) & (g2070) & (!g2071) & (!g2074) & (!g2125)) + ((g2079) & (!g2104) & (g2070) & (g2071) & (!g2074) & (!g2125)) + ((g2079) & (g2104) & (!g2070) & (!g2071) & (!g2074) & (!g2125)) + ((g2079) & (g2104) & (!g2070) & (!g2071) & (g2074) & (g2125)) + ((g2079) & (g2104) & (!g2070) & (g2071) & (g2074) & (!g2125)) + ((g2079) & (g2104) & (!g2070) & (g2071) & (g2074) & (g2125)) + ((g2079) & (g2104) & (g2070) & (!g2071) & (g2074) & (!g2125)) + ((g2079) & (g2104) & (g2070) & (!g2071) & (g2074) & (g2125)) + ((g2079) & (g2104) & (g2070) & (g2071) & (g2074) & (!g2125)) + ((g2079) & (g2104) & (g2070) & (g2071) & (g2074) & (g2125)));
	assign g3147 = (((!g3145) & (g3146) & (!sk[66]) & (!g2081)) + ((!g3145) & (g3146) & (!sk[66]) & (g2081)) + ((!g3145) & (g3146) & (sk[66]) & (g2081)) + ((g3145) & (!g3146) & (!sk[66]) & (!g2081)) + ((g3145) & (!g3146) & (!sk[66]) & (g2081)) + ((g3145) & (!g3146) & (sk[66]) & (!g2081)) + ((g3145) & (g3146) & (!sk[66]) & (!g2081)) + ((g3145) & (g3146) & (!sk[66]) & (g2081)) + ((g3145) & (g3146) & (sk[66]) & (!g2081)) + ((g3145) & (g3146) & (sk[66]) & (g2081)));
	assign g3148 = (((!g3149) & (!sk[67]) & (g3150)) + ((!g3149) & (sk[67]) & (!g3150)) + ((g3149) & (!sk[67]) & (g3150)));
	assign g3149 = (((!g2764) & (!sk[68]) & (g3151)) + ((!g2764) & (sk[68]) & (g3151)) + ((g2764) & (!sk[68]) & (g3151)));
	assign g3150 = (((!g2764) & (!sk[69]) & (g3154)) + ((g2764) & (!sk[69]) & (g3154)) + ((g2764) & (sk[69]) & (g3154)));
	assign g3151 = (((!sk[70]) & (!g3152) & (g3153)) + ((!sk[70]) & (g3152) & (g3153)) + ((sk[70]) & (!g3152) & (!g3153)));
	assign g3152 = (((!sk[71]) & (!g2356) & (g3157)) + ((!sk[71]) & (g2356) & (g3157)) + ((sk[71]) & (!g2356) & (g3157)));
	assign g3153 = (((!sk[72]) & (!g2356) & (g3158)) + ((!sk[72]) & (g2356) & (g3158)) + ((sk[72]) & (g2356) & (g3158)));
	assign g3154 = (((!g3155) & (!sk[73]) & (g3156)) + ((!g3155) & (sk[73]) & (!g3156)) + ((g3155) & (!sk[73]) & (g3156)));
	assign g3155 = (((!sk[74]) & (!g2356) & (g3159)) + ((!sk[74]) & (g2356) & (g3159)) + ((sk[74]) & (!g2356) & (g3159)));
	assign g3156 = (((!sk[75]) & (!g2356) & (g3160)) + ((!sk[75]) & (g2356) & (g3160)) + ((sk[75]) & (g2356) & (g3160)));
	assign g3157 = (((!sk[76]) & (!g2768) & (!g2766) & (!g2028) & (g2843)) + ((!sk[76]) & (!g2768) & (!g2766) & (g2028) & (g2843)) + ((!sk[76]) & (!g2768) & (g2766) & (!g2028) & (!g2843)) + ((!sk[76]) & (!g2768) & (g2766) & (!g2028) & (g2843)) + ((!sk[76]) & (!g2768) & (g2766) & (g2028) & (!g2843)) + ((!sk[76]) & (!g2768) & (g2766) & (g2028) & (g2843)) + ((!sk[76]) & (g2768) & (!g2766) & (!g2028) & (!g2843)) + ((!sk[76]) & (g2768) & (!g2766) & (!g2028) & (g2843)) + ((!sk[76]) & (g2768) & (!g2766) & (g2028) & (!g2843)) + ((!sk[76]) & (g2768) & (!g2766) & (g2028) & (g2843)) + ((!sk[76]) & (g2768) & (g2766) & (!g2028) & (!g2843)) + ((!sk[76]) & (g2768) & (g2766) & (!g2028) & (g2843)) + ((!sk[76]) & (g2768) & (g2766) & (g2028) & (!g2843)) + ((!sk[76]) & (g2768) & (g2766) & (g2028) & (g2843)) + ((sk[76]) & (!g2768) & (g2766) & (g2028) & (g2843)) + ((sk[76]) & (g2768) & (!g2766) & (g2028) & (g2843)) + ((sk[76]) & (g2768) & (g2766) & (g2028) & (g2843)));
	assign g3158 = (((!g1955) & (!sk[77]) & (g2843)) + ((g1955) & (!sk[77]) & (g2843)) + ((g1955) & (sk[77]) & (g2843)));
	assign g3159 = (((!g2768) & (!g2766) & (!g2028) & (!sk[78]) & (g2843)) + ((!g2768) & (!g2766) & (!g2028) & (sk[78]) & (!g2843)) + ((!g2768) & (!g2766) & (!g2028) & (sk[78]) & (g2843)) + ((!g2768) & (!g2766) & (g2028) & (!sk[78]) & (g2843)) + ((!g2768) & (!g2766) & (g2028) & (sk[78]) & (!g2843)) + ((!g2768) & (g2766) & (!g2028) & (!sk[78]) & (!g2843)) + ((!g2768) & (g2766) & (!g2028) & (!sk[78]) & (g2843)) + ((!g2768) & (g2766) & (!g2028) & (sk[78]) & (!g2843)) + ((!g2768) & (g2766) & (!g2028) & (sk[78]) & (g2843)) + ((!g2768) & (g2766) & (g2028) & (!sk[78]) & (!g2843)) + ((!g2768) & (g2766) & (g2028) & (!sk[78]) & (g2843)) + ((!g2768) & (g2766) & (g2028) & (sk[78]) & (!g2843)) + ((!g2768) & (g2766) & (g2028) & (sk[78]) & (g2843)) + ((g2768) & (!g2766) & (!g2028) & (!sk[78]) & (!g2843)) + ((g2768) & (!g2766) & (!g2028) & (!sk[78]) & (g2843)) + ((g2768) & (!g2766) & (!g2028) & (sk[78]) & (!g2843)) + ((g2768) & (!g2766) & (!g2028) & (sk[78]) & (g2843)) + ((g2768) & (!g2766) & (g2028) & (!sk[78]) & (!g2843)) + ((g2768) & (!g2766) & (g2028) & (!sk[78]) & (g2843)) + ((g2768) & (!g2766) & (g2028) & (sk[78]) & (!g2843)) + ((g2768) & (!g2766) & (g2028) & (sk[78]) & (g2843)) + ((g2768) & (g2766) & (!g2028) & (!sk[78]) & (!g2843)) + ((g2768) & (g2766) & (!g2028) & (!sk[78]) & (g2843)) + ((g2768) & (g2766) & (!g2028) & (sk[78]) & (!g2843)) + ((g2768) & (g2766) & (!g2028) & (sk[78]) & (g2843)) + ((g2768) & (g2766) & (g2028) & (!sk[78]) & (!g2843)) + ((g2768) & (g2766) & (g2028) & (!sk[78]) & (g2843)) + ((g2768) & (g2766) & (g2028) & (sk[78]) & (!g2843)) + ((g2768) & (g2766) & (g2028) & (sk[78]) & (g2843)));
	assign g3160 = (((!sk[79]) & (!g1955) & (g2843)) + ((!sk[79]) & (g1955) & (g2843)) + ((sk[79]) & (!g1955) & (!g2843)) + ((sk[79]) & (g1955) & (!g2843)) + ((sk[79]) & (g1955) & (g2843)));
	assign g3161 = (((!g3162) & (!sk[80]) & (g3163)) + ((!g3162) & (sk[80]) & (!g3163)) + ((g3162) & (!sk[80]) & (g3163)));
	assign g3162 = (((!sk[81]) & (!g2746) & (g3164)) + ((!sk[81]) & (g2746) & (g3164)) + ((sk[81]) & (!g2746) & (g3164)));
	assign g3163 = (((!g2746) & (!sk[82]) & (g3167)) + ((g2746) & (!sk[82]) & (g3167)) + ((g2746) & (sk[82]) & (g3167)));
	assign g3164 = (((!sk[83]) & (!g3165) & (g3166)) + ((!sk[83]) & (g3165) & (g3166)) + ((sk[83]) & (!g3165) & (!g3166)));
	assign g3165 = (((!sk[84]) & (!g2356) & (g3170)) + ((!sk[84]) & (g2356) & (g3170)) + ((sk[84]) & (!g2356) & (g3170)));
	assign g3166 = (((!sk[85]) & (!g2356) & (g3171)) + ((!sk[85]) & (g2356) & (g3171)) + ((sk[85]) & (g2356) & (g3171)));
	assign g3167 = (((!g3168) & (!sk[86]) & (g3169)) + ((!g3168) & (sk[86]) & (!g3169)) + ((g3168) & (!sk[86]) & (g3169)));
	assign g3168 = (((!g2356) & (!sk[87]) & (g3172)) + ((!g2356) & (sk[87]) & (g3172)) + ((g2356) & (!sk[87]) & (g3172)));
	assign g3169 = (((!sk[88]) & (!g2356) & (g3173)) + ((!sk[88]) & (g2356) & (g3173)) + ((sk[88]) & (g2356) & (g3173)));
	assign g3170 = (((!sk[89]) & (!g2749) & (!g2747) & (!g2028) & (g2843)) + ((!sk[89]) & (!g2749) & (!g2747) & (g2028) & (g2843)) + ((!sk[89]) & (!g2749) & (g2747) & (!g2028) & (!g2843)) + ((!sk[89]) & (!g2749) & (g2747) & (!g2028) & (g2843)) + ((!sk[89]) & (!g2749) & (g2747) & (g2028) & (!g2843)) + ((!sk[89]) & (!g2749) & (g2747) & (g2028) & (g2843)) + ((!sk[89]) & (g2749) & (!g2747) & (!g2028) & (!g2843)) + ((!sk[89]) & (g2749) & (!g2747) & (!g2028) & (g2843)) + ((!sk[89]) & (g2749) & (!g2747) & (g2028) & (!g2843)) + ((!sk[89]) & (g2749) & (!g2747) & (g2028) & (g2843)) + ((!sk[89]) & (g2749) & (g2747) & (!g2028) & (!g2843)) + ((!sk[89]) & (g2749) & (g2747) & (!g2028) & (g2843)) + ((!sk[89]) & (g2749) & (g2747) & (g2028) & (!g2843)) + ((!sk[89]) & (g2749) & (g2747) & (g2028) & (g2843)) + ((sk[89]) & (!g2749) & (g2747) & (g2028) & (g2843)) + ((sk[89]) & (g2749) & (!g2747) & (g2028) & (g2843)) + ((sk[89]) & (g2749) & (g2747) & (g2028) & (g2843)));
	assign g3171 = (((!g1942) & (!sk[90]) & (g2843)) + ((g1942) & (!sk[90]) & (g2843)) + ((g1942) & (sk[90]) & (g2843)));
	assign g3172 = (((!sk[91]) & (!g2749) & (!g2747) & (!g2028) & (g2843)) + ((!sk[91]) & (!g2749) & (!g2747) & (g2028) & (g2843)) + ((!sk[91]) & (!g2749) & (g2747) & (!g2028) & (!g2843)) + ((!sk[91]) & (!g2749) & (g2747) & (!g2028) & (g2843)) + ((!sk[91]) & (!g2749) & (g2747) & (g2028) & (!g2843)) + ((!sk[91]) & (!g2749) & (g2747) & (g2028) & (g2843)) + ((!sk[91]) & (g2749) & (!g2747) & (!g2028) & (!g2843)) + ((!sk[91]) & (g2749) & (!g2747) & (!g2028) & (g2843)) + ((!sk[91]) & (g2749) & (!g2747) & (g2028) & (!g2843)) + ((!sk[91]) & (g2749) & (!g2747) & (g2028) & (g2843)) + ((!sk[91]) & (g2749) & (g2747) & (!g2028) & (!g2843)) + ((!sk[91]) & (g2749) & (g2747) & (!g2028) & (g2843)) + ((!sk[91]) & (g2749) & (g2747) & (g2028) & (!g2843)) + ((!sk[91]) & (g2749) & (g2747) & (g2028) & (g2843)) + ((sk[91]) & (!g2749) & (!g2747) & (!g2028) & (!g2843)) + ((sk[91]) & (!g2749) & (!g2747) & (!g2028) & (g2843)) + ((sk[91]) & (!g2749) & (!g2747) & (g2028) & (!g2843)) + ((sk[91]) & (!g2749) & (g2747) & (!g2028) & (!g2843)) + ((sk[91]) & (!g2749) & (g2747) & (!g2028) & (g2843)) + ((sk[91]) & (!g2749) & (g2747) & (g2028) & (!g2843)) + ((sk[91]) & (!g2749) & (g2747) & (g2028) & (g2843)) + ((sk[91]) & (g2749) & (!g2747) & (!g2028) & (!g2843)) + ((sk[91]) & (g2749) & (!g2747) & (!g2028) & (g2843)) + ((sk[91]) & (g2749) & (!g2747) & (g2028) & (!g2843)) + ((sk[91]) & (g2749) & (!g2747) & (g2028) & (g2843)) + ((sk[91]) & (g2749) & (g2747) & (!g2028) & (!g2843)) + ((sk[91]) & (g2749) & (g2747) & (!g2028) & (g2843)) + ((sk[91]) & (g2749) & (g2747) & (g2028) & (!g2843)) + ((sk[91]) & (g2749) & (g2747) & (g2028) & (g2843)));
	assign g3173 = (((!sk[92]) & (!g1942) & (g2843)) + ((!sk[92]) & (g1942) & (g2843)) + ((sk[92]) & (!g1942) & (!g2843)) + ((sk[92]) & (g1942) & (!g2843)) + ((sk[92]) & (g1942) & (g2843)));
	assign g3174 = (((!g3175) & (!sk[93]) & (g3176)) + ((!g3175) & (sk[93]) & (!g3176)) + ((g3175) & (!sk[93]) & (g3176)));
	assign g3175 = (((!g2691) & (!sk[94]) & (g3177)) + ((!g2691) & (sk[94]) & (g3177)) + ((g2691) & (!sk[94]) & (g3177)));
	assign g3176 = (((!g2691) & (!sk[95]) & (g3180)) + ((g2691) & (!sk[95]) & (g3180)) + ((g2691) & (sk[95]) & (g3180)));
	assign g3177 = (((!g3178) & (!sk[96]) & (g3179)) + ((!g3178) & (sk[96]) & (!g3179)) + ((g3178) & (!sk[96]) & (g3179)));
	assign g3178 = (((!g2356) & (!sk[97]) & (g3183)) + ((!g2356) & (sk[97]) & (g3183)) + ((g2356) & (!sk[97]) & (g3183)));
	assign g3179 = (((!g2356) & (!sk[98]) & (g3184)) + ((g2356) & (!sk[98]) & (g3184)) + ((g2356) & (sk[98]) & (g3184)));
	assign g3180 = (((!sk[99]) & (!g3181) & (g3182)) + ((!sk[99]) & (g3181) & (g3182)) + ((sk[99]) & (!g3181) & (!g3182)));
	assign g3181 = (((!g2356) & (!sk[100]) & (g3185)) + ((!g2356) & (sk[100]) & (g3185)) + ((g2356) & (!sk[100]) & (g3185)));
	assign g3182 = (((!g2356) & (!sk[101]) & (g3186)) + ((g2356) & (!sk[101]) & (g3186)) + ((g2356) & (sk[101]) & (g3186)));
	assign g3183 = (((!sk[102]) & (!g2697) & (!g2695) & (!g2028) & (g2843)) + ((!sk[102]) & (!g2697) & (!g2695) & (g2028) & (g2843)) + ((!sk[102]) & (!g2697) & (g2695) & (!g2028) & (!g2843)) + ((!sk[102]) & (!g2697) & (g2695) & (!g2028) & (g2843)) + ((!sk[102]) & (!g2697) & (g2695) & (g2028) & (!g2843)) + ((!sk[102]) & (!g2697) & (g2695) & (g2028) & (g2843)) + ((!sk[102]) & (g2697) & (!g2695) & (!g2028) & (!g2843)) + ((!sk[102]) & (g2697) & (!g2695) & (!g2028) & (g2843)) + ((!sk[102]) & (g2697) & (!g2695) & (g2028) & (!g2843)) + ((!sk[102]) & (g2697) & (!g2695) & (g2028) & (g2843)) + ((!sk[102]) & (g2697) & (g2695) & (!g2028) & (!g2843)) + ((!sk[102]) & (g2697) & (g2695) & (!g2028) & (g2843)) + ((!sk[102]) & (g2697) & (g2695) & (g2028) & (!g2843)) + ((!sk[102]) & (g2697) & (g2695) & (g2028) & (g2843)) + ((sk[102]) & (!g2697) & (g2695) & (g2028) & (g2843)) + ((sk[102]) & (g2697) & (!g2695) & (g2028) & (g2843)) + ((sk[102]) & (g2697) & (g2695) & (g2028) & (g2843)));
	assign g3184 = (((!g1902) & (!sk[103]) & (g2843)) + ((g1902) & (!sk[103]) & (g2843)) + ((g1902) & (sk[103]) & (g2843)));
	assign g3185 = (((!g2697) & (!sk[104]) & (!g2695) & (!g2028) & (g2843)) + ((!g2697) & (!sk[104]) & (!g2695) & (g2028) & (g2843)) + ((!g2697) & (!sk[104]) & (g2695) & (!g2028) & (!g2843)) + ((!g2697) & (!sk[104]) & (g2695) & (!g2028) & (g2843)) + ((!g2697) & (!sk[104]) & (g2695) & (g2028) & (!g2843)) + ((!g2697) & (!sk[104]) & (g2695) & (g2028) & (g2843)) + ((!g2697) & (sk[104]) & (!g2695) & (!g2028) & (!g2843)) + ((!g2697) & (sk[104]) & (!g2695) & (!g2028) & (g2843)) + ((!g2697) & (sk[104]) & (!g2695) & (g2028) & (!g2843)) + ((!g2697) & (sk[104]) & (g2695) & (!g2028) & (!g2843)) + ((!g2697) & (sk[104]) & (g2695) & (!g2028) & (g2843)) + ((!g2697) & (sk[104]) & (g2695) & (g2028) & (!g2843)) + ((!g2697) & (sk[104]) & (g2695) & (g2028) & (g2843)) + ((g2697) & (!sk[104]) & (!g2695) & (!g2028) & (!g2843)) + ((g2697) & (!sk[104]) & (!g2695) & (!g2028) & (g2843)) + ((g2697) & (!sk[104]) & (!g2695) & (g2028) & (!g2843)) + ((g2697) & (!sk[104]) & (!g2695) & (g2028) & (g2843)) + ((g2697) & (!sk[104]) & (g2695) & (!g2028) & (!g2843)) + ((g2697) & (!sk[104]) & (g2695) & (!g2028) & (g2843)) + ((g2697) & (!sk[104]) & (g2695) & (g2028) & (!g2843)) + ((g2697) & (!sk[104]) & (g2695) & (g2028) & (g2843)) + ((g2697) & (sk[104]) & (!g2695) & (!g2028) & (!g2843)) + ((g2697) & (sk[104]) & (!g2695) & (!g2028) & (g2843)) + ((g2697) & (sk[104]) & (!g2695) & (g2028) & (!g2843)) + ((g2697) & (sk[104]) & (!g2695) & (g2028) & (g2843)) + ((g2697) & (sk[104]) & (g2695) & (!g2028) & (!g2843)) + ((g2697) & (sk[104]) & (g2695) & (!g2028) & (g2843)) + ((g2697) & (sk[104]) & (g2695) & (g2028) & (!g2843)) + ((g2697) & (sk[104]) & (g2695) & (g2028) & (g2843)));
	assign g3186 = (((!g1902) & (!sk[105]) & (g2843)) + ((!g1902) & (sk[105]) & (!g2843)) + ((g1902) & (!sk[105]) & (g2843)) + ((g1902) & (sk[105]) & (!g2843)) + ((g1902) & (sk[105]) & (g2843)));
	assign g3187 = (((!sk[106]) & (!g3188) & (g3189)) + ((!sk[106]) & (g3188) & (g3189)) + ((sk[106]) & (!g3188) & (!g3189)));
	assign g3188 = (((!sk[107]) & (!g2654) & (g3190)) + ((!sk[107]) & (g2654) & (g3190)) + ((sk[107]) & (!g2654) & (g3190)));
	assign g3189 = (((!sk[108]) & (!g2654) & (g3193)) + ((!sk[108]) & (g2654) & (g3193)) + ((sk[108]) & (g2654) & (g3193)));
	assign g3190 = (((!g3191) & (!sk[109]) & (g3192)) + ((!g3191) & (sk[109]) & (!g3192)) + ((g3191) & (!sk[109]) & (g3192)));
	assign g3191 = (((!g2356) & (!sk[110]) & (g3196)) + ((!g2356) & (sk[110]) & (g3196)) + ((g2356) & (!sk[110]) & (g3196)));
	assign g3192 = (((!g2356) & (!sk[111]) & (g3197)) + ((g2356) & (!sk[111]) & (g3197)) + ((g2356) & (sk[111]) & (g3197)));
	assign g3193 = (((!sk[112]) & (!g3194) & (g3195)) + ((!sk[112]) & (g3194) & (g3195)) + ((sk[112]) & (!g3194) & (!g3195)));
	assign g3194 = (((!g2356) & (!sk[113]) & (g3198)) + ((!g2356) & (sk[113]) & (g3198)) + ((g2356) & (!sk[113]) & (g3198)));
	assign g3195 = (((!g2356) & (!sk[114]) & (g3199)) + ((g2356) & (!sk[114]) & (g3199)) + ((g2356) & (sk[114]) & (g3199)));
	assign g3196 = (((!g2658) & (!sk[115]) & (!g2656) & (!g2028) & (g2843)) + ((!g2658) & (!sk[115]) & (!g2656) & (g2028) & (g2843)) + ((!g2658) & (!sk[115]) & (g2656) & (!g2028) & (!g2843)) + ((!g2658) & (!sk[115]) & (g2656) & (!g2028) & (g2843)) + ((!g2658) & (!sk[115]) & (g2656) & (g2028) & (!g2843)) + ((!g2658) & (!sk[115]) & (g2656) & (g2028) & (g2843)) + ((!g2658) & (sk[115]) & (g2656) & (g2028) & (g2843)) + ((g2658) & (!sk[115]) & (!g2656) & (!g2028) & (!g2843)) + ((g2658) & (!sk[115]) & (!g2656) & (!g2028) & (g2843)) + ((g2658) & (!sk[115]) & (!g2656) & (g2028) & (!g2843)) + ((g2658) & (!sk[115]) & (!g2656) & (g2028) & (g2843)) + ((g2658) & (!sk[115]) & (g2656) & (!g2028) & (!g2843)) + ((g2658) & (!sk[115]) & (g2656) & (!g2028) & (g2843)) + ((g2658) & (!sk[115]) & (g2656) & (g2028) & (!g2843)) + ((g2658) & (!sk[115]) & (g2656) & (g2028) & (g2843)) + ((g2658) & (sk[115]) & (!g2656) & (g2028) & (g2843)) + ((g2658) & (sk[115]) & (g2656) & (g2028) & (g2843)));
	assign g3197 = (((!g1876) & (!sk[116]) & (g2843)) + ((g1876) & (!sk[116]) & (g2843)) + ((g1876) & (sk[116]) & (g2843)));
	assign g3198 = (((!g2658) & (!sk[117]) & (!g2656) & (!g2028) & (g2843)) + ((!g2658) & (!sk[117]) & (!g2656) & (g2028) & (g2843)) + ((!g2658) & (!sk[117]) & (g2656) & (!g2028) & (!g2843)) + ((!g2658) & (!sk[117]) & (g2656) & (!g2028) & (g2843)) + ((!g2658) & (!sk[117]) & (g2656) & (g2028) & (!g2843)) + ((!g2658) & (!sk[117]) & (g2656) & (g2028) & (g2843)) + ((!g2658) & (sk[117]) & (!g2656) & (!g2028) & (!g2843)) + ((!g2658) & (sk[117]) & (!g2656) & (!g2028) & (g2843)) + ((!g2658) & (sk[117]) & (!g2656) & (g2028) & (!g2843)) + ((!g2658) & (sk[117]) & (g2656) & (!g2028) & (!g2843)) + ((!g2658) & (sk[117]) & (g2656) & (!g2028) & (g2843)) + ((!g2658) & (sk[117]) & (g2656) & (g2028) & (!g2843)) + ((!g2658) & (sk[117]) & (g2656) & (g2028) & (g2843)) + ((g2658) & (!sk[117]) & (!g2656) & (!g2028) & (!g2843)) + ((g2658) & (!sk[117]) & (!g2656) & (!g2028) & (g2843)) + ((g2658) & (!sk[117]) & (!g2656) & (g2028) & (!g2843)) + ((g2658) & (!sk[117]) & (!g2656) & (g2028) & (g2843)) + ((g2658) & (!sk[117]) & (g2656) & (!g2028) & (!g2843)) + ((g2658) & (!sk[117]) & (g2656) & (!g2028) & (g2843)) + ((g2658) & (!sk[117]) & (g2656) & (g2028) & (!g2843)) + ((g2658) & (!sk[117]) & (g2656) & (g2028) & (g2843)) + ((g2658) & (sk[117]) & (!g2656) & (!g2028) & (!g2843)) + ((g2658) & (sk[117]) & (!g2656) & (!g2028) & (g2843)) + ((g2658) & (sk[117]) & (!g2656) & (g2028) & (!g2843)) + ((g2658) & (sk[117]) & (!g2656) & (g2028) & (g2843)) + ((g2658) & (sk[117]) & (g2656) & (!g2028) & (!g2843)) + ((g2658) & (sk[117]) & (g2656) & (!g2028) & (g2843)) + ((g2658) & (sk[117]) & (g2656) & (g2028) & (!g2843)) + ((g2658) & (sk[117]) & (g2656) & (g2028) & (g2843)));
	assign g3199 = (((!sk[118]) & (!g1876) & (g2843)) + ((!sk[118]) & (g1876) & (g2843)) + ((sk[118]) & (!g1876) & (!g2843)) + ((sk[118]) & (g1876) & (!g2843)) + ((sk[118]) & (g1876) & (g2843)));
	assign g3200 = (((!g3201) & (!sk[119]) & (g3202)) + ((!g3201) & (sk[119]) & (!g3202)) + ((g3201) & (!sk[119]) & (g3202)));
	assign g3201 = (((!sk[120]) & (!g2599) & (g3203)) + ((!sk[120]) & (g2599) & (g3203)) + ((sk[120]) & (!g2599) & (g3203)));
	assign g3202 = (((!sk[121]) & (!g2599) & (g3206)) + ((!sk[121]) & (g2599) & (g3206)) + ((sk[121]) & (g2599) & (g3206)));
	assign g3203 = (((!sk[122]) & (!g3204) & (g3205)) + ((!sk[122]) & (g3204) & (g3205)) + ((sk[122]) & (!g3204) & (!g3205)));
	assign g3204 = (((!g2356) & (!sk[123]) & (g3209)) + ((!g2356) & (sk[123]) & (g3209)) + ((g2356) & (!sk[123]) & (g3209)));
	assign g3205 = (((!sk[124]) & (!g2356) & (g3210)) + ((!sk[124]) & (g2356) & (g3210)) + ((sk[124]) & (g2356) & (g3210)));
	assign g3206 = (((!sk[125]) & (!g3207) & (g3208)) + ((!sk[125]) & (g3207) & (g3208)) + ((sk[125]) & (!g3207) & (!g3208)));
	assign g3207 = (((!g2356) & (!sk[126]) & (g3211)) + ((!g2356) & (sk[126]) & (g3211)) + ((g2356) & (!sk[126]) & (g3211)));
	assign g3208 = (((!g2356) & (!sk[127]) & (g3212)) + ((g2356) & (!sk[127]) & (g3212)) + ((g2356) & (sk[127]) & (g3212)));
	assign g3209 = (((!g2606) & (!g2604) & (!sk[0]) & (!g2028) & (g2843)) + ((!g2606) & (!g2604) & (!sk[0]) & (g2028) & (g2843)) + ((!g2606) & (g2604) & (!sk[0]) & (!g2028) & (!g2843)) + ((!g2606) & (g2604) & (!sk[0]) & (!g2028) & (g2843)) + ((!g2606) & (g2604) & (!sk[0]) & (g2028) & (!g2843)) + ((!g2606) & (g2604) & (!sk[0]) & (g2028) & (g2843)) + ((!g2606) & (g2604) & (sk[0]) & (g2028) & (g2843)) + ((g2606) & (!g2604) & (!sk[0]) & (!g2028) & (!g2843)) + ((g2606) & (!g2604) & (!sk[0]) & (!g2028) & (g2843)) + ((g2606) & (!g2604) & (!sk[0]) & (g2028) & (!g2843)) + ((g2606) & (!g2604) & (!sk[0]) & (g2028) & (g2843)) + ((g2606) & (!g2604) & (sk[0]) & (g2028) & (g2843)) + ((g2606) & (g2604) & (!sk[0]) & (!g2028) & (!g2843)) + ((g2606) & (g2604) & (!sk[0]) & (!g2028) & (g2843)) + ((g2606) & (g2604) & (!sk[0]) & (g2028) & (!g2843)) + ((g2606) & (g2604) & (!sk[0]) & (g2028) & (g2843)) + ((g2606) & (g2604) & (sk[0]) & (g2028) & (g2843)));
	assign g3210 = (((!sk[1]) & (!g1837) & (g2843)) + ((!sk[1]) & (g1837) & (g2843)) + ((sk[1]) & (g1837) & (g2843)));
	assign g3211 = (((!g2606) & (!g2604) & (!g2028) & (!sk[2]) & (g2843)) + ((!g2606) & (!g2604) & (!g2028) & (sk[2]) & (!g2843)) + ((!g2606) & (!g2604) & (!g2028) & (sk[2]) & (g2843)) + ((!g2606) & (!g2604) & (g2028) & (!sk[2]) & (g2843)) + ((!g2606) & (!g2604) & (g2028) & (sk[2]) & (!g2843)) + ((!g2606) & (g2604) & (!g2028) & (!sk[2]) & (!g2843)) + ((!g2606) & (g2604) & (!g2028) & (!sk[2]) & (g2843)) + ((!g2606) & (g2604) & (!g2028) & (sk[2]) & (!g2843)) + ((!g2606) & (g2604) & (!g2028) & (sk[2]) & (g2843)) + ((!g2606) & (g2604) & (g2028) & (!sk[2]) & (!g2843)) + ((!g2606) & (g2604) & (g2028) & (!sk[2]) & (g2843)) + ((!g2606) & (g2604) & (g2028) & (sk[2]) & (!g2843)) + ((!g2606) & (g2604) & (g2028) & (sk[2]) & (g2843)) + ((g2606) & (!g2604) & (!g2028) & (!sk[2]) & (!g2843)) + ((g2606) & (!g2604) & (!g2028) & (!sk[2]) & (g2843)) + ((g2606) & (!g2604) & (!g2028) & (sk[2]) & (!g2843)) + ((g2606) & (!g2604) & (!g2028) & (sk[2]) & (g2843)) + ((g2606) & (!g2604) & (g2028) & (!sk[2]) & (!g2843)) + ((g2606) & (!g2604) & (g2028) & (!sk[2]) & (g2843)) + ((g2606) & (!g2604) & (g2028) & (sk[2]) & (!g2843)) + ((g2606) & (!g2604) & (g2028) & (sk[2]) & (g2843)) + ((g2606) & (g2604) & (!g2028) & (!sk[2]) & (!g2843)) + ((g2606) & (g2604) & (!g2028) & (!sk[2]) & (g2843)) + ((g2606) & (g2604) & (!g2028) & (sk[2]) & (!g2843)) + ((g2606) & (g2604) & (!g2028) & (sk[2]) & (g2843)) + ((g2606) & (g2604) & (g2028) & (!sk[2]) & (!g2843)) + ((g2606) & (g2604) & (g2028) & (!sk[2]) & (g2843)) + ((g2606) & (g2604) & (g2028) & (sk[2]) & (!g2843)) + ((g2606) & (g2604) & (g2028) & (sk[2]) & (g2843)));
	assign g3212 = (((!sk[3]) & (!g1837) & (g2843)) + ((!sk[3]) & (g1837) & (g2843)) + ((sk[3]) & (!g1837) & (!g2843)) + ((sk[3]) & (g1837) & (!g2843)) + ((sk[3]) & (g1837) & (g2843)));
	assign g3213 = (((!g3214) & (!sk[4]) & (g3215)) + ((!g3214) & (sk[4]) & (!g3215)) + ((g3214) & (!sk[4]) & (g3215)));
	assign g3214 = (((!g2584) & (!sk[5]) & (g3216)) + ((!g2584) & (sk[5]) & (g3216)) + ((g2584) & (!sk[5]) & (g3216)));
	assign g3215 = (((!g2584) & (!sk[6]) & (g3219)) + ((g2584) & (!sk[6]) & (g3219)) + ((g2584) & (sk[6]) & (g3219)));
	assign g3216 = (((!g3217) & (!sk[7]) & (g3218)) + ((!g3217) & (sk[7]) & (!g3218)) + ((g3217) & (!sk[7]) & (g3218)));
	assign g3217 = (((!sk[8]) & (!g2356) & (g3222)) + ((!sk[8]) & (g2356) & (g3222)) + ((sk[8]) & (!g2356) & (g3222)));
	assign g3218 = (((!sk[9]) & (!g2356) & (g3223)) + ((!sk[9]) & (g2356) & (g3223)) + ((sk[9]) & (g2356) & (g3223)));
	assign g3219 = (((!g3220) & (!sk[10]) & (g3221)) + ((!g3220) & (sk[10]) & (!g3221)) + ((g3220) & (!sk[10]) & (g3221)));
	assign g3220 = (((!sk[11]) & (!g2356) & (g3224)) + ((!sk[11]) & (g2356) & (g3224)) + ((sk[11]) & (!g2356) & (g3224)));
	assign g3221 = (((!g2356) & (!sk[12]) & (g3225)) + ((g2356) & (!sk[12]) & (g3225)) + ((g2356) & (sk[12]) & (g3225)));
	assign g3222 = (((!g2588) & (!g2586) & (!sk[13]) & (!g2028) & (g2843)) + ((!g2588) & (!g2586) & (!sk[13]) & (g2028) & (g2843)) + ((!g2588) & (g2586) & (!sk[13]) & (!g2028) & (!g2843)) + ((!g2588) & (g2586) & (!sk[13]) & (!g2028) & (g2843)) + ((!g2588) & (g2586) & (!sk[13]) & (g2028) & (!g2843)) + ((!g2588) & (g2586) & (!sk[13]) & (g2028) & (g2843)) + ((!g2588) & (g2586) & (sk[13]) & (g2028) & (g2843)) + ((g2588) & (!g2586) & (!sk[13]) & (!g2028) & (!g2843)) + ((g2588) & (!g2586) & (!sk[13]) & (!g2028) & (g2843)) + ((g2588) & (!g2586) & (!sk[13]) & (g2028) & (!g2843)) + ((g2588) & (!g2586) & (!sk[13]) & (g2028) & (g2843)) + ((g2588) & (!g2586) & (sk[13]) & (g2028) & (g2843)) + ((g2588) & (g2586) & (!sk[13]) & (!g2028) & (!g2843)) + ((g2588) & (g2586) & (!sk[13]) & (!g2028) & (g2843)) + ((g2588) & (g2586) & (!sk[13]) & (g2028) & (!g2843)) + ((g2588) & (g2586) & (!sk[13]) & (g2028) & (g2843)) + ((g2588) & (g2586) & (sk[13]) & (g2028) & (g2843)));
	assign g3223 = (((!g1824) & (!sk[14]) & (g2843)) + ((g1824) & (!sk[14]) & (g2843)) + ((g1824) & (sk[14]) & (g2843)));
	assign g3224 = (((!g2588) & (!g2586) & (!sk[15]) & (!g2028) & (g2843)) + ((!g2588) & (!g2586) & (!sk[15]) & (g2028) & (g2843)) + ((!g2588) & (!g2586) & (sk[15]) & (!g2028) & (!g2843)) + ((!g2588) & (!g2586) & (sk[15]) & (!g2028) & (g2843)) + ((!g2588) & (!g2586) & (sk[15]) & (g2028) & (!g2843)) + ((!g2588) & (g2586) & (!sk[15]) & (!g2028) & (!g2843)) + ((!g2588) & (g2586) & (!sk[15]) & (!g2028) & (g2843)) + ((!g2588) & (g2586) & (!sk[15]) & (g2028) & (!g2843)) + ((!g2588) & (g2586) & (!sk[15]) & (g2028) & (g2843)) + ((!g2588) & (g2586) & (sk[15]) & (!g2028) & (!g2843)) + ((!g2588) & (g2586) & (sk[15]) & (!g2028) & (g2843)) + ((!g2588) & (g2586) & (sk[15]) & (g2028) & (!g2843)) + ((!g2588) & (g2586) & (sk[15]) & (g2028) & (g2843)) + ((g2588) & (!g2586) & (!sk[15]) & (!g2028) & (!g2843)) + ((g2588) & (!g2586) & (!sk[15]) & (!g2028) & (g2843)) + ((g2588) & (!g2586) & (!sk[15]) & (g2028) & (!g2843)) + ((g2588) & (!g2586) & (!sk[15]) & (g2028) & (g2843)) + ((g2588) & (!g2586) & (sk[15]) & (!g2028) & (!g2843)) + ((g2588) & (!g2586) & (sk[15]) & (!g2028) & (g2843)) + ((g2588) & (!g2586) & (sk[15]) & (g2028) & (!g2843)) + ((g2588) & (!g2586) & (sk[15]) & (g2028) & (g2843)) + ((g2588) & (g2586) & (!sk[15]) & (!g2028) & (!g2843)) + ((g2588) & (g2586) & (!sk[15]) & (!g2028) & (g2843)) + ((g2588) & (g2586) & (!sk[15]) & (g2028) & (!g2843)) + ((g2588) & (g2586) & (!sk[15]) & (g2028) & (g2843)) + ((g2588) & (g2586) & (sk[15]) & (!g2028) & (!g2843)) + ((g2588) & (g2586) & (sk[15]) & (!g2028) & (g2843)) + ((g2588) & (g2586) & (sk[15]) & (g2028) & (!g2843)) + ((g2588) & (g2586) & (sk[15]) & (g2028) & (g2843)));
	assign g3225 = (((!g1824) & (!sk[16]) & (g2843)) + ((!g1824) & (sk[16]) & (!g2843)) + ((g1824) & (!sk[16]) & (g2843)) + ((g1824) & (sk[16]) & (!g2843)) + ((g1824) & (sk[16]) & (g2843)));
	assign g3226 = (((!g3227) & (!sk[17]) & (g3228)) + ((!g3227) & (sk[17]) & (!g3228)) + ((g3227) & (!sk[17]) & (g3228)));
	assign g3227 = (((!g2521) & (!sk[18]) & (g3229)) + ((!g2521) & (sk[18]) & (g3229)) + ((g2521) & (!sk[18]) & (g3229)));
	assign g3228 = (((!g2521) & (!sk[19]) & (g3232)) + ((g2521) & (!sk[19]) & (g3232)) + ((g2521) & (sk[19]) & (g3232)));
	assign g3229 = (((!g3230) & (!sk[20]) & (g3231)) + ((!g3230) & (sk[20]) & (!g3231)) + ((g3230) & (!sk[20]) & (g3231)));
	assign g3230 = (((!g2356) & (!sk[21]) & (g3235)) + ((!g2356) & (sk[21]) & (g3235)) + ((g2356) & (!sk[21]) & (g3235)));
	assign g3231 = (((!sk[22]) & (!g2356) & (g3236)) + ((!sk[22]) & (g2356) & (g3236)) + ((sk[22]) & (g2356) & (g3236)));
	assign g3232 = (((!sk[23]) & (!g3233) & (g3234)) + ((!sk[23]) & (g3233) & (g3234)) + ((sk[23]) & (!g3233) & (!g3234)));
	assign g3233 = (((!sk[24]) & (!g2356) & (g3237)) + ((!sk[24]) & (g2356) & (g3237)) + ((sk[24]) & (!g2356) & (g3237)));
	assign g3234 = (((!g2356) & (!sk[25]) & (g3238)) + ((g2356) & (!sk[25]) & (g3238)) + ((g2356) & (sk[25]) & (g3238)));
	assign g3235 = (((!sk[26]) & (!g2525) & (!g2522) & (!g2028) & (g2843)) + ((!sk[26]) & (!g2525) & (!g2522) & (g2028) & (g2843)) + ((!sk[26]) & (!g2525) & (g2522) & (!g2028) & (!g2843)) + ((!sk[26]) & (!g2525) & (g2522) & (!g2028) & (g2843)) + ((!sk[26]) & (!g2525) & (g2522) & (g2028) & (!g2843)) + ((!sk[26]) & (!g2525) & (g2522) & (g2028) & (g2843)) + ((!sk[26]) & (g2525) & (!g2522) & (!g2028) & (!g2843)) + ((!sk[26]) & (g2525) & (!g2522) & (!g2028) & (g2843)) + ((!sk[26]) & (g2525) & (!g2522) & (g2028) & (!g2843)) + ((!sk[26]) & (g2525) & (!g2522) & (g2028) & (g2843)) + ((!sk[26]) & (g2525) & (g2522) & (!g2028) & (!g2843)) + ((!sk[26]) & (g2525) & (g2522) & (!g2028) & (g2843)) + ((!sk[26]) & (g2525) & (g2522) & (g2028) & (!g2843)) + ((!sk[26]) & (g2525) & (g2522) & (g2028) & (g2843)) + ((sk[26]) & (!g2525) & (g2522) & (g2028) & (g2843)) + ((sk[26]) & (g2525) & (!g2522) & (g2028) & (g2843)) + ((sk[26]) & (g2525) & (g2522) & (g2028) & (g2843)));
	assign g3236 = (((!g1785) & (!sk[27]) & (g2843)) + ((g1785) & (!sk[27]) & (g2843)) + ((g1785) & (sk[27]) & (g2843)));
	assign g3237 = (((!g2525) & (!g2522) & (!sk[28]) & (!g2028) & (g2843)) + ((!g2525) & (!g2522) & (!sk[28]) & (g2028) & (g2843)) + ((!g2525) & (!g2522) & (sk[28]) & (!g2028) & (!g2843)) + ((!g2525) & (!g2522) & (sk[28]) & (!g2028) & (g2843)) + ((!g2525) & (!g2522) & (sk[28]) & (g2028) & (!g2843)) + ((!g2525) & (g2522) & (!sk[28]) & (!g2028) & (!g2843)) + ((!g2525) & (g2522) & (!sk[28]) & (!g2028) & (g2843)) + ((!g2525) & (g2522) & (!sk[28]) & (g2028) & (!g2843)) + ((!g2525) & (g2522) & (!sk[28]) & (g2028) & (g2843)) + ((!g2525) & (g2522) & (sk[28]) & (!g2028) & (!g2843)) + ((!g2525) & (g2522) & (sk[28]) & (!g2028) & (g2843)) + ((!g2525) & (g2522) & (sk[28]) & (g2028) & (!g2843)) + ((!g2525) & (g2522) & (sk[28]) & (g2028) & (g2843)) + ((g2525) & (!g2522) & (!sk[28]) & (!g2028) & (!g2843)) + ((g2525) & (!g2522) & (!sk[28]) & (!g2028) & (g2843)) + ((g2525) & (!g2522) & (!sk[28]) & (g2028) & (!g2843)) + ((g2525) & (!g2522) & (!sk[28]) & (g2028) & (g2843)) + ((g2525) & (!g2522) & (sk[28]) & (!g2028) & (!g2843)) + ((g2525) & (!g2522) & (sk[28]) & (!g2028) & (g2843)) + ((g2525) & (!g2522) & (sk[28]) & (g2028) & (!g2843)) + ((g2525) & (!g2522) & (sk[28]) & (g2028) & (g2843)) + ((g2525) & (g2522) & (!sk[28]) & (!g2028) & (!g2843)) + ((g2525) & (g2522) & (!sk[28]) & (!g2028) & (g2843)) + ((g2525) & (g2522) & (!sk[28]) & (g2028) & (!g2843)) + ((g2525) & (g2522) & (!sk[28]) & (g2028) & (g2843)) + ((g2525) & (g2522) & (sk[28]) & (!g2028) & (!g2843)) + ((g2525) & (g2522) & (sk[28]) & (!g2028) & (g2843)) + ((g2525) & (g2522) & (sk[28]) & (g2028) & (!g2843)) + ((g2525) & (g2522) & (sk[28]) & (g2028) & (g2843)));
	assign g3238 = (((!sk[29]) & (!g1785) & (g2843)) + ((!sk[29]) & (g1785) & (g2843)) + ((sk[29]) & (!g1785) & (!g2843)) + ((sk[29]) & (g1785) & (!g2843)) + ((sk[29]) & (g1785) & (g2843)));
	assign g3239 = (((!sk[30]) & (!g3240) & (g3241)) + ((!sk[30]) & (g3240) & (g3241)) + ((sk[30]) & (!g3240) & (!g3241)));
	assign g3240 = (((!sk[31]) & (!g2474) & (g3242)) + ((!sk[31]) & (g2474) & (g3242)) + ((sk[31]) & (!g2474) & (g3242)));
	assign g3241 = (((!g2474) & (!sk[32]) & (g3245)) + ((g2474) & (!sk[32]) & (g3245)) + ((g2474) & (sk[32]) & (g3245)));
	assign g3242 = (((!g3243) & (!sk[33]) & (g3244)) + ((!g3243) & (sk[33]) & (!g3244)) + ((g3243) & (!sk[33]) & (g3244)));
	assign g3243 = (((!sk[34]) & (!g2356) & (g3248)) + ((!sk[34]) & (g2356) & (g3248)) + ((sk[34]) & (!g2356) & (g3248)));
	assign g3244 = (((!g2356) & (!sk[35]) & (g3249)) + ((g2356) & (!sk[35]) & (g3249)) + ((g2356) & (sk[35]) & (g3249)));
	assign g3245 = (((!g3246) & (!sk[36]) & (g3247)) + ((!g3246) & (sk[36]) & (!g3247)) + ((g3246) & (!sk[36]) & (g3247)));
	assign g3246 = (((!sk[37]) & (!g2356) & (g3250)) + ((!sk[37]) & (g2356) & (g3250)) + ((sk[37]) & (!g2356) & (g3250)));
	assign g3247 = (((!g2356) & (!sk[38]) & (g3251)) + ((g2356) & (!sk[38]) & (g3251)) + ((g2356) & (sk[38]) & (g3251)));
	assign g3248 = (((!g2478) & (!sk[39]) & (!g2475) & (!g2028) & (g2843)) + ((!g2478) & (!sk[39]) & (!g2475) & (g2028) & (g2843)) + ((!g2478) & (!sk[39]) & (g2475) & (!g2028) & (!g2843)) + ((!g2478) & (!sk[39]) & (g2475) & (!g2028) & (g2843)) + ((!g2478) & (!sk[39]) & (g2475) & (g2028) & (!g2843)) + ((!g2478) & (!sk[39]) & (g2475) & (g2028) & (g2843)) + ((!g2478) & (sk[39]) & (g2475) & (g2028) & (g2843)) + ((g2478) & (!sk[39]) & (!g2475) & (!g2028) & (!g2843)) + ((g2478) & (!sk[39]) & (!g2475) & (!g2028) & (g2843)) + ((g2478) & (!sk[39]) & (!g2475) & (g2028) & (!g2843)) + ((g2478) & (!sk[39]) & (!g2475) & (g2028) & (g2843)) + ((g2478) & (!sk[39]) & (g2475) & (!g2028) & (!g2843)) + ((g2478) & (!sk[39]) & (g2475) & (!g2028) & (g2843)) + ((g2478) & (!sk[39]) & (g2475) & (g2028) & (!g2843)) + ((g2478) & (!sk[39]) & (g2475) & (g2028) & (g2843)) + ((g2478) & (sk[39]) & (!g2475) & (g2028) & (g2843)) + ((g2478) & (sk[39]) & (g2475) & (g2028) & (g2843)));
	assign g3249 = (((!sk[40]) & (!g1759) & (g2843)) + ((!sk[40]) & (g1759) & (g2843)) + ((sk[40]) & (g1759) & (g2843)));
	assign g3250 = (((!sk[41]) & (!g2478) & (!g2475) & (!g2028) & (g2843)) + ((!sk[41]) & (!g2478) & (!g2475) & (g2028) & (g2843)) + ((!sk[41]) & (!g2478) & (g2475) & (!g2028) & (!g2843)) + ((!sk[41]) & (!g2478) & (g2475) & (!g2028) & (g2843)) + ((!sk[41]) & (!g2478) & (g2475) & (g2028) & (!g2843)) + ((!sk[41]) & (!g2478) & (g2475) & (g2028) & (g2843)) + ((!sk[41]) & (g2478) & (!g2475) & (!g2028) & (!g2843)) + ((!sk[41]) & (g2478) & (!g2475) & (!g2028) & (g2843)) + ((!sk[41]) & (g2478) & (!g2475) & (g2028) & (!g2843)) + ((!sk[41]) & (g2478) & (!g2475) & (g2028) & (g2843)) + ((!sk[41]) & (g2478) & (g2475) & (!g2028) & (!g2843)) + ((!sk[41]) & (g2478) & (g2475) & (!g2028) & (g2843)) + ((!sk[41]) & (g2478) & (g2475) & (g2028) & (!g2843)) + ((!sk[41]) & (g2478) & (g2475) & (g2028) & (g2843)) + ((sk[41]) & (!g2478) & (!g2475) & (!g2028) & (!g2843)) + ((sk[41]) & (!g2478) & (!g2475) & (!g2028) & (g2843)) + ((sk[41]) & (!g2478) & (!g2475) & (g2028) & (!g2843)) + ((sk[41]) & (!g2478) & (g2475) & (!g2028) & (!g2843)) + ((sk[41]) & (!g2478) & (g2475) & (!g2028) & (g2843)) + ((sk[41]) & (!g2478) & (g2475) & (g2028) & (!g2843)) + ((sk[41]) & (!g2478) & (g2475) & (g2028) & (g2843)) + ((sk[41]) & (g2478) & (!g2475) & (!g2028) & (!g2843)) + ((sk[41]) & (g2478) & (!g2475) & (!g2028) & (g2843)) + ((sk[41]) & (g2478) & (!g2475) & (g2028) & (!g2843)) + ((sk[41]) & (g2478) & (!g2475) & (g2028) & (g2843)) + ((sk[41]) & (g2478) & (g2475) & (!g2028) & (!g2843)) + ((sk[41]) & (g2478) & (g2475) & (!g2028) & (g2843)) + ((sk[41]) & (g2478) & (g2475) & (g2028) & (!g2843)) + ((sk[41]) & (g2478) & (g2475) & (g2028) & (g2843)));
	assign g3251 = (((!sk[42]) & (!g1759) & (g2843)) + ((!sk[42]) & (g1759) & (g2843)) + ((sk[42]) & (!g1759) & (!g2843)) + ((sk[42]) & (g1759) & (!g2843)) + ((sk[42]) & (g1759) & (g2843)));
	assign g3252 = (((!g3253) & (!sk[43]) & (g3254)) + ((!g3253) & (sk[43]) & (!g3254)) + ((g3253) & (!sk[43]) & (g3254)));
	assign g3253 = (((!sk[44]) & (!g107) & (g3255)) + ((!sk[44]) & (g107) & (g3255)) + ((sk[44]) & (!g107) & (g3255)));
	assign g3254 = (((!sk[45]) & (!g107) & (g3258)) + ((!sk[45]) & (g107) & (g3258)) + ((sk[45]) & (g107) & (g3258)));
	assign g3255 = (((!sk[46]) & (!g3256) & (g3257)) + ((!sk[46]) & (g3256) & (g3257)) + ((sk[46]) & (!g3256) & (!g3257)));
	assign g3256 = (((!sk[47]) & (!g2034) & (g3261)) + ((!sk[47]) & (g2034) & (g3261)) + ((sk[47]) & (!g2034) & (g3261)));
	assign g3257 = (((!sk[48]) & (!g2034) & (g3262)) + ((!sk[48]) & (g2034) & (g3262)) + ((sk[48]) & (g2034) & (g3262)));
	assign g3258 = (((!g3259) & (!sk[49]) & (g3260)) + ((!g3259) & (sk[49]) & (!g3260)) + ((g3259) & (!sk[49]) & (g3260)));
	assign g3259 = (((!sk[50]) & (!g2034) & (g3263)) + ((!sk[50]) & (g2034) & (g3263)) + ((sk[50]) & (!g2034) & (g3263)));
	assign g3260 = (((!sk[51]) & (!g2034) & (g3264)) + ((!sk[51]) & (g2034) & (g3264)) + ((sk[51]) & (g2034) & (g3264)));
	assign g3261 = (((!sk[52]) & (!g2033) & (!g2823) & (!g2824) & (g1544)) + ((!sk[52]) & (!g2033) & (!g2823) & (g2824) & (g1544)) + ((!sk[52]) & (!g2033) & (g2823) & (!g2824) & (!g1544)) + ((!sk[52]) & (!g2033) & (g2823) & (!g2824) & (g1544)) + ((!sk[52]) & (!g2033) & (g2823) & (g2824) & (!g1544)) + ((!sk[52]) & (!g2033) & (g2823) & (g2824) & (g1544)) + ((!sk[52]) & (g2033) & (!g2823) & (!g2824) & (!g1544)) + ((!sk[52]) & (g2033) & (!g2823) & (!g2824) & (g1544)) + ((!sk[52]) & (g2033) & (!g2823) & (g2824) & (!g1544)) + ((!sk[52]) & (g2033) & (!g2823) & (g2824) & (g1544)) + ((!sk[52]) & (g2033) & (g2823) & (!g2824) & (!g1544)) + ((!sk[52]) & (g2033) & (g2823) & (!g2824) & (g1544)) + ((!sk[52]) & (g2033) & (g2823) & (g2824) & (!g1544)) + ((!sk[52]) & (g2033) & (g2823) & (g2824) & (g1544)) + ((sk[52]) & (!g2033) & (!g2823) & (g2824) & (!g1544)) + ((sk[52]) & (!g2033) & (!g2823) & (g2824) & (g1544)) + ((sk[52]) & (!g2033) & (g2823) & (g2824) & (!g1544)) + ((sk[52]) & (!g2033) & (g2823) & (g2824) & (g1544)) + ((sk[52]) & (g2033) & (!g2823) & (!g2824) & (g1544)) + ((sk[52]) & (g2033) & (!g2823) & (g2824) & (g1544)) + ((sk[52]) & (g2033) & (g2823) & (!g2824) & (!g1544)) + ((sk[52]) & (g2033) & (g2823) & (g2824) & (!g1544)));
	assign g3262 = (((!sk[53]) & (!g2033) & (g1994)) + ((!sk[53]) & (g2033) & (g1994)) + ((sk[53]) & (!g2033) & (g1994)));
	assign g3263 = (((!sk[54]) & (!g2033) & (!g2823) & (!g2824) & (g1544)) + ((!sk[54]) & (!g2033) & (!g2823) & (g2824) & (g1544)) + ((!sk[54]) & (!g2033) & (g2823) & (!g2824) & (!g1544)) + ((!sk[54]) & (!g2033) & (g2823) & (!g2824) & (g1544)) + ((!sk[54]) & (!g2033) & (g2823) & (g2824) & (!g1544)) + ((!sk[54]) & (!g2033) & (g2823) & (g2824) & (g1544)) + ((!sk[54]) & (g2033) & (!g2823) & (!g2824) & (!g1544)) + ((!sk[54]) & (g2033) & (!g2823) & (!g2824) & (g1544)) + ((!sk[54]) & (g2033) & (!g2823) & (g2824) & (!g1544)) + ((!sk[54]) & (g2033) & (!g2823) & (g2824) & (g1544)) + ((!sk[54]) & (g2033) & (g2823) & (!g2824) & (!g1544)) + ((!sk[54]) & (g2033) & (g2823) & (!g2824) & (g1544)) + ((!sk[54]) & (g2033) & (g2823) & (g2824) & (!g1544)) + ((!sk[54]) & (g2033) & (g2823) & (g2824) & (g1544)) + ((sk[54]) & (!g2033) & (!g2823) & (g2824) & (!g1544)) + ((sk[54]) & (!g2033) & (!g2823) & (g2824) & (g1544)) + ((sk[54]) & (!g2033) & (g2823) & (g2824) & (!g1544)) + ((sk[54]) & (!g2033) & (g2823) & (g2824) & (g1544)) + ((sk[54]) & (g2033) & (!g2823) & (!g2824) & (!g1544)) + ((sk[54]) & (g2033) & (!g2823) & (g2824) & (!g1544)) + ((sk[54]) & (g2033) & (g2823) & (!g2824) & (g1544)) + ((sk[54]) & (g2033) & (g2823) & (g2824) & (g1544)));
	assign g3264 = (((!sk[55]) & (!g2033) & (g1994)) + ((!sk[55]) & (g2033) & (g1994)) + ((sk[55]) & (!g2033) & (g1994)));
	assign g3265 = (((!sk[56]) & (!g3266) & (g3267)) + ((!sk[56]) & (g3266) & (g3267)) + ((sk[56]) & (!g3266) & (!g3267)));
	assign g3266 = (((!g2774) & (!sk[57]) & (g3268)) + ((!g2774) & (sk[57]) & (g3268)) + ((g2774) & (!sk[57]) & (g3268)));
	assign g3267 = (((!g2774) & (!sk[58]) & (g3271)) + ((g2774) & (!sk[58]) & (g3271)) + ((g2774) & (sk[58]) & (g3271)));
	assign g3268 = (((!g3269) & (!sk[59]) & (g3270)) + ((!g3269) & (sk[59]) & (!g3270)) + ((g3269) & (!sk[59]) & (g3270)));
	assign g3269 = (((!g2125) & (!sk[60]) & (g3274)) + ((!g2125) & (sk[60]) & (g3274)) + ((g2125) & (!sk[60]) & (g3274)));
	assign g3270 = (((!g2125) & (!sk[61]) & (g3275)) + ((g2125) & (!sk[61]) & (g3275)) + ((g2125) & (sk[61]) & (g3275)));
	assign g3271 = (((!sk[62]) & (!g3272) & (g3273)) + ((!sk[62]) & (g3272) & (g3273)) + ((sk[62]) & (!g3272) & (!g3273)));
	assign g3272 = (((!g2125) & (!sk[63]) & (g3276)) + ((!g2125) & (sk[63]) & (g3276)) + ((g2125) & (!sk[63]) & (g3276)));
	assign g3273 = (((!g2125) & (!sk[64]) & (g3277)) + ((g2125) & (!sk[64]) & (g3277)) + ((g2125) & (sk[64]) & (g3277)));
	assign g3274 = (((!g2771) & (!g2098) & (!sk[65]) & (!g2772) & (g2081)) + ((!g2771) & (!g2098) & (!sk[65]) & (g2772) & (g2081)) + ((!g2771) & (!g2098) & (sk[65]) & (g2772) & (!g2081)) + ((!g2771) & (g2098) & (!sk[65]) & (!g2772) & (!g2081)) + ((!g2771) & (g2098) & (!sk[65]) & (!g2772) & (g2081)) + ((!g2771) & (g2098) & (!sk[65]) & (g2772) & (!g2081)) + ((!g2771) & (g2098) & (!sk[65]) & (g2772) & (g2081)) + ((!g2771) & (g2098) & (sk[65]) & (!g2772) & (!g2081)) + ((g2771) & (!g2098) & (!sk[65]) & (!g2772) & (!g2081)) + ((g2771) & (!g2098) & (!sk[65]) & (!g2772) & (g2081)) + ((g2771) & (!g2098) & (!sk[65]) & (g2772) & (!g2081)) + ((g2771) & (!g2098) & (!sk[65]) & (g2772) & (g2081)) + ((g2771) & (!g2098) & (sk[65]) & (!g2772) & (!g2081)) + ((g2771) & (g2098) & (!sk[65]) & (!g2772) & (!g2081)) + ((g2771) & (g2098) & (!sk[65]) & (!g2772) & (g2081)) + ((g2771) & (g2098) & (!sk[65]) & (g2772) & (!g2081)) + ((g2771) & (g2098) & (!sk[65]) & (g2772) & (g2081)) + ((g2771) & (g2098) & (sk[65]) & (g2772) & (!g2081)));
	assign g3275 = (((!g2771) & (!sk[66]) & (!g2098) & (!g2777) & (g2081)) + ((!g2771) & (!sk[66]) & (!g2098) & (g2777) & (g2081)) + ((!g2771) & (!sk[66]) & (g2098) & (!g2777) & (!g2081)) + ((!g2771) & (!sk[66]) & (g2098) & (!g2777) & (g2081)) + ((!g2771) & (!sk[66]) & (g2098) & (g2777) & (!g2081)) + ((!g2771) & (!sk[66]) & (g2098) & (g2777) & (g2081)) + ((!g2771) & (sk[66]) & (!g2098) & (g2777) & (!g2081)) + ((!g2771) & (sk[66]) & (g2098) & (g2777) & (!g2081)) + ((g2771) & (!sk[66]) & (!g2098) & (!g2777) & (!g2081)) + ((g2771) & (!sk[66]) & (!g2098) & (!g2777) & (g2081)) + ((g2771) & (!sk[66]) & (!g2098) & (g2777) & (!g2081)) + ((g2771) & (!sk[66]) & (!g2098) & (g2777) & (g2081)) + ((g2771) & (!sk[66]) & (g2098) & (!g2777) & (!g2081)) + ((g2771) & (!sk[66]) & (g2098) & (!g2777) & (g2081)) + ((g2771) & (!sk[66]) & (g2098) & (g2777) & (!g2081)) + ((g2771) & (!sk[66]) & (g2098) & (g2777) & (g2081)) + ((g2771) & (sk[66]) & (!g2098) & (g2777) & (!g2081)) + ((g2771) & (sk[66]) & (g2098) & (!g2777) & (g2081)) + ((g2771) & (sk[66]) & (g2098) & (g2777) & (!g2081)) + ((g2771) & (sk[66]) & (g2098) & (g2777) & (g2081)));
	assign g3276 = (((!g2771) & (!g2098) & (!g2772) & (!sk[67]) & (g2081)) + ((!g2771) & (!g2098) & (!g2772) & (sk[67]) & (g2081)) + ((!g2771) & (!g2098) & (g2772) & (!sk[67]) & (g2081)) + ((!g2771) & (!g2098) & (g2772) & (sk[67]) & (!g2081)) + ((!g2771) & (!g2098) & (g2772) & (sk[67]) & (g2081)) + ((!g2771) & (g2098) & (!g2772) & (!sk[67]) & (!g2081)) + ((!g2771) & (g2098) & (!g2772) & (!sk[67]) & (g2081)) + ((!g2771) & (g2098) & (!g2772) & (sk[67]) & (!g2081)) + ((!g2771) & (g2098) & (!g2772) & (sk[67]) & (g2081)) + ((!g2771) & (g2098) & (g2772) & (!sk[67]) & (!g2081)) + ((!g2771) & (g2098) & (g2772) & (!sk[67]) & (g2081)) + ((!g2771) & (g2098) & (g2772) & (sk[67]) & (g2081)) + ((g2771) & (!g2098) & (!g2772) & (!sk[67]) & (!g2081)) + ((g2771) & (!g2098) & (!g2772) & (!sk[67]) & (g2081)) + ((g2771) & (!g2098) & (!g2772) & (sk[67]) & (!g2081)) + ((g2771) & (!g2098) & (!g2772) & (sk[67]) & (g2081)) + ((g2771) & (!g2098) & (g2772) & (!sk[67]) & (!g2081)) + ((g2771) & (!g2098) & (g2772) & (!sk[67]) & (g2081)) + ((g2771) & (!g2098) & (g2772) & (sk[67]) & (g2081)) + ((g2771) & (g2098) & (!g2772) & (!sk[67]) & (!g2081)) + ((g2771) & (g2098) & (!g2772) & (!sk[67]) & (g2081)) + ((g2771) & (g2098) & (!g2772) & (sk[67]) & (g2081)) + ((g2771) & (g2098) & (g2772) & (!sk[67]) & (!g2081)) + ((g2771) & (g2098) & (g2772) & (!sk[67]) & (g2081)) + ((g2771) & (g2098) & (g2772) & (sk[67]) & (!g2081)) + ((g2771) & (g2098) & (g2772) & (sk[67]) & (g2081)));
	assign g3277 = (((!sk[68]) & (!g2771) & (!g2098) & (!g2777) & (g2081)) + ((!sk[68]) & (!g2771) & (!g2098) & (g2777) & (g2081)) + ((!sk[68]) & (!g2771) & (g2098) & (!g2777) & (!g2081)) + ((!sk[68]) & (!g2771) & (g2098) & (!g2777) & (g2081)) + ((!sk[68]) & (!g2771) & (g2098) & (g2777) & (!g2081)) + ((!sk[68]) & (!g2771) & (g2098) & (g2777) & (g2081)) + ((!sk[68]) & (g2771) & (!g2098) & (!g2777) & (!g2081)) + ((!sk[68]) & (g2771) & (!g2098) & (!g2777) & (g2081)) + ((!sk[68]) & (g2771) & (!g2098) & (g2777) & (!g2081)) + ((!sk[68]) & (g2771) & (!g2098) & (g2777) & (g2081)) + ((!sk[68]) & (g2771) & (g2098) & (!g2777) & (!g2081)) + ((!sk[68]) & (g2771) & (g2098) & (!g2777) & (g2081)) + ((!sk[68]) & (g2771) & (g2098) & (g2777) & (!g2081)) + ((!sk[68]) & (g2771) & (g2098) & (g2777) & (g2081)) + ((sk[68]) & (!g2771) & (!g2098) & (g2777) & (!g2081)) + ((sk[68]) & (!g2771) & (g2098) & (g2777) & (!g2081)) + ((sk[68]) & (g2771) & (!g2098) & (g2777) & (!g2081)) + ((sk[68]) & (g2771) & (g2098) & (!g2777) & (g2081)) + ((sk[68]) & (g2771) & (g2098) & (g2777) & (!g2081)) + ((sk[68]) & (g2771) & (g2098) & (g2777) & (g2081)));
	assign g3278 = (((!g3279) & (!sk[69]) & (g3280)) + ((!g3279) & (sk[69]) & (!g3280)) + ((g3279) & (!sk[69]) & (g3280)));
	assign g3279 = (((!g75) & (!sk[70]) & (g3281)) + ((!g75) & (sk[70]) & (g3281)) + ((g75) & (!sk[70]) & (g3281)));
	assign g3280 = (((!sk[71]) & (!g75) & (g3284)) + ((!sk[71]) & (g75) & (g3284)) + ((sk[71]) & (g75) & (g3284)));
	assign g3281 = (((!g3282) & (!sk[72]) & (g3283)) + ((!g3282) & (sk[72]) & (!g3283)) + ((g3282) & (!sk[72]) & (g3283)));
	assign g3282 = (((!sk[73]) & (!g2280) & (g2763)) + ((!sk[73]) & (g2280) & (g2763)) + ((sk[73]) & (!g2280) & (g2763)));
	assign g3283 = (((!sk[74]) & (!g2091) & (g2280)) + ((!sk[74]) & (g2091) & (g2280)) + ((sk[74]) & (g2091) & (g2280)));
	assign g3284 = (((!sk[75]) & (!g3285) & (g3286)) + ((!sk[75]) & (g3285) & (g3286)) + ((sk[75]) & (!g3285) & (!g3286)));
	assign g3285 = (((!g2280) & (!sk[76]) & (g3287)) + ((!g2280) & (sk[76]) & (g3287)) + ((g2280) & (!sk[76]) & (g3287)));
	assign g3286 = (((!g2280) & (!sk[77]) & (g3288)) + ((g2280) & (!sk[77]) & (g3288)) + ((g2280) & (sk[77]) & (g3288)));
	assign g3287 = (((!dmem_dat_ix27x) & (!g2127) & (sk[78]) & (g2550)) + ((!dmem_dat_ix27x) & (g2127) & (!sk[78]) & (!g2550)) + ((!dmem_dat_ix27x) & (g2127) & (!sk[78]) & (g2550)) + ((!dmem_dat_ix27x) & (g2127) & (sk[78]) & (g2550)) + ((dmem_dat_ix27x) & (!g2127) & (!sk[78]) & (!g2550)) + ((dmem_dat_ix27x) & (!g2127) & (!sk[78]) & (g2550)) + ((dmem_dat_ix27x) & (!g2127) & (sk[78]) & (g2550)) + ((dmem_dat_ix27x) & (g2127) & (!sk[78]) & (!g2550)) + ((dmem_dat_ix27x) & (g2127) & (!sk[78]) & (g2550)) + ((dmem_dat_ix27x) & (g2127) & (sk[78]) & (!g2550)) + ((dmem_dat_ix27x) & (g2127) & (sk[78]) & (g2550)));
	assign g3288 = (((!sk[79]) & (!dmem_dat_ix27x) & (g2127) & (!g2550)) + ((!sk[79]) & (!dmem_dat_ix27x) & (g2127) & (g2550)) + ((!sk[79]) & (dmem_dat_ix27x) & (!g2127) & (!g2550)) + ((!sk[79]) & (dmem_dat_ix27x) & (!g2127) & (g2550)) + ((!sk[79]) & (dmem_dat_ix27x) & (g2127) & (!g2550)) + ((!sk[79]) & (dmem_dat_ix27x) & (g2127) & (g2550)) + ((sk[79]) & (!dmem_dat_ix27x) & (!g2127) & (g2550)) + ((sk[79]) & (!dmem_dat_ix27x) & (g2127) & (g2550)) + ((sk[79]) & (dmem_dat_ix27x) & (!g2127) & (g2550)) + ((sk[79]) & (dmem_dat_ix27x) & (g2127) & (!g2550)) + ((sk[79]) & (dmem_dat_ix27x) & (g2127) & (g2550)));
	assign g3289 = (((!g3290) & (!sk[80]) & (g3291)) + ((!g3290) & (sk[80]) & (!g3291)) + ((g3290) & (!sk[80]) & (g3291)));
	assign g3290 = (((!g2752) & (!sk[81]) & (g3292)) + ((!g2752) & (sk[81]) & (g3292)) + ((g2752) & (!sk[81]) & (g3292)));
	assign g3291 = (((!sk[82]) & (!g2752) & (g3295)) + ((!sk[82]) & (g2752) & (g3295)) + ((sk[82]) & (g2752) & (g3295)));
	assign g3292 = (((!g3293) & (!sk[83]) & (g3294)) + ((!g3293) & (sk[83]) & (!g3294)) + ((g3293) & (!sk[83]) & (g3294)));
	assign g3293 = (((!sk[84]) & (!g2125) & (g3298)) + ((!sk[84]) & (g2125) & (g3298)) + ((sk[84]) & (!g2125) & (g3298)));
	assign g3294 = (((!sk[85]) & (!g2125) & (g3299)) + ((!sk[85]) & (g2125) & (g3299)) + ((sk[85]) & (g2125) & (g3299)));
	assign g3295 = (((!sk[86]) & (!g3296) & (g3297)) + ((!sk[86]) & (g3296) & (g3297)) + ((sk[86]) & (!g3296) & (!g3297)));
	assign g3296 = (((!g2125) & (!sk[87]) & (g3300)) + ((!g2125) & (sk[87]) & (g3300)) + ((g2125) & (!sk[87]) & (g3300)));
	assign g3297 = (((!sk[88]) & (!g2125) & (g3301)) + ((!sk[88]) & (g2125) & (g3301)) + ((sk[88]) & (g2125) & (g3301)));
	assign g3298 = (((!g2738) & (!sk[89]) & (g2081) & (!g2737)) + ((!g2738) & (!sk[89]) & (g2081) & (g2737)) + ((g2738) & (!sk[89]) & (!g2081) & (!g2737)) + ((g2738) & (!sk[89]) & (!g2081) & (g2737)) + ((g2738) & (!sk[89]) & (g2081) & (!g2737)) + ((g2738) & (!sk[89]) & (g2081) & (g2737)) + ((g2738) & (sk[89]) & (g2081) & (g2737)));
	assign g3299 = (((!g2081) & (g2758) & (!sk[90]) & (!g2759)) + ((!g2081) & (g2758) & (!sk[90]) & (g2759)) + ((!g2081) & (g2758) & (sk[90]) & (!g2759)) + ((!g2081) & (g2758) & (sk[90]) & (g2759)) + ((g2081) & (!g2758) & (!sk[90]) & (!g2759)) + ((g2081) & (!g2758) & (!sk[90]) & (g2759)) + ((g2081) & (!g2758) & (sk[90]) & (g2759)) + ((g2081) & (g2758) & (!sk[90]) & (!g2759)) + ((g2081) & (g2758) & (!sk[90]) & (g2759)) + ((g2081) & (g2758) & (sk[90]) & (g2759)));
	assign g3300 = (((!g2738) & (!g2081) & (sk[91]) & (!g2737)) + ((!g2738) & (!g2081) & (sk[91]) & (g2737)) + ((!g2738) & (g2081) & (!sk[91]) & (!g2737)) + ((!g2738) & (g2081) & (!sk[91]) & (g2737)) + ((!g2738) & (g2081) & (sk[91]) & (!g2737)) + ((!g2738) & (g2081) & (sk[91]) & (g2737)) + ((g2738) & (!g2081) & (!sk[91]) & (!g2737)) + ((g2738) & (!g2081) & (!sk[91]) & (g2737)) + ((g2738) & (!g2081) & (sk[91]) & (!g2737)) + ((g2738) & (!g2081) & (sk[91]) & (g2737)) + ((g2738) & (g2081) & (!sk[91]) & (!g2737)) + ((g2738) & (g2081) & (!sk[91]) & (g2737)) + ((g2738) & (g2081) & (sk[91]) & (!g2737)));
	assign g3301 = (((!g2081) & (!sk[92]) & (g2758) & (!g2759)) + ((!g2081) & (!sk[92]) & (g2758) & (g2759)) + ((!g2081) & (sk[92]) & (g2758) & (!g2759)) + ((!g2081) & (sk[92]) & (g2758) & (g2759)) + ((g2081) & (!sk[92]) & (!g2758) & (!g2759)) + ((g2081) & (!sk[92]) & (!g2758) & (g2759)) + ((g2081) & (!sk[92]) & (g2758) & (!g2759)) + ((g2081) & (!sk[92]) & (g2758) & (g2759)) + ((g2081) & (sk[92]) & (!g2758) & (g2759)) + ((g2081) & (sk[92]) & (g2758) & (g2759)));
	assign g3302 = (((!g3303) & (!sk[93]) & (g3304)) + ((!g3303) & (sk[93]) & (!g3304)) + ((g3303) & (!sk[93]) & (g3304)));
	assign g3303 = (((!g75) & (!sk[94]) & (g3305)) + ((!g75) & (sk[94]) & (g3305)) + ((g75) & (!sk[94]) & (g3305)));
	assign g3304 = (((!sk[95]) & (!g75) & (g3308)) + ((!sk[95]) & (g75) & (g3308)) + ((sk[95]) & (g75) & (g3308)));
	assign g3305 = (((!g3306) & (!sk[96]) & (g3307)) + ((!g3306) & (sk[96]) & (!g3307)) + ((g3306) & (!sk[96]) & (g3307)));
	assign g3306 = (((!sk[97]) & (!g2280) & (g2745)) + ((!sk[97]) & (g2280) & (g2745)) + ((sk[97]) & (!g2280) & (g2745)));
	assign g3307 = (((!g2090) & (!sk[98]) & (g2280)) + ((g2090) & (!sk[98]) & (g2280)) + ((g2090) & (sk[98]) & (g2280)));
	assign g3308 = (((!g3309) & (!sk[99]) & (g3310)) + ((!g3309) & (sk[99]) & (!g3310)) + ((g3309) & (!sk[99]) & (g3310)));
	assign g3309 = (((!g2280) & (!sk[100]) & (g3311)) + ((!g2280) & (sk[100]) & (g3311)) + ((g2280) & (!sk[100]) & (g3311)));
	assign g3310 = (((!sk[101]) & (!g2280) & (g3312)) + ((!sk[101]) & (g2280) & (g3312)) + ((sk[101]) & (g2280) & (g3312)));
	assign g3311 = (((!sk[102]) & (!dmem_dat_ix26x) & (g2127) & (!g2550)) + ((!sk[102]) & (!dmem_dat_ix26x) & (g2127) & (g2550)) + ((!sk[102]) & (dmem_dat_ix26x) & (!g2127) & (!g2550)) + ((!sk[102]) & (dmem_dat_ix26x) & (!g2127) & (g2550)) + ((!sk[102]) & (dmem_dat_ix26x) & (g2127) & (!g2550)) + ((!sk[102]) & (dmem_dat_ix26x) & (g2127) & (g2550)) + ((sk[102]) & (!dmem_dat_ix26x) & (!g2127) & (g2550)) + ((sk[102]) & (!dmem_dat_ix26x) & (g2127) & (g2550)) + ((sk[102]) & (dmem_dat_ix26x) & (!g2127) & (g2550)) + ((sk[102]) & (dmem_dat_ix26x) & (g2127) & (!g2550)) + ((sk[102]) & (dmem_dat_ix26x) & (g2127) & (g2550)));
	assign g3312 = (((!dmem_dat_ix26x) & (!g2127) & (sk[103]) & (g2550)) + ((!dmem_dat_ix26x) & (g2127) & (!sk[103]) & (!g2550)) + ((!dmem_dat_ix26x) & (g2127) & (!sk[103]) & (g2550)) + ((!dmem_dat_ix26x) & (g2127) & (sk[103]) & (g2550)) + ((dmem_dat_ix26x) & (!g2127) & (!sk[103]) & (!g2550)) + ((dmem_dat_ix26x) & (!g2127) & (!sk[103]) & (g2550)) + ((dmem_dat_ix26x) & (!g2127) & (sk[103]) & (g2550)) + ((dmem_dat_ix26x) & (g2127) & (!sk[103]) & (!g2550)) + ((dmem_dat_ix26x) & (g2127) & (!sk[103]) & (g2550)) + ((dmem_dat_ix26x) & (g2127) & (sk[103]) & (!g2550)) + ((dmem_dat_ix26x) & (g2127) & (sk[103]) & (g2550)));
	assign g3313 = (((!sk[104]) & (!g3314) & (g3315)) + ((!sk[104]) & (g3314) & (g3315)) + ((sk[104]) & (!g3314) & (!g3315)));
	assign g3314 = (((!g2738) & (!sk[105]) & (g3316)) + ((!g2738) & (sk[105]) & (g3316)) + ((g2738) & (!sk[105]) & (g3316)));
	assign g3315 = (((!sk[106]) & (!g2738) & (g3319)) + ((!sk[106]) & (g2738) & (g3319)) + ((sk[106]) & (g2738) & (g3319)));
	assign g3316 = (((!g3317) & (!sk[107]) & (g3318)) + ((!g3317) & (sk[107]) & (!g3318)) + ((g3317) & (!sk[107]) & (g3318)));
	assign g3317 = (((!g2125) & (!sk[108]) & (g2737)) + ((!g2125) & (sk[108]) & (g2737)) + ((g2125) & (!sk[108]) & (g2737)));
	assign g3318 = (((!g2125) & (!sk[109]) & (g3322)) + ((g2125) & (!sk[109]) & (g3322)) + ((g2125) & (sk[109]) & (g3322)));
	assign g3319 = (((!sk[110]) & (!g3320) & (g3321)) + ((!sk[110]) & (g3320) & (g3321)) + ((sk[110]) & (!g3320) & (!g3321)));
	assign g3320 = (((!g2125) & (!sk[111]) & (g3323)) + ((!g2125) & (sk[111]) & (g3323)) + ((g2125) & (!sk[111]) & (g3323)));
	assign g3321 = (((!sk[112]) & (!g2125) & (g3324)) + ((!sk[112]) & (g2125) & (g3324)) + ((sk[112]) & (g2125) & (g3324)));
	assign g3322 = (((!g2734) & (!sk[113]) & (!g2081) & (!g2090) & (g2741)) + ((!g2734) & (!sk[113]) & (!g2081) & (g2090) & (g2741)) + ((!g2734) & (!sk[113]) & (g2081) & (!g2090) & (!g2741)) + ((!g2734) & (!sk[113]) & (g2081) & (!g2090) & (g2741)) + ((!g2734) & (!sk[113]) & (g2081) & (g2090) & (!g2741)) + ((!g2734) & (!sk[113]) & (g2081) & (g2090) & (g2741)) + ((!g2734) & (sk[113]) & (!g2081) & (!g2090) & (g2741)) + ((!g2734) & (sk[113]) & (!g2081) & (g2090) & (g2741)) + ((g2734) & (!sk[113]) & (!g2081) & (!g2090) & (!g2741)) + ((g2734) & (!sk[113]) & (!g2081) & (!g2090) & (g2741)) + ((g2734) & (!sk[113]) & (!g2081) & (g2090) & (!g2741)) + ((g2734) & (!sk[113]) & (!g2081) & (g2090) & (g2741)) + ((g2734) & (!sk[113]) & (g2081) & (!g2090) & (!g2741)) + ((g2734) & (!sk[113]) & (g2081) & (!g2090) & (g2741)) + ((g2734) & (!sk[113]) & (g2081) & (g2090) & (!g2741)) + ((g2734) & (!sk[113]) & (g2081) & (g2090) & (g2741)) + ((g2734) & (sk[113]) & (!g2081) & (!g2090) & (g2741)) + ((g2734) & (sk[113]) & (!g2081) & (g2090) & (g2741)) + ((g2734) & (sk[113]) & (g2081) & (g2090) & (!g2741)) + ((g2734) & (sk[113]) & (g2081) & (g2090) & (g2741)));
	assign g3323 = (((!sk[114]) & (!g2081) & (g2737)) + ((!sk[114]) & (g2081) & (g2737)) + ((sk[114]) & (!g2081) & (g2737)) + ((sk[114]) & (g2081) & (!g2737)));
	assign g3324 = (((!g2734) & (!g2081) & (!g2090) & (!sk[115]) & (g2741)) + ((!g2734) & (!g2081) & (!g2090) & (sk[115]) & (g2741)) + ((!g2734) & (!g2081) & (g2090) & (!sk[115]) & (g2741)) + ((!g2734) & (!g2081) & (g2090) & (sk[115]) & (g2741)) + ((!g2734) & (g2081) & (!g2090) & (!sk[115]) & (!g2741)) + ((!g2734) & (g2081) & (!g2090) & (!sk[115]) & (g2741)) + ((!g2734) & (g2081) & (g2090) & (!sk[115]) & (!g2741)) + ((!g2734) & (g2081) & (g2090) & (!sk[115]) & (g2741)) + ((g2734) & (!g2081) & (!g2090) & (!sk[115]) & (!g2741)) + ((g2734) & (!g2081) & (!g2090) & (!sk[115]) & (g2741)) + ((g2734) & (!g2081) & (!g2090) & (sk[115]) & (g2741)) + ((g2734) & (!g2081) & (g2090) & (!sk[115]) & (!g2741)) + ((g2734) & (!g2081) & (g2090) & (!sk[115]) & (g2741)) + ((g2734) & (!g2081) & (g2090) & (sk[115]) & (g2741)) + ((g2734) & (g2081) & (!g2090) & (!sk[115]) & (!g2741)) + ((g2734) & (g2081) & (!g2090) & (!sk[115]) & (g2741)) + ((g2734) & (g2081) & (g2090) & (!sk[115]) & (!g2741)) + ((g2734) & (g2081) & (g2090) & (!sk[115]) & (g2741)) + ((g2734) & (g2081) & (g2090) & (sk[115]) & (!g2741)) + ((g2734) & (g2081) & (g2090) & (sk[115]) & (g2741)));
	assign g3325 = (((!sk[116]) & (!g3326) & (g3327)) + ((!sk[116]) & (g3326) & (g3327)) + ((sk[116]) & (!g3326) & (!g3327)));
	assign g3326 = (((!g75) & (!sk[117]) & (g3328)) + ((!g75) & (sk[117]) & (g3328)) + ((g75) & (!sk[117]) & (g3328)));
	assign g3327 = (((!sk[118]) & (!g75) & (g3331)) + ((!sk[118]) & (g75) & (g3331)) + ((sk[118]) & (g75) & (g3331)));
	assign g3328 = (((!g3329) & (!sk[119]) & (g3330)) + ((!g3329) & (sk[119]) & (!g3330)) + ((g3329) & (!sk[119]) & (g3330)));
	assign g3329 = (((!sk[120]) & (!g2280) & (g2726)) + ((!sk[120]) & (g2280) & (g2726)) + ((sk[120]) & (!g2280) & (g2726)));
	assign g3330 = (((!sk[121]) & (!g2089) & (g2280)) + ((!sk[121]) & (g2089) & (g2280)) + ((sk[121]) & (g2089) & (g2280)));
	assign g3331 = (((!g3332) & (!sk[122]) & (g3333)) + ((!g3332) & (sk[122]) & (!g3333)) + ((g3332) & (!sk[122]) & (g3333)));
	assign g3332 = (((!g2280) & (!sk[123]) & (g3334)) + ((!g2280) & (sk[123]) & (g3334)) + ((g2280) & (!sk[123]) & (g3334)));
	assign g3333 = (((!g2280) & (!sk[124]) & (g3335)) + ((g2280) & (!sk[124]) & (g3335)) + ((g2280) & (sk[124]) & (g3335)));
	assign g3334 = (((!dmem_dat_ix25x) & (!g2127) & (sk[125]) & (g2550)) + ((!dmem_dat_ix25x) & (g2127) & (!sk[125]) & (!g2550)) + ((!dmem_dat_ix25x) & (g2127) & (!sk[125]) & (g2550)) + ((!dmem_dat_ix25x) & (g2127) & (sk[125]) & (g2550)) + ((dmem_dat_ix25x) & (!g2127) & (!sk[125]) & (!g2550)) + ((dmem_dat_ix25x) & (!g2127) & (!sk[125]) & (g2550)) + ((dmem_dat_ix25x) & (!g2127) & (sk[125]) & (g2550)) + ((dmem_dat_ix25x) & (g2127) & (!sk[125]) & (!g2550)) + ((dmem_dat_ix25x) & (g2127) & (!sk[125]) & (g2550)) + ((dmem_dat_ix25x) & (g2127) & (sk[125]) & (!g2550)) + ((dmem_dat_ix25x) & (g2127) & (sk[125]) & (g2550)));
	assign g3335 = (((!dmem_dat_ix25x) & (!sk[126]) & (g2127) & (!g2550)) + ((!dmem_dat_ix25x) & (!sk[126]) & (g2127) & (g2550)) + ((!dmem_dat_ix25x) & (sk[126]) & (!g2127) & (g2550)) + ((!dmem_dat_ix25x) & (sk[126]) & (g2127) & (g2550)) + ((dmem_dat_ix25x) & (!sk[126]) & (!g2127) & (!g2550)) + ((dmem_dat_ix25x) & (!sk[126]) & (!g2127) & (g2550)) + ((dmem_dat_ix25x) & (!sk[126]) & (g2127) & (!g2550)) + ((dmem_dat_ix25x) & (!sk[126]) & (g2127) & (g2550)) + ((dmem_dat_ix25x) & (sk[126]) & (!g2127) & (g2550)) + ((dmem_dat_ix25x) & (sk[126]) & (g2127) & (!g2550)) + ((dmem_dat_ix25x) & (sk[126]) & (g2127) & (g2550)));
	assign g3336 = (((!g3337) & (!sk[127]) & (g3338)) + ((!g3337) & (sk[127]) & (!g3338)) + ((g3337) & (!sk[127]) & (g3338)));
	assign g3337 = (((!g2718) & (!sk[0]) & (g3339)) + ((!g2718) & (sk[0]) & (g3339)) + ((g2718) & (!sk[0]) & (g3339)));
	assign g3338 = (((!g2718) & (!sk[1]) & (g3342)) + ((g2718) & (!sk[1]) & (g3342)) + ((g2718) & (sk[1]) & (g3342)));
	assign g3339 = (((!g3340) & (!sk[2]) & (g3341)) + ((!g3340) & (sk[2]) & (!g3341)) + ((g3340) & (!sk[2]) & (g3341)));
	assign g3340 = (((!sk[3]) & (!g2125) & (g3345)) + ((!sk[3]) & (g2125) & (g3345)) + ((sk[3]) & (!g2125) & (g3345)));
	assign g3341 = (((!g2125) & (!sk[4]) & (g3346)) + ((g2125) & (!sk[4]) & (g3346)) + ((g2125) & (sk[4]) & (g3346)));
	assign g3342 = (((!g3343) & (!sk[5]) & (g3344)) + ((!g3343) & (sk[5]) & (!g3344)) + ((g3343) & (!sk[5]) & (g3344)));
	assign g3343 = (((!g2125) & (!sk[6]) & (g3347)) + ((!g2125) & (sk[6]) & (g3347)) + ((g2125) & (!sk[6]) & (g3347)));
	assign g3344 = (((!sk[7]) & (!g2125) & (g3348)) + ((!sk[7]) & (g2125) & (g3348)) + ((sk[7]) & (g2125) & (g3348)));
	assign g3345 = (((!sk[8]) & (!g2081) & (g2717)) + ((!sk[8]) & (g2081) & (g2717)) + ((sk[8]) & (!g2081) & (g2717)));
	assign g3346 = (((!g2715) & (!g2081) & (!sk[9]) & (!g2089) & (g2722)) + ((!g2715) & (!g2081) & (!sk[9]) & (g2089) & (g2722)) + ((!g2715) & (!g2081) & (sk[9]) & (!g2089) & (g2722)) + ((!g2715) & (!g2081) & (sk[9]) & (g2089) & (g2722)) + ((!g2715) & (g2081) & (!sk[9]) & (!g2089) & (!g2722)) + ((!g2715) & (g2081) & (!sk[9]) & (!g2089) & (g2722)) + ((!g2715) & (g2081) & (!sk[9]) & (g2089) & (!g2722)) + ((!g2715) & (g2081) & (!sk[9]) & (g2089) & (g2722)) + ((g2715) & (!g2081) & (!sk[9]) & (!g2089) & (!g2722)) + ((g2715) & (!g2081) & (!sk[9]) & (!g2089) & (g2722)) + ((g2715) & (!g2081) & (!sk[9]) & (g2089) & (!g2722)) + ((g2715) & (!g2081) & (!sk[9]) & (g2089) & (g2722)) + ((g2715) & (!g2081) & (sk[9]) & (!g2089) & (g2722)) + ((g2715) & (!g2081) & (sk[9]) & (g2089) & (g2722)) + ((g2715) & (g2081) & (!sk[9]) & (!g2089) & (!g2722)) + ((g2715) & (g2081) & (!sk[9]) & (!g2089) & (g2722)) + ((g2715) & (g2081) & (!sk[9]) & (g2089) & (!g2722)) + ((g2715) & (g2081) & (!sk[9]) & (g2089) & (g2722)) + ((g2715) & (g2081) & (sk[9]) & (g2089) & (!g2722)) + ((g2715) & (g2081) & (sk[9]) & (g2089) & (g2722)));
	assign g3347 = (((!g2081) & (!sk[10]) & (g2717)) + ((!g2081) & (sk[10]) & (g2717)) + ((g2081) & (!sk[10]) & (g2717)) + ((g2081) & (sk[10]) & (!g2717)) + ((g2081) & (sk[10]) & (g2717)));
	assign g3348 = (((!g2715) & (!g2081) & (!sk[11]) & (!g2089) & (g2722)) + ((!g2715) & (!g2081) & (!sk[11]) & (g2089) & (g2722)) + ((!g2715) & (!g2081) & (sk[11]) & (!g2089) & (g2722)) + ((!g2715) & (!g2081) & (sk[11]) & (g2089) & (g2722)) + ((!g2715) & (g2081) & (!sk[11]) & (!g2089) & (!g2722)) + ((!g2715) & (g2081) & (!sk[11]) & (!g2089) & (g2722)) + ((!g2715) & (g2081) & (!sk[11]) & (g2089) & (!g2722)) + ((!g2715) & (g2081) & (!sk[11]) & (g2089) & (g2722)) + ((g2715) & (!g2081) & (!sk[11]) & (!g2089) & (!g2722)) + ((g2715) & (!g2081) & (!sk[11]) & (!g2089) & (g2722)) + ((g2715) & (!g2081) & (!sk[11]) & (g2089) & (!g2722)) + ((g2715) & (!g2081) & (!sk[11]) & (g2089) & (g2722)) + ((g2715) & (!g2081) & (sk[11]) & (!g2089) & (g2722)) + ((g2715) & (!g2081) & (sk[11]) & (g2089) & (g2722)) + ((g2715) & (g2081) & (!sk[11]) & (!g2089) & (!g2722)) + ((g2715) & (g2081) & (!sk[11]) & (!g2089) & (g2722)) + ((g2715) & (g2081) & (!sk[11]) & (g2089) & (!g2722)) + ((g2715) & (g2081) & (!sk[11]) & (g2089) & (g2722)) + ((g2715) & (g2081) & (sk[11]) & (g2089) & (!g2722)) + ((g2715) & (g2081) & (sk[11]) & (g2089) & (g2722)));
	assign g3349 = (((!g3350) & (!sk[12]) & (g3351)) + ((!g3350) & (sk[12]) & (!g3351)) + ((g3350) & (!sk[12]) & (g3351)));
	assign g3350 = (((!g75) & (!sk[13]) & (g3352)) + ((!g75) & (sk[13]) & (g3352)) + ((g75) & (!sk[13]) & (g3352)));
	assign g3351 = (((!sk[14]) & (!g75) & (g3355)) + ((!sk[14]) & (g75) & (g3355)) + ((sk[14]) & (g75) & (g3355)));
	assign g3352 = (((!g3353) & (!sk[15]) & (g3354)) + ((!g3353) & (sk[15]) & (!g3354)) + ((g3353) & (!sk[15]) & (g3354)));
	assign g3353 = (((!g2280) & (!sk[16]) & (g2709)) + ((!g2280) & (sk[16]) & (g2709)) + ((g2280) & (!sk[16]) & (g2709)));
	assign g3354 = (((!sk[17]) & (!g2088) & (g2280)) + ((!sk[17]) & (g2088) & (g2280)) + ((sk[17]) & (g2088) & (g2280)));
	assign g3355 = (((!g3356) & (!sk[18]) & (g3357)) + ((!g3356) & (sk[18]) & (!g3357)) + ((g3356) & (!sk[18]) & (g3357)));
	assign g3356 = (((!sk[19]) & (!g2280) & (g3358)) + ((!sk[19]) & (g2280) & (g3358)) + ((sk[19]) & (!g2280) & (g3358)));
	assign g3357 = (((!g2280) & (!sk[20]) & (g3359)) + ((g2280) & (!sk[20]) & (g3359)) + ((g2280) & (sk[20]) & (g3359)));
	assign g3358 = (((!sk[21]) & (!dmem_dat_ix24x) & (g2127) & (!g2550)) + ((!sk[21]) & (!dmem_dat_ix24x) & (g2127) & (g2550)) + ((!sk[21]) & (dmem_dat_ix24x) & (!g2127) & (!g2550)) + ((!sk[21]) & (dmem_dat_ix24x) & (!g2127) & (g2550)) + ((!sk[21]) & (dmem_dat_ix24x) & (g2127) & (!g2550)) + ((!sk[21]) & (dmem_dat_ix24x) & (g2127) & (g2550)) + ((sk[21]) & (!dmem_dat_ix24x) & (!g2127) & (g2550)) + ((sk[21]) & (!dmem_dat_ix24x) & (g2127) & (g2550)) + ((sk[21]) & (dmem_dat_ix24x) & (!g2127) & (g2550)) + ((sk[21]) & (dmem_dat_ix24x) & (g2127) & (!g2550)) + ((sk[21]) & (dmem_dat_ix24x) & (g2127) & (g2550)));
	assign g3359 = (((!sk[22]) & (!dmem_dat_ix24x) & (g2127) & (!g2550)) + ((!sk[22]) & (!dmem_dat_ix24x) & (g2127) & (g2550)) + ((!sk[22]) & (dmem_dat_ix24x) & (!g2127) & (!g2550)) + ((!sk[22]) & (dmem_dat_ix24x) & (!g2127) & (g2550)) + ((!sk[22]) & (dmem_dat_ix24x) & (g2127) & (!g2550)) + ((!sk[22]) & (dmem_dat_ix24x) & (g2127) & (g2550)) + ((sk[22]) & (!dmem_dat_ix24x) & (!g2127) & (g2550)) + ((sk[22]) & (!dmem_dat_ix24x) & (g2127) & (g2550)) + ((sk[22]) & (dmem_dat_ix24x) & (!g2127) & (g2550)) + ((sk[22]) & (dmem_dat_ix24x) & (g2127) & (!g2550)) + ((sk[22]) & (dmem_dat_ix24x) & (g2127) & (g2550)));
	assign g3360 = (((!sk[23]) & (!g3361) & (g3362)) + ((!sk[23]) & (g3361) & (g3362)) + ((sk[23]) & (!g3361) & (!g3362)));
	assign g3361 = (((!g2701) & (!sk[24]) & (g3363)) + ((!g2701) & (sk[24]) & (g3363)) + ((g2701) & (!sk[24]) & (g3363)));
	assign g3362 = (((!sk[25]) & (!g2701) & (g3366)) + ((!sk[25]) & (g2701) & (g3366)) + ((sk[25]) & (g2701) & (g3366)));
	assign g3363 = (((!sk[26]) & (!g3364) & (g3365)) + ((!sk[26]) & (g3364) & (g3365)) + ((sk[26]) & (!g3364) & (!g3365)));
	assign g3364 = (((!sk[27]) & (!g2125) & (g3369)) + ((!sk[27]) & (g2125) & (g3369)) + ((sk[27]) & (!g2125) & (g3369)));
	assign g3365 = (((!g2125) & (!sk[28]) & (g3370)) + ((g2125) & (!sk[28]) & (g3370)) + ((g2125) & (sk[28]) & (g3370)));
	assign g3366 = (((!sk[29]) & (!g3367) & (g3368)) + ((!sk[29]) & (g3367) & (g3368)) + ((sk[29]) & (!g3367) & (!g3368)));
	assign g3367 = (((!g2125) & (!sk[30]) & (g3371)) + ((!g2125) & (sk[30]) & (g3371)) + ((g2125) & (!sk[30]) & (g3371)));
	assign g3368 = (((!sk[31]) & (!g2125) & (g3372)) + ((!sk[31]) & (g2125) & (g3372)) + ((sk[31]) & (g2125) & (g3372)));
	assign g3369 = (((!sk[32]) & (!g2081) & (g2700)) + ((!sk[32]) & (g2081) & (g2700)) + ((sk[32]) & (!g2081) & (g2700)));
	assign g3370 = (((!g2699) & (!sk[33]) & (!g2081) & (!g2088) & (g2705)) + ((!g2699) & (!sk[33]) & (!g2081) & (g2088) & (g2705)) + ((!g2699) & (!sk[33]) & (g2081) & (!g2088) & (!g2705)) + ((!g2699) & (!sk[33]) & (g2081) & (!g2088) & (g2705)) + ((!g2699) & (!sk[33]) & (g2081) & (g2088) & (!g2705)) + ((!g2699) & (!sk[33]) & (g2081) & (g2088) & (g2705)) + ((!g2699) & (sk[33]) & (!g2081) & (!g2088) & (g2705)) + ((!g2699) & (sk[33]) & (!g2081) & (g2088) & (g2705)) + ((g2699) & (!sk[33]) & (!g2081) & (!g2088) & (!g2705)) + ((g2699) & (!sk[33]) & (!g2081) & (!g2088) & (g2705)) + ((g2699) & (!sk[33]) & (!g2081) & (g2088) & (!g2705)) + ((g2699) & (!sk[33]) & (!g2081) & (g2088) & (g2705)) + ((g2699) & (!sk[33]) & (g2081) & (!g2088) & (!g2705)) + ((g2699) & (!sk[33]) & (g2081) & (!g2088) & (g2705)) + ((g2699) & (!sk[33]) & (g2081) & (g2088) & (!g2705)) + ((g2699) & (!sk[33]) & (g2081) & (g2088) & (g2705)) + ((g2699) & (sk[33]) & (!g2081) & (!g2088) & (g2705)) + ((g2699) & (sk[33]) & (!g2081) & (g2088) & (g2705)) + ((g2699) & (sk[33]) & (g2081) & (g2088) & (!g2705)) + ((g2699) & (sk[33]) & (g2081) & (g2088) & (g2705)));
	assign g3371 = (((!sk[34]) & (!g2081) & (g2700)) + ((!sk[34]) & (g2081) & (g2700)) + ((sk[34]) & (!g2081) & (g2700)) + ((sk[34]) & (g2081) & (!g2700)) + ((sk[34]) & (g2081) & (g2700)));
	assign g3372 = (((!g2699) & (!g2081) & (!sk[35]) & (!g2088) & (g2705)) + ((!g2699) & (!g2081) & (!sk[35]) & (g2088) & (g2705)) + ((!g2699) & (!g2081) & (sk[35]) & (!g2088) & (g2705)) + ((!g2699) & (!g2081) & (sk[35]) & (g2088) & (g2705)) + ((!g2699) & (g2081) & (!sk[35]) & (!g2088) & (!g2705)) + ((!g2699) & (g2081) & (!sk[35]) & (!g2088) & (g2705)) + ((!g2699) & (g2081) & (!sk[35]) & (g2088) & (!g2705)) + ((!g2699) & (g2081) & (!sk[35]) & (g2088) & (g2705)) + ((g2699) & (!g2081) & (!sk[35]) & (!g2088) & (!g2705)) + ((g2699) & (!g2081) & (!sk[35]) & (!g2088) & (g2705)) + ((g2699) & (!g2081) & (!sk[35]) & (g2088) & (!g2705)) + ((g2699) & (!g2081) & (!sk[35]) & (g2088) & (g2705)) + ((g2699) & (!g2081) & (sk[35]) & (!g2088) & (g2705)) + ((g2699) & (!g2081) & (sk[35]) & (g2088) & (g2705)) + ((g2699) & (g2081) & (!sk[35]) & (!g2088) & (!g2705)) + ((g2699) & (g2081) & (!sk[35]) & (!g2088) & (g2705)) + ((g2699) & (g2081) & (!sk[35]) & (g2088) & (!g2705)) + ((g2699) & (g2081) & (!sk[35]) & (g2088) & (g2705)) + ((g2699) & (g2081) & (sk[35]) & (g2088) & (!g2705)) + ((g2699) & (g2081) & (sk[35]) & (g2088) & (g2705)));
	assign g3373 = (((!sk[36]) & (!g3374) & (g3375)) + ((!sk[36]) & (g3374) & (g3375)) + ((sk[36]) & (!g3374) & (!g3375)));
	assign g3374 = (((!g75) & (!sk[37]) & (g3376)) + ((!g75) & (sk[37]) & (g3376)) + ((g75) & (!sk[37]) & (g3376)));
	assign g3375 = (((!g75) & (!sk[38]) & (g3379)) + ((g75) & (!sk[38]) & (g3379)) + ((g75) & (sk[38]) & (g3379)));
	assign g3376 = (((!sk[39]) & (!g3377) & (g3378)) + ((!sk[39]) & (g3377) & (g3378)) + ((sk[39]) & (!g3377) & (!g3378)));
	assign g3377 = (((!g2280) & (!sk[40]) & (g2690)) + ((!g2280) & (sk[40]) & (g2690)) + ((g2280) & (!sk[40]) & (g2690)));
	assign g3378 = (((!g2096) & (!sk[41]) & (g2280)) + ((g2096) & (!sk[41]) & (g2280)) + ((g2096) & (sk[41]) & (g2280)));
	assign g3379 = (((!sk[42]) & (!g3380) & (g3381)) + ((!sk[42]) & (g3380) & (g3381)) + ((sk[42]) & (!g3380) & (!g3381)));
	assign g3380 = (((!g2280) & (!sk[43]) & (g3382)) + ((!g2280) & (sk[43]) & (g3382)) + ((g2280) & (!sk[43]) & (g3382)));
	assign g3381 = (((!g2280) & (!sk[44]) & (g3383)) + ((g2280) & (!sk[44]) & (g3383)) + ((g2280) & (sk[44]) & (g3383)));
	assign g3382 = (((!dmem_dat_ix23x) & (!g2127) & (sk[45]) & (g2550)) + ((!dmem_dat_ix23x) & (g2127) & (!sk[45]) & (!g2550)) + ((!dmem_dat_ix23x) & (g2127) & (!sk[45]) & (g2550)) + ((!dmem_dat_ix23x) & (g2127) & (sk[45]) & (g2550)) + ((dmem_dat_ix23x) & (!g2127) & (!sk[45]) & (!g2550)) + ((dmem_dat_ix23x) & (!g2127) & (!sk[45]) & (g2550)) + ((dmem_dat_ix23x) & (!g2127) & (sk[45]) & (g2550)) + ((dmem_dat_ix23x) & (g2127) & (!sk[45]) & (!g2550)) + ((dmem_dat_ix23x) & (g2127) & (!sk[45]) & (g2550)) + ((dmem_dat_ix23x) & (g2127) & (sk[45]) & (!g2550)) + ((dmem_dat_ix23x) & (g2127) & (sk[45]) & (g2550)));
	assign g3383 = (((!dmem_dat_ix23x) & (!g2127) & (sk[46]) & (g2550)) + ((!dmem_dat_ix23x) & (g2127) & (!sk[46]) & (!g2550)) + ((!dmem_dat_ix23x) & (g2127) & (!sk[46]) & (g2550)) + ((!dmem_dat_ix23x) & (g2127) & (sk[46]) & (g2550)) + ((dmem_dat_ix23x) & (!g2127) & (!sk[46]) & (!g2550)) + ((dmem_dat_ix23x) & (!g2127) & (!sk[46]) & (g2550)) + ((dmem_dat_ix23x) & (!g2127) & (sk[46]) & (g2550)) + ((dmem_dat_ix23x) & (g2127) & (!sk[46]) & (!g2550)) + ((dmem_dat_ix23x) & (g2127) & (!sk[46]) & (g2550)) + ((dmem_dat_ix23x) & (g2127) & (sk[46]) & (!g2550)) + ((dmem_dat_ix23x) & (g2127) & (sk[46]) & (g2550)));
	assign g3384 = (((!g3385) & (!sk[47]) & (g3386)) + ((!g3385) & (sk[47]) & (!g3386)) + ((g3385) & (!sk[47]) & (g3386)));
	assign g3385 = (((!sk[48]) & (!g2683) & (g3387)) + ((!sk[48]) & (g2683) & (g3387)) + ((sk[48]) & (!g2683) & (g3387)));
	assign g3386 = (((!g2683) & (!sk[49]) & (g3390)) + ((g2683) & (!sk[49]) & (g3390)) + ((g2683) & (sk[49]) & (g3390)));
	assign g3387 = (((!g3388) & (!sk[50]) & (g3389)) + ((!g3388) & (sk[50]) & (!g3389)) + ((g3388) & (!sk[50]) & (g3389)));
	assign g3388 = (((!g2125) & (!sk[51]) & (g3393)) + ((!g2125) & (sk[51]) & (g3393)) + ((g2125) & (!sk[51]) & (g3393)));
	assign g3389 = (((!sk[52]) & (!g2125) & (g3394)) + ((!sk[52]) & (g2125) & (g3394)) + ((sk[52]) & (g2125) & (g3394)));
	assign g3390 = (((!sk[53]) & (!g3391) & (g3392)) + ((!sk[53]) & (g3391) & (g3392)) + ((sk[53]) & (!g3391) & (!g3392)));
	assign g3391 = (((!sk[54]) & (!g2125) & (g3395)) + ((!sk[54]) & (g2125) & (g3395)) + ((sk[54]) & (!g2125) & (g3395)));
	assign g3392 = (((!sk[55]) & (!g2125) & (g3396)) + ((!sk[55]) & (g2125) & (g3396)) + ((sk[55]) & (g2125) & (g3396)));
	assign g3393 = (((!g2680) & (!g2096) & (!g2681) & (!sk[56]) & (g2081)) + ((!g2680) & (!g2096) & (g2681) & (!sk[56]) & (g2081)) + ((!g2680) & (!g2096) & (g2681) & (sk[56]) & (!g2081)) + ((!g2680) & (g2096) & (!g2681) & (!sk[56]) & (!g2081)) + ((!g2680) & (g2096) & (!g2681) & (!sk[56]) & (g2081)) + ((!g2680) & (g2096) & (!g2681) & (sk[56]) & (!g2081)) + ((!g2680) & (g2096) & (g2681) & (!sk[56]) & (!g2081)) + ((!g2680) & (g2096) & (g2681) & (!sk[56]) & (g2081)) + ((g2680) & (!g2096) & (!g2681) & (!sk[56]) & (!g2081)) + ((g2680) & (!g2096) & (!g2681) & (!sk[56]) & (g2081)) + ((g2680) & (!g2096) & (!g2681) & (sk[56]) & (!g2081)) + ((g2680) & (!g2096) & (g2681) & (!sk[56]) & (!g2081)) + ((g2680) & (!g2096) & (g2681) & (!sk[56]) & (g2081)) + ((g2680) & (g2096) & (!g2681) & (!sk[56]) & (!g2081)) + ((g2680) & (g2096) & (!g2681) & (!sk[56]) & (g2081)) + ((g2680) & (g2096) & (g2681) & (!sk[56]) & (!g2081)) + ((g2680) & (g2096) & (g2681) & (!sk[56]) & (g2081)) + ((g2680) & (g2096) & (g2681) & (sk[56]) & (!g2081)));
	assign g3394 = (((!g2680) & (!g2096) & (!sk[57]) & (!g2686) & (g2081)) + ((!g2680) & (!g2096) & (!sk[57]) & (g2686) & (g2081)) + ((!g2680) & (!g2096) & (sk[57]) & (g2686) & (!g2081)) + ((!g2680) & (g2096) & (!sk[57]) & (!g2686) & (!g2081)) + ((!g2680) & (g2096) & (!sk[57]) & (!g2686) & (g2081)) + ((!g2680) & (g2096) & (!sk[57]) & (g2686) & (!g2081)) + ((!g2680) & (g2096) & (!sk[57]) & (g2686) & (g2081)) + ((!g2680) & (g2096) & (sk[57]) & (g2686) & (!g2081)) + ((g2680) & (!g2096) & (!sk[57]) & (!g2686) & (!g2081)) + ((g2680) & (!g2096) & (!sk[57]) & (!g2686) & (g2081)) + ((g2680) & (!g2096) & (!sk[57]) & (g2686) & (!g2081)) + ((g2680) & (!g2096) & (!sk[57]) & (g2686) & (g2081)) + ((g2680) & (!g2096) & (sk[57]) & (g2686) & (!g2081)) + ((g2680) & (g2096) & (!sk[57]) & (!g2686) & (!g2081)) + ((g2680) & (g2096) & (!sk[57]) & (!g2686) & (g2081)) + ((g2680) & (g2096) & (!sk[57]) & (g2686) & (!g2081)) + ((g2680) & (g2096) & (!sk[57]) & (g2686) & (g2081)) + ((g2680) & (g2096) & (sk[57]) & (!g2686) & (g2081)) + ((g2680) & (g2096) & (sk[57]) & (g2686) & (!g2081)) + ((g2680) & (g2096) & (sk[57]) & (g2686) & (g2081)));
	assign g3395 = (((!g2680) & (!g2096) & (!sk[58]) & (!g2681) & (g2081)) + ((!g2680) & (!g2096) & (!sk[58]) & (g2681) & (g2081)) + ((!g2680) & (!g2096) & (sk[58]) & (!g2681) & (g2081)) + ((!g2680) & (!g2096) & (sk[58]) & (g2681) & (!g2081)) + ((!g2680) & (!g2096) & (sk[58]) & (g2681) & (g2081)) + ((!g2680) & (g2096) & (!sk[58]) & (!g2681) & (!g2081)) + ((!g2680) & (g2096) & (!sk[58]) & (!g2681) & (g2081)) + ((!g2680) & (g2096) & (!sk[58]) & (g2681) & (!g2081)) + ((!g2680) & (g2096) & (!sk[58]) & (g2681) & (g2081)) + ((!g2680) & (g2096) & (sk[58]) & (!g2681) & (!g2081)) + ((!g2680) & (g2096) & (sk[58]) & (!g2681) & (g2081)) + ((!g2680) & (g2096) & (sk[58]) & (g2681) & (g2081)) + ((g2680) & (!g2096) & (!sk[58]) & (!g2681) & (!g2081)) + ((g2680) & (!g2096) & (!sk[58]) & (!g2681) & (g2081)) + ((g2680) & (!g2096) & (!sk[58]) & (g2681) & (!g2081)) + ((g2680) & (!g2096) & (!sk[58]) & (g2681) & (g2081)) + ((g2680) & (!g2096) & (sk[58]) & (!g2681) & (!g2081)) + ((g2680) & (!g2096) & (sk[58]) & (!g2681) & (g2081)) + ((g2680) & (!g2096) & (sk[58]) & (g2681) & (g2081)) + ((g2680) & (g2096) & (!sk[58]) & (!g2681) & (!g2081)) + ((g2680) & (g2096) & (!sk[58]) & (!g2681) & (g2081)) + ((g2680) & (g2096) & (!sk[58]) & (g2681) & (!g2081)) + ((g2680) & (g2096) & (!sk[58]) & (g2681) & (g2081)) + ((g2680) & (g2096) & (sk[58]) & (!g2681) & (g2081)) + ((g2680) & (g2096) & (sk[58]) & (g2681) & (!g2081)) + ((g2680) & (g2096) & (sk[58]) & (g2681) & (g2081)));
	assign g3396 = (((!g2680) & (!sk[59]) & (!g2096) & (!g2686) & (g2081)) + ((!g2680) & (!sk[59]) & (!g2096) & (g2686) & (g2081)) + ((!g2680) & (!sk[59]) & (g2096) & (!g2686) & (!g2081)) + ((!g2680) & (!sk[59]) & (g2096) & (!g2686) & (g2081)) + ((!g2680) & (!sk[59]) & (g2096) & (g2686) & (!g2081)) + ((!g2680) & (!sk[59]) & (g2096) & (g2686) & (g2081)) + ((!g2680) & (sk[59]) & (!g2096) & (g2686) & (!g2081)) + ((!g2680) & (sk[59]) & (g2096) & (g2686) & (!g2081)) + ((g2680) & (!sk[59]) & (!g2096) & (!g2686) & (!g2081)) + ((g2680) & (!sk[59]) & (!g2096) & (!g2686) & (g2081)) + ((g2680) & (!sk[59]) & (!g2096) & (g2686) & (!g2081)) + ((g2680) & (!sk[59]) & (!g2096) & (g2686) & (g2081)) + ((g2680) & (!sk[59]) & (g2096) & (!g2686) & (!g2081)) + ((g2680) & (!sk[59]) & (g2096) & (!g2686) & (g2081)) + ((g2680) & (!sk[59]) & (g2096) & (g2686) & (!g2081)) + ((g2680) & (!sk[59]) & (g2096) & (g2686) & (g2081)) + ((g2680) & (sk[59]) & (!g2096) & (g2686) & (!g2081)) + ((g2680) & (sk[59]) & (g2096) & (!g2686) & (g2081)) + ((g2680) & (sk[59]) & (g2096) & (g2686) & (!g2081)) + ((g2680) & (sk[59]) & (g2096) & (g2686) & (g2081)));
	assign g3397 = (((!sk[60]) & (!g3398) & (g3399)) + ((!sk[60]) & (g3398) & (g3399)) + ((sk[60]) & (!g3398) & (!g3399)));
	assign g3398 = (((!sk[61]) & (!g75) & (g3400)) + ((!sk[61]) & (g75) & (g3400)) + ((sk[61]) & (!g75) & (g3400)));
	assign g3399 = (((!g75) & (!sk[62]) & (g3403)) + ((g75) & (!sk[62]) & (g3403)) + ((g75) & (sk[62]) & (g3403)));
	assign g3400 = (((!sk[63]) & (!g3401) & (g3402)) + ((!sk[63]) & (g3401) & (g3402)) + ((sk[63]) & (!g3401) & (!g3402)));
	assign g3401 = (((!g2280) & (!sk[64]) & (g2672)) + ((!g2280) & (sk[64]) & (g2672)) + ((g2280) & (!sk[64]) & (g2672)));
	assign g3402 = (((!g2095) & (!sk[65]) & (g2280)) + ((g2095) & (!sk[65]) & (g2280)) + ((g2095) & (sk[65]) & (g2280)));
	assign g3403 = (((!sk[66]) & (!g3404) & (g3405)) + ((!sk[66]) & (g3404) & (g3405)) + ((sk[66]) & (!g3404) & (!g3405)));
	assign g3404 = (((!sk[67]) & (!g2280) & (g3406)) + ((!sk[67]) & (g2280) & (g3406)) + ((sk[67]) & (!g2280) & (g3406)));
	assign g3405 = (((!g2280) & (!sk[68]) & (g3407)) + ((g2280) & (!sk[68]) & (g3407)) + ((g2280) & (sk[68]) & (g3407)));
	assign g3406 = (((!dmem_dat_ix22x) & (!g2127) & (sk[69]) & (g2550)) + ((!dmem_dat_ix22x) & (g2127) & (!sk[69]) & (!g2550)) + ((!dmem_dat_ix22x) & (g2127) & (!sk[69]) & (g2550)) + ((!dmem_dat_ix22x) & (g2127) & (sk[69]) & (g2550)) + ((dmem_dat_ix22x) & (!g2127) & (!sk[69]) & (!g2550)) + ((dmem_dat_ix22x) & (!g2127) & (!sk[69]) & (g2550)) + ((dmem_dat_ix22x) & (!g2127) & (sk[69]) & (g2550)) + ((dmem_dat_ix22x) & (g2127) & (!sk[69]) & (!g2550)) + ((dmem_dat_ix22x) & (g2127) & (!sk[69]) & (g2550)) + ((dmem_dat_ix22x) & (g2127) & (sk[69]) & (!g2550)) + ((dmem_dat_ix22x) & (g2127) & (sk[69]) & (g2550)));
	assign g3407 = (((!dmem_dat_ix22x) & (!sk[70]) & (g2127) & (!g2550)) + ((!dmem_dat_ix22x) & (!sk[70]) & (g2127) & (g2550)) + ((!dmem_dat_ix22x) & (sk[70]) & (!g2127) & (g2550)) + ((!dmem_dat_ix22x) & (sk[70]) & (g2127) & (g2550)) + ((dmem_dat_ix22x) & (!sk[70]) & (!g2127) & (!g2550)) + ((dmem_dat_ix22x) & (!sk[70]) & (!g2127) & (g2550)) + ((dmem_dat_ix22x) & (!sk[70]) & (g2127) & (!g2550)) + ((dmem_dat_ix22x) & (!sk[70]) & (g2127) & (g2550)) + ((dmem_dat_ix22x) & (sk[70]) & (!g2127) & (g2550)) + ((dmem_dat_ix22x) & (sk[70]) & (g2127) & (!g2550)) + ((dmem_dat_ix22x) & (sk[70]) & (g2127) & (g2550)));
	assign g3408 = (((!g3409) & (!sk[71]) & (g3410)) + ((!g3409) & (sk[71]) & (!g3410)) + ((g3409) & (!sk[71]) & (g3410)));
	assign g3409 = (((!sk[72]) & (!g2662) & (g3411)) + ((!sk[72]) & (g2662) & (g3411)) + ((sk[72]) & (!g2662) & (g3411)));
	assign g3410 = (((!g2662) & (!sk[73]) & (g3414)) + ((g2662) & (!sk[73]) & (g3414)) + ((g2662) & (sk[73]) & (g3414)));
	assign g3411 = (((!sk[74]) & (!g3412) & (g3413)) + ((!sk[74]) & (g3412) & (g3413)) + ((sk[74]) & (!g3412) & (!g3413)));
	assign g3412 = (((!g2125) & (!sk[75]) & (g2661)) + ((!g2125) & (sk[75]) & (g2661)) + ((g2125) & (!sk[75]) & (g2661)));
	assign g3413 = (((!g2125) & (!sk[76]) & (g3417)) + ((g2125) & (!sk[76]) & (g3417)) + ((g2125) & (sk[76]) & (g3417)));
	assign g3414 = (((!sk[77]) & (!g3415) & (g3416)) + ((!sk[77]) & (g3415) & (g3416)) + ((sk[77]) & (!g3415) & (!g3416)));
	assign g3415 = (((!sk[78]) & (!g2125) & (g3418)) + ((!sk[78]) & (g2125) & (g3418)) + ((sk[78]) & (!g2125) & (g3418)));
	assign g3416 = (((!sk[79]) & (!g2125) & (g3419)) + ((!sk[79]) & (g2125) & (g3419)) + ((sk[79]) & (g2125) & (g3419)));
	assign g3417 = (((!g2660) & (!sk[80]) & (!g2081) & (!g2095) & (g2668)) + ((!g2660) & (!sk[80]) & (!g2081) & (g2095) & (g2668)) + ((!g2660) & (!sk[80]) & (g2081) & (!g2095) & (!g2668)) + ((!g2660) & (!sk[80]) & (g2081) & (!g2095) & (g2668)) + ((!g2660) & (!sk[80]) & (g2081) & (g2095) & (!g2668)) + ((!g2660) & (!sk[80]) & (g2081) & (g2095) & (g2668)) + ((!g2660) & (sk[80]) & (!g2081) & (!g2095) & (g2668)) + ((!g2660) & (sk[80]) & (!g2081) & (g2095) & (g2668)) + ((g2660) & (!sk[80]) & (!g2081) & (!g2095) & (!g2668)) + ((g2660) & (!sk[80]) & (!g2081) & (!g2095) & (g2668)) + ((g2660) & (!sk[80]) & (!g2081) & (g2095) & (!g2668)) + ((g2660) & (!sk[80]) & (!g2081) & (g2095) & (g2668)) + ((g2660) & (!sk[80]) & (g2081) & (!g2095) & (!g2668)) + ((g2660) & (!sk[80]) & (g2081) & (!g2095) & (g2668)) + ((g2660) & (!sk[80]) & (g2081) & (g2095) & (!g2668)) + ((g2660) & (!sk[80]) & (g2081) & (g2095) & (g2668)) + ((g2660) & (sk[80]) & (!g2081) & (!g2095) & (g2668)) + ((g2660) & (sk[80]) & (!g2081) & (g2095) & (g2668)) + ((g2660) & (sk[80]) & (g2081) & (g2095) & (!g2668)) + ((g2660) & (sk[80]) & (g2081) & (g2095) & (g2668)));
	assign g3418 = (((!g2081) & (!sk[81]) & (g2661)) + ((!g2081) & (sk[81]) & (g2661)) + ((g2081) & (!sk[81]) & (g2661)) + ((g2081) & (sk[81]) & (!g2661)));
	assign g3419 = (((!sk[82]) & (!g2660) & (!g2081) & (!g2095) & (g2668)) + ((!sk[82]) & (!g2660) & (!g2081) & (g2095) & (g2668)) + ((!sk[82]) & (!g2660) & (g2081) & (!g2095) & (!g2668)) + ((!sk[82]) & (!g2660) & (g2081) & (!g2095) & (g2668)) + ((!sk[82]) & (!g2660) & (g2081) & (g2095) & (!g2668)) + ((!sk[82]) & (!g2660) & (g2081) & (g2095) & (g2668)) + ((!sk[82]) & (g2660) & (!g2081) & (!g2095) & (!g2668)) + ((!sk[82]) & (g2660) & (!g2081) & (!g2095) & (g2668)) + ((!sk[82]) & (g2660) & (!g2081) & (g2095) & (!g2668)) + ((!sk[82]) & (g2660) & (!g2081) & (g2095) & (g2668)) + ((!sk[82]) & (g2660) & (g2081) & (!g2095) & (!g2668)) + ((!sk[82]) & (g2660) & (g2081) & (!g2095) & (g2668)) + ((!sk[82]) & (g2660) & (g2081) & (g2095) & (!g2668)) + ((!sk[82]) & (g2660) & (g2081) & (g2095) & (g2668)) + ((sk[82]) & (!g2660) & (!g2081) & (!g2095) & (g2668)) + ((sk[82]) & (!g2660) & (!g2081) & (g2095) & (g2668)) + ((sk[82]) & (g2660) & (!g2081) & (!g2095) & (g2668)) + ((sk[82]) & (g2660) & (!g2081) & (g2095) & (g2668)) + ((sk[82]) & (g2660) & (g2081) & (g2095) & (!g2668)) + ((sk[82]) & (g2660) & (g2081) & (g2095) & (g2668)));
	assign g3420 = (((!g3421) & (!sk[83]) & (g3422)) + ((!g3421) & (sk[83]) & (!g3422)) + ((g3421) & (!sk[83]) & (g3422)));
	assign g3421 = (((!g75) & (!sk[84]) & (g3423)) + ((!g75) & (sk[84]) & (g3423)) + ((g75) & (!sk[84]) & (g3423)));
	assign g3422 = (((!sk[85]) & (!g75) & (g3426)) + ((!sk[85]) & (g75) & (g3426)) + ((sk[85]) & (g75) & (g3426)));
	assign g3423 = (((!g3424) & (!sk[86]) & (g3425)) + ((!g3424) & (sk[86]) & (!g3425)) + ((g3424) & (!sk[86]) & (g3425)));
	assign g3424 = (((!g2280) & (!sk[87]) & (g2653)) + ((!g2280) & (sk[87]) & (g2653)) + ((g2280) & (!sk[87]) & (g2653)));
	assign g3425 = (((!sk[88]) & (!g2094) & (g2280)) + ((!sk[88]) & (g2094) & (g2280)) + ((sk[88]) & (g2094) & (g2280)));
	assign g3426 = (((!g3427) & (!sk[89]) & (g3428)) + ((!g3427) & (sk[89]) & (!g3428)) + ((g3427) & (!sk[89]) & (g3428)));
	assign g3427 = (((!g2280) & (!sk[90]) & (g3429)) + ((!g2280) & (sk[90]) & (g3429)) + ((g2280) & (!sk[90]) & (g3429)));
	assign g3428 = (((!sk[91]) & (!g2280) & (g3430)) + ((!sk[91]) & (g2280) & (g3430)) + ((sk[91]) & (g2280) & (g3430)));
	assign g3429 = (((!dmem_dat_ix21x) & (!sk[92]) & (g2127) & (!g2550)) + ((!dmem_dat_ix21x) & (!sk[92]) & (g2127) & (g2550)) + ((!dmem_dat_ix21x) & (sk[92]) & (!g2127) & (g2550)) + ((!dmem_dat_ix21x) & (sk[92]) & (g2127) & (g2550)) + ((dmem_dat_ix21x) & (!sk[92]) & (!g2127) & (!g2550)) + ((dmem_dat_ix21x) & (!sk[92]) & (!g2127) & (g2550)) + ((dmem_dat_ix21x) & (!sk[92]) & (g2127) & (!g2550)) + ((dmem_dat_ix21x) & (!sk[92]) & (g2127) & (g2550)) + ((dmem_dat_ix21x) & (sk[92]) & (!g2127) & (g2550)) + ((dmem_dat_ix21x) & (sk[92]) & (g2127) & (!g2550)) + ((dmem_dat_ix21x) & (sk[92]) & (g2127) & (g2550)));
	assign g3430 = (((!dmem_dat_ix21x) & (!sk[93]) & (g2127) & (!g2550)) + ((!dmem_dat_ix21x) & (!sk[93]) & (g2127) & (g2550)) + ((!dmem_dat_ix21x) & (sk[93]) & (!g2127) & (g2550)) + ((!dmem_dat_ix21x) & (sk[93]) & (g2127) & (g2550)) + ((dmem_dat_ix21x) & (!sk[93]) & (!g2127) & (!g2550)) + ((dmem_dat_ix21x) & (!sk[93]) & (!g2127) & (g2550)) + ((dmem_dat_ix21x) & (!sk[93]) & (g2127) & (!g2550)) + ((dmem_dat_ix21x) & (!sk[93]) & (g2127) & (g2550)) + ((dmem_dat_ix21x) & (sk[93]) & (!g2127) & (g2550)) + ((dmem_dat_ix21x) & (sk[93]) & (g2127) & (!g2550)) + ((dmem_dat_ix21x) & (sk[93]) & (g2127) & (g2550)));
	assign g3431 = (((!g3432) & (!sk[94]) & (g3433)) + ((!g3432) & (sk[94]) & (!g3433)) + ((g3432) & (!sk[94]) & (g3433)));
	assign g3432 = (((!g2646) & (!sk[95]) & (g3434)) + ((!g2646) & (sk[95]) & (g3434)) + ((g2646) & (!sk[95]) & (g3434)));
	assign g3433 = (((!sk[96]) & (!g2646) & (g3437)) + ((!sk[96]) & (g2646) & (g3437)) + ((sk[96]) & (g2646) & (g3437)));
	assign g3434 = (((!sk[97]) & (!g3435) & (g3436)) + ((!sk[97]) & (g3435) & (g3436)) + ((sk[97]) & (!g3435) & (!g3436)));
	assign g3435 = (((!sk[98]) & (!g2125) & (g3440)) + ((!sk[98]) & (g2125) & (g3440)) + ((sk[98]) & (!g2125) & (g3440)));
	assign g3436 = (((!sk[99]) & (!g2125) & (g3441)) + ((!sk[99]) & (g2125) & (g3441)) + ((sk[99]) & (g2125) & (g3441)));
	assign g3437 = (((!g3438) & (!sk[100]) & (g3439)) + ((!g3438) & (sk[100]) & (!g3439)) + ((g3438) & (!sk[100]) & (g3439)));
	assign g3438 = (((!sk[101]) & (!g2125) & (g3442)) + ((!sk[101]) & (g2125) & (g3442)) + ((sk[101]) & (!g2125) & (g3442)));
	assign g3439 = (((!sk[102]) & (!g2125) & (g3443)) + ((!sk[102]) & (g2125) & (g3443)) + ((sk[102]) & (g2125) & (g3443)));
	assign g3440 = (((!sk[103]) & (!g2081) & (g2645)) + ((!sk[103]) & (g2081) & (g2645)) + ((sk[103]) & (!g2081) & (g2645)));
	assign g3441 = (((!g2642) & (!sk[104]) & (!g2081) & (!g2094) & (g2649)) + ((!g2642) & (!sk[104]) & (!g2081) & (g2094) & (g2649)) + ((!g2642) & (!sk[104]) & (g2081) & (!g2094) & (!g2649)) + ((!g2642) & (!sk[104]) & (g2081) & (!g2094) & (g2649)) + ((!g2642) & (!sk[104]) & (g2081) & (g2094) & (!g2649)) + ((!g2642) & (!sk[104]) & (g2081) & (g2094) & (g2649)) + ((!g2642) & (sk[104]) & (!g2081) & (!g2094) & (g2649)) + ((!g2642) & (sk[104]) & (!g2081) & (g2094) & (g2649)) + ((g2642) & (!sk[104]) & (!g2081) & (!g2094) & (!g2649)) + ((g2642) & (!sk[104]) & (!g2081) & (!g2094) & (g2649)) + ((g2642) & (!sk[104]) & (!g2081) & (g2094) & (!g2649)) + ((g2642) & (!sk[104]) & (!g2081) & (g2094) & (g2649)) + ((g2642) & (!sk[104]) & (g2081) & (!g2094) & (!g2649)) + ((g2642) & (!sk[104]) & (g2081) & (!g2094) & (g2649)) + ((g2642) & (!sk[104]) & (g2081) & (g2094) & (!g2649)) + ((g2642) & (!sk[104]) & (g2081) & (g2094) & (g2649)) + ((g2642) & (sk[104]) & (!g2081) & (!g2094) & (g2649)) + ((g2642) & (sk[104]) & (!g2081) & (g2094) & (g2649)) + ((g2642) & (sk[104]) & (g2081) & (g2094) & (!g2649)) + ((g2642) & (sk[104]) & (g2081) & (g2094) & (g2649)));
	assign g3442 = (((!g2081) & (!sk[105]) & (g2645)) + ((!g2081) & (sk[105]) & (g2645)) + ((g2081) & (!sk[105]) & (g2645)) + ((g2081) & (sk[105]) & (!g2645)) + ((g2081) & (sk[105]) & (g2645)));
	assign g3443 = (((!sk[106]) & (!g2642) & (!g2081) & (!g2094) & (g2649)) + ((!sk[106]) & (!g2642) & (!g2081) & (g2094) & (g2649)) + ((!sk[106]) & (!g2642) & (g2081) & (!g2094) & (!g2649)) + ((!sk[106]) & (!g2642) & (g2081) & (!g2094) & (g2649)) + ((!sk[106]) & (!g2642) & (g2081) & (g2094) & (!g2649)) + ((!sk[106]) & (!g2642) & (g2081) & (g2094) & (g2649)) + ((!sk[106]) & (g2642) & (!g2081) & (!g2094) & (!g2649)) + ((!sk[106]) & (g2642) & (!g2081) & (!g2094) & (g2649)) + ((!sk[106]) & (g2642) & (!g2081) & (g2094) & (!g2649)) + ((!sk[106]) & (g2642) & (!g2081) & (g2094) & (g2649)) + ((!sk[106]) & (g2642) & (g2081) & (!g2094) & (!g2649)) + ((!sk[106]) & (g2642) & (g2081) & (!g2094) & (g2649)) + ((!sk[106]) & (g2642) & (g2081) & (g2094) & (!g2649)) + ((!sk[106]) & (g2642) & (g2081) & (g2094) & (g2649)) + ((sk[106]) & (!g2642) & (!g2081) & (!g2094) & (g2649)) + ((sk[106]) & (!g2642) & (!g2081) & (g2094) & (g2649)) + ((sk[106]) & (g2642) & (!g2081) & (!g2094) & (g2649)) + ((sk[106]) & (g2642) & (!g2081) & (g2094) & (g2649)) + ((sk[106]) & (g2642) & (g2081) & (g2094) & (!g2649)) + ((sk[106]) & (g2642) & (g2081) & (g2094) & (g2649)));
	assign g3444 = (((!g3445) & (!sk[107]) & (g3446)) + ((!g3445) & (sk[107]) & (!g3446)) + ((g3445) & (!sk[107]) & (g3446)));
	assign g3445 = (((!sk[108]) & (!g75) & (g3447)) + ((!sk[108]) & (g75) & (g3447)) + ((sk[108]) & (!g75) & (g3447)));
	assign g3446 = (((!sk[109]) & (!g75) & (g3450)) + ((!sk[109]) & (g75) & (g3450)) + ((sk[109]) & (g75) & (g3450)));
	assign g3447 = (((!g3448) & (!sk[110]) & (g3449)) + ((!g3448) & (sk[110]) & (!g3449)) + ((g3448) & (!sk[110]) & (g3449)));
	assign g3448 = (((!g2280) & (!sk[111]) & (g2635)) + ((!g2280) & (sk[111]) & (g2635)) + ((g2280) & (!sk[111]) & (g2635)));
	assign g3449 = (((!sk[112]) & (!g2093) & (g2280)) + ((!sk[112]) & (g2093) & (g2280)) + ((sk[112]) & (g2093) & (g2280)));
	assign g3450 = (((!g3451) & (!sk[113]) & (g3452)) + ((!g3451) & (sk[113]) & (!g3452)) + ((g3451) & (!sk[113]) & (g3452)));
	assign g3451 = (((!sk[114]) & (!g2280) & (g3453)) + ((!sk[114]) & (g2280) & (g3453)) + ((sk[114]) & (!g2280) & (g3453)));
	assign g3452 = (((!g2280) & (!sk[115]) & (g3454)) + ((g2280) & (!sk[115]) & (g3454)) + ((g2280) & (sk[115]) & (g3454)));
	assign g3453 = (((!sk[116]) & (!dmem_dat_ix20x) & (g2127) & (!g2550)) + ((!sk[116]) & (!dmem_dat_ix20x) & (g2127) & (g2550)) + ((!sk[116]) & (dmem_dat_ix20x) & (!g2127) & (!g2550)) + ((!sk[116]) & (dmem_dat_ix20x) & (!g2127) & (g2550)) + ((!sk[116]) & (dmem_dat_ix20x) & (g2127) & (!g2550)) + ((!sk[116]) & (dmem_dat_ix20x) & (g2127) & (g2550)) + ((sk[116]) & (!dmem_dat_ix20x) & (!g2127) & (g2550)) + ((sk[116]) & (!dmem_dat_ix20x) & (g2127) & (g2550)) + ((sk[116]) & (dmem_dat_ix20x) & (!g2127) & (g2550)) + ((sk[116]) & (dmem_dat_ix20x) & (g2127) & (!g2550)) + ((sk[116]) & (dmem_dat_ix20x) & (g2127) & (g2550)));
	assign g3454 = (((!dmem_dat_ix20x) & (!g2127) & (sk[117]) & (g2550)) + ((!dmem_dat_ix20x) & (g2127) & (!sk[117]) & (!g2550)) + ((!dmem_dat_ix20x) & (g2127) & (!sk[117]) & (g2550)) + ((!dmem_dat_ix20x) & (g2127) & (sk[117]) & (g2550)) + ((dmem_dat_ix20x) & (!g2127) & (!sk[117]) & (!g2550)) + ((dmem_dat_ix20x) & (!g2127) & (!sk[117]) & (g2550)) + ((dmem_dat_ix20x) & (!g2127) & (sk[117]) & (g2550)) + ((dmem_dat_ix20x) & (g2127) & (!sk[117]) & (!g2550)) + ((dmem_dat_ix20x) & (g2127) & (!sk[117]) & (g2550)) + ((dmem_dat_ix20x) & (g2127) & (sk[117]) & (!g2550)) + ((dmem_dat_ix20x) & (g2127) & (sk[117]) & (g2550)));
	assign g3455 = (((!sk[118]) & (!g3456) & (g3457)) + ((!sk[118]) & (g3456) & (g3457)) + ((sk[118]) & (!g3456) & (!g3457)));
	assign g3456 = (((!sk[119]) & (!g2626) & (g3458)) + ((!sk[119]) & (g2626) & (g3458)) + ((sk[119]) & (!g2626) & (g3458)));
	assign g3457 = (((!g2626) & (!sk[120]) & (g3461)) + ((g2626) & (!sk[120]) & (g3461)) + ((g2626) & (sk[120]) & (g3461)));
	assign g3458 = (((!sk[121]) & (!g3459) & (g3460)) + ((!sk[121]) & (g3459) & (g3460)) + ((sk[121]) & (!g3459) & (!g3460)));
	assign g3459 = (((!sk[122]) & (!g2125) & (g3464)) + ((!sk[122]) & (g2125) & (g3464)) + ((sk[122]) & (!g2125) & (g3464)));
	assign g3460 = (((!g2125) & (!sk[123]) & (g3465)) + ((g2125) & (!sk[123]) & (g3465)) + ((g2125) & (sk[123]) & (g3465)));
	assign g3461 = (((!sk[124]) & (!g3462) & (g3463)) + ((!sk[124]) & (g3462) & (g3463)) + ((sk[124]) & (!g3462) & (!g3463)));
	assign g3462 = (((!sk[125]) & (!g2125) & (g3466)) + ((!sk[125]) & (g2125) & (g3466)) + ((sk[125]) & (!g2125) & (g3466)));
	assign g3463 = (((!g2125) & (!sk[126]) & (g3467)) + ((g2125) & (!sk[126]) & (g3467)) + ((g2125) & (sk[126]) & (g3467)));
	assign g3464 = (((!g2610) & (g2081) & (!sk[127]) & (!g2609)) + ((!g2610) & (g2081) & (!sk[127]) & (g2609)) + ((g2610) & (!g2081) & (!sk[127]) & (!g2609)) + ((g2610) & (!g2081) & (!sk[127]) & (g2609)) + ((g2610) & (g2081) & (!sk[127]) & (!g2609)) + ((g2610) & (g2081) & (!sk[127]) & (g2609)) + ((g2610) & (g2081) & (sk[127]) & (g2609)));
	assign g3465 = (((!g2081) & (g2630) & (!sk[0]) & (!g2631)) + ((!g2081) & (g2630) & (!sk[0]) & (g2631)) + ((!g2081) & (g2630) & (sk[0]) & (!g2631)) + ((!g2081) & (g2630) & (sk[0]) & (g2631)) + ((g2081) & (!g2630) & (!sk[0]) & (!g2631)) + ((g2081) & (!g2630) & (!sk[0]) & (g2631)) + ((g2081) & (!g2630) & (sk[0]) & (g2631)) + ((g2081) & (g2630) & (!sk[0]) & (!g2631)) + ((g2081) & (g2630) & (!sk[0]) & (g2631)) + ((g2081) & (g2630) & (sk[0]) & (g2631)));
	assign g3466 = (((!g2610) & (!sk[1]) & (g2081) & (!g2609)) + ((!g2610) & (!sk[1]) & (g2081) & (g2609)) + ((!g2610) & (sk[1]) & (!g2081) & (!g2609)) + ((!g2610) & (sk[1]) & (!g2081) & (g2609)) + ((!g2610) & (sk[1]) & (g2081) & (!g2609)) + ((!g2610) & (sk[1]) & (g2081) & (g2609)) + ((g2610) & (!sk[1]) & (!g2081) & (!g2609)) + ((g2610) & (!sk[1]) & (!g2081) & (g2609)) + ((g2610) & (!sk[1]) & (g2081) & (!g2609)) + ((g2610) & (!sk[1]) & (g2081) & (g2609)) + ((g2610) & (sk[1]) & (!g2081) & (!g2609)) + ((g2610) & (sk[1]) & (!g2081) & (g2609)) + ((g2610) & (sk[1]) & (g2081) & (!g2609)));
	assign g3467 = (((!g2081) & (g2630) & (!sk[2]) & (!g2631)) + ((!g2081) & (g2630) & (!sk[2]) & (g2631)) + ((!g2081) & (g2630) & (sk[2]) & (!g2631)) + ((!g2081) & (g2630) & (sk[2]) & (g2631)) + ((g2081) & (!g2630) & (!sk[2]) & (!g2631)) + ((g2081) & (!g2630) & (!sk[2]) & (g2631)) + ((g2081) & (!g2630) & (sk[2]) & (g2631)) + ((g2081) & (g2630) & (!sk[2]) & (!g2631)) + ((g2081) & (g2630) & (!sk[2]) & (g2631)) + ((g2081) & (g2630) & (sk[2]) & (g2631)));
	assign g3468 = (((!g3469) & (!sk[3]) & (g3470)) + ((!g3469) & (sk[3]) & (!g3470)) + ((g3469) & (!sk[3]) & (g3470)));
	assign g3469 = (((!sk[4]) & (!g75) & (g3471)) + ((!sk[4]) & (g75) & (g3471)) + ((sk[4]) & (!g75) & (g3471)));
	assign g3470 = (((!g75) & (!sk[5]) & (g3474)) + ((g75) & (!sk[5]) & (g3474)) + ((g75) & (sk[5]) & (g3474)));
	assign g3471 = (((!g3472) & (!sk[6]) & (g3473)) + ((!g3472) & (sk[6]) & (!g3473)) + ((g3472) & (!sk[6]) & (g3473)));
	assign g3472 = (((!g2280) & (!sk[7]) & (g2618)) + ((!g2280) & (sk[7]) & (g2618)) + ((g2280) & (!sk[7]) & (g2618)));
	assign g3473 = (((!sk[8]) & (!g2086) & (g2280)) + ((!sk[8]) & (g2086) & (g2280)) + ((sk[8]) & (g2086) & (g2280)));
	assign g3474 = (((!g3475) & (!sk[9]) & (g3476)) + ((!g3475) & (sk[9]) & (!g3476)) + ((g3475) & (!sk[9]) & (g3476)));
	assign g3475 = (((!sk[10]) & (!g2280) & (g3477)) + ((!sk[10]) & (g2280) & (g3477)) + ((sk[10]) & (!g2280) & (g3477)));
	assign g3476 = (((!g2280) & (!sk[11]) & (g3478)) + ((g2280) & (!sk[11]) & (g3478)) + ((g2280) & (sk[11]) & (g3478)));
	assign g3477 = (((!sk[12]) & (!dmem_dat_ix19x) & (g2127) & (!g2550)) + ((!sk[12]) & (!dmem_dat_ix19x) & (g2127) & (g2550)) + ((!sk[12]) & (dmem_dat_ix19x) & (!g2127) & (!g2550)) + ((!sk[12]) & (dmem_dat_ix19x) & (!g2127) & (g2550)) + ((!sk[12]) & (dmem_dat_ix19x) & (g2127) & (!g2550)) + ((!sk[12]) & (dmem_dat_ix19x) & (g2127) & (g2550)) + ((sk[12]) & (!dmem_dat_ix19x) & (!g2127) & (g2550)) + ((sk[12]) & (!dmem_dat_ix19x) & (g2127) & (g2550)) + ((sk[12]) & (dmem_dat_ix19x) & (!g2127) & (g2550)) + ((sk[12]) & (dmem_dat_ix19x) & (g2127) & (!g2550)) + ((sk[12]) & (dmem_dat_ix19x) & (g2127) & (g2550)));
	assign g3478 = (((!sk[13]) & (!dmem_dat_ix19x) & (g2127) & (!g2550)) + ((!sk[13]) & (!dmem_dat_ix19x) & (g2127) & (g2550)) + ((!sk[13]) & (dmem_dat_ix19x) & (!g2127) & (!g2550)) + ((!sk[13]) & (dmem_dat_ix19x) & (!g2127) & (g2550)) + ((!sk[13]) & (dmem_dat_ix19x) & (g2127) & (!g2550)) + ((!sk[13]) & (dmem_dat_ix19x) & (g2127) & (g2550)) + ((sk[13]) & (!dmem_dat_ix19x) & (!g2127) & (g2550)) + ((sk[13]) & (!dmem_dat_ix19x) & (g2127) & (g2550)) + ((sk[13]) & (dmem_dat_ix19x) & (!g2127) & (g2550)) + ((sk[13]) & (dmem_dat_ix19x) & (g2127) & (!g2550)) + ((sk[13]) & (dmem_dat_ix19x) & (g2127) & (g2550)));
	assign g3479 = (((!g3480) & (!sk[14]) & (g3481)) + ((!g3480) & (sk[14]) & (!g3481)) + ((g3480) & (!sk[14]) & (g3481)));
	assign g3480 = (((!g2610) & (!sk[15]) & (g3482)) + ((!g2610) & (sk[15]) & (g3482)) + ((g2610) & (!sk[15]) & (g3482)));
	assign g3481 = (((!sk[16]) & (!g2610) & (g3485)) + ((!sk[16]) & (g2610) & (g3485)) + ((sk[16]) & (g2610) & (g3485)));
	assign g3482 = (((!g3483) & (!sk[17]) & (g3484)) + ((!g3483) & (sk[17]) & (!g3484)) + ((g3483) & (!sk[17]) & (g3484)));
	assign g3483 = (((!g2125) & (!sk[18]) & (g2609)) + ((!g2125) & (sk[18]) & (g2609)) + ((g2125) & (!sk[18]) & (g2609)));
	assign g3484 = (((!g2125) & (!sk[19]) & (g3488)) + ((g2125) & (!sk[19]) & (g3488)) + ((g2125) & (sk[19]) & (g3488)));
	assign g3485 = (((!sk[20]) & (!g3486) & (g3487)) + ((!sk[20]) & (g3486) & (g3487)) + ((sk[20]) & (!g3486) & (!g3487)));
	assign g3486 = (((!g2125) & (!sk[21]) & (g3489)) + ((!g2125) & (sk[21]) & (g3489)) + ((g2125) & (!sk[21]) & (g3489)));
	assign g3487 = (((!g2125) & (!sk[22]) & (g3490)) + ((g2125) & (!sk[22]) & (g3490)) + ((g2125) & (sk[22]) & (g3490)));
	assign g3488 = (((!sk[23]) & (!g2608) & (!g2081) & (!g2086) & (g2614)) + ((!sk[23]) & (!g2608) & (!g2081) & (g2086) & (g2614)) + ((!sk[23]) & (!g2608) & (g2081) & (!g2086) & (!g2614)) + ((!sk[23]) & (!g2608) & (g2081) & (!g2086) & (g2614)) + ((!sk[23]) & (!g2608) & (g2081) & (g2086) & (!g2614)) + ((!sk[23]) & (!g2608) & (g2081) & (g2086) & (g2614)) + ((!sk[23]) & (g2608) & (!g2081) & (!g2086) & (!g2614)) + ((!sk[23]) & (g2608) & (!g2081) & (!g2086) & (g2614)) + ((!sk[23]) & (g2608) & (!g2081) & (g2086) & (!g2614)) + ((!sk[23]) & (g2608) & (!g2081) & (g2086) & (g2614)) + ((!sk[23]) & (g2608) & (g2081) & (!g2086) & (!g2614)) + ((!sk[23]) & (g2608) & (g2081) & (!g2086) & (g2614)) + ((!sk[23]) & (g2608) & (g2081) & (g2086) & (!g2614)) + ((!sk[23]) & (g2608) & (g2081) & (g2086) & (g2614)) + ((sk[23]) & (!g2608) & (!g2081) & (!g2086) & (g2614)) + ((sk[23]) & (!g2608) & (!g2081) & (g2086) & (g2614)) + ((sk[23]) & (g2608) & (!g2081) & (!g2086) & (g2614)) + ((sk[23]) & (g2608) & (!g2081) & (g2086) & (g2614)) + ((sk[23]) & (g2608) & (g2081) & (g2086) & (!g2614)) + ((sk[23]) & (g2608) & (g2081) & (g2086) & (g2614)));
	assign g3489 = (((!g2081) & (!sk[24]) & (g2609)) + ((!g2081) & (sk[24]) & (g2609)) + ((g2081) & (!sk[24]) & (g2609)) + ((g2081) & (sk[24]) & (!g2609)));
	assign g3490 = (((!g2608) & (!g2081) & (!g2086) & (!sk[25]) & (g2614)) + ((!g2608) & (!g2081) & (!g2086) & (sk[25]) & (g2614)) + ((!g2608) & (!g2081) & (g2086) & (!sk[25]) & (g2614)) + ((!g2608) & (!g2081) & (g2086) & (sk[25]) & (g2614)) + ((!g2608) & (g2081) & (!g2086) & (!sk[25]) & (!g2614)) + ((!g2608) & (g2081) & (!g2086) & (!sk[25]) & (g2614)) + ((!g2608) & (g2081) & (g2086) & (!sk[25]) & (!g2614)) + ((!g2608) & (g2081) & (g2086) & (!sk[25]) & (g2614)) + ((g2608) & (!g2081) & (!g2086) & (!sk[25]) & (!g2614)) + ((g2608) & (!g2081) & (!g2086) & (!sk[25]) & (g2614)) + ((g2608) & (!g2081) & (!g2086) & (sk[25]) & (g2614)) + ((g2608) & (!g2081) & (g2086) & (!sk[25]) & (!g2614)) + ((g2608) & (!g2081) & (g2086) & (!sk[25]) & (g2614)) + ((g2608) & (!g2081) & (g2086) & (sk[25]) & (g2614)) + ((g2608) & (g2081) & (!g2086) & (!sk[25]) & (!g2614)) + ((g2608) & (g2081) & (!g2086) & (!sk[25]) & (g2614)) + ((g2608) & (g2081) & (g2086) & (!sk[25]) & (!g2614)) + ((g2608) & (g2081) & (g2086) & (!sk[25]) & (g2614)) + ((g2608) & (g2081) & (g2086) & (sk[25]) & (!g2614)) + ((g2608) & (g2081) & (g2086) & (sk[25]) & (g2614)));
	assign g3491 = (((!g3492) & (!sk[26]) & (g3493)) + ((!g3492) & (sk[26]) & (!g3493)) + ((g3492) & (!sk[26]) & (g3493)));
	assign g3492 = (((!sk[27]) & (!g75) & (g3494)) + ((!sk[27]) & (g75) & (g3494)) + ((sk[27]) & (!g75) & (g3494)));
	assign g3493 = (((!sk[28]) & (!g75) & (g3497)) + ((!sk[28]) & (g75) & (g3497)) + ((sk[28]) & (g75) & (g3497)));
	assign g3494 = (((!sk[29]) & (!g3495) & (g3496)) + ((!sk[29]) & (g3495) & (g3496)) + ((sk[29]) & (!g3495) & (!g3496)));
	assign g3495 = (((!sk[30]) & (!g2280) & (g2598)) + ((!sk[30]) & (g2280) & (g2598)) + ((sk[30]) & (!g2280) & (g2598)));
	assign g3496 = (((!sk[31]) & (!g2085) & (g2280)) + ((!sk[31]) & (g2085) & (g2280)) + ((sk[31]) & (g2085) & (g2280)));
	assign g3497 = (((!sk[32]) & (!g3498) & (g3499)) + ((!sk[32]) & (g3498) & (g3499)) + ((sk[32]) & (!g3498) & (!g3499)));
	assign g3498 = (((!sk[33]) & (!g2280) & (g3500)) + ((!sk[33]) & (g2280) & (g3500)) + ((sk[33]) & (!g2280) & (g3500)));
	assign g3499 = (((!g2280) & (!sk[34]) & (g3501)) + ((g2280) & (!sk[34]) & (g3501)) + ((g2280) & (sk[34]) & (g3501)));
	assign g3500 = (((!dmem_dat_ix18x) & (!sk[35]) & (g2127) & (!g2550)) + ((!dmem_dat_ix18x) & (!sk[35]) & (g2127) & (g2550)) + ((!dmem_dat_ix18x) & (sk[35]) & (!g2127) & (g2550)) + ((!dmem_dat_ix18x) & (sk[35]) & (g2127) & (g2550)) + ((dmem_dat_ix18x) & (!sk[35]) & (!g2127) & (!g2550)) + ((dmem_dat_ix18x) & (!sk[35]) & (!g2127) & (g2550)) + ((dmem_dat_ix18x) & (!sk[35]) & (g2127) & (!g2550)) + ((dmem_dat_ix18x) & (!sk[35]) & (g2127) & (g2550)) + ((dmem_dat_ix18x) & (sk[35]) & (!g2127) & (g2550)) + ((dmem_dat_ix18x) & (sk[35]) & (g2127) & (!g2550)) + ((dmem_dat_ix18x) & (sk[35]) & (g2127) & (g2550)));
	assign g3501 = (((!dmem_dat_ix18x) & (!sk[36]) & (g2127) & (!g2550)) + ((!dmem_dat_ix18x) & (!sk[36]) & (g2127) & (g2550)) + ((!dmem_dat_ix18x) & (sk[36]) & (!g2127) & (g2550)) + ((!dmem_dat_ix18x) & (sk[36]) & (g2127) & (g2550)) + ((dmem_dat_ix18x) & (!sk[36]) & (!g2127) & (!g2550)) + ((dmem_dat_ix18x) & (!sk[36]) & (!g2127) & (g2550)) + ((dmem_dat_ix18x) & (!sk[36]) & (g2127) & (!g2550)) + ((dmem_dat_ix18x) & (!sk[36]) & (g2127) & (g2550)) + ((dmem_dat_ix18x) & (sk[36]) & (!g2127) & (g2550)) + ((dmem_dat_ix18x) & (sk[36]) & (g2127) & (!g2550)) + ((dmem_dat_ix18x) & (sk[36]) & (g2127) & (g2550)));
	assign g3502 = (((!g3503) & (!sk[37]) & (g3504)) + ((!g3503) & (sk[37]) & (!g3504)) + ((g3503) & (!sk[37]) & (g3504)));
	assign g3503 = (((!g3142) & (!sk[38]) & (g3505)) + ((!g3142) & (sk[38]) & (g3505)) + ((g3142) & (!sk[38]) & (g3505)));
	assign g3504 = (((!g3142) & (!sk[39]) & (g3508)) + ((g3142) & (!sk[39]) & (g3508)) + ((g3142) & (sk[39]) & (g3508)));
	assign g3505 = (((!g3506) & (!sk[40]) & (g3507)) + ((!g3506) & (sk[40]) & (!g3507)) + ((g3506) & (!sk[40]) & (g3507)));
	assign g3506 = (((!sk[41]) & (!g2125) & (g3511)) + ((!sk[41]) & (g2125) & (g3511)) + ((sk[41]) & (!g2125) & (g3511)));
	assign g3507 = (((!g2125) & (!sk[42]) & (g3512)) + ((g2125) & (!sk[42]) & (g3512)) + ((g2125) & (sk[42]) & (g3512)));
	assign g3508 = (((!sk[43]) & (!g3509) & (g3510)) + ((!sk[43]) & (g3509) & (g3510)) + ((sk[43]) & (!g3509) & (!g3510)));
	assign g3509 = (((!g2125) & (!sk[44]) & (g3513)) + ((!g2125) & (sk[44]) & (g3513)) + ((g2125) & (!sk[44]) & (g3513)));
	assign g3510 = (((!g2125) & (!sk[45]) & (g3514)) + ((g2125) & (!sk[45]) & (g3514)) + ((g2125) & (sk[45]) & (g3514)));
	assign g3511 = (((!sk[46]) & (!g2590) & (!g2085) & (!g2591) & (g2081)) + ((!sk[46]) & (!g2590) & (!g2085) & (g2591) & (g2081)) + ((!sk[46]) & (!g2590) & (g2085) & (!g2591) & (!g2081)) + ((!sk[46]) & (!g2590) & (g2085) & (!g2591) & (g2081)) + ((!sk[46]) & (!g2590) & (g2085) & (g2591) & (!g2081)) + ((!sk[46]) & (!g2590) & (g2085) & (g2591) & (g2081)) + ((!sk[46]) & (g2590) & (!g2085) & (!g2591) & (!g2081)) + ((!sk[46]) & (g2590) & (!g2085) & (!g2591) & (g2081)) + ((!sk[46]) & (g2590) & (!g2085) & (g2591) & (!g2081)) + ((!sk[46]) & (g2590) & (!g2085) & (g2591) & (g2081)) + ((!sk[46]) & (g2590) & (g2085) & (!g2591) & (!g2081)) + ((!sk[46]) & (g2590) & (g2085) & (!g2591) & (g2081)) + ((!sk[46]) & (g2590) & (g2085) & (g2591) & (!g2081)) + ((!sk[46]) & (g2590) & (g2085) & (g2591) & (g2081)) + ((sk[46]) & (!g2590) & (!g2085) & (g2591) & (!g2081)) + ((sk[46]) & (!g2590) & (g2085) & (!g2591) & (!g2081)) + ((sk[46]) & (g2590) & (!g2085) & (!g2591) & (!g2081)) + ((sk[46]) & (g2590) & (g2085) & (g2591) & (!g2081)));
	assign g3512 = (((!g2590) & (!sk[47]) & (!g2085) & (!g2594) & (g2081)) + ((!g2590) & (!sk[47]) & (!g2085) & (g2594) & (g2081)) + ((!g2590) & (!sk[47]) & (g2085) & (!g2594) & (!g2081)) + ((!g2590) & (!sk[47]) & (g2085) & (!g2594) & (g2081)) + ((!g2590) & (!sk[47]) & (g2085) & (g2594) & (!g2081)) + ((!g2590) & (!sk[47]) & (g2085) & (g2594) & (g2081)) + ((!g2590) & (sk[47]) & (!g2085) & (g2594) & (!g2081)) + ((!g2590) & (sk[47]) & (g2085) & (g2594) & (!g2081)) + ((g2590) & (!sk[47]) & (!g2085) & (!g2594) & (!g2081)) + ((g2590) & (!sk[47]) & (!g2085) & (!g2594) & (g2081)) + ((g2590) & (!sk[47]) & (!g2085) & (g2594) & (!g2081)) + ((g2590) & (!sk[47]) & (!g2085) & (g2594) & (g2081)) + ((g2590) & (!sk[47]) & (g2085) & (!g2594) & (!g2081)) + ((g2590) & (!sk[47]) & (g2085) & (!g2594) & (g2081)) + ((g2590) & (!sk[47]) & (g2085) & (g2594) & (!g2081)) + ((g2590) & (!sk[47]) & (g2085) & (g2594) & (g2081)) + ((g2590) & (sk[47]) & (!g2085) & (g2594) & (!g2081)) + ((g2590) & (sk[47]) & (g2085) & (!g2594) & (g2081)) + ((g2590) & (sk[47]) & (g2085) & (g2594) & (!g2081)) + ((g2590) & (sk[47]) & (g2085) & (g2594) & (g2081)));
	assign g3513 = (((!g2590) & (!sk[48]) & (!g2085) & (!g2591) & (g2081)) + ((!g2590) & (!sk[48]) & (!g2085) & (g2591) & (g2081)) + ((!g2590) & (!sk[48]) & (g2085) & (!g2591) & (!g2081)) + ((!g2590) & (!sk[48]) & (g2085) & (!g2591) & (g2081)) + ((!g2590) & (!sk[48]) & (g2085) & (g2591) & (!g2081)) + ((!g2590) & (!sk[48]) & (g2085) & (g2591) & (g2081)) + ((!g2590) & (sk[48]) & (!g2085) & (!g2591) & (g2081)) + ((!g2590) & (sk[48]) & (!g2085) & (g2591) & (!g2081)) + ((!g2590) & (sk[48]) & (!g2085) & (g2591) & (g2081)) + ((!g2590) & (sk[48]) & (g2085) & (!g2591) & (!g2081)) + ((!g2590) & (sk[48]) & (g2085) & (!g2591) & (g2081)) + ((!g2590) & (sk[48]) & (g2085) & (g2591) & (g2081)) + ((g2590) & (!sk[48]) & (!g2085) & (!g2591) & (!g2081)) + ((g2590) & (!sk[48]) & (!g2085) & (!g2591) & (g2081)) + ((g2590) & (!sk[48]) & (!g2085) & (g2591) & (!g2081)) + ((g2590) & (!sk[48]) & (!g2085) & (g2591) & (g2081)) + ((g2590) & (!sk[48]) & (g2085) & (!g2591) & (!g2081)) + ((g2590) & (!sk[48]) & (g2085) & (!g2591) & (g2081)) + ((g2590) & (!sk[48]) & (g2085) & (g2591) & (!g2081)) + ((g2590) & (!sk[48]) & (g2085) & (g2591) & (g2081)) + ((g2590) & (sk[48]) & (!g2085) & (!g2591) & (!g2081)) + ((g2590) & (sk[48]) & (!g2085) & (!g2591) & (g2081)) + ((g2590) & (sk[48]) & (!g2085) & (g2591) & (g2081)) + ((g2590) & (sk[48]) & (g2085) & (!g2591) & (g2081)) + ((g2590) & (sk[48]) & (g2085) & (g2591) & (!g2081)) + ((g2590) & (sk[48]) & (g2085) & (g2591) & (g2081)));
	assign g3514 = (((!g2590) & (!g2085) & (!sk[49]) & (!g2594) & (g2081)) + ((!g2590) & (!g2085) & (!sk[49]) & (g2594) & (g2081)) + ((!g2590) & (!g2085) & (sk[49]) & (g2594) & (!g2081)) + ((!g2590) & (g2085) & (!sk[49]) & (!g2594) & (!g2081)) + ((!g2590) & (g2085) & (!sk[49]) & (!g2594) & (g2081)) + ((!g2590) & (g2085) & (!sk[49]) & (g2594) & (!g2081)) + ((!g2590) & (g2085) & (!sk[49]) & (g2594) & (g2081)) + ((!g2590) & (g2085) & (sk[49]) & (g2594) & (!g2081)) + ((g2590) & (!g2085) & (!sk[49]) & (!g2594) & (!g2081)) + ((g2590) & (!g2085) & (!sk[49]) & (!g2594) & (g2081)) + ((g2590) & (!g2085) & (!sk[49]) & (g2594) & (!g2081)) + ((g2590) & (!g2085) & (!sk[49]) & (g2594) & (g2081)) + ((g2590) & (!g2085) & (sk[49]) & (g2594) & (!g2081)) + ((g2590) & (g2085) & (!sk[49]) & (!g2594) & (!g2081)) + ((g2590) & (g2085) & (!sk[49]) & (!g2594) & (g2081)) + ((g2590) & (g2085) & (!sk[49]) & (g2594) & (!g2081)) + ((g2590) & (g2085) & (!sk[49]) & (g2594) & (g2081)) + ((g2590) & (g2085) & (sk[49]) & (!g2594) & (g2081)) + ((g2590) & (g2085) & (sk[49]) & (g2594) & (!g2081)) + ((g2590) & (g2085) & (sk[49]) & (g2594) & (g2081)));
	assign g3515 = (((!g3516) & (!sk[50]) & (g3517)) + ((!g3516) & (sk[50]) & (!g3517)) + ((g3516) & (!sk[50]) & (g3517)));
	assign g3516 = (((!sk[51]) & (!g75) & (g3518)) + ((!sk[51]) & (g75) & (g3518)) + ((sk[51]) & (!g75) & (g3518)));
	assign g3517 = (((!sk[52]) & (!g75) & (g3521)) + ((!sk[52]) & (g75) & (g3521)) + ((sk[52]) & (g75) & (g3521)));
	assign g3518 = (((!g3519) & (!sk[53]) & (g3520)) + ((!g3519) & (sk[53]) & (!g3520)) + ((g3519) & (!sk[53]) & (g3520)));
	assign g3519 = (((!g2280) & (!sk[54]) & (g2583)) + ((!g2280) & (sk[54]) & (g2583)) + ((g2280) & (!sk[54]) & (g2583)));
	assign g3520 = (((!g2084) & (!sk[55]) & (g2280)) + ((g2084) & (!sk[55]) & (g2280)) + ((g2084) & (sk[55]) & (g2280)));
	assign g3521 = (((!g3522) & (!sk[56]) & (g3523)) + ((!g3522) & (sk[56]) & (!g3523)) + ((g3522) & (!sk[56]) & (g3523)));
	assign g3522 = (((!g2280) & (!sk[57]) & (g3524)) + ((!g2280) & (sk[57]) & (g3524)) + ((g2280) & (!sk[57]) & (g3524)));
	assign g3523 = (((!g2280) & (!sk[58]) & (g3525)) + ((g2280) & (!sk[58]) & (g3525)) + ((g2280) & (sk[58]) & (g3525)));
	assign g3524 = (((!sk[59]) & (!dmem_dat_ix17x) & (g2127) & (!g2550)) + ((!sk[59]) & (!dmem_dat_ix17x) & (g2127) & (g2550)) + ((!sk[59]) & (dmem_dat_ix17x) & (!g2127) & (!g2550)) + ((!sk[59]) & (dmem_dat_ix17x) & (!g2127) & (g2550)) + ((!sk[59]) & (dmem_dat_ix17x) & (g2127) & (!g2550)) + ((!sk[59]) & (dmem_dat_ix17x) & (g2127) & (g2550)) + ((sk[59]) & (!dmem_dat_ix17x) & (!g2127) & (g2550)) + ((sk[59]) & (!dmem_dat_ix17x) & (g2127) & (g2550)) + ((sk[59]) & (dmem_dat_ix17x) & (!g2127) & (g2550)) + ((sk[59]) & (dmem_dat_ix17x) & (g2127) & (!g2550)) + ((sk[59]) & (dmem_dat_ix17x) & (g2127) & (g2550)));
	assign g3525 = (((!sk[60]) & (!dmem_dat_ix17x) & (g2127) & (!g2550)) + ((!sk[60]) & (!dmem_dat_ix17x) & (g2127) & (g2550)) + ((!sk[60]) & (dmem_dat_ix17x) & (!g2127) & (!g2550)) + ((!sk[60]) & (dmem_dat_ix17x) & (!g2127) & (g2550)) + ((!sk[60]) & (dmem_dat_ix17x) & (g2127) & (!g2550)) + ((!sk[60]) & (dmem_dat_ix17x) & (g2127) & (g2550)) + ((sk[60]) & (!dmem_dat_ix17x) & (!g2127) & (g2550)) + ((sk[60]) & (!dmem_dat_ix17x) & (g2127) & (g2550)) + ((sk[60]) & (dmem_dat_ix17x) & (!g2127) & (g2550)) + ((sk[60]) & (dmem_dat_ix17x) & (g2127) & (!g2550)) + ((sk[60]) & (dmem_dat_ix17x) & (g2127) & (g2550)));
	assign g3526 = (((!sk[61]) & (!g3527) & (g3528)) + ((!sk[61]) & (g3527) & (g3528)) + ((sk[61]) & (!g3527) & (!g3528)));
	assign g3527 = (((!g2571) & (!sk[62]) & (g3529)) + ((!g2571) & (sk[62]) & (g3529)) + ((g2571) & (!sk[62]) & (g3529)));
	assign g3528 = (((!g2571) & (!sk[63]) & (g3532)) + ((g2571) & (!sk[63]) & (g3532)) + ((g2571) & (sk[63]) & (g3532)));
	assign g3529 = (((!sk[64]) & (!g3530) & (g3531)) + ((!sk[64]) & (g3530) & (g3531)) + ((sk[64]) & (!g3530) & (!g3531)));
	assign g3530 = (((!sk[65]) & (!g2125) & (g3535)) + ((!sk[65]) & (g2125) & (g3535)) + ((sk[65]) & (!g2125) & (g3535)));
	assign g3531 = (((!sk[66]) & (!g2125) & (g3536)) + ((!sk[66]) & (g2125) & (g3536)) + ((sk[66]) & (g2125) & (g3536)));
	assign g3532 = (((!g3533) & (!sk[67]) & (g3534)) + ((!g3533) & (sk[67]) & (!g3534)) + ((g3533) & (!sk[67]) & (g3534)));
	assign g3533 = (((!sk[68]) & (!g2125) & (g3537)) + ((!sk[68]) & (g2125) & (g3537)) + ((sk[68]) & (!g2125) & (g3537)));
	assign g3534 = (((!sk[69]) & (!g2125) & (g3538)) + ((!sk[69]) & (g2125) & (g3538)) + ((sk[69]) & (g2125) & (g3538)));
	assign g3535 = (((!g2555) & (!sk[70]) & (g2081) & (!g2554)) + ((!g2555) & (!sk[70]) & (g2081) & (g2554)) + ((g2555) & (!sk[70]) & (!g2081) & (!g2554)) + ((g2555) & (!sk[70]) & (!g2081) & (g2554)) + ((g2555) & (!sk[70]) & (g2081) & (!g2554)) + ((g2555) & (!sk[70]) & (g2081) & (g2554)) + ((g2555) & (sk[70]) & (g2081) & (g2554)));
	assign g3536 = (((!sk[71]) & (!g2081) & (g2578) & (!g2579)) + ((!sk[71]) & (!g2081) & (g2578) & (g2579)) + ((!sk[71]) & (g2081) & (!g2578) & (!g2579)) + ((!sk[71]) & (g2081) & (!g2578) & (g2579)) + ((!sk[71]) & (g2081) & (g2578) & (!g2579)) + ((!sk[71]) & (g2081) & (g2578) & (g2579)) + ((sk[71]) & (!g2081) & (g2578) & (!g2579)) + ((sk[71]) & (!g2081) & (g2578) & (g2579)) + ((sk[71]) & (g2081) & (!g2578) & (g2579)) + ((sk[71]) & (g2081) & (g2578) & (g2579)));
	assign g3537 = (((!sk[72]) & (!g2555) & (g2081) & (!g2554)) + ((!sk[72]) & (!g2555) & (g2081) & (g2554)) + ((!sk[72]) & (g2555) & (!g2081) & (!g2554)) + ((!sk[72]) & (g2555) & (!g2081) & (g2554)) + ((!sk[72]) & (g2555) & (g2081) & (!g2554)) + ((!sk[72]) & (g2555) & (g2081) & (g2554)) + ((sk[72]) & (!g2555) & (!g2081) & (!g2554)) + ((sk[72]) & (!g2555) & (!g2081) & (g2554)) + ((sk[72]) & (!g2555) & (g2081) & (!g2554)) + ((sk[72]) & (!g2555) & (g2081) & (g2554)) + ((sk[72]) & (g2555) & (!g2081) & (!g2554)) + ((sk[72]) & (g2555) & (!g2081) & (g2554)) + ((sk[72]) & (g2555) & (g2081) & (!g2554)));
	assign g3538 = (((!g2081) & (!sk[73]) & (g2578) & (!g2579)) + ((!g2081) & (!sk[73]) & (g2578) & (g2579)) + ((!g2081) & (sk[73]) & (g2578) & (!g2579)) + ((!g2081) & (sk[73]) & (g2578) & (g2579)) + ((g2081) & (!sk[73]) & (!g2578) & (!g2579)) + ((g2081) & (!sk[73]) & (!g2578) & (g2579)) + ((g2081) & (!sk[73]) & (g2578) & (!g2579)) + ((g2081) & (!sk[73]) & (g2578) & (g2579)) + ((g2081) & (sk[73]) & (!g2578) & (g2579)) + ((g2081) & (sk[73]) & (g2578) & (g2579)));
	assign g3539 = (((!g3540) & (!sk[74]) & (g3541)) + ((!g3540) & (sk[74]) & (!g3541)) + ((g3540) & (!sk[74]) & (g3541)));
	assign g3540 = (((!g75) & (!sk[75]) & (g3542)) + ((!g75) & (sk[75]) & (g3542)) + ((g75) & (!sk[75]) & (g3542)));
	assign g3541 = (((!sk[76]) & (!g75) & (g3545)) + ((!sk[76]) & (g75) & (g3545)) + ((sk[76]) & (g75) & (g3545)));
	assign g3542 = (((!g3543) & (!sk[77]) & (g3544)) + ((!g3543) & (sk[77]) & (!g3544)) + ((g3543) & (!sk[77]) & (g3544)));
	assign g3543 = (((!g2280) & (!sk[78]) & (g2562)) + ((!g2280) & (sk[78]) & (g2562)) + ((g2280) & (!sk[78]) & (g2562)));
	assign g3544 = (((!g2083) & (!sk[79]) & (g2280)) + ((g2083) & (!sk[79]) & (g2280)) + ((g2083) & (sk[79]) & (g2280)));
	assign g3545 = (((!g3546) & (!sk[80]) & (g3547)) + ((!g3546) & (sk[80]) & (!g3547)) + ((g3546) & (!sk[80]) & (g3547)));
	assign g3546 = (((!sk[81]) & (!g2280) & (g3548)) + ((!sk[81]) & (g2280) & (g3548)) + ((sk[81]) & (!g2280) & (g3548)));
	assign g3547 = (((!g2280) & (!sk[82]) & (g3549)) + ((g2280) & (!sk[82]) & (g3549)) + ((g2280) & (sk[82]) & (g3549)));
	assign g3548 = (((!dmem_dat_ix16x) & (!sk[83]) & (g2127) & (!g2550)) + ((!dmem_dat_ix16x) & (!sk[83]) & (g2127) & (g2550)) + ((!dmem_dat_ix16x) & (sk[83]) & (!g2127) & (g2550)) + ((!dmem_dat_ix16x) & (sk[83]) & (g2127) & (g2550)) + ((dmem_dat_ix16x) & (!sk[83]) & (!g2127) & (!g2550)) + ((dmem_dat_ix16x) & (!sk[83]) & (!g2127) & (g2550)) + ((dmem_dat_ix16x) & (!sk[83]) & (g2127) & (!g2550)) + ((dmem_dat_ix16x) & (!sk[83]) & (g2127) & (g2550)) + ((dmem_dat_ix16x) & (sk[83]) & (!g2127) & (g2550)) + ((dmem_dat_ix16x) & (sk[83]) & (g2127) & (!g2550)) + ((dmem_dat_ix16x) & (sk[83]) & (g2127) & (g2550)));
	assign g3549 = (((!dmem_dat_ix16x) & (!g2127) & (sk[84]) & (g2550)) + ((!dmem_dat_ix16x) & (g2127) & (!sk[84]) & (!g2550)) + ((!dmem_dat_ix16x) & (g2127) & (!sk[84]) & (g2550)) + ((!dmem_dat_ix16x) & (g2127) & (sk[84]) & (g2550)) + ((dmem_dat_ix16x) & (!g2127) & (!sk[84]) & (!g2550)) + ((dmem_dat_ix16x) & (!g2127) & (!sk[84]) & (g2550)) + ((dmem_dat_ix16x) & (!g2127) & (sk[84]) & (g2550)) + ((dmem_dat_ix16x) & (g2127) & (!sk[84]) & (!g2550)) + ((dmem_dat_ix16x) & (g2127) & (!sk[84]) & (g2550)) + ((dmem_dat_ix16x) & (g2127) & (sk[84]) & (!g2550)) + ((dmem_dat_ix16x) & (g2127) & (sk[84]) & (g2550)));
	assign g3550 = (((!sk[85]) & (!g3551) & (g3552)) + ((!sk[85]) & (g3551) & (g3552)) + ((sk[85]) & (!g3551) & (!g3552)));
	assign g3551 = (((!g2555) & (!sk[86]) & (g3553)) + ((!g2555) & (sk[86]) & (g3553)) + ((g2555) & (!sk[86]) & (g3553)));
	assign g3552 = (((!sk[87]) & (!g2555) & (g3556)) + ((!sk[87]) & (g2555) & (g3556)) + ((sk[87]) & (g2555) & (g3556)));
	assign g3553 = (((!sk[88]) & (!g3554) & (g3555)) + ((!sk[88]) & (g3554) & (g3555)) + ((sk[88]) & (!g3554) & (!g3555)));
	assign g3554 = (((!g2125) & (!sk[89]) & (g2554)) + ((!g2125) & (sk[89]) & (g2554)) + ((g2125) & (!sk[89]) & (g2554)));
	assign g3555 = (((!g2125) & (!sk[90]) & (g3559)) + ((g2125) & (!sk[90]) & (g3559)) + ((g2125) & (sk[90]) & (g3559)));
	assign g3556 = (((!g3557) & (!sk[91]) & (g3558)) + ((!g3557) & (sk[91]) & (!g3558)) + ((g3557) & (!sk[91]) & (g3558)));
	assign g3557 = (((!sk[92]) & (!g2125) & (g3560)) + ((!sk[92]) & (g2125) & (g3560)) + ((sk[92]) & (!g2125) & (g3560)));
	assign g3558 = (((!sk[93]) & (!g2125) & (g3561)) + ((!sk[93]) & (g2125) & (g3561)) + ((sk[93]) & (g2125) & (g3561)));
	assign g3559 = (((!g2551) & (!g2081) & (!sk[94]) & (!g2083) & (g2558)) + ((!g2551) & (!g2081) & (!sk[94]) & (g2083) & (g2558)) + ((!g2551) & (!g2081) & (sk[94]) & (!g2083) & (g2558)) + ((!g2551) & (!g2081) & (sk[94]) & (g2083) & (g2558)) + ((!g2551) & (g2081) & (!sk[94]) & (!g2083) & (!g2558)) + ((!g2551) & (g2081) & (!sk[94]) & (!g2083) & (g2558)) + ((!g2551) & (g2081) & (!sk[94]) & (g2083) & (!g2558)) + ((!g2551) & (g2081) & (!sk[94]) & (g2083) & (g2558)) + ((g2551) & (!g2081) & (!sk[94]) & (!g2083) & (!g2558)) + ((g2551) & (!g2081) & (!sk[94]) & (!g2083) & (g2558)) + ((g2551) & (!g2081) & (!sk[94]) & (g2083) & (!g2558)) + ((g2551) & (!g2081) & (!sk[94]) & (g2083) & (g2558)) + ((g2551) & (!g2081) & (sk[94]) & (!g2083) & (g2558)) + ((g2551) & (!g2081) & (sk[94]) & (g2083) & (g2558)) + ((g2551) & (g2081) & (!sk[94]) & (!g2083) & (!g2558)) + ((g2551) & (g2081) & (!sk[94]) & (!g2083) & (g2558)) + ((g2551) & (g2081) & (!sk[94]) & (g2083) & (!g2558)) + ((g2551) & (g2081) & (!sk[94]) & (g2083) & (g2558)) + ((g2551) & (g2081) & (sk[94]) & (g2083) & (!g2558)) + ((g2551) & (g2081) & (sk[94]) & (g2083) & (g2558)));
	assign g3560 = (((!g2081) & (!sk[95]) & (g2554)) + ((!g2081) & (sk[95]) & (g2554)) + ((g2081) & (!sk[95]) & (g2554)) + ((g2081) & (sk[95]) & (!g2554)));
	assign g3561 = (((!g2551) & (!sk[96]) & (!g2081) & (!g2083) & (g2558)) + ((!g2551) & (!sk[96]) & (!g2081) & (g2083) & (g2558)) + ((!g2551) & (!sk[96]) & (g2081) & (!g2083) & (!g2558)) + ((!g2551) & (!sk[96]) & (g2081) & (!g2083) & (g2558)) + ((!g2551) & (!sk[96]) & (g2081) & (g2083) & (!g2558)) + ((!g2551) & (!sk[96]) & (g2081) & (g2083) & (g2558)) + ((!g2551) & (sk[96]) & (!g2081) & (!g2083) & (g2558)) + ((!g2551) & (sk[96]) & (!g2081) & (g2083) & (g2558)) + ((g2551) & (!sk[96]) & (!g2081) & (!g2083) & (!g2558)) + ((g2551) & (!sk[96]) & (!g2081) & (!g2083) & (g2558)) + ((g2551) & (!sk[96]) & (!g2081) & (g2083) & (!g2558)) + ((g2551) & (!sk[96]) & (!g2081) & (g2083) & (g2558)) + ((g2551) & (!sk[96]) & (g2081) & (!g2083) & (!g2558)) + ((g2551) & (!sk[96]) & (g2081) & (!g2083) & (g2558)) + ((g2551) & (!sk[96]) & (g2081) & (g2083) & (!g2558)) + ((g2551) & (!sk[96]) & (g2081) & (g2083) & (g2558)) + ((g2551) & (sk[96]) & (!g2081) & (!g2083) & (g2558)) + ((g2551) & (sk[96]) & (!g2081) & (g2083) & (g2558)) + ((g2551) & (sk[96]) & (g2081) & (g2083) & (!g2558)) + ((g2551) & (sk[96]) & (g2081) & (g2083) & (g2558)));
	assign g3562 = (((!g3563) & (!sk[97]) & (g3564)) + ((!g3563) & (sk[97]) & (!g3564)) + ((g3563) & (!sk[97]) & (g3564)));
	assign g3563 = (((!g2531) & (!sk[98]) & (g3565)) + ((!g2531) & (sk[98]) & (g3565)) + ((g2531) & (!sk[98]) & (g3565)));
	assign g3564 = (((!sk[99]) & (!g2531) & (g3568)) + ((!sk[99]) & (g2531) & (g3568)) + ((sk[99]) & (g2531) & (g3568)));
	assign g3565 = (((!sk[100]) & (!g3566) & (g3567)) + ((!sk[100]) & (g3566) & (g3567)) + ((sk[100]) & (!g3566) & (!g3567)));
	assign g3566 = (((!sk[101]) & (!g2125) & (g3571)) + ((!sk[101]) & (g2125) & (g3571)) + ((sk[101]) & (!g2125) & (g3571)));
	assign g3567 = (((!g2125) & (!sk[102]) & (g3572)) + ((g2125) & (!sk[102]) & (g3572)) + ((g2125) & (sk[102]) & (g3572)));
	assign g3568 = (((!sk[103]) & (!g3569) & (g3570)) + ((!sk[103]) & (g3569) & (g3570)) + ((sk[103]) & (!g3569) & (!g3570)));
	assign g3569 = (((!sk[104]) & (!g2125) & (g3573)) + ((!sk[104]) & (g2125) & (g3573)) + ((sk[104]) & (!g2125) & (g3573)));
	assign g3570 = (((!sk[105]) & (!g2125) & (g3574)) + ((!sk[105]) & (g2125) & (g3574)) + ((sk[105]) & (g2125) & (g3574)));
	assign g3571 = (((!g2081) & (!sk[106]) & (g2530)) + ((!g2081) & (sk[106]) & (g2530)) + ((g2081) & (!sk[106]) & (g2530)));
	assign g3572 = (((!g2529) & (!g2081) & (!g2121) & (!sk[107]) & (g2535)) + ((!g2529) & (!g2081) & (!g2121) & (sk[107]) & (g2535)) + ((!g2529) & (!g2081) & (g2121) & (!sk[107]) & (g2535)) + ((!g2529) & (!g2081) & (g2121) & (sk[107]) & (g2535)) + ((!g2529) & (g2081) & (!g2121) & (!sk[107]) & (!g2535)) + ((!g2529) & (g2081) & (!g2121) & (!sk[107]) & (g2535)) + ((!g2529) & (g2081) & (g2121) & (!sk[107]) & (!g2535)) + ((!g2529) & (g2081) & (g2121) & (!sk[107]) & (g2535)) + ((g2529) & (!g2081) & (!g2121) & (!sk[107]) & (!g2535)) + ((g2529) & (!g2081) & (!g2121) & (!sk[107]) & (g2535)) + ((g2529) & (!g2081) & (!g2121) & (sk[107]) & (g2535)) + ((g2529) & (!g2081) & (g2121) & (!sk[107]) & (!g2535)) + ((g2529) & (!g2081) & (g2121) & (!sk[107]) & (g2535)) + ((g2529) & (!g2081) & (g2121) & (sk[107]) & (g2535)) + ((g2529) & (g2081) & (!g2121) & (!sk[107]) & (!g2535)) + ((g2529) & (g2081) & (!g2121) & (!sk[107]) & (g2535)) + ((g2529) & (g2081) & (g2121) & (!sk[107]) & (!g2535)) + ((g2529) & (g2081) & (g2121) & (!sk[107]) & (g2535)) + ((g2529) & (g2081) & (g2121) & (sk[107]) & (!g2535)) + ((g2529) & (g2081) & (g2121) & (sk[107]) & (g2535)));
	assign g3573 = (((!g2081) & (!sk[108]) & (g2530)) + ((!g2081) & (sk[108]) & (g2530)) + ((g2081) & (!sk[108]) & (g2530)) + ((g2081) & (sk[108]) & (!g2530)) + ((g2081) & (sk[108]) & (g2530)));
	assign g3574 = (((!g2529) & (!g2081) & (!g2121) & (!sk[109]) & (g2535)) + ((!g2529) & (!g2081) & (!g2121) & (sk[109]) & (g2535)) + ((!g2529) & (!g2081) & (g2121) & (!sk[109]) & (g2535)) + ((!g2529) & (!g2081) & (g2121) & (sk[109]) & (g2535)) + ((!g2529) & (g2081) & (!g2121) & (!sk[109]) & (!g2535)) + ((!g2529) & (g2081) & (!g2121) & (!sk[109]) & (g2535)) + ((!g2529) & (g2081) & (g2121) & (!sk[109]) & (!g2535)) + ((!g2529) & (g2081) & (g2121) & (!sk[109]) & (g2535)) + ((g2529) & (!g2081) & (!g2121) & (!sk[109]) & (!g2535)) + ((g2529) & (!g2081) & (!g2121) & (!sk[109]) & (g2535)) + ((g2529) & (!g2081) & (!g2121) & (sk[109]) & (g2535)) + ((g2529) & (!g2081) & (g2121) & (!sk[109]) & (!g2535)) + ((g2529) & (!g2081) & (g2121) & (!sk[109]) & (g2535)) + ((g2529) & (!g2081) & (g2121) & (sk[109]) & (g2535)) + ((g2529) & (g2081) & (!g2121) & (!sk[109]) & (!g2535)) + ((g2529) & (g2081) & (!g2121) & (!sk[109]) & (g2535)) + ((g2529) & (g2081) & (g2121) & (!sk[109]) & (!g2535)) + ((g2529) & (g2081) & (g2121) & (!sk[109]) & (g2535)) + ((g2529) & (g2081) & (g2121) & (sk[109]) & (!g2535)) + ((g2529) & (g2081) & (g2121) & (sk[109]) & (g2535)));
	assign g3575 = (((!g3576) & (!sk[110]) & (g3577)) + ((!g3576) & (sk[110]) & (!g3577)) + ((g3576) & (!sk[110]) & (g3577)));
	assign g3576 = (((!sk[111]) & (!g2508) & (g3578)) + ((!sk[111]) & (g2508) & (g3578)) + ((sk[111]) & (!g2508) & (g3578)));
	assign g3577 = (((!sk[112]) & (!g2508) & (g3581)) + ((!sk[112]) & (g2508) & (g3581)) + ((sk[112]) & (g2508) & (g3581)));
	assign g3578 = (((!g3579) & (!sk[113]) & (g3580)) + ((!g3579) & (sk[113]) & (!g3580)) + ((g3579) & (!sk[113]) & (g3580)));
	assign g3579 = (((!sk[114]) & (!g2125) & (g3584)) + ((!sk[114]) & (g2125) & (g3584)) + ((sk[114]) & (!g2125) & (g3584)));
	assign g3580 = (((!g2125) & (!sk[115]) & (g3585)) + ((g2125) & (!sk[115]) & (g3585)) + ((g2125) & (sk[115]) & (g3585)));
	assign g3581 = (((!g3582) & (!sk[116]) & (g3583)) + ((!g3582) & (sk[116]) & (!g3583)) + ((g3582) & (!sk[116]) & (g3583)));
	assign g3582 = (((!sk[117]) & (!g2125) & (g3586)) + ((!sk[117]) & (g2125) & (g3586)) + ((sk[117]) & (!g2125) & (g3586)));
	assign g3583 = (((!sk[118]) & (!g2125) & (g3587)) + ((!sk[118]) & (g2125) & (g3587)) + ((sk[118]) & (g2125) & (g3587)));
	assign g3584 = (((!g2485) & (g2081) & (!sk[119]) & (!g2484)) + ((!g2485) & (g2081) & (!sk[119]) & (g2484)) + ((g2485) & (!g2081) & (!sk[119]) & (!g2484)) + ((g2485) & (!g2081) & (!sk[119]) & (g2484)) + ((g2485) & (g2081) & (!sk[119]) & (!g2484)) + ((g2485) & (g2081) & (!sk[119]) & (g2484)) + ((g2485) & (g2081) & (sk[119]) & (g2484)));
	assign g3585 = (((!sk[120]) & (!g2081) & (g2512) & (!g2513)) + ((!sk[120]) & (!g2081) & (g2512) & (g2513)) + ((!sk[120]) & (g2081) & (!g2512) & (!g2513)) + ((!sk[120]) & (g2081) & (!g2512) & (g2513)) + ((!sk[120]) & (g2081) & (g2512) & (!g2513)) + ((!sk[120]) & (g2081) & (g2512) & (g2513)) + ((sk[120]) & (!g2081) & (g2512) & (!g2513)) + ((sk[120]) & (!g2081) & (g2512) & (g2513)) + ((sk[120]) & (g2081) & (!g2512) & (g2513)) + ((sk[120]) & (g2081) & (g2512) & (g2513)));
	assign g3586 = (((!g2485) & (!g2081) & (sk[121]) & (!g2484)) + ((!g2485) & (!g2081) & (sk[121]) & (g2484)) + ((!g2485) & (g2081) & (!sk[121]) & (!g2484)) + ((!g2485) & (g2081) & (!sk[121]) & (g2484)) + ((!g2485) & (g2081) & (sk[121]) & (!g2484)) + ((!g2485) & (g2081) & (sk[121]) & (g2484)) + ((g2485) & (!g2081) & (!sk[121]) & (!g2484)) + ((g2485) & (!g2081) & (!sk[121]) & (g2484)) + ((g2485) & (!g2081) & (sk[121]) & (!g2484)) + ((g2485) & (!g2081) & (sk[121]) & (g2484)) + ((g2485) & (g2081) & (!sk[121]) & (!g2484)) + ((g2485) & (g2081) & (!sk[121]) & (g2484)) + ((g2485) & (g2081) & (sk[121]) & (!g2484)));
	assign g3587 = (((!g2081) & (!sk[122]) & (g2512) & (!g2513)) + ((!g2081) & (!sk[122]) & (g2512) & (g2513)) + ((!g2081) & (sk[122]) & (g2512) & (!g2513)) + ((!g2081) & (sk[122]) & (g2512) & (g2513)) + ((g2081) & (!sk[122]) & (!g2512) & (!g2513)) + ((g2081) & (!sk[122]) & (!g2512) & (g2513)) + ((g2081) & (!sk[122]) & (g2512) & (!g2513)) + ((g2081) & (!sk[122]) & (g2512) & (g2513)) + ((g2081) & (sk[122]) & (!g2512) & (g2513)) + ((g2081) & (sk[122]) & (g2512) & (g2513)));
	assign g3588 = (((!sk[123]) & (!g3589) & (g3590)) + ((!sk[123]) & (g3589) & (g3590)) + ((sk[123]) & (!g3589) & (!g3590)));
	assign g3589 = (((!sk[124]) & (!g2485) & (g3591)) + ((!sk[124]) & (g2485) & (g3591)) + ((sk[124]) & (!g2485) & (g3591)));
	assign g3590 = (((!g2485) & (!sk[125]) & (g3594)) + ((g2485) & (!sk[125]) & (g3594)) + ((g2485) & (sk[125]) & (g3594)));
	assign g3591 = (((!sk[126]) & (!g3592) & (g3593)) + ((!sk[126]) & (g3592) & (g3593)) + ((sk[126]) & (!g3592) & (!g3593)));
	assign g3592 = (((!g2125) & (!sk[127]) & (g3597)) + ((!g2125) & (sk[127]) & (g3597)) + ((g2125) & (!sk[127]) & (g3597)));
	assign g3593 = (((!g2125) & (!sk[0]) & (g3598)) + ((g2125) & (!sk[0]) & (g3598)) + ((g2125) & (sk[0]) & (g3598)));
	assign g3594 = (((!sk[1]) & (!g3595) & (g3596)) + ((!sk[1]) & (g3595) & (g3596)) + ((sk[1]) & (!g3595) & (!g3596)));
	assign g3595 = (((!g2125) & (!sk[2]) & (g3599)) + ((!g2125) & (sk[2]) & (g3599)) + ((g2125) & (!sk[2]) & (g3599)));
	assign g3596 = (((!g2125) & (!sk[3]) & (g3600)) + ((g2125) & (!sk[3]) & (g3600)) + ((g2125) & (sk[3]) & (g3600)));
	assign g3597 = (((!g2482) & (!sk[4]) & (g2119) & (!g2483)) + ((!g2482) & (!sk[4]) & (g2119) & (g2483)) + ((!g2482) & (sk[4]) & (!g2119) & (g2483)) + ((!g2482) & (sk[4]) & (g2119) & (!g2483)) + ((g2482) & (!sk[4]) & (!g2119) & (!g2483)) + ((g2482) & (!sk[4]) & (!g2119) & (g2483)) + ((g2482) & (!sk[4]) & (g2119) & (!g2483)) + ((g2482) & (!sk[4]) & (g2119) & (g2483)) + ((g2482) & (sk[4]) & (!g2119) & (!g2483)) + ((g2482) & (sk[4]) & (g2119) & (g2483)));
	assign g3598 = (((!sk[5]) & (!g2482) & (!g2119) & (!g2488) & (g2081)) + ((!sk[5]) & (!g2482) & (!g2119) & (g2488) & (g2081)) + ((!sk[5]) & (!g2482) & (g2119) & (!g2488) & (!g2081)) + ((!sk[5]) & (!g2482) & (g2119) & (!g2488) & (g2081)) + ((!sk[5]) & (!g2482) & (g2119) & (g2488) & (!g2081)) + ((!sk[5]) & (!g2482) & (g2119) & (g2488) & (g2081)) + ((!sk[5]) & (g2482) & (!g2119) & (!g2488) & (!g2081)) + ((!sk[5]) & (g2482) & (!g2119) & (!g2488) & (g2081)) + ((!sk[5]) & (g2482) & (!g2119) & (g2488) & (!g2081)) + ((!sk[5]) & (g2482) & (!g2119) & (g2488) & (g2081)) + ((!sk[5]) & (g2482) & (g2119) & (!g2488) & (!g2081)) + ((!sk[5]) & (g2482) & (g2119) & (!g2488) & (g2081)) + ((!sk[5]) & (g2482) & (g2119) & (g2488) & (!g2081)) + ((!sk[5]) & (g2482) & (g2119) & (g2488) & (g2081)) + ((sk[5]) & (!g2482) & (!g2119) & (g2488) & (!g2081)) + ((sk[5]) & (!g2482) & (g2119) & (g2488) & (!g2081)) + ((sk[5]) & (g2482) & (!g2119) & (g2488) & (!g2081)) + ((sk[5]) & (g2482) & (g2119) & (!g2488) & (g2081)) + ((sk[5]) & (g2482) & (g2119) & (g2488) & (!g2081)) + ((sk[5]) & (g2482) & (g2119) & (g2488) & (g2081)));
	assign g3599 = (((!g2482) & (!g2119) & (!sk[6]) & (!g2483) & (g2081)) + ((!g2482) & (!g2119) & (!sk[6]) & (g2483) & (g2081)) + ((!g2482) & (!g2119) & (sk[6]) & (!g2483) & (g2081)) + ((!g2482) & (!g2119) & (sk[6]) & (g2483) & (!g2081)) + ((!g2482) & (g2119) & (!sk[6]) & (!g2483) & (!g2081)) + ((!g2482) & (g2119) & (!sk[6]) & (!g2483) & (g2081)) + ((!g2482) & (g2119) & (!sk[6]) & (g2483) & (!g2081)) + ((!g2482) & (g2119) & (!sk[6]) & (g2483) & (g2081)) + ((!g2482) & (g2119) & (sk[6]) & (!g2483) & (!g2081)) + ((!g2482) & (g2119) & (sk[6]) & (g2483) & (g2081)) + ((g2482) & (!g2119) & (!sk[6]) & (!g2483) & (!g2081)) + ((g2482) & (!g2119) & (!sk[6]) & (!g2483) & (g2081)) + ((g2482) & (!g2119) & (!sk[6]) & (g2483) & (!g2081)) + ((g2482) & (!g2119) & (!sk[6]) & (g2483) & (g2081)) + ((g2482) & (!g2119) & (sk[6]) & (!g2483) & (!g2081)) + ((g2482) & (!g2119) & (sk[6]) & (g2483) & (g2081)) + ((g2482) & (g2119) & (!sk[6]) & (!g2483) & (!g2081)) + ((g2482) & (g2119) & (!sk[6]) & (!g2483) & (g2081)) + ((g2482) & (g2119) & (!sk[6]) & (g2483) & (!g2081)) + ((g2482) & (g2119) & (!sk[6]) & (g2483) & (g2081)) + ((g2482) & (g2119) & (sk[6]) & (!g2483) & (g2081)) + ((g2482) & (g2119) & (sk[6]) & (g2483) & (!g2081)));
	assign g3600 = (((!g2482) & (!g2119) & (!sk[7]) & (!g2488) & (g2081)) + ((!g2482) & (!g2119) & (!sk[7]) & (g2488) & (g2081)) + ((!g2482) & (!g2119) & (sk[7]) & (g2488) & (!g2081)) + ((!g2482) & (g2119) & (!sk[7]) & (!g2488) & (!g2081)) + ((!g2482) & (g2119) & (!sk[7]) & (!g2488) & (g2081)) + ((!g2482) & (g2119) & (!sk[7]) & (g2488) & (!g2081)) + ((!g2482) & (g2119) & (!sk[7]) & (g2488) & (g2081)) + ((!g2482) & (g2119) & (sk[7]) & (g2488) & (!g2081)) + ((g2482) & (!g2119) & (!sk[7]) & (!g2488) & (!g2081)) + ((g2482) & (!g2119) & (!sk[7]) & (!g2488) & (g2081)) + ((g2482) & (!g2119) & (!sk[7]) & (g2488) & (!g2081)) + ((g2482) & (!g2119) & (!sk[7]) & (g2488) & (g2081)) + ((g2482) & (!g2119) & (sk[7]) & (g2488) & (!g2081)) + ((g2482) & (g2119) & (!sk[7]) & (!g2488) & (!g2081)) + ((g2482) & (g2119) & (!sk[7]) & (!g2488) & (g2081)) + ((g2482) & (g2119) & (!sk[7]) & (g2488) & (!g2081)) + ((g2482) & (g2119) & (!sk[7]) & (g2488) & (g2081)) + ((g2482) & (g2119) & (sk[7]) & (!g2488) & (g2081)) + ((g2482) & (g2119) & (sk[7]) & (g2488) & (!g2081)) + ((g2482) & (g2119) & (sk[7]) & (g2488) & (g2081)));
	assign g3601 = (((!g3602) & (!sk[8]) & (g3603)) + ((!g3602) & (sk[8]) & (!g3603)) + ((g3602) & (!sk[8]) & (g3603)));
	assign g3602 = (((!g2459) & (!sk[9]) & (g3604)) + ((!g2459) & (sk[9]) & (g3604)) + ((g2459) & (!sk[9]) & (g3604)));
	assign g3603 = (((!sk[10]) & (!g2459) & (g3607)) + ((!sk[10]) & (g2459) & (g3607)) + ((sk[10]) & (g2459) & (g3607)));
	assign g3604 = (((!sk[11]) & (!g3605) & (g3606)) + ((!sk[11]) & (g3605) & (g3606)) + ((sk[11]) & (!g3605) & (!g3606)));
	assign g3605 = (((!g2125) & (!sk[12]) & (g3610)) + ((!g2125) & (sk[12]) & (g3610)) + ((g2125) & (!sk[12]) & (g3610)));
	assign g3606 = (((!sk[13]) & (!g2125) & (g3611)) + ((!sk[13]) & (g2125) & (g3611)) + ((sk[13]) & (g2125) & (g3611)));
	assign g3607 = (((!g3608) & (!sk[14]) & (g3609)) + ((!g3608) & (sk[14]) & (!g3609)) + ((g3608) & (!sk[14]) & (g3609)));
	assign g3608 = (((!g2125) & (!sk[15]) & (g3612)) + ((!g2125) & (sk[15]) & (g3612)) + ((g2125) & (!sk[15]) & (g3612)));
	assign g3609 = (((!sk[16]) & (!g2125) & (g3613)) + ((!sk[16]) & (g2125) & (g3613)) + ((sk[16]) & (g2125) & (g3613)));
	assign g3610 = (((!g2081) & (!sk[17]) & (g2458)) + ((!g2081) & (sk[17]) & (g2458)) + ((g2081) & (!sk[17]) & (g2458)));
	assign g3611 = (((!g2457) & (!sk[18]) & (!g2081) & (!g2118) & (g2466)) + ((!g2457) & (!sk[18]) & (!g2081) & (g2118) & (g2466)) + ((!g2457) & (!sk[18]) & (g2081) & (!g2118) & (!g2466)) + ((!g2457) & (!sk[18]) & (g2081) & (!g2118) & (g2466)) + ((!g2457) & (!sk[18]) & (g2081) & (g2118) & (!g2466)) + ((!g2457) & (!sk[18]) & (g2081) & (g2118) & (g2466)) + ((!g2457) & (sk[18]) & (!g2081) & (!g2118) & (g2466)) + ((!g2457) & (sk[18]) & (!g2081) & (g2118) & (g2466)) + ((g2457) & (!sk[18]) & (!g2081) & (!g2118) & (!g2466)) + ((g2457) & (!sk[18]) & (!g2081) & (!g2118) & (g2466)) + ((g2457) & (!sk[18]) & (!g2081) & (g2118) & (!g2466)) + ((g2457) & (!sk[18]) & (!g2081) & (g2118) & (g2466)) + ((g2457) & (!sk[18]) & (g2081) & (!g2118) & (!g2466)) + ((g2457) & (!sk[18]) & (g2081) & (!g2118) & (g2466)) + ((g2457) & (!sk[18]) & (g2081) & (g2118) & (!g2466)) + ((g2457) & (!sk[18]) & (g2081) & (g2118) & (g2466)) + ((g2457) & (sk[18]) & (!g2081) & (!g2118) & (g2466)) + ((g2457) & (sk[18]) & (!g2081) & (g2118) & (g2466)) + ((g2457) & (sk[18]) & (g2081) & (g2118) & (!g2466)) + ((g2457) & (sk[18]) & (g2081) & (g2118) & (g2466)));
	assign g3612 = (((!sk[19]) & (!g2081) & (g2458)) + ((!sk[19]) & (g2081) & (g2458)) + ((sk[19]) & (!g2081) & (g2458)) + ((sk[19]) & (g2081) & (!g2458)) + ((sk[19]) & (g2081) & (g2458)));
	assign g3613 = (((!sk[20]) & (!g2457) & (!g2081) & (!g2118) & (g2466)) + ((!sk[20]) & (!g2457) & (!g2081) & (g2118) & (g2466)) + ((!sk[20]) & (!g2457) & (g2081) & (!g2118) & (!g2466)) + ((!sk[20]) & (!g2457) & (g2081) & (!g2118) & (g2466)) + ((!sk[20]) & (!g2457) & (g2081) & (g2118) & (!g2466)) + ((!sk[20]) & (!g2457) & (g2081) & (g2118) & (g2466)) + ((!sk[20]) & (g2457) & (!g2081) & (!g2118) & (!g2466)) + ((!sk[20]) & (g2457) & (!g2081) & (!g2118) & (g2466)) + ((!sk[20]) & (g2457) & (!g2081) & (g2118) & (!g2466)) + ((!sk[20]) & (g2457) & (!g2081) & (g2118) & (g2466)) + ((!sk[20]) & (g2457) & (g2081) & (!g2118) & (!g2466)) + ((!sk[20]) & (g2457) & (g2081) & (!g2118) & (g2466)) + ((!sk[20]) & (g2457) & (g2081) & (g2118) & (!g2466)) + ((!sk[20]) & (g2457) & (g2081) & (g2118) & (g2466)) + ((sk[20]) & (!g2457) & (!g2081) & (!g2118) & (g2466)) + ((sk[20]) & (!g2457) & (!g2081) & (g2118) & (g2466)) + ((sk[20]) & (g2457) & (!g2081) & (!g2118) & (g2466)) + ((sk[20]) & (g2457) & (!g2081) & (g2118) & (g2466)) + ((sk[20]) & (g2457) & (g2081) & (g2118) & (!g2466)) + ((sk[20]) & (g2457) & (g2081) & (g2118) & (g2466)));
	assign g3614 = (((!sk[21]) & (!g3615) & (g3616)) + ((!sk[21]) & (g3615) & (g3616)) + ((sk[21]) & (!g3615) & (!g3616)));
	assign g3615 = (((!sk[22]) & (!g2443) & (g3617)) + ((!sk[22]) & (g2443) & (g3617)) + ((sk[22]) & (!g2443) & (g3617)));
	assign g3616 = (((!sk[23]) & (!g2443) & (g3620)) + ((!sk[23]) & (g2443) & (g3620)) + ((sk[23]) & (g2443) & (g3620)));
	assign g3617 = (((!g3618) & (!sk[24]) & (g3619)) + ((!g3618) & (sk[24]) & (!g3619)) + ((g3618) & (!sk[24]) & (g3619)));
	assign g3618 = (((!g2125) & (!sk[25]) & (g3623)) + ((!g2125) & (sk[25]) & (g3623)) + ((g2125) & (!sk[25]) & (g3623)));
	assign g3619 = (((!sk[26]) & (!g2125) & (g3624)) + ((!sk[26]) & (g2125) & (g3624)) + ((sk[26]) & (g2125) & (g3624)));
	assign g3620 = (((!sk[27]) & (!g3621) & (g3622)) + ((!sk[27]) & (g3621) & (g3622)) + ((sk[27]) & (!g3621) & (!g3622)));
	assign g3621 = (((!g2125) & (!sk[28]) & (g3625)) + ((!g2125) & (sk[28]) & (g3625)) + ((g2125) & (!sk[28]) & (g3625)));
	assign g3622 = (((!sk[29]) & (!g2125) & (g3626)) + ((!sk[29]) & (g2125) & (g3626)) + ((sk[29]) & (g2125) & (g3626)));
	assign g3623 = (((!g2420) & (g2081) & (!sk[30]) & (!g2419)) + ((!g2420) & (g2081) & (!sk[30]) & (g2419)) + ((g2420) & (!g2081) & (!sk[30]) & (!g2419)) + ((g2420) & (!g2081) & (!sk[30]) & (g2419)) + ((g2420) & (g2081) & (!sk[30]) & (!g2419)) + ((g2420) & (g2081) & (!sk[30]) & (g2419)) + ((g2420) & (g2081) & (sk[30]) & (g2419)));
	assign g3624 = (((!g2081) & (!sk[31]) & (g2446) & (!g2447)) + ((!g2081) & (!sk[31]) & (g2446) & (g2447)) + ((!g2081) & (sk[31]) & (g2446) & (!g2447)) + ((!g2081) & (sk[31]) & (g2446) & (g2447)) + ((g2081) & (!sk[31]) & (!g2446) & (!g2447)) + ((g2081) & (!sk[31]) & (!g2446) & (g2447)) + ((g2081) & (!sk[31]) & (g2446) & (!g2447)) + ((g2081) & (!sk[31]) & (g2446) & (g2447)) + ((g2081) & (sk[31]) & (!g2446) & (g2447)) + ((g2081) & (sk[31]) & (g2446) & (g2447)));
	assign g3625 = (((!sk[32]) & (!g2420) & (g2081) & (!g2419)) + ((!sk[32]) & (!g2420) & (g2081) & (g2419)) + ((!sk[32]) & (g2420) & (!g2081) & (!g2419)) + ((!sk[32]) & (g2420) & (!g2081) & (g2419)) + ((!sk[32]) & (g2420) & (g2081) & (!g2419)) + ((!sk[32]) & (g2420) & (g2081) & (g2419)) + ((sk[32]) & (!g2420) & (!g2081) & (!g2419)) + ((sk[32]) & (!g2420) & (!g2081) & (g2419)) + ((sk[32]) & (!g2420) & (g2081) & (!g2419)) + ((sk[32]) & (!g2420) & (g2081) & (g2419)) + ((sk[32]) & (g2420) & (!g2081) & (!g2419)) + ((sk[32]) & (g2420) & (!g2081) & (g2419)) + ((sk[32]) & (g2420) & (g2081) & (!g2419)));
	assign g3626 = (((!g2081) & (g2446) & (!sk[33]) & (!g2447)) + ((!g2081) & (g2446) & (!sk[33]) & (g2447)) + ((!g2081) & (g2446) & (sk[33]) & (!g2447)) + ((!g2081) & (g2446) & (sk[33]) & (g2447)) + ((g2081) & (!g2446) & (!sk[33]) & (!g2447)) + ((g2081) & (!g2446) & (!sk[33]) & (g2447)) + ((g2081) & (!g2446) & (sk[33]) & (g2447)) + ((g2081) & (g2446) & (!sk[33]) & (!g2447)) + ((g2081) & (g2446) & (!sk[33]) & (g2447)) + ((g2081) & (g2446) & (sk[33]) & (g2447)));
	assign g3627 = (((!sk[34]) & (!g3628) & (g3629)) + ((!sk[34]) & (g3628) & (g3629)) + ((sk[34]) & (!g3628) & (!g3629)));
	assign g3628 = (((!g2356) & (!sk[35]) & (g3630)) + ((!g2356) & (sk[35]) & (g3630)) + ((g2356) & (!sk[35]) & (g3630)));
	assign g3629 = (((!sk[36]) & (!g2356) & (g3633)) + ((!sk[36]) & (g2356) & (g3633)) + ((sk[36]) & (g2356) & (g3633)));
	assign g3630 = (((!g3631) & (!sk[37]) & (g3632)) + ((!g3631) & (sk[37]) & (!g3632)) + ((g3631) & (!sk[37]) & (g3632)));
	assign g3631 = (((!g123) & (!sk[38]) & (g3636)) + ((!g123) & (sk[38]) & (g3636)) + ((g123) & (!sk[38]) & (g3636)));
	assign g3632 = (((!sk[39]) & (!g123) & (g2379)) + ((!sk[39]) & (g123) & (g2379)) + ((sk[39]) & (g123) & (g2379)));
	assign g3633 = (((!sk[40]) & (!g3634) & (g3635)) + ((!sk[40]) & (g3634) & (g3635)) + ((sk[40]) & (!g3634) & (!g3635)));
	assign g3634 = (((!g123) & (!sk[41]) & (g3637)) + ((!g123) & (sk[41]) & (g3637)) + ((g123) & (!sk[41]) & (g3637)));
	assign g3635 = (((!g123) & (!sk[42]) & (g2379)) + ((g123) & (!sk[42]) & (g2379)) + ((g123) & (sk[42]) & (g2379)));
	assign g3636 = (((!g2022) & (!sk[43]) & (g2435)) + ((!g2022) & (sk[43]) & (g2435)) + ((g2022) & (!sk[43]) & (g2435)));
	assign g3637 = (((!g2436) & (!g2028) & (!g2022) & (!sk[44]) & (g2435)) + ((!g2436) & (!g2028) & (!g2022) & (sk[44]) & (g2435)) + ((!g2436) & (!g2028) & (g2022) & (!sk[44]) & (g2435)) + ((!g2436) & (g2028) & (!g2022) & (!sk[44]) & (!g2435)) + ((!g2436) & (g2028) & (!g2022) & (!sk[44]) & (g2435)) + ((!g2436) & (g2028) & (!g2022) & (sk[44]) & (g2435)) + ((!g2436) & (g2028) & (g2022) & (!sk[44]) & (!g2435)) + ((!g2436) & (g2028) & (g2022) & (!sk[44]) & (g2435)) + ((!g2436) & (g2028) & (g2022) & (sk[44]) & (g2435)) + ((g2436) & (!g2028) & (!g2022) & (!sk[44]) & (!g2435)) + ((g2436) & (!g2028) & (!g2022) & (!sk[44]) & (g2435)) + ((g2436) & (!g2028) & (!g2022) & (sk[44]) & (g2435)) + ((g2436) & (!g2028) & (g2022) & (!sk[44]) & (!g2435)) + ((g2436) & (!g2028) & (g2022) & (!sk[44]) & (g2435)) + ((g2436) & (!g2028) & (g2022) & (sk[44]) & (!g2435)) + ((g2436) & (!g2028) & (g2022) & (sk[44]) & (g2435)) + ((g2436) & (g2028) & (!g2022) & (!sk[44]) & (!g2435)) + ((g2436) & (g2028) & (!g2022) & (!sk[44]) & (g2435)) + ((g2436) & (g2028) & (!g2022) & (sk[44]) & (g2435)) + ((g2436) & (g2028) & (g2022) & (!sk[44]) & (!g2435)) + ((g2436) & (g2028) & (g2022) & (!sk[44]) & (g2435)) + ((g2436) & (g2028) & (g2022) & (sk[44]) & (g2435)));
	assign g3638 = (((!g3639) & (!sk[45]) & (g3640)) + ((!g3639) & (sk[45]) & (!g3640)) + ((g3639) & (!sk[45]) & (g3640)));
	assign g3639 = (((!sk[46]) & (!g2420) & (g3641)) + ((!sk[46]) & (g2420) & (g3641)) + ((sk[46]) & (!g2420) & (g3641)));
	assign g3640 = (((!sk[47]) & (!g2420) & (g3644)) + ((!sk[47]) & (g2420) & (g3644)) + ((sk[47]) & (g2420) & (g3644)));
	assign g3641 = (((!sk[48]) & (!g3642) & (g3643)) + ((!sk[48]) & (g3642) & (g3643)) + ((sk[48]) & (!g3642) & (!g3643)));
	assign g3642 = (((!g2125) & (!sk[49]) & (g2419)) + ((!g2125) & (sk[49]) & (g2419)) + ((g2125) & (!sk[49]) & (g2419)));
	assign g3643 = (((!sk[50]) & (!g2125) & (g3647)) + ((!sk[50]) & (g2125) & (g3647)) + ((sk[50]) & (g2125) & (g3647)));
	assign g3644 = (((!g3645) & (!sk[51]) & (g3646)) + ((!g3645) & (sk[51]) & (!g3646)) + ((g3645) & (!sk[51]) & (g3646)));
	assign g3645 = (((!sk[52]) & (!g2125) & (g3648)) + ((!sk[52]) & (g2125) & (g3648)) + ((sk[52]) & (!g2125) & (g3648)));
	assign g3646 = (((!sk[53]) & (!g2125) & (g3649)) + ((!sk[53]) & (g2125) & (g3649)) + ((sk[53]) & (g2125) & (g3649)));
	assign g3647 = (((!g2418) & (!g2081) & (!g2110) & (!sk[54]) & (g2424)) + ((!g2418) & (!g2081) & (!g2110) & (sk[54]) & (g2424)) + ((!g2418) & (!g2081) & (g2110) & (!sk[54]) & (g2424)) + ((!g2418) & (!g2081) & (g2110) & (sk[54]) & (g2424)) + ((!g2418) & (g2081) & (!g2110) & (!sk[54]) & (!g2424)) + ((!g2418) & (g2081) & (!g2110) & (!sk[54]) & (g2424)) + ((!g2418) & (g2081) & (g2110) & (!sk[54]) & (!g2424)) + ((!g2418) & (g2081) & (g2110) & (!sk[54]) & (g2424)) + ((g2418) & (!g2081) & (!g2110) & (!sk[54]) & (!g2424)) + ((g2418) & (!g2081) & (!g2110) & (!sk[54]) & (g2424)) + ((g2418) & (!g2081) & (!g2110) & (sk[54]) & (g2424)) + ((g2418) & (!g2081) & (g2110) & (!sk[54]) & (!g2424)) + ((g2418) & (!g2081) & (g2110) & (!sk[54]) & (g2424)) + ((g2418) & (!g2081) & (g2110) & (sk[54]) & (g2424)) + ((g2418) & (g2081) & (!g2110) & (!sk[54]) & (!g2424)) + ((g2418) & (g2081) & (!g2110) & (!sk[54]) & (g2424)) + ((g2418) & (g2081) & (g2110) & (!sk[54]) & (!g2424)) + ((g2418) & (g2081) & (g2110) & (!sk[54]) & (g2424)) + ((g2418) & (g2081) & (g2110) & (sk[54]) & (!g2424)) + ((g2418) & (g2081) & (g2110) & (sk[54]) & (g2424)));
	assign g3648 = (((!g2081) & (!sk[55]) & (g2419)) + ((!g2081) & (sk[55]) & (g2419)) + ((g2081) & (!sk[55]) & (g2419)) + ((g2081) & (sk[55]) & (!g2419)));
	assign g3649 = (((!sk[56]) & (!g2418) & (!g2081) & (!g2110) & (g2424)) + ((!sk[56]) & (!g2418) & (!g2081) & (g2110) & (g2424)) + ((!sk[56]) & (!g2418) & (g2081) & (!g2110) & (!g2424)) + ((!sk[56]) & (!g2418) & (g2081) & (!g2110) & (g2424)) + ((!sk[56]) & (!g2418) & (g2081) & (g2110) & (!g2424)) + ((!sk[56]) & (!g2418) & (g2081) & (g2110) & (g2424)) + ((!sk[56]) & (g2418) & (!g2081) & (!g2110) & (!g2424)) + ((!sk[56]) & (g2418) & (!g2081) & (!g2110) & (g2424)) + ((!sk[56]) & (g2418) & (!g2081) & (g2110) & (!g2424)) + ((!sk[56]) & (g2418) & (!g2081) & (g2110) & (g2424)) + ((!sk[56]) & (g2418) & (g2081) & (!g2110) & (!g2424)) + ((!sk[56]) & (g2418) & (g2081) & (!g2110) & (g2424)) + ((!sk[56]) & (g2418) & (g2081) & (g2110) & (!g2424)) + ((!sk[56]) & (g2418) & (g2081) & (g2110) & (g2424)) + ((sk[56]) & (!g2418) & (!g2081) & (!g2110) & (g2424)) + ((sk[56]) & (!g2418) & (!g2081) & (g2110) & (g2424)) + ((sk[56]) & (g2418) & (!g2081) & (!g2110) & (g2424)) + ((sk[56]) & (g2418) & (!g2081) & (g2110) & (g2424)) + ((sk[56]) & (g2418) & (g2081) & (g2110) & (!g2424)) + ((sk[56]) & (g2418) & (g2081) & (g2110) & (g2424)));
	assign g3650 = (((!sk[57]) & (!g3651) & (g3652)) + ((!sk[57]) & (g3651) & (g3652)) + ((sk[57]) & (!g3651) & (!g3652)));
	assign g3651 = (((!sk[58]) & (!g2394) & (g3653)) + ((!sk[58]) & (g2394) & (g3653)) + ((sk[58]) & (!g2394) & (g3653)));
	assign g3652 = (((!g2394) & (!sk[59]) & (g3656)) + ((g2394) & (!sk[59]) & (g3656)) + ((g2394) & (sk[59]) & (g3656)));
	assign g3653 = (((!g3654) & (!sk[60]) & (g3655)) + ((!g3654) & (sk[60]) & (!g3655)) + ((g3654) & (!sk[60]) & (g3655)));
	assign g3654 = (((!sk[61]) & (!g2125) & (g3659)) + ((!sk[61]) & (g2125) & (g3659)) + ((sk[61]) & (!g2125) & (g3659)));
	assign g3655 = (((!sk[62]) & (!g2125) & (g3660)) + ((!sk[62]) & (g2125) & (g3660)) + ((sk[62]) & (g2125) & (g3660)));
	assign g3656 = (((!sk[63]) & (!g3657) & (g3658)) + ((!sk[63]) & (g3657) & (g3658)) + ((sk[63]) & (!g3657) & (!g3658)));
	assign g3657 = (((!g2125) & (!sk[64]) & (g3661)) + ((!g2125) & (sk[64]) & (g3661)) + ((g2125) & (!sk[64]) & (g3661)));
	assign g3658 = (((!g2125) & (!sk[65]) & (g3662)) + ((g2125) & (!sk[65]) & (g3662)) + ((g2125) & (sk[65]) & (g3662)));
	assign g3659 = (((!sk[66]) & (!g2081) & (g2393)) + ((!sk[66]) & (g2081) & (g2393)) + ((sk[66]) & (!g2081) & (g2393)));
	assign g3660 = (((!g2391) & (!g2081) & (!sk[67]) & (!g2109) & (g2398)) + ((!g2391) & (!g2081) & (!sk[67]) & (g2109) & (g2398)) + ((!g2391) & (!g2081) & (sk[67]) & (!g2109) & (g2398)) + ((!g2391) & (!g2081) & (sk[67]) & (g2109) & (g2398)) + ((!g2391) & (g2081) & (!sk[67]) & (!g2109) & (!g2398)) + ((!g2391) & (g2081) & (!sk[67]) & (!g2109) & (g2398)) + ((!g2391) & (g2081) & (!sk[67]) & (g2109) & (!g2398)) + ((!g2391) & (g2081) & (!sk[67]) & (g2109) & (g2398)) + ((g2391) & (!g2081) & (!sk[67]) & (!g2109) & (!g2398)) + ((g2391) & (!g2081) & (!sk[67]) & (!g2109) & (g2398)) + ((g2391) & (!g2081) & (!sk[67]) & (g2109) & (!g2398)) + ((g2391) & (!g2081) & (!sk[67]) & (g2109) & (g2398)) + ((g2391) & (!g2081) & (sk[67]) & (!g2109) & (g2398)) + ((g2391) & (!g2081) & (sk[67]) & (g2109) & (g2398)) + ((g2391) & (g2081) & (!sk[67]) & (!g2109) & (!g2398)) + ((g2391) & (g2081) & (!sk[67]) & (!g2109) & (g2398)) + ((g2391) & (g2081) & (!sk[67]) & (g2109) & (!g2398)) + ((g2391) & (g2081) & (!sk[67]) & (g2109) & (g2398)) + ((g2391) & (g2081) & (sk[67]) & (g2109) & (!g2398)) + ((g2391) & (g2081) & (sk[67]) & (g2109) & (g2398)));
	assign g3661 = (((!sk[68]) & (!g2081) & (g2393)) + ((!sk[68]) & (g2081) & (g2393)) + ((sk[68]) & (!g2081) & (g2393)) + ((sk[68]) & (g2081) & (!g2393)) + ((sk[68]) & (g2081) & (g2393)));
	assign g3662 = (((!g2391) & (!g2081) & (!g2109) & (!sk[69]) & (g2398)) + ((!g2391) & (!g2081) & (!g2109) & (sk[69]) & (g2398)) + ((!g2391) & (!g2081) & (g2109) & (!sk[69]) & (g2398)) + ((!g2391) & (!g2081) & (g2109) & (sk[69]) & (g2398)) + ((!g2391) & (g2081) & (!g2109) & (!sk[69]) & (!g2398)) + ((!g2391) & (g2081) & (!g2109) & (!sk[69]) & (g2398)) + ((!g2391) & (g2081) & (g2109) & (!sk[69]) & (!g2398)) + ((!g2391) & (g2081) & (g2109) & (!sk[69]) & (g2398)) + ((g2391) & (!g2081) & (!g2109) & (!sk[69]) & (!g2398)) + ((g2391) & (!g2081) & (!g2109) & (!sk[69]) & (g2398)) + ((g2391) & (!g2081) & (!g2109) & (sk[69]) & (g2398)) + ((g2391) & (!g2081) & (g2109) & (!sk[69]) & (!g2398)) + ((g2391) & (!g2081) & (g2109) & (!sk[69]) & (g2398)) + ((g2391) & (!g2081) & (g2109) & (sk[69]) & (g2398)) + ((g2391) & (g2081) & (!g2109) & (!sk[69]) & (!g2398)) + ((g2391) & (g2081) & (!g2109) & (!sk[69]) & (g2398)) + ((g2391) & (g2081) & (g2109) & (!sk[69]) & (!g2398)) + ((g2391) & (g2081) & (g2109) & (!sk[69]) & (g2398)) + ((g2391) & (g2081) & (g2109) & (sk[69]) & (!g2398)) + ((g2391) & (g2081) & (g2109) & (sk[69]) & (g2398)));
	assign g3663 = (((!g3664) & (!sk[70]) & (g3665)) + ((!g3664) & (sk[70]) & (!g3665)) + ((g3664) & (!sk[70]) & (g3665)));
	assign g3664 = (((!sk[71]) & (!g2368) & (g3666)) + ((!sk[71]) & (g2368) & (g3666)) + ((sk[71]) & (!g2368) & (g3666)));
	assign g3665 = (((!sk[72]) & (!g2368) & (g3669)) + ((!sk[72]) & (g2368) & (g3669)) + ((sk[72]) & (g2368) & (g3669)));
	assign g3666 = (((!sk[73]) & (!g3667) & (g3668)) + ((!sk[73]) & (g3667) & (g3668)) + ((sk[73]) & (!g3667) & (!g3668)));
	assign g3667 = (((!g2125) & (!sk[74]) & (g3672)) + ((!g2125) & (sk[74]) & (g3672)) + ((g2125) & (!sk[74]) & (g3672)));
	assign g3668 = (((!sk[75]) & (!g2125) & (g3673)) + ((!sk[75]) & (g2125) & (g3673)) + ((sk[75]) & (g2125) & (g3673)));
	assign g3669 = (((!sk[76]) & (!g3670) & (g3671)) + ((!sk[76]) & (g3670) & (g3671)) + ((sk[76]) & (!g3670) & (!g3671)));
	assign g3670 = (((!sk[77]) & (!g2125) & (g3674)) + ((!sk[77]) & (g2125) & (g3674)) + ((sk[77]) & (!g2125) & (g3674)));
	assign g3671 = (((!sk[78]) & (!g2125) & (g3675)) + ((!sk[78]) & (g2125) & (g3675)) + ((sk[78]) & (g2125) & (g3675)));
	assign g3672 = (((!g2365) & (!g2108) & (!g2366) & (!sk[79]) & (g2081)) + ((!g2365) & (!g2108) & (g2366) & (!sk[79]) & (g2081)) + ((!g2365) & (!g2108) & (g2366) & (sk[79]) & (!g2081)) + ((!g2365) & (g2108) & (!g2366) & (!sk[79]) & (!g2081)) + ((!g2365) & (g2108) & (!g2366) & (!sk[79]) & (g2081)) + ((!g2365) & (g2108) & (!g2366) & (sk[79]) & (!g2081)) + ((!g2365) & (g2108) & (g2366) & (!sk[79]) & (!g2081)) + ((!g2365) & (g2108) & (g2366) & (!sk[79]) & (g2081)) + ((g2365) & (!g2108) & (!g2366) & (!sk[79]) & (!g2081)) + ((g2365) & (!g2108) & (!g2366) & (!sk[79]) & (g2081)) + ((g2365) & (!g2108) & (!g2366) & (sk[79]) & (!g2081)) + ((g2365) & (!g2108) & (g2366) & (!sk[79]) & (!g2081)) + ((g2365) & (!g2108) & (g2366) & (!sk[79]) & (g2081)) + ((g2365) & (g2108) & (!g2366) & (!sk[79]) & (!g2081)) + ((g2365) & (g2108) & (!g2366) & (!sk[79]) & (g2081)) + ((g2365) & (g2108) & (g2366) & (!sk[79]) & (!g2081)) + ((g2365) & (g2108) & (g2366) & (!sk[79]) & (g2081)) + ((g2365) & (g2108) & (g2366) & (sk[79]) & (!g2081)));
	assign g3673 = (((!g2365) & (!g2108) & (!sk[80]) & (!g2371) & (g2081)) + ((!g2365) & (!g2108) & (!sk[80]) & (g2371) & (g2081)) + ((!g2365) & (!g2108) & (sk[80]) & (g2371) & (!g2081)) + ((!g2365) & (g2108) & (!sk[80]) & (!g2371) & (!g2081)) + ((!g2365) & (g2108) & (!sk[80]) & (!g2371) & (g2081)) + ((!g2365) & (g2108) & (!sk[80]) & (g2371) & (!g2081)) + ((!g2365) & (g2108) & (!sk[80]) & (g2371) & (g2081)) + ((!g2365) & (g2108) & (sk[80]) & (g2371) & (!g2081)) + ((g2365) & (!g2108) & (!sk[80]) & (!g2371) & (!g2081)) + ((g2365) & (!g2108) & (!sk[80]) & (!g2371) & (g2081)) + ((g2365) & (!g2108) & (!sk[80]) & (g2371) & (!g2081)) + ((g2365) & (!g2108) & (!sk[80]) & (g2371) & (g2081)) + ((g2365) & (!g2108) & (sk[80]) & (g2371) & (!g2081)) + ((g2365) & (g2108) & (!sk[80]) & (!g2371) & (!g2081)) + ((g2365) & (g2108) & (!sk[80]) & (!g2371) & (g2081)) + ((g2365) & (g2108) & (!sk[80]) & (g2371) & (!g2081)) + ((g2365) & (g2108) & (!sk[80]) & (g2371) & (g2081)) + ((g2365) & (g2108) & (sk[80]) & (!g2371) & (g2081)) + ((g2365) & (g2108) & (sk[80]) & (g2371) & (!g2081)) + ((g2365) & (g2108) & (sk[80]) & (g2371) & (g2081)));
	assign g3674 = (((!sk[81]) & (!g2365) & (!g2108) & (!g2366) & (g2081)) + ((!sk[81]) & (!g2365) & (!g2108) & (g2366) & (g2081)) + ((!sk[81]) & (!g2365) & (g2108) & (!g2366) & (!g2081)) + ((!sk[81]) & (!g2365) & (g2108) & (!g2366) & (g2081)) + ((!sk[81]) & (!g2365) & (g2108) & (g2366) & (!g2081)) + ((!sk[81]) & (!g2365) & (g2108) & (g2366) & (g2081)) + ((!sk[81]) & (g2365) & (!g2108) & (!g2366) & (!g2081)) + ((!sk[81]) & (g2365) & (!g2108) & (!g2366) & (g2081)) + ((!sk[81]) & (g2365) & (!g2108) & (g2366) & (!g2081)) + ((!sk[81]) & (g2365) & (!g2108) & (g2366) & (g2081)) + ((!sk[81]) & (g2365) & (g2108) & (!g2366) & (!g2081)) + ((!sk[81]) & (g2365) & (g2108) & (!g2366) & (g2081)) + ((!sk[81]) & (g2365) & (g2108) & (g2366) & (!g2081)) + ((!sk[81]) & (g2365) & (g2108) & (g2366) & (g2081)) + ((sk[81]) & (!g2365) & (!g2108) & (!g2366) & (g2081)) + ((sk[81]) & (!g2365) & (!g2108) & (g2366) & (!g2081)) + ((sk[81]) & (!g2365) & (!g2108) & (g2366) & (g2081)) + ((sk[81]) & (!g2365) & (g2108) & (!g2366) & (!g2081)) + ((sk[81]) & (!g2365) & (g2108) & (!g2366) & (g2081)) + ((sk[81]) & (!g2365) & (g2108) & (g2366) & (g2081)) + ((sk[81]) & (g2365) & (!g2108) & (!g2366) & (!g2081)) + ((sk[81]) & (g2365) & (!g2108) & (!g2366) & (g2081)) + ((sk[81]) & (g2365) & (!g2108) & (g2366) & (g2081)) + ((sk[81]) & (g2365) & (g2108) & (!g2366) & (g2081)) + ((sk[81]) & (g2365) & (g2108) & (g2366) & (!g2081)) + ((sk[81]) & (g2365) & (g2108) & (g2366) & (g2081)));
	assign g3675 = (((!sk[82]) & (!g2365) & (!g2108) & (!g2371) & (g2081)) + ((!sk[82]) & (!g2365) & (!g2108) & (g2371) & (g2081)) + ((!sk[82]) & (!g2365) & (g2108) & (!g2371) & (!g2081)) + ((!sk[82]) & (!g2365) & (g2108) & (!g2371) & (g2081)) + ((!sk[82]) & (!g2365) & (g2108) & (g2371) & (!g2081)) + ((!sk[82]) & (!g2365) & (g2108) & (g2371) & (g2081)) + ((!sk[82]) & (g2365) & (!g2108) & (!g2371) & (!g2081)) + ((!sk[82]) & (g2365) & (!g2108) & (!g2371) & (g2081)) + ((!sk[82]) & (g2365) & (!g2108) & (g2371) & (!g2081)) + ((!sk[82]) & (g2365) & (!g2108) & (g2371) & (g2081)) + ((!sk[82]) & (g2365) & (g2108) & (!g2371) & (!g2081)) + ((!sk[82]) & (g2365) & (g2108) & (!g2371) & (g2081)) + ((!sk[82]) & (g2365) & (g2108) & (g2371) & (!g2081)) + ((!sk[82]) & (g2365) & (g2108) & (g2371) & (g2081)) + ((sk[82]) & (!g2365) & (!g2108) & (g2371) & (!g2081)) + ((sk[82]) & (!g2365) & (g2108) & (g2371) & (!g2081)) + ((sk[82]) & (g2365) & (!g2108) & (g2371) & (!g2081)) + ((sk[82]) & (g2365) & (g2108) & (!g2371) & (g2081)) + ((sk[82]) & (g2365) & (g2108) & (g2371) & (!g2081)) + ((sk[82]) & (g2365) & (g2108) & (g2371) & (g2081)));
	assign g3676 = (((!g3677) & (!sk[83]) & (g3678)) + ((!g3677) & (sk[83]) & (!g3678)) + ((g3677) & (!sk[83]) & (g3678)));
	assign g3677 = (((!sk[84]) & (!g2131) & (g3679)) + ((!sk[84]) & (g2131) & (g3679)) + ((sk[84]) & (!g2131) & (g3679)));
	assign g3678 = (((!sk[85]) & (!g2131) & (g3682)) + ((!sk[85]) & (g2131) & (g3682)) + ((sk[85]) & (g2131) & (g3682)));
	assign g3679 = (((!sk[86]) & (!g3680) & (g3681)) + ((!sk[86]) & (g3680) & (g3681)) + ((sk[86]) & (!g3680) & (!g3681)));
	assign g3680 = (((!sk[87]) & (!g75) & (g3687)) + ((!sk[87]) & (g75) & (g3687)) + ((sk[87]) & (!g75) & (g3687)));
	assign g3681 = (((!sk[88]) & (!g75) & (g3685)) + ((!sk[88]) & (g75) & (g3685)) + ((sk[88]) & (g75) & (g3685)));
	assign g3682 = (((!sk[89]) & (!g3683) & (g3684)) + ((!sk[89]) & (g3683) & (g3684)) + ((sk[89]) & (!g3683) & (!g3684)));
	assign g3683 = (((!g75) & (!sk[90]) & (g3687)) + ((!g75) & (sk[90]) & (g3687)) + ((g75) & (!sk[90]) & (g3687)));
	assign g3684 = (((!g75) & (!sk[91]) & (g3686)) + ((g75) & (!sk[91]) & (g3686)) + ((g75) & (sk[91]) & (g3686)));
	assign g3685 = (((!g2127) & (!g2339) & (!dmem_dat_ix7x) & (!sk[92]) & (g2338)) + ((!g2127) & (!g2339) & (!dmem_dat_ix7x) & (sk[92]) & (g2338)) + ((!g2127) & (!g2339) & (dmem_dat_ix7x) & (!sk[92]) & (g2338)) + ((!g2127) & (!g2339) & (dmem_dat_ix7x) & (sk[92]) & (g2338)) + ((!g2127) & (g2339) & (!dmem_dat_ix7x) & (!sk[92]) & (!g2338)) + ((!g2127) & (g2339) & (!dmem_dat_ix7x) & (!sk[92]) & (g2338)) + ((!g2127) & (g2339) & (!dmem_dat_ix7x) & (sk[92]) & (!g2338)) + ((!g2127) & (g2339) & (!dmem_dat_ix7x) & (sk[92]) & (g2338)) + ((!g2127) & (g2339) & (dmem_dat_ix7x) & (!sk[92]) & (!g2338)) + ((!g2127) & (g2339) & (dmem_dat_ix7x) & (!sk[92]) & (g2338)) + ((!g2127) & (g2339) & (dmem_dat_ix7x) & (sk[92]) & (!g2338)) + ((!g2127) & (g2339) & (dmem_dat_ix7x) & (sk[92]) & (g2338)) + ((g2127) & (!g2339) & (!dmem_dat_ix7x) & (!sk[92]) & (!g2338)) + ((g2127) & (!g2339) & (!dmem_dat_ix7x) & (!sk[92]) & (g2338)) + ((g2127) & (!g2339) & (!dmem_dat_ix7x) & (sk[92]) & (g2338)) + ((g2127) & (!g2339) & (dmem_dat_ix7x) & (!sk[92]) & (!g2338)) + ((g2127) & (!g2339) & (dmem_dat_ix7x) & (!sk[92]) & (g2338)) + ((g2127) & (!g2339) & (dmem_dat_ix7x) & (sk[92]) & (!g2338)) + ((g2127) & (!g2339) & (dmem_dat_ix7x) & (sk[92]) & (g2338)) + ((g2127) & (g2339) & (!dmem_dat_ix7x) & (!sk[92]) & (!g2338)) + ((g2127) & (g2339) & (!dmem_dat_ix7x) & (!sk[92]) & (g2338)) + ((g2127) & (g2339) & (!dmem_dat_ix7x) & (sk[92]) & (!g2338)) + ((g2127) & (g2339) & (!dmem_dat_ix7x) & (sk[92]) & (g2338)) + ((g2127) & (g2339) & (dmem_dat_ix7x) & (!sk[92]) & (!g2338)) + ((g2127) & (g2339) & (dmem_dat_ix7x) & (!sk[92]) & (g2338)) + ((g2127) & (g2339) & (dmem_dat_ix7x) & (sk[92]) & (!g2338)) + ((g2127) & (g2339) & (dmem_dat_ix7x) & (sk[92]) & (g2338)));
	assign g3686 = (((!sk[93]) & (!g2127) & (g2339) & (!dmem_dat_ix7x)) + ((!sk[93]) & (!g2127) & (g2339) & (dmem_dat_ix7x)) + ((!sk[93]) & (g2127) & (!g2339) & (!dmem_dat_ix7x)) + ((!sk[93]) & (g2127) & (!g2339) & (dmem_dat_ix7x)) + ((!sk[93]) & (g2127) & (g2339) & (!dmem_dat_ix7x)) + ((!sk[93]) & (g2127) & (g2339) & (dmem_dat_ix7x)) + ((sk[93]) & (!g2127) & (g2339) & (!dmem_dat_ix7x)) + ((sk[93]) & (!g2127) & (g2339) & (dmem_dat_ix7x)) + ((sk[93]) & (g2127) & (!g2339) & (dmem_dat_ix7x)) + ((sk[93]) & (g2127) & (g2339) & (!dmem_dat_ix7x)) + ((sk[93]) & (g2127) & (g2339) & (dmem_dat_ix7x)));
	assign g3687 = (((!sk[94]) & (!g3688) & (g3689)) + ((!sk[94]) & (g3688) & (g3689)) + ((sk[94]) & (!g3688) & (!g3689)));
	assign g3688 = (((!sk[95]) & (!g2116) & (g3690)) + ((!sk[95]) & (g2116) & (g3690)) + ((sk[95]) & (!g2116) & (g3690)));
	assign g3689 = (((!g2116) & (!sk[96]) & (g3693)) + ((g2116) & (!sk[96]) & (g3693)) + ((g2116) & (sk[96]) & (g3693)));
	assign g3690 = (((!g3691) & (!sk[97]) & (g3692)) + ((!g3691) & (sk[97]) & (!g3692)) + ((g3691) & (!sk[97]) & (g3692)));
	assign g3691 = (((!sk[98]) & (!g2264) & (g3696)) + ((!sk[98]) & (g2264) & (g3696)) + ((sk[98]) & (!g2264) & (g3696)));
	assign g3692 = (((!g2264) & (!sk[99]) & (g3697)) + ((g2264) & (!sk[99]) & (g3697)) + ((g2264) & (sk[99]) & (g3697)));
	assign g3693 = (((!sk[100]) & (!g3694) & (g3695)) + ((!sk[100]) & (g3694) & (g3695)) + ((sk[100]) & (!g3694) & (!g3695)));
	assign g3694 = (((!g2264) & (!sk[101]) & (g3698)) + ((!g2264) & (sk[101]) & (g3698)) + ((g2264) & (!sk[101]) & (g3698)));
	assign g3695 = (((!sk[102]) & (!g2264) & (g3699)) + ((!sk[102]) & (g2264) & (g3699)) + ((sk[102]) & (g2264) & (g3699)));
	assign g3696 = (((!g2340) & (!sk[103]) & (!g2124) & (!g2354) & (g2280)) + ((!g2340) & (!sk[103]) & (!g2124) & (g2354) & (g2280)) + ((!g2340) & (!sk[103]) & (g2124) & (!g2354) & (!g2280)) + ((!g2340) & (!sk[103]) & (g2124) & (!g2354) & (g2280)) + ((!g2340) & (!sk[103]) & (g2124) & (g2354) & (!g2280)) + ((!g2340) & (!sk[103]) & (g2124) & (g2354) & (g2280)) + ((!g2340) & (sk[103]) & (!g2124) & (g2354) & (!g2280)) + ((g2340) & (!sk[103]) & (!g2124) & (!g2354) & (!g2280)) + ((g2340) & (!sk[103]) & (!g2124) & (!g2354) & (g2280)) + ((g2340) & (!sk[103]) & (!g2124) & (g2354) & (!g2280)) + ((g2340) & (!sk[103]) & (!g2124) & (g2354) & (g2280)) + ((g2340) & (!sk[103]) & (g2124) & (!g2354) & (!g2280)) + ((g2340) & (!sk[103]) & (g2124) & (!g2354) & (g2280)) + ((g2340) & (!sk[103]) & (g2124) & (g2354) & (!g2280)) + ((g2340) & (!sk[103]) & (g2124) & (g2354) & (g2280)) + ((g2340) & (sk[103]) & (!g2124) & (g2354) & (!g2280)) + ((g2340) & (sk[103]) & (g2124) & (!g2354) & (!g2280)) + ((g2340) & (sk[103]) & (g2124) & (g2354) & (!g2280)));
	assign g3697 = (((!g2340) & (!sk[104]) & (!g2124) & (!g3700) & (g2280)) + ((!g2340) & (!sk[104]) & (!g2124) & (g3700) & (g2280)) + ((!g2340) & (!sk[104]) & (g2124) & (!g3700) & (!g2280)) + ((!g2340) & (!sk[104]) & (g2124) & (!g3700) & (g2280)) + ((!g2340) & (!sk[104]) & (g2124) & (g3700) & (!g2280)) + ((!g2340) & (!sk[104]) & (g2124) & (g3700) & (g2280)) + ((!g2340) & (sk[104]) & (!g2124) & (g3700) & (!g2280)) + ((g2340) & (!sk[104]) & (!g2124) & (!g3700) & (!g2280)) + ((g2340) & (!sk[104]) & (!g2124) & (!g3700) & (g2280)) + ((g2340) & (!sk[104]) & (!g2124) & (g3700) & (!g2280)) + ((g2340) & (!sk[104]) & (!g2124) & (g3700) & (g2280)) + ((g2340) & (!sk[104]) & (g2124) & (!g3700) & (!g2280)) + ((g2340) & (!sk[104]) & (g2124) & (!g3700) & (g2280)) + ((g2340) & (!sk[104]) & (g2124) & (g3700) & (!g2280)) + ((g2340) & (!sk[104]) & (g2124) & (g3700) & (g2280)) + ((g2340) & (sk[104]) & (!g2124) & (g3700) & (!g2280)) + ((g2340) & (sk[104]) & (g2124) & (!g3700) & (!g2280)) + ((g2340) & (sk[104]) & (g2124) & (g3700) & (!g2280)));
	assign g3698 = (((!g2124) & (!sk[105]) & (g2354) & (!g2280)) + ((!g2124) & (!sk[105]) & (g2354) & (g2280)) + ((!g2124) & (sk[105]) & (!g2354) & (g2280)) + ((!g2124) & (sk[105]) & (g2354) & (!g2280)) + ((!g2124) & (sk[105]) & (g2354) & (g2280)) + ((g2124) & (!sk[105]) & (!g2354) & (!g2280)) + ((g2124) & (!sk[105]) & (!g2354) & (g2280)) + ((g2124) & (!sk[105]) & (g2354) & (!g2280)) + ((g2124) & (!sk[105]) & (g2354) & (g2280)) + ((g2124) & (sk[105]) & (!g2354) & (!g2280)) + ((g2124) & (sk[105]) & (!g2354) & (g2280)) + ((g2124) & (sk[105]) & (g2354) & (!g2280)) + ((g2124) & (sk[105]) & (g2354) & (g2280)));
	assign g3699 = (((!g2340) & (!g2124) & (!sk[106]) & (!g3700) & (g2280)) + ((!g2340) & (!g2124) & (!sk[106]) & (g3700) & (g2280)) + ((!g2340) & (!g2124) & (sk[106]) & (!g3700) & (g2280)) + ((!g2340) & (!g2124) & (sk[106]) & (g3700) & (!g2280)) + ((!g2340) & (!g2124) & (sk[106]) & (g3700) & (g2280)) + ((!g2340) & (g2124) & (!sk[106]) & (!g3700) & (!g2280)) + ((!g2340) & (g2124) & (!sk[106]) & (!g3700) & (g2280)) + ((!g2340) & (g2124) & (!sk[106]) & (g3700) & (!g2280)) + ((!g2340) & (g2124) & (!sk[106]) & (g3700) & (g2280)) + ((!g2340) & (g2124) & (sk[106]) & (!g3700) & (!g2280)) + ((!g2340) & (g2124) & (sk[106]) & (!g3700) & (g2280)) + ((!g2340) & (g2124) & (sk[106]) & (g3700) & (!g2280)) + ((!g2340) & (g2124) & (sk[106]) & (g3700) & (g2280)) + ((g2340) & (!g2124) & (!sk[106]) & (!g3700) & (!g2280)) + ((g2340) & (!g2124) & (!sk[106]) & (!g3700) & (g2280)) + ((g2340) & (!g2124) & (!sk[106]) & (g3700) & (!g2280)) + ((g2340) & (!g2124) & (!sk[106]) & (g3700) & (g2280)) + ((g2340) & (!g2124) & (sk[106]) & (!g3700) & (g2280)) + ((g2340) & (!g2124) & (sk[106]) & (g3700) & (!g2280)) + ((g2340) & (!g2124) & (sk[106]) & (g3700) & (g2280)) + ((g2340) & (g2124) & (!sk[106]) & (!g3700) & (!g2280)) + ((g2340) & (g2124) & (!sk[106]) & (!g3700) & (g2280)) + ((g2340) & (g2124) & (!sk[106]) & (g3700) & (!g2280)) + ((g2340) & (g2124) & (!sk[106]) & (g3700) & (g2280)) + ((g2340) & (g2124) & (sk[106]) & (!g3700) & (g2280)) + ((g2340) & (g2124) & (sk[106]) & (g3700) & (g2280)));
	assign g3700 = (((!g3701) & (!sk[107]) & (g3702)) + ((!g3701) & (sk[107]) & (!g3702)) + ((g3701) & (!sk[107]) & (g3702)));
	assign g3701 = (((!sk[108]) & (!g2342) & (g3703)) + ((!sk[108]) & (g2342) & (g3703)) + ((sk[108]) & (!g2342) & (g3703)));
	assign g3702 = (((!g2342) & (!sk[109]) & (g3706)) + ((g2342) & (!sk[109]) & (g3706)) + ((g2342) & (sk[109]) & (g3706)));
	assign g3703 = (((!sk[110]) & (!g3704) & (g3705)) + ((!sk[110]) & (g3704) & (g3705)) + ((sk[110]) & (!g3704) & (!g3705)));
	assign g3704 = (((!g2125) & (!sk[111]) & (g2341)) + ((!g2125) & (sk[111]) & (g2341)) + ((g2125) & (!sk[111]) & (g2341)));
	assign g3705 = (((!sk[112]) & (!g2125) & (g3709)) + ((!sk[112]) & (g2125) & (g3709)) + ((sk[112]) & (g2125) & (g3709)));
	assign g3706 = (((!sk[113]) & (!g3707) & (g3708)) + ((!sk[113]) & (g3707) & (g3708)) + ((sk[113]) & (!g3707) & (!g3708)));
	assign g3707 = (((!g2125) & (!sk[114]) & (g3710)) + ((!g2125) & (sk[114]) & (g3710)) + ((g2125) & (!sk[114]) & (g3710)));
	assign g3708 = (((!g2125) & (!sk[115]) & (g3711)) + ((g2125) & (!sk[115]) & (g3711)) + ((g2125) & (sk[115]) & (g3711)));
	assign g3709 = (((!sk[116]) & (!g2340) & (!g2081) & (!g2116) & (g2349)) + ((!sk[116]) & (!g2340) & (!g2081) & (g2116) & (g2349)) + ((!sk[116]) & (!g2340) & (g2081) & (!g2116) & (!g2349)) + ((!sk[116]) & (!g2340) & (g2081) & (!g2116) & (g2349)) + ((!sk[116]) & (!g2340) & (g2081) & (g2116) & (!g2349)) + ((!sk[116]) & (!g2340) & (g2081) & (g2116) & (g2349)) + ((!sk[116]) & (g2340) & (!g2081) & (!g2116) & (!g2349)) + ((!sk[116]) & (g2340) & (!g2081) & (!g2116) & (g2349)) + ((!sk[116]) & (g2340) & (!g2081) & (g2116) & (!g2349)) + ((!sk[116]) & (g2340) & (!g2081) & (g2116) & (g2349)) + ((!sk[116]) & (g2340) & (g2081) & (!g2116) & (!g2349)) + ((!sk[116]) & (g2340) & (g2081) & (!g2116) & (g2349)) + ((!sk[116]) & (g2340) & (g2081) & (g2116) & (!g2349)) + ((!sk[116]) & (g2340) & (g2081) & (g2116) & (g2349)) + ((sk[116]) & (!g2340) & (!g2081) & (!g2116) & (g2349)) + ((sk[116]) & (!g2340) & (!g2081) & (g2116) & (g2349)) + ((sk[116]) & (g2340) & (!g2081) & (!g2116) & (g2349)) + ((sk[116]) & (g2340) & (!g2081) & (g2116) & (g2349)) + ((sk[116]) & (g2340) & (g2081) & (g2116) & (!g2349)) + ((sk[116]) & (g2340) & (g2081) & (g2116) & (g2349)));
	assign g3710 = (((!sk[117]) & (!g2081) & (g2341)) + ((!sk[117]) & (g2081) & (g2341)) + ((sk[117]) & (!g2081) & (g2341)) + ((sk[117]) & (g2081) & (!g2341)));
	assign g3711 = (((!g2340) & (!g2081) & (!g2116) & (!sk[118]) & (g2349)) + ((!g2340) & (!g2081) & (!g2116) & (sk[118]) & (g2349)) + ((!g2340) & (!g2081) & (g2116) & (!sk[118]) & (g2349)) + ((!g2340) & (!g2081) & (g2116) & (sk[118]) & (g2349)) + ((!g2340) & (g2081) & (!g2116) & (!sk[118]) & (!g2349)) + ((!g2340) & (g2081) & (!g2116) & (!sk[118]) & (g2349)) + ((!g2340) & (g2081) & (g2116) & (!sk[118]) & (!g2349)) + ((!g2340) & (g2081) & (g2116) & (!sk[118]) & (g2349)) + ((g2340) & (!g2081) & (!g2116) & (!sk[118]) & (!g2349)) + ((g2340) & (!g2081) & (!g2116) & (!sk[118]) & (g2349)) + ((g2340) & (!g2081) & (!g2116) & (sk[118]) & (g2349)) + ((g2340) & (!g2081) & (g2116) & (!sk[118]) & (!g2349)) + ((g2340) & (!g2081) & (g2116) & (!sk[118]) & (g2349)) + ((g2340) & (!g2081) & (g2116) & (sk[118]) & (g2349)) + ((g2340) & (g2081) & (!g2116) & (!sk[118]) & (!g2349)) + ((g2340) & (g2081) & (!g2116) & (!sk[118]) & (g2349)) + ((g2340) & (g2081) & (g2116) & (!sk[118]) & (!g2349)) + ((g2340) & (g2081) & (g2116) & (!sk[118]) & (g2349)) + ((g2340) & (g2081) & (g2116) & (sk[118]) & (!g2349)) + ((g2340) & (g2081) & (g2116) & (sk[118]) & (g2349)));
	assign g3712 = (((!g3713) & (!sk[119]) & (g3714)) + ((!g3713) & (sk[119]) & (!g3714)) + ((g3713) & (!sk[119]) & (g3714)));
	assign g3713 = (((!g2316) & (!sk[120]) & (g3715)) + ((!g2316) & (sk[120]) & (g3715)) + ((g2316) & (!sk[120]) & (g3715)));
	assign g3714 = (((!sk[121]) & (!g2316) & (g3718)) + ((!sk[121]) & (g2316) & (g3718)) + ((sk[121]) & (g2316) & (g3718)));
	assign g3715 = (((!g3716) & (!sk[122]) & (g3717)) + ((!g3716) & (sk[122]) & (!g3717)) + ((g3716) & (!sk[122]) & (g3717)));
	assign g3716 = (((!g2125) & (!sk[123]) & (g3721)) + ((!g2125) & (sk[123]) & (g3721)) + ((g2125) & (!sk[123]) & (g3721)));
	assign g3717 = (((!sk[124]) & (!g2125) & (g3722)) + ((!sk[124]) & (g2125) & (g3722)) + ((sk[124]) & (g2125) & (g3722)));
	assign g3718 = (((!g3719) & (!sk[125]) & (g3720)) + ((!g3719) & (sk[125]) & (!g3720)) + ((g3719) & (!sk[125]) & (g3720)));
	assign g3719 = (((!g2125) & (!sk[126]) & (g3723)) + ((!g2125) & (sk[126]) & (g3723)) + ((g2125) & (!sk[126]) & (g3723)));
	assign g3720 = (((!g2125) & (!sk[127]) & (g3724)) + ((g2125) & (!sk[127]) & (g3724)) + ((g2125) & (sk[127]) & (g3724)));
	assign g3721 = (((!sk[0]) & (!g2081) & (g2315)) + ((!sk[0]) & (g2081) & (g2315)) + ((sk[0]) & (!g2081) & (g2315)));
	assign g3722 = (((!g2312) & (!g2081) & (!g2115) & (!sk[1]) & (g2319)) + ((!g2312) & (!g2081) & (!g2115) & (sk[1]) & (g2319)) + ((!g2312) & (!g2081) & (g2115) & (!sk[1]) & (g2319)) + ((!g2312) & (!g2081) & (g2115) & (sk[1]) & (g2319)) + ((!g2312) & (g2081) & (!g2115) & (!sk[1]) & (!g2319)) + ((!g2312) & (g2081) & (!g2115) & (!sk[1]) & (g2319)) + ((!g2312) & (g2081) & (g2115) & (!sk[1]) & (!g2319)) + ((!g2312) & (g2081) & (g2115) & (!sk[1]) & (g2319)) + ((g2312) & (!g2081) & (!g2115) & (!sk[1]) & (!g2319)) + ((g2312) & (!g2081) & (!g2115) & (!sk[1]) & (g2319)) + ((g2312) & (!g2081) & (!g2115) & (sk[1]) & (g2319)) + ((g2312) & (!g2081) & (g2115) & (!sk[1]) & (!g2319)) + ((g2312) & (!g2081) & (g2115) & (!sk[1]) & (g2319)) + ((g2312) & (!g2081) & (g2115) & (sk[1]) & (g2319)) + ((g2312) & (g2081) & (!g2115) & (!sk[1]) & (!g2319)) + ((g2312) & (g2081) & (!g2115) & (!sk[1]) & (g2319)) + ((g2312) & (g2081) & (g2115) & (!sk[1]) & (!g2319)) + ((g2312) & (g2081) & (g2115) & (!sk[1]) & (g2319)) + ((g2312) & (g2081) & (g2115) & (sk[1]) & (!g2319)) + ((g2312) & (g2081) & (g2115) & (sk[1]) & (g2319)));
	assign g3723 = (((!g2081) & (!sk[2]) & (g2315)) + ((!g2081) & (sk[2]) & (g2315)) + ((g2081) & (!sk[2]) & (g2315)) + ((g2081) & (sk[2]) & (!g2315)) + ((g2081) & (sk[2]) & (g2315)));
	assign g3724 = (((!g2312) & (!g2081) & (!sk[3]) & (!g2115) & (g2319)) + ((!g2312) & (!g2081) & (!sk[3]) & (g2115) & (g2319)) + ((!g2312) & (!g2081) & (sk[3]) & (!g2115) & (g2319)) + ((!g2312) & (!g2081) & (sk[3]) & (g2115) & (g2319)) + ((!g2312) & (g2081) & (!sk[3]) & (!g2115) & (!g2319)) + ((!g2312) & (g2081) & (!sk[3]) & (!g2115) & (g2319)) + ((!g2312) & (g2081) & (!sk[3]) & (g2115) & (!g2319)) + ((!g2312) & (g2081) & (!sk[3]) & (g2115) & (g2319)) + ((g2312) & (!g2081) & (!sk[3]) & (!g2115) & (!g2319)) + ((g2312) & (!g2081) & (!sk[3]) & (!g2115) & (g2319)) + ((g2312) & (!g2081) & (!sk[3]) & (g2115) & (!g2319)) + ((g2312) & (!g2081) & (!sk[3]) & (g2115) & (g2319)) + ((g2312) & (!g2081) & (sk[3]) & (!g2115) & (g2319)) + ((g2312) & (!g2081) & (sk[3]) & (g2115) & (g2319)) + ((g2312) & (g2081) & (!sk[3]) & (!g2115) & (!g2319)) + ((g2312) & (g2081) & (!sk[3]) & (!g2115) & (g2319)) + ((g2312) & (g2081) & (!sk[3]) & (g2115) & (!g2319)) + ((g2312) & (g2081) & (!sk[3]) & (g2115) & (g2319)) + ((g2312) & (g2081) & (sk[3]) & (g2115) & (!g2319)) + ((g2312) & (g2081) & (sk[3]) & (g2115) & (g2319)));
	assign g3725 = (((!sk[4]) & (!g3726) & (g3727)) + ((!sk[4]) & (g3726) & (g3727)) + ((sk[4]) & (!g3726) & (!g3727)));
	assign g3726 = (((!sk[5]) & (!g2290) & (g3728)) + ((!sk[5]) & (g2290) & (g3728)) + ((sk[5]) & (!g2290) & (g3728)));
	assign g3727 = (((!sk[6]) & (!g2290) & (g3731)) + ((!sk[6]) & (g2290) & (g3731)) + ((sk[6]) & (g2290) & (g3731)));
	assign g3728 = (((!sk[7]) & (!g3729) & (g3730)) + ((!sk[7]) & (g3729) & (g3730)) + ((sk[7]) & (!g3729) & (!g3730)));
	assign g3729 = (((!sk[8]) & (!g2125) & (g3734)) + ((!sk[8]) & (g2125) & (g3734)) + ((sk[8]) & (!g2125) & (g3734)));
	assign g3730 = (((!g2125) & (!sk[9]) & (g3735)) + ((g2125) & (!sk[9]) & (g3735)) + ((g2125) & (sk[9]) & (g3735)));
	assign g3731 = (((!g3732) & (!sk[10]) & (g3733)) + ((!g3732) & (sk[10]) & (!g3733)) + ((g3732) & (!sk[10]) & (g3733)));
	assign g3732 = (((!g2125) & (!sk[11]) & (g3736)) + ((!g2125) & (sk[11]) & (g3736)) + ((g2125) & (!sk[11]) & (g3736)));
	assign g3733 = (((!g2125) & (!sk[12]) & (g3737)) + ((g2125) & (!sk[12]) & (g3737)) + ((g2125) & (sk[12]) & (g3737)));
	assign g3734 = (((!g2267) & (!sk[13]) & (g2081) & (!g2266)) + ((!g2267) & (!sk[13]) & (g2081) & (g2266)) + ((g2267) & (!sk[13]) & (!g2081) & (!g2266)) + ((g2267) & (!sk[13]) & (!g2081) & (g2266)) + ((g2267) & (!sk[13]) & (g2081) & (!g2266)) + ((g2267) & (!sk[13]) & (g2081) & (g2266)) + ((g2267) & (sk[13]) & (g2081) & (g2266)));
	assign g3735 = (((!sk[14]) & (!g2081) & (g2294) & (!g2295)) + ((!sk[14]) & (!g2081) & (g2294) & (g2295)) + ((!sk[14]) & (g2081) & (!g2294) & (!g2295)) + ((!sk[14]) & (g2081) & (!g2294) & (g2295)) + ((!sk[14]) & (g2081) & (g2294) & (!g2295)) + ((!sk[14]) & (g2081) & (g2294) & (g2295)) + ((sk[14]) & (!g2081) & (g2294) & (!g2295)) + ((sk[14]) & (!g2081) & (g2294) & (g2295)) + ((sk[14]) & (g2081) & (!g2294) & (g2295)) + ((sk[14]) & (g2081) & (g2294) & (g2295)));
	assign g3736 = (((!g2267) & (!sk[15]) & (g2081) & (!g2266)) + ((!g2267) & (!sk[15]) & (g2081) & (g2266)) + ((!g2267) & (sk[15]) & (!g2081) & (!g2266)) + ((!g2267) & (sk[15]) & (!g2081) & (g2266)) + ((!g2267) & (sk[15]) & (g2081) & (!g2266)) + ((!g2267) & (sk[15]) & (g2081) & (g2266)) + ((g2267) & (!sk[15]) & (!g2081) & (!g2266)) + ((g2267) & (!sk[15]) & (!g2081) & (g2266)) + ((g2267) & (!sk[15]) & (g2081) & (!g2266)) + ((g2267) & (!sk[15]) & (g2081) & (g2266)) + ((g2267) & (sk[15]) & (!g2081) & (!g2266)) + ((g2267) & (sk[15]) & (!g2081) & (g2266)) + ((g2267) & (sk[15]) & (g2081) & (!g2266)));
	assign g3737 = (((!sk[16]) & (!g2081) & (g2294) & (!g2295)) + ((!sk[16]) & (!g2081) & (g2294) & (g2295)) + ((!sk[16]) & (g2081) & (!g2294) & (!g2295)) + ((!sk[16]) & (g2081) & (!g2294) & (g2295)) + ((!sk[16]) & (g2081) & (g2294) & (!g2295)) + ((!sk[16]) & (g2081) & (g2294) & (g2295)) + ((sk[16]) & (!g2081) & (g2294) & (!g2295)) + ((sk[16]) & (!g2081) & (g2294) & (g2295)) + ((sk[16]) & (g2081) & (!g2294) & (g2295)) + ((sk[16]) & (g2081) & (g2294) & (g2295)));
	assign g3738 = (((!g3739) & (!sk[17]) & (g3740)) + ((!g3739) & (sk[17]) & (!g3740)) + ((g3739) & (!sk[17]) & (g3740)));
	assign g3739 = (((!g2267) & (!sk[18]) & (g3741)) + ((!g2267) & (sk[18]) & (g3741)) + ((g2267) & (!sk[18]) & (g3741)));
	assign g3740 = (((!g2267) & (!sk[19]) & (g3744)) + ((g2267) & (!sk[19]) & (g3744)) + ((g2267) & (sk[19]) & (g3744)));
	assign g3741 = (((!sk[20]) & (!g3742) & (g3743)) + ((!sk[20]) & (g3742) & (g3743)) + ((sk[20]) & (!g3742) & (!g3743)));
	assign g3742 = (((!g2125) & (!sk[21]) & (g3747)) + ((!g2125) & (sk[21]) & (g3747)) + ((g2125) & (!sk[21]) & (g3747)));
	assign g3743 = (((!g2125) & (!sk[22]) & (g3748)) + ((g2125) & (!sk[22]) & (g3748)) + ((g2125) & (sk[22]) & (g3748)));
	assign g3744 = (((!sk[23]) & (!g3745) & (g3746)) + ((!sk[23]) & (g3745) & (g3746)) + ((sk[23]) & (!g3745) & (!g3746)));
	assign g3745 = (((!g2125) & (!sk[24]) & (g3749)) + ((!g2125) & (sk[24]) & (g3749)) + ((g2125) & (!sk[24]) & (g3749)));
	assign g3746 = (((!sk[25]) & (!g2125) & (g3750)) + ((!sk[25]) & (g2125) & (g3750)) + ((sk[25]) & (g2125) & (g3750)));
	assign g3747 = (((!sk[26]) & (!g2113) & (g2073) & (!g2265)) + ((!sk[26]) & (!g2113) & (g2073) & (g2265)) + ((!sk[26]) & (g2113) & (!g2073) & (!g2265)) + ((!sk[26]) & (g2113) & (!g2073) & (g2265)) + ((!sk[26]) & (g2113) & (g2073) & (!g2265)) + ((!sk[26]) & (g2113) & (g2073) & (g2265)) + ((sk[26]) & (!g2113) & (!g2073) & (g2265)) + ((sk[26]) & (!g2113) & (g2073) & (!g2265)) + ((sk[26]) & (g2113) & (!g2073) & (!g2265)) + ((sk[26]) & (g2113) & (g2073) & (g2265)));
	assign g3748 = (((!g2113) & (!sk[27]) & (!g2073) & (!g2271) & (g2081)) + ((!g2113) & (!sk[27]) & (!g2073) & (g2271) & (g2081)) + ((!g2113) & (!sk[27]) & (g2073) & (!g2271) & (!g2081)) + ((!g2113) & (!sk[27]) & (g2073) & (!g2271) & (g2081)) + ((!g2113) & (!sk[27]) & (g2073) & (g2271) & (!g2081)) + ((!g2113) & (!sk[27]) & (g2073) & (g2271) & (g2081)) + ((!g2113) & (sk[27]) & (!g2073) & (g2271) & (!g2081)) + ((!g2113) & (sk[27]) & (g2073) & (g2271) & (!g2081)) + ((g2113) & (!sk[27]) & (!g2073) & (!g2271) & (!g2081)) + ((g2113) & (!sk[27]) & (!g2073) & (!g2271) & (g2081)) + ((g2113) & (!sk[27]) & (!g2073) & (g2271) & (!g2081)) + ((g2113) & (!sk[27]) & (!g2073) & (g2271) & (g2081)) + ((g2113) & (!sk[27]) & (g2073) & (!g2271) & (!g2081)) + ((g2113) & (!sk[27]) & (g2073) & (!g2271) & (g2081)) + ((g2113) & (!sk[27]) & (g2073) & (g2271) & (!g2081)) + ((g2113) & (!sk[27]) & (g2073) & (g2271) & (g2081)) + ((g2113) & (sk[27]) & (!g2073) & (g2271) & (!g2081)) + ((g2113) & (sk[27]) & (g2073) & (!g2271) & (g2081)) + ((g2113) & (sk[27]) & (g2073) & (g2271) & (!g2081)) + ((g2113) & (sk[27]) & (g2073) & (g2271) & (g2081)));
	assign g3749 = (((!g2113) & (!g2073) & (!g2265) & (!sk[28]) & (g2081)) + ((!g2113) & (!g2073) & (!g2265) & (sk[28]) & (g2081)) + ((!g2113) & (!g2073) & (g2265) & (!sk[28]) & (g2081)) + ((!g2113) & (!g2073) & (g2265) & (sk[28]) & (!g2081)) + ((!g2113) & (g2073) & (!g2265) & (!sk[28]) & (!g2081)) + ((!g2113) & (g2073) & (!g2265) & (!sk[28]) & (g2081)) + ((!g2113) & (g2073) & (!g2265) & (sk[28]) & (!g2081)) + ((!g2113) & (g2073) & (g2265) & (!sk[28]) & (!g2081)) + ((!g2113) & (g2073) & (g2265) & (!sk[28]) & (g2081)) + ((!g2113) & (g2073) & (g2265) & (sk[28]) & (g2081)) + ((g2113) & (!g2073) & (!g2265) & (!sk[28]) & (!g2081)) + ((g2113) & (!g2073) & (!g2265) & (!sk[28]) & (g2081)) + ((g2113) & (!g2073) & (!g2265) & (sk[28]) & (!g2081)) + ((g2113) & (!g2073) & (g2265) & (!sk[28]) & (!g2081)) + ((g2113) & (!g2073) & (g2265) & (!sk[28]) & (g2081)) + ((g2113) & (!g2073) & (g2265) & (sk[28]) & (g2081)) + ((g2113) & (g2073) & (!g2265) & (!sk[28]) & (!g2081)) + ((g2113) & (g2073) & (!g2265) & (!sk[28]) & (g2081)) + ((g2113) & (g2073) & (!g2265) & (sk[28]) & (g2081)) + ((g2113) & (g2073) & (g2265) & (!sk[28]) & (!g2081)) + ((g2113) & (g2073) & (g2265) & (!sk[28]) & (g2081)) + ((g2113) & (g2073) & (g2265) & (sk[28]) & (!g2081)));
	assign g3750 = (((!g2113) & (!sk[29]) & (!g2073) & (!g2271) & (g2081)) + ((!g2113) & (!sk[29]) & (!g2073) & (g2271) & (g2081)) + ((!g2113) & (!sk[29]) & (g2073) & (!g2271) & (!g2081)) + ((!g2113) & (!sk[29]) & (g2073) & (!g2271) & (g2081)) + ((!g2113) & (!sk[29]) & (g2073) & (g2271) & (!g2081)) + ((!g2113) & (!sk[29]) & (g2073) & (g2271) & (g2081)) + ((!g2113) & (sk[29]) & (!g2073) & (g2271) & (!g2081)) + ((!g2113) & (sk[29]) & (g2073) & (g2271) & (!g2081)) + ((g2113) & (!sk[29]) & (!g2073) & (!g2271) & (!g2081)) + ((g2113) & (!sk[29]) & (!g2073) & (!g2271) & (g2081)) + ((g2113) & (!sk[29]) & (!g2073) & (g2271) & (!g2081)) + ((g2113) & (!sk[29]) & (!g2073) & (g2271) & (g2081)) + ((g2113) & (!sk[29]) & (g2073) & (!g2271) & (!g2081)) + ((g2113) & (!sk[29]) & (g2073) & (!g2271) & (g2081)) + ((g2113) & (!sk[29]) & (g2073) & (g2271) & (!g2081)) + ((g2113) & (!sk[29]) & (g2073) & (g2271) & (g2081)) + ((g2113) & (sk[29]) & (!g2073) & (g2271) & (!g2081)) + ((g2113) & (sk[29]) & (g2073) & (!g2271) & (g2081)) + ((g2113) & (sk[29]) & (g2073) & (g2271) & (!g2081)) + ((g2113) & (sk[29]) & (g2073) & (g2271) & (g2081)));
	assign g3751 = (((!sk[30]) & (!g3752) & (g3753)) + ((!sk[30]) & (g3752) & (g3753)) + ((sk[30]) & (!g3752) & (!g3753)));
	assign g3752 = (((!g2240) & (!sk[31]) & (g3754)) + ((!g2240) & (sk[31]) & (g3754)) + ((g2240) & (!sk[31]) & (g3754)));
	assign g3753 = (((!sk[32]) & (!g2240) & (g3757)) + ((!sk[32]) & (g2240) & (g3757)) + ((sk[32]) & (g2240) & (g3757)));
	assign g3754 = (((!g3755) & (!sk[33]) & (g3756)) + ((!g3755) & (sk[33]) & (!g3756)) + ((g3755) & (!sk[33]) & (g3756)));
	assign g3755 = (((!g2125) & (!sk[34]) & (g3760)) + ((!g2125) & (sk[34]) & (g3760)) + ((g2125) & (!sk[34]) & (g3760)));
	assign g3756 = (((!sk[35]) & (!g2125) & (g3761)) + ((!sk[35]) & (g2125) & (g3761)) + ((sk[35]) & (g2125) & (g3761)));
	assign g3757 = (((!g3758) & (!sk[36]) & (g3759)) + ((!g3758) & (sk[36]) & (!g3759)) + ((g3758) & (!sk[36]) & (g3759)));
	assign g3758 = (((!g2125) & (!sk[37]) & (g3762)) + ((!g2125) & (sk[37]) & (g3762)) + ((g2125) & (!sk[37]) & (g3762)));
	assign g3759 = (((!g2125) & (!sk[38]) & (g3763)) + ((g2125) & (!sk[38]) & (g3763)) + ((g2125) & (sk[38]) & (g3763)));
	assign g3760 = (((!g2106) & (!sk[39]) & (g2076) & (!g2238)) + ((!g2106) & (!sk[39]) & (g2076) & (g2238)) + ((!g2106) & (sk[39]) & (!g2076) & (g2238)) + ((!g2106) & (sk[39]) & (g2076) & (!g2238)) + ((g2106) & (!sk[39]) & (!g2076) & (!g2238)) + ((g2106) & (!sk[39]) & (!g2076) & (g2238)) + ((g2106) & (!sk[39]) & (g2076) & (!g2238)) + ((g2106) & (!sk[39]) & (g2076) & (g2238)) + ((g2106) & (sk[39]) & (!g2076) & (!g2238)) + ((g2106) & (sk[39]) & (g2076) & (g2238)));
	assign g3761 = (((!g2106) & (!g2076) & (!g3143) & (!sk[40]) & (g2081)) + ((!g2106) & (!g2076) & (g3143) & (!sk[40]) & (g2081)) + ((!g2106) & (!g2076) & (g3143) & (sk[40]) & (!g2081)) + ((!g2106) & (g2076) & (!g3143) & (!sk[40]) & (!g2081)) + ((!g2106) & (g2076) & (!g3143) & (!sk[40]) & (g2081)) + ((!g2106) & (g2076) & (g3143) & (!sk[40]) & (!g2081)) + ((!g2106) & (g2076) & (g3143) & (!sk[40]) & (g2081)) + ((!g2106) & (g2076) & (g3143) & (sk[40]) & (!g2081)) + ((g2106) & (!g2076) & (!g3143) & (!sk[40]) & (!g2081)) + ((g2106) & (!g2076) & (!g3143) & (!sk[40]) & (g2081)) + ((g2106) & (!g2076) & (g3143) & (!sk[40]) & (!g2081)) + ((g2106) & (!g2076) & (g3143) & (!sk[40]) & (g2081)) + ((g2106) & (!g2076) & (g3143) & (sk[40]) & (!g2081)) + ((g2106) & (g2076) & (!g3143) & (!sk[40]) & (!g2081)) + ((g2106) & (g2076) & (!g3143) & (!sk[40]) & (g2081)) + ((g2106) & (g2076) & (!g3143) & (sk[40]) & (g2081)) + ((g2106) & (g2076) & (g3143) & (!sk[40]) & (!g2081)) + ((g2106) & (g2076) & (g3143) & (!sk[40]) & (g2081)) + ((g2106) & (g2076) & (g3143) & (sk[40]) & (!g2081)) + ((g2106) & (g2076) & (g3143) & (sk[40]) & (g2081)));
	assign g3762 = (((!g2106) & (!g2076) & (!g2238) & (!sk[41]) & (g2081)) + ((!g2106) & (!g2076) & (!g2238) & (sk[41]) & (g2081)) + ((!g2106) & (!g2076) & (g2238) & (!sk[41]) & (g2081)) + ((!g2106) & (!g2076) & (g2238) & (sk[41]) & (!g2081)) + ((!g2106) & (g2076) & (!g2238) & (!sk[41]) & (!g2081)) + ((!g2106) & (g2076) & (!g2238) & (!sk[41]) & (g2081)) + ((!g2106) & (g2076) & (!g2238) & (sk[41]) & (!g2081)) + ((!g2106) & (g2076) & (g2238) & (!sk[41]) & (!g2081)) + ((!g2106) & (g2076) & (g2238) & (!sk[41]) & (g2081)) + ((!g2106) & (g2076) & (g2238) & (sk[41]) & (g2081)) + ((g2106) & (!g2076) & (!g2238) & (!sk[41]) & (!g2081)) + ((g2106) & (!g2076) & (!g2238) & (!sk[41]) & (g2081)) + ((g2106) & (!g2076) & (!g2238) & (sk[41]) & (!g2081)) + ((g2106) & (!g2076) & (g2238) & (!sk[41]) & (!g2081)) + ((g2106) & (!g2076) & (g2238) & (!sk[41]) & (g2081)) + ((g2106) & (!g2076) & (g2238) & (sk[41]) & (g2081)) + ((g2106) & (g2076) & (!g2238) & (!sk[41]) & (!g2081)) + ((g2106) & (g2076) & (!g2238) & (!sk[41]) & (g2081)) + ((g2106) & (g2076) & (!g2238) & (sk[41]) & (g2081)) + ((g2106) & (g2076) & (g2238) & (!sk[41]) & (!g2081)) + ((g2106) & (g2076) & (g2238) & (!sk[41]) & (g2081)) + ((g2106) & (g2076) & (g2238) & (sk[41]) & (!g2081)));
	assign g3763 = (((!g2106) & (!g2076) & (!sk[42]) & (!g3143) & (g2081)) + ((!g2106) & (!g2076) & (!sk[42]) & (g3143) & (g2081)) + ((!g2106) & (!g2076) & (sk[42]) & (g3143) & (!g2081)) + ((!g2106) & (g2076) & (!sk[42]) & (!g3143) & (!g2081)) + ((!g2106) & (g2076) & (!sk[42]) & (!g3143) & (g2081)) + ((!g2106) & (g2076) & (!sk[42]) & (g3143) & (!g2081)) + ((!g2106) & (g2076) & (!sk[42]) & (g3143) & (g2081)) + ((!g2106) & (g2076) & (sk[42]) & (g3143) & (!g2081)) + ((g2106) & (!g2076) & (!sk[42]) & (!g3143) & (!g2081)) + ((g2106) & (!g2076) & (!sk[42]) & (!g3143) & (g2081)) + ((g2106) & (!g2076) & (!sk[42]) & (g3143) & (!g2081)) + ((g2106) & (!g2076) & (!sk[42]) & (g3143) & (g2081)) + ((g2106) & (!g2076) & (sk[42]) & (g3143) & (!g2081)) + ((g2106) & (g2076) & (!sk[42]) & (!g3143) & (!g2081)) + ((g2106) & (g2076) & (!sk[42]) & (!g3143) & (g2081)) + ((g2106) & (g2076) & (!sk[42]) & (g3143) & (!g2081)) + ((g2106) & (g2076) & (!sk[42]) & (g3143) & (g2081)) + ((g2106) & (g2076) & (sk[42]) & (!g3143) & (g2081)) + ((g2106) & (g2076) & (sk[42]) & (g3143) & (!g2081)) + ((g2106) & (g2076) & (sk[42]) & (g3143) & (g2081)));
	assign g3764 = (((!sk[43]) & (!g3765) & (g3766)) + ((!sk[43]) & (g3765) & (g3766)) + ((sk[43]) & (!g3765) & (!g3766)));
	assign g3765 = (((!g2214) & (!sk[44]) & (g3767)) + ((!g2214) & (sk[44]) & (g3767)) + ((g2214) & (!sk[44]) & (g3767)));
	assign g3766 = (((!sk[45]) & (!g2214) & (g3770)) + ((!sk[45]) & (g2214) & (g3770)) + ((sk[45]) & (g2214) & (g3770)));
	assign g3767 = (((!sk[46]) & (!g3768) & (g3769)) + ((!sk[46]) & (g3768) & (g3769)) + ((sk[46]) & (!g3768) & (!g3769)));
	assign g3768 = (((!sk[47]) & (!g2125) & (g3773)) + ((!sk[47]) & (g2125) & (g3773)) + ((sk[47]) & (!g2125) & (g3773)));
	assign g3769 = (((!sk[48]) & (!g2125) & (g3774)) + ((!sk[48]) & (g2125) & (g3774)) + ((sk[48]) & (g2125) & (g3774)));
	assign g3770 = (((!sk[49]) & (!g3771) & (g3772)) + ((!sk[49]) & (g3771) & (g3772)) + ((sk[49]) & (!g3771) & (!g3772)));
	assign g3771 = (((!sk[50]) & (!g2125) & (g3775)) + ((!sk[50]) & (g2125) & (g3775)) + ((sk[50]) & (!g2125) & (g3775)));
	assign g3772 = (((!g2125) & (!sk[51]) & (g3776)) + ((g2125) & (!sk[51]) & (g3776)) + ((g2125) & (sk[51]) & (g3776)));
	assign g3773 = (((!g2081) & (!sk[52]) & (g2213)) + ((!g2081) & (sk[52]) & (g2213)) + ((g2081) & (!sk[52]) & (g2213)));
	assign g3774 = (((!g2105) & (!g2081) & (!g2077) & (!sk[53]) & (g3144)) + ((!g2105) & (!g2081) & (!g2077) & (sk[53]) & (g3144)) + ((!g2105) & (!g2081) & (g2077) & (!sk[53]) & (g3144)) + ((!g2105) & (!g2081) & (g2077) & (sk[53]) & (g3144)) + ((!g2105) & (g2081) & (!g2077) & (!sk[53]) & (!g3144)) + ((!g2105) & (g2081) & (!g2077) & (!sk[53]) & (g3144)) + ((!g2105) & (g2081) & (g2077) & (!sk[53]) & (!g3144)) + ((!g2105) & (g2081) & (g2077) & (!sk[53]) & (g3144)) + ((g2105) & (!g2081) & (!g2077) & (!sk[53]) & (!g3144)) + ((g2105) & (!g2081) & (!g2077) & (!sk[53]) & (g3144)) + ((g2105) & (!g2081) & (!g2077) & (sk[53]) & (g3144)) + ((g2105) & (!g2081) & (g2077) & (!sk[53]) & (!g3144)) + ((g2105) & (!g2081) & (g2077) & (!sk[53]) & (g3144)) + ((g2105) & (!g2081) & (g2077) & (sk[53]) & (g3144)) + ((g2105) & (g2081) & (!g2077) & (!sk[53]) & (!g3144)) + ((g2105) & (g2081) & (!g2077) & (!sk[53]) & (g3144)) + ((g2105) & (g2081) & (g2077) & (!sk[53]) & (!g3144)) + ((g2105) & (g2081) & (g2077) & (!sk[53]) & (g3144)) + ((g2105) & (g2081) & (g2077) & (sk[53]) & (!g3144)) + ((g2105) & (g2081) & (g2077) & (sk[53]) & (g3144)));
	assign g3775 = (((!g2081) & (!sk[54]) & (g2213)) + ((!g2081) & (sk[54]) & (g2213)) + ((g2081) & (!sk[54]) & (g2213)) + ((g2081) & (sk[54]) & (!g2213)) + ((g2081) & (sk[54]) & (g2213)));
	assign g3776 = (((!g2105) & (!sk[55]) & (!g2081) & (!g2077) & (g3144)) + ((!g2105) & (!sk[55]) & (!g2081) & (g2077) & (g3144)) + ((!g2105) & (!sk[55]) & (g2081) & (!g2077) & (!g3144)) + ((!g2105) & (!sk[55]) & (g2081) & (!g2077) & (g3144)) + ((!g2105) & (!sk[55]) & (g2081) & (g2077) & (!g3144)) + ((!g2105) & (!sk[55]) & (g2081) & (g2077) & (g3144)) + ((!g2105) & (sk[55]) & (!g2081) & (!g2077) & (g3144)) + ((!g2105) & (sk[55]) & (!g2081) & (g2077) & (g3144)) + ((g2105) & (!sk[55]) & (!g2081) & (!g2077) & (!g3144)) + ((g2105) & (!sk[55]) & (!g2081) & (!g2077) & (g3144)) + ((g2105) & (!sk[55]) & (!g2081) & (g2077) & (!g3144)) + ((g2105) & (!sk[55]) & (!g2081) & (g2077) & (g3144)) + ((g2105) & (!sk[55]) & (g2081) & (!g2077) & (!g3144)) + ((g2105) & (!sk[55]) & (g2081) & (!g2077) & (g3144)) + ((g2105) & (!sk[55]) & (g2081) & (g2077) & (!g3144)) + ((g2105) & (!sk[55]) & (g2081) & (g2077) & (g3144)) + ((g2105) & (sk[55]) & (!g2081) & (!g2077) & (g3144)) + ((g2105) & (sk[55]) & (!g2081) & (g2077) & (g3144)) + ((g2105) & (sk[55]) & (g2081) & (g2077) & (!g3144)) + ((g2105) & (sk[55]) & (g2081) & (g2077) & (g3144)));
	assign g3777 = (((!g3778) & (!sk[56]) & (g3779)) + ((!g3778) & (sk[56]) & (!g3779)) + ((g3778) & (!sk[56]) & (g3779)));
	assign g3778 = (((!sk[57]) & (!g2130) & (g3780)) + ((!sk[57]) & (g2130) & (g3780)) + ((sk[57]) & (!g2130) & (g3780)));
	assign g3779 = (((!g2130) & (!sk[58]) & (g3783)) + ((g2130) & (!sk[58]) & (g3783)) + ((g2130) & (sk[58]) & (g3783)));
	assign g3780 = (((!g3781) & (!sk[59]) & (g3782)) + ((!g3781) & (sk[59]) & (!g3782)) + ((g3781) & (!sk[59]) & (g3782)));
	assign g3781 = (((!sk[60]) & (!g75) & (g2126)) + ((!sk[60]) & (g75) & (g2126)) + ((sk[60]) & (!g75) & (g2126)));
	assign g3782 = (((!sk[61]) & (!g75) & (g3786)) + ((!sk[61]) & (g75) & (g3786)) + ((sk[61]) & (g75) & (g3786)));
	assign g3783 = (((!sk[62]) & (!g3784) & (g3785)) + ((!sk[62]) & (g3784) & (g3785)) + ((sk[62]) & (!g3784) & (!g3785)));
	assign g3784 = (((!g75) & (!sk[63]) & (g2126)) + ((!g75) & (sk[63]) & (g2126)) + ((g75) & (!sk[63]) & (g2126)));
	assign g3785 = (((!sk[64]) & (!g75) & (g3787)) + ((!sk[64]) & (g75) & (g3787)) + ((sk[64]) & (g75) & (g3787)));
	assign g3786 = (((!g2127) & (g2133) & (!sk[65]) & (!dmem_dat_ix0x)) + ((!g2127) & (g2133) & (!sk[65]) & (dmem_dat_ix0x)) + ((!g2127) & (g2133) & (sk[65]) & (!dmem_dat_ix0x)) + ((!g2127) & (g2133) & (sk[65]) & (dmem_dat_ix0x)) + ((g2127) & (!g2133) & (!sk[65]) & (!dmem_dat_ix0x)) + ((g2127) & (!g2133) & (!sk[65]) & (dmem_dat_ix0x)) + ((g2127) & (!g2133) & (sk[65]) & (dmem_dat_ix0x)) + ((g2127) & (g2133) & (!sk[65]) & (!dmem_dat_ix0x)) + ((g2127) & (g2133) & (!sk[65]) & (dmem_dat_ix0x)) + ((g2127) & (g2133) & (sk[65]) & (!dmem_dat_ix0x)) + ((g2127) & (g2133) & (sk[65]) & (dmem_dat_ix0x)));
	assign g3787 = (((!g2127) & (!g2133) & (!sk[66]) & (!dmem_dat_ix0x) & (g2131)) + ((!g2127) & (!g2133) & (!sk[66]) & (dmem_dat_ix0x) & (g2131)) + ((!g2127) & (!g2133) & (sk[66]) & (!dmem_dat_ix0x) & (!g2131)) + ((!g2127) & (!g2133) & (sk[66]) & (dmem_dat_ix0x) & (!g2131)) + ((!g2127) & (g2133) & (!sk[66]) & (!dmem_dat_ix0x) & (!g2131)) + ((!g2127) & (g2133) & (!sk[66]) & (!dmem_dat_ix0x) & (g2131)) + ((!g2127) & (g2133) & (!sk[66]) & (dmem_dat_ix0x) & (!g2131)) + ((!g2127) & (g2133) & (!sk[66]) & (dmem_dat_ix0x) & (g2131)) + ((!g2127) & (g2133) & (sk[66]) & (!dmem_dat_ix0x) & (!g2131)) + ((!g2127) & (g2133) & (sk[66]) & (!dmem_dat_ix0x) & (g2131)) + ((!g2127) & (g2133) & (sk[66]) & (dmem_dat_ix0x) & (!g2131)) + ((!g2127) & (g2133) & (sk[66]) & (dmem_dat_ix0x) & (g2131)) + ((g2127) & (!g2133) & (!sk[66]) & (!dmem_dat_ix0x) & (!g2131)) + ((g2127) & (!g2133) & (!sk[66]) & (!dmem_dat_ix0x) & (g2131)) + ((g2127) & (!g2133) & (!sk[66]) & (dmem_dat_ix0x) & (!g2131)) + ((g2127) & (!g2133) & (!sk[66]) & (dmem_dat_ix0x) & (g2131)) + ((g2127) & (!g2133) & (sk[66]) & (!dmem_dat_ix0x) & (!g2131)) + ((g2127) & (!g2133) & (sk[66]) & (dmem_dat_ix0x) & (!g2131)) + ((g2127) & (!g2133) & (sk[66]) & (dmem_dat_ix0x) & (g2131)) + ((g2127) & (g2133) & (!sk[66]) & (!dmem_dat_ix0x) & (!g2131)) + ((g2127) & (g2133) & (!sk[66]) & (!dmem_dat_ix0x) & (g2131)) + ((g2127) & (g2133) & (!sk[66]) & (dmem_dat_ix0x) & (!g2131)) + ((g2127) & (g2133) & (!sk[66]) & (dmem_dat_ix0x) & (g2131)) + ((g2127) & (g2133) & (sk[66]) & (!dmem_dat_ix0x) & (!g2131)) + ((g2127) & (g2133) & (sk[66]) & (!dmem_dat_ix0x) & (g2131)) + ((g2127) & (g2133) & (sk[66]) & (dmem_dat_ix0x) & (!g2131)) + ((g2127) & (g2133) & (sk[66]) & (dmem_dat_ix0x) & (g2131)));
	assign g3788 = (((!g3789) & (!sk[67]) & (g3790)) + ((!g3789) & (sk[67]) & (!g3790)) + ((g3789) & (!sk[67]) & (g3790)));
	assign g3789 = (((!g2103) & (!sk[68]) & (g3791)) + ((!g2103) & (sk[68]) & (g3791)) + ((g2103) & (!sk[68]) & (g3791)));
	assign g3790 = (((!g2103) & (!sk[69]) & (g3794)) + ((g2103) & (!sk[69]) & (g3794)) + ((g2103) & (sk[69]) & (g3794)));
	assign g3791 = (((!g3792) & (!sk[70]) & (g3793)) + ((!g3792) & (sk[70]) & (!g3793)) + ((g3792) & (!sk[70]) & (g3793)));
	assign g3792 = (((!sk[71]) & (!g2080) & (g3797)) + ((!sk[71]) & (g2080) & (g3797)) + ((sk[71]) & (!g2080) & (g3797)));
	assign g3793 = (((!sk[72]) & (!g2080) & (g3798)) + ((!sk[72]) & (g2080) & (g3798)) + ((sk[72]) & (g2080) & (g3798)));
	assign g3794 = (((!sk[73]) & (!g3795) & (g3796)) + ((!sk[73]) & (g3795) & (g3796)) + ((sk[73]) & (!g3795) & (!g3796)));
	assign g3795 = (((!g2080) & (!sk[74]) & (g3799)) + ((!g2080) & (sk[74]) & (g3799)) + ((g2080) & (!sk[74]) & (g3799)));
	assign g3796 = (((!sk[75]) & (!g2080) & (g3800)) + ((!sk[75]) & (g2080) & (g3800)) + ((sk[75]) & (g2080) & (g3800)));
	assign g3797 = (((!sk[76]) & (!g2073) & (g2123)) + ((!sk[76]) & (g2073) & (g2123)) + ((sk[76]) & (!g2073) & (g2123)));
	assign g3798 = (((!g2070) & (!sk[77]) & (g2071) & (!g2081)) + ((!g2070) & (!sk[77]) & (g2071) & (g2081)) + ((!g2070) & (sk[77]) & (g2071) & (!g2081)) + ((g2070) & (!sk[77]) & (!g2071) & (!g2081)) + ((g2070) & (!sk[77]) & (!g2071) & (g2081)) + ((g2070) & (!sk[77]) & (g2071) & (!g2081)) + ((g2070) & (!sk[77]) & (g2071) & (g2081)) + ((g2070) & (sk[77]) & (!g2071) & (!g2081)) + ((g2070) & (sk[77]) & (g2071) & (g2081)));
	assign g3799 = (((!g2073) & (!sk[78]) & (g2123)) + ((!g2073) & (sk[78]) & (g2123)) + ((g2073) & (!sk[78]) & (g2123)) + ((g2073) & (sk[78]) & (!g2123)) + ((g2073) & (sk[78]) & (g2123)));
	assign g3800 = (((!g2070) & (!sk[79]) & (g2071) & (!g2081)) + ((!g2070) & (!sk[79]) & (g2071) & (g2081)) + ((!g2070) & (sk[79]) & (g2071) & (!g2081)) + ((g2070) & (!sk[79]) & (!g2071) & (!g2081)) + ((g2070) & (!sk[79]) & (!g2071) & (g2081)) + ((g2070) & (!sk[79]) & (g2071) & (!g2081)) + ((g2070) & (!sk[79]) & (g2071) & (g2081)) + ((g2070) & (sk[79]) & (!g2071) & (!g2081)) + ((g2070) & (sk[79]) & (g2071) & (g2081)));
	assign g3801 = (((!sk[80]) & (!g3802) & (g3803)) + ((!sk[80]) & (g3802) & (g3803)) + ((sk[80]) & (!g3802) & (!g3803)));
	assign g3802 = (((!sk[81]) & (!g2079) & (g3804)) + ((!sk[81]) & (g2079) & (g3804)) + ((sk[81]) & (!g2079) & (g3804)));
	assign g3803 = (((!sk[82]) & (!g2079) & (g3807)) + ((!sk[82]) & (g2079) & (g3807)) + ((sk[82]) & (g2079) & (g3807)));
	assign g3804 = (((!g3805) & (!sk[83]) & (g3806)) + ((!g3805) & (sk[83]) & (!g3806)) + ((g3805) & (!sk[83]) & (g3806)));
	assign g3805 = (((!g2080) & (!sk[84]) & (g3810)) + ((!g2080) & (sk[84]) & (g3810)) + ((g2080) & (!sk[84]) & (g3810)));
	assign g3806 = (((!g2080) & (!sk[85]) & (g3811)) + ((g2080) & (!sk[85]) & (g3811)) + ((g2080) & (sk[85]) & (g3811)));
	assign g3807 = (((!g3808) & (!sk[86]) & (g3809)) + ((!g3808) & (sk[86]) & (!g3809)) + ((g3808) & (!sk[86]) & (g3809)));
	assign g3808 = (((!sk[87]) & (!g2080) & (g3812)) + ((!sk[87]) & (g2080) & (g3812)) + ((sk[87]) & (!g2080) & (g3812)));
	assign g3809 = (((!g2080) & (!sk[88]) & (g3813)) + ((g2080) & (!sk[88]) & (g3813)) + ((g2080) & (sk[88]) & (g3813)));
	assign g3810 = (((!sk[89]) & (!g2078) & (!g2081) & (!g2073) & (g2070)) + ((!sk[89]) & (!g2078) & (!g2081) & (g2073) & (g2070)) + ((!sk[89]) & (!g2078) & (g2081) & (!g2073) & (!g2070)) + ((!sk[89]) & (!g2078) & (g2081) & (!g2073) & (g2070)) + ((!sk[89]) & (!g2078) & (g2081) & (g2073) & (!g2070)) + ((!sk[89]) & (!g2078) & (g2081) & (g2073) & (g2070)) + ((!sk[89]) & (g2078) & (!g2081) & (!g2073) & (!g2070)) + ((!sk[89]) & (g2078) & (!g2081) & (!g2073) & (g2070)) + ((!sk[89]) & (g2078) & (!g2081) & (g2073) & (!g2070)) + ((!sk[89]) & (g2078) & (!g2081) & (g2073) & (g2070)) + ((!sk[89]) & (g2078) & (g2081) & (!g2073) & (!g2070)) + ((!sk[89]) & (g2078) & (g2081) & (!g2073) & (g2070)) + ((!sk[89]) & (g2078) & (g2081) & (g2073) & (!g2070)) + ((!sk[89]) & (g2078) & (g2081) & (g2073) & (g2070)) + ((sk[89]) & (!g2078) & (!g2081) & (!g2073) & (g2070)) + ((sk[89]) & (!g2078) & (!g2081) & (g2073) & (g2070)) + ((sk[89]) & (g2078) & (!g2081) & (!g2073) & (g2070)) + ((sk[89]) & (g2078) & (!g2081) & (g2073) & (g2070)) + ((sk[89]) & (g2078) & (g2081) & (!g2073) & (!g2070)) + ((sk[89]) & (g2078) & (g2081) & (!g2073) & (g2070)));
	assign g3811 = (((!sk[90]) & (!g2071) & (g2070)) + ((!sk[90]) & (g2071) & (g2070)) + ((sk[90]) & (!g2071) & (g2070)) + ((sk[90]) & (g2071) & (!g2070)));
	assign g3812 = (((!g2078) & (!g2081) & (!g2073) & (!sk[91]) & (g2070)) + ((!g2078) & (!g2081) & (!g2073) & (sk[91]) & (g2070)) + ((!g2078) & (!g2081) & (g2073) & (!sk[91]) & (g2070)) + ((!g2078) & (!g2081) & (g2073) & (sk[91]) & (g2070)) + ((!g2078) & (g2081) & (!g2073) & (!sk[91]) & (!g2070)) + ((!g2078) & (g2081) & (!g2073) & (!sk[91]) & (g2070)) + ((!g2078) & (g2081) & (g2073) & (!sk[91]) & (!g2070)) + ((!g2078) & (g2081) & (g2073) & (!sk[91]) & (g2070)) + ((g2078) & (!g2081) & (!g2073) & (!sk[91]) & (!g2070)) + ((g2078) & (!g2081) & (!g2073) & (!sk[91]) & (g2070)) + ((g2078) & (!g2081) & (!g2073) & (sk[91]) & (g2070)) + ((g2078) & (!g2081) & (g2073) & (!sk[91]) & (!g2070)) + ((g2078) & (!g2081) & (g2073) & (!sk[91]) & (g2070)) + ((g2078) & (!g2081) & (g2073) & (sk[91]) & (g2070)) + ((g2078) & (g2081) & (!g2073) & (!sk[91]) & (!g2070)) + ((g2078) & (g2081) & (!g2073) & (!sk[91]) & (g2070)) + ((g2078) & (g2081) & (!g2073) & (sk[91]) & (!g2070)) + ((g2078) & (g2081) & (!g2073) & (sk[91]) & (g2070)) + ((g2078) & (g2081) & (g2073) & (!sk[91]) & (!g2070)) + ((g2078) & (g2081) & (g2073) & (!sk[91]) & (g2070)));
	assign g3813 = (((!sk[92]) & (!g2081) & (g2071) & (!g2070)) + ((!sk[92]) & (!g2081) & (g2071) & (g2070)) + ((!sk[92]) & (g2081) & (!g2071) & (!g2070)) + ((!sk[92]) & (g2081) & (!g2071) & (g2070)) + ((!sk[92]) & (g2081) & (g2071) & (!g2070)) + ((!sk[92]) & (g2081) & (g2071) & (g2070)) + ((sk[92]) & (!g2081) & (!g2071) & (g2070)) + ((sk[92]) & (!g2081) & (g2071) & (!g2070)) + ((sk[92]) & (g2081) & (!g2071) & (!g2070)) + ((sk[92]) & (g2081) & (g2071) & (g2070)));
	assign g3814 = (((!g3815) & (!sk[93]) & (g3816)) + ((!g3815) & (sk[93]) & (!g3816)) + ((g3815) & (!sk[93]) & (g3816)));
	assign g3815 = (((!sk[94]) & (!g75) & (g3817)) + ((!sk[94]) & (g75) & (g3817)) + ((sk[94]) & (!g75) & (g3817)));
	assign g3816 = (((!g75) & (!sk[95]) & (g3820)) + ((g75) & (!sk[95]) & (g3820)) + ((g75) & (sk[95]) & (g3820)));
	assign g3817 = (((!g3818) & (!sk[96]) & (g3819)) + ((!g3818) & (sk[96]) & (!g3819)) + ((g3818) & (!sk[96]) & (g3819)));
	assign g3818 = (((!g67) & (!sk[97]) & (g3821)) + ((!g67) & (sk[97]) & (g3821)) + ((g67) & (!sk[97]) & (g3821)));
	assign g3819 = (((!sk[98]) & (!g67) & (g3822)) + ((!sk[98]) & (g67) & (g3822)) + ((sk[98]) & (g67) & (g3822)));
	assign g3820 = (((!g67) & (!sk[99]) & (dmem_ack_i)) + ((g67) & (!sk[99]) & (dmem_ack_i)) + ((g67) & (sk[99]) & (!dmem_ack_i)));
	assign g3821 = (((!g128) & (!g74) & (!g2010) & (!sk[100]) & (g129)) + ((!g128) & (!g74) & (g2010) & (!sk[100]) & (g129)) + ((!g128) & (g74) & (!g2010) & (!sk[100]) & (!g129)) + ((!g128) & (g74) & (!g2010) & (!sk[100]) & (g129)) + ((!g128) & (g74) & (g2010) & (!sk[100]) & (!g129)) + ((!g128) & (g74) & (g2010) & (!sk[100]) & (g129)) + ((g128) & (!g74) & (!g2010) & (!sk[100]) & (!g129)) + ((g128) & (!g74) & (!g2010) & (!sk[100]) & (g129)) + ((g128) & (!g74) & (g2010) & (!sk[100]) & (!g129)) + ((g128) & (!g74) & (g2010) & (!sk[100]) & (g129)) + ((g128) & (!g74) & (g2010) & (sk[100]) & (!g129)) + ((g128) & (g74) & (!g2010) & (!sk[100]) & (!g129)) + ((g128) & (g74) & (!g2010) & (!sk[100]) & (g129)) + ((g128) & (g74) & (g2010) & (!sk[100]) & (!g129)) + ((g128) & (g74) & (g2010) & (!sk[100]) & (g129)));
	assign g3822 = (((!sk[101]) & (!dmem_ack_i) & (g129)) + ((!sk[101]) & (dmem_ack_i) & (g129)) + ((sk[101]) & (!dmem_ack_i) & (!g129)) + ((sk[101]) & (!dmem_ack_i) & (g129)) + ((sk[101]) & (dmem_ack_i) & (!g129)));
	assign g3823 = (((!sk[102]) & (!g3824) & (g3825)) + ((!sk[102]) & (g3824) & (g3825)) + ((sk[102]) & (!g3824) & (!g3825)));
	assign g3824 = (((!sk[103]) & (!g1229) & (g3826)) + ((!sk[103]) & (g1229) & (g3826)) + ((sk[103]) & (!g1229) & (g3826)));
	assign g3825 = (((!sk[104]) & (!g1229) & (g3829)) + ((!sk[104]) & (g1229) & (g3829)) + ((sk[104]) & (g1229) & (g3829)));
	assign g3826 = (((!sk[105]) & (!g3827) & (g3828)) + ((!sk[105]) & (g3827) & (g3828)) + ((sk[105]) & (!g3827) & (!g3828)));
	assign g3827 = (((!g679) & (!sk[106]) & (g3832)) + ((!g679) & (sk[106]) & (g3832)) + ((g679) & (!sk[106]) & (g3832)));
	assign g3828 = (((!g679) & (!sk[107]) & (g3833)) + ((g679) & (!sk[107]) & (g3833)) + ((g679) & (sk[107]) & (g3833)));
	assign g3829 = (((!sk[108]) & (!g3830) & (g3831)) + ((!sk[108]) & (g3830) & (g3831)) + ((sk[108]) & (!g3830) & (!g3831)));
	assign g3830 = (((!sk[109]) & (!g679) & (g3834)) + ((!sk[109]) & (g679) & (g3834)) + ((sk[109]) & (!g679) & (g3834)));
	assign g3831 = (((!sk[110]) & (!g679) & (g3835)) + ((!sk[110]) & (g679) & (g3835)) + ((sk[110]) & (g679) & (g3835)));
	assign g3832 = (((!g1319) & (!sk[111]) & (!g1231) & (!g107) & (g1274)) + ((!g1319) & (!sk[111]) & (!g1231) & (g107) & (g1274)) + ((!g1319) & (!sk[111]) & (g1231) & (!g107) & (!g1274)) + ((!g1319) & (!sk[111]) & (g1231) & (!g107) & (g1274)) + ((!g1319) & (!sk[111]) & (g1231) & (g107) & (!g1274)) + ((!g1319) & (!sk[111]) & (g1231) & (g107) & (g1274)) + ((!g1319) & (sk[111]) & (!g1231) & (g107) & (g1274)) + ((!g1319) & (sk[111]) & (g1231) & (g107) & (!g1274)) + ((!g1319) & (sk[111]) & (g1231) & (g107) & (g1274)) + ((g1319) & (!sk[111]) & (!g1231) & (!g107) & (!g1274)) + ((g1319) & (!sk[111]) & (!g1231) & (!g107) & (g1274)) + ((g1319) & (!sk[111]) & (!g1231) & (g107) & (!g1274)) + ((g1319) & (!sk[111]) & (!g1231) & (g107) & (g1274)) + ((g1319) & (!sk[111]) & (g1231) & (!g107) & (!g1274)) + ((g1319) & (!sk[111]) & (g1231) & (!g107) & (g1274)) + ((g1319) & (!sk[111]) & (g1231) & (g107) & (!g1274)) + ((g1319) & (!sk[111]) & (g1231) & (g107) & (g1274)));
	assign g3833 = (((!g1319) & (!sk[112]) & (!g1231) & (!g867) & (g1274)) + ((!g1319) & (!sk[112]) & (!g1231) & (g867) & (g1274)) + ((!g1319) & (!sk[112]) & (g1231) & (!g867) & (!g1274)) + ((!g1319) & (!sk[112]) & (g1231) & (!g867) & (g1274)) + ((!g1319) & (!sk[112]) & (g1231) & (g867) & (!g1274)) + ((!g1319) & (!sk[112]) & (g1231) & (g867) & (g1274)) + ((!g1319) & (sk[112]) & (!g1231) & (g867) & (g1274)) + ((!g1319) & (sk[112]) & (g1231) & (g867) & (!g1274)) + ((!g1319) & (sk[112]) & (g1231) & (g867) & (g1274)) + ((g1319) & (!sk[112]) & (!g1231) & (!g867) & (!g1274)) + ((g1319) & (!sk[112]) & (!g1231) & (!g867) & (g1274)) + ((g1319) & (!sk[112]) & (!g1231) & (g867) & (!g1274)) + ((g1319) & (!sk[112]) & (!g1231) & (g867) & (g1274)) + ((g1319) & (!sk[112]) & (g1231) & (!g867) & (!g1274)) + ((g1319) & (!sk[112]) & (g1231) & (!g867) & (g1274)) + ((g1319) & (!sk[112]) & (g1231) & (g867) & (!g1274)) + ((g1319) & (!sk[112]) & (g1231) & (g867) & (g1274)));
	assign g3834 = (((!g1319) & (!sk[113]) & (!g1231) & (!g107) & (g1274)) + ((!g1319) & (!sk[113]) & (!g1231) & (g107) & (g1274)) + ((!g1319) & (!sk[113]) & (g1231) & (!g107) & (!g1274)) + ((!g1319) & (!sk[113]) & (g1231) & (!g107) & (g1274)) + ((!g1319) & (!sk[113]) & (g1231) & (g107) & (!g1274)) + ((!g1319) & (!sk[113]) & (g1231) & (g107) & (g1274)) + ((!g1319) & (sk[113]) & (!g1231) & (g107) & (!g1274)) + ((!g1319) & (sk[113]) & (!g1231) & (g107) & (g1274)) + ((!g1319) & (sk[113]) & (g1231) & (g107) & (!g1274)) + ((!g1319) & (sk[113]) & (g1231) & (g107) & (g1274)) + ((g1319) & (!sk[113]) & (!g1231) & (!g107) & (!g1274)) + ((g1319) & (!sk[113]) & (!g1231) & (!g107) & (g1274)) + ((g1319) & (!sk[113]) & (!g1231) & (g107) & (!g1274)) + ((g1319) & (!sk[113]) & (!g1231) & (g107) & (g1274)) + ((g1319) & (!sk[113]) & (g1231) & (!g107) & (!g1274)) + ((g1319) & (!sk[113]) & (g1231) & (!g107) & (g1274)) + ((g1319) & (!sk[113]) & (g1231) & (g107) & (!g1274)) + ((g1319) & (!sk[113]) & (g1231) & (g107) & (g1274)) + ((g1319) & (sk[113]) & (g1231) & (!g107) & (g1274)));
	assign g3835 = (((!g1319) & (!g1231) & (!sk[114]) & (!g867) & (g1274)) + ((!g1319) & (!g1231) & (!sk[114]) & (g867) & (g1274)) + ((!g1319) & (!g1231) & (sk[114]) & (g867) & (!g1274)) + ((!g1319) & (!g1231) & (sk[114]) & (g867) & (g1274)) + ((!g1319) & (g1231) & (!sk[114]) & (!g867) & (!g1274)) + ((!g1319) & (g1231) & (!sk[114]) & (!g867) & (g1274)) + ((!g1319) & (g1231) & (!sk[114]) & (g867) & (!g1274)) + ((!g1319) & (g1231) & (!sk[114]) & (g867) & (g1274)) + ((!g1319) & (g1231) & (sk[114]) & (g867) & (!g1274)) + ((!g1319) & (g1231) & (sk[114]) & (g867) & (g1274)) + ((g1319) & (!g1231) & (!sk[114]) & (!g867) & (!g1274)) + ((g1319) & (!g1231) & (!sk[114]) & (!g867) & (g1274)) + ((g1319) & (!g1231) & (!sk[114]) & (g867) & (!g1274)) + ((g1319) & (!g1231) & (!sk[114]) & (g867) & (g1274)) + ((g1319) & (g1231) & (!sk[114]) & (!g867) & (!g1274)) + ((g1319) & (g1231) & (!sk[114]) & (!g867) & (g1274)) + ((g1319) & (g1231) & (!sk[114]) & (g867) & (!g1274)) + ((g1319) & (g1231) & (!sk[114]) & (g867) & (g1274)) + ((g1319) & (g1231) & (sk[114]) & (!g867) & (g1274)));
	assign g3836 = (((!sk[115]) & (!g3837) & (g3838)) + ((!sk[115]) & (g3837) & (g3838)) + ((sk[115]) & (!g3837) & (!g3838)));
	assign g3837 = (((!g1004) & (!sk[116]) & (g3839)) + ((!g1004) & (sk[116]) & (g3839)) + ((g1004) & (!sk[116]) & (g3839)));
	assign g3838 = (((!sk[117]) & (!g1004) & (g3842)) + ((!sk[117]) & (g1004) & (g3842)) + ((sk[117]) & (g1004) & (g3842)));
	assign g3839 = (((!g3840) & (!sk[118]) & (g3841)) + ((!g3840) & (sk[118]) & (!g3841)) + ((g3840) & (!sk[118]) & (g3841)));
	assign g3840 = (((!g679) & (!sk[119]) & (g3845)) + ((!g679) & (sk[119]) & (g3845)) + ((g679) & (!sk[119]) & (g3845)));
	assign g3841 = (((!sk[120]) & (!g679) & (g3846)) + ((!sk[120]) & (g679) & (g3846)) + ((sk[120]) & (g679) & (g3846)));
	assign g3842 = (((!sk[121]) & (!g3843) & (g3844)) + ((!sk[121]) & (g3843) & (g3844)) + ((sk[121]) & (!g3843) & (!g3844)));
	assign g3843 = (((!sk[122]) & (!g679) & (g3847)) + ((!sk[122]) & (g679) & (g3847)) + ((sk[122]) & (!g679) & (g3847)));
	assign g3844 = (((!g679) & (!sk[123]) & (g3848)) + ((g679) & (!sk[123]) & (g3848)) + ((g679) & (sk[123]) & (g3848)));
	assign g3845 = (((!g1094) & (!g1006) & (!g107) & (!sk[124]) & (g1049)) + ((!g1094) & (!g1006) & (g107) & (!sk[124]) & (g1049)) + ((!g1094) & (!g1006) & (g107) & (sk[124]) & (g1049)) + ((!g1094) & (g1006) & (!g107) & (!sk[124]) & (!g1049)) + ((!g1094) & (g1006) & (!g107) & (!sk[124]) & (g1049)) + ((!g1094) & (g1006) & (g107) & (!sk[124]) & (!g1049)) + ((!g1094) & (g1006) & (g107) & (!sk[124]) & (g1049)) + ((!g1094) & (g1006) & (g107) & (sk[124]) & (!g1049)) + ((!g1094) & (g1006) & (g107) & (sk[124]) & (g1049)) + ((g1094) & (!g1006) & (!g107) & (!sk[124]) & (!g1049)) + ((g1094) & (!g1006) & (!g107) & (!sk[124]) & (g1049)) + ((g1094) & (!g1006) & (g107) & (!sk[124]) & (!g1049)) + ((g1094) & (!g1006) & (g107) & (!sk[124]) & (g1049)) + ((g1094) & (g1006) & (!g107) & (!sk[124]) & (!g1049)) + ((g1094) & (g1006) & (!g107) & (!sk[124]) & (g1049)) + ((g1094) & (g1006) & (g107) & (!sk[124]) & (!g1049)) + ((g1094) & (g1006) & (g107) & (!sk[124]) & (g1049)));
	assign g3846 = (((!g1094) & (!g1006) & (!sk[125]) & (!g867) & (g1049)) + ((!g1094) & (!g1006) & (!sk[125]) & (g867) & (g1049)) + ((!g1094) & (!g1006) & (sk[125]) & (g867) & (g1049)) + ((!g1094) & (g1006) & (!sk[125]) & (!g867) & (!g1049)) + ((!g1094) & (g1006) & (!sk[125]) & (!g867) & (g1049)) + ((!g1094) & (g1006) & (!sk[125]) & (g867) & (!g1049)) + ((!g1094) & (g1006) & (!sk[125]) & (g867) & (g1049)) + ((!g1094) & (g1006) & (sk[125]) & (g867) & (!g1049)) + ((!g1094) & (g1006) & (sk[125]) & (g867) & (g1049)) + ((g1094) & (!g1006) & (!sk[125]) & (!g867) & (!g1049)) + ((g1094) & (!g1006) & (!sk[125]) & (!g867) & (g1049)) + ((g1094) & (!g1006) & (!sk[125]) & (g867) & (!g1049)) + ((g1094) & (!g1006) & (!sk[125]) & (g867) & (g1049)) + ((g1094) & (g1006) & (!sk[125]) & (!g867) & (!g1049)) + ((g1094) & (g1006) & (!sk[125]) & (!g867) & (g1049)) + ((g1094) & (g1006) & (!sk[125]) & (g867) & (!g1049)) + ((g1094) & (g1006) & (!sk[125]) & (g867) & (g1049)));
	assign g3847 = (((!g1094) & (!g1006) & (!g107) & (!sk[126]) & (g1049)) + ((!g1094) & (!g1006) & (g107) & (!sk[126]) & (g1049)) + ((!g1094) & (!g1006) & (g107) & (sk[126]) & (!g1049)) + ((!g1094) & (!g1006) & (g107) & (sk[126]) & (g1049)) + ((!g1094) & (g1006) & (!g107) & (!sk[126]) & (!g1049)) + ((!g1094) & (g1006) & (!g107) & (!sk[126]) & (g1049)) + ((!g1094) & (g1006) & (g107) & (!sk[126]) & (!g1049)) + ((!g1094) & (g1006) & (g107) & (!sk[126]) & (g1049)) + ((!g1094) & (g1006) & (g107) & (sk[126]) & (!g1049)) + ((!g1094) & (g1006) & (g107) & (sk[126]) & (g1049)) + ((g1094) & (!g1006) & (!g107) & (!sk[126]) & (!g1049)) + ((g1094) & (!g1006) & (!g107) & (!sk[126]) & (g1049)) + ((g1094) & (!g1006) & (g107) & (!sk[126]) & (!g1049)) + ((g1094) & (!g1006) & (g107) & (!sk[126]) & (g1049)) + ((g1094) & (g1006) & (!g107) & (!sk[126]) & (!g1049)) + ((g1094) & (g1006) & (!g107) & (!sk[126]) & (g1049)) + ((g1094) & (g1006) & (!g107) & (sk[126]) & (g1049)) + ((g1094) & (g1006) & (g107) & (!sk[126]) & (!g1049)) + ((g1094) & (g1006) & (g107) & (!sk[126]) & (g1049)));
	assign g3848 = (((!g1094) & (!sk[127]) & (!g1006) & (!g867) & (g1049)) + ((!g1094) & (!sk[127]) & (!g1006) & (g867) & (g1049)) + ((!g1094) & (!sk[127]) & (g1006) & (!g867) & (!g1049)) + ((!g1094) & (!sk[127]) & (g1006) & (!g867) & (g1049)) + ((!g1094) & (!sk[127]) & (g1006) & (g867) & (!g1049)) + ((!g1094) & (!sk[127]) & (g1006) & (g867) & (g1049)) + ((!g1094) & (sk[127]) & (!g1006) & (g867) & (!g1049)) + ((!g1094) & (sk[127]) & (!g1006) & (g867) & (g1049)) + ((!g1094) & (sk[127]) & (g1006) & (g867) & (!g1049)) + ((!g1094) & (sk[127]) & (g1006) & (g867) & (g1049)) + ((g1094) & (!sk[127]) & (!g1006) & (!g867) & (!g1049)) + ((g1094) & (!sk[127]) & (!g1006) & (!g867) & (g1049)) + ((g1094) & (!sk[127]) & (!g1006) & (g867) & (!g1049)) + ((g1094) & (!sk[127]) & (!g1006) & (g867) & (g1049)) + ((g1094) & (!sk[127]) & (g1006) & (!g867) & (!g1049)) + ((g1094) & (!sk[127]) & (g1006) & (!g867) & (g1049)) + ((g1094) & (!sk[127]) & (g1006) & (g867) & (!g1049)) + ((g1094) & (!sk[127]) & (g1006) & (g867) & (g1049)) + ((g1094) & (sk[127]) & (g1006) & (!g867) & (g1049)));
	assign g3849 = (((!g3850) & (!sk[0]) & (g3851)) + ((!g3850) & (sk[0]) & (!g3851)) + ((g3850) & (!sk[0]) & (g3851)));
	assign g3850 = (((!g586) & (!sk[1]) & (g3852)) + ((!g586) & (sk[1]) & (g3852)) + ((g586) & (!sk[1]) & (g3852)));
	assign g3851 = (((!g586) & (!sk[2]) & (g3855)) + ((g586) & (!sk[2]) & (g3855)) + ((g586) & (sk[2]) & (g3855)));
	assign g3852 = (((!sk[3]) & (!g3853) & (g3854)) + ((!sk[3]) & (g3853) & (g3854)) + ((sk[3]) & (!g3853) & (!g3854)));
	assign g3853 = (((!sk[4]) & (!g126) & (g587)) + ((!sk[4]) & (g126) & (g587)) + ((sk[4]) & (!g126) & (g587)));
	assign g3854 = (((!sk[5]) & (!g126) & (g3858)) + ((!sk[5]) & (g126) & (g3858)) + ((sk[5]) & (g126) & (g3858)));
	assign g3855 = (((!g3856) & (!sk[6]) & (g3857)) + ((!g3856) & (sk[6]) & (!g3857)) + ((g3856) & (!sk[6]) & (g3857)));
	assign g3856 = (((!g126) & (!sk[7]) & (g587)) + ((!g126) & (sk[7]) & (g587)) + ((g126) & (!sk[7]) & (g587)));
	assign g3857 = (((!g126) & (!sk[8]) & (g3859)) + ((g126) & (!sk[8]) & (g3859)) + ((g126) & (sk[8]) & (g3859)));
	assign g3858 = (((!g542) & (!g91) & (!g584) & (!sk[9]) & (g629)) + ((!g542) & (!g91) & (!g584) & (sk[9]) & (g629)) + ((!g542) & (!g91) & (g584) & (!sk[9]) & (g629)) + ((!g542) & (!g91) & (g584) & (sk[9]) & (g629)) + ((!g542) & (g91) & (!g584) & (!sk[9]) & (!g629)) + ((!g542) & (g91) & (!g584) & (!sk[9]) & (g629)) + ((!g542) & (g91) & (!g584) & (sk[9]) & (g629)) + ((!g542) & (g91) & (g584) & (!sk[9]) & (!g629)) + ((!g542) & (g91) & (g584) & (!sk[9]) & (g629)) + ((!g542) & (g91) & (g584) & (sk[9]) & (!g629)) + ((g542) & (!g91) & (!g584) & (!sk[9]) & (!g629)) + ((g542) & (!g91) & (!g584) & (!sk[9]) & (g629)) + ((g542) & (!g91) & (!g584) & (sk[9]) & (g629)) + ((g542) & (!g91) & (g584) & (!sk[9]) & (!g629)) + ((g542) & (!g91) & (g584) & (!sk[9]) & (g629)) + ((g542) & (!g91) & (g584) & (sk[9]) & (!g629)) + ((g542) & (g91) & (!g584) & (!sk[9]) & (!g629)) + ((g542) & (g91) & (!g584) & (!sk[9]) & (g629)) + ((g542) & (g91) & (!g584) & (sk[9]) & (!g629)) + ((g542) & (g91) & (g584) & (!sk[9]) & (!g629)) + ((g542) & (g91) & (g584) & (!sk[9]) & (g629)) + ((g542) & (g91) & (g584) & (sk[9]) & (!g629)));
	assign g3859 = (((!g542) & (!g91) & (!sk[10]) & (!g584) & (g629)) + ((!g542) & (!g91) & (!sk[10]) & (g584) & (g629)) + ((!g542) & (!g91) & (sk[10]) & (!g584) & (!g629)) + ((!g542) & (!g91) & (sk[10]) & (g584) & (!g629)) + ((!g542) & (g91) & (!sk[10]) & (!g584) & (!g629)) + ((!g542) & (g91) & (!sk[10]) & (!g584) & (g629)) + ((!g542) & (g91) & (!sk[10]) & (g584) & (!g629)) + ((!g542) & (g91) & (!sk[10]) & (g584) & (g629)) + ((!g542) & (g91) & (sk[10]) & (!g584) & (!g629)) + ((!g542) & (g91) & (sk[10]) & (g584) & (g629)) + ((g542) & (!g91) & (!sk[10]) & (!g584) & (!g629)) + ((g542) & (!g91) & (!sk[10]) & (!g584) & (g629)) + ((g542) & (!g91) & (!sk[10]) & (g584) & (!g629)) + ((g542) & (!g91) & (!sk[10]) & (g584) & (g629)) + ((g542) & (!g91) & (sk[10]) & (!g584) & (!g629)) + ((g542) & (!g91) & (sk[10]) & (g584) & (g629)) + ((g542) & (g91) & (!sk[10]) & (!g584) & (!g629)) + ((g542) & (g91) & (!sk[10]) & (!g584) & (g629)) + ((g542) & (g91) & (!sk[10]) & (g584) & (!g629)) + ((g542) & (g91) & (!sk[10]) & (g584) & (g629)) + ((g542) & (g91) & (sk[10]) & (!g584) & (g629)) + ((g542) & (g91) & (sk[10]) & (g584) & (g629)));
	assign g3860 = (((!g3861) & (!sk[11]) & (g3862)) + ((!g3861) & (sk[11]) & (!g3862)) + ((g3861) & (!sk[11]) & (g3862)));
	assign g3861 = (((!g495) & (!sk[12]) & (g3863)) + ((!g495) & (sk[12]) & (g3863)) + ((g495) & (!sk[12]) & (g3863)));
	assign g3862 = (((!sk[13]) & (!g495) & (g3866)) + ((!sk[13]) & (g495) & (g3866)) + ((sk[13]) & (g495) & (g3866)));
	assign g3863 = (((!sk[14]) & (!g3864) & (g3865)) + ((!sk[14]) & (g3864) & (g3865)) + ((sk[14]) & (!g3864) & (!g3865)));
	assign g3864 = (((!g126) & (!sk[15]) & (g453)) + ((!g126) & (sk[15]) & (g453)) + ((g126) & (!sk[15]) & (g453)));
	assign g3865 = (((!g126) & (!sk[16]) & (g3869)) + ((g126) & (!sk[16]) & (g3869)) + ((g126) & (sk[16]) & (g3869)));
	assign g3866 = (((!g3867) & (!sk[17]) & (g3868)) + ((!g3867) & (sk[17]) & (!g3868)) + ((g3867) & (!sk[17]) & (g3868)));
	assign g3867 = (((!g126) & (!sk[18]) & (g453)) + ((!g126) & (sk[18]) & (g453)) + ((g126) & (!sk[18]) & (g453)));
	assign g3868 = (((!g126) & (!sk[19]) & (g3870)) + ((g126) & (!sk[19]) & (g3870)) + ((g126) & (sk[19]) & (g3870)));
	assign g3869 = (((!sk[20]) & (!g451) & (!g409) & (!g85) & (g86)) + ((!sk[20]) & (!g451) & (!g409) & (g85) & (g86)) + ((!sk[20]) & (!g451) & (g409) & (!g85) & (!g86)) + ((!sk[20]) & (!g451) & (g409) & (!g85) & (g86)) + ((!sk[20]) & (!g451) & (g409) & (g85) & (!g86)) + ((!sk[20]) & (!g451) & (g409) & (g85) & (g86)) + ((!sk[20]) & (g451) & (!g409) & (!g85) & (!g86)) + ((!sk[20]) & (g451) & (!g409) & (!g85) & (g86)) + ((!sk[20]) & (g451) & (!g409) & (g85) & (!g86)) + ((!sk[20]) & (g451) & (!g409) & (g85) & (g86)) + ((!sk[20]) & (g451) & (g409) & (!g85) & (!g86)) + ((!sk[20]) & (g451) & (g409) & (!g85) & (g86)) + ((!sk[20]) & (g451) & (g409) & (g85) & (!g86)) + ((!sk[20]) & (g451) & (g409) & (g85) & (g86)) + ((sk[20]) & (!g451) & (!g409) & (g85) & (!g86)) + ((sk[20]) & (!g451) & (!g409) & (g85) & (g86)) + ((sk[20]) & (!g451) & (g409) & (!g85) & (g86)) + ((sk[20]) & (!g451) & (g409) & (g85) & (!g86)) + ((sk[20]) & (g451) & (!g409) & (!g85) & (g86)) + ((sk[20]) & (g451) & (!g409) & (g85) & (!g86)) + ((sk[20]) & (g451) & (g409) & (!g85) & (!g86)) + ((sk[20]) & (g451) & (g409) & (!g85) & (g86)));
	assign g3870 = (((!g451) & (!sk[21]) & (!g409) & (!g85) & (g86)) + ((!g451) & (!sk[21]) & (!g409) & (g85) & (g86)) + ((!g451) & (!sk[21]) & (g409) & (!g85) & (!g86)) + ((!g451) & (!sk[21]) & (g409) & (!g85) & (g86)) + ((!g451) & (!sk[21]) & (g409) & (g85) & (!g86)) + ((!g451) & (!sk[21]) & (g409) & (g85) & (g86)) + ((!g451) & (sk[21]) & (!g409) & (!g85) & (!g86)) + ((!g451) & (sk[21]) & (!g409) & (!g85) & (g86)) + ((!g451) & (sk[21]) & (g409) & (!g85) & (!g86)) + ((!g451) & (sk[21]) & (g409) & (g85) & (g86)) + ((g451) & (!sk[21]) & (!g409) & (!g85) & (!g86)) + ((g451) & (!sk[21]) & (!g409) & (!g85) & (g86)) + ((g451) & (!sk[21]) & (!g409) & (g85) & (!g86)) + ((g451) & (!sk[21]) & (!g409) & (g85) & (g86)) + ((g451) & (!sk[21]) & (g409) & (!g85) & (!g86)) + ((g451) & (!sk[21]) & (g409) & (!g85) & (g86)) + ((g451) & (!sk[21]) & (g409) & (g85) & (!g86)) + ((g451) & (!sk[21]) & (g409) & (g85) & (g86)) + ((g451) & (sk[21]) & (!g409) & (!g85) & (!g86)) + ((g451) & (sk[21]) & (!g409) & (g85) & (g86)) + ((g451) & (sk[21]) & (g409) & (g85) & (!g86)) + ((g451) & (sk[21]) & (g409) & (g85) & (g86)));
	assign g3871 = (((!g3872) & (!sk[22]) & (g3873)) + ((!g3872) & (sk[22]) & (!g3873)) + ((g3872) & (!sk[22]) & (g3873)));
	assign g3872 = (((!sk[23]) & (!g364) & (g3874)) + ((!sk[23]) & (g364) & (g3874)) + ((sk[23]) & (!g364) & (g3874)));
	assign g3873 = (((!sk[24]) & (!g364) & (g3877)) + ((!sk[24]) & (g364) & (g3877)) + ((sk[24]) & (g364) & (g3877)));
	assign g3874 = (((!sk[25]) & (!g3875) & (g3876)) + ((!sk[25]) & (g3875) & (g3876)) + ((sk[25]) & (!g3875) & (!g3876)));
	assign g3875 = (((!g126) & (!sk[26]) & (g365)) + ((!g126) & (sk[26]) & (g365)) + ((g126) & (!sk[26]) & (g365)));
	assign g3876 = (((!sk[27]) & (!g126) & (g3880)) + ((!sk[27]) & (g126) & (g3880)) + ((sk[27]) & (g126) & (g3880)));
	assign g3877 = (((!sk[28]) & (!g3878) & (g3879)) + ((!sk[28]) & (g3878) & (g3879)) + ((sk[28]) & (!g3878) & (!g3879)));
	assign g3878 = (((!g126) & (!sk[29]) & (g365)) + ((!g126) & (sk[29]) & (g365)) + ((g126) & (!sk[29]) & (g365)));
	assign g3879 = (((!sk[30]) & (!g126) & (g3881)) + ((!sk[30]) & (g126) & (g3881)) + ((sk[30]) & (g126) & (g3881)));
	assign g3880 = (((!g320) & (!g318) & (!sk[31]) & (!g362) & (g407)) + ((!g320) & (!g318) & (!sk[31]) & (g362) & (g407)) + ((!g320) & (!g318) & (sk[31]) & (!g362) & (g407)) + ((!g320) & (!g318) & (sk[31]) & (g362) & (g407)) + ((!g320) & (g318) & (!sk[31]) & (!g362) & (!g407)) + ((!g320) & (g318) & (!sk[31]) & (!g362) & (g407)) + ((!g320) & (g318) & (!sk[31]) & (g362) & (!g407)) + ((!g320) & (g318) & (!sk[31]) & (g362) & (g407)) + ((!g320) & (g318) & (sk[31]) & (!g362) & (g407)) + ((!g320) & (g318) & (sk[31]) & (g362) & (!g407)) + ((g320) & (!g318) & (!sk[31]) & (!g362) & (!g407)) + ((g320) & (!g318) & (!sk[31]) & (!g362) & (g407)) + ((g320) & (!g318) & (!sk[31]) & (g362) & (!g407)) + ((g320) & (!g318) & (!sk[31]) & (g362) & (g407)) + ((g320) & (!g318) & (sk[31]) & (!g362) & (g407)) + ((g320) & (!g318) & (sk[31]) & (g362) & (!g407)) + ((g320) & (g318) & (!sk[31]) & (!g362) & (!g407)) + ((g320) & (g318) & (!sk[31]) & (!g362) & (g407)) + ((g320) & (g318) & (!sk[31]) & (g362) & (!g407)) + ((g320) & (g318) & (!sk[31]) & (g362) & (g407)) + ((g320) & (g318) & (sk[31]) & (!g362) & (!g407)) + ((g320) & (g318) & (sk[31]) & (g362) & (!g407)));
	assign g3881 = (((!g320) & (!sk[32]) & (!g318) & (!g362) & (g407)) + ((!g320) & (!sk[32]) & (!g318) & (g362) & (g407)) + ((!g320) & (!sk[32]) & (g318) & (!g362) & (!g407)) + ((!g320) & (!sk[32]) & (g318) & (!g362) & (g407)) + ((!g320) & (!sk[32]) & (g318) & (g362) & (!g407)) + ((!g320) & (!sk[32]) & (g318) & (g362) & (g407)) + ((!g320) & (sk[32]) & (!g318) & (!g362) & (!g407)) + ((!g320) & (sk[32]) & (!g318) & (g362) & (!g407)) + ((!g320) & (sk[32]) & (g318) & (!g362) & (!g407)) + ((!g320) & (sk[32]) & (g318) & (g362) & (g407)) + ((g320) & (!sk[32]) & (!g318) & (!g362) & (!g407)) + ((g320) & (!sk[32]) & (!g318) & (!g362) & (g407)) + ((g320) & (!sk[32]) & (!g318) & (g362) & (!g407)) + ((g320) & (!sk[32]) & (!g318) & (g362) & (g407)) + ((g320) & (!sk[32]) & (g318) & (!g362) & (!g407)) + ((g320) & (!sk[32]) & (g318) & (!g362) & (g407)) + ((g320) & (!sk[32]) & (g318) & (g362) & (!g407)) + ((g320) & (!sk[32]) & (g318) & (g362) & (g407)) + ((g320) & (sk[32]) & (!g318) & (!g362) & (!g407)) + ((g320) & (sk[32]) & (!g318) & (g362) & (g407)) + ((g320) & (sk[32]) & (g318) & (!g362) & (g407)) + ((g320) & (sk[32]) & (g318) & (g362) & (g407)));
	assign g3882 = (((!sk[33]) & (!g3883) & (g3884)) + ((!sk[33]) & (g3883) & (g3884)) + ((sk[33]) & (!g3883) & (!g3884)));
	assign g3883 = (((!g317) & (!sk[34]) & (g3885)) + ((!g317) & (sk[34]) & (g3885)) + ((g317) & (!sk[34]) & (g3885)));
	assign g3884 = (((!sk[35]) & (!g317) & (g3888)) + ((!sk[35]) & (g317) & (g3888)) + ((sk[35]) & (g317) & (g3888)));
	assign g3885 = (((!g3886) & (!sk[36]) & (g3887)) + ((!g3886) & (sk[36]) & (!g3887)) + ((g3886) & (!sk[36]) & (g3887)));
	assign g3886 = (((!sk[37]) & (!g126) & (g275)) + ((!sk[37]) & (g126) & (g275)) + ((sk[37]) & (!g126) & (g275)));
	assign g3887 = (((!sk[38]) & (!g126) & (g3891)) + ((!sk[38]) & (g126) & (g3891)) + ((sk[38]) & (g126) & (g3891)));
	assign g3888 = (((!sk[39]) & (!g3889) & (g3890)) + ((!sk[39]) & (g3889) & (g3890)) + ((sk[39]) & (!g3889) & (!g3890)));
	assign g3889 = (((!g126) & (!sk[40]) & (g275)) + ((!g126) & (sk[40]) & (g275)) + ((g126) & (!sk[40]) & (g275)));
	assign g3890 = (((!g126) & (!sk[41]) & (g3892)) + ((g126) & (!sk[41]) & (g3892)) + ((g126) & (sk[41]) & (g3892)));
	assign g3891 = (((!sk[42]) & (!g273) & (!g231) & (!g90) & (g87)) + ((!sk[42]) & (!g273) & (!g231) & (g90) & (g87)) + ((!sk[42]) & (!g273) & (g231) & (!g90) & (!g87)) + ((!sk[42]) & (!g273) & (g231) & (!g90) & (g87)) + ((!sk[42]) & (!g273) & (g231) & (g90) & (!g87)) + ((!sk[42]) & (!g273) & (g231) & (g90) & (g87)) + ((!sk[42]) & (g273) & (!g231) & (!g90) & (!g87)) + ((!sk[42]) & (g273) & (!g231) & (!g90) & (g87)) + ((!sk[42]) & (g273) & (!g231) & (g90) & (!g87)) + ((!sk[42]) & (g273) & (!g231) & (g90) & (g87)) + ((!sk[42]) & (g273) & (g231) & (!g90) & (!g87)) + ((!sk[42]) & (g273) & (g231) & (!g90) & (g87)) + ((!sk[42]) & (g273) & (g231) & (g90) & (!g87)) + ((!sk[42]) & (g273) & (g231) & (g90) & (g87)) + ((sk[42]) & (!g273) & (!g231) & (g90) & (!g87)) + ((sk[42]) & (!g273) & (!g231) & (g90) & (g87)) + ((sk[42]) & (!g273) & (g231) & (!g90) & (g87)) + ((sk[42]) & (!g273) & (g231) & (g90) & (!g87)) + ((sk[42]) & (g273) & (!g231) & (!g90) & (g87)) + ((sk[42]) & (g273) & (!g231) & (g90) & (!g87)) + ((sk[42]) & (g273) & (g231) & (!g90) & (!g87)) + ((sk[42]) & (g273) & (g231) & (!g90) & (g87)));
	assign g3892 = (((!g273) & (!g231) & (!g90) & (!sk[43]) & (g87)) + ((!g273) & (!g231) & (!g90) & (sk[43]) & (!g87)) + ((!g273) & (!g231) & (!g90) & (sk[43]) & (g87)) + ((!g273) & (!g231) & (g90) & (!sk[43]) & (g87)) + ((!g273) & (g231) & (!g90) & (!sk[43]) & (!g87)) + ((!g273) & (g231) & (!g90) & (!sk[43]) & (g87)) + ((!g273) & (g231) & (!g90) & (sk[43]) & (!g87)) + ((!g273) & (g231) & (g90) & (!sk[43]) & (!g87)) + ((!g273) & (g231) & (g90) & (!sk[43]) & (g87)) + ((!g273) & (g231) & (g90) & (sk[43]) & (g87)) + ((g273) & (!g231) & (!g90) & (!sk[43]) & (!g87)) + ((g273) & (!g231) & (!g90) & (!sk[43]) & (g87)) + ((g273) & (!g231) & (!g90) & (sk[43]) & (!g87)) + ((g273) & (!g231) & (g90) & (!sk[43]) & (!g87)) + ((g273) & (!g231) & (g90) & (!sk[43]) & (g87)) + ((g273) & (!g231) & (g90) & (sk[43]) & (g87)) + ((g273) & (g231) & (!g90) & (!sk[43]) & (!g87)) + ((g273) & (g231) & (!g90) & (!sk[43]) & (g87)) + ((g273) & (g231) & (g90) & (!sk[43]) & (!g87)) + ((g273) & (g231) & (g90) & (!sk[43]) & (g87)) + ((g273) & (g231) & (g90) & (sk[43]) & (!g87)) + ((g273) & (g231) & (g90) & (sk[43]) & (g87)));
	assign gnd = ();
	assign vcc = ();

endmodule