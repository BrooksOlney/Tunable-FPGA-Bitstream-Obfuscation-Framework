module ks_apex2_qmap_map (clk, sk, in, outreg);

	wire i_36_;
	wire i_34_;
	wire i_28_;
	wire i_29_;
	wire i_35_;
	wire i_27_;
	wire i_23_;
	wire i_24_;
	wire i_16_;
	wire i_13_;
	wire i_7_;
	wire i_8_;
	wire i_12_;
	wire i_6_;
	wire i_2_;
	wire i_4_;
	wire i_5_;
	wire i_9_;
	wire i_17_;
	wire i_11_;
	wire i_19_;
	wire i_3_;
	wire i_18_;
	wire i_14_;
	wire i_10_;
	wire i_32_;
	wire i_1_;
	wire i_31_;
	wire i_30_;
	wire i_21_;
	wire i_26_;
	wire i_25_;
	wire i_22_;
	wire i_33_;
	wire i_20_;
	wire i_0_;
	wire i_37_;
	wire i_38_;
	wire o_0_;
	wire o_1_;
	wire o_2_;

	
input [13:0] in;
reg [13:0] inreg;
input clk;
output reg [7:0] outreg;
wire [7:0] out;
	
always@(posedge clk)
begin
	inreg <= in;
	outreg <= out;
end


	input [127 : 0] sk /* synthesis noprune */;
	
	assign {i_36_, i_34_, i_28_, i_29_, i_35_, i_27_, i_23_, i_24_, i_16_, i_13_, i_7_, i_8_, i_12_, i_6_, i_2_, i_4_, i_5_, i_9_, i_17_, i_11_, i_19_, i_3_, i_18_, i_14_, i_10_, i_32_, i_1_, i_31_, i_30_, i_21_, i_26_, i_25_, i_22_, i_33_, i_20_, i_0_, i_37_, i_38_} =  inreg;
	assign out={o_0_, o_1_, o_2_};

	wire g427, g661, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19;
	wire g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40;
	wire g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57, g58, g59, g60, g61;
	wire g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g79, g80, g81, g82;
	wire g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101, g102, g103;
	wire g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124;
	wire g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145;
	wire g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166;
	wire g167, g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183, g712, g184, g185, g186;
	wire g187, g188, g189, g190, g191, g192, g193, g194, g195, g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207;
	wire g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219, g220, g702, g221, g222, g223, g224, g225, g226, g227;
	wire g228, g229, g230, g231, g232, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242, g243, g244, g245, g247, g248, g249;
	wire g250, g251, g252, g253, g254, g255, g256, g257, g258, g259, g260, g261, g262, g263, g264, g265, g266, g267, g268, g269, g270;
	wire g271, g272, g273, g274, g275, g276, g277, g278, g279, g280, g281, g282, g283, g284, g285, g286, g287, g288, g289, g290, g291;
	wire g292, g293, g294, g295, g296, g297, g298, g299, g300, g301, g302, g303, g304, g305, g306, g307, g308, g309, g310, g311, g312;
	wire g313, g314, g315, g316, g317, g318, g319, g320, g321, g322, g323, g324, g325, g326, g327, g328, g329, g330, g331, g332, g333;
	wire g334, g335, g336, g337, g338, g339, g340, g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351, g352, g353, g354;
	wire g355, g356, g357, g358, g359, g360, g361, g362, g363, g364, g365, g366, g367, g368, g369, g370, g371, g372, g373, g374, g375;
	wire g376, g377, g378, g379, g380, g381, g382, g383, g384, g385, g386, g387, g388, g389, g390, g391, g392, g393, g394, g395, g396;
	wire g397, g398, g399, g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410, g411, g412, g413, g414, g415, g416, g417;
	wire g418, g419, g420, g421, g422, g423, g424, g425, g426, g428, g429, g430, g431, g432, g433, g434, g435, g436, g437, g438, g439;
	wire g440, g441, g442, g443, g444, g445, g446, g447, g448, g449, g450, g451, g452, g453, g454, g455, g456, g457, g458, g459, g460;
	wire g461, g462, g463, g464, g465, g466, g467, g468, g469, g470, g471, g472, g473, g474, g475, g696, g476, g477, g478, g479, g480;
	wire g481, g482, g483, g484, g485, g486, g487, g488, g489, g490, g491, g492, g493, g494, g495, g496, g497, g498, g499, g500, g501;
	wire g502, g503, g504, g505, g506, g507, g508, g509, g510, g511, g512, g513, g514, g515, g516, g517, g518, g519, g520, g521, g522;
	wire g523, g524, g525, g526, g527, g528, g529, g530, g531, g532, g533, g534, g535, g536, g537, g538, g539, g540, g541, g542, g543;
	wire g544, g545, g546, g547, g548, g549, g550, g551, g552, g553, g554, g555, g556, g557, g558, g559, g560, g561, g562, g563, g564;
	wire g565, g566, g567, g568, g569, g570, g571, g572, g573, g574, g575, g576, g577, g578, g579, g580, g685, g581, g582, g583, g584;
	wire g585, g586, g587, g588, g589, g590, g591, g592, g593, g594, g595, g596, g597, g598, g599, g600, g601, g602, g603, g604, g605;
	wire g606, g607, g608, g609, g610, g611, g612, g613, g614, g615, g616, g617, g618, g619, g620, g621, g672, g622, g623, g624, g625;
	wire g626, g627, g628, g629, g630, g631, g632, g633, g634, g635, g636, g637, g638, g639, g640, g641, g642, g643, g644, g645, g646;
	wire g647, g648, g649, g662, g650, g651, g652, g653, g654, g655, g656, g657, g658, g659, g660, g663, g664, g665, g666, g669, g667;
	wire g668, g670, g671, g673, g674, g675, g678, g676, g677, g681, g682, g679, g680, g683, g684, g686, g687, g688, g691, g689, g690;
	wire g693, g694, g692, g695, g697, g698, g699, g700, g701, g703, g704, g705, g706, g709, g707, g708, g710, g711, g713, g714, g715;
	wire g716, g717, g718;

	assign o_1_ = (((sk[0]) & (!g427)));
	assign o_2_ = (((sk[1]) & (!g661)));
	assign g1 = (((i_28_) & (!sk[2]) & (i_29_)) + ((!i_28_) & (sk[2]) & (!i_29_)));
	assign g2 = (((!sk[3]) & (i_34_) & (i_35_)) + ((sk[3]) & (!i_34_) & (i_35_)));
	assign g3 = (((!sk[4]) & (!i_27_) & (i_28_) & (i_23_)) + ((sk[4]) & (!i_27_) & (!i_28_) & (!i_23_)));
	assign g4 = (((!sk[5]) & (g2) & (!g3) & (i_29_)) + ((sk[5]) & (g2) & (g3) & (!i_29_)));
	assign g5 = (((i_24_) & (sk[6]) & (!i_27_) & (!i_23_)) + ((!i_24_) & (sk[6]) & (i_27_) & (!i_23_)) + ((i_24_) & (!sk[6]) & (!i_27_) & (i_23_)) + ((!i_24_) & (sk[6]) & (!i_27_) & (i_23_)));
	assign g6 = (((!sk[7]) & (!i_34_) & (!g1) & (!g4) & (g5)) + ((!sk[7]) & (!i_34_) & (!g1) & (!g4) & (g5)) + ((!sk[7]) & (i_34_) & (!g1) & (g4) & (!g5)) + ((sk[7]) & (!i_34_) & (!g1) & (!g4) & (!g5)) + ((sk[7]) & (!i_34_) & (!g1) & (!g4) & (!g5)));
	assign g7 = (((!sk[8]) & (!i_7_) & (i_8_)) + ((sk[8]) & (!i_7_) & (!i_8_)));
	assign g8 = (((i_2_) & (!sk[9]) & (!i_4_) & (i_5_)) + ((!i_2_) & (sk[9]) & (!i_4_) & (!i_5_)));
	assign g9 = (((i_12_) & (!i_6_) & (!sk[10]) & (g8)) + ((!i_12_) & (!i_6_) & (sk[10]) & (g8)));
	assign g10 = (((!sk[11]) & (!i_2_) & (!i_9_) & (!i_6_) & (i_4_) & (!i_5_)) + ((!sk[11]) & (i_2_) & (!i_9_) & (!i_6_) & (!i_4_) & (i_5_)) + ((sk[11]) & (!i_2_) & (!i_9_) & (!i_6_) & (!i_4_) & (!i_5_)));
	assign g11 = (((g7) & (!sk[12]) & (g10)) + ((!g7) & (!sk[12]) & (g10)));
	assign g12 = (((!i_11_) & (!sk[13]) & (i_19_)) + ((!i_11_) & (sk[13]) & (!i_19_)));
	assign g13 = (((!sk[14]) & (!i_17_) & (g12)) + ((!sk[14]) & (!i_17_) & (g12)));
	assign g14 = (((i_6_) & (!i_4_) & (!sk[15]) & (i_5_)) + ((!i_6_) & (!i_4_) & (sk[15]) & (!i_5_)));
	assign g15 = (((i_17_) & (!i_9_) & (!sk[16]) & (i_18_)) + ((!i_17_) & (!i_9_) & (sk[16]) & (!i_18_)));
	assign g16 = (((!sk[17]) & (!i_2_) & (!i_7_) & (!i_3_) & (g14) & (!g15)) + ((!sk[17]) & (i_2_) & (!i_7_) & (!i_3_) & (!g14) & (g15)) + ((!sk[17]) & (!i_2_) & (!i_7_) & (i_3_) & (g14) & (g15)));
	assign g17 = (((!i_16_) & (!i_8_) & (!sk[18]) & (!g11) & (g13) & (!g16)) + ((!i_16_) & (!i_8_) & (!sk[18]) & (g11) & (g13) & (!g16)) + ((i_16_) & (!i_8_) & (!sk[18]) & (!g11) & (!g13) & (g16)) + ((!i_16_) & (!i_8_) & (sk[18]) & (!g11) & (!g13) & (g16)));
	assign g18 = (((!i_16_) & (!i_13_) & (!g7) & (!sk[19]) & (g9) & (!g17)) + ((!i_16_) & (!i_13_) & (!g7) & (sk[19]) & (!g9) & (g17)) + ((i_16_) & (!i_13_) & (!g7) & (!sk[19]) & (!g9) & (g17)) + ((!i_16_) & (!i_13_) & (g7) & (!sk[19]) & (g9) & (!g17)));
	assign g19 = (((!sk[20]) & (!i_27_) & (i_28_)) + ((sk[20]) & (!i_27_) & (!i_28_)));
	assign g20 = (((!sk[21]) & (!i_24_) & (g19)) + ((!sk[21]) & (!i_24_) & (g19)));
	assign g21 = (((!sk[22]) & (!g20) & (i_29_)) + ((sk[22]) & (g20) & (!i_29_)));
	assign g22 = (((!sk[23]) & (!i_13_) & (i_14_)) + ((!sk[23]) & (i_13_) & (i_14_)));
	assign g23 = (((i_16_) & (!i_17_) & (!sk[24]) & (i_23_)) + ((!i_16_) & (!i_17_) & (sk[24]) & (!i_23_)));
	assign g24 = (((!i_13_) & (!sk[25]) & (i_10_)) + ((!i_13_) & (!sk[25]) & (i_10_)));
	assign g25 = (((!sk[26]) & (!g11) & (g24)) + ((sk[26]) & (g11) & (!g24)));
	assign g26 = (((g22) & (!g23) & (!sk[27]) & (g25)) + ((!g22) & (g23) & (sk[27]) & (g25)));
	assign g27 = (((!i_16_) & (!sk[28]) & (!i_13_) & (!i_14_) & (i_10_)) + ((i_16_) & (!sk[28]) & (!i_13_) & (i_14_) & (!i_10_)) + ((!i_16_) & (sk[28]) & (!i_13_) & (!i_14_) & (!i_10_)) + ((!i_16_) & (sk[28]) & (i_13_) & (!i_14_) & (!i_10_)));
	assign g28 = (((sk[29]) & (!i_16_) & (!i_13_) & (!i_14_)) + ((!sk[29]) & (i_16_) & (!i_13_) & (i_14_)) + ((sk[29]) & (!i_16_) & (!i_13_) & (!i_14_)));
	assign g29 = (((i_2_) & (!g14) & (!sk[30]) & (i_1_)) + ((!i_2_) & (g14) & (sk[30]) & (!i_1_)));
	assign g30 = (((!g28) & (!i_7_) & (!i_8_) & (!sk[31]) & (g29)) + ((g28) & (!i_7_) & (i_8_) & (!sk[31]) & (!g29)) + ((g28) & (!i_7_) & (!i_8_) & (!sk[31]) & (g29)));
	assign g31 = (((i_7_) & (!sk[32]) & (!i_9_) & (i_6_)) + ((!i_7_) & (sk[32]) & (!i_9_) & (!i_6_)));
	assign g32 = (((g8) & (!sk[33]) & (g31)) + ((!g8) & (!sk[33]) & (g31)));
	assign g33 = (((!i_24_) & (!sk[34]) & (i_23_)) + ((!i_24_) & (sk[34]) & (!i_23_)));
	assign g34 = (((i_27_) & (!sk[35]) & (!i_28_) & (i_29_)) + ((!i_27_) & (sk[35]) & (!i_28_) & (!i_29_)));
	assign g35 = (((i_17_) & (!g33) & (!sk[36]) & (g34)) + ((!i_17_) & (g33) & (sk[36]) & (g34)));
	assign g36 = (((!i_32_) & (!g27) & (!sk[37]) & (!g30) & (g32) & (!g35)) + ((i_32_) & (!g27) & (!sk[37]) & (!g30) & (!g32) & (g35)) + ((!i_32_) & (!g27) & (sk[37]) & (g30) & (!g32) & (g35)) + ((!i_32_) & (g27) & (!sk[37]) & (!g30) & (g32) & (g35)));
	assign g37 = (((!sk[38]) & (!i_32_) & (g1)) + ((!sk[38]) & (!i_32_) & (g1)));
	assign g38 = (((i_27_) & (!i_17_) & (!sk[39]) & (i_23_)) + ((!i_27_) & (!i_17_) & (sk[39]) & (!i_23_)));
	assign g39 = (((!g37) & (!g27) & (!sk[40]) & (!g32) & (g38)) + ((g37) & (!g27) & (!sk[40]) & (g32) & (!g38)) + ((g37) & (g27) & (!sk[40]) & (g32) & (g38)));
	assign g40 = (((!i_34_) & (!i_35_) & (!g34) & (!sk[41]) & (g26) & (!g39)) + ((!i_34_) & (!i_35_) & (!g34) & (sk[41]) & (!g26) & (!g39)) + ((i_34_) & (!i_35_) & (!g34) & (!sk[41]) & (!g26) & (g39)) + ((!i_34_) & (!i_35_) & (!g34) & (sk[41]) & (!g26) & (!g39)) + ((!i_34_) & (!i_35_) & (!g34) & (!sk[41]) & (g26) & (!g39)));
	assign g41 = (((!sk[42]) & (!i_17_) & (!g28) & (!i_7_) & (g29)) + ((!sk[42]) & (i_17_) & (!g28) & (i_7_) & (!g29)) + ((!sk[42]) & (!i_17_) & (g28) & (!i_7_) & (g29)));
	assign g42 = (((!g5) & (!sk[43]) & (g37)) + ((!g5) & (!sk[43]) & (g37)));
	assign g43 = (((!sk[44]) & (i_34_) & (!g41) & (g42)) + ((sk[44]) & (i_34_) & (!g41) & (!g42)) + ((!sk[44]) & (i_34_) & (!g41) & (g42)));
	assign g44 = (((!sk[45]) & (!g21) & (!g26) & (!g36) & (g40) & (!g43)) + ((sk[45]) & (!g21) & (!g26) & (g36) & (!g40) & (!g43)) + ((!sk[45]) & (g21) & (!g26) & (!g36) & (!g40) & (g43)) + ((sk[45]) & (!g21) & (!g26) & (!g36) & (!g40) & (!g43)) + ((!sk[45]) & (g21) & (g26) & (!g36) & (!g40) & (g43)));
	assign g45 = (((!i_16_) & (!sk[46]) & (i_13_)) + ((!i_16_) & (sk[46]) & (!i_13_)));
	assign g46 = (((!i_2_) & (!sk[47]) & (i_8_)) + ((!i_2_) & (sk[47]) & (!i_8_)));
	assign g47 = (((!i_3_) & (!g14) & (!sk[48]) & (!g15) & (g46)) + ((i_3_) & (!g14) & (!sk[48]) & (g15) & (!g46)) + ((i_3_) & (g14) & (!sk[48]) & (g15) & (g46)));
	assign g48 = (((i_9_) & (!sk[49]) & (!i_6_) & (i_8_)) + ((!i_9_) & (sk[49]) & (!i_6_) & (!i_8_)));
	assign g49 = (((g8) & (!sk[50]) & (g48)) + ((!g8) & (!sk[50]) & (g48)));
	assign g50 = (((!i_23_) & (!g45) & (!g13) & (g47) & (!sk[51]) & (!g49)) + ((!i_23_) & (g45) & (!g13) & (g47) & (!sk[51]) & (!g49)) + ((i_23_) & (!g45) & (!g13) & (!g47) & (!sk[51]) & (g49)) + ((!i_23_) & (g45) & (g13) & (!g47) & (sk[51]) & (g49)));
	assign g51 = (((!sk[52]) & (!i_8_) & (g9)) + ((!sk[52]) & (!i_8_) & (g9)));
	assign g52 = (((!i_23_) & (!sk[53]) & (!g28) & (!i_31_) & (g50) & (!g51)) + ((!i_23_) & (sk[53]) & (!g28) & (!i_31_) & (!g50) & (!g51)) + ((!i_23_) & (sk[53]) & (!g28) & (i_31_) & (!g50) & (!g51)) + ((!i_23_) & (sk[53]) & (!g28) & (!i_31_) & (!g50) & (!g51)) + ((i_23_) & (!sk[53]) & (!g28) & (!i_31_) & (!g50) & (g51)));
	assign g53 = (((!i_17_) & (!sk[54]) & (g45)) + ((!i_17_) & (!sk[54]) & (g45)));
	assign g54 = (((!i_16_) & (!sk[55]) & (i_14_)) + ((!i_16_) & (sk[55]) & (!i_14_)));
	assign g55 = (((!sk[56]) & (!i_17_) & (g54)) + ((!sk[56]) & (!i_17_) & (g54)));
	assign g56 = (((!i_13_) & (!g53) & (!sk[57]) & (!g10) & (i_10_) & (!g55)) + ((i_13_) & (!g53) & (!sk[57]) & (!g10) & (!i_10_) & (g55)) + ((i_13_) & (!g53) & (!sk[57]) & (g10) & (!i_10_) & (g55)) + ((!i_13_) & (g53) & (sk[57]) & (g10) & (!i_10_) & (!g55)));
	assign g57 = (((!i_32_) & (!sk[58]) & (i_31_)) + ((!i_32_) & (sk[58]) & (!i_31_)));
	assign g58 = (((g29) & (!sk[59]) & (g23)) + ((!g29) & (!sk[59]) & (g23)));
	assign g59 = (((!sk[60]) & (!g20) & (!g22) & (!g57) & (i_29_) & (!g58)) + ((!sk[60]) & (g20) & (!g22) & (!g57) & (!i_29_) & (g58)) + ((!sk[60]) & (g20) & (!g22) & (g57) & (!i_29_) & (g58)));
	assign g60 = (((!i_31_) & (!sk[61]) & (g1)) + ((!i_31_) & (!sk[61]) & (g1)));
	assign g61 = (((!i_17_) & (!g28) & (!sk[62]) & (!i_8_) & (g29)) + ((i_17_) & (!g28) & (!sk[62]) & (i_8_) & (!g29)) + ((!i_17_) & (g28) & (!sk[62]) & (!i_8_) & (g29)));
	assign g62 = (((!g5) & (!g27) & (g60) & (g61) & (!g49) & (!g35)) + ((!g5) & (g27) & (!g60) & (!g61) & (g49) & (g35)));
	assign g63 = (((!g42) & (!g56) & (!sk[64]) & (!g59) & (g62)) + ((g42) & (!g56) & (!sk[64]) & (g59) & (!g62)) + ((!g42) & (!g56) & (sk[64]) & (!g59) & (!g62)) + ((!g42) & (!g56) & (sk[64]) & (!g59) & (!g62)));
	assign g64 = (((!i_34_) & (!i_35_) & (!sk[65]) & (!g52) & (g21) & (!g63)) + ((i_34_) & (!i_35_) & (!sk[65]) & (!g52) & (!g21) & (g63)) + ((i_34_) & (!i_35_) & (!sk[65]) & (!g52) & (g21) & (!g63)) + ((i_34_) & (!i_35_) & (sk[65]) & (!g52) & (!g21) & (!g63)));
	assign g65 = (((!i_35_) & (!sk[66]) & (i_32_)) + ((!i_35_) & (sk[66]) & (!i_32_)));
	assign g66 = (((i_34_) & (!sk[67]) & (g65)) + ((!i_34_) & (!sk[67]) & (g65)));
	assign g67 = (((!sk[68]) & (!i_2_) & (!i_9_) & (!i_3_) & (g14)) + ((!sk[68]) & (i_2_) & (!i_9_) & (i_3_) & (!g14)) + ((!sk[68]) & (!i_2_) & (!i_9_) & (i_3_) & (g14)));
	assign g68 = (((g33) & (!i_18_) & (!i_11_) & (!i_19_) & (g67) & (!g10)) + ((g33) & (!i_18_) & (!i_11_) & (!i_19_) & (!g67) & (g10)));
	assign g69 = (((!sk[70]) & (!g53) & (g68)) + ((!sk[70]) & (g53) & (g68)));
	assign g70 = (((!i_30_) & (!sk[71]) & (i_32_)) + ((i_30_) & (sk[71]) & (!i_32_)));
	assign g71 = (((!sk[72]) & (!i_24_) & (i_26_)) + ((sk[72]) & (i_24_) & (!i_26_)));
	assign g72 = (((!i_27_) & (!sk[73]) & (!i_23_) & (!i_21_) & (g71)) + ((i_27_) & (!sk[73]) & (!i_23_) & (i_21_) & (!g71)) + ((!i_27_) & (sk[73]) & (!i_23_) & (!i_21_) & (!g71)));
	assign g73 = (((i_12_) & (!g22) & (!sk[74]) & (i_7_)) + ((!i_12_) & (!g22) & (sk[74]) & (!i_7_)));
	assign g74 = (((i_16_) & (!sk[75]) & (!g72) & (g73)) + ((!i_16_) & (sk[75]) & (g72) & (g73)));
	assign g75 = (((!sk[76]) & (i_28_) & (!g70) & (g74)) + ((sk[76]) & (!i_28_) & (!g70) & (g74)));
	assign g76 = (((!i_24_) & (!i_34_) & (!sk[77]) & (!i_35_) & (i_32_) & (!g34)) + ((i_24_) & (!i_34_) & (!sk[77]) & (!i_35_) & (!i_32_) & (g34)) + ((!i_24_) & (i_34_) & (sk[77]) & (!i_35_) & (!i_32_) & (g34)) + ((!i_24_) & (!i_34_) & (sk[77]) & (i_35_) & (!i_32_) & (g34)));
	assign g77 = (((!i_7_) & (!sk[78]) & (g9)) + ((!i_7_) & (!sk[78]) & (g9)));
	assign g78 = (((g13) & (!sk[79]) & (g32)) + ((!g13) & (!sk[79]) & (g32)));
	assign g79 = (((!i_23_) & (!g45) & (!g77) & (g16) & (!sk[80]) & (!g78)) + ((!i_23_) & (g45) & (!g77) & (g16) & (!sk[80]) & (!g78)) + ((i_23_) & (!g45) & (!g77) & (!g16) & (!sk[80]) & (g78)) + ((!i_23_) & (g45) & (g77) & (!g16) & (sk[80]) & (!g78)) + ((!i_23_) & (g45) & (!g77) & (!g16) & (sk[80]) & (g78)));
	assign g80 = (((!g66) & (!g34) & (!g69) & (!g75) & (!g76) & (!g79)) + ((!g66) & (!g34) & (!g69) & (!g75) & (!g76) & (!g79)) + ((!g66) & (!g34) & (!g69) & (!g75) & (!g76) & (!g79)) + ((!g66) & (!g34) & (!g69) & (!g75) & (!g76) & (!g79)) + ((!g66) & (!g34) & (!g69) & (!g75) & (!g76) & (!g79)) + ((!g66) & (!g34) & (!g69) & (!g75) & (!g76) & (!g79)));
	assign g81 = (((!i_28_) & (!i_17_) & (!g72) & (!sk[82]) & (g30)) + ((i_28_) & (!i_17_) & (g72) & (!sk[82]) & (!g30)) + ((!i_28_) & (!i_17_) & (g72) & (!sk[82]) & (g30)));
	assign g82 = (((i_28_) & (!sk[83]) & (!g2) & (i_29_)) + ((!i_28_) & (sk[83]) & (g2) & (!i_29_)));
	assign g83 = (((g30) & (!sk[84]) & (!g38) & (g82)) + ((g30) & (!sk[84]) & (g38) & (g82)));
	assign g84 = (((!sk[85]) & (i_28_) & (!i_30_) & (i_29_)) + ((sk[85]) & (!i_28_) & (!i_30_) & (!i_29_)));
	assign g85 = (((!i_34_) & (!g57) & (!g33) & (!sk[86]) & (g84)) + ((i_34_) & (!g57) & (g33) & (!sk[86]) & (!g84)) + ((i_34_) & (g57) & (g33) & (!sk[86]) & (g84)));
	assign g86 = (((!sk[87]) & (!i_31_) & (g70)) + ((sk[87]) & (i_31_) & (!g70)));
	assign g87 = (((!sk[88]) & (!i_7_) & (!g85) & (!g82) & (g86)) + ((sk[88]) & (!i_7_) & (g85) & (!g82) & (!g86)) + ((!sk[88]) & (i_7_) & (!g85) & (g82) & (!g86)) + ((sk[88]) & (!i_7_) & (!g85) & (g82) & (!g86)));
	assign g88 = (((!i_28_) & (!sk[89]) & (i_29_)) + ((!i_28_) & (!sk[89]) & (i_29_)));
	assign g89 = (((!sk[90]) & (!i_32_) & (g88)) + ((!sk[90]) & (!i_32_) & (g88)));
	assign g90 = (((i_16_) & (!i_27_) & (sk[91]) & (!i_23_)) + ((!i_16_) & (i_27_) & (sk[91]) & (!i_23_)) + ((i_16_) & (!i_27_) & (!sk[91]) & (i_23_)) + ((!i_16_) & (!i_27_) & (sk[91]) & (i_23_)));
	assign g91 = (((!g2) & (!i_32_) & (!g84) & (!sk[92]) & (g90)) + ((g2) & (!i_32_) & (g84) & (!sk[92]) & (!g90)) + ((g2) & (!i_32_) & (g84) & (!sk[92]) & (!g90)));
	assign g92 = (((!g14) & (!g73) & (!g74) & (g89) & (!sk[93]) & (!g91)) + ((g14) & (!g73) & (g74) & (g89) & (!sk[93]) & (!g91)) + ((!g14) & (g73) & (!g74) & (!g89) & (sk[93]) & (g91)) + ((g14) & (!g73) & (!g74) & (!g89) & (!sk[93]) & (g91)));
	assign g93 = (((i_24_) & (!sk[94]) & (!i_23_) & (i_26_)) + ((!i_24_) & (sk[94]) & (!i_23_) & (!i_26_)));
	assign g94 = (((g19) & (!g93) & (!sk[95]) & (i_30_)) + ((g19) & (g93) & (sk[95]) & (!i_30_)));
	assign g95 = (((!i_17_) & (!i_21_) & (!i_2_) & (!sk[96]) & (g94) & (!g28)) + ((i_17_) & (!i_21_) & (!i_2_) & (!sk[96]) & (!g94) & (g28)) + ((!i_17_) & (!i_21_) & (!i_2_) & (!sk[96]) & (g94) & (g28)));
	assign g96 = (((!i_30_) & (!sk[97]) & (i_31_)) + ((!i_30_) & (sk[97]) & (!i_31_)));
	assign g97 = (((!sk[98]) & (i_28_) & (!i_29_) & (g96)) + ((sk[98]) & (!i_28_) & (!i_29_) & (g96)));
	assign g98 = (((!sk[99]) & (!g33) & (g97)) + ((!sk[99]) & (g33) & (g97)));
	assign g99 = (((!i_7_) & (!sk[100]) & (!i_32_) & (!g95) & (g66) & (!g98)) + ((!i_7_) & (!sk[100]) & (!i_32_) & (!g95) & (g66) & (g98)) + ((i_7_) & (!sk[100]) & (!i_32_) & (!g95) & (!g66) & (g98)) + ((!i_7_) & (sk[100]) & (!i_32_) & (g95) & (!g66) & (!g98)));
	assign g100 = (((!sk[101]) & (!g93) & (g34)) + ((!sk[101]) & (g93) & (g34)));
	assign g101 = (((!sk[102]) & (!g19) & (i_26_)) + ((sk[102]) & (g19) & (!i_26_)));
	assign g102 = (((!i_21_) & (!g33) & (!sk[103]) & (!g100) & (g101)) + ((i_21_) & (!g33) & (!sk[103]) & (g100) & (!g101)) + ((!i_21_) & (!g33) & (sk[103]) & (!g100) & (!g101)) + ((i_21_) & (!g33) & (!sk[103]) & (!g100) & (g101)) + ((!i_21_) & (!g33) & (!sk[103]) & (!g100) & (g101)));
	assign g103 = (((!i_32_) & (!g4) & (!sk[104]) & (!g102) & (g41)) + ((i_32_) & (!g4) & (!sk[104]) & (g102) & (!g41)) + ((!i_32_) & (g4) & (!sk[104]) & (!g102) & (g41)) + ((!i_32_) & (!g4) & (!sk[104]) & (!g102) & (g41)));
	assign g104 = (((!g83) & (!sk[105]) & (!g87) & (!g92) & (g99) & (!g103)) + ((g83) & (!sk[105]) & (!g87) & (!g92) & (!g99) & (g103)) + ((!g83) & (sk[105]) & (!g87) & (!g92) & (!g99) & (!g103)));
	assign g105 = (((g88) & (!sk[106]) & (!g7) & (g27)) + ((g88) & (!sk[106]) & (g7) & (g27)));
	assign g106 = (((!i_17_) & (!i_9_) & (!sk[107]) & (!g14) & (g72) & (!g105)) + ((i_17_) & (!i_9_) & (!sk[107]) & (!g14) & (!g72) & (g105)) + ((!i_17_) & (!i_9_) & (!sk[107]) & (g14) & (g72) & (g105)));
	assign g107 = (((!sk[108]) & (!i_23_) & (g54)) + ((!sk[108]) & (!i_23_) & (g54)));
	assign g108 = (((!sk[109]) & (!i_27_) & (g71)) + ((sk[109]) & (i_27_) & (!g71)));
	assign g109 = (((!i_23_) & (!g28) & (!g37) & (!sk[110]) & (g77) & (!g108)) + ((i_23_) & (!g28) & (!g37) & (!sk[110]) & (!g77) & (g108)) + ((!i_23_) & (g28) & (g37) & (!sk[110]) & (g77) & (!g108)));
	assign g110 = (((!sk[111]) & (!g7) & (!g54) & (!g6) & (g9)) + ((!sk[111]) & (g7) & (!g54) & (g6) & (!g9)) + ((!sk[111]) & (g7) & (g54) & (!g6) & (g9)));
	assign g111 = (((i_27_) & (!sk[112]) & (!g93) & (g88)) + ((!i_27_) & (sk[112]) & (g93) & (g88)));
	assign g112 = (((!i_3_) & (!i_18_) & (g14) & (!sk[113]) & (g12)) + ((!i_3_) & (!i_18_) & (!g14) & (!sk[113]) & (g12)) + ((i_3_) & (!i_18_) & (g14) & (!sk[113]) & (!g12)) + ((i_3_) & (!i_18_) & (g14) & (!sk[113]) & (!g12)));
	assign g113 = (((!g111) & (!i_9_) & (!g112) & (!sk[114]) & (g53)) + ((g111) & (!i_9_) & (g112) & (!sk[114]) & (!g53)) + ((g111) & (!i_9_) & (g112) & (!sk[114]) & (g53)));
	assign g114 = (((!i_21_) & (!g28) & (g7) & (!g9) & (!g100) & (g113)) + ((!i_21_) & (g28) & (g7) & (g9) & (g100) & (!g113)));
	assign g115 = (((!g77) & (!g76) & (!g107) & (!g109) & (!g110) & (!g114)) + ((!g77) & (!g76) & (!g107) & (!g109) & (!g110) & (!g114)) + ((!g77) & (!g76) & (!g107) & (!g109) & (!g110) & (!g114)));
	assign g116 = (((!g80) & (!g81) & (!sk[117]) & (!g104) & (g106) & (!g115)) + ((g80) & (!g81) & (!sk[117]) & (!g104) & (!g106) & (g115)) + ((g80) & (!g81) & (!sk[117]) & (g104) & (!g106) & (g115)));
	assign g117 = (((!g6) & (!g18) & (!g44) & (!sk[118]) & (g64) & (!g116)) + ((g6) & (!g18) & (!g44) & (!sk[118]) & (!g64) & (g116)) + ((g6) & (!g18) & (!g44) & (!sk[118]) & (!g64) & (g116)) + ((!g6) & (!g18) & (!g44) & (sk[118]) & (!g64) & (g116)));
	assign g118 = (((!i_35_) & (!sk[119]) & (i_36_)) + ((!i_35_) & (!sk[119]) & (i_36_)));
	assign g119 = (((!i_32_) & (!sk[120]) & (g118)) + ((!i_32_) & (!sk[120]) & (g118)));
	assign g120 = (((!g22) & (!sk[121]) & (!g108) & (!g60) & (g58)) + ((g22) & (!sk[121]) & (!g108) & (g60) & (!g58)) + ((!g22) & (!sk[121]) & (!g108) & (g60) & (g58)));
	assign g121 = (((!i_28_) & (!sk[122]) & (g71)) + ((!i_28_) & (sk[122]) & (!g71)));
	assign g122 = (((!i_34_) & (!sk[123]) & (!i_29_) & (!g96) & (g121)) + ((i_34_) & (!sk[123]) & (!i_29_) & (g96) & (!g121)) + ((!i_34_) & (!sk[123]) & (!i_29_) & (g96) & (g121)));
	assign g123 = (((!g100) & (!sk[124]) & (!g56) & (!g119) & (g120) & (!g122)) + ((!g100) & (!sk[124]) & (!g56) & (g119) & (g120) & (!g122)) + ((g100) & (!sk[124]) & (!g56) & (!g119) & (!g120) & (g122)) + ((!g100) & (sk[124]) & (!g56) & (g119) & (!g120) & (g122)) + ((g100) & (sk[124]) & (g56) & (g119) & (!g120) & (!g122)));
	assign g124 = (((!g95) & (!sk[125]) & (!i_31_) & (!i_8_) & (g102) & (!g61)) + ((g95) & (!sk[125]) & (!i_31_) & (!i_8_) & (!g102) & (g61)) + ((g95) & (sk[125]) & (!i_31_) & (!i_8_) & (!g102) & (!g61)) + ((!g95) & (sk[125]) & (!i_31_) & (!i_8_) & (!g102) & (g61)));
	assign g125 = (((!i_16_) & (!sk[126]) & (!g22) & (!g33) & (g9)) + ((i_16_) & (!sk[126]) & (!g22) & (g33) & (!g9)) + ((!i_16_) & (!sk[126]) & (!g22) & (g33) & (g9)));
	assign g126 = (((!i_34_) & (!sk[127]) & (!g57) & (!g34) & (g125)) + ((i_34_) & (!sk[127]) & (!g57) & (g34) & (!g125)) + ((i_34_) & (!sk[127]) & (g57) & (g34) & (g125)));
	assign g127 = (((!g1) & (!sk[0]) & (!g108) & (!g50) & (g124) & (!g126)) + ((g1) & (!sk[0]) & (!g108) & (!g50) & (!g124) & (g126)) + ((!g1) & (sk[0]) & (!g108) & (!g50) & (!g124) & (!g126)) + ((!g1) & (sk[0]) & (g108) & (!g50) & (!g124) & (!g126)) + ((!g1) & (sk[0]) & (!g108) & (!g50) & (!g124) & (!g126)));
	assign g128 = (((!sk[1]) & (!i_7_) & (i_10_)) + ((!sk[1]) & (i_7_) & (i_10_)));
	assign g129 = (((!i_17_) & (!i_12_) & (!sk[2]) & (!i_13_) & (g54) & (!g128)) + ((i_17_) & (!i_12_) & (!sk[2]) & (!i_13_) & (!g54) & (g128)) + ((!i_17_) & (!i_12_) & (!sk[2]) & (i_13_) & (g54) & (g128)) + ((!i_17_) & (!i_12_) & (!sk[2]) & (i_13_) & (g54) & (g128)));
	assign g130 = (((!i_27_) & (!sk[3]) & (g88)) + ((!i_27_) & (!sk[3]) & (g88)));
	assign g131 = (((!sk[4]) & (g33) & (!g130) & (i_22_)) + ((!sk[4]) & (g33) & (g130) & (i_22_)));
	assign g132 = (((i_33_) & (!sk[5]) & (g57)) + ((!i_33_) & (!sk[5]) & (g57)));
	assign g133 = (((!sk[6]) & (g33) & (!g84) & (g132)) + ((!sk[6]) & (g33) & (g84) & (g132)));
	assign g134 = (((!sk[7]) & (i_17_) & (!i_12_) & (g54)) + ((sk[7]) & (!i_17_) & (!i_12_) & (g54)) + ((!sk[7]) & (i_17_) & (!i_12_) & (g54)));
	assign g135 = (((!i_12_) & (!g45) & (i_25_) & (!g131) & (g133) & (!g134)) + ((!i_12_) & (!g45) & (!i_25_) & (g131) & (!g133) & (g134)) + ((!i_12_) & (g45) & (!i_25_) & (g131) & (!g133) & (!g134)));
	assign g136 = (((!i_28_) & (!i_31_) & (!sk[9]) & (!i_29_) & (g5)) + ((i_28_) & (!i_31_) & (!sk[9]) & (i_29_) & (!g5)) + ((!i_28_) & (i_31_) & (sk[9]) & (!i_29_) & (!g5)));
	assign g137 = (((!sk[10]) & (i_21_) & (!i_30_) & (g33)) + ((!sk[10]) & (i_21_) & (!i_30_) & (g33)));
	assign g138 = (((!i_28_) & (i_14_) & (!g132) & (!i_25_) & (g133) & (!g137)) + ((!i_28_) & (i_14_) & (g132) & (!i_25_) & (!g133) & (g137)) + ((!i_28_) & (!i_14_) & (g132) & (i_25_) & (!g133) & (g137)));
	assign g139 = (((!i_34_) & (!g129) & (!g135) & (!sk[12]) & (g136) & (!g138)) + ((i_34_) & (!g129) & (!g135) & (!sk[12]) & (!g136) & (g138)) + ((i_34_) & (!g129) & (g135) & (sk[12]) & (!g136) & (!g138)) + ((i_34_) & (g129) & (!g135) & (!sk[12]) & (g136) & (!g138)));
	assign g140 = (((!sk[13]) & (!i_24_) & (!i_28_) & (!i_26_) & (i_30_)) + ((!sk[13]) & (i_24_) & (!i_28_) & (i_26_) & (!i_30_)) + ((sk[13]) & (!i_24_) & (!i_28_) & (!i_26_) & (!i_30_)));
	assign g141 = (((!i_33_) & (!i_28_) & (!g2) & (!sk[14]) & (g86)) + ((i_33_) & (!i_28_) & (g2) & (!sk[14]) & (!g86)) + ((i_33_) & (!i_28_) & (g2) & (!sk[14]) & (!g86)));
	assign g142 = (((!sk[15]) & (!i_34_) & (!g132) & (!g140) & (g141)) + ((sk[15]) & (!i_34_) & (!g132) & (!g140) & (!g141)) + ((sk[15]) & (!i_34_) & (!g132) & (!g140) & (!g141)) + ((!sk[15]) & (i_34_) & (!g132) & (g140) & (!g141)));
	assign g143 = (((i_33_) & (!sk[16]) & (!g2) & (g1)) + ((i_33_) & (!sk[16]) & (g2) & (g1)));
	assign g144 = (((!i_34_) & (!sk[17]) & (!g71) & (!g84) & (g132)) + ((i_34_) & (!sk[17]) & (!g71) & (g84) & (!g132)) + ((!i_34_) & (!sk[17]) & (!g71) & (g84) & (g132)));
	assign g145 = (((g86) & (!g143) & (!sk[18]) & (g144)) + ((g86) & (!g143) & (sk[18]) & (!g144)) + ((!g86) & (!g143) & (sk[18]) & (!g144)));
	assign g146 = (((!sk[19]) & (!i_14_) & (!i_21_) & (!g142) & (i_25_) & (!g145)) + ((!sk[19]) & (!i_14_) & (!i_21_) & (!g142) & (i_25_) & (!g145)) + ((!sk[19]) & (!i_14_) & (i_21_) & (!g142) & (i_25_) & (!g145)) + ((!sk[19]) & (i_14_) & (!i_21_) & (!g142) & (!i_25_) & (g145)) + ((sk[19]) & (i_14_) & (!i_21_) & (!g142) & (!i_25_) & (!g145)) + ((!sk[19]) & (i_14_) & (i_21_) & (!g142) & (!i_25_) & (g145)));
	assign g147 = (((!sk[20]) & (g2) & (!g86) & (i_22_)) + ((!sk[20]) & (g2) & (!g86) & (i_22_)));
	assign g148 = (((!i_34_) & (i_35_) & (!g71) & (!i_30_) & (!i_32_) & (!i_31_)) + ((!i_34_) & (!i_35_) & (!g71) & (!i_30_) & (!i_32_) & (!i_31_)));
	assign g149 = (((!sk[22]) & (!i_21_) & (!g88) & (!i_20_) & (g147) & (!g148)) + ((!sk[22]) & (!i_21_) & (g88) & (!i_20_) & (g147) & (!g148)) + ((!sk[22]) & (i_21_) & (!g88) & (!i_20_) & (!g147) & (g148)) + ((sk[22]) & (!i_21_) & (g88) & (i_20_) & (!g147) & (g148)));
	assign g150 = (((!i_17_) & (sk[23]) & (!i_12_) & (g45)) + ((i_17_) & (!sk[23]) & (!i_12_) & (g45)) + ((!i_17_) & (sk[23]) & (!i_12_) & (g45)));
	assign g151 = (((g33) & (i_29_) & (g101) & (g55) & (i_22_) & (!g150)) + ((g33) & (i_29_) & (g101) & (!g55) & (i_22_) & (g150)));
	assign g152 = (((!i_12_) & (!sk[25]) & (g28)) + ((!i_12_) & (!sk[25]) & (g28)));
	assign g153 = (((!sk[26]) & (!i_21_) & (!i_2_) & (!g111) & (g152) & (!i_20_)) + ((!sk[26]) & (i_21_) & (!i_2_) & (!g111) & (!g152) & (i_20_)) + ((!sk[26]) & (!i_21_) & (i_2_) & (g111) & (g152) & (!i_20_)));
	assign g154 = (((!i_34_) & (!i_23_) & (!i_26_) & (g88) & (!sk[27]) & (!i_22_)) + ((i_34_) & (!i_23_) & (!i_26_) & (!g88) & (!sk[27]) & (i_22_)) + ((i_34_) & (!i_23_) & (!i_26_) & (g88) & (!sk[27]) & (i_22_)) + ((!i_34_) & (!i_23_) & (!i_26_) & (g88) & (!sk[27]) & (i_22_)));
	assign g155 = (((!sk[28]) & (!i_24_) & (!i_30_) & (!g57) & (g153) & (!g154)) + ((sk[28]) & (!i_24_) & (i_30_) & (!g57) & (!g153) & (!g154)) + ((sk[28]) & (!i_24_) & (!i_30_) & (!g57) & (!g153) & (!g154)) + ((sk[28]) & (!i_24_) & (!i_30_) & (!g57) & (!g153) & (!g154)) + ((!sk[28]) & (i_24_) & (!i_30_) & (!g57) & (!g153) & (g154)));
	assign g156 = (((!i_34_) & (!g53) & (!g131) & (!sk[29]) & (g151) & (!g155)) + ((i_34_) & (!g53) & (!g131) & (!sk[29]) & (!g151) & (g155)) + ((!i_34_) & (!g53) & (!g131) & (sk[29]) & (!g151) & (g155)) + ((!i_34_) & (!g53) & (!g131) & (sk[29]) & (!g151) & (g155)) + ((!i_34_) & (!g53) & (!g131) & (sk[29]) & (!g151) & (g155)));
	assign g157 = (((!sk[30]) & (i_17_) & (!i_12_) & (g28)) + ((sk[30]) & (!i_17_) & (!i_12_) & (g28)) + ((!sk[30]) & (i_17_) & (!i_12_) & (g28)));
	assign g158 = (((!i_16_) & (!i_12_) & (!i_13_) & (i_14_) & (!g90) & (!g38)) + ((!i_16_) & (!i_12_) & (!i_13_) & (i_14_) & (!g90) & (g38)));
	assign g159 = (((i_21_) & (!i_22_) & (!sk[32]) & (i_20_)) + ((!i_21_) & (!i_22_) & (sk[32]) & (i_20_)));
	assign g160 = (((!g111) & (g143) & (!sk[33]) & (!g157) & (g158) & (!g159)) + ((!g111) & (!g143) & (!sk[33]) & (!g157) & (g158) & (!g159)) + ((g111) & (!g143) & (!sk[33]) & (!g157) & (!g158) & (g159)) + ((g111) & (!g143) & (!sk[33]) & (g157) & (!g158) & (g159)));
	assign g161 = (((!sk[34]) & (!i_16_) & (!i_36_) & (!g33) & (g70) & (!g73)) + ((!sk[34]) & (i_16_) & (!i_36_) & (!g33) & (!g70) & (g73)) + ((sk[34]) & (!i_16_) & (i_36_) & (g33) & (!g70) & (g73)));
	assign g162 = (((g33) & (!i_8_) & (!sk[35]) & (g157)) + ((g33) & (!i_8_) & (!sk[35]) & (g157)));
	assign g163 = (((i_34_) & (!g96) & (g34) & (g161) & (!g118) & (!g162)) + ((i_34_) & (g96) & (g34) & (!g161) & (g118) & (g162)));
	assign g164 = (((i_33_) & (!sk[37]) & (i_25_)) + ((!i_33_) & (!sk[37]) & (i_25_)));
	assign g165 = (((!sk[38]) & (!g134) & (g164)) + ((!sk[38]) & (g134) & (g164)));
	assign g166 = (((!i_27_) & (!sk[39]) & (!i_28_) & (!i_31_) & (g129) & (!g165)) + ((i_27_) & (!sk[39]) & (!i_28_) & (!i_31_) & (!g129) & (g165)) + ((!i_27_) & (!sk[39]) & (!i_28_) & (i_31_) & (g129) & (!g165)) + ((!i_27_) & (sk[39]) & (!i_28_) & (!i_31_) & (!g129) & (g165)));
	assign g167 = (((!i_24_) & (!i_34_) & (!i_35_) & (i_23_) & (!sk[40]) & (!i_21_)) + ((i_24_) & (!i_34_) & (!i_35_) & (!i_23_) & (!sk[40]) & (i_21_)) + ((!i_24_) & (i_34_) & (!i_35_) & (!i_23_) & (sk[40]) & (i_21_)) + ((!i_24_) & (!i_34_) & (i_35_) & (!i_23_) & (sk[40]) & (i_21_)));
	assign g168 = (((!i_27_) & (!i_28_) & (!g93) & (!sk[41]) & (i_31_) & (!g4)) + ((!i_27_) & (!i_28_) & (!g93) & (!sk[41]) & (i_31_) & (g4)) + ((i_27_) & (!i_28_) & (!g93) & (!sk[41]) & (!i_31_) & (g4)) + ((!i_27_) & (!i_28_) & (g93) & (!sk[41]) & (i_31_) & (!g4)));
	assign g169 = (((!i_16_) & (i_33_) & (!i_17_) & (!i_12_) & (!i_13_) & (i_14_)) + ((!i_16_) & (i_33_) & (!i_17_) & (!i_12_) & (!i_13_) & (i_14_)));
	assign g170 = (((!g20) & (!i_34_) & (!i_35_) & (!sk[43]) & (i_21_)) + ((g20) & (!i_34_) & (i_35_) & (!sk[43]) & (!i_21_)) + ((g20) & (i_34_) & (!i_35_) & (!sk[43]) & (i_21_)) + ((!g20) & (!i_34_) & (i_35_) & (!sk[43]) & (i_21_)));
	assign g171 = (((!g3) & (!g168) & (!g129) & (g169) & (!sk[44]) & (!g170)) + ((!g3) & (g168) & (g129) & (!g169) & (sk[44]) & (!g170)) + ((g3) & (!g168) & (!g129) & (g169) & (!sk[44]) & (g170)) + ((g3) & (!g168) & (!g129) & (!g169) & (!sk[44]) & (g170)));
	assign g172 = (((!g160) & (!g163) & (!g166) & (g167) & (!sk[45]) & (!g171)) + ((g160) & (!g163) & (!g166) & (!g167) & (!sk[45]) & (g171)) + ((!g160) & (!g163) & (!g166) & (!g167) & (sk[45]) & (!g171)) + ((!g160) & (!g163) & (!g166) & (!g167) & (sk[45]) & (!g171)));
	assign g173 = (((!i_3_) & (!i_18_) & (!i_4_) & (i_5_) & (!sk[46]) & (!g31)) + ((i_3_) & (!i_18_) & (!i_4_) & (!i_5_) & (!sk[46]) & (g31)) + ((i_3_) & (!i_18_) & (!i_4_) & (!i_5_) & (!sk[46]) & (g31)));
	assign g174 = (((!sk[47]) & (!i_7_) & (!i_9_) & (!g14) & (g12)) + ((!sk[47]) & (i_7_) & (!i_9_) & (g14) & (!g12)) + ((!sk[47]) & (!i_7_) & (!i_9_) & (g14) & (g12)));
	assign g175 = (((!sk[48]) & (!i_36_) & (!g89) & (!g173) & (g174)) + ((!sk[48]) & (i_36_) & (!g89) & (g173) & (!g174)) + ((!sk[48]) & (i_36_) & (g89) & (g173) & (!g174)) + ((!sk[48]) & (i_36_) & (g89) & (!g173) & (g174)));
	assign g176 = (((!i_2_) & (!sk[49]) & (!g14) & (!i_8_) & (g118)) + ((i_2_) & (!sk[49]) & (!g14) & (i_8_) & (!g118)) + ((!i_2_) & (sk[49]) & (!g14) & (!i_8_) & (!g118)) + ((!i_2_) & (!sk[49]) & (!g14) & (!i_8_) & (g118)) + ((!i_2_) & (!sk[49]) & (!g14) & (i_8_) & (g118)));
	assign g177 = (((!g88) & (!i_9_) & (!sk[50]) & (!g12) & (g176)) + ((g88) & (!i_9_) & (!sk[50]) & (g12) & (!g176)) + ((g88) & (!i_9_) & (!sk[50]) & (g12) & (!g176)));
	assign g178 = (((!i_4_) & (!i_5_) & (!g48) & (!sk[51]) & (g118)) + ((i_4_) & (!i_5_) & (g48) & (!sk[51]) & (!g118)) + ((!i_4_) & (!i_5_) & (g48) & (!sk[51]) & (g118)));
	assign g179 = (((!i_2_) & (g88) & (!i_9_) & (i_3_) & (!i_18_) & (g178)) + ((i_2_) & (g88) & (!i_9_) & (i_3_) & (!i_18_) & (!g178)));
	assign g180 = (((!g53) & (!g72) & (!g175) & (!sk[53]) & (g177) & (!g179)) + ((g53) & (g72) & (!g175) & (!sk[53]) & (g177) & (!g179)) + ((g53) & (g72) & (!g175) & (!sk[53]) & (!g177) & (g179)) + ((g53) & (!g72) & (!g175) & (!sk[53]) & (!g177) & (g179)) + ((g53) & (g72) & (g175) & (sk[53]) & (!g177) & (!g179)));
	assign g181 = (((!sk[54]) & (!i_24_) & (!i_34_) & (!i_35_) & (i_26_)) + ((!sk[54]) & (i_24_) & (!i_34_) & (i_35_) & (!i_26_)) + ((sk[54]) & (i_24_) & (!i_34_) & (!i_35_) & (!i_26_)) + ((!sk[54]) & (!i_24_) & (!i_34_) & (!i_35_) & (i_26_)) + ((!sk[54]) & (i_24_) & (i_34_) & (i_35_) & (!i_26_)));
	assign g182 = (((!i_27_) & (!sk[55]) & (!i_36_) & (!g84) & (g181)) + ((i_27_) & (!sk[55]) & (!i_36_) & (g84) & (!g181)) + ((!i_27_) & (sk[55]) & (i_36_) & (g84) & (!g181)));
	assign g183 = (((!i_23_) & (!i_7_) & (!i_8_) & (!sk[56]) & (g152) & (!g182)) + ((!i_23_) & (i_7_) & (!i_8_) & (!sk[56]) & (g152) & (!g182)) + ((i_23_) & (!i_7_) & (!i_8_) & (!sk[56]) & (!g152) & (g182)) + ((!i_23_) & (!i_7_) & (!i_8_) & (!sk[56]) & (g152) & (g182)));
	assign g184 = (((!i_7_) & (!sk[57]) & (!i_9_) & (!g712) & (g180) & (!g183)) + ((i_7_) & (!sk[57]) & (!i_9_) & (!g712) & (!g180) & (g183)) + ((!i_7_) & (sk[57]) & (!i_9_) & (!g712) & (!g180) & (!g183)) + ((i_7_) & (!sk[57]) & (i_9_) & (!g712) & (!g180) & (g183)) + ((i_7_) & (!sk[57]) & (!i_9_) & (g712) & (!g180) & (g183)));
	assign g185 = (((!g146) & (!g149) & (!sk[58]) & (!g156) & (g172) & (!g184)) + ((g146) & (!g149) & (!sk[58]) & (!g156) & (!g172) & (g184)) + ((!g146) & (!g149) & (!sk[58]) & (g156) & (g172) & (g184)));
	assign g186 = (((!g118) & (!sk[59]) & (!g123) & (!g127) & (g139) & (!g185)) + ((g118) & (!sk[59]) & (!g123) & (!g127) & (!g139) & (g185)) + ((!g118) & (sk[59]) & (!g123) & (!g127) & (!g139) & (g185)) + ((!g118) & (sk[59]) & (!g123) & (g127) & (!g139) & (g185)));
	assign g187 = (((!sk[60]) & (!g27) & (!g30) & (!g49) & (g118)) + ((!sk[60]) & (g27) & (!g30) & (g49) & (!g118)) + ((sk[60]) & (!g27) & (!g30) & (!g49) & (!g118)) + ((sk[60]) & (!g27) & (!g30) & (!g49) & (!g118)) + ((sk[60]) & (!g27) & (!g30) & (!g49) & (!g118)));
	assign g188 = (((!sk[61]) & (i_17_) & (!i_36_) & (g33)) + ((sk[61]) & (!i_17_) & (i_36_) & (g33)));
	assign g189 = (((!i_29_) & (!g69) & (!g119) & (g187) & (!sk[62]) & (!g188)) + ((i_29_) & (!g69) & (!g119) & (!g187) & (!sk[62]) & (g188)) + ((!i_29_) & (g69) & (g119) & (!g187) & (sk[62]) & (!g188)) + ((!i_29_) & (!g69) & (!g119) & (!g187) & (sk[62]) & (g188)));
	assign g190 = (((i_3_) & (!sk[63]) & (!g14) & (g15)) + ((i_3_) & (!sk[63]) & (g14) & (g15)));
	assign g191 = (((!i_16_) & (!i_17_) & (!i_13_) & (i_14_) & (!sk[64]) & (!i_10_)) + ((i_16_) & (!i_17_) & (!i_13_) & (!i_14_) & (!sk[64]) & (i_10_)) + ((!i_16_) & (!i_17_) & (i_13_) & (!i_14_) & (sk[64]) & (!i_10_)) + ((!i_16_) & (!i_17_) & (!i_13_) & (!i_14_) & (sk[64]) & (!i_10_)));
	assign g192 = (((!i_31_) & (!g14) & (!sk[65]) & (!g119) & (g152)) + ((i_31_) & (!g14) & (!sk[65]) & (g119) & (!g152)) + ((!i_31_) & (g14) & (!sk[65]) & (g119) & (g152)));
	assign g193 = (((!i_36_) & (!i_7_) & (!sk[66]) & (!i_32_) & (g14)) + ((i_36_) & (!i_7_) & (!sk[66]) & (i_32_) & (!g14)) + ((i_36_) & (!i_7_) & (!sk[66]) & (!i_32_) & (g14)));
	assign g194 = (((!i_9_) & (!sk[67]) & (!g14) & (!g45) & (g13) & (!g119)) + ((i_9_) & (!sk[67]) & (!g14) & (!g45) & (!g13) & (g119)) + ((!i_9_) & (!sk[67]) & (g14) & (g45) & (g13) & (g119)));
	assign g195 = (((i_9_) & (!g176) & (!g191) & (!g192) & (!g193) & (!g194)) + ((!i_9_) & (!g176) & (!g191) & (!g192) & (!g193) & (!g194)) + ((!i_9_) & (g176) & (!g191) & (!g192) & (!g193) & (!g194)));
	assign g196 = (((!i_29_) & (!g45) & (!sk[69]) & (!g119) & (g190) & (!g195)) + ((i_29_) & (!g45) & (!sk[69]) & (!g119) & (!g190) & (g195)) + ((i_29_) & (!g45) & (sk[69]) & (!g119) & (!g190) & (!g195)) + ((i_29_) & (g45) & (!sk[69]) & (g119) & (g190) & (!g195)));
	assign g197 = (((!sk[70]) & (!i_30_) & (g7)) + ((!sk[70]) & (!i_30_) & (g7)));
	assign g198 = (((!i_17_) & (!i_36_) & (!i_2_) & (g28) & (!sk[71]) & (!g197)) + ((i_17_) & (!i_36_) & (!i_2_) & (!g28) & (!sk[71]) & (g197)) + ((!i_17_) & (i_36_) & (!i_2_) & (g28) & (!sk[71]) & (g197)));
	assign g199 = (((!g86) & (!g118) & (!sk[72]) & (!g152) & (g198)) + ((!g86) & (!g118) & (sk[72]) & (!g152) & (!g198)) + ((!g86) & (!g118) & (sk[72]) & (!g152) & (!g198)) + ((g86) & (!g118) & (!sk[72]) & (g152) & (!g198)));
	assign g200 = (((!i_21_) & (!sk[73]) & (!g33) & (!g189) & (g196) & (!g199)) + ((i_21_) & (sk[73]) & (!g33) & (!g189) & (!g196) & (!g199)) + ((!i_21_) & (sk[73]) & (!g33) & (!g189) & (!g196) & (!g199)) + ((i_21_) & (!sk[73]) & (!g33) & (!g189) & (!g196) & (g199)) + ((!i_21_) & (sk[73]) & (!g33) & (!g189) & (!g196) & (g199)));
	assign g201 = (((!g57) & (!i_29_) & (!g96) & (g125) & (!sk[74]) & (!g162)) + ((g57) & (!i_29_) & (!g96) & (g125) & (!sk[74]) & (!g162)) + ((g57) & (!i_29_) & (!g96) & (!g125) & (!sk[74]) & (g162)) + ((!g57) & (!i_29_) & (g96) & (!g125) & (sk[74]) & (g162)));
	assign g202 = (((!i_12_) & (!g33) & (!i_29_) & (!sk[75]) & (g54) & (!i_22_)) + ((i_12_) & (!g33) & (!i_29_) & (!sk[75]) & (!g54) & (i_22_)) + ((!i_12_) & (g33) & (i_29_) & (!sk[75]) & (g54) & (i_22_)));
	assign g203 = (((!i_29_) & (!g161) & (!sk[76]) & (!g118) & (g201) & (!g202)) + ((i_29_) & (!g161) & (!sk[76]) & (!g118) & (!g201) & (g202)) + ((i_29_) & (!g161) & (sk[76]) & (!g118) & (!g201) & (!g202)) + ((!i_29_) & (!g161) & (sk[76]) & (!g118) & (!g201) & (!g202)) + ((i_29_) & (!g161) & (!sk[76]) & (!g118) & (g201) & (!g202)) + ((!i_29_) & (!g161) & (!sk[76]) & (!g118) & (g201) & (!g202)));
	assign g204 = (((!sk[77]) & (!g2) & (!i_21_) & (!g130) & (i_22_) & (!i_20_)) + ((!sk[77]) & (g2) & (!i_21_) & (g130) & (i_22_) & (!i_20_)) + ((!sk[77]) & (g2) & (!i_21_) & (!g130) & (!i_22_) & (i_20_)) + ((!sk[77]) & (g2) & (!i_21_) & (g130) & (!i_22_) & (i_20_)));
	assign g205 = (((!i_24_) & (!i_27_) & (!i_28_) & (i_29_) & (!g86) & (!g157)) + ((!i_24_) & (!i_27_) & (!i_28_) & (i_29_) & (!g86) & (g157)));
	assign g206 = (((!i_34_) & (!i_21_) & (!i_20_) & (!sk[79]) & (g205)) + ((i_34_) & (!i_21_) & (i_20_) & (!sk[79]) & (!g205)) + ((i_34_) & (!i_21_) & (i_20_) & (!sk[79]) & (g205)));
	assign g207 = (((i_34_) & (!sk[80]) & (!g34) & (g101)) + ((!i_34_) & (sk[80]) & (!g34) & (!g101)) + ((!i_34_) & (sk[80]) & (!g34) & (!g101)));
	assign g208 = (((!sk[81]) & (!i_33_) & (!i_24_) & (!i_13_) & (i_14_) & (!i_25_)) + ((!sk[81]) & (i_33_) & (!i_24_) & (!i_13_) & (!i_14_) & (i_25_)) + ((!sk[81]) & (i_33_) & (!i_24_) & (!i_13_) & (i_14_) & (!i_25_)) + ((!sk[81]) & (i_33_) & (!i_24_) & (!i_13_) & (!i_14_) & (i_25_)));
	assign g209 = (((!sk[82]) & (!i_16_) & (!i_17_) & (!i_12_) & (g207) & (!g208)) + ((!sk[82]) & (i_16_) & (!i_17_) & (!i_12_) & (!g207) & (g208)) + ((sk[82]) & (!i_16_) & (!i_17_) & (!i_12_) & (!g207) & (g208)) + ((sk[82]) & (!i_16_) & (!i_17_) & (!i_12_) & (!g207) & (g208)));
	assign g210 = (((!i_3_) & (!sk[83]) & (!i_18_) & (!i_11_) & (i_19_) & (!g128)) + ((i_3_) & (!sk[83]) & (!i_18_) & (!i_11_) & (!i_19_) & (g128)) + ((i_3_) & (!sk[83]) & (!i_18_) & (!i_11_) & (!i_19_) & (g128)) + ((!i_3_) & (sk[83]) & (!i_18_) & (!i_11_) & (!i_19_) & (g128)));
	assign g211 = (((!i_27_) & (!i_28_) & (!g2) & (i_31_) & (!sk[84]) & (!i_29_)) + ((i_27_) & (!i_28_) & (!g2) & (!i_31_) & (!sk[84]) & (i_29_)) + ((!i_27_) & (!i_28_) & (g2) & (i_31_) & (!sk[84]) & (!i_29_)));
	assign g212 = (((!g150) & (!sk[85]) & (!g209) & (!g210) & (g211)) + ((g150) & (!sk[85]) & (!g209) & (g210) & (!g211)) + ((!g150) & (sk[85]) & (!g209) & (!g210) & (!g211)) + ((!g150) & (sk[85]) & (!g209) & (!g210) & (!g211)) + ((!g150) & (sk[85]) & (!g209) & (!g210) & (!g211)));
	assign g213 = (((!g28) & (!g108) & (!sk[86]) & (!g60) & (g51) & (!g118)) + ((g28) & (!g108) & (!sk[86]) & (!g60) & (!g51) & (g118)) + ((g28) & (!g108) & (!sk[86]) & (g60) & (g51) & (g118)));
	assign g214 = (((!i_27_) & (!g2) & (!sk[87]) & (!g1) & (g165) & (!g213)) + ((i_27_) & (!g2) & (!sk[87]) & (!g1) & (!g165) & (g213)) + ((!i_27_) & (!g2) & (sk[87]) & (!g1) & (!g165) & (!g213)) + ((i_27_) & (!g2) & (!sk[87]) & (!g1) & (g165) & (!g213)) + ((!i_27_) & (!g2) & (!sk[87]) & (!g1) & (g165) & (!g213)) + ((!i_27_) & (!g2) & (!sk[87]) & (!g1) & (g165) & (!g213)));
	assign g215 = (((!sk[88]) & (!g157) & (!g204) & (!g206) & (g212) & (!g214)) + ((!sk[88]) & (g157) & (!g204) & (!g206) & (!g212) & (g214)) + ((!sk[88]) & (!g157) & (!g204) & (!g206) & (g212) & (g214)) + ((!sk[88]) & (!g157) & (!g204) & (!g206) & (g212) & (g214)));
	assign g216 = (((!i_23_) & (!g101) & (!sk[89]) & (!g200) & (g203) & (!g215)) + ((i_23_) & (!g101) & (sk[89]) & (!g200) & (!g203) & (!g215)) + ((i_23_) & (!g101) & (!sk[89]) & (g200) & (g203) & (!g215)) + ((!i_23_) & (!g101) & (sk[89]) & (!g200) & (!g203) & (g215)) + ((i_23_) & (!g101) & (!sk[89]) & (!g200) & (!g203) & (g215)) + ((!i_23_) & (!g101) & (!sk[89]) & (g200) & (g203) & (g215)));
	assign g217 = (((!g2) & (!i_32_) & (!sk[90]) & (!g84) & (g38)) + ((g2) & (!i_32_) & (!sk[90]) & (g84) & (!g38)) + ((g2) & (!i_32_) & (!sk[90]) & (g84) & (g38)));
	assign g218 = (((!i_17_) & (!g33) & (!i_29_) & (!sk[91]) & (g70) & (!g101)) + ((i_17_) & (!g33) & (!i_29_) & (!sk[91]) & (!g70) & (g101)) + ((!i_17_) & (g33) & (!i_29_) & (sk[91]) & (!g70) & (g101)));
	assign g219 = (((!i_34_) & (!g70) & (!g35) & (g217) & (!sk[92]) & (!g218)) + ((i_34_) & (!g70) & (!g35) & (!g217) & (!sk[92]) & (g218)) + ((!i_34_) & (!g70) & (!g35) & (!g217) & (sk[92]) & (!g218)) + ((!i_34_) & (g70) & (!g35) & (!g217) & (sk[92]) & (!g218)) + ((!i_34_) & (!g70) & (!g35) & (!g217) & (sk[92]) & (!g218)));
	assign g220 = (((!sk[93]) & (!g19) & (!i_30_) & (!g130) & (g14)) + ((!sk[93]) & (!g19) & (!i_30_) & (g130) & (g14)) + ((sk[93]) & (g19) & (!i_30_) & (!g130) & (!g14)) + ((!sk[93]) & (g19) & (!i_30_) & (g130) & (!g14)));
	assign g221 = (((!i_12_) & (!i_7_) & (!sk[94]) & (!i_9_) & (g702)) + ((i_12_) & (!i_7_) & (!sk[94]) & (i_9_) & (!g702)) + ((!i_12_) & (i_7_) & (!sk[94]) & (!i_9_) & (g702)));
	assign g222 = (((!i_12_) & (!i_21_) & (!i_36_) & (!sk[95]) & (g93) & (!g7)) + ((i_12_) & (!i_21_) & (!i_36_) & (!sk[95]) & (!g93) & (g7)) + ((!i_12_) & (!i_21_) & (i_36_) & (!sk[95]) & (g93) & (g7)));
	assign g223 = (((!i_28_) & (!sk[96]) & (g96)) + ((!i_28_) & (!sk[96]) & (g96)));
	assign g224 = (((!sk[97]) & (!i_2_) & (!g88) & (!g119) & (i_0_) & (!g223)) + ((!sk[97]) & (!i_2_) & (g88) & (!g119) & (i_0_) & (!g223)) + ((!sk[97]) & (i_2_) & (!g88) & (!g119) & (!i_0_) & (g223)) + ((sk[97]) & (!i_2_) & (!g88) & (g119) & (!i_0_) & (g223)));
	assign g225 = (((g7) & (!sk[98]) & (!g23) & (g182)) + ((g7) & (!sk[98]) & (g23) & (g182)));
	assign g226 = (((i_12_) & (!sk[99]) & (!g88) & (i_0_)) + ((!i_12_) & (sk[99]) & (g88) & (i_0_)));
	assign g227 = (((!i_17_) & (!g72) & (!g224) & (!sk[100]) & (g225) & (!g226)) + ((!i_17_) & (!g72) & (!g224) & (sk[100]) & (!g225) & (!g226)) + ((i_17_) & (!g72) & (!g224) & (!sk[100]) & (!g225) & (g226)) + ((i_17_) & (!g72) & (!g224) & (sk[100]) & (!g225) & (!g226)) + ((!i_17_) & (!g72) & (!g224) & (sk[100]) & (!g225) & (!g226)));
	assign g228 = (((!sk[101]) & (!g220) & (!g221) & (!g222) & (g227)) + ((!sk[101]) & (g220) & (!g221) & (g222) & (!g227)) + ((!sk[101]) & (!g220) & (!g221) & (!g222) & (g227)) + ((!sk[101]) & (!g220) & (!g221) & (!g222) & (g227)));
	assign g229 = (((!i_16_) & (!sk[102]) & (!i_36_) & (!i_7_) & (g219) & (!g228)) + ((i_16_) & (!sk[102]) & (!i_36_) & (!i_7_) & (!g219) & (g228)) + ((!i_16_) & (sk[102]) & (!i_36_) & (!i_7_) & (!g219) & (!g228)) + ((!i_16_) & (sk[102]) & (i_36_) & (!i_7_) & (!g219) & (!g228)));
	assign g230 = (((i_16_) & (!sk[103]) & (!i_17_) & (g702)) + ((!i_16_) & (sk[103]) & (!i_17_) & (g702)));
	assign g231 = (((!i_7_) & (!sk[104]) & (!i_9_) & (!g23) & (g230) & (!g712)) + ((i_7_) & (!sk[104]) & (!i_9_) & (!g23) & (g230) & (!g712)) + ((i_7_) & (!sk[104]) & (!i_9_) & (!g23) & (!g230) & (g712)) + ((i_7_) & (sk[104]) & (!i_9_) & (g23) & (!g230) & (!g712)));
	assign g232 = (((!i_28_) & (!i_12_) & (!i_30_) & (!i_31_) & (!i_29_) & (!g14)) + ((!i_28_) & (!i_12_) & (!i_30_) & (!i_31_) & (i_29_) & (g14)));
	assign g233 = (((!i_23_) & (!i_8_) & (!g108) & (!sk[106]) & (g118) & (!g232)) + ((i_23_) & (!i_8_) & (!g108) & (!sk[106]) & (!g118) & (g232)) + ((!i_23_) & (!i_8_) & (!g108) & (!sk[106]) & (g118) & (g232)));
	assign g234 = (((!sk[107]) & (!g111) & (!i_9_) & (!g14) & (g24)) + ((!sk[107]) & (g111) & (!i_9_) & (g14) & (!g24)) + ((!sk[107]) & (g111) & (!i_9_) & (g14) & (!g24)));
	assign g235 = (((g19) & (!g93) & (!sk[108]) & (i_31_)) + ((g19) & (g93) & (sk[108]) & (!i_31_)));
	assign g236 = (((!sk[109]) & (!i_17_) & (!g29) & (!g119) & (g234) & (!g235)) + ((!sk[109]) & (!i_17_) & (!g29) & (g119) & (g234) & (!g235)) + ((!sk[109]) & (i_17_) & (!g29) & (!g119) & (!g234) & (g235)) + ((sk[109]) & (!i_17_) & (g29) & (g119) & (!g234) & (g235)));
	assign g237 = (((!i_16_) & (!i_21_) & (!g233) & (!sk[110]) & (g236)) + ((i_16_) & (!i_21_) & (g233) & (!sk[110]) & (!g236)) + ((!i_16_) & (!i_21_) & (!g233) & (!sk[110]) & (g236)) + ((!i_16_) & (!i_21_) & (g233) & (sk[110]) & (!g236)));
	assign g238 = (((!i_3_) & (!i_18_) & (!i_11_) & (i_19_) & (!sk[111]) & (!g128)) + ((!i_3_) & (!i_18_) & (!i_11_) & (!i_19_) & (sk[111]) & (!g128)) + ((i_3_) & (!i_18_) & (!i_11_) & (!i_19_) & (!sk[111]) & (g128)) + ((i_3_) & (!i_18_) & (!i_11_) & (!i_19_) & (!sk[111]) & (g128)) + ((!i_3_) & (!i_18_) & (!i_11_) & (!i_19_) & (sk[111]) & (g128)));
	assign g239 = (((!i_31_) & (!g33) & (!sk[112]) & (!i_18_) & (i_19_) & (!g207)) + ((i_31_) & (!g33) & (!sk[112]) & (!i_18_) & (!i_19_) & (g207)) + ((i_31_) & (g33) & (sk[112]) & (!i_18_) & (!i_19_) & (!g207)) + ((i_31_) & (g33) & (!sk[112]) & (!i_18_) & (i_19_) & (!g207)));
	assign g240 = (((!i_24_) & (i_34_) & (!i_35_) & (g3) & (i_21_) & (i_31_)) + ((!i_24_) & (!i_34_) & (i_35_) & (g3) & (i_21_) & (i_31_)));
	assign g241 = (((!sk[114]) & (i_3_) & (!i_11_) & (g128)) + ((!sk[114]) & (i_3_) & (!i_11_) & (g128)));
	assign g242 = (((!g33) & (g238) & (!g239) & (!sk[115]) & (g240) & (!g241)) + ((!g33) & (!g238) & (!g239) & (!sk[115]) & (g240) & (!g241)) + ((!g33) & (!g238) & (g239) & (sk[115]) & (!g240) & (g241)) + ((g33) & (!g238) & (!g239) & (!sk[115]) & (!g240) & (g241)) + ((g33) & (g238) & (g239) & (sk[115]) & (!g240) & (!g241)));
	assign g243 = (((!i_16_) & (!i_17_) & (!sk[116]) & (!i_12_) & (i_13_)) + ((i_16_) & (!i_17_) & (!sk[116]) & (i_12_) & (!i_13_)) + ((!i_16_) & (!i_17_) & (sk[116]) & (!i_12_) & (!i_13_)) + ((!i_16_) & (!i_17_) & (sk[116]) & (!i_12_) & (!i_13_)));
	assign g244 = (((!i_3_) & (!i_11_) & (!sk[117]) & (!g128) & (g242) & (!g243)) + ((i_3_) & (!i_11_) & (!sk[117]) & (!g128) & (!g242) & (g243)) + ((i_3_) & (!i_11_) & (!sk[117]) & (g128) & (g242) & (g243)) + ((!i_3_) & (!i_11_) & (!sk[117]) & (g128) & (g242) & (g243)));
	assign g245 = (((!g22) & (!sk[118]) & (!g229) & (!g231) & (g237) & (!g244)) + ((g22) & (!sk[118]) & (!g229) & (!g231) & (!g237) & (g244)) + ((g22) & (sk[118]) & (!g229) & (!g231) & (!g237) & (!g244)) + ((!g22) & (sk[118]) & (!g229) & (!g231) & (!g237) & (!g244)) + ((g22) & (!sk[118]) & (g229) & (!g231) & (!g237) & (g244)));
	assign o_0_ = (((!i_36_) & (!g117) & (!g186) & (!g216) & (sk[119]) & (!g245)) + ((!i_36_) & (!g117) & (!g186) & (g216) & (!sk[119]) & (!g245)) + ((!i_36_) & (!g117) & (!g186) & (!g216) & (sk[119]) & (!g245)) + ((!i_36_) & (!g117) & (!g186) & (!g216) & (sk[119]) & (!g245)) + ((i_36_) & (!g117) & (!g186) & (!g216) & (!sk[119]) & (g245)) + ((i_36_) & (!g117) & (!g186) & (!g216) & (!sk[119]) & (g245)));
	assign g247 = (((!i_23_) & (!sk[120]) & (!g45) & (!g50) & (g51)) + ((i_23_) & (!sk[120]) & (!g45) & (g50) & (!g51)) + ((!i_23_) & (sk[120]) & (!g45) & (!g50) & (!g51)) + ((i_23_) & (!sk[120]) & (!g45) & (!g50) & (g51)) + ((!i_23_) & (!sk[120]) & (!g45) & (!g50) & (g51)));
	assign g248 = (((i_4_) & (!sk[121]) & (!i_5_) & (i_0_)) + ((!i_4_) & (sk[121]) & (!i_5_) & (!i_0_)));
	assign g249 = (((!g54) & (!sk[122]) & (g24)) + ((g54) & (sk[122]) & (!g24)));
	assign g250 = (((!i_33_) & (!sk[123]) & (!g45) & (!i_10_) & (g249)) + ((i_33_) & (sk[123]) & (!g45) & (!i_10_) & (!g249)) + ((!i_33_) & (sk[123]) & (!g45) & (!i_10_) & (!g249)) + ((!i_33_) & (sk[123]) & (!g45) & (i_10_) & (!g249)) + ((i_33_) & (!sk[123]) & (!g45) & (i_10_) & (!g249)));
	assign g251 = (((!i_17_) & (!i_23_) & (!sk[124]) & (!i_20_) & (i_37_)) + ((i_17_) & (!i_23_) & (!sk[124]) & (i_20_) & (!i_37_)) + ((!i_17_) & (!i_23_) & (!sk[124]) & (!i_20_) & (i_37_)));
	assign g252 = (((!sk[125]) & (!g31) & (!g89) & (!g248) & (g250) & (!g251)) + ((!sk[125]) & (g31) & (!g89) & (!g248) & (!g250) & (g251)) + ((!sk[125]) & (g31) & (g89) & (g248) & (!g250) & (g251)));
	assign g253 = (((!i_17_) & (!i_23_) & (!sk[126]) & (!g88) & (i_20_)) + ((i_17_) & (!i_23_) & (!sk[126]) & (g88) & (!i_20_)) + ((!i_17_) & (!i_23_) & (sk[126]) & (g88) & (!i_20_)));
	assign g254 = (((!i_35_) & (!sk[127]) & (i_37_)) + ((!i_35_) & (!sk[127]) & (i_37_)));
	assign g255 = (((!i_33_) & (!sk[0]) & (!g45) & (!i_10_) & (g254)) + ((i_33_) & (!sk[0]) & (!g45) & (i_10_) & (!g254)) + ((!i_33_) & (!sk[0]) & (g45) & (!i_10_) & (g254)));
	assign g256 = (((!g48) & (!g254) & (!g249) & (!sk[1]) & (g248) & (!g255)) + ((g48) & (!g254) & (!g249) & (!sk[1]) & (!g248) & (g255)) + ((g48) & (g254) & (g249) & (!sk[1]) & (g248) & (!g255)) + ((g48) & (g254) & (!g249) & (!sk[1]) & (g248) & (g255)));
	assign g257 = (((!i_2_) & (!g28) & (g253) & (!sk[2]) & (g256)) + ((!i_2_) & (!g28) & (!g253) & (!sk[2]) & (g256)) + ((i_2_) & (g28) & (g253) & (!sk[2]) & (!g256)) + ((i_2_) & (!g28) & (g253) & (!sk[2]) & (!g256)));
	assign g258 = (((!i_23_) & (!i_21_) & (!g88) & (!sk[3]) & (i_22_) & (!g157)) + ((i_23_) & (!i_21_) & (!g88) & (!sk[3]) & (!i_22_) & (g157)) + ((!i_23_) & (i_21_) & (g88) & (sk[3]) & (!i_22_) & (g157)));
	assign g259 = (((!sk[4]) & (!i_33_) & (!i_13_) & (!i_14_) & (g254)) + ((!sk[4]) & (!i_33_) & (!i_13_) & (!i_14_) & (g254)) + ((!sk[4]) & (i_33_) & (!i_13_) & (i_14_) & (!g254)) + ((!sk[4]) & (!i_33_) & (!i_13_) & (!i_14_) & (g254)));
	assign g260 = (((!i_16_) & (!i_23_) & (!sk[5]) & (!i_20_) & (g259)) + ((i_16_) & (!i_23_) & (!sk[5]) & (i_20_) & (!g259)) + ((!i_16_) & (!i_23_) & (!sk[5]) & (!i_20_) & (g259)));
	assign g261 = (((!sk[6]) & (!i_17_) & (!i_12_) & (!i_23_) & (i_20_) & (!i_0_)) + ((!sk[6]) & (i_17_) & (!i_12_) & (!i_23_) & (!i_20_) & (i_0_)) + ((sk[6]) & (!i_17_) & (!i_12_) & (!i_23_) & (!i_20_) & (!i_0_)) + ((sk[6]) & (!i_17_) & (!i_12_) & (!i_23_) & (!i_20_) & (!i_0_)));
	assign g262 = (((!i_28_) & (!g70) & (!g258) & (!sk[7]) & (g260) & (!g261)) + ((!i_28_) & (!g70) & (!g258) & (sk[7]) & (!g260) & (!g261)) + ((i_28_) & (!g70) & (!g258) & (!sk[7]) & (!g260) & (g261)) + ((i_28_) & (!g70) & (!g258) & (!sk[7]) & (g260) & (!g261)) + ((!i_28_) & (g70) & (!g258) & (!sk[7]) & (g260) & (!g261)) + ((!i_28_) & (!g70) & (!g258) & (!sk[7]) & (g260) & (!g261)));
	assign g263 = (((!sk[8]) & (g14) & (!i_1_) & (i_0_)) + ((sk[8]) & (g14) & (!i_1_) & (!i_0_)));
	assign g264 = (((!i_7_) & (!sk[9]) & (!i_8_) & (!i_37_) & (g263) & (!g253)) + ((i_7_) & (!sk[9]) & (!i_8_) & (!i_37_) & (!g263) & (g253)) + ((!i_7_) & (!sk[9]) & (!i_8_) & (i_37_) & (g263) & (g253)));
	assign g265 = (((!i_33_) & (!g45) & (!sk[10]) & (!g54) & (g264)) + ((!i_33_) & (!g45) & (!sk[10]) & (g54) & (g264)) + ((i_33_) & (!g45) & (!sk[10]) & (g54) & (!g264)) + ((!i_33_) & (g45) & (!sk[10]) & (!g54) & (g264)));
	assign g266 = (((!i_33_) & (!i_13_) & (!i_14_) & (g37) & (g58) & (g254)) + ((!i_33_) & (!i_13_) & (!i_14_) & (g37) & (g58) & (g254)));
	assign g267 = (((!i_33_) & (!i_17_) & (!sk[12]) & (!g28) & (g54) & (!g254)) + ((i_33_) & (!i_17_) & (!sk[12]) & (!g28) & (!g54) & (g254)) + ((!i_33_) & (!i_17_) & (!sk[12]) & (g28) & (g54) & (g254)) + ((!i_33_) & (!i_17_) & (sk[12]) & (g28) & (!g54) & (g254)));
	assign g268 = (((!i_23_) & (!i_9_) & (!g89) & (i_20_) & (!sk[13]) & (!g267)) + ((i_23_) & (!i_9_) & (!g89) & (!i_20_) & (!sk[13]) & (g267)) + ((!i_23_) & (!i_9_) & (g89) & (!i_20_) & (sk[13]) & (g267)));
	assign g269 = (((!sk[14]) & (!i_3_) & (!i_18_) & (!g14) & (i_0_)) + ((!sk[14]) & (i_3_) & (!i_18_) & (g14) & (!i_0_)) + ((!sk[14]) & (i_3_) & (!i_18_) & (g14) & (!i_0_)));
	assign g270 = (((!i_6_) & (!sk[15]) & (!g12) & (!g248) & (g268) & (!g269)) + ((!i_6_) & (!sk[15]) & (!g12) & (!g248) & (g268) & (g269)) + ((i_6_) & (!sk[15]) & (!g12) & (!g248) & (!g268) & (g269)) + ((!i_6_) & (!sk[15]) & (g12) & (g248) & (g268) & (!g269)));
	assign g271 = (((!g257) & (!g262) & (!g265) & (!sk[16]) & (g266) & (!g270)) + ((g257) & (!g262) & (!g265) & (!sk[16]) & (!g266) & (g270)) + ((!g257) & (g262) & (!g265) & (sk[16]) & (!g266) & (!g270)));
	assign g272 = (((i_33_) & (!sk[17]) & (!g1) & (g254)) + ((!i_33_) & (sk[17]) & (g1) & (g254)));
	assign g273 = (((!sk[18]) & (!g13) & (!g107) & (!g47) & (g49) & (!g51)) + ((sk[18]) & (!g13) & (g107) & (g47) & (!g49) & (!g51)) + ((!sk[18]) & (g13) & (g107) & (!g47) & (g49) & (!g51)) + ((!sk[18]) & (g13) & (!g107) & (!g47) & (!g49) & (g51)) + ((sk[18]) & (!g13) & (g107) & (!g47) & (!g49) & (g51)));
	assign g274 = (((!i_12_) & (!i_6_) & (!sk[19]) & (!g248) & (g260)) + ((i_12_) & (!i_6_) & (!sk[19]) & (g248) & (!g260)) + ((!i_12_) & (!i_6_) & (!sk[19]) & (g248) & (g260)));
	assign g275 = (((!sk[20]) & (!g1) & (!g89) & (!g254) & (g273) & (!g274)) + ((!sk[20]) & (g1) & (!g89) & (g254) & (g273) & (!g274)) + ((!sk[20]) & (g1) & (!g89) & (!g254) & (!g273) & (g274)) + ((sk[20]) & (!g1) & (g89) & (!g254) & (!g273) & (g274)));
	assign g276 = (((!g247) & (!g252) & (!sk[21]) & (!g271) & (g272) & (!g275)) + ((g247) & (!g252) & (!sk[21]) & (!g271) & (!g272) & (g275)) + ((!g247) & (!g252) & (sk[21]) & (g271) & (!g272) & (!g275)) + ((g247) & (!g252) & (!sk[21]) & (g271) & (g272) & (!g275)));
	assign g277 = (((!sk[22]) & (i_33_) & (!i_34_) & (i_32_)) + ((sk[22]) & (!i_33_) & (i_34_) & (!i_32_)));
	assign g278 = (((!i_16_) & (!i_13_) & (!sk[23]) & (!g33) & (g9) & (!g69)) + ((i_16_) & (!i_13_) & (!sk[23]) & (!g33) & (!g9) & (g69)) + ((!i_16_) & (!i_13_) & (sk[23]) & (!g33) & (!g9) & (!g69)) + ((i_16_) & (!i_13_) & (!sk[23]) & (!g33) & (g9) & (!g69)) + ((!i_16_) & (i_13_) & (!sk[23]) & (!g33) & (g9) & (!g69)) + ((!i_16_) & (!i_13_) & (!sk[23]) & (!g33) & (g9) & (!g69)));
	assign g279 = (((!sk[24]) & (i_33_) & (!g2) & (i_37_)) + ((sk[24]) & (!i_33_) & (g2) & (i_37_)));
	assign g280 = (((!i_16_) & (!i_17_) & (!i_12_) & (!i_13_) & (!i_23_) & (g7)) + ((!i_16_) & (!i_17_) & (!i_12_) & (!i_13_) & (!i_23_) & (g7)));
	assign g281 = (((!i_16_) & (!sk[26]) & (!i_34_) & (!i_12_) & (i_13_) & (!g33)) + ((i_16_) & (!sk[26]) & (!i_34_) & (!i_12_) & (!i_13_) & (g33)) + ((!i_16_) & (sk[26]) & (i_34_) & (!i_12_) & (!i_13_) & (g33)));
	assign g282 = (((!i_33_) & (!i_8_) & (!g254) & (!sk[27]) & (g281)) + ((i_33_) & (!i_8_) & (g254) & (!sk[27]) & (!g281)) + ((!i_33_) & (!i_8_) & (g254) & (!sk[27]) & (g281)));
	assign g283 = (((!i_30_) & (!g279) & (!g280) & (!sk[28]) & (g282)) + ((!i_30_) & (!g279) & (!g280) & (!sk[28]) & (g282)) + ((i_30_) & (!g279) & (g280) & (!sk[28]) & (!g282)) + ((!i_30_) & (g279) & (g280) & (sk[28]) & (!g282)));
	assign g284 = (((!sk[29]) & (!g93) & (!g53) & (!g10) & (i_10_) & (!i_37_)) + ((!sk[29]) & (g93) & (!g53) & (!g10) & (!i_10_) & (i_37_)) + ((!sk[29]) & (g93) & (g53) & (g10) & (!i_10_) & (i_37_)));
	assign g285 = (((!i_13_) & (!i_10_) & (!sk[30]) & (!g11) & (g23)) + ((i_13_) & (!i_10_) & (!sk[30]) & (g11) & (!g23)) + ((!i_13_) & (!i_10_) & (!sk[30]) & (g11) & (g23)));
	assign g286 = (((!sk[31]) & (i_33_) & (!i_32_) & (i_37_)) + ((sk[31]) & (!i_33_) & (!i_32_) & (i_37_)));
	assign g287 = (((!g93) & (!i_30_) & (!i_31_) & (!sk[32]) & (g150) & (!g286)) + ((g93) & (!i_30_) & (!i_31_) & (!sk[32]) & (!g150) & (g286)) + ((g93) & (!i_30_) & (i_31_) & (!sk[32]) & (g150) & (g286)));
	assign g288 = (((!sk[33]) & (!i_33_) & (!g93) & (!g55) & (g254)) + ((!sk[33]) & (i_33_) & (!g93) & (g55) & (!g254)) + ((!sk[33]) & (!i_33_) & (g93) & (!g55) & (g254)) + ((!sk[33]) & (!i_33_) & (g93) & (g55) & (g254)));
	assign g289 = (((!g61) & (!g279) & (!g285) & (g287) & (!sk[34]) & (!g288)) + ((g61) & (!g279) & (!g285) & (!g287) & (!sk[34]) & (g288)) + ((!g61) & (!g279) & (!g285) & (!g287) & (sk[34]) & (!g288)) + ((!g61) & (!g279) & (!g285) & (!g287) & (sk[34]) & (!g288)) + ((!g61) & (!g279) & (!g285) & (!g287) & (sk[34]) & (!g288)) + ((!g61) & (!g279) & (!g285) & (!g287) & (sk[34]) & (!g288)));
	assign g290 = (((!i_33_) & (!g65) & (!g283) & (!sk[35]) & (g284) & (!g289)) + ((i_33_) & (!g65) & (!g283) & (!sk[35]) & (!g284) & (g289)) + ((i_33_) & (!g65) & (!g283) & (!sk[35]) & (!g284) & (g289)) + ((!i_33_) & (!g65) & (!g283) & (sk[35]) & (!g284) & (g289)) + ((!i_33_) & (!g65) & (!g283) & (!sk[35]) & (g284) & (g289)));
	assign g291 = (((i_32_) & (!sk[36]) & (!g79) & (g279)) + ((!i_32_) & (sk[36]) & (g79) & (g279)));
	assign g292 = (((!g254) & (!g277) & (!sk[37]) & (!g278) & (g290) & (!g291)) + ((g254) & (!g277) & (!sk[37]) & (!g278) & (!g290) & (g291)) + ((!g254) & (!g277) & (!sk[37]) & (!g278) & (g290) & (!g291)) + ((!g254) & (!g277) & (!sk[37]) & (!g278) & (g290) & (!g291)) + ((!g254) & (!g277) & (!sk[37]) & (g278) & (g290) & (!g291)));
	assign g293 = (((!i_27_) & (!g71) & (!g1) & (g276) & (!sk[38]) & (!g292)) + ((i_27_) & (!g71) & (!g1) & (!g276) & (!sk[38]) & (g292)) + ((!i_27_) & (!g71) & (!g1) & (!g276) & (sk[38]) & (!g292)) + ((!i_27_) & (!g71) & (g1) & (!g276) & (sk[38]) & (!g292)));
	assign g294 = (((!sk[39]) & (!i_7_) & (g29)) + ((!sk[39]) & (!i_7_) & (g29)));
	assign g295 = (((g32) & (!sk[40]) & (g249)) + ((!g32) & (!sk[40]) & (g249)));
	assign g296 = (((!sk[41]) & (g45) & (!i_8_) & (g294)) + ((!sk[41]) & (g45) & (!i_8_) & (g294)));
	assign g297 = (((!i_33_) & (!g2) & (!sk[42]) & (!i_32_) & (g1) & (!i_37_)) + ((i_33_) & (!g2) & (!sk[42]) & (!i_32_) & (!g1) & (i_37_)) + ((!i_33_) & (g2) & (!sk[42]) & (!i_32_) & (g1) & (i_37_)) + ((!i_33_) & (g2) & (!sk[42]) & (!i_32_) & (g1) & (i_37_)));
	assign g298 = (((!i_33_) & (!g37) & (!g295) & (!sk[43]) & (g296) & (!g297)) + ((i_33_) & (!g37) & (!g295) & (!sk[43]) & (!g296) & (g297)) + ((!i_33_) & (!g37) & (!g295) & (!sk[43]) & (g296) & (g297)) + ((!i_33_) & (!g37) & (g295) & (!sk[43]) & (g296) & (g297)) + ((!i_33_) & (g37) & (g295) & (sk[43]) & (!g296) & (g297)));
	assign g299 = (((!g2) & (!g1) & (!sk[44]) & (!g54) & (i_37_)) + ((g2) & (!g1) & (!sk[44]) & (g54) & (!i_37_)) + ((g2) & (g1) & (!sk[44]) & (g54) & (i_37_)));
	assign g300 = (((!i_8_) & (!sk[45]) & (!g294) & (!g38) & (g298) & (!g299)) + ((!i_8_) & (!sk[45]) & (!g294) & (g38) & (g298) & (!g299)) + ((i_8_) & (!sk[45]) & (!g294) & (!g38) & (!g298) & (g299)) + ((!i_8_) & (sk[45]) & (g294) & (g38) & (!g298) & (g299)));
	assign g301 = (((!i_33_) & (!i_17_) & (!g45) & (!sk[46]) & (i_8_) & (!g294)) + ((i_33_) & (!i_17_) & (!g45) & (!sk[46]) & (!i_8_) & (g294)) + ((!i_33_) & (!i_17_) & (g45) & (sk[46]) & (!i_8_) & (g294)) + ((!i_33_) & (!i_17_) & (g45) & (!sk[46]) & (i_8_) & (g294)));
	assign g302 = (((!g53) & (!g42) & (!g35) & (!sk[47]) & (g296) & (!g301)) + ((g53) & (g42) & (!g35) & (!sk[47]) & (!g296) & (g301)) + ((g53) & (!g42) & (!g35) & (!sk[47]) & (!g296) & (g301)) + ((!g53) & (!g42) & (g35) & (!sk[47]) & (g296) & (g301)) + ((!g53) & (g42) & (g35) & (sk[47]) & (!g296) & (g301)));
	assign g303 = (((!sk[48]) & (!i_8_) & (!g294) & (!g42) & (g55) & (!g35)) + ((!sk[48]) & (!i_8_) & (g294) & (g42) & (g55) & (!g35)) + ((!sk[48]) & (i_8_) & (!g294) & (!g42) & (!g55) & (g35)) + ((!sk[48]) & (!i_8_) & (g294) & (!g42) & (g55) & (g35)));
	assign g304 = (((!sk[49]) & (!i_33_) & (!i_7_) & (!g57) & (g33) & (!g84)) + ((!sk[49]) & (i_33_) & (!i_7_) & (!g57) & (!g33) & (g84)) + ((!sk[49]) & (!i_33_) & (!i_7_) & (g57) & (g33) & (g84)));
	assign g305 = (((!sk[50]) & (!i_33_) & (!i_30_) & (!g21) & (g304) & (!g280)) + ((sk[50]) & (!i_33_) & (i_30_) & (!g21) & (!g304) & (!g280)) + ((sk[50]) & (!i_33_) & (!i_30_) & (!g21) & (!g304) & (!g280)) + ((sk[50]) & (!i_33_) & (!i_30_) & (!g21) & (!g304) & (!g280)) + ((!sk[50]) & (i_33_) & (!i_30_) & (!g21) & (!g304) & (g280)));
	assign g306 = (((!sk[51]) & (!i_34_) & (!i_37_) & (!g302) & (g303) & (!g305)) + ((!sk[51]) & (i_34_) & (i_37_) & (!g302) & (g303) & (!g305)) + ((!sk[51]) & (i_34_) & (!i_37_) & (!g302) & (!g303) & (g305)) + ((sk[51]) & (i_34_) & (i_37_) & (!g302) & (!g303) & (!g305)) + ((!sk[51]) & (i_34_) & (i_37_) & (g302) & (!g303) & (g305)));
	assign g307 = (((!g142) & (!i_25_) & (!g144) & (!sk[52]) & (i_20_)) + ((!g142) & (i_25_) & (g144) & (sk[52]) & (!i_20_)) + ((g142) & (!i_25_) & (g144) & (!sk[52]) & (!i_20_)) + ((!g142) & (i_25_) & (!g144) & (!sk[52]) & (i_20_)));
	assign g308 = (((!i_13_) & (!sk[53]) & (!g10) & (!i_10_) & (g55)) + ((i_13_) & (!sk[53]) & (!g10) & (i_10_) & (!g55)) + ((i_13_) & (!sk[53]) & (g10) & (!i_10_) & (g55)) + ((!i_13_) & (!sk[53]) & (g10) & (!i_10_) & (g55)));
	assign g309 = (((i_34_) & (g42) & (!g21) & (g254) & (g308) & (!g273)) + ((i_34_) & (!g42) & (g21) & (g254) & (!g308) & (g273)));
	assign g310 = (((!i_24_) & (!i_34_) & (!sk[55]) & (!i_35_) & (g34) & (!i_37_)) + ((i_24_) & (!i_34_) & (!sk[55]) & (!i_35_) & (!g34) & (i_37_)) + ((!i_24_) & (i_34_) & (!sk[55]) & (!i_35_) & (g34) & (i_37_)) + ((!i_24_) & (!i_34_) & (!sk[55]) & (i_35_) & (g34) & (i_37_)));
	assign g311 = (((!i_34_) & (!i_29_) & (!sk[56]) & (!g34) & (g101) & (!g254)) + ((i_34_) & (!i_29_) & (!sk[56]) & (!g34) & (!g101) & (g254)) + ((i_34_) & (!i_29_) & (!sk[56]) & (g34) & (!g101) & (g254)) + ((!i_34_) & (!i_29_) & (!sk[56]) & (!g34) & (g101) & (g254)));
	assign g312 = (((!i_16_) & (!i_17_) & (!i_12_) & (!i_14_) & (g33) & (!i_8_)) + ((!i_16_) & (!i_17_) & (!i_12_) & (!i_14_) & (g33) & (!i_8_)));
	assign g313 = (((!sk[58]) & (i_12_) & (!g7) & (g107)) + ((sk[58]) & (!i_12_) & (g7) & (g107)));
	assign g314 = (((!sk[59]) & (!i_30_) & (!g310) & (!g311) & (g312) & (!g313)) + ((!sk[59]) & (!i_30_) & (!g310) & (g311) & (g312) & (!g313)) + ((!sk[59]) & (i_30_) & (!g310) & (!g311) & (!g312) & (g313)) + ((sk[59]) & (!i_30_) & (g310) & (!g311) & (!g312) & (g313)));
	assign g315 = (((!sk[60]) & (!i_32_) & (!i_29_) & (!g101) & (g254)) + ((!sk[60]) & (i_32_) & (!i_29_) & (g101) & (!g254)) + ((!sk[60]) & (!i_32_) & (!i_29_) & (g101) & (g254)));
	assign g316 = (((!g66) & (!g34) & (!i_37_) & (!sk[61]) & (g315)) + ((g66) & (!g34) & (i_37_) & (!sk[61]) & (!g315)) + ((!g66) & (!g34) & (!i_37_) & (sk[61]) & (!g315)) + ((!g66) & (!g34) & (!i_37_) & (sk[61]) & (!g315)) + ((g66) & (!g34) & (i_37_) & (!sk[61]) & (!g315)));
	assign g317 = (((!i_16_) & (!sk[62]) & (!i_14_) & (!g33) & (g9)) + ((i_16_) & (!sk[62]) & (!i_14_) & (g33) & (!g9)) + ((!i_16_) & (!sk[62]) & (!i_14_) & (g33) & (g9)));
	assign g318 = (((!g68) & (!sk[63]) & (!g55) & (!g314) & (g316) & (!g317)) + ((!g68) & (!sk[63]) & (!g55) & (!g314) & (g316) & (!g317)) + ((g68) & (!sk[63]) & (!g55) & (!g314) & (!g316) & (g317)) + ((!g68) & (sk[63]) & (!g55) & (!g314) & (!g316) & (!g317)) + ((!g68) & (sk[63]) & (!g55) & (!g314) & (!g316) & (!g317)));
	assign g319 = (((!g300) & (!g306) & (!g307) & (!sk[64]) & (g309) & (!g318)) + ((g300) & (!g306) & (!g307) & (!sk[64]) & (!g309) & (g318)) + ((!g300) & (!g306) & (!g307) & (sk[64]) & (!g309) & (g318)));
	assign g320 = (((!sk[65]) & (!i_33_) & (!i_17_) & (!i_12_) & (g45) & (!g54)) + ((!sk[65]) & (!i_33_) & (!i_17_) & (!i_12_) & (g45) & (!g54)) + ((!sk[65]) & (!i_33_) & (!i_17_) & (!i_12_) & (g45) & (!g54)) + ((!sk[65]) & (i_33_) & (!i_17_) & (!i_12_) & (!g45) & (g54)) + ((sk[65]) & (!i_33_) & (!i_17_) & (!i_12_) & (!g45) & (g54)) + ((sk[65]) & (!i_33_) & (!i_17_) & (!i_12_) & (!g45) & (g54)));
	assign g321 = (((!sk[66]) & (!i_31_) & (!g84) & (!g5) & (g320)) + ((!sk[66]) & (i_31_) & (!g84) & (g5) & (!g320)) + ((!sk[66]) & (i_31_) & (g84) & (!g5) & (g320)));
	assign g322 = (((i_34_) & (!g35) & (!g295) & (!sk[67]) & (g321)) + ((!i_34_) & (!g35) & (!g295) & (!sk[67]) & (g321)) + ((i_34_) & (g35) & (g295) & (!sk[67]) & (!g321)) + ((i_34_) & (!g35) & (g295) & (!sk[67]) & (!g321)));
	assign g323 = (((i_16_) & (!sk[68]) & (!i_17_) & (i_20_)) + ((!i_16_) & (sk[68]) & (!i_17_) & (!i_20_)));
	assign g324 = (((!g19) & (!i_14_) & (!sk[69]) & (!i_7_) & (i_0_) & (!g323)) + ((g19) & (!i_14_) & (!sk[69]) & (!i_7_) & (!i_0_) & (g323)) + ((g19) & (!i_14_) & (!sk[69]) & (!i_7_) & (!i_0_) & (g323)));
	assign g325 = (((!i_31_) & (!sk[70]) & (!g34) & (!g134) & (g324)) + ((i_31_) & (!sk[70]) & (!g34) & (g134) & (!g324)) + ((!i_31_) & (sk[70]) & (!g34) & (!g134) & (!g324)) + ((!i_31_) & (sk[70]) & (!g34) & (!g134) & (!g324)) + ((i_31_) & (!sk[70]) & (!g34) & (g134) & (!g324)));
	assign g326 = (((!sk[71]) & (!g111) & (!g13) & (!g31) & (i_20_) & (!g248)) + ((!sk[71]) & (g111) & (!g13) & (!g31) & (!i_20_) & (g248)) + ((!sk[71]) & (g111) & (g13) & (g31) & (!i_20_) & (g248)));
	assign g327 = (((g111) & (!g190) & (!sk[72]) & (i_20_)) + ((g111) & (g190) & (sk[72]) & (!i_20_)));
	assign g328 = (((i_7_) & (!i_0_) & (!sk[73]) & (g327)) + ((!i_7_) & (!i_0_) & (sk[73]) & (g327)));
	assign g329 = (((!i_12_) & (!i_7_) & (!g130) & (i_6_) & (!sk[74]) & (!g248)) + ((i_12_) & (!i_7_) & (!g130) & (!i_6_) & (!sk[74]) & (g248)) + ((!i_12_) & (!i_7_) & (g130) & (!i_6_) & (sk[74]) & (g248)));
	assign g330 = (((!g19) & (!i_12_) & (!i_30_) & (i_7_) & (!sk[75]) & (!i_0_)) + ((g19) & (!i_12_) & (!i_30_) & (!i_7_) & (!sk[75]) & (i_0_)) + ((g19) & (!i_12_) & (!i_30_) & (!i_7_) & (sk[75]) & (!i_0_)));
	assign g331 = (((!sk[76]) & (!g93) & (!i_20_) & (!g329) & (g330)) + ((!sk[76]) & (g93) & (!i_20_) & (g329) & (!g330)) + ((!sk[76]) & (g93) & (!i_20_) & (g329) & (!g330)) + ((!sk[76]) & (g93) & (!i_20_) & (!g329) & (g330)));
	assign g332 = (((g54) & (!sk[77]) & (!g326) & (g328) & (!g331)) + ((g54) & (!sk[77]) & (!g326) & (!g328) & (g331)) + ((!g54) & (!sk[77]) & (!g326) & (!g328) & (g331)) + ((g54) & (sk[77]) & (g326) & (!g328) & (!g331)));
	assign g333 = (((!g93) & (!i_30_) & (!sk[78]) & (!g325) & (g332)) + ((!g93) & (!i_30_) & (sk[78]) & (!g325) & (!g332)) + ((!g93) & (i_30_) & (sk[78]) & (!g325) & (!g332)) + ((g93) & (!i_30_) & (!sk[78]) & (g325) & (!g332)));
	assign g334 = (((!i_29_) & (!sk[79]) & (i_20_)) + ((i_29_) & (sk[79]) & (!i_20_)));
	assign g335 = (((!i_9_) & (!sk[80]) & (i_6_)) + ((!i_9_) & (sk[80]) & (!i_6_)));
	assign g336 = (((g335) & (!sk[81]) & (!i_10_) & (g248)) + ((g335) & (!sk[81]) & (!i_10_) & (g248)));
	assign g337 = (((!i_33_) & (!sk[82]) & (!g53) & (!g254) & (g336)) + ((i_33_) & (!sk[82]) & (!g53) & (g254) & (!g336)) + ((!i_33_) & (!sk[82]) & (g53) & (g254) & (g336)));
	assign g338 = (((!g335) & (!g24) & (!sk[83]) & (!g254) & (g248)) + ((g335) & (!g24) & (!sk[83]) & (g254) & (!g248)) + ((g335) & (!g24) & (!sk[83]) & (g254) & (g248)));
	assign g339 = (((!i_7_) & (!i_37_) & (!sk[84]) & (!g263) & (g338)) + ((!i_7_) & (!i_37_) & (sk[84]) & (!g263) & (!g338)) + ((!i_7_) & (!i_37_) & (sk[84]) & (!g263) & (!g338)) + ((i_7_) & (!i_37_) & (!sk[84]) & (g263) & (!g338)));
	assign g340 = (((g33) & (g101) & (!g55) & (g334) & (g337) & (!g339)) + ((g33) & (g101) & (g55) & (g334) & (!g337) & (!g339)));
	assign g341 = (((!g2) & (!i_7_) & (!g29) & (!sk[86]) & (i_37_)) + ((g2) & (!i_7_) & (g29) & (!sk[86]) & (!i_37_)) + ((g2) & (!i_7_) & (g29) & (!sk[86]) & (i_37_)));
	assign g342 = (((!g3) & (!i_29_) & (!g55) & (!sk[87]) & (g341)) + ((g3) & (!i_29_) & (g55) & (!sk[87]) & (!g341)) + ((g3) & (!i_29_) & (g55) & (!sk[87]) & (g341)));
	assign g343 = (((!i_14_) & (!g111) & (!sk[88]) & (!g254) & (g263) & (!g323)) + ((i_14_) & (!g111) & (!sk[88]) & (!g254) & (!g263) & (g323)) + ((!i_14_) & (g111) & (!sk[88]) & (g254) & (g263) & (g323)));
	assign g344 = (((!i_14_) & (i_21_) & (!g84) & (g88) & (g223) & (!g254)) + ((!i_14_) & (i_21_) & (!g84) & (!g88) & (g223) & (g254)) + ((!i_14_) & (!i_21_) & (g84) & (!g88) & (g223) & (g254)));
	assign g345 = (((!i_34_) & (!sk[90]) & (!g71) & (!g342) & (g343) & (!g344)) + ((i_34_) & (!sk[90]) & (!g71) & (!g342) & (!g343) & (g344)) + ((!i_34_) & (sk[90]) & (g71) & (!g342) & (!g343) & (!g344)) + ((!i_34_) & (sk[90]) & (!g71) & (!g342) & (!g343) & (!g344)) + ((i_34_) & (!sk[90]) & (!g71) & (!g342) & (!g343) & (g344)));
	assign g346 = (((!g100) & (!sk[91]) & (!g254) & (!g308) & (g340) & (!g345)) + ((g100) & (!sk[91]) & (!g254) & (!g308) & (!g340) & (g345)) + ((!g100) & (sk[91]) & (!g254) & (!g308) & (!g340) & (g345)) + ((!g100) & (sk[91]) & (!g254) & (!g308) & (!g340) & (g345)) + ((!g100) & (sk[91]) & (!g254) & (!g308) & (!g340) & (g345)));
	assign g347 = (((!g53) & (!g10) & (!sk[92]) & (!i_10_) & (g42)) + ((g53) & (!g10) & (!sk[92]) & (i_10_) & (!g42)) + ((g53) & (g10) & (!sk[92]) & (!i_10_) & (g42)));
	assign g348 = (((!g45) & (!sk[93]) & (!i_10_) & (!g49) & (g35)) + ((g45) & (!sk[93]) & (!i_10_) & (g49) & (!g35)) + ((g45) & (!sk[93]) & (!i_10_) & (g49) & (g35)));
	assign g349 = (((!i_33_) & (!sk[94]) & (!i_34_) & (!i_35_) & (g347) & (!g348)) + ((i_33_) & (!sk[94]) & (!i_34_) & (!i_35_) & (!g347) & (g348)) + ((!i_33_) & (!sk[94]) & (i_34_) & (!i_35_) & (g347) & (!g348)) + ((!i_33_) & (sk[94]) & (i_34_) & (!i_35_) & (!g347) & (g348)));
	assign g350 = (((g77) & (!sk[95]) & (!g16) & (!g78) & (g107)) + ((!g77) & (!sk[95]) & (!g16) & (!g78) & (g107)) + ((!g77) & (!sk[95]) & (g16) & (!g78) & (g107)) + ((!g77) & (!sk[95]) & (!g16) & (g78) & (g107)) + ((g77) & (!sk[95]) & (!g16) & (g78) & (!g107)));
	assign g351 = (((!g197) & (!sk[96]) & (!i_20_) & (!i_0_) & (g320)) + ((g197) & (!sk[96]) & (!i_20_) & (i_0_) & (!g320)) + ((g197) & (!sk[96]) & (!i_20_) & (!i_0_) & (g320)));
	assign g352 = (((!sk[97]) & (!i_33_) & (!i_34_) & (!g21) & (g285)) + ((!sk[97]) & (i_33_) & (!i_34_) & (g21) & (!g285)) + ((!sk[97]) & (!i_33_) & (i_34_) & (g21) & (g285)));
	assign g353 = (((!sk[98]) & (!i_33_) & (!g2) & (!g37) & (g38)) + ((!sk[98]) & (i_33_) & (!g2) & (g37) & (!g38)) + ((!sk[98]) & (!i_33_) & (g2) & (g37) & (g38)));
	assign g354 = (((g45) & (!i_10_) & (g32) & (!g35) & (!g277) & (g353)) + ((g45) & (!i_10_) & (g32) & (g35) & (g277) & (!g353)));
	assign g355 = (((!g33) & (!g101) & (!g351) & (!sk[100]) & (g352) & (!g354)) + ((g33) & (!g101) & (!g351) & (!sk[100]) & (!g352) & (g354)) + ((!g33) & (!g101) & (!g351) & (sk[100]) & (!g352) & (!g354)) + ((!g33) & (!g101) & (!g351) & (sk[100]) & (!g352) & (!g354)) + ((!g33) & (!g101) & (!g351) & (sk[100]) & (!g352) & (!g354)));
	assign g356 = (((!g76) & (!g110) & (!sk[101]) & (!g349) & (g350) & (!g355)) + ((g76) & (!g110) & (!sk[101]) & (!g349) & (!g350) & (g355)) + ((!g76) & (!g110) & (sk[101]) & (!g349) & (!g350) & (g355)) + ((!g76) & (!g110) & (sk[101]) & (!g349) & (!g350) & (g355)));
	assign g357 = (((!i_32_) & (!i_37_) & (!g322) & (!g333) & (!g346) & (!g356)) + ((!i_32_) & (i_37_) & (!g322) & (!g333) & (!g346) & (!g356)) + ((!i_32_) & (i_37_) & (g322) & (!g333) & (!g346) & (!g356)) + ((!i_32_) & (i_37_) & (!g322) & (!g333) & (!g346) & (!g356)));
	assign g358 = (((g23) & (!sk[103]) & (g310)) + ((!g23) & (!sk[103]) & (g310)));
	assign g359 = (((!g7) & (!g335) & (!sk[104]) & (!g248) & (g323)) + ((g7) & (!g335) & (!sk[104]) & (g248) & (!g323)) + ((g7) & (g335) & (!sk[104]) & (g248) & (g323)));
	assign g360 = (((!g2) & (!i_7_) & (!sk[105]) & (!i_32_) & (g97)) + ((g2) & (!i_7_) & (!sk[105]) & (i_32_) & (!g97)) + ((g2) & (!i_7_) & (!sk[105]) & (!i_32_) & (g97)));
	assign g361 = (((!g111) & (!g24) & (!sk[106]) & (!g359) & (g360)) + ((g111) & (!g24) & (!sk[106]) & (g359) & (!g360)) + ((!g111) & (!g24) & (sk[106]) & (!g359) & (!g360)) + ((!g111) & (!g24) & (sk[106]) & (!g359) & (!g360)) + ((g111) & (g24) & (!sk[106]) & (g359) & (!g360)));
	assign g362 = (((!g6) & (!sk[107]) & (!g17) & (!i_37_) & (g361)) + ((!g6) & (sk[107]) & (!g17) & (i_37_) & (!g361)) + ((g6) & (!sk[107]) & (!g17) & (i_37_) & (!g361)) + ((!g6) & (!sk[107]) & (g17) & (i_37_) & (g361)));
	assign g363 = (((!sk[108]) & (i_10_) & (!g11) & (g197)) + ((sk[108]) & (i_10_) & (!g11) & (!g197)) + ((sk[108]) & (!i_10_) & (!g11) & (!g197)));
	assign g364 = (((!i_24_) & (!i_34_) & (!i_23_) & (g1) & (!sk[109]) & (!i_37_)) + ((i_24_) & (!i_34_) & (!i_23_) & (!g1) & (!sk[109]) & (i_37_)) + ((!i_24_) & (i_34_) & (!i_23_) & (g1) & (!sk[109]) & (i_37_)));
	assign g365 = (((!i_7_) & (!sk[110]) & (!g85) & (!g86) & (g254) & (!g364)) + ((!i_7_) & (!sk[110]) & (g85) & (!g86) & (g254) & (!g364)) + ((i_7_) & (!sk[110]) & (!g85) & (!g86) & (!g254) & (g364)) + ((!i_7_) & (sk[110]) & (!g85) & (!g86) & (!g254) & (g364)));
	assign g366 = (((!i_14_) & (!sk[111]) & (!g358) & (!g362) & (g363) & (!g365)) + ((!i_14_) & (sk[111]) & (!g358) & (g362) & (!g363) & (!g365)) + ((!i_14_) & (sk[111]) & (!g358) & (!g362) & (!g363) & (g365)) + ((i_14_) & (!sk[111]) & (!g358) & (!g362) & (!g363) & (g365)) + ((!i_14_) & (sk[111]) & (g358) & (!g362) & (!g363) & (!g365)));
	assign g367 = (((!sk[112]) & (i_33_) & (!i_32_) & (i_29_)) + ((sk[112]) & (!i_33_) & (!i_32_) & (!i_29_)));
	assign g368 = (((!sk[113]) & (!i_24_) & (!i_23_) & (!i_30_) & (i_8_)) + ((!sk[113]) & (i_24_) & (!i_23_) & (i_30_) & (!i_8_)) + ((sk[113]) & (!i_24_) & (!i_23_) & (!i_30_) & (!i_8_)));
	assign g369 = (((!sk[114]) & (!i_33_) & (!i_29_) & (!g243) & (g368)) + ((!sk[114]) & (i_33_) & (!i_29_) & (g243) & (!g368)) + ((!sk[114]) & (!i_33_) & (!i_29_) & (g243) & (g368)));
	assign g370 = (((!sk[115]) & (g254) & (!g367) & (g369) & (!g278)) + ((!sk[115]) & (!g254) & (!g367) & (!g369) & (g278)) + ((sk[115]) & (g254) & (g367) & (!g369) & (!g278)));
	assign g371 = (((i_3_) & (!i_18_) & (!sk[116]) & (g12)) + ((!i_3_) & (!i_18_) & (sk[116]) & (!g12)) + ((!i_3_) & (i_18_) & (sk[116]) & (!g12)));
	assign g372 = (((i_17_) & (!sk[117]) & (!i_9_) & (g371)) + ((!i_17_) & (sk[117]) & (!i_9_) & (!g371)));
	assign g373 = (((!i_16_) & (!i_7_) & (!sk[118]) & (!i_8_) & (i_0_) & (!i_37_)) + ((i_16_) & (!i_7_) & (!sk[118]) & (!i_8_) & (!i_0_) & (i_37_)) + ((!i_16_) & (!i_7_) & (sk[118]) & (!i_8_) & (!i_0_) & (i_37_)));
	assign g374 = (((!i_33_) & (!i_13_) & (!i_14_) & (!sk[119]) & (g14) & (!g373)) + ((i_33_) & (!i_13_) & (!i_14_) & (!sk[119]) & (!g14) & (g373)) + ((!i_33_) & (!i_13_) & (!i_14_) & (!sk[119]) & (g14) & (g373)) + ((!i_33_) & (!i_13_) & (!i_14_) & (!sk[119]) & (g14) & (g373)));
	assign g375 = (((!i_7_) & (!sk[120]) & (!g53) & (!g286) & (g263)) + ((i_7_) & (!sk[120]) & (!g53) & (g286) & (!g263)) + ((!i_7_) & (!sk[120]) & (g53) & (g286) & (g263)));
	assign g376 = (((!i_29_) & (!i_8_) & (!g263) & (!sk[121]) & (g267) & (!g375)) + ((i_29_) & (!i_8_) & (!g263) & (!sk[121]) & (!g267) & (g375)) + ((i_29_) & (!i_8_) & (!g263) & (sk[121]) & (!g267) & (!g375)) + ((i_29_) & (i_8_) & (!g263) & (!sk[121]) & (g267) & (!g375)) + ((i_29_) & (!i_8_) & (!g263) & (!sk[121]) & (g267) & (!g375)));
	assign g377 = (((i_17_) & (!sk[122]) & (!g33) & (g49)) + ((!i_17_) & (sk[122]) & (g33) & (g49)));
	assign g378 = (((!sk[123]) & (!g33) & (!i_29_) & (!i_20_) & (g377) & (!g255)) + ((!sk[123]) & (g33) & (!i_29_) & (!i_20_) & (!g377) & (g255)) + ((!sk[123]) & (!g33) & (!i_29_) & (!i_20_) & (g377) & (g255)) + ((sk[123]) & (g33) & (i_29_) & (!i_20_) & (!g377) & (!g255)));
	assign g379 = (((!sk[124]) & (!i_12_) & (!g372) & (!g374) & (g376) & (!g378)) + ((sk[124]) & (!i_12_) & (!g372) & (!g374) & (!g376) & (g378)) + ((!sk[124]) & (i_12_) & (!g372) & (!g374) & (!g376) & (g378)) + ((!sk[124]) & (!i_12_) & (!g372) & (g374) & (g376) & (g378)) + ((!sk[124]) & (!i_12_) & (g372) & (g374) & (g376) & (g378)));
	assign g380 = (((!g101) & (!g202) & (!sk[125]) & (!g366) & (g370) & (!g379)) + ((!g101) & (!g202) & (sk[125]) & (!g366) & (!g370) & (!g379)) + ((g101) & (!g202) & (!sk[125]) & (!g366) & (!g370) & (g379)) + ((!g101) & (!g202) & (sk[125]) & (!g366) & (!g370) & (!g379)));
	assign g381 = (((!g45) & (!g286) & (!g326) & (!sk[126]) & (g328) & (!g331)) + ((g45) & (g286) & (!g326) & (!sk[126]) & (g328) & (!g331)) + ((g45) & (g286) & (!g326) & (!sk[126]) & (!g328) & (g331)) + ((g45) & (!g286) & (!g326) & (!sk[126]) & (!g328) & (g331)) + ((g45) & (g286) & (g326) & (sk[126]) & (!g328) & (!g331)));
	assign g382 = (((!sk[127]) & (!i_34_) & (!i_13_) & (!g58) & (g254)) + ((!sk[127]) & (i_34_) & (!i_13_) & (g58) & (!g254)) + ((!sk[127]) & (i_34_) & (!i_13_) & (g58) & (g254)));
	assign g383 = (((g20) & (i_34_) & (g79) & (i_37_) & (g367) & (!g382)) + ((g20) & (i_34_) & (!g79) & (i_37_) & (g367) & (g382)));
	assign g384 = (((!i_34_) & (!g53) & (!i_8_) & (!sk[1]) & (g29) & (!g254)) + ((i_34_) & (!g53) & (!i_8_) & (!sk[1]) & (!g29) & (g254)) + ((i_34_) & (g53) & (!i_8_) & (!sk[1]) & (g29) & (g254)));
	assign g385 = (((!sk[2]) & (i_33_) & (!i_34_) & (g5)) + ((sk[2]) & (!i_33_) & (i_34_) & (!g5)));
	assign g386 = (((!g1) & (!g18) & (!i_37_) & (!sk[3]) & (g384) & (!g385)) + ((g1) & (!g18) & (!i_37_) & (!sk[3]) & (!g384) & (g385)) + ((g1) & (g18) & (i_37_) & (!sk[3]) & (!g384) & (g385)) + ((g1) & (!g18) & (i_37_) & (!sk[3]) & (g384) & (g385)));
	assign g387 = (((!i_33_) & (!g7) & (!sk[4]) & (!g65) & (g263) & (!g336)) + ((!i_33_) & (!g7) & (!sk[4]) & (g65) & (g263) & (!g336)) + ((i_33_) & (!g7) & (!sk[4]) & (!g65) & (!g263) & (g336)) + ((!i_33_) & (g7) & (sk[4]) & (!g65) & (!g263) & (g336)));
	assign g388 = (((!g94) & (!i_7_) & (!sk[5]) & (!i_0_) & (g286)) + ((g94) & (!i_7_) & (!sk[5]) & (i_0_) & (!g286)) + ((g94) & (!i_7_) & (!sk[5]) & (!i_0_) & (g286)));
	assign g389 = (((!g111) & (!i_37_) & (!g387) & (!sk[6]) & (g388)) + ((g111) & (!i_37_) & (g387) & (!sk[6]) & (!g388)) + ((!g111) & (!i_37_) & (!g387) & (sk[6]) & (!g388)) + ((!g111) & (!i_37_) & (!g387) & (sk[6]) & (!g388)) + ((g111) & (!i_37_) & (g387) & (!sk[6]) & (!g388)));
	assign g390 = (((!i_33_) & (!g54) & (!g152) & (i_20_) & (!sk[7]) & (!g254)) + ((i_33_) & (!g54) & (!g152) & (!i_20_) & (!sk[7]) & (g254)) + ((!i_33_) & (!g54) & (g152) & (!i_20_) & (sk[7]) & (g254)) + ((!i_33_) & (g54) & (g152) & (!i_20_) & (sk[7]) & (g254)));
	assign g391 = (((!i_33_) & (!g28) & (!sk[8]) & (!g54) & (g48) & (!g254)) + ((i_33_) & (!g28) & (!sk[8]) & (!g54) & (!g48) & (g254)) + ((!i_33_) & (g28) & (!sk[8]) & (!g54) & (g48) & (g254)) + ((!i_33_) & (g28) & (!sk[8]) & (g54) & (g48) & (g254)));
	assign g392 = (((!g111) & (!g13) & (!i_20_) & (!sk[9]) & (g391)) + ((g111) & (!g13) & (i_20_) & (!sk[9]) & (!g391)) + ((g111) & (g13) & (!i_20_) & (!sk[9]) & (g391)));
	assign g393 = (((!sk[10]) & (!g111) & (!i_6_) & (!i_8_) & (g390) & (!g392)) + ((!sk[10]) & (g111) & (!i_6_) & (!i_8_) & (!g390) & (g392)) + ((sk[10]) & (!g111) & (!i_6_) & (!i_8_) & (!g390) & (!g392)) + ((!sk[10]) & (!g111) & (!i_6_) & (!i_8_) & (g390) & (!g392)) + ((!sk[10]) & (!g111) & (i_6_) & (!i_8_) & (g390) & (!g392)) + ((!sk[10]) & (!g111) & (!i_6_) & (i_8_) & (g390) & (!g392)));
	assign g394 = (((!sk[11]) & (!i_13_) & (!g248) & (!g323) & (g389) & (!g393)) + ((!sk[11]) & (i_13_) & (!g248) & (!g323) & (!g389) & (g393)) + ((sk[11]) & (!i_13_) & (g248) & (!g323) & (!g389) & (!g393)) + ((sk[11]) & (!i_13_) & (!g248) & (g323) & (!g389) & (!g393)));
	assign g395 = (((!sk[12]) & (!i_33_) & (!g45) & (!i_8_) & (g35) & (!g254)) + ((!sk[12]) & (i_33_) & (!g45) & (!i_8_) & (!g35) & (g254)) + ((!sk[12]) & (!i_33_) & (g45) & (!i_8_) & (g35) & (g254)));
	assign g396 = (((!i_28_) & (!g33) & (!g132) & (!sk[13]) & (i_25_) & (!i_20_)) + ((i_28_) & (!g33) & (!g132) & (!sk[13]) & (!i_25_) & (i_20_)) + ((!i_28_) & (g33) & (g132) & (!sk[13]) & (i_25_) & (i_20_)));
	assign g397 = (((!sk[14]) & (!i_34_) & (!i_30_) & (!g395) & (g396)) + ((!sk[14]) & (i_34_) & (!i_30_) & (g395) & (!g396)) + ((!sk[14]) & (i_34_) & (!i_30_) & (g395) & (!g396)) + ((!sk[14]) & (i_34_) & (!i_30_) & (!g395) & (g396)));
	assign g398 = (((!i_34_) & (!sk[15]) & (!i_35_) & (!i_21_) & (i_29_) & (!i_22_)) + ((i_34_) & (!sk[15]) & (!i_35_) & (i_21_) & (i_29_) & (!i_22_)) + ((!i_34_) & (!sk[15]) & (i_35_) & (i_21_) & (i_29_) & (!i_22_)) + ((i_34_) & (!sk[15]) & (!i_35_) & (!i_21_) & (!i_29_) & (i_22_)) + ((!i_34_) & (!sk[15]) & (i_35_) & (!i_21_) & (i_29_) & (i_22_)));
	assign g399 = (((!i_24_) & (!i_34_) & (!i_26_) & (!sk[16]) & (i_22_)) + ((i_24_) & (!i_34_) & (!i_26_) & (sk[16]) & (!i_22_)) + ((!i_24_) & (!i_34_) & (i_26_) & (sk[16]) & (!i_22_)) + ((!i_24_) & (i_34_) & (i_26_) & (!sk[16]) & (i_22_)) + ((i_24_) & (!i_34_) & (i_26_) & (!sk[16]) & (!i_22_)));
	assign g400 = (((!i_21_) & (!sk[17]) & (!i_29_) & (!i_20_) & (g399)) + ((i_21_) & (!sk[17]) & (!i_29_) & (i_20_) & (!g399)) + ((!i_21_) & (!sk[17]) & (i_29_) & (!i_20_) & (g399)));
	assign g401 = (((!i_24_) & (!i_34_) & (!sk[18]) & (!i_35_) & (i_26_) & (!g157)) + ((i_24_) & (!i_34_) & (!sk[18]) & (!i_35_) & (!i_26_) & (g157)) + ((!i_24_) & (!i_34_) & (sk[18]) & (!i_35_) & (!i_26_) & (g157)) + ((!i_24_) & (!i_34_) & (sk[18]) & (i_35_) & (!i_26_) & (g157)) + ((!i_24_) & (i_34_) & (!sk[18]) & (!i_35_) & (i_26_) & (g157)));
	assign g402 = (((!g3) & (!sk[19]) & (!g164) & (!g398) & (g400) & (!g401)) + ((g3) & (!sk[19]) & (!g164) & (!g398) & (!g400) & (g401)) + ((g3) & (!sk[19]) & (g164) & (!g398) & (!g400) & (g401)) + ((g3) & (!sk[19]) & (!g164) & (g398) & (!g400) & (g401)));
	assign g403 = (((!g2) & (!sk[20]) & (!i_21_) & (!g88) & (i_22_)) + ((g2) & (!sk[20]) & (!i_21_) & (g88) & (!i_22_)) + ((g2) & (!sk[20]) & (i_21_) & (g88) & (!i_22_)) + ((g2) & (!sk[20]) & (!i_21_) & (g88) & (i_22_)));
	assign g404 = (((!i_7_) & (!sk[21]) & (!g1) & (!g279) & (g403)) + ((!i_7_) & (sk[21]) & (!g1) & (!g279) & (!g403)) + ((!i_7_) & (sk[21]) & (!g1) & (!g279) & (!g403)) + ((i_7_) & (!sk[21]) & (!g1) & (g279) & (!g403)));
	assign g405 = (((!g86) & (!sk[22]) & (!g143) & (!i_25_) & (g404)) + ((g86) & (!sk[22]) & (!g143) & (i_25_) & (!g404)) + ((!g86) & (sk[22]) & (!g143) & (!i_25_) & (!g404)) + ((!g86) & (!sk[22]) & (g143) & (i_25_) & (g404)));
	assign g406 = (((!i_33_) & (!g28) & (!sk[23]) & (!g54) & (g254)) + ((i_33_) & (!g28) & (!sk[23]) & (g54) & (!g254)) + ((!i_33_) & (g28) & (!sk[23]) & (!g54) & (g254)) + ((!i_33_) & (g28) & (!sk[23]) & (g54) & (g254)));
	assign g407 = (((!i_8_) & (!i_0_) & (!g327) & (!sk[24]) & (g406)) + ((i_8_) & (!i_0_) & (g327) & (!sk[24]) & (!g406)) + ((!i_8_) & (!i_0_) & (g327) & (!sk[24]) & (g406)));
	assign g408 = (((g94) & (!i_8_) & (!i_0_) & (!g323) & (g390) & (!g259)) + ((g94) & (!i_8_) & (!i_0_) & (g323) & (!g390) & (g259)));
	assign g409 = (((!i_24_) & (!i_34_) & (!i_35_) & (i_26_) & (!sk[26]) & (!g334)) + ((!i_24_) & (!i_34_) & (!i_35_) & (!i_26_) & (sk[26]) & (!g334)) + ((i_24_) & (!i_34_) & (!i_35_) & (!i_26_) & (!sk[26]) & (g334)) + ((!i_24_) & (!i_34_) & (i_35_) & (!i_26_) & (sk[26]) & (!g334)) + ((!i_24_) & (i_34_) & (!i_35_) & (!i_26_) & (sk[26]) & (!g334)));
	assign g410 = (((!g3) & (!i_7_) & (!sk[27]) & (!i_31_) & (g157) & (!g409)) + ((g3) & (!i_7_) & (!sk[27]) & (!i_31_) & (!g157) & (g409)) + ((g3) & (i_7_) & (!sk[27]) & (i_31_) & (g157) & (g409)));
	assign g411 = (((!i_34_) & (!g57) & (!g88) & (!sk[28]) & (g137) & (!g410)) + ((i_34_) & (!g57) & (!g88) & (!sk[28]) & (!g137) & (g410)) + ((!i_34_) & (!g57) & (!g88) & (sk[28]) & (!g137) & (!g410)) + ((!i_34_) & (!g57) & (!g88) & (!sk[28]) & (g137) & (!g410)) + ((!i_34_) & (!g57) & (!g88) & (!sk[28]) & (g137) & (!g410)) + ((!i_34_) & (!g57) & (!g88) & (!sk[28]) & (g137) & (!g410)));
	assign g412 = (((!sk[29]) & (i_13_) & (!i_14_) & (g11)) + ((!sk[29]) & (i_13_) & (!i_14_) & (g11)));
	assign g413 = (((!g358) & (!sk[30]) & (!g311) & (!g377) & (g249) & (!g412)) + ((g358) & (!sk[30]) & (!g311) & (!g377) & (!g249) & (g412)) + ((!g358) & (!sk[30]) & (g311) & (g377) & (g249) & (!g412)));
	assign g414 = (((!g405) & (!g407) & (!sk[31]) & (!g408) & (g411) & (!g413)) + ((g405) & (!g407) & (!sk[31]) & (!g408) & (!g411) & (g413)) + ((!g405) & (!g407) & (!sk[31]) & (!g408) & (g411) & (!g413)));
	assign g415 = (((!i_34_) & (!g135) & (g156) & (!g397) & (!g402) & (g414)) + ((!i_34_) & (!g135) & (g156) & (!g397) & (!g402) & (g414)));
	assign g416 = (((i_14_) & (!sk[33]) & (!i_32_) & (g58)) + ((!i_14_) & (sk[33]) & (!i_32_) & (g58)));
	assign g417 = (((!sk[34]) & (!i_33_) & (!i_34_) & (!g21) & (g247) & (!g416)) + ((!sk[34]) & (i_33_) & (!i_34_) & (!g21) & (!g247) & (g416)) + ((sk[34]) & (!i_33_) & (i_34_) & (g21) & (!g247) & (!g416)) + ((sk[34]) & (!i_33_) & (i_34_) & (g21) & (!g247) & (g416)));
	assign g418 = (((!i_34_) & (!g1) & (!i_8_) & (g5) & (!sk[35]) & (!g29)) + ((i_34_) & (!g1) & (!i_8_) & (!g5) & (!sk[35]) & (g29)) + ((i_34_) & (g1) & (!i_8_) & (!g5) & (!sk[35]) & (g29)));
	assign g419 = (((g98) & (!sk[36]) & (!g55) & (g277) & (!g418)) + ((!g98) & (!sk[36]) & (!g55) & (!g277) & (g418)) + ((!g98) & (!sk[36]) & (g55) & (!g277) & (g418)));
	assign g420 = (((!i_33_) & (!i_32_) & (!sk[37]) & (!g122) & (g419)) + ((!i_33_) & (i_32_) & (sk[37]) & (!g122) & (!g419)) + ((!i_33_) & (!i_32_) & (sk[37]) & (!g122) & (!g419)) + ((i_33_) & (!i_32_) & (!sk[37]) & (g122) & (!g419)));
	assign g421 = (((!i_33_) & (!sk[38]) & (!g2) & (!i_32_) & (g150) & (!g134)) + ((i_33_) & (!sk[38]) & (!g2) & (!i_32_) & (!g150) & (g134)) + ((!i_33_) & (!sk[38]) & (g2) & (!i_32_) & (g150) & (!g134)) + ((!i_33_) & (sk[38]) & (g2) & (!i_32_) & (!g150) & (g134)));
	assign g422 = (((!sk[39]) & (!i_30_) & (!i_31_) & (!i_29_) & (i_37_) & (!g421)) + ((!sk[39]) & (i_30_) & (!i_31_) & (!i_29_) & (!i_37_) & (g421)) + ((!sk[39]) & (!i_30_) & (i_31_) & (!i_29_) & (i_37_) & (g421)));
	assign g423 = (((g53) & (g367) & (!sk[40]) & (g341)) + ((g53) & (!g367) & (!sk[40]) & (g341)));
	assign g424 = (((!i_29_) & (!g18) & (!g279) & (!sk[41]) & (g422) & (!g423)) + ((i_29_) & (!g18) & (!g279) & (!sk[41]) & (!g422) & (g423)) + ((i_29_) & (!g18) & (!g279) & (sk[41]) & (!g422) & (!g423)) + ((!i_29_) & (!g18) & (!g279) & (sk[41]) & (!g422) & (!g423)) + ((!i_29_) & (!g18) & (!g279) & (sk[41]) & (!g422) & (!g423)));
	assign g425 = (((!g3) & (!g254) & (!sk[42]) & (!g417) & (g420) & (!g424)) + ((!g3) & (!g254) & (sk[42]) & (!g417) & (!g420) & (!g424)) + ((!g3) & (!g254) & (!sk[42]) & (!g417) & (g420) & (!g424)) + ((g3) & (!g254) & (!sk[42]) & (!g417) & (!g420) & (g424)) + ((!g3) & (!g254) & (!sk[42]) & (!g417) & (g420) & (g424)) + ((!g3) & (!g254) & (sk[42]) & (!g417) & (!g420) & (g424)));
	assign g426 = (((!g381) & (!g383) & (!g386) & (!g394) & (g415) & (g425)));
	assign g427 = (((!sk[44]) & (!g293) & (!g319) & (!g357) & (g380) & (!g426)) + ((!sk[44]) & (g293) & (!g319) & (!g357) & (!g380) & (g426)) + ((!sk[44]) & (!g293) & (g319) & (!g357) & (g380) & (g426)));
	assign g428 = (((!i_35_) & (!sk[45]) & (i_38_)) + ((!i_35_) & (!sk[45]) & (i_38_)));
	assign g429 = (((!sk[46]) & (!i_33_) & (g428)) + ((!sk[46]) & (!i_33_) & (g428)));
	assign g430 = (((!i_9_) & (!i_8_) & (!g9) & (i_10_) & (!sk[47]) & (!g29)) + ((i_9_) & (!i_8_) & (!g9) & (!i_10_) & (!sk[47]) & (g29)) + ((i_9_) & (!i_8_) & (!g9) & (!i_10_) & (!sk[47]) & (g29)) + ((i_9_) & (!i_8_) & (g9) & (!i_10_) & (sk[47]) & (!g29)));
	assign g431 = (((!i_33_) & (!sk[48]) & (!i_7_) & (!g70) & (i_38_)) + ((i_33_) & (!sk[48]) & (!i_7_) & (g70) & (!i_38_)) + ((!i_33_) & (!sk[48]) & (!i_7_) & (!g70) & (i_38_)));
	assign g432 = (((!i_2_) & (!sk[49]) & (!i_8_) & (!g96) & (g429) & (!g431)) + ((!i_2_) & (sk[49]) & (!i_8_) & (!g96) & (!g429) & (g431)) + ((i_2_) & (!sk[49]) & (!i_8_) & (!g96) & (!g429) & (g431)) + ((!i_2_) & (!sk[49]) & (!i_8_) & (g96) & (g429) & (!g431)));
	assign g433 = (((!sk[50]) & (!i_33_) & (!g57) & (!g9) & (g29) & (!g428)) + ((!sk[50]) & (i_33_) & (!g57) & (!g9) & (!g29) & (g428)) + ((!sk[50]) & (!i_33_) & (g57) & (!g9) & (g29) & (g428)) + ((sk[50]) & (!i_33_) & (g57) & (g9) & (!g29) & (g428)));
	assign g434 = (((!i_23_) & (!sk[51]) & (!i_29_) & (!g157) & (g433)) + ((i_23_) & (!sk[51]) & (!i_29_) & (g157) & (!g433)) + ((!i_23_) & (sk[51]) & (!i_29_) & (!g157) & (!g433)) + ((!i_23_) & (sk[51]) & (!i_29_) & (g157) & (!g433)));
	assign g435 = (((!sk[52]) & (!i_31_) & (g428)) + ((!sk[52]) & (!i_31_) & (g428)));
	assign g436 = (((!i_2_) & (!i_7_) & (!i_9_) & (i_3_) & (!i_18_) & (g14)));
	assign g437 = (((g12) & (!g32) & (!sk[54]) & (g436)) + ((!g12) & (!g32) & (sk[54]) & (!g436)) + ((!g12) & (!g32) & (sk[54]) & (!g436)));
	assign g438 = (((i_32_) & (sk[55]) & (!g25) & (!g437)) + ((i_32_) & (!sk[55]) & (!g25) & (g437)) + ((!i_32_) & (sk[55]) & (!g25) & (g437)));
	assign g439 = (((!i_9_) & (!i_3_) & (!sk[56]) & (!i_18_) & (g14) & (!g46)) + ((i_9_) & (!i_3_) & (!sk[56]) & (!i_18_) & (!g14) & (g46)) + ((!i_9_) & (i_3_) & (!sk[56]) & (!i_18_) & (g14) & (g46)));
	assign g440 = (((!sk[57]) & (g12) & (!g49) & (g439)) + ((sk[57]) & (!g12) & (!g49) & (!g439)) + ((sk[57]) & (!g12) & (!g49) & (!g439)));
	assign g441 = (((!i_33_) & (!sk[58]) & (!i_38_) & (!g435) & (g438) & (!g440)) + ((i_33_) & (!sk[58]) & (!i_38_) & (!g435) & (!g438) & (g440)) + ((!i_33_) & (sk[58]) & (i_38_) & (!g435) & (!g438) & (!g440)) + ((!i_33_) & (sk[58]) & (!i_38_) & (g435) & (!g438) & (!g440)));
	assign g442 = (((g121) & (!g429) & (!g430) & (g432) & (!g434) & (!g441)) + ((g121) & (!g429) & (!g430) & (!g432) & (!g434) & (!g441)) + ((g121) & (!g429) & (!g430) & (!g432) & (!g434) & (g441)) + ((g121) & (g429) & (g430) & (!g432) & (!g434) & (!g441)));
	assign g443 = (((!g71) & (!sk[60]) & (i_25_)) + ((!g71) & (sk[60]) & (!i_25_)));
	assign g444 = (((i_35_) & (!sk[61]) & (!i_31_) & (g438) & (!g440)) + ((!i_35_) & (!sk[61]) & (!i_31_) & (!g438) & (g440)) + ((!i_35_) & (!sk[61]) & (!i_31_) & (g438) & (g440)) + ((!i_35_) & (sk[61]) & (i_31_) & (g438) & (!g440)));
	assign g445 = (((!i_32_) & (!i_31_) & (!sk[62]) & (!g9) & (g29) & (!g428)) + ((i_32_) & (!i_31_) & (!sk[62]) & (!g9) & (!g29) & (g428)) + ((!i_32_) & (!i_31_) & (!sk[62]) & (!g9) & (g29) & (g428)) + ((!i_32_) & (!i_31_) & (sk[62]) & (g9) & (!g29) & (g428)));
	assign g446 = (((!i_2_) & (!i_7_) & (!g70) & (i_38_) & (!sk[63]) & (!g445)) + ((i_2_) & (!i_7_) & (!g70) & (!i_38_) & (!sk[63]) & (g445)) + ((!i_2_) & (!i_7_) & (!g70) & (!i_38_) & (sk[63]) & (!g445)) + ((i_2_) & (!i_7_) & (!g70) & (!i_38_) & (sk[63]) & (!g445)) + ((!i_2_) & (i_7_) & (!g70) & (!i_38_) & (sk[63]) & (!g445)) + ((!i_2_) & (!i_7_) & (g70) & (!i_38_) & (sk[63]) & (!g445)));
	assign g447 = (((!g46) & (!g223) & (!g428) & (!sk[64]) & (g430) & (!g446)) + ((g46) & (!g223) & (!g428) & (!sk[64]) & (!g430) & (g446)) + ((!g46) & (!g223) & (!g428) & (sk[64]) & (!g430) & (g446)) + ((!g46) & (!g223) & (!g428) & (sk[64]) & (!g430) & (g446)) + ((!g46) & (!g223) & (!g428) & (sk[64]) & (!g430) & (g446)));
	assign g448 = (((!sk[65]) & (!i_28_) & (!i_38_) & (!g443) & (g444) & (!g447)) + ((!sk[65]) & (i_28_) & (!i_38_) & (!g443) & (!g444) & (g447)) + ((sk[65]) & (!i_28_) & (!i_38_) & (g443) & (!g444) & (!g447)) + ((sk[65]) & (!i_28_) & (i_38_) & (g443) & (!g444) & (!g447)));
	assign g449 = (((!sk[66]) & (!i_18_) & (!i_11_) & (!i_19_) & (g67) & (!g10)) + ((!sk[66]) & (!i_18_) & (!i_11_) & (!i_19_) & (g67) & (!g10)) + ((!sk[66]) & (i_18_) & (!i_11_) & (!i_19_) & (!g67) & (g10)) + ((sk[66]) & (!i_18_) & (!i_11_) & (!i_19_) & (!g67) & (g10)));
	assign g450 = (((!i_32_) & (!i_25_) & (!sk[67]) & (!g449) & (g435)) + ((i_32_) & (!i_25_) & (!sk[67]) & (g449) & (!g435)) + ((!i_32_) & (!i_25_) & (!sk[67]) & (g449) & (g435)));
	assign g451 = (((!i_7_) & (!sk[68]) & (!i_8_) & (!g9) & (g29)) + ((i_7_) & (!sk[68]) & (!i_8_) & (g9) & (!g29)) + ((!i_7_) & (!sk[68]) & (!i_8_) & (!g9) & (g29)) + ((!i_7_) & (sk[68]) & (!i_8_) & (g9) & (!g29)));
	assign g452 = (((!i_9_) & (!sk[69]) & (!g65) & (!g9) & (i_10_)) + ((i_9_) & (!sk[69]) & (!g65) & (g9) & (!i_10_)) + ((i_9_) & (!sk[69]) & (g65) & (g9) & (!i_10_)));
	assign g453 = (((!i_33_) & (!i_31_) & (!sk[70]) & (!g65) & (g449)) + ((i_33_) & (!i_31_) & (!sk[70]) & (g65) & (!g449)) + ((!i_33_) & (!i_31_) & (!sk[70]) & (g65) & (g449)));
	assign g454 = (((!g164) & (!i_38_) & (!g451) & (g452) & (!sk[71]) & (!g453)) + ((!g164) & (i_38_) & (!g451) & (g452) & (!sk[71]) & (!g453)) + ((!g164) & (i_38_) & (!g451) & (!g452) & (sk[71]) & (g453)) + ((g164) & (!i_38_) & (!g451) & (!g452) & (!sk[71]) & (g453)) + ((!g164) & (i_38_) & (g451) & (!g452) & (sk[71]) & (!g453)));
	assign g455 = (((sk[72]) & (!i_8_) & (g9) & (!g29)) + ((!sk[72]) & (i_8_) & (!g9) & (g29)) + ((sk[72]) & (!i_8_) & (!g9) & (g29)));
	assign g456 = (((!sk[73]) & (i_13_) & (!i_9_) & (i_18_)) + ((sk[73]) & (!i_13_) & (i_9_) & (i_18_)));
	assign g457 = (((i_11_) & (!sk[74]) & (!g455) & (g456)) + ((i_11_) & (!sk[74]) & (g455) & (g456)));
	assign g458 = (((!i_12_) & (i_9_) & (!i_3_) & (g14) & (!i_1_) & (g46)) + ((!i_12_) & (i_9_) & (!i_3_) & (g14) & (!i_1_) & (g46)));
	assign g459 = (((!sk[76]) & (i_13_) & (!i_11_) & (g458)) + ((sk[76]) & (!i_13_) & (i_11_) & (g458)));
	assign g460 = (((!i_33_) & (!i_30_) & (!i_32_) & (!sk[77]) & (i_31_) & (!i_25_)) + ((i_33_) & (!i_30_) & (!i_32_) & (!sk[77]) & (!i_31_) & (i_25_)) + ((!i_33_) & (!i_30_) & (!i_32_) & (sk[77]) & (!i_31_) & (!i_25_)) + ((!i_33_) & (!i_30_) & (!i_32_) & (sk[77]) & (!i_31_) & (!i_25_)));
	assign g461 = (((!i_2_) & (!g164) & (g428) & (g457) & (!g459) & (!g460)) + ((!i_2_) & (!g164) & (g428) & (!g457) & (g459) & (!g460)) + ((!i_2_) & (!g164) & (g428) & (!g457) & (!g459) & (g460)));
	assign g462 = (((!i_24_) & (!i_28_) & (!i_26_) & (g450) & (!g454) & (!g461)) + ((!i_24_) & (!i_28_) & (!i_26_) & (!g450) & (g454) & (!g461)) + ((!i_24_) & (!i_28_) & (!i_26_) & (!g450) & (!g454) & (g461)));
	assign g463 = (((!i_32_) & (!sk[80]) & (!g223) & (!g443) & (g428)) + ((i_32_) & (!sk[80]) & (!g223) & (g443) & (!g428)) + ((!i_32_) & (!sk[80]) & (g223) & (g443) & (g428)));
	assign g464 = (((!i_12_) & (!g86) & (!g121) & (g429) & (!sk[81]) & (!g463)) + ((i_12_) & (!g86) & (!g121) & (!g429) & (!sk[81]) & (g463)) + ((i_12_) & (!g86) & (g121) & (g429) & (!sk[81]) & (!g463)));
	assign g465 = (((!i_35_) & (!i_31_) & (!i_8_) & (!sk[82]) & (i_38_)) + ((i_35_) & (!i_31_) & (i_8_) & (!sk[82]) & (!i_38_)) + ((!i_35_) & (!i_31_) & (!i_8_) & (!sk[82]) & (i_38_)));
	assign g466 = (((!sk[83]) & (!i_7_) & (!i_32_) & (!g335) & (i_38_) & (!g465)) + ((!sk[83]) & (i_7_) & (!i_32_) & (!g335) & (!i_38_) & (g465)) + ((sk[83]) & (!i_7_) & (!i_32_) & (g335) & (!i_38_) & (g465)) + ((!sk[83]) & (!i_7_) & (!i_32_) & (g335) & (i_38_) & (!g465)));
	assign g467 = (((!i_28_) & (!i_26_) & (!sk[84]) & (!i_25_) & (g466)) + ((i_28_) & (!i_26_) & (!sk[84]) & (i_25_) & (!g466)) + ((!i_28_) & (!i_26_) & (!sk[84]) & (!i_25_) & (g466)));
	assign g468 = (((!sk[85]) & (!i_28_) & (!i_26_) & (!i_31_) & (g48)) + ((!sk[85]) & (i_28_) & (!i_26_) & (i_31_) & (!g48)) + ((!sk[85]) & (!i_28_) & (!i_26_) & (!i_31_) & (g48)));
	assign g469 = (((!i_28_) & (!i_26_) & (!sk[86]) & (!i_32_) & (g31)) + ((i_28_) & (!i_26_) & (!sk[86]) & (i_32_) & (!g31)) + ((!i_28_) & (!i_26_) & (!sk[86]) & (!i_32_) & (g31)));
	assign g470 = (((!i_33_) & (!i_35_) & (!sk[87]) & (!i_38_) & (g468) & (!g469)) + ((i_33_) & (!i_35_) & (!sk[87]) & (!i_38_) & (!g468) & (g469)) + ((!i_33_) & (!i_35_) & (!sk[87]) & (i_38_) & (g468) & (!g469)) + ((!i_33_) & (!i_35_) & (sk[87]) & (i_38_) & (!g468) & (g469)));
	assign g471 = (((!i_24_) & (!sk[88]) & (!g8) & (!g467) & (g470)) + ((i_24_) & (!sk[88]) & (!g8) & (g467) & (!g470)) + ((!i_24_) & (!sk[88]) & (g8) & (!g467) & (g470)) + ((!i_24_) & (sk[88]) & (g8) & (g467) & (!g470)));
	assign g472 = (((!i_35_) & (!sk[89]) & (!i_30_) & (!i_32_) & (i_38_)) + ((i_35_) & (!sk[89]) & (!i_30_) & (i_32_) & (!i_38_)) + ((!i_35_) & (!sk[89]) & (!i_30_) & (!i_32_) & (i_38_)));
	assign g473 = (((!sk[90]) & (!i_33_) & (!i_28_) & (!g71) & (i_25_) & (!g472)) + ((!sk[90]) & (i_33_) & (!i_28_) & (!g71) & (!i_25_) & (g472)) + ((sk[90]) & (!i_33_) & (!i_28_) & (!g71) & (!i_25_) & (g472)) + ((sk[90]) & (!i_33_) & (!i_28_) & (!g71) & (!i_25_) & (g472)));
	assign g474 = (((i_13_) & (!i_3_) & (!sk[91]) & (i_11_)) + ((!i_13_) & (!i_3_) & (sk[91]) & (i_11_)));
	assign g475 = (((i_2_) & (!sk[92]) & (!i_9_) & (g473) & (!g474)) + ((!i_2_) & (!sk[92]) & (!i_9_) & (!g473) & (g474)) + ((!i_2_) & (sk[92]) & (!i_9_) & (!g473) & (!g474)) + ((!i_2_) & (!sk[92]) & (!i_9_) & (!g473) & (g474)) + ((!i_2_) & (!sk[92]) & (!i_9_) & (!g473) & (g474)));
	assign g476 = (((!i_13_) & (!i_9_) & (!g160) & (!g464) & (!g471) & (g696)) + ((!i_13_) & (!i_9_) & (!g160) & (!g464) & (!g471) & (g696)) + ((!i_13_) & (!i_9_) & (!g160) & (!g464) & (!g471) & (g696)) + ((!i_13_) & (!i_9_) & (!g160) & (!g464) & (!g471) & (g696)));
	assign g477 = (((i_22_) & (!g160) & (!g442) & (!g448) & (!g462) & (!g476)) + ((!i_22_) & (!g160) & (!g442) & (!g448) & (!g462) & (g476)));
	assign g478 = (((!i_24_) & (!sk[95]) & (i_25_)) + ((!i_24_) & (sk[95]) & (!i_25_)));
	assign g479 = (((!i_33_) & (!i_28_) & (!i_32_) & (!sk[96]) & (i_29_) & (!i_25_)) + ((i_33_) & (!i_28_) & (!i_32_) & (!sk[96]) & (!i_29_) & (i_25_)) + ((!i_33_) & (!i_28_) & (!i_32_) & (sk[96]) & (!i_29_) & (!i_25_)) + ((!i_33_) & (!i_28_) & (!i_32_) & (sk[96]) & (!i_29_) & (!i_25_)));
	assign g480 = (((!i_24_) & (!i_30_) & (!g1) & (g7) & (!sk[97]) & (!i_25_)) + ((i_24_) & (!i_30_) & (!g1) & (!g7) & (!sk[97]) & (i_25_)) + ((!i_24_) & (!i_30_) & (g1) & (g7) & (!sk[97]) & (!i_25_)));
	assign g481 = (((!i_24_) & (!g32) & (!g24) & (!sk[98]) & (g479) & (!g480)) + ((i_24_) & (!g32) & (!g24) & (!sk[98]) & (!g479) & (g480)) + ((!i_24_) & (!g32) & (!g24) & (sk[98]) & (!g479) & (!g480)) + ((i_24_) & (!g32) & (!g24) & (!sk[98]) & (g479) & (!g480)) + ((!i_24_) & (!g32) & (!g24) & (!sk[98]) & (g479) & (!g480)) + ((!i_24_) & (!g32) & (g24) & (!sk[98]) & (g479) & (!g480)));
	assign g482 = (((!i_33_) & (!i_24_) & (!sk[99]) & (!g1) & (g25) & (!g481)) + ((i_33_) & (!i_24_) & (!sk[99]) & (!g1) & (!g25) & (g481)) + ((!i_33_) & (!i_24_) & (sk[99]) & (!g1) & (!g25) & (g481)) + ((!i_33_) & (i_24_) & (!sk[99]) & (!g1) & (g25) & (g481)) + ((!i_33_) & (!i_24_) & (!sk[99]) & (!g1) & (g25) & (g481)));
	assign g483 = (((!sk[100]) & (!i_7_) & (!i_32_) & (!g84) & (g478) & (!g482)) + ((!sk[100]) & (i_7_) & (!i_32_) & (!g84) & (!g478) & (g482)) + ((sk[100]) & (!i_7_) & (!i_32_) & (!g84) & (!g478) & (g482)) + ((!sk[100]) & (!i_7_) & (i_32_) & (!g84) & (g478) & (g482)) + ((!sk[100]) & (!i_7_) & (!i_32_) & (!g84) & (g478) & (g482)));
	assign g484 = (((!i_24_) & (!g12) & (!g32) & (!sk[101]) & (g436)) + ((!i_24_) & (!g12) & (!g32) & (!sk[101]) & (g436)) + ((i_24_) & (!g12) & (g32) & (!sk[101]) & (!g436)) + ((!i_24_) & (g12) & (g32) & (sk[101]) & (!g436)));
	assign g485 = (((!sk[102]) & (!g37) & (g484)) + ((!sk[102]) & (g37) & (g484)));
	assign g486 = (((g12) & (!sk[103]) & (!i_8_) & (g11) & (!g436)) + ((!g12) & (!sk[103]) & (!i_8_) & (!g11) & (g436)) + ((!g12) & (!sk[103]) & (!i_8_) & (!g11) & (g436)));
	assign g487 = (((!i_24_) & (!i_30_) & (!g1) & (!sk[104]) & (g7) & (!g486)) + ((i_24_) & (!i_30_) & (!g1) & (!sk[104]) & (!g7) & (g486)) + ((!i_24_) & (!i_30_) & (g1) & (!sk[104]) & (g7) & (!g486)) + ((!i_24_) & (!i_30_) & (g1) & (sk[104]) & (!g7) & (g486)));
	assign g488 = (((!sk[105]) & (!i_24_) & (i_28_)) + ((sk[105]) & (!i_24_) & (!i_28_)));
	assign g489 = (((!i_7_) & (!i_29_) & (!sk[106]) & (!g70) & (g488)) + ((i_7_) & (!i_29_) & (!sk[106]) & (g70) & (!g488)) + ((!i_7_) & (!i_29_) & (!sk[106]) & (!g70) & (g488)));
	assign g490 = (((!i_33_) & (i_38_) & (!g483) & (!g485) & (!g487) & (!g489)) + ((!i_33_) & (i_38_) & (!g483) & (g485) & (!g487) & (!g489)) + ((!i_33_) & (i_38_) & (!g483) & (!g485) & (g487) & (!g489)) + ((!i_33_) & (i_38_) & (!g483) & (!g485) & (!g487) & (g489)));
	assign g491 = (((!sk[108]) & (i_24_) & (!i_9_) & (i_10_)) + ((sk[108]) & (!i_24_) & (i_9_) & (!i_10_)));
	assign g492 = (((i_30_) & (!i_32_) & (!sk[109]) & (g428)) + ((!i_30_) & (!i_32_) & (sk[109]) & (g428)));
	assign g493 = (((!g1) & (!sk[110]) & (!i_25_) & (!g491) & (g492)) + ((g1) & (!sk[110]) & (!i_25_) & (g491) & (!g492)) + ((g1) & (!sk[110]) & (!i_25_) & (g491) & (g492)));
	assign g494 = (((!sk[111]) & (!i_28_) & (g478)) + ((!sk[111]) & (!i_28_) & (g478)));
	assign g495 = (((!sk[112]) & (i_9_) & (!i_8_) & (i_10_)) + ((sk[112]) & (i_9_) & (!i_8_) & (!i_10_)));
	assign g496 = (((!i_30_) & (!i_29_) & (!g428) & (!sk[113]) & (g494) & (!g495)) + ((i_30_) & (!i_29_) & (!g428) & (!sk[113]) & (!g494) & (g495)) + ((!i_30_) & (!i_29_) & (g428) & (!sk[113]) & (g494) & (g495)));
	assign g497 = (((!g84) & (!g478) & (!g465) & (g493) & (!sk[114]) & (!g496)) + ((g84) & (!g478) & (!g465) & (!g493) & (!sk[114]) & (g496)) + ((!g84) & (!g478) & (!g465) & (!g493) & (sk[114]) & (!g496)) + ((!g84) & (!g478) & (!g465) & (!g493) & (sk[114]) & (!g496)) + ((!g84) & (!g478) & (!g465) & (!g493) & (sk[114]) & (!g496)));
	assign g498 = (((!i_24_) & (!sk[115]) & (!g12) & (!g49) & (g439)) + ((!i_24_) & (!sk[115]) & (!g12) & (!g49) & (g439)) + ((i_24_) & (!sk[115]) & (!g12) & (g49) & (!g439)) + ((!i_24_) & (sk[115]) & (g12) & (g49) & (!g439)));
	assign g499 = (((!sk[116]) & (!i_24_) & (!i_35_) & (!i_31_) & (g25) & (!g498)) + ((!sk[116]) & (!i_24_) & (!i_35_) & (!i_31_) & (g25) & (!g498)) + ((!sk[116]) & (i_24_) & (!i_35_) & (!i_31_) & (!g25) & (g498)) + ((sk[116]) & (!i_24_) & (!i_35_) & (!i_31_) & (!g25) & (g498)));
	assign g500 = (((!sk[117]) & (g1) & (!i_25_) & (i_38_)) + ((!sk[117]) & (g1) & (!i_25_) & (i_38_)));
	assign g501 = (((i_29_) & (!g494) & (!sk[118]) & (g435)) + ((!i_29_) & (g494) & (sk[118]) & (g435)));
	assign g502 = (((!i_24_) & (!g60) & (!sk[119]) & (!g429) & (g455) & (!g501)) + ((!i_24_) & (!g60) & (!sk[119]) & (!g429) & (g455) & (g501)) + ((i_24_) & (!g60) & (!sk[119]) & (!g429) & (!g455) & (g501)) + ((!i_24_) & (g60) & (!sk[119]) & (g429) & (g455) & (!g501)));
	assign g503 = (((!sk[120]) & (!i_32_) & (!g484) & (!g499) & (g500) & (!g502)) + ((!sk[120]) & (i_32_) & (!g484) & (!g499) & (!g500) & (g502)) + ((sk[120]) & (!i_32_) & (!g484) & (!g499) & (!g500) & (!g502)) + ((!sk[120]) & (i_32_) & (!g484) & (!g499) & (g500) & (!g502)) + ((!sk[120]) & (!i_32_) & (!g484) & (!g499) & (g500) & (!g502)));
	assign g504 = (((!sk[121]) & (!i_24_) & (!i_17_) & (!i_12_) & (g22)) + ((!sk[121]) & (!i_24_) & (!i_17_) & (!i_12_) & (g22)) + ((!sk[121]) & (i_24_) & (!i_17_) & (i_12_) & (!g22)) + ((sk[121]) & (!i_24_) & (i_17_) & (i_12_) & (!g22)));
	assign g505 = (((!sk[122]) & (!i_28_) & (!i_31_) & (!i_29_) & (g504)) + ((!sk[122]) & (i_28_) & (!i_31_) & (i_29_) & (!g504)) + ((!sk[122]) & (!i_28_) & (i_31_) & (!i_29_) & (g504)));
	assign g506 = (((!i_24_) & (!i_30_) & (!g1) & (g429) & (!sk[123]) & (!g495)) + ((i_24_) & (!i_30_) & (!g1) & (!g429) & (!sk[123]) & (g495)) + ((!i_24_) & (!i_30_) & (g1) & (g429) & (!sk[123]) & (g495)));
	assign g507 = (((!i_17_) & (!sk[124]) & (!i_12_) & (!g22) & (g86)) + ((!i_17_) & (!sk[124]) & (!i_12_) & (g22) & (g86)) + ((i_17_) & (!sk[124]) & (!i_12_) & (g22) & (!g86)) + ((i_17_) & (!sk[124]) & (i_12_) & (!g22) & (g86)));
	assign g508 = (((!sk[125]) & (!i_23_) & (!i_22_) & (!g488) & (g507)) + ((!sk[125]) & (i_23_) & (!i_22_) & (g488) & (!g507)) + ((!sk[125]) & (i_23_) & (i_22_) & (g488) & (!g507)) + ((!sk[125]) & (!i_23_) & (i_22_) & (g488) & (g507)));
	assign g509 = (((!i_14_) & (!g133) & (!sk[126]) & (!g505) & (g506) & (!g508)) + ((i_14_) & (!g133) & (!sk[126]) & (!g505) & (!g506) & (g508)) + ((!i_14_) & (!g133) & (sk[126]) & (!g505) & (!g506) & (!g508)) + ((!i_14_) & (!g133) & (sk[126]) & (!g505) & (!g506) & (!g508)));
	assign g510 = (((!i_34_) & (!g490) & (!g497) & (g503) & (!sk[127]) & (!g509)) + ((i_34_) & (g490) & (!g497) & (!g503) & (!sk[127]) & (g509)) + ((i_34_) & (!g490) & (!g497) & (!g503) & (!sk[127]) & (g509)) + ((i_34_) & (!g490) & (!g497) & (!g503) & (!sk[127]) & (g509)) + ((i_34_) & (!g490) & (!g497) & (!g503) & (sk[127]) & (!g509)));
	assign g511 = (((i_30_) & (!g121) & (!sk[0]) & (g495)) + ((!i_30_) & (g121) & (sk[0]) & (g495)));
	assign g512 = (((i_34_) & (!i_26_) & (!sk[1]) & (g488)) + ((!i_34_) & (!i_26_) & (sk[1]) & (g488)));
	assign g513 = (((!i_33_) & (!i_29_) & (!g457) & (!g459) & (g511) & (!g512)) + ((!i_33_) & (!i_29_) & (g457) & (!g459) & (!g511) & (g512)) + ((!i_33_) & (!i_29_) & (!g457) & (g459) & (!g511) & (g512)));
	assign g514 = (((!i_13_) & (!i_11_) & (!g478) & (!sk[3]) & (g457) & (!g458)) + ((!i_13_) & (!i_11_) & (g478) & (!sk[3]) & (g457) & (!g458)) + ((i_13_) & (!i_11_) & (!g478) & (!sk[3]) & (!g457) & (g458)) + ((!i_13_) & (i_11_) & (g478) & (sk[3]) & (!g457) & (g458)));
	assign g515 = (((!i_34_) & (!i_26_) & (!i_29_) & (!sk[4]) & (i_22_)) + ((i_34_) & (!i_26_) & (!i_29_) & (sk[4]) & (!i_22_)) + ((i_34_) & (!i_26_) & (i_29_) & (!sk[4]) & (!i_22_)) + ((!i_34_) & (!i_26_) & (!i_29_) & (sk[4]) & (!i_22_)) + ((!i_34_) & (!i_26_) & (!i_29_) & (!sk[4]) & (i_22_)));
	assign g516 = (((!i_13_) & (!i_19_) & (!g488) & (!sk[5]) & (g458)) + ((i_13_) & (!i_19_) & (g488) & (!sk[5]) & (!g458)) + ((!i_13_) & (i_19_) & (g488) & (!sk[5]) & (g458)));
	assign g517 = (((!i_13_) & (!i_18_) & (!sk[6]) & (!i_19_) & (g488)) + ((i_13_) & (!i_18_) & (!sk[6]) & (i_19_) & (!g488)) + ((!i_13_) & (i_18_) & (!sk[6]) & (i_19_) & (g488)));
	assign g518 = (((!i_9_) & (!i_8_) & (!g9) & (g29) & (!sk[7]) & (!g517)) + ((i_9_) & (!i_8_) & (!g9) & (!g29) & (!sk[7]) & (g517)) + ((i_9_) & (!i_8_) & (g9) & (!g29) & (!sk[7]) & (g517)) + ((i_9_) & (!i_8_) & (!g9) & (g29) & (!sk[7]) & (g517)));
	assign g519 = (((!g164) & (!sk[8]) & (!g515) & (!g516) & (g518)) + ((g164) & (!sk[8]) & (!g515) & (g516) & (!g518)) + ((!g164) & (!sk[8]) & (g515) & (!g516) & (g518)) + ((!g164) & (sk[8]) & (g515) & (g516) & (!g518)));
	assign g520 = (((!i_26_) & (!sk[9]) & (!i_29_) & (!i_22_) & (g488)) + ((i_26_) & (!sk[9]) & (!i_29_) & (i_22_) & (!g488)) + ((!i_26_) & (!sk[9]) & (!i_29_) & (!i_22_) & (g488)) + ((!i_26_) & (!sk[9]) & (!i_29_) & (!i_22_) & (g488)));
	assign g521 = (((!i_31_) & (!sk[10]) & (!i_25_) & (!g520) & (g455)) + ((i_31_) & (!sk[10]) & (!i_25_) & (g520) & (!g455)) + ((!i_31_) & (!sk[10]) & (!i_25_) & (g520) & (g455)));
	assign g522 = (((!sk[11]) & (!g84) & (!g277) & (!g443) & (g491) & (!g495)) + ((!sk[11]) & (g84) & (g277) & (!g443) & (g491) & (!g495)) + ((!sk[11]) & (g84) & (!g277) & (!g443) & (!g491) & (g495)) + ((!sk[11]) & (g84) & (!g277) & (g443) & (!g491) & (g495)));
	assign g523 = (((!sk[12]) & (!i_34_) & (!i_26_) & (!i_29_) & (g488)) + ((!sk[12]) & (i_34_) & (!i_26_) & (i_29_) & (!g488)) + ((!sk[12]) & (i_34_) & (!i_26_) & (!i_29_) & (g488)) + ((!sk[12]) & (!i_34_) & (!i_26_) & (!i_29_) & (g488)));
	assign g524 = (((!i_12_) & (!sk[13]) & (!i_2_) & (!g14) & (i_1_)) + ((i_12_) & (!sk[13]) & (!i_2_) & (g14) & (!i_1_)) + ((!i_12_) & (sk[13]) & (!i_2_) & (g14) & (!i_1_)) + ((!i_12_) & (sk[13]) & (!i_2_) & (g14) & (!i_1_)));
	assign g525 = (((!g57) & (!g164) & (!sk[14]) & (!g523) & (g524)) + ((g57) & (!g164) & (!sk[14]) & (g523) & (!g524)) + ((g57) & (!g164) & (!sk[14]) & (g523) & (g524)));
	assign g526 = (((!i_9_) & (i_8_) & (!sk[15]) & (!g9) & (g70) & (!g29)) + ((!i_9_) & (!i_8_) & (!sk[15]) & (!g9) & (g70) & (!g29)) + ((i_9_) & (!i_8_) & (!sk[15]) & (!g9) & (!g70) & (g29)) + ((!i_9_) & (!i_8_) & (!sk[15]) & (!g9) & (g70) & (!g29)) + ((!i_9_) & (!i_8_) & (!sk[15]) & (!g9) & (g70) & (!g29)));
	assign g527 = (((i_28_) & (!sk[16]) & (!i_26_) & (g478)) + ((!i_28_) & (sk[16]) & (!i_26_) & (g478)));
	assign g528 = (((!i_29_) & (!sk[17]) & (!i_9_) & (!i_10_) & (g527)) + ((i_29_) & (!sk[17]) & (!i_9_) & (i_10_) & (!g527)) + ((!i_29_) & (!sk[17]) & (i_9_) & (!i_10_) & (g527)));
	assign g529 = (((!g521) & (!g522) & (!g525) & (g526) & (!sk[18]) & (!g528)) + ((g521) & (!g522) & (!g525) & (!g526) & (!sk[18]) & (g528)) + ((!g521) & (!g522) & (!g525) & (g526) & (!sk[18]) & (!g528)) + ((!g521) & (!g522) & (!g525) & (!g526) & (sk[18]) & (!g528)));
	assign g530 = (((!sk[19]) & (!i_34_) & (!g1) & (!g514) & (g519) & (!g529)) + ((!sk[19]) & (i_34_) & (!g1) & (!g514) & (!g519) & (g529)) + ((sk[19]) & (!i_34_) & (!g1) & (!g514) & (!g519) & (g529)) + ((!sk[19]) & (i_34_) & (!g1) & (!g514) & (!g519) & (g529)) + ((!sk[19]) & (i_34_) & (!g1) & (!g514) & (!g519) & (g529)));
	assign g531 = (((i_24_) & (!i_30_) & (i_32_) & (!g7) & (!g484) & (!g499)) + ((!i_24_) & (i_30_) & (i_32_) & (!g7) & (!g484) & (!g499)) + ((!i_24_) & (!i_30_) & (i_32_) & (!g7) & (!g484) & (!g499)) + ((i_24_) & (!i_30_) & (!i_32_) & (!g7) & (!g484) & (!g499)) + ((!i_24_) & (i_30_) & (!i_32_) & (!g7) & (!g484) & (!g499)) + ((!i_24_) & (!i_30_) & (!i_32_) & (!g7) & (!g484) & (!g499)));
	assign g532 = (((i_33_) & (!i_34_) & (!sk[21]) & (g428)) + ((!i_33_) & (i_34_) & (sk[21]) & (g428)));
	assign g533 = (((!i_33_) & (!sk[22]) & (!i_26_) & (!g84) & (g65) & (!i_38_)) + ((i_33_) & (!sk[22]) & (!i_26_) & (!g84) & (!g65) & (i_38_)) + ((!i_33_) & (!sk[22]) & (!i_26_) & (g84) & (g65) & (i_38_)));
	assign g534 = (((!g1) & (!sk[23]) & (!g70) & (!g532) & (g533)) + ((g1) & (!sk[23]) & (!g70) & (g532) & (!g533)) + ((!g1) & (sk[23]) & (!g70) & (!g532) & (!g533)) + ((!g1) & (sk[23]) & (!g70) & (!g532) & (!g533)) + ((g1) & (!sk[23]) & (g70) & (g532) & (!g533)));
	assign g535 = (((!sk[24]) & (!i_26_) & (g1)) + ((!sk[24]) & (!i_26_) & (g1)));
	assign g536 = (((!g84) & (!g66) & (!sk[25]) & (!i_38_) & (g535) & (!g492)) + ((!g84) & (!g66) & (!sk[25]) & (!i_38_) & (g535) & (g492)) + ((g84) & (!g66) & (!sk[25]) & (!i_38_) & (!g535) & (g492)) + ((g84) & (g66) & (sk[25]) & (i_38_) & (!g535) & (!g492)));
	assign g537 = (((!sk[26]) & (!g478) & (g536)) + ((!sk[26]) & (g478) & (g536)));
	assign g538 = (((!i_24_) & (!i_11_) & (!sk[27]) & (!g456) & (g534) & (!g537)) + ((i_24_) & (!i_11_) & (!sk[27]) & (!g456) & (!g534) & (g537)) + ((!i_24_) & (i_11_) & (sk[27]) & (g456) & (!g534) & (!g537)) + ((!i_24_) & (i_11_) & (sk[27]) & (g456) & (!g534) & (g537)));
	assign g539 = (((!i_28_) & (!i_26_) & (!sk[28]) & (!i_29_) & (i_25_) & (!i_38_)) + ((i_28_) & (!i_26_) & (!sk[28]) & (!i_29_) & (!i_25_) & (i_38_)) + ((!i_28_) & (!i_26_) & (sk[28]) & (!i_29_) & (!i_25_) & (i_38_)));
	assign g540 = (((!g428) & (!g513) & (!g530) & (g531) & (!g538) & (!g539)) + ((!g428) & (!g513) & (!g530) & (!g531) & (!g538) & (!g539)) + ((!g428) & (!g513) & (g530) & (g531) & (!g538) & (!g539)) + ((!g428) & (!g513) & (g530) & (!g531) & (!g538) & (!g539)));
	assign g541 = (((!i_24_) & (i_9_) & (!i_8_) & (g9) & (!i_10_) & (!g29)) + ((!i_24_) & (i_9_) & (!i_8_) & (!g9) & (!i_10_) & (g29)));
	assign g542 = (((!sk[31]) & (!i_33_) & (!g428) & (!g541) & (g514)) + ((!sk[31]) & (!i_33_) & (g428) & (!g541) & (g514)) + ((!sk[31]) & (i_33_) & (!g428) & (g541) & (!g514)) + ((sk[31]) & (!i_33_) & (g428) & (g541) & (!g514)));
	assign g543 = (((!sk[32]) & (!i_9_) & (!g9) & (!i_10_) & (g29)) + ((!sk[32]) & (i_9_) & (!g9) & (i_10_) & (!g29)) + ((!sk[32]) & (i_9_) & (!g9) & (!i_10_) & (g29)) + ((sk[32]) & (i_9_) & (g9) & (!i_10_) & (!g29)));
	assign g544 = (((i_32_) & (!g428) & (!sk[33]) & (g543)) + ((!i_32_) & (g428) & (sk[33]) & (g543)));
	assign g545 = (((!i_30_) & (!i_32_) & (!i_8_) & (!sk[34]) & (g449) & (!g435)) + ((i_30_) & (!i_32_) & (!i_8_) & (!sk[34]) & (!g449) & (g435)) + ((!i_30_) & (!i_32_) & (!i_8_) & (!sk[34]) & (g449) & (g435)) + ((!i_30_) & (!i_32_) & (!i_8_) & (sk[34]) & (!g449) & (g435)));
	assign g546 = (((!g8) & (!g24) & (g478) & (!g466) & (g544) & (!g545)) + ((!g8) & (!g24) & (g478) & (!g466) & (!g544) & (g545)) + ((g8) & (!g24) & (g478) & (g466) & (!g544) & (!g545)));
	assign g547 = (((!sk[36]) & (!i_33_) & (!i_38_) & (!g472) & (g491) & (!g531)) + ((!sk[36]) & (!i_33_) & (!i_38_) & (g472) & (g491) & (!g531)) + ((!sk[36]) & (i_33_) & (!i_38_) & (!g472) & (!g491) & (g531)) + ((sk[36]) & (!i_33_) & (i_38_) & (!g472) & (!g491) & (!g531)));
	assign g548 = (((!sk[37]) & (!i_28_) & (!i_26_) & (!i_30_) & (i_22_) & (!g478)) + ((!sk[37]) & (i_28_) & (!i_26_) & (!i_30_) & (!i_22_) & (g478)) + ((sk[37]) & (!i_28_) & (!i_26_) & (!i_30_) & (!i_22_) & (g478)));
	assign g549 = (((i_33_) & (!sk[38]) & (!g71) & (g428)) + ((!i_33_) & (sk[38]) & (!g71) & (g428)));
	assign g550 = (((!i_22_) & (!g223) & (g548) & (g435) & (!sk[39]) & (!g549)) + ((!i_22_) & (!g223) & (!g548) & (g435) & (!sk[39]) & (!g549)) + ((i_22_) & (!g223) & (!g548) & (!g435) & (!sk[39]) & (g549)) + ((!i_22_) & (g223) & (!g548) & (!g435) & (sk[39]) & (g549)));
	assign g551 = (((!i_33_) & (!sk[40]) & (!i_25_) & (!i_22_) & (i_38_)) + ((i_33_) & (!sk[40]) & (!i_25_) & (i_22_) & (!i_38_)) + ((!i_33_) & (!sk[40]) & (!i_25_) & (!i_22_) & (i_38_)) + ((!i_33_) & (!sk[40]) & (!i_25_) & (!i_22_) & (i_38_)));
	assign g552 = (((!i_26_) & (!i_30_) & (!i_7_) & (!i_32_) & (g488) & (g551)));
	assign g553 = (((!sk[42]) & (i_8_) & (!g550) & (g552)) + ((sk[42]) & (i_8_) & (!g550) & (!g552)) + ((sk[42]) & (!i_8_) & (!g550) & (!g552)));
	assign g554 = (((!i_33_) & (!sk[43]) & (!i_12_) & (!i_25_) & (i_22_) & (!i_38_)) + ((i_33_) & (!sk[43]) & (!i_12_) & (!i_25_) & (!i_22_) & (i_38_)) + ((!i_33_) & (sk[43]) & (i_12_) & (!i_25_) & (!i_22_) & (i_38_)) + ((!i_33_) & (sk[43]) & (i_12_) & (!i_25_) & (!i_22_) & (i_38_)));
	assign g555 = (((!i_24_) & (!i_28_) & (!sk[44]) & (!i_26_) & (g197) & (!g554)) + ((i_24_) & (!i_28_) & (!sk[44]) & (!i_26_) & (!g197) & (g554)) + ((!i_24_) & (!i_28_) & (!sk[44]) & (!i_26_) & (g197) & (g554)));
	assign g556 = (((!i_13_) & (!i_18_) & (!sk[45]) & (!i_19_) & (g555)) + ((i_13_) & (!i_18_) & (!sk[45]) & (i_19_) & (!g555)) + ((!i_13_) & (i_18_) & (!sk[45]) & (i_19_) & (g555)));
	assign g557 = (((i_22_) & (!g474) & (!sk[46]) & (g464)) + ((!i_22_) & (g474) & (sk[46]) & (g464)));
	assign g558 = (((!i_12_) & (!i_13_) & (!sk[47]) & (!i_18_) & (i_11_)) + ((i_12_) & (!i_13_) & (!sk[47]) & (i_18_) & (!i_11_)) + ((i_12_) & (!i_13_) & (!sk[47]) & (i_18_) & (i_11_)));
	assign g559 = (((!sk[48]) & (!i_10_) & (!g553) & (!g556) & (g557) & (!g558)) + ((!sk[48]) & (i_10_) & (!g553) & (!g556) & (g557) & (!g558)) + ((sk[48]) & (i_10_) & (!g553) & (g556) & (!g557) & (!g558)) + ((!sk[48]) & (i_10_) & (!g553) & (!g556) & (!g557) & (g558)) + ((!sk[48]) & (i_10_) & (!g553) & (!g556) & (!g557) & (g558)));
	assign g560 = (((!g57) & (!i_29_) & (!i_8_) & (!sk[49]) & (g96) & (!g449)) + ((!g57) & (!i_29_) & (!i_8_) & (!sk[49]) & (g96) & (!g449)) + ((g57) & (!i_29_) & (!i_8_) & (!sk[49]) & (!g96) & (g449)) + ((g57) & (!i_29_) & (!i_8_) & (!sk[49]) & (!g96) & (g449)));
	assign g561 = (((!sk[50]) & (!i_34_) & (g428)) + ((!sk[50]) & (i_34_) & (g428)));
	assign g562 = (((g479) & (!sk[51]) & (!g561) & (g543)) + ((g479) & (!sk[51]) & (g561) & (g543)));
	assign g563 = (((!sk[52]) & (!i_16_) & (!i_27_) & (!i_32_) & (g96)) + ((!sk[52]) & (!i_16_) & (!i_27_) & (!i_32_) & (g96)) + ((sk[52]) & (!i_16_) & (!i_27_) & (!i_32_) & (!g96)) + ((!sk[52]) & (i_16_) & (!i_27_) & (i_32_) & (!g96)));
	assign g564 = (((!i_28_) & (i_34_) & (i_23_) & (!i_29_) & (!i_22_) & (!g563)) + ((!i_28_) & (i_34_) & (!i_23_) & (!i_29_) & (!i_22_) & (!g563)) + ((!i_28_) & (i_34_) & (!i_23_) & (!i_29_) & (i_22_) & (!g563)));
	assign g565 = (((!i_24_) & (!i_28_) & (!g532) & (!g560) & (g562) & (!g564)) + ((!i_24_) & (!i_28_) & (!g532) & (!g560) & (!g562) & (g564)) + ((!i_24_) & (!i_28_) & (g532) & (g560) & (!g562) & (!g564)));
	assign g566 = (((!g535) & (!g542) & (!g546) & (!g547) & (!g559) & (!g565)) + ((!g535) & (!g542) & (!g546) & (!g547) & (!g559) & (!g565)));
	assign g567 = (((!i_13_) & (!i_3_) & (!sk[56]) & (!i_19_) & (i_22_)) + ((i_13_) & (!i_3_) & (!sk[56]) & (i_19_) & (!i_22_)) + ((!i_13_) & (!i_3_) & (sk[56]) & (i_19_) & (!i_22_)));
	assign g568 = (((!i_13_) & (!i_18_) & (!g12) & (!sk[57]) & (i_22_)) + ((i_13_) & (!i_18_) & (g12) & (!sk[57]) & (!i_22_)) + ((!i_13_) & (i_18_) & (!g12) & (sk[57]) & (!i_22_)));
	assign g569 = (((!g567) & (!sk[58]) & (g568)) + ((!g567) & (sk[58]) & (!g568)));
	assign g570 = (((i_12_) & (!g473) & (!sk[59]) & (g552) & (!g569)) + ((!i_12_) & (!g473) & (!sk[59]) & (!g552) & (g569)) + ((i_12_) & (g473) & (sk[59]) & (!g552) & (!g569)));
	assign g571 = (((!i_12_) & (!i_2_) & (!sk[60]) & (!i_22_) & (g474) & (!g568)) + ((i_12_) & (!i_2_) & (!sk[60]) & (!i_22_) & (g474) & (!g568)) + ((!i_12_) & (!i_2_) & (sk[60]) & (!i_22_) & (!g474) & (g568)) + ((i_12_) & (!i_2_) & (!sk[60]) & (!i_22_) & (!g474) & (g568)));
	assign g572 = (((!sk[61]) & (!i_28_) & (!g70) & (!g527) & (g549) & (!g492)) + ((!sk[61]) & (!i_28_) & (!g70) & (!g527) & (g549) & (!g492)) + ((!sk[61]) & (i_28_) & (!g70) & (!g527) & (!g549) & (g492)) + ((sk[61]) & (!i_28_) & (!g70) & (g527) & (!g549) & (g492)));
	assign g573 = (((!i_12_) & (!i_2_) & (!i_10_) & (!sk[62]) & (i_22_) & (!g572)) + ((i_12_) & (!i_2_) & (!i_10_) & (!sk[62]) & (!i_22_) & (g572)) + ((i_12_) & (!i_2_) & (!i_10_) & (!sk[62]) & (!i_22_) & (g572)) + ((!i_12_) & (!i_2_) & (!i_10_) & (sk[62]) & (!i_22_) & (g572)));
	assign g574 = (((!i_35_) & (!i_26_) & (!i_30_) & (!sk[63]) & (g488) & (!g551)) + ((i_35_) & (!i_26_) & (!i_30_) & (!sk[63]) & (!g488) & (g551)) + ((!i_35_) & (!i_26_) & (!i_30_) & (!sk[63]) & (g488) & (g551)));
	assign g575 = (((!i_13_) & (!sk[64]) & (!i_3_) & (!i_19_) & (g46) & (!g574)) + ((i_13_) & (!sk[64]) & (!i_3_) & (!i_19_) & (!g46) & (g574)) + ((!i_13_) & (!sk[64]) & (!i_3_) & (i_19_) & (g46) & (g574)));
	assign g576 = (((!g473) & (!g555) & (!sk[65]) & (!g571) & (g573) & (!g575)) + ((g473) & (!g555) & (!sk[65]) & (!g571) & (!g573) & (g575)) + ((!g473) & (!g555) & (sk[65]) & (!g571) & (!g573) & (!g575)) + ((!g473) & (!g555) & (sk[65]) & (!g571) & (!g573) & (!g575)));
	assign g577 = (((!sk[66]) & (!i_24_) & (!i_19_) & (!i_25_) & (g534) & (!g536)) + ((!sk[66]) & (i_24_) & (!i_19_) & (!i_25_) & (!g534) & (g536)) + ((sk[66]) & (!i_24_) & (i_19_) & (!i_25_) & (!g534) & (!g536)) + ((!sk[66]) & (!i_24_) & (i_19_) & (!i_25_) & (g534) & (g536)));
	assign g578 = (((!i_24_) & (!g474) & (!g534) & (!sk[67]) & (g537)) + ((i_24_) & (!g474) & (g534) & (!sk[67]) & (!g537)) + ((!i_24_) & (g474) & (!g534) & (!sk[67]) & (g537)) + ((!i_24_) & (g474) & (!g534) & (sk[67]) & (!g537)));
	assign g579 = (((!i_13_) & (!sk[68]) & (!i_3_) & (!g577) & (g578)) + ((!i_13_) & (sk[68]) & (i_3_) & (!g577) & (!g578)) + ((!i_13_) & (sk[68]) & (!i_3_) & (!g577) & (!g578)) + ((i_13_) & (!sk[68]) & (!i_3_) & (g577) & (!g578)));
	assign g580 = (((!sk[69]) & (i_33_) & (!g71) & (i_38_)) + ((sk[69]) & (!i_33_) & (!g71) & (i_38_)));
	assign g581 = (((!g37) & (!g31) & (!g48) & (!sk[70]) & (g580) & (!g685)) + ((g37) & (g31) & (!g48) & (!sk[70]) & (g580) & (!g685)) + ((g37) & (!g31) & (!g48) & (!sk[70]) & (!g580) & (g685)) + ((!g37) & (!g31) & (g48) & (sk[70]) & (!g580) & (!g685)));
	assign g582 = (((!i_32_) & (!sk[71]) & (!i_31_) & (!i_25_) & (g520) & (!g428)) + ((i_32_) & (!sk[71]) & (!i_31_) & (!i_25_) & (!g520) & (g428)) + ((!i_32_) & (!sk[71]) & (!i_31_) & (!i_25_) & (g520) & (g428)));
	assign g583 = (((!i_33_) & (!i_34_) & (!sk[72]) & (!g121) & (g428) & (!g494)) + ((!i_33_) & (i_34_) & (!sk[72]) & (!g121) & (g428) & (!g494)) + ((!i_33_) & (!i_34_) & (!sk[72]) & (g121) & (g428) & (!g494)) + ((i_33_) & (!i_34_) & (!sk[72]) & (!g121) & (!g428) & (g494)) + ((!i_33_) & (i_34_) & (!sk[72]) & (!g121) & (g428) & (g494)));
	assign g584 = (((!i_26_) & (!i_25_) & (!sk[73]) & (!g488) & (g583)) + ((i_26_) & (!i_25_) & (!sk[73]) & (g488) & (!g583)) + ((!i_26_) & (!i_25_) & (!sk[73]) & (g488) & (g583)) + ((!i_26_) & (!i_25_) & (!sk[73]) & (g488) & (g583)));
	assign g585 = (((!sk[74]) & (!i_33_) & (!i_24_) & (!g57) & (g1) & (!g561)) + ((!sk[74]) & (i_33_) & (!i_24_) & (!g57) & (!g1) & (g561)) + ((!sk[74]) & (!i_33_) & (!i_24_) & (g57) & (g1) & (g561)));
	assign g586 = (((!sk[75]) & (!i_28_) & (!g57) & (!i_22_) & (g549) & (!g585)) + ((!sk[75]) & (i_28_) & (!g57) & (!i_22_) & (!g549) & (g585)) + ((sk[75]) & (!i_28_) & (!g57) & (!i_22_) & (!g549) & (!g585)) + ((!sk[75]) & (i_28_) & (!g57) & (!i_22_) & (g549) & (!g585)) + ((!sk[75]) & (!i_28_) & (!g57) & (!i_22_) & (g549) & (!g585)) + ((!sk[75]) & (!i_28_) & (!g57) & (i_22_) & (g549) & (!g585)));
	assign g587 = (((!g57) & (!i_29_) & (!g582) & (g584) & (!sk[76]) & (!g586)) + ((g57) & (!i_29_) & (!g582) & (!g584) & (!sk[76]) & (g586)) + ((!g57) & (!i_29_) & (!g582) & (!g584) & (sk[76]) & (g586)) + ((!g57) & (i_29_) & (!g582) & (!g584) & (sk[76]) & (g586)) + ((!g57) & (!i_29_) & (!g582) & (!g584) & (sk[76]) & (g586)));
	assign g588 = (((!g8) & (!g335) & (!g24) & (!sk[77]) & (g581) & (!g587)) + ((g8) & (!g335) & (!g24) & (!sk[77]) & (g581) & (!g587)) + ((g8) & (!g335) & (!g24) & (!sk[77]) & (!g581) & (g587)) + ((g8) & (g335) & (!g24) & (sk[77]) & (!g581) & (!g587)));
	assign g589 = (((!i_9_) & (!g570) & (!g576) & (g579) & (!sk[78]) & (!g588)) + ((i_9_) & (!g570) & (!g576) & (!g579) & (!sk[78]) & (g588)) + ((!i_9_) & (!g570) & (!g576) & (!g579) & (sk[78]) & (!g588)) + ((!i_9_) & (!g570) & (g576) & (g579) & (!sk[78]) & (!g588)));
	assign g590 = (((!i_16_) & (!sk[79]) & (!i_33_) & (!i_34_) & (g33) & (!g34)) + ((i_16_) & (!sk[79]) & (!i_33_) & (!i_34_) & (!g33) & (g34)) + ((!i_16_) & (!sk[79]) & (i_33_) & (i_34_) & (g33) & (g34)));
	assign g591 = (((!i_33_) & (!i_34_) & (!i_14_) & (g45) & (!sk[80]) & (!g35)) + ((i_33_) & (!i_34_) & (!i_14_) & (!g45) & (!sk[80]) & (g35)) + ((i_33_) & (i_34_) & (i_14_) & (g45) & (!sk[80]) & (g35)));
	assign g592 = (((!i_12_) & (!sk[81]) & (!i_13_) & (!i_14_) & (g590) & (!g591)) + ((i_12_) & (!sk[81]) & (!i_13_) & (!i_14_) & (!g590) & (g591)) + ((!i_12_) & (sk[81]) & (!i_13_) & (!i_14_) & (!g590) & (!g591)) + ((i_12_) & (!sk[81]) & (!i_13_) & (!i_14_) & (g590) & (!g591)) + ((!i_12_) & (!sk[81]) & (i_13_) & (!i_14_) & (g590) & (!g591)) + ((!i_12_) & (!sk[81]) & (!i_13_) & (!i_14_) & (g590) & (!g591)));
	assign g593 = (((i_7_) & (!sk[82]) & (!g70) & (g451)) + ((i_7_) & (sk[82]) & (!g70) & (!g451)) + ((!i_7_) & (sk[82]) & (g70) & (!g451)));
	assign g594 = (((!g66) & (!g60) & (g478) & (!g449) & (g535) & (!g593)) + ((g66) & (g60) & (g478) & (g449) & (!g535) & (!g593)));
	assign g595 = (((!i_26_) & (!i_29_) & (!i_22_) & (!sk[84]) & (g478)) + ((i_26_) & (!i_29_) & (i_22_) & (!sk[84]) & (!g478)) + ((!i_26_) & (i_29_) & (!i_22_) & (sk[84]) & (!g478)) + ((i_26_) & (i_29_) & (!i_22_) & (!sk[84]) & (g478)) + ((!i_26_) & (i_29_) & (i_22_) & (!sk[84]) & (g478)));
	assign g596 = (((!i_7_) & (!i_32_) & (!sk[85]) & (!g9) & (g29)) + ((i_7_) & (!i_32_) & (!sk[85]) & (g9) & (!g29)) + ((!i_7_) & (!i_32_) & (!sk[85]) & (!g9) & (g29)) + ((!i_7_) & (!i_32_) & (sk[85]) & (g9) & (!g29)));
	assign g597 = (((!i_28_) & (!sk[86]) & (!i_34_) & (!i_35_) & (i_26_) & (!g164)) + ((i_28_) & (!sk[86]) & (!i_34_) & (!i_35_) & (!i_26_) & (g164)) + ((!i_28_) & (sk[86]) & (!i_34_) & (!i_35_) & (!i_26_) & (!g164)) + ((!i_28_) & (!sk[86]) & (i_34_) & (!i_35_) & (i_26_) & (!g164)) + ((!i_28_) & (!sk[86]) & (!i_34_) & (i_35_) & (i_26_) & (!g164)));
	assign g598 = (((!i_24_) & (!g2) & (!sk[87]) & (!g595) & (g596) & (!g597)) + ((i_24_) & (!g2) & (!sk[87]) & (!g595) & (!g596) & (g597)) + ((!i_24_) & (!g2) & (!sk[87]) & (!g595) & (g596) & (g597)) + ((!i_24_) & (g2) & (!sk[87]) & (!g595) & (g596) & (g597)));
	assign g599 = (((!i_33_) & (!sk[88]) & (!i_34_) & (!i_29_) & (g96)) + ((i_33_) & (!sk[88]) & (!i_34_) & (i_29_) & (!g96)) + ((!i_33_) & (!sk[88]) & (!i_34_) & (!i_29_) & (g96)) + ((!i_33_) & (!sk[88]) & (i_34_) & (!i_29_) & (g96)));
	assign g600 = (((!i_33_) & (!i_34_) & (!sk[89]) & (!g65) & (g121) & (!g494)) + ((!i_33_) & (!i_34_) & (!sk[89]) & (g65) & (g121) & (!g494)) + ((i_33_) & (!i_34_) & (!sk[89]) & (!g65) & (!g121) & (g494)) + ((!i_33_) & (!i_34_) & (!sk[89]) & (g65) & (g121) & (g494)) + ((!i_33_) & (i_34_) & (sk[89]) & (g65) & (!g121) & (!g494)) + ((!i_33_) & (i_34_) & (sk[89]) & (g65) & (!g121) & (g494)));
	assign g601 = (((!i_26_) & (!i_25_) & (!sk[90]) & (!g488) & (g599) & (!g600)) + ((i_26_) & (!i_25_) & (!sk[90]) & (!g488) & (!g599) & (g600)) + ((!i_26_) & (!i_25_) & (!sk[90]) & (g488) & (g599) & (g600)) + ((!i_26_) & (!i_25_) & (!sk[90]) & (g488) & (g599) & (g600)));
	assign g602 = (((!i_33_) & (!g71) & (!g65) & (g60) & (!sk[91]) & (!g449)) + ((i_33_) & (!g71) & (!g65) & (!g60) & (!sk[91]) & (g449)) + ((!i_33_) & (!g71) & (g65) & (g60) & (!sk[91]) & (g449)));
	assign g603 = (((!g2) & (!sk[92]) & (!g84) & (!g7) & (i_25_)) + ((g2) & (!sk[92]) & (!g84) & (g7) & (!i_25_)) + ((g2) & (!sk[92]) & (g84) & (g7) & (!i_25_)));
	assign g604 = (((i_33_) & (!sk[93]) & (!g2) & (g1)) + ((!i_33_) & (sk[93]) & (g2) & (g1)));
	assign g605 = (((!i_2_) & (!sk[94]) & (!i_30_) & (!g7) & (g604) & (!g548)) + ((!i_2_) & (!sk[94]) & (!i_30_) & (g7) & (g604) & (!g548)) + ((i_2_) & (!sk[94]) & (!i_30_) & (!g7) & (!g604) & (g548)) + ((!i_2_) & (sk[94]) & (!i_30_) & (g7) & (!g604) & (g548)));
	assign g606 = (((!g2) & (!sk[95]) & (!g479) & (!g437) & (g603) & (!g605)) + ((g2) & (!sk[95]) & (!g479) & (!g437) & (!g603) & (g605)) + ((!g2) & (sk[95]) & (!g479) & (!g437) & (!g603) & (!g605)) + ((!g2) & (sk[95]) & (!g479) & (!g437) & (!g603) & (!g605)) + ((!g2) & (sk[95]) & (!g479) & (g437) & (!g603) & (!g605)));
	assign g607 = (((!sk[96]) & (!g592) & (!g598) & (!g601) & (g602) & (!g606)) + ((!sk[96]) & (g592) & (!g598) & (!g601) & (!g602) & (g606)) + ((!sk[96]) & (g592) & (!g598) & (!g601) & (!g602) & (g606)));
	assign g608 = (((!i_32_) & (!sk[97]) & (!g1) & (!g11) & (g32)) + ((i_32_) & (!sk[97]) & (!g1) & (g11) & (!g32)) + ((!i_32_) & (sk[97]) & (g1) & (g11) & (!g32)) + ((!i_32_) & (!sk[97]) & (g1) & (!g11) & (g32)));
	assign g609 = (((!i_33_) & (!g2) & (!sk[98]) & (!g24) & (g608)) + ((i_33_) & (!g2) & (!sk[98]) & (g24) & (!g608)) + ((!i_33_) & (g2) & (!sk[98]) & (!g24) & (g608)));
	assign g610 = (((!i_32_) & (!g11) & (!sk[99]) & (!g32) & (g24)) + ((i_32_) & (!g11) & (!sk[99]) & (g32) & (!g24)) + ((!i_32_) & (g11) & (sk[99]) & (!g32) & (!g24)) + ((!i_32_) & (!g11) & (sk[99]) & (g32) & (!g24)));
	assign g611 = (((!sk[100]) & (i_34_) & (!g1) & (g478)) + ((!sk[100]) & (i_34_) & (g1) & (g478)));
	assign g612 = (((!g82) & (!i_25_) & (g451) & (g604) & (!g610) & (!g611)) + ((!g82) & (!i_25_) & (g451) & (!g604) & (!g610) & (g611)) + ((g82) & (!i_25_) & (g451) & (!g604) & (!g610) & (!g611)) + ((g82) & (!i_25_) & (!g451) & (!g604) & (g610) & (!g611)));
	assign g613 = (((!i_33_) & (!g451) & (!g523) & (g609) & (!sk[102]) & (!g612)) + ((i_33_) & (!g451) & (!g523) & (!g609) & (!sk[102]) & (g612)) + ((i_33_) & (!g451) & (!g523) & (!g609) & (sk[102]) & (!g612)) + ((!i_33_) & (!g451) & (!g523) & (!g609) & (sk[102]) & (!g612)) + ((!i_33_) & (!g451) & (!g523) & (!g609) & (sk[102]) & (!g612)));
	assign g614 = (((!g2) & (!sk[103]) & (!i_7_) & (!g1) & (g70)) + ((g2) & (!sk[103]) & (!i_7_) & (g1) & (!g70)) + ((g2) & (!sk[103]) & (!i_7_) & (g1) & (!g70)));
	assign g615 = (((!i_34_) & (!sk[104]) & (!i_26_) & (!i_29_) & (i_22_) & (!g494)) + ((i_34_) & (!sk[104]) & (!i_26_) & (!i_29_) & (!i_22_) & (g494)) + ((i_34_) & (!sk[104]) & (!i_26_) & (!i_29_) & (!i_22_) & (g494)) + ((!i_34_) & (sk[104]) & (!i_26_) & (!i_29_) & (!i_22_) & (g494)));
	assign g616 = (((!g2) & (!g1) & (!g164) & (g486) & (!g443) & (g615)) + ((!g2) & (g1) & (!g164) & (g486) & (g443) & (!g615)) + ((g2) & (g1) & (!g164) & (g486) & (!g443) & (!g615)));
	assign g617 = (((!i_33_) & (!i_25_) & (!sk[106]) & (!g614) & (g616)) + ((i_33_) & (!i_25_) & (!sk[106]) & (g614) & (!g616)) + ((!i_33_) & (!i_25_) & (sk[106]) & (!g614) & (!g616)) + ((i_33_) & (i_25_) & (!sk[106]) & (g614) & (!g616)));
	assign g618 = (((!i_38_) & (g592) & (!g594) & (!g607) & (!g613) & (!g617)) + ((!i_38_) & (!g592) & (!g594) & (g607) & (g613) & (g617)));
	assign g619 = (((!sk[108]) & (g1) & (!g541) & (g561)) + ((!sk[108]) & (g1) & (g541) & (g561)));
	assign g620 = (((!i_12_) & (!sk[109]) & (!i_9_) & (!i_8_) & (g550)) + ((i_12_) & (!sk[109]) & (!i_9_) & (i_8_) & (!g550)) + ((i_12_) & (!sk[109]) & (i_9_) & (!i_8_) & (g550)));
	assign g621 = (((!g108) & (!g164) & (!g258) & (!sk[110]) & (g619) & (!g620)) + ((g108) & (!g164) & (!g258) & (!sk[110]) & (!g619) & (g620)) + ((g108) & (!g164) & (!g258) & (sk[110]) & (!g619) & (!g620)) + ((!g108) & (!g164) & (!g258) & (sk[110]) & (!g619) & (!g620)) + ((g108) & (g164) & (!g258) & (!sk[110]) & (g619) & (!g620)) + ((!g108) & (g164) & (!g258) & (!sk[110]) & (g619) & (!g620)));
	assign g622 = (((!sk[111]) & (!i_28_) & (!i_22_) & (!g672) & (g621)) + ((!sk[111]) & (i_28_) & (!i_22_) & (!g672) & (g621)) + ((!sk[111]) & (!i_28_) & (!i_22_) & (!g672) & (g621)) + ((!sk[111]) & (!i_28_) & (!i_22_) & (!g672) & (g621)) + ((!sk[111]) & (i_28_) & (!i_22_) & (g672) & (!g621)));
	assign g623 = (((!sk[112]) & (i_24_) & (!g70) & (g498)) + ((sk[112]) & (i_24_) & (!g70) & (!g498)) + ((sk[112]) & (!i_24_) & (g70) & (!g498)));
	assign g624 = (((!g60) & (g456) & (!sk[113]) & (!g532) & (g577) & (!g623)) + ((!g60) & (!g456) & (!sk[113]) & (!g532) & (g577) & (!g623)) + ((g60) & (!g456) & (!sk[113]) & (!g532) & (!g577) & (g623)) + ((g60) & (!g456) & (sk[113]) & (g532) & (!g577) & (!g623)));
	assign g625 = (((!sk[114]) & (!i_12_) & (!i_13_) & (!i_18_) & (i_19_) & (!i_10_)) + ((!sk[114]) & (i_12_) & (!i_13_) & (!i_18_) & (!i_19_) & (i_10_)) + ((!sk[114]) & (i_12_) & (!i_13_) & (i_18_) & (i_19_) & (i_10_)));
	assign g626 = (((!i_10_) & (!g464) & (!g553) & (!sk[115]) & (g569) & (!g625)) + ((!i_10_) & (!g464) & (!g553) & (sk[115]) & (!g569) & (g625)) + ((i_10_) & (!g464) & (!g553) & (!sk[115]) & (!g569) & (g625)) + ((i_10_) & (g464) & (!g553) & (sk[115]) & (!g569) & (!g625)));
	assign g627 = (((!i_34_) & (!g1) & (!g70) & (!sk[116]) & (g504)) + ((i_34_) & (!g1) & (g70) & (!sk[116]) & (!g504)) + ((i_34_) & (g1) & (g70) & (!sk[116]) & (g504)));
	assign g628 = (((!i_14_) & (!sk[117]) & (!g86) & (!g143) & (g627)) + ((i_14_) & (!sk[117]) & (!g86) & (g143) & (!g627)) + ((!i_14_) & (sk[117]) & (!g86) & (!g143) & (!g627)) + ((!i_14_) & (sk[117]) & (!g86) & (!g143) & (!g627)) + ((i_14_) & (!sk[117]) & (g86) & (g143) & (!g627)));
	assign g629 = (((!i_24_) & (!i_28_) & (!i_26_) & (!sk[118]) & (g65) & (!i_10_)) + ((i_24_) & (!i_28_) & (!i_26_) & (!sk[118]) & (!g65) & (i_10_)) + ((!i_24_) & (!i_28_) & (!i_26_) & (!sk[118]) & (g65) & (!i_10_)));
	assign g630 = (((!sk[119]) & (!i_9_) & (!g29) & (!g551) & (g629)) + ((!sk[119]) & (i_9_) & (!g29) & (g551) & (!g629)) + ((!sk[119]) & (i_9_) & (g29) & (g551) & (g629)));
	assign g631 = (((!i_7_) & (!i_3_) & (!i_18_) & (i_11_) & (!i_19_) & (!i_8_)) + ((!i_7_) & (!i_3_) & (i_18_) & (i_11_) & (!i_19_) & (!i_8_)) + ((!i_7_) & (!i_3_) & (!i_18_) & (!i_11_) & (i_19_) & (!i_8_)));
	assign g632 = (((!i_12_) & (!g24) & (!sk[121]) & (!g140) & (g551) & (!g631)) + ((i_12_) & (!g24) & (!sk[121]) & (!g140) & (!g551) & (g631)) + ((i_12_) & (g24) & (!sk[121]) & (g140) & (g551) & (g631)));
	assign g633 = (((!i_12_) & (!i_2_) & (!i_22_) & (!sk[122]) & (g495)) + ((i_12_) & (!i_2_) & (i_22_) & (!sk[122]) & (!g495)) + ((i_12_) & (!i_2_) & (!i_22_) & (!sk[122]) & (g495)) + ((!i_12_) & (!i_2_) & (!i_22_) & (!sk[122]) & (g495)));
	assign g634 = (((!sk[123]) & (!i_33_) & (!g140) & (!i_25_) & (g428) & (!g633)) + ((!sk[123]) & (i_33_) & (!g140) & (!i_25_) & (!g428) & (g633)) + ((!sk[123]) & (!i_33_) & (g140) & (!i_25_) & (g428) & (g633)) + ((!sk[123]) & (!i_33_) & (g140) & (!i_25_) & (g428) & (g633)));
	assign g635 = (((!sk[124]) & (!g90) & (!g70) & (!g121) & (g634)) + ((!sk[124]) & (g90) & (!g70) & (g121) & (!g634)) + ((sk[124]) & (!g90) & (!g70) & (!g121) & (!g634)) + ((sk[124]) & (!g90) & (!g70) & (!g121) & (!g634)) + ((!sk[124]) & (g90) & (!g70) & (g121) & (!g634)));
	assign g636 = (((!i_12_) & (!i_2_) & (!g12) & (i_8_) & (!sk[125]) & (!g456)) + ((i_12_) & (!i_2_) & (!g12) & (!i_8_) & (!sk[125]) & (g456)) + ((i_12_) & (!i_2_) & (!g12) & (!i_8_) & (!sk[125]) & (g456)) + ((!i_12_) & (!i_2_) & (!g12) & (!i_8_) & (sk[125]) & (g456)));
	assign g637 = (((!i_9_) & (!g46) & (!g474) & (!sk[126]) & (g574) & (!g636)) + ((!i_9_) & (!g46) & (!g474) & (!sk[126]) & (g574) & (g636)) + ((i_9_) & (!g46) & (!g474) & (!sk[126]) & (!g574) & (g636)) + ((i_9_) & (g46) & (g474) & (!sk[126]) & (g574) & (!g636)));
	assign g638 = (((!i_13_) & (!sk[127]) & (!i_9_) & (!g164) & (g488) & (!g428)) + ((i_13_) & (!sk[127]) & (!i_9_) & (!g164) & (!g488) & (g428)) + ((!i_13_) & (!sk[127]) & (i_9_) & (!g164) & (g488) & (g428)));
	assign g639 = (((!i_34_) & (!i_26_) & (!i_30_) & (i_29_) & (!sk[0]) & (!i_8_)) + ((i_34_) & (!i_26_) & (!i_30_) & (!i_29_) & (!sk[0]) & (i_8_)) + ((i_34_) & (!i_26_) & (!i_30_) & (!i_29_) & (sk[0]) & (!i_8_)) + ((!i_34_) & (!i_26_) & (!i_30_) & (!i_29_) & (sk[0]) & (!i_8_)));
	assign g640 = (((!sk[1]) & (!i_34_) & (!i_26_) & (!i_32_) & (i_29_) & (!i_22_)) + ((!sk[1]) & (i_34_) & (!i_26_) & (!i_32_) & (!i_29_) & (i_22_)) + ((sk[1]) & (i_34_) & (!i_26_) & (!i_32_) & (!i_29_) & (!i_22_)) + ((sk[1]) & (!i_34_) & (!i_26_) & (!i_32_) & (!i_29_) & (!i_22_)) + ((!sk[1]) & (!i_34_) & (!i_26_) & (!i_32_) & (i_29_) & (!i_22_)));
	assign g641 = (((!sk[2]) & (!g371) & (!g524) & (!g638) & (g639) & (!g640)) + ((!sk[2]) & (g371) & (!g524) & (g638) & (g639) & (!g640)) + ((!sk[2]) & (g371) & (!g524) & (!g638) & (!g639) & (g640)) + ((!sk[2]) & (g371) & (g524) & (g638) & (!g639) & (g640)));
	assign g642 = (((!i_33_) & (!g486) & (!g520) & (i_38_) & (!sk[3]) & (!g641)) + ((i_33_) & (!g486) & (!g520) & (!i_38_) & (!sk[3]) & (g641)) + ((!i_33_) & (!g486) & (!g520) & (!i_38_) & (sk[3]) & (!g641)) + ((i_33_) & (!g486) & (!g520) & (!i_38_) & (sk[3]) & (!g641)) + ((!i_33_) & (!g486) & (!g520) & (!i_38_) & (sk[3]) & (!g641)) + ((!i_33_) & (!g486) & (!g520) & (!i_38_) & (sk[3]) & (!g641)));
	assign g643 = (((!g630) & (!sk[4]) & (!g632) & (!g635) & (g637) & (!g642)) + ((g630) & (!sk[4]) & (!g632) & (!g635) & (!g637) & (g642)) + ((!g630) & (sk[4]) & (!g632) & (g635) & (!g637) & (g642)));
	assign g644 = (((!i_31_) & (!sk[5]) & (!g520) & (!g429) & (g455)) + ((i_31_) & (!sk[5]) & (!g520) & (g429) & (!g455)) + ((!i_31_) & (!sk[5]) & (g520) & (g429) & (g455)));
	assign g645 = (((!sk[6]) & (g37) & (!g549) & (g543)) + ((!sk[6]) & (g37) & (g549) & (g543)));
	assign g646 = (((!i_28_) & (!i_2_) & (!i_22_) & (!g197) & (g596) & (g580)) + ((!i_28_) & (!i_2_) & (!i_22_) & (g197) & (!g596) & (g580)));
	assign g647 = (((!i_2_) & (!i_9_) & (!sk[8]) & (!g473) & (g567)) + ((i_2_) & (!i_9_) & (!sk[8]) & (g473) & (!g567)) + ((!i_2_) & (i_9_) & (!sk[8]) & (g473) & (g567)));
	assign g648 = (((!sk[9]) & (!i_27_) & (!g71) & (!g88) & (i_22_)) + ((!sk[9]) & (i_27_) & (!g71) & (g88) & (!i_22_)) + ((!sk[9]) & (i_27_) & (!g71) & (g88) & (!i_22_)));
	assign g649 = (((!sk[10]) & (!i_33_) & (!i_14_) & (!g121) & (g647) & (!g648)) + ((!sk[10]) & (i_33_) & (!i_14_) & (!g121) & (!g647) & (g648)) + ((sk[10]) & (!i_33_) & (!i_14_) & (!g121) & (!g647) & (!g648)) + ((sk[10]) & (!i_33_) & (!i_14_) & (!g121) & (!g647) & (!g648)) + ((sk[10]) & (!i_33_) & (!i_14_) & (!g121) & (!g647) & (!g648)));
	assign g650 = (((!g644) & (!g645) & (!g662) & (g646) & (!sk[11]) & (!g649)) + ((g644) & (!g645) & (!g662) & (!g646) & (!sk[11]) & (g649)) + ((!g644) & (!g645) & (!g662) & (!g646) & (sk[11]) & (g649)));
	assign g651 = (((!i_7_) & (!sk[12]) & (!i_32_) & (!g443) & (g435) & (!g580)) + ((!i_7_) & (!sk[12]) & (!i_32_) & (g443) & (g435) & (!g580)) + ((i_7_) & (!sk[12]) & (!i_32_) & (!g443) & (!g435) & (g580)) + ((!i_7_) & (sk[12]) & (!i_32_) & (!g443) & (!g435) & (g580)));
	assign g652 = (((!i_33_) & (!g71) & (!sk[13]) & (!g84) & (g465) & (!g651)) + ((i_33_) & (!g71) & (!sk[13]) & (!g84) & (!g465) & (g651)) + ((!i_33_) & (!g71) & (sk[13]) & (g84) & (!g465) & (g651)) + ((!i_33_) & (!g71) & (!sk[13]) & (g84) & (g465) & (!g651)));
	assign g653 = (((!sk[14]) & (g2) & (!i_29_) & (i_22_)) + ((sk[14]) & (g2) & (!i_29_) & (!i_22_)));
	assign g654 = (((!i_28_) & (!i_26_) & (!g504) & (g507) & (!sk[15]) & (!g653)) + ((!i_28_) & (!i_26_) & (!g504) & (g507) & (!sk[15]) & (g653)) + ((i_28_) & (!i_26_) & (!g504) & (!g507) & (!sk[15]) & (g653)) + ((!i_28_) & (!i_26_) & (g504) & (g507) & (!sk[15]) & (!g653)));
	assign g655 = (((!i_10_) & (!i_22_) & (!g471) & (!sk[16]) & (g652) & (!g654)) + ((i_10_) & (!i_22_) & (!g471) & (!sk[16]) & (!g652) & (g654)) + ((i_10_) & (!i_22_) & (!g471) & (sk[16]) & (!g652) & (!g654)) + ((!i_10_) & (i_22_) & (!g471) & (sk[16]) & (!g652) & (!g654)) + ((!i_10_) & (!i_22_) & (!g471) & (sk[16]) & (!g652) & (!g654)));
	assign g656 = (((!i_9_) & (!sk[17]) & (!i_3_) & (!i_8_) & (g574)) + ((i_9_) & (!sk[17]) & (!i_3_) & (i_8_) & (!g574)) + ((i_9_) & (!sk[17]) & (!i_3_) & (!i_8_) & (g574)));
	assign g657 = (((i_3_) & (!i_8_) & (!i_10_) & (!g550) & (!g552) & (!g656)) + ((!i_3_) & (!i_8_) & (!i_10_) & (!g550) & (!g552) & (!g656)) + ((!i_3_) & (i_8_) & (!i_10_) & (!g550) & (!g552) & (!g656)) + ((!i_3_) & (!i_8_) & (!i_10_) & (!g550) & (!g552) & (!g656)));
	assign g658 = (((!i_12_) & (!i_13_) & (!sk[19]) & (!i_11_) & (i_19_) & (!g657)) + ((i_12_) & (!i_13_) & (!sk[19]) & (!i_11_) & (!i_19_) & (g657)) + ((i_12_) & (!i_13_) & (!sk[19]) & (!i_11_) & (i_19_) & (!g657)) + ((i_12_) & (!i_13_) & (sk[19]) & (i_11_) & (!i_19_) & (!g657)));
	assign g659 = (((!g628) & (!sk[20]) & (!g643) & (!g650) & (g655) & (!g658)) + ((g628) & (!sk[20]) & (!g643) & (!g650) & (!g655) & (g658)) + ((g628) & (!sk[20]) & (g643) & (g650) & (g655) & (!g658)));
	assign g660 = (((!g618) & (!g622) & (!sk[21]) & (!g624) & (g626) & (!g659)) + ((g618) & (!g622) & (!sk[21]) & (!g624) & (!g626) & (g659)) + ((g618) & (g622) & (!sk[21]) & (!g624) & (!g626) & (g659)));
	assign g661 = (((g477) & (!g510) & (g540) & (g566) & (g589) & (g660)));
	assign g662 = (((!sk[23]) & (!g663) & (g664)) + ((sk[23]) & (!g663) & (!g664)));
	assign g663 = (((!sk[24]) & (!g2) & (g665)) + ((!sk[24]) & (!g2) & (g665)));
	assign g664 = (((!sk[25]) & (!g2) & (g666)) + ((!sk[25]) & (g2) & (g666)));
	assign g665 = (((i_31_) & (!sk[26]) & (g669)) + ((!i_31_) & (!sk[26]) & (g669)));
	assign g666 = (((!g667) & (!sk[27]) & (g668)) + ((!g667) & (sk[27]) & (!g668)));
	assign g667 = (((!i_31_) & (!sk[28]) & (g670)) + ((!i_31_) & (!sk[28]) & (g670)));
	assign g668 = (((!sk[29]) & (!i_31_) & (g671)) + ((!sk[29]) & (i_31_) & (g671)));
	assign g669 = (((g90) & (!sk[30]) & (!g71) & (i_28_)) + ((g90) & (sk[30]) & (!g71) & (!i_28_)));
	assign g670 = (((!g90) & (!sk[31]) & (!i_29_) & (!g70) & (i_28_)) + ((g90) & (!sk[31]) & (!i_29_) & (g70) & (!i_28_)) + ((g90) & (!sk[31]) & (!i_29_) & (g70) & (!i_28_)));
	assign g671 = (((!g90) & (!i_29_) & (!sk[32]) & (!g71) & (i_28_)) + ((g90) & (!i_29_) & (!sk[32]) & (g71) & (!i_28_)) + ((g90) & (!i_29_) & (sk[32]) & (!g71) & (!i_28_)) + ((g90) & (!i_29_) & (!sk[32]) & (g71) & (!i_28_)));
	assign g672 = (((!g673) & (!sk[33]) & (g674)) + ((!g673) & (sk[33]) & (!g674)));
	assign g673 = (((!sk[34]) & (!g90) & (g675)) + ((!sk[34]) & (!g90) & (g675)));
	assign g674 = (((!sk[35]) & (!g90) & (g678)) + ((!sk[35]) & (g90) & (g678)));
	assign g675 = (((!sk[36]) & (!g676) & (g677)) + ((sk[36]) & (!g676) & (!g677)));
	assign g676 = (((!sk[37]) & (!i_34_) & (g681)) + ((!sk[37]) & (!i_34_) & (g681)));
	assign g677 = (((i_34_) & (!sk[38]) & (g682)) + ((!i_34_) & (!sk[38]) & (g682)));
	assign g678 = (((!sk[39]) & (!g679) & (g680)) + ((sk[39]) & (!g679) & (!g680)));
	assign g679 = (((!sk[40]) & (!i_34_) & (g683)) + ((!sk[40]) & (!i_34_) & (g683)));
	assign g680 = (((!sk[41]) & (!i_34_) & (g684)) + ((!sk[41]) & (i_34_) & (g684)));
	assign g681 = (((i_14_) & (i_33_) & (!sk[42]) & (i_35_)) + ((i_14_) & (!i_33_) & (!sk[42]) & (i_35_)));
	assign g682 = (((!sk[43]) & (i_14_) & (!i_33_) & (i_24_)) + ((sk[43]) & (i_14_) & (i_33_) & (!i_24_)));
	assign g683 = (((!i_14_) & (!i_33_) & (!sk[44]) & (!g86) & (i_35_)) + ((!i_14_) & (!i_33_) & (!sk[44]) & (g86) & (i_35_)) + ((i_14_) & (!i_33_) & (!sk[44]) & (g86) & (!i_35_)) + ((i_14_) & (i_33_) & (!sk[44]) & (!g86) & (i_35_)));
	assign g684 = (((i_14_) & (!i_33_) & (!sk[45]) & (i_24_)) + ((i_14_) & (i_33_) & (sk[45]) & (!i_24_)));
	assign g685 = (((!g686) & (!sk[46]) & (g687)) + ((!g686) & (sk[46]) & (!g687)));
	assign g686 = (((!i_33_) & (!sk[47]) & (g688)) + ((!i_33_) & (!sk[47]) & (g688)));
	assign g687 = (((!sk[48]) & (!i_33_) & (g691)) + ((!sk[48]) & (i_33_) & (g691)));
	assign g688 = (((!sk[49]) & (!g689) & (g690)) + ((sk[49]) & (!g689) & (!g690)));
	assign g689 = (((!i_34_) & (!sk[50]) & (g693)) + ((!i_34_) & (!sk[50]) & (g693)));
	assign g690 = (((i_34_) & (!sk[51]) & (g694)) + ((!i_34_) & (!sk[51]) & (g694)));
	assign g691 = (((!sk[52]) & (!i_34_) & (g692)) + ((sk[52]) & (i_34_) & (!g692)));
	assign g692 = (((i_34_) & (!sk[53]) & (g695)) + ((!i_34_) & (!sk[53]) & (g695)));
	assign g693 = (((!g428) & (!sk[54]) & (!g60) & (!i_26_) & (i_24_)) + ((!g428) & (sk[54]) & (!g60) & (!i_26_) & (!i_24_)) + ((!g428) & (sk[54]) & (!g60) & (!i_26_) & (!i_24_)) + ((g428) & (!sk[54]) & (!g60) & (i_26_) & (!i_24_)));
	assign g694 = (((!g428) & (sk[55]) & (!g60) & (!i_24_)) + ((!g428) & (sk[55]) & (!g60) & (!i_24_)) + ((g428) & (!sk[55]) & (!g60) & (i_24_)));
	assign g695 = (((!sk[56]) & (!g428) & (!g60) & (!i_25_) & (i_24_)) + ((sk[56]) & (!g428) & (!g60) & (!i_25_) & (!i_24_)) + ((sk[56]) & (!g428) & (!g60) & (!i_25_) & (!i_24_)) + ((!sk[56]) & (g428) & (!g60) & (i_25_) & (!i_24_)));
	assign g696 = (((!sk[57]) & (!g475) & (g697)) + ((!sk[57]) & (g475) & (g697)));
	assign g697 = (((!sk[58]) & (!g698) & (g699)) + ((sk[58]) & (!g698) & (!g699)));
	assign g698 = (((!i_34_) & (!sk[59]) & (g700)) + ((!i_34_) & (!sk[59]) & (g700)));
	assign g699 = (((!sk[60]) & (!i_34_) & (g701)) + ((!sk[60]) & (i_34_) & (g701)));
	assign g700 = (((sk[61]) & (!i_20_) & (!g88) & (!i_35_) & (!i_21_)) + ((!sk[61]) & (!i_20_) & (!g88) & (!i_35_) & (i_21_)) + ((!sk[61]) & (i_20_) & (!g88) & (i_35_) & (!i_21_)) + ((sk[61]) & (!i_20_) & (!g88) & (!i_35_) & (!i_21_)) + ((sk[61]) & (!i_20_) & (!g88) & (!i_35_) & (!i_21_)));
	assign g701 = (((!i_20_) & (!g88) & (sk[62]) & (!i_24_) & (!i_21_)) + ((i_20_) & (!g88) & (!sk[62]) & (i_24_) & (!i_21_)) + ((!i_20_) & (!g88) & (!sk[62]) & (!i_24_) & (i_21_)) + ((!i_20_) & (!g88) & (sk[62]) & (!i_24_) & (!i_21_)) + ((!i_20_) & (!g88) & (!sk[62]) & (i_24_) & (i_21_)));
	assign g702 = (((!sk[63]) & (!g703) & (g704)) + ((sk[63]) & (!g703) & (!g704)));
	assign g703 = (((!sk[64]) & (!g3) & (g705)) + ((!sk[64]) & (!g3) & (g705)));
	assign g704 = (((!sk[65]) & (!g3) & (g706)) + ((!sk[65]) & (g3) & (g706)));
	assign g705 = (((i_34_) & (!sk[66]) & (g709)) + ((!i_34_) & (!sk[66]) & (g709)));
	assign g706 = (((!g707) & (!sk[67]) & (g708)) + ((!g707) & (sk[67]) & (!g708)));
	assign g707 = (((!i_34_) & (!sk[68]) & (g710)) + ((!i_34_) & (!sk[68]) & (g710)));
	assign g708 = (((!sk[69]) & (!i_34_) & (g711)) + ((!sk[69]) & (i_34_) & (g711)));
	assign g709 = (((!sk[70]) & (!g5) & (!i_31_) & (!i_28_) & (i_21_)) + ((!sk[70]) & (g5) & (!i_31_) & (i_28_) & (!i_21_)) + ((!sk[70]) & (!g5) & (i_31_) & (!i_28_) & (i_21_)));
	assign g710 = (((i_31_) & (i_35_) & (!sk[71]) & (i_21_)) + ((i_31_) & (!i_35_) & (!sk[71]) & (i_21_)));
	assign g711 = (((!g5) & (!sk[72]) & (!i_31_) & (!i_28_) & (i_21_)) + ((g5) & (!sk[72]) & (!i_31_) & (i_28_) & (!i_21_)) + ((!g5) & (!sk[72]) & (i_31_) & (!i_28_) & (i_21_)));
	assign g712 = (((!sk[73]) & (!i_31_) & (g713)) + ((sk[73]) & (i_31_) & (!g713)));
	assign g713 = (((i_31_) & (!sk[74]) & (g714)) + ((!i_31_) & (!sk[74]) & (g714)));
	assign g714 = (((!sk[75]) & (!g715) & (g716)) + ((sk[75]) & (!g715) & (!g716)));
	assign g715 = (((!sk[76]) & (!i_34_) & (g717)) + ((!sk[76]) & (!i_34_) & (g717)));
	assign g716 = (((!sk[77]) & (!i_34_) & (g718)) + ((!sk[77]) & (i_34_) & (g718)));
	assign g717 = (((!g108) & (!sk[78]) & (!g34) & (!i_35_) & (i_28_)) + ((!g108) & (!sk[78]) & (!g34) & (!i_35_) & (i_28_)) + ((!g108) & (!sk[78]) & (!g34) & (!i_35_) & (i_28_)) + ((g108) & (!sk[78]) & (!g34) & (i_35_) & (!i_28_)) + ((g108) & (sk[78]) & (!g34) & (!i_35_) & (!i_28_)) + ((g108) & (!sk[78]) & (!g34) & (i_35_) & (!i_28_)));
	assign g718 = (((g108) & (sk[79]) & (!g21) & (!i_28_)) + ((g108) & (!sk[79]) & (!g21) & (i_28_)) + ((!g108) & (sk[79]) & (!g21) & (i_28_)));

endmodule