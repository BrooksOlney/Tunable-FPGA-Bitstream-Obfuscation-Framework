module ks_alu4x8xv (i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_, o_1_, o_2_, o_0_, o_7_, o_5_, o_6_, o_3_, o_4_);

	input i_9_;
	input i_10_;
	input i_7_;
	input i_8_;
	input i_5_;
	input i_6_;
	input i_3_;
	input i_13_;
	input i_4_;
	input i_12_;
	input i_1_;
	input i_11_;
	input i_2_;
	input i_0_;
	output o_1_;
	output o_2_;
	output o_0_;
	output o_7_;
	output o_5_;
	output o_6_;
	output o_3_;
	output o_4_;

	wire [15 : 0] sk /* synthesis noprune */;

	lut_sub lut_3 ({sk[0], i_9_, i_10_, i_8_, i_3_, i_13_, i_4_, i_12_, i_11_}, o_1_);
	defparam lut_3.LUT_SIZE = 9;
	defparam lut_3.mask = 512'h33ff33ff33ff33ff3fff3fff3fff3fffffffffffffffffffffffffffffffffffa5aa0f00c3cc0f00a5aaf0ffc3cc0f00a5aa0f00c3ccf0ffa5aaf0ffc3ccf0ff;

	lut_sub lut_30 ({sk[1], n_n878, x6520x, x6521x, n_n872, x6529x}, o_2_);
	defparam lut_30.LUT_SIZE = 6;
	defparam lut_30.mask = 64'h1115ffff7fffffff;

	lut_sub lut_36 ({sk[2], i_9_, i_10_, i_8_, i_3_, i_2_, x327x, x6536x, x6537x}, o_0_);
	defparam lut_36.LUT_SIZE = 9;
	defparam lut_36.mask = 512'h33ff33ff33ff33ff3fff3fff3fff3fffffffffffffffffffffffffffffffffff77777777777777777f7f7f7f77777777777777777777ffff7fffffff77ffffff;

	lut_sub lut_43 ({sk[3], x6830x, x6704x, x6705x, x6792x, n_n1231, n_n1233}, o_7_);
	defparam lut_43.LUT_SIZE = 7;
	defparam lut_43.mask = 128'h0303ffffffffffff7fffffffffffffff;

	lut_sub lut_50 ({sk[4], x6950x, n_n1119, n_n1107, n_n1114, x6947x}, o_5_);
	defparam lut_50.LUT_SIZE = 6;
	defparam lut_50.mask = 64'h1115ffff7fffffff;

	lut_sub lut_56 ({sk[5], n_n1185, x6975x, x6991x, x6992x, n_n1187, x6999x}, o_6_);
	defparam lut_56.LUT_SIZE = 7;
	defparam lut_56.mask = 128'h0303ffffffffffff7fffffffffffffff;

	lut_sub lut_63 ({sk[6], n_n908, n_n906, x7065x, x7075x}, o_3_);
	defparam lut_63.LUT_SIZE = 5;
	defparam lut_63.mask = 32'h07ff7fff;

	lut_sub lut_68 ({sk[7], i_7_, x7341x, x7245x, x711x, x7179x, n_n986, x7242x, x7337x}, o_4_);
	defparam lut_68.LUT_SIZE = 9;
	defparam lut_68.mask = 512'h33ff33ff33ff33ff3fff3fff3fff3fffffffffffffffffffffffffffffffffff7fff7fffffffffffffffffffffffffff7fffffffffffffffffffffffffffffff;

	lut_sub lut_76 ({sk[8], i_8_, i_11_, x384x, x385x, x1822x, x1826x, x7983x}, n_n878);
	defparam lut_76.LUT_SIZE = 8;
	defparam lut_76.mask = 256'h3333ffff3333ffffffffffffffffffffbfbfbfbfbfffffffbfbfbfbfbfbfffff;

	lut_sub lut_82 ({sk[9], i_10_, i_6_, i_3_, i_1_, i_2_, i_0_, x665x, x7982x}, x6520x);
	defparam lut_82.LUT_SIZE = 9;
	defparam lut_82.mask = 512'h33ff33ff33ff33ff3fff3fff3fff3fffffffffffffffffffffffffffffffffffaaaaaaabaaaaaaafaaaaaaabaaaaaaafaaaaafafaaaaafafaaaaaaabaaaaaaaf;

	lut_sub lut_87 ({sk[10], i_11_, x663x, x6513x, x1805x, x1814x, x6505x, x7981x}, x6521x);
	defparam lut_87.LUT_SIZE = 8;
	defparam lut_87.mask = 256'h3333ffff3333ffffffffffffffffffffbfffffffbfffffffbfffffffffffffff;

	lut_sub lut_94 ({sk[11], i_9_, i_10_, i_5_, i_12_, i_1_, x683x, x6526x, x6527x}, n_n872);
	defparam lut_94.LUT_SIZE = 9;
	defparam lut_94.mask = 512'h33ff33ff33ff33ff3fff3fff3fff3fffffffffffffffffffffffffffffffffff7777777777777f7f7777777777777f7f7777777777777f7f7777777777777fff;

	lut_sub lut_99 ({sk[12], i_5_, x648x, x1832x, x1841x, x6491x, x6496x, x7980x}, x6529x);
	defparam lut_99.LUT_SIZE = 8;
	defparam lut_99.mask = 256'h3333ffff3333ffffffffffffffffffffbfffffffffffffffbfffffffbfffffff;

	lut_sub lut_106 ({sk[13], i_6_, i_3_, i_2_, i_0_}, x327x);
	defparam lut_106.LUT_SIZE = 5;
	defparam lut_106.mask = 32'h07ff0100;

	lut_sub lut_108 ({sk[14], i_9_, i_10_, i_8_, i_5_, i_6_, i_3_, i_1_, i_0_}, x6536x);
	defparam lut_108.LUT_SIZE = 9;
	defparam lut_108.mask = 512'h33ff33ff33ff33ff3fff3fff3fff3fffffffffffffffffffffffffffffffffff00000000000000003f0f3f0f3300330000005555000055553f3f7f7f33337777;

	lut_sub lut_113 ({sk[15], i_9_, i_10_, i_7_, i_5_, i_6_, i_1_, i_2_, i_0_}, x6537x);
	defparam lut_113.LUT_SIZE = 9;
	defparam lut_113.mask = 512'h33ff33ff33ff33ff3fff3fff3fff3fffffffffffffffffffffffffffffffffff00000000000000007777333355550000000f000f333f333f777f333f777f333f;

	lut_sub lut_118 ({sk[0], n_n1226, n_n1223, x6823x, x6824x, x6825x}, x6830x);
	defparam lut_118.LUT_SIZE = 6;
	defparam lut_118.mask = 64'h7777777f7fffffff;

	lut_sub lut_124 ({sk[1], n_n1250, x1623x, x6652x, x6658x, x6659x, x1595x, x6666x}, x6704x);
	defparam lut_124.LUT_SIZE = 8;
	defparam lut_124.mask = 256'h333333333333ffffffffffffffffffff7fffffffffffffffffffffffffffffff;

	lut_sub lut_132 ({sk[2], n_n1248, x1584x, x6678x, x1570x, x6683x, x1547x, x1564x, x6693x}, x6705x);
	defparam lut_132.LUT_SIZE = 9;
	defparam lut_132.mask = 512'h0055ffff035fffff0055ffff035fffff0055ffff035fffff0055ffff035fffff7fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;

	lut_sub lut_141 ({sk[3], i_8_, x6730x, x6731x, x1511x, x6738x, x575x, x6789x}, x6792x);
	defparam lut_141.LUT_SIZE = 8;
	defparam lut_141.mask = 256'h333333333333ffffffffffffffffffff7fffffffffffffff5fffffffffffffff;

	lut_sub lut_148 ({sk[4], i_9_, i_13_, i_11_, x477x, x6746x, n_n1259, x523x, x6758x}, n_n1231);
	defparam lut_148.LUT_SIZE = 9;
	defparam lut_148.mask = 512'h0055ffff035fffff0055ffff035fffff0055ffff035fffff0055ffff035fffff5fff5fff7fffffff5fff5fff5fff5fff5fff5fff5fff5fff5fff5fff5fff5fff;

	lut_sub lut_154 ({sk[5], i_7_, i_6_, n_n1265, x6766x, x6767x, x611x, x6779x, x6780x}, n_n1233);
	defparam lut_154.LUT_SIZE = 9;
	defparam lut_154.mask = 512'h0055ffff035fffff0055ffff035fffff0055ffff035fffff0055ffff035fffff7fffffffffffffff77ffffffffffffff77ffffffffffffff77ffffffffffffff;

	lut_sub lut_161 ({sk[6], i_6_, n_n1121, x6841x, x6869x, x444x, n_n1116, n_n1118}, x6950x);
	defparam lut_161.LUT_SIZE = 8;
	defparam lut_161.mask = 256'h333333333333ffffffffffffffffffff7fffffffffffffff77ffffffffffffff;

	lut_sub lut_168 ({sk[7], i_6_, n_n787, x448x, x1355x, x1356x, x1351x, x1352x, x1354x}, n_n1119);
	defparam lut_168.LUT_SIZE = 9;
	defparam lut_168.mask = 512'h0055ffff035fffff0055ffff035fffff0055ffff035fffff0055ffff035fffff7f7f7f7f7f7f7f7f7f7f7f7fffffffff7fffffff7fffffff7fffffff7fffffff;

	lut_sub lut_175 ({sk[8], x6891x, x6892x, n_n1129, n_n1123, x6919x, n_n1128, x6935x}, n_n1107);
	defparam lut_175.LUT_SIZE = 8;
	defparam lut_175.mask = 256'h333333333333ffffffffffffffffffff7fffffffffffffffffffffffffffffff;

	lut_sub lut_183 ({sk[9], i_6_, x313x, x9x, x43x, x371x, x1198x, x1199x, x1194x}, n_n1114);
	defparam lut_183.LUT_SIZE = 9;
	defparam lut_183.mask = 512'h0055ffff035fffff0055ffff035fffff0055ffff035fffff0055ffff035fffff7f7f7fff7f7f7fff7f7f7fffffffffff555555ff555555ff555555ffffffffff;

	lut_sub lut_189 ({sk[10], i_6_, i_13_, i_1_, x340x, x632x, x1191x, x7975x}, x6947x);
	defparam lut_189.LUT_SIZE = 8;
	defparam lut_189.mask = 256'h0fff0fff3fff3fff0fff0fff3fff3fffbbbbbfffbbbbbbff00000fff000000ff;

	lut_sub lut_194 ({sk[11], i_7_, i_3_, i_4_, i_2_, n_n816, x6965x, x625x, x1156x}, n_n1185);
	defparam lut_194.LUT_SIZE = 9;
	defparam lut_194.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff00007f7f00ff7fff00005f5f00005f5f00007f7f00007f7f00005f5f00005f5f;

	lut_sub lut_199 ({sk[12], i_7_, i_8_, x369x, x617x, x1139x, x1141x, x6969x, x6970x}, x6975x);
	defparam lut_199.LUT_SIZE = 9;
	defparam lut_199.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff7fffffffffffffff7fffffff7fffffff7fff7fff7fff7fff7fff7fff7fff7fff;

	lut_sub lut_206 ({sk[13], i_3_, i_2_, n_n592, x614x, x1107x, x1110x, x6978x, x6979x}, x6991x);
	defparam lut_206.LUT_SIZE = 9;
	defparam lut_206.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff7fffffff7fffffff7fff7fff7fff7fff7fffffff7fffffff7fff7fffffffffff;

	lut_sub lut_213 ({sk[14], i_3_, i_2_, n_n638, x367x, x1108x, x6986x, x7974x}, x6992x);
	defparam lut_213.LUT_SIZE = 8;
	defparam lut_213.mask = 256'h0fff0fff3fff3fff0fff0fff3fff3fff3f3f3f3f3fff3fffbfbfbfbfbfffffff;

	lut_sub lut_219 ({sk[15], i_7_, i_3_, i_2_, n_n764, n_n570, x630x, x629x, x628x}, n_n1187);
	defparam lut_219.LUT_SIZE = 9;
	defparam lut_219.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff33333333333333ff33333333333333335f5f5f5f0f0f0fff5f5f5f5f0f0f0f0f;

	lut_sub lut_224 ({sk[0], i_13_, i_12_, i_11_, x600x, x1167x, x7972x, x7988x}, x6999x);
	defparam lut_224.LUT_SIZE = 8;
	defparam lut_224.mask = 256'h0fff0fff3fff3fff0fff0fff3fff3fffdfdfdfdfdfdfdfffdfdfdfdfdfdfdfdf;

	lut_sub lut_229 ({sk[1], i_10_, i_7_, i_8_, n_n791, x659x, x7004x, x7005x, x7007x}, n_n908);
	defparam lut_229.LUT_SIZE = 9;
	defparam lut_229.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff7fffffff7f7f7f7f7fff7fff7f7f7f7f55555555555555555555555555555555;

	lut_sub lut_235 ({sk[2], i_9_, i_10_, i_8_, i_3_, i_12_, n_n914, n_n913, x696x}, n_n906);
	defparam lut_235.LUT_SIZE = 9;
	defparam lut_235.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff7f3f7f3fff3f7f3f7f3f7f3f7f3f7f3f7f3f7f3f7f3f7f3f7f3f7f3f7f3f7f3f;

	lut_sub lut_240 ({sk[3], i_12_, n_n911, n_n910, n_n918, x678x, x7039x, x7062x}, x7065x);
	defparam lut_240.LUT_SIZE = 8;
	defparam lut_240.mask = 256'h0fff0fff3fff3fff0fff0fff3fff3fff7fffffffffffffff77ffffffffffffff;

	lut_sub lut_247 ({sk[4], i_8_, i_11_, x274x, x378x, x971x, x7986x}, x7075x);
	defparam lut_247.LUT_SIZE = 7;
	defparam lut_247.mask = 128'h0f0f5f5f0f0fffff7fff7f7f7f7f7f7f;

	lut_sub lut_252 ({sk[5], n_n959, n_n961, x7321x, x7335x, x7964x}, x7341x);
	defparam lut_252.LUT_SIZE = 6;
	defparam lut_252.mask = 64'h5fffffffbfffffff;

	lut_sub lut_258 ({sk[6], i_3_, n_n988, n_n991, x687x, x7192x, x7233x, x7197x, x7231x}, x7245x);
	defparam lut_258.LUT_SIZE = 9;
	defparam lut_258.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff7fff7fffffffffffffffffffffffffff7fffffffffffffffffffffffffffffff;

	lut_sub lut_266 ({sk[7], i_9_, i_5_, i_6_, i_12_, i_11_, i_0_, x21x, x712x}, x711x);
	defparam lut_266.LUT_SIZE = 9;
	defparam lut_266.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff0000550000005500000055000000550000005500000055000000550000005703;

	lut_sub lut_269 ({sk[8], i_7_, i_4_, i_12_, i_11_, n_n826, x708x, x10x, x710x}, x7179x);
	defparam lut_269.LUT_SIZE = 9;
	defparam lut_269.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff00550f5f0055005500000f0f0000000000770077007700770000000000000000;

	lut_sub lut_273 ({sk[9], x357x, x731x, x730x, x729x, x7199x, x7200x, x247x, x248x}, n_n986);
	defparam lut_273.LUT_SIZE = 9;
	defparam lut_273.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff7777777777ff77ff7f7f7f7f7fff7fff7777ffff77ffffff7f7fffff7fffffff;

	lut_sub lut_279 ({sk[10], i_4_, i_1_, n_n213, x744x, x742x, x7235x, x7236x, x200x}, x7242x);
	defparam lut_279.LUT_SIZE = 9;
	defparam lut_279.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff575757575757ffff57ff57ff57ffffff57575757575757575757575757575757;

	lut_sub lut_284 ({sk[11], n_n972, n_n977, n_n984, x7161x, x7162x, x7167x, x7168x}, x7337x);
	defparam lut_284.LUT_SIZE = 8;
	defparam lut_284.mask = 256'h0fff0fff3fff3fff0fff0fff3fff3fff7fffffffffffffffffffffffffffffff;

	lut_sub lut_292 ({sk[12], i_13_, i_12_, i_11_, x460x, x6587x, n_n1244, x466x, x6604x}, n_n1226);
	defparam lut_292.LUT_SIZE = 9;
	defparam lut_292.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff5fff5fff5fff5fff5fff5fff5fff5fff7fffffff5fffffff7fff7fff5fff5fff;

	lut_sub lut_298 ({sk[13], i_9_, i_10_, x6815x, x585x, x598x}, n_n1223);
	defparam lut_298.LUT_SIZE = 6;
	defparam lut_298.mask = 64'h5fffffff0f0f0f7f;

	lut_sub lut_302 ({sk[14], i_9_, i_11_, x1766x, x1723x, x421x, x457x, x6552x, x6576x}, x6823x);
	defparam lut_302.LUT_SIZE = 9;
	defparam lut_302.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff7777ffffffffffff7777ffffffffffff77ffffffffffffff7fffffffffffffff;

	lut_sub lut_309 ({sk[15], x1676x, x6617x, x1662x, x6627x, x6715x, x6716x}, x6824x);
	defparam lut_309.LUT_SIZE = 7;
	defparam lut_309.mask = 128'h0f0f5f5f0f0fffff7fffffffffffffff;

	lut_sub lut_316 ({sk[0], i_10_, i_11_, n_n1245, x6567x, x583x, x581x, x6805x}, x6825x);
	defparam lut_316.LUT_SIZE = 8;
	defparam lut_316.mask = 256'h0fff0fff3fff3fff0fff0fff3fff3fff55ffffff55ffffff5fffffff7fffffff;

	lut_sub lut_322 ({sk[1], i_6_, i_4_, i_11_, n_n761, x441x, x438x, x437x, x1376x}, n_n1121);
	defparam lut_322.LUT_SIZE = 9;
	defparam lut_322.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff5555555555555f5f5555555555557f7f555555ff55555f5f555555ff55557f7f;

	lut_sub lut_327 ({sk[2], i_6_, n_n675, n_n849, x1369x, x442x, x295x, x1362x, x6836x}, x6841x);
	defparam lut_327.LUT_SIZE = 9;
	defparam lut_327.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff3333333333ff33ff7777777777ff77ff3333ffff33ffffff7f7fffff7fffffff;

	lut_sub lut_333 ({sk[3], i_6_, x295x, x1324x, x6865x, x475x, x1314x, x1315x, x1316x}, x6869x);
	defparam lut_333.LUT_SIZE = 9;
	defparam lut_333.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff7f7fffffffffffff7fffffffffffffff7f7f7f7f7f7f7f7f7fff7fff7fff7fff;

	lut_sub lut_340 ({sk[4], i_3_, i_13_, i_4_, i_12_, i_1_, i_11_, n_n764, x1371x}, x444x);
	defparam lut_340.LUT_SIZE = 9;
	defparam lut_340.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff5755555557555755555555555555555555555555575557555555555555555555;

	lut_sub lut_344 ({sk[5], n_n849, x370x, n_n810, x470x, x1340x, x1341x, x1342x, x1344x}, n_n1116);
	defparam lut_344.LUT_SIZE = 9;
	defparam lut_344.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff7fff7fff7fff7fff7fffffff7fffffff7fff7fffffffffff7fffffffffffffff;

	lut_sub lut_351 ({sk[6], i_6_, n_n273, x45x, x371x, x1332x, x1333x, x471x, x1328x}, n_n1118);
	defparam lut_351.LUT_SIZE = 9;
	defparam lut_351.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff555555555555ffff777777777777ffff5fff5fff5fffffff7fff7fff7fffffff;

	lut_sub lut_357 ({sk[7], i_10_, n_n761, x7107x, x7108x, x670x, x7113x, x674x, x7116x}, n_n959);
	defparam lut_357.LUT_SIZE = 9;
	defparam lut_357.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff7f7fffffffffffff7fffffffffffffff5f5fffffffffffff5fffffffffffffff;

	lut_sub lut_364 ({sk[8], i_9_, i_13_, i_11_, n_n979, x858x, x7141x, x721x, x7149x}, n_n961);
	defparam lut_364.LUT_SIZE = 9;
	defparam lut_364.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffff5fffffff7fffffff5fffffff5fffffff5fffffff5fffffff5fffffff5fffffff;

	lut_sub lut_370 ({sk[9], n_n1001, n_n1000, x7262x, n_n998, x7311x, x7308x}, x7321x);
	defparam lut_370.LUT_SIZE = 7;
	defparam lut_370.mask = 128'h0f0f5f5f0f0fffff7fffffffffffffff;

	lut_sub lut_377 ({sk[10], i_5_, i_0_, n_n971, n_n970, x7331x, x758x}, x7335x);
	defparam lut_377.LUT_SIZE = 7;
	defparam lut_377.mask = 128'h0f0f5f5f0f0fffff3fff7fff3fff3fff;

	lut_sub lut_382 ({sk[11], i_13_, i_12_, n_n978, x7125x, n_n994, n_n996, x714x, x7318x}, x7964x);
	defparam lut_382.LUT_SIZE = 9;
	defparam lut_382.mask = 512'h5f5f5f5fffffffffffffffffffffffff5f5f5f5fffffffffffffffffffffffffa0000000000000008000000000000000a000000000000000a000000000000000;

	lut_sub lut_386 ({sk[12], i_3_, i_4_}, x21x);
	defparam lut_386.LUT_SIZE = 3;
	defparam lut_386.mask = 8'h52;

	lut_sub lut_388 ({sk[13], i_5_, i_6_, i_3_, i_2_}, x384x);
	defparam lut_388.LUT_SIZE = 5;
	defparam lut_388.mask = 32'h0f5f1000;

	lut_sub lut_390 ({sk[14], i_5_, i_6_, i_2_}, x385x);
	defparam lut_390.LUT_SIZE = 4;
	defparam lut_390.mask = 16'h7740;

	lut_sub lut_392 ({sk[15], i_9_, i_7_, i_6_, i_12_, i_2_, i_0_}, x1822x);
	defparam lut_392.LUT_SIZE = 7;
	defparam lut_392.mask = 128'h0f0f5f5f0f0fffff0000000000000001;

	lut_sub lut_394 ({sk[0], i_10_, i_5_, i_6_, i_1_, i_11_}, x1826x);
	defparam lut_394.LUT_SIZE = 6;
	defparam lut_394.mask = 64'h00ff1fff00001000;

	lut_sub lut_396 ({sk[1], i_10_, i_7_, i_8_, i_6_, i_3_, i_12_, i_2_, i_0_}, x7983x);
	defparam lut_396.LUT_SIZE = 9;
	defparam lut_396.mask = 512'h5555555555ff55ff55555555fffffffffffffffffffffffffffffffffffffffffffffffefffffefefffffffafffffafafffffefefffffefefffffffafffffafa;

	lut_sub lut_403 ({sk[2], i_9_, i_10_, i_7_, i_8_, i_12_, i_11_}, x665x);
	defparam lut_403.LUT_SIZE = 7;
	defparam lut_403.mask = 128'h555555ffffffffff5353ff5353ffffff;

	lut_sub lut_408 ({sk[3], i_7_, i_8_, i_3_, i_12_, i_1_, i_11_, i_0_}, x7982x);
	defparam lut_408.LUT_SIZE = 8;
	defparam lut_408.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5ffffffefefefefffffefefffffffffffefffe;

	lut_sub lut_416 ({sk[4], i_7_, i_6_, i_3_, i_12_, i_2_, i_0_}, x663x);
	defparam lut_416.LUT_SIZE = 7;
	defparam lut_416.mask = 128'h555555ffffffffff0f5f0f0f0f1f0f0f;

	lut_sub lut_420 ({sk[5], i_7_, i_8_, i_6_, i_3_, i_12_, i_1_, i_11_, i_0_}, x6513x);
	defparam lut_420.LUT_SIZE = 9;
	defparam lut_420.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff1111111100000000000000000000000000000005000000050005000500050005;

	lut_sub lut_424 ({sk[6], i_9_, i_10_, i_7_, i_8_, i_6_, i_11_, i_2_, i_0_}, x1805x);
	defparam lut_424.LUT_SIZE = 9;
	defparam lut_424.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0100000001000000010001000100000001000000010001000100010001000100;

	lut_sub lut_428 ({sk[7], i_7_, i_8_, i_5_, i_6_, i_3_, i_11_}, x1814x);
	defparam lut_428.LUT_SIZE = 7;
	defparam lut_428.mask = 128'h555555ffffffffff5000100000000000;

	lut_sub lut_431 ({sk[8], i_9_, i_10_, i_6_, i_1_, i_0_}, x6505x);
	defparam lut_431.LUT_SIZE = 6;
	defparam lut_431.mask = 64'h00ff1fff00000155;

	lut_sub lut_434 ({sk[9], i_9_, i_10_, i_7_, i_5_, i_6_, i_11_, i_2_, i_0_}, x7981x);
	defparam lut_434.LUT_SIZE = 9;
	defparam lut_434.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffffffffffffffffffffa8aaffffaaaaffffffffaaaafcffaaaaa8aaaaaaa8aaaaaa;

	lut_sub lut_446 ({sk[10], i_9_, i_7_, i_8_, i_6_, i_3_, i_1_, i_2_}, x683x);
	defparam lut_446.LUT_SIZE = 8;
	defparam lut_446.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff01010101010101010101010101773377;

	lut_sub lut_451 ({sk[11], i_10_, i_7_, i_5_, i_6_, i_3_, i_12_, i_1_}, x6526x);
	defparam lut_451.LUT_SIZE = 8;
	defparam lut_451.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000000000001010000110000001101;

	lut_sub lut_454 ({sk[12], i_9_, i_7_, i_5_, i_12_, i_1_, i_11_, i_2_}, x6527x);
	defparam lut_454.LUT_SIZE = 8;
	defparam lut_454.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000000000000000000000000000007;

	lut_sub lut_457 ({sk[13], i_9_, i_8_}, x18x);
	defparam lut_457.LUT_SIZE = 3;
	defparam lut_457.mask = 8'h51;

	lut_sub lut_459 ({sk[14], i_3_, i_2_, i_0_}, n_n818);
	defparam lut_459.LUT_SIZE = 4;
	defparam lut_459.mask = 16'h5501;

	lut_sub lut_461 ({sk[15], i_1_, i_2_, i_0_}, n_n833);
	defparam lut_461.LUT_SIZE = 4;
	defparam lut_461.mask = 16'h5504;

	lut_sub lut_463 ({sk[0], i_9_, i_10_, i_7_, i_8_, i_6_, i_13_, i_12_, i_11_}, x423x);
	defparam lut_463.LUT_SIZE = 9;
	defparam lut_463.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000000a000000080000000000000000000;

	lut_sub lut_466 ({sk[1], i_10_, i_7_, i_8_, i_6_, i_13_, i_12_}, x6548x);
	defparam lut_466.LUT_SIZE = 7;
	defparam lut_466.mask = 128'h555555ffffffffff0000008000000000;

	lut_sub lut_468 ({sk[2], i_9_, i_10_, i_7_, i_8_, i_6_, i_13_, i_12_, i_11_}, x7985x);
	defparam lut_468.LUT_SIZE = 9;
	defparam lut_468.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffffffffffffffffffffff5fffffff7fffffffffffffffffffffffffffffffffffff;

	lut_sub lut_488 ({sk[3], i_9_, i_5_, i_3_, i_4_, n_n833, x423x, x6548x, x7985x}, x1766x);
	defparam lut_488.LUT_SIZE = 9;
	defparam lut_488.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff00000000000f00000000000000aa000000000000003f00000000000000aa0000;

	lut_sub lut_492 ({sk[4], i_13_, i_12_}, n_n665);
	defparam lut_492.LUT_SIZE = 3;
	defparam lut_492.mask = 8'h52;

	lut_sub lut_494 ({sk[5], i_9_, i_10_, i_8_, i_13_, i_11_}, x337x);
	defparam lut_494.LUT_SIZE = 6;
	defparam lut_494.mask = 64'h00ff1fff00000020;

	lut_sub lut_496 ({sk[6], i_9_, i_10_, i_8_, i_5_, i_6_, i_2_, i_0_}, x1746x);
	defparam lut_496.LUT_SIZE = 8;
	defparam lut_496.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000000000000000000000000000103;

	lut_sub lut_499 ({sk[7], i_7_, i_5_, i_6_, i_1_, i_2_, i_0_}, x433x);
	defparam lut_499.LUT_SIZE = 7;
	defparam lut_499.mask = 128'h555555ffffffffffeec0aa80ccc08880;

	lut_sub lut_505 ({sk[8], i_7_, i_5_, i_1_, i_0_}, x6558x);
	defparam lut_505.LUT_SIZE = 5;
	defparam lut_505.mask = 32'h57573100;

	lut_sub lut_508 ({sk[9], i_10_, i_8_, i_11_, n_n665, x337x, x1746x, x433x, x6558x}, n_n1245);
	defparam lut_508.LUT_SIZE = 9;
	defparam lut_508.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff00550f5f00550f5f00550f5f00550f5f00553f7f00550f5f00550f5f00550f5f;

	lut_sub lut_512 ({sk[10], i_9_, i_10_, i_7_, i_8_, i_6_, i_1_, i_11_, i_0_}, x1757x);
	defparam lut_512.LUT_SIZE = 9;
	defparam lut_512.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000808800000000000085dd;

	lut_sub lut_517 ({sk[11], i_9_, i_7_, i_8_, i_13_, i_11_}, x353x);
	defparam lut_517.LUT_SIZE = 6;
	defparam lut_517.mask = 64'h00ff1fff00000200;

	lut_sub lut_519 ({sk[12], i_9_, i_8_, i_5_, i_6_, i_1_, i_11_, i_2_, i_0_}, x1738x);
	defparam lut_519.LUT_SIZE = 9;
	defparam lut_519.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff00000000000000000000000000000000000000000000000080008080c000c0c0;

	lut_sub lut_524 ({sk[13], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x434x);
	defparam lut_524.LUT_SIZE = 7;
	defparam lut_524.mask = 128'h555555ffffffffff0000000800000004;

	lut_sub lut_527 ({sk[14], i_9_, i_7_, i_8_, i_5_, i_6_, i_1_, i_11_}, x6555x);
	defparam lut_527.LUT_SIZE = 8;
	defparam lut_527.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff0000000000000000000000000000008f;

	lut_sub lut_530 ({sk[15], i_9_, i_10_, i_7_, i_8_, i_5_, i_1_, i_2_, i_0_}, x7978x);
	defparam lut_530.LUT_SIZE = 9;
	defparam lut_530.mask = 512'h5555555555ff55ff55555555fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffefcfffffef0;

	lut_sub lut_538 ({sk[0], i_13_, i_12_, x1757x, x353x, x1738x, x434x, x6555x, x7978x}, x6567x);
	defparam lut_538.LUT_SIZE = 9;
	defparam lut_538.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff00000f0f00000f0f00000f0f00000f0fbbffbfffffffffff00000f0f00000f0f;

	lut_sub lut_544 ({sk[1], i_5_, i_3_, i_4_}, n_n541);
	defparam lut_544.LUT_SIZE = 4;
	defparam lut_544.mask = 16'h5520;

	lut_sub lut_546 ({sk[2], i_9_, i_7_, i_8_}, n_n638);
	defparam lut_546.LUT_SIZE = 4;
	defparam lut_546.mask = 16'h5501;

	lut_sub lut_548 ({sk[3], i_3_, i_4_, i_1_, i_2_}, x298x);
	defparam lut_548.LUT_SIZE = 5;
	defparam lut_548.mask = 32'h57570040;

	lut_sub lut_550 ({sk[4], i_3_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_}, x306x);
	defparam lut_550.LUT_SIZE = 8;
	defparam lut_550.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000000000000000020000000000000;

	lut_sub lut_552 ({sk[5], i_10_, i_6_, i_13_, i_12_, i_1_, i_11_, i_2_, i_0_}, x459x);
	defparam lut_552.LUT_SIZE = 9;
	defparam lut_552.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff1c0c000000000000100000000000000000000000000000000000000000000000;

	lut_sub lut_555 ({sk[6], i_10_, i_5_, i_6_, i_13_, i_12_, i_11_}, x6572x);
	defparam lut_555.LUT_SIZE = 7;
	defparam lut_555.mask = 128'h555555ffffffffff0040000000000000;

	lut_sub lut_557 ({sk[7], i_5_, i_6_, i_3_, i_4_, i_12_, i_1_, i_2_}, x1728x);
	defparam lut_557.LUT_SIZE = 8;
	defparam lut_557.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000000000000000000000000001000;

	lut_sub lut_559 ({sk[8], i_6_, n_n541, n_n638, x298x, x306x, x459x, x6572x, x1728x}, x1723x);
	defparam lut_559.LUT_SIZE = 9;
	defparam lut_559.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0000000055557777000000005f5f7f7f0000000055ff77ff000000005fff7fff;

	lut_sub lut_564 ({sk[9], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_, n_n592, n_n597}, x460x);
	defparam lut_564.LUT_SIZE = 9;
	defparam lut_564.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0000000000000500000000000503000000000000000000300000000050300000;

	lut_sub lut_571 ({sk[10], i_9_, i_5_, i_13_, n_n844, n_n832, n_n1574, x6581x, x6583x}, x6587x);
	defparam lut_571.LUT_SIZE = 9;
	defparam lut_571.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0f0f0f0f0f0f5f5f0f0f0f0f0f0f5f5f0f0f0f0f0f0f5f5f0f3f0f3f0f3f5f7f;

	lut_sub lut_575 ({sk[11], n_n665, x337x, x465x, x464x, x1702x, n_n597, x6588x, x6590x}, n_n1244);
	defparam lut_575.LUT_SIZE = 9;
	defparam lut_575.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff000033330000333300003333ffffffff05ff37ff05ff37ff05ff37ffffffffff;

	lut_sub lut_580 ({sk[12], i_9_, i_7_, i_8_, x469x, x467x, x6598x, x6599x, x1691x}, x466x);
	defparam lut_580.LUT_SIZE = 9;
	defparam lut_580.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff5757575757575757575757575757575757ff57ff575757575757ffff57575757;

	lut_sub lut_585 ({sk[13], i_9_, i_10_, i_13_, i_12_, i_11_, n_n844, x391x, x6596x}, x6604x);
	defparam lut_585.LUT_SIZE = 9;
	defparam lut_585.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0357000000000000000000000000000003030000000000000000000000000000;

	lut_sub lut_588 ({sk[14], i_7_, i_8_, i_6_}, n_n748);
	defparam lut_588.LUT_SIZE = 4;
	defparam lut_588.mask = 16'h5510;

	lut_sub lut_590 ({sk[15], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x409x);
	defparam lut_590.LUT_SIZE = 7;
	defparam lut_590.mask = 128'h555555ffffffffff0000000000000002;

	lut_sub lut_592 ({sk[0], i_9_, i_13_, i_12_, i_11_}, x284x);
	defparam lut_592.LUT_SIZE = 5;
	defparam lut_592.mask = 32'h57574000;

	lut_sub lut_594 ({sk[1], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x484x);
	defparam lut_594.LUT_SIZE = 7;
	defparam lut_594.mask = 128'h555555ffffffffff0800000004000000;

	lut_sub lut_597 ({sk[2], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x6613x);
	defparam lut_597.LUT_SIZE = 7;
	defparam lut_597.mask = 128'h555555ffffffffff0000400000000000;

	lut_sub lut_599 ({sk[3], i_5_, i_3_, i_4_, n_n748, x409x, x284x, x484x, x6613x}, x1676x);
	defparam lut_599.LUT_SIZE = 9;
	defparam lut_599.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff000f030f00000303000003030000030305050707000003030000030300000303;

	lut_sub lut_603 ({sk[4], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x391x);
	defparam lut_603.LUT_SIZE = 7;
	defparam lut_603.mask = 128'h555555ffffffffff0000800000000000;

	lut_sub lut_605 ({sk[5], i_10_, i_7_, i_8_, i_6_, i_13_, i_12_, i_11_}, x482x);
	defparam lut_605.LUT_SIZE = 8;
	defparam lut_605.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff000000000000a0c00000000000000000;

	lut_sub lut_608 ({sk[6], i_13_, i_12_, i_1_, i_11_, i_2_, i_0_}, x6607x);
	defparam lut_608.LUT_SIZE = 7;
	defparam lut_608.mask = 128'h555555ffffffffff0000200000000000;

	lut_sub lut_610 ({sk[7], i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x6608x);
	defparam lut_610.LUT_SIZE = 8;
	defparam lut_610.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000000000000000000000000000020;

	lut_sub lut_612 ({sk[8], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x6609x);
	defparam lut_612.LUT_SIZE = 7;
	defparam lut_612.mask = 128'h555555ffffffffff0000000000000001;

	lut_sub lut_614 ({sk[9], i_9_, i_5_, i_3_, i_13_, i_4_, i_12_}, x6610x);
	defparam lut_614.LUT_SIZE = 7;
	defparam lut_614.mask = 128'h555555ffffffffff0000800000000000;

	lut_sub lut_616 ({sk[10], i_9_, i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x6611x);
	defparam lut_616.LUT_SIZE = 8;
	defparam lut_616.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000000000000000000100000000000;

	lut_sub lut_618 ({sk[11], i_13_, i_12_, i_1_, i_11_, i_2_, i_0_}, x6612x);
	defparam lut_618.LUT_SIZE = 7;
	defparam lut_618.mask = 128'h555555ffffffffff0800000000000000;

	lut_sub lut_620 ({sk[12], x391x, x482x, x6607x, x6608x, x6609x, x6610x, x6611x, x6612x}, x6617x);
	defparam lut_620.LUT_SIZE = 9;
	defparam lut_620.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff000f000f000fffff333f333f333fffff555f555f555fffff777f777f777fffff;

	lut_sub lut_625 ({sk[13], i_7_, i_8_, i_6_}, n_n746);
	defparam lut_625.LUT_SIZE = 4;
	defparam lut_625.mask = 16'h5520;

	lut_sub lut_627 ({sk[14], i_9_, i_10_, i_13_, i_12_, i_11_}, x282x);
	defparam lut_627.LUT_SIZE = 6;
	defparam lut_627.mask = 64'h00ff1fff40000000;

	lut_sub lut_629 ({sk[15], i_8_, i_5_, i_6_, i_3_, i_4_, i_2_}, x1669x);
	defparam lut_629.LUT_SIZE = 7;
	defparam lut_629.mask = 128'h555555ffffffffff0000000040000000;

	lut_sub lut_631 ({sk[0], i_7_, i_8_, i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x7979x);
	defparam lut_631.LUT_SIZE = 9;
	defparam lut_631.mask = 512'h5555555555ff55ff55555555fffffffffffffffffffffffffffffffffffffffffffffffffffffffff0fffffffafffffffffffffffffffffffcffffffffffffff;

	lut_sub lut_639 ({sk[1], i_3_, i_4_, i_0_, n_n746, x282x, x1669x, x7979x}, x1662x);
	defparam lut_639.LUT_SIZE = 8;
	defparam lut_639.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff0b0b0b0f0b0b0b0b0b0b0b0b0b0b0b0b;

	lut_sub lut_643 ({sk[2], i_1_, i_2_, i_0_}, n_n844);
	defparam lut_643.LUT_SIZE = 4;
	defparam lut_643.mask = 16'h5501;

	lut_sub lut_645 ({sk[3], i_7_, i_8_, i_6_}, n_n756);
	defparam lut_645.LUT_SIZE = 4;
	defparam lut_645.mask = 16'h5502;

	lut_sub lut_647 ({sk[4], i_10_, i_13_, i_12_, i_11_}, x294x);
	defparam lut_647.LUT_SIZE = 5;
	defparam lut_647.mask = 32'h57574000;

	lut_sub lut_649 ({sk[5], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x501x);
	defparam lut_649.LUT_SIZE = 7;
	defparam lut_649.mask = 128'h555555ffffffffff2000000010000000;

	lut_sub lut_652 ({sk[6], i_9_, i_10_, i_8_, i_3_, i_13_, i_12_}, x6619x);
	defparam lut_652.LUT_SIZE = 7;
	defparam lut_652.mask = 128'h555555ffffffffff0080000000000000;

	lut_sub lut_654 ({sk[7], i_4_, n_n844, x391x, n_n756, x284x, x294x, x501x, x6619x}, x6627x);
	defparam lut_654.LUT_SIZE = 9;
	defparam lut_654.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff000000330f0f0f3f555555775f5f5f7f000000330f0f0f3f000000330f0f0f3f;

	lut_sub lut_658 ({sk[8], i_3_, i_13_, i_12_, i_11_, n_n835, x1637x, x499x, x1634x}, n_n1250);
	defparam lut_658.LUT_SIZE = 9;
	defparam lut_658.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff5f5f55555f5f55557fff55555f5f55555f5f55555f5f55557f7f55555f5f5555;

	lut_sub lut_663 ({sk[9], i_5_, i_3_, i_4_, n_n725, n_n837, x520x, x1629x, x6648x}, x1623x);
	defparam lut_663.LUT_SIZE = 9;
	defparam lut_663.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000033773f7f000000000000000000000000;

	lut_sub lut_667 ({sk[10], i_9_, i_0_, x303x, n_n837, x6650x, x518x, x517x, x6643x}, x6652x);
	defparam lut_667.LUT_SIZE = 9;
	defparam lut_667.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff111111ff111111ff111111ff1f1f1fff1111111111111111111111111f1f1f1f;

	lut_sub lut_671 ({sk[11], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_, x6650x, x6654x}, x6658x);
	defparam lut_671.LUT_SIZE = 9;
	defparam lut_671.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0500000000000000000000000000000000050000300000050000000000000000;

	lut_sub lut_676 ({sk[12], n_n725, n_n832, n_n837, n_n710, x541x, x6655x, x6656x, x6657x}, x6659x);
	defparam lut_676.LUT_SIZE = 9;
	defparam lut_676.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff00000000000033330000555500007777000000000f0f3f3f00ff55ff0fff7fff;

	lut_sub lut_681 ({sk[13], i_13_, i_12_, i_11_, n_n844, n_n710, x546x, x6662x, x1605x}, x1595x);
	defparam lut_681.LUT_SIZE = 9;
	defparam lut_681.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff00005f7f00005577000055770000557700005577000055770000557700005577;

	lut_sub lut_685 ({sk[14], i_7_, i_8_, i_6_, n_n849, n_n755, x405x, x544x, x543x}, x6666x);
	defparam lut_685.LUT_SIZE = 9;
	defparam lut_685.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0f0f0f0f00330033000000000000555500000000000000000000000000000000;

	lut_sub lut_689 ({sk[15], i_7_, i_13_, i_11_, x18x, x455x, x454x, x453x, x6631x}, n_n1248);
	defparam lut_689.LUT_SIZE = 9;
	defparam lut_689.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0055005500550055005533770055005500550f5f00550f5f00550f5f00550f5f;

	lut_sub lut_693 ({sk[0], i_9_, i_10_, i_5_, i_6_, i_11_, n_n761, n_n672, x6674x}, x1584x);
	defparam lut_693.LUT_SIZE = 9;
	defparam lut_693.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0007000500050007000500050005000700070005000500050005000500050005;

	lut_sub lut_697 ({sk[1], i_3_, x17x, x266x, n_n835, x399x, x480x, x6670x, x6672x}, x6678x);
	defparam lut_697.LUT_SIZE = 9;
	defparam lut_697.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff030303035757575703ffffff57ffffff030303035757575703ff03ff57ff57ff;

	lut_sub lut_702 ({sk[2], i_10_, i_5_, i_3_, i_13_, i_4_, i_12_, x573x, x572x}, x1570x);
	defparam lut_702.LUT_SIZE = 9;
	defparam lut_702.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0005000000000000000300000000000000000000000000000000000000000000;

	lut_sub lut_705 ({sk[3], x313x, x17x, x266x, n_n752, x6679x, x121x, x404x, x570x}, x6683x);
	defparam lut_705.LUT_SIZE = 9;
	defparam lut_705.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff00000f0f55555f5f00ff0fff55ff5fff33333f3f77777f7f33ff3fff77ff7fff;

	lut_sub lut_710 ({sk[4], i_3_, i_13_, i_12_, n_n651, x550x, x1552x, x6697x, x1554x}, x1547x);
	defparam lut_710.LUT_SIZE = 9;
	defparam lut_710.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff00000000000000005fff7fff0000000000000000000000005f5f7f7f00000000;

	lut_sub lut_715 ({sk[5], i_10_, i_13_, i_12_, i_11_, x28x, n_n710, x6689x, x108x}, x1564x);
	defparam lut_715.LUT_SIZE = 9;
	defparam lut_715.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff000000000000777f000000000000000000000000000077770000000000000000;

	lut_sub lut_719 ({sk[6], x274x, x313x, x17x, x266x, n_n678, x6684x, x6685x, x6686x}, x6693x);
	defparam lut_719.LUT_SIZE = 9;
	defparam lut_719.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff000f555f000f555f333f777f333f777f000f555fffffffff333f777fffffffff;

	lut_sub lut_724 ({sk[7], i_1_, i_0_}, x377x);
	defparam lut_724.LUT_SIZE = 3;
	defparam lut_724.mask = 8'h58;

	lut_sub lut_726 ({sk[8], i_7_, i_8_, i_6_}, n_n843);
	defparam lut_726.LUT_SIZE = 4;
	defparam lut_726.mask = 16'h5580;

	lut_sub lut_728 ({sk[9], i_5_, i_3_, i_13_, i_4_, i_12_}, x302x);
	defparam lut_728.LUT_SIZE = 6;
	defparam lut_728.mask = 64'h00ff1fff00800000;

	lut_sub lut_730 ({sk[10], i_9_, i_7_, i_8_, i_5_, i_6_}, x6706x);
	defparam lut_730.LUT_SIZE = 6;
	defparam lut_730.mask = 64'h00ff1fff20000000;

	lut_sub lut_732 ({sk[11], i_10_, i_3_, i_13_, i_4_, i_12_, i_1_, i_11_, i_2_}, x6707x);
	defparam lut_732.LUT_SIZE = 9;
	defparam lut_732.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000040000000000000;

	lut_sub lut_734 ({sk[12], i_10_, i_7_, i_8_, i_6_, i_11_}, x6710x);
	defparam lut_734.LUT_SIZE = 6;
	defparam lut_734.mask = 64'h00ff1fff00001000;

	lut_sub lut_736 ({sk[13], i_10_, i_5_, i_3_, i_13_, i_4_, i_12_, i_11_}, x6711x);
	defparam lut_736.LUT_SIZE = 8;
	defparam lut_736.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000000000000000000000000002000;

	lut_sub lut_738 ({sk[14], i_2_, x377x, n_n843, x302x, x6706x, x6707x, x6710x, x6711x}, x6715x);
	defparam lut_738.LUT_SIZE = 9;
	defparam lut_738.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff000f000f000f000f000f000f000f000f000f000f000f000f000f333f555f777f;

	lut_sub lut_742 ({sk[15], i_5_, i_3_, i_4_}, n_n538);
	defparam lut_742.LUT_SIZE = 4;
	defparam lut_742.mask = 16'h5502;

	lut_sub lut_744 ({sk[0], i_9_, i_10_, i_7_, i_8_, i_6_, i_13_, i_12_, i_11_}, x568x);
	defparam lut_744.LUT_SIZE = 9;
	defparam lut_744.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0000000000000000a0c000000000000000000000000000000000000000000000;

	lut_sub lut_748 ({sk[1], i_9_, i_10_, i_7_, i_5_, i_6_, i_3_, i_1_, i_0_}, x567x);
	defparam lut_748.LUT_SIZE = 9;
	defparam lut_748.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff000000000000000000000000000000000000000000000000000000000005030f;

	lut_sub lut_752 ({sk[2], i_13_, i_12_, i_1_, i_2_, i_0_, n_n538, x568x, x567x}, x6716x);
	defparam lut_752.LUT_SIZE = 9;
	defparam lut_752.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0000000300000000000000030000000055555557555555550000000300000000;

	lut_sub lut_755 ({sk[3], i_10_, i_4_, n_n853, x6718x, x394x, x6719x, x6720x, x6724x}, x6730x);
	defparam lut_755.LUT_SIZE = 9;
	defparam lut_755.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0303030357ff57ff0303030357ffffff0303030303ff03ff0303030303ffffff;

	lut_sub lut_760 ({sk[4], n_n2368, x322x, x336x, x420x, x6721x, x6722x, x6723x, x6725x}, x6731x);
	defparam lut_760.LUT_SIZE = 9;
	defparam lut_760.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff000000ff0f0f0fff333333ff3f3f3fff555555ff5f5f5fff777777ff7f7f7fff;

	lut_sub lut_765 ({sk[5], i_9_, i_7_, i_8_, i_6_, i_4_, i_0_, n_n816, x451x}, x1511x);
	defparam lut_765.LUT_SIZE = 9;
	defparam lut_765.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0057005500000000000000000000000000000000000000000000000000000000;

	lut_sub lut_768 ({sk[6], i_6_, i_4_, i_1_, i_0_, n_n792, n_n853, x70x, x450x}, x6738x);
	defparam lut_768.LUT_SIZE = 9;
	defparam lut_768.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff3377337733773377337f3377337f33773377337733773377337f337733773377;

	lut_sub lut_773 ({sk[7], i_5_, i_6_, i_1_, i_2_, i_0_, n_n816, x9x, x266x}, x575x);
	defparam lut_773.LUT_SIZE = 9;
	defparam lut_773.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0000030300000303000000000000030300005557000055570000000000005557;

	lut_sub lut_780 ({sk[8], i_7_, i_13_, i_4_, i_1_, i_0_, n_n816, x574x, x6786x}, x6789x);
	defparam lut_780.LUT_SIZE = 9;
	defparam lut_780.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0303030303570303030303030303030300000000005500000000000000000000;

	lut_sub lut_783 ({sk[9], n_n835, x307x, x272x, x46x, x115x, x302x, x6808x, x6810x}, x6815x);
	defparam lut_783.LUT_SIZE = 9;
	defparam lut_783.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff00ff00ff00ffffff00ff00ff00ffffff05ff05ff05ffffff37ff37ff37ffffff;

	lut_sub lut_788 ({sk[10], i_13_, i_12_, i_11_, n_n847, x292x, x588x, x587x, x586x}, x585x);
	defparam lut_788.LUT_SIZE = 9;
	defparam lut_788.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff000055550000555500005555000055553fff7fff33ff77ff0fff5fff00ff55ff;

	lut_sub lut_793 ({sk[11], i_5_, i_6_, i_13_, i_12_, i_11_, n_n818, x272x, x384x}, x598x);
	defparam lut_793.LUT_SIZE = 9;
	defparam lut_793.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff000000005f005f00000000005f0f5500333300007f335f00333300007f3f5500;

	lut_sub lut_798 ({sk[12], i_13_, i_12_}, n_n761);
	defparam lut_798.LUT_SIZE = 3;
	defparam lut_798.mask = 8'h54;

	lut_sub lut_800 ({sk[13], i_10_, i_7_, i_8_, i_3_, i_1_, i_2_}, x441x);
	defparam lut_800.LUT_SIZE = 7;
	defparam lut_800.mask = 128'h555555ffffffffffc888000088880000;

	lut_sub lut_803 ({sk[14], i_9_, i_10_, i_7_, i_8_, i_3_, i_4_, i_1_, i_2_}, x438x);
	defparam lut_803.LUT_SIZE = 9;
	defparam lut_803.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0c000c080c000c08000008080c000c080c000c00000000000000000000000000;

	lut_sub lut_807 ({sk[15], i_9_, i_10_, i_7_, i_8_, i_3_, i_1_, i_2_}, x437x);
	defparam lut_807.LUT_SIZE = 8;
	defparam lut_807.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffffcc8080cc808080cccc80808080808080;

	lut_sub lut_811 ({sk[0], i_10_, i_8_, i_13_, i_4_, i_12_, i_1_, i_11_, i_2_}, x1376x);
	defparam lut_811.LUT_SIZE = 9;
	defparam lut_811.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0000002000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_813 ({sk[1], i_3_, i_1_, i_2_}, n_n675);
	defparam lut_813.LUT_SIZE = 4;
	defparam lut_813.mask = 16'h5580;

	lut_sub lut_815 ({sk[2], i_10_, i_13_, i_12_}, n_n849);
	defparam lut_815.LUT_SIZE = 4;
	defparam lut_815.mask = 16'h5540;

	lut_sub lut_817 ({sk[3], i_10_, i_7_, i_8_, i_13_, i_4_, i_12_, i_1_}, x1369x);
	defparam lut_817.LUT_SIZE = 8;
	defparam lut_817.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff02000000000000000000000000000000;

	lut_sub lut_819 ({sk[4], i_7_, i_8_, i_6_, i_3_, i_4_, i_1_, i_2_}, x442x);
	defparam lut_819.LUT_SIZE = 8;
	defparam lut_819.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000c0800000c000000080800000000;

	lut_sub lut_822 ({sk[5], i_13_, i_4_, i_12_}, x295x);
	defparam lut_822.LUT_SIZE = 4;
	defparam lut_822.mask = 16'h5510;

	lut_sub lut_824 ({sk[6], i_7_, i_6_, i_13_, i_12_, i_1_, i_11_, i_2_}, x1362x);
	defparam lut_824.LUT_SIZE = 8;
	defparam lut_824.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000000000000002000000000000000;

	lut_sub lut_826 ({sk[7], i_8_, i_6_, i_13_, i_12_, i_11_}, x6836x);
	defparam lut_826.LUT_SIZE = 6;
	defparam lut_826.mask = 64'h00ff1fff00200000;

	lut_sub lut_828 ({sk[8], i_13_, i_11_}, n_n787);
	defparam lut_828.LUT_SIZE = 3;
	defparam lut_828.mask = 8'h54;

	lut_sub lut_830 ({sk[9], i_9_, i_7_, i_8_, i_3_, i_4_, i_1_, i_2_}, x448x);
	defparam lut_830.LUT_SIZE = 8;
	defparam lut_830.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff080008080c000c080800080008000800;

	lut_sub lut_834 ({sk[10], i_9_, i_7_, i_8_, i_3_, i_13_, i_1_, i_11_}, x1355x);
	defparam lut_834.LUT_SIZE = 8;
	defparam lut_834.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000000200000000000000000000000;

	lut_sub lut_836 ({sk[11], i_9_, i_7_, i_13_, i_12_, i_1_, i_11_, i_2_}, x1356x);
	defparam lut_836.LUT_SIZE = 8;
	defparam lut_836.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff08080000080000000000000000000000;

	lut_sub lut_839 ({sk[12], i_9_, i_7_, i_6_, i_3_, i_13_, i_12_, i_1_, i_11_}, x1351x);
	defparam lut_839.LUT_SIZE = 9;
	defparam lut_839.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0000000000000000000000002000000000000000000000000000000000000000;

	lut_sub lut_841 ({sk[13], i_9_, i_8_, i_6_, i_3_, i_13_, i_12_, i_1_, i_2_}, x1352x);
	defparam lut_841.LUT_SIZE = 9;
	defparam lut_841.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0000000000000000000000002000000000000000000000000000000000000000;

	lut_sub lut_843 ({sk[14], i_9_, i_7_, i_6_, i_13_, i_12_, i_1_, i_2_}, x1354x);
	defparam lut_843.LUT_SIZE = 8;
	defparam lut_843.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000000000020000000000000000000;

	lut_sub lut_845 ({sk[15], i_9_, i_10_, i_8_, i_3_, i_13_, i_12_, i_11_}, x1324x);
	defparam lut_845.LUT_SIZE = 8;
	defparam lut_845.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00004000000000000000000000000000;

	lut_sub lut_847 ({sk[0], i_9_, i_10_, i_7_, i_13_, i_4_, i_12_, i_11_, i_2_}, x6865x);
	defparam lut_847.LUT_SIZE = 9;
	defparam lut_847.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0033000020330000000000000000000000000000202000000000000000000000;

	lut_sub lut_850 ({sk[1], i_9_, i_7_, i_8_, i_6_, i_3_, i_2_}, x475x);
	defparam lut_850.LUT_SIZE = 7;
	defparam lut_850.mask = 128'h555555ffffffffff000a0c0f00000000;

	lut_sub lut_854 ({sk[2], i_10_, i_7_, i_8_, i_6_, i_3_, i_13_, i_12_, i_11_}, x1314x);
	defparam lut_854.LUT_SIZE = 9;
	defparam lut_854.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0000000040000000000000000000000000000000000000000000000000000000;

	lut_sub lut_856 ({sk[3], i_9_, i_6_, i_3_, i_13_, i_4_, i_12_, i_2_}, x1315x);
	defparam lut_856.LUT_SIZE = 8;
	defparam lut_856.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff00000000020000000000000000000000;

	lut_sub lut_858 ({sk[4], i_10_, i_8_, i_6_, i_3_, i_13_, i_12_, i_11_, i_2_}, x1316x);
	defparam lut_858.LUT_SIZE = 9;
	defparam lut_858.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0000000000000000200000000000000000000000000000000000000000000000;

	lut_sub lut_860 ({sk[5], i_9_, i_10_, i_7_, i_3_, i_12_, i_1_, n_n1126, x6887x}, x6891x);
	defparam lut_860.LUT_SIZE = 9;
	defparam lut_860.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff333337373333373733333737333337373333373733333737333337373333373f;

	lut_sub lut_864 ({sk[6], i_3_, x1294x, x491x, x1293x, x1295x, x1296x, x6889x}, x6892x);
	defparam lut_864.LUT_SIZE = 8;
	defparam lut_864.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5fffff7fff7fffffffffff7fffffffffffffff;

	lut_sub lut_871 ({sk[7], i_4_, i_12_, i_1_, i_11_, x298x, x504x, x1268x, x6894x}, n_n1129);
	defparam lut_871.LUT_SIZE = 9;
	defparam lut_871.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff77ff77777fff7f7f777777777f7f7f7f77ff777777ff77777777777777777777;

	lut_sub lut_876 ({sk[8], i_6_, i_3_, i_1_, n_n311, n_n592, x508x, x1256x, x6904x}, n_n1123);
	defparam lut_876.LUT_SIZE = 9;
	defparam lut_876.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff7f7f7f7f7f7f7f7f7f7f7f7f7f7f7f7f7777777777777777777777ff77777777;

	lut_sub lut_881 ({sk[9], x1246x, x1247x, x6909x, x7976x, x7989x}, x6919x);
	defparam lut_881.LUT_SIZE = 6;
	defparam lut_881.mask = 64'h00ff1fffdfffffff;

	lut_sub lut_887 ({sk[10], i_9_, i_8_, i_6_, i_12_, n_n346, x554x, x1219x, x1220x}, n_n1128);
	defparam lut_887.LUT_SIZE = 9;
	defparam lut_887.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff7f7f7f7f777777777f7f7f7f777777777f7f7f7f777777777f7f7f7f777777ff;

	lut_sub lut_892 ({sk[11], i_6_, i_3_, i_4_, i_1_, i_11_, i_2_, x604x, x603x}, x6935x);
	defparam lut_892.LUT_SIZE = 9;
	defparam lut_892.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff00000000000000005f5577770000000000000000000000005555777700000000;

	lut_sub lut_896 ({sk[12], i_10_, i_13_, i_12_, i_11_}, x313x);
	defparam lut_896.LUT_SIZE = 5;
	defparam lut_896.mask = 32'h57571000;

	lut_sub lut_898 ({sk[13], i_9_, i_4_}, x9x);
	defparam lut_898.LUT_SIZE = 3;
	defparam lut_898.mask = 8'h54;

	lut_sub lut_900 ({sk[14], i_10_, i_7_, i_8_, i_6_, i_3_, i_2_}, x43x);
	defparam lut_900.LUT_SIZE = 7;
	defparam lut_900.mask = 128'h555555ffffffffffe0c0a00000000000;

	lut_sub lut_903 ({sk[15], i_13_, i_4_, i_1_}, x371x);
	defparam lut_903.LUT_SIZE = 4;
	defparam lut_903.mask = 16'h5510;

	lut_sub lut_905 ({sk[0], i_10_, i_7_, i_8_, i_3_, i_13_, i_4_, i_1_, i_11_}, x1198x);
	defparam lut_905.LUT_SIZE = 9;
	defparam lut_905.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff2300030000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_908 ({sk[1], i_10_, i_8_, i_3_, i_13_, i_4_, i_12_, i_1_, i_2_}, x1199x);
	defparam lut_908.LUT_SIZE = 9;
	defparam lut_908.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0022000000000000202200000000000000000000000000000000000000000000;

	lut_sub lut_911 ({sk[2], i_10_, i_8_, i_6_, i_3_, i_13_, i_1_, i_11_, i_2_}, x1194x);
	defparam lut_911.LUT_SIZE = 9;
	defparam lut_911.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff0800000000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_913 ({sk[3], i_9_, i_10_, i_13_, i_4_}, x340x);
	defparam lut_913.LUT_SIZE = 5;
	defparam lut_913.mask = 32'h57574000;

	lut_sub lut_915 ({sk[4], i_9_, i_10_, i_7_, i_8_, i_3_, i_12_, i_11_, i_2_}, x632x);
	defparam lut_915.LUT_SIZE = 9;
	defparam lut_915.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffffcc88f888cc00f000000000000000000000000000000000000000000000000000;

	lut_sub lut_919 ({sk[5], i_10_, i_7_, i_8_, i_3_, i_13_, i_12_, i_1_, i_11_}, x1191x);
	defparam lut_919.LUT_SIZE = 9;
	defparam lut_919.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff2000000030000000000000000000000000000000000000000000000000000000;

	lut_sub lut_922 ({sk[6], i_10_, i_7_, i_13_, i_12_, i_1_, i_11_, i_2_}, x7975x);
	defparam lut_922.LUT_SIZE = 8;
	defparam lut_922.mask = 256'h5f5f5fff5f5fffff5f5f5fff5f5ffffff7f7fffff5ffffffffffffffffffffff;

	lut_sub lut_930 ({sk[7], i_10_, i_13_, i_11_}, n_n816);
	defparam lut_930.LUT_SIZE = 4;
	defparam lut_930.mask = 16'h5540;

	lut_sub lut_932 ({sk[8], i_9_, i_10_, i_8_, i_3_, i_13_, i_4_, i_12_, i_11_}, x6965x);
	defparam lut_932.LUT_SIZE = 9;
	defparam lut_932.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffffaf000f008f000f00000000000000000000000000000000000000000000000000;

	lut_sub lut_936 ({sk[9], i_10_, i_7_, i_8_, i_13_, i_12_, i_11_}, x625x);
	defparam lut_936.LUT_SIZE = 7;
	defparam lut_936.mask = 128'h555555ffffffffffa0c0000000000000;

	lut_sub lut_940 ({sk[10], i_9_, i_10_, i_7_, i_8_, i_3_, i_13_, i_4_, i_12_}, x1156x);
	defparam lut_940.LUT_SIZE = 9;
	defparam lut_940.mask = 512'h5555555555ff55ff55555555ffffffffffffffffffffffffffffffffffffffff3030a0000000a000000000000000000030300000000000000000000000000000;

	lut_sub lut_943 ({sk[11], i_10_, i_13_, i_4_, i_11_}, x369x);
	defparam lut_943.LUT_SIZE = 5;
	defparam lut_943.mask = 32'h57571000;

	lut_sub lut_945 ({sk[12], i_9_, i_10_, i_8_, i_3_, i_13_, i_4_, i_12_, i_11_}, x617x);
	defparam lut_945.LUT_SIZE = 9;
	defparam lut_945.mask = 512'h5f5fffff5f5fffffffffffffffffffff5f5fffff5f5fffffffffffffffffffff0500050045000500000000000000000000000000440000000000000000000000;

	lut_sub lut_948 ({sk[13], i_9_, i_7_, i_8_, i_3_, i_13_, i_4_, i_11_, i_2_}, x1139x);
	defparam lut_948.LUT_SIZE = 9;
	defparam lut_948.mask = 512'h5f5fffff5f5fffffffffffffffffffff5f5fffff5f5fffffffffffffffffffff0000000000000000450000000500000000000000000000000000000000000000;

	lut_sub lut_951 ({sk[14], i_9_, i_7_, i_8_, i_3_, i_13_, i_4_, i_12_, i_11_}, x1141x);
	defparam lut_951.LUT_SIZE = 9;
	defparam lut_951.mask = 512'h5f5fffff5f5fffffffffffffffffffff5f5fffff5f5fffffffffffffffffffff0000000000000000230000000300000000000000000000000000000000000000;

	lut_sub lut_954 ({sk[15], i_9_, i_10_, i_7_, i_3_, i_13_, i_4_, i_12_, i_2_}, x6969x);
	defparam lut_954.LUT_SIZE = 9;
	defparam lut_954.mask = 512'h5f5fffff5f5fffffffffffffffffffff5f5fffff5f5fffffffffffffffffffff0500000003000300000000000000000005000000000000000000000000000000;

	lut_sub lut_957 ({sk[0], i_9_, i_10_, i_7_, i_8_, i_13_, i_4_, i_12_, i_11_}, x6970x);
	defparam lut_957.LUT_SIZE = 9;
	defparam lut_957.mask = 512'h5f5fffff5f5fffffffffffffffffffff5f5fffff5f5fffffffffffffffffffff0100010001000300000000000000030000000000000000000000000000000000;

	lut_sub lut_960 ({sk[1], i_10_, i_7_, i_8_}, n_n592);
	defparam lut_960.LUT_SIZE = 4;
	defparam lut_960.mask = 16'h5508;

	lut_sub lut_962 ({sk[2], i_10_, i_7_, i_8_, i_3_, i_13_, i_12_, i_11_}, x614x);
	defparam lut_962.LUT_SIZE = 8;
	defparam lut_962.mask = 256'h7777777777777777ffffffffffffffff08080808080808080888080808cc0808;

	lut_sub lut_966 ({sk[3], i_10_, i_7_, i_8_, i_4_, i_12_, i_11_, i_2_}, x1107x);
	defparam lut_966.LUT_SIZE = 8;
	defparam lut_966.mask = 256'h7777777777777777ffffffffffffffff000008000000000000000c0000000000;

	lut_sub lut_969 ({sk[4], i_9_, i_10_, i_7_, i_3_, i_12_}, x1110x);
	defparam lut_969.LUT_SIZE = 6;
	defparam lut_969.mask = 64'h3333ffff00000002;

	lut_sub lut_971 ({sk[5], i_9_, i_10_, i_7_, i_8_, i_13_, i_4_, i_12_, i_2_}, x6978x);
	defparam lut_971.LUT_SIZE = 9;
	defparam lut_971.mask = 512'h5f5fffff5f5fffffffffffffffffffff5f5fffff5f5fffffffffffffffffffff0000000000880088000000000088008800000000008800880000101000881098;

	lut_sub lut_974 ({sk[6], i_9_, i_10_, i_7_, i_8_, i_3_, i_13_, i_11_, i_2_}, x6979x);
	defparam lut_974.LUT_SIZE = 9;
	defparam lut_974.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff000000000000000000cc000000000000000000000505050500cc000005050505;

	lut_sub lut_977 ({sk[7], i_9_, i_10_, i_13_}, x367x);
	defparam lut_977.LUT_SIZE = 4;
	defparam lut_977.mask = 16'h1f01;

	lut_sub lut_979 ({sk[8], i_9_, i_10_, i_7_, i_8_, i_4_, i_12_, i_11_, i_2_}, x1108x);
	defparam lut_979.LUT_SIZE = 9;
	defparam lut_979.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff0000000000000000000005000000000000000000000005001100050011000500;

	lut_sub lut_983 ({sk[9], i_9_, i_10_, i_7_, i_13_, i_12_, i_11_, i_2_}, x6986x);
	defparam lut_983.LUT_SIZE = 8;
	defparam lut_983.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffff0088000000dd00000088000000dd00c0;

	lut_sub lut_988 ({sk[10], i_9_, i_10_, i_7_, i_8_, i_12_, i_11_, i_2_}, x7974x);
	defparam lut_988.LUT_SIZE = 8;
	defparam lut_988.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffffffffffffffffffffff77ff0f22222a0a;

	lut_sub lut_997 ({sk[11], i_9_, i_7_, i_8_}, n_n764);
	defparam lut_997.LUT_SIZE = 4;
	defparam lut_997.mask = 16'h1f10;

	lut_sub lut_999 ({sk[12], i_13_, i_12_}, n_n570);
	defparam lut_999.LUT_SIZE = 3;
	defparam lut_999.mask = 8'h38;

	lut_sub lut_1001 ({sk[13], i_9_, i_8_, i_3_, i_13_, i_4_, i_12_, i_11_, i_2_}, x630x);
	defparam lut_1001.LUT_SIZE = 9;
	defparam lut_1001.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff404a000000000000405f000000550000000a000000000000000a000000000000;

	lut_sub lut_1005 ({sk[14], i_9_, i_8_, i_3_, i_13_, i_4_, i_12_, i_11_, i_2_}, x629x);
	defparam lut_1005.LUT_SIZE = 9;
	defparam lut_1005.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff0022000000000000202200000022000000220000000000002022000000000000;

	lut_sub lut_1009 ({sk[15], i_10_, i_8_, i_3_, i_13_, i_4_, i_12_, i_11_}, x628x);
	defparam lut_1009.LUT_SIZE = 8;
	defparam lut_1009.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffff23000300000000002200000000000000;

	lut_sub lut_1012 ({sk[0], i_4_, i_1_, i_0_}, n_n791);
	defparam lut_1012.LUT_SIZE = 4;
	defparam lut_1012.mask = 16'h1f08;

	lut_sub lut_1014 ({sk[1], i_5_, i_4_, i_1_, i_2_, i_0_}, x659x);
	defparam lut_1014.LUT_SIZE = 6;
	defparam lut_1014.mask = 64'h0000ffff00c00080;

	lut_sub lut_1017 ({sk[2], i_7_, i_5_, i_6_, i_3_, i_4_, i_12_, i_1_}, x7004x);
	defparam lut_1017.LUT_SIZE = 8;
	defparam lut_1017.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffff0a008a88000000000000888800000000;

	lut_sub lut_1020 ({sk[3], i_7_, i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x7005x);
	defparam lut_1020.LUT_SIZE = 8;
	defparam lut_1020.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffff00e0000000a0000000c0000000000000;

	lut_sub lut_1023 ({sk[4], i_9_, i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x7007x);
	defparam lut_1023.LUT_SIZE = 8;
	defparam lut_1023.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffff0080000000c000000080000000800000;

	lut_sub lut_1026 ({sk[5], i_8_, i_12_, n_n764, x274x, x407x, x7043x, x690x, x7042x}, n_n914);
	defparam lut_1026.LUT_SIZE = 9;
	defparam lut_1026.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff5fff5fff7fff7fff00ff00ff33ff33ff5fffffff7fffffff00ff00ff33ff33ff;

	lut_sub lut_1032 ({sk[6], i_9_, i_10_, i_11_, x392x, x275x, x693x, x1012x, x7047x}, n_n913);
	defparam lut_1032.LUT_SIZE = 9;
	defparam lut_1032.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff7fffffff7777ffff7f7fffff7777ffff7f7fffff7777ffff7f7fffff7777ffff;

	lut_sub lut_1038 ({sk[7], i_6_, i_3_, i_1_, i_0_, n_n764, x7052x, x1004x, x1007x}, x696x);
	defparam lut_1038.LUT_SIZE = 9;
	defparam lut_1038.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff7f7f7f7f7f7f7f7f7f7f7f7f7f7f7f7fffff7f7f7fff7f7fffff7f7f7f7f7f7f;

	lut_sub lut_1044 ({sk[8], i_10_, i_7_, i_8_, i_11_, x41x, x1081x, x7009x, x1075x}, n_n911);
	defparam lut_1044.LUT_SIZE = 9;
	defparam lut_1044.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff7fff55557f7f55557f7f55557f7f55557f7f55557f7f55557f7f55557f7f5555;

	lut_sub lut_1049 ({sk[9], i_5_, i_3_, i_1_, i_11_, n_n792, x7017x, x7018x, x7019x}, n_n910);
	defparam lut_1049.LUT_SIZE = 9;
	defparam lut_1049.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff7fff55557f7f55557f7f55557f7f55557f7f55557f7f55557f7f55557f7f5555;

	lut_sub lut_1054 ({sk[10], i_5_, i_4_, x336x, n_n699, n_n678, x676x, x7028x, x7029x}, n_n918);
	defparam lut_1054.LUT_SIZE = 9;
	defparam lut_1054.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff777777ff777777ff7f7f7fffffffffff777777ff777777ff7f7f7fff7f7f7fff;

	lut_sub lut_1060 ({sk[11], i_9_, i_7_, i_6_, i_1_, i_2_, i_0_, x679x, x1041x}, x678x);
	defparam lut_1060.LUT_SIZE = 9;
	defparam lut_1060.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff7575757555555555f5757575f555f5557575757555555555f5757575f5555555;

	lut_sub lut_1065 ({sk[12], x406x, x7021x, x7038x, x7970x, x7987x}, x7039x);
	defparam lut_1065.LUT_SIZE = 6;
	defparam lut_1065.mask = 64'h0000ffffdfffffff;

	lut_sub lut_1071 ({sk[13], i_5_, i_12_, i_11_, i_0_, x984x, x985x, x986x, x987x}, x7062x);
	defparam lut_1071.LUT_SIZE = 9;
	defparam lut_1071.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffffffff7fff7fff7fffffff7fff7fff7fffffff7fff7fff7fff7fff7fff7fff7fff;

	lut_sub lut_1078 ({sk[14], i_10_, i_5_, i_3_, i_1_, i_2_}, x274x);
	defparam lut_1078.LUT_SIZE = 6;
	defparam lut_1078.mask = 64'h0000ffff80000000;

	lut_sub lut_1080 ({sk[15], i_10_, i_7_, i_8_}, n_n792);
	defparam lut_1080.LUT_SIZE = 4;
	defparam lut_1080.mask = 16'h1f80;

	lut_sub lut_1082 ({sk[0], i_10_, i_7_, i_8_, i_5_, i_4_, i_1_}, x378x);
	defparam lut_1082.LUT_SIZE = 7;
	defparam lut_1082.mask = 128'h1f5f1f5f1f5f1f5f2000000000000000;

	lut_sub lut_1084 ({sk[1], i_9_, i_10_, i_13_, i_12_, i_11_}, x305x);
	defparam lut_1084.LUT_SIZE = 6;
	defparam lut_1084.mask = 64'h0000ffff80000000;

	lut_sub lut_1086 ({sk[2], i_10_, i_7_, i_8_, i_5_, i_3_, i_13_, i_12_, i_11_}, x964x);
	defparam lut_1086.LUT_SIZE = 9;
	defparam lut_1086.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffffa0000000c0000000e0c00000c0c0000000000000000000000000000000000000;

	lut_sub lut_1090 ({sk[3], i_10_, i_7_, i_5_, i_3_, i_13_, i_4_, i_11_}, x7080x);
	defparam lut_1090.LUT_SIZE = 8;
	defparam lut_1090.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffffb0a00000300000000000000000000000;

	lut_sub lut_1093 ({sk[4], i_9_, i_10_, i_6_, i_13_, i_12_, i_1_, i_11_, i_0_}, x959x);
	defparam lut_1093.LUT_SIZE = 9;
	defparam lut_1093.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff4040000050000000000000000000000000000000000000000000000000000000;

	lut_sub lut_1096 ({sk[5], i_10_, i_7_, i_5_, i_6_, i_13_, i_12_, i_2_, i_0_}, x960x);
	defparam lut_1096.LUT_SIZE = 9;
	defparam lut_1096.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff0000000000000000400000000000000000000000000000000000000000000000;

	lut_sub lut_1098 ({sk[6], i_1_, i_2_, i_0_, x305x, x964x, x7080x, x959x, x960x}, n_n971);
	defparam lut_1098.LUT_SIZE = 9;
	defparam lut_1098.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff777777777fffffff777777777777ffff77777777777777777777777777777777;

	lut_sub lut_1104 ({sk[7], i_10_, i_13_, i_12_}, n_n575);
	defparam lut_1104.LUT_SIZE = 4;
	defparam lut_1104.mask = 16'h1f80;

	lut_sub lut_1106 ({sk[8], i_5_, i_6_, i_3_, i_2_, i_0_}, x413x);
	defparam lut_1106.LUT_SIZE = 6;
	defparam lut_1106.mask = 64'h0000ffff40000000;

	lut_sub lut_1108 ({sk[9], i_7_, i_8_, i_5_, i_6_, i_3_, i_2_, i_0_}, x534x);
	defparam lut_1108.LUT_SIZE = 8;
	defparam lut_1108.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffff55000000500000004400000040000000;

	lut_sub lut_1113 ({sk[10], i_10_, i_7_, i_8_, i_6_, i_13_, i_12_, i_11_}, x533x);
	defparam lut_1113.LUT_SIZE = 8;
	defparam lut_1113.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffffa000c000000000000000000000000000;

	lut_sub lut_1116 ({sk[11], i_8_, i_5_, i_6_, i_3_, i_11_, i_2_, i_0_}, x532x);
	defparam lut_1116.LUT_SIZE = 8;
	defparam lut_1116.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffff40400000000000004440000000000000;

	lut_sub lut_1119 ({sk[12], i_5_, i_3_, i_0_}, x7083x);
	defparam lut_1119.LUT_SIZE = 4;
	defparam lut_1119.mask = 16'h1f40;

	lut_sub lut_1121 ({sk[13], i_10_, i_13_, i_4_}, x7085x);
	defparam lut_1121.LUT_SIZE = 4;
	defparam lut_1121.mask = 16'h1f40;

	lut_sub lut_1123 ({sk[14], i_10_, i_8_, i_13_, i_11_}, x7086x);
	defparam lut_1123.LUT_SIZE = 5;
	defparam lut_1123.mask = 32'h11ff8000;

	lut_sub lut_1125 ({sk[15], n_n575, x413x, x534x, x533x, x532x, x7083x, x7085x, x7086x}, n_n970);
	defparam lut_1125.LUT_SIZE = 9;
	defparam lut_1125.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff00000f0f33333f3f55555f5f77777f7f00ff0fff33ff3fff55ff5fff77ff7fff;

	lut_sub lut_1130 ({sk[0], i_9_, i_10_, i_13_, i_12_, i_11_}, x303x);
	defparam lut_1130.LUT_SIZE = 6;
	defparam lut_1130.mask = 64'h0000ffff20000000;

	lut_sub lut_1132 ({sk[1], i_7_, i_8_, i_3_, i_2_}, x536x);
	defparam lut_1132.LUT_SIZE = 5;
	defparam lut_1132.mask = 32'h11ffeac0;

	lut_sub lut_1135 ({sk[2], i_9_, i_10_, i_8_, i_3_, i_13_, i_12_, i_11_}, x44x);
	defparam lut_1135.LUT_SIZE = 8;
	defparam lut_1135.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffffa0008000000000000000000000000000;

	lut_sub lut_1138 ({sk[3], i_9_, i_10_, i_7_, i_8_, i_3_, i_12_, i_11_, i_2_}, x538x);
	defparam lut_1138.LUT_SIZE = 9;
	defparam lut_1138.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff8888f888a0a0f0a0000000000000000000000000000000000000000000000000;

	lut_sub lut_1142 ({sk[4], i_9_, i_10_, i_13_, i_4_, i_12_, i_11_, i_2_}, x7092x);
	defparam lut_1142.LUT_SIZE = 8;
	defparam lut_1142.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffff80ff0000000000000000000000000000;

	lut_sub lut_1145 ({sk[5], i_5_, i_13_, i_0_, x303x, x536x, x44x, x538x, x7092x}, n_n972);
	defparam lut_1145.LUT_SIZE = 9;
	defparam lut_1145.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff000000007f7f7f7f000000005f5f5f5f000000ff7f7f7fff000000ff5f5f5fff;

	lut_sub lut_1150 ({sk[6], i_5_, i_6_, i_2_}, n_n624);
	defparam lut_1150.LUT_SIZE = 4;
	defparam lut_1150.mask = 16'h1f02;

	lut_sub lut_1152 ({sk[7], i_9_, i_7_, i_8_, i_13_, i_4_, i_12_, i_11_}, x580x);
	defparam lut_1152.LUT_SIZE = 8;
	defparam lut_1152.mask = 256'h5f5f5f5fffffffff5f5f5f5fffffffffaa00af0088008f000000000000000000;

	lut_sub lut_1156 ({sk[8], i_9_, i_8_, i_13_, i_4_, i_12_, i_11_}, x579x);
	defparam lut_1156.LUT_SIZE = 7;
	defparam lut_1156.mask = 128'h1f5f1f5f1f5f1f5faf00cf0000000000;

	lut_sub lut_1160 ({sk[9], i_9_, i_7_, i_8_, i_6_, i_13_, i_4_, i_12_, i_2_}, x578x);
	defparam lut_1160.LUT_SIZE = 9;
	defparam lut_1160.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff00000000000000000000880000008f0000000000000000000000000000000000;

	lut_sub lut_1163 ({sk[10], i_9_, i_7_, i_5_, i_13_, i_1_, i_11_, i_2_, i_0_}, x925x);
	defparam lut_1163.LUT_SIZE = 9;
	defparam lut_1163.mask = 512'h3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff3f3fffff0000000040000000000000000000000000000000000000000000000000000000;

	lut_sub lut_1165 ({sk[11], i_5_, i_6_, i_3_, i_2_, i_0_}, x7097x);
	defparam lut_1165.LUT_SIZE = 6;
	defparam lut_1165.mask = 64'h0000ffff00000040;

	lut_sub lut_1167 ({sk[12], i_5_, i_0_, n_n624, x580x, x579x, x578x, x925x, x7097x}, n_n978);
	defparam lut_1167.LUT_SIZE = 9;
	defparam lut_1167.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff3377337733773377337733773377ffff33773377337733773f7f3f7f3f7fffff;

	lut_sub lut_1172 ({sk[13], i_5_, i_6_, i_1_, n_n787, x9x, n_n849, x294x, x666x}, x7107x);
	defparam lut_1172.LUT_SIZE = 9;
	defparam lut_1172.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff00005555000055553333777700005555000f555f000f555f000f555f000f555f;

	lut_sub lut_1176 ({sk[14], i_5_, i_6_, i_3_, i_1_, n_n816, x70x, x667x, x7103x}, x7108x);
	defparam lut_1176.LUT_SIZE = 9;
	defparam lut_1176.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff5f7f5f7f0f3f0f3f5f7f0f3f0f3f0f3f0f3f0f3f0f3f0f3f0f3f0f3f0f3f0f3f;

	lut_sub lut_1181 ({sk[15], i_9_, i_8_, i_5_, i_6_, i_4_, i_2_, n_n277, x7967x}, x670x);
	defparam lut_1181.LUT_SIZE = 9;
	defparam lut_1181.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffffaaaaaaaaaaaababaaaaaaaaaaaaabafaaaaaaaaaaaaababaaaaaaaaaaaaababa;

	lut_sub lut_1185 ({sk[0], i_10_, i_8_, i_5_, i_13_, i_12_, i_11_, n_n675, x669x}, x7113x);
	defparam lut_1185.LUT_SIZE = 9;
	defparam lut_1185.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff0050000000500000035000000050000000500000005000000050000000500000;

	lut_sub lut_1188 ({sk[1], i_7_, i_5_, i_6_, i_1_, i_11_, i_2_, n_n570, x317x}, x674x);
	defparam lut_1188.LUT_SIZE = 9;
	defparam lut_1188.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff0010001000100010001000100010001000300030003000100010001000100010;

	lut_sub lut_1192 ({sk[2], i_5_, n_n816, x9x, x29x, x19x, x282x, x671x, x893x}, x7116x);
	defparam lut_1192.LUT_SIZE = 9;
	defparam lut_1192.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff555f5f5f555f5f5f777f7f7fffffffff55555555555555557777777777777777;

	lut_sub lut_1198 ({sk[3], i_13_, i_12_, i_11_}, n_n716);
	defparam lut_1198.LUT_SIZE = 4;
	defparam lut_1198.mask = 16'h5f20;

	lut_sub lut_1200 ({sk[4], i_9_, i_13_, i_11_}, n_n719);
	defparam lut_1200.LUT_SIZE = 4;
	defparam lut_1200.mask = 16'h5f80;

	lut_sub lut_1202 ({sk[5], i_7_, i_8_, i_6_}, n_n837);
	defparam lut_1202.LUT_SIZE = 4;
	defparam lut_1202.mask = 16'h5f04;

	lut_sub lut_1204 ({sk[6], i_9_, i_8_, i_5_, i_6_, i_3_, i_1_, i_2_}, x713x);
	defparam lut_1204.LUT_SIZE = 8;
	defparam lut_1204.mask = 256'h00ff33ff33ff33ff55ff77ff77ff77ff000080a0000000000000000000000000;

	lut_sub lut_1207 ({sk[7], i_9_, i_5_, i_6_, i_13_, i_12_, i_1_, i_0_}, x882x);
	defparam lut_1207.LUT_SIZE = 8;
	defparam lut_1207.mask = 256'h00ff33ff33ff33ff55ff77ff77ff77ff00000000000040000000000000000000;

	lut_sub lut_1209 ({sk[8], i_5_, i_3_, i_0_, n_n716, n_n719, n_n837, x713x, x882x}, x7125x);
	defparam lut_1209.LUT_SIZE = 9;
	defparam lut_1209.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff5555777755557777555577775555777755557777555f777f5555777755557777;

	lut_sub lut_1213 ({sk[9], n_n838, x26x, x284x, x875x, x7129x, x873x, x874x, x637x}, n_n979);
	defparam lut_1213.LUT_SIZE = 9;
	defparam lut_1213.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff00000000555555553f3f3f3f7f7f7f7f00ffffff55ffffff3fffffff7fffffff;

	lut_sub lut_1219 ({sk[10], i_8_, i_5_, i_11_, n_n761, x37x, n_n835, x763x, x864x}, x858x);
	defparam lut_1219.LUT_SIZE = 9;
	defparam lut_1219.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff0000000000000000555f777f555f555f00000000000000005555777755555555;

	lut_sub lut_1223 ({sk[11], x37x, x13x, x19x, x405x, x361x, x861x, x862x, x7131x}, x7141x);
	defparam lut_1223.LUT_SIZE = 9;
	defparam lut_1223.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff0000ffff00ffffff3f3fffff3fffffff5555ffff55ffffff7f7fffff7fffffff;

	lut_sub lut_1229 ({sk[12], i_7_, i_8_, i_5_, i_4_, i_1_, i_0_, x722x, x7146x}, x721x);
	defparam lut_1229.LUT_SIZE = 9;
	defparam lut_1229.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff5555777755555555555577775555555555557777555555555555f77755555555;

	lut_sub lut_1233 ({sk[13], i_7_, i_5_, i_0_, n_n819, x301x, x284x, x361x, x7143x}, x7149x);
	defparam lut_1233.LUT_SIZE = 9;
	defparam lut_1233.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff050505ff050505050505050505050505373737ff373737373737373737373737;

	lut_sub lut_1237 ({sk[14], i_9_, i_8_, i_13_, i_4_, i_12_, i_11_}, x735x);
	defparam lut_1237.LUT_SIZE = 7;
	defparam lut_1237.mask = 128'h0f3fffff3f3fffffaf00cf0000000000;

	lut_sub lut_1241 ({sk[15], i_9_, i_7_, i_8_, i_13_, i_4_, i_12_, i_1_, i_11_}, x802x);
	defparam lut_1241.LUT_SIZE = 9;
	defparam lut_1241.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff80800000808000008080000080cc000000000000000000000000000000000000;

	lut_sub lut_1244 ({sk[0], i_9_, i_7_, i_8_, i_6_, i_3_, i_13_, i_12_, i_11_}, x803x);
	defparam lut_1244.LUT_SIZE = 9;
	defparam lut_1244.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff0000000000000000000080000000c00000000000000000000000000000000000;

	lut_sub lut_1247 ({sk[1], i_9_, i_7_, i_5_, i_6_, i_3_, i_13_, i_4_, i_0_}, x798x);
	defparam lut_1247.LUT_SIZE = 9;
	defparam lut_1247.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff0000000000000000000000000000100000000000000000000000000000000000;

	lut_sub lut_1249 ({sk[2], i_7_, i_5_, i_3_, i_1_, i_0_}, x7174x);
	defparam lut_1249.LUT_SIZE = 6;
	defparam lut_1249.mask = 64'h33773f7f00000040;

	lut_sub lut_1251 ({sk[3], i_9_, i_5_, i_6_, i_13_, i_1_, i_11_, i_0_}, x800x);
	defparam lut_1251.LUT_SIZE = 8;
	defparam lut_1251.mask = 256'h00ff33ff33ff33ff55ff77ff77ff77ff00000000400000000000000000000000;

	lut_sub lut_1253 ({sk[4], i_5_, i_0_, x735x, x802x, x803x, x798x, x7174x, x800x}, n_n977);
	defparam lut_1253.LUT_SIZE = 9;
	defparam lut_1253.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff5f5f5f5f7f7f7f7f5f5f5f5f7f7f7f7f5f5f5f5f7f7f7f7f5fffffff7fffffff;

	lut_sub lut_1259 ({sk[5], x272x, x591x, x590x, x7208x, x7209x, x7210x, x238x, x7211x}, n_n988);
	defparam lut_1259.LUT_SIZE = 9;
	defparam lut_1259.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff777777ff777777ff7f7f7fff7f7f7fff777777ffffffffff7f7f7fffffffffff;

	lut_sub lut_1265 ({sk[6], i_8_, i_4_, x657x, x772x, x773x, x776x, x7968x}, n_n991);
	defparam lut_1265.LUT_SIZE = 8;
	defparam lut_1265.mask = 256'h00ff33ff33ff33ff55ff77ff77ff77ffbfffbfff0fff0fffbfffffff0fff0fff;

	lut_sub lut_1271 ({sk[7], i_9_, i_10_, i_5_, i_12_, i_11_, i_0_, n_n752, x411x}, x687x);
	defparam lut_1271.LUT_SIZE = 9;
	defparam lut_1271.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff5555555555555555555555555555555555557555555555555555775755555555;

	lut_sub lut_1275 ({sk[8], i_9_, i_3_, i_12_, i_2_, i_0_, x686x, x7189x, x368x}, x7192x);
	defparam lut_1275.LUT_SIZE = 9;
	defparam lut_1275.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff55555555555555555555555f5555555f55555555555555555555555f5555777f;

	lut_sub lut_1279 ({sk[9], n_n541, x22x, x115x, x737x, x736x, x739x, x225x, x7218x}, x7233x);
	defparam lut_1279.LUT_SIZE = 9;
	defparam lut_1279.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff33337777ffffffff3f3f7f7fffffffff33ff77ffffffffff3fff7fffffffffff;

	lut_sub lut_1285 ({sk[10], i_6_, i_4_, i_2_, i_0_, x355x, x717x, x716x, x255x}, x7197x);
	defparam lut_1285.LUT_SIZE = 9;
	defparam lut_1285.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff5f5f5f5f7f7f7f7f55555555555555555f5f5fff7f7f7fff555555ff555555ff;

	lut_sub lut_1290 ({sk[11], i_5_, i_6_, i_4_, n_n818, n_n213, x218x, x212x, x213x}, x7231x);
	defparam lut_1290.LUT_SIZE = 9;
	defparam lut_1290.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff7f7f7fff777777777f7f7f7f777777777f7f7f7f777777777f7f7f7f77777777;

	lut_sub lut_1295 ({sk[12], i_9_, i_10_, i_1_, x557x, x46x, x276x, x190x, x7251x}, n_n1001);
	defparam lut_1295.LUT_SIZE = 9;
	defparam lut_1295.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff7777777777ff77ff7777ffff77ffffff7777777777ff77ff7777ffff7fffffff;

	lut_sub lut_1301 ({sk[13], i_10_, i_7_, i_12_, i_11_, x560x, x559x, x174x, x175x}, n_n1000);
	defparam lut_1301.LUT_SIZE = 9;
	defparam lut_1301.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff77ff77ff7777777777ff77ff777777777fff77ff7f7f777777ff77ff77777777;

	lut_sub lut_1306 ({sk[14], i_9_, i_10_, i_1_, i_11_, i_0_, x565x, x563x, x161x}, x7262x);
	defparam lut_1306.LUT_SIZE = 9;
	defparam lut_1306.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff55555555555555555555555555555555555555555f5f5f5f555577775fff7fff;

	lut_sub lut_1311 ({sk[15], i_8_, x597x, x596x, x127x, x128x, x7284x, x130x, x7289x}, n_n998);
	defparam lut_1311.LUT_SIZE = 9;
	defparam lut_1311.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff77ffffffffffffff7fffffffffffffff77ffffff77ffffff7fffffff7fffffff;

	lut_sub lut_1318 ({sk[0], i_10_, i_8_, i_11_, x359x, x705x, x7300x, x750x, x88x}, x7311x);
	defparam lut_1318.LUT_SIZE = 9;
	defparam lut_1318.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff7f7f7f7f7f7f7f7f5f5f5f5f5f5f5f5f7f7fffff7fff7fff5f5f5f5f5fff5fff;

	lut_sub lut_1324 ({sk[1], i_10_, i_7_, i_8_, i_3_, x749x, x87x, x7965x}, x7308x);
	defparam lut_1324.LUT_SIZE = 8;
	defparam lut_1324.mask = 256'h00ff33ff33ff33ff55ff77ff77ff77ff3333333333333333333f3333bbbf3333;

	lut_sub lut_1328 ({sk[2], i_10_, i_7_, i_8_, i_5_, i_13_, i_4_, i_12_, i_11_}, x757x);
	defparam lut_1328.LUT_SIZE = 9;
	defparam lut_1328.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffffaf000000cf000000000000000000000000000000000000000000000000000000;

	lut_sub lut_1332 ({sk[3], i_10_, i_8_, i_5_, i_13_, i_4_, i_1_, i_2_, i_0_}, x40x);
	defparam lut_1332.LUT_SIZE = 9;
	defparam lut_1332.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff0040000000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_1334 ({sk[4], i_10_, i_5_, i_6_, i_13_, i_1_, i_11_, i_0_}, x48x);
	defparam lut_1334.LUT_SIZE = 8;
	defparam lut_1334.mask = 256'h00ff33ff33ff33ff55ff77ff77ff77ff40000000000000000000000000000000;

	lut_sub lut_1336 ({sk[5], i_3_, i_1_, i_0_, x313x, x9x, x757x, x40x, x48x}, x7331x);
	defparam lut_1336.LUT_SIZE = 9;
	defparam lut_1336.mask = 512'h00ffffff00ffffff00ffffff00ffffff00ffffff33ffffff55ffffff77ffffff777777ff7f7f7fff777777ff777777ff777777ff777777ff777777ff777777ff;

	lut_sub lut_1341 ({sk[6], i_13_, i_12_, i_11_}, n_n853);
	defparam lut_1341.LUT_SIZE = 4;
	defparam lut_1341.mask = 16'h5f10;

	lut_sub lut_1343 ({sk[7], i_9_, i_10_, i_13_, i_4_, i_12_, i_11_}, n_n2368);
	defparam lut_1343.LUT_SIZE = 7;
	defparam lut_1343.mask = 128'h0f3fffff3f3fffff0100000000000000;

	lut_sub lut_1345 ({sk[8], i_13_, i_4_, i_12_, i_11_}, x17x);
	defparam lut_1345.LUT_SIZE = 5;
	defparam lut_1345.mask = 32'h55ff0100;

	lut_sub lut_1347 ({sk[9], i_10_, i_13_, i_4_, i_12_}, x37x);
	defparam lut_1347.LUT_SIZE = 5;
	defparam lut_1347.mask = 32'h55ff1000;

	lut_sub lut_1349 ({sk[10], i_10_, i_8_, i_1_, i_2_, i_0_}, x6718x);
	defparam lut_1349.LUT_SIZE = 6;
	defparam lut_1349.mask = 64'h33773f7f80000000;

	lut_sub lut_1351 ({sk[11], i_10_, i_12_, i_11_}, n_n822);
	defparam lut_1351.LUT_SIZE = 4;
	defparam lut_1351.mask = 16'h5f10;

	lut_sub lut_1353 ({sk[12], i_9_, i_10_, i_13_, i_4_, i_12_, i_11_}, x266x);
	defparam lut_1353.LUT_SIZE = 7;
	defparam lut_1353.mask = 128'h0f3fffff3f3fffff0100000000000000;

	lut_sub lut_1355 ({sk[13], i_9_, i_8_, i_5_, i_6_}, x322x);
	defparam lut_1355.LUT_SIZE = 5;
	defparam lut_1355.mask = 32'h33ff0100;

	lut_sub lut_1357 ({sk[14], i_10_, i_8_, i_6_, i_2_}, x336x);
	defparam lut_1357.LUT_SIZE = 5;
	defparam lut_1357.mask = 32'h33ff8000;

	lut_sub lut_1359 ({sk[15], i_10_, i_8_, i_6_, i_4_, i_2_, i_0_}, x394x);
	defparam lut_1359.LUT_SIZE = 7;
	defparam lut_1359.mask = 128'h55ff55ff55ff55ff0800000000000000;

	lut_sub lut_1361 ({sk[0], i_1_, i_2_, i_0_}, n_n838);
	defparam lut_1361.LUT_SIZE = 4;
	defparam lut_1361.mask = 16'h7740;

	lut_sub lut_1363 ({sk[1], i_6_, i_1_, i_2_, i_0_}, x420x);
	defparam lut_1363.LUT_SIZE = 5;
	defparam lut_1363.mask = 32'h33ff4440;

	lut_sub lut_1366 ({sk[2], i_5_, i_4_, i_1_}, x6719x);
	defparam lut_1366.LUT_SIZE = 4;
	defparam lut_1366.mask = 16'h7710;

	lut_sub lut_1368 ({sk[3], i_9_, i_10_, i_7_, i_8_, i_13_, i_11_}, x6720x);
	defparam lut_1368.LUT_SIZE = 7;
	defparam lut_1368.mask = 128'h55ff55ff55ff55ff4000000000000000;

	lut_sub lut_1370 ({sk[4], i_8_, i_5_, i_4_, i_1_, i_2_}, x6724x);
	defparam lut_1370.LUT_SIZE = 6;
	defparam lut_1370.mask = 64'h3f3f3f3f08000000;

	lut_sub lut_1372 ({sk[5], i_9_, i_10_, i_8_, i_13_, i_4_, i_12_, i_11_}, x6721x);
	defparam lut_1372.LUT_SIZE = 8;
	defparam lut_1372.mask = 256'h55ff7fff55ff7fff55ff7fff55ff7fff01000000000000000000000000000000;

	lut_sub lut_1374 ({sk[6], i_5_, i_13_, i_4_, i_12_, i_11_}, x6722x);
	defparam lut_1374.LUT_SIZE = 6;
	defparam lut_1374.mask = 64'h3f3f3f3f01000000;

	lut_sub lut_1376 ({sk[7], i_10_, i_13_, i_4_, i_12_, i_2_}, x6723x);
	defparam lut_1376.LUT_SIZE = 6;
	defparam lut_1376.mask = 64'h3f3f3f3f01000000;

	lut_sub lut_1378 ({sk[8], i_8_, i_1_, i_2_}, x6725x);
	defparam lut_1378.LUT_SIZE = 4;
	defparam lut_1378.mask = 16'h7701;

	lut_sub lut_1380 ({sk[9], i_1_, i_2_, i_0_}, n_n835);
	defparam lut_1380.LUT_SIZE = 4;
	defparam lut_1380.mask = 16'h7780;

	lut_sub lut_1382 ({sk[10], i_10_, i_13_, i_12_, i_11_}, n_n725);
	defparam lut_1382.LUT_SIZE = 5;
	defparam lut_1382.mask = 32'h33ff2000;

	lut_sub lut_1384 ({sk[11], i_10_, i_1_, i_2_, i_0_, n_n538, n_n748, n_n716, n_n746}, x421x);
	defparam lut_1384.LUT_SIZE = 9;
	defparam lut_1384.mask = 512'h00ff00ffffffffff55ff55ffffffffff00ff00ffffffffff55ff55ffffffffff0003000000000000001100000000000000030000000000000000000000000000;

	lut_sub lut_1387 ({sk[12], i_7_, i_2_}, x29x);
	defparam lut_1387.LUT_SIZE = 3;
	defparam lut_1387.mask = 8'h12;

	lut_sub lut_1389 ({sk[13], i_8_, i_3_, i_13_, i_12_, i_1_, i_11_, i_2_}, x1371x);
	defparam lut_1389.LUT_SIZE = 8;
	defparam lut_1389.mask = 256'h5555ffff5555ffff5555ffffffffffff00000000000000002000000000000000;

	lut_sub lut_1391 ({sk[14], i_9_, i_7_, i_6_}, n_n819);
	defparam lut_1391.LUT_SIZE = 4;
	defparam lut_1391.mask = 16'h5710;

	lut_sub lut_1393 ({sk[15], i_3_, i_1_, i_2_}, n_n273);
	defparam lut_1393.LUT_SIZE = 4;
	defparam lut_1393.mask = 16'h5720;

	lut_sub lut_1395 ({sk[0], i_1_, i_2_, i_0_}, n_n847);
	defparam lut_1395.LUT_SIZE = 4;
	defparam lut_1395.mask = 16'h5720;

	lut_sub lut_1397 ({sk[1], i_7_, i_6_}, x28x);
	defparam lut_1397.LUT_SIZE = 3;
	defparam lut_1397.mask = 8'h18;

	lut_sub lut_1399 ({sk[2], i_10_, i_11_}, n_n213);
	defparam lut_1399.LUT_SIZE = 3;
	defparam lut_1399.mask = 8'h11;

	lut_sub lut_1401 ({sk[3], i_12_, i_11_}, n_n311);
	defparam lut_1401.LUT_SIZE = 3;
	defparam lut_1401.mask = 8'h14;

	lut_sub lut_1403 ({sk[4], i_5_, i_6_}, x13x);
	defparam lut_1403.LUT_SIZE = 3;
	defparam lut_1403.mask = 8'h12;

	lut_sub lut_1405 ({sk[5], i_7_, i_8_, i_5_}, n_n185);
	defparam lut_1405.LUT_SIZE = 4;
	defparam lut_1405.mask = 16'h5702;

	lut_sub lut_1407 ({sk[6], i_3_, i_1_, i_0_}, n_n826);
	defparam lut_1407.LUT_SIZE = 4;
	defparam lut_1407.mask = 16'h5701;

	lut_sub lut_1409 ({sk[7], i_10_, i_7_, i_6_}, n_n699);
	defparam lut_1409.LUT_SIZE = 4;
	defparam lut_1409.mask = 16'h5780;

	lut_sub lut_1411 ({sk[8], i_3_, i_4_, i_0_}, n_n678);
	defparam lut_1411.LUT_SIZE = 4;
	defparam lut_1411.mask = 16'h5720;

	lut_sub lut_1413 ({sk[9], i_5_, i_6_}, x26x);
	defparam lut_1413.LUT_SIZE = 3;
	defparam lut_1413.mask = 8'h14;

	lut_sub lut_1415 ({sk[10], i_13_, i_4_, i_11_}, x370x);
	defparam lut_1415.LUT_SIZE = 4;
	defparam lut_1415.mask = 16'h5710;

	lut_sub lut_1417 ({sk[11], i_10_, i_7_, i_8_, i_5_, i_6_, i_13_, i_4_, i_11_}, x70x);
	defparam lut_1417.LUT_SIZE = 9;
	defparam lut_1417.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff1000000000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_1419 ({sk[12], i_9_, i_5_, i_13_, i_4_, i_12_, i_1_, i_11_}, x450x);
	defparam lut_1419.LUT_SIZE = 8;
	defparam lut_1419.mask = 256'h5555ffff5555ffff5555ffffffffffff00050000000100000004000000000000;

	lut_sub lut_1422 ({sk[13], i_10_, i_5_, i_6_, i_13_, i_12_, i_1_, i_11_, i_0_}, x451x);
	defparam lut_1422.LUT_SIZE = 9;
	defparam lut_1422.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff0101000001010000013300000103000000000000000000000000000000000000;

	lut_sub lut_1426 ({sk[14], i_8_, i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x455x);
	defparam lut_1426.LUT_SIZE = 8;
	defparam lut_1426.mask = 256'h5555ffff5555ffff5555ffffffffffff00000000000000000100100000002000;

	lut_sub lut_1430 ({sk[15], i_5_, i_6_, i_3_, i_13_, i_1_, i_11_, i_2_, i_0_}, x454x);
	defparam lut_1430.LUT_SIZE = 9;
	defparam lut_1430.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff0000000000002000000000000000002000000000000010000000000000000011;

	lut_sub lut_1435 ({sk[0], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x453x);
	defparam lut_1435.LUT_SIZE = 7;
	defparam lut_1435.mask = 128'h0037ffff0037ffff0080000000400000;

	lut_sub lut_1438 ({sk[1], i_10_, i_7_, i_13_, i_12_}, x6631x);
	defparam lut_1438.LUT_SIZE = 5;
	defparam lut_1438.mask = 32'h333f0020;

	lut_sub lut_1440 ({sk[2], i_7_, i_8_, i_6_}, n_n752);
	defparam lut_1440.LUT_SIZE = 4;
	defparam lut_1440.mask = 16'h5701;

	lut_sub lut_1442 ({sk[3], i_9_, i_5_, i_3_, i_4_}, x307x);
	defparam lut_1442.LUT_SIZE = 5;
	defparam lut_1442.mask = 32'h333f0002;

	lut_sub lut_1444 ({sk[4], i_13_, i_12_, i_1_, i_2_, i_0_, n_n541, n_n752, n_n756}, x457x);
	defparam lut_1444.LUT_SIZE = 9;
	defparam lut_1444.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff0500030000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_1447 ({sk[5], i_7_, i_8_, i_6_}, n_n832);
	defparam lut_1447.LUT_SIZE = 4;
	defparam lut_1447.mask = 16'h5708;

	lut_sub lut_1449 ({sk[6], i_9_, i_10_, i_13_, i_12_, i_11_}, n_n1574);
	defparam lut_1449.LUT_SIZE = 6;
	defparam lut_1449.mask = 64'h115511ff00000008;

	lut_sub lut_1451 ({sk[7], i_10_, i_7_, i_8_}, n_n597);
	defparam lut_1451.LUT_SIZE = 4;
	defparam lut_1451.mask = 16'h5702;

	lut_sub lut_1453 ({sk[8], i_3_, i_13_, i_1_, i_11_, i_2_, i_0_}, x6581x);
	defparam lut_1453.LUT_SIZE = 7;
	defparam lut_1453.mask = 128'h0037ffff0037ffff0000100000000000;

	lut_sub lut_1455 ({sk[9], i_10_, i_7_, i_8_, i_5_, i_6_, i_3_}, x6583x);
	defparam lut_1455.LUT_SIZE = 7;
	defparam lut_1455.mask = 128'h0037ffff0037ffff0000000040000000;

	lut_sub lut_1457 ({sk[10], i_7_, i_5_, i_6_, i_1_, i_2_, i_0_}, x465x);
	defparam lut_1457.LUT_SIZE = 7;
	defparam lut_1457.mask = 128'h0037ffff0037ffff7703550133031101;

	lut_sub lut_1463 ({sk[11], i_5_, i_6_, i_13_, i_12_, i_1_, i_0_}, x464x);
	defparam lut_1463.LUT_SIZE = 7;
	defparam lut_1463.mask = 128'h0037ffff0037ffff00ff008000800080;

	lut_sub lut_1466 ({sk[12], i_10_, i_7_, i_8_, i_5_, i_1_, i_11_}, x1702x);
	defparam lut_1466.LUT_SIZE = 7;
	defparam lut_1466.mask = 128'h0037ffff0037ffff0000000080000000;

	lut_sub lut_1468 ({sk[13], i_10_, i_7_, i_8_, i_11_}, x6588x);
	defparam lut_1468.LUT_SIZE = 5;
	defparam lut_1468.mask = 32'h333f0080;

	lut_sub lut_1470 ({sk[14], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x6590x);
	defparam lut_1470.LUT_SIZE = 7;
	defparam lut_1470.mask = 128'h0037ffff0037ffff0000000000080000;

	lut_sub lut_1472 ({sk[15], i_8_, i_3_}, x19x);
	defparam lut_1472.LUT_SIZE = 3;
	defparam lut_1472.mask = 8'h12;

	lut_sub lut_1474 ({sk[0], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x469x);
	defparam lut_1474.LUT_SIZE = 7;
	defparam lut_1474.mask = 128'h0037ffff0037ffff2000000000000100;

	lut_sub lut_1477 ({sk[1], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x467x);
	defparam lut_1477.LUT_SIZE = 7;
	defparam lut_1477.mask = 128'h0037ffff0037ffff0000080040000400;

	lut_sub lut_1481 ({sk[2], i_8_, i_5_, i_3_}, x6598x);
	defparam lut_1481.LUT_SIZE = 4;
	defparam lut_1481.mask = 16'h5780;

	lut_sub lut_1483 ({sk[3], i_9_, i_7_, i_6_, i_1_, i_2_, i_0_}, x6599x);
	defparam lut_1483.LUT_SIZE = 7;
	defparam lut_1483.mask = 128'h0037ffff0037ffff0000000000000002;

	lut_sub lut_1485 ({sk[4], i_7_, i_8_, i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x1691x);
	defparam lut_1485.LUT_SIZE = 9;
	defparam lut_1485.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff8000000000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_1487 ({sk[5], i_3_, i_4_, i_2_}, n_n672);
	defparam lut_1487.LUT_SIZE = 4;
	defparam lut_1487.mask = 16'h5720;

	lut_sub lut_1489 ({sk[6], i_9_, i_6_, i_4_}, n_n810);
	defparam lut_1489.LUT_SIZE = 4;
	defparam lut_1489.mask = 16'h5710;

	lut_sub lut_1491 ({sk[7], i_9_, i_10_, i_7_, i_12_, i_2_}, x407x);
	defparam lut_1491.LUT_SIZE = 6;
	defparam lut_1491.mask = 64'h115511ff08000000;

	lut_sub lut_1493 ({sk[8], i_10_, i_7_, i_8_, i_6_, i_3_, i_2_}, x470x);
	defparam lut_1493.LUT_SIZE = 7;
	defparam lut_1493.mask = 128'h0037ffff0037fffff0c0a00000000000;

	lut_sub lut_1497 ({sk[9], i_9_, i_10_, i_3_, i_13_, i_12_, i_1_, i_11_, i_2_}, x1340x);
	defparam lut_1497.LUT_SIZE = 9;
	defparam lut_1497.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff0c00000008000000000000000000000000000000000000000000000000000000;

	lut_sub lut_1500 ({sk[10], i_9_, i_10_, i_8_, i_6_, i_3_, i_13_, i_12_, i_11_}, x1341x);
	defparam lut_1500.LUT_SIZE = 9;
	defparam lut_1500.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff0000200000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_1502 ({sk[11], i_10_, i_6_, i_3_, i_13_, i_4_, i_11_, i_2_}, x1342x);
	defparam lut_1502.LUT_SIZE = 8;
	defparam lut_1502.mask = 256'h5555ffff5555ffff5555ffffffffffff02000000000000000000000000000000;

	lut_sub lut_1504 ({sk[12], i_9_, i_10_, i_7_, i_13_, i_12_, i_1_, i_2_}, x1344x);
	defparam lut_1504.LUT_SIZE = 8;
	defparam lut_1504.mask = 256'h5555ffff5555ffff5555ffffffffffff00002000000000000000000000000000;

	lut_sub lut_1506 ({sk[13], i_9_, i_7_, i_8_, i_6_, i_3_, i_2_}, x45x);
	defparam lut_1506.LUT_SIZE = 7;
	defparam lut_1506.mask = 128'h0037ffff0037ffff000a0c0e00000000;

	lut_sub lut_1509 ({sk[14], i_9_, i_7_, i_8_, i_3_, i_13_, i_4_, i_12_, i_1_}, x1332x);
	defparam lut_1509.LUT_SIZE = 9;
	defparam lut_1509.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff0000000000000000000000004500050000000000000000000000000000000000;

	lut_sub lut_1512 ({sk[15], i_9_, i_7_, i_8_, i_3_, i_13_, i_12_, i_11_, i_2_}, x1333x);
	defparam lut_1512.LUT_SIZE = 9;
	defparam lut_1512.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff08000800080008000c0000000000000000000000000000000000000000000000;

	lut_sub lut_1515 ({sk[0], i_9_, i_8_, i_6_, i_13_, i_4_, i_11_}, x471x);
	defparam lut_1515.LUT_SIZE = 7;
	defparam lut_1515.mask = 128'h0037ffff0037ffff00b0003000000000;

	lut_sub lut_1518 ({sk[1], i_9_, i_8_, i_6_, i_3_, i_13_, i_12_, i_11_, i_2_}, x1328x);
	defparam lut_1518.LUT_SIZE = 9;
	defparam lut_1518.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff0000000008000000000000000000000000000000000000000000000000000000;

	lut_sub lut_1520 ({sk[2], i_13_, i_12_, i_11_, i_2_}, x301x);
	defparam lut_1520.LUT_SIZE = 5;
	defparam lut_1520.mask = 32'h333f2000;

	lut_sub lut_1522 ({sk[3], i_4_, i_1_, i_2_}, n_n346);
	defparam lut_1522.LUT_SIZE = 4;
	defparam lut_1522.mask = 16'h5710;

	lut_sub lut_1524 ({sk[4], i_9_, i_13_, i_11_}, n_n755);
	defparam lut_1524.LUT_SIZE = 4;
	defparam lut_1524.mask = 16'h5740;

	lut_sub lut_1526 ({sk[5], i_5_, i_3_, i_4_}, n_n846);
	defparam lut_1526.LUT_SIZE = 4;
	defparam lut_1526.mask = 16'h5701;

	lut_sub lut_1528 ({sk[6], i_9_, i_8_, i_5_, i_4_, i_1_, i_2_}, x406x);
	defparam lut_1528.LUT_SIZE = 7;
	defparam lut_1528.mask = 128'h0037ffff0037ffff0000000800000000;

	lut_sub lut_1530 ({sk[7], i_9_, i_8_, i_5_, i_6_, i_4_, i_1_, i_2_, i_0_}, x478x);
	defparam lut_1530.LUT_SIZE = 9;
	defparam lut_1530.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff00000000000000000080008800c000c800000000000000000000000000000000;

	lut_sub lut_1534 ({sk[8], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_, n_n752, n_n756}, x477x);
	defparam lut_1534.LUT_SIZE = 9;
	defparam lut_1534.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff0000000000000000000000000050003000000000000000000000000000050000;

	lut_sub lut_1538 ({sk[9], i_9_, i_13_, i_1_, i_2_, i_0_}, x6740x);
	defparam lut_1538.LUT_SIZE = 6;
	defparam lut_1538.mask = 64'h115511ff01000000;

	lut_sub lut_1540 ({sk[10], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x6741x);
	defparam lut_1540.LUT_SIZE = 7;
	defparam lut_1540.mask = 128'h0037ffff0037ffff0000000000000001;

	lut_sub lut_1542 ({sk[11], i_13_, i_4_, i_12_, i_11_, i_2_}, x6742x);
	defparam lut_1542.LUT_SIZE = 6;
	defparam lut_1542.mask = 64'h115511ff00020000;

	lut_sub lut_1544 ({sk[12], i_9_, i_7_, i_8_, i_1_, i_0_}, x6743x);
	defparam lut_1544.LUT_SIZE = 6;
	defparam lut_1544.mask = 64'h115511ff00010000;

	lut_sub lut_1546 ({sk[13], n_n853, x37x, x322x, x478x, x6740x, x6741x, x6742x, x6743x}, x6746x);
	defparam lut_1546.LUT_SIZE = 9;
	defparam lut_1546.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff000f000f333f333f555f555f777f777f000fffff333fffff555fffff777fffff;

	lut_sub lut_1551 ({sk[14], i_3_, i_13_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_}, x113x);
	defparam lut_1551.LUT_SIZE = 9;
	defparam lut_1551.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff0000000000000800000000000000000000000000000000000000000000000000;

	lut_sub lut_1553 ({sk[15], i_10_, i_6_, i_3_, i_2_, i_0_}, x399x);
	defparam lut_1553.LUT_SIZE = 6;
	defparam lut_1553.mask = 64'h115511ff80000000;

	lut_sub lut_1555 ({sk[0], i_9_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_}, x6674x);
	defparam lut_1555.LUT_SIZE = 9;
	defparam lut_1555.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff000000000088000000c0000000c8000000000000000000000000000000000000;

	lut_sub lut_1558 ({sk[1], i_5_, i_6_, i_3_, i_2_, i_0_}, x480x);
	defparam lut_1558.LUT_SIZE = 6;
	defparam lut_1558.mask = 64'h115511ffc0008000;

	lut_sub lut_1561 ({sk[2], i_10_, i_13_, i_12_, i_11_}, x6670x);
	defparam lut_1561.LUT_SIZE = 5;
	defparam lut_1561.mask = 32'h333f0008;

	lut_sub lut_1563 ({sk[3], i_6_, i_3_, i_2_, i_0_}, x6672x);
	defparam lut_1563.LUT_SIZE = 5;
	defparam lut_1563.mask = 32'h333f4000;

	lut_sub lut_1565 ({sk[4], i_9_, i_13_, i_12_}, n_n550);
	defparam lut_1565.LUT_SIZE = 4;
	defparam lut_1565.mask = 16'h5780;

	lut_sub lut_1567 ({sk[5], i_9_, i_10_, i_6_, i_13_, i_12_, i_1_, i_11_}, n_n1126);
	defparam lut_1567.LUT_SIZE = 8;
	defparam lut_1567.mask = 256'h5555ffff5555ffff5555ffffffffffff008800c000bb00c0008800f300bb00f3;

	lut_sub lut_1577 ({sk[6], i_4_, i_1_}, x22x);
	defparam lut_1577.LUT_SIZE = 3;
	defparam lut_1577.mask = 8'h14;

	lut_sub lut_1579 ({sk[7], i_9_, i_10_, i_7_, i_8_, i_6_, i_4_, i_1_, i_11_}, x1294x);
	defparam lut_1579.LUT_SIZE = 9;
	defparam lut_1579.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff0000000000000000100000000000000000100000000000001010000000000000;

	lut_sub lut_1583 ({sk[8], i_9_, i_10_, i_7_, i_8_, i_6_, i_12_, i_11_}, x6887x);
	defparam lut_1583.LUT_SIZE = 8;
	defparam lut_1583.mask = 256'h5555ffff5555ffff5555ffffffffffff00000000000000000005000000050030;

	lut_sub lut_1586 ({sk[9], i_9_, i_10_, i_7_, i_8_, i_6_, i_12_, i_11_}, x491x);
	defparam lut_1586.LUT_SIZE = 8;
	defparam lut_1586.mask = 256'h5555ffff5555ffff5555ffffffffffff00000000000000000004000000042020;

	lut_sub lut_1589 ({sk[10], i_9_, i_8_, i_6_, i_4_, i_12_, i_1_, i_11_, i_2_}, x1293x);
	defparam lut_1589.LUT_SIZE = 9;
	defparam lut_1589.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff0000000010000000000000000000000000000000110000000000000000000000;

	lut_sub lut_1592 ({sk[11], i_9_, i_7_, i_8_, i_6_, i_4_, i_12_, i_1_, i_11_}, x1295x);
	defparam lut_1592.LUT_SIZE = 9;
	defparam lut_1592.mask = 512'h000000ff000000ffffffffffffffffffffffffffffffffffffffffffffffffff0000400000000000000000000000000000005000000000000000000000000000;

	lut_sub lut_1595 ({sk[12], i_9_, i_10_, i_8_, i_6_, i_4_, i_1_, i_11_, i_2_}, x1296x);
	defparam lut_1595.LUT_SIZE = 9;
	defparam lut_1595.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000010000000000000000000100000000000100010000000000;

	lut_sub lut_1598 ({sk[13], i_10_, i_7_, i_6_, i_12_, i_1_, i_11_, i_2_}, x6889x);
	defparam lut_1598.LUT_SIZE = 8;
	defparam lut_1598.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000000004545500000000000;

	lut_sub lut_1603 ({sk[14], i_9_, i_8_, i_4_}, x318x);
	defparam lut_1603.LUT_SIZE = 4;
	defparam lut_1603.mask = 16'h0f10;

	lut_sub lut_1605 ({sk[15], i_10_, i_5_, i_13_, i_4_, i_12_, i_1_, i_11_}, x1493x);
	defparam lut_1605.LUT_SIZE = 8;
	defparam lut_1605.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000700000000000000040000;

	lut_sub lut_1608 ({sk[0], i_9_, i_8_, i_5_, i_6_, i_1_, i_2_, i_0_}, x494x);
	defparam lut_1608.LUT_SIZE = 8;
	defparam lut_1608.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000001103130000000000000000;

	lut_sub lut_1611 ({sk[1], i_10_, i_13_, i_12_, i_1_, i_2_, i_0_}, x6747x);
	defparam lut_1611.LUT_SIZE = 7;
	defparam lut_1611.mask = 128'h0f0fffffffffffff0001000000000000;

	lut_sub lut_1613 ({sk[2], i_5_, i_6_, i_13_, i_4_, i_12_, i_1_, i_11_, i_0_}, x6749x);
	defparam lut_1613.LUT_SIZE = 9;
	defparam lut_1613.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff000000200000000000000020000000000000002000000000000000ff00000000;

	lut_sub lut_1616 ({sk[3], i_10_, i_6_, i_13_, i_4_, i_12_, i_11_, i_0_}, x6750x);
	defparam lut_1616.LUT_SIZE = 8;
	defparam lut_1616.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000700000000000000020000;

	lut_sub lut_1619 ({sk[4], n_n764, x37x, x318x, x1493x, x494x, x6747x, x6749x, x6750x}, n_n1259);
	defparam lut_1619.LUT_SIZE = 9;
	defparam lut_1619.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff000000000f0f0f0f00ff00ff0fff0fff7777ffff7f7fffff77ffffff7fffffff;

	lut_sub lut_1625 ({sk[5], i_9_, i_5_, i_6_, i_3_, i_13_, i_12_, i_2_, i_0_}, x1637x);
	defparam lut_1625.LUT_SIZE = 9;
	defparam lut_1625.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000008000000000000000c00000;

	lut_sub lut_1628 ({sk[6], i_9_, i_7_, i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x499x);
	defparam lut_1628.LUT_SIZE = 9;
	defparam lut_1628.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000c000c000a000aa00f000ff00;

	lut_sub lut_1634 ({sk[7], i_10_, i_5_, i_3_, i_13_, i_12_, i_1_, i_11_, i_2_}, x1634x);
	defparam lut_1634.LUT_SIZE = 9;
	defparam lut_1634.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000008000000000000000000000000000;

	lut_sub lut_1636 ({sk[8], i_3_, i_4_, i_1_, i_2_}, x272x);
	defparam lut_1636.LUT_SIZE = 5;
	defparam lut_1636.mask = 32'h5fff0010;

	lut_sub lut_1638 ({sk[9], i_9_, i_10_, i_6_, i_12_, i_11_}, x504x);
	defparam lut_1638.LUT_SIZE = 6;
	defparam lut_1638.mask = 64'h77ff77ff00100011;

	lut_sub lut_1641 ({sk[10], i_9_, i_6_, i_3_, i_4_, i_12_, i_1_, i_11_, i_2_}, x1268x);
	defparam lut_1641.LUT_SIZE = 9;
	defparam lut_1641.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000005000000000000000000000000003000055070000;

	lut_sub lut_1646 ({sk[11], i_10_, i_6_, i_3_, i_4_, i_1_, i_11_, i_2_}, x6894x);
	defparam lut_1646.LUT_SIZE = 8;
	defparam lut_1646.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000000000000450000000000;

	lut_sub lut_1649 ({sk[12], i_9_, i_8_, i_12_}, x270x);
	defparam lut_1649.LUT_SIZE = 4;
	defparam lut_1649.mask = 16'h0f01;

	lut_sub lut_1651 ({sk[13], i_10_, i_7_, i_8_, i_3_, i_12_, i_1_, i_11_, i_2_}, x508x);
	defparam lut_1651.LUT_SIZE = 9;
	defparam lut_1651.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000004547000000000000454f00000000;

	lut_sub lut_1656 ({sk[14], i_10_, i_8_, i_6_, i_3_, i_12_, i_1_, i_11_, i_2_}, x1256x);
	defparam lut_1656.LUT_SIZE = 9;
	defparam lut_1656.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000004000000050000000000000000000;

	lut_sub lut_1659 ({sk[15], i_9_, i_10_, i_8_, i_6_, i_3_, i_12_, i_1_, i_11_}, x6904x);
	defparam lut_1659.LUT_SIZE = 9;
	defparam lut_1659.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000010001000100010001;

	lut_sub lut_1662 ({sk[0], i_9_, i_10_, i_7_, i_6_, i_3_, i_12_, i_1_, i_11_}, x1246x);
	defparam lut_1662.LUT_SIZE = 9;
	defparam lut_1662.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000011005100000000;

	lut_sub lut_1665 ({sk[1], i_9_, i_7_, i_8_, i_6_, i_3_, i_12_, i_1_, i_11_}, x1247x);
	defparam lut_1665.LUT_SIZE = 9;
	defparam lut_1665.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000080003;

	lut_sub lut_1668 ({sk[2], i_9_, i_8_, i_6_, i_3_, i_12_, i_1_, i_11_, i_2_}, x6909x);
	defparam lut_1668.LUT_SIZE = 9;
	defparam lut_1668.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000404000005505;

	lut_sub lut_1673 ({sk[3], i_10_, i_7_, i_8_, i_6_, i_3_, i_12_, i_1_, i_11_}, x7976x);
	defparam lut_1673.LUT_SIZE = 9;
	defparam lut_1673.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeefffffffffffffff5ffffffffffff;

	lut_sub lut_1685 ({sk[4], i_9_, i_10_, i_7_, i_6_, i_12_, i_1_, i_11_, i_2_}, x7989x);
	defparam lut_1685.LUT_SIZE = 9;
	defparam lut_1685.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000404055054545550545455505;

	lut_sub lut_1700 ({sk[5], i_5_, i_3_, i_4_}, n_n710);
	defparam lut_1700.LUT_SIZE = 4;
	defparam lut_1700.mask = 16'h0f40;

	lut_sub lut_1702 ({sk[6], i_5_, i_3_, i_13_, i_4_, i_12_, i_11_}, x6650x);
	defparam lut_1702.LUT_SIZE = 7;
	defparam lut_1702.mask = 128'h0f0fffffffffffff0000000020000000;

	lut_sub lut_1704 ({sk[7], i_7_, i_8_, i_6_, i_3_, i_4_, i_1_}, x518x);
	defparam lut_1704.LUT_SIZE = 7;
	defparam lut_1704.mask = 128'h0f0fffffffffffff0000000040c00000;

	lut_sub lut_1707 ({sk[8], i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x517x);
	defparam lut_1707.LUT_SIZE = 8;
	defparam lut_1707.mask = 256'h0fffffff0fffffff0fffffff0fffffff80800000000000008000000000000000;

	lut_sub lut_1710 ({sk[9], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x520x);
	defparam lut_1710.LUT_SIZE = 7;
	defparam lut_1710.mask = 128'h0f0fffffffffffff0220000000000000;

	lut_sub lut_1713 ({sk[10], i_9_, i_10_, i_7_, i_8_, i_13_, i_12_, i_1_, i_11_}, x1629x);
	defparam lut_1713.LUT_SIZE = 9;
	defparam lut_1713.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000002000000000000000000000000000000000000000000000000000000;

	lut_sub lut_1715 ({sk[11], i_9_, i_13_, i_1_, i_11_, i_2_, i_0_}, x6648x);
	defparam lut_1715.LUT_SIZE = 7;
	defparam lut_1715.mask = 128'h0f0fffffffffffff0010000000000000;

	lut_sub lut_1717 ({sk[12], i_10_, i_13_, i_1_, i_11_, i_2_, i_0_}, x6643x);
	defparam lut_1717.LUT_SIZE = 7;
	defparam lut_1717.mask = 128'h0f0fffffffffffff0010000000000000;

	lut_sub lut_1719 ({sk[13], i_9_, i_10_, i_8_, i_3_, i_11_}, x392x);
	defparam lut_1719.LUT_SIZE = 6;
	defparam lut_1719.mask = 64'h77ff77ff80000000;

	lut_sub lut_1721 ({sk[14], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_, n_n748, n_n746}, x523x);
	defparam lut_1721.LUT_SIZE = 9;
	defparam lut_1721.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000005000300000000000000000000000000005000300;

	lut_sub lut_1726 ({sk[15], i_8_, i_5_, i_6_, i_3_, i_0_}, x522x);
	defparam lut_1726.LUT_SIZE = 6;
	defparam lut_1726.mask = 64'h77ff77ff040c0000;

	lut_sub lut_1729 ({sk[0], i_5_, i_13_, i_4_, i_12_, i_1_, i_2_, i_0_}, x521x);
	defparam lut_1729.LUT_SIZE = 8;
	defparam lut_1729.mask = 256'h0fffffff0fffffff0fffffff0fffffff01010000000000000103000000000000;

	lut_sub lut_1732 ({sk[1], i_4_, i_2_, x303x, x392x, x522x, x521x, x6753x, x6754x}, x6758x);
	defparam lut_1732.LUT_SIZE = 9;
	defparam lut_1732.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff11111f1f11111f1f11111f1f11ff1fff11111f1f11111f1f11111f1f11111f1f;

	lut_sub lut_1736 ({sk[2], i_7_, i_2_}, x275x);
	defparam lut_1736.LUT_SIZE = 3;
	defparam lut_1736.mask = 8'h58;

	lut_sub lut_1738 ({sk[3], i_10_, i_7_, i_8_}, n_n651);
	defparam lut_1738.LUT_SIZE = 4;
	defparam lut_1738.mask = 16'h0f01;

	lut_sub lut_1740 ({sk[4], i_9_, i_5_, i_3_, i_13_, i_4_, i_11_}, x6654x);
	defparam lut_1740.LUT_SIZE = 7;
	defparam lut_1740.mask = 128'h0f0fffffffffffff0000100000000000;

	lut_sub lut_1742 ({sk[5], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x541x);
	defparam lut_1742.LUT_SIZE = 7;
	defparam lut_1742.mask = 128'h0f0fffffffffffff0400000008000000;

	lut_sub lut_1745 ({sk[6], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x6655x);
	defparam lut_1745.LUT_SIZE = 7;
	defparam lut_1745.mask = 128'h0f0fffffffffffff4000000000000000;

	lut_sub lut_1747 ({sk[7], i_9_, i_13_, i_1_, i_11_, i_2_, i_0_}, x6656x);
	defparam lut_1747.LUT_SIZE = 7;
	defparam lut_1747.mask = 128'h0f0fffffffffffff0002000000000000;

	lut_sub lut_1749 ({sk[8], i_9_, i_13_, i_1_, i_11_, i_2_, i_0_}, x6657x);
	defparam lut_1749.LUT_SIZE = 7;
	defparam lut_1749.mask = 128'h0f0fffffffffffff0200000000000000;

	lut_sub lut_1751 ({sk[9], i_5_, i_3_, i_13_, i_4_, i_1_, i_11_, i_2_, i_0_}, x405x);
	defparam lut_1751.LUT_SIZE = 9;
	defparam lut_1751.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000080000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_1753 ({sk[10], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x544x);
	defparam lut_1753.LUT_SIZE = 7;
	defparam lut_1753.mask = 128'h0f0fffffffffffff0008000000040000;

	lut_sub lut_1756 ({sk[11], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x543x);
	defparam lut_1756.LUT_SIZE = 7;
	defparam lut_1756.mask = 128'h0f0fffffffffffff0010000000200000;

	lut_sub lut_1759 ({sk[12], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x573x);
	defparam lut_1759.LUT_SIZE = 7;
	defparam lut_1759.mask = 128'h0f0fffffffffffff0000020000000800;

	lut_sub lut_1762 ({sk[13], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x572x);
	defparam lut_1762.LUT_SIZE = 7;
	defparam lut_1762.mask = 128'h0f0fffffffffffff0000000000000440;

	lut_sub lut_1765 ({sk[14], i_10_, i_7_, i_3_, i_1_, i_0_}, x6679x);
	defparam lut_1765.LUT_SIZE = 6;
	defparam lut_1765.mask = 64'h77ff77ff80000000;

	lut_sub lut_1767 ({sk[15], i_5_, i_3_, i_13_, i_4_, i_12_, i_1_, i_2_, i_0_}, x121x);
	defparam lut_1767.LUT_SIZE = 9;
	defparam lut_1767.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000080000000000000000000000000;

	lut_sub lut_1769 ({sk[0], i_7_, i_5_, i_3_, i_4_, i_1_}, x404x);
	defparam lut_1769.LUT_SIZE = 6;
	defparam lut_1769.mask = 64'h77ff77ff20000000;

	lut_sub lut_1771 ({sk[1], i_7_, i_6_, i_3_, i_1_, i_0_}, x570x);
	defparam lut_1771.LUT_SIZE = 6;
	defparam lut_1771.mask = 64'h77ff77ff50400000;

	lut_sub lut_1774 ({sk[2], i_10_, i_7_, i_6_, i_13_, i_12_, i_11_}, x6684x);
	defparam lut_1774.LUT_SIZE = 7;
	defparam lut_1774.mask = 128'h0f0fffffffffffff1000000000000000;

	lut_sub lut_1776 ({sk[3], i_9_, i_7_, i_5_, i_6_, i_3_, i_4_, i_1_, i_0_}, x6689x);
	defparam lut_1776.LUT_SIZE = 9;
	defparam lut_1776.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff000000000000000000000a000c000f0000000000000000000000000000000000;

	lut_sub lut_1780 ({sk[4], i_10_, i_7_, i_8_, i_4_, i_12_, i_1_, i_11_, i_2_}, x554x);
	defparam lut_1780.LUT_SIZE = 9;
	defparam lut_1780.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff00000000004000000000000000400000000000000045000000000000004f0000;

	lut_sub lut_1785 ({sk[5], i_9_, i_10_, i_7_, i_8_, i_6_, i_4_, i_12_, i_1_}, x1219x);
	defparam lut_1785.LUT_SIZE = 9;
	defparam lut_1785.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000100000000000001010;

	lut_sub lut_1788 ({sk[6], i_10_, i_7_, i_8_, i_6_, i_4_, i_12_, i_1_, i_11_}, x1220x);
	defparam lut_1788.LUT_SIZE = 9;
	defparam lut_1788.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff000000000000000000000000080000000000000000000000000000000a000000;

	lut_sub lut_1791 ({sk[7], i_7_, i_5_, i_6_, i_12_, i_1_, i_11_, i_2_, i_0_}, x557x);
	defparam lut_1791.LUT_SIZE = 9;
	defparam lut_1791.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0011001100110011020200000000000000000000000000000000000000000000;

	lut_sub lut_1794 ({sk[8], i_9_, i_10_, i_5_, i_12_, i_11_}, x46x);
	defparam lut_1794.LUT_SIZE = 6;
	defparam lut_1794.mask = 64'h77ff77ff000000a8;

	lut_sub lut_1797 ({sk[9], i_5_, i_12_}, x276x);
	defparam lut_1797.LUT_SIZE = 3;
	defparam lut_1797.mask = 8'h52;

	lut_sub lut_1799 ({sk[10], i_9_, i_10_, i_3_, i_12_, i_11_, i_2_, i_0_}, x190x);
	defparam lut_1799.LUT_SIZE = 8;
	defparam lut_1799.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000000000000000000010005;

	lut_sub lut_1802 ({sk[11], i_10_, i_7_, i_5_, i_6_, i_12_, i_11_, i_2_, i_0_}, x7251x);
	defparam lut_1802.LUT_SIZE = 9;
	defparam lut_1802.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000001010001000000000000000000000000;

	lut_sub lut_1805 ({sk[12], i_10_, i_7_, i_5_, i_6_, i_1_, i_11_, i_2_, i_0_}, x560x);
	defparam lut_1805.LUT_SIZE = 9;
	defparam lut_1805.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000a0002000aa002200a0000000aa0000;

	lut_sub lut_1810 ({sk[13], i_5_, i_6_, i_12_, i_1_, i_2_}, x559x);
	defparam lut_1810.LUT_SIZE = 6;
	defparam lut_1810.mask = 64'h77ff77ff11150000;

	lut_sub lut_1813 ({sk[14], i_10_, i_7_, i_5_, i_6_, i_12_, i_2_, i_0_}, x174x);
	defparam lut_1813.LUT_SIZE = 8;
	defparam lut_1813.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000000000001000000000000;

	lut_sub lut_1815 ({sk[15], i_10_, i_5_, i_6_, i_1_, i_11_, i_0_}, x175x);
	defparam lut_1815.LUT_SIZE = 7;
	defparam lut_1815.mask = 128'h0f0fffffffffffff000000000d000000;

	lut_sub lut_1818 ({sk[0], i_5_, i_6_, i_12_, i_11_, i_0_}, x565x);
	defparam lut_1818.LUT_SIZE = 6;
	defparam lut_1818.mask = 64'h77ff77ff008800f5;

	lut_sub lut_1823 ({sk[1], i_5_, i_6_, i_12_, i_2_, i_0_}, x563x);
	defparam lut_1823.LUT_SIZE = 6;
	defparam lut_1823.mask = 64'h77ff77ff11003100;

	lut_sub lut_1826 ({sk[2], i_9_, i_10_, i_5_, i_6_, i_12_, i_11_, i_2_, i_0_}, x161x);
	defparam lut_1826.LUT_SIZE = 9;
	defparam lut_1826.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000003100000011;

	lut_sub lut_1829 ({sk[3], i_5_, i_3_, i_4_}, n_n851);
	defparam lut_1829.LUT_SIZE = 4;
	defparam lut_1829.mask = 16'h0f10;

	lut_sub lut_1831 ({sk[4], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x610x);
	defparam lut_1831.LUT_SIZE = 7;
	defparam lut_1831.mask = 128'h0f0fffffffffffff0220000008800000;

	lut_sub lut_1836 ({sk[5], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x609x);
	defparam lut_1836.LUT_SIZE = 7;
	defparam lut_1836.mask = 128'h0f0fffffffffffff0010000004400000;

	lut_sub lut_1840 ({sk[6], i_10_, i_13_, i_1_, i_2_, i_0_}, x6768x);
	defparam lut_1840.LUT_SIZE = 6;
	defparam lut_1840.mask = 64'h77ff77ff01000000;

	lut_sub lut_1842 ({sk[7], n_n2368, n_n849, n_n843, n_n846, n_n851, x610x, x609x, x6768x}, n_n1265);
	defparam lut_1842.LUT_SIZE = 9;
	defparam lut_1842.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff000000000055005500330f3f00770f7fffffffffffffffffffffffffffffffff;

	lut_sub lut_1847 ({sk[8], i_10_, i_13_, i_11_, x327x, x9x, x37x, x606x, x384x}, x6766x);
	defparam lut_1847.LUT_SIZE = 9;
	defparam lut_1847.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff03030303035703ff030303030303030303030303030303030303030303030303;

	lut_sub lut_1851 ({sk[9], x313x, x9x, n_n849, x266x, x6764x, x287x, x6762x, x6763x}, x6767x);
	defparam lut_1851.LUT_SIZE = 9;
	defparam lut_1851.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000555500ff55ff000055550fff5fff0000555500ff55ff333377773fff7fff;

	lut_sub lut_1856 ({sk[10], i_9_, i_5_, i_3_, i_13_, i_4_, i_0_, n_n816, n_n822}, x611x);
	defparam lut_1856.LUT_SIZE = 9;
	defparam lut_1856.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000330033000000000057000300000000000000000000000000000000;

	lut_sub lut_1860 ({sk[11], i_7_, i_6_, i_3_, i_1_, i_2_, x313x, x9x, x402x}, x6779x);
	defparam lut_1860.LUT_SIZE = 9;
	defparam lut_1860.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000555500005555000055550003555700000000000000000000000000030003;

	lut_sub lut_1863 ({sk[12], i_10_, i_13_, i_12_, i_11_, x9x, x292x, x359x, x612x}, x6780x);
	defparam lut_1863.LUT_SIZE = 9;
	defparam lut_1863.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff000f003f555f557f000000000000000000000000000000000000000000000000;

	lut_sub lut_1867 ({sk[13], i_9_, i_5_, i_3_, i_4_, i_1_, i_0_}, x574x);
	defparam lut_1867.LUT_SIZE = 7;
	defparam lut_1867.mask = 128'h0f0fffffffffffff0003000100000000;

	lut_sub lut_1870 ({sk[14], i_5_, i_3_, i_4_, i_12_, i_1_, i_2_, i_0_}, x584x);
	defparam lut_1870.LUT_SIZE = 8;
	defparam lut_1870.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000010100000000000002000000;

	lut_sub lut_1873 ({sk[15], i_9_, i_7_, i_8_, i_6_, i_2_}, x6800x);
	defparam lut_1873.LUT_SIZE = 6;
	defparam lut_1873.mask = 64'h77ff77ff20000000;

	lut_sub lut_1875 ({sk[0], i_9_, i_7_, i_8_, i_6_, i_13_, i_12_}, x6802x);
	defparam lut_1875.LUT_SIZE = 7;
	defparam lut_1875.mask = 128'h0f0fffffffffffff0000080000000000;

	lut_sub lut_1877 ({sk[1], i_11_, n_n761, n_n833, n_n538, n_n843, x584x, x6800x, x6802x}, x583x);
	defparam lut_1877.LUT_SIZE = 9;
	defparam lut_1877.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff000f000f000f555f000f333f000f777f000f000f000f555f000f000f000f555f;

	lut_sub lut_1881 ({sk[2], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x6796x);
	defparam lut_1881.LUT_SIZE = 7;
	defparam lut_1881.mask = 128'h0f0fffffffffffff0000080000000000;

	lut_sub lut_1883 ({sk[3], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x6798x);
	defparam lut_1883.LUT_SIZE = 7;
	defparam lut_1883.mask = 128'h0f0fffffffffffff0000000000004000;

	lut_sub lut_1885 ({sk[4], i_7_, i_8_, i_6_, n_n835, n_n550, x302x, x6796x, x6798x}, x581x);
	defparam lut_1885.LUT_SIZE = 9;
	defparam lut_1885.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000550f5f003300330000000000000000;

	lut_sub lut_1889 ({sk[5], i_9_, i_10_, i_3_, i_4_, i_1_, i_2_, i_0_}, x115x);
	defparam lut_1889.LUT_SIZE = 8;
	defparam lut_1889.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000000000000000000000100;

	lut_sub lut_1891 ({sk[6], i_10_, i_7_, i_6_, i_13_, i_12_, i_11_}, x6808x);
	defparam lut_1891.LUT_SIZE = 7;
	defparam lut_1891.mask = 128'h0f0fffffffffffff0000000000200000;

	lut_sub lut_1893 ({sk[7], i_9_, i_10_, i_7_, i_6_, i_11_}, x6810x);
	defparam lut_1893.LUT_SIZE = 6;
	defparam lut_1893.mask = 64'h77ff77ff00000004;

	lut_sub lut_1895 ({sk[8], i_3_, i_1_, i_2_, i_0_}, x292x);
	defparam lut_1895.LUT_SIZE = 5;
	defparam lut_1895.mask = 32'h5fff0001;

	lut_sub lut_1897 ({sk[9], i_7_, i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x588x);
	defparam lut_1897.LUT_SIZE = 8;
	defparam lut_1897.mask = 256'h0fffffff0fffffff0fffffff0fffffff00ff000f005500050003000300000000;

	lut_sub lut_1903 ({sk[10], i_7_, i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x587x);
	defparam lut_1903.LUT_SIZE = 8;
	defparam lut_1903.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000300330005000500070037;

	lut_sub lut_1907 ({sk[11], i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_11_}, x586x);
	defparam lut_1907.LUT_SIZE = 8;
	defparam lut_1907.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000040000000200000000000;

	lut_sub lut_1910 ({sk[12], i_9_, i_7_, i_5_, i_6_}, x591x);
	defparam lut_1910.LUT_SIZE = 5;
	defparam lut_1910.mask = 32'h5fff0405;

	lut_sub lut_1913 ({sk[13], i_9_, i_10_, i_5_, i_12_, i_11_}, x590x);
	defparam lut_1913.LUT_SIZE = 6;
	defparam lut_1913.mask = 64'h77ff77ff00a00cac;

	lut_sub lut_1916 ({sk[14], i_10_, i_12_, i_11_, i_0_}, x7208x);
	defparam lut_1916.LUT_SIZE = 5;
	defparam lut_1916.mask = 32'h5fff080c;

	lut_sub lut_1919 ({sk[15], i_7_, i_5_, i_6_, i_3_, i_4_}, x7209x);
	defparam lut_1919.LUT_SIZE = 6;
	defparam lut_1919.mask = 64'h77ff77ff00000200;

	lut_sub lut_1921 ({sk[0], i_10_, i_3_, i_4_, i_12_, i_0_}, x7210x);
	defparam lut_1921.LUT_SIZE = 6;
	defparam lut_1921.mask = 64'h77ff77ff00000010;

	lut_sub lut_1923 ({sk[1], i_9_, i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x238x);
	defparam lut_1923.LUT_SIZE = 8;
	defparam lut_1923.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000000000000000000000100;

	lut_sub lut_1925 ({sk[2], i_5_, i_3_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_}, x7211x);
	defparam lut_1925.LUT_SIZE = 9;
	defparam lut_1925.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000002000000000000000000000000000000022000000000000;

	lut_sub lut_1928 ({sk[3], i_9_, i_10_, i_7_, i_8_, i_2_}, x597x);
	defparam lut_1928.LUT_SIZE = 6;
	defparam lut_1928.mask = 64'h77ff77ff0044004f;

	lut_sub lut_1931 ({sk[4], i_10_, i_5_, i_6_, i_3_, i_12_, i_11_, i_2_, i_0_}, x596x);
	defparam lut_1931.LUT_SIZE = 9;
	defparam lut_1931.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000005000000150000000000000000;

	lut_sub lut_1934 ({sk[5], i_10_, i_8_, i_5_, i_3_, i_12_, i_1_, i_2_, i_0_}, x127x);
	defparam lut_1934.LUT_SIZE = 9;
	defparam lut_1934.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000002000000000000000000;

	lut_sub lut_1936 ({sk[6], i_10_, i_7_, i_8_, i_5_, i_3_, i_1_, i_11_, i_0_}, x128x);
	defparam lut_1936.LUT_SIZE = 9;
	defparam lut_1936.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000010000000000000000000000000000;

	lut_sub lut_1938 ({sk[7], i_5_, i_6_, i_3_, i_12_, i_11_}, x7284x);
	defparam lut_1938.LUT_SIZE = 6;
	defparam lut_1938.mask = 64'h77ff77ff00020000;

	lut_sub lut_1940 ({sk[8], i_9_, i_10_, i_7_, i_5_, i_6_, i_3_, i_12_, i_11_}, x130x);
	defparam lut_1940.LUT_SIZE = 9;
	defparam lut_1940.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000040000000000;

	lut_sub lut_1942 ({sk[9], i_9_, i_10_, i_7_, i_6_, i_3_, i_12_, i_11_, i_0_}, x7289x);
	defparam lut_1942.LUT_SIZE = 9;
	defparam lut_1942.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000011000000000005;

	lut_sub lut_1945 ({sk[10], i_9_, i_7_, i_11_}, n_n277);
	defparam lut_1945.LUT_SIZE = 4;
	defparam lut_1945.mask = 16'h0f80;

	lut_sub lut_1947 ({sk[11], i_9_, i_8_, i_3_, i_4_, i_2_}, x600x);
	defparam lut_1947.LUT_SIZE = 6;
	defparam lut_1947.mask = 64'h77ff77ff20222020;

	lut_sub lut_1950 ({sk[12], i_9_, i_10_, i_7_, i_6_, i_12_, i_11_}, x604x);
	defparam lut_1950.LUT_SIZE = 7;
	defparam lut_1950.mask = 128'h0f0fffffffffffff0000503005035533;

	lut_sub lut_1955 ({sk[13], i_9_, i_10_, i_7_, i_6_, i_12_, i_1_, i_11_}, x603x);
	defparam lut_1955.LUT_SIZE = 8;
	defparam lut_1955.mask = 256'h0fffffff0fffffff0fffffff0fffffff0040080000400a000050080000500a00;

	lut_sub lut_1960 ({sk[14], i_9_, i_7_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_}, x6764x);
	defparam lut_1960.LUT_SIZE = 9;
	defparam lut_1960.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000010001000000000001000f00000000000000000000000000000000;

	lut_sub lut_1963 ({sk[15], i_9_, i_7_, i_5_, i_6_, i_3_, i_1_, i_0_}, x606x);
	defparam lut_1963.LUT_SIZE = 8;
	defparam lut_1963.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000503070000000000000000;

	lut_sub lut_1966 ({sk[0], i_7_, i_3_, i_1_, i_0_}, x287x);
	defparam lut_1966.LUT_SIZE = 5;
	defparam lut_1966.mask = 32'h5fff0001;

	lut_sub lut_1968 ({sk[1], i_7_, i_6_, i_3_}, x6762x);
	defparam lut_1968.LUT_SIZE = 4;
	defparam lut_1968.mask = 16'h0f01;

	lut_sub lut_1970 ({sk[2], i_5_, i_6_, i_3_, i_2_}, x6763x);
	defparam lut_1970.LUT_SIZE = 5;
	defparam lut_1970.mask = 32'h5fff0010;

	lut_sub lut_1972 ({sk[3], i_5_, i_3_, i_1_, i_2_}, x359x);
	defparam lut_1972.LUT_SIZE = 5;
	defparam lut_1972.mask = 32'h5fff0100;

	lut_sub lut_1974 ({sk[4], i_9_, i_10_, i_5_, i_3_, i_13_, i_4_, i_12_, i_11_}, x402x);
	defparam lut_1974.LUT_SIZE = 9;
	defparam lut_1974.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000100000000000000000000000000000000000000000000000000;

	lut_sub lut_1976 ({sk[5], i_9_, i_5_, i_6_, i_3_, i_4_, i_2_, i_0_}, x612x);
	defparam lut_1976.LUT_SIZE = 8;
	defparam lut_1976.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000001000000030000000000000000;

	lut_sub lut_1979 ({sk[6], i_9_, i_10_, i_8_, i_4_, i_12_, i_2_}, x355x);
	defparam lut_1979.LUT_SIZE = 7;
	defparam lut_1979.mask = 128'h0f0fffffffffffff0000000000000010;

	lut_sub lut_1981 ({sk[7], i_9_, i_8_, i_5_, i_3_, i_13_, i_4_, i_12_, i_11_}, x875x);
	defparam lut_1981.LUT_SIZE = 9;
	defparam lut_1981.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff00000000aa00000000000000cf000f0000000000000000000000000000000000;

	lut_sub lut_1985 ({sk[8], i_9_, i_7_, i_5_, i_3_, i_13_, i_4_, i_12_}, x7129x);
	defparam lut_1985.LUT_SIZE = 8;
	defparam lut_1985.mask = 256'h0fffffff0fffffff0fffffff0fffffff000030000000b0a00000000000000000;

	lut_sub lut_1988 ({sk[9], i_9_, i_7_, i_3_, i_13_, i_4_, i_11_, i_0_}, x873x);
	defparam lut_1988.LUT_SIZE = 8;
	defparam lut_1988.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000020000000000000000000000;

	lut_sub lut_1990 ({sk[10], i_13_, i_12_, i_1_, i_11_, i_0_}, x874x);
	defparam lut_1990.LUT_SIZE = 6;
	defparam lut_1990.mask = 64'h77ff77ff20000000;

	lut_sub lut_1992 ({sk[11], i_7_, i_8_, i_5_, i_6_, i_3_, i_1_, i_0_}, x637x);
	defparam lut_1992.LUT_SIZE = 8;
	defparam lut_1992.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000000000000000080a00000;

	lut_sub lut_1995 ({sk[12], i_6_, i_3_, i_1_, i_0_}, x41x);
	defparam lut_1995.LUT_SIZE = 5;
	defparam lut_1995.mask = 32'h5fffa080;

	lut_sub lut_1998 ({sk[13], i_9_, i_10_, i_8_, i_6_, i_3_, i_2_, i_0_}, x1081x);
	defparam lut_1998.LUT_SIZE = 8;
	defparam lut_1998.mask = 256'h0fffffff0fffffff0fffffff0fffffff80800000008000008000000000000000;

	lut_sub lut_2001 ({sk[14], i_7_, i_8_, i_6_, i_3_, i_1_, i_2_, i_0_}, x7009x);
	defparam lut_2001.LUT_SIZE = 8;
	defparam lut_2001.mask = 256'h0fffffff0fffffff0fffffff0fffffffa0a08080a0a08080a0a08000a0a00000;

	lut_sub lut_2005 ({sk[15], i_9_, i_10_, i_7_, i_6_, i_11_, i_2_, i_0_}, x1075x);
	defparam lut_2005.LUT_SIZE = 8;
	defparam lut_2005.mask = 256'h0fffffff0fffffff0fffffff0fffffff80800000008000008000000000000000;

	lut_sub lut_2008 ({sk[0], i_9_, i_10_, i_8_, i_5_, i_6_, i_3_, i_1_, i_2_}, x7017x);
	defparam lut_2008.LUT_SIZE = 9;
	defparam lut_2008.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffffcc008080cc0000000000808000000000cc000000cc0000000000000000000000;

	lut_sub lut_2011 ({sk[1], i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_1_, i_0_}, x7018x);
	defparam lut_2011.LUT_SIZE = 9;
	defparam lut_2011.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000cc000000cc0080a0cce00000cc0000000000000000000000000000000000;

	lut_sub lut_2016 ({sk[2], i_9_, i_10_, i_7_, i_5_, i_1_, i_11_, i_2_}, x7019x);
	defparam lut_2016.LUT_SIZE = 8;
	defparam lut_2016.mask = 256'h0fffffff0fffffff0fffffff0fffffff80800000008000008000000000000000;

	lut_sub lut_2019 ({sk[3], i_9_, i_10_, i_7_, i_8_, i_3_, i_1_, i_11_, i_2_}, x648x);
	defparam lut_2019.LUT_SIZE = 9;
	defparam lut_2019.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0101000101010001010100010101000101010001010101010303030303030303;

	lut_sub lut_2024 ({sk[4], i_9_, i_10_, i_5_, i_12_, i_1_, i_11_, i_2_, i_0_}, x657x);
	defparam lut_2024.LUT_SIZE = 9;
	defparam lut_2024.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000002000000000000000310000000000000020000000000000003100000011;

	lut_sub lut_2028 ({sk[5], i_10_, i_8_, i_5_, i_4_, i_12_, i_1_, i_11_, i_2_}, x772x);
	defparam lut_2028.LUT_SIZE = 9;
	defparam lut_2028.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000004000000000000;

	lut_sub lut_2030 ({sk[6], i_9_, i_8_, i_5_, i_4_, i_12_, i_1_, i_2_, i_0_}, x773x);
	defparam lut_2030.LUT_SIZE = 9;
	defparam lut_2030.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000010000;

	lut_sub lut_2032 ({sk[7], i_10_, i_7_, i_8_, i_5_, i_6_, i_12_, i_11_}, x776x);
	defparam lut_2032.LUT_SIZE = 8;
	defparam lut_2032.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000000000000000000000200;

	lut_sub lut_2034 ({sk[8], i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_12_, i_0_}, x7968x);
	defparam lut_2034.LUT_SIZE = 9;
	defparam lut_2034.mask = 512'h555555ffffffffffffffffffffffffff555555fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffffffffffffffefffffffffffffefe;

	lut_sub lut_2042 ({sk[9], i_7_, i_8_, i_5_, i_3_, i_4_, i_1_, i_2_}, x667x);
	defparam lut_2042.LUT_SIZE = 8;
	defparam lut_2042.mask = 256'h0fffffff0fffffff0fffffff0fffffff0c0800000c0000000808000000000000;

	lut_sub lut_2045 ({sk[10], i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_}, x666x);
	defparam lut_2045.LUT_SIZE = 9;
	defparam lut_2045.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff3222000030000000000000000000000000000000000000000000000000000000;

	lut_sub lut_2048 ({sk[11], i_10_, i_7_, i_8_, i_13_, i_12_, i_11_}, x7103x);
	defparam lut_2048.LUT_SIZE = 7;
	defparam lut_2048.mask = 128'h0f0fffffffffffff0040000000000000;

	lut_sub lut_2050 ({sk[12], i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_}, x7967x);
	defparam lut_2050.LUT_SIZE = 9;
	defparam lut_2050.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffffffffffffffffffffffffdfcfffffddcdffffffffffffffffffffffffffffffff;

	lut_sub lut_2058 ({sk[13], i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_1_}, x669x);
	defparam lut_2058.LUT_SIZE = 8;
	defparam lut_2058.mask = 256'h0fffffff0fffffff0fffffff0fffffff00a000a000ac00a00000000000000000;

	lut_sub lut_2062 ({sk[14], i_8_, i_5_, i_6_, i_3_}, x317x);
	defparam lut_2062.LUT_SIZE = 5;
	defparam lut_2062.mask = 32'h5fff0080;

	lut_sub lut_2064 ({sk[15], i_5_, i_6_, i_3_, i_4_, i_1_, i_2_}, x671x);
	defparam lut_2064.LUT_SIZE = 7;
	defparam lut_2064.mask = 128'h0f0fffffffffffff0a00080000000000;

	lut_sub lut_2067 ({sk[0], i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_2_, i_0_}, x676x);
	defparam lut_2067.LUT_SIZE = 9;
	defparam lut_2067.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffffff00aa0080008000800080008000800000000000000000000000000000000000;

	lut_sub lut_2071 ({sk[1], i_9_, i_10_, i_8_, i_6_, i_4_, i_2_, i_0_}, x7028x);
	defparam lut_2071.LUT_SIZE = 8;
	defparam lut_2071.mask = 256'h0fffffff0fffffff0fffffff0fffffff0f0f0f0f000000000800000000000000;

	lut_sub lut_2074 ({sk[2], i_10_, i_7_, i_5_, i_6_, i_3_, i_4_, i_2_}, x7029x);
	defparam lut_2074.LUT_SIZE = 8;
	defparam lut_2074.mask = 256'h0fffffff0fffffff0fffffff0fffffff30000000200000000000000000000000;

	lut_sub lut_2077 ({sk[3], i_9_, i_7_, i_3_, i_4_, i_1_, i_0_}, x108x);
	defparam lut_2077.LUT_SIZE = 7;
	defparam lut_2077.mask = 128'h0f0fffffffffffff0000080000000000;

	lut_sub lut_2079 ({sk[4], i_10_, i_7_, i_8_, i_3_, i_2_}, x679x);
	defparam lut_2079.LUT_SIZE = 6;
	defparam lut_2079.mask = 64'h77ff77ff0caa0000;

	lut_sub lut_2082 ({sk[5], i_9_, i_10_, i_7_, i_8_, i_3_, i_1_, i_0_}, x1041x);
	defparam lut_2082.LUT_SIZE = 8;
	defparam lut_2082.mask = 256'h0fffffff0fffffff0fffffff0fffffff00800080000000800080000000000000;

	lut_sub lut_2085 ({sk[6], i_9_, i_7_, i_6_, i_3_, i_4_, i_2_, i_0_}, x7021x);
	defparam lut_2085.LUT_SIZE = 8;
	defparam lut_2085.mask = 256'h0fffffff0fffffff0fffffff0fffffff0000080000000a000000000000000000;

	lut_sub lut_2088 ({sk[7], i_9_, i_7_, i_8_, i_5_, i_3_, i_4_, i_1_, i_0_}, x7038x);
	defparam lut_2088.LUT_SIZE = 9;
	defparam lut_2088.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff000000000000000008000c0008000c0c00000000000000000000000000000000;

	lut_sub lut_2092 ({sk[8], i_9_, i_7_, i_8_, i_6_, i_4_, i_1_, i_2_, i_0_}, x7970x);
	defparam lut_2092.LUT_SIZE = 9;
	defparam lut_2092.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffffffffffffff7fff77ffffffffff5fff57ffffffffffffffffffffffffffffffff;

	lut_sub lut_2100 ({sk[9], i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_2_}, x7987x);
	defparam lut_2100.LUT_SIZE = 9;
	defparam lut_2100.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000002000000022000000300000003200000000000000000000000000000000;

	lut_sub lut_2106 ({sk[10], i_9_, i_8_, i_5_, i_12_, i_1_, i_11_, i_2_, i_0_}, x411x);
	defparam lut_2106.LUT_SIZE = 9;
	defparam lut_2106.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000020002000200000;

	lut_sub lut_2109 ({sk[11], i_9_, i_10_, i_8_, i_5_, i_6_, i_12_}, x686x);
	defparam lut_2109.LUT_SIZE = 7;
	defparam lut_2109.mask = 128'h0f0fffffffffffff0000000000010011;

	lut_sub lut_2112 ({sk[12], i_8_, i_5_, i_6_, i_11_, i_0_}, x7189x);
	defparam lut_2112.LUT_SIZE = 6;
	defparam lut_2112.mask = 64'h77ff77ff00000800;

	lut_sub lut_2114 ({sk[13], i_9_, i_8_, i_5_, i_3_, i_12_, i_1_, i_2_, i_0_}, x368x);
	defparam lut_2114.LUT_SIZE = 9;
	defparam lut_2114.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000301;

	lut_sub lut_2117 ({sk[14], i_9_, i_10_, i_8_, i_5_, i_6_, i_3_, i_2_}, x7043x);
	defparam lut_2117.LUT_SIZE = 8;
	defparam lut_2117.mask = 256'h0fffffff0fffffff0fffffff0fffffff00008008000000080000800000000000;

	lut_sub lut_2120 ({sk[15], i_5_, i_6_, i_3_, i_4_, i_12_, i_1_, i_0_}, x690x);
	defparam lut_2120.LUT_SIZE = 8;
	defparam lut_2120.mask = 256'h0fffffff0fffffff0fffffff0fffffff0000000000aa00aac0c00000c0ff00ff;

	lut_sub lut_2124 ({sk[0], i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_1_, i_2_}, x7042x);
	defparam lut_2124.LUT_SIZE = 9;
	defparam lut_2124.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000008080000000aa000080aa00000000000000000000000000000000;

	lut_sub lut_2127 ({sk[1], i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_2_}, x693x);
	defparam lut_2127.LUT_SIZE = 8;
	defparam lut_2127.mask = 256'h0fffffff0fffffff0fffffff0fffffff00080000000c00000000000000000000;

	lut_sub lut_2130 ({sk[2], i_9_, i_10_, i_7_, i_5_, i_6_, i_12_, i_1_, i_2_}, x1012x);
	defparam lut_2130.LUT_SIZE = 9;
	defparam lut_2130.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff00000000a0808080000000000000808000000000a08000000000000000000000;

	lut_sub lut_2134 ({sk[3], i_9_, i_10_, i_7_, i_5_, i_6_, i_11_, i_2_}, x7047x);
	defparam lut_2134.LUT_SIZE = 8;
	defparam lut_2134.mask = 256'h0fffffff0fffffff0fffffff0fffffff80080000000800008000000000000000;

	lut_sub lut_2137 ({sk[4], i_10_, i_8_, i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x7052x);
	defparam lut_2137.LUT_SIZE = 9;
	defparam lut_2137.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff00000000aaaaaaaa88008000aaaaaaaa00000000aaaaaaaa80008000aaaaaaaa;

	lut_sub lut_2141 ({sk[5], i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_1_}, x1004x);
	defparam lut_2141.LUT_SIZE = 8;
	defparam lut_2141.mask = 256'h0fffffff0fffffff0fffffff0fffffff0000c800000000000000000000000000;

	lut_sub lut_2144 ({sk[6], i_9_, i_8_, i_6_, i_3_, i_2_, i_0_}, x1007x);
	defparam lut_2144.LUT_SIZE = 7;
	defparam lut_2144.mask = 128'h0f0fffffffffffff0000008000000000;

	lut_sub lut_2146 ({sk[7], i_9_, i_10_, i_3_, i_12_, i_1_, i_11_, i_0_}, x700x);
	defparam lut_2146.LUT_SIZE = 8;
	defparam lut_2146.mask = 256'h0fffffff0fffffff0fffffff0fffffff0000000000000000000000080000000d;

	lut_sub lut_2149 ({sk[8], i_7_, i_5_, i_3_, i_1_, i_11_, i_0_}, x699x);
	defparam lut_2149.LUT_SIZE = 7;
	defparam lut_2149.mask = 128'h0f0fffffffffffff0000001100000015;

	lut_sub lut_2152 ({sk[9], i_9_, i_8_, i_5_, i_6_, i_3_, i_12_, i_11_, i_2_}, x150x);
	defparam lut_2152.LUT_SIZE = 9;
	defparam lut_2152.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000100000;

	lut_sub lut_2154 ({sk[10], i_9_, i_7_, i_5_, i_6_, i_12_, i_11_, i_2_, i_0_}, x151x);
	defparam lut_2154.LUT_SIZE = 9;
	defparam lut_2154.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000010011;

	lut_sub lut_2157 ({sk[11], i_9_, i_8_, i_5_, i_6_, i_3_, i_11_, i_2_, i_0_}, x152x);
	defparam lut_2157.LUT_SIZE = 9;
	defparam lut_2157.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000010000;

	lut_sub lut_2159 ({sk[12], i_9_, i_10_, i_8_, i_5_, i_3_, i_1_, i_2_, i_0_}, x153x);
	defparam lut_2159.LUT_SIZE = 9;
	defparam lut_2159.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000010000;

	lut_sub lut_2161 ({sk[13], n_n185, x270x, x700x, x699x, x150x, x151x, x152x, x153x}, n_n994);
	defparam lut_2161.LUT_SIZE = 9;
	defparam lut_2161.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff7fff7fff7fff7fff7fffffff7fffffff7fff7fffffffffff7fffffffffffffff;

	lut_sub lut_2168 ({sk[14], i_5_, i_6_, i_3_, i_1_}, x704x);
	defparam lut_2168.LUT_SIZE = 5;
	defparam lut_2168.mask = 32'h5fff0031;

	lut_sub lut_2171 ({sk[15], i_7_, i_8_, i_5_, i_6_, i_3_, i_1_, i_0_}, x703x);
	defparam lut_2171.LUT_SIZE = 8;
	defparam lut_2171.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000005010000000000000000;

	lut_sub lut_2174 ({sk[0], i_9_, i_7_, i_8_, i_12_, i_11_}, x7274x);
	defparam lut_2174.LUT_SIZE = 6;
	defparam lut_2174.mask = 64'h77ff77ff00000400;

	lut_sub lut_2176 ({sk[1], i_9_, i_7_, i_5_, i_6_, i_12_, i_11_, i_2_, i_0_}, x139x);
	defparam lut_2176.LUT_SIZE = 9;
	defparam lut_2176.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000003010000;

	lut_sub lut_2179 ({sk[2], i_9_, i_5_, i_13_, i_12_, i_11_, i_0_}, x7966x);
	defparam lut_2179.LUT_SIZE = 7;
	defparam lut_2179.mask = 128'h0f0fffffffffffffff7fff5fff7fff0a;

	lut_sub lut_2186 ({sk[3], i_9_, i_11_, x704x, x703x, x7274x, x139x, x7966x}, n_n996);
	defparam lut_2186.LUT_SIZE = 8;
	defparam lut_2186.mask = 256'h0fffffff0fffffff0fffffff0fffffffbbbbbfbfbbbbbfbfbbbbbfbfbbffbfff;

	lut_sub lut_2191 ({sk[4], i_7_, i_8_, i_5_, i_6_, i_3_, i_12_, i_1_, i_0_}, x705x);
	defparam lut_2191.LUT_SIZE = 9;
	defparam lut_2191.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0055000000a00020000000000000000000000000000000000000000000000000;

	lut_sub lut_2195 ({sk[5], i_9_, i_10_, i_5_, i_13_, i_12_, i_11_, i_0_}, x7300x);
	defparam lut_2195.LUT_SIZE = 8;
	defparam lut_2195.mask = 256'h0fffffff0fffffff0fffffff0fffffff0088000000dd0000008800f000dd00f5;

	lut_sub lut_2202 ({sk[6], i_10_, i_5_, i_3_, i_4_, i_1_, i_0_}, x712x);
	defparam lut_2202.LUT_SIZE = 7;
	defparam lut_2202.mask = 128'h0f0fffffffffffff0020000000300000;

	lut_sub lut_2205 ({sk[7], i_9_, i_5_, i_3_, i_4_, i_1_, i_0_}, x708x);
	defparam lut_2205.LUT_SIZE = 7;
	defparam lut_2205.mask = 128'h0f0fffffffffffff0000002000000030;

	lut_sub lut_2208 ({sk[8], i_9_, i_10_, i_5_, i_12_}, x10x);
	defparam lut_2208.LUT_SIZE = 5;
	defparam lut_2208.mask = 32'h5fff0405;

	lut_sub lut_2211 ({sk[9], i_9_, i_10_, i_7_, i_5_, i_12_, i_11_}, x710x);
	defparam lut_2211.LUT_SIZE = 7;
	defparam lut_2211.mask = 128'h0f0fffffffffffff0000500000035003;

	lut_sub lut_2214 ({sk[10], i_9_, i_7_, i_5_, i_3_, i_4_, i_1_, i_11_, i_2_}, x7122x);
	defparam lut_2214.LUT_SIZE = 9;
	defparam lut_2214.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000080a080800000000000a0000000000000000000000000000000000000;

	lut_sub lut_2217 ({sk[11], i_9_, i_5_, i_6_, i_4_, n_n764, n_n672, x406x, x7122x}, x714x);
	defparam lut_2217.LUT_SIZE = 9;
	defparam lut_2217.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff7777777777777777777777777f7f7fff777777777777777777777777777777ff;

	lut_sub lut_2222 ({sk[12], i_9_, i_10_, i_5_, i_12_, i_11_, i_0_}, x717x);
	defparam lut_2222.LUT_SIZE = 7;
	defparam lut_2222.mask = 128'h0f0fffffffffffff0000010000010101;

	lut_sub lut_2226 ({sk[13], i_9_, i_10_, i_8_, i_5_, i_6_, i_12_, i_11_, i_0_}, x716x);
	defparam lut_2226.LUT_SIZE = 9;
	defparam lut_2226.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff000000000008000000000000000d0000000000000008000500000000000d0005;

	lut_sub lut_2231 ({sk[14], i_10_, i_7_, i_8_, i_6_, i_3_, i_1_, i_2_, i_0_}, x763x);
	defparam lut_2231.LUT_SIZE = 9;
	defparam lut_2231.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffffa888a00088880000000000000000000000000000000000000000000000000000;

	lut_sub lut_2234 ({sk[15], i_10_, i_7_, i_8_, i_13_, i_4_, i_12_, i_1_, i_0_}, x864x);
	defparam lut_2234.LUT_SIZE = 9;
	defparam lut_2234.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0008000000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_2236 ({sk[0], i_5_, i_13_, i_12_, i_1_, i_11_, i_2_, i_0_}, x361x);
	defparam lut_2236.LUT_SIZE = 8;
	defparam lut_2236.mask = 256'h0fffffff0fffffff0fffffff0fffffff08000000000000000000000000000000;

	lut_sub lut_2238 ({sk[1], i_10_, i_7_, i_3_, i_13_, i_4_, i_12_, i_0_}, x861x);
	defparam lut_2238.LUT_SIZE = 8;
	defparam lut_2238.mask = 256'h0fffffff0fffffff0fffffff0fffffff02000000000000000000000000000000;

	lut_sub lut_2240 ({sk[2], i_13_, i_12_, i_1_, i_11_, i_0_}, x862x);
	defparam lut_2240.LUT_SIZE = 6;
	defparam lut_2240.mask = 64'h77ff77ff00800000;

	lut_sub lut_2242 ({sk[3], i_7_, i_5_, i_3_, i_1_, i_0_}, x7131x);
	defparam lut_2242.LUT_SIZE = 6;
	defparam lut_2242.mask = 64'h77ff77ff00800000;

	lut_sub lut_2244 ({sk[4], i_7_, i_8_, i_6_, i_3_, i_1_, i_2_, i_0_}, x722x);
	defparam lut_2244.LUT_SIZE = 8;
	defparam lut_2244.mask = 256'h0fffffff0fffffff0fffffff0fffffff0000000080808080a000a000a080aaaa;

	lut_sub lut_2248 ({sk[5], i_8_, i_5_, i_6_, i_3_, i_4_, i_2_, i_0_}, x7146x);
	defparam lut_2248.LUT_SIZE = 8;
	defparam lut_2248.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000800000000000000080800000000;

	lut_sub lut_2251 ({sk[6], i_9_, i_10_, i_5_, i_4_, i_12_, i_11_, i_0_}, x756x);
	defparam lut_2251.LUT_SIZE = 8;
	defparam lut_2251.mask = 256'h0fffffff0fffffff0fffffff0fffffff00002000110020000000310011003100;

	lut_sub lut_2255 ({sk[7], i_9_, i_8_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_}, x755x);
	defparam lut_2255.LUT_SIZE = 9;
	defparam lut_2255.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000880000008000800088008800000000000000000000000000000000;

	lut_sub lut_2259 ({sk[8], i_9_, i_7_, i_8_, i_5_, i_6_, i_4_, i_12_, i_11_}, x834x);
	defparam lut_2259.LUT_SIZE = 9;
	defparam lut_2259.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000004000000000000000000000000000;

	lut_sub lut_2261 ({sk[9], i_9_, i_7_, i_8_, i_6_, i_0_}, x7153x);
	defparam lut_2261.LUT_SIZE = 6;
	defparam lut_2261.mask = 64'h77ff77ff00020000;

	lut_sub lut_2263 ({sk[10], i_4_, n_n853, n_n843, x113x, x756x, x755x, x834x, x7153x}, n_n984);
	defparam lut_2263.LUT_SIZE = 9;
	defparam lut_2263.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff3333ffff33ffffff3f3fffff3fffffff3333ffff33ffffff7f7fffff7fffffff;

	lut_sub lut_2269 ({sk[11], i_6_, i_0_}, x271x);
	defparam lut_2269.LUT_SIZE = 3;
	defparam lut_2269.mask = 8'h58;

	lut_sub lut_2271 ({sk[12], i_4_, n_n792, n_n853, x6718x, n_n699, n_n678, n_n791, x271x}, x7161x);
	defparam lut_2271.LUT_SIZE = 9;
	defparam lut_2271.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff00000000000f000f00000000333f333f00000000000fffff00000000777fffff;

	lut_sub lut_2276 ({sk[13], i_4_, n_n764, n_n853, x394x, n_n791, x399x, x6679x, x108x}, x7162x);
	defparam lut_2276.LUT_SIZE = 9;
	defparam lut_2276.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff000000005555ffff0000000055ffffff000000007f7fffff000000007fffffff;

	lut_sub lut_2282 ({sk[14], i_10_, i_7_, i_8_, i_6_, i_3_, i_1_, i_2_, i_0_}, x725x);
	defparam lut_2282.LUT_SIZE = 9;
	defparam lut_2282.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff8880808080808080880080000000000080808080808080808000800000000000;

	lut_sub lut_2286 ({sk[15], i_10_, i_8_, i_3_, i_13_, i_4_, i_12_, i_2_, i_0_}, x723x);
	defparam lut_2286.LUT_SIZE = 9;
	defparam lut_2286.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0008000000080000000800000000000000000000000000000000000000000000;

	lut_sub lut_2289 ({sk[0], i_8_, i_5_}, x357x);
	defparam lut_2289.LUT_SIZE = 3;
	defparam lut_2289.mask = 8'h54;

	lut_sub lut_2291 ({sk[1], i_9_, i_10_, i_5_, i_6_, i_11_}, x731x);
	defparam lut_2291.LUT_SIZE = 6;
	defparam lut_2291.mask = 64'h77ff77ff00400444;

	lut_sub lut_2294 ({sk[2], i_9_, i_5_, i_3_, i_4_, i_0_}, x730x);
	defparam lut_2294.LUT_SIZE = 6;
	defparam lut_2294.mask = 64'h77ff77ff0008000c;

	lut_sub lut_2297 ({sk[3], i_9_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_}, x729x);
	defparam lut_2297.LUT_SIZE = 8;
	defparam lut_2297.mask = 256'h0fffffff0fffffff0fffffff0fffffff00020000000000000003000100000000;

	lut_sub lut_2301 ({sk[4], i_7_, i_6_, i_12_, i_11_}, x7199x);
	defparam lut_2301.LUT_SIZE = 5;
	defparam lut_2301.mask = 32'h5fff4000;

	lut_sub lut_2303 ({sk[5], i_7_, i_3_, i_4_, i_0_}, x7200x);
	defparam lut_2303.LUT_SIZE = 5;
	defparam lut_2303.mask = 32'h5fff0400;

	lut_sub lut_2305 ({sk[6], i_9_, i_7_, i_5_, i_3_, i_4_, i_1_, i_11_, i_0_}, x247x);
	defparam lut_2305.LUT_SIZE = 9;
	defparam lut_2305.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000001000000000000000000;

	lut_sub lut_2307 ({sk[7], i_10_, i_8_, i_5_, i_4_, i_1_, i_11_, i_2_, i_0_}, x248x);
	defparam lut_2307.LUT_SIZE = 9;
	defparam lut_2307.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000010000000000000000000000000000;

	lut_sub lut_2309 ({sk[8], i_9_, i_10_, i_5_, i_6_, i_12_, i_11_}, x737x);
	defparam lut_2309.LUT_SIZE = 7;
	defparam lut_2309.mask = 128'h0f0fffffffffffff0000030000530353;

	lut_sub lut_2314 ({sk[9], i_10_, i_6_, i_12_, i_1_, i_11_, i_2_, i_0_}, x736x);
	defparam lut_2314.LUT_SIZE = 8;
	defparam lut_2314.mask = 256'h0fffffff0fffffff0fffffff0fffffff00200020002020200031003100312031;

	lut_sub lut_2318 ({sk[10], i_9_, i_10_, i_7_, i_8_, i_5_, i_12_, i_11_, i_0_}, x739x);
	defparam lut_2318.LUT_SIZE = 9;
	defparam lut_2318.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff00000000000008000000000000000d0000000000000008050000000000000d05;

	lut_sub lut_2324 ({sk[11], i_7_, i_8_, i_5_, i_6_, i_12_, i_11_, i_0_}, x218x);
	defparam lut_2324.LUT_SIZE = 8;
	defparam lut_2324.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000000000000000000080000;

	lut_sub lut_2326 ({sk[12], i_10_, i_5_, i_6_, i_3_, i_4_, i_12_, i_11_, i_2_}, x225x);
	defparam lut_2326.LUT_SIZE = 9;
	defparam lut_2326.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000004000000000000000000;

	lut_sub lut_2328 ({sk[13], i_3_, i_4_, i_2_, i_0_}, x7218x);
	defparam lut_2328.LUT_SIZE = 5;
	defparam lut_2328.mask = 32'h5fff0010;

	lut_sub lut_2330 ({sk[14], i_9_, i_7_, i_8_, i_5_, i_6_, i_2_, i_0_}, x744x);
	defparam lut_2330.LUT_SIZE = 8;
	defparam lut_2330.mask = 256'h0fffffff0fffffff0fffffff0fffffff10000000100000005050000010000000;

	lut_sub lut_2333 ({sk[15], i_9_, i_10_, i_7_, i_8_, i_5_, i_12_, i_11_, i_0_}, x742x);
	defparam lut_2333.LUT_SIZE = 9;
	defparam lut_2333.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0020000000000000112000000000000000310000000000001131000000000000;

	lut_sub lut_2338 ({sk[0], i_10_, i_5_, i_6_, i_3_, i_12_, i_11_, i_2_, i_0_}, x750x);
	defparam lut_2338.LUT_SIZE = 9;
	defparam lut_2338.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000101000000000000020000000000;

	lut_sub lut_2341 ({sk[1], i_5_, i_12_, i_1_, i_11_, i_2_, i_0_}, x749x);
	defparam lut_2341.LUT_SIZE = 7;
	defparam lut_2341.mask = 128'h0f0fffffffffffff0031001100200000;

	lut_sub lut_2344 ({sk[2], i_10_, i_7_, i_8_, i_5_, i_3_, i_12_, i_1_, i_0_}, x88x);
	defparam lut_2344.LUT_SIZE = 9;
	defparam lut_2344.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000001000000000000;

	lut_sub lut_2346 ({sk[3], i_10_, i_5_, i_12_, i_11_, i_0_}, x754x);
	defparam lut_2346.LUT_SIZE = 6;
	defparam lut_2346.mask = 64'h77ff77ff08000d00;

	lut_sub lut_2349 ({sk[4], i_7_, i_8_, i_3_, i_12_, i_2_}, x753x);
	defparam lut_2349.LUT_SIZE = 6;
	defparam lut_2349.mask = 64'h77ff77ff00031113;

	lut_sub lut_2352 ({sk[5], i_10_, i_7_, i_6_, i_3_, i_13_, i_12_, i_11_, i_2_}, x59x);
	defparam lut_2352.LUT_SIZE = 9;
	defparam lut_2352.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffffc800880000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_2355 ({sk[6], i_10_, i_7_, i_8_, i_13_, i_4_, i_1_}, x58x);
	defparam lut_2355.LUT_SIZE = 7;
	defparam lut_2355.mask = 128'h0f0fffffffffffff2000000000000000;

	lut_sub lut_2357 ({sk[7], i_10_, i_6_, i_13_, i_12_, i_1_, i_11_, x59x, x58x}, x758x);
	defparam lut_2357.LUT_SIZE = 9;
	defparam lut_2357.mask = 512'h555555ffffffffffffffffffffffffff555555fffffffffffffffffffffffffff777777777777777ff7777777777777777777777777777777777777777777777;

	lut_sub lut_2362 ({sk[8], i_9_, i_10_, i_7_, i_5_, i_6_, i_3_, i_4_}, x546x);
	defparam lut_2362.LUT_SIZE = 8;
	defparam lut_2362.mask = 256'h0fffffff0fffffff0fffffff0fffffff80000008000000088000000000000000;

	lut_sub lut_2365 ({sk[9], i_10_, i_7_, i_8_, i_5_, i_6_, i_1_, i_2_, i_0_}, x550x);
	defparam lut_2365.LUT_SIZE = 9;
	defparam lut_2365.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000002000000000000400800;

	lut_sub lut_2369 ({sk[10], i_9_, i_7_, i_6_, i_2_}, x7313x);
	defparam lut_2369.LUT_SIZE = 5;
	defparam lut_2369.mask = 32'h5fff0001;

	lut_sub lut_2371 ({sk[11], i_9_, i_10_, i_7_, i_5_, i_1_, i_2_, i_0_}, x66x);
	defparam lut_2371.LUT_SIZE = 8;
	defparam lut_2371.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000000000000000000000100;

	lut_sub lut_2373 ({sk[12], i_9_, i_7_, i_5_, i_12_, i_1_, i_11_, i_2_, i_0_}, x67x);
	defparam lut_2373.LUT_SIZE = 9;
	defparam lut_2373.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000020002000330011;

	lut_sub lut_2378 ({sk[13], i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_12_, i_0_}, x87x);
	defparam lut_2378.LUT_SIZE = 9;
	defparam lut_2378.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000001000000000000;

	lut_sub lut_2380 ({sk[14], i_5_, i_6_, i_12_, i_11_}, x7235x);
	defparam lut_2380.LUT_SIZE = 5;
	defparam lut_2380.mask = 32'h5fff0040;

	lut_sub lut_2382 ({sk[15], i_9_, i_8_, i_4_, i_2_, i_0_}, x7236x);
	defparam lut_2382.LUT_SIZE = 6;
	defparam lut_2382.mask = 64'h77ff77ff20003000;

	lut_sub lut_2385 ({sk[0], i_9_, i_8_, i_5_, i_6_, i_4_, i_11_, i_2_, i_0_}, x200x);
	defparam lut_2385.LUT_SIZE = 9;
	defparam lut_2385.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000010000000000000000000000;

	lut_sub lut_2387 ({sk[1], i_5_, i_6_, i_3_, i_4_, i_12_, i_11_, i_2_, i_0_}, x212x);
	defparam lut_2387.LUT_SIZE = 9;
	defparam lut_2387.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000020000000000000000000000;

	lut_sub lut_2389 ({sk[2], i_9_, i_5_, i_6_, i_3_, i_4_, i_12_, i_11_, i_2_}, x213x);
	defparam lut_2389.LUT_SIZE = 9;
	defparam lut_2389.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000100000000000;

	lut_sub lut_2391 ({sk[3], i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_12_, i_0_}, x255x);
	defparam lut_2391.LUT_SIZE = 9;
	defparam lut_2391.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000000001;

	lut_sub lut_2393 ({sk[4], i_8_, i_5_, i_6_, i_3_, i_2_, i_0_}, x7143x);
	defparam lut_2393.LUT_SIZE = 7;
	defparam lut_2393.mask = 128'h0f0fffffffffffff0000000000800000;

	lut_sub lut_2395 ({sk[5], i_10_, i_8_, i_5_, i_6_, i_13_, i_4_, i_11_, i_2_}, x893x);
	defparam lut_2395.LUT_SIZE = 9;
	defparam lut_2395.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0200000000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_2397 ({sk[6], i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_12_}, x971x);
	defparam lut_2397.LUT_SIZE = 8;
	defparam lut_2397.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000000080000000000000000;

	lut_sub lut_2399 ({sk[7], i_10_, i_8_, i_5_, i_6_, i_3_, i_11_, i_2_}, x984x);
	defparam lut_2399.LUT_SIZE = 8;
	defparam lut_2399.mask = 256'h0fffffff0fffffff0fffffff0fffffff80000000000000000000000000000000;

	lut_sub lut_2401 ({sk[8], i_9_, i_7_, i_5_, i_6_, i_3_, i_12_, i_11_}, x985x);
	defparam lut_2401.LUT_SIZE = 8;
	defparam lut_2401.mask = 256'h0fffffff0fffffff0fffffff0fffffff00000000000000800000000000000000;

	lut_sub lut_2403 ({sk[9], i_9_, i_10_, i_5_, i_6_, i_3_, i_12_, i_11_, i_2_}, x986x);
	defparam lut_2403.LUT_SIZE = 9;
	defparam lut_2403.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffffc080c080c080c080000000000000000080800000000000000000000000000000;

	lut_sub lut_2407 ({sk[10], i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_12_, i_11_}, x987x);
	defparam lut_2407.LUT_SIZE = 9;
	defparam lut_2407.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffffa000000080000000000000000000000000000000000000000000000000000000;

	lut_sub lut_2410 ({sk[11], i_10_, i_8_, i_13_, i_4_, i_12_, i_11_, i_2_}, x1167x);
	defparam lut_2410.LUT_SIZE = 8;
	defparam lut_2410.mask = 256'h0fffffff0fffffff0fffffff0fffffff00020000000000000000000000000000;

	lut_sub lut_2412 ({sk[12], i_9_, i_10_, i_7_, i_8_, i_12_, i_11_}, x6786x);
	defparam lut_2412.LUT_SIZE = 7;
	defparam lut_2412.mask = 128'h0f0fffffffffffff1000000000000000;

	lut_sub lut_2414 ({sk[13], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x6753x);
	defparam lut_2414.LUT_SIZE = 7;
	defparam lut_2414.mask = 128'h0f0fffffffffffff0010000000000000;

	lut_sub lut_2416 ({sk[14], i_10_, i_5_, i_3_, i_13_, i_4_, i_12_, i_11_}, x6754x);
	defparam lut_2416.LUT_SIZE = 8;
	defparam lut_2416.mask = 256'h0fffffff0fffffff0fffffff0fffffff20000000000000000000000000000000;

	lut_sub lut_2418 ({sk[15], i_7_, i_8_, i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x1552x);
	defparam lut_2418.LUT_SIZE = 9;
	defparam lut_2418.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000000000000000000000008000;

	lut_sub lut_2420 ({sk[0], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x6697x);
	defparam lut_2420.LUT_SIZE = 7;
	defparam lut_2420.mask = 128'h0f0fffffffffffff0400000000000000;

	lut_sub lut_2422 ({sk[1], i_10_, i_7_, i_5_, i_6_, i_3_, i_1_, i_11_, i_0_}, x1554x);
	defparam lut_2422.LUT_SIZE = 9;
	defparam lut_2422.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff00000000000000000000000000000000cc00c000880080000000000000000000;

	lut_sub lut_2427 ({sk[2], i_9_, i_7_, i_3_, i_4_, i_1_}, x6685x);
	defparam lut_2427.LUT_SIZE = 6;
	defparam lut_2427.mask = 64'h77ff77ff00200000;

	lut_sub lut_2429 ({sk[3], i_3_, i_1_, i_2_, i_0_}, x6686x);
	defparam lut_2429.LUT_SIZE = 5;
	defparam lut_2429.mask = 32'h5fff4000;

	lut_sub lut_2431 ({sk[4], i_10_, i_7_, i_8_, i_6_, i_13_, i_12_}, x6662x);
	defparam lut_2431.LUT_SIZE = 7;
	defparam lut_2431.mask = 128'h0f0fffffffffffff0040000000000000;

	lut_sub lut_2433 ({sk[5], i_9_, i_10_, i_3_, i_13_, i_4_, i_12_, i_11_}, x1605x);
	defparam lut_2433.LUT_SIZE = 8;
	defparam lut_2433.mask = 256'h0fffffff0fffffff0fffffff0fffffff80000000000000000000000000000000;

	lut_sub lut_2435 ({sk[6], i_8_, i_6_, i_3_, i_4_, i_2_, i_0_}, x6596x);
	defparam lut_2435.LUT_SIZE = 7;
	defparam lut_2435.mask = 128'h0f0fffffffffffff0000000010000000;

	lut_sub lut_2437 ({sk[7], i_9_, i_10_, i_5_, i_3_, i_13_, i_4_, i_12_, i_11_}, x6541x);
	defparam lut_2437.LUT_SIZE = 9;
	defparam lut_2437.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000002000000000000000000000000000;

	lut_sub lut_2439 ({sk[8], i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_12_, i_2_}, x1832x);
	defparam lut_2439.LUT_SIZE = 9;
	defparam lut_2439.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000100000001000100010000000100000001000000010001000100010001;

	lut_sub lut_2443 ({sk[9], i_10_, i_7_, i_8_, i_5_, i_3_, i_1_, i_11_, i_2_}, x1841x);
	defparam lut_2443.LUT_SIZE = 9;
	defparam lut_2443.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0303000000030000000000000000000003030000010300000000000000000000;

	lut_sub lut_2447 ({sk[10], i_9_, i_8_, i_5_, i_6_, i_12_, i_1_, i_11_, i_2_}, x6491x);
	defparam lut_2447.LUT_SIZE = 9;
	defparam lut_2447.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000005000500000303000000000000030300050005;

	lut_sub lut_2450 ({sk[11], i_10_, i_7_, i_5_, i_6_, i_3_, i_12_, i_1_, i_2_}, x6496x);
	defparam lut_2450.LUT_SIZE = 9;
	defparam lut_2450.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000005000000000000000500000000010101050000000000000005;

	lut_sub lut_2453 ({sk[12], i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_12_, i_1_}, x7980x);
	defparam lut_2453.LUT_SIZE = 9;
	defparam lut_2453.mask = 512'h555555ffffffffffffffffffffffffff555555fffffffffffffffffffffffffffffffffffffffffffffffffcffffeeccffffffeeffffffeeffffffecffffeecc;

	lut_sub lut_2463 ({sk[13], i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_11_}, x7984x);
	defparam lut_2463.LUT_SIZE = 9;
	defparam lut_2463.mask = 512'h555555ffffffffffffffffffffffffff555555fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7ffffffffffffffffffffffff;

	lut_sub lut_2484 ({sk[14], i_13_, i_12_, i_1_, i_2_, i_0_, n_n748, x6541x, x7984x}, x6552x);
	defparam lut_2484.LUT_SIZE = 9;
	defparam lut_2484.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0003000000000000aa0300000000000000030000000000000003000000000000;

	lut_sub lut_2487 ({sk[15], i_9_, i_5_, i_1_, i_11_, i_2_, i_0_, x21x, n_n752}, x6576x);
	defparam lut_2487.LUT_SIZE = 9;
	defparam lut_2487.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000000000000001000000000000000010001;

	lut_sub lut_2490 ({sk[0], i_10_, i_7_, i_8_, i_5_, i_6_, i_11_, x272x, x306x}, x6805x);
	defparam lut_2490.LUT_SIZE = 9;
	defparam lut_2490.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000075005500000000000000000000000000;

	lut_sub lut_2493 ({sk[1], i_9_, i_10_, i_7_, i_8_, i_4_, i_12_, i_11_, i_2_}, x7972x);
	defparam lut_2493.LUT_SIZE = 9;
	defparam lut_2493.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffffffffffffdfffffffeefffeffdfffffffffffffffcefffeffeefffeffcefffeff;

	lut_sub lut_2504 ({sk[2], i_9_, i_10_, i_7_, i_3_, i_4_, i_12_, i_11_, i_2_}, x7988x);
	defparam lut_2504.LUT_SIZE = 9;
	defparam lut_2504.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff000088000000a0000000dd000000a000000088000000f5000000dd000000f500;

	lut_sub lut_2512 ({sk[3], i_9_, i_10_, i_5_, i_6_, i_12_, i_1_, i_11_, i_2_}, x7986x);
	defparam lut_2512.LUT_SIZE = 9;
	defparam lut_2512.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffffc0c0f000c0c0f80000000000c000f800c000c000000000000000000000000000;

	lut_sub lut_2525 ({sk[4], i_5_, i_13_, i_12_, i_11_, n_n819, n_n678, x121x, x725x}, x7167x);
	defparam lut_2525.LUT_SIZE = 9;
	defparam lut_2525.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff333333333333333f3333333333333333333333337777333f3333333333333333;

	lut_sub lut_2529 ({sk[5], i_5_, i_6_, i_3_, i_0_, x37x, n_n725, n_n843, x723x}, x7168x);
	defparam lut_2529.LUT_SIZE = 9;
	defparam lut_2529.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff0000000000000000000000000000000057775555557755550333000000330000;

	lut_sub lut_2533 ({sk[6], i_5_, i_6_, i_3_, i_12_, i_1_, i_11_}, x7965x);
	defparam lut_2533.LUT_SIZE = 7;
	defparam lut_2533.mask = 128'h0f0ffffffffffffffffdfff5ffffffff;

	lut_sub lut_2547 ({sk[7], i_9_, i_0_, n_n213, x754x, x753x, x7313x, x66x, x67x}, x7318x);
	defparam lut_2547.LUT_SIZE = 9;
	defparam lut_2547.mask = 512'h555555ffffffffffffffffffffffffff555555ffffffffffffffffffffffffff77777f7f77777f7f77777f7f77777f7f77777f7f77777f7f77777f7f77ff7fff;


endmodule