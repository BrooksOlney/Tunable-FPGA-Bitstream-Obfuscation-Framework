module pdcx6xv (i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, i_13_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_, i_15_, o_1_, o_19_, o_2_, o_0_, o_29_, o_39_, o_38_, o_25_, o_12_, o_37_, o_26_, o_11_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_, o_16_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_30_, o_20_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

	input i_9_;
	input i_10_;
	input i_7_;
	input i_8_;
	input i_5_;
	input i_6_;
	input i_14_;
	input i_3_;
	input i_13_;
	input i_4_;
	input i_12_;
	input i_1_;
	input i_11_;
	input i_2_;
	input i_0_;
	input i_15_;
	output o_1_;
	output o_19_;
	output o_2_;
	output o_0_;
	output o_29_;
	output o_39_;
	output o_38_;
	output o_25_;
	output o_12_;
	output o_37_;
	output o_26_;
	output o_11_;
	output o_36_;
	output o_27_;
	output o_14_;
	output o_35_;
	output o_28_;
	output o_13_;
	output o_34_;
	output o_21_;
	output o_16_;
	output o_33_;
	output o_22_;
	output o_15_;
	output o_32_;
	output o_23_;
	output o_18_;
	output o_31_;
	output o_24_;
	output o_17_;
	output o_30_;
	output o_20_;
	output o_10_;
	output o_9_;
	output o_7_;
	output o_8_;
	output o_5_;
	output o_6_;
	output o_3_;
	output o_4_;

	wire [2993 : 0] sk /* synthesis noprune */;

	lut_sub lut_3 ({sk[0], n_n5231, x507x, x19375x, x24150x}, o_1_);
	defparam lut_3.LUT_SIZE = 5;
	defparam lut_3.mask = 32'h55ffbfff;

	lut_sub lut_8 ({sk[1], n_n5231, n_n3619, n_n3621, x19589x, x19590x, x19591x}, o_19_);
	defparam lut_8.LUT_SIZE = 7;
	defparam lut_8.mask = 128'h05ff05ffffffffff7fffffffffffffff;

	lut_sub lut_15 ({sk[2], n_n5231, x5464x, x19600x, x19602x}, o_2_);
	defparam lut_15.LUT_SIZE = 5;
	defparam lut_15.mask = 32'h55ff7fff;

	lut_sub lut_20 ({sk[3], n_n5231, x5457x, x19610x, x19619x, x19620x}, o_0_);
	defparam lut_20.LUT_SIZE = 6;
	defparam lut_20.mask = 64'h777777777fffffff;

	lut_sub lut_26 ({sk[4], n_n5231, n_n4442, n_n4440, n_n4441, n_n4439, x19644x}, o_29_);
	defparam lut_26.LUT_SIZE = 7;
	defparam lut_26.mask = 128'h05ff05ffffffffff7fffffffffffffff;

	lut_sub lut_33 ({sk[5], i_7_, i_6_, i_4_, n_n5231, x260x, x259x}, o_39_);
	defparam lut_33.LUT_SIZE = 7;
	defparam lut_33.mask = 128'h05ff05ffffffffff0f0f3f7f0f0f0f0f;

	lut_sub lut_37 ({sk[6], i_7_, i_6_, i_4_, n_n5231, x260x, x259x}, o_38_);
	defparam lut_37.LUT_SIZE = 7;
	defparam lut_37.mask = 128'h05ff05ffffffffff0f0f0f0f3f7f0f0f;

	lut_sub lut_41 ({sk[7], n_n5231, x19736x, n_n4307, n_n4308, x19766x}, o_25_);
	defparam lut_41.LUT_SIZE = 6;
	defparam lut_41.mask = 64'h5555ffff7fffffff;

	lut_sub lut_47 ({sk[8], n_n5231, n_n2570, x19821x}, o_12_);
	defparam lut_47.LUT_SIZE = 4;
	defparam lut_47.mask = 16'h117f;

	lut_sub lut_51 ({sk[9], n_n5231, x19830x, x19835x, x5140x, x19837x, x24141x}, o_37_);
	defparam lut_51.LUT_SIZE = 7;
	defparam lut_51.mask = 128'h11551177ffffffffbfffffffffffffff;

	lut_sub lut_58 ({sk[10], n_n5231, n_n227, x5130x, x1814x, x19843x, x24176x}, o_26_);
	defparam lut_58.LUT_SIZE = 7;
	defparam lut_58.mask = 128'h11551177ffffffffbbffbfffffffffff;

	lut_sub lut_64 ({sk[11], n_n5231, x19850x, n_n2547, x19859x, x24177x}, o_11_);
	defparam lut_64.LUT_SIZE = 6;
	defparam lut_64.mask = 64'h5555ffffbfffffff;

	lut_sub lut_70 ({sk[12], n_n5231, x19890x, x19891x, n_n4720, n_n4718, x19990x}, o_36_);
	defparam lut_70.LUT_SIZE = 7;
	defparam lut_70.mask = 128'h11551177ffffffff7fffffffffffffff;

	lut_sub lut_77 ({sk[13], i_7_, i_6_, n_n5231, n_n264, n_n120}, o_27_);
	defparam lut_77.LUT_SIZE = 6;
	defparam lut_77.mask = 64'h5555ffff0f0f0f1f;

	lut_sub lut_80 ({sk[14], n_n5231, n_n153, x583x, x450x, x261x, x20003x}, o_14_);
	defparam lut_80.LUT_SIZE = 7;
	defparam lut_80.mask = 128'h11551177ffffffff5fff7fffffffffff;

	lut_sub lut_86 ({sk[15], n_n5231, n_n152, n_n4705, x20008x, x1704x, x20012x}, o_35_);
	defparam lut_86.LUT_SIZE = 7;
	defparam lut_86.mask = 128'h11551177ffffffff5fff7fffffffffff;

	lut_sub lut_92 ({sk[16], n_n5231, n_n4413, n_n4415, n_n4416, n_n4418, x20033x}, o_28_);
	defparam lut_92.LUT_SIZE = 7;
	defparam lut_92.mask = 128'h11551177ffffffff7fffffffffffffff;

	lut_sub lut_99 ({sk[17], n_n5231, n_n5240}, o_13_);
	defparam lut_99.LUT_SIZE = 3;
	defparam lut_99.mask = 8'h17;

	lut_sub lut_102 ({sk[18], n_n5231, n_n4530, x20245x}, o_34_);
	defparam lut_102.LUT_SIZE = 4;
	defparam lut_102.mask = 16'h117f;

	lut_sub lut_106 ({sk[19], n_n5231, n_n3892, x20353x, n_n3918, n_n3919}, o_21_);
	defparam lut_106.LUT_SIZE = 6;
	defparam lut_106.mask = 64'h5555ffff7fffffff;

	lut_sub lut_112 ({sk[20], n_n5231, x20571x, n_n2792, n_n2793, x20626x}, o_16_);
	defparam lut_112.LUT_SIZE = 6;
	defparam lut_112.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_118 ({sk[21], n_n5231, n_n4512, x20635x, x20636x, n_n4508, x20647x}, o_33_);
	defparam lut_118.LUT_SIZE = 7;
	defparam lut_118.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_125 ({sk[22], n_n5231, x392x, x490x, x735x, x822x, x20659x}, o_22_);
	defparam lut_125.LUT_SIZE = 7;
	defparam lut_125.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_132 ({sk[23], i_2_, i_0_, n_n5247, x535x, n_n4495, x450x}, o_15_);
	defparam lut_132.LUT_SIZE = 7;
	defparam lut_132.mask = 128'h5555ffff5555ffff7fff7fffffff7fff;

	lut_sub lut_138 ({sk[24], n_n5231, x20672x}, o_32_);
	defparam lut_138.LUT_SIZE = 3;
	defparam lut_138.mask = 8'h57;

	lut_sub lut_141 ({sk[25], n_n5231, n_n4194, x20753x}, o_23_);
	defparam lut_141.LUT_SIZE = 4;
	defparam lut_141.mask = 16'h557f;

	lut_sub lut_145 ({sk[26], n_n5231, n_n3361, n_n3360, x20913x, x20914x}, o_18_);
	defparam lut_145.LUT_SIZE = 6;
	defparam lut_145.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_151 ({sk[27], n_n5231, x935x, x758x, x923x, x3945x, x20920x}, o_31_);
	defparam lut_151.LUT_SIZE = 7;
	defparam lut_151.mask = 128'h5555ffff5555ffff77ff7fffffffffff;

	lut_sub lut_157 ({sk[28], n_n5231, x20924x}, o_24_);
	defparam lut_157.LUT_SIZE = 3;
	defparam lut_157.mask = 8'h57;

	lut_sub lut_160 ({sk[29], x21156x, x21063x, x21064x, n_n3093, x21129x, x21130x}, o_17_);
	defparam lut_160.LUT_SIZE = 7;
	defparam lut_160.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_167 ({sk[30], n_n5231, x21179x}, o_30_);
	defparam lut_167.LUT_SIZE = 3;
	defparam lut_167.mask = 8'h57;

	lut_sub lut_170 ({sk[31], n_n5231, n_n3892, n_n3890, n_n3896, x21292x}, o_20_);
	defparam lut_170.LUT_SIZE = 6;
	defparam lut_170.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_176 ({sk[32], n_n5231, x21359x, x21319x, x21320x, n_n2428, x21364x}, o_10_);
	defparam lut_176.LUT_SIZE = 7;
	defparam lut_176.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_183 ({sk[33], n_n5231, n_n2058, x21618x, x21619x, x21620x}, o_9_);
	defparam lut_183.LUT_SIZE = 6;
	defparam lut_183.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_189 ({sk[34], n_n5231, n_n148, n_n106, n_n126, x3242x, x21631x}, o_7_);
	defparam lut_189.LUT_SIZE = 7;
	defparam lut_189.mask = 128'h5555ffff5555ffff777f7f7fffffffff;

	lut_sub lut_195 ({sk[35], n_n5231, x21881x, n_n1680, x21880x, x21904x}, o_8_);
	defparam lut_195.LUT_SIZE = 6;
	defparam lut_195.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_201 ({sk[36], n_n5231, x22334x, x22331x}, o_5_);
	defparam lut_201.LUT_SIZE = 4;
	defparam lut_201.mask = 16'h557f;

	lut_sub lut_205 ({sk[37], i_3_, i_1_, i_2_, i_0_, n_n5247}, o_6_);
	defparam lut_205.LUT_SIZE = 6;
	defparam lut_205.mask = 64'h3f3f3f3f5555dd55;

	lut_sub lut_209 ({sk[38], n_n5231, x22588x, n_n341, x22583x, x24074x}, o_3_);
	defparam lut_209.LUT_SIZE = 6;
	defparam lut_209.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_215 ({sk[39], n_n5231, x22827x, n_n732, x22826x, x22847x}, o_4_);
	defparam lut_215.LUT_SIZE = 6;
	defparam lut_215.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_221 ({sk[40], n_n5007, n_n5005, n_n5004, x19357x, n_n5006, x19359x}, n_n5231);
	defparam lut_221.LUT_SIZE = 7;
	defparam lut_221.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_228 ({sk[41], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, x507x);
	defparam lut_228.LUT_SIZE = 7;
	defparam lut_228.mask = 128'h5555ffff5555ffff0010101010101000;

	lut_sub lut_235 ({sk[42], n_n139, x19365x, n_n111, x251x, x54x, x19373x}, x19375x);
	defparam lut_235.LUT_SIZE = 7;
	defparam lut_235.mask = 128'h5555ffff5555ffff5555ffff7fffffff;

	lut_sub lut_241 ({sk[43], n_n139, n_n152, x48x, n_n110, x54x, x19369x}, x24150x);
	defparam lut_241.LUT_SIZE = 7;
	defparam lut_241.mask = 128'h5555ffff5555ffffaaaa8080a0008000;

	lut_sub lut_246 ({sk[44], n_n3638, x19399x, x19420x, x19421x}, n_n3619);
	defparam lut_246.LUT_SIZE = 5;
	defparam lut_246.mask = 32'h0f0f7fff;

	lut_sub lut_251 ({sk[45], x19530x, x832x, x19504x, x19505x, x19523x}, n_n3621);
	defparam lut_251.LUT_SIZE = 6;
	defparam lut_251.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_257 ({sk[46], x19435x, x19436x, x19456x, x19453x, x19454x}, x19589x);
	defparam lut_257.LUT_SIZE = 6;
	defparam lut_257.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_263 ({sk[47], x19481x, x19546x, x19547x, n_n3686, x19477x, x19478x}, x19590x);
	defparam lut_263.LUT_SIZE = 7;
	defparam lut_263.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_270 ({sk[48], x19573x, x19574x, x19586x, x19582x, x19583x, x19587x}, x19591x);
	defparam lut_270.LUT_SIZE = 7;
	defparam lut_270.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_277 ({sk[49], n_n281, x913x, x921x, n_n208, x907x, x914x}, x5464x);
	defparam lut_277.LUT_SIZE = 7;
	defparam lut_277.mask = 128'h5555ffff5555ffff000000000007000f;

	lut_sub lut_281 ({sk[50], i_7_, i_6_, x364x, n_n118, n_n264, n_n116}, x19600x);
	defparam lut_281.LUT_SIZE = 7;
	defparam lut_281.mask = 128'h5555ffff5555ffff13ff13ff13ff13ff;

	lut_sub lut_291 ({sk[51], i_9_, i_10_, x48x, n_n110, n_n124, x819x}, x19602x);
	defparam lut_291.LUT_SIZE = 7;
	defparam lut_291.mask = 128'h5555ffff5555ffff7777577757775777;

	lut_sub lut_296 ({sk[52], x921x, n_n283, n_n107, x250x, x283x, x19607x}, x5457x);
	defparam lut_296.LUT_SIZE = 7;
	defparam lut_296.mask = 128'h5555ffff5555ffff0000000000007fff;

	lut_sub lut_301 ({sk[53], x48x, n_n110, n_n124, x364x, n_n5769, x54x}, x19610x);
	defparam lut_301.LUT_SIZE = 7;
	defparam lut_301.mask = 128'h5555ffff5555ffff3f7f3fff3fff3fff;

	lut_sub lut_307 ({sk[54], n_n151, n_n5671, n_n148, n_n5678, x396x, x583x}, x19619x);
	defparam lut_307.LUT_SIZE = 7;
	defparam lut_307.mask = 128'h5555ffff5555ffff5f7fffff7f7fffff;

	lut_sub lut_313 ({sk[55], n_n124, n_n163, x582x, x294x, n_n108, x5444x}, x19620x);
	defparam lut_313.LUT_SIZE = 7;
	defparam lut_313.mask = 128'h5555ffff5555ffff55ff55ff7fffffff;

	lut_sub lut_319 ({sk[56], x19627x, n_n271, x896x, x54x, x609x}, n_n4442);
	defparam lut_319.LUT_SIZE = 6;
	defparam lut_319.mask = 64'h3f3f3f3f5557ffff;

	lut_sub lut_323 ({sk[57], n_n139, n_n124, n_n127, n_n111, n_n132, x54x}, n_n4440);
	defparam lut_323.LUT_SIZE = 7;
	defparam lut_323.mask = 128'h5555ffff5555ffff115f5f5f1f5f5f5f;

	lut_sub lut_330 ({sk[58], n_n130, n_n121, n_n111, n_n122, n_n132, x54x}, n_n4441);
	defparam lut_330.LUT_SIZE = 7;
	defparam lut_330.mask = 128'h5555ffff5555ffff053f55ff557f55ff;

	lut_sub lut_337 ({sk[59], i_7_, i_6_, n_n139, x19639x, x924x, x54x}, n_n4439);
	defparam lut_337.LUT_SIZE = 7;
	defparam lut_337.mask = 128'h5555ffff5555ffff0f5f0f5f0f5f3f7f;

	lut_sub lut_341 ({sk[60], i_7_, i_6_, x927x, x929x, x19643x, x24167x}, x19644x);
	defparam lut_341.LUT_SIZE = 7;
	defparam lut_341.mask = 128'h5555ffff5555ffffbbbbbbbbbfbfbfff;

	lut_sub lut_347 ({sk[61], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x260x);
	defparam lut_347.LUT_SIZE = 7;
	defparam lut_347.mask = 128'h5555ffff5555ffff0000000800000000;

	lut_sub lut_349 ({sk[62], i_5_, i_3_, i_1_, i_2_, i_0_}, x259x);
	defparam lut_349.LUT_SIZE = 6;
	defparam lut_349.mask = 64'h3f3f3f3f00000008;

	lut_sub lut_351 ({sk[63], x19723x, x19724x, x19727x, x19728x, x19732x, x19733x}, x19736x);
	defparam lut_351.LUT_SIZE = 7;
	defparam lut_351.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_358 ({sk[64], x5341x, x19686x, n_n4316, x473x, x19694x, x19697x}, n_n4307);
	defparam lut_358.LUT_SIZE = 7;
	defparam lut_358.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_365 ({sk[65], x19703x, x19704x, x19709x, x19710x, x19717x}, n_n4308);
	defparam lut_365.LUT_SIZE = 6;
	defparam lut_365.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_371 ({sk[66], x19677x, x19678x, x513x, x551x, x19761x, x19762x}, x19766x);
	defparam lut_371.LUT_SIZE = 7;
	defparam lut_371.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_378 ({sk[67], x19778x, x19779x, x19793x, x19794x, x19810x, x19811x}, n_n2570);
	defparam lut_378.LUT_SIZE = 7;
	defparam lut_378.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_385 ({sk[68], n_n2, x5161x, x137x, x132x, x5153x, x19819x}, x19821x);
	defparam lut_385.LUT_SIZE = 7;
	defparam lut_385.mask = 128'h5555ffff5555ffff7777ffff7fffffff;

	lut_sub lut_391 ({sk[69], n_n5671, n_n5678, x582x, n_n121, x1359x, x5144x}, x19830x);
	defparam lut_391.LUT_SIZE = 7;
	defparam lut_391.mask = 128'h5555ffff5555ffff57ffffffffffffff;

	lut_sub lut_397 ({sk[70], i_9_, i_10_, x48x, n_n110, n_n124, x5139x}, x19835x);
	defparam lut_397.LUT_SIZE = 7;
	defparam lut_397.mask = 128'h5555ffff5555ffff7777577757775777;

	lut_sub lut_402 ({sk[71], x48x, n_n110, n_n108, n_n122, x103x, x54x}, x5140x);
	defparam lut_402.LUT_SIZE = 7;
	defparam lut_402.mask = 128'h5555ffff5555ffff070f0f0f0f0f0f0f;

	lut_sub lut_408 ({sk[72], i_7_, i_8_, i_6_, x48x, n_n165, n_n284}, x19837x);
	defparam lut_408.LUT_SIZE = 7;
	defparam lut_408.mask = 128'h5555ffff5555ffff0100000011001100;

	lut_sub lut_411 ({sk[73], x364x, x819x, x583x, x318x, x758x, x757x}, x24141x);
	defparam lut_411.LUT_SIZE = 7;
	defparam lut_411.mask = 128'h5555ffff5555ffff8000000000000000;

	lut_sub lut_413 ({sk[74], i_7_, i_8_, i_6_, x909x}, n_n227);
	defparam lut_413.LUT_SIZE = 5;
	defparam lut_413.mask = 32'h0f0f1000;

	lut_sub lut_415 ({sk[75], i_14_, i_13_, i_12_, x902x, n_n227}, x5130x);
	defparam lut_415.LUT_SIZE = 6;
	defparam lut_415.mask = 64'h3f3f3f3f00001110;

	lut_sub lut_419 ({sk[76], i_14_, i_13_, i_12_, i_15_, n_n259, x275x}, x1814x);
	defparam lut_419.LUT_SIZE = 7;
	defparam lut_419.mask = 128'h5555ffff5555ffff5577555575577575;

	lut_sub lut_427 ({sk[77], n_n208, x909x, n_n228, x902x, n_n227, x897x}, x19843x);
	defparam lut_427.LUT_SIZE = 7;
	defparam lut_427.mask = 128'h5555ffff5555ffff0013001300130057;

	lut_sub lut_431 ({sk[78], n_n9, n_n207, x480x, x262x, n_n3550, x1813x}, x24176x);
	defparam lut_431.LUT_SIZE = 7;
	defparam lut_431.mask = 128'h5555ffff5555ffffcc008000cc000000;

	lut_sub lut_434 ({sk[79], n_n281, x907x, n_n265, x101x, n_n62, x598x}, x19850x);
	defparam lut_434.LUT_SIZE = 7;
	defparam lut_434.mask = 128'h5555ffff5555ffff557f557f557f55ff;

	lut_sub lut_439 ({sk[80], x916x, n_n271, x124x, n_n3513, x1729x, x24152x}, n_n2547);
	defparam lut_439.LUT_SIZE = 7;
	defparam lut_439.mask = 128'h5555ffff5555ffffafafafafafafbfff;

	lut_sub lut_444 ({sk[81], x916x, n_n271, x400x, x157x, x156x, x19857x}, x19859x);
	defparam lut_444.LUT_SIZE = 7;
	defparam lut_444.mask = 128'h5555ffff5555ffff5555555555557fff;

	lut_sub lut_449 ({sk[82], n_n268, n_n3246, x206x, n_n240, n_n59, x1326x}, x24177x);
	defparam lut_449.LUT_SIZE = 7;
	defparam lut_449.mask = 128'h5555ffff5555ffffffff000080000000;

	lut_sub lut_452 ({sk[83], x909x, n_n261, x156x, x24140x, x24174x}, x19890x);
	defparam lut_452.LUT_SIZE = 6;
	defparam lut_452.mask = 64'h3f3f3f3feeeeeeef;

	lut_sub lut_456 ({sk[84], x19882x, x19883x, x19876x, x19877x, x24139x}, x19891x);
	defparam lut_456.LUT_SIZE = 6;
	defparam lut_456.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_462 ({sk[85], x19896x, x19897x, x19900x, x19901x, x19904x, x19905x}, n_n4720);
	defparam lut_462.LUT_SIZE = 7;
	defparam lut_462.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_469 ({sk[86], x19982x, x19946x, x19947x, n_n4744, x19968x}, n_n4718);
	defparam lut_469.LUT_SIZE = 6;
	defparam lut_469.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_475 ({sk[87], x19872x, x19873x, x19921x, x19922x, x19987x}, x19990x);
	defparam lut_475.LUT_SIZE = 6;
	defparam lut_475.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_481 ({sk[88], i_5_, i_3_, i_4_}, n_n264);
	defparam lut_481.LUT_SIZE = 4;
	defparam lut_481.mask = 16'h5508;

	lut_sub lut_483 ({sk[89], i_1_, i_2_, i_0_}, n_n120);
	defparam lut_483.LUT_SIZE = 4;
	defparam lut_483.mask = 16'h5504;

	lut_sub lut_485 ({sk[90], i_7_, i_6_}, n_n153);
	defparam lut_485.LUT_SIZE = 3;
	defparam lut_485.mask = 8'h51;

	lut_sub lut_487 ({sk[91], i_7_, i_5_, i_6_, i_3_, i_4_, n_n118}, x583x);
	defparam lut_487.LUT_SIZE = 7;
	defparam lut_487.mask = 128'h5555ffff5555ffff4040404040404040;

	lut_sub lut_496 ({sk[92], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, x450x);
	defparam lut_496.LUT_SIZE = 7;
	defparam lut_496.mask = 128'h5555ffff5555ffff5555151555151515;

	lut_sub lut_509 ({sk[93], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x261x);
	defparam lut_509.LUT_SIZE = 7;
	defparam lut_509.mask = 128'h5555ffff5555ffff0000000000100000;

	lut_sub lut_511 ({sk[94], i_3_, x535x, n_n118, n_n4495, n_n5668, x859x}, x20003x);
	defparam lut_511.LUT_SIZE = 7;
	defparam lut_511.mask = 128'h5555ffff5555ffff7f7fffff7fffffff;

	lut_sub lut_517 ({sk[95], i_7_, i_8_, i_6_, x917x}, n_n152);
	defparam lut_517.LUT_SIZE = 5;
	defparam lut_517.mask = 32'h0f0f4000;

	lut_sub lut_519 ({sk[96], n_n110, n_n124, x20007x, n_n111, n_n108, n_n132}, n_n4705);
	defparam lut_519.LUT_SIZE = 7;
	defparam lut_519.mask = 128'h5555ffff5555ffff15ff3fff55ffffff;

	lut_sub lut_527 ({sk[97], n_n139, x913x, n_n127, n_n220, x914x, x905x}, x20008x);
	defparam lut_527.LUT_SIZE = 7;
	defparam lut_527.mask = 128'h5555ffff5555ffff0000000f07070f0f;

	lut_sub lut_532 ({sk[98], i_9_, i_10_, i_11_, i_15_, n_n220}, x1704x);
	defparam lut_532.LUT_SIZE = 6;
	defparam lut_532.mask = 64'h3f3f3f3fff404040;

	lut_sub lut_537 ({sk[99], n_n110, n_n121, n_n111, n_n128, n_n122, x20011x}, x20012x);
	defparam lut_537.LUT_SIZE = 7;
	defparam lut_537.mask = 128'h5555ffff5555ffff557f557f7f7fffff;

	lut_sub lut_544 ({sk[100], n_n139, n_n152, x48x, n_n110, x289x, x260x}, n_n4413);
	defparam lut_544.LUT_SIZE = 7;
	defparam lut_544.mask = 128'h5555ffff5555ffff11111fff11ff1fff;

	lut_sub lut_549 ({sk[101], x48x, n_n110, n_n130, n_n121, n_n122, n_n132}, n_n4415);
	defparam lut_549.LUT_SIZE = 7;
	defparam lut_549.mask = 128'h5555ffff5555ffff00007f7f3fff7fff;

	lut_sub lut_556 ({sk[102], x48x, n_n110, n_n130, n_n128, x20021x, x4892x}, n_n4416);
	defparam lut_556.LUT_SIZE = 7;
	defparam lut_556.mask = 128'h5555ffff5555ffff77777fff7f7f7fff;

	lut_sub lut_562 ({sk[103], i_7_, i_6_, x919x, x920x, x20027x, x261x}, n_n4418);
	defparam lut_562.LUT_SIZE = 7;
	defparam lut_562.mask = 128'h5555ffff5555ffff3fff77ff33333333;

	lut_sub lut_568 ({sk[104], n_n139, x48x, n_n110, n_n132, x1076x, x20032x}, x20033x);
	defparam lut_568.LUT_SIZE = 7;
	defparam lut_568.mask = 128'h5555ffff5555ffff55777f7f55ff7fff;

	lut_sub lut_574 ({sk[105], x20054x, x20055x, n_n2656, n_n2657, n_n2659, x20113x}, n_n5240);
	defparam lut_574.LUT_SIZE = 7;
	defparam lut_574.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_581 ({sk[106], x20209x, x20210x, n_n4556, x20232x, x20233x, x20240x}, n_n4530);
	defparam lut_581.LUT_SIZE = 7;
	defparam lut_581.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_588 ({sk[107], n_n4548, x20130x, x20147x, x20148x, n_n4532, n_n4531}, x20245x);
	defparam lut_588.LUT_SIZE = 7;
	defparam lut_588.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_595 ({sk[108], n_n3901, n_n3925, n_n3923, x20295x, x24134x}, n_n3892);
	defparam lut_595.LUT_SIZE = 6;
	defparam lut_595.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_601 ({sk[109], n_n108, n_n53, x676x, x298x, x20350x, x24196x}, x20353x);
	defparam lut_601.LUT_SIZE = 7;
	defparam lut_601.mask = 128'h5555ffff5555ffffbfffbfffbfffffff;

	lut_sub lut_607 ({sk[110], n_n48, x213x, n_n3974, n_n4090, x20328x, x20330x}, n_n3918);
	defparam lut_607.LUT_SIZE = 7;
	defparam lut_607.mask = 128'h5555ffff5555ffff7fff7fff7fffffff;

	lut_sub lut_613 ({sk[111], x475x, n_n6879, x474x, x20341x, x20339x}, n_n3919);
	defparam lut_613.LUT_SIZE = 6;
	defparam lut_613.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_619 ({sk[112], n_n2798, n_n2817, n_n2796, x24199x}, x20571x);
	defparam lut_619.LUT_SIZE = 5;
	defparam lut_619.mask = 32'h0f0fbfff;

	lut_sub lut_624 ({sk[113], x20452x, x20453x, n_n2801, x20482x, x20483x}, n_n2792);
	defparam lut_624.LUT_SIZE = 6;
	defparam lut_624.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_630 ({sk[114], x20553x, n_n2803, x20544x, x20545x}, n_n2793);
	defparam lut_630.LUT_SIZE = 5;
	defparam lut_630.mask = 32'h0f0f7fff;

	lut_sub lut_635 ({sk[115], x20590x, x20591x, n_n2795, n_n2840, n_n2839, x20622x}, x20626x);
	defparam lut_635.LUT_SIZE = 7;
	defparam lut_635.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_642 ({sk[116], n_n133, n_n121, x20630x, n_n135, n_n132, n_n107}, n_n4512);
	defparam lut_642.LUT_SIZE = 7;
	defparam lut_642.mask = 128'h5555ffff5555ffff11ff1fff11ffffff;

	lut_sub lut_647 ({sk[117], i_7_, i_5_, i_6_, i_3_, i_4_, n_n118}, x20635x);
	defparam lut_647.LUT_SIZE = 7;
	defparam lut_647.mask = 128'h5555ffff5555ffff5000400000000000;

	lut_sub lut_651 ({sk[118], i_7_, i_6_, n_n264, n_n116, x261x, x4238x}, x20636x);
	defparam lut_651.LUT_SIZE = 7;
	defparam lut_651.mask = 128'h5555ffff5555ffff77775555555f5555;

	lut_sub lut_655 ({sk[119], n_n133, n_n135, n_n132, n_n107, x1784x, x20639x}, n_n4508);
	defparam lut_655.LUT_SIZE = 7;
	defparam lut_655.mask = 128'h5555ffff5555ffff575777ff77ff77ff;

	lut_sub lut_662 ({sk[120], i_7_, i_6_, x936x, n_n128, x216x, x24151x}, x20647x);
	defparam lut_662.LUT_SIZE = 7;
	defparam lut_662.mask = 128'h5555ffff5555ffffabffabababffabab;

	lut_sub lut_667 ({sk[121], i_7_, i_8_, i_6_, x915x, n_n54, n_n105}, x392x);
	defparam lut_667.LUT_SIZE = 7;
	defparam lut_667.mask = 128'h5555ffff5555ffff0000000000030005;

	lut_sub lut_670 ({sk[122], i_7_, i_8_, i_6_, x915x, n_n258, x899x}, x490x);
	defparam lut_670.LUT_SIZE = 7;
	defparam lut_670.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_672 ({sk[123], i_7_, i_8_, i_6_, x915x, n_n258, x897x}, x735x);
	defparam lut_672.LUT_SIZE = 7;
	defparam lut_672.mask = 128'h5555ffff5555ffff0000000000000001;

	lut_sub lut_674 ({sk[124], i_7_, i_8_, i_6_, x915x, n_n258, x901x}, x822x);
	defparam lut_674.LUT_SIZE = 7;
	defparam lut_674.mask = 128'h5555ffff5555ffff0000000000000001;

	lut_sub lut_676 ({sk[125], n_n255, n_n4186, x559x, n_n258, x912x, x902x}, x20659x);
	defparam lut_676.LUT_SIZE = 7;
	defparam lut_676.mask = 128'h5555ffff5555ffff00ffffff07ffffff;

	lut_sub lut_681 ({sk[126], n_n5007, n_n5005, n_n5004, x19357x, n_n5006, x20662x}, n_n5247);
	defparam lut_681.LUT_SIZE = 7;
	defparam lut_681.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_688 ({sk[127], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, x535x);
	defparam lut_688.LUT_SIZE = 7;
	defparam lut_688.mask = 128'h5555ffff5555ffff0000000000004040;

	lut_sub lut_691 ({sk[128], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, n_n4495);
	defparam lut_691.LUT_SIZE = 7;
	defparam lut_691.mask = 128'h5555ffff5555ffff0000404000400000;

	lut_sub lut_695 ({sk[129], i_7_, i_5_, i_6_, i_3_, i_4_, n_n165}, x20672x);
	defparam lut_695.LUT_SIZE = 7;
	defparam lut_695.mask = 128'h5555ffff5555ffff0000010050510001;

	lut_sub lut_703 ({sk[130], n_n4219, x20718x, x20733x, x20734x, x20741x, x20742x}, n_n4194);
	defparam lut_703.LUT_SIZE = 7;
	defparam lut_703.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_710 ({sk[131], x513x, n_n4211, x20686x, n_n4197, x20748x, x20749x}, x20753x);
	defparam lut_710.LUT_SIZE = 7;
	defparam lut_710.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_717 ({sk[132], x811x, x20771x, x20782x, x20783x, x20786x, x20787x}, n_n3361);
	defparam lut_717.LUT_SIZE = 7;
	defparam lut_717.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_724 ({sk[133], x832x, x20836x, n_n3367, x20856x, x20857x}, n_n3360);
	defparam lut_724.LUT_SIZE = 6;
	defparam lut_724.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_730 ({sk[134], x20872x, x20873x, x20895x, x20896x}, x20913x);
	defparam lut_730.LUT_SIZE = 5;
	defparam lut_730.mask = 32'h0f0f7fff;

	lut_sub lut_735 ({sk[135], n_n3375, x20805x, x20817x, x20818x, x20910x, x20911x}, x20914x);
	defparam lut_735.LUT_SIZE = 7;
	defparam lut_735.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_742 ({sk[136], i_7_, i_8_, i_6_, x260x}, x935x);
	defparam lut_742.LUT_SIZE = 5;
	defparam lut_742.mask = 32'h0f0f4000;

	lut_sub lut_744 ({sk[137], i_9_, i_10_, i_7_, i_8_, i_6_, x910x}, x758x);
	defparam lut_744.LUT_SIZE = 7;
	defparam lut_744.mask = 128'h5555ffff5555ffff0000400000000000;

	lut_sub lut_746 ({sk[138], i_9_, i_10_}, x923x);
	defparam lut_746.LUT_SIZE = 3;
	defparam lut_746.mask = 8'h52;

	lut_sub lut_748 ({sk[139], i_9_, i_10_, x921x, n_n124, n_n283, n_n122}, x3945x);
	defparam lut_748.LUT_SIZE = 7;
	defparam lut_748.mask = 128'h5555ffff5555ffff5f7f000000000000;

	lut_sub lut_752 ({sk[140], i_9_, i_10_, x260x, n_n273, n_n283, x910x}, x20920x);
	defparam lut_752.LUT_SIZE = 7;
	defparam lut_752.mask = 128'h5555ffff5555ffff050f003311110000;

	lut_sub lut_757 ({sk[141], x295x, n_n106, x396x, n_n132, x299x, x251x}, x20924x);
	defparam lut_757.LUT_SIZE = 7;
	defparam lut_757.mask = 128'h5555ffff5555ffff070707ff0f0f0fff;

	lut_sub lut_762 ({sk[142], n_n5231, x20944x, x20945x, x21149x, x24118x}, x21156x);
	defparam lut_762.LUT_SIZE = 6;
	defparam lut_762.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_768 ({sk[143], x21004x, n_n3123, x21002x, x21003x, x21061x}, x21063x);
	defparam lut_768.LUT_SIZE = 6;
	defparam lut_768.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_774 ({sk[144], x21036x, x21037x, x21054x, x21055x}, x21064x);
	defparam lut_774.LUT_SIZE = 5;
	defparam lut_774.mask = 32'h0f0f7fff;

	lut_sub lut_779 ({sk[145], x21122x, x21095x, x21116x, x21117x, n_n3132, n_n3133}, n_n3093);
	defparam lut_779.LUT_SIZE = 7;
	defparam lut_779.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_786 ({sk[146], n_n5, n_n197, x411x, x1926x, x21126x, x21128x}, x21129x);
	defparam lut_786.LUT_SIZE = 7;
	defparam lut_786.mask = 128'h5555ffff5555ffff77ff77ff7fffffff;

	lut_sub lut_792 ({sk[147], x20971x, x20972x, n_n3116, x24198x}, x21130x);
	defparam lut_792.LUT_SIZE = 5;
	defparam lut_792.mask = 32'h0f0fbfff;

	lut_sub lut_797 ({sk[148], n_n4464, n_n4471, x21162x, x21161x, x21173x, x21178x}, x21179x);
	defparam lut_797.LUT_SIZE = 7;
	defparam lut_797.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_804 ({sk[149], n_n3895, x21243x, x21244x, x24116x, x24117x, x24202x}, n_n3890);
	defparam lut_804.LUT_SIZE = 7;
	defparam lut_804.mask = 128'h5555ffff5555fffffeffffffffffffff;

	lut_sub lut_811 ({sk[150], n_n4, n_n3, x21291x, x1461x, x1460x, x21288x}, n_n3896);
	defparam lut_811.LUT_SIZE = 7;
	defparam lut_811.mask = 128'h5555ffff5555ffff55ff5fff77ff7fff;

	lut_sub lut_816 ({sk[151], x21186x, x21264x, n_n3918, n_n3919, n_n3914, n_n3915}, x21292x);
	defparam lut_816.LUT_SIZE = 7;
	defparam lut_816.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_823 ({sk[152], n_n56, n_n2433, x21330x, x21331x, x1848x, x21356x}, x21359x);
	defparam lut_823.LUT_SIZE = 7;
	defparam lut_823.mask = 128'h5555ffff5555ffff5fffffff7fffffff;

	lut_sub lut_829 ({sk[153], n_n57, n_n56, n_n54, x51x, x1245x, x1244x}, x21319x);
	defparam lut_829.LUT_SIZE = 7;
	defparam lut_829.mask = 128'h5555ffff5555ffff000033ff5f5f7fff;

	lut_sub lut_834 ({sk[154], x21312x, x21303x, x24112x, x24113x}, x21320x);
	defparam lut_834.LUT_SIZE = 5;
	defparam lut_834.mask = 32'h0f0fefff;

	lut_sub lut_839 ({sk[155], n_n2434, n_n2436, x21351x}, n_n2428);
	defparam lut_839.LUT_SIZE = 4;
	defparam lut_839.mask = 16'h557f;

	lut_sub lut_843 ({sk[156], n_n271, x909x, n_n2440, x159x, x21361x, x21362x}, x21364x);
	defparam lut_843.LUT_SIZE = 7;
	defparam lut_843.mask = 128'h5555ffff5555ffff55ff55ff55ff7fff;

	lut_sub lut_848 ({sk[157], x21514x, x21470x, x21471x, x21507x, x21508x}, n_n2058);
	defparam lut_848.LUT_SIZE = 6;
	defparam lut_848.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_854 ({sk[158], n_n5, n_n2062, n_n2081, n_n2080, x1487x, x21556x}, x21618x);
	defparam lut_854.LUT_SIZE = 7;
	defparam lut_854.mask = 128'h5555ffff5555ffff5fffffff7fffffff;

	lut_sub lut_860 ({sk[159], x21588x, x21589x, x21613x, n_n2154, x621x, x21611x}, x21619x);
	defparam lut_860.LUT_SIZE = 7;
	defparam lut_860.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_867 ({sk[160], x21396x, x21397x, n_n2061, x21616x}, x21620x);
	defparam lut_867.LUT_SIZE = 5;
	defparam lut_867.mask = 32'h0f0f7fff;

	lut_sub lut_872 ({sk[161], i_14_, i_13_, i_12_, x914x}, n_n148);
	defparam lut_872.LUT_SIZE = 5;
	defparam lut_872.mask = 32'h0f0f4000;

	lut_sub lut_874 ({sk[162], i_14_, i_13_, i_12_, x907x}, n_n106);
	defparam lut_874.LUT_SIZE = 5;
	defparam lut_874.mask = 32'h0f0f4000;

	lut_sub lut_876 ({sk[163], i_1_, i_2_, i_0_, n_n284, n_n273}, n_n126);
	defparam lut_876.LUT_SIZE = 6;
	defparam lut_876.mask = 64'h3f3f3f3f00001000;

	lut_sub lut_878 ({sk[164], i_9_, i_10_, x921x, n_n283, x299x, x251x}, x3242x);
	defparam lut_878.LUT_SIZE = 7;
	defparam lut_878.mask = 128'h5555ffff5555ffff000f000700070007;

	lut_sub lut_882 ({sk[165], i_7_, i_6_, n_n118, n_n284, n_n116, x21630x}, x21631x);
	defparam lut_882.LUT_SIZE = 7;
	defparam lut_882.mask = 128'h5555ffff5555ffff5757575f575f575f;

	lut_sub lut_891 ({sk[166], x21739x, x21740x, x21768x, x21769x, n_n1688, n_n1687}, x21881x);
	defparam lut_891.LUT_SIZE = 7;
	defparam lut_891.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_898 ({sk[167], n_n1685, x21673x, x21674x, n_n1703, n_n1704, x21709x}, n_n1680);
	defparam lut_898.LUT_SIZE = 7;
	defparam lut_898.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_905 ({sk[168], n_n1781, n_n1782, x21856x, n_n1692, x21853x}, x21880x);
	defparam lut_905.LUT_SIZE = 6;
	defparam lut_905.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_911 ({sk[169], n_n1730, n_n1729, x21900x, x21903x}, x21904x);
	defparam lut_911.LUT_SIZE = 5;
	defparam lut_911.mask = 32'h0f0f7fff;

	lut_sub lut_916 ({sk[170], n_n1083, x22324x, x22325x, x22326x, x22327x, x22330x}, x22334x);
	defparam lut_916.LUT_SIZE = 7;
	defparam lut_916.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_923 ({sk[171], x21950x, n_n1089, n_n1157, x21920x, x21928x, x21925x}, x22331x);
	defparam lut_923.LUT_SIZE = 7;
	defparam lut_923.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_930 ({sk[172], n_n342, x22465x, x22466x, n_n345, x22504x, x22505x}, x22588x);
	defparam lut_930.LUT_SIZE = 7;
	defparam lut_930.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_937 ({sk[173], x833x, n_n359, n_n409, n_n360, x22579x}, n_n341);
	defparam lut_937.LUT_SIZE = 6;
	defparam lut_937.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_943 ({sk[174], x22394x, x22421x, x22422x, x22391x, x22392x}, x22583x);
	defparam lut_943.LUT_SIZE = 6;
	defparam lut_943.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_949 ({sk[175], n_n338, n_n381, n_n340, n_n354, x22545x, x22592x}, x24074x);
	defparam lut_949.LUT_SIZE = 7;
	defparam lut_949.mask = 128'h5555ffff5555ffff8000000000000000;

	lut_sub lut_951 ({sk[176], n_n743, n_n742, x22670x, x22671x, n_n739}, x22827x);
	defparam lut_951.LUT_SIZE = 6;
	defparam lut_951.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_957 ({sk[177], x22815x, x22812x, x22813x, x22821x, x24071x}, n_n732);
	defparam lut_957.LUT_SIZE = 6;
	defparam lut_957.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_963 ({sk[178], x22717x, x22744x, x22745x, x22714x, x22715x}, x22826x);
	defparam lut_963.LUT_SIZE = 6;
	defparam lut_963.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_969 ({sk[179], n_n783, n_n781, x22843x, x22846x}, x22847x);
	defparam lut_969.LUT_SIZE = 5;
	defparam lut_969.mask = 32'h0f0f7fff;

	lut_sub lut_974 ({sk[180], n_n5020, n_n5019, x19230x}, n_n5007);
	defparam lut_974.LUT_SIZE = 4;
	defparam lut_974.mask = 16'h557f;

	lut_sub lut_978 ({sk[181], x5959x, x19243x, x5957x, x19250x, x19260x, x19261x}, n_n5005);
	defparam lut_978.LUT_SIZE = 7;
	defparam lut_978.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_985 ({sk[182], n_n5030, x19323x, x5861x, x19331x, x5849x, x19339x}, n_n5004);
	defparam lut_985.LUT_SIZE = 7;
	defparam lut_985.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_992 ({sk[183], n_n5029, x5876x, x19315x, x19349x, x19355x}, x19357x);
	defparam lut_992.LUT_SIZE = 6;
	defparam lut_992.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_998 ({sk[184], x19277x, x19278x, n_n5017, n_n5048, x19303x}, n_n5006);
	defparam lut_998.LUT_SIZE = 6;
	defparam lut_998.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_1004 ({sk[185], i_3_, i_1_, i_2_, i_0_}, x19359x);
	defparam lut_1004.LUT_SIZE = 5;
	defparam lut_1004.mask = 32'h0f0f23a7;

	lut_sub lut_1009 ({sk[186], x915x, n_n261, x160x, x4847x, x1152x, x20053x}, x20054x);
	defparam lut_1009.LUT_SIZE = 7;
	defparam lut_1009.mask = 128'h5555ffff5555ffff5f5f5f5f5f5f7fff;

	lut_sub lut_1014 ({sk[187], n_n2676, x20041x, x20047x, x20048x, x20040x}, x20055x);
	defparam lut_1014.LUT_SIZE = 6;
	defparam lut_1014.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_1020 ({sk[188], n_n100, x20061x, x20062x, x1662x, x20068x, x20073x}, n_n2656);
	defparam lut_1020.LUT_SIZE = 7;
	defparam lut_1020.mask = 128'h5555ffff5555ffff77ffffff7fffffff;

	lut_sub lut_1026 ({sk[189], n_n94, x112x, x877x, n_n2667, x20081x, x24138x}, n_n2657);
	defparam lut_1026.LUT_SIZE = 7;
	defparam lut_1026.mask = 128'h5555ffff5555ffffbfffbfffbfffffff;

	lut_sub lut_1032 ({sk[190], n_n6820, x382x, n_n2713, x493x, n_n2673, x20104x}, n_n2659);
	defparam lut_1032.LUT_SIZE = 7;
	defparam lut_1032.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_1039 ({sk[191], n_n94, n_n6835, x50x, n_n2702, n_n2671, x20111x}, x20113x);
	defparam lut_1039.LUT_SIZE = 7;
	defparam lut_1039.mask = 128'h5555ffff5555ffff7f7fffff7fffffff;

	lut_sub lut_1045 ({sk[192], i_3_, i_1_, i_2_, i_0_}, x20662x);
	defparam lut_1045.LUT_SIZE = 5;
	defparam lut_1045.mask = 32'h0f0f0105;

	lut_sub lut_1048 ({sk[193], i_1_, i_2_, i_0_}, n_n165);
	defparam lut_1048.LUT_SIZE = 4;
	defparam lut_1048.mask = 16'h5508;

	lut_sub lut_1050 ({sk[194], i_14_, i_13_, i_12_, x913x, x911x}, x295x);
	defparam lut_1050.LUT_SIZE = 6;
	defparam lut_1050.mask = 64'h3f3f3f3f50303000;

	lut_sub lut_1054 ({sk[195], i_7_, i_8_, i_6_, n_n165, n_n284}, x396x);
	defparam lut_1054.LUT_SIZE = 6;
	defparam lut_1054.mask = 64'h3f3f3f3f00110000;

	lut_sub lut_1057 ({sk[196], i_7_, i_8_, i_6_, x896x}, n_n132);
	defparam lut_1057.LUT_SIZE = 5;
	defparam lut_1057.mask = 32'h0f0f4000;

	lut_sub lut_1059 ({sk[197], i_14_, i_13_, i_12_, x914x, x912x}, x299x);
	defparam lut_1059.LUT_SIZE = 6;
	defparam lut_1059.mask = 64'h3f3f3f3f50303000;

	lut_sub lut_1063 ({sk[198], i_14_, i_13_, i_12_, x905x, x899x}, x251x);
	defparam lut_1063.LUT_SIZE = 6;
	defparam lut_1063.mask = 64'h3f3f3f3f50303000;

	lut_sub lut_1067 ({sk[199], n_n1, n_n2, n_n3155, x1027x, x1026x, x20941x}, x20944x);
	defparam lut_1067.LUT_SIZE = 7;
	defparam lut_1067.mask = 128'h5555ffff5555ffff55ff77ff5fff7fff;

	lut_sub lut_1072 ({sk[200], x20931x, x20932x, x20936x, x20937x}, x20945x);
	defparam lut_1072.LUT_SIZE = 5;
	defparam lut_1072.mask = 32'h0f0f7fff;

	lut_sub lut_1077 ({sk[201], n_n4, x111x, x21136x, n_n3229, x21147x, x24119x}, x21149x);
	defparam lut_1077.LUT_SIZE = 7;
	defparam lut_1077.mask = 128'h5555ffff5555ffffbfffbfffbfffffff;

	lut_sub lut_1083 ({sk[202], n_n4, n_n3140, n_n3138, x1021x, x21140x, x21151x}, x24118x);
	defparam lut_1083.LUT_SIZE = 7;
	defparam lut_1083.mask = 128'h5555ffff5555ffff8800000080000000;

	lut_sub lut_1086 ({sk[203], x48x, n_n124, x364x, n_n122, x21167x, x21166x}, n_n4464);
	defparam lut_1086.LUT_SIZE = 7;
	defparam lut_1086.mask = 128'h5555ffff5555ffff77ff77ff7fffffff;

	lut_sub lut_1092 ({sk[204], x48x, n_n110, n_n121, n_n111, n_n122, x54x}, n_n4471);
	defparam lut_1092.LUT_SIZE = 7;
	defparam lut_1092.mask = 128'h5555ffff5555ffff135733ff13ff33ff;

	lut_sub lut_1099 ({sk[205], x48x, n_n110, n_n130, n_n111, n_n128, x54x}, x21162x);
	defparam lut_1099.LUT_SIZE = 7;
	defparam lut_1099.mask = 128'h5555ffff5555ffff135733ff13ff33ff;

	lut_sub lut_1106 ({sk[206], x759x, x831x, n_n5682, x4972x, x871x, x886x}, x21161x);
	defparam lut_1106.LUT_SIZE = 7;
	defparam lut_1106.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_1113 ({sk[207], n_n153, x583x, n_n4495, x859x, x261x, x21171x}, x21173x);
	defparam lut_1113.LUT_SIZE = 7;
	defparam lut_1113.mask = 128'h5555ffff5555ffff5fffffff7fffffff;

	lut_sub lut_1119 ({sk[208], x917x, x48x, n_n272, n_n283, n_n111, x24149x}, x21178x);
	defparam lut_1119.LUT_SIZE = 7;
	defparam lut_1119.mask = 128'h5555ffff5555ffffaaaaaaaaabffafff;

	lut_sub lut_1124 ({sk[209], x22063x, x22096x, x22099x, x22100x, x24094x}, n_n1083);
	defparam lut_1124.LUT_SIZE = 6;
	defparam lut_1124.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_1130 ({sk[210], x22177x, n_n1102, x22174x, x22175x}, x22324x);
	defparam lut_1130.LUT_SIZE = 5;
	defparam lut_1130.mask = 32'h0f0f7fff;

	lut_sub lut_1135 ({sk[211], x22229x, x22230x, x22253x, x22254x}, x22325x);
	defparam lut_1135.LUT_SIZE = 5;
	defparam lut_1135.mask = 32'h0f0f7fff;

	lut_sub lut_1140 ({sk[212], n_n1099, x22303x, x22300x, x22301x}, x22326x);
	defparam lut_1140.LUT_SIZE = 5;
	defparam lut_1140.mask = 32'h0f0f7fff;

	lut_sub lut_1145 ({sk[213], n_n1095, x22150x, x22151x, n_n1100}, x22327x);
	defparam lut_1145.LUT_SIZE = 5;
	defparam lut_1145.mask = 32'h0f0f7fff;

	lut_sub lut_1150 ({sk[214], n_n1091, x2825x, x21981x, n_n1115, x21990x, x21991x}, x22330x);
	defparam lut_1150.LUT_SIZE = 7;
	defparam lut_1150.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_1157 ({sk[215], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x917x);
	defparam lut_1157.LUT_SIZE = 7;
	defparam lut_1157.mask = 128'h5555ffff5555ffff0008000000000000;

	lut_sub lut_1159 ({sk[216], i_7_, i_8_, i_6_, x917x}, n_n139);
	defparam lut_1159.LUT_SIZE = 5;
	defparam lut_1159.mask = 32'h0f0f1000;

	lut_sub lut_1161 ({sk[217], i_14_, i_13_, i_12_}, n_n281);
	defparam lut_1161.LUT_SIZE = 4;
	defparam lut_1161.mask = 16'h5580;

	lut_sub lut_1163 ({sk[218], i_9_, i_10_, i_11_, i_15_}, x913x);
	defparam lut_1163.LUT_SIZE = 5;
	defparam lut_1163.mask = 32'h0f0f0800;

	lut_sub lut_1165 ({sk[219], i_14_, i_13_, i_12_, x913x}, n_n151);
	defparam lut_1165.LUT_SIZE = 5;
	defparam lut_1165.mask = 32'h0f0f4000;

	lut_sub lut_1167 ({sk[220], i_7_, i_6_}, n_n155);
	defparam lut_1167.LUT_SIZE = 3;
	defparam lut_1167.mask = 8'h58;

	lut_sub lut_1169 ({sk[221], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x927x);
	defparam lut_1169.LUT_SIZE = 7;
	defparam lut_1169.mask = 128'h5555ffff5555ffff0040000000000000;

	lut_sub lut_1171 ({sk[222], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x918x);
	defparam lut_1171.LUT_SIZE = 7;
	defparam lut_1171.mask = 128'h5555ffff5555ffff0010000000000000;

	lut_sub lut_1173 ({sk[223], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x929x);
	defparam lut_1173.LUT_SIZE = 7;
	defparam lut_1173.mask = 128'h5555ffff5555ffff0000000000400000;

	lut_sub lut_1175 ({sk[224], i_7_, i_6_, x918x, x929x, x261x}, n_n312);
	defparam lut_1175.LUT_SIZE = 6;
	defparam lut_1175.mask = 64'h3f3f3f3f5f5f5f7f;

	lut_sub lut_1185 ({sk[225], i_9_, i_10_}, n_n163);
	defparam lut_1185.LUT_SIZE = 3;
	defparam lut_1185.mask = 8'h58;

	lut_sub lut_1187 ({sk[226], i_7_, i_8_, i_6_, x917x, n_n148, n_n163}, x19365x);
	defparam lut_1187.LUT_SIZE = 7;
	defparam lut_1187.mask = 128'h5555ffff5555ffff0005030300000000;

	lut_sub lut_1191 ({sk[227], i_14_, i_13_, i_12_, x913x, x911x}, x48x);
	defparam lut_1191.LUT_SIZE = 6;
	defparam lut_1191.mask = 64'h3f3f3f3f50003000;

	lut_sub lut_1194 ({sk[228], i_7_, i_8_, i_6_, x917x, x48x}, n_n4476);
	defparam lut_1194.LUT_SIZE = 6;
	defparam lut_1194.mask = 64'h3f3f3f3f10003030;

	lut_sub lut_1197 ({sk[229], i_9_, i_10_, i_11_, i_15_}, x914x);
	defparam lut_1197.LUT_SIZE = 5;
	defparam lut_1197.mask = 32'h0f0f0080;

	lut_sub lut_1199 ({sk[230], i_9_, i_10_, i_11_, i_15_}, x912x);
	defparam lut_1199.LUT_SIZE = 5;
	defparam lut_1199.mask = 32'h0f0f0040;

	lut_sub lut_1201 ({sk[231], i_14_, i_13_, i_12_, x913x, x914x, x912x}, x211x);
	defparam lut_1201.LUT_SIZE = 7;
	defparam lut_1201.mask = 128'h5555ffff5555ffff55000f0033000000;

	lut_sub lut_1205 ({sk[232], i_9_, i_10_, i_11_, i_15_}, x911x);
	defparam lut_1205.LUT_SIZE = 5;
	defparam lut_1205.mask = 32'h0f0f0400;

	lut_sub lut_1207 ({sk[233], i_14_, i_13_, i_12_, x913x}, n_n110);
	defparam lut_1207.LUT_SIZE = 5;
	defparam lut_1207.mask = 32'h0f0f0400;

	lut_sub lut_1209 ({sk[234], i_1_, i_2_, i_0_}, n_n116);
	defparam lut_1209.LUT_SIZE = 4;
	defparam lut_1209.mask = 16'h5540;

	lut_sub lut_1211 ({sk[235], i_7_, i_8_, i_6_, x917x}, n_n142);
	defparam lut_1211.LUT_SIZE = 5;
	defparam lut_1211.mask = 32'h0f0f0400;

	lut_sub lut_1213 ({sk[236], i_7_, i_8_, i_6_, x917x}, n_n136);
	defparam lut_1213.LUT_SIZE = 5;
	defparam lut_1213.mask = 32'h0f0f0100;

	lut_sub lut_1215 ({sk[237], i_7_, i_8_, i_6_, x915x}, n_n255);
	defparam lut_1215.LUT_SIZE = 5;
	defparam lut_1215.mask = 32'h0f0f0010;

	lut_sub lut_1217 ({sk[238], i_7_, i_8_, i_6_, x915x}, n_n241);
	defparam lut_1217.LUT_SIZE = 5;
	defparam lut_1217.mask = 32'h0f0f0001;

	lut_sub lut_1219 ({sk[239], i_14_, i_13_, i_12_, x897x}, n_n103);
	defparam lut_1219.LUT_SIZE = 5;
	defparam lut_1219.mask = 32'h0f0f0010;

	lut_sub lut_1221 ({sk[240], i_14_, i_13_, i_12_, x902x}, n_n31);
	defparam lut_1221.LUT_SIZE = 5;
	defparam lut_1221.mask = 32'h0f0f0010;

	lut_sub lut_1223 ({sk[241], i_14_, i_13_, i_12_, x915x, x898x, n_n261}, x524x);
	defparam lut_1223.LUT_SIZE = 7;
	defparam lut_1223.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_1225 ({sk[242], n_n255, x392x, n_n241, n_n103, n_n31, x524x}, x19380x);
	defparam lut_1225.LUT_SIZE = 7;
	defparam lut_1225.mask = 128'h5555ffff5555ffff555fffff777fffff;

	lut_sub lut_1230 ({sk[243], i_7_, i_8_, i_6_}, n_n273);
	defparam lut_1230.LUT_SIZE = 4;
	defparam lut_1230.mask = 16'h5520;

	lut_sub lut_1232 ({sk[244], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x909x);
	defparam lut_1232.LUT_SIZE = 7;
	defparam lut_1232.mask = 128'h5555ffff5555ffff0000000000800000;

	lut_sub lut_1234 ({sk[245], i_14_, i_13_, i_12_, x906x}, n_n45);
	defparam lut_1234.LUT_SIZE = 5;
	defparam lut_1234.mask = 32'h0f0f0040;

	lut_sub lut_1236 ({sk[246], i_7_, i_8_, i_6_, x909x, n_n200, n_n101}, x372x);
	defparam lut_1236.LUT_SIZE = 7;
	defparam lut_1236.mask = 128'h5555ffff5555ffff0500030000000000;

	lut_sub lut_1239 ({sk[247], i_7_, i_8_, i_6_, x909x, n_n279, x904x}, x875x);
	defparam lut_1239.LUT_SIZE = 7;
	defparam lut_1239.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_1241 ({sk[248], x19380x, n_n273, x909x, n_n45, x372x, x875x}, n_n863);
	defparam lut_1241.LUT_SIZE = 7;
	defparam lut_1241.mask = 128'h5555ffff5555ffff7777777fffffffff;

	lut_sub lut_1246 ({sk[249], x916x, n_n271, n_n59, n_n3418, n_n3417, x597x}, n_n3638);
	defparam lut_1246.LUT_SIZE = 7;
	defparam lut_1246.mask = 128'h5555ffff5555ffff7f7f7f7f7f7f7fff;

	lut_sub lut_1251 ({sk[250], x19390x, x19391x, x19393x, x19396x, x19397x}, x19399x);
	defparam lut_1251.LUT_SIZE = 6;
	defparam lut_1251.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_1257 ({sk[251], n_n208, x916x, n_n3, n_n3408, x1556x, x1555x}, x19420x);
	defparam lut_1257.LUT_SIZE = 7;
	defparam lut_1257.mask = 128'h5555ffff5555ffff0f3f0f3f0f3f5f7f;

	lut_sub lut_1261 ({sk[252], x19405x, x19406x, x19413x, x19414x}, x19421x);
	defparam lut_1261.LUT_SIZE = 5;
	defparam lut_1261.mask = 32'h0f0f7fff;

	lut_sub lut_1266 ({sk[253], n_n1, n_n2, x170x, n_n22, x49x, x46x}, n_n2597);
	defparam lut_1266.LUT_SIZE = 7;
	defparam lut_1266.mask = 128'h5555ffff5555ffff000033ff5f5f7fff;

	lut_sub lut_1271 ({sk[254], x915x, n_n273, n_n283, n_n22, x92x, x1953x}, n_n2598);
	defparam lut_1271.LUT_SIZE = 7;
	defparam lut_1271.mask = 128'h5555ffff5555ffff00000000000f777f;

	lut_sub lut_1275 ({sk[255], n_n1, n_n2, n_n9, x1899x, x70x, x1591x}, x19433x);
	defparam lut_1275.LUT_SIZE = 7;
	defparam lut_1275.mask = 128'h5555ffff5555ffff00005f5f33ff7fff;

	lut_sub lut_1280 ({sk[256], n_n2597, n_n2598, x19433x}, x19435x);
	defparam lut_1280.LUT_SIZE = 4;
	defparam lut_1280.mask = 16'h557f;

	lut_sub lut_1284 ({sk[257], x915x, n_n273, n_n283, x176x, x44x, x1867x}, n_n3424);
	defparam lut_1284.LUT_SIZE = 7;
	defparam lut_1284.mask = 128'h5555ffff5555ffff0000000000553f7f;

	lut_sub lut_1288 ({sk[258], n_n1, n_n2, n_n76, x163x, x207x, x56x}, x812x);
	defparam lut_1288.LUT_SIZE = 7;
	defparam lut_1288.mask = 128'h5555ffff5555ffff000055553fff7fff;

	lut_sub lut_1293 ({sk[259], i_7_, i_8_, i_6_, x915x, x1873x, x1858x}, x19427x);
	defparam lut_1293.LUT_SIZE = 7;
	defparam lut_1293.mask = 128'h5555ffff5555ffff0300050000000000;

	lut_sub lut_1296 ({sk[260], n_n1, n_n2, n_n42, x68x, x45x, x171x}, x19426x);
	defparam lut_1296.LUT_SIZE = 7;
	defparam lut_1296.mask = 128'h5555ffff5555ffff00007f7f00ff7fff;

	lut_sub lut_1301 ({sk[261], n_n1, n_n2, n_n12, n_n76, x209x, x1879x}, x19431x);
	defparam lut_1301.LUT_SIZE = 7;
	defparam lut_1301.mask = 128'h5555ffff5555ffff00005f5f33ff7fff;

	lut_sub lut_1306 ({sk[262], n_n3424, x812x, x19427x, x19426x, x19431x}, x19436x);
	defparam lut_1306.LUT_SIZE = 6;
	defparam lut_1306.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_1312 ({sk[263], n_n1, n_n2, x81x, n_n95, x179x, x98x}, x19440x);
	defparam lut_1312.LUT_SIZE = 7;
	defparam lut_1312.mask = 128'h5555ffff5555ffff000077ff3f3f7fff;

	lut_sub lut_1318 ({sk[264], n_n281, n_n208, x916x, x648x, x908x, x866x}, x19445x);
	defparam lut_1318.LUT_SIZE = 7;
	defparam lut_1318.mask = 128'h5555ffff5555ffff5f5f5f5f5f5f5f7f;

	lut_sub lut_1322 ({sk[265], n_n4, x476x, n_n1356, x5683x, x5682x, x1787x}, x19446x);
	defparam lut_1322.LUT_SIZE = 7;
	defparam lut_1322.mask = 128'h5555ffff5555ffff3fffffff7fffffff;

	lut_sub lut_1328 ({sk[266], x915x, n_n273, n_n283, x81x, n_n42, x43x}, x19438x);
	defparam lut_1328.LUT_SIZE = 7;
	defparam lut_1328.mask = 128'h5555ffff5555ffff0000000000770f7f;

	lut_sub lut_1332 ({sk[267], x915x, n_n273, x204x, x43x, x98x}, x19439x);
	defparam lut_1332.LUT_SIZE = 6;
	defparam lut_1332.mask = 64'h3f3f3f3f0000007f;

	lut_sub lut_1336 ({sk[268], x19440x, x19445x, x19446x, x19438x, x19439x}, x19456x);
	defparam lut_1336.LUT_SIZE = 6;
	defparam lut_1336.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_1342 ({sk[269], i_7_, i_8_, i_6_, x909x, x1799x, x1798x}, n_n3448);
	defparam lut_1342.LUT_SIZE = 7;
	defparam lut_1342.mask = 128'h5555ffff5555ffff0000000005000300;

	lut_sub lut_1345 ({sk[270], n_n4, x166x, n_n94, n_n77, x156x, x257x}, x19467x);
	defparam lut_1345.LUT_SIZE = 7;
	defparam lut_1345.mask = 128'h5555ffff5555ffff007700770f7fffff;

	lut_sub lut_1350 ({sk[271], x909x, x173x, n_n261, n_n263, x539x, x199x}, x19472x);
	defparam lut_1350.LUT_SIZE = 7;
	defparam lut_1350.mask = 128'h5555ffff5555ffff3333333333773fff;

	lut_sub lut_1355 ({sk[272], n_n208, x916x, x374x, n_n30, x466x, x455x}, x19465x);
	defparam lut_1355.LUT_SIZE = 7;
	defparam lut_1355.mask = 128'h5555ffff5555ffff77ff77ff77ff7fff;

	lut_sub lut_1360 ({sk[273], n_n208, x916x, n_n93, n_n6814, x1942x, x471x}, x19466x);
	defparam lut_1360.LUT_SIZE = 7;
	defparam lut_1360.mask = 128'h5555ffff5555ffff5f5f5f5f5f5f7fff;

	lut_sub lut_1365 ({sk[274], n_n6, n_n5, x208x, x165x, n_n59, x167x}, x19471x);
	defparam lut_1365.LUT_SIZE = 7;
	defparam lut_1365.mask = 128'h5555ffff5555ffff00007f7f00ff7fff;

	lut_sub lut_1370 ({sk[275], n_n3448, x19467x, x19472x, x19465x, x19466x, x19471x}, x19481x);
	defparam lut_1370.LUT_SIZE = 7;
	defparam lut_1370.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_1377 ({sk[276], x909x, n_n263, x166x, x389x, x708x}, n_n4773);
	defparam lut_1377.LUT_SIZE = 6;
	defparam lut_1377.mask = 64'h3f3f3f3f7777777f;

	lut_sub lut_1381 ({sk[277], i_7_, i_8_, i_6_, x909x, x224x, x1908x}, n_n4772);
	defparam lut_1381.LUT_SIZE = 7;
	defparam lut_1381.mask = 128'h5555ffff5555ffff0000000005000300;

	lut_sub lut_1384 ({sk[278], i_7_, i_8_, i_6_, x909x, x153x, x1895x}, x19485x);
	defparam lut_1384.LUT_SIZE = 7;
	defparam lut_1384.mask = 128'h5555ffff5555ffff0000000000000700;

	lut_sub lut_1387 ({sk[279], n_n5, x904x, n_n225, x77x, x190x, n_n4770}, x19527x);
	defparam lut_1387.LUT_SIZE = 7;
	defparam lut_1387.mask = 128'h5555ffff5555ffff555555557f7f7fff;

	lut_sub lut_1392 ({sk[280], n_n6, n_n5, x190x, x1554x, x1553x, x1747x}, x24143x);
	defparam lut_1392.LUT_SIZE = 7;
	defparam lut_1392.mask = 128'h5555ffff5555ffffffffcccca0008000;

	lut_sub lut_1397 ({sk[281], n_n4773, n_n4772, x19485x, x19527x, x24143x}, x19530x);
	defparam lut_1397.LUT_SIZE = 6;
	defparam lut_1397.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_1403 ({sk[282], n_n48, n_n53, x1280x, x1559x, x19509x, x19513x}, x832x);
	defparam lut_1403.LUT_SIZE = 7;
	defparam lut_1403.mask = 128'h5555ffff5555ffff777777ff7f7f7fff;

	lut_sub lut_1408 ({sk[283], n_n53, n_n76, n_n6858, x478x, x1948x, x19503x}, x19504x);
	defparam lut_1408.LUT_SIZE = 7;
	defparam lut_1408.mask = 128'h5555ffff5555ffff5fff5fff7fffffff;

	lut_sub lut_1414 ({sk[284], n_n4774, x19489x, x19490x, x5607x, x19495x}, x19505x);
	defparam lut_1414.LUT_SIZE = 6;
	defparam lut_1414.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_1420 ({sk[285], n_n48, n_n95, x473x, x298x, x19520x, x19519x}, x19523x);
	defparam lut_1420.LUT_SIZE = 7;
	defparam lut_1420.mask = 128'h5555ffff5555ffff7fff7fff7fffffff;

	lut_sub lut_1426 ({sk[286], i_7_, i_8_, i_6_, x909x}, n_n56);
	defparam lut_1426.LUT_SIZE = 5;
	defparam lut_1426.mask = 32'h0f0f0010;

	lut_sub lut_1428 ({sk[287], i_14_, i_13_, i_12_, x908x, x902x}, x163x);
	defparam lut_1428.LUT_SIZE = 6;
	defparam lut_1428.mask = 64'h3f3f3f3f05053000;

	lut_sub lut_1432 ({sk[288], i_14_, i_13_, i_12_, i_15_, x908x, n_n270}, x207x);
	defparam lut_1432.LUT_SIZE = 7;
	defparam lut_1432.mask = 128'h5555ffff5555ffff0533005000000000;

	lut_sub lut_1436 ({sk[289], n_n271, n_n220, x909x, x904x, x204x}, x788x);
	defparam lut_1436.LUT_SIZE = 6;
	defparam lut_1436.mask = 64'h3f3f3f3f00000507;

	lut_sub lut_1439 ({sk[290], n_n57, n_n56, x170x, n_n22, x49x, x46x}, n_n3708);
	defparam lut_1439.LUT_SIZE = 7;
	defparam lut_1439.mask = 128'h5555ffff5555ffff000033ff5f5f7fff;

	lut_sub lut_1444 ({sk[291], n_n57, n_n56, n_n76, x1861x, x70x, x1761x}, x24160x);
	defparam lut_1444.LUT_SIZE = 7;
	defparam lut_1444.mask = 128'h5555ffff5555ffffffffaa00c0c08000;

	lut_sub lut_1449 ({sk[292], n_n56, x163x, x207x, x788x, n_n3708, x24160x}, x19546x);
	defparam lut_1449.LUT_SIZE = 7;
	defparam lut_1449.mask = 128'h5555ffff5555ffffbfbfbfbfbfffffff;

	lut_sub lut_1455 ({sk[293], i_7_, i_8_, i_6_, x909x, x176x, x465x}, n_n4781);
	defparam lut_1455.LUT_SIZE = 7;
	defparam lut_1455.mask = 128'h5555ffff5555ffff5555555555555557;

	lut_sub lut_1458 ({sk[294], i_7_, i_8_, i_6_, x909x, x179x, n_n4677}, x19533x);
	defparam lut_1458.LUT_SIZE = 7;
	defparam lut_1458.mask = 128'h5555ffff5555ffff5555555555555557;

	lut_sub lut_1461 ({sk[295], n_n57, n_n56, x45x, x43x, x171x, x98x}, x19534x);
	defparam lut_1461.LUT_SIZE = 7;
	defparam lut_1461.mask = 128'h5555ffff5555ffff000033ff5f5f7fff;

	lut_sub lut_1466 ({sk[296], i_7_, i_8_, i_6_, x909x, n_n22, x1441x}, n_n3709);
	defparam lut_1466.LUT_SIZE = 7;
	defparam lut_1466.mask = 128'h5555ffff5555ffff0000000000030005;

	lut_sub lut_1469 ({sk[297], n_n57, n_n56, n_n76, x163x, x207x, x56x}, n_n3711);
	defparam lut_1469.LUT_SIZE = 7;
	defparam lut_1469.mask = 128'h5555ffff5555ffff000055553fff7fff;

	lut_sub lut_1474 ({sk[298], n_n4781, x19533x, x19534x, n_n3709, n_n3711}, x19547x);
	defparam lut_1474.LUT_SIZE = 6;
	defparam lut_1474.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_1480 ({sk[299], i_7_, i_8_, i_6_, x915x}, n_n100);
	defparam lut_1480.LUT_SIZE = 5;
	defparam lut_1480.mask = 32'h0f0f0004;

	lut_sub lut_1482 ({sk[300], i_7_, i_8_, i_6_, x915x}, n_n94);
	defparam lut_1482.LUT_SIZE = 5;
	defparam lut_1482.mask = 32'h0f0f0040;

	lut_sub lut_1484 ({sk[301], i_14_, i_13_, i_12_, i_15_, n_n270}, x181x);
	defparam lut_1484.LUT_SIZE = 6;
	defparam lut_1484.mask = 64'h3f3f3f3f11040000;

	lut_sub lut_1488 ({sk[302], i_14_, i_13_, i_12_, x915x, n_n261, x908x}, x5529x);
	defparam lut_1488.LUT_SIZE = 7;
	defparam lut_1488.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_1491 ({sk[303], i_14_, i_13_, i_12_, i_15_, n_n275, x903x}, x1800x);
	defparam lut_1491.LUT_SIZE = 7;
	defparam lut_1491.mask = 128'h5555ffff5555ffff0055555503000330;

	lut_sub lut_1498 ({sk[304], n_n103, n_n100, n_n94, x181x, x5529x, x1800x}, x19554x);
	defparam lut_1498.LUT_SIZE = 7;
	defparam lut_1498.mask = 128'h5555ffff5555ffff33773f7f33ff3fff;

	lut_sub lut_1503 ({sk[305], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x915x);
	defparam lut_1503.LUT_SIZE = 7;
	defparam lut_1503.mask = 128'h5555ffff5555ffff0080000000000000;

	lut_sub lut_1505 ({sk[306], i_7_, i_8_, i_6_}, n_n261);
	defparam lut_1505.LUT_SIZE = 4;
	defparam lut_1505.mask = 16'h5502;

	lut_sub lut_1507 ({sk[307], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x91x);
	defparam lut_1507.LUT_SIZE = 7;
	defparam lut_1507.mask = 128'h5555ffff5555ffff0000000001000104;

	lut_sub lut_1511 ({sk[308], i_9_, i_10_, i_11_, i_15_, n_n258, x44x}, x121x);
	defparam lut_1511.LUT_SIZE = 7;
	defparam lut_1511.mask = 128'h5555ffff5555ffff5555555555555575;

	lut_sub lut_1514 ({sk[309], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1903x);
	defparam lut_1514.LUT_SIZE = 7;
	defparam lut_1514.mask = 128'h5555ffff5555ffff0101000504000400;

	lut_sub lut_1521 ({sk[310], x40x, n_n100, n_n94, x1860x, n_n15, x1801x}, x19572x);
	defparam lut_1521.LUT_SIZE = 7;
	defparam lut_1521.mask = 128'h5555ffff5555ffff005f337f005fffff;

	lut_sub lut_1526 ({sk[311], x915x, n_n261, x91x, x121x, x1903x, x19572x}, x19573x);
	defparam lut_1526.LUT_SIZE = 7;
	defparam lut_1526.mask = 128'h5555ffff5555ffff5555555555557fff;

	lut_sub lut_1531 ({sk[312], n_n281, x146x, x908x, n_n100, n_n59, x156x}, x19560x);
	defparam lut_1531.LUT_SIZE = 7;
	defparam lut_1531.mask = 128'h5555ffff5555ffff07070f0f070f0f0f;

	lut_sub lut_1536 ({sk[313], x146x, n_n94, x121x, x137x, n_n3481, x132x}, x19561x);
	defparam lut_1536.LUT_SIZE = 7;
	defparam lut_1536.mask = 128'h5555ffff5555ffff33337fff3333ffff;

	lut_sub lut_1542 ({sk[314], n_n266, n_n271, x909x, x81x, n_n95, x98x}, x19564x);
	defparam lut_1542.LUT_SIZE = 7;
	defparam lut_1542.mask = 128'h5555ffff5555ffff0000005f0033007f;

	lut_sub lut_1546 ({sk[315], n_n57, n_n56, x204x, x179x, n_n4681, x43x}, x19565x);
	defparam lut_1546.LUT_SIZE = 7;
	defparam lut_1546.mask = 128'h5555ffff5555ffff33337f7f33ff7fff;

	lut_sub lut_1551 ({sk[316], n_n281, x915x, n_n263, x908x, x370x}, x19566x);
	defparam lut_1551.LUT_SIZE = 6;
	defparam lut_1551.mask = 64'h3f3f3f3f55555557;

	lut_sub lut_1554 ({sk[317], x19560x, x19561x, x19564x, x19565x, x19566x}, x19574x);
	defparam lut_1554.LUT_SIZE = 6;
	defparam lut_1554.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_1560 ({sk[318], i_14_, i_13_, i_12_, i_15_, n_n267}, x94x);
	defparam lut_1560.LUT_SIZE = 6;
	defparam lut_1560.mask = 64'h3f3f3f3f00014040;

	lut_sub lut_1564 ({sk[319], i_14_, i_13_, i_12_, x904x}, x77x);
	defparam lut_1564.LUT_SIZE = 5;
	defparam lut_1564.mask = 32'h0f0f1400;

	lut_sub lut_1567 ({sk[320], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1321x);
	defparam lut_1567.LUT_SIZE = 7;
	defparam lut_1567.mask = 128'h5555ffff5555ffff0101000505000504;

	lut_sub lut_1577 ({sk[321], i_14_, i_13_, i_12_, i_15_, x900x, n_n267}, x1934x);
	defparam lut_1577.LUT_SIZE = 7;
	defparam lut_1577.mask = 128'h5555ffff5555ffff0000000005330550;

	lut_sub lut_1582 ({sk[322], n_n100, x94x, n_n94, x77x, x1321x, x1934x}, x19586x);
	defparam lut_1582.LUT_SIZE = 7;
	defparam lut_1582.mask = 128'h5555ffff5555ffff005500ff3f7f3fff;

	lut_sub lut_1587 ({sk[323], x51x, n_n105, n_n100, x94x, x599x, x138x}, x19582x);
	defparam lut_1587.LUT_SIZE = 7;
	defparam lut_1587.mask = 128'h5555ffff5555ffff337f33ff33ff33ff;

	lut_sub lut_1593 ({sk[324], x915x, n_n261, n_n263, x108x, x1943x, x1369x}, x19583x);
	defparam lut_1593.LUT_SIZE = 7;
	defparam lut_1593.mask = 128'h5555ffff5555ffff0000000000770f7f;

	lut_sub lut_1597 ({sk[325], x19586x, x19582x, x19583x}, x811x);
	defparam lut_1597.LUT_SIZE = 4;
	defparam lut_1597.mask = 16'h557f;

	lut_sub lut_1601 ({sk[326], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x921x);
	defparam lut_1601.LUT_SIZE = 7;
	defparam lut_1601.mask = 128'h5555ffff5555ffff0800000000000000;

	lut_sub lut_1603 ({sk[327], i_5_, i_3_, i_4_}, n_n284);
	defparam lut_1603.LUT_SIZE = 4;
	defparam lut_1603.mask = 16'h5580;

	lut_sub lut_1605 ({sk[328], i_7_, i_8_, i_6_, n_n165, n_n284}, n_n124);
	defparam lut_1605.LUT_SIZE = 6;
	defparam lut_1605.mask = 64'h3f3f3f3f01000000;

	lut_sub lut_1607 ({sk[329], i_7_, i_8_, i_6_}, n_n208);
	defparam lut_1607.LUT_SIZE = 4;
	defparam lut_1607.mask = 16'h5510;

	lut_sub lut_1609 ({sk[330], i_7_, i_6_}, x289x);
	defparam lut_1609.LUT_SIZE = 3;
	defparam lut_1609.mask = 8'h57;

	lut_sub lut_1613 ({sk[331], i_7_, i_6_, i_1_, i_2_, i_0_, n_n284}, x364x);
	defparam lut_1613.LUT_SIZE = 7;
	defparam lut_1613.mask = 128'h5555ffff5555ffff0000000000000040;

	lut_sub lut_1615 ({sk[332], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, n_n5671);
	defparam lut_1615.LUT_SIZE = 7;
	defparam lut_1615.mask = 128'h5555ffff5555ffff0000000000000040;

	lut_sub lut_1617 ({sk[333], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, n_n5672);
	defparam lut_1617.LUT_SIZE = 7;
	defparam lut_1617.mask = 128'h5555ffff5555ffff0000000000004000;

	lut_sub lut_1619 ({sk[334], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, n_n5674);
	defparam lut_1619.LUT_SIZE = 7;
	defparam lut_1619.mask = 128'h5555ffff5555ffff0000400000000000;

	lut_sub lut_1621 ({sk[335], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, n_n5673);
	defparam lut_1621.LUT_SIZE = 7;
	defparam lut_1621.mask = 128'h5555ffff5555ffff0000004000000000;

	lut_sub lut_1623 ({sk[336], i_14_, i_13_, i_12_}, n_n220);
	defparam lut_1623.LUT_SIZE = 4;
	defparam lut_1623.mask = 16'h5520;

	lut_sub lut_1625 ({sk[337], i_9_, i_10_, i_11_, i_15_}, x905x);
	defparam lut_1625.LUT_SIZE = 5;
	defparam lut_1625.mask = 32'h0f0f0008;

	lut_sub lut_1627 ({sk[338], i_14_, i_13_, i_12_, x905x, x899x}, x103x);
	defparam lut_1627.LUT_SIZE = 6;
	defparam lut_1627.mask = 64'h3f3f3f3f50003000;

	lut_sub lut_1630 ({sk[339], i_14_, i_13_, i_12_, x914x, x912x}, x54x);
	defparam lut_1630.LUT_SIZE = 6;
	defparam lut_1630.mask = 64'h3f3f3f3f50003000;

	lut_sub lut_1633 ({sk[340], n_n124, n_n220, x914x, x905x, x103x, x54x}, x819x);
	defparam lut_1633.LUT_SIZE = 7;
	defparam lut_1633.mask = 128'h5555ffff5555ffff0000000077777fff;

	lut_sub lut_1638 ({sk[341], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x919x);
	defparam lut_1638.LUT_SIZE = 7;
	defparam lut_1638.mask = 128'h5555ffff5555ffff0000000010000000;

	lut_sub lut_1640 ({sk[342], i_1_, i_2_, i_0_}, n_n118);
	defparam lut_1640.LUT_SIZE = 4;
	defparam lut_1640.mask = 16'h5510;

	lut_sub lut_1642 ({sk[343], i_9_, i_10_, i_11_, i_15_}, x907x);
	defparam lut_1642.LUT_SIZE = 5;
	defparam lut_1642.mask = 32'h0f0f8000;

	lut_sub lut_1644 ({sk[344], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x936x);
	defparam lut_1644.LUT_SIZE = 7;
	defparam lut_1644.mask = 128'h5555ffff5555ffff4000000000000000;

	lut_sub lut_1646 ({sk[345], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, n_n5678);
	defparam lut_1646.LUT_SIZE = 7;
	defparam lut_1646.mask = 128'h5555ffff5555ffff4000000000000000;

	lut_sub lut_1648 ({sk[346], i_7_, i_8_, i_6_}, n_n283);
	defparam lut_1648.LUT_SIZE = 4;
	defparam lut_1648.mask = 16'h5580;

	lut_sub lut_1650 ({sk[347], i_14_, i_13_, i_12_, x899x}, n_n107);
	defparam lut_1650.LUT_SIZE = 5;
	defparam lut_1650.mask = 32'h0f0f4000;

	lut_sub lut_1652 ({sk[348], i_14_, i_13_, i_12_, x905x}, x250x);
	defparam lut_1652.LUT_SIZE = 5;
	defparam lut_1652.mask = 32'h0f0f0440;

	lut_sub lut_1655 ({sk[349], i_14_, i_13_, i_12_, x913x, x912x}, x283x);
	defparam lut_1655.LUT_SIZE = 6;
	defparam lut_1655.mask = 64'h3f3f3f3f50303000;

	lut_sub lut_1659 ({sk[350], i_9_, i_10_, n_n133, n_n220, x914x, n_n279}, x19607x);
	defparam lut_1659.LUT_SIZE = 7;
	defparam lut_1659.mask = 128'h5555ffff5555ffffffff13ff13ff13ff;

	lut_sub lut_1664 ({sk[351], i_7_, i_6_, i_1_, i_2_, i_0_, n_n284}, n_n5769);
	defparam lut_1664.LUT_SIZE = 7;
	defparam lut_1664.mask = 128'h5555ffff5555ffff0000000000400000;

	lut_sub lut_1666 ({sk[352], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, x582x);
	defparam lut_1666.LUT_SIZE = 7;
	defparam lut_1666.mask = 128'h5555ffff5555ffff0040404040404000;

	lut_sub lut_1673 ({sk[353], i_9_, i_10_, i_11_, i_15_, n_n220}, x266x);
	defparam lut_1673.LUT_SIZE = 6;
	defparam lut_1673.mask = 64'h3f3f3f3fff000040;

	lut_sub lut_1676 ({sk[354], i_9_, i_10_, i_11_, i_15_}, x899x);
	defparam lut_1676.LUT_SIZE = 5;
	defparam lut_1676.mask = 32'h0f0f0004;

	lut_sub lut_1678 ({sk[355], i_14_, i_13_, i_12_, x914x, x905x, x899x}, x294x);
	defparam lut_1678.LUT_SIZE = 7;
	defparam lut_1678.mask = 128'h5555ffff5555ffff55000f0033000000;

	lut_sub lut_1682 ({sk[356], i_7_, i_6_}, n_n272);
	defparam lut_1682.LUT_SIZE = 3;
	defparam lut_1682.mask = 8'h52;

	lut_sub lut_1684 ({sk[357], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x924x);
	defparam lut_1684.LUT_SIZE = 7;
	defparam lut_1684.mask = 128'h5555ffff5555ffff0000000000000008;

	lut_sub lut_1686 ({sk[358], i_14_, i_13_, i_12_, n_n130, x914x}, x831x);
	defparam lut_1686.LUT_SIZE = 6;
	defparam lut_1686.mask = 64'h3f3f3f3f00100000;

	lut_sub lut_1688 ({sk[359], i_9_, i_10_, i_7_, i_8_, i_6_, x260x}, n_n5693);
	defparam lut_1688.LUT_SIZE = 7;
	defparam lut_1688.mask = 128'h5555ffff5555ffff0400000000000000;

	lut_sub lut_1690 ({sk[360], i_9_, i_10_, i_7_, i_8_, i_6_, x910x}, x318x);
	defparam lut_1690.LUT_SIZE = 7;
	defparam lut_1690.mask = 128'h5555ffff5555ffff0400000040000000;

	lut_sub lut_1693 ({sk[361], i_7_, i_6_, x924x, x831x, n_n5693, x318x}, x19627x);
	defparam lut_1693.LUT_SIZE = 7;
	defparam lut_1693.mask = 128'h5555ffff5555ffff7f7f7f7f7f7f7fff;

	lut_sub lut_1698 ({sk[362], i_7_, i_8_, i_6_}, n_n271);
	defparam lut_1698.LUT_SIZE = 4;
	defparam lut_1698.mask = 16'h5504;

	lut_sub lut_1700 ({sk[363], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x896x);
	defparam lut_1700.LUT_SIZE = 7;
	defparam lut_1700.mask = 128'h5555ffff5555ffff0000000000080000;

	lut_sub lut_1702 ({sk[364], i_9_, i_10_, n_n220, n_n128, x935x, x914x}, x609x);
	defparam lut_1702.LUT_SIZE = 7;
	defparam lut_1702.mask = 128'h5555ffff5555ffff0005000533370005;

	lut_sub lut_1705 ({sk[365], i_1_, i_2_, i_0_, n_n284, n_n283}, n_n127);
	defparam lut_1705.LUT_SIZE = 6;
	defparam lut_1705.mask = 64'h3f3f3f3f00001000;

	lut_sub lut_1707 ({sk[366], i_14_, i_13_, i_12_, x914x}, n_n111);
	defparam lut_1707.LUT_SIZE = 5;
	defparam lut_1707.mask = 32'h0f0f0400;

	lut_sub lut_1709 ({sk[367], i_7_, i_8_, i_6_, x896x}, n_n130);
	defparam lut_1709.LUT_SIZE = 5;
	defparam lut_1709.mask = 32'h0f0f1000;

	lut_sub lut_1711 ({sk[368], i_1_, i_2_, i_0_, n_n264, n_n271}, n_n121);
	defparam lut_1711.LUT_SIZE = 6;
	defparam lut_1711.mask = 64'h3f3f3f3f00001000;

	lut_sub lut_1713 ({sk[369], i_7_, i_8_, i_6_, n_n165, n_n264}, n_n122);
	defparam lut_1713.LUT_SIZE = 6;
	defparam lut_1713.mask = 64'h3f3f3f3f01000000;

	lut_sub lut_1715 ({sk[370], i_7_, i_6_, n_n152, x924x, n_n111, x54x}, x19639x);
	defparam lut_1715.LUT_SIZE = 7;
	defparam lut_1715.mask = 128'h5555ffff5555ffff00770f7f0f7f0077;

	lut_sub lut_1720 ({sk[371], i_7_, i_6_}, x116x);
	defparam lut_1720.LUT_SIZE = 3;
	defparam lut_1720.mask = 8'h53;

	lut_sub lut_1723 ({sk[372], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x920x);
	defparam lut_1723.LUT_SIZE = 7;
	defparam lut_1723.mask = 128'h5555ffff5555ffff1000000000000000;

	lut_sub lut_1725 ({sk[373], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x111x);
	defparam lut_1725.LUT_SIZE = 7;
	defparam lut_1725.mask = 128'h5555ffff5555ffff0000000010004040;

	lut_sub lut_1729 ({sk[374], i_14_, i_13_, i_12_, x903x, x897x}, x92x);
	defparam lut_1729.LUT_SIZE = 6;
	defparam lut_1729.mask = 64'h3f3f3f3f05053000;

	lut_sub lut_1733 ({sk[375], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x147x);
	defparam lut_1733.LUT_SIZE = 7;
	defparam lut_1733.mask = 128'h5555ffff5555ffff0000000001000404;

	lut_sub lut_1737 ({sk[376], i_14_, i_13_, i_12_, x903x, x897x}, x46x);
	defparam lut_1737.LUT_SIZE = 6;
	defparam lut_1737.mask = 64'h3f3f3f3f53030000;

	lut_sub lut_1741 ({sk[377], x909x, n_n261, x111x, x92x, x147x, x46x}, x19659x);
	defparam lut_1741.LUT_SIZE = 7;
	defparam lut_1741.mask = 128'h5555ffff5555ffff0000000000007fff;

	lut_sub lut_1746 ({sk[378], i_7_, i_8_, i_6_, x909x}, n_n5);
	defparam lut_1746.LUT_SIZE = 5;
	defparam lut_1746.mask = 32'h0f0f0040;

	lut_sub lut_1748 ({sk[379], i_14_, i_13_, i_12_, x908x}, n_n76);
	defparam lut_1748.LUT_SIZE = 5;
	defparam lut_1748.mask = 32'h0f0f0400;

	lut_sub lut_1750 ({sk[380], i_14_, i_13_, i_12_, x902x}, x49x);
	defparam lut_1750.LUT_SIZE = 5;
	defparam lut_1750.mask = 32'h0f0f0014;

	lut_sub lut_1753 ({sk[381], i_7_, i_8_, i_6_, n_n220, x909x, x903x}, x5388x);
	defparam lut_1753.LUT_SIZE = 7;
	defparam lut_1753.mask = 128'h5555ffff5555ffff0000000000000100;

	lut_sub lut_1755 ({sk[382], i_7_, i_8_, i_6_, x909x, x82x}, x5385x);
	defparam lut_1755.LUT_SIZE = 6;
	defparam lut_1755.mask = 64'h3f3f3f3f00000010;

	lut_sub lut_1757 ({sk[383], i_14_, i_13_, i_12_, i_15_, x908x, n_n270}, x1017x);
	defparam lut_1757.LUT_SIZE = 7;
	defparam lut_1757.mask = 128'h5555ffff5555ffff0537005555005050;

	lut_sub lut_1767 ({sk[384], n_n5, n_n76, x49x, x5388x, x5385x, x1017x}, x19660x);
	defparam lut_1767.LUT_SIZE = 7;
	defparam lut_1767.mask = 128'h5555ffff5555ffff3f3f3f3f7fffffff;

	lut_sub lut_1773 ({sk[385], i_7_, i_8_, i_6_, x909x}, n_n6);
	defparam lut_1773.LUT_SIZE = 5;
	defparam lut_1773.mask = 32'h0f0f0004;

	lut_sub lut_1775 ({sk[386], i_14_, i_13_, i_12_, i_15_, n_n247, n_n137}, x1082x);
	defparam lut_1775.LUT_SIZE = 7;
	defparam lut_1775.mask = 128'h5555ffff5555ffff5353507373535370;

	lut_sub lut_1786 ({sk[387], i_14_, i_13_, i_12_, i_15_, n_n253, x45x}, x1081x);
	defparam lut_1786.LUT_SIZE = 7;
	defparam lut_1786.mask = 128'h5555ffff5555ffff5775757555555555;

	lut_sub lut_1792 ({sk[388], n_n6, n_n5, n_n111, n_n6582, x1894x, x85x}, x19665x);
	defparam lut_1792.LUT_SIZE = 7;
	defparam lut_1792.mask = 128'h5555ffff5555ffff0f0f7f7f0fff7fff;

	lut_sub lut_1797 ({sk[389], i_14_, i_13_, i_12_, i_15_, n_n253, n_n267}, x1087x);
	defparam lut_1797.LUT_SIZE = 7;
	defparam lut_1797.mask = 128'h5555ffff5555ffff0555005557037370;

	lut_sub lut_1812 ({sk[390], n_n6, n_n5, x1082x, x1081x, x19665x, x1087x}, x19677x);
	defparam lut_1812.LUT_SIZE = 7;
	defparam lut_1812.mask = 128'h5555ffff5555ffff33337f7f33ff7fff;

	lut_sub lut_1817 ({sk[391], n_n271, x909x, n_n261, x632x, x171x, x1273x}, n_n4330);
	defparam lut_1817.LUT_SIZE = 7;
	defparam lut_1817.mask = 128'h5555ffff5555ffff0f0f0f3f0f0f5f7f;

	lut_sub lut_1821 ({sk[392], n_n266, x909x, n_n261, x45x, x1085x, x71x}, x19672x);
	defparam lut_1821.LUT_SIZE = 7;
	defparam lut_1821.mask = 128'h5555ffff5555ffff0000005f0000337f;

	lut_sub lut_1825 ({sk[393], n_n271, x909x, x225x, x130x, x19670x}, x19671x);
	defparam lut_1825.LUT_SIZE = 6;
	defparam lut_1825.mask = 64'h3f3f3f3f5555557f;

	lut_sub lut_1829 ({sk[394], x909x, n_n261, n_n263, x81x, n_n42, x1088x}, x19676x);
	defparam lut_1829.LUT_SIZE = 7;
	defparam lut_1829.mask = 128'h5555ffff5555ffff0000000000337f7f;

	lut_sub lut_1834 ({sk[395], n_n4330, x19672x, x19671x, x19676x}, x19678x);
	defparam lut_1834.LUT_SIZE = 5;
	defparam lut_1834.mask = 32'h0f0f7fff;

	lut_sub lut_1839 ({sk[396], i_9_, i_10_}, n_n274);
	defparam lut_1839.LUT_SIZE = 3;
	defparam lut_1839.mask = 8'h54;

	lut_sub lut_1841 ({sk[397], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x183x);
	defparam lut_1841.LUT_SIZE = 7;
	defparam lut_1841.mask = 128'h5555ffff5555ffff0000100000400010;

	lut_sub lut_1845 ({sk[398], i_7_, i_8_, i_6_, x183x, x909x}, n_n4807);
	defparam lut_1845.LUT_SIZE = 6;
	defparam lut_1845.mask = 64'h3f3f3f3f00000010;

	lut_sub lut_1847 ({sk[399], i_14_, i_13_, i_12_, x908x}, n_n60);
	defparam lut_1847.LUT_SIZE = 5;
	defparam lut_1847.mask = 32'h0f0f4000;

	lut_sub lut_1849 ({sk[400], i_14_, i_13_, i_12_, x905x, x899x}, x118x);
	defparam lut_1849.LUT_SIZE = 6;
	defparam lut_1849.mask = 64'h3f3f3f3f00000305;

	lut_sub lut_1852 ({sk[401], i_7_, i_8_, i_6_, x909x, n_n60, x118x}, x541x);
	defparam lut_1852.LUT_SIZE = 7;
	defparam lut_1852.mask = 128'h5555ffff5555ffff0000000003000500;

	lut_sub lut_1855 ({sk[402], i_14_, i_13_, i_12_, x913x, x911x}, x218x);
	defparam lut_1855.LUT_SIZE = 6;
	defparam lut_1855.mask = 64'h3f3f3f3f30500300;

	lut_sub lut_1859 ({sk[403], i_14_, i_13_, i_12_, x905x, x899x}, x72x);
	defparam lut_1859.LUT_SIZE = 6;
	defparam lut_1859.mask = 64'h3f3f3f3f30500000;

	lut_sub lut_1862 ({sk[404], i_14_, i_13_, i_12_, x911x}, n_n206);
	defparam lut_1862.LUT_SIZE = 5;
	defparam lut_1862.mask = 32'h0f0f0001;

	lut_sub lut_1864 ({sk[405], n_n6, x541x, n_n5, x218x, x72x, n_n206}, n_n4223);
	defparam lut_1864.LUT_SIZE = 7;
	defparam lut_1864.mask = 128'h5555ffff5555ffff005fffff337fffff;

	lut_sub lut_1869 ({sk[406], i_14_, i_13_, i_12_, x902x, x63x}, x146x);
	defparam lut_1869.LUT_SIZE = 6;
	defparam lut_1869.mask = 64'h3f3f3f3f55555557;

	lut_sub lut_1872 ({sk[407], i_14_, i_13_, i_12_, x897x}, n_n59);
	defparam lut_1872.LUT_SIZE = 5;
	defparam lut_1872.mask = 32'h0f0f0001;

	lut_sub lut_1874 ({sk[408], i_14_, i_13_, i_12_, x903x, x897x}, x156x);
	defparam lut_1874.LUT_SIZE = 6;
	defparam lut_1874.mask = 64'h3f3f3f3f30500300;

	lut_sub lut_1878 ({sk[409], i_14_, i_13_, i_12_, x903x, x897x}, x132x);
	defparam lut_1878.LUT_SIZE = 6;
	defparam lut_1878.mask = 64'h3f3f3f3f30500000;

	lut_sub lut_1881 ({sk[410], n_n6, n_n5, x146x, n_n59, x156x, x132x}, n_n4224);
	defparam lut_1881.LUT_SIZE = 7;
	defparam lut_1881.mask = 128'h5555ffff5555ffff000055ff3f3f7fff;

	lut_sub lut_1886 ({sk[411], n_n57, n_n56, n_n4959, x166x, x180x, x254x}, x19723x);
	defparam lut_1886.LUT_SIZE = 7;
	defparam lut_1886.mask = 128'h5555ffff5555ffff00ff55ff3fff7fff;

	lut_sub lut_1891 ({sk[412], n_n57, x219x, x189x, n_n4955, n_n4956, x5288x}, x19724x);
	defparam lut_1891.LUT_SIZE = 7;
	defparam lut_1891.mask = 128'h5555ffff5555ffff7f7f7f7f7fffffff;

	lut_sub lut_1897 ({sk[413], n_n266, x909x, n_n4948, n_n4952, x157x, x5284x}, x19727x);
	defparam lut_1897.LUT_SIZE = 7;
	defparam lut_1897.mask = 128'h5555ffff5555ffff5fff5fff5fff7fff;

	lut_sub lut_1902 ({sk[414], n_n57, x200x, x277x, n_n4950, n_n4947, x112x}, x19728x);
	defparam lut_1902.LUT_SIZE = 7;
	defparam lut_1902.mask = 128'h5555ffff5555ffff3f3f3f3f7fffffff;

	lut_sub lut_1908 ({sk[415], n_n57, n_n56, n_n4970, x166x, x99x, x41x}, x19732x);
	defparam lut_1908.LUT_SIZE = 7;
	defparam lut_1908.mask = 128'h5555ffff5555ffff00ff0fff77ff7fff;

	lut_sub lut_1913 ({sk[416], n_n57, n_n56, x153x, x180x, x224x, n_n4967}, x19733x);
	defparam lut_1913.LUT_SIZE = 7;
	defparam lut_1913.mask = 128'h5555ffff5555ffff55557fff77777fff;

	lut_sub lut_1919 ({sk[417], i_7_, i_8_, i_6_}, n_n263);
	defparam lut_1919.LUT_SIZE = 4;
	defparam lut_1919.mask = 16'h5508;

	lut_sub lut_1921 ({sk[418], n_n151, x909x, n_n261, n_n263, x72x, x118x}, x390x);
	defparam lut_1921.LUT_SIZE = 7;
	defparam lut_1921.mask = 128'h5555ffff5555ffff00000707000007ff;

	lut_sub lut_1925 ({sk[419], i_14_, i_13_, i_12_, i_15_, x900x, n_n267}, x176x);
	defparam lut_1925.LUT_SIZE = 7;
	defparam lut_1925.mask = 128'h5555ffff5555ffff0000050000500033;

	lut_sub lut_1929 ({sk[420], n_n6, n_n5, x186x, x90x, x733x, x258x}, x19743x);
	defparam lut_1929.LUT_SIZE = 7;
	defparam lut_1929.mask = 128'h5555ffff5555ffff333377ff3f3f7fff;

	lut_sub lut_1934 ({sk[421], n_n6, x60x, x5260x, x79x, n_n70, x1893x}, x19747x);
	defparam lut_1934.LUT_SIZE = 7;
	defparam lut_1934.mask = 128'h5555ffff5555ffff00ff00ff7fffffff;

	lut_sub lut_1940 ({sk[422], n_n6, n_n5, n_n108, x125x, x60x, x1880x}, x19748x);
	defparam lut_1940.LUT_SIZE = 7;
	defparam lut_1940.mask = 128'h5555ffff5555ffff000077770fff7fff;

	lut_sub lut_1945 ({sk[423], n_n6, n_n5, n_n65, n_n4826, x125x, x44x}, x24172x);
	defparam lut_1945.LUT_SIZE = 7;
	defparam lut_1945.mask = 128'h5555ffff5555fffff0f0c000a0a08000;

	lut_sub lut_1950 ({sk[424], n_n6, x176x, x19743x, x19747x, x19748x, x24172x}, x513x);
	defparam lut_1950.LUT_SIZE = 7;
	defparam lut_1950.mask = 128'h5555ffff5555ffffbfffbfffbfffffff;

	lut_sub lut_1956 ({sk[425], n_n6, n_n5, n_n111, x49x, x131x, x1884x}, x19753x);
	defparam lut_1956.LUT_SIZE = 7;
	defparam lut_1956.mask = 128'h5555ffff5555ffff000055ff3f3f7fff;

	lut_sub lut_1961 ({sk[426], n_n6, n_n5, n_n32, x92x, x207x, x1876x}, x19754x);
	defparam lut_1961.LUT_SIZE = 7;
	defparam lut_1961.mask = 128'h5555ffff5555ffff00000fff77777fff;

	lut_sub lut_1966 ({sk[427], n_n6, n_n5, x55x, x56x, x1919x, x1944x}, x19755x);
	defparam lut_1966.LUT_SIZE = 7;
	defparam lut_1966.mask = 128'h5555ffff5555ffff000033ff5f5f7fff;

	lut_sub lut_1971 ({sk[428], n_n6, n_n5, n_n76, x1937x, x1945x, x1921x}, x19756x);
	defparam lut_1971.LUT_SIZE = 7;
	defparam lut_1971.mask = 128'h5555ffff5555ffff000077770fff7fff;

	lut_sub lut_1976 ({sk[429], x19753x, x19754x, x19755x, x19756x}, x551x);
	defparam lut_1976.LUT_SIZE = 5;
	defparam lut_1976.mask = 32'h0f0f7fff;

	lut_sub lut_1981 ({sk[430], i_7_, i_8_, i_6_, x915x}, n_n1);
	defparam lut_1981.LUT_SIZE = 5;
	defparam lut_1981.mask = 32'h0f0f0400;

	lut_sub lut_1983 ({sk[431], i_7_, i_8_, i_6_, x915x}, n_n2);
	defparam lut_1983.LUT_SIZE = 5;
	defparam lut_1983.mask = 32'h0f0f4000;

	lut_sub lut_1985 ({sk[432], x915x, n_n273, n_n283, x1623x, x1624x, x19776x}, x19778x);
	defparam lut_1985.LUT_SIZE = 7;
	defparam lut_1985.mask = 128'h5555ffff5555ffff5555555555775f7f;

	lut_sub lut_1989 ({sk[433], n_n2597, n_n2598, x812x, x19770x, x24157x}, x19779x);
	defparam lut_1989.LUT_SIZE = 6;
	defparam lut_1989.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_1995 ({sk[434], n_n2589, x5185x, x19791x}, x19793x);
	defparam lut_1995.LUT_SIZE = 4;
	defparam lut_1995.mask = 16'h557f;

	lut_sub lut_1999 ({sk[435], x19785x, x19787x, x19788x, x24142x}, x19794x);
	defparam lut_1999.LUT_SIZE = 5;
	defparam lut_1999.mask = 32'h0f0fbfff;

	lut_sub lut_2004 ({sk[436], n_n106, n_n2, n_n3162, x591x, x1925x, x1627x}, x19810x);
	defparam lut_2004.LUT_SIZE = 7;
	defparam lut_2004.mask = 128'h5555ffff5555ffff0fff7fff0fffffff;

	lut_sub lut_2010 ({sk[437], x19798x, x19804x, x19805x, x19796x, x19797x}, x19811x);
	defparam lut_2010.LUT_SIZE = 6;
	defparam lut_2010.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_2016 ({sk[438], i_9_, i_10_, i_11_, i_15_}, x908x);
	defparam lut_2016.LUT_SIZE = 5;
	defparam lut_2016.mask = 32'h0f0f0020;

	lut_sub lut_2018 ({sk[439], n_n281, x915x, n_n273, x908x, n_n59, x156x}, x5161x);
	defparam lut_2018.LUT_SIZE = 7;
	defparam lut_2018.mask = 128'h5555ffff5555ffff000000770000007f;

	lut_sub lut_2022 ({sk[440], i_7_, i_8_, i_6_, n_n281, x915x, x908x}, x5159x);
	defparam lut_2022.LUT_SIZE = 7;
	defparam lut_2022.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_2024 ({sk[441], i_14_, i_13_, i_12_, i_15_, n_n247, n_n242}, x1359x);
	defparam lut_2024.LUT_SIZE = 7;
	defparam lut_2024.mask = 128'h5555ffff5555ffff0700700070000000;

	lut_sub lut_2031 ({sk[442], i_9_, i_10_, n_n122}, x5144x);
	defparam lut_2031.LUT_SIZE = 4;
	defparam lut_2031.mask = 16'h5540;

	lut_sub lut_2033 ({sk[443], x913x, x266x, x294x, n_n127, n_n220, x54x}, x5139x);
	defparam lut_2033.LUT_SIZE = 7;
	defparam lut_2033.mask = 128'h5555ffff5555ffff050f0f0f070f0f0f;

	lut_sub lut_2038 ({sk[444], i_14_, i_13_, i_12_, x911x}, n_n133);
	defparam lut_2038.LUT_SIZE = 5;
	defparam lut_2038.mask = 32'h0f0f4000;

	lut_sub lut_2040 ({sk[445], i_7_, i_8_, i_6_}, n_n266);
	defparam lut_2040.LUT_SIZE = 4;
	defparam lut_2040.mask = 16'h5501;

	lut_sub lut_2042 ({sk[446], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x916x);
	defparam lut_2042.LUT_SIZE = 7;
	defparam lut_2042.mask = 128'h5555ffff5555ffff8000000000000000;

	lut_sub lut_2044 ({sk[447], i_7_, i_8_, i_6_, x916x}, n_n265);
	defparam lut_2044.LUT_SIZE = 5;
	defparam lut_2044.mask = 32'h0f0f0001;

	lut_sub lut_2046 ({sk[448], i_7_, i_8_, i_6_, x916x}, n_n268);
	defparam lut_2046.LUT_SIZE = 5;
	defparam lut_2046.mask = 32'h0f0f0010;

	lut_sub lut_2048 ({sk[449], i_14_, i_13_, i_12_, x916x, n_n271, x912x}, n_n3246);
	defparam lut_2048.LUT_SIZE = 7;
	defparam lut_2048.mask = 128'h5555ffff5555ffff0101000100000000;

	lut_sub lut_2052 ({sk[450], i_14_, i_13_, i_12_, x907x, x901x}, x101x);
	defparam lut_2052.LUT_SIZE = 6;
	defparam lut_2052.mask = 64'h3f3f3f3f00000305;

	lut_sub lut_2055 ({sk[451], i_14_, i_13_, i_12_, x901x}, n_n62);
	defparam lut_2055.LUT_SIZE = 5;
	defparam lut_2055.mask = 32'h0f0f0400;

	lut_sub lut_2057 ({sk[452], i_14_, i_13_, i_12_, x916x, n_n271, x914x}, x598x);
	defparam lut_2057.LUT_SIZE = 7;
	defparam lut_2057.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_2059 ({sk[453], i_14_, i_13_, i_12_, x903x}, x124x);
	defparam lut_2059.LUT_SIZE = 5;
	defparam lut_2059.mask = 32'h0f0f0045;

	lut_sub lut_2063 ({sk[454], n_n281, x916x, n_n271, x911x, x84x}, n_n3513);
	defparam lut_2063.LUT_SIZE = 6;
	defparam lut_2063.mask = 64'h3f3f3f3f00050007;

	lut_sub lut_2066 ({sk[455], i_14_, i_13_, i_12_, i_15_, n_n242, x19851x}, x1729x);
	defparam lut_2066.LUT_SIZE = 7;
	defparam lut_2066.mask = 128'h5555ffff5555ffff5575757577577775;

	lut_sub lut_2077 ({sk[456], i_7_, i_8_, i_6_, x916x, x212x, x277x}, x24152x);
	defparam lut_2077.LUT_SIZE = 7;
	defparam lut_2077.mask = 128'h5555ffff5555fffffffffffffffcfffa;

	lut_sub lut_2084 ({sk[457], i_14_, i_13_, i_12_, x907x}, n_n33);
	defparam lut_2084.LUT_SIZE = 5;
	defparam lut_2084.mask = 32'h0f0f0100;

	lut_sub lut_2086 ({sk[458], i_14_, i_13_, i_12_, x907x}, x78x);
	defparam lut_2086.LUT_SIZE = 5;
	defparam lut_2086.mask = 32'h0f0f1400;

	lut_sub lut_2089 ({sk[459], i_14_, i_13_, i_12_, x907x}, x268x);
	defparam lut_2089.LUT_SIZE = 5;
	defparam lut_2089.mask = 32'h0f0f1500;

	lut_sub lut_2093 ({sk[460], i_9_, i_10_, i_11_}, n_n242);
	defparam lut_2093.LUT_SIZE = 4;
	defparam lut_2093.mask = 16'h5520;

	lut_sub lut_2095 ({sk[461], i_14_, i_13_, i_12_, i_15_, x911x, n_n242}, x400x);
	defparam lut_2095.LUT_SIZE = 7;
	defparam lut_2095.mask = 128'h5555ffff5555ffff5000050000000033;

	lut_sub lut_2099 ({sk[462], i_7_, i_5_, i_6_, i_3_, i_4_, n_n165}, n_n5796);
	defparam lut_2099.LUT_SIZE = 7;
	defparam lut_2099.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_2101 ({sk[463], i_7_, i_8_, i_6_, x909x, x72x, n_n206}, n_n4809);
	defparam lut_2101.LUT_SIZE = 7;
	defparam lut_2101.mask = 128'h5555ffff5555ffff0000000005000300;

	lut_sub lut_2104 ({sk[464], i_14_, i_13_, i_12_, x906x}, x153x);
	defparam lut_2104.LUT_SIZE = 5;
	defparam lut_2104.mask = 32'h0f0f1500;

	lut_sub lut_2108 ({sk[465], i_14_, i_13_, i_12_, i_15_, x914x, n_n137}, x189x);
	defparam lut_2108.LUT_SIZE = 7;
	defparam lut_2108.mask = 128'h5555ffff5555ffff5050505073505073;

	lut_sub lut_2112 ({sk[466], i_7_, i_8_, i_6_, x909x, x99x, x1907x}, n_n4770);
	defparam lut_2112.LUT_SIZE = 7;
	defparam lut_2112.mask = 128'h5555ffff5555ffff0000000007000000;

	lut_sub lut_2115 ({sk[467], n_n6, x153x, x189x, n_n4770, n_n4773, n_n4772}, x19872x);
	defparam lut_2115.LUT_SIZE = 7;
	defparam lut_2115.mask = 128'h5555ffff5555ffff7f7f7f7f7fffffff;

	lut_sub lut_2121 ({sk[468], i_14_, i_13_, i_12_, x900x, x906x}, x1895x);
	defparam lut_2121.LUT_SIZE = 6;
	defparam lut_2121.mask = 64'h3f3f3f3f33035055;

	lut_sub lut_2128 ({sk[469], n_n6, n_n5, x904x, n_n225, x219x, x77x}, x616x);
	defparam lut_2128.LUT_SIZE = 7;
	defparam lut_2128.mask = 128'h5555ffff5555ffff0000555f3333777f;

	lut_sub lut_2132 ({sk[470], x909x, n_n261, x99x, x632x, x1911x}, n_n4774);
	defparam lut_2132.LUT_SIZE = 6;
	defparam lut_2132.mask = 64'h3f3f3f3f3333337f;

	lut_sub lut_2136 ({sk[471], n_n6, n_n111, x131x, x5376x, x19862x, x1859x}, x19865x);
	defparam lut_2136.LUT_SIZE = 7;
	defparam lut_2136.mask = 128'h5555ffff5555ffff3f3f3f3f7fffffff;

	lut_sub lut_2142 ({sk[472], n_n6, n_n5, n_n32, x1894x, x205x, x1876x}, x19866x);
	defparam lut_2142.LUT_SIZE = 7;
	defparam lut_2142.mask = 128'h5555ffff5555ffff00003fff55557fff;

	lut_sub lut_2147 ({sk[473], n_n6, x1895x, x616x, n_n4774, x19865x, x19866x}, x19873x);
	defparam lut_2147.LUT_SIZE = 7;
	defparam lut_2147.mask = 128'h5555ffff5555ffff7fff7fff7fffffff;

	lut_sub lut_2153 ({sk[474], x541x, n_n5, n_n4815, x522x, x265x, x137x}, x24140x);
	defparam lut_2153.LUT_SIZE = 7;
	defparam lut_2153.mask = 128'h5555ffff5555fffff000800000000000;

	lut_sub lut_2156 ({sk[475], n_n6, n_n5, x146x, x498x, n_n59, x132x}, x24174x);
	defparam lut_2156.LUT_SIZE = 7;
	defparam lut_2156.mask = 128'h5555ffff5555fffff0f0a000c0c08000;

	lut_sub lut_2161 ({sk[476], n_n110, n_n5, x125x, x90x, x5259x, x155x}, x19882x);
	defparam lut_2161.LUT_SIZE = 7;
	defparam lut_2161.mask = 128'h5555ffff5555ffff33337fff3333ffff;

	lut_sub lut_2167 ({sk[477], n_n110, n_n6, n_n5, x90x, x1893x, x1922x}, x19883x);
	defparam lut_2167.LUT_SIZE = 7;
	defparam lut_2167.mask = 128'h5555ffff5555ffff00553f7f0055ffff;

	lut_sub lut_2172 ({sk[478], x909x, n_n65, n_n261, n_n263, n_n11, x44x}, x19876x);
	defparam lut_2172.LUT_SIZE = 7;
	defparam lut_2172.mask = 128'h5555ffff5555ffff0000000005770f7f;

	lut_sub lut_2177 ({sk[479], n_n12, x909x, n_n261, n_n263, x265x, x70x}, x19877x);
	defparam lut_2177.LUT_SIZE = 7;
	defparam lut_2177.mask = 128'h5555ffff5555ffff00000537000005ff;

	lut_sub lut_2181 ({sk[480], n_n5, x186x, n_n4826, n_n4823, x258x, x293x}, x24139x);
	defparam lut_2181.LUT_SIZE = 7;
	defparam lut_2181.mask = 128'h5555ffff5555fffff000f00080000000;

	lut_sub lut_2184 ({sk[481], n_n6, x82x, x111x, x79x, n_n70, x5386x}, x19896x);
	defparam lut_2184.LUT_SIZE = 7;
	defparam lut_2184.mask = 128'h5555ffff5555ffff555555557fffffff;

	lut_sub lut_2190 ({sk[482], n_n6, n_n5, n_n108, x125x, x60x, x1075x}, x19897x);
	defparam lut_2190.LUT_SIZE = 7;
	defparam lut_2190.mask = 128'h5555ffff5555ffff000077770fff7fff;

	lut_sub lut_2195 ({sk[483], n_n6, n_n5, n_n111, x49x, x207x, x1945x}, x19900x);
	defparam lut_2195.LUT_SIZE = 7;
	defparam lut_2195.mask = 128'h5555ffff5555ffff000055ff3f3f7fff;

	lut_sub lut_2200 ({sk[484], n_n6, n_n5, x136x, x55x, x1937x, x1944x}, x19901x);
	defparam lut_2200.LUT_SIZE = 7;
	defparam lut_2200.mask = 128'h5555ffff5555ffff00000fff77777fff;

	lut_sub lut_2205 ({sk[485], n_n6, n_n5, n_n4846, x92x, x56x, x1919x}, x19904x);
	defparam lut_2205.LUT_SIZE = 7;
	defparam lut_2205.mask = 128'h5555ffff5555ffff00ff5fff33ff7fff;

	lut_sub lut_2210 ({sk[486], n_n6, n_n5, n_n76, x1920x, x147x, x1921x}, x19905x);
	defparam lut_2210.LUT_SIZE = 7;
	defparam lut_2210.mask = 128'h5555ffff5555ffff000055553fff7fff;

	lut_sub lut_2215 ({sk[487], i_7_, i_8_, i_6_, x909x}, n_n57);
	defparam lut_2215.LUT_SIZE = 5;
	defparam lut_2215.mask = 32'h0f0f0001;

	lut_sub lut_2217 ({sk[488], i_7_, i_8_, i_6_, x909x, n_n228, x912x}, x5022x);
	defparam lut_2217.LUT_SIZE = 7;
	defparam lut_2217.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_2219 ({sk[489], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x113x);
	defparam lut_2219.LUT_SIZE = 7;
	defparam lut_2219.mask = 128'h5555ffff5555ffff4000100000000000;

	lut_sub lut_2222 ({sk[490], n_n106, n_n266, n_n271, x101x, x909x, x293x}, x884x);
	defparam lut_2222.LUT_SIZE = 7;
	defparam lut_2222.mask = 128'h5555ffff5555ffff0011031300330333;

	lut_sub lut_2226 ({sk[491], n_n266, n_n271, x146x, x909x, x265x, x393x}, x19918x);
	defparam lut_2226.LUT_SIZE = 7;
	defparam lut_2226.mask = 128'h5555ffff5555ffff55555757555f575f;

	lut_sub lut_2230 ({sk[492], n_n266, x909x, x265x, x5019x, n_n11, n_n60}, x24181x);
	defparam lut_2230.LUT_SIZE = 7;
	defparam lut_2230.mask = 128'h5555ffff5555fffff0f0f0f0f0f08000;

	lut_sub lut_2234 ({sk[493], n_n57, x5022x, x113x, x884x, x19918x, x24181x}, x19921x);
	defparam lut_2234.LUT_SIZE = 7;
	defparam lut_2234.mask = 128'h5555ffff5555ffffbfbfffffbfffffff;

	lut_sub lut_2240 ({sk[494], n_n151, x183x, n_n266, n_n271, x909x, x118x}, x709x);
	defparam lut_2240.LUT_SIZE = 7;
	defparam lut_2240.mask = 128'h5555ffff5555ffff0101013301330133;

	lut_sub lut_2244 ({sk[495], n_n57, n_n56, x878x, n_n59, x156x, x132x}, x19910x);
	defparam lut_2244.LUT_SIZE = 7;
	defparam lut_2244.mask = 128'h5555ffff5555ffff00ff55ff3fff7fff;

	lut_sub lut_2249 ({sk[496], n_n155, x924x, x218x, x146x, n_n56, x72x}, x19909x);
	defparam lut_2249.LUT_SIZE = 7;
	defparam lut_2249.mask = 128'h5555ffff5555ffff133313331333ffff;

	lut_sub lut_2254 ({sk[497], n_n110, n_n266, n_n271, x909x, x90x, x82x}, x19913x);
	defparam lut_2254.LUT_SIZE = 7;
	defparam lut_2254.mask = 128'h5555ffff5555ffff0005030700050f0f;

	lut_sub lut_2258 ({sk[498], n_n108, n_n57, n_n56, x111x, x1898x, x70x}, x19914x);
	defparam lut_2258.LUT_SIZE = 7;
	defparam lut_2258.mask = 128'h5555ffff5555ffff003f557f00ff55ff;

	lut_sub lut_2263 ({sk[499], x709x, x19910x, n_n4781, x19909x, x19913x, x19914x}, x19922x);
	defparam lut_2263.LUT_SIZE = 7;
	defparam lut_2263.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_2270 ({sk[500], n_n57, n_n56, x219x, x189x, x277x, x112x}, x19926x);
	defparam lut_2270.LUT_SIZE = 7;
	defparam lut_2270.mask = 128'h5555ffff5555ffff00000fff77777fff;

	lut_sub lut_2275 ({sk[501], x268x, n_n57, n_n56, x200x, x157x, n_n4940}, x19927x);
	defparam lut_2275.LUT_SIZE = 7;
	defparam lut_2275.mask = 128'h5555ffff5555ffff55775f7f55ffffff;

	lut_sub lut_2281 ({sk[502], n_n266, n_n271, x909x, n_n4959, x166x, x180x}, x19973x);
	defparam lut_2281.LUT_SIZE = 7;
	defparam lut_2281.mask = 128'h5555ffff5555ffff0f0f0f7f0f3f0f7f;

	lut_sub lut_2286 ({sk[503], n_n57, n_n56, x180x, x224x, x254x, x1683x}, x19974x);
	defparam lut_2286.LUT_SIZE = 7;
	defparam lut_2286.mask = 128'h5555ffff5555ffff000077770fff7fff;

	lut_sub lut_2291 ({sk[504], n_n266, x909x, n_n4952, x219x, x189x, x157x}, x19978x);
	defparam lut_2291.LUT_SIZE = 7;
	defparam lut_2291.mask = 128'h5555ffff5555ffff00ff00ff00ff7fff;

	lut_sub lut_2296 ({sk[505], n_n56, n_n4948, x99x, n_n4955, n_n4950, x112x}, x19979x);
	defparam lut_2296.LUT_SIZE = 7;
	defparam lut_2296.mask = 128'h5555ffff5555ffff3f3fffff7fffffff;

	lut_sub lut_2302 ({sk[506], x19926x, x19927x, x19973x, x19974x, x19978x, x19979x}, x19982x);
	defparam lut_2302.LUT_SIZE = 7;
	defparam lut_2302.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_2309 ({sk[507], n_n271, x909x, x163x, x763x, x19943x, x19944x}, x19946x);
	defparam lut_2309.LUT_SIZE = 7;
	defparam lut_2309.mask = 128'h5555ffff5555ffff7f7f7f7f7f7f7fff;

	lut_sub lut_2314 ({sk[508], x19930x, x19931x, x19937x, x19932x, x19933x}, x19947x);
	defparam lut_2314.LUT_SIZE = 6;
	defparam lut_2314.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_2320 ({sk[509], i_7_, i_6_, x917x, x4962x, x4958x, x24180x}, n_n4744);
	defparam lut_2320.LUT_SIZE = 7;
	defparam lut_2320.mask = 128'h5555ffff5555ffffbfbfbfbfbfbfbfff;

	lut_sub lut_2325 ({sk[510], x19953x, x19954x, x19965x, x19966x}, x19968x);
	defparam lut_2325.LUT_SIZE = 5;
	defparam lut_2325.mask = 32'h0f0f7fff;

	lut_sub lut_2330 ({sk[511], i_7_, i_5_, i_6_, i_3_, i_4_, n_n118}, n_n5668);
	defparam lut_2330.LUT_SIZE = 7;
	defparam lut_2330.mask = 128'h5555ffff5555ffff1000000000000000;

	lut_sub lut_2332 ({sk[512], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, x879x);
	defparam lut_2332.LUT_SIZE = 7;
	defparam lut_2332.mask = 128'h5555ffff5555ffff4040001040001010;

	lut_sub lut_2339 ({sk[513], i_7_, i_5_, i_6_, i_3_, i_4_, n_n118}, x859x);
	defparam lut_2339.LUT_SIZE = 7;
	defparam lut_2339.mask = 128'h5555ffff5555ffff0010101010101000;

	lut_sub lut_2346 ({sk[514], x921x, n_n283, n_n220, n_n122, x914x, x905x}, x20007x);
	defparam lut_2346.LUT_SIZE = 7;
	defparam lut_2346.mask = 128'h5555ffff5555ffff0005000500050077;

	lut_sub lut_2350 ({sk[515], i_14_, i_13_, i_12_, x905x}, n_n108);
	defparam lut_2350.LUT_SIZE = 5;
	defparam lut_2350.mask = 32'h0f0f0400;

	lut_sub lut_2352 ({sk[516], i_14_, i_13_, i_12_, n_n121, x914x}, x759x);
	defparam lut_2352.LUT_SIZE = 6;
	defparam lut_2352.mask = 64'h3f3f3f3f00100000;

	lut_sub lut_2354 ({sk[517], i_7_, i_8_, i_6_, x896x}, n_n128);
	defparam lut_2354.LUT_SIZE = 5;
	defparam lut_2354.mask = 32'h0f0f0010;

	lut_sub lut_2356 ({sk[518], n_n281, x913x, n_n56, n_n258, x709x, n_n150}, n_n4251);
	defparam lut_2356.LUT_SIZE = 7;
	defparam lut_2356.mask = 128'h5555ffff5555ffff3377337f337733ff;

	lut_sub lut_2361 ({sk[519], i_7_, i_8_, i_6_, x146x, x909x}, n_n4892);
	defparam lut_2361.LUT_SIZE = 6;
	defparam lut_2361.mask = 64'h3f3f3f3f00000100;

	lut_sub lut_2363 ({sk[520], n_n271, x909x, n_n258, n_n228, x903x, x897x}, x5019x);
	defparam lut_2363.LUT_SIZE = 7;
	defparam lut_2363.mask = 128'h5555ffff5555ffff0000000000000537;

	lut_sub lut_2366 ({sk[521], i_7_, i_8_, i_6_, n_n281, x909x, x908x}, x5020x);
	defparam lut_2366.LUT_SIZE = 7;
	defparam lut_2366.mask = 128'h5555ffff5555ffff0000000000000001;

	lut_sub lut_2368 ({sk[522], n_n266, n_n271, x909x, n_n59, x156x, x132x}, x488x);
	defparam lut_2368.LUT_SIZE = 7;
	defparam lut_2368.mask = 128'h5555ffff5555ffff00000055003f007f;

	lut_sub lut_2372 ({sk[523], n_n266, n_n271, x909x, n_n60, n_n206, x1870x}, x878x);
	defparam lut_2372.LUT_SIZE = 7;
	defparam lut_2372.mask = 128'h5555ffff5555ffff0000003f0055007f;

	lut_sub lut_2376 ({sk[524], n_n4251, n_n4892, x5019x, x5020x, x488x, x878x}, n_n4548);
	defparam lut_2376.LUT_SIZE = 7;
	defparam lut_2376.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_2383 ({sk[525], n_n266, x909x, x176x, n_n228, x912x, x393x}, n_n4256);
	defparam lut_2383.LUT_SIZE = 7;
	defparam lut_2383.mask = 128'h5555ffff5555ffff55555555555557ff;

	lut_sub lut_2387 ({sk[526], x909x, n_n258, n_n261, x389x, x900x, x174x}, x20127x);
	defparam lut_2387.LUT_SIZE = 7;
	defparam lut_2387.mask = 128'h5555ffff5555ffff0f0f0f0f0f5f0f7f;

	lut_sub lut_2391 ({sk[527], n_n6, n_n5, n_n6524, x1905x, x1613x, x4763x}, x20128x);
	defparam lut_2391.LUT_SIZE = 7;
	defparam lut_2391.mask = 128'h5555ffff5555ffff55ff77ff5fff7fff;

	lut_sub lut_2396 ({sk[528], n_n57, x265x, x5022x, x734x, x113x, x884x}, x24188x);
	defparam lut_2396.LUT_SIZE = 7;
	defparam lut_2396.mask = 128'h5555ffff5555ffffa000a00080000000;

	lut_sub lut_2399 ({sk[529], n_n4256, x20127x, x20128x, x24188x}, x20130x);
	defparam lut_2399.LUT_SIZE = 5;
	defparam lut_2399.mask = 32'h0f0fbfff;

	lut_sub lut_2404 ({sk[530], n_n6, n_n5, n_n41, x115x, x77x, x174x}, n_n3180);
	defparam lut_2404.LUT_SIZE = 7;
	defparam lut_2404.mask = 128'h5555ffff5555ffff000077770fff7fff;

	lut_sub lut_2409 ({sk[531], i_14_, i_13_, i_12_, i_15_, n_n267}, x1760x);
	defparam lut_2409.LUT_SIZE = 6;
	defparam lut_2409.mask = 64'h3f3f3f3f11055054;

	lut_sub lut_2419 ({sk[532], x909x, n_n54, x51x, n_n261, n_n263, x1928x}, x20145x);
	defparam lut_2419.LUT_SIZE = 7;
	defparam lut_2419.mask = 128'h5555ffff5555ffff00000000111f333f;

	lut_sub lut_2423 ({sk[533], x909x, n_n261, n_n3180, x1760x, x20145x}, x20147x);
	defparam lut_2423.LUT_SIZE = 6;
	defparam lut_2423.mask = 64'h3f3f3f3f5f5f5f7f;

	lut_sub lut_2427 ({sk[534], n_n111, x909x, n_n261, x213x, n_n6582, x222x}, x317x);
	defparam lut_2427.LUT_SIZE = 7;
	defparam lut_2427.mask = 128'h5555ffff5555ffff3333337f333333ff;

	lut_sub lut_2432 ({sk[535], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x1611x);
	defparam lut_2432.LUT_SIZE = 7;
	defparam lut_2432.mask = 128'h5555ffff5555ffff3305005555055550;

	lut_sub lut_2443 ({sk[536], n_n6, n_n5, x115x, x141x, x181x, x222x}, x20142x);
	defparam lut_2443.LUT_SIZE = 7;
	defparam lut_2443.mask = 128'h5555ffff5555ffff000055ff3f3f7fff;

	lut_sub lut_2448 ({sk[537], n_n6, x78x, n_n5, n_n41, x67x, x213x}, x20141x);
	defparam lut_2448.LUT_SIZE = 7;
	defparam lut_2448.mask = 128'h5555ffff5555ffff007f007f007fffff;

	lut_sub lut_2453 ({sk[538], n_n6, n_n104, x4743x, x1927x, x221x, x20136x}, x24137x);
	defparam lut_2453.LUT_SIZE = 7;
	defparam lut_2453.mask = 128'h5555ffff5555ffffff00ff0080000000;

	lut_sub lut_2456 ({sk[539], n_n5, x317x, x1611x, x20142x, x20141x, x24137x}, x20148x);
	defparam lut_2456.LUT_SIZE = 7;
	defparam lut_2456.mask = 128'h5555ffff5555ffffbfbfffffbfffffff;

	lut_sub lut_2462 ({sk[540], n_n197, x909x, n_n261, x4716x, x411x, x1946x}, x20153x);
	defparam lut_2462.LUT_SIZE = 7;
	defparam lut_2462.mask = 128'h5555ffff5555ffff3f3f3f7f3f3f3fff;

	lut_sub lut_2467 ({sk[541], n_n6, n_n5, x188x, x141x, x181x, x1778x}, x20154x);
	defparam lut_2467.LUT_SIZE = 7;
	defparam lut_2467.mask = 128'h5555ffff5555ffff00007f7f00ff7fff;

	lut_sub lut_2472 ({sk[542], n_n197, x909x, n_n261, n_n263, x62x, x1926x}, x20157x);
	defparam lut_2472.LUT_SIZE = 7;
	defparam lut_2472.mask = 128'h5555ffff5555ffff0000053700000f3f;

	lut_sub lut_2476 ({sk[543], x909x, n_n261, n_n263, x62x, x1781x, x1780x}, x20158x);
	defparam lut_2476.LUT_SIZE = 7;
	defparam lut_2476.mask = 128'h5555ffff5555ffff00000000003f557f;

	lut_sub lut_2480 ({sk[544], x909x, n_n258, n_n261, x40x, x897x, x1904x}, x20164x);
	defparam lut_2480.LUT_SIZE = 7;
	defparam lut_2480.mask = 128'h5555ffff5555ffff00000000005f007f;

	lut_sub lut_2484 ({sk[545], n_n6, n_n5, n_n103, x593x, x91x, x1782x}, x20165x);
	defparam lut_2484.LUT_SIZE = 7;
	defparam lut_2484.mask = 128'h5555ffff5555ffff0f0f5fff3f3f7fff;

	lut_sub lut_2489 ({sk[546], x20153x, x20154x, x20157x, x20158x, x20164x, x20165x}, n_n4532);
	defparam lut_2489.LUT_SIZE = 7;
	defparam lut_2489.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_2496 ({sk[547], n_n220, x911x, x909x, x159x, n_n261, x225x}, x20168x);
	defparam lut_2496.LUT_SIZE = 7;
	defparam lut_2496.mask = 128'h5555ffff5555ffff0013001300130033;

	lut_sub lut_2500 ({sk[548], n_n281, x913x, x183x, x390x, x909x, n_n263}, x20169x);
	defparam lut_2500.LUT_SIZE = 7;
	defparam lut_2500.mask = 128'h5555ffff5555ffff0f1f0f1f0f1f1f1f;

	lut_sub lut_2504 ({sk[549], n_n6, n_n5, x523x, x208x, n_n59, n_n3803}, x20176x);
	defparam lut_2504.LUT_SIZE = 7;
	defparam lut_2504.mask = 128'h5555ffff5555ffff55ff7fff5fff7fff;

	lut_sub lut_2510 ({sk[550], n_n6, n_n5, x199x, n_n63, x20173x, x24136x}, x20177x);
	defparam lut_2510.LUT_SIZE = 7;
	defparam lut_2510.mask = 128'h5555ffff5555ffff0000aaaa3fffbfff;

	lut_sub lut_2515 ({sk[551], n_n5, x101x, n_n12, x176x, x121x, n_n15}, x4680x);
	defparam lut_2515.LUT_SIZE = 7;
	defparam lut_2515.mask = 128'h5555ffff5555ffff000000007fffffff;

	lut_sub lut_2521 ({sk[552], x909x, n_n261, n_n263, x1325x, x1324x, x1827x}, x20183x);
	defparam lut_2521.LUT_SIZE = 7;
	defparam lut_2521.mask = 128'h5555ffff5555ffff0000000000335f7f;

	lut_sub lut_2525 ({sk[553], x20168x, x20169x, x20176x, x20177x, x4680x, x20183x}, n_n4531);
	defparam lut_2525.LUT_SIZE = 7;
	defparam lut_2525.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_2532 ({sk[554], n_n271, x909x, n_n3204, x1885x, x1761x, x20204x}, x20209x);
	defparam lut_2532.LUT_SIZE = 7;
	defparam lut_2532.mask = 128'h5555ffff5555ffff55ff55ff55ff7fff;

	lut_sub lut_2537 ({sk[555], x20200x, x20201x, n_n3711, x20205x}, x20210x);
	defparam lut_2537.LUT_SIZE = 5;
	defparam lut_2537.mask = 32'h0f0f7fff;

	lut_sub lut_2542 ({sk[556], n_n266, x909x, x179x, n_n4677, x20220x, x20219x}, n_n4556);
	defparam lut_2542.LUT_SIZE = 7;
	defparam lut_2542.mask = 128'h5555ffff5555ffff7f7f7f7f7f7f7fff;

	lut_sub lut_2547 ({sk[557], n_n4259, x465x, n_n3708, x20227x}, x20232x);
	defparam lut_2547.LUT_SIZE = 5;
	defparam lut_2547.mask = 32'h0f0f7fff;

	lut_sub lut_2552 ({sk[558], x682x, n_n4261, x721x, n_n3709, x24178x}, x20233x);
	defparam lut_2552.LUT_SIZE = 6;
	defparam lut_2552.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_2558 ({sk[559], n_n4598, n_n4596, x20215x, x20214x, x20238x}, x20240x);
	defparam lut_2558.LUT_SIZE = 6;
	defparam lut_2558.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_2564 ({sk[560], n_n48, n_n105, x94x, x108x, n_n4183, x571x}, x20304x);
	defparam lut_2564.LUT_SIZE = 7;
	defparam lut_2564.mask = 128'h5555ffff5555ffff777777777fffffff;

	lut_sub lut_2570 ({sk[561], n_n53, x407x, x457x, x77x, x1233x, x20300x}, x20305x);
	defparam lut_2570.LUT_SIZE = 7;
	defparam lut_2570.mask = 128'h5555ffff5555ffff55ffffff7fffffff;

	lut_sub lut_2576 ({sk[562], n_n104, n_n41, n_n48, n_n53, x67x, x1433x}, x20312x);
	defparam lut_2576.LUT_SIZE = 7;
	defparam lut_2576.mask = 128'h5555ffff5555ffff07070f0f0fff0fff;

	lut_sub lut_2582 ({sk[563], n_n258, x898x, x51x, n_n48, x619x, x1366x}, x20318x);
	defparam lut_2582.LUT_SIZE = 7;
	defparam lut_2582.mask = 128'h5555ffff5555ffff373f373f373f3f3f;

	lut_sub lut_2587 ({sk[564], i_7_, i_8_, i_6_, x922x, x1367x, x1434x}, x24135x);
	defparam lut_2587.LUT_SIZE = 7;
	defparam lut_2587.mask = 128'h5555ffff5555fffffafffcffffffffff;

	lut_sub lut_2594 ({sk[565], x20304x, x20305x, x20312x, x20318x, x24135x}, n_n3901);
	defparam lut_2594.LUT_SIZE = 6;
	defparam lut_2594.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_2600 ({sk[566], n_n48, x368x, n_n6505, x483x, x20253x, x24189x}, n_n3925);
	defparam lut_2600.LUT_SIZE = 7;
	defparam lut_2600.mask = 128'h5555ffff5555ffffbfffbfffbfffffff;

	lut_sub lut_2606 ({sk[567], n_n31, n_n48, x4600x, x864x, n_n4073, x20263x}, n_n3923);
	defparam lut_2606.LUT_SIZE = 7;
	defparam lut_2606.mask = 128'h5555ffff5555ffff7fff7fff7fffffff;

	lut_sub lut_2612 ({sk[568], n_n3978, x20282x, x4557x, x20288x, n_n3980}, x20295x);
	defparam lut_2612.LUT_SIZE = 6;
	defparam lut_2612.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_2618 ({sk[569], n_n48, x20290x, x20291x, x20269x, x20270x, x20293x}, x24134x);
	defparam lut_2618.LUT_SIZE = 7;
	defparam lut_2618.mask = 128'h5555ffff5555ffff8080808080000000;

	lut_sub lut_2621 ({sk[570], i_7_, i_8_, i_6_, x922x}, n_n53);
	defparam lut_2621.LUT_SIZE = 5;
	defparam lut_2621.mask = 32'h0f0f0400;

	lut_sub lut_2623 ({sk[571], n_n273, x905x, n_n258, x922x, x899x, n_n228}, x676x);
	defparam lut_2623.LUT_SIZE = 7;
	defparam lut_2623.mask = 128'h5555ffff5555ffff000000000101010f;

	lut_sub lut_2626 ({sk[572], i_7_, i_8_, i_6_, x922x, x869x, x1852x}, x298x);
	defparam lut_2626.LUT_SIZE = 7;
	defparam lut_2626.mask = 128'h5555ffff5555ffff3333373333333333;

	lut_sub lut_2629 ({sk[573], n_n273, x922x, n_n60, x373x, x626x, x865x}, x20350x);
	defparam lut_2629.LUT_SIZE = 7;
	defparam lut_2629.mask = 128'h5555ffff5555ffff7f7f7f7f7f7f7fff;

	lut_sub lut_2634 ({sk[574], n_n53, x111x, n_n6878, x475x, x406x, x695x}, x24196x);
	defparam lut_2634.LUT_SIZE = 7;
	defparam lut_2634.mask = 128'h5555ffff5555ffff8000800080000000;

	lut_sub lut_2637 ({sk[575], i_7_, i_8_, i_6_, x916x}, n_n4);
	defparam lut_2637.LUT_SIZE = 5;
	defparam lut_2637.mask = 32'h0f0f0100;

	lut_sub lut_2639 ({sk[576], i_14_, i_13_, i_12_, x914x, x912x}, x95x);
	defparam lut_2639.LUT_SIZE = 6;
	defparam lut_2639.mask = 64'h3f3f3f3f00500300;

	lut_sub lut_2642 ({sk[577], i_14_, i_13_, i_12_}, n_n228);
	defparam lut_2642.LUT_SIZE = 4;
	defparam lut_2642.mask = 16'h5501;

	lut_sub lut_2644 ({sk[578], i_9_, i_10_, i_11_, i_15_, x95x, n_n228}, x206x);
	defparam lut_2644.LUT_SIZE = 7;
	defparam lut_2644.mask = 128'h5555ffff5555ffff3333333337333333;

	lut_sub lut_2647 ({sk[579], i_9_, i_10_, i_11_, i_15_}, x900x);
	defparam lut_2647.LUT_SIZE = 5;
	defparam lut_2647.mask = 32'h0f0f0100;

	lut_sub lut_2649 ({sk[580], i_14_, i_13_, i_12_, x900x}, n_n64);
	defparam lut_2649.LUT_SIZE = 5;
	defparam lut_2649.mask = 32'h0f0f0400;

	lut_sub lut_2651 ({sk[581], i_14_, i_13_, i_12_, n_n208, x916x, x900x}, n_n7402);
	defparam lut_2651.LUT_SIZE = 7;
	defparam lut_2651.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_2653 ({sk[582], i_9_, i_10_, i_11_, i_15_}, x906x);
	defparam lut_2653.LUT_SIZE = 5;
	defparam lut_2653.mask = 32'h0f0f0200;

	lut_sub lut_2655 ({sk[583], i_14_, i_13_, i_12_, x906x}, n_n13);
	defparam lut_2655.LUT_SIZE = 5;
	defparam lut_2655.mask = 32'h0f0f0010;

	lut_sub lut_2657 ({sk[584], n_n2876, n_n2875, n_n2820, x20374x, x20381x, x20382x}, n_n2798);
	defparam lut_2657.LUT_SIZE = 7;
	defparam lut_2657.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_2664 ({sk[585], n_n4, x20399x, n_n876, x20403x, x117x, x20398x}, n_n2817);
	defparam lut_2664.LUT_SIZE = 7;
	defparam lut_2664.mask = 128'h5555ffff5555ffff5fffffff7fffffff;

	lut_sub lut_2670 ({sk[586], x4319x, x20562x, x24130x, x24131x}, n_n2796);
	defparam lut_2670.LUT_SIZE = 5;
	defparam lut_2670.mask = 32'h0f0fefff;

	lut_sub lut_2675 ({sk[587], n_n3964, x736x, x20392x, x876x, x533x, x20410x}, x24199x);
	defparam lut_2675.LUT_SIZE = 7;
	defparam lut_2675.mask = 128'h5555ffff5555ffff8000000000000000;

	lut_sub lut_2677 ({sk[588], i_14_, i_13_, i_12_, n_n208, x916x, x899x}, x485x);
	defparam lut_2677.LUT_SIZE = 7;
	defparam lut_2677.mask = 128'h5555ffff5555ffff0000000000010100;

	lut_sub lut_2680 ({sk[589], i_7_, i_8_, i_6_, x916x, x374x, x1959x}, x867x);
	defparam lut_2680.LUT_SIZE = 7;
	defparam lut_2680.mask = 128'h5555ffff5555ffff3333333733333333;

	lut_sub lut_2683 ({sk[590], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1466x);
	defparam lut_2683.LUT_SIZE = 7;
	defparam lut_2683.mask = 128'h5555ffff5555ffff0104440400000000;

	lut_sub lut_2689 ({sk[591], n_n4, n_n76, x92x, x80x, n_n7306, x1941x}, x24154x);
	defparam lut_2689.LUT_SIZE = 7;
	defparam lut_2689.mask = 128'h5555ffff5555ffffcccccccc80000000;

	lut_sub lut_2692 ({sk[592], n_n208, x916x, x485x, x867x, x1466x, x24154x}, x20590x);
	defparam lut_2692.LUT_SIZE = 7;
	defparam lut_2692.mask = 128'h5555ffff5555ffffafffafffafffbfff;

	lut_sub lut_2697 ({sk[593], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x93x);
	defparam lut_2697.LUT_SIZE = 7;
	defparam lut_2697.mask = 128'h5555ffff5555ffff0010001040000000;

	lut_sub lut_2701 ({sk[594], n_n208, x916x, x905x, n_n256, x1854x}, x378x);
	defparam lut_2701.LUT_SIZE = 6;
	defparam lut_2701.mask = 64'h3f3f3f3f00000057;

	lut_sub lut_2704 ({sk[595], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1883x);
	defparam lut_2704.LUT_SIZE = 7;
	defparam lut_2704.mask = 128'h5555ffff5555ffff0010001050105040;

	lut_sub lut_2713 ({sk[596], n_n111, n_n4, x136x, x85x, x98x, x24204x}, x4304x);
	defparam lut_2713.LUT_SIZE = 7;
	defparam lut_2713.mask = 128'h5555ffff5555ffff00007fff0000ffff;

	lut_sub lut_2719 ({sk[597], n_n4, n_n65, n_n7355, x44x, x111x, x1693x}, x20583x);
	defparam lut_2719.LUT_SIZE = 7;
	defparam lut_2719.mask = 128'h5555ffff5555ffff00ff00ff7fffffff;

	lut_sub lut_2725 ({sk[598], n_n4, x93x, x378x, x1883x, x4304x, x20583x}, x20591x);
	defparam lut_2725.LUT_SIZE = 7;
	defparam lut_2725.mask = 128'h5555ffff5555ffff77ff77ff7fffffff;

	lut_sub lut_2731 ({sk[599], n_n1, x218x, x72x, x133x, x113x, x24124x}, x4281x);
	defparam lut_2731.LUT_SIZE = 7;
	defparam lut_2731.mask = 128'h5555ffff5555ffff00000000bfffffff;

	lut_sub lut_2737 ({sk[600], n_n1, n_n265, x200x, x209x, x277x, x112x}, x20600x);
	defparam lut_2737.LUT_SIZE = 7;
	defparam lut_2737.mask = 128'h5555ffff5555ffff000077ff0f0f7fff;

	lut_sub lut_2742 ({sk[601], n_n1, x206x, x410x, x186x, x354x, x440x}, x4276x);
	defparam lut_2742.LUT_SIZE = 7;
	defparam lut_2742.mask = 128'h5555ffff5555ffff000000007fffffff;

	lut_sub lut_2748 ({sk[602], x915x, n_n273, n_n108, x90x, x155x, x1864x}, x20606x);
	defparam lut_2748.LUT_SIZE = 7;
	defparam lut_2748.mask = 128'h5555ffff5555ffff0000000000007fff;

	lut_sub lut_2753 ({sk[603], n_n106, n_n265, x268x, n_n4, x101x, x1924x}, x20611x);
	defparam lut_2753.LUT_SIZE = 7;
	defparam lut_2753.mask = 128'h5555ffff5555ffff050537ff0505ffff;

	lut_sub lut_2758 ({sk[604], n_n4, n_n95, x68x, x1283x, x455x, x605x}, x20612x);
	defparam lut_2758.LUT_SIZE = 7;
	defparam lut_2758.mask = 128'h5555ffff5555ffff777777777fffffff;

	lut_sub lut_2764 ({sk[605], x4281x, x20600x, x4276x, x20606x, x20611x, x20612x}, n_n2795);
	defparam lut_2764.LUT_SIZE = 7;
	defparam lut_2764.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_2771 ({sk[606], i_14_, i_13_, i_12_, x902x}, n_n9);
	defparam lut_2771.LUT_SIZE = 5;
	defparam lut_2771.mask = 32'h0f0f0001;

	lut_sub lut_2773 ({sk[607], i_15_, n_n208, x916x, n_n220, n_n61, n_n270}, x648x);
	defparam lut_2773.LUT_SIZE = 7;
	defparam lut_2773.mask = 128'h5555ffff5555ffff0000003300000037;

	lut_sub lut_2776 ({sk[608], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1525x);
	defparam lut_2776.LUT_SIZE = 7;
	defparam lut_2776.mask = 128'h5555ffff5555ffff4000110000040001;

	lut_sub lut_2782 ({sk[609], n_n208, x916x, n_n9, x648x, n_n60, x1525x}, n_n2840);
	defparam lut_2782.LUT_SIZE = 7;
	defparam lut_2782.mask = 128'h5555ffff5555ffff0f0f0f0f0f0f7fff;

	lut_sub lut_2787 ({sk[610], i_14_, i_13_, i_12_, x903x}, n_n7);
	defparam lut_2787.LUT_SIZE = 5;
	defparam lut_2787.mask = 32'h0f0f4000;

	lut_sub lut_2789 ({sk[611], i_7_, i_8_, i_6_, x916x, x905x, n_n258}, n_n7441);
	defparam lut_2789.LUT_SIZE = 7;
	defparam lut_2789.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_2791 ({sk[612], i_7_, i_8_, i_6_, x916x, x899x, n_n228}, n_n7440);
	defparam lut_2791.LUT_SIZE = 7;
	defparam lut_2791.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_2793 ({sk[613], n_n281, n_n208, x916x, n_n220, x905x, x899x}, x446x);
	defparam lut_2793.LUT_SIZE = 7;
	defparam lut_2793.mask = 128'h5555ffff5555ffff0000000500000037;

	lut_sub lut_2796 ({sk[614], i_14_, i_13_, i_12_, x913x, x911x}, x1541x);
	defparam lut_2796.LUT_SIZE = 6;
	defparam lut_2796.mask = 64'h3f3f3f3f30500305;

	lut_sub lut_2801 ({sk[615], n_n4, n_n7, n_n7441, n_n7440, x446x, x1541x}, n_n2839);
	defparam lut_2801.LUT_SIZE = 7;
	defparam lut_2801.mask = 128'h5555ffff5555ffff3fff3fff7fffffff;

	lut_sub lut_2807 ({sk[616], i_9_, i_10_, i_11_, i_15_}, x901x);
	defparam lut_2807.LUT_SIZE = 5;
	defparam lut_2807.mask = 32'h0f0f4000;

	lut_sub lut_2809 ({sk[617], i_14_, i_13_, i_12_, x907x, x914x, x901x}, x410x);
	defparam lut_2809.LUT_SIZE = 7;
	defparam lut_2809.mask = 128'h5555ffff5555ffff33000000000f0055;

	lut_sub lut_2813 ({sk[618], i_14_, i_13_, i_12_, x906x}, n_n12);
	defparam lut_2813.LUT_SIZE = 5;
	defparam lut_2813.mask = 32'h0f0f4000;

	lut_sub lut_2815 ({sk[619], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, n_n5682);
	defparam lut_2815.LUT_SIZE = 7;
	defparam lut_2815.mask = 128'h5555ffff5555ffff0000100000000000;

	lut_sub lut_2817 ({sk[620], n_n281, n_n130, n_n122, x911x, x899x, x912x}, x20630x);
	defparam lut_2817.LUT_SIZE = 7;
	defparam lut_2817.mask = 128'h5555ffff5555ffff00000000007f7f7f;

	lut_sub lut_2824 ({sk[621], i_14_, i_13_, i_12_, x912x}, n_n135);
	defparam lut_2824.LUT_SIZE = 5;
	defparam lut_2824.mask = 32'h0f0f4000;

	lut_sub lut_2826 ({sk[622], i_7_, i_5_, i_6_, i_3_, i_4_, n_n118}, x4238x);
	defparam lut_2826.LUT_SIZE = 7;
	defparam lut_2826.mask = 128'h5555ffff5555ffff0000000050005000;

	lut_sub lut_2831 ({sk[623], i_7_, i_8_, i_6_, x917x, n_n165, n_n284}, x1784x);
	defparam lut_2831.LUT_SIZE = 7;
	defparam lut_2831.mask = 128'h5555ffff5555ffff1f1f000000000000;

	lut_sub lut_2836 ({sk[624], i_9_, i_10_, i_7_, i_8_, i_6_, x917x}, x20639x);
	defparam lut_2836.LUT_SIZE = 7;
	defparam lut_2836.mask = 128'h5555ffff5555ffff5000000000000000;

	lut_sub lut_2839 ({sk[625], i_9_, i_10_, i_11_, i_15_, n_n281}, x216x);
	defparam lut_2839.LUT_SIZE = 6;
	defparam lut_2839.mask = 64'h3f3f3f3f00101000;

	lut_sub lut_2842 ({sk[626], i_14_, i_13_, i_12_, x913x, n_n273, x909x}, x515x);
	defparam lut_2842.LUT_SIZE = 7;
	defparam lut_2842.mask = 128'h5555ffff5555ffff0000000001000000;

	lut_sub lut_2844 ({sk[627], i_7_, i_8_, i_6_, x909x, x905x, n_n279}, x569x);
	defparam lut_2844.LUT_SIZE = 7;
	defparam lut_2844.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_2846 ({sk[628], i_14_, i_13_, i_12_, x907x, n_n273, x909x}, x872x);
	defparam lut_2846.LUT_SIZE = 7;
	defparam lut_2846.mask = 128'h5555ffff5555ffff0000000001000000;

	lut_sub lut_2848 ({sk[629], i_7_, i_8_, i_6_, x914x, x909x, n_n279}, x894x);
	defparam lut_2848.LUT_SIZE = 7;
	defparam lut_2848.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_2850 ({sk[630], x372x, x515x, x569x, x872x, x875x, x894x}, n_n4186);
	defparam lut_2850.LUT_SIZE = 7;
	defparam lut_2850.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_2857 ({sk[631], i_14_, i_13_, i_12_, x898x}, n_n54);
	defparam lut_2857.LUT_SIZE = 5;
	defparam lut_2857.mask = 32'h0f0f0010;

	lut_sub lut_2859 ({sk[632], i_14_, i_13_, i_12_, x900x}, n_n105);
	defparam lut_2859.LUT_SIZE = 5;
	defparam lut_2859.mask = 32'h0f0f0010;

	lut_sub lut_2861 ({sk[633], i_14_, i_13_, i_12_, x899x}, n_n197);
	defparam lut_2861.LUT_SIZE = 5;
	defparam lut_2861.mask = 32'h0f0f0010;

	lut_sub lut_2863 ({sk[634], i_14_, i_13_, i_12_}, n_n258);
	defparam lut_2863.LUT_SIZE = 4;
	defparam lut_2863.mask = 16'h5504;

	lut_sub lut_2865 ({sk[635], i_7_, i_8_, i_6_, x909x}, n_n177);
	defparam lut_2865.LUT_SIZE = 5;
	defparam lut_2865.mask = 32'h0f0f0400;

	lut_sub lut_2867 ({sk[636], x915x, n_n266, x911x, n_n258, n_n45, n_n177}, x559x);
	defparam lut_2867.LUT_SIZE = 7;
	defparam lut_2867.mask = 128'h5555ffff5555ffff111111111111111f;

	lut_sub lut_2870 ({sk[637], i_9_, i_10_, i_11_, i_15_}, x897x);
	defparam lut_2870.LUT_SIZE = 5;
	defparam lut_2870.mask = 32'h0f0f1000;

	lut_sub lut_2872 ({sk[638], i_14_, i_13_, i_12_, x901x}, n_n104);
	defparam lut_2872.LUT_SIZE = 5;
	defparam lut_2872.mask = 32'h0f0f0010;

	lut_sub lut_2874 ({sk[639], i_9_, i_10_, i_11_, i_15_}, x902x);
	defparam lut_2874.LUT_SIZE = 5;
	defparam lut_2874.mask = 32'h0f0f0010;

	lut_sub lut_2876 ({sk[640], i_14_, i_13_, i_12_, x912x}, n_n41);
	defparam lut_2876.LUT_SIZE = 5;
	defparam lut_2876.mask = 32'h0f0f0010;

	lut_sub lut_2878 ({sk[641], i_14_, i_13_, i_12_, x898x}, x99x);
	defparam lut_2878.LUT_SIZE = 5;
	defparam lut_2878.mask = 32'h0f0f5100;

	lut_sub lut_2882 ({sk[642], x909x, n_n261, n_n263, x224x, x904x, n_n225}, x708x);
	defparam lut_2882.LUT_SIZE = 7;
	defparam lut_2882.mask = 128'h5555ffff5555ffff00000000000f111f;

	lut_sub lut_2885 ({sk[643], n_n6, n_n5796, x5037x, x389x, x632x, x1911x}, x20675x);
	defparam lut_2885.LUT_SIZE = 7;
	defparam lut_2885.mask = 128'h5555ffff5555ffff3fffffff7fffffff;

	lut_sub lut_2891 ({sk[644], x909x, n_n261, n_n4251, x99x, x708x, x20675x}, n_n4211);
	defparam lut_2891.LUT_SIZE = 7;
	defparam lut_2891.mask = 128'h5555ffff5555ffff77ff77ff77ff7fff;

	lut_sub lut_2896 ({sk[645], n_n6, n_n5, x153x, x166x, x224x, x1895x}, x20680x);
	defparam lut_2896.LUT_SIZE = 7;
	defparam lut_2896.mask = 128'h5555ffff5555ffff00000f0f77ff7fff;

	lut_sub lut_2901 ({sk[646], n_n266, n_n271, x909x, x734x, n_n60, x137x}, x20682x);
	defparam lut_2901.LUT_SIZE = 7;
	defparam lut_2901.mask = 128'h5555ffff5555ffff0f0f0f5f0f3f0f7f;

	lut_sub lut_2905 ({sk[647], n_n5, x1907x, x1908x, n_n4892, x5021x, x5022x}, x24123x);
	defparam lut_2905.LUT_SIZE = 7;
	defparam lut_2905.mask = 128'h5555ffff5555ffff8080808080000000;

	lut_sub lut_2908 ({sk[648], x20680x, x488x, x878x, x20682x, x24123x}, x20686x);
	defparam lut_2908.LUT_SIZE = 6;
	defparam lut_2908.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_2914 ({sk[649], n_n111, x909x, n_n261, x5376x, x189x, x616x}, x20689x);
	defparam lut_2914.LUT_SIZE = 7;
	defparam lut_2914.mask = 128'h5555ffff5555ffff5f5f5f7f5f5f5fff;

	lut_sub lut_2919 ({sk[650], n_n6, n_n5, x99x, x19862x, x1894x, x1859x}, x20690x);
	defparam lut_2919.LUT_SIZE = 7;
	defparam lut_2919.mask = 128'h5555ffff5555ffff0f0f3fff5f5f7fff;

	lut_sub lut_2924 ({sk[651], x19753x, x19754x, x19755x, x19756x, x20689x, x20690x}, n_n4197);
	defparam lut_2924.LUT_SIZE = 7;
	defparam lut_2924.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_2931 ({sk[652], n_n56, n_n4959, x254x, n_n4960, n_n4952, x20710x}, n_n4219);
	defparam lut_2931.LUT_SIZE = 7;
	defparam lut_2931.mask = 128'h5555ffff5555ffff7f7fffff7fffffff;

	lut_sub lut_2937 ({sk[653], x20703x, x20704x, n_n4280, n_n4279, x20715x}, x20718x);
	defparam lut_2937.LUT_SIZE = 6;
	defparam lut_2937.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_2943 ({sk[654], x562x, x4998x, x555x, n_n4261, n_n4256, x465x}, x20733x);
	defparam lut_2943.LUT_SIZE = 7;
	defparam lut_2943.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_2950 ({sk[655], n_n4259, x721x, x20729x, x24187x}, x20734x);
	defparam lut_2950.LUT_SIZE = 5;
	defparam lut_2950.mask = 32'h0f0fbfff;

	lut_sub lut_2955 ({sk[656], n_n57, x165x, n_n4941, n_n4942, n_n4938, x20740x}, x20741x);
	defparam lut_2955.LUT_SIZE = 7;
	defparam lut_2955.mask = 128'h5555ffff5555ffff7fff7fff7fffffff;

	lut_sub lut_2961 ({sk[657], x20698x, x20723x, x20724x, x20696x, x20697x}, x20742x);
	defparam lut_2961.LUT_SIZE = 6;
	defparam lut_2961.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_2967 ({sk[658], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x910x);
	defparam lut_2967.LUT_SIZE = 7;
	defparam lut_2967.mask = 128'h5555ffff5555ffff0000080000000000;

	lut_sub lut_2969 ({sk[659], i_14_, i_13_, i_12_, n_n3, x904x}, n_n7407);
	defparam lut_2969.LUT_SIZE = 6;
	defparam lut_2969.mask = 64'h3f3f3f3f10000000;

	lut_sub lut_2971 ({sk[660], i_14_, i_13_, i_12_, n_n3, x898x, x904x}, x409x);
	defparam lut_2971.LUT_SIZE = 7;
	defparam lut_2971.mask = 128'h5555ffff5555ffff0000030000050000;

	lut_sub lut_2974 ({sk[661], i_14_, i_13_, i_12_, n_n3, x914x, x912x}, x3937x);
	defparam lut_2974.LUT_SIZE = 7;
	defparam lut_2974.mask = 128'h5555ffff5555ffff0000000000030005;

	lut_sub lut_2977 ({sk[662], n_n148, n_n4, x206x, n_n7407, x409x, x3937x}, n_n3140);
	defparam lut_2977.LUT_SIZE = 7;
	defparam lut_2977.mask = 128'h5555ffff5555ffff7f7f7fff7f7fffff;

	lut_sub lut_2983 ({sk[663], i_7_, i_8_, i_6_, x916x, n_n228, x902x}, n_n7424);
	defparam lut_2983.LUT_SIZE = 7;
	defparam lut_2983.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_2985 ({sk[664], i_7_, i_8_, i_6_, x916x}, n_n3);
	defparam lut_2985.LUT_SIZE = 5;
	defparam lut_2985.mask = 32'h0f0f1000;

	lut_sub lut_2987 ({sk[665], i_7_, i_8_, i_6_, n_n281, x916x, x908x}, x439x);
	defparam lut_2987.LUT_SIZE = 7;
	defparam lut_2987.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_2989 ({sk[666], i_14_, i_13_, i_12_, x908x}, n_n61);
	defparam lut_2989.LUT_SIZE = 5;
	defparam lut_2989.mask = 32'h0f0f0010;

	lut_sub lut_2991 ({sk[667], i_9_, i_10_, i_11_}, n_n270);
	defparam lut_2991.LUT_SIZE = 4;
	defparam lut_2991.mask = 16'h5504;

	lut_sub lut_2993 ({sk[668], x915x, n_n273, n_n283, n_n108, x82x, x1932x}, n_n3155);
	defparam lut_2993.LUT_SIZE = 7;
	defparam lut_2993.mask = 128'h5555ffff5555ffff0000000000770f7f;

	lut_sub lut_2997 ({sk[669], i_14_, i_13_, i_12_, i_15_, n_n247, x44x}, x1027x);
	defparam lut_2997.LUT_SIZE = 7;
	defparam lut_2997.mask = 128'h5555ffff5555ffff7555575555755557;

	lut_sub lut_3003 ({sk[670], i_14_, i_13_, i_12_, i_15_, x160x, n_n253}, x1026x);
	defparam lut_3003.LUT_SIZE = 7;
	defparam lut_3003.mask = 128'h5555ffff5555ffff7333373333733337;

	lut_sub lut_3009 ({sk[671], x915x, n_n273, n_n283, n_n108, x258x, x70x}, x20941x);
	defparam lut_3009.LUT_SIZE = 7;
	defparam lut_3009.mask = 128'h5555ffff5555ffff00000000003f557f;

	lut_sub lut_3013 ({sk[672], n_n1, x5159x, x209x, x739x, x1023x, x118x}, x20931x);
	defparam lut_3013.LUT_SIZE = 7;
	defparam lut_3013.mask = 128'h5555ffff5555ffff0f0fffff7fffffff;

	lut_sub lut_3019 ({sk[673], n_n2, n_n268, n_n3246, x146x, x20928x, x1326x}, x20932x);
	defparam lut_3019.LUT_SIZE = 7;
	defparam lut_3019.mask = 128'h5555ffff5555ffff00ff55ff3fff7fff;

	lut_sub lut_3024 ({sk[674], x916x, n_n271, n_n3, x1025x, x45x, x171x}, x20936x);
	defparam lut_3024.LUT_SIZE = 7;
	defparam lut_3024.mask = 128'h5555ffff5555ffff0077007700770f7f;

	lut_sub lut_3028 ({sk[675], n_n4, n_n3, n_n95, x68x, x1283x, x598x}, x20937x);
	defparam lut_3028.LUT_SIZE = 7;
	defparam lut_3028.mask = 128'h5555ffff5555ffff55555f5f7fff7fff;

	lut_sub lut_3034 ({sk[676], i_14_, i_13_, i_12_, x905x, x899x}, x159x);
	defparam lut_3034.LUT_SIZE = 6;
	defparam lut_3034.mask = 64'h3f3f3f3f30500300;

	lut_sub lut_3038 ({sk[677], i_7_, i_6_, x916x, n_n226, n_n7441}, x24209x);
	defparam lut_3038.LUT_SIZE = 6;
	defparam lut_3038.mask = 64'h3f3f3f3faaa8aaaa;

	lut_sub lut_3043 ({sk[678], n_n281, n_n3, x159x, x908x, x446x, x24209x}, n_n3138);
	defparam lut_3043.LUT_SIZE = 7;
	defparam lut_3043.mask = 128'h5555ffff5555ffffbbbbbbffbbbbbfff;

	lut_sub lut_3048 ({sk[679], n_n4, n_n3, n_n76, x485x, x80x, n_n7306}, x21136x);
	defparam lut_3048.LUT_SIZE = 7;
	defparam lut_3048.mask = 128'h5555ffff5555ffff5f5f5fff7fff7fff;

	lut_sub lut_3054 ({sk[680], n_n208, x916x, n_n220, n_n3, x905x, x70x}, n_n3229);
	defparam lut_3054.LUT_SIZE = 7;
	defparam lut_3054.mask = 128'h5555ffff5555ffff0003000300035557;

	lut_sub lut_3057 ({sk[681], n_n208, x916x, n_n3, n_n70, x1240x, x1854x}, x21147x);
	defparam lut_3057.LUT_SIZE = 7;
	defparam lut_3057.mask = 128'h5555ffff5555ffff0033003300335f7f;

	lut_sub lut_3061 ({sk[682], n_n3, n_n7355, x867x, x979x, n_n15, x742x}, x24119x);
	defparam lut_3061.LUT_SIZE = 7;
	defparam lut_3061.mask = 128'h5555ffff5555ffffaa00000080000000;

	lut_sub lut_3064 ({sk[683], i_14_, i_13_, i_12_, x914x, x912x}, x184x);
	defparam lut_3064.LUT_SIZE = 6;
	defparam lut_3064.mask = 64'h3f3f3f3f30500000;

	lut_sub lut_3067 ({sk[684], i_14_, i_13_, i_12_, i_15_, x908x, n_n270}, x63x);
	defparam lut_3067.LUT_SIZE = 7;
	defparam lut_3067.mask = 128'h5555ffff5555ffff0000050000330000;

	lut_sub lut_3070 ({sk[685], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x953x);
	defparam lut_3070.LUT_SIZE = 7;
	defparam lut_3070.mask = 128'h5555ffff5555ffff4000110000040001;

	lut_sub lut_3076 ({sk[686], n_n139, x48x, n_n110, n_n127, x299x, x1844x}, x21167x);
	defparam lut_3076.LUT_SIZE = 7;
	defparam lut_3076.mask = 128'h5555ffff5555ffff030f0f0f575f5f5f;

	lut_sub lut_3081 ({sk[687], x211x, x48x, n_n124, n_n5769, n_n111, n_n132}, x21166x);
	defparam lut_3081.LUT_SIZE = 7;
	defparam lut_3081.mask = 128'h5555ffff5555ffff1f3f5f7f5fff5fff;

	lut_sub lut_3088 ({sk[688], i_14_, i_13_, i_12_, n_n208, x916x, x905x}, n_n7355);
	defparam lut_3088.LUT_SIZE = 7;
	defparam lut_3088.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_3090 ({sk[689], i_14_, i_13_, i_12_, n_n283, x914x, x922x}, x373x);
	defparam lut_3090.LUT_SIZE = 7;
	defparam lut_3090.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_3092 ({sk[690], i_7_, i_8_, i_6_, x916x, x111x}, n_n3506);
	defparam lut_3092.LUT_SIZE = 6;
	defparam lut_3092.mask = 64'h3f3f3f3f00010000;

	lut_sub lut_3094 ({sk[691], n_n4, n_n76, x485x, x80x, n_n7306, x455x}, x21183x);
	defparam lut_3094.LUT_SIZE = 7;
	defparam lut_3094.mask = 128'h5555ffff5555ffff77ff77ff7fffffff;

	lut_sub lut_3100 ({sk[692], n_n7355, x867x, x373x, n_n3506, x378x, x21183x}, x21186x);
	defparam lut_3100.LUT_SIZE = 7;
	defparam lut_3100.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_3107 ({sk[693], x21228x, x21229x, x533x, n_n3909, x21233x, x21234x}, n_n3895);
	defparam lut_3107.LUT_SIZE = 7;
	defparam lut_3107.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_3114 ({sk[694], n_n3, n_n59, x156x, x21189x, x21239x, x21240x}, x21243x);
	defparam lut_3114.LUT_SIZE = 7;
	defparam lut_3114.mask = 128'h5555ffff5555ffff7f7f7f7f7fffffff;

	lut_sub lut_3120 ({sk[695], n_n3929, n_n3406, n_n3932, x21201x, x21200x}, x21244x);
	defparam lut_3120.LUT_SIZE = 6;
	defparam lut_3120.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_3126 ({sk[696], n_n208, x916x, n_n3, x1502x, x1524x, x1523x}, x24116x);
	defparam lut_3126.LUT_SIZE = 7;
	defparam lut_3126.mask = 128'h5555ffff5555ffffffc0ffc0ffc0aa80;

	lut_sub lut_3133 ({sk[697], n_n3, n_n216, x333x, n_n2986, n_n7344, x1436x}, x24117x);
	defparam lut_3133.LUT_SIZE = 7;
	defparam lut_3133.mask = 128'h5555ffff5555ffffc000c00080000000;

	lut_sub lut_3136 ({sk[698], n_n4, n_n103, n_n876, x3678x, x1435x, x117x}, x24202x);
	defparam lut_3136.LUT_SIZE = 7;
	defparam lut_3136.mask = 128'h5555ffff5555fffff000f00080000000;

	lut_sub lut_3139 ({sk[699], n_n208, x916x, n_n220, x906x, x5762x, x98x}, x19390x);
	defparam lut_3139.LUT_SIZE = 7;
	defparam lut_3139.mask = 128'h5555ffff5555ffff333333333333777f;

	lut_sub lut_3143 ({sk[700], n_n208, x916x, n_n3, x45x, x171x, x1924x}, x19391x);
	defparam lut_3143.LUT_SIZE = 7;
	defparam lut_3143.mask = 128'h5555ffff5555ffff003f003f003f557f;

	lut_sub lut_3147 ({sk[701], x439x, x648x, x557x, n_n7440, n_n7442}, x21263x);
	defparam lut_3147.LUT_SIZE = 6;
	defparam lut_3147.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_3153 ({sk[702], x19390x, x19391x, x21263x}, x21264x);
	defparam lut_3153.LUT_SIZE = 4;
	defparam lut_3153.mask = 16'h557f;

	lut_sub lut_3157 ({sk[703], x916x, n_n271, x136x, x50x, x377x, x24115x}, x3626x);
	defparam lut_3157.LUT_SIZE = 7;
	defparam lut_3157.mask = 128'h5555ffff5555ffff000000000000bfff;

	lut_sub lut_3162 ({sk[704], n_n110, n_n268, n_n22, x779x, x55x, x1480x}, x21283x);
	defparam lut_3162.LUT_SIZE = 7;
	defparam lut_3162.mask = 128'h5555ffff5555ffff0f0f7fff0f0fffff;

	lut_sub lut_3168 ({sk[705], x916x, n_n271, n_n240, x160x, n_n147, n_n59}, x3629x);
	defparam lut_3168.LUT_SIZE = 7;
	defparam lut_3168.mask = 128'h5555ffff5555ffff0000000000007fff;

	lut_sub lut_3173 ({sk[706], n_n106, n_n265, n_n4, n_n54, n_n62, x598x}, x21270x);
	defparam lut_3173.LUT_SIZE = 7;
	defparam lut_3173.mask = 128'h5555ffff5555ffff555f777f555fffff;

	lut_sub lut_3178 ({sk[707], i_7_, i_8_, i_6_, x916x, x101x, x1481x}, x24114x);
	defparam lut_3178.LUT_SIZE = 7;
	defparam lut_3178.mask = 128'h5555ffff5555fffffffffffffffffff8;

	lut_sub lut_3184 ({sk[708], x3626x, x21283x, x3629x, x21270x, x24114x}, x21291x);
	defparam lut_3184.LUT_SIZE = 6;
	defparam lut_3184.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_3190 ({sk[709], i_14_, i_13_, i_12_, i_15_, n_n267, x138x}, x1461x);
	defparam lut_3190.LUT_SIZE = 7;
	defparam lut_3190.mask = 128'h5555ffff5555ffff5575755777557775;

	lut_sub lut_3200 ({sk[710], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1460x);
	defparam lut_3200.LUT_SIZE = 7;
	defparam lut_3200.mask = 128'h5555ffff5555ffff0101000505000504;

	lut_sub lut_3210 ({sk[711], n_n208, x916x, n_n3, n_n105, n_n896, x77x}, x21288x);
	defparam lut_3210.LUT_SIZE = 7;
	defparam lut_3210.mask = 128'h5555ffff5555ffff333f333f333f7f7f;

	lut_sub lut_3215 ({sk[712], i_14_, i_13_, i_12_, x899x}, n_n226);
	defparam lut_3215.LUT_SIZE = 5;
	defparam lut_3215.mask = 32'h0f0f0001;

	lut_sub lut_3217 ({sk[713], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1155x);
	defparam lut_3217.LUT_SIZE = 7;
	defparam lut_3217.mask = 128'h5555ffff5555ffff4000100000400010;

	lut_sub lut_3222 ({sk[714], n_n151, x183x, n_n57, n_n56, n_n226, x1155x}, n_n2440);
	defparam lut_3222.LUT_SIZE = 7;
	defparam lut_3222.mask = 128'h5555ffff5555ffff03570f5f0f5f0f5f;

	lut_sub lut_3227 ({sk[715], n_n197, n_n57, n_n56, x62x, x481x, x1789x}, n_n2433);
	defparam lut_3227.LUT_SIZE = 7;
	defparam lut_3227.mask = 128'h5555ffff5555ffff337f7f7f33ff7fff;

	lut_sub lut_3234 ({sk[716], n_n281, n_n266, x206x, x914x, x909x, x1807x}, x21330x);
	defparam lut_3234.LUT_SIZE = 7;
	defparam lut_3234.mask = 128'h5555ffff5555ffff0000113300001333;

	lut_sub lut_3238 ({sk[717], i_7_, i_8_, i_6_, x909x, n_n2442, x1808x}, x21331x);
	defparam lut_3238.LUT_SIZE = 7;
	defparam lut_3238.mask = 128'h5555ffff5555ffff3333333333373333;

	lut_sub lut_3241 ({sk[718], i_14_, i_13_, i_12_, i_15_, x176x, n_n259}, x1848x);
	defparam lut_3241.LUT_SIZE = 7;
	defparam lut_3241.mask = 128'h5555ffff5555ffff3777737777337773;

	lut_sub lut_3254 ({sk[719], n_n12, n_n57, n_n56, x121x, n_n15, x1764x}, x21356x);
	defparam lut_3254.LUT_SIZE = 7;
	defparam lut_3254.mask = 128'h5555ffff5555ffff003f7f7f00ff7fff;

	lut_sub lut_3261 ({sk[720], i_14_, i_13_, i_12_, x908x, x902x}, x199x);
	defparam lut_3261.LUT_SIZE = 6;
	defparam lut_3261.mask = 64'h3f3f3f3f00000305;

	lut_sub lut_3264 ({sk[721], i_14_, i_13_, i_12_, i_15_, x199x, n_n270}, x21361x);
	defparam lut_3264.LUT_SIZE = 7;
	defparam lut_3264.mask = 128'h5555ffff5555ffff7333373333333333;

	lut_sub lut_3268 ({sk[722], i_9_, i_10_, i_11_, i_15_}, x903x);
	defparam lut_3268.LUT_SIZE = 5;
	defparam lut_3268.mask = 32'h0f0f2000;

	lut_sub lut_3270 ({sk[723], i_14_, i_13_, i_12_}, n_n279);
	defparam lut_3270.LUT_SIZE = 4;
	defparam lut_3270.mask = 16'h5508;

	lut_sub lut_3272 ({sk[724], i_14_, i_13_, i_12_, x903x}, x40x);
	defparam lut_3272.LUT_SIZE = 5;
	defparam lut_3272.mask = 32'h0f0f1400;

	lut_sub lut_3275 ({sk[725], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x150x);
	defparam lut_3275.LUT_SIZE = 7;
	defparam lut_3275.mask = 128'h5555ffff5555ffff0100000404000000;

	lut_sub lut_3279 ({sk[726], n_n4, n_n279, x40x, x899x, x150x, x897x}, x21372x);
	defparam lut_3279.LUT_SIZE = 7;
	defparam lut_3279.mask = 128'h5555ffff5555ffff0000000033ff7fff;

	lut_sub lut_3284 ({sk[727], i_14_, i_13_, i_12_, x905x, x899x}, x307x);
	defparam lut_3284.LUT_SIZE = 6;
	defparam lut_3284.mask = 64'h3f3f3f3f50033000;

	lut_sub lut_3288 ({sk[728], i_14_, i_13_, i_12_, n_n208, x916x, x905x}, x333x);
	defparam lut_3288.LUT_SIZE = 7;
	defparam lut_3288.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_3291 ({sk[729], i_14_, i_13_, i_12_, x913x, x911x}, x987x);
	defparam lut_3291.LUT_SIZE = 6;
	defparam lut_3291.mask = 64'h3f3f3f3f50037000;

	lut_sub lut_3296 ({sk[730], i_14_, i_13_, i_12_, i_15_, x21371x, n_n270}, x989x);
	defparam lut_3296.LUT_SIZE = 7;
	defparam lut_3296.mask = 128'h5555ffff5555ffff3773737373333333;

	lut_sub lut_3303 ({sk[731], n_n4, n_n3, x307x, x333x, x987x, x989x}, x21373x);
	defparam lut_3303.LUT_SIZE = 7;
	defparam lut_3303.mask = 128'h5555ffff5555ffff0f0f7f7f0fff7fff;

	lut_sub lut_3308 ({sk[732], n_n208, x916x, n_n220, x908x, n_n256, x24158x}, n_n2104);
	defparam lut_3308.LUT_SIZE = 7;
	defparam lut_3308.mask = 128'h5555ffff5555ffffaaaaaaaaaaaaabaf;

	lut_sub lut_3312 ({sk[733], i_14_, i_13_, i_12_, i_15_, n_n247, x1037x}, x1036x);
	defparam lut_3312.LUT_SIZE = 7;
	defparam lut_3312.mask = 128'h5555ffff5555ffff5755557577555555;

	lut_sub lut_3318 ({sk[734], i_14_, i_13_, i_12_, n_n3, x904x}, x476x);
	defparam lut_3318.LUT_SIZE = 6;
	defparam lut_3318.mask = 64'h3f3f3f3f01100000;

	lut_sub lut_3321 ({sk[735], i_14_, i_13_, i_12_, i_15_, n_n253, n_n267}, x1040x);
	defparam lut_3321.LUT_SIZE = 7;
	defparam lut_3321.mask = 128'h5555ffff5555ffff0700007075000000;

	lut_sub lut_3329 ({sk[736], i_14_, i_13_, i_12_, n_n4, x914x, x1037x}, x3530x);
	defparam lut_3329.LUT_SIZE = 7;
	defparam lut_3329.mask = 128'h5555ffff5555ffff0507070505050505;

	lut_sub lut_3333 ({sk[737], n_n3, n_n2104, x1036x, x476x, x1040x, x3530x}, x21396x);
	defparam lut_3333.LUT_SIZE = 7;
	defparam lut_3333.mask = 128'h5555ffff5555ffff5f5fffff7fffffff;

	lut_sub lut_3339 ({sk[738], n_n106, n_n265, n_n4, n_n186, x598x, x3526x}, n_n2110);
	defparam lut_3339.LUT_SIZE = 7;
	defparam lut_3339.mask = 128'h5555ffff5555ffff777f777f777fffff;

	lut_sub lut_3344 ({sk[739], n_n265, x252x, n_n32, x765x, x934x, x205x}, x21387x);
	defparam lut_3344.LUT_SIZE = 7;
	defparam lut_3344.mask = 128'h5555ffff5555ffff3f3f3f3f7fffffff;

	lut_sub lut_3350 ({sk[740], x916x, n_n271, x90x, x329x, x46x, x327x}, x3521x);
	defparam lut_3350.LUT_SIZE = 7;
	defparam lut_3350.mask = 128'h5555ffff5555ffff0000000000007fff;

	lut_sub lut_3355 ({sk[741], n_n4, n_n3, x51x, n_n93, x467x, x1041x}, x21395x);
	defparam lut_3355.LUT_SIZE = 7;
	defparam lut_3355.mask = 128'h5555ffff5555ffff333333ff7f7f7fff;

	lut_sub lut_3360 ({sk[742], n_n2110, x21387x, x3521x, x21395x}, x21397x);
	defparam lut_3360.LUT_SIZE = 5;
	defparam lut_3360.mask = 32'h0f0f7fff;

	lut_sub lut_3365 ({sk[743], i_14_, i_13_, i_12_, x905x}, n_n145);
	defparam lut_3365.LUT_SIZE = 5;
	defparam lut_3365.mask = 32'h0f0f4000;

	lut_sub lut_3367 ({sk[744], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x157x);
	defparam lut_3367.LUT_SIZE = 7;
	defparam lut_3367.mask = 128'h5555ffff5555ffff0040404000000000;

	lut_sub lut_3371 ({sk[745], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x21414x);
	defparam lut_3371.LUT_SIZE = 7;
	defparam lut_3371.mask = 128'h5555ffff5555ffff0144444405000000;

	lut_sub lut_3381 ({sk[746], i_14_, i_13_, i_12_, i_15_, n_n282, n_n270}, x1102x);
	defparam lut_3381.LUT_SIZE = 7;
	defparam lut_3381.mask = 128'h5555ffff5555ffff0770707077000000;

	lut_sub lut_3394 ({sk[747], i_14_, i_13_, i_12_, x914x, x912x}, x330x);
	defparam lut_3394.LUT_SIZE = 6;
	defparam lut_3394.mask = 64'h3f3f3f3f50007000;

	lut_sub lut_3398 ({sk[748], n_n1, n_n2, x157x, x21414x, x1102x, x330x}, x21415x);
	defparam lut_3398.LUT_SIZE = 7;
	defparam lut_3398.mask = 128'h5555ffff5555ffff00005fff33337fff;

	lut_sub lut_3403 ({sk[749], i_7_, i_8_, i_6_, x915x}, x135x);
	defparam lut_3403.LUT_SIZE = 5;
	defparam lut_3403.mask = 32'h0f0f4400;

	lut_sub lut_3406 ({sk[750], x915x, n_n273, n_n268, n_n145, x264x, x24104x}, n_n2113);
	defparam lut_3406.LUT_SIZE = 7;
	defparam lut_3406.mask = 128'h5555ffff5555ffffaabbaabbaabbafbf;

	lut_sub lut_3410 ({sk[751], x915x, n_n273, n_n283, x21401x, x21402x, x1097x}, n_n2075);
	defparam lut_3410.LUT_SIZE = 7;
	defparam lut_3410.mask = 128'h5555ffff5555ffff0000000000553f7f;

	lut_sub lut_3414 ({sk[752], n_n1, n_n2, x1101x, x21407x, x281x, x338x}, x21409x);
	defparam lut_3414.LUT_SIZE = 7;
	defparam lut_3414.mask = 128'h5555ffff5555ffff000077ff0fff7fff;

	lut_sub lut_3420 ({sk[753], n_n12, x21415x, x135x, n_n2113, n_n2075, x21409x}, n_n2061);
	defparam lut_3420.LUT_SIZE = 7;
	defparam lut_3420.mask = 128'h5555ffff5555ffff7f7fffff7fffffff;

	lut_sub lut_3426 ({sk[754], x915x, n_n273, n_n283, x1159x, x21422x, x24109x}, n_n2077);
	defparam lut_3426.LUT_SIZE = 7;
	defparam lut_3426.mask = 128'h5555ffff5555ffff0000000000bb0fbf;

	lut_sub lut_3430 ({sk[755], n_n208, x916x, n_n279, x900x, x333x, x467x}, n_n2129);
	defparam lut_3430.LUT_SIZE = 7;
	defparam lut_3430.mask = 128'h5555ffff5555ffff777777777777777f;

	lut_sub lut_3434 ({sk[756], n_n4, n_n12, n_n7407, x466x, x476x, n_n7443}, x21431x);
	defparam lut_3434.LUT_SIZE = 7;
	defparam lut_3434.mask = 128'h5555ffff5555ffff7fff7fff7fffffff;

	lut_sub lut_3440 ({sk[757], n_n208, x916x, n_n109, x79x, x296x, x21430x}, x21432x);
	defparam lut_3440.LUT_SIZE = 7;
	defparam lut_3440.mask = 128'h5555ffff5555ffff5555555555557fff;

	lut_sub lut_3445 ({sk[758], x915x, n_n273, n_n6868, n_n6856, n_n2274, x1162x}, x21438x);
	defparam lut_3445.LUT_SIZE = 7;
	defparam lut_3445.mask = 128'h5555ffff5555ffff3fff3fff3fff7fff;

	lut_sub lut_3450 ({sk[759], n_n106, n_n2, x78x, n_n2272, x1029x, x24108x}, x21439x);
	defparam lut_3450.LUT_SIZE = 7;
	defparam lut_3450.mask = 128'h5555ffff5555ffffafafbfffafafffff;

	lut_sub lut_3456 ({sk[760], n_n2077, n_n2129, x21431x, x21432x, x21438x, x21439x}, n_n2062);
	defparam lut_3456.LUT_SIZE = 7;
	defparam lut_3456.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_3463 ({sk[761], x915x, n_n263, x119x, x167x, x21477x, x21479x}, n_n2095);
	defparam lut_3463.LUT_SIZE = 7;
	defparam lut_3463.mask = 128'h5555ffff5555ffff5555555555557fff;

	lut_sub lut_3468 ({sk[762], i_7_, i_8_, i_6_, x915x, x1416x, x330x}, n_n2097);
	defparam lut_3468.LUT_SIZE = 7;
	defparam lut_3468.mask = 128'h5555ffff5555ffff0000000003000700;

	lut_sub lut_3472 ({sk[763], i_14_, i_13_, i_12_, i_15_, n_n282, n_n247}, x1418x);
	defparam lut_3472.LUT_SIZE = 7;
	defparam lut_3472.mask = 128'h5555ffff5555ffff0370707033000000;

	lut_sub lut_3482 ({sk[764], n_n280, n_n100, n_n32, x391x, x1417x, x24111x}, x21511x);
	defparam lut_3482.LUT_SIZE = 7;
	defparam lut_3482.mask = 128'h5555ffff5555ffffafafbfffafafffff;

	lut_sub lut_3488 ({sk[765], x915x, n_n263, n_n2095, n_n2097, x1418x, x21511x}, x21514x);
	defparam lut_3488.LUT_SIZE = 7;
	defparam lut_3488.mask = 128'h5555ffff5555ffff5fff5fff5fff7fff;

	lut_sub lut_3493 ({sk[766], n_n56, x520x, n_n2169, x205x, x21464x, x24186x}, x21470x);
	defparam lut_3493.LUT_SIZE = 7;
	defparam lut_3493.mask = 128'h5555ffff5555ffff55ffffff7fffffff;

	lut_sub lut_3499 ({sk[767], n_n2172, x21453x, x21462x, x21463x, x21452x}, x21471x);
	defparam lut_3499.LUT_SIZE = 6;
	defparam lut_3499.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_3505 ({sk[768], n_n2166, x21504x, x21505x}, x21507x);
	defparam lut_3505.LUT_SIZE = 4;
	defparam lut_3505.mask = 16'h557f;

	lut_sub lut_3509 ({sk[769], n_n2162, x21493x, n_n2159, n_n2158, x21492x, x21498x}, x21508x);
	defparam lut_3509.LUT_SIZE = 7;
	defparam lut_3509.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_3516 ({sk[770], n_n148, n_n4, n_n3, n_n7, n_n60, n_n7443}, x24210x);
	defparam lut_3516.LUT_SIZE = 7;
	defparam lut_3516.mask = 128'h5555ffff5555ffffaa80a080aa000000;

	lut_sub lut_3520 ({sk[771], n_n208, n_n106, x916x, n_n3, n_n60, x24210x}, x21525x);
	defparam lut_3520.LUT_SIZE = 7;
	defparam lut_3520.mask = 128'h5555ffff5555ffffaaaaafafaabbafff;

	lut_sub lut_3525 ({sk[772], i_14_, i_13_, i_12_, i_15_, n_n247, n_n267}, x1512x);
	defparam lut_3525.LUT_SIZE = 7;
	defparam lut_3525.mask = 128'h5555ffff5555ffff0750507077000000;

	lut_sub lut_3536 ({sk[773], n_n6, n_n5, x389x, x253x, x1285x, x1511x}, x21587x);
	defparam lut_3536.LUT_SIZE = 7;
	defparam lut_3536.mask = 128'h5555ffff5555ffff00ff77ff0fff7fff;

	lut_sub lut_3541 ({sk[774], i_7_, i_8_, i_6_, x909x, x1512x, x21587x}, x21588x);
	defparam lut_3541.LUT_SIZE = 7;
	defparam lut_3541.mask = 128'h5555ffff5555ffff5555555555555755;

	lut_sub lut_3544 ({sk[775], n_n106, n_n145, n_n48, n_n53, n_n60, x21564x}, n_n2148);
	defparam lut_3544.LUT_SIZE = 7;
	defparam lut_3544.mask = 128'h5555ffff5555ffff57575f5f5fff5fff;

	lut_sub lut_3550 ({sk[776], x909x, n_n279, n_n261, x902x, x296x, x21575x}, n_n2140);
	defparam lut_3550.LUT_SIZE = 7;
	defparam lut_3550.mask = 128'h5555ffff5555ffff555555555577557f;

	lut_sub lut_3554 ({sk[777], n_n151, n_n273, n_n283, x922x, x376x, x21571x}, x21572x);
	defparam lut_3554.LUT_SIZE = 7;
	defparam lut_3554.mask = 128'h5555ffff5555ffff77777777777f7f7f;

	lut_sub lut_3559 ({sk[778], n_n6, x78x, n_n279, x901x, x267x, x873x}, x21580x);
	defparam lut_3559.LUT_SIZE = 7;
	defparam lut_3559.mask = 128'h5555ffff5555ffff55555555777fffff;

	lut_sub lut_3564 ({sk[779], n_n5, x373x, x462x, x492x, x21568x, x1510x}, x24106x);
	defparam lut_3564.LUT_SIZE = 7;
	defparam lut_3564.mask = 128'h5555ffff5555ffffc000000080000000;

	lut_sub lut_3567 ({sk[780], n_n2148, n_n2140, x21572x, x21580x, x24106x}, x21589x);
	defparam lut_3567.LUT_SIZE = 6;
	defparam lut_3567.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_3573 ({sk[781], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x922x);
	defparam lut_3573.LUT_SIZE = 7;
	defparam lut_3573.mask = 128'h5555ffff5555ffff0000000080000000;

	lut_sub lut_3575 ({sk[782], i_14_, i_13_, i_12_, i_15_, x901x, n_n247}, x1469x);
	defparam lut_3575.LUT_SIZE = 7;
	defparam lut_3575.mask = 128'h5555ffff5555ffff0550505077000000;

	lut_sub lut_3583 ({sk[783], n_n283, x922x, x456x, x1092x, x21603x, x286x}, x21606x);
	defparam lut_3583.LUT_SIZE = 7;
	defparam lut_3583.mask = 128'h5555ffff5555ffff77ff77ff77ff7fff;

	lut_sub lut_3588 ({sk[784], x905x, n_n279, n_n48, n_n53, x899x, x1508x}, x21607x);
	defparam lut_3588.LUT_SIZE = 7;
	defparam lut_3588.mask = 128'h5555ffff5555ffff0555057705550f7f;

	lut_sub lut_3593 ({sk[785], n_n283, x922x, x464x, x376x, x21595x, x1470x}, x24105x);
	defparam lut_3593.LUT_SIZE = 7;
	defparam lut_3593.mask = 128'h5555ffff5555ffffc000c000c0008000;

	lut_sub lut_3597 ({sk[786], n_n273, x922x, x1469x, x21606x, x21607x, x24105x}, x21613x);
	defparam lut_3597.LUT_SIZE = 7;
	defparam lut_3597.mask = 128'h5555ffff5555ffffbfbfbfbfbfbfbfff;

	lut_sub lut_3602 ({sk[787], i_7_, i_6_, i_1_, i_2_, i_0_, n_n284}, n_n5660);
	defparam lut_3602.LUT_SIZE = 7;
	defparam lut_3602.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_3604 ({sk[788], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, x880x);
	defparam lut_3604.LUT_SIZE = 7;
	defparam lut_3604.mask = 128'h5555ffff5555ffff0000000040400000;

	lut_sub lut_3607 ({sk[789], i_7_, i_8_, i_6_, x916x, n_n222, x902x}, n_n7297);
	defparam lut_3607.LUT_SIZE = 7;
	defparam lut_3607.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_3609 ({sk[790], i_14_, i_13_, i_12_, x908x, x902x}, x249x);
	defparam lut_3609.LUT_SIZE = 6;
	defparam lut_3609.mask = 64'h3f3f3f3f05050030;

	lut_sub lut_3613 ({sk[791], i_14_, i_13_, i_12_, x914x, x912x}, x263x);
	defparam lut_3613.LUT_SIZE = 6;
	defparam lut_3613.mask = 64'h3f3f3f3f50300000;

	lut_sub lut_3616 ({sk[792], i_14_, i_13_, i_12_, i_15_, x912x, n_n137}, x313x);
	defparam lut_3616.LUT_SIZE = 7;
	defparam lut_3616.mask = 128'h5555ffff5555ffff5073507350505050;

	lut_sub lut_3620 ({sk[793], n_n4, n_n3, n_n7297, x249x, x263x, x313x}, n_n1730);
	defparam lut_3620.LUT_SIZE = 7;
	defparam lut_3620.mask = 128'h5555ffff5555ffff00ff77ff0fff7fff;

	lut_sub lut_3625 ({sk[794], i_14_, i_13_, i_12_, x897x}, n_n25);
	defparam lut_3625.LUT_SIZE = 5;
	defparam lut_3625.mask = 32'h0f0f0004;

	lut_sub lut_3627 ({sk[795], n_n281, n_n208, x916x, n_n220, x908x, x902x}, x641x);
	defparam lut_3627.LUT_SIZE = 7;
	defparam lut_3627.mask = 128'h5555ffff5555ffff0000000300000057;

	lut_sub lut_3630 ({sk[796], i_14_, i_13_, i_12_, i_15_, n_n275, x228x}, x1732x);
	defparam lut_3630.LUT_SIZE = 7;
	defparam lut_3630.mask = 128'h5555ffff5555ffff5557555755557755;

	lut_sub lut_3636 ({sk[797], n_n208, x916x, n_n3, n_n25, x641x, x1732x}, n_n1729);
	defparam lut_3636.LUT_SIZE = 7;
	defparam lut_3636.mask = 128'h5555ffff5555ffff3377337733773f7f;

	lut_sub lut_3640 ({sk[798], n_n266, x909x, x379x, x21736x, x21737x, x24103x}, x21739x);
	defparam lut_3640.LUT_SIZE = 7;
	defparam lut_3640.mask = 128'h5555ffff5555ffffbfbfbfbfbfbfbfff;

	lut_sub lut_3645 ({sk[799], n_n1787, n_n1788, n_n1791, x21719x, x21718x, x21727x}, x21740x);
	defparam lut_3645.LUT_SIZE = 7;
	defparam lut_3645.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_3652 ({sk[800], n_n57, n_n56, x180x, x99x, n_n6046, x24166x}, x21768x);
	defparam lut_3652.LUT_SIZE = 7;
	defparam lut_3652.mask = 128'h5555ffff5555ffffbbbbbbffbfffbfff;

	lut_sub lut_3658 ({sk[801], n_n100, x1597x, x21752x, x21759x, x21760x, x3066x}, x21769x);
	defparam lut_3658.LUT_SIZE = 7;
	defparam lut_3658.mask = 128'h5555ffff5555ffff7fff7fff7fffffff;

	lut_sub lut_3664 ({sk[802], x21779x, x21792x, x21800x, n_n1773, x24099x}, n_n1688);
	defparam lut_3664.LUT_SIZE = 6;
	defparam lut_3664.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_3670 ({sk[803], x21808x, x21809x, x21817x, x21825x, n_n1761, x21816x}, n_n1687);
	defparam lut_3670.LUT_SIZE = 7;
	defparam lut_3670.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_3677 ({sk[804], i_7_, i_8_, i_6_, x916x, n_n222, x899x}, n_n7345);
	defparam lut_3677.LUT_SIZE = 7;
	defparam lut_3677.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_3679 ({sk[805], i_14_, i_13_, i_12_, x903x, x897x, x279x}, x1749x);
	defparam lut_3679.LUT_SIZE = 7;
	defparam lut_3679.mask = 128'h5555ffff5555ffff77555f5555555555;

	lut_sub lut_3683 ({sk[806], i_14_, i_13_, i_12_, x908x, x902x}, x1748x);
	defparam lut_3683.LUT_SIZE = 6;
	defparam lut_3683.mask = 64'h3f3f3f3f05050070;

	lut_sub lut_3688 ({sk[807], n_n281, n_n208, x916x, n_n220, x905x, x899x}, x622x);
	defparam lut_3688.LUT_SIZE = 7;
	defparam lut_3688.mask = 128'h5555ffff5555ffff0000000300000057;

	lut_sub lut_3691 ({sk[808], n_n4, n_n3, n_n7345, x1749x, x1748x, x622x}, x21885x);
	defparam lut_3691.LUT_SIZE = 7;
	defparam lut_3691.mask = 128'h5555ffff5555ffff55ff77ff5fff7fff;

	lut_sub lut_3696 ({sk[809], i_14_, i_13_, i_12_, i_15_, n_n242, x230x}, x1821x);
	defparam lut_3696.LUT_SIZE = 7;
	defparam lut_3696.mask = 128'h5555ffff5555ffff5757755755557755;

	lut_sub lut_3704 ({sk[810], i_14_, i_13_, i_12_, i_15_, n_n242, n_n259}, x1820x);
	defparam lut_3704.LUT_SIZE = 7;
	defparam lut_3704.mask = 128'h5555ffff5555ffff0007000700007300;

	lut_sub lut_3712 ({sk[811], i_7_, i_8_, i_6_, x916x, x1821x, x1820x}, x21886x);
	defparam lut_3712.LUT_SIZE = 7;
	defparam lut_3712.mask = 128'h5555ffff5555ffff0003000500000000;

	lut_sub lut_3715 ({sk[812], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x248x);
	defparam lut_3715.LUT_SIZE = 7;
	defparam lut_3715.mask = 128'h5555ffff5555ffff0010001000004000;

	lut_sub lut_3719 ({sk[813], i_14_, i_13_, i_12_, x907x, x901x}, x154x);
	defparam lut_3719.LUT_SIZE = 6;
	defparam lut_3719.mask = 64'h3f3f3f3f50300000;

	lut_sub lut_3722 ({sk[814], i_9_, i_10_, i_11_}, n_n282);
	defparam lut_3722.LUT_SIZE = 4;
	defparam lut_3722.mask = 16'h5580;

	lut_sub lut_3724 ({sk[815], i_14_, i_13_, i_12_, i_15_, x154x, n_n282}, x957x);
	defparam lut_3724.LUT_SIZE = 7;
	defparam lut_3724.mask = 128'h5555ffff5555ffff3337333733337733;

	lut_sub lut_3730 ({sk[816], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, n_n137);
	defparam lut_3730.LUT_SIZE = 7;
	defparam lut_3730.mask = 128'h5555ffff5555ffff0000000000080000;

	lut_sub lut_3732 ({sk[817], i_15_, n_n137}, n_n88);
	defparam lut_3732.LUT_SIZE = 3;
	defparam lut_3732.mask = 8'h51;

	lut_sub lut_3734 ({sk[818], n_n208, x916x, x374x, n_n7306, x141x, n_n1346}, x21935x);
	defparam lut_3734.LUT_SIZE = 7;
	defparam lut_3734.mask = 128'h5555ffff5555ffff5fff5fff5fff7fff;

	lut_sub lut_3739 ({sk[819], n_n208, x916x, n_n41, x93x, x476x, n_n1356}, x21941x);
	defparam lut_3739.LUT_SIZE = 7;
	defparam lut_3739.mask = 128'h5555ffff5555ffff7777777777777fff;

	lut_sub lut_3744 ({sk[820], n_n208, x916x, n_n258, x897x, x3678x, x1390x}, x21946x);
	defparam lut_3744.LUT_SIZE = 7;
	defparam lut_3744.mask = 128'h5555ffff5555ffff333333333333777f;

	lut_sub lut_3748 ({sk[821], n_n4, n_n3, n_n76, x92x, x56x, x1391x}, x21947x);
	defparam lut_3748.LUT_SIZE = 7;
	defparam lut_3748.mask = 128'h5555ffff5555ffff000077770fff7fff;

	lut_sub lut_3753 ({sk[822], n_n4, n_n3, x1491x, x1490x, x1493x, x1492x}, x24085x);
	defparam lut_3753.LUT_SIZE = 7;
	defparam lut_3753.mask = 128'h5555ffff5555ffffffffc0c0aa008000;

	lut_sub lut_3758 ({sk[823], x21935x, x21941x, x21946x, x21947x, x24085x}, x21950x);
	defparam lut_3758.LUT_SIZE = 6;
	defparam lut_3758.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_3764 ({sk[824], i_14_, i_13_, i_12_, i_15_, n_n282, n_n270}, x991x);
	defparam lut_3764.LUT_SIZE = 7;
	defparam lut_3764.mask = 128'h5555ffff5555ffff0333300770057570;

	lut_sub lut_3779 ({sk[825], n_n1, n_n2, x93x, n_n32, x990x, x85x}, x21956x);
	defparam lut_3779.LUT_SIZE = 7;
	defparam lut_3779.mask = 128'h5555ffff5555ffff00003fff55557fff;

	lut_sub lut_3784 ({sk[826], x915x, n_n273, n_n283, x93x, x1053x, x1052x}, n_n1118);
	defparam lut_3784.LUT_SIZE = 7;
	defparam lut_3784.mask = 128'h5555ffff5555ffff0000000000335f7f;

	lut_sub lut_3788 ({sk[827], i_14_, i_13_, i_12_, i_15_, n_n275, x431x}, x1425x);
	defparam lut_3788.LUT_SIZE = 7;
	defparam lut_3788.mask = 128'h5555ffff5555ffff5775755555577775;

	lut_sub lut_3797 ({sk[828], n_n1, n_n2, n_n76, x92x, x56x, x1424x}, x21968x);
	defparam lut_3797.LUT_SIZE = 7;
	defparam lut_3797.mask = 128'h5555ffff5555ffff000077770fff7fff;

	lut_sub lut_3802 ({sk[829], n_n1, x991x, x21956x, n_n1118, x1425x, x21968x}, n_n1091);
	defparam lut_3802.LUT_SIZE = 7;
	defparam lut_3802.mask = 128'h5555ffff5555ffff5fff5fff7fffffff;

	lut_sub lut_3808 ({sk[830], n_n265, n_n268, x124x, x212x, x1454x, x1453x}, n_n1112);
	defparam lut_3808.LUT_SIZE = 7;
	defparam lut_3808.mask = 128'h5555ffff5555ffff00003fff55557fff;

	lut_sub lut_3813 ({sk[831], x907x, n_n266, x916x, n_n3246, n_n220, x24211x}, x22007x);
	defparam lut_3813.LUT_SIZE = 7;
	defparam lut_3813.mask = 128'h5555ffff5555ffffafafafafafafafbf;

	lut_sub lut_3817 ({sk[832], n_n208, n_n266, x916x, n_n62, x68x, x1471x}, n_n1176);
	defparam lut_3817.LUT_SIZE = 7;
	defparam lut_3817.mask = 128'h5555ffff5555ffff0000000f0077007f;

	lut_sub lut_3821 ({sk[833], n_n4, x518x, x94x, x77x, x3635x, x455x}, x22012x);
	defparam lut_3821.LUT_SIZE = 7;
	defparam lut_3821.mask = 128'h5555ffff5555ffff7777ffff7fffffff;

	lut_sub lut_3827 ({sk[834], n_n268, n_n3, n_n1173, x1428x, x22003x, x22004x}, x24084x);
	defparam lut_3827.LUT_SIZE = 7;
	defparam lut_3827.mask = 128'h5555ffff5555ffffff00f00088008000;

	lut_sub lut_3832 ({sk[835], n_n1112, x22007x, n_n1176, x22012x, x24084x}, n_n1089);
	defparam lut_3832.LUT_SIZE = 6;
	defparam lut_3832.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_3838 ({sk[836], n_n1204, x22041x, n_n1208, x22054x, x22040x, x22053x}, x22063x);
	defparam lut_3838.LUT_SIZE = 7;
	defparam lut_3838.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_3845 ({sk[837], n_n1215, n_n1212, x22076x, x22088x, x22075x, x22087x}, x22096x);
	defparam lut_3845.LUT_SIZE = 7;
	defparam lut_3845.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_3852 ({sk[838], n_n6, n_n5, n_n1217, x1209x, x1208x, x22097x}, x22099x);
	defparam lut_3852.LUT_SIZE = 7;
	defparam lut_3852.mask = 128'h5555ffff5555ffff55ff77ff5fff7fff;

	lut_sub lut_3857 ({sk[839], x22020x, x22021x, x2777x, x22031x}, x22100x);
	defparam lut_3857.LUT_SIZE = 5;
	defparam lut_3857.mask = 32'h0f0f7fff;

	lut_sub lut_3862 ({sk[840], n_n1, n_n1173, n_n1210, x1388x, x22061x, x22093x}, x24094x);
	defparam lut_3862.LUT_SIZE = 7;
	defparam lut_3862.mask = 128'h5555ffff5555ffff8800000080000000;

	lut_sub lut_3865 ({sk[841], i_14_, i_13_, i_12_, x913x}, n_n240);
	defparam lut_3865.LUT_SIZE = 5;
	defparam lut_3865.mask = 32'h0f0f0010;

	lut_sub lut_3867 ({sk[842], n_n4, n_n3, n_n70, x1211x, x1210x, x743x}, x22338x);
	defparam lut_3867.LUT_SIZE = 7;
	defparam lut_3867.mask = 128'h5555ffff5555ffff555577775fff7fff;

	lut_sub lut_3872 ({sk[843], n_n208, x916x, n_n3, x1214x, x22336x, x1212x}, x22339x);
	defparam lut_3872.LUT_SIZE = 7;
	defparam lut_3872.mask = 128'h5555ffff5555ffff003f003f003f557f;

	lut_sub lut_3876 ({sk[844], n_n3, n_n7224, x518x, x904x, n_n256, x833x}, x22348x);
	defparam lut_3876.LUT_SIZE = 7;
	defparam lut_3876.mask = 128'h5555ffff5555ffff55ffffff57ffffff;

	lut_sub lut_3881 ({sk[845], n_n4, n_n3, n_n7306, x1218x, x320x, x1257x}, x22357x);
	defparam lut_3881.LUT_SIZE = 7;
	defparam lut_3881.mask = 128'h5555ffff5555ffff00ff55ff3fff7fff;

	lut_sub lut_3886 ({sk[846], n_n4, n_n3, x1216x, x1215x, x642x, x1217x}, x24076x);
	defparam lut_3886.LUT_SIZE = 7;
	defparam lut_3886.mask = 128'h5555ffff5555ffffcccc8080cc008000;

	lut_sub lut_3891 ({sk[847], x22338x, x22339x, x22348x, x22357x, x24076x}, n_n338);
	defparam lut_3891.LUT_SIZE = 6;
	defparam lut_3891.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_3897 ({sk[848], i_14_, i_13_, i_12_, x905x}, n_n257);
	defparam lut_3897.LUT_SIZE = 5;
	defparam lut_3897.mask = 32'h0f0f0010;

	lut_sub lut_3899 ({sk[849], i_14_, i_13_, i_12_, x913x}, n_n67);
	defparam lut_3899.LUT_SIZE = 5;
	defparam lut_3899.mask = 32'h0f0f1000;

	lut_sub lut_3901 ({sk[850], i_14_, i_13_, i_12_, x904x}, n_n252);
	defparam lut_3901.LUT_SIZE = 5;
	defparam lut_3901.mask = 32'h0f0f0010;

	lut_sub lut_3903 ({sk[851], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x308x);
	defparam lut_3903.LUT_SIZE = 7;
	defparam lut_3903.mask = 128'h5555ffff5555ffff0010000040004000;

	lut_sub lut_3907 ({sk[852], i_14_, i_13_, i_12_, i_15_, x906x, n_n259}, x22364x);
	defparam lut_3907.LUT_SIZE = 7;
	defparam lut_3907.mask = 128'h5555ffff5555ffff0050000000370050;

	lut_sub lut_3912 ({sk[853], n_n4, n_n3, n_n67, n_n252, x308x, x22364x}, n_n381);
	defparam lut_3912.LUT_SIZE = 7;
	defparam lut_3912.mask = 128'h5555ffff5555ffff000077770fff7fff;

	lut_sub lut_3917 ({sk[854], x22432x, x22433x, x22440x, n_n418, x24173x}, n_n342);
	defparam lut_3917.LUT_SIZE = 6;
	defparam lut_3917.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_3923 ({sk[855], n_n273, x922x, n_n439, x1128x, x22463x}, x22465x);
	defparam lut_3923.LUT_SIZE = 6;
	defparam lut_3923.mask = 64'h3f3f3f3f5f5f5f7f;

	lut_sub lut_3927 ({sk[856], x22447x, n_n442, n_n438, n_n443, x22446x, x22457x}, x22466x);
	defparam lut_3927.LUT_SIZE = 7;
	defparam lut_3927.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_3934 ({sk[857], x2309x, x22470x, n_n372, x22481x}, n_n345);
	defparam lut_3934.LUT_SIZE = 5;
	defparam lut_3934.mask = 32'h0f0f7fff;

	lut_sub lut_3939 ({sk[858], x915x, n_n261, n_n464, x1261x, x22502x}, x22504x);
	defparam lut_3939.LUT_SIZE = 6;
	defparam lut_3939.mask = 64'h3f3f3f3f5f5f5f7f;

	lut_sub lut_3943 ({sk[859], x22487x, x22493x, n_n467, x22492x, x24081x}, x22505x);
	defparam lut_3943.LUT_SIZE = 6;
	defparam lut_3943.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_3949 ({sk[860], i_9_, i_10_, i_11_, i_15_, n_n225}, x126x);
	defparam lut_3949.LUT_SIZE = 6;
	defparam lut_3949.mask = 64'h3f3f3f3f50000000;

	lut_sub lut_3952 ({sk[861], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x177x);
	defparam lut_3952.LUT_SIZE = 7;
	defparam lut_3952.mask = 128'h5555ffff5555ffff0000000010001040;

	lut_sub lut_3956 ({sk[862], n_n208, x916x, n_n104, n_n3, x126x, x177x}, n_n783);
	defparam lut_3956.LUT_SIZE = 7;
	defparam lut_3956.mask = 128'h5555ffff5555ffff07070707070757ff;

	lut_sub lut_3961 ({sk[863], i_14_, i_13_, i_12_, i_15_, n_n270}, x88x);
	defparam lut_3961.LUT_SIZE = 6;
	defparam lut_3961.mask = 64'h3f3f3f3f00001004;

	lut_sub lut_3964 ({sk[864], i_9_, i_10_, i_11_, i_15_, n_n225}, x114x);
	defparam lut_3964.LUT_SIZE = 6;
	defparam lut_3964.mask = 64'h3f3f3f3f00000500;

	lut_sub lut_3967 ({sk[865], i_14_, i_13_, i_12_, i_15_, n_n275, x897x}, x1300x);
	defparam lut_3967.LUT_SIZE = 7;
	defparam lut_3967.mask = 128'h5555ffff5555ffff0000000003550330;

	lut_sub lut_3972 ({sk[866], n_n4, n_n3, x88x, x114x, n_n7297, x1300x}, n_n781);
	defparam lut_3972.LUT_SIZE = 7;
	defparam lut_3972.mask = 128'h5555ffff5555ffff333377773fff7fff;

	lut_sub lut_3977 ({sk[867], i_14_, i_13_, i_12_, x911x}, n_n216);
	defparam lut_3977.LUT_SIZE = 5;
	defparam lut_3977.mask = 32'h0f0f0010;

	lut_sub lut_3979 ({sk[868], i_9_, i_10_, i_11_, i_15_, n_n225}, x128x);
	defparam lut_3979.LUT_SIZE = 6;
	defparam lut_3979.mask = 64'h3f3f3f3f00000050;

	lut_sub lut_3982 ({sk[869], i_7_, i_8_, i_6_, x916x, n_n258, x899x}, n_n7344);
	defparam lut_3982.LUT_SIZE = 7;
	defparam lut_3982.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_3984 ({sk[870], i_14_, i_13_, i_12_, n_n4, x905x, x899x}, n_n876);
	defparam lut_3984.LUT_SIZE = 7;
	defparam lut_3984.mask = 128'h5555ffff5555ffff0000000005000503;

	lut_sub lut_3988 ({sk[871], n_n4, n_n3, n_n216, x128x, n_n7344, n_n876}, x22602x);
	defparam lut_3988.LUT_SIZE = 7;
	defparam lut_3988.mask = 128'h5555ffff5555ffff777777ff7fff7fff;

	lut_sub lut_3994 ({sk[872], i_9_, i_10_, i_11_, i_15_, n_n225}, x120x);
	defparam lut_3994.LUT_SIZE = 6;
	defparam lut_3994.mask = 64'h3f3f3f3f05000000;

	lut_sub lut_3997 ({sk[873], i_14_, i_13_, i_12_, x91x, x903x, x897x}, x1256x);
	defparam lut_3997.LUT_SIZE = 7;
	defparam lut_3997.mask = 128'h5555ffff5555ffff0f0f0f7f0f5f0f0f;

	lut_sub lut_4002 ({sk[874], i_14_, i_13_, i_12_, i_15_, n_n242, n_n270}, x1635x);
	defparam lut_4002.LUT_SIZE = 7;
	defparam lut_4002.mask = 128'h5555ffff5555ffff0000007707000770;

	lut_sub lut_4013 ({sk[875], n_n4, n_n31, n_n3, x120x, x1256x, x1635x}, x22603x);
	defparam lut_4013.LUT_SIZE = 7;
	defparam lut_4013.mask = 128'h5555ffff5555ffff005f00ff337f33ff;

	lut_sub lut_4018 ({sk[876], x22611x, x22612x, x22620x, x22621x, x22625x, x22626x}, n_n743);
	defparam lut_4018.LUT_SIZE = 7;
	defparam lut_4018.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_4025 ({sk[877], x22640x, n_n838, x22644x, x22645x, x24213x}, n_n742);
	defparam lut_4025.LUT_SIZE = 6;
	defparam lut_4025.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_4031 ({sk[878], n_n863, n_n100, n_n94, x1934x, x1396x, x22667x}, x22670x);
	defparam lut_4031.LUT_SIZE = 7;
	defparam lut_4031.mask = 128'h5555ffff5555ffff555f777fffffffff;

	lut_sub lut_4036 ({sk[879], n_n855, x22655x, x22662x, x22663x, x22654x}, x22671x);
	defparam lut_4036.LUT_SIZE = 6;
	defparam lut_4036.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_4042 ({sk[880], x22678x, x22679x, x22685x, x22686x, x22691x, x22692x}, n_n739);
	defparam lut_4042.LUT_SIZE = 7;
	defparam lut_4042.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_4049 ({sk[881], i_7_, i_8_, i_6_, x916x, x900x, n_n228}, n_n7400);
	defparam lut_4049.LUT_SIZE = 7;
	defparam lut_4049.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_4051 ({sk[882], i_14_, i_13_, i_12_, x898x}, n_n15);
	defparam lut_4051.LUT_SIZE = 5;
	defparam lut_4051.mask = 32'h0f0f0001;

	lut_sub lut_4053 ({sk[883], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x109x);
	defparam lut_4053.LUT_SIZE = 7;
	defparam lut_4053.mask = 128'h5555ffff5555ffff0000000010001040;

	lut_sub lut_4057 ({sk[884], i_14_, i_13_, i_12_, i_15_, x900x, n_n259}, x22834x);
	defparam lut_4057.LUT_SIZE = 7;
	defparam lut_4057.mask = 128'h5555ffff5555ffff0000005500050033;

	lut_sub lut_4062 ({sk[885], i_7_, i_8_, i_6_, x916x, x901x, n_n228}, x505x);
	defparam lut_4062.LUT_SIZE = 7;
	defparam lut_4062.mask = 128'h5555ffff5555ffff0001000100000000;

	lut_sub lut_4065 ({sk[886], n_n3, n_n7400, n_n15, x109x, x22834x, x505x}, x22839x);
	defparam lut_4065.LUT_SIZE = 7;
	defparam lut_4065.mask = 128'h5555ffff5555ffff5555ffff7fffffff;

	lut_sub lut_4071 ({sk[887], i_14_, i_13_, i_12_}, n_n225);
	defparam lut_4071.LUT_SIZE = 4;
	defparam lut_4071.mask = 16'h5510;

	lut_sub lut_4073 ({sk[888], i_9_, i_10_, i_11_}, n_n247);
	defparam lut_4073.LUT_SIZE = 4;
	defparam lut_4073.mask = 16'h5508;

	lut_sub lut_4075 ({sk[889], i_14_, i_13_, i_12_, x914x, x912x}, x368x);
	defparam lut_4075.LUT_SIZE = 6;
	defparam lut_4075.mask = 64'h3f3f3f3f00005003;

	lut_sub lut_4078 ({sk[890], i_14_, i_13_, i_12_, i_15_, n_n247, x368x}, x115x);
	defparam lut_4078.LUT_SIZE = 7;
	defparam lut_4078.mask = 128'h5555ffff5555ffff5555555555555755;

	lut_sub lut_4081 ({sk[891], i_14_, i_13_, i_12_, x914x, x115x, x912x}, x960x);
	defparam lut_4081.LUT_SIZE = 7;
	defparam lut_4081.mask = 128'h5555ffff5555ffff3333337f33773333;

	lut_sub lut_4086 ({sk[892], i_7_, i_8_, i_6_, x909x}, n_n189);
	defparam lut_4086.LUT_SIZE = 5;
	defparam lut_4086.mask = 32'h0f0f4000;

	lut_sub lut_4088 ({sk[893], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x24216x);
	defparam lut_4088.LUT_SIZE = 7;
	defparam lut_4088.mask = 128'h5555ffff5555ffff00000000dd1d1515;

	lut_sub lut_4094 ({sk[894], i_9_, i_10_, i_11_, i_15_, n_n279, x24216x}, x961x);
	defparam lut_4094.LUT_SIZE = 7;
	defparam lut_4094.mask = 128'h5555ffff5555ffff5555555557575555;

	lut_sub lut_4098 ({sk[895], i_9_, i_10_, i_14_, i_13_, i_12_}, x24147x);
	defparam lut_4098.LUT_SIZE = 6;
	defparam lut_4098.mask = 64'h3f3f3f3fff04ffff;

	lut_sub lut_4102 ({sk[896], i_9_, i_10_, i_11_, i_15_, n_n258, x24147x}, x964x);
	defparam lut_4102.LUT_SIZE = 7;
	defparam lut_4102.mask = 128'h5555ffff5555ffffaabababaaaaaaaaa;

	lut_sub lut_4107 ({sk[897], i_9_, i_10_, i_14_, i_13_, i_12_}, x24146x);
	defparam lut_4107.LUT_SIZE = 6;
	defparam lut_4107.mask = 64'h3f3f3f3fffff04ff;

	lut_sub lut_4111 ({sk[898], i_9_, i_10_, i_11_, i_15_, n_n258, x24146x}, x967x);
	defparam lut_4111.LUT_SIZE = 7;
	defparam lut_4111.mask = 128'h5555ffff5555ffffffffffffbabaaaaa;

	lut_sub lut_4116 ({sk[899], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19198x);
	defparam lut_4116.LUT_SIZE = 7;
	defparam lut_4116.mask = 128'h5555ffff5555ffffffcf000000000000;

	lut_sub lut_4123 ({sk[900], i_9_, i_10_, i_11_, i_15_, n_n258, x19198x}, x970x);
	defparam lut_4123.LUT_SIZE = 7;
	defparam lut_4123.mask = 128'h5555ffff5555ffff75555555ffffffff;

	lut_sub lut_4127 ({sk[901], i_7_, i_6_, x915x}, x5923x);
	defparam lut_4127.LUT_SIZE = 4;
	defparam lut_4127.mask = 16'h5510;

	lut_sub lut_4129 ({sk[902], n_n255, n_n241, x964x, x967x, x970x, x5923x}, n_n5020);
	defparam lut_4129.LUT_SIZE = 7;
	defparam lut_4129.mask = 128'h5555ffff5555ffff555577ff5f5f7fff;

	lut_sub lut_4134 ({sk[903], i_14_, i_13_, i_12_}, n_n222);
	defparam lut_4134.LUT_SIZE = 4;
	defparam lut_4134.mask = 16'h5502;

	lut_sub lut_4136 ({sk[904], i_9_, i_10_, i_11_, i_15_}, x898x);
	defparam lut_4136.LUT_SIZE = 5;
	defparam lut_4136.mask = 32'h0f0f0001;

	lut_sub lut_4138 ({sk[905], i_7_, i_8_, i_6_, x909x, n_n222, x898x}, n_n6036);
	defparam lut_4138.LUT_SIZE = 7;
	defparam lut_4138.mask = 128'h5555ffff5555ffff0000000000000001;

	lut_sub lut_4140 ({sk[906], i_7_, i_8_, i_6_, x909x, n_n258, x898x}, n_n6035);
	defparam lut_4140.LUT_SIZE = 7;
	defparam lut_4140.mask = 128'h5555ffff5555ffff0000000000000001;

	lut_sub lut_4142 ({sk[907], i_14_, i_13_, i_12_, x898x}, n_n186);
	defparam lut_4142.LUT_SIZE = 5;
	defparam lut_4142.mask = 32'h0f0f0040;

	lut_sub lut_4144 ({sk[908], i_14_, i_13_, i_12_, n_n266, x909x, x898x}, n_n4970);
	defparam lut_4144.LUT_SIZE = 7;
	defparam lut_4144.mask = 128'h5555ffff5555ffff0000000001010100;

	lut_sub lut_4148 ({sk[909], i_14_, i_13_, i_12_, x906x}, x51x);
	defparam lut_4148.LUT_SIZE = 5;
	defparam lut_4148.mask = 32'h0f0f1400;

	lut_sub lut_4151 ({sk[910], i_14_, i_13_, i_12_, n_n266, x909x, x906x}, n_n4959);
	defparam lut_4151.LUT_SIZE = 7;
	defparam lut_4151.mask = 128'h5555ffff5555ffff0001010100000000;

	lut_sub lut_4155 ({sk[911], i_14_, i_13_, i_12_, x901x}, n_n280);
	defparam lut_4155.LUT_SIZE = 5;
	defparam lut_4155.mask = 32'h0f0f4000;

	lut_sub lut_4157 ({sk[912], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x64x);
	defparam lut_4157.LUT_SIZE = 7;
	defparam lut_4157.mask = 128'h5555ffff5555ffff0010001000000000;

	lut_sub lut_4160 ({sk[913], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x200x);
	defparam lut_4160.LUT_SIZE = 7;
	defparam lut_4160.mask = 128'h5555ffff5555ffff3305000500000000;

	lut_sub lut_4164 ({sk[914], i_14_, i_13_, i_12_, n_n56, x64x, x901x}, n_n4948);
	defparam lut_4164.LUT_SIZE = 7;
	defparam lut_4164.mask = 128'h5555ffff5555ffff0703030303030303;

	lut_sub lut_4167 ({sk[915], i_14_, i_13_, i_12_, i_15_, n_n270}, x170x);
	defparam lut_4167.LUT_SIZE = 6;
	defparam lut_4167.mask = 64'h3f3f3f3f00001044;

	lut_sub lut_4171 ({sk[916], i_14_, i_13_, i_12_, x900x}, n_n65);
	defparam lut_4171.LUT_SIZE = 5;
	defparam lut_4171.mask = 32'h0f0f0001;

	lut_sub lut_4173 ({sk[917], i_9_, i_10_, i_11_}, n_n267);
	defparam lut_4173.LUT_SIZE = 4;
	defparam lut_4173.mask = 16'h5510;

	lut_sub lut_4175 ({sk[918], i_14_, i_13_, i_12_, i_15_, n_n267}, x186x);
	defparam lut_4175.LUT_SIZE = 6;
	defparam lut_4175.mask = 64'h3f3f3f3f40100400;

	lut_sub lut_4179 ({sk[919], i_9_, i_10_, i_11_, i_15_}, x904x);
	defparam lut_4179.LUT_SIZE = 5;
	defparam lut_4179.mask = 32'h0f0f0002;

	lut_sub lut_4181 ({sk[920], i_14_, i_13_, i_12_, x898x, x904x}, x173x);
	defparam lut_4181.LUT_SIZE = 6;
	defparam lut_4181.mask = 64'h3f3f3f3f00300503;

	lut_sub lut_4185 ({sk[921], i_14_, i_13_, i_12_, i_15_, x173x, n_n267}, x972x);
	defparam lut_4185.LUT_SIZE = 7;
	defparam lut_4185.mask = 128'h5555ffff5555ffff7333373333333333;

	lut_sub lut_4189 ({sk[922], i_14_, i_13_, i_12_, x907x, x905x, x113x}, x19685x);
	defparam lut_4189.LUT_SIZE = 7;
	defparam lut_4189.mask = 128'h5555ffff5555ffff55777777555f5555;

	lut_sub lut_4195 ({sk[923], i_9_, i_10_, i_11_}, n_n253);
	defparam lut_4195.LUT_SIZE = 4;
	defparam lut_4195.mask = 16'h5501;

	lut_sub lut_4197 ({sk[924], i_14_, i_13_, i_12_, i_15_, n_n247, n_n253}, x974x);
	defparam lut_4197.LUT_SIZE = 7;
	defparam lut_4197.mask = 128'h5555ffff5555ffff7000070000700007;

	lut_sub lut_4206 ({sk[925], i_14_, i_13_, i_12_, x901x}, n_n63);
	defparam lut_4206.LUT_SIZE = 5;
	defparam lut_4206.mask = 32'h0f0f0001;

	lut_sub lut_4208 ({sk[926], i_14_, i_13_, i_12_, x900x, x906x}, x246x);
	defparam lut_4208.LUT_SIZE = 6;
	defparam lut_4208.mask = 64'h3f3f3f3f00000503;

	lut_sub lut_4211 ({sk[927], n_n281, n_n56, x19685x, x904x, n_n63, x246x}, x5341x);
	defparam lut_4211.LUT_SIZE = 7;
	defparam lut_4211.mask = 128'h5555ffff5555ffff000077ff00007fff;

	lut_sub lut_4216 ({sk[928], n_n57, n_n56, n_n65, x186x, x972x, x974x}, x19686x);
	defparam lut_4216.LUT_SIZE = 7;
	defparam lut_4216.mask = 128'h5555ffff5555ffff000033335fff7fff;

	lut_sub lut_4221 ({sk[929], i_14_, i_13_, i_12_, x898x, x904x}, x70x);
	defparam lut_4221.LUT_SIZE = 6;
	defparam lut_4221.mask = 64'h3f3f3f3f00000503;

	lut_sub lut_4224 ({sk[930], i_7_, i_8_, i_6_, n_n108, x909x, x70x}, n_n4826);
	defparam lut_4224.LUT_SIZE = 7;
	defparam lut_4224.mask = 128'h5555ffff5555ffff0000000003001100;

	lut_sub lut_4227 ({sk[931], i_9_, i_10_}, n_n269);
	defparam lut_4227.LUT_SIZE = 3;
	defparam lut_4227.mask = 8'h51;

	lut_sub lut_4229 ({sk[932], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x125x);
	defparam lut_4229.LUT_SIZE = 7;
	defparam lut_4229.mask = 128'h5555ffff5555ffff0010001040000000;

	lut_sub lut_4233 ({sk[933], i_7_, i_8_, i_6_, x909x, x176x}, n_n4823);
	defparam lut_4233.LUT_SIZE = 6;
	defparam lut_4233.mask = 64'h3f3f3f3f00000010;

	lut_sub lut_4235 ({sk[934], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x90x);
	defparam lut_4235.LUT_SIZE = 7;
	defparam lut_4235.mask = 128'h5555ffff5555ffff1040004000000000;

	lut_sub lut_4239 ({sk[935], i_14_, i_13_, i_12_, i_15_, x899x, n_n259}, x1922x);
	defparam lut_4239.LUT_SIZE = 7;
	defparam lut_4239.mask = 128'h5555ffff5555ffff0000000005337350;

	lut_sub lut_4245 ({sk[936], i_7_, i_8_, i_6_, n_n110, x909x, x1922x}, x733x);
	defparam lut_4245.LUT_SIZE = 7;
	defparam lut_4245.mask = 128'h5555ffff5555ffff0000000011000300;

	lut_sub lut_4248 ({sk[937], i_9_, i_10_, i_11_}, n_n259);
	defparam lut_4248.LUT_SIZE = 4;
	defparam lut_4248.mask = 16'h5502;

	lut_sub lut_4250 ({sk[938], i_14_, i_13_, i_12_, i_15_, x905x, n_n259}, x258x);
	defparam lut_4250.LUT_SIZE = 7;
	defparam lut_4250.mask = 128'h5555ffff5555ffff0533005000000000;

	lut_sub lut_4254 ({sk[939], i_7_, i_8_, i_6_, x146x, x909x}, n_n4815);
	defparam lut_4254.LUT_SIZE = 6;
	defparam lut_4254.mask = 64'h3f3f3f3f00000010;

	lut_sub lut_4256 ({sk[940], i_7_, i_8_, i_6_, n_n281, x909x, x908x}, x522x);
	defparam lut_4256.LUT_SIZE = 7;
	defparam lut_4256.mask = 128'h5555ffff5555ffff0000000000000100;

	lut_sub lut_4258 ({sk[941], i_14_, i_13_, i_12_, x914x, x912x}, x265x);
	defparam lut_4258.LUT_SIZE = 6;
	defparam lut_4258.mask = 64'h3f3f3f3f30500300;

	lut_sub lut_4262 ({sk[942], i_9_, i_10_, i_11_, i_15_, n_n220, x101x}, x293x);
	defparam lut_4262.LUT_SIZE = 7;
	defparam lut_4262.mask = 128'h5555ffff5555ffff5755555555555555;

	lut_sub lut_4265 ({sk[943], i_14_, i_13_, i_12_, x912x}, n_n11);
	defparam lut_4265.LUT_SIZE = 5;
	defparam lut_4265.mask = 32'h0f0f0001;

	lut_sub lut_4267 ({sk[944], n_n106, n_n6, n_n5, x101x, n_n11, x113x}, x498x);
	defparam lut_4267.LUT_SIZE = 7;
	defparam lut_4267.mask = 128'h5555ffff5555ffff00335f7f00ff5fff;

	lut_sub lut_4272 ({sk[945], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, n_n138);
	defparam lut_4272.LUT_SIZE = 7;
	defparam lut_4272.mask = 128'h5555ffff5555ffff0000000800000000;

	lut_sub lut_4274 ({sk[946], i_9_, i_10_, i_11_, i_15_, n_n258, n_n138}, x60x);
	defparam lut_4274.LUT_SIZE = 7;
	defparam lut_4274.mask = 128'h5555ffff5555ffff0505070505050505;

	lut_sub lut_4277 ({sk[947], i_7_, i_8_, i_6_, x909x, x60x}, x5259x);
	defparam lut_4277.LUT_SIZE = 6;
	defparam lut_4277.mask = 64'h3f3f3f3f00000010;

	lut_sub lut_4279 ({sk[948], i_14_, i_13_, i_12_, x913x, x909x, n_n263}, x5260x);
	defparam lut_4279.LUT_SIZE = 7;
	defparam lut_4279.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_4281 ({sk[949], i_14_, i_13_, i_12_, x906x}, x166x);
	defparam lut_4281.LUT_SIZE = 5;
	defparam lut_4281.mask = 32'h0f0f0045;

	lut_sub lut_4285 ({sk[950], i_14_, i_13_, i_12_, x900x}, x180x);
	defparam lut_4285.LUT_SIZE = 5;
	defparam lut_4285.mask = 32'h0f0f5100;

	lut_sub lut_4289 ({sk[951], i_14_, i_13_, i_12_, x900x}, x224x);
	defparam lut_4289.LUT_SIZE = 5;
	defparam lut_4289.mask = 32'h0f0f0054;

	lut_sub lut_4293 ({sk[952], i_7_, i_8_, i_6_, x909x, x224x}, n_n4966);
	defparam lut_4293.LUT_SIZE = 6;
	defparam lut_4293.mask = 64'h3f3f3f3f00000100;

	lut_sub lut_4295 ({sk[953], i_14_, i_13_, i_12_, n_n266, x909x, x904x}, x484x);
	defparam lut_4295.LUT_SIZE = 7;
	defparam lut_4295.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_4298 ({sk[954], i_14_, i_13_, i_12_, n_n266, x909x, x904x}, n_n4967);
	defparam lut_4298.LUT_SIZE = 7;
	defparam lut_4298.mask = 128'h5555ffff5555ffff0001010100000000;

	lut_sub lut_4302 ({sk[955], i_14_, i_13_, i_12_, x904x}, x41x);
	defparam lut_4302.LUT_SIZE = 5;
	defparam lut_4302.mask = 32'h0f0f0045;

	lut_sub lut_4306 ({sk[956], n_n266, n_n271, x909x, x166x, x99x, x41x}, x20703x);
	defparam lut_4306.LUT_SIZE = 7;
	defparam lut_4306.mask = 128'h5555ffff5555ffff0000000f007f007f;

	lut_sub lut_4311 ({sk[957], n_n57, n_n56, x153x, x180x, x224x, n_n4967}, x20704x);
	defparam lut_4311.LUT_SIZE = 7;
	defparam lut_4311.mask = 128'h5555ffff5555ffff55557fff77777fff;

	lut_sub lut_4317 ({sk[958], i_14_, i_13_, i_12_, x911x}, n_n150);
	defparam lut_4317.LUT_SIZE = 5;
	defparam lut_4317.mask = 32'h0f0f0400;

	lut_sub lut_4319 ({sk[959], i_7_, i_8_, i_6_, x909x, x72x}, x5037x);
	defparam lut_4319.LUT_SIZE = 6;
	defparam lut_4319.mask = 64'h3f3f3f3f00000100;

	lut_sub lut_4321 ({sk[960], i_14_, i_13_, i_12_, x898x}, n_n50);
	defparam lut_4321.LUT_SIZE = 5;
	defparam lut_4321.mask = 32'h0f0f4000;

	lut_sub lut_4323 ({sk[961], i_14_, i_13_, i_12_, x909x, n_n261, x904x}, x389x);
	defparam lut_4323.LUT_SIZE = 7;
	defparam lut_4323.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_4326 ({sk[962], i_14_, i_13_, i_12_, x909x, x898x, n_n261}, x632x);
	defparam lut_4326.LUT_SIZE = 7;
	defparam lut_4326.mask = 128'h5555ffff5555ffff0000000000010100;

	lut_sub lut_4329 ({sk[963], i_14_, i_13_, i_12_, x898x, x904x}, x1911x);
	defparam lut_4329.LUT_SIZE = 6;
	defparam lut_4329.mask = 64'h3f3f3f3f00007055;

	lut_sub lut_4334 ({sk[964], i_14_, i_13_, i_12_, x906x}, x76x);
	defparam lut_4334.LUT_SIZE = 5;
	defparam lut_4334.mask = 32'h0f0f0005;

	lut_sub lut_4337 ({sk[965], i_14_, i_13_, i_12_, i_15_, n_n267}, x81x);
	defparam lut_4337.LUT_SIZE = 6;
	defparam lut_4337.mask = 64'h3f3f3f3f00000110;

	lut_sub lut_4340 ({sk[966], i_14_, i_13_, i_12_, x900x}, n_n93);
	defparam lut_4340.LUT_SIZE = 5;
	defparam lut_4340.mask = 32'h0f0f0040;

	lut_sub lut_4342 ({sk[967], i_14_, i_13_, i_12_, x898x, x904x}, x1907x);
	defparam lut_4342.LUT_SIZE = 6;
	defparam lut_4342.mask = 64'h3f3f3f3f00007375;

	lut_sub lut_4349 ({sk[968], i_14_, i_13_, i_12_, x900x, x906x}, x1908x);
	defparam lut_4349.LUT_SIZE = 6;
	defparam lut_4349.mask = 64'h3f3f3f3f37570000;

	lut_sub lut_4356 ({sk[969], i_7_, i_8_, i_6_, x909x, x113x}, x5021x);
	defparam lut_4356.LUT_SIZE = 6;
	defparam lut_4356.mask = 64'h3f3f3f3f00000001;

	lut_sub lut_4358 ({sk[970], i_7_, i_8_, i_6_, x146x, x909x, x265x}, x734x);
	defparam lut_4358.LUT_SIZE = 7;
	defparam lut_4358.mask = 128'h5555ffff5555ffff0000000000110003;

	lut_sub lut_4361 ({sk[971], i_14_, i_13_, i_12_, x905x, x899x}, x1870x);
	defparam lut_4361.LUT_SIZE = 6;
	defparam lut_4361.mask = 64'h3f3f3f3f30500305;

	lut_sub lut_4366 ({sk[972], i_7_, i_8_, i_6_, x922x}, n_n48);
	defparam lut_4366.LUT_SIZE = 5;
	defparam lut_4366.mask = 32'h0f0f4000;

	lut_sub lut_4368 ({sk[973], i_14_, i_13_, i_12_, x906x}, n_n42);
	defparam lut_4368.LUT_SIZE = 5;
	defparam lut_4368.mask = 32'h0f0f0400;

	lut_sub lut_4370 ({sk[974], i_7_, i_8_, i_6_, n_n258, x922x, x900x}, x619x);
	defparam lut_4370.LUT_SIZE = 7;
	defparam lut_4370.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_4372 ({sk[975], i_14_, i_13_, i_12_, x903x}, n_n73);
	defparam lut_4372.LUT_SIZE = 5;
	defparam lut_4372.mask = 32'h0f0f1000;

	lut_sub lut_4374 ({sk[976], i_14_, i_13_, i_12_, x903x}, n_n22);
	defparam lut_4374.LUT_SIZE = 5;
	defparam lut_4374.mask = 32'h0f0f0400;

	lut_sub lut_4376 ({sk[977], i_7_, i_8_, i_6_, x922x, x40x}, x4600x);
	defparam lut_4376.LUT_SIZE = 6;
	defparam lut_4376.mask = 64'h3f3f3f3f00100000;

	lut_sub lut_4378 ({sk[978], i_14_, i_13_, i_12_, n_n273, x922x, x899x}, n_n6860);
	defparam lut_4378.LUT_SIZE = 7;
	defparam lut_4378.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_4380 ({sk[979], i_14_, i_13_, i_12_, x901x}, n_n84);
	defparam lut_4380.LUT_SIZE = 5;
	defparam lut_4380.mask = 32'h0f0f0040;

	lut_sub lut_4382 ({sk[980], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x89x);
	defparam lut_4382.LUT_SIZE = 7;
	defparam lut_4382.mask = 128'h5555ffff5555ffff0000000010000040;

	lut_sub lut_4385 ({sk[981], n_n273, n_n222, x922x, x901x, x89x}, n_n4094);
	defparam lut_4385.LUT_SIZE = 6;
	defparam lut_4385.mask = 64'h3f3f3f3f00000507;

	lut_sub lut_4388 ({sk[982], i_7_, i_8_, i_6_, x916x, n_n258, x900x}, n_n7224);
	defparam lut_4388.LUT_SIZE = 7;
	defparam lut_4388.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_4390 ({sk[983], i_7_, i_8_, i_6_, x916x, n_n222, x900x}, n_n7225);
	defparam lut_4390.LUT_SIZE = 7;
	defparam lut_4390.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_4392 ({sk[984], i_14_, i_13_, i_12_, x914x}, x67x);
	defparam lut_4392.LUT_SIZE = 5;
	defparam lut_4392.mask = 32'h0f0f1400;

	lut_sub lut_4395 ({sk[985], i_14_, i_13_, i_12_, n_n283, x922x, x901x}, x623x);
	defparam lut_4395.LUT_SIZE = 7;
	defparam lut_4395.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_4397 ({sk[986], i_9_, i_10_, i_11_, n_n261, x922x}, x407x);
	defparam lut_4397.LUT_SIZE = 6;
	defparam lut_4397.mask = 64'h3f3f3f3f10000000;

	lut_sub lut_4399 ({sk[987], i_9_, i_10_, i_11_, n_n263, x922x}, x457x);
	defparam lut_4399.LUT_SIZE = 6;
	defparam lut_4399.mask = 64'h3f3f3f3f00001000;

	lut_sub lut_4401 ({sk[988], i_7_, i_8_, i_6_, n_n104, x922x, n_n282}, x20333x);
	defparam lut_4401.LUT_SIZE = 7;
	defparam lut_4401.mask = 128'h5555ffff5555ffff0000030000001100;

	lut_sub lut_4404 ({sk[989], i_14_, i_13_, i_12_, n_n273, x922x, x908x}, n_n6872);
	defparam lut_4404.LUT_SIZE = 7;
	defparam lut_4404.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_4406 ({sk[990], i_14_, i_13_, i_12_, n_n273, x905x, x922x}, n_n6871);
	defparam lut_4406.LUT_SIZE = 7;
	defparam lut_4406.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_4408 ({sk[991], i_14_, i_13_, i_12_}, n_n256);
	defparam lut_4408.LUT_SIZE = 4;
	defparam lut_4408.mask = 16'h5540;

	lut_sub lut_4410 ({sk[992], i_7_, i_8_, i_6_, x905x, x922x, n_n256}, n_n6870);
	defparam lut_4410.LUT_SIZE = 7;
	defparam lut_4410.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_4412 ({sk[993], i_14_, i_13_, i_12_, n_n273, x905x, x922x}, x456x);
	defparam lut_4412.LUT_SIZE = 7;
	defparam lut_4412.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_4415 ({sk[994], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x117x);
	defparam lut_4415.LUT_SIZE = 7;
	defparam lut_4415.mask = 128'h5555ffff5555ffff0000001040004000;

	lut_sub lut_4419 ({sk[995], i_14_, i_13_, i_12_, i_15_, n_n53, n_n259}, x286x);
	defparam lut_4419.LUT_SIZE = 7;
	defparam lut_4419.mask = 128'h5555ffff5555ffff0100001000000000;

	lut_sub lut_4422 ({sk[996], n_n273, x922x, x899x, n_n256, x117x, x286x}, x864x);
	defparam lut_4422.LUT_SIZE = 7;
	defparam lut_4422.mask = 128'h5555ffff5555ffff555555555555777f;

	lut_sub lut_4426 ({sk[997], n_n273, n_n258, x922x, x456x, x864x, x908x}, n_n3964);
	defparam lut_4426.LUT_SIZE = 7;
	defparam lut_4426.mask = 128'h5555ffff5555ffff3f3f3f3f3f3f3f7f;

	lut_sub lut_4430 ({sk[998], i_7_, i_8_, i_6_, x916x, n_n228, x906x}, x518x);
	defparam lut_4430.LUT_SIZE = 7;
	defparam lut_4430.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_4432 ({sk[999], i_14_, i_13_, i_12_, n_n4, x900x, x906x}, n_n896);
	defparam lut_4432.LUT_SIZE = 7;
	defparam lut_4432.mask = 128'h5555ffff5555ffff0000000003000305;

	lut_sub lut_4436 ({sk[1000], i_14_, i_13_, i_12_, x904x}, n_n95);
	defparam lut_4436.LUT_SIZE = 5;
	defparam lut_4436.mask = 32'h0f0f0400;

	lut_sub lut_4438 ({sk[1001], i_7_, i_8_, i_6_, n_n220, x909x, x904x}, n_n6046);
	defparam lut_4438.LUT_SIZE = 7;
	defparam lut_4438.mask = 128'h5555ffff5555ffff0000000000000001;

	lut_sub lut_4440 ({sk[1002], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x106x);
	defparam lut_4440.LUT_SIZE = 7;
	defparam lut_4440.mask = 128'h5555ffff5555ffff1040004000000000;

	lut_sub lut_4444 ({sk[1003], i_14_, i_13_, i_12_, i_15_, x902x, n_n270}, x1861x);
	defparam lut_4444.LUT_SIZE = 7;
	defparam lut_4444.mask = 128'h5555ffff5555ffff0000000005337350;

	lut_sub lut_4450 ({sk[1004], i_14_, i_13_, i_12_, n_n271, x914x, x909x}, x520x);
	defparam lut_4450.LUT_SIZE = 7;
	defparam lut_4450.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_4452 ({sk[1005], n_n266, n_n271, x909x, x106x, x1861x, x520x}, n_n3204);
	defparam lut_4452.LUT_SIZE = 7;
	defparam lut_4452.mask = 128'h5555ffff5555ffff5555555f5577557f;

	lut_sub lut_4456 ({sk[1006], i_14_, i_13_, i_12_, x914x}, n_n246);
	defparam lut_4456.LUT_SIZE = 5;
	defparam lut_4456.mask = 32'h0f0f0010;

	lut_sub lut_4458 ({sk[1007], i_14_, i_13_, i_12_, x914x, x912x}, x160x);
	defparam lut_4458.LUT_SIZE = 6;
	defparam lut_4458.mask = 64'h3f3f3f3f00000305;

	lut_sub lut_4461 ({sk[1008], i_14_, i_13_, i_12_, n_n3, x898x}, n_n7406);
	defparam lut_4461.LUT_SIZE = 6;
	defparam lut_4461.mask = 64'h3f3f3f3f00100000;

	lut_sub lut_4463 ({sk[1009], i_14_, i_13_, i_12_, n_n3, x904x}, n_n7405);
	defparam lut_4463.LUT_SIZE = 6;
	defparam lut_4463.mask = 64'h3f3f3f3f00000100;

	lut_sub lut_4465 ({sk[1010], i_14_, i_13_, i_12_, n_n266, x909x, x905x}, n_n6190);
	defparam lut_4465.LUT_SIZE = 7;
	defparam lut_4465.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_4467 ({sk[1011], i_14_, i_13_, i_12_, n_n271, x909x, x905x}, x720x);
	defparam lut_4467.LUT_SIZE = 7;
	defparam lut_4467.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_4469 ({sk[1012], i_14_, i_13_, i_12_, x898x}, n_n14);
	defparam lut_4469.LUT_SIZE = 5;
	defparam lut_4469.mask = 32'h0f0f0400;

	lut_sub lut_4471 ({sk[1013], i_14_, i_13_, i_12_, x898x, x904x}, x44x);
	defparam lut_4471.LUT_SIZE = 6;
	defparam lut_4471.mask = 64'h3f3f3f3f50300000;

	lut_sub lut_4474 ({sk[1014], i_14_, i_13_, i_12_, x899x}, x82x);
	defparam lut_4474.LUT_SIZE = 5;
	defparam lut_4474.mask = 32'h0f0f0014;

	lut_sub lut_4477 ({sk[1015], i_14_, i_13_, i_12_, x898x, x121x}, x1897x);
	defparam lut_4477.LUT_SIZE = 6;
	defparam lut_4477.mask = 64'h3f3f3f3f55555557;

	lut_sub lut_4480 ({sk[1016], i_7_, i_8_, i_6_, x909x, x111x}, x636x);
	defparam lut_4480.LUT_SIZE = 6;
	defparam lut_4480.mask = 64'h3f3f3f3f00000100;

	lut_sub lut_4482 ({sk[1017], i_14_, i_13_, i_12_, i_15_, x905x, n_n259}, x1898x);
	defparam lut_4482.LUT_SIZE = 7;
	defparam lut_4482.mask = 128'h5555ffff5555ffff0537005550000000;

	lut_sub lut_4489 ({sk[1018], x206x, n_n57, x258x, x720x, x44x, x70x}, x21070x);
	defparam lut_4489.LUT_SIZE = 7;
	defparam lut_4489.mask = 128'h5555ffff5555ffff0f0f7fff0f0fffff;

	lut_sub lut_4495 ({sk[1019], n_n56, n_n6190, x82x, x1897x, x111x, x1898x}, x21071x);
	defparam lut_4495.LUT_SIZE = 7;
	defparam lut_4495.mask = 128'h5555ffff5555ffff0000ffff7fffffff;

	lut_sub lut_4501 ({sk[1020], i_14_, i_13_, i_12_, x909x, n_n263, x904x}, x539x);
	defparam lut_4501.LUT_SIZE = 7;
	defparam lut_4501.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_4503 ({sk[1021], i_14_, i_13_, i_12_, i_15_, n_n247, x160x}, x977x);
	defparam lut_4503.LUT_SIZE = 7;
	defparam lut_4503.mask = 128'h5555ffff5555ffff7555575555555555;

	lut_sub lut_4507 ({sk[1022], n_n281, x909x, n_n263, x904x, n_n228, x912x}, x20950x);
	defparam lut_4507.LUT_SIZE = 7;
	defparam lut_4507.mask = 128'h5555ffff5555ffff000000110000001f;

	lut_sub lut_4510 ({sk[1023], x909x, x173x, n_n261, n_n263, x977x, x20950x}, n_n3172);
	defparam lut_4510.LUT_SIZE = 7;
	defparam lut_4510.mask = 128'h5555ffff5555ffff5555555555775f7f;

	lut_sub lut_4514 ({sk[1024], i_14_, i_13_, i_12_, x909x, n_n261, x899x}, x523x);
	defparam lut_4514.LUT_SIZE = 7;
	defparam lut_4514.mask = 128'h5555ffff5555ffff0000000000000001;

	lut_sub lut_4516 ({sk[1025], i_14_, i_13_, i_12_, x908x, x902x}, x208x);
	defparam lut_4516.LUT_SIZE = 6;
	defparam lut_4516.mask = 64'h3f3f3f3f30500000;

	lut_sub lut_4519 ({sk[1026], i_14_, i_13_, i_12_, x905x, x899x}, x314x);
	defparam lut_4519.LUT_SIZE = 6;
	defparam lut_4519.mask = 64'h3f3f3f3f00500305;

	lut_sub lut_4523 ({sk[1027], i_14_, i_13_, i_12_, i_15_, x199x, n_n259}, x978x);
	defparam lut_4523.LUT_SIZE = 7;
	defparam lut_4523.mask = 128'h5555ffff5555ffff3333373333733337;

	lut_sub lut_4528 ({sk[1028], x146x, x909x, n_n261, n_n263, x265x, x978x}, x20956x);
	defparam lut_4528.LUT_SIZE = 7;
	defparam lut_4528.mask = 128'h5555ffff5555ffff00000707000007ff;

	lut_sub lut_4532 ({sk[1029], i_14_, i_13_, i_12_, n_n3, x908x}, x3762x);
	defparam lut_4532.LUT_SIZE = 6;
	defparam lut_4532.mask = 64'h3f3f3f3f00100000;

	lut_sub lut_4534 ({sk[1030], i_14_, i_13_, i_12_, n_n208, x916x, x902x}, x374x);
	defparam lut_4534.LUT_SIZE = 7;
	defparam lut_4534.mask = 128'h5555ffff5555ffff0000000000010100;

	lut_sub lut_4537 ({sk[1031], i_14_, i_13_, i_12_, i_15_, x163x, n_n270}, x1959x);
	defparam lut_4537.LUT_SIZE = 7;
	defparam lut_4537.mask = 128'h5555ffff5555ffff3333333337337373;

	lut_sub lut_4542 ({sk[1032], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x979x);
	defparam lut_4542.LUT_SIZE = 7;
	defparam lut_4542.mask = 128'h5555ffff5555ffff0105400505010504;

	lut_sub lut_4555 ({sk[1033], i_14_, i_13_, i_12_, i_15_, n_n270}, x80x);
	defparam lut_4555.LUT_SIZE = 6;
	defparam lut_4555.mask = 64'h3f3f3f3f10040000;

	lut_sub lut_4558 ({sk[1034], i_7_, i_8_, i_6_, x916x, x908x, n_n256}, n_n7306);
	defparam lut_4558.LUT_SIZE = 7;
	defparam lut_4558.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_4560 ({sk[1035], i_14_, i_13_, i_12_, i_15_, n_n247, n_n137}, x136x);
	defparam lut_4560.LUT_SIZE = 7;
	defparam lut_4560.mask = 128'h5555ffff5555ffff5050505053505070;

	lut_sub lut_4564 ({sk[1036], i_14_, i_13_, i_12_, i_15_, x912x, n_n137}, x55x);
	defparam lut_4564.LUT_SIZE = 7;
	defparam lut_4564.mask = 128'h5555ffff5555ffff0505050505370505;

	lut_sub lut_4567 ({sk[1037], i_14_, i_13_, i_12_, i_15_, n_n247, x55x}, x980x);
	defparam lut_4567.LUT_SIZE = 7;
	defparam lut_4567.mask = 128'h5555ffff5555ffff5775557557557575;

	lut_sub lut_4575 ({sk[1038], i_14_, i_13_, i_12_, i_15_, x902x, n_n270}, x1858x);
	defparam lut_4575.LUT_SIZE = 7;
	defparam lut_4575.mask = 128'h5555ffff5555ffff0000000005337350;

	lut_sub lut_4581 ({sk[1039], n_n1, n_n2, n_n111, x93x, x163x, x1858x}, x20962x);
	defparam lut_4581.LUT_SIZE = 7;
	defparam lut_4581.mask = 128'h5555ffff5555ffff000000ff7f7f7fff;

	lut_sub lut_4586 ({sk[1040], n_n1, n_n2, n_n111, x106x, x93x, x980x}, x20963x);
	defparam lut_4586.LUT_SIZE = 7;
	defparam lut_4586.mask = 128'h5555ffff5555ffff000077770fff7fff;

	lut_sub lut_4591 ({sk[1041], i_14_, i_13_, i_12_, i_15_, x905x, n_n259}, x1923x);
	defparam lut_4591.LUT_SIZE = 7;
	defparam lut_4591.mask = 128'h5555ffff5555ffff0537005550000000;

	lut_sub lut_4598 ({sk[1042], i_7_, i_8_, i_6_, x915x, x111x, x1923x}, n_n2860);
	defparam lut_4598.LUT_SIZE = 7;
	defparam lut_4598.mask = 128'h5555ffff5555ffff0000070000000000;

	lut_sub lut_4601 ({sk[1043], i_14_, i_13_, i_12_, x908x, x902x, x80x}, x1899x);
	defparam lut_4601.LUT_SIZE = 7;
	defparam lut_4601.mask = 128'h5555ffff5555ffff557f55775f555555;

	lut_sub lut_4607 ({sk[1044], i_14_, i_13_, i_12_, i_15_, x908x, n_n270}, x1949x);
	defparam lut_4607.LUT_SIZE = 7;
	defparam lut_4607.mask = 128'h5555ffff5555ffff0533335000000000;

	lut_sub lut_4612 ({sk[1045], x915x, n_n273, n_n283, x170x, x1949x, x49x}, x20965x);
	defparam lut_4612.LUT_SIZE = 7;
	defparam lut_4612.mask = 128'h5555ffff5555ffff00000000005f337f;

	lut_sub lut_4616 ({sk[1046], i_14_, i_13_, i_12_, x898x, x904x}, x45x);
	defparam lut_4616.LUT_SIZE = 6;
	defparam lut_4616.mask = 64'h3f3f3f3f03035000;

	lut_sub lut_4620 ({sk[1047], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x204x);
	defparam lut_4620.LUT_SIZE = 7;
	defparam lut_4620.mask = 128'h5555ffff5555ffff0104000400000000;

	lut_sub lut_4624 ({sk[1048], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x171x);
	defparam lut_4624.LUT_SIZE = 7;
	defparam lut_4624.mask = 128'h5555ffff5555ffff0000000001000404;

	lut_sub lut_4628 ({sk[1049], x915x, n_n273, x45x, x204x, x171x}, n_n3162);
	defparam lut_4628.LUT_SIZE = 6;
	defparam lut_4628.mask = 64'h3f3f3f3f0000007f;

	lut_sub lut_4632 ({sk[1050], i_14_, i_13_, i_12_, x898x}, x68x);
	defparam lut_4632.LUT_SIZE = 5;
	defparam lut_4632.mask = 32'h0f0f0014;

	lut_sub lut_4635 ({sk[1051], i_14_, i_13_, i_12_, i_15_, x904x, n_n253}, x1873x);
	defparam lut_4635.LUT_SIZE = 7;
	defparam lut_4635.mask = 128'h5555ffff5555ffff0550335000000000;

	lut_sub lut_4640 ({sk[1052], i_15_, n_n258, x912x, x136x, n_n137}, x1947x);
	defparam lut_4640.LUT_SIZE = 6;
	defparam lut_4640.mask = 64'h3f3f3f3f333f777f;

	lut_sub lut_4644 ({sk[1053], n_n1, n_n2, n_n95, x68x, x45x, x171x}, x20968x);
	defparam lut_4644.LUT_SIZE = 7;
	defparam lut_4644.mask = 128'h5555ffff5555ffff00007f7f00ff7fff;

	lut_sub lut_4649 ({sk[1054], n_n1, n_n2, n_n3162, x1873x, x1947x, x20968x}, x20971x);
	defparam lut_4649.LUT_SIZE = 7;
	defparam lut_4649.mask = 128'h5555ffff5555ffff55ff5fff77ff7fff;

	lut_sub lut_4654 ({sk[1055], x915x, n_n273, n_n283, n_n76, x82x, x1899x}, x20964x);
	defparam lut_4654.LUT_SIZE = 7;
	defparam lut_4654.mask = 128'h5555ffff5555ffff00000000005f337f;

	lut_sub lut_4658 ({sk[1056], x20962x, x20963x, n_n2860, x20965x, x20964x}, x20972x);
	defparam lut_4658.LUT_SIZE = 6;
	defparam lut_4658.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_4664 ({sk[1057], i_14_, i_13_, i_12_, x907x}, n_n10);
	defparam lut_4664.LUT_SIZE = 5;
	defparam lut_4664.mask = 32'h0f0f0010;

	lut_sub lut_4666 ({sk[1058], i_14_, i_13_, i_12_, x907x, x915x, n_n261}, n_n6843);
	defparam lut_4666.LUT_SIZE = 7;
	defparam lut_4666.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_4668 ({sk[1059], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x84x);
	defparam lut_4668.LUT_SIZE = 7;
	defparam lut_4668.mask = 128'h5555ffff5555ffff0010001000000000;

	lut_sub lut_4671 ({sk[1060], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x155x);
	defparam lut_4671.LUT_SIZE = 7;
	defparam lut_4671.mask = 128'h5555ffff5555ffff0010001040000000;

	lut_sub lut_4675 ({sk[1061], i_14_, i_13_, i_12_, n_n273, x922x, x899x}, n_n6868);
	defparam lut_4675.LUT_SIZE = 7;
	defparam lut_4675.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_4677 ({sk[1062], i_14_, i_13_, i_12_, i_15_, x913x, n_n242}, x983x);
	defparam lut_4677.LUT_SIZE = 7;
	defparam lut_4677.mask = 128'h5555ffff5555ffff0533335055000000;

	lut_sub lut_4684 ({sk[1063], i_14_, i_13_, i_12_, x913x}, x62x);
	defparam lut_4684.LUT_SIZE = 5;
	defparam lut_4684.mask = 32'h0f0f1400;

	lut_sub lut_4687 ({sk[1064], i_14_, i_13_, i_12_, x899x}, n_n223);
	defparam lut_4687.LUT_SIZE = 5;
	defparam lut_4687.mask = 32'h0f0f0040;

	lut_sub lut_4689 ({sk[1065], x909x, n_n261, n_n263, x983x, x62x, n_n223}, n_n2136);
	defparam lut_4689.LUT_SIZE = 7;
	defparam lut_4689.mask = 128'h5555ffff5555ffff0000000000770f7f;

	lut_sub lut_4693 ({sk[1066], i_14_, i_13_, i_12_, x907x}, n_n35);
	defparam lut_4693.LUT_SIZE = 5;
	defparam lut_4693.mask = 32'h0f0f0040;

	lut_sub lut_4695 ({sk[1067], i_9_, i_10_, i_11_, i_15_, n_n279}, x252x);
	defparam lut_4695.LUT_SIZE = 6;
	defparam lut_4695.mask = 64'h3f3f3f3f50000000;

	lut_sub lut_4698 ({sk[1068], i_14_, i_13_, i_12_, x912x}, n_n179);
	defparam lut_4698.LUT_SIZE = 5;
	defparam lut_4698.mask = 32'h0f0f0040;

	lut_sub lut_4700 ({sk[1069], i_14_, i_13_, i_12_, x914x}, n_n113);
	defparam lut_4700.LUT_SIZE = 5;
	defparam lut_4700.mask = 32'h0f0f0040;

	lut_sub lut_4702 ({sk[1070], i_9_, i_10_, i_11_, i_15_, n_n279}, x329x);
	defparam lut_4702.LUT_SIZE = 6;
	defparam lut_4702.mask = 64'h3f3f3f3f00005000;

	lut_sub lut_4705 ({sk[1071], i_14_, i_13_, i_12_, n_n266, x914x, x909x}, x538x);
	defparam lut_4705.LUT_SIZE = 7;
	defparam lut_4705.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_4707 ({sk[1072], n_n266, n_n271, n_n111, x909x, n_n95, x106x}, x21444x);
	defparam lut_4707.LUT_SIZE = 7;
	defparam lut_4707.mask = 128'h5555ffff5555ffff00000303050f070f;

	lut_sub lut_4711 ({sk[1073], n_n266, n_n271, x909x, x252x, x329x, x21444x}, n_n2169);
	defparam lut_4711.LUT_SIZE = 7;
	defparam lut_4711.mask = 128'h5555ffff5555ffff5555555f5577557f;

	lut_sub lut_4715 ({sk[1074], i_7_, i_8_, i_6_, x909x}, x164x);
	defparam lut_4715.LUT_SIZE = 5;
	defparam lut_4715.mask = 32'h0f0f0044;

	lut_sub lut_4718 ({sk[1075], i_14_, i_13_, i_12_, x905x}, x83x);
	defparam lut_4718.LUT_SIZE = 5;
	defparam lut_4718.mask = 32'h0f0f1400;

	lut_sub lut_4721 ({sk[1076], i_7_, i_8_, i_6_, n_n281, x909x, x904x}, x21528x);
	defparam lut_4721.LUT_SIZE = 7;
	defparam lut_4721.mask = 128'h5555ffff5555ffff0000000001000100;

	lut_sub lut_4724 ({sk[1077], i_7_, i_8_, i_6_, n_n12, x909x, x21528x}, x21529x);
	defparam lut_4724.LUT_SIZE = 7;
	defparam lut_4724.mask = 128'h5555ffff5555ffff5555555557555755;

	lut_sub lut_4728 ({sk[1078], n_n148, n_n6, n_n5, n_n7, n_n60, x21532x}, x21533x);
	defparam lut_4728.LUT_SIZE = 7;
	defparam lut_4728.mask = 128'h5555ffff5555ffff557f5f7f55ffffff;

	lut_sub lut_4735 ({sk[1079], n_n5, n_n2136, x307x, x83x, x21529x, x21533x}, n_n2081);
	defparam lut_4735.LUT_SIZE = 7;
	defparam lut_4735.mask = 128'h5555ffff5555ffff7777ffff7fffffff;

	lut_sub lut_4741 ({sk[1080], i_14_, i_13_, i_12_, x905x}, n_n109);
	defparam lut_4741.LUT_SIZE = 5;
	defparam lut_4741.mask = 32'h0f0f0040;

	lut_sub lut_4743 ({sk[1081], i_14_, i_13_, i_12_, x905x, x899x}, x79x);
	defparam lut_4743.LUT_SIZE = 6;
	defparam lut_4743.mask = 64'h3f3f3f3f50030000;

	lut_sub lut_4746 ({sk[1082], i_14_, i_13_, i_12_, x911x}, n_n204);
	defparam lut_4746.LUT_SIZE = 5;
	defparam lut_4746.mask = 32'h0f0f0040;

	lut_sub lut_4748 ({sk[1083], i_9_, i_10_, i_11_}, n_n275);
	defparam lut_4748.LUT_SIZE = 4;
	defparam lut_4748.mask = 16'h5540;

	lut_sub lut_4750 ({sk[1084], i_14_, i_13_, i_12_, i_15_, x902x, n_n275}, x21371x);
	defparam lut_4750.LUT_SIZE = 7;
	defparam lut_4750.mask = 128'h5555ffff5555ffff0550505073000000;

	lut_sub lut_4757 ({sk[1085], i_14_, i_13_, i_12_, x912x}, n_n147);
	defparam lut_4757.LUT_SIZE = 5;
	defparam lut_4757.mask = 32'h0f0f0400;

	lut_sub lut_4759 ({sk[1086], i_14_, i_13_, i_12_, x915x, n_n263, x912x}, n_n6847);
	defparam lut_4759.LUT_SIZE = 7;
	defparam lut_4759.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_4761 ({sk[1087], i_14_, i_13_, i_12_, n_n273, x922x, x901x}, n_n6500);
	defparam lut_4761.LUT_SIZE = 7;
	defparam lut_4761.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_4763 ({sk[1088], i_14_, i_13_, i_12_, x907x}, n_n32);
	defparam lut_4763.LUT_SIZE = 5;
	defparam lut_4763.mask = 32'h0f0f0400;

	lut_sub lut_4765 ({sk[1089], i_7_, i_8_, i_6_, x907x, n_n220, x922x}, n_n6503);
	defparam lut_4765.LUT_SIZE = 7;
	defparam lut_4765.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_4767 ({sk[1090], i_14_, i_13_, i_12_, x902x}, n_n80);
	defparam lut_4767.LUT_SIZE = 5;
	defparam lut_4767.mask = 32'h0f0f0004;

	lut_sub lut_4769 ({sk[1091], i_7_, i_8_, i_6_, n_n220, x909x, x906x}, x5379x);
	defparam lut_4769.LUT_SIZE = 7;
	defparam lut_4769.mask = 128'h5555ffff5555ffff0000000001000000;

	lut_sub lut_4771 ({sk[1092], i_14_, i_13_, i_12_, x909x, n_n263, x908x}, x4716x);
	defparam lut_4771.LUT_SIZE = 7;
	defparam lut_4771.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_4774 ({sk[1093], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x990x);
	defparam lut_4774.LUT_SIZE = 7;
	defparam lut_4774.mask = 128'h5555ffff5555ffff1040400000105040;

	lut_sub lut_4782 ({sk[1094], i_14_, i_13_, i_12_, x901x}, x85x);
	defparam lut_4782.LUT_SIZE = 5;
	defparam lut_4782.mask = 32'h0f0f0014;

	lut_sub lut_4785 ({sk[1095], i_14_, i_13_, i_12_, n_n3, x911x}, x664x);
	defparam lut_4785.LUT_SIZE = 6;
	defparam lut_4785.mask = 64'h3f3f3f3f00000100;

	lut_sub lut_4787 ({sk[1096], i_14_, i_13_, i_12_, i_15_, n_n270, x182x}, x431x);
	defparam lut_4787.LUT_SIZE = 7;
	defparam lut_4787.mask = 128'h5555ffff5555ffff5755555555555555;

	lut_sub lut_4790 ({sk[1097], i_14_, i_13_, i_12_, i_15_, n_n242, x431x}, x993x);
	defparam lut_4790.LUT_SIZE = 7;
	defparam lut_4790.mask = 128'h5555ffff5555ffff5777755775557775;

	lut_sub lut_4801 ({sk[1098], i_9_, i_10_, i_11_, i_15_, x60x, n_n228}, x337x);
	defparam lut_4801.LUT_SIZE = 7;
	defparam lut_4801.mask = 128'h5555ffff5555ffff3333733333333333;

	lut_sub lut_4804 ({sk[1099], i_14_, i_13_, i_12_, i_15_, x337x, n_n259}, x992x);
	defparam lut_4804.LUT_SIZE = 7;
	defparam lut_4804.mask = 128'h5555ffff5555ffff3737333773337373;

	lut_sub lut_4812 ({sk[1100], n_n4, x485x, x3762x, x333x, x664x, x992x}, x21911x);
	defparam lut_4812.LUT_SIZE = 7;
	defparam lut_4812.mask = 128'h5555ffff5555ffff3fffffff7fffffff;

	lut_sub lut_4818 ({sk[1101], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x131x);
	defparam lut_4818.LUT_SIZE = 7;
	defparam lut_4818.mask = 128'h5555ffff5555ffff0010001040000000;

	lut_sub lut_4822 ({sk[1102], i_14_, i_13_, i_12_, i_15_, n_n247, n_n137}, x213x);
	defparam lut_4822.LUT_SIZE = 7;
	defparam lut_4822.mask = 128'h5555ffff5555ffff5050505370505050;

	lut_sub lut_4826 ({sk[1103], i_14_, i_13_, i_12_, i_15_, n_n282, n_n270}, x995x);
	defparam lut_4826.LUT_SIZE = 7;
	defparam lut_4826.mask = 128'h5555ffff5555ffff0735300550007370;

	lut_sub lut_4839 ({sk[1104], i_14_, i_13_, i_12_, x914x, x55x}, x303x);
	defparam lut_4839.LUT_SIZE = 6;
	defparam lut_4839.mask = 64'h3f3f3f3f55555557;

	lut_sub lut_4842 ({sk[1105], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x994x);
	defparam lut_4842.LUT_SIZE = 7;
	defparam lut_4842.mask = 128'h5555ffff5555ffff1050000000101040;

	lut_sub lut_4849 ({sk[1106], n_n6, n_n5, n_n111, x49x, x131x, x995x}, x22107x);
	defparam lut_4849.LUT_SIZE = 7;
	defparam lut_4849.mask = 128'h5555ffff5555ffff000000ff7f7f7fff;

	lut_sub lut_4854 ({sk[1107], i_7_, i_8_, i_6_, x914x, x909x, n_n256}, n_n6582);
	defparam lut_4854.LUT_SIZE = 7;
	defparam lut_4854.mask = 128'h5555ffff5555ffff0000000000000100;

	lut_sub lut_4856 ({sk[1108], i_7_, i_8_, i_6_, x909x, x85x}, x5376x);
	defparam lut_4856.LUT_SIZE = 6;
	defparam lut_4856.mask = 64'h3f3f3f3f00001000;

	lut_sub lut_4858 ({sk[1109], i_7_, i_8_, i_6_, x78x, x909x}, x4743x);
	defparam lut_4858.LUT_SIZE = 6;
	defparam lut_4858.mask = 64'h3f3f3f3f00001000;

	lut_sub lut_4860 ({sk[1110], i_14_, i_13_, i_12_, i_15_, n_n282, n_n253}, x997x);
	defparam lut_4860.LUT_SIZE = 7;
	defparam lut_4860.mask = 128'h5555ffff5555ffff0757500770003030;

	lut_sub lut_4873 ({sk[1111], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x996x);
	defparam lut_4873.LUT_SIZE = 7;
	defparam lut_4873.mask = 128'h5555ffff5555ffff1010001040105040;

	lut_sub lut_4882 ({sk[1112], n_n6, n_n111, n_n104, n_n6582, x5376x, x4743x}, x22112x);
	defparam lut_4882.LUT_SIZE = 7;
	defparam lut_4882.mask = 128'h5555ffff5555ffff7f7f7f7f7fffffff;

	lut_sub lut_4888 ({sk[1113], i_7_, i_8_, i_6_, x909x, n_n22, x49x}, n_n4846);
	defparam lut_4888.LUT_SIZE = 7;
	defparam lut_4888.mask = 128'h5555ffff5555ffff0000000005000300;

	lut_sub lut_4891 ({sk[1114], i_14_, i_13_, i_12_, x909x, n_n261, x908x}, x593x);
	defparam lut_4891.LUT_SIZE = 7;
	defparam lut_4891.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_4894 ({sk[1115], i_14_, i_13_, i_12_, i_15_, n_n275, x897x}, x999x);
	defparam lut_4894.LUT_SIZE = 7;
	defparam lut_4894.mask = 128'h5555ffff5555ffff0333000330557530;

	lut_sub lut_4904 ({sk[1116], i_14_, i_13_, i_12_, i_15_, x908x, n_n275}, x998x);
	defparam lut_4904.LUT_SIZE = 7;
	defparam lut_4904.mask = 128'h5555ffff5555ffff0550500033007773;

	lut_sub lut_4914 ({sk[1117], n_n103, x909x, n_n263, n_n4846, x92x, x593x}, x22117x);
	defparam lut_4914.LUT_SIZE = 7;
	defparam lut_4914.mask = 128'h5555ffff5555ffff5f5f5f7f5f5f5fff;

	lut_sub lut_4919 ({sk[1118], i_7_, i_8_, i_6_, x909x, x999x, x998x}, x22118x);
	defparam lut_4919.LUT_SIZE = 7;
	defparam lut_4919.mask = 128'h5555ffff5555ffff0000000005000300;

	lut_sub lut_4922 ({sk[1119], n_n6, n_n5, x213x, x994x, x997x, x996x}, x24089x);
	defparam lut_4922.LUT_SIZE = 7;
	defparam lut_4922.mask = 128'h5555ffff5555ffffffffc000aaaa8000;

	lut_sub lut_4927 ({sk[1120], x22107x, x22112x, x22117x, x22118x, x24089x}, n_n1095);
	defparam lut_4927.LUT_SIZE = 6;
	defparam lut_4927.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_4933 ({sk[1121], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1056x);
	defparam lut_4933.LUT_SIZE = 7;
	defparam lut_4933.mask = 128'h5555ffff5555ffff0001000104000504;

	lut_sub lut_4940 ({sk[1122], i_14_, i_13_, i_12_, n_n283, x914x, x922x}, x22125x);
	defparam lut_4940.LUT_SIZE = 7;
	defparam lut_4940.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_4943 ({sk[1123], x909x, n_n261, n_n48, x213x, x1056x, x22125x}, x22130x);
	defparam lut_4943.LUT_SIZE = 7;
	defparam lut_4943.mask = 128'h5555ffff5555ffff555f555f555f777f;

	lut_sub lut_4947 ({sk[1124], i_14_, i_13_, i_12_, x907x, x911x}, x1057x);
	defparam lut_4947.LUT_SIZE = 6;
	defparam lut_4947.mask = 64'h3f3f3f3f00500033;

	lut_sub lut_4951 ({sk[1125], n_n273, n_n283, n_n222, x922x, x901x, x223x}, x24190x);
	defparam lut_4951.LUT_SIZE = 7;
	defparam lut_4951.mask = 128'h5555ffff5555fffffffffafafffcfaf8;

	lut_sub lut_4959 ({sk[1126], n_n273, x922x, x457x, x20333x, x1057x, x24190x}, x22142x);
	defparam lut_4959.LUT_SIZE = 7;
	defparam lut_4959.mask = 128'h5555ffff5555ffffafffafffafffbfff;

	lut_sub lut_4964 ({sk[1127], i_7_, i_8_, i_6_, x909x, n_n258, x898x}, x748x);
	defparam lut_4964.LUT_SIZE = 7;
	defparam lut_4964.mask = 128'h5555ffff5555ffff0000000001000000;

	lut_sub lut_4966 ({sk[1128], i_14_, i_13_, i_12_, i_15_, n_n253, n_n267}, x1001x);
	defparam lut_4966.LUT_SIZE = 7;
	defparam lut_4966.mask = 128'h5555ffff5555ffff0555000550057770;

	lut_sub lut_4979 ({sk[1129], i_14_, i_13_, i_12_, x898x, x900x, x906x}, x1000x);
	defparam lut_4979.LUT_SIZE = 7;
	defparam lut_4979.mask = 128'h5555ffff5555ffff3f33003355005555;

	lut_sub lut_4987 ({sk[1130], n_n6, x51x, x389x, x81x, x5379x, x748x}, x22148x);
	defparam lut_4987.LUT_SIZE = 7;
	defparam lut_4987.mask = 128'h5555ffff5555ffff77ff77ff7fffffff;

	lut_sub lut_4993 ({sk[1131], x909x, n_n261, n_n263, x1001x, x1000x, x22148x}, x22150x);
	defparam lut_4993.LUT_SIZE = 7;
	defparam lut_4993.mask = 128'h5555ffff5555ffff55555555555f777f;

	lut_sub lut_4997 ({sk[1132], n_n280, n_n53, x131x, x461x, x376x, x2687x}, n_n1240);
	defparam lut_4997.LUT_SIZE = 7;
	defparam lut_4997.mask = 128'h5555ffff5555ffff7f7f7fff7f7fffff;

	lut_sub lut_5003 ({sk[1133], n_n48, n_n53, n_n6879, x679x, x1338x, x1337x}, n_n1242);
	defparam lut_5003.LUT_SIZE = 7;
	defparam lut_5003.mask = 128'h5555ffff5555ffff0fff3fff5fff7fff;

	lut_sub lut_5008 ({sk[1134], n_n48, n_n6517, n_n6520, x50x, x22134x, x22136x}, n_n1243);
	defparam lut_5008.LUT_SIZE = 7;
	defparam lut_5008.mask = 128'h5555ffff5555ffff77ffffff7fffffff;

	lut_sub lut_5014 ({sk[1135], n_n6524, n_n6517, n_n6520, n_n6511, n_n6512, x631x}, x22129x);
	defparam lut_5014.LUT_SIZE = 7;
	defparam lut_5014.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_5021 ({sk[1136], x22130x, x22142x, n_n1240, n_n1242, n_n1243, x22129x}, x22151x);
	defparam lut_5021.LUT_SIZE = 7;
	defparam lut_5021.mask = 128'h5555ffff5555ffff7fffffffffffffff;

	lut_sub lut_5028 ({sk[1137], i_14_, i_13_, i_12_, x897x}, x56x);
	defparam lut_5028.LUT_SIZE = 5;
	defparam lut_5028.mask = 32'h0f0f0014;

	lut_sub lut_5031 ({sk[1138], i_7_, i_8_, i_6_, x922x, x56x}, x5627x);
	defparam lut_5031.LUT_SIZE = 6;
	defparam lut_5031.mask = 64'h3f3f3f3f00100000;

	lut_sub lut_5033 ({sk[1139], i_14_, i_13_, i_12_, i_15_, n_n242, n_n259}, x1489x);
	defparam lut_5033.LUT_SIZE = 7;
	defparam lut_5033.mask = 128'h5555ffff5555ffff0000000550007370;

	lut_sub lut_5041 ({sk[1140], i_14_, i_13_, i_12_, i_15_, x902x, n_n242}, x1488x);
	defparam lut_5041.LUT_SIZE = 7;
	defparam lut_5041.mask = 128'h5555ffff5555ffff3705000550005050;

	lut_sub lut_5049 ({sk[1141], i_7_, i_8_, i_6_, x922x, x1489x, x1488x}, x22159x);
	defparam lut_5049.LUT_SIZE = 7;
	defparam lut_5049.mask = 128'h5555ffff5555ffff0500030000000000;

	lut_sub lut_5052 ({sk[1142], i_14_, i_13_, i_12_, i_15_, n_n267}, x73x);
	defparam lut_5052.LUT_SIZE = 6;
	defparam lut_5052.mask = 64'h3f3f3f3f00100400;

	lut_sub lut_5055 ({sk[1143], i_14_, i_13_, i_12_, i_15_, x907x, n_n259}, x22167x);
	defparam lut_5055.LUT_SIZE = 7;
	defparam lut_5055.mask = 128'h5555ffff5555ffff0000500550335000;

	lut_sub lut_5061 ({sk[1144], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x22166x);
	defparam lut_5061.LUT_SIZE = 7;
	defparam lut_5061.mask = 128'h5555ffff5555ffff0050010000040000;

	lut_sub lut_5066 ({sk[1145], n_n283, x922x, n_n107, x73x, x22167x, x22166x}, x2638x);
	defparam lut_5066.LUT_SIZE = 7;
	defparam lut_5066.mask = 128'h5555ffff5555ffff0000000000007fff;

	lut_sub lut_5071 ({sk[1146], i_14_, i_13_, i_12_, x913x, x911x}, x324x);
	defparam lut_5071.LUT_SIZE = 6;
	defparam lut_5071.mask = 64'h3f3f3f3f53300000;

	lut_sub lut_5075 ({sk[1147], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1533x);
	defparam lut_5075.LUT_SIZE = 7;
	defparam lut_5075.mask = 128'h5555ffff5555ffff0000005353000053;

	lut_sub lut_5082 ({sk[1148], n_n283, x905x, x922x, x82x, n_n228}, x24208x);
	defparam lut_5082.LUT_SIZE = 6;
	defparam lut_5082.mask = 64'h3f3f3f3ffffffcf8;

	lut_sub lut_5087 ({sk[1149], n_n273, x922x, x155x, x324x, x1533x, x24208x}, x22169x);
	defparam lut_5087.LUT_SIZE = 7;
	defparam lut_5087.mask = 128'h5555ffff5555ffffaaaaaaaaaaaabfff;

	lut_sub lut_5092 ({sk[1150], i_14_, i_13_, i_12_, i_15_, x902x, n_n270}, x22170x);
	defparam lut_5092.LUT_SIZE = 7;
	defparam lut_5092.mask = 128'h5555ffff5555ffff0000000000007350;

	lut_sub lut_5096 ({sk[1151], i_14_, i_13_, i_12_, i_15_, n_n275, x22170x}, x1003x);
	defparam lut_5096.LUT_SIZE = 7;
	defparam lut_5096.mask = 128'h5555ffff5555ffff5777555775577775;

	lut_sub lut_5107 ({sk[1152], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x212x);
	defparam lut_5107.LUT_SIZE = 7;
	defparam lut_5107.mask = 128'h5555ffff5555ffff0101000100000000;

	lut_sub lut_5111 ({sk[1153], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1002x);
	defparam lut_5111.LUT_SIZE = 7;
	defparam lut_5111.mask = 128'h5555ffff5555ffff0101000104000404;

	lut_sub lut_5118 ({sk[1154], n_n108, n_n216, x60x, n_n48, n_n53, x62x}, x22156x);
	defparam lut_5118.LUT_SIZE = 7;
	defparam lut_5118.mask = 128'h5555ffff5555ffff050f373f373f373f;

	lut_sub lut_5123 ({sk[1155], n_n6870, n_n6868, n_n6867, x406x, x621x}, x22157x);
	defparam lut_5123.LUT_SIZE = 6;
	defparam lut_5123.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_5129 ({sk[1156], x22159x, x2638x, x22169x, x22156x, x22157x}, x22177x);
	defparam lut_5129.LUT_SIZE = 6;
	defparam lut_5129.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_5135 ({sk[1157], i_14_, i_13_, i_12_, x914x}, n_n87);
	defparam lut_5135.LUT_SIZE = 5;
	defparam lut_5135.mask = 32'h0f0f0001;

	lut_sub lut_5137 ({sk[1158], i_14_, i_13_, i_12_, x908x}, n_n77);
	defparam lut_5137.LUT_SIZE = 5;
	defparam lut_5137.mask = 32'h0f0f0100;

	lut_sub lut_5139 ({sk[1159], i_14_, i_13_, i_12_, i_15_, x902x, n_n270}, x1860x);
	defparam lut_5139.LUT_SIZE = 7;
	defparam lut_5139.mask = 128'h5555ffff5555ffff0000000005053350;

	lut_sub lut_5144 ({sk[1160], i_14_, i_13_, i_12_, x915x, n_n261, x899x}, x552x);
	defparam lut_5144.LUT_SIZE = 7;
	defparam lut_5144.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5146 ({sk[1161], n_n197, n_n100, n_n94, x114x, x120x, x1860x}, n_n855);
	defparam lut_5146.LUT_SIZE = 7;
	defparam lut_5146.mask = 128'h5555ffff5555ffff005f337f005fffff;

	lut_sub lut_5151 ({sk[1162], i_7_, i_8_, i_6_, x915x, x912x, n_n225}, n_n6834);
	defparam lut_5151.LUT_SIZE = 7;
	defparam lut_5151.mask = 128'h5555ffff5555ffff0000000001000000;

	lut_sub lut_5153 ({sk[1163], i_14_, i_13_, i_12_, x915x, n_n261, x902x}, x881x);
	defparam lut_5153.LUT_SIZE = 7;
	defparam lut_5153.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5155 ({sk[1164], i_9_, i_10_, i_11_, i_15_, x91x, n_n225}, x1007x);
	defparam lut_5155.LUT_SIZE = 7;
	defparam lut_5155.mask = 128'h5555ffff5555ffff3377333373333333;

	lut_sub lut_5160 ({sk[1165], i_14_, i_13_, i_12_, i_15_, x902x, n_n270}, x201x);
	defparam lut_5160.LUT_SIZE = 7;
	defparam lut_5160.mask = 128'h5555ffff5555ffff0000000005003350;

	lut_sub lut_5164 ({sk[1166], x915x, n_n261, n_n263, x114x, x1007x, x201x}, x22655x);
	defparam lut_5164.LUT_SIZE = 7;
	defparam lut_5164.mask = 128'h5555ffff5555ffff0000000000335f7f;

	lut_sub lut_5168 ({sk[1167], i_14_, i_13_, i_12_, x907x, x901x}, x301x);
	defparam lut_5168.LUT_SIZE = 6;
	defparam lut_5168.mask = 64'h3f3f3f3f00070003;

	lut_sub lut_5172 ({sk[1168], i_14_, i_13_, i_12_, n_n283, x922x, x912x}, n_n6504);
	defparam lut_5172.LUT_SIZE = 7;
	defparam lut_5172.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5174 ({sk[1169], i_7_, i_8_, i_6_, i_15_, x922x, n_n137}, n_n6505);
	defparam lut_5174.LUT_SIZE = 7;
	defparam lut_5174.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_5176 ({sk[1170], i_15_, n_n283, n_n258, x922x, x912x, n_n137}, x461x);
	defparam lut_5176.LUT_SIZE = 7;
	defparam lut_5176.mask = 128'h5555ffff5555ffff0000000300000507;

	lut_sub lut_5179 ({sk[1171], i_14_, i_13_, i_12_, x914x, x912x}, x304x);
	defparam lut_5179.LUT_SIZE = 6;
	defparam lut_5179.mask = 64'h3f3f3f3f00070003;

	lut_sub lut_5183 ({sk[1172], n_n48, n_n53, n_n179, x301x, x461x, x304x}, n_n824);
	defparam lut_5183.LUT_SIZE = 7;
	defparam lut_5183.mask = 128'h5555ffff5555ffff33333f3f77ff7fff;

	lut_sub lut_5188 ({sk[1173], i_7_, i_8_, i_6_, x909x, n_n258, x898x}, n_n6524);
	defparam lut_5188.LUT_SIZE = 7;
	defparam lut_5188.mask = 128'h5555ffff5555ffff0000000000000100;

	lut_sub lut_5190 ({sk[1174], i_7_, i_8_, i_6_, x922x, x901x, n_n228}, x495x);
	defparam lut_5190.LUT_SIZE = 7;
	defparam lut_5190.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_5192 ({sk[1175], i_14_, i_13_, i_12_, i_15_, n_n267}, x108x);
	defparam lut_5192.LUT_SIZE = 6;
	defparam lut_5192.mask = 64'h3f3f3f3f00001014;

	lut_sub lut_5196 ({sk[1176], x909x, n_n258, n_n261, x900x, x108x}, x670x);
	defparam lut_5196.LUT_SIZE = 6;
	defparam lut_5196.mask = 64'h3f3f3f3f00000507;

	lut_sub lut_5199 ({sk[1177], i_14_, i_13_, i_12_, x900x, x906x, x108x}, x1010x);
	defparam lut_5199.LUT_SIZE = 7;
	defparam lut_5199.mask = 128'h5555ffff5555ffff5555557f555f5555;

	lut_sub lut_5204 ({sk[1178], i_9_, i_10_, i_11_, i_15_, n_n225}, x134x);
	defparam lut_5204.LUT_SIZE = 6;
	defparam lut_5204.mask = 64'h3f3f3f3f00000005;

	lut_sub lut_5207 ({sk[1179], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x202x);
	defparam lut_5207.LUT_SIZE = 7;
	defparam lut_5207.mask = 128'h5555ffff5555ffff0000000001000104;

	lut_sub lut_5211 ({sk[1180], x909x, n_n261, n_n263, x1010x, x134x, x202x}, x22723x);
	defparam lut_5211.LUT_SIZE = 7;
	defparam lut_5211.mask = 128'h5555ffff5555ffff00000000000f777f;

	lut_sub lut_5215 ({sk[1181], i_13_, i_12_}, n_n254);
	defparam lut_5215.LUT_SIZE = 3;
	defparam lut_5215.mask = 8'h51;

	lut_sub lut_5217 ({sk[1182], i_7_, i_8_, i_6_, x909x}, n_n207);
	defparam lut_5217.LUT_SIZE = 5;
	defparam lut_5217.mask = 32'h0f0f0100;

	lut_sub lut_5219 ({sk[1183], i_13_, i_12_}, n_n278);
	defparam lut_5219.LUT_SIZE = 3;
	defparam lut_5219.mask = 8'h52;

	lut_sub lut_5221 ({sk[1184], i_9_, i_10_, i_12_, i_11_}, n_n149);
	defparam lut_5221.LUT_SIZE = 5;
	defparam lut_5221.mask = 32'h0f0f0200;

	lut_sub lut_5223 ({sk[1185], i_14_, i_13_, i_12_, x902x}, n_n30);
	defparam lut_5223.LUT_SIZE = 5;
	defparam lut_5223.mask = 32'h0f0f0040;

	lut_sub lut_5225 ({sk[1186], i_14_, i_13_, i_12_, x899x}, n_n144);
	defparam lut_5225.LUT_SIZE = 5;
	defparam lut_5225.mask = 32'h0f0f0400;

	lut_sub lut_5227 ({sk[1187], i_14_, i_13_, i_12_, x901x}, n_n34);
	defparam lut_5227.LUT_SIZE = 5;
	defparam lut_5227.mask = 32'h0f0f1000;

	lut_sub lut_5229 ({sk[1188], i_14_, i_13_, i_12_, x897x}, n_n171);
	defparam lut_5229.LUT_SIZE = 5;
	defparam lut_5229.mask = 32'h0f0f0040;

	lut_sub lut_5231 ({sk[1189], i_14_, i_13_, i_12_, x905x}, n_n21);
	defparam lut_5231.LUT_SIZE = 5;
	defparam lut_5231.mask = 32'h0f0f0001;

	lut_sub lut_5233 ({sk[1190], i_14_, i_13_, i_12_, x911x}, n_n17);
	defparam lut_5233.LUT_SIZE = 5;
	defparam lut_5233.mask = 32'h0f0f1000;

	lut_sub lut_5235 ({sk[1191], i_14_, i_13_, i_12_, x903x}, n_n236);
	defparam lut_5235.LUT_SIZE = 5;
	defparam lut_5235.mask = 32'h0f0f0010;

	lut_sub lut_5237 ({sk[1192], i_14_, i_13_, i_12_, x904x}, n_n102);
	defparam lut_5237.LUT_SIZE = 5;
	defparam lut_5237.mask = 32'h0f0f0040;

	lut_sub lut_5239 ({sk[1193], i_14_, i_13_, i_12_, x903x}, n_n200);
	defparam lut_5239.LUT_SIZE = 5;
	defparam lut_5239.mask = 32'h0f0f0040;

	lut_sub lut_5241 ({sk[1194], i_14_, i_13_, i_12_, x905x}, n_n70);
	defparam lut_5241.LUT_SIZE = 5;
	defparam lut_5241.mask = 32'h0f0f1000;

	lut_sub lut_5243 ({sk[1195], i_7_, i_8_, i_6_, x915x, n_n256, x897x}, n_n6814);
	defparam lut_5243.LUT_SIZE = 7;
	defparam lut_5243.mask = 128'h5555ffff5555ffff0000000001000000;

	lut_sub lut_5245 ({sk[1196], i_14_, i_13_, i_12_, n_n273, x922x, x902x}, n_n6856);
	defparam lut_5245.LUT_SIZE = 7;
	defparam lut_5245.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_5247 ({sk[1197], i_7_, i_8_, i_6_, x922x, x899x, n_n256}, n_n6867);
	defparam lut_5247.LUT_SIZE = 7;
	defparam lut_5247.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_5249 ({sk[1198], i_7_, i_8_, i_6_, x922x, n_n228, x902x}, n_n6878);
	defparam lut_5249.LUT_SIZE = 7;
	defparam lut_5249.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_5251 ({sk[1199], i_14_, i_13_, i_12_, x904x}, n_n52);
	defparam lut_5251.LUT_SIZE = 5;
	defparam lut_5251.mask = 32'h0f0f0004;

	lut_sub lut_5253 ({sk[1200], i_14_, i_13_, i_12_, x899x}, n_n71);
	defparam lut_5253.LUT_SIZE = 5;
	defparam lut_5253.mask = 32'h0f0f0100;

	lut_sub lut_5255 ({sk[1201], i_14_, i_13_, i_12_, x902x}, n_n8);
	defparam lut_5255.LUT_SIZE = 5;
	defparam lut_5255.mask = 32'h0f0f0400;

	lut_sub lut_5257 ({sk[1202], i_14_, i_13_, i_12_, x904x}, n_n98);
	defparam lut_5257.LUT_SIZE = 5;
	defparam lut_5257.mask = 32'h0f0f0001;

	lut_sub lut_5259 ({sk[1203], i_7_, i_8_, i_6_}, x19206x);
	defparam lut_5259.LUT_SIZE = 4;
	defparam lut_5259.mask = 16'h552a;

	lut_sub lut_5262 ({sk[1204], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x5918x);
	defparam lut_5262.LUT_SIZE = 7;
	defparam lut_5262.mask = 128'h5555ffff5555ffff0888000000000000;

	lut_sub lut_5265 ({sk[1205], i_9_, i_10_, i_12_, i_11_}, x19205x);
	defparam lut_5265.LUT_SIZE = 5;
	defparam lut_5265.mask = 32'h0f0f7fff;

	lut_sub lut_5270 ({sk[1206], n_n281, n_n283, x901x, x19206x, x5918x, x19205x}, x1011x);
	defparam lut_5270.LUT_SIZE = 7;
	defparam lut_5270.mask = 128'h5555ffff5555ffff0f0f7f7f0f0f7fff;

	lut_sub lut_5275 ({sk[1207], i_9_, i_10_, i_11_, i_15_, n_n281, n_n279}, x284x);
	defparam lut_5275.LUT_SIZE = 7;
	defparam lut_5275.mask = 128'h5555ffff5555ffff0000000000ff3500;

	lut_sub lut_5279 ({sk[1208], i_9_, i_10_, i_11_, i_15_, n_n281, n_n279}, x282x);
	defparam lut_5279.LUT_SIZE = 7;
	defparam lut_5279.mask = 128'h5555ffff5555ffff000000ff35000000;

	lut_sub lut_5283 ({sk[1209], i_14_, i_13_, i_12_, i_15_, n_n247, x282x}, x19316x);
	defparam lut_5283.LUT_SIZE = 7;
	defparam lut_5283.mask = 128'h5555ffff5555ffff5577577755777777;

	lut_sub lut_5288 ({sk[1210], i_7_, i_8_, i_6_, x921x, x284x, x19316x}, n_n5030);
	defparam lut_5288.LUT_SIZE = 7;
	defparam lut_5288.mask = 128'h5555ffff5555ffff0007000000000000;

	lut_sub lut_5291 ({sk[1211], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19208x);
	defparam lut_5291.LUT_SIZE = 7;
	defparam lut_5291.mask = 128'h5555ffff5555ffff000000000000ffcf;

	lut_sub lut_5298 ({sk[1212], x915x, n_n271, x905x, n_n258, x904x, x19208x}, x5909x);
	defparam lut_5298.LUT_SIZE = 7;
	defparam lut_5298.mask = 128'h5555ffff5555ffff000000000000575f;

	lut_sub lut_5302 ({sk[1213], i_14_, i_13_, i_12_, x898x}, x254x);
	defparam lut_5302.LUT_SIZE = 5;
	defparam lut_5302.mask = 32'h0f0f0054;

	lut_sub lut_5306 ({sk[1214], i_14_, i_13_, i_12_, x902x}, x165x);
	defparam lut_5306.LUT_SIZE = 5;
	defparam lut_5306.mask = 32'h0f0f5100;

	lut_sub lut_5310 ({sk[1215], i_7_, i_8_, i_6_, n_n220, x909x, x908x}, x5386x);
	defparam lut_5310.LUT_SIZE = 7;
	defparam lut_5310.mask = 128'h5555ffff5555ffff0000000001000000;

	lut_sub lut_5312 ({sk[1216], i_14_, i_13_, i_12_, x903x, x897x}, x1920x);
	defparam lut_5312.LUT_SIZE = 6;
	defparam lut_5312.mask = 64'h3f3f3f3f57073000;

	lut_sub lut_5319 ({sk[1217], i_7_, i_8_, i_6_, x909x, x180x}, n_n4960);
	defparam lut_5319.LUT_SIZE = 6;
	defparam lut_5319.mask = 64'h3f3f3f3f00000001;

	lut_sub lut_5321 ({sk[1218], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x87x);
	defparam lut_5321.LUT_SIZE = 7;
	defparam lut_5321.mask = 128'h5555ffff5555ffff1010000000000000;

	lut_sub lut_5324 ({sk[1219], n_n266, x909x, x912x, n_n225, x87x}, n_n4952);
	defparam lut_5324.LUT_SIZE = 6;
	defparam lut_5324.mask = 64'h3f3f3f3f00000057;

	lut_sub lut_5327 ({sk[1220], i_14_, i_13_, i_12_, i_15_, x912x, n_n137}, x219x);
	defparam lut_5327.LUT_SIZE = 7;
	defparam lut_5327.mask = 128'h5555ffff5555ffff0505050537370505;

	lut_sub lut_5331 ({sk[1221], i_14_, i_13_, i_12_, n_n271, x909x, x904x}, x497x);
	defparam lut_5331.LUT_SIZE = 7;
	defparam lut_5331.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_5334 ({sk[1222], i_14_, i_13_, i_12_, n_n271, x909x, x904x}, n_n4955);
	defparam lut_5334.LUT_SIZE = 7;
	defparam lut_5334.mask = 128'h5555ffff5555ffff0001010100000000;

	lut_sub lut_5338 ({sk[1223], i_7_, i_8_, i_6_, x909x, x99x}, n_n4956);
	defparam lut_5338.LUT_SIZE = 6;
	defparam lut_5338.mask = 64'h3f3f3f3f00000100;

	lut_sub lut_5340 ({sk[1224], i_7_, i_8_, i_6_, x909x, x41x}, x5288x);
	defparam lut_5340.LUT_SIZE = 6;
	defparam lut_5340.mask = 64'h3f3f3f3f00000100;

	lut_sub lut_5342 ({sk[1225], n_n57, x219x, x189x, n_n4955, n_n4956, x5288x}, x20710x);
	defparam lut_5342.LUT_SIZE = 7;
	defparam lut_5342.mask = 128'h5555ffff5555ffff7f7f7f7f7fffffff;

	lut_sub lut_5348 ({sk[1226], i_7_, i_6_, i_4_, n_n6582, x259x}, x19862x);
	defparam lut_5348.LUT_SIZE = 6;
	defparam lut_5348.mask = 64'h3f3f3f3f37333333;

	lut_sub lut_5351 ({sk[1227], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1894x);
	defparam lut_5351.LUT_SIZE = 7;
	defparam lut_5351.mask = 128'h5555ffff5555ffff0010001050004040;

	lut_sub lut_5358 ({sk[1228], i_14_, i_13_, i_12_, n_n273, x922x, x899x}, n_n6875);
	defparam lut_5358.LUT_SIZE = 7;
	defparam lut_5358.mask = 128'h5555ffff5555ffff0000000000000001;

	lut_sub lut_5360 ({sk[1229], i_7_, i_8_, i_6_, x916x, n_n258, x908x}, n_n7425);
	defparam lut_5360.LUT_SIZE = 7;
	defparam lut_5360.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_5362 ({sk[1230], i_7_, i_8_, i_6_, n_n222, x922x, x899x}, n_n6861);
	defparam lut_5362.LUT_SIZE = 7;
	defparam lut_5362.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_5364 ({sk[1231], n_n273, x905x, n_n279, x922x, x899x, n_n228}, x4598x);
	defparam lut_5364.LUT_SIZE = 7;
	defparam lut_5364.mask = 128'h5555ffff5555ffff0000000000030507;

	lut_sub lut_5367 ({sk[1232], n_n273, n_n222, x922x, x899x, x4598x}, n_n4073);
	defparam lut_5367.LUT_SIZE = 6;
	defparam lut_5367.mask = 64'h3f3f3f3f55555557;

	lut_sub lut_5370 ({sk[1233], i_14_, i_13_, i_12_, n_n273, x922x, x899x}, n_n6876);
	defparam lut_5370.LUT_SIZE = 7;
	defparam lut_5370.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_5372 ({sk[1234], n_n281, n_n273, n_n220, x905x, x922x, x899x}, x475x);
	defparam lut_5372.LUT_SIZE = 7;
	defparam lut_5372.mask = 128'h5555ffff5555ffff0000001100000313;

	lut_sub lut_5375 ({sk[1235], i_7_, i_8_, i_6_, n_n281, x922x, x908x}, x438x);
	defparam lut_5375.LUT_SIZE = 7;
	defparam lut_5375.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_5377 ({sk[1236], n_n273, n_n220, x922x, x899x, n_n228, x902x}, x20386x);
	defparam lut_5377.LUT_SIZE = 7;
	defparam lut_5377.mask = 128'h5555ffff5555ffff0000000000030057;

	lut_sub lut_5380 ({sk[1237], i_14_, i_13_, i_12_, x904x}, n_n49);
	defparam lut_5380.LUT_SIZE = 5;
	defparam lut_5380.mask = 32'h0f0f1000;

	lut_sub lut_5382 ({sk[1238], i_14_, i_13_, i_12_, n_n3, x900x}, x3635x);
	defparam lut_5382.LUT_SIZE = 6;
	defparam lut_5382.mask = 64'h3f3f3f3f00000100;

	lut_sub lut_5384 ({sk[1239], i_14_, i_13_, i_12_, x915x, n_n263, x908x}, x3776x);
	defparam lut_5384.LUT_SIZE = 7;
	defparam lut_5384.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_5387 ({sk[1240], i_7_, i_8_, i_6_, n_n220, x909x, x908x}, x562x);
	defparam lut_5387.LUT_SIZE = 7;
	defparam lut_5387.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5389 ({sk[1241], i_7_, i_8_, i_6_, x909x, x82x}, x4998x);
	defparam lut_5389.LUT_SIZE = 6;
	defparam lut_5389.mask = 64'h3f3f3f3f00000001;

	lut_sub lut_5391 ({sk[1242], i_7_, i_8_, i_6_, x909x, x207x}, n_n4924);
	defparam lut_5391.LUT_SIZE = 6;
	defparam lut_5391.mask = 64'h3f3f3f3f00000100;

	lut_sub lut_5393 ({sk[1243], i_7_, i_8_, i_6_, x909x, x163x, x207x}, x555x);
	defparam lut_5393.LUT_SIZE = 7;
	defparam lut_5393.mask = 128'h5555ffff5555ffff0000000000070000;

	lut_sub lut_5396 ({sk[1244], i_7_, i_8_, i_6_, x909x, x125x, x111x}, x682x);
	defparam lut_5396.LUT_SIZE = 7;
	defparam lut_5396.mask = 128'h5555ffff5555ffff0000000000000007;

	lut_sub lut_5399 ({sk[1245], n_n57, n_n56, n_n76, x82x, x163x, x207x}, x21075x);
	defparam lut_5399.LUT_SIZE = 7;
	defparam lut_5399.mask = 128'h5555ffff5555ffff000077ff7fff7fff;

	lut_sub lut_5407 ({sk[1246], i_14_, i_13_, i_12_, x915x, x914x, n_n263}, x500x);
	defparam lut_5407.LUT_SIZE = 7;
	defparam lut_5407.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5409 ({sk[1247], i_7_, i_8_, i_6_, x915x, x912x, n_n256}, n_n6835);
	defparam lut_5409.LUT_SIZE = 7;
	defparam lut_5409.mask = 128'h5555ffff5555ffff0000000001000000;

	lut_sub lut_5411 ({sk[1248], i_14_, i_13_, i_12_, x915x, n_n263, x912x}, x686x);
	defparam lut_5411.LUT_SIZE = 7;
	defparam lut_5411.mask = 128'h5555ffff5555ffff0001000100000000;

	lut_sub lut_5414 ({sk[1249], i_15_, x915x, x914x, n_n263, n_n228, n_n137}, x825x);
	defparam lut_5414.LUT_SIZE = 7;
	defparam lut_5414.mask = 128'h5555ffff5555ffff0000050700000003;

	lut_sub lut_5417 ({sk[1250], n_n88, n_n228, x912x, n_n94, x500x, x686x}, x24120x);
	defparam lut_5417.LUT_SIZE = 7;
	defparam lut_5417.mask = 128'h5555ffff5555ffff8888888080808080;

	lut_sub lut_5421 ({sk[1251], n_n208, x916x, n_n31, n_n6847, x825x, x24120x}, n_n3167);
	defparam lut_5421.LUT_SIZE = 7;
	defparam lut_5421.mask = 128'h5555ffff5555ffffbfbfbfbfbfbfbfff;

	lut_sub lut_5426 ({sk[1252], i_14_, i_13_, i_12_, x915x, n_n263, x912x}, n_n6830);
	defparam lut_5426.LUT_SIZE = 7;
	defparam lut_5426.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5428 ({sk[1253], i_7_, i_8_, i_6_, x909x}, x278x);
	defparam lut_5428.LUT_SIZE = 5;
	defparam lut_5428.mask = 32'h0f0f1100;

	lut_sub lut_5431 ({sk[1254], i_14_, i_13_, i_12_, x902x, n_n227}, x655x);
	defparam lut_5431.LUT_SIZE = 6;
	defparam lut_5431.mask = 64'h3f3f3f3f00010000;

	lut_sub lut_5433 ({sk[1255], i_7_, i_8_, i_6_, x909x, x905x, n_n256}, x685x);
	defparam lut_5433.LUT_SIZE = 7;
	defparam lut_5433.mask = 128'h5555ffff5555ffff0001000000000000;

	lut_sub lut_5435 ({sk[1256], i_14_, i_13_, i_12_, i_15_, n_n259, n_n270}, x1019x);
	defparam lut_5435.LUT_SIZE = 7;
	defparam lut_5435.mask = 128'h5555ffff5555ffff0003005035073570;

	lut_sub lut_5446 ({sk[1257], i_7_, i_8_, i_6_, x909x, x1019x}, x3870x);
	defparam lut_5446.LUT_SIZE = 6;
	defparam lut_5446.mask = 64'h3f3f3f3f01000000;

	lut_sub lut_5448 ({sk[1258], i_14_, i_13_, i_12_, n_n3, x904x}, x19389x);
	defparam lut_5448.LUT_SIZE = 6;
	defparam lut_5448.mask = 64'h3f3f3f3f01100000;

	lut_sub lut_5451 ({sk[1259], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x71x);
	defparam lut_5451.LUT_SIZE = 7;
	defparam lut_5451.mask = 128'h5555ffff5555ffff0100000400000000;

	lut_sub lut_5454 ({sk[1260], i_14_, i_13_, i_12_, n_n3, x904x, x71x}, x557x);
	defparam lut_5454.LUT_SIZE = 7;
	defparam lut_5454.mask = 128'h5555ffff5555ffff0507070505050505;

	lut_sub lut_5458 ({sk[1261], i_14_, i_13_, i_12_, i_15_, n_n247, x55x}, x1022x);
	defparam lut_5458.LUT_SIZE = 7;
	defparam lut_5458.mask = 128'h5555ffff5555ffff5775557557557575;

	lut_sub lut_5466 ({sk[1262], i_14_, i_13_, i_12_, i_15_, n_n247, x55x}, x1021x);
	defparam lut_5466.LUT_SIZE = 7;
	defparam lut_5466.mask = 128'h5555ffff5555ffff5775757557557575;

	lut_sub lut_5475 ({sk[1263], n_n4, n_n3, x93x, x19389x, x1022x, x71x}, x21140x);
	defparam lut_5475.LUT_SIZE = 7;
	defparam lut_5475.mask = 128'h5555ffff5555ffff0f0f7fff0fff7fff;

	lut_sub lut_5481 ({sk[1264], i_14_, i_13_, i_12_, i_15_, x908x, n_n270}, x209x);
	defparam lut_5481.LUT_SIZE = 7;
	defparam lut_5481.mask = 128'h5555ffff5555ffff3300050000330000;

	lut_sub lut_5485 ({sk[1265], i_7_, i_8_, i_6_, x915x, x899x, n_n228}, x739x);
	defparam lut_5485.LUT_SIZE = 7;
	defparam lut_5485.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_5487 ({sk[1266], i_14_, i_13_, i_12_, i_15_, x159x, n_n247}, x20928x);
	defparam lut_5487.LUT_SIZE = 7;
	defparam lut_5487.mask = 128'h5555ffff5555ffff7333373333333333;

	lut_sub lut_5491 ({sk[1267], i_14_, i_13_, i_12_, x905x, x899x, x902x}, x1023x);
	defparam lut_5491.LUT_SIZE = 7;
	defparam lut_5491.mask = 128'h5555ffff5555ffff0f00330000000055;

	lut_sub lut_5495 ({sk[1268], i_14_, i_13_, i_12_, i_15_, n_n247, x189x}, x1326x);
	defparam lut_5495.LUT_SIZE = 7;
	defparam lut_5495.mask = 128'h5555ffff5555ffff5555555557575755;

	lut_sub lut_5500 ({sk[1269], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1283x);
	defparam lut_5500.LUT_SIZE = 7;
	defparam lut_5500.mask = 128'h5555ffff5555ffff0105000505000404;

	lut_sub lut_5510 ({sk[1270], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x1025x);
	defparam lut_5510.LUT_SIZE = 7;
	defparam lut_5510.mask = 128'h5555ffff5555ffff0040504000400010;

	lut_sub lut_5517 ({sk[1271], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1932x);
	defparam lut_5517.LUT_SIZE = 7;
	defparam lut_5517.mask = 128'h5555ffff5555ffff0010001050004040;

	lut_sub lut_5524 ({sk[1272], i_7_, i_8_, i_6_, x915x, n_n220, x905x}, x5204x);
	defparam lut_5524.LUT_SIZE = 7;
	defparam lut_5524.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_5526 ({sk[1273], i_7_, i_8_, i_6_, x915x, x258x}, n_n3520);
	defparam lut_5526.LUT_SIZE = 6;
	defparam lut_5526.mask = 64'h3f3f3f3f10000000;

	lut_sub lut_5528 ({sk[1274], i_14_, i_13_, i_12_, x907x}, n_n81);
	defparam lut_5528.LUT_SIZE = 5;
	defparam lut_5528.mask = 32'h0f0f1000;

	lut_sub lut_5530 ({sk[1275], i_7_, i_8_, i_6_, x907x, x915x, n_n256}, n_n6829);
	defparam lut_5530.LUT_SIZE = 7;
	defparam lut_5530.mask = 128'h5555ffff5555ffff0000000000000100;

	lut_sub lut_5532 ({sk[1276], n_n281, x907x, n_n273, x922x, x901x, n_n225}, x470x);
	defparam lut_5532.LUT_SIZE = 7;
	defparam lut_5532.mask = 128'h5555ffff5555ffff0000000500030007;

	lut_sub lut_5535 ({sk[1277], i_9_, i_10_, i_11_, i_15_, x79x, n_n256}, x188x);
	defparam lut_5535.LUT_SIZE = 7;
	defparam lut_5535.mask = 128'h5555ffff5555ffff3333333333333733;

	lut_sub lut_5538 ({sk[1278], i_7_, i_8_, i_6_, x916x, x188x}, n_n2986);
	defparam lut_5538.LUT_SIZE = 6;
	defparam lut_5538.mask = 64'h3f3f3f3f00010000;

	lut_sub lut_5540 ({sk[1279], i_14_, i_13_, i_12_, n_n273, x914x, x922x}, x561x);
	defparam lut_5540.LUT_SIZE = 7;
	defparam lut_5540.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_5542 ({sk[1280], n_n281, x914x, n_n48, n_n53, x908x, x903x}, x21564x);
	defparam lut_5542.LUT_SIZE = 7;
	defparam lut_5542.mask = 128'h5555ffff5555ffff0000000005770fff;

	lut_sub lut_5548 ({sk[1281], i_14_, i_13_, i_12_, n_n273, x905x, x922x}, n_n2272);
	defparam lut_5548.LUT_SIZE = 7;
	defparam lut_5548.mask = 128'h5555ffff5555ffff0001010100000000;

	lut_sub lut_5552 ({sk[1282], i_14_, i_13_, i_12_, x907x, x901x}, x267x);
	defparam lut_5552.LUT_SIZE = 6;
	defparam lut_5552.mask = 64'h3f3f3f3f50033000;

	lut_sub lut_5556 ({sk[1283], i_14_, i_13_, i_12_, x907x, x901x}, x1029x);
	defparam lut_5556.LUT_SIZE = 6;
	defparam lut_5556.mask = 64'h3f3f3f3f50037000;

	lut_sub lut_5561 ({sk[1284], i_9_, i_10_, i_11_, i_15_, n_n279}, x264x);
	defparam lut_5561.LUT_SIZE = 6;
	defparam lut_5561.mask = 64'h3f3f3f3f05000000;

	lut_sub lut_5564 ({sk[1285], n_n151, n_n1, n_n2, n_n7, n_n145, n_n60}, x24104x);
	defparam lut_5564.LUT_SIZE = 7;
	defparam lut_5564.mask = 128'h5555ffff5555ffffff80f080ff000000;

	lut_sub lut_5568 ({sk[1286], i_14_, i_13_, i_12_, x908x}, n_n101);
	defparam lut_5568.LUT_SIZE = 5;
	defparam lut_5568.mask = 32'h0f0f0040;

	lut_sub lut_5570 ({sk[1287], i_14_, i_13_, i_12_, i_15_, x908x, n_n270}, x296x);
	defparam lut_5570.LUT_SIZE = 7;
	defparam lut_5570.mask = 128'h5555ffff5555ffff0500005033000000;

	lut_sub lut_5574 ({sk[1288], i_14_, i_13_, i_12_, n_n208, x916x, x908x}, x466x);
	defparam lut_5574.LUT_SIZE = 7;
	defparam lut_5574.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_5577 ({sk[1289], n_n4, n_n3, x67x, n_n30, n_n171, x296x}, x24158x);
	defparam lut_5577.LUT_SIZE = 7;
	defparam lut_5577.mask = 128'h5555ffff5555ffffffffcc00a0a08000;

	lut_sub lut_5582 ({sk[1290], n_n57, n_n56, n_n76, x264x, x207x, x46x}, n_n2166);
	defparam lut_5582.LUT_SIZE = 7;
	defparam lut_5582.mask = 128'h5555ffff5555ffff00005f5f33ff7fff;

	lut_sub lut_5587 ({sk[1291], i_14_, i_13_, i_12_, x909x, x905x, n_n261}, x411x);
	defparam lut_5587.LUT_SIZE = 7;
	defparam lut_5587.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_5590 ({sk[1292], i_14_, i_13_, i_12_, x913x, x911x}, x1034x);
	defparam lut_5590.LUT_SIZE = 6;
	defparam lut_5590.mask = 64'h3f3f3f3f50037000;

	lut_sub lut_5595 ({sk[1293], i_14_, i_13_, i_12_, i_15_, x907x, n_n282}, x1037x);
	defparam lut_5595.LUT_SIZE = 7;
	defparam lut_5595.mask = 128'h5555ffff5555ffff0533335055000000;

	lut_sub lut_5602 ({sk[1294], n_n281, x913x, n_n268, n_n111, x106x, x903x}, x3526x);
	defparam lut_5602.LUT_SIZE = 7;
	defparam lut_5602.mask = 128'h5555ffff5555ffff003f003f007f00ff;

	lut_sub lut_5607 ({sk[1295], i_14_, i_13_, i_12_, x913x, x916x, n_n271}, x765x);
	defparam lut_5607.LUT_SIZE = 7;
	defparam lut_5607.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_5609 ({sk[1296], i_7_, i_8_, i_6_, x907x, x916x, n_n220}, x779x);
	defparam lut_5609.LUT_SIZE = 7;
	defparam lut_5609.mask = 128'h5555ffff5555ffff0000000000000001;

	lut_sub lut_5611 ({sk[1297], i_7_, i_8_, i_6_, x916x, n_n220, x903x}, x934x);
	defparam lut_5611.LUT_SIZE = 7;
	defparam lut_5611.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5613 ({sk[1298], i_14_, i_13_, i_12_, x907x, x901x}, x205x);
	defparam lut_5613.LUT_SIZE = 6;
	defparam lut_5613.mask = 64'h3f3f3f3f53030000;

	lut_sub lut_5617 ({sk[1299], i_14_, i_13_, i_12_, x900x, x906x}, x149x);
	defparam lut_5617.LUT_SIZE = 6;
	defparam lut_5617.mask = 64'h3f3f3f3f30055000;

	lut_sub lut_5621 ({sk[1300], n_n208, x916x, n_n3, n_n186, x51x, x149x}, x467x);
	defparam lut_5621.LUT_SIZE = 7;
	defparam lut_5621.mask = 128'h5555ffff5555ffff000f000f000f777f;

	lut_sub lut_5625 ({sk[1301], i_14_, i_13_, i_12_, i_15_, n_n247, n_n253}, x1041x);
	defparam lut_5625.LUT_SIZE = 7;
	defparam lut_5625.mask = 128'h5555ffff5555ffff0750507073000000;

	lut_sub lut_5635 ({sk[1302], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x279x);
	defparam lut_5635.LUT_SIZE = 7;
	defparam lut_5635.mask = 128'h5555ffff5555ffff0001000100000400;

	lut_sub lut_5639 ({sk[1303], i_14_, i_13_, i_12_, x903x, x897x}, x228x);
	defparam lut_5639.LUT_SIZE = 6;
	defparam lut_5639.mask = 64'h3f3f3f3f50300000;

	lut_sub lut_5642 ({sk[1304], i_14_, i_13_, i_12_, i_15_, n_n275, x228x}, x1042x);
	defparam lut_5642.LUT_SIZE = 7;
	defparam lut_5642.mask = 128'h5555ffff5555ffff5557555755557755;

	lut_sub lut_5648 ({sk[1305], n_n48, n_n53, n_n76, n_n25, n_n6856, x1042x}, n_n1779);
	defparam lut_5648.LUT_SIZE = 7;
	defparam lut_5648.mask = 128'h5555ffff5555ffff33333fff77777fff;

	lut_sub lut_5653 ({sk[1306], i_14_, i_13_, i_12_, x897x}, n_n58);
	defparam lut_5653.LUT_SIZE = 5;
	defparam lut_5653.mask = 32'h0f0f0400;

	lut_sub lut_5655 ({sk[1307], i_7_, i_8_, i_6_, i_15_, x915x, n_n138}, n_n6818);
	defparam lut_5655.LUT_SIZE = 7;
	defparam lut_5655.mask = 128'h5555ffff5555ffff0000000001000000;

	lut_sub lut_5657 ({sk[1308], i_14_, i_13_, i_12_, x913x, x915x, n_n263}, n_n6823);
	defparam lut_5657.LUT_SIZE = 7;
	defparam lut_5657.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_5659 ({sk[1309], i_7_, i_8_, i_6_, x915x, x911x, n_n225}, n_n6820);
	defparam lut_5659.LUT_SIZE = 7;
	defparam lut_5659.mask = 128'h5555ffff5555ffff0000000001000000;

	lut_sub lut_5661 ({sk[1310], i_14_, i_13_, i_12_, x915x, x911x, n_n263}, x696x);
	defparam lut_5661.LUT_SIZE = 7;
	defparam lut_5661.mask = 128'h5555ffff5555ffff0100000100000000;

	lut_sub lut_5664 ({sk[1311], x913x, n_n220, n_n94, x897x, x686x, n_n6818}, x21689x);
	defparam lut_5664.LUT_SIZE = 7;
	defparam lut_5664.mask = 128'h5555ffff5555ffff7777777f777777ff;

	lut_sub lut_5669 ({sk[1312], i_15_, x915x, n_n263, n_n137, x696x, x21689x}, n_n1757);
	defparam lut_5669.LUT_SIZE = 7;
	defparam lut_5669.mask = 128'h5555ffff5555ffff7777777f7777777f;

	lut_sub lut_5674 ({sk[1313], i_14_, i_13_, i_12_, n_n208, x909x, x905x}, x480x);
	defparam lut_5674.LUT_SIZE = 7;
	defparam lut_5674.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5676 ({sk[1314], i_7_, i_8_, i_6_, x913x, x909x, n_n256}, x700x);
	defparam lut_5676.LUT_SIZE = 7;
	defparam lut_5676.mask = 128'h5555ffff5555ffff0000000100000000;

	lut_sub lut_5678 ({sk[1315], i_14_, i_13_, i_12_, i_15_, x913x, n_n259}, x1043x);
	defparam lut_5678.LUT_SIZE = 7;
	defparam lut_5678.mask = 128'h5555ffff5555ffff0005000050375050;

	lut_sub lut_5685 ({sk[1316], n_n227, x685x, x480x, x700x, x1043x}, n_n1215);
	defparam lut_5685.LUT_SIZE = 6;
	defparam lut_5685.mask = 64'h3f3f3f3f3fff7fff;

	lut_sub lut_5690 ({sk[1317], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x142x);
	defparam lut_5690.LUT_SIZE = 7;
	defparam lut_5690.mask = 128'h5555ffff5555ffff0000000040004040;

	lut_sub lut_5694 ({sk[1318], i_14_, i_13_, i_12_, x915x, n_n263, x899x}, x566x);
	defparam lut_5694.LUT_SIZE = 7;
	defparam lut_5694.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5696 ({sk[1319], i_14_, i_13_, i_12_, i_15_, n_n242, n_n259}, x1045x);
	defparam lut_5696.LUT_SIZE = 7;
	defparam lut_5696.mask = 128'h5555ffff5555ffff0033000000035570;

	lut_sub lut_5704 ({sk[1320], i_14_, i_13_, i_12_, i_15_, x905x, n_n259}, x355x);
	defparam lut_5704.LUT_SIZE = 7;
	defparam lut_5704.mask = 128'h5555ffff5555ffff0533500000000000;

	lut_sub lut_5708 ({sk[1321], i_14_, i_13_, i_12_, i_15_, n_n242, x355x}, x1044x);
	defparam lut_5708.LUT_SIZE = 7;
	defparam lut_5708.mask = 128'h5555ffff5555ffff5757555755575755;

	lut_sub lut_5715 ({sk[1322], i_14_, i_13_, i_12_, i_15_, n_n242, n_n138}, x514x);
	defparam lut_5715.LUT_SIZE = 7;
	defparam lut_5715.mask = 128'h5555ffff5555ffff5050505070505050;

	lut_sub lut_5718 ({sk[1323], n_n100, n_n94, n_n6820, x142x, x1045x, x514x}, x22184x);
	defparam lut_5718.LUT_SIZE = 7;
	defparam lut_5718.mask = 128'h5555ffff5555ffff00ff77ff0fff7fff;

	lut_sub lut_5723 ({sk[1324], i_15_, n_n281, x911x, n_n94, n_n138, n_n6823}, x24182x);
	defparam lut_5723.LUT_SIZE = 7;
	defparam lut_5723.mask = 128'h5555ffff5555ffffaaaaaaa0a8a8a8a0;

	lut_sub lut_5729 ({sk[1325], x915x, n_n261, x62x, x566x, x1044x, x24182x}, x22185x);
	defparam lut_5729.LUT_SIZE = 7;
	defparam lut_5729.mask = 128'h5555ffff5555ffffafafafafafafbfff;

	lut_sub lut_5734 ({sk[1326], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1046x);
	defparam lut_5734.LUT_SIZE = 7;
	defparam lut_5734.mask = 128'h5555ffff5555ffff0105000104010504;

	lut_sub lut_5744 ({sk[1327], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x223x);
	defparam lut_5744.LUT_SIZE = 7;
	defparam lut_5744.mask = 128'h5555ffff5555ffff0000100000400000;

	lut_sub lut_5747 ({sk[1328], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1048x);
	defparam lut_5747.LUT_SIZE = 7;
	defparam lut_5747.mask = 128'h5555ffff5555ffff0053000000005300;

	lut_sub lut_5752 ({sk[1329], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1047x);
	defparam lut_5752.LUT_SIZE = 7;
	defparam lut_5752.mask = 128'h5555ffff5555ffff0053500000530000;

	lut_sub lut_5758 ({sk[1330], i_14_, i_13_, i_12_, x913x, x911x}, x75x);
	defparam lut_5758.LUT_SIZE = 6;
	defparam lut_5758.mask = 64'h3f3f3f3f00500300;

	lut_sub lut_5761 ({sk[1331], i_9_, i_10_, i_11_, n_n261, x922x}, x579x);
	defparam lut_5761.LUT_SIZE = 6;
	defparam lut_5761.mask = 64'h3f3f3f3f00100000;

	lut_sub lut_5763 ({sk[1332], i_9_, i_10_, i_11_, n_n263, x922x}, x764x);
	defparam lut_5763.LUT_SIZE = 6;
	defparam lut_5763.mask = 64'h3f3f3f3f00000010;

	lut_sub lut_5765 ({sk[1333], i_14_, i_13_, i_12_, i_15_, x911x, n_n259}, x1049x);
	defparam lut_5765.LUT_SIZE = 7;
	defparam lut_5765.mask = 128'h5555ffff5555ffff0000370000500000;

	lut_sub lut_5769 ({sk[1334], n_n57, n_n261, x922x, n_n282, x457x, x75x}, x24091x);
	defparam lut_5769.LUT_SIZE = 7;
	defparam lut_5769.mask = 128'h5555ffff5555ffffccccccc088888880;

	lut_sub lut_5776 ({sk[1335], n_n271, x909x, x579x, x764x, x1049x, x24091x}, x22264x);
	defparam lut_5776.LUT_SIZE = 7;
	defparam lut_5776.mask = 128'h5555ffff5555ffffafffafffafffbfff;

	lut_sub lut_5781 ({sk[1336], n_n57, n_n56, n_n53, x1046x, x1048x, x1047x}, x22265x);
	defparam lut_5781.LUT_SIZE = 7;
	defparam lut_5781.mask = 128'h5555ffff5555ffff000f555f333f777f;

	lut_sub lut_5785 ({sk[1337], i_14_, i_13_, i_12_, i_15_, x902x, n_n242}, x1051x);
	defparam lut_5785.LUT_SIZE = 7;
	defparam lut_5785.mask = 128'h5555ffff5555ffff3777003750055550;

	lut_sub lut_5798 ({sk[1338], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1050x);
	defparam lut_5798.LUT_SIZE = 7;
	defparam lut_5798.mask = 128'h5555ffff5555ffff1000000000005040;

	lut_sub lut_5803 ({sk[1339], x909x, n_n261, x60x, x5260x, x411x, x1050x}, x22020x);
	defparam lut_5803.LUT_SIZE = 7;
	defparam lut_5803.mask = 128'h5555ffff5555ffff3f3f3f3f3f3f7fff;

	lut_sub lut_5808 ({sk[1340], n_n6, n_n5, n_n197, x125x, x4716x, x1051x}, x22021x);
	defparam lut_5808.LUT_SIZE = 7;
	defparam lut_5808.mask = 128'h5555ffff5555ffff333377773fff7fff;

	lut_sub lut_5813 ({sk[1341], i_14_, i_13_, i_12_, i_15_, n_n282, n_n253}, x1053x);
	defparam lut_5813.LUT_SIZE = 7;
	defparam lut_5813.mask = 128'h5555ffff5555ffff0777500770037370;

	lut_sub lut_5831 ({sk[1342], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x1052x);
	defparam lut_5831.LUT_SIZE = 7;
	defparam lut_5831.mask = 128'h5555ffff5555ffff1040400000105040;

	lut_sub lut_5839 ({sk[1343], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x123x);
	defparam lut_5839.LUT_SIZE = 7;
	defparam lut_5839.mask = 128'h5555ffff5555ffff0000000040004040;

	lut_sub lut_5843 ({sk[1344], i_14_, i_13_, i_12_, x899x}, x100x);
	defparam lut_5843.LUT_SIZE = 5;
	defparam lut_5843.mask = 32'h0f0f5100;

	lut_sub lut_5847 ({sk[1345], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x42x);
	defparam lut_5847.LUT_SIZE = 7;
	defparam lut_5847.mask = 128'h5555ffff5555ffff0000000000004040;

	lut_sub lut_5850 ({sk[1346], i_14_, i_13_, i_12_, x905x, x899x, x42x}, x1054x);
	defparam lut_5850.LUT_SIZE = 7;
	defparam lut_5850.mask = 128'h5555ffff5555ffff777755775f555555;

	lut_sub lut_5856 ({sk[1347], n_n208, x916x, n_n3, x83x, n_n252, x1054x}, n_n1159);
	defparam lut_5856.LUT_SIZE = 7;
	defparam lut_5856.mask = 128'h5555ffff5555ffff005f005f005f337f;

	lut_sub lut_5860 ({sk[1348], i_14_, i_13_, i_12_, i_15_, n_n242, n_n138}, x97x);
	defparam lut_5860.LUT_SIZE = 7;
	defparam lut_5860.mask = 128'h5555ffff5555ffff5050505370505050;

	lut_sub lut_5864 ({sk[1349], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1055x);
	defparam lut_5864.LUT_SIZE = 7;
	defparam lut_5864.mask = 128'h5555ffff5555ffff1050001040004000;

	lut_sub lut_5871 ({sk[1350], x913x, n_n220, n_n4, n_n3, x82x, x1055x}, n_n1160);
	defparam lut_5871.LUT_SIZE = 7;
	defparam lut_5871.mask = 128'h5555ffff5555ffff03570357035703ff;

	lut_sub lut_5875 ({sk[1351], i_14_, i_13_, i_12_, x907x, n_n273, x922x}, n_n6517);
	defparam lut_5875.LUT_SIZE = 7;
	defparam lut_5875.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5877 ({sk[1352], i_14_, i_13_, i_12_, x907x, n_n273, x922x}, x376x);
	defparam lut_5877.LUT_SIZE = 7;
	defparam lut_5877.mask = 128'h5555ffff5555ffff0001010000000000;

	lut_sub lut_5880 ({sk[1353], i_7_, i_8_, i_6_, x914x, x922x, n_n228}, x2687x);
	defparam lut_5880.LUT_SIZE = 7;
	defparam lut_5880.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_5882 ({sk[1354], i_7_, i_8_, i_6_, x914x, n_n258, x922x}, n_n6520);
	defparam lut_5882.LUT_SIZE = 7;
	defparam lut_5882.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_5884 ({sk[1355], i_7_, i_8_, i_6_, x922x, x912x, n_n256}, n_n6511);
	defparam lut_5884.LUT_SIZE = 7;
	defparam lut_5884.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_5886 ({sk[1356], i_14_, i_13_, i_12_, n_n283, x922x, x912x}, n_n6512);
	defparam lut_5886.LUT_SIZE = 7;
	defparam lut_5886.mask = 128'h5555ffff5555ffff0100000000000000;

	lut_sub lut_5888 ({sk[1357], i_14_, i_13_, i_12_, n_n283, x922x, x912x}, x629x);
	defparam lut_5888.LUT_SIZE = 7;
	defparam lut_5888.mask = 128'h5555ffff5555ffff0101000000000000;

	lut_sub lut_5891 ({sk[1358], i_14_, i_13_, i_12_, n_n283, x922x, x912x}, n_n6521);
	defparam lut_5891.LUT_SIZE = 7;
	defparam lut_5891.mask = 128'h5555ffff5555ffff0000010000000000;

	lut_sub lut_5893 ({sk[1359], n_n273, n_n283, n_n220, x922x, x901x, x912x}, x631x);
	defparam lut_5893.LUT_SIZE = 7;
	defparam lut_5893.mask = 128'h5555ffff5555ffff0000000500030007;

	lut_sub lut_5896 ({sk[1360], i_14_, i_13_, i_12_, n_n273, x905x, x922x}, n_n6879);
	defparam lut_5896.LUT_SIZE = 7;
	defparam lut_5896.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5898 ({sk[1361], i_8_, n_n155, n_n220, x922x, x902x, n_n6876}, x679x);
	defparam lut_5898.LUT_SIZE = 7;
	defparam lut_5898.mask = 128'h5555ffff5555ffff5555555755555555;

	lut_sub lut_5901 ({sk[1362], i_14_, i_13_, i_12_, x913x, x903x, x897x}, x1338x);
	defparam lut_5901.LUT_SIZE = 7;
	defparam lut_5901.mask = 128'h5555ffff5555ffff00005500003f0000;

	lut_sub lut_5905 ({sk[1363], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1337x);
	defparam lut_5905.LUT_SIZE = 7;
	defparam lut_5905.mask = 128'h5555ffff5555ffff0000530000500000;

	lut_sub lut_5909 ({sk[1364], i_14_, i_13_, i_12_, x903x, x897x}, x50x);
	defparam lut_5909.LUT_SIZE = 6;
	defparam lut_5909.mask = 64'h3f3f3f3f00500300;

	lut_sub lut_5912 ({sk[1365], n_n273, n_n220, n_n258, x922x, x908x, x902x}, x22134x);
	defparam lut_5912.LUT_SIZE = 7;
	defparam lut_5912.mask = 128'h5555ffff5555ffff0000000000030507;

	lut_sub lut_5915 ({sk[1366], i_8_, n_n155, n_n220, x922x, x901x, n_n6521}, x22136x);
	defparam lut_5915.LUT_SIZE = 7;
	defparam lut_5915.mask = 128'h5555ffff5555ffff5555555755555557;

	lut_sub lut_5919 ({sk[1367], i_14_, i_13_, i_12_, x914x, x115x, x912x}, x1059x);
	defparam lut_5919.LUT_SIZE = 7;
	defparam lut_5919.mask = 128'h5555ffff5555ffff3333337f33773333;

	lut_sub lut_5924 ({sk[1368], n_n208, x916x, n_n104, n_n3, x134x, x1059x}, n_n784);
	defparam lut_5924.LUT_SIZE = 7;
	defparam lut_5924.mask = 128'h5555ffff5555ffff030f030f030f575f;

	lut_sub lut_5928 ({sk[1369], i_7_, i_8_, i_6_, x915x}, x168x);
	defparam lut_5928.LUT_SIZE = 5;
	defparam lut_5928.mask = 32'h0f0f0044;

	lut_sub lut_5931 ({sk[1370], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1060x);
	defparam lut_5931.LUT_SIZE = 7;
	defparam lut_5931.mask = 128'h5555ffff5555ffff0000005010001041;

	lut_sub lut_5938 ({sk[1371], i_15_, x915x, x911x, n_n279, n_n263, n_n138}, x381x);
	defparam lut_5938.LUT_SIZE = 7;
	defparam lut_5938.mask = 128'h5555ffff5555ffff0000000300001113;

	lut_sub lut_5941 ({sk[1372], x913x, x915x, n_n263, n_n228, n_n204, n_n6818}, n_n1058);
	defparam lut_5941.LUT_SIZE = 7;
	defparam lut_5941.mask = 128'h5555ffff5555ffff555555775555557f;

	lut_sub lut_5945 ({sk[1373], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x107x);
	defparam lut_5945.LUT_SIZE = 7;
	defparam lut_5945.mask = 128'h5555ffff5555ffff0000000010001040;

	lut_sub lut_5949 ({sk[1374], i_14_, i_13_, i_12_, x915x, x911x, n_n263}, x567x);
	defparam lut_5949.LUT_SIZE = 7;
	defparam lut_5949.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5951 ({sk[1375], x913x, x915x, x911x, n_n263, n_n225}, x697x);
	defparam lut_5951.LUT_SIZE = 6;
	defparam lut_5951.mask = 64'h3f3f3f3f00010011;

	lut_sub lut_5954 ({sk[1376], i_9_, i_10_, i_11_, i_15_, n_n225}, x161x);
	defparam lut_5954.LUT_SIZE = 6;
	defparam lut_5954.mask = 64'h3f3f3f3f00500000;

	lut_sub lut_5957 ({sk[1377], n_n100, x566x, x109x, n_n1058, x107x, x567x}, x22611x);
	defparam lut_5957.LUT_SIZE = 7;
	defparam lut_5957.mask = 128'h5555ffff5555ffff5f5fffff7fffffff;

	lut_sub lut_5963 ({sk[1378], n_n216, n_n100, n_n15, x697x, x128x, x161x}, x24163x);
	defparam lut_5963.LUT_SIZE = 7;
	defparam lut_5963.mask = 128'h5555ffff5555fffff0f08000f0f00000;

	lut_sub lut_5966 ({sk[1379], x915x, n_n65, n_n261, n_n263, x1060x, x24163x}, x22612x);
	defparam lut_5966.LUT_SIZE = 7;
	defparam lut_5966.mask = 128'h5555ffff5555ffffaaaaaaaaababafff;

	lut_sub lut_5971 ({sk[1380], i_14_, i_13_, i_12_, n_n273, x922x, x901x}, x516x);
	defparam lut_5971.LUT_SIZE = 7;
	defparam lut_5971.mask = 128'h5555ffff5555ffff0000000000010100;

	lut_sub lut_5974 ({sk[1381], n_n48, n_n53, x899x, n_n228, x902x, x516x}, x22728x);
	defparam lut_5974.LUT_SIZE = 7;
	defparam lut_5974.mask = 128'h5555ffff5555ffff5555555f575f575f;

	lut_sub lut_5979 ({sk[1382], n_n48, n_n53, n_n84, n_n206, n_n59, x22728x}, n_n825);
	defparam lut_5979.LUT_SIZE = 7;
	defparam lut_5979.mask = 128'h5555ffff5555ffff55557fff5f5f7fff;

	lut_sub lut_5985 ({sk[1383], i_14_, i_13_, i_12_, n_n283, x922x, x899x}, x752x);
	defparam lut_5985.LUT_SIZE = 7;
	defparam lut_5985.mask = 128'h5555ffff5555ffff0000000000010000;

	lut_sub lut_5987 ({sk[1384], i_9_, i_10_, i_14_, i_11_, i_15_, n_n254}, x1065x);
	defparam lut_5987.LUT_SIZE = 7;
	defparam lut_5987.mask = 128'h5555ffff5555ffff0000500000100001;

	lut_sub lut_5992 ({sk[1385], i_9_, i_10_, i_14_, i_11_, i_15_, n_n254}, x22729x);
	defparam lut_5992.LUT_SIZE = 7;
	defparam lut_5992.mask = 128'h5555ffff5555ffff0001000000105000;

	lut_sub lut_5997 ({sk[1386], n_n197, n_n48, n_n53, x901x, x900x, n_n228}, x22732x);
	defparam lut_5997.LUT_SIZE = 7;
	defparam lut_5997.mask = 128'h5555ffff5555ffff001515150015ffff;

	lut_sub lut_6003 ({sk[1387], n_n283, x922x, x109x, x22729x, x22732x}, x22734x);
	defparam lut_6003.LUT_SIZE = 6;
	defparam lut_6003.mask = 64'h3f3f3f3f5555557f;

	lut_sub lut_6007 ({sk[1388], i_9_, i_10_, i_11_, i_15_, n_n256}, x110x);
	defparam lut_6007.LUT_SIZE = 6;
	defparam lut_6007.mask = 64'h3f3f3f3f00500000;

	lut_sub lut_6010 ({sk[1389], i_14_, i_13_, i_12_, i_15_, n_n259, x187x}, x1643x);
	defparam lut_6010.LUT_SIZE = 7;
	defparam lut_6010.mask = 128'h5555ffff5555ffff5555555575557575;

	lut_sub lut_6015 ({sk[1390], n_n197, n_n100, n_n94, n_n252, x110x, x1643x}, n_n458);
	defparam lut_6015.LUT_SIZE = 7;
	defparam lut_6015.mask = 128'h5555ffff5555ffff00553f7f00ff3fff;

	lut_sub lut_6020 ({sk[1391], x907x, x915x, x911x, n_n258, n_n261, x142x}, x22371x);
	defparam lut_6020.LUT_SIZE = 7;
	defparam lut_6020.mask = 128'h5555ffff5555ffff0000111300001313;

	lut_sub lut_6024 ({sk[1392], n_n13, n_n61, n_n246, n_n100, x168x, x22371x}, x22372x);
	defparam lut_6024.LUT_SIZE = 7;
	defparam lut_6024.mask = 128'h5555ffff5555ffff555f5f5f777f7f7f;

	lut_sub lut_6029 ({sk[1393], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x357x);
	defparam lut_6029.LUT_SIZE = 7;
	defparam lut_6029.mask = 128'h5555ffff5555ffff0000000000010004;

	lut_sub lut_6032 ({sk[1394], i_14_, i_13_, i_12_, i_15_, n_n267, x22377x}, x1758x);
	defparam lut_6032.LUT_SIZE = 7;
	defparam lut_6032.mask = 128'h5555ffff5555ffff5555555575575555;

	lut_sub lut_6036 ({sk[1395], n_n57, n_n56, n_n222, x904x, x357x, x1758x}, n_n454);
	defparam lut_6036.LUT_SIZE = 7;
	defparam lut_6036.mask = 128'h5555ffff5555ffff0000333f5555777f;

	lut_sub lut_6040 ({sk[1396], i_14_, i_13_, i_12_, x904x}, x486x);
	defparam lut_6040.LUT_SIZE = 5;
	defparam lut_6040.mask = 32'h0f0f0005;

	lut_sub lut_6043 ({sk[1397], n_n257, n_n61, n_n6035, n_n100, n_n94, n_n236}, x22381x);
	defparam lut_6043.LUT_SIZE = 7;
	defparam lut_6043.mask = 128'h5555ffff5555ffff05ff37ff3fff3fff;

	lut_sub lut_6049 ({sk[1398], n_n266, x909x, n_n240, x168x, x486x, x22381x}, x22382x);
	defparam lut_6049.LUT_SIZE = 7;
	defparam lut_6049.mask = 128'h5555ffff5555ffff555f555f555f777f;

	lut_sub lut_6053 ({sk[1399], i_9_, i_10_, i_11_, i_15_, n_n256}, x175x);
	defparam lut_6053.LUT_SIZE = 6;
	defparam lut_6053.mask = 64'h3f3f3f3f00000005;

	lut_sub lut_6056 ({sk[1400], i_14_, i_13_, i_12_, x900x, x906x}, x1756x);
	defparam lut_6056.LUT_SIZE = 6;
	defparam lut_6056.mask = 64'h3f3f3f3f07005355;

	lut_sub lut_6063 ({sk[1401], n_n57, n_n56, n_n102, n_n454, x175x, x1756x}, x22383x);
	defparam lut_6063.LUT_SIZE = 7;
	defparam lut_6063.mask = 128'h5555ffff5555ffff0f0f5f5f3fff7fff;

	lut_sub lut_6068 ({sk[1402], i_14_, i_13_, i_12_, x908x}, x140x);
	defparam lut_6068.LUT_SIZE = 5;
	defparam lut_6068.mask = 32'h55ff0045;

	lut_sub lut_6072 ({sk[1403], i_7_, i_8_, i_6_, x915x, x140x}, n_n2738);
	defparam lut_6072.LUT_SIZE = 6;
	defparam lut_6072.mask = 64'h7777777700001000;

	lut_sub lut_6074 ({sk[1404], i_14_, i_13_, i_12_, i_15_, n_n275, n_n259}, x1070x);
	defparam lut_6074.LUT_SIZE = 7;
	defparam lut_6074.mask = 128'h57ff57ff57ff57ff0077000070007070;

	lut_sub lut_6085 ({sk[1405], i_9_, i_10_, i_11_, i_15_, n_n256}, x182x);
	defparam lut_6085.LUT_SIZE = 6;
	defparam lut_6085.mask = 64'h7777777700000500;

	lut_sub lut_6088 ({sk[1406], n_n10, n_n94, n_n252, x142x, x110x, x403x}, x2430x);
	defparam lut_6088.LUT_SIZE = 7;
	defparam lut_6088.mask = 128'h57ff57ff57ff57ff00007fff0000ffff;

	lut_sub lut_6094 ({sk[1407], n_n458, x22372x, x22382x, x22383x, x2430x}, x22394x);
	defparam lut_6094.LUT_SIZE = 6;
	defparam lut_6094.mask = 64'h777777777fffffff;

	lut_sub lut_6100 ({sk[1408], i_14_, i_13_, i_12_, x915x, n_n263, x903x}, n_n6813);
	defparam lut_6100.LUT_SIZE = 7;
	defparam lut_6100.mask = 128'h57ff57ff57ff57ff0000000001000000;

	lut_sub lut_6102 ({sk[1409], i_14_, i_13_, i_12_, x907x, x915x, n_n261}, n_n6826);
	defparam lut_6102.LUT_SIZE = 7;
	defparam lut_6102.mask = 128'h57ff57ff57ff57ff0000000000000001;

	lut_sub lut_6104 ({sk[1410], i_14_, i_13_, i_12_, x905x}, n_n72);
	defparam lut_6104.LUT_SIZE = 5;
	defparam lut_6104.mask = 32'h55ff0004;

	lut_sub lut_6106 ({sk[1411], i_14_, i_13_, i_12_, x914x}, n_n85);
	defparam lut_6106.LUT_SIZE = 5;
	defparam lut_6106.mask = 32'h55ff0100;

	lut_sub lut_6108 ({sk[1412], i_14_, i_13_, i_12_, i_11_, x908x, n_n269}, x19267x);
	defparam lut_6108.LUT_SIZE = 7;
	defparam lut_6108.mask = 128'h57ff57ff57ff57ff5050505050005073;

	lut_sub lut_6113 ({sk[1413], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19265x);
	defparam lut_6113.LUT_SIZE = 7;
	defparam lut_6113.mask = 128'h57ff57ff57ff57ff0400000001000000;

	lut_sub lut_6116 ({sk[1414], i_9_, i_10_, i_11_, i_15_, n_n258, x19265x}, x19268x);
	defparam lut_6116.LUT_SIZE = 7;
	defparam lut_6116.mask = 128'h57ff57ff57ff57ffff555555555557ff;

	lut_sub lut_6121 ({sk[1415], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x5845x);
	defparam lut_6121.LUT_SIZE = 7;
	defparam lut_6121.mask = 128'h57ff57ff57ff57ff0888000000000000;

	lut_sub lut_6124 ({sk[1416], i_14_, i_13_, i_12_, i_11_, x899x, n_n269}, x435x);
	defparam lut_6124.LUT_SIZE = 7;
	defparam lut_6124.mask = 128'h57ff57ff57ff57ff0050335000505050;

	lut_sub lut_6128 ({sk[1417], i_9_, i_10_, i_12_, i_11_}, x287x);
	defparam lut_6128.LUT_SIZE = 5;
	defparam lut_6128.mask = 32'h55ff7000;

	lut_sub lut_6131 ({sk[1418], n_n281, x921x, n_n208, x901x, x5845x, x287x}, x5844x);
	defparam lut_6131.LUT_SIZE = 7;
	defparam lut_6131.mask = 128'h57ff57ff57ff57ff000000770000007f;

	lut_sub lut_6135 ({sk[1419], i_9_, i_10_, i_11_, n_n124, x435x, x5844x}, n_n5029);
	defparam lut_6135.LUT_SIZE = 7;
	defparam lut_6135.mask = 128'h57ff57ff57ff57ff575757575757575f;

	lut_sub lut_6139 ({sk[1420], i_14_, i_13_, i_12_, x901x}, x277x);
	defparam lut_6139.LUT_SIZE = 5;
	defparam lut_6139.mask = 32'h55ff0054;

	lut_sub lut_6143 ({sk[1421], i_14_, i_13_, i_12_, n_n271, x909x, x901x}, n_n4950);
	defparam lut_6143.LUT_SIZE = 7;
	defparam lut_6143.mask = 128'h111fffff111fffff0000000001010100;

	lut_sub lut_6147 ({sk[1422], i_14_, i_13_, i_12_, i_15_, n_n242, n_n270}, x1075x);
	defparam lut_6147.LUT_SIZE = 7;
	defparam lut_6147.mask = 128'h111fffff111fffff0555005557007070;

	lut_sub lut_6160 ({sk[1423], i_7_, i_8_, i_6_, n_n165, n_n284}, x1076x);
	defparam lut_6160.LUT_SIZE = 6;
	defparam lut_6160.mask = 64'h7f7f7f7f11000000;

	lut_sub lut_6163 ({sk[1424], i_14_, i_13_, i_12_, x905x, x899x}, x1273x);
	defparam lut_6163.LUT_SIZE = 6;
	defparam lut_6163.mask = 64'h7f7f7f7f30500305;

	lut_sub lut_6168 ({sk[1425], i_14_, i_13_, i_12_, x913x, x911x, x905x}, x1085x);
	defparam lut_6168.LUT_SIZE = 7;
	defparam lut_6168.mask = 128'h111fffff111fffff5f003300000f0033;

	lut_sub lut_6174 ({sk[1426], i_14_, i_13_, i_12_, x913x, x911x}, x225x);
	defparam lut_6174.LUT_SIZE = 6;
	defparam lut_6174.mask = 64'h7f7f7f7f00000305;

	lut_sub lut_6177 ({sk[1427], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x130x);
	defparam lut_6177.LUT_SIZE = 7;
	defparam lut_6177.mask = 128'h111fffff111fffff4000100000000000;

	lut_sub lut_6180 ({sk[1428], i_14_, i_13_, i_12_, i_15_, n_n267}, x1088x);
	defparam lut_6180.LUT_SIZE = 6;
	defparam lut_6180.mask = 64'h7f7f7f7f15055044;

	lut_sub lut_6190 ({sk[1429], i_7_, i_8_, i_6_, x922x, x908x, n_n256}, n_n6858);
	defparam lut_6190.LUT_SIZE = 7;
	defparam lut_6190.mask = 128'h111fffff111fffff0000010000000000;

	lut_sub lut_6192 ({sk[1430], i_14_, i_13_, i_12_, i_15_, n_n270}, x141x);
	defparam lut_6192.LUT_SIZE = 6;
	defparam lut_6192.mask = 64'h7f7f7f7f00014040;

	lut_sub lut_6196 ({sk[1431], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1913x);
	defparam lut_6196.LUT_SIZE = 7;
	defparam lut_6196.mask = 128'h111fffff111fffff0010001040004000;

	lut_sub lut_6201 ({sk[1432], n_n273, x922x, n_n6504, x470x, x376x, x1913x}, n_n3974);
	defparam lut_6201.LUT_SIZE = 7;
	defparam lut_6201.mask = 128'h111fffff111fffff3fff3fff3fff7fff;

	lut_sub lut_6206 ({sk[1433], i_15_, n_n283, x922x, x368x, n_n137}, n_n4090);
	defparam lut_6206.LUT_SIZE = 6;
	defparam lut_6206.mask = 64'h7f7f7f7f00030007;

	lut_sub lut_6209 ({sk[1434], i_14_, i_13_, i_12_, n_n283, x914x, x922x}, x462x);
	defparam lut_6209.LUT_SIZE = 7;
	defparam lut_6209.mask = 128'h111fffff111fffff0001010000000000;

	lut_sub lut_6212 ({sk[1435], n_n281, n_n283, x914x, x922x, x912x, n_n225}, x464x);
	defparam lut_6212.LUT_SIZE = 7;
	defparam lut_6212.mask = 128'h111fffff111fffff0000000500000307;

	lut_sub lut_6215 ({sk[1436], i_14_, i_13_, i_12_, x907x, n_n273, x922x}, x492x);
	defparam lut_6215.LUT_SIZE = 7;
	defparam lut_6215.mask = 128'h111fffff111fffff0100000000000000;

	lut_sub lut_6217 ({sk[1437], n_n281, x907x, n_n258, n_n53, n_n6520, n_n6511}, x20328x);
	defparam lut_6217.LUT_SIZE = 7;
	defparam lut_6217.mask = 128'h111fffff111fffff7777777f77777f7f;

	lut_sub lut_6222 ({sk[1438], n_n48, n_n11, x495x, x631x, x462x, x464x}, x20330x);
	defparam lut_6222.LUT_SIZE = 7;
	defparam lut_6222.mask = 128'h111fffff111fffff7fff7fff7fffffff;

	lut_sub lut_6228 ({sk[1439], n_n151, n_n226, n_n48, n_n53, x225x, x130x}, x474x);
	defparam lut_6228.LUT_SIZE = 7;
	defparam lut_6228.mask = 128'h111fffff111fffff070707ff07ff07ff;

	lut_sub lut_6233 ({sk[1440], i_14_, i_13_, i_12_, i_15_, x199x, n_n270}, x20335x);
	defparam lut_6233.LUT_SIZE = 7;
	defparam lut_6233.mask = 128'h111fffff111fffff7333373333333333;

	lut_sub lut_6237 ({sk[1441], n_n226, n_n7, n_n222, n_n53, x901x, x89x}, x24193x);
	defparam lut_6237.LUT_SIZE = 7;
	defparam lut_6237.mask = 128'h111fffff111fffff05070f0f0f0f0f0f;

	lut_sub lut_6246 ({sk[1442], x183x, n_n283, x922x, x20335x, x24193x}, x20341x);
	defparam lut_6246.LUT_SIZE = 6;
	defparam lut_6246.mask = 64'h7f7f7f7f5557555f;

	lut_sub lut_6250 ({sk[1443], n_n283, x159x, n_n263, x922x, n_n247, x20333x}, x20339x);
	defparam lut_6250.LUT_SIZE = 7;
	defparam lut_6250.mask = 128'h111fffff111fffff5557555755575f5f;

	lut_sub lut_6254 ({sk[1444], i_14_, i_13_, i_12_, i_15_, x79x, n_n259}, x1854x);
	defparam lut_6254.LUT_SIZE = 7;
	defparam lut_6254.mask = 128'h111fffff111fffff3337333773333333;

	lut_sub lut_6259 ({sk[1445], i_14_, i_13_, i_12_, n_n208, x916x, x900x}, x455x);
	defparam lut_6259.LUT_SIZE = 7;
	defparam lut_6259.mask = 128'h111fffff111fffff0000000000010100;

	lut_sub lut_6262 ({sk[1446], i_14_, i_13_, i_12_, x900x, x906x}, x179x);
	defparam lut_6262.LUT_SIZE = 6;
	defparam lut_6262.mask = 64'h7f7f7f7f00003055;

	lut_sub lut_6266 ({sk[1447], n_n226, x159x, n_n48, n_n60, x475x, x676x}, n_n3184);
	defparam lut_6266.LUT_SIZE = 7;
	defparam lut_6266.mask = 128'h111fffff111fffff777f77ff77ff77ff;

	lut_sub lut_6272 ({sk[1448], n_n208, x916x, n_n258, x899x, x466x, x181x}, x20399x);
	defparam lut_6272.LUT_SIZE = 7;
	defparam lut_6272.mask = 128'h111fffff111fffff333333333333777f;

	lut_sub lut_6276 ({sk[1449], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1915x);
	defparam lut_6276.LUT_SIZE = 7;
	defparam lut_6276.mask = 128'h111fffff111fffff0000000001010104;

	lut_sub lut_6281 ({sk[1450], n_n208, x916x, n_n3, x333x, x188x, x1915x}, x20987x);
	defparam lut_6281.LUT_SIZE = 7;
	defparam lut_6281.mask = 128'h111fffff111fffff0f5f0f5f0f5f3f7f;

	lut_sub lut_6285 ({sk[1451], n_n208, x916x, n_n222, x88x, x902x, x141x}, x20398x);
	defparam lut_6285.LUT_SIZE = 7;
	defparam lut_6285.mask = 128'h111fffff111fffff0000000000005f7f;

	lut_sub lut_6289 ({sk[1452], n_n4, x20399x, x20987x, n_n876, x117x, x20398x}, n_n3116);
	defparam lut_6289.LUT_SIZE = 7;
	defparam lut_6289.mask = 128'h111fffff111fffff5fffffff7fffffff;

	lut_sub lut_6295 ({sk[1453], i_14_, i_13_, i_12_, n_n208, x916x, x899x}, n_n7442);
	defparam lut_6295.LUT_SIZE = 7;
	defparam lut_6295.mask = 128'h111fffff111fffff0000010000000000;

	lut_sub lut_6297 ({sk[1454], i_14_, i_13_, i_12_, n_n208, x916x, x905x}, n_n7443);
	defparam lut_6297.LUT_SIZE = 7;
	defparam lut_6297.mask = 128'h111fffff111fffff0100000000000000;

	lut_sub lut_6299 ({sk[1455], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x174x);
	defparam lut_6299.LUT_SIZE = 7;
	defparam lut_6299.mask = 128'h111fffff111fffff0101000400000000;

	lut_sub lut_6303 ({sk[1456], i_14_, i_13_, i_12_, x898x, x904x, x174x}, x21296x);
	defparam lut_6303.LUT_SIZE = 7;
	defparam lut_6303.mask = 128'h111fffff111fffff555555555f555577;

	lut_sub lut_6307 ({sk[1457], i_14_, i_13_, i_12_, i_15_, n_n253, x21296x}, x1090x);
	defparam lut_6307.LUT_SIZE = 7;
	defparam lut_6307.mask = 128'h111fffff111fffff5555555775557555;

	lut_sub lut_6312 ({sk[1458], n_n273, n_n283, x909x, n_n279, x904x, x906x}, x386x);
	defparam lut_6312.LUT_SIZE = 7;
	defparam lut_6312.mask = 128'h111fffff111fffff0000000300050007;

	lut_sub lut_6315 ({sk[1459], i_14_, i_13_, i_12_, i_15_, n_n267}, x1091x);
	defparam lut_6315.LUT_SIZE = 6;
	defparam lut_6315.mask = 64'h7f7f7f7f00015154;

	lut_sub lut_6323 ({sk[1460], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1092x);
	defparam lut_6323.LUT_SIZE = 7;
	defparam lut_6323.mask = 128'h111fffff111fffff1440404040000000;

	lut_sub lut_6330 ({sk[1461], n_n281, n_n273, n_n283, x922x, x904x, x906x}, x21603x);
	defparam lut_6330.LUT_SIZE = 7;
	defparam lut_6330.mask = 128'h111fffff111fffff0000000000050707;

	lut_sub lut_6334 ({sk[1462], i_9_, i_10_, i_11_, i_15_, n_n279}, x413x);
	defparam lut_6334.LUT_SIZE = 6;
	defparam lut_6334.mask = 64'h7f7f7f7f00000050;

	lut_sub lut_6337 ({sk[1463], n_n110, n_n57, n_n56, x90x, x258x, x413x}, n_n2162);
	defparam lut_6337.LUT_SIZE = 7;
	defparam lut_6337.mask = 128'h111fffff111fffff00770f7f0077ffff;

	lut_sub lut_6342 ({sk[1464], i_9_, i_10_, i_11_, i_15_, n_n279}, x327x);
	defparam lut_6342.LUT_SIZE = 6;
	defparam lut_6342.mask = 64'h7f7f7f7f00500000;

	lut_sub lut_6345 ({sk[1465], i_14_, i_13_, i_12_, x913x, n_n271, x909x}, x783x);
	defparam lut_6345.LUT_SIZE = 7;
	defparam lut_6345.mask = 128'h111fffff111fffff0000010000000000;

	lut_sub lut_6347 ({sk[1466], i_9_, i_10_, i_11_, i_15_, n_n281}, x1096x);
	defparam lut_6347.LUT_SIZE = 6;
	defparam lut_6347.mask = 64'h7f7f7f7f00040004;

	lut_sub lut_6350 ({sk[1467], n_n106, n_n57, n_n56, x90x, x327x, x1096x}, x24214x);
	defparam lut_6350.LUT_SIZE = 7;
	defparam lut_6350.mask = 128'h111fffff111fffff003f777f00ffffff;

	lut_sub lut_6366 ({sk[1468], x913x, n_n220, n_n57, n_n56, x905x, x24214x}, x21493x);
	defparam lut_6366.LUT_SIZE = 7;
	defparam lut_6366.mask = 128'h111fffff111fffff5555557755555f7f;

	lut_sub lut_6370 ({sk[1469], i_9_, i_10_, i_11_, i_15_, n_n281, n_n279}, x21401x);
	defparam lut_6370.LUT_SIZE = 7;
	defparam lut_6370.mask = 128'h111fffff111fffff0000570000005700;

	lut_sub lut_6377 ({sk[1470], i_14_, i_13_, i_12_, i_15_, x905x, n_n275}, x21402x);
	defparam lut_6377.LUT_SIZE = 7;
	defparam lut_6377.mask = 128'h111fffff111fffff0573737355000000;

	lut_sub lut_6387 ({sk[1471], i_14_, i_13_, i_12_, i_15_, n_n242, n_n270}, x1097x);
	defparam lut_6387.LUT_SIZE = 7;
	defparam lut_6387.mask = 128'h111fffff111fffff0770707077000000;

	lut_sub lut_6400 ({sk[1472], i_9_, i_10_, i_11_, i_15_, n_n281}, x1101x);
	defparam lut_6400.LUT_SIZE = 6;
	defparam lut_6400.mask = 64'h7f7f7f7f40004004;

	lut_sub lut_6404 ({sk[1473], i_14_, i_13_, i_12_, x913x, x908x}, x21407x);
	defparam lut_6404.LUT_SIZE = 6;
	defparam lut_6404.mask = 64'h7f7f7f7f53330000;

	lut_sub lut_6409 ({sk[1474], i_14_, i_13_, i_12_, x905x}, x281x);
	defparam lut_6409.LUT_SIZE = 5;
	defparam lut_6409.mask = 32'h7f7f1500;

	lut_sub lut_6413 ({sk[1475], i_14_, i_13_, i_12_, x905x, x899x}, x338x);
	defparam lut_6413.LUT_SIZE = 6;
	defparam lut_6413.mask = 64'h7f7f7f7f50007000;

	lut_sub lut_6417 ({sk[1476], i_14_, i_13_, i_12_, x915x, x911x, n_n263}, x722x);
	defparam lut_6417.LUT_SIZE = 7;
	defparam lut_6417.mask = 128'h111fffff111fffff0000010000000000;

	lut_sub lut_6419 ({sk[1477], n_n208, x916x, n_n222, x899x, x249x, x722x}, x21693x);
	defparam lut_6419.LUT_SIZE = 7;
	defparam lut_6419.mask = 128'h111fffff111fffff555555555555777f;

	lut_sub lut_6423 ({sk[1478], x907x, x915x, n_n220, n_n258, n_n261, x901x}, x645x);
	defparam lut_6423.LUT_SIZE = 7;
	defparam lut_6423.mask = 128'h111fffff111fffff0000001100000313;

	lut_sub lut_6426 ({sk[1479], i_14_, i_13_, i_12_, x903x, x63x}, x1104x);
	defparam lut_6426.LUT_SIZE = 6;
	defparam lut_6426.mask = 64'h7f7f7f7f55555755;

	lut_sub lut_6429 ({sk[1480], i_14_, i_13_, i_12_, i_15_, n_n259, n_n267}, x22210x);
	defparam lut_6429.LUT_SIZE = 7;
	defparam lut_6429.mask = 128'h111fffff111fffff0003050330500000;

	lut_sub lut_6435 ({sk[1481], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1105x);
	defparam lut_6435.LUT_SIZE = 7;
	defparam lut_6435.mask = 128'h111fffff111fffff0000005353000053;

	lut_sub lut_6442 ({sk[1482], i_14_, i_13_, i_12_, x907x, x901x, x220x}, x22209x);
	defparam lut_6442.LUT_SIZE = 7;
	defparam lut_6442.mask = 128'h111fffff111fffff55557755555f5555;

	lut_sub lut_6446 ({sk[1483], x915x, n_n263, x355x, x22210x, x22209x}, x2594x);
	defparam lut_6446.LUT_SIZE = 6;
	defparam lut_6446.mask = 64'h7f7f7f7f0000007f;

	lut_sub lut_6450 ({sk[1484], x915x, n_n220, n_n263, x912x, x500x, x50x}, x24093x);
	defparam lut_6450.LUT_SIZE = 7;
	defparam lut_6450.mask = 128'h111fffff111fffffcccccccccc88cc80;

	lut_sub lut_6455 ({sk[1485], x915x, n_n261, x645x, x1104x, x1105x, x24093x}, x22212x);
	defparam lut_6455.LUT_SIZE = 7;
	defparam lut_6455.mask = 128'h111fffff111fffffaaffaaffaaffbfff;

	lut_sub lut_6460 ({sk[1486], i_9_, i_10_, i_11_, i_15_, n_n256}, x144x);
	defparam lut_6460.LUT_SIZE = 6;
	defparam lut_6460.mask = 64'h7f7f7f7f50000000;

	lut_sub lut_6463 ({sk[1487], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1107x);
	defparam lut_6463.LUT_SIZE = 7;
	defparam lut_6463.mask = 128'h111fffff111fffff0050001040004000;

	lut_sub lut_6469 ({sk[1488], n_n273, n_n280, x922x, n_n32, x461x, x1107x}, n_n1255);
	defparam lut_6469.LUT_SIZE = 7;
	defparam lut_6469.mask = 128'h111fffff111fffff33333333337f33ff;

	lut_sub lut_6474 ({sk[1489], i_14_, i_13_, i_12_, n_n273, x922x, x902x}, n_n6848);
	defparam lut_6474.LUT_SIZE = 7;
	defparam lut_6474.mask = 128'h111fffff111fffff0000000000010000;

	lut_sub lut_6476 ({sk[1490], i_14_, i_13_, i_12_, n_n273, x922x, x908x}, x479x);
	defparam lut_6476.LUT_SIZE = 7;
	defparam lut_6476.mask = 128'h111fffff111fffff0001010000000000;

	lut_sub lut_6479 ({sk[1491], n_n273, n_n222, x922x, x908x, x902x}, x656x);
	defparam lut_6479.LUT_SIZE = 6;
	defparam lut_6479.mask = 64'h7f7f7f7f00000007;

	lut_sub lut_6482 ({sk[1492], i_14_, i_13_, i_12_, x908x, x902x}, x1109x);
	defparam lut_6482.LUT_SIZE = 6;
	defparam lut_6482.mask = 64'h7f7f7f7f05053003;

	lut_sub lut_6487 ({sk[1493], n_n53, n_n6856, x629x, x462x, n_n6848, x1109x}, x22287x);
	defparam lut_6487.LUT_SIZE = 7;
	defparam lut_6487.mask = 128'h111fffff111fffff3fffffff7fffffff;

	lut_sub lut_6493 ({sk[1494], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1110x);
	defparam lut_6493.LUT_SIZE = 7;
	defparam lut_6493.mask = 128'h111fffff111fffff0350000053000000;

	lut_sub lut_6498 ({sk[1495], n_n4, n_n3, x648x, n_n62, n_n10, x1110x}, n_n1157);
	defparam lut_6498.LUT_SIZE = 7;
	defparam lut_6498.mask = 128'h111fffff111fffff00ff77ff3fff7fff;

	lut_sub lut_6504 ({sk[1496], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1112x);
	defparam lut_6504.LUT_SIZE = 7;
	defparam lut_6504.mask = 128'h111fffff111fffff0003530000535300;

	lut_sub lut_6512 ({sk[1497], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1111x);
	defparam lut_6512.LUT_SIZE = 7;
	defparam lut_6512.mask = 128'h111fffff111fffff0053530000000000;

	lut_sub lut_6517 ({sk[1498], n_n4, n_n3, n_n7441, n_n7442, x1112x, x1111x}, x21920x);
	defparam lut_6517.LUT_SIZE = 7;
	defparam lut_6517.mask = 128'h111fffff111fffff0fff3fff5fff7fff;

	lut_sub lut_6522 ({sk[1499], i_15_, x915x, x914x, n_n279, n_n263, n_n137}, x3786x);
	defparam lut_6522.LUT_SIZE = 7;
	defparam lut_6522.mask = 128'h111fffff111fffff0000111300000003;

	lut_sub lut_6525 ({sk[1500], i_14_, i_13_, i_12_, x908x, x902x}, x1933x);
	defparam lut_6525.LUT_SIZE = 6;
	defparam lut_6525.mask = 64'h7f7f7f7f55053033;

	lut_sub lut_6532 ({sk[1501], x915x, n_n261, x49x, n_n6834, x3786x, x1933x}, x22193x);
	defparam lut_6532.LUT_SIZE = 7;
	defparam lut_6532.mask = 128'h111fffff111fffff3f3f3f3f3f3f7fff;

	lut_sub lut_6537 ({sk[1502], i_14_, i_13_, i_12_, i_15_, n_n275, n_n259}, x1114x);
	defparam lut_6537.LUT_SIZE = 7;
	defparam lut_6537.mask = 128'h111fffff111fffff0337300770037770;

	lut_sub lut_6554 ({sk[1503], i_14_, i_13_, i_12_, x915x, n_n263, x902x}, x2601x);
	defparam lut_6554.LUT_SIZE = 7;
	defparam lut_6554.mask = 128'h111fffff111fffff0101000100010100;

	lut_sub lut_6560 ({sk[1504], n_n197, n_n100, x3776x, n_n2738, x1114x, x2601x}, x22201x);
	defparam lut_6560.LUT_SIZE = 7;
	defparam lut_6560.mask = 128'h111fffff111fffff5fff7fff5fffffff;

	lut_sub lut_6566 ({sk[1505], n_n94, n_n6814, n_n6813, x257x, x1333x, x22187x}, n_n1295);
	defparam lut_6566.LUT_SIZE = 7;
	defparam lut_6566.mask = 128'h111fffff111fffff55ffffff7fffffff;

	lut_sub lut_6572 ({sk[1506], n_n111, n_n135, n_n103, n_n94, x688x, x5529x}, x22192x);
	defparam lut_6572.LUT_SIZE = 7;
	defparam lut_6572.mask = 128'h111fffff111fffff777f7f7f7f7f7f7f;

	lut_sub lut_6578 ({sk[1507], x22184x, x22185x, x22193x, x22201x, n_n1295, x22192x}, n_n1102);
	defparam lut_6578.LUT_SIZE = 7;
	defparam lut_6578.mask = 128'h111fffff111fffff7fffffffffffffff;

	lut_sub lut_6585 ({sk[1508], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1168x);
	defparam lut_6585.LUT_SIZE = 7;
	defparam lut_6585.mask = 128'h111fffff111fffff0003530000005300;

	lut_sub lut_6591 ({sk[1509], i_14_, i_13_, i_12_, i_15_, n_n267}, x1167x);
	defparam lut_6591.LUT_SIZE = 6;
	defparam lut_6591.mask = 64'h7f7f7f7f00014154;

	lut_sub lut_6598 ({sk[1510], x915x, n_n271, x909x, n_n261, x1168x, x1167x}, x22220x);
	defparam lut_6598.LUT_SIZE = 7;
	defparam lut_6598.mask = 128'h111fffff111fffff0000005503030357;

	lut_sub lut_6601 ({sk[1511], i_7_, i_8_, i_6_, x909x, x81x, n_n42}, n_n4681);
	defparam lut_6601.LUT_SIZE = 7;
	defparam lut_6601.mask = 128'h111fffff111fffff0000000000050003;

	lut_sub lut_6604 ({sk[1512], i_14_, i_13_, i_12_, i_15_, x900x, n_n267}, x300x);
	defparam lut_6604.LUT_SIZE = 7;
	defparam lut_6604.mask = 128'h111fffff111fffff3373000000000000;

	lut_sub lut_6608 ({sk[1513], i_14_, i_13_, i_12_, i_15_, n_n253, x300x}, x1115x);
	defparam lut_6608.LUT_SIZE = 7;
	defparam lut_6608.mask = 128'h111fffff111fffff5755555555557775;

	lut_sub lut_6614 ({sk[1514], n_n57, n_n56, n_n54, x51x, x81x, n_n42}, x22225x);
	defparam lut_6614.LUT_SIZE = 7;
	defparam lut_6614.mask = 128'h111fffff111fffff000055ff3f3f7fff;

	lut_sub lut_6619 ({sk[1515], n_n57, n_n56, x166x, x303x, x497x, x1115x}, x22228x);
	defparam lut_6619.LUT_SIZE = 7;
	defparam lut_6619.mask = 128'h111fffff111fffff333377773fff7fff;

	lut_sub lut_6624 ({sk[1516], n_n271, x909x, n_n4960, x45x, x22225x, x22228x}, x22229x);
	defparam lut_6624.LUT_SIZE = 7;
	defparam lut_6624.mask = 128'h111fffff111fffff77ff77ff77ff7fff;

	lut_sub lut_6629 ({sk[1517], n_n57, n_n6036, n_n6035, x45x, x486x, x2589x}, n_n1284);
	defparam lut_6629.LUT_SIZE = 7;
	defparam lut_6629.mask = 128'h111fffff111fffff55ffffff7fffffff;

	lut_sub lut_6635 ({sk[1518], n_n57, x484x, n_n50, n_n94, x722x, x1166x}, x22219x);
	defparam lut_6635.LUT_SIZE = 7;
	defparam lut_6635.mask = 128'h111fffff111fffff3737ffff37ffffff;

	lut_sub lut_6640 ({sk[1519], x2594x, x22212x, x22220x, n_n1284, x22219x}, x22230x);
	defparam lut_6640.LUT_SIZE = 6;
	defparam lut_6640.mask = 64'h7f7f7f7f7fffffff;

	lut_sub lut_6646 ({sk[1520], i_7_, i_8_, i_6_, x915x, n_n41, n_n216}, x22242x);
	defparam lut_6646.LUT_SIZE = 7;
	defparam lut_6646.mask = 128'h111fffff111fffff0000000000030005;

	lut_sub lut_6649 ({sk[1521], i_8_, n_n153, x915x, x822x, n_n258, x899x}, x22240x);
	defparam lut_6649.LUT_SIZE = 7;
	defparam lut_6649.mask = 128'h111fffff111fffff0f0f0f1f0f0f0f0f;

	lut_sub lut_6652 ({sk[1522], x907x, n_n273, n_n283, x914x, x909x, n_n279}, x22241x);
	defparam lut_6652.LUT_SIZE = 7;
	defparam lut_6652.mask = 128'h111fffff111fffff0001000100011111;

	lut_sub lut_6655 ({sk[1523], x515x, x569x, x524x, x22242x, x22240x, x22241x}, x22246x);
	defparam lut_6655.LUT_SIZE = 7;
	defparam lut_6655.mask = 128'h111fffff111fffff7fffffffffffffff;

	lut_sub lut_6662 ({sk[1524], i_14_, i_13_, i_12_, x915x, x898x, n_n263}, x599x);
	defparam lut_6662.LUT_SIZE = 7;
	defparam lut_6662.mask = 128'h111fffff111fffff0000000000010000;

	lut_sub lut_6664 ({sk[1525], i_14_, i_13_, i_12_, x900x, x906x}, x1936x);
	defparam lut_6664.LUT_SIZE = 6;
	defparam lut_6664.mask = 64'h7f7f7f7f33035055;

	lut_sub lut_6671 ({sk[1526], i_14_, i_13_, i_12_, i_15_, x906x, n_n253}, x1117x);
	defparam lut_6671.LUT_SIZE = 7;
	defparam lut_6671.mask = 128'h111fffff111fffff0555730550005550;

	lut_sub lut_6682 ({sk[1527], i_14_, i_13_, i_12_, i_15_, n_n247, n_n267}, x1116x);
	defparam lut_6682.LUT_SIZE = 7;
	defparam lut_6682.mask = 128'h111fffff111fffff0000000330073730;

	lut_sub lut_6691 ({sk[1528], x915x, n_n54, x51x, n_n261, n_n263, x1936x}, x22251x);
	defparam lut_6691.LUT_SIZE = 7;
	defparam lut_6691.mask = 128'h111fffff111fffff00000000050f373f;

	lut_sub lut_6695 ({sk[1529], x915x, n_n261, n_n263, x1117x, x1116x, x22251x}, x22253x);
	defparam lut_6695.LUT_SIZE = 7;
	defparam lut_6695.mask = 128'h111fffff111fffff55555555555f777f;

	lut_sub lut_6699 ({sk[1530], i_14_, i_13_, i_12_, x915x, n_n261, x901x}, n_n6824);
	defparam lut_6699.LUT_SIZE = 7;
	defparam lut_6699.mask = 128'h111fffff111fffff0000000000010000;

	lut_sub lut_6701 ({sk[1531], i_7_, i_8_, i_6_, x915x, x112x}, x798x);
	defparam lut_6701.LUT_SIZE = 6;
	defparam lut_6701.mask = 64'h7f7f7f7f00001000;

	lut_sub lut_6703 ({sk[1532], n_n100, n_n94, n_n87, x548x, x1292x, x22231x}, n_n1298);
	defparam lut_6703.LUT_SIZE = 7;
	defparam lut_6703.mask = 128'h111fffff111fffff5f5f5fff7f7f7fff;

	lut_sub lut_6708 ({sk[1533], n_n100, n_n94, x1294x, x1293x, x1386x, x1385x}, x24092x);
	defparam lut_6708.LUT_SIZE = 7;
	defparam lut_6708.mask = 128'h111fffff111fffffffffcc00a0a08000;

	lut_sub lut_6713 ({sk[1534], n_n6826, x22246x, n_n6824, x798x, n_n1298, x24092x}, x22254x);
	defparam lut_6713.LUT_SIZE = 7;
	defparam lut_6713.mask = 128'h111fffff111fffffbfffffffffffffff;

	lut_sub lut_6720 ({sk[1535], i_14_, i_13_, i_12_, i_15_, x911x, n_n242}, x1901x);
	defparam lut_6720.LUT_SIZE = 7;
	defparam lut_6720.mask = 128'h111fffff111fffff0000000005330550;

	lut_sub lut_6725 ({sk[1536], i_14_, i_13_, i_12_, x907x, x901x, x177x}, x1119x);
	defparam lut_6725.LUT_SIZE = 7;
	defparam lut_6725.mask = 128'h111fffff111fffff5555557f55775577;

	lut_sub lut_6731 ({sk[1537], i_14_, i_13_, i_12_, x898x, x904x}, x356x);
	defparam lut_6731.LUT_SIZE = 6;
	defparam lut_6731.mask = 64'h7f7f7f7f00070005;

	lut_sub lut_6735 ({sk[1538], x915x, x911x, n_n261, n_n263, x899x, n_n228}, x22613x);
	defparam lut_6735.LUT_SIZE = 7;
	defparam lut_6735.mask = 128'h111fffff111fffff0000000001010555;

	lut_sub lut_6739 ({sk[1539], i_9_, i_10_, i_11_, i_15_, n_n225}, x139x);
	defparam lut_6739.LUT_SIZE = 6;
	defparam lut_6739.mask = 64'h7f7f7f7f00050000;

	lut_sub lut_6742 ({sk[1540], i_14_, i_13_, i_12_, x900x, x906x}, x335x);
	defparam lut_6742.LUT_SIZE = 6;
	defparam lut_6742.mask = 64'h7f7f7f7f00070005;

	lut_sub lut_6746 ({sk[1541], n_n228, x912x, x902x, n_n100, n_n94, x897x}, x22618x);
	defparam lut_6746.LUT_SIZE = 7;
	defparam lut_6746.mask = 128'h111fffff111fffff00000000153f3f3f;

	lut_sub lut_6753 ({sk[1542], i_7_, i_8_, i_6_, x909x, x224x, x22618x}, x22620x);
	defparam lut_6753.LUT_SIZE = 7;
	defparam lut_6753.mask = 128'h111fffff111fffff5555555555575557;

	lut_sub lut_6757 ({sk[1543], i_7_, i_8_, i_6_, x909x, x335x}, x2138x);
	defparam lut_6757.LUT_SIZE = 6;
	defparam lut_6757.mask = 64'h7f7f7f7f00000100;

	lut_sub lut_6759 ({sk[1544], x915x, n_n261, n_n263, x899x, x901x, n_n228}, x22616x);
	defparam lut_6759.LUT_SIZE = 7;
	defparam lut_6759.mask = 128'h111fffff111fffff0000000000111515;

	lut_sub lut_6763 ({sk[1545], n_n57, n_n4970, x356x, x22613x, x2138x, x22616x}, x22621x);
	defparam lut_6763.LUT_SIZE = 7;
	defparam lut_6763.mask = 128'h111fffff111fffff7f7fffff7fffffff;

	lut_sub lut_6769 ({sk[1546], i_14_, i_13_, i_12_, i_15_, x902x, n_n270}, x1918x);
	defparam lut_6769.LUT_SIZE = 7;
	defparam lut_6769.mask = 128'h111fffff111fffff0000000005053350;

	lut_sub lut_6774 ({sk[1547], x909x, n_n261, n_n263, x120x, x91x, x1918x}, n_n816);
	defparam lut_6774.LUT_SIZE = 7;
	defparam lut_6774.mask = 128'h111fffff111fffff0000000000553f7f;

	lut_sub lut_6778 ({sk[1548], n_n53, n_n6860, x142x, x123x, x752x, x110x}, x22400x);
	defparam lut_6778.LUT_SIZE = 7;
	defparam lut_6778.mask = 128'h111fffff111fffff3333ffff7fffffff;

	lut_sub lut_6784 ({sk[1549], n_n273, x905x, x922x, x899x, n_n256}, x624x);
	defparam lut_6784.LUT_SIZE = 6;
	defparam lut_6784.mask = 64'h7f7f7f7f00000105;

	lut_sub lut_6787 ({sk[1550], i_9_, i_10_, i_11_, i_15_, n_n256, x142x}, x1496x);
	defparam lut_6787.LUT_SIZE = 7;
	defparam lut_6787.mask = 128'h111fffff111fffff5555775555555555;

	lut_sub lut_6791 ({sk[1551], i_14_, i_13_, i_12_, i_15_, n_n259, n_n270}, x1498x);
	defparam lut_6791.LUT_SIZE = 7;
	defparam lut_6791.mask = 128'h111fffff111fffff0055000070007070;

	lut_sub lut_6800 ({sk[1552], n_n216, n_n48, n_n53, x624x, x1496x, x1498x}, x22401x);
	defparam lut_6800.LUT_SIZE = 7;
	defparam lut_6800.mask = 128'h111fffff111fffff0f0f7f7f0fffffff;

	lut_sub lut_6806 ({sk[1553], i_14_, i_13_, i_12_, x907x, x914x, x904x}, x1739x);
	defparam lut_6806.LUT_SIZE = 7;
	defparam lut_6806.mask = 128'h111fffff111fffff000000000f770f0f;

	lut_sub lut_6812 ({sk[1554], n_n53, x457x, x20333x, n_n6504, x144x, x1739x}, x22412x);
	defparam lut_6812.LUT_SIZE = 7;
	defparam lut_6812.mask = 128'h111fffff111fffff0fffffff7fffffff;

	lut_sub lut_6818 ({sk[1555], n_n283, x914x, x922x, x912x, n_n256, x189x}, x630x);
	defparam lut_6818.LUT_SIZE = 7;
	defparam lut_6818.mask = 128'h111fffff111fffff0000000000570077;

	lut_sub lut_6822 ({sk[1556], i_14_, i_13_, i_12_, i_15_, x900x, n_n267}, x1124x);
	defparam lut_6822.LUT_SIZE = 7;
	defparam lut_6822.mask = 128'h111fffff111fffff0055000050335050;

	lut_sub lut_6829 ({sk[1557], i_14_, i_13_, i_12_, i_15_, n_n253, x1124x}, x1123x);
	defparam lut_6829.LUT_SIZE = 7;
	defparam lut_6829.mask = 128'h111fffff111fffff5557555575557555;

	lut_sub lut_6834 ({sk[1558], x909x, n_n261, n_n263, x1124x, x1123x, x357x}, x22420x);
	defparam lut_6834.LUT_SIZE = 7;
	defparam lut_6834.mask = 128'h111fffff111fffff00000000005f337f;

	lut_sub lut_6838 ({sk[1559], n_n6, n_n6524, n_n98, n_n49, n_n6517, n_n6520}, x24155x);
	defparam lut_6838.LUT_SIZE = 7;
	defparam lut_6838.mask = 128'h111fffff111fffff8888000080000000;

	lut_sub lut_6841 ({sk[1560], x630x, x22420x, x24155x}, x22421x);
	defparam lut_6841.LUT_SIZE = 4;
	defparam lut_6841.mask = 16'h33bf;

	lut_sub lut_6845 ({sk[1561], n_n240, n_n61, n_n48, n_n53, n_n6520, x22406x}, n_n431);
	defparam lut_6845.LUT_SIZE = 7;
	defparam lut_6845.mask = 128'h111fffff111fffff77777f7f7fff7fff;

	lut_sub lut_6851 ({sk[1562], x907x, n_n258, n_n48, n_n53, x906x, x1738x}, x22411x);
	defparam lut_6851.LUT_SIZE = 7;
	defparam lut_6851.mask = 128'h111fffff111fffff0055037700550f7f;

	lut_sub lut_6856 ({sk[1563], x22400x, x22401x, x22412x, n_n431, x22411x}, x22422x);
	defparam lut_6856.LUT_SIZE = 6;
	defparam lut_6856.mask = 64'h7f7f7f7f7fffffff;

	lut_sub lut_6862 ({sk[1564], i_14_, i_13_, i_12_, i_15_, n_n247, x233x}, x1700x);
	defparam lut_6862.LUT_SIZE = 7;
	defparam lut_6862.mask = 128'h111fffff111fffff5557555575577575;

	lut_sub lut_6869 ({sk[1565], x914x, x909x, n_n261, n_n256, x1700x}, x22432x);
	defparam lut_6869.LUT_SIZE = 6;
	defparam lut_6869.mask = 64'h7f7f7f7f00050007;

	lut_sub lut_6872 ({sk[1566], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x359x);
	defparam lut_6872.LUT_SIZE = 7;
	defparam lut_6872.mask = 128'h111fffff111fffff0010000040004000;

	lut_sub lut_6876 ({sk[1567], i_14_, i_13_, i_12_, i_15_, x907x, n_n282}, x1608x);
	defparam lut_6876.LUT_SIZE = 7;
	defparam lut_6876.mask = 128'h111fffff111fffff0037000050005000;

	lut_sub lut_6881 ({sk[1568], i_14_, i_13_, i_12_, x914x, x912x}, x351x);
	defparam lut_6881.LUT_SIZE = 6;
	defparam lut_6881.mask = 64'h7f7f7f7f00000503;

	lut_sub lut_6884 ({sk[1569], i_14_, i_13_, i_12_, i_15_, n_n282, n_n253}, x1701x);
	defparam lut_6884.LUT_SIZE = 7;
	defparam lut_6884.mask = 128'h111fffff111fffff0077000070037030;

	lut_sub lut_6895 ({sk[1570], n_n6, n_n5, x359x, x1608x, x351x, x1701x}, x22433x);
	defparam lut_6895.LUT_SIZE = 7;
	defparam lut_6895.mask = 128'h111fffff111fffff000077ff0f0f7fff;

	lut_sub lut_6900 ({sk[1571], i_14_, i_13_, i_12_, i_15_, n_n275, n_n270}, x1126x);
	defparam lut_6900.LUT_SIZE = 7;
	defparam lut_6900.mask = 128'h111fffff111fffff0077000070057050;

	lut_sub lut_6911 ({sk[1572], i_14_, i_13_, i_12_, x905x, x899x}, x306x);
	defparam lut_6911.LUT_SIZE = 6;
	defparam lut_6911.mask = 64'h7f7f7f7f00000503;

	lut_sub lut_6914 ({sk[1573], i_14_, i_13_, i_12_, i_15_, n_n275, x306x}, x1125x);
	defparam lut_6914.LUT_SIZE = 7;
	defparam lut_6914.mask = 128'h111fffff111fffff5577555575577575;

	lut_sub lut_6922 ({sk[1574], i_14_, i_13_, i_12_, i_15_, n_n270, x276x}, x1645x);
	defparam lut_6922.LUT_SIZE = 7;
	defparam lut_6922.mask = 128'h111fffff111fffff5577555575557555;

	lut_sub lut_6928 ({sk[1575], i_14_, i_13_, i_12_, x914x, x903x, x897x}, x1644x);
	defparam lut_6928.LUT_SIZE = 7;
	defparam lut_6928.mask = 128'h111fffff111fffff000f000000550033;

	lut_sub lut_6932 ({sk[1576], n_n6, n_n5, x1126x, x1125x, x1645x, x1644x}, x22440x);
	defparam lut_6932.LUT_SIZE = 7;
	defparam lut_6932.mask = 128'h111fffff111fffff000055ff3f3f7fff;

	lut_sub lut_6937 ({sk[1577], n_n6, n_n5, n_n246, n_n70, x308x, x1649x}, n_n418);
	defparam lut_6937.LUT_SIZE = 7;
	defparam lut_6937.mask = 128'h111fffff111fffff00007f7f55ff7fff;

	lut_sub lut_6943 ({sk[1578], n_n6, n_n5, n_n70, x1652x, x1651x, x306x}, x24173x);
	defparam lut_6943.LUT_SIZE = 7;
	defparam lut_6943.mask = 128'h111fffff111fffffffffa0a0cc008000;

	lut_sub lut_6948 ({sk[1579], i_7_, i_8_, i_6_, x922x, x902x, n_n256}, x578x);
	defparam lut_6948.LUT_SIZE = 7;
	defparam lut_6948.mask = 128'h111fffff111fffff0000010000000000;

	lut_sub lut_6950 ({sk[1580], i_14_, i_13_, i_12_, x903x, x897x}, x1518x);
	defparam lut_6950.LUT_SIZE = 6;
	defparam lut_6950.mask = 64'h7f7f7f7f07003033;

	lut_sub lut_6956 ({sk[1581], n_n31, n_n48, n_n53, n_n6858, x578x, x1518x}, x22447x);
	defparam lut_6956.LUT_SIZE = 7;
	defparam lut_6956.mask = 128'h111fffff111fffff3f7f7f7f3f7fffff;

	lut_sub lut_6962 ({sk[1582], i_14_, i_13_, i_12_, x907x}, x112x);
	defparam lut_6962.LUT_SIZE = 5;
	defparam lut_6962.mask = 32'h7f7f0045;

	lut_sub lut_6966 ({sk[1583], n_n273, n_n283, n_n104, x922x, x144x, x112x}, n_n439);
	defparam lut_6966.LUT_SIZE = 7;
	defparam lut_6966.mask = 128'h111fffff111fffff00000707050f070f;

	lut_sub lut_6971 ({sk[1584], i_9_, i_10_, i_11_, i_15_, n_n256}, x229x);
	defparam lut_6971.LUT_SIZE = 6;
	defparam lut_6971.mask = 64'h7f7f7f7f00050000;

	lut_sub lut_6974 ({sk[1585], i_7_, i_8_, i_6_, x922x, n_n105, x175x}, x22454x);
	defparam lut_6974.LUT_SIZE = 7;
	defparam lut_6974.mask = 128'h111fffff111fffff0300070000000000;

	lut_sub lut_6978 ({sk[1586], n_n283, x166x, x922x, x229x, x22454x}, n_n442);
	defparam lut_6978.LUT_SIZE = 6;
	defparam lut_6978.mask = 64'h7f7f7f7f5555575f;

	lut_sub lut_6982 ({sk[1587], i_14_, i_13_, i_12_, n_n273, x922x, x912x}, x677x);
	defparam lut_6982.LUT_SIZE = 7;
	defparam lut_6982.mask = 128'h111fffff111fffff0000000000010000;

	lut_sub lut_6984 ({sk[1588], i_14_, i_13_, i_12_, i_15_, n_n247, n_n267}, x1128x);
	defparam lut_6984.LUT_SIZE = 7;
	defparam lut_6984.mask = 128'h111fffff111fffff0077000070007070;

	lut_sub lut_6995 ({sk[1589], n_n104, n_n54, n_n48, x677x, x41x, x175x}, x22463x);
	defparam lut_6995.LUT_SIZE = 7;
	defparam lut_6995.mask = 128'h111fffff111fffff0f7f0fff0fff0fff;

	lut_sub lut_7001 ({sk[1590], n_n273, x922x, n_n6504, x144x, n_n6848, x630x}, n_n438);
	defparam lut_7001.LUT_SIZE = 7;
	defparam lut_7001.mask = 128'h111fffff111fffff77ff77ff77ff7fff;

	lut_sub lut_7006 ({sk[1591], n_n56, n_n257, x407x, x457x, n_n4183, x2328x}, n_n443);
	defparam lut_7006.LUT_SIZE = 7;
	defparam lut_7006.mask = 128'h111fffff111fffff7fff7fff7fffffff;

	lut_sub lut_7012 ({sk[1592], i_7_, i_8_, i_6_, n_n103, x922x, x140x}, x22446x);
	defparam lut_7012.LUT_SIZE = 7;
	defparam lut_7012.mask = 128'h111fffff111fffff0300130000000000;

	lut_sub lut_7016 ({sk[1593], x914x, n_n56, n_n258, x908x, x2319x, x2321x}, x22457x);
	defparam lut_7016.LUT_SIZE = 7;
	defparam lut_7016.mask = 128'h111fffff111fffff7777777f777777ff;

	lut_sub lut_7021 ({sk[1594], i_14_, i_13_, i_12_, x915x, n_n263, x903x}, n_n6812);
	defparam lut_7021.LUT_SIZE = 7;
	defparam lut_7021.mask = 128'h111fffff111fffff0000000000000100;

	lut_sub lut_7023 ({sk[1595], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x5905x);
	defparam lut_7023.LUT_SIZE = 7;
	defparam lut_7023.mask = 128'h111fffff111fffff5554000000000000;

	lut_sub lut_7027 ({sk[1596], i_9_, i_10_, i_11_, i_15_, n_n228, x5905x}, x1130x);
	defparam lut_7027.LUT_SIZE = 7;
	defparam lut_7027.mask = 128'h111fffff111fffffff7555ff55555555;

	lut_sub lut_7032 ({sk[1597], i_14_, i_13_, i_12_, x911x, n_n242, n_n207}, x5900x);
	defparam lut_7032.LUT_SIZE = 7;
	defparam lut_7032.mask = 128'h111fffff111fffff0000001105000005;

	lut_sub lut_7036 ({sk[1598], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19218x);
	defparam lut_7036.LUT_SIZE = 7;
	defparam lut_7036.mask = 128'h111fffff111fffff000000001000df55;

	lut_sub lut_7042 ({sk[1599], i_14_, i_13_, i_12_, x899x, x908x, x19218x}, x1132x);
	defparam lut_7042.LUT_SIZE = 7;
	defparam lut_7042.mask = 128'h111fffff111fffff555555555f775f5f;

	lut_sub lut_7048 ({sk[1600], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19221x);
	defparam lut_7048.LUT_SIZE = 7;
	defparam lut_7048.mask = 128'h111fffff111fffff0000aa8a44000000;

	lut_sub lut_7054 ({sk[1601], i_14_, i_13_, i_12_, x911x, n_n247, x908x}, x19222x);
	defparam lut_7054.LUT_SIZE = 7;
	defparam lut_7054.mask = 128'h111fffff111fffff33333333773f7733;

	lut_sub lut_7059 ({sk[1602], n_n227, x1130x, x5900x, x1132x, x19221x, x19222x}, n_n5019);
	defparam lut_7059.LUT_SIZE = 7;
	defparam lut_7059.mask = 128'h111fffff111fffff00ff00ff7fffffff;

	lut_sub lut_7065 ({sk[1603], i_14_, i_13_, i_12_, x897x}, x190x);
	defparam lut_7065.LUT_SIZE = 5;
	defparam lut_7065.mask = 32'h7f7f0054;

	lut_sub lut_7069 ({sk[1604], i_7_, i_8_, i_6_, x909x, x189x}, n_n4941);
	defparam lut_7069.LUT_SIZE = 6;
	defparam lut_7069.mask = 64'h7f7f7f7f00000100;

	lut_sub lut_7071 ({sk[1605], i_7_, i_8_, i_6_, x909x, x219x}, n_n4942);
	defparam lut_7071.LUT_SIZE = 6;
	defparam lut_7071.mask = 64'h7f7f7f7f00000100;

	lut_sub lut_7073 ({sk[1606], i_7_, i_8_, i_6_, x268x, x909x}, n_n4947);
	defparam lut_7073.LUT_SIZE = 6;
	defparam lut_7073.mask = 64'h7f7f7f7f00000100;

	lut_sub lut_7075 ({sk[1607], n_n271, x909x, x912x, n_n225, x87x}, n_n4940);
	defparam lut_7075.LUT_SIZE = 6;
	defparam lut_7075.mask = 64'h7f7f7f7f00000057;

	lut_sub lut_7078 ({sk[1608], i_7_, i_8_, i_6_, x909x, x157x}, x5325x);
	defparam lut_7078.LUT_SIZE = 6;
	defparam lut_7078.mask = 64'h7f7f7f7f00000100;

	lut_sub lut_7080 ({sk[1609], n_n153, x260x, n_n283, n_n5693, n_n274, x910x}, x20021x);
	defparam lut_7080.LUT_SIZE = 7;
	defparam lut_7080.mask = 128'h111fffff111fffff0f1f0f3f0f1fffff;

	lut_sub lut_7085 ({sk[1610], i_9_, i_10_, i_7_, i_8_, i_6_, x910x}, x4892x);
	defparam lut_7085.LUT_SIZE = 7;
	defparam lut_7085.mask = 128'h111fffff111fffff0400000000000000;

	lut_sub lut_7087 ({sk[1611], i_7_, i_6_, n_n5673, x920x, x918x, x261x}, x20027x);
	defparam lut_7087.LUT_SIZE = 7;
	defparam lut_7087.mask = 128'h111fffff111fffff77ff3fff00ff00ff;

	lut_sub lut_7093 ({sk[1612], i_14_, i_13_, i_12_, x911x, n_n57, x84x}, n_n4394);
	defparam lut_7093.LUT_SIZE = 7;
	defparam lut_7093.mask = 128'h111fffff111fffff1311111111111111;

	lut_sub lut_7096 ({sk[1613], i_14_, i_13_, i_12_, i_15_, n_n242, n_n259}, x1138x);
	defparam lut_7096.LUT_SIZE = 7;
	defparam lut_7096.mask = 128'h111fffff111fffff0737303755055550;

	lut_sub lut_7112 ({sk[1614], i_14_, i_13_, i_12_, i_15_, x911x, n_n138}, x217x);
	defparam lut_7112.LUT_SIZE = 7;
	defparam lut_7112.mask = 128'h111fffff111fffff0505050537370505;

	lut_sub lut_7116 ({sk[1615], i_14_, i_13_, i_12_, i_15_, n_n242, x217x}, x1137x);
	defparam lut_7116.LUT_SIZE = 7;
	defparam lut_7116.mask = 128'h111fffff111fffff5575757575557575;

	lut_sub lut_7124 ({sk[1616], n_n266, n_n271, x909x, n_n4394, x1138x, x1137x}, n_n4316);
	defparam lut_7124.LUT_SIZE = 7;
	defparam lut_7124.mask = 128'h111fffff111fffff0f0f0f3f0f5f0f7f;

	lut_sub lut_7128 ({sk[1617], i_14_, i_13_, i_12_, x903x, x897x}, x133x);
	defparam lut_7128.LUT_SIZE = 6;
	defparam lut_7128.mask = 64'h7f7f7f7f00500305;

	lut_sub lut_7132 ({sk[1618], i_14_, i_13_, i_12_, x903x, x897x}, x137x);
	defparam lut_7132.LUT_SIZE = 6;
	defparam lut_7132.mask = 64'h7f7f7f7f00000305;

	lut_sub lut_7135 ({sk[1619], n_n266, n_n271, x909x, n_n7, x133x, x137x}, x473x);
	defparam lut_7135.LUT_SIZE = 7;
	defparam lut_7135.mask = 128'h111fffff111fffff0000003f0055007f;

	lut_sub lut_7139 ({sk[1620], i_14_, i_13_, i_12_, i_15_, n_n282, x314x}, x1140x);
	defparam lut_7139.LUT_SIZE = 7;
	defparam lut_7139.mask = 128'h111fffff111fffff7555575555755557;

	lut_sub lut_7145 ({sk[1621], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x1139x);
	defparam lut_7145.LUT_SIZE = 7;
	defparam lut_7145.mask = 128'h111fffff111fffff0400010000440010;

	lut_sub lut_7151 ({sk[1622], n_n266, n_n271, n_n9, x184x, x909x, x209x}, x19694x);
	defparam lut_7151.LUT_SIZE = 7;
	defparam lut_7151.mask = 128'h111fffff111fffff0000030311331333;

	lut_sub lut_7155 ({sk[1623], n_n9, n_n57, n_n56, x1140x, x1139x, x132x}, x19697x);
	defparam lut_7155.LUT_SIZE = 7;
	defparam lut_7155.mask = 128'h111fffff111fffff00335f7f00ff5fff;

	lut_sub lut_7160 ({sk[1624], i_14_, i_13_, i_12_, n_n266, x909x, x897x}, n_n4930);
	defparam lut_7160.LUT_SIZE = 7;
	defparam lut_7160.mask = 128'h111fffff111fffff0000000001010100;

	lut_sub lut_7164 ({sk[1625], n_n139, n_n124, n_n127, n_n132, n_n107, x250x}, n_n4280);
	defparam lut_7164.LUT_SIZE = 7;
	defparam lut_7164.mask = 128'h111fffff111fffff0377777757777777;

	lut_sub lut_7171 ({sk[1626], i_7_, i_6_, n_n139, n_n281, x924x, x899x}, x20712x);
	defparam lut_7171.LUT_SIZE = 7;
	defparam lut_7171.mask = 128'h111fffff111fffff3337000500050005;

	lut_sub lut_7174 ({sk[1627], x917x, n_n283, n_n108, n_n4970, x103x, x20712x}, n_n4279);
	defparam lut_7174.LUT_SIZE = 7;
	defparam lut_7174.mask = 128'h111fffff111fffff5f5f5f5f5f5f7fff;

	lut_sub lut_7179 ({sk[1628], n_n273, n_n220, x922x, n_n60, x902x, x133x}, x20274x);
	defparam lut_7179.LUT_SIZE = 7;
	defparam lut_7179.mask = 128'h111fffff111fffff00000000005f007f;

	lut_sub lut_7183 ({sk[1629], n_n283, x922x, n_n228, x897x, x156x, x20274x}, n_n3978);
	defparam lut_7183.LUT_SIZE = 7;
	defparam lut_7183.mask = 128'h111fffff111fffff555555555555777f;

	lut_sub lut_7187 ({sk[1630], i_7_, i_8_, i_6_, x916x, x78x, n_n41}, n_n1346);
	defparam lut_7187.LUT_SIZE = 7;
	defparam lut_7187.mask = 128'h111fffff111fffff0005000300000000;

	lut_sub lut_7190 ({sk[1631], n_n208, x916x, n_n222, x88x, x902x}, n_n884);
	defparam lut_7190.LUT_SIZE = 6;
	defparam lut_7190.mask = 64'h7f7f7f7f00000037;

	lut_sub lut_7193 ({sk[1632], i_14_, i_13_, i_12_, i_15_, n_n247, x897x}, x1144x);
	defparam lut_7193.LUT_SIZE = 7;
	defparam lut_7193.mask = 128'h111fffff111fffff0333303333553330;

	lut_sub lut_7206 ({sk[1633], n_n208, x916x, n_n31, x466x, x141x, n_n1346}, x21228x);
	defparam lut_7206.LUT_SIZE = 7;
	defparam lut_7206.mask = 128'h111fffff111fffff5f5f5f5f5f5f7fff;

	lut_sub lut_7211 ({sk[1634], n_n4, n_n3, x88x, n_n7297, x181x, x1144x}, x21229x);
	defparam lut_7211.LUT_SIZE = 7;
	defparam lut_7211.mask = 128'h111fffff111fffff0f0f5f5f3fff7fff;

	lut_sub lut_7216 ({sk[1635], i_14_, i_13_, i_12_, x905x, x188x}, x1145x);
	defparam lut_7216.LUT_SIZE = 6;
	defparam lut_7216.mask = 64'h7f7f7f7f57755555;

	lut_sub lut_7220 ({sk[1636], x915x, n_n261, n_n263, x121x, n_n15, x1145x}, n_n3212);
	defparam lut_7220.LUT_SIZE = 7;
	defparam lut_7220.mask = 128'h111fffff111fffff0000000000553f7f;

	lut_sub lut_7224 ({sk[1637], i_7_, i_8_, i_6_, n_n220, x922x, x904x}, x741x);
	defparam lut_7224.LUT_SIZE = 7;
	defparam lut_7224.mask = 128'h111fffff111fffff0100000000000000;

	lut_sub lut_7226 ({sk[1638], n_n273, n_n220, n_n258, x922x, x908x, x902x}, x626x);
	defparam lut_7226.LUT_SIZE = 7;
	defparam lut_7226.mask = 128'h111fffff111fffff0000000000030507;

	lut_sub lut_7229 ({sk[1639], i_7_, i_8_, i_6_, x915x, x68x}, x591x);
	defparam lut_7229.LUT_SIZE = 6;
	defparam lut_7229.mask = 64'h7f7f7f7f00100000;

	lut_sub lut_7231 ({sk[1640], i_15_, n_n273, x922x, n_n270, n_n225, n_n6856}, x478x);
	defparam lut_7231.LUT_SIZE = 7;
	defparam lut_7231.mask = 128'h111fffff111fffff5555555755555555;

	lut_sub lut_7234 ({sk[1641], n_n273, n_n258, x922x, x899x, x902x, n_n256}, x20387x);
	defparam lut_7234.LUT_SIZE = 7;
	defparam lut_7234.mask = 128'h111fffff111fffff000000000011001f;

	lut_sub lut_7237 ({sk[1642], n_n6861, x4598x, x479x, x478x, x20387x}, x736x);
	defparam lut_7237.LUT_SIZE = 6;
	defparam lut_7237.mask = 64'h7f7f7f7f7fffffff;

	lut_sub lut_7243 ({sk[1643], n_n6878, x475x, x438x, x20386x, n_n6879, x591x}, x20392x);
	defparam lut_7243.LUT_SIZE = 7;
	defparam lut_7243.mask = 128'h111fffff111fffff7fffffffffffffff;

	lut_sub lut_7250 ({sk[1644], n_n281, n_n208, x916x, n_n220, x908x, x902x}, x20394x);
	defparam lut_7250.LUT_SIZE = 7;
	defparam lut_7250.mask = 128'h111fffff111fffff0000000500000037;

	lut_sub lut_7253 ({sk[1645], i_14_, i_13_, i_12_, n_n3, x898x}, x349x);
	defparam lut_7253.LUT_SIZE = 6;
	defparam lut_7253.mask = 64'h7f7f7f7f00000001;

	lut_sub lut_7255 ({sk[1646], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1914x);
	defparam lut_7255.LUT_SIZE = 7;
	defparam lut_7255.mask = 128'h111fffff111fffff0101000504000400;

	lut_sub lut_7262 ({sk[1647], i_14_, i_13_, i_12_, n_n273, x922x, x902x}, x20247x);
	defparam lut_7262.LUT_SIZE = 7;
	defparam lut_7262.mask = 128'h111fffff111fffff0000000000010100;

	lut_sub lut_7265 ({sk[1648], i_7_, i_8_, i_6_, x88x, x922x, x20247x}, x483x);
	defparam lut_7265.LUT_SIZE = 7;
	defparam lut_7265.mask = 128'h111fffff111fffff5555575555555555;

	lut_sub lut_7268 ({sk[1649], n_n273, n_n7441, x88x, x922x, x141x, x20247x}, x876x);
	defparam lut_7268.LUT_SIZE = 7;
	defparam lut_7268.mask = 128'h111fffff111fffff5555ffff575fffff;

	lut_sub lut_7273 ({sk[1650], n_n148, x206x, n_n48, n_n53, n_n15, x1192x}, x21004x);
	defparam lut_7273.LUT_SIZE = 7;
	defparam lut_7273.mask = 128'h111fffff111fffff00770f7f0f7f0f7f;

	lut_sub lut_7278 ({sk[1651], n_n48, n_n6511, n_n3184, x1909x, x21013x, x21014x}, n_n3123);
	defparam lut_7278.LUT_SIZE = 7;
	defparam lut_7278.mask = 128'h111fffff111fffff77ffffff7fffffff;

	lut_sub lut_7284 ({sk[1652], n_n273, n_n283, n_n108, x922x, x82x, x70x}, x21002x);
	defparam lut_7284.LUT_SIZE = 7;
	defparam lut_7284.mask = 128'h111fffff111fffff0000030f050f070f;

	lut_sub lut_7289 ({sk[1653], n_n273, n_n283, x922x, x44x, x463x, x1938x}, x21003x);
	defparam lut_7289.LUT_SIZE = 7;
	defparam lut_7289.mask = 128'h111fffff111fffff33333377333f337f;

	lut_sub lut_7293 ({sk[1654], x406x, x865x, x21058x, x24156x}, x21061x);
	defparam lut_7293.LUT_SIZE = 5;
	defparam lut_7293.mask = 32'h7f7fbfff;

	lut_sub lut_7298 ({sk[1655], n_n6, n_n5, x1918x, x1868x, x21032x, x21034x}, x21036x);
	defparam lut_7298.LUT_SIZE = 7;
	defparam lut_7298.mask = 128'h111fffff111fffff777777ff7f7f7fff;

	lut_sub lut_7303 ({sk[1656], n_n3180, x317x, x21019x, n_n2890, x21028x, x21027x}, x21037x);
	defparam lut_7303.LUT_SIZE = 7;
	defparam lut_7303.mask = 128'h111fffff111fffff7fffffffffffffff;

	lut_sub lut_7310 ({sk[1657], n_n273, x922x, x869x, x1881x, x1852x, x21052x}, x21054x);
	defparam lut_7310.LUT_SIZE = 7;
	defparam lut_7310.mask = 128'h111fffff111fffff55ff55ff55ff7fff;

	lut_sub lut_7315 ({sk[1658], x21039x, x21040x, x781x, x21044x, x21045x, x21046x}, x21055x);
	defparam lut_7315.LUT_SIZE = 7;
	defparam lut_7315.mask = 128'h111fffff111fffff7fffffffffffffff;

	lut_sub lut_7322 ({sk[1659], n_n266, n_n271, x909x, x106x, x1885x, x1902x}, x21119x);
	defparam lut_7322.LUT_SIZE = 7;
	defparam lut_7322.mask = 128'h111fffff111fffff00000033005f007f;

	lut_sub lut_7326 ({sk[1660], n_n56, x170x, n_n3204, x49x, x538x, x682x}, x24122x);
	defparam lut_7326.LUT_SIZE = 7;
	defparam lut_7326.mask = 128'h111fffff111fffff8800880080000000;

	lut_sub lut_7329 ({sk[1661], x21070x, x21071x, x21075x, x21119x, x24122x}, x21122x);
	defparam lut_7329.LUT_SIZE = 6;
	defparam lut_7329.mask = 64'h7f7f7f7fbfffffff;

	lut_sub lut_7335 ({sk[1662], n_n197, n_n94, n_n3212, x1910x, x701x, n_n2926}, x21095x);
	defparam lut_7335.LUT_SIZE = 7;
	defparam lut_7335.mask = 128'h111fffff111fffff77ff7fff77ffffff;

	lut_sub lut_7341 ({sk[1663], n_n54, n_n94, n_n3722, n_n3221, x1943x, x821x}, x21116x);
	defparam lut_7341.LUT_SIZE = 7;
	defparam lut_7341.mask = 128'h111fffff111fffff5fff7fff5fffffff;

	lut_sub lut_7347 ({sk[1664], n_n100, x21101x, x21102x, x383x, x1896x, x21106x}, x21117x);
	defparam lut_7347.LUT_SIZE = 7;
	defparam lut_7347.mask = 128'h111fffff111fffff5fffffff7fffffff;

	lut_sub lut_7353 ({sk[1665], n_n266, x909x, x204x, x370x, x21080x, x24161x}, n_n3132);
	defparam lut_7353.LUT_SIZE = 7;
	defparam lut_7353.mask = 128'h111fffff111fffffbfbfbfbfbfbfbfff;

	lut_sub lut_7358 ({sk[1666], x184x, n_n100, x654x, n_n3209, x21090x, x24165x}, n_n3133);
	defparam lut_7358.LUT_SIZE = 7;
	defparam lut_7358.mask = 128'h111fffff111fffffbfffbfffbfffffff;

	lut_sub lut_7364 ({sk[1667], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1926x);
	defparam lut_7364.LUT_SIZE = 7;
	defparam lut_7364.mask = 128'h111fffff111fffff0000001050005040;

	lut_sub lut_7371 ({sk[1668], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1146x);
	defparam lut_7371.LUT_SIZE = 7;
	defparam lut_7371.mask = 128'h111fffff111fffff4000100000040001;

	lut_sub lut_7376 ({sk[1669], i_14_, i_13_, i_12_, i_15_, x907x, n_n282}, x290x);
	defparam lut_7376.LUT_SIZE = 7;
	defparam lut_7376.mask = 128'h111fffff111fffff5000050000330000;

	lut_sub lut_7380 ({sk[1670], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1147x);
	defparam lut_7380.LUT_SIZE = 7;
	defparam lut_7380.mask = 128'h111fffff111fffff4000100000440001;

	lut_sub lut_7386 ({sk[1671], i_14_, i_13_, i_12_, i_15_, n_n275, x209x}, x1588x);
	defparam lut_7386.LUT_SIZE = 7;
	defparam lut_7386.mask = 128'h111fffff111fffff5555555555755557;

	lut_sub lut_7390 ({sk[1672], x915x, n_n7, n_n261, n_n263, x133x, x1588x}, n_n2676);
	defparam lut_7390.LUT_SIZE = 7;
	defparam lut_7390.mask = 128'h111fffff111fffff0000000003570f5f;

	lut_sub lut_7394 ({sk[1673], i_14_, i_13_, i_12_, x907x, x915x, n_n261}, x528x);
	defparam lut_7394.LUT_SIZE = 7;
	defparam lut_7394.mask = 128'h111fffff111fffff0100000000000000;

	lut_sub lut_7396 ({sk[1674], i_7_, i_8_, i_6_, n_n106, x915x, x160x}, n_n2702);
	defparam lut_7396.LUT_SIZE = 7;
	defparam lut_7396.mask = 128'h111fffff111fffff0000000011000300;

	lut_sub lut_7399 ({sk[1675], i_7_, i_8_, i_6_, x915x, x901x, n_n228}, x601x);
	defparam lut_7399.LUT_SIZE = 7;
	defparam lut_7399.mask = 128'h111fffff111fffff0000000000000100;

	lut_sub lut_7401 ({sk[1676], n_n281, x915x, n_n220, x914x, n_n263, x912x}, x654x);
	defparam lut_7401.LUT_SIZE = 7;
	defparam lut_7401.mask = 128'h111fffff111fffff0000001100000313;

	lut_sub lut_7404 ({sk[1677], n_n9, x314x, n_n100, n_n2702, x654x, x132x}, x20041x);
	defparam lut_7404.LUT_SIZE = 7;
	defparam lut_7404.mask = 128'h111fffff111fffff3f7f3fff3fff3fff;

	lut_sub lut_7410 ({sk[1678], i_14_, i_13_, i_12_, x913x, x915x, n_n263}, n_n2398);
	defparam lut_7410.LUT_SIZE = 7;
	defparam lut_7410.mask = 128'h111fffff111fffff0001010100000000;

	lut_sub lut_7414 ({sk[1679], i_14_, i_13_, i_12_, i_15_, x899x, n_n259}, x227x);
	defparam lut_7414.LUT_SIZE = 7;
	defparam lut_7414.mask = 128'h111fffff111fffff0000000005333300;

	lut_sub lut_7418 ({sk[1680], i_14_, i_13_, i_12_, x905x, x899x, x42x}, x1151x);
	defparam lut_7418.LUT_SIZE = 7;
	defparam lut_7418.mask = 128'h111fffff111fffff777755777f777755;

	lut_sub lut_7427 ({sk[1681], i_14_, i_13_, i_12_, i_15_, n_n242, x217x}, x1150x);
	defparam lut_7427.LUT_SIZE = 7;
	defparam lut_7427.mask = 128'h111fffff111fffff5777757755555555;

	lut_sub lut_7435 ({sk[1682], i_14_, i_13_, i_12_, x915x, x911x, n_n263}, x20045x);
	defparam lut_7435.LUT_SIZE = 7;
	defparam lut_7435.mask = 128'h111fffff111fffff0101000100000000;

	lut_sub lut_7439 ({sk[1683], x915x, n_n261, x142x, n_n2398, x20045x}, x20047x);
	defparam lut_7439.LUT_SIZE = 6;
	defparam lut_7439.mask = 64'h7f7f7f7f7777777f;

	lut_sub lut_7443 ({sk[1684], i_7_, i_8_, i_6_, x915x, x1151x, x1150x}, x20048x);
	defparam lut_7443.LUT_SIZE = 7;
	defparam lut_7443.mask = 128'h111fffff111fffff0000000003000500;

	lut_sub lut_7446 ({sk[1685], i_14_, i_13_, i_12_, x915x, n_n263, x904x}, x4847x);
	defparam lut_7446.LUT_SIZE = 7;
	defparam lut_7446.mask = 128'h111fffff111fffff0100000000000000;

	lut_sub lut_7448 ({sk[1686], i_14_, i_13_, i_12_, x901x, x900x, x906x}, x20050x);
	defparam lut_7448.LUT_SIZE = 7;
	defparam lut_7448.mask = 128'h111fffff111fffff000000000055003f;

	lut_sub lut_7452 ({sk[1687], i_14_, i_13_, i_12_, x907x, x905x, x113x}, x20051x);
	defparam lut_7452.LUT_SIZE = 7;
	defparam lut_7452.mask = 128'h111fffff111fffff55777777555f5555;

	lut_sub lut_7458 ({sk[1688], i_14_, i_13_, i_12_, i_15_, x184x, n_n253}, x1152x);
	defparam lut_7458.LUT_SIZE = 7;
	defparam lut_7458.mask = 128'h111fffff111fffff7333373333733337;

	lut_sub lut_7464 ({sk[1689], n_n100, n_n94, x20050x, x20051x, x1763x, x1762x}, x20053x);
	defparam lut_7464.LUT_SIZE = 7;
	defparam lut_7464.mask = 128'h111fffff111fffff00003fff55557fff;

	lut_sub lut_7469 ({sk[1690], n_n228, x902x, n_n94, x209x, x645x, x601x}, x20040x);
	defparam lut_7469.LUT_SIZE = 7;
	defparam lut_7469.mask = 128'h111fffff111fffff777f777f777f77ff;

	lut_sub lut_7474 ({sk[1691], i_9_, i_10_, i_11_, i_15_, n_n279, n_n225}, x1157x);
	defparam lut_7474.LUT_SIZE = 7;
	defparam lut_7474.mask = 128'h111fffff111fffff0053300000000000;

	lut_sub lut_7478 ({sk[1692], n_n208, x909x, n_n145, n_n263, x700x, x1157x}, x21539x);
	defparam lut_7478.LUT_SIZE = 7;
	defparam lut_7478.mask = 128'h111fffff111fffff3333333f3333777f;

	lut_sub lut_7482 ({sk[1693], n_n151, x164x, n_n77, n_n227, n_n30, x21539x}, n_n2133);
	defparam lut_7482.LUT_SIZE = 7;
	defparam lut_7482.mask = 128'h111fffff111fffff575f575f575fffff;

	lut_sub lut_7487 ({sk[1694], i_14_, i_13_, i_12_, x913x, x911x, n_n94}, x388x);
	defparam lut_7487.LUT_SIZE = 7;
	defparam lut_7487.mask = 128'h111fffff111fffff1100000500000000;

	lut_sub lut_7490 ({sk[1695], i_14_, i_13_, i_12_, x903x, x897x}, x257x);
	defparam lut_7490.LUT_SIZE = 6;
	defparam lut_7490.mask = 64'h7f7f7f7f53300000;

	lut_sub lut_7494 ({sk[1696], x911x, x905x, n_n279, n_n94, n_n227, x257x}, x21543x);
	defparam lut_7494.LUT_SIZE = 7;
	defparam lut_7494.mask = 128'h111fffff111fffff05050537050f053f;

	lut_sub lut_7498 ({sk[1697], i_14_, i_13_, i_12_, x915x, n_n261, x901x}, x382x);
	defparam lut_7498.LUT_SIZE = 7;
	defparam lut_7498.mask = 128'h111fffff111fffff0000000001000000;

	lut_sub lut_7500 ({sk[1698], i_7_, i_8_, i_6_, x907x, x915x, n_n225}, x892x);
	defparam lut_7500.LUT_SIZE = 7;
	defparam lut_7500.mask = 128'h111fffff111fffff0000000000000100;

	lut_sub lut_7502 ({sk[1699], i_14_, i_13_, i_12_, x907x, x915x, n_n261}, x391x);
	defparam lut_7502.LUT_SIZE = 7;
	defparam lut_7502.mask = 128'h111fffff111fffff0001000100000000;

	lut_sub lut_7505 ({sk[1700], n_n151, n_n7, n_n100, n_n35, n_n94, x382x}, x24107x);
	defparam lut_7505.LUT_SIZE = 7;
	defparam lut_7505.mask = 128'h111fffff111fffffaaa0888088808880;

	lut_sub lut_7510 ({sk[1701], n_n4, n_n30, n_n6823, x528x, x391x, x24107x}, x21549x);
	defparam lut_7510.LUT_SIZE = 7;
	defparam lut_7510.mask = 128'h111fffff111fffffbfffbfffbfffffff;

	lut_sub lut_7516 ({sk[1702], x685x, n_n6813, n_n2133, x388x, x21543x, x21549x}, n_n2080);
	defparam lut_7516.LUT_SIZE = 7;
	defparam lut_7516.mask = 128'h111fffff111fffff7fffffffffffffff;

	lut_sub lut_7523 ({sk[1703], i_14_, i_13_, i_12_, i_15_, n_n247, n_n267}, x1159x);
	defparam lut_7523.LUT_SIZE = 7;
	defparam lut_7523.mask = 128'h111fffff111fffff0770707077000000;

	lut_sub lut_7536 ({sk[1704], i_14_, i_13_, i_12_, x904x, x906x}, x21422x);
	defparam lut_7536.LUT_SIZE = 6;
	defparam lut_7536.mask = 64'h7f7f7f7f07770000;

	lut_sub lut_7543 ({sk[1705], i_9_, i_10_, i_11_, i_15_, n_n281, n_n279}, x24109x);
	defparam lut_7543.LUT_SIZE = 7;
	defparam lut_7543.mask = 128'h111fffff111fffffa8ffffa8ffffffa8;

	lut_sub lut_7550 ({sk[1706], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x253x);
	defparam lut_7550.LUT_SIZE = 7;
	defparam lut_7550.mask = 128'h111fffff111fffff0100000404000000;

	lut_sub lut_7554 ({sk[1707], i_14_, i_13_, i_12_, n_n273, x922x, x908x}, n_n2274);
	defparam lut_7554.LUT_SIZE = 7;
	defparam lut_7554.mask = 128'h111fffff111fffff0001010100000000;

	lut_sub lut_7558 ({sk[1708], i_9_, i_10_, i_11_, i_15_, n_n279}, x369x);
	defparam lut_7558.LUT_SIZE = 6;
	defparam lut_7558.mask = 64'h7f7f7f7f00000500;

	lut_sub lut_7561 ({sk[1709], i_14_, i_13_, i_12_, x898x, x904x}, x1162x);
	defparam lut_7561.LUT_SIZE = 6;
	defparam lut_7561.mask = 64'h7f7f7f7f35557000;

	lut_sub lut_7568 ({sk[1710], i_14_, i_13_, i_12_, x903x, x897x}, x1165x);
	defparam lut_7568.LUT_SIZE = 6;
	defparam lut_7568.mask = 64'h7f7f7f7f00050053;

	lut_sub lut_7572 ({sk[1711], i_14_, i_13_, i_12_, i_15_, x911x, n_n259}, x1164x);
	defparam lut_7572.LUT_SIZE = 7;
	defparam lut_7572.mask = 128'h111fffff111fffff0000370000500000;

	lut_sub lut_7576 ({sk[1712], i_7_, i_8_, i_6_, x909x, x75x}, x2782x);
	defparam lut_7576.LUT_SIZE = 6;
	defparam lut_7576.mask = 64'h7f7f7f7f00000010;

	lut_sub lut_7578 ({sk[1713], n_n5, n_n103, n_n207, x1165x, x1164x, x2782x}, n_n1217);
	defparam lut_7578.LUT_SIZE = 7;
	defparam lut_7578.mask = 128'h111fffff111fffff555f55ff777f77ff;

	lut_sub lut_7583 ({sk[1714], i_7_, i_8_, i_6_, x915x, x223x}, x2589x);
	defparam lut_7583.LUT_SIZE = 6;
	defparam lut_7583.mask = 64'h7f7f7f7f00001000;

	lut_sub lut_7585 ({sk[1715], i_14_, i_13_, i_12_, x913x, x63x}, x1166x);
	defparam lut_7585.LUT_SIZE = 6;
	defparam lut_7585.mask = 64'h7f7f7f7f55555755;

	lut_sub lut_7588 ({sk[1716], i_14_, i_13_, i_12_, i_15_, n_n282, n_n253}, x1170x);
	defparam lut_7588.LUT_SIZE = 7;
	defparam lut_7588.mask = 128'h111fffff111fffff0777300330003330;

	lut_sub lut_7601 ({sk[1717], i_14_, i_13_, i_12_, i_15_, x907x, n_n247}, x1169x);
	defparam lut_7601.LUT_SIZE = 7;
	defparam lut_7601.mask = 128'h111fffff111fffff0505000550005073;

	lut_sub lut_7609 ({sk[1718], n_n53, x67x, x623x, x516x, x55x, x741x}, x22294x);
	defparam lut_7609.LUT_SIZE = 7;
	defparam lut_7609.mask = 128'h111fffff111fffff5fff5fff7fffffff;

	lut_sub lut_7615 ({sk[1719], i_7_, i_8_, i_6_, x922x, x1170x, x1169x}, x22295x);
	defparam lut_7615.LUT_SIZE = 7;
	defparam lut_7615.mask = 128'h111fffff111fffff0300050000000000;

	lut_sub lut_7618 ({sk[1720], i_14_, i_13_, i_12_, x907x, x64x, x901x}, x1925x);
	defparam lut_7618.LUT_SIZE = 7;
	defparam lut_7618.mask = 128'h111fffff111fffff773333333f333f3f;

	lut_sub lut_7624 ({sk[1721], x915x, n_n283, x85x, n_n6879, x1925x}, n_n1204);
	defparam lut_7624.LUT_SIZE = 6;
	defparam lut_7624.mask = 64'h7f7f7f7f3333337f;

	lut_sub lut_7628 ({sk[1722], n_n273, x905x, n_n279, x922x, x899x, n_n225}, x4509x);
	defparam lut_7628.LUT_SIZE = 7;
	defparam lut_7628.mask = 128'h111fffff111fffff000000000101010f;

	lut_sub lut_7631 ({sk[1723], i_14_, i_13_, i_12_, x907x, x915x, n_n283}, x2761x);
	defparam lut_7631.LUT_SIZE = 7;
	defparam lut_7631.mask = 128'h111fffff111fffff0001010000010000;

	lut_sub lut_7635 ({sk[1724], i_14_, i_13_, i_12_, n_n273, x922x, x899x}, x22035x);
	defparam lut_7635.LUT_SIZE = 7;
	defparam lut_7635.mask = 128'h111fffff111fffff0100010000000000;

	lut_sub lut_7638 ({sk[1725], n_n1, n_n6867, x41x, x4509x, x2761x, x22035x}, x22041x);
	defparam lut_7638.LUT_SIZE = 7;
	defparam lut_7638.mask = 128'h111fffff111fffff7f7fffff7fffffff;

	lut_sub lut_7644 ({sk[1726], i_7_, i_8_, i_6_, x909x, x62x}, x4708x);
	defparam lut_7644.LUT_SIZE = 6;
	defparam lut_7644.mask = 64'h7f7f7f7f00000010;

	lut_sub lut_7646 ({sk[1727], i_14_, i_13_, i_12_, i_15_, x911x, n_n253}, x22028x);
	defparam lut_7646.LUT_SIZE = 7;
	defparam lut_7646.mask = 128'h111fffff111fffff3333053300500000;

	lut_sub lut_7652 ({sk[1728], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x220x);
	defparam lut_7652.LUT_SIZE = 7;
	defparam lut_7652.mask = 128'h111fffff111fffff0000010000040000;

	lut_sub lut_7655 ({sk[1729], i_14_, i_13_, i_12_, x900x, x906x, x220x}, x22025x);
	defparam lut_7655.LUT_SIZE = 7;
	defparam lut_7655.mask = 128'h111fffff111fffff55555f5555775555;

	lut_sub lut_7659 ({sk[1730], i_14_, i_13_, i_12_, i_15_, x905x, n_n259}, x22026x);
	defparam lut_7659.LUT_SIZE = 7;
	defparam lut_7659.mask = 128'h111fffff111fffff0533500000005550;

	lut_sub lut_7666 ({sk[1731], x909x, n_n261, n_n246, x142x, x73x, x22028x}, x2777x);
	defparam lut_7666.LUT_SIZE = 7;
	defparam lut_7666.mask = 128'h111fffff111fffff0000000000007fff;

	lut_sub lut_7671 ({sk[1732], n_n5, n_n197, x125x, x4708x, x22025x, x22026x}, x22031x);
	defparam lut_7671.LUT_SIZE = 7;
	defparam lut_7671.mask = 128'h111fffff111fffff0f0f0f0f7fffffff;

	lut_sub lut_7677 ({sk[1733], i_14_, i_13_, i_12_, n_n266, x909x, x905x}, x481x);
	defparam lut_7677.LUT_SIZE = 7;
	defparam lut_7677.mask = 128'h111fffff111fffff0001010000000000;

	lut_sub lut_7680 ({sk[1734], n_n57, x125x, x60x, x783x, n_n4394, x481x}, x22270x);
	defparam lut_7680.LUT_SIZE = 7;
	defparam lut_7680.mask = 128'h111fffff111fffff7f7f7f7f7fffffff;

	lut_sub lut_7686 ({sk[1735], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1336x);
	defparam lut_7686.LUT_SIZE = 7;
	defparam lut_7686.mask = 128'h111fffff111fffff1050001040105040;

	lut_sub lut_7696 ({sk[1736], i_14_, i_13_, i_12_, i_15_, x899x, n_n242}, x1335x);
	defparam lut_7696.LUT_SIZE = 7;
	defparam lut_7696.mask = 128'h111fffff111fffff3300000050005050;

	lut_sub lut_7701 ({sk[1737], n_n197, n_n57, n_n56, x62x, x1336x, x1335x}, x22271x);
	defparam lut_7701.LUT_SIZE = 7;
	defparam lut_7701.mask = 128'h111fffff111fffff00335f7f00ff5fff;

	lut_sub lut_7706 ({sk[1738], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x22275x);
	defparam lut_7706.LUT_SIZE = 7;
	defparam lut_7706.mask = 128'h111fffff111fffff0010001040005040;

	lut_sub lut_7713 ({sk[1739], n_n271, x909x, x355x, x22275x, x22274x}, x2521x);
	defparam lut_7713.LUT_SIZE = 6;
	defparam lut_7713.mask = 64'h7f7f7f7f0000007f;

	lut_sub lut_7717 ({sk[1740], n_n57, n_n56, n_n246, n_n147, x291x, x24090x}, x22277x);
	defparam lut_7717.LUT_SIZE = 7;
	defparam lut_7717.mask = 128'h111fffff111fffff00003fffaaaabfff;

	lut_sub lut_7722 ({sk[1741], x22264x, x22265x, x22270x, x22271x, x2521x, x22277x}, n_n1099);
	defparam lut_7722.LUT_SIZE = 7;
	defparam lut_7722.mask = 128'h111fffff111fffff7fffffffffffffff;

	lut_sub lut_7729 ({sk[1742], i_7_, i_8_, i_6_, n_n220, x922x, x904x}, x5574x);
	defparam lut_7729.LUT_SIZE = 7;
	defparam lut_7729.mask = 128'h111fffff111fffff0000010000000000;

	lut_sub lut_7731 ({sk[1743], i_14_, i_13_, i_12_, x900x, x906x}, x43x);
	defparam lut_7731.LUT_SIZE = 6;
	defparam lut_7731.mask = 64'h7f7f7f7f03035000;

	lut_sub lut_7735 ({sk[1744], i_14_, i_13_, i_12_, i_15_, n_n253, n_n267}, x1177x);
	defparam lut_7735.LUT_SIZE = 7;
	defparam lut_7735.mask = 128'h111fffff111fffff0505000770037370;

	lut_sub lut_7748 ({sk[1745], i_14_, i_13_, i_12_, i_15_, n_n267}, x416x);
	defparam lut_7748.LUT_SIZE = 6;
	defparam lut_7748.mask = 64'h7f7f7f7f14400000;

	lut_sub lut_7752 ({sk[1746], n_n48, x912x, n_n225, x189x, x479x, x656x}, x22286x);
	defparam lut_7752.LUT_SIZE = 7;
	defparam lut_7752.mask = 128'h111fffff111fffff777777777f7f7fff;

	lut_sub lut_7757 ({sk[1747], n_n1255, x22287x, x22294x, x22295x, x22286x}, x22303x);
	defparam lut_7757.LUT_SIZE = 6;
	defparam lut_7757.mask = 64'h7f7f7f7f7fffffff;

	lut_sub lut_7763 ({sk[1748], i_7_, i_8_, i_6_, x78x, x909x}, x3598x);
	defparam lut_7763.LUT_SIZE = 6;
	defparam lut_7763.mask = 64'h7f7f7f7f00000100;

	lut_sub lut_7765 ({sk[1749], i_14_, i_13_, i_12_, n_n266, x909x, x901x}, x3599x);
	defparam lut_7765.LUT_SIZE = 7;
	defparam lut_7765.mask = 128'h111fffff111fffff0000000000010000;

	lut_sub lut_7767 ({sk[1750], i_7_, i_8_, i_6_, x909x, x85x}, x4663x);
	defparam lut_7767.LUT_SIZE = 6;
	defparam lut_7767.mask = 64'h7f7f7f7f00000100;

	lut_sub lut_7769 ({sk[1751], i_7_, i_8_, i_6_, x909x, x112x}, x5284x);
	defparam lut_7769.LUT_SIZE = 6;
	defparam lut_7769.mask = 64'h7f7f7f7f00000100;

	lut_sub lut_7771 ({sk[1752], n_n4948, x538x, x3598x, x3599x, x4663x, x5284x}, x22308x);
	defparam lut_7771.LUT_SIZE = 7;
	defparam lut_7771.mask = 128'h111fffff111fffff7fffffffffffffff;

	lut_sub lut_7778 ({sk[1753], i_14_, i_13_, i_12_, n_n266, x909x, x908x}, x3569x);
	defparam lut_7778.LUT_SIZE = 7;
	defparam lut_7778.mask = 128'h111fffff111fffff0001010000000000;

	lut_sub lut_7781 ({sk[1754], n_n103, n_n57, n_n56, x49x, x165x, x140x}, x24212x);
	defparam lut_7781.LUT_SIZE = 7;
	defparam lut_7781.mask = 128'h111fffff111fffffffff8080ff008000;

	lut_sub lut_7786 ({sk[1755], n_n271, n_n220, x914x, x909x, x3569x, x24212x}, x22314x);
	defparam lut_7786.LUT_SIZE = 7;
	defparam lut_7786.mask = 128'h111fffff111fffffbbbbbbbbbbbbbbbf;

	lut_sub lut_7790 ({sk[1756], i_14_, i_13_, i_12_, n_n271, x909x, x908x}, x3567x);
	defparam lut_7790.LUT_SIZE = 7;
	defparam lut_7790.mask = 128'h111fffff111fffff0001010000000000;

	lut_sub lut_7793 ({sk[1757], i_14_, i_13_, i_12_, i_15_, n_n275, n_n259}, x1179x);
	defparam lut_7793.LUT_SIZE = 7;
	defparam lut_7793.mask = 128'h111fffff111fffff0333000330037770;

	lut_sub lut_7806 ({sk[1758], i_14_, i_13_, i_12_, x908x, x903x, x897x}, x1178x);
	defparam lut_7806.LUT_SIZE = 7;
	defparam lut_7806.mask = 128'h111fffff111fffff553333000f000f0f;

	lut_sub lut_7813 ({sk[1759], n_n266, n_n271, x909x, n_n22, x49x, x1178x}, x22319x);
	defparam lut_7813.LUT_SIZE = 7;
	defparam lut_7813.mask = 128'h111fffff111fffff00000077000f007f;

	lut_sub lut_7817 ({sk[1760], n_n197, n_n57, n_n56, x165x, x3567x, x1179x}, x22320x);
	defparam lut_7817.LUT_SIZE = 7;
	defparam lut_7817.mask = 128'h111fffff111fffff333f777f333fffff;

	lut_sub lut_7822 ({sk[1761], i_7_, i_8_, i_6_, x909x, x1513x, x1516x}, x24088x);
	defparam lut_7822.LUT_SIZE = 7;
	defparam lut_7822.mask = 128'h111fffff111ffffffffffffffffafffc;

	lut_sub lut_7829 ({sk[1762], x22308x, x22314x, x22319x, x22320x, x24088x}, n_n1100);
	defparam lut_7829.LUT_SIZE = 6;
	defparam lut_7829.mask = 64'h7f7f7f7fbfffffff;

	lut_sub lut_7835 ({sk[1763], i_14_, i_13_, i_12_, n_n273, x922x, x899x}, x406x);
	defparam lut_7835.LUT_SIZE = 7;
	defparam lut_7835.mask = 128'h111fffff111fffff0000000000010100;

	lut_sub lut_7838 ({sk[1764], i_14_, i_13_, i_12_, n_n273, x922x, x899x}, n_n952);
	defparam lut_7838.LUT_SIZE = 7;
	defparam lut_7838.mask = 128'h111fffff111fffff0000000001010100;

	lut_sub lut_7842 ({sk[1765], n_n6, n_n5, n_n104, n_n41, x126x, x177x}, n_n819);
	defparam lut_7842.LUT_SIZE = 7;
	defparam lut_7842.mask = 128'h111fffff111fffff00003f3f77ff7fff;

	lut_sub lut_7848 ({sk[1766], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x6020x);
	defparam lut_7848.LUT_SIZE = 7;
	defparam lut_7848.mask = 128'h111fffff111fffff5000000000000000;

	lut_sub lut_7851 ({sk[1767], i_9_, i_10_, i_11_, i_15_, n_n258, x6020x}, x19272x);
	defparam lut_7851.LUT_SIZE = 7;
	defparam lut_7851.mask = 128'h111fffff111fffff557555ff55555555;

	lut_sub lut_7855 ({sk[1768], i_14_, i_13_, i_12_, i_15_, n_n242, x903x}, x19273x);
	defparam lut_7855.LUT_SIZE = 7;
	defparam lut_7855.mask = 128'h111fffff111fffff3300330055005700;

	lut_sub lut_7861 ({sk[1769], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19276x);
	defparam lut_7861.LUT_SIZE = 7;
	defparam lut_7861.mask = 128'h111fffff111fffff000000000000ea2a;

	lut_sub lut_7866 ({sk[1770], i_9_, i_10_, i_11_, n_n208, x909x, n_n254}, x6008x);
	defparam lut_7866.LUT_SIZE = 7;
	defparam lut_7866.mask = 128'h111fffff111fffff0000000003020000;

	lut_sub lut_7869 ({sk[1771], n_n189, x898x, n_n279, x899x, x19276x, x6008x}, x19277x);
	defparam lut_7869.LUT_SIZE = 7;
	defparam lut_7869.mask = 128'h111fffff111fffff55555555777f77ff;

	lut_sub lut_7874 ({sk[1772], n_n208, x909x, x19267x, x19268x, x19272x, x19273x}, x19278x);
	defparam lut_7874.LUT_SIZE = 7;
	defparam lut_7874.mask = 128'h111fffff111fffff0000000000007fff;

	lut_sub lut_7879 ({sk[1773], i_9_, i_10_, i_11_}, x328x);
	defparam lut_7879.LUT_SIZE = 4;
	defparam lut_7879.mask = 16'h3307;

	lut_sub lut_7882 ({sk[1774], i_9_, i_10_, i_11_, n_n266, x916x, n_n271}, x19226x);
	defparam lut_7882.LUT_SIZE = 7;
	defparam lut_7882.mask = 128'h0f0fffffffffffff1103031303131313;

	lut_sub lut_7890 ({sk[1775], i_9_, i_7_, i_8_, i_6_, x922x}, x24145x);
	defparam lut_7890.LUT_SIZE = 6;
	defparam lut_7890.mask = 64'h555fffffeeaeeeea;

	lut_sub lut_7897 ({sk[1776], x916x, x1011x, x5909x, x19226x, x24145x}, x19230x);
	defparam lut_7897.LUT_SIZE = 6;
	defparam lut_7897.mask = 64'h555fffffbfbfbfff;

	lut_sub lut_7902 ({sk[1777], i_14_, i_13_, i_12_, n_n266, x909x, x902x}, n_n4938);
	defparam lut_7902.LUT_SIZE = 7;
	defparam lut_7902.mask = 128'h0f0fffffffffffff0000000001010100;

	lut_sub lut_7906 ({sk[1778], i_14_, i_13_, i_12_, x908x}, x167x);
	defparam lut_7906.LUT_SIZE = 5;
	defparam lut_7906.mask = 32'h0fff1500;

	lut_sub lut_7910 ({sk[1779], i_7_, i_8_, i_6_, x909x, x167x}, x5000x);
	defparam lut_7910.LUT_SIZE = 6;
	defparam lut_7910.mask = 64'h555fffff00000001;

	lut_sub lut_7912 ({sk[1780], i_14_, i_13_, i_12_, x903x}, x119x);
	defparam lut_7912.LUT_SIZE = 5;
	defparam lut_7912.mask = 32'h3f3f1500;

	lut_sub lut_7916 ({sk[1781], i_7_, i_8_, i_6_, x909x, n_n4930, x119x}, x761x);
	defparam lut_7916.LUT_SIZE = 7;
	defparam lut_7916.mask = 128'h33ffffff33ffffff3333333333373333;

	lut_sub lut_7919 ({sk[1782], n_n266, x909x, x165x, x140x, x761x}, x19930x);
	defparam lut_7919.LUT_SIZE = 6;
	defparam lut_7919.mask = 64'h77ff77ff5555557f;

	lut_sub lut_7923 ({sk[1783], n_n56, x124x, x212x, x190x, n_n4938, x5000x}, x19931x);
	defparam lut_7923.LUT_SIZE = 7;
	defparam lut_7923.mask = 128'h33ffffff33ffffff777777777fffffff;

	lut_sub lut_7929 ({sk[1784], i_7_, i_8_, i_6_, x909x, x119x}, x763x);
	defparam lut_7929.LUT_SIZE = 6;
	defparam lut_7929.mask = 64'h77ff77ff00000001;

	lut_sub lut_7931 ({sk[1785], n_n266, n_n271, x909x, x124x, x212x, n_n4930}, x20698x);
	defparam lut_7931.LUT_SIZE = 7;
	defparam lut_7931.mask = 128'h33ffffff33ffffff5555557f5577557f;

	lut_sub lut_7936 ({sk[1786], n_n273, n_n258, x898x, x922x, x579x, x764x}, n_n4183);
	defparam lut_7936.LUT_SIZE = 7;
	defparam lut_7936.mask = 128'h33ffffff33ffffff777777777777777f;

	lut_sub lut_7940 ({sk[1787], i_14_, i_13_, i_12_, i_15_, x898x, n_n267}, x1190x);
	defparam lut_7940.LUT_SIZE = 7;
	defparam lut_7940.mask = 128'h33ffffff33ffffff5000050000500037;

	lut_sub lut_7946 ({sk[1788], i_14_, i_13_, i_12_, i_15_, n_n267, x246x}, x1189x);
	defparam lut_7946.LUT_SIZE = 7;
	defparam lut_7946.mask = 128'h33ffffff33ffffff7555575555555555;

	lut_sub lut_7950 ({sk[1789], i_7_, i_8_, i_6_, x915x, x1190x, x1189x}, n_n3481);
	defparam lut_7950.LUT_SIZE = 7;
	defparam lut_7950.mask = 128'h33ffffff33ffffff0000000003000500;

	lut_sub lut_7953 ({sk[1790], i_7_, i_8_, i_6_, x206x, x922x}, n_n4160);
	defparam lut_7953.LUT_SIZE = 6;
	defparam lut_7953.mask = 64'h77ff77ff00100000;

	lut_sub lut_7955 ({sk[1791], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x1886x);
	defparam lut_7955.LUT_SIZE = 7;
	defparam lut_7955.mask = 128'h33ffffff33ffffff1050405040004000;

	lut_sub lut_7964 ({sk[1792], i_14_, i_13_, i_12_, i_15_, n_n247, x368x}, x1929x);
	defparam lut_7964.LUT_SIZE = 7;
	defparam lut_7964.mask = 128'h33ffffff33ffffff5555555555575755;

	lut_sub lut_7968 ({sk[1793], i_7_, i_8_, i_6_, x915x, x77x}, x768x);
	defparam lut_7968.LUT_SIZE = 6;
	defparam lut_7968.mask = 64'h77ff77ff00001000;

	lut_sub lut_7970 ({sk[1794], i_14_, i_13_, i_12_, i_15_, n_n247, n_n253}, x1191x);
	defparam lut_7970.LUT_SIZE = 7;
	defparam lut_7970.mask = 128'h33ffffff33ffffff0705007000000000;

	lut_sub lut_7976 ({sk[1795], n_n88, n_n94, x368x, n_n6834, x3786x, x1191x}, x21101x);
	defparam lut_7976.LUT_SIZE = 7;
	defparam lut_7976.mask = 128'h33ffffff33ffffff3f3f7fff3f3fffff;

	lut_sub lut_7982 ({sk[1796], n_n100, n_n6835, n_n6830, x1886x, x1929x, x768x}, x21102x);
	defparam lut_7982.LUT_SIZE = 7;
	defparam lut_7982.mask = 128'h33ffffff33ffffff55ffffff7fffffff;

	lut_sub lut_7988 ({sk[1797], i_15_, n_n283, x922x, n_n247, n_n246, n_n228}, x463x);
	defparam lut_7988.LUT_SIZE = 7;
	defparam lut_7988.mask = 128'h33ffffff33ffffff0000003300000037;

	lut_sub lut_7991 ({sk[1798], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1938x);
	defparam lut_7991.LUT_SIZE = 7;
	defparam lut_7991.mask = 128'h33ffffff33ffffff0010001050004040;

	lut_sub lut_7998 ({sk[1799], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1192x);
	defparam lut_7998.LUT_SIZE = 7;
	defparam lut_7998.mask = 128'h33ffffff33ffffff1440014000040000;

	lut_sub lut_8005 ({sk[1800], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x1909x);
	defparam lut_8005.LUT_SIZE = 7;
	defparam lut_8005.mask = 128'h33ffffff33ffffff0000001050004040;

	lut_sub lut_8011 ({sk[1801], n_n273, x922x, n_n60, x373x, n_n6521, x626x}, x21013x);
	defparam lut_8011.LUT_SIZE = 7;
	defparam lut_8011.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_8016 ({sk[1802], n_n41, x146x, n_n48, x457x, n_n6505, n_n6878}, x21014x);
	defparam lut_8016.LUT_SIZE = 7;
	defparam lut_8016.mask = 128'h33ffffff33ffffff7f7f7fff7fff7fff;

	lut_sub lut_8022 ({sk[1803], i_14_, i_13_, i_12_, i_15_, x902x, n_n270}, x1868x);
	defparam lut_8022.LUT_SIZE = 7;
	defparam lut_8022.mask = 128'h33ffffff33ffffff0000000005053350;

	lut_sub lut_8027 ({sk[1804], x909x, n_n261, n_n263, x67x, x593x, x181x}, x21032x);
	defparam lut_8027.LUT_SIZE = 7;
	defparam lut_8027.mask = 128'h33ffffff33ffffff33333333333f777f;

	lut_sub lut_8031 ({sk[1805], n_n6, n_n5, n_n197, x4716x, x141x, x181x}, x21034x);
	defparam lut_8031.LUT_SIZE = 7;
	defparam lut_8031.mask = 128'h33ffffff33ffffff0f0f7f7f3fff7fff;

	lut_sub lut_8037 ({sk[1806], n_n41, x909x, x115x, n_n263, x213x, x222x}, x21019x);
	defparam lut_8037.LUT_SIZE = 7;
	defparam lut_8037.mask = 128'h33ffffff33ffffff0000070f00000f0f;

	lut_sub lut_8042 ({sk[1807], i_7_, i_8_, i_6_, x909x, x174x, x1905x}, n_n2890);
	defparam lut_8042.LUT_SIZE = 7;
	defparam lut_8042.mask = 128'h33ffffff33ffffff0000000000000700;

	lut_sub lut_8045 ({sk[1808], x909x, n_n54, n_n263, n_n6521, x1928x, x21022x}, x21028x);
	defparam lut_8045.LUT_SIZE = 7;
	defparam lut_8045.mask = 128'h33ffffff33ffffff5f5f5f5f5f7f5fff;

	lut_sub lut_8050 ({sk[1809], x389x, n_n6524, x373x, x464x, x463x}, x21027x);
	defparam lut_8050.LUT_SIZE = 6;
	defparam lut_8050.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_8056 ({sk[1810], i_14_, i_13_, i_12_, n_n273, x922x, x902x}, x869x);
	defparam lut_8056.LUT_SIZE = 7;
	defparam lut_8056.mask = 128'h33ffffff33ffffff0000000000010100;

	lut_sub lut_8059 ({sk[1811], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x1881x);
	defparam lut_8059.LUT_SIZE = 7;
	defparam lut_8059.mask = 128'h33ffffff33ffffff1050405040000000;

	lut_sub lut_8067 ({sk[1812], i_14_, i_13_, i_12_, i_15_, x163x, n_n270}, x1852x);
	defparam lut_8067.LUT_SIZE = 7;
	defparam lut_8067.mask = 128'h33ffffff33ffffff3333333337337373;

	lut_sub lut_8072 ({sk[1813], i_14_, i_13_, i_12_, i_15_, n_n48, n_n247}, x21052x);
	defparam lut_8072.LUT_SIZE = 7;
	defparam lut_8072.mask = 128'h33ffffff33ffffff0111101111011110;

	lut_sub lut_8085 ({sk[1814], n_n48, n_n53, n_n95, x136x, x68x, x204x}, x21039x);
	defparam lut_8085.LUT_SIZE = 7;
	defparam lut_8085.mask = 128'h33ffffff33ffffff00000fff77777fff;

	lut_sub lut_8090 ({sk[1815], n_n48, n_n53, n_n95, x55x, x1280x, x1917x}, x21040x);
	defparam lut_8090.LUT_SIZE = 7;
	defparam lut_8090.mask = 128'h33ffffff33ffffff00003f3f55ff7fff;

	lut_sub lut_8095 ({sk[1816], n_n271, x909x, x159x, n_n53, x68x, x764x}, x781x);
	defparam lut_8095.LUT_SIZE = 7;
	defparam lut_8095.mask = 128'h33ffffff33ffffff57575757575757ff;

	lut_sub lut_8099 ({sk[1817], n_n148, n_n266, n_n271, x146x, x909x, n_n226}, x21044x);
	defparam lut_8099.LUT_SIZE = 7;
	defparam lut_8099.mask = 128'h33ffffff33ffffff0013001300133333;

	lut_sub lut_8103 ({sk[1818], n_n266, n_n271, n_n9, x184x, x909x, x209x}, x21045x);
	defparam lut_8103.LUT_SIZE = 7;
	defparam lut_8103.mask = 128'h33ffffff33ffffff0000030311331333;

	lut_sub lut_8107 ({sk[1819], n_n57, n_n56, x160x, n_n60, x1870x, x3821x}, x21046x);
	defparam lut_8107.LUT_SIZE = 7;
	defparam lut_8107.mask = 128'h33ffffff33ffffff55555fff77777fff;

	lut_sub lut_8112 ({sk[1820], i_14_, i_13_, i_12_, n_n273, x922x, x908x}, x20344x);
	defparam lut_8112.LUT_SIZE = 7;
	defparam lut_8112.mask = 128'h33ffffff33ffffff0001010000000000;

	lut_sub lut_8115 ({sk[1821], n_n273, n_n220, x922x, x908x, n_n256, x478x}, x695x);
	defparam lut_8115.LUT_SIZE = 7;
	defparam lut_8115.mask = 128'h33ffffff33ffffff555555555557555f;

	lut_sub lut_8119 ({sk[1822], i_14_, i_13_, i_12_, i_15_, x908x, n_n270}, x1930x);
	defparam lut_8119.LUT_SIZE = 7;
	defparam lut_8119.mask = 128'h33ffffff33ffffff0533335000000000;

	lut_sub lut_8124 ({sk[1823], n_n273, x922x, n_n70, n_n6867, x4509x, x286x}, x865x);
	defparam lut_8124.LUT_SIZE = 7;
	defparam lut_8124.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_8129 ({sk[1824], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1910x);
	defparam lut_8129.LUT_SIZE = 7;
	defparam lut_8129.mask = 128'h33ffffff33ffffff0000001050005040;

	lut_sub lut_8136 ({sk[1825], i_7_, i_8_, i_6_, x915x, x83x}, x701x);
	defparam lut_8136.LUT_SIZE = 6;
	defparam lut_8136.mask = 64'h77ff77ff00000010;

	lut_sub lut_8138 ({sk[1826], x915x, n_n261, x188x, x109x, x117x}, n_n2926);
	defparam lut_8138.LUT_SIZE = 6;
	defparam lut_8138.mask = 64'h77ff77ff0000007f;

	lut_sub lut_8142 ({sk[1827], i_7_, i_8_, i_6_, x915x, x1321x}, n_n3722);
	defparam lut_8142.LUT_SIZE = 6;
	defparam lut_8142.mask = 64'h77ff77ff00000010;

	lut_sub lut_8144 ({sk[1828], n_n255, n_n197, x569x, x524x, x21109x, x24121x}, n_n3221);
	defparam lut_8144.LUT_SIZE = 7;
	defparam lut_8144.mask = 128'h33ffffff33ffffffbfffbfffbfffffff;

	lut_sub lut_8150 ({sk[1829], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1943x);
	defparam lut_8150.LUT_SIZE = 7;
	defparam lut_8150.mask = 128'h33ffffff33ffffff0000000105000504;

	lut_sub lut_8157 ({sk[1830], i_7_, i_8_, i_6_, x915x, x77x}, x821x);
	defparam lut_8157.LUT_SIZE = 6;
	defparam lut_8157.mask = 64'h77ff77ff00000010;

	lut_sub lut_8159 ({sk[1831], x915x, n_n258, n_n261, x902x, x1855x}, x383x);
	defparam lut_8159.LUT_SIZE = 6;
	defparam lut_8159.mask = 64'h77ff77ff00000507;

	lut_sub lut_8162 ({sk[1832], i_14_, i_13_, i_12_, i_15_, x908x, n_n270}, x1896x);
	defparam lut_8162.LUT_SIZE = 7;
	defparam lut_8162.mask = 128'h33ffffff33ffffff0537335000000000;

	lut_sub lut_8168 ({sk[1833], x915x, n_n263, x1860x, x552x, x3776x, x1238x}, x21106x);
	defparam lut_8168.LUT_SIZE = 7;
	defparam lut_8168.mask = 128'h33ffffff33ffffff3f3f3f3f3f3f7fff;

	lut_sub lut_8173 ({sk[1834], i_14_, i_13_, i_12_, i_15_, n_n247, x55x}, x1885x);
	defparam lut_8173.LUT_SIZE = 7;
	defparam lut_8173.mask = 128'h33ffffff33ffffff5557555777557575;

	lut_sub lut_8181 ({sk[1835], i_15_, x915x, n_n258, n_n263, x912x, n_n137}, x548x);
	defparam lut_8181.LUT_SIZE = 7;
	defparam lut_8181.mask = 128'h33ffffff33ffffff0000000300000507;

	lut_sub lut_8184 ({sk[1836], i_7_, i_8_, i_6_, x907x, x915x, n_n220}, x774x);
	defparam lut_8184.LUT_SIZE = 7;
	defparam lut_8184.mask = 128'h33ffffff33ffffff0000000000000100;

	lut_sub lut_8186 ({sk[1837], i_14_, i_13_, i_12_, x912x, x189x, x157x}, x1194x);
	defparam lut_8186.LUT_SIZE = 7;
	defparam lut_8186.mask = 128'h33ffffff33ffffff7f7777777f777777;

	lut_sub lut_8191 ({sk[1838], i_14_, i_13_, i_12_, x908x, x902x, n_n100}, x20061x);
	defparam lut_8191.LUT_SIZE = 7;
	defparam lut_8191.mask = 128'h33ffffff33ffffff1115051515111505;

	lut_sub lut_8204 ({sk[1839], n_n94, x686x, x391x, x548x, x774x, x1194x}, x20062x);
	defparam lut_8204.LUT_SIZE = 7;
	defparam lut_8204.mask = 128'h33ffffff33ffffff3fffffff7fffffff;

	lut_sub lut_8210 ({sk[1840], x915x, n_n261, n_n263, n_n144, n_n150, n_n58}, x24101x);
	defparam lut_8210.LUT_SIZE = 7;
	defparam lut_8210.mask = 128'h33ffffff33ffffffffffffffff808080;

	lut_sub lut_8214 ({sk[1841], n_n57, n_n6036, n_n94, n_n52, n_n8, x24101x}, n_n1798);
	defparam lut_8214.LUT_SIZE = 7;
	defparam lut_8214.mask = 128'h33ffffff33ffffffaabbffffafbfffff;

	lut_sub lut_8219 ({sk[1842], i_9_, i_10_, i_11_, i_15_, n_n220}, x1199x);
	defparam lut_8219.LUT_SIZE = 6;
	defparam lut_8219.mask = 64'h77ff77ff00010001;

	lut_sub lut_8222 ({sk[1843], n_n108, n_n57, n_n56, n_n147, x100x, x1199x}, n_n1787);
	defparam lut_8222.LUT_SIZE = 7;
	defparam lut_8222.mask = 128'h33ffffff33ffffff00775f7f00ff5fff;

	lut_sub lut_8228 ({sk[1844], i_14_, i_13_, i_12_, i_15_, n_n275, x228x}, x1201x);
	defparam lut_8228.LUT_SIZE = 7;
	defparam lut_8228.mask = 128'h33ffffff33ffffff5557555755557755;

	lut_sub lut_8234 ({sk[1845], i_14_, i_13_, i_12_, x908x, x902x}, x230x);
	defparam lut_8234.LUT_SIZE = 6;
	defparam lut_8234.mask = 64'h77ff77ff50300000;

	lut_sub lut_8237 ({sk[1846], i_14_, i_13_, i_12_, x908x, x902x, x897x}, x1200x);
	defparam lut_8237.LUT_SIZE = 7;
	defparam lut_8237.mask = 128'h33ffffff33ffffff33000f0000005500;

	lut_sub lut_8241 ({sk[1847], i_14_, i_13_, i_12_, i_15_, n_n282, n_n247}, x21639x);
	defparam lut_8241.LUT_SIZE = 7;
	defparam lut_8241.mask = 128'h33ffffff33ffffff0505500300003300;

	lut_sub lut_8248 ({sk[1848], i_14_, i_13_, i_12_, i_15_, n_n282, n_n253}, x1564x);
	defparam lut_8248.LUT_SIZE = 7;
	defparam lut_8248.mask = 128'h33ffffff33ffffff0707700700007700;

	lut_sub lut_8261 ({sk[1849], i_9_, i_10_, i_11_, i_15_, n_n225, n_n137}, x428x);
	defparam lut_8261.LUT_SIZE = 7;
	defparam lut_8261.mask = 128'h33ffffff33ffffff5555555557555555;

	lut_sub lut_8265 ({sk[1850], i_14_, i_13_, i_12_, i_15_, x900x, n_n267}, x21638x);
	defparam lut_8265.LUT_SIZE = 7;
	defparam lut_8265.mask = 128'h33ffffff33ffffff3333500500005500;

	lut_sub lut_8272 ({sk[1851], n_n1, n_n2, x21639x, x1564x, x428x, x21638x}, n_n1701);
	defparam lut_8272.LUT_SIZE = 7;
	defparam lut_8272.mask = 128'h33ffffff33ffffff00000f0f77ff7fff;

	lut_sub lut_8277 ({sk[1852], i_14_, i_13_, i_12_, x905x, x899x}, x237x);
	defparam lut_8277.LUT_SIZE = 6;
	defparam lut_8277.mask = 64'h77ff77ff55300000;

	lut_sub lut_8281 ({sk[1853], i_9_, i_10_, i_11_, i_15_, n_n138, n_n225}, x857x);
	defparam lut_8281.LUT_SIZE = 7;
	defparam lut_8281.mask = 128'h33ffffff33ffffff3333373333333333;

	lut_sub lut_8285 ({sk[1854], i_14_, i_13_, i_12_, i_15_, n_n270, x379x}, x21642x);
	defparam lut_8285.LUT_SIZE = 7;
	defparam lut_8285.mask = 128'h33ffffff33ffffff5757755755555555;

	lut_sub lut_8291 ({sk[1855], i_14_, i_13_, i_12_, i_15_, n_n242, x240x}, x21641x);
	defparam lut_8291.LUT_SIZE = 7;
	defparam lut_8291.mask = 128'h33ffffff33ffffff5757755555555555;

	lut_sub lut_8296 ({sk[1856], n_n1, n_n2, x237x, x857x, x21642x, x21641x}, n_n1699);
	defparam lut_8296.LUT_SIZE = 7;
	defparam lut_8296.mask = 128'h33ffffff33ffffff00007f7f5fff7fff;

	lut_sub lut_8303 ({sk[1857], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x21646x);
	defparam lut_8303.LUT_SIZE = 7;
	defparam lut_8303.mask = 128'h33ffffff33ffffff1111440000000000;

	lut_sub lut_8310 ({sk[1858], i_14_, i_13_, i_12_, i_15_, n_n275, n_n270}, x21647x);
	defparam lut_8310.LUT_SIZE = 7;
	defparam lut_8310.mask = 128'h33ffffff33ffffff0505500700007700;

	lut_sub lut_8320 ({sk[1859], i_14_, i_13_, i_12_, i_15_, n_n247, n_n275}, x1202x);
	defparam lut_8320.LUT_SIZE = 7;
	defparam lut_8320.mask = 128'h33ffffff33ffffff0707700700007700;

	lut_sub lut_8333 ({sk[1860], x915x, n_n273, n_n283, x21646x, x21647x, x1202x}, x21648x);
	defparam lut_8333.LUT_SIZE = 7;
	defparam lut_8333.mask = 128'h33ffffff33ffffff0000000000553f7f;

	lut_sub lut_8337 ({sk[1861], n_n1701, n_n1699, x21648x}, n_n1685);
	defparam lut_8337.LUT_SIZE = 4;
	defparam lut_8337.mask = 16'h777f;

	lut_sub lut_8341 ({sk[1862], i_9_, i_10_, i_11_, i_15_, n_n222}, x426x);
	defparam lut_8341.LUT_SIZE = 6;
	defparam lut_8341.mask = 64'h77ff77ff05000000;

	lut_sub lut_8344 ({sk[1863], n_n2, n_n268, n_n220, x899x, x212x, x903x}, x21653x);
	defparam lut_8344.LUT_SIZE = 7;
	defparam lut_8344.mask = 128'h33ffffff33ffffff00003377000f337f;

	lut_sub lut_8348 ({sk[1864], i_15_, x916x, n_n271, n_n138, x426x, x21653x}, n_n1738);
	defparam lut_8348.LUT_SIZE = 7;
	defparam lut_8348.mask = 128'h33ffffff33ffffff5555557f5555557f;

	lut_sub lut_8353 ({sk[1865], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x158x);
	defparam lut_8353.LUT_SIZE = 7;
	defparam lut_8353.mask = 128'h33ffffff33ffffff0000000000005000;

	lut_sub lut_8356 ({sk[1866], i_14_, i_13_, i_12_, i_15_, n_n253, x226x}, x1812x);
	defparam lut_8356.LUT_SIZE = 7;
	defparam lut_8356.mask = 128'h33ffffff33ffffff5557555755557755;

	lut_sub lut_8362 ({sk[1867], n_n208, n_n266, x916x, x200x, x158x, x1812x}, x21666x);
	defparam lut_8362.LUT_SIZE = 7;
	defparam lut_8362.mask = 128'h33ffffff33ffffff0000003f0055007f;

	lut_sub lut_8366 ({sk[1868], i_14_, i_13_, i_12_, n_n3, x898x, x904x}, x690x);
	defparam lut_8366.LUT_SIZE = 7;
	defparam lut_8366.mask = 128'h33ffffff33ffffff0300050000000000;

	lut_sub lut_8369 ({sk[1869], i_14_, i_13_, i_12_, x900x, x906x}, x270x);
	defparam lut_8369.LUT_SIZE = 6;
	defparam lut_8369.mask = 64'h77ff77ff30500000;

	lut_sub lut_8372 ({sk[1870], i_14_, i_13_, i_12_, x898x, x904x}, x129x);
	defparam lut_8372.LUT_SIZE = 6;
	defparam lut_8372.mask = 64'h77ff77ff03030050;

	lut_sub lut_8376 ({sk[1871], n_n4, n_n3, n_n222, x898x, x270x, x129x}, x835x);
	defparam lut_8376.LUT_SIZE = 7;
	defparam lut_8376.mask = 128'h33ffffff33ffffff0000555f3333777f;

	lut_sub lut_8380 ({sk[1872], i_14_, i_13_, i_12_, i_15_, x906x, n_n267}, x21668x);
	defparam lut_8380.LUT_SIZE = 7;
	defparam lut_8380.mask = 128'h33ffffff33ffffff0000000500003300;

	lut_sub lut_8383 ({sk[1873], i_14_, i_13_, i_12_, x900x, x21668x}, x151x);
	defparam lut_8383.LUT_SIZE = 6;
	defparam lut_8383.mask = 64'h77ff77ff57555555;

	lut_sub lut_8386 ({sk[1874], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x1628x);
	defparam lut_8386.LUT_SIZE = 7;
	defparam lut_8386.mask = 128'h33ffffff33ffffff0005000500007300;

	lut_sub lut_8391 ({sk[1875], n_n3, n_n7225, x690x, x835x, x151x, x270x}, x21672x);
	defparam lut_8391.LUT_SIZE = 7;
	defparam lut_8391.mask = 128'h33ffffff33ffffff0fffffff7fffffff;

	lut_sub lut_8397 ({sk[1876], i_15_, n_n111, n_n135, n_n137, x151x, x313x}, x24097x);
	defparam lut_8397.LUT_SIZE = 7;
	defparam lut_8397.mask = 128'h33ffffff33ffffff8800000080000000;

	lut_sub lut_8400 ({sk[1877], n_n208, x916x, n_n3, x1628x, x21672x, x24097x}, x21673x);
	defparam lut_8400.LUT_SIZE = 7;
	defparam lut_8400.mask = 128'h33ffffff33ffffff333f333f333fbbbf;

	lut_sub lut_8404 ({sk[1878], n_n2, n_n220, x898x, x901x, x237x, x21651x}, n_n1740);
	defparam lut_8404.LUT_SIZE = 7;
	defparam lut_8404.mask = 128'h33ffffff33ffffff5555555577777fff;

	lut_sub lut_8409 ({sk[1879], n_n266, x916x, n_n271, n_n3246, n_n32, x1731x}, n_n1736);
	defparam lut_8409.LUT_SIZE = 7;
	defparam lut_8409.mask = 128'h33ffffff33ffffff0f0f0f5f0f0f3f7f;

	lut_sub lut_8413 ({sk[1880], n_n2, n_n220, x912x, x902x, x3201x, x3203x}, x21656x);
	defparam lut_8413.LUT_SIZE = 7;
	defparam lut_8413.mask = 128'h33ffffff33ffffff7777777777777fff;

	lut_sub lut_8418 ({sk[1881], n_n110, n_n268, n_n147, x605x, n_n3513, x3192x}, x21665x);
	defparam lut_8418.LUT_SIZE = 7;
	defparam lut_8418.mask = 128'h33ffffff33ffffff7f7f7fff7f7fffff;

	lut_sub lut_8424 ({sk[1882], n_n1738, x21666x, n_n1740, n_n1736, x21656x, x21665x}, x21674x);
	defparam lut_8424.LUT_SIZE = 7;
	defparam lut_8424.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_8431 ({sk[1883], i_14_, i_13_, i_12_, i_15_, n_n259, n_n267}, x1793x);
	defparam lut_8431.LUT_SIZE = 7;
	defparam lut_8431.mask = 128'h33ffffff33ffffff0007000700007000;

	lut_sub lut_8438 ({sk[1884], n_n4, n_n7225, n_n8, x690x, x622x, x1793x}, x21684x);
	defparam lut_8438.LUT_SIZE = 7;
	defparam lut_8438.mask = 128'h33ffffff33ffffff3f3fffff7fffffff;

	lut_sub lut_8444 ({sk[1885], n_n273, n_n7402, x922x, n_n76, n_n7406, n_n6856}, x21679x);
	defparam lut_8444.LUT_SIZE = 7;
	defparam lut_8444.mask = 128'h33ffffff33ffffff7777ffff777fffff;

	lut_sub lut_8449 ({sk[1886], n_n53, x902x, n_n256, n_n225, n_n7442, x656x}, x21680x);
	defparam lut_8449.LUT_SIZE = 7;
	defparam lut_8449.mask = 128'h33ffffff33ffffff7777777777777fff;

	lut_sub lut_8454 ({sk[1887], x835x, x21684x, x21679x, x21680x}, n_n1703);
	defparam lut_8454.LUT_SIZE = 5;
	defparam lut_8454.mask = 32'h3f3f7fff;

	lut_sub lut_8459 ({sk[1888], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x143x);
	defparam lut_8459.LUT_SIZE = 7;
	defparam lut_8459.mask = 128'h33ffffff33ffffff0010000000004000;

	lut_sub lut_8462 ({sk[1889], i_15_, n_n207, n_n138, n_n17, n_n6814, x3143x}, x24096x);
	defparam lut_8462.LUT_SIZE = 7;
	defparam lut_8462.mask = 128'h33ffffff33ffffff8888800088888080;

	lut_sub lut_8466 ({sk[1890], x902x, n_n227, n_n225, n_n6812, x143x, x24096x}, x21697x);
	defparam lut_8466.LUT_SIZE = 7;
	defparam lut_8466.mask = 128'h33ffffff33ffffffafafbfbfafafbfff;

	lut_sub lut_8471 ({sk[1891], n_n6847, n_n1757, n_n7297, x641x, x21693x, x21697x}, n_n1704);
	defparam lut_8471.LUT_SIZE = 7;
	defparam lut_8471.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_8478 ({sk[1892], n_n273, x905x, n_n222, x922x, x899x, n_n225}, x3128x);
	defparam lut_8478.LUT_SIZE = 7;
	defparam lut_8478.mask = 128'h33ffffff33ffffff000000000101010f;

	lut_sub lut_8481 ({sk[1893], n_n2, n_n222, x901x, n_n6871, n_n6876, x3128x}, x21704x);
	defparam lut_8481.LUT_SIZE = 7;
	defparam lut_8481.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_8486 ({sk[1894], n_n53, n_n6868, n_n6867, n_n8, n_n6861, x21704x}, n_n1752);
	defparam lut_8486.LUT_SIZE = 7;
	defparam lut_8486.mask = 128'h33ffffff33ffffff77ffffff7fffffff;

	lut_sub lut_8492 ({sk[1895], i_14_, i_13_, i_12_, i_15_, x900x, n_n267}, x21706x);
	defparam lut_8492.LUT_SIZE = 7;
	defparam lut_8492.mask = 128'h33ffffff33ffffff3333500500005500;

	lut_sub lut_8499 ({sk[1896], i_14_, i_13_, i_12_, i_15_, n_n282, x21706x}, x1207x);
	defparam lut_8499.LUT_SIZE = 7;
	defparam lut_8499.mask = 128'h33ffffff33ffffff5757755755557555;

	lut_sub lut_8506 ({sk[1897], i_14_, i_13_, i_12_, x898x, x904x}, x363x);
	defparam lut_8506.LUT_SIZE = 6;
	defparam lut_8506.mask = 64'h77ff77ff33500000;

	lut_sub lut_8510 ({sk[1898], i_14_, i_13_, i_12_, i_15_, n_n253, x363x}, x1206x);
	defparam lut_8510.LUT_SIZE = 7;
	defparam lut_8510.mask = 128'h33ffffff33ffffff5555555755557755;

	lut_sub lut_8515 ({sk[1899], n_n1, n_n2, n_n62, n_n1752, x1207x, x1206x}, x21709x);
	defparam lut_8515.LUT_SIZE = 7;
	defparam lut_8515.mask = 128'h33ffffff33ffffff0f0f3fff5f5f7fff;

	lut_sub lut_8520 ({sk[1900], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1209x);
	defparam lut_8520.LUT_SIZE = 7;
	defparam lut_8520.mask = 128'h33ffffff33ffffff0053000000005300;

	lut_sub lut_8525 ({sk[1901], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1208x);
	defparam lut_8525.LUT_SIZE = 7;
	defparam lut_8525.mask = 128'h33ffffff33ffffff0053500000530000;

	lut_sub lut_8531 ({sk[1902], i_14_, i_13_, i_12_, n_n3, x898x}, n_n1356);
	defparam lut_8531.LUT_SIZE = 6;
	defparam lut_8531.mask = 64'h77ff77ff11010000;

	lut_sub lut_8535 ({sk[1903], n_n208, x916x, n_n258, x908x, x906x}, x22043x);
	defparam lut_8535.LUT_SIZE = 6;
	defparam lut_8535.mask = 64'h77ff77ff00000007;

	lut_sub lut_8538 ({sk[1904], n_n208, x916x, n_n220, x899x, x902x}, x22044x);
	defparam lut_8538.LUT_SIZE = 6;
	defparam lut_8538.mask = 64'h77ff77ff00000007;

	lut_sub lut_8541 ({sk[1905], n_n3, x99x, n_n95, n_n49, x22043x, x22044x}, n_n1208);
	defparam lut_8541.LUT_SIZE = 7;
	defparam lut_8541.mask = 128'h33ffffff33ffffff777777777fffffff;

	lut_sub lut_8547 ({sk[1906], i_7_, i_8_, i_6_, x922x, x140x}, n_n639);
	defparam lut_8547.LUT_SIZE = 6;
	defparam lut_8547.mask = 64'h77ff77ff00100000;

	lut_sub lut_8549 ({sk[1907], i_14_, i_13_, i_12_, n_n273, x922x, x902x}, x694x);
	defparam lut_8549.LUT_SIZE = 7;
	defparam lut_8549.mask = 128'h33ffffff33ffffff0101000100000000;

	lut_sub lut_8553 ({sk[1908], n_n7402, n_n7441, n_n6860, n_n6861, n_n639, x694x}, x22054x);
	defparam lut_8553.LUT_SIZE = 7;
	defparam lut_8553.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_8560 ({sk[1909], i_14_, i_13_, i_12_, x903x, x897x}, x365x);
	defparam lut_8560.LUT_SIZE = 6;
	defparam lut_8560.mask = 64'h77ff77ff00055003;

	lut_sub lut_8564 ({sk[1910], i_7_, i_8_, i_6_, x916x, x56x}, x680x);
	defparam lut_8564.LUT_SIZE = 6;
	defparam lut_8564.mask = 64'h77ff77ff00000100;

	lut_sub lut_8566 ({sk[1911], i_7_, i_8_, i_6_, x915x, x899x, n_n228}, x22775x);
	defparam lut_8566.LUT_SIZE = 7;
	defparam lut_8566.mask = 128'h33ffffff33ffffff0100010000000000;

	lut_sub lut_8569 ({sk[1912], n_n268, x135x, n_n206, x56x, x365x, x22775x}, n_n790);
	defparam lut_8569.LUT_SIZE = 7;
	defparam lut_8569.mask = 128'h33ffffff33ffffff555555ff7f7f7fff;

	lut_sub lut_8574 ({sk[1913], i_14_, i_13_, i_12_, x903x, x897x}, x1211x);
	defparam lut_8574.LUT_SIZE = 6;
	defparam lut_8574.mask = 64'h77ff77ff07003030;

	lut_sub lut_8579 ({sk[1914], i_14_, i_13_, i_12_, x908x, x902x}, x276x);
	defparam lut_8579.LUT_SIZE = 6;
	defparam lut_8579.mask = 64'h77ff77ff00000503;

	lut_sub lut_8582 ({sk[1915], i_14_, i_13_, i_12_, x908x, x902x}, x312x);
	defparam lut_8582.LUT_SIZE = 6;
	defparam lut_8582.mask = 64'h77ff77ff05003030;

	lut_sub lut_8586 ({sk[1916], i_14_, i_13_, i_12_, x908x, x902x}, x1210x);
	defparam lut_8586.LUT_SIZE = 6;
	defparam lut_8586.mask = 64'h77ff77ff05003533;

	lut_sub lut_8592 ({sk[1917], n_n208, x916x, x905x, n_n258, x899x, n_n228}, x743x);
	defparam lut_8592.LUT_SIZE = 7;
	defparam lut_8592.mask = 128'h33ffffff33ffffff0000000000000357;

	lut_sub lut_8595 ({sk[1918], i_14_, i_13_, i_12_, i_15_, n_n242, n_n138}, x1214x);
	defparam lut_8595.LUT_SIZE = 7;
	defparam lut_8595.mask = 128'h33ffffff33ffffff5053505070535070;

	lut_sub lut_8601 ({sk[1919], i_9_, i_10_, i_11_, i_15_, n_n256}, x22336x);
	defparam lut_8601.LUT_SIZE = 6;
	defparam lut_8601.mask = 64'h77ff77ff00400400;

	lut_sub lut_8604 ({sk[1920], i_14_, i_13_, i_12_, i_15_, n_n242, n_n259}, x1212x);
	defparam lut_8604.LUT_SIZE = 7;
	defparam lut_8604.mask = 128'h33ffffff33ffffff0007000070037030;

	lut_sub lut_8613 ({sk[1921], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1956x);
	defparam lut_8613.LUT_SIZE = 7;
	defparam lut_8613.mask = 128'h33ffffff33ffffff0001000004010404;

	lut_sub lut_8619 ({sk[1922], n_n208, x916x, n_n3, x906x, n_n256, x1956x}, x833x);
	defparam lut_8619.LUT_SIZE = 7;
	defparam lut_8619.mask = 128'h33ffffff33ffffff0055005500550357;

	lut_sub lut_8622 ({sk[1923], i_14_, i_13_, i_12_, x900x, x906x}, x244x);
	defparam lut_8622.LUT_SIZE = 6;
	defparam lut_8622.mask = 64'h77ff77ff03005050;

	lut_sub lut_8626 ({sk[1924], i_14_, i_13_, i_12_, i_15_, n_n247, x244x}, x1216x);
	defparam lut_8626.LUT_SIZE = 7;
	defparam lut_8626.mask = 128'h33ffffff33ffffff5577555575577575;

	lut_sub lut_8634 ({sk[1925], i_14_, i_13_, i_12_, i_15_, n_n282, n_n267}, x1215x);
	defparam lut_8634.LUT_SIZE = 7;
	defparam lut_8634.mask = 128'h33ffffff33ffffff0057000070037030;

	lut_sub lut_8644 ({sk[1926], n_n208, x916x, n_n258, x908x, n_n228, x902x}, x642x);
	defparam lut_8644.LUT_SIZE = 7;
	defparam lut_8644.mask = 128'h33ffffff33ffffff0000000000000357;

	lut_sub lut_8647 ({sk[1927], i_14_, i_13_, i_12_, i_15_, n_n282, x312x}, x1218x);
	defparam lut_8647.LUT_SIZE = 7;
	defparam lut_8647.mask = 128'h33ffffff33ffffff5577555575577575;

	lut_sub lut_8655 ({sk[1928], i_14_, i_13_, i_12_, i_15_, x907x, n_n247}, x1217x);
	defparam lut_8655.LUT_SIZE = 7;
	defparam lut_8655.mask = 128'h33ffffff33ffffff0077000050055050;

	lut_sub lut_8663 ({sk[1929], n_n139, x435x, x19241x, x19240x}, x5959x);
	defparam lut_8663.LUT_SIZE = 5;
	defparam lut_8663.mask = 32'h3f3f007f;

	lut_sub lut_8667 ({sk[1930], x917x, n_n208, x19235x, x19236x, x5960x}, x19243x);
	defparam lut_8667.LUT_SIZE = 6;
	defparam lut_8667.mask = 64'h77ff77ff5555557f;

	lut_sub lut_8671 ({sk[1931], n_n281, n_n142, x911x, x19249x, x19233x, x331x}, x5957x);
	defparam lut_8671.LUT_SIZE = 7;
	defparam lut_8671.mask = 128'h33ffffff33ffffff00007f7f00007fff;

	lut_sub lut_8676 ({sk[1932], x917x, n_n139, n_n283, x19245x, x19246x, x1268x}, x19250x);
	defparam lut_8676.LUT_SIZE = 7;
	defparam lut_8676.mask = 128'h33ffffff33ffffff00005555003f557f;

	lut_sub lut_8680 ({sk[1933], n_n281, n_n130, n_n132, x905x, x285x, x19256x}, x19260x);
	defparam lut_8680.LUT_SIZE = 7;
	defparam lut_8680.mask = 128'h33ffffff33ffffff0077007700770f7f;

	lut_sub lut_8684 ({sk[1934], i_8_, n_n155, x896x, x1271x, x412x, x19252x}, x19261x);
	defparam lut_8684.LUT_SIZE = 7;
	defparam lut_8684.mask = 128'h33ffffff33ffffff000f007f000f00ff;

	lut_sub lut_8689 ({sk[1935], x921x, n_n124, n_n273, x19321x, x19322x, x1399x}, x19323x);
	defparam lut_8689.LUT_SIZE = 7;
	defparam lut_8689.mask = 128'h33ffffff33ffffff00005555003f557f;

	lut_sub lut_8693 ({sk[1936], n_n130, x19329x, x19327x, x19328x}, x5861x);
	defparam lut_8693.LUT_SIZE = 5;
	defparam lut_8693.mask = 32'h3f3f007f;

	lut_sub lut_8697 ({sk[1937], i_7_, i_8_, i_6_, x896x, x398x, x19324x}, x19331x);
	defparam lut_8697.LUT_SIZE = 7;
	defparam lut_8697.mask = 128'h33ffffff33ffffff0000000f00070000;

	lut_sub lut_8701 ({sk[1938], x921x, n_n283, x184x, x19336x, x398x, x196x}, x5849x);
	defparam lut_8701.LUT_SIZE = 7;
	defparam lut_8701.mask = 128'h33ffffff33ffffff0000000000007fff;

	lut_sub lut_8706 ({sk[1939], n_n127, n_n266, x896x, x5855x, x1458x, x5848x}, x19339x);
	defparam lut_8706.LUT_SIZE = 7;
	defparam lut_8706.mask = 128'h33ffffff33ffffff5f5f5fff7f7f7fff;

	lut_sub lut_8711 ({sk[1940], n_n281, x913x, n_n122, x19314x, x196x, x215x}, x5876x);
	defparam lut_8711.LUT_SIZE = 7;
	defparam lut_8711.mask = 128'h33ffffff33ffffff007f007f007f00ff;

	lut_sub lut_8716 ({sk[1941], n_n121, x19309x, x398x, x5874x, x19308x}, x19315x);
	defparam lut_8716.LUT_SIZE = 6;
	defparam lut_8716.mask = 64'h77ff77ff33337fff;

	lut_sub lut_8721 ({sk[1942], x921x, n_n208, n_n122, x412x, x1500x, x19344x}, x19349x);
	defparam lut_8721.LUT_SIZE = 7;
	defparam lut_8721.mask = 128'h33ffffff33ffffff005f005f005f337f;

	lut_sub lut_8725 ({sk[1943], i_6_, i_1_, i_2_, i_0_, n_n264, x1887x}, x19355x);
	defparam lut_8725.LUT_SIZE = 7;
	defparam lut_8725.mask = 128'h33ffffff33ffffff0000350000000500;

	lut_sub lut_8728 ({sk[1944], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19284x);
	defparam lut_8728.LUT_SIZE = 7;
	defparam lut_8728.mask = 128'h33ffffff33ffffffcc0c000000000000;

	lut_sub lut_8733 ({sk[1945], i_9_, i_10_, i_12_, i_11_}, x5999x);
	defparam lut_8733.LUT_SIZE = 5;
	defparam lut_8733.mask = 32'h3f3f3100;

	lut_sub lut_8737 ({sk[1946], n_n279, x901x, x897x, x19284x, x5999x}, x1220x);
	defparam lut_8737.LUT_SIZE = 6;
	defparam lut_8737.mask = 64'h77ff77ff77777fff;

	lut_sub lut_8742 ({sk[1947], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x5994x);
	defparam lut_8742.LUT_SIZE = 7;
	defparam lut_8742.mask = 128'h33ffffff33ffffff0000cc0c00000000;

	lut_sub lut_8747 ({sk[1948], x911x, n_n279, x900x, n_n149, x5994x}, x1224x);
	defparam lut_8747.LUT_SIZE = 6;
	defparam lut_8747.mask = 64'h77ff77ff777f77ff;

	lut_sub lut_8752 ({sk[1949], i_9_, i_10_, i_12_, i_11_}, x1223x);
	defparam lut_8752.LUT_SIZE = 5;
	defparam lut_8752.mask = 32'h3f3fff20;

	lut_sub lut_8755 ({sk[1950], n_n189, x961x, n_n177, x1220x, x1224x, x1223x}, n_n5017);
	defparam lut_8755.LUT_SIZE = 7;
	defparam lut_8755.mask = 128'h33ffffff33ffffff003f003f557fffff;

	lut_sub lut_8760 ({sk[1951], i_14_, i_13_, i_12_, x912x, n_n137}, x285x);
	defparam lut_8760.LUT_SIZE = 6;
	defparam lut_8760.mask = 64'h77ff77ff55757555;

	lut_sub lut_8764 ({sk[1952], i_14_, i_13_, i_12_, x911x, n_n138, x285x}, x19314x);
	defparam lut_8764.LUT_SIZE = 7;
	defparam lut_8764.mask = 128'h33ffffff33ffffff77777f777f777777;

	lut_sub lut_8769 ({sk[1953], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x397x);
	defparam lut_8769.LUT_SIZE = 7;
	defparam lut_8769.mask = 128'h33ffffff33ffffff0000777f00000000;

	lut_sub lut_8773 ({sk[1954], i_15_, n_n281, n_n163, n_n279, n_n247, x397x}, x19309x);
	defparam lut_8773.LUT_SIZE = 7;
	defparam lut_8773.mask = 128'h33ffffff33ffffff55ff77ff57ff57ff;

	lut_sub lut_8778 ({sk[1955], i_9_, i_10_, i_12_, i_11_}, x196x);
	defparam lut_8778.LUT_SIZE = 5;
	defparam lut_8778.mask = 32'h3f3f0070;

	lut_sub lut_8781 ({sk[1956], i_9_, i_10_, i_12_, i_11_}, x215x);
	defparam lut_8781.LUT_SIZE = 5;
	defparam lut_8781.mask = 32'h3f3f0700;

	lut_sub lut_8784 ({sk[1957], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x398x);
	defparam lut_8784.LUT_SIZE = 7;
	defparam lut_8784.mask = 128'h33ffffff33ffffff4000100010000000;

	lut_sub lut_8788 ({sk[1958], i_7_, i_8_, i_6_, n_n165, n_n264}, x5874x);
	defparam lut_8788.LUT_SIZE = 6;
	defparam lut_8788.mask = 64'h77ff77ff00010001;

	lut_sub lut_8791 ({sk[1959], i_9_, i_10_, i_11_, i_15_, n_n220, x19237x}, x19308x);
	defparam lut_8791.LUT_SIZE = 7;
	defparam lut_8791.mask = 128'h33ffffff33ffffff5555555557ffffff;

	lut_sub lut_8796 ({sk[1960], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1893x);
	defparam lut_8796.LUT_SIZE = 7;
	defparam lut_8796.mask = 128'h33ffffff33ffffff0010001050004040;

	lut_sub lut_8803 ({sk[1961], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x122x);
	defparam lut_8803.LUT_SIZE = 7;
	defparam lut_8803.mask = 128'h33ffffff33ffffff0000000010004040;

	lut_sub lut_8807 ({sk[1962], n_n271, x909x, x60x, n_n6190, x155x, x122x}, n_n4261);
	defparam lut_8807.LUT_SIZE = 7;
	defparam lut_8807.mask = 128'h33ffffff33ffffff0f0f0f0f0f0f7fff;

	lut_sub lut_8812 ({sk[1963], n_n5796, n_n130, n_n122, n_n132, n_n107, x250x}, x20715x);
	defparam lut_8812.LUT_SIZE = 7;
	defparam lut_8812.mask = 128'h33ffffff33ffffff05777777ffffffff;

	lut_sub lut_8819 ({sk[1964], n_n266, x268x, x909x, x200x, n_n4948, n_n4950}, x20723x);
	defparam lut_8819.LUT_SIZE = 7;
	defparam lut_8819.mask = 128'h33ffffff33ffffff77777777777f77ff;

	lut_sub lut_8824 ({sk[1965], x268x, n_n57, n_n56, x157x, x277x, x112x}, x20724x);
	defparam lut_8824.LUT_SIZE = 7;
	defparam lut_8824.mask = 128'h33ffffff33ffffff00557f7f00ff7fff;

	lut_sub lut_8830 ({sk[1966], n_n266, n_n271, x909x, n_n65, x186x, x44x}, x465x);
	defparam lut_8830.LUT_SIZE = 7;
	defparam lut_8830.mask = 128'h33ffffff33ffffff0000003f0055007f;

	lut_sub lut_8834 ({sk[1967], n_n110, n_n57, n_n56, x90x, x82x, x155x}, n_n4259);
	defparam lut_8834.LUT_SIZE = 7;
	defparam lut_8834.mask = 128'h33ffffff33ffffff00335f7f0033ffff;

	lut_sub lut_8839 ({sk[1968], n_n110, n_n57, n_n56, x90x, x60x, x122x}, x721x);
	defparam lut_8839.LUT_SIZE = 7;
	defparam lut_8839.mask = 128'h33ffffff33ffffff000f777f00ff77ff;

	lut_sub lut_8844 ({sk[1969], n_n266, x909x, x258x, x720x, x682x, x70x}, x20729x);
	defparam lut_8844.LUT_SIZE = 7;
	defparam lut_8844.mask = 128'h33ffffff33ffffff3f3f3f3f3f3f7fff;

	lut_sub lut_8849 ({sk[1970], n_n57, n_n56, x265x, x111x, x1898x, x884x}, x24187x);
	defparam lut_8849.LUT_SIZE = 7;
	defparam lut_8849.mask = 128'h33ffffff33ffffffaaaa8080aa008000;

	lut_sub lut_8854 ({sk[1971], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1233x);
	defparam lut_8854.LUT_SIZE = 7;
	defparam lut_8854.mask = 128'h33ffffff33ffffff0101000505000504;

	lut_sub lut_8864 ({sk[1972], i_9_, i_10_, i_11_, n_n261, n_n263, x922x}, x309x);
	defparam lut_8864.LUT_SIZE = 7;
	defparam lut_8864.mask = 128'h33ffffff33ffffff0000000500000011;

	lut_sub lut_8867 ({sk[1973], i_9_, i_10_, i_11_, n_n261, x922x}, x571x);
	defparam lut_8867.LUT_SIZE = 6;
	defparam lut_8867.mask = 64'h77ff77ff01000000;

	lut_sub lut_8869 ({sk[1974], i_7_, i_8_, i_6_, n_n258, x922x, x900x}, x665x);
	defparam lut_8869.LUT_SIZE = 7;
	defparam lut_8869.mask = 128'h33ffffff33ffffff0100000000000000;

	lut_sub lut_8871 ({sk[1975], i_7_, i_8_, i_6_, x922x, n_n270}, x737x);
	defparam lut_8871.LUT_SIZE = 6;
	defparam lut_8871.mask = 64'h77ff77ff00001000;

	lut_sub lut_8873 ({sk[1976], i_9_, i_10_, i_8_, i_11_, n_n272, x922x}, x20300x);
	defparam lut_8873.LUT_SIZE = 7;
	defparam lut_8873.mask = 128'h33ffffff33ffffff0000000101000100;

	lut_sub lut_8877 ({sk[1977], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x105x);
	defparam lut_8877.LUT_SIZE = 7;
	defparam lut_8877.mask = 128'h33ffffff33ffffff1010004000000000;

	lut_sub lut_8881 ({sk[1978], x915x, n_n261, n_n263, x97x, x1910x, x105x}, x20774x);
	defparam lut_8881.LUT_SIZE = 7;
	defparam lut_8881.mask = 128'h33ffffff33ffffff0000000000335f7f;

	lut_sub lut_8885 ({sk[1979], n_n226, x159x, x208x, x314x, n_n100, n_n94}, n_n3209);
	defparam lut_8885.LUT_SIZE = 7;
	defparam lut_8885.mask = 128'h33ffffff33ffffff0555377737773777;

	lut_sub lut_8890 ({sk[1980], i_14_, i_13_, i_12_, i_15_, n_n270}, x1855x);
	defparam lut_8890.LUT_SIZE = 6;
	defparam lut_8890.mask = 64'h77ff77ff00015054;

	lut_sub lut_8897 ({sk[1981], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x1238x);
	defparam lut_8897.LUT_SIZE = 7;
	defparam lut_8897.mask = 128'h33ffffff33ffffff0141400504000400;

	lut_sub lut_8906 ({sk[1982], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x222x);
	defparam lut_8906.LUT_SIZE = 7;
	defparam lut_8906.mask = 128'h33ffffff33ffffff1010004000000000;

	lut_sub lut_8910 ({sk[1983], i_14_, i_13_, i_12_, x914x, x909x, n_n261}, x873x);
	defparam lut_8910.LUT_SIZE = 7;
	defparam lut_8910.mask = 128'h33ffffff33ffffff0001010000000000;

	lut_sub lut_8913 ({sk[1984], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1905x);
	defparam lut_8913.LUT_SIZE = 7;
	defparam lut_8913.mask = 128'h33ffffff33ffffff0000000105000504;

	lut_sub lut_8920 ({sk[1985], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1928x);
	defparam lut_8920.LUT_SIZE = 7;
	defparam lut_8920.mask = 128'h33ffffff33ffffff0000000105000504;

	lut_sub lut_8927 ({sk[1986], i_14_, i_13_, i_12_, n_n283, x914x, x922x}, x21022x);
	defparam lut_8927.LUT_SIZE = 7;
	defparam lut_8927.mask = 128'h33ffffff33ffffff0001010000000000;

	lut_sub lut_8930 ({sk[1987], i_7_, i_8_, i_6_, x916x, x44x}, x742x);
	defparam lut_8930.LUT_SIZE = 6;
	defparam lut_8930.mask = 64'h77ff77ff00010000;

	lut_sub lut_8932 ({sk[1988], i_14_, i_13_, i_12_, i_15_, x905x, n_n259}, x1240x);
	defparam lut_8932.LUT_SIZE = 7;
	defparam lut_8932.mask = 128'h33ffffff33ffffff0537005555055550;

	lut_sub lut_8944 ({sk[1989], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x232x);
	defparam lut_8944.LUT_SIZE = 7;
	defparam lut_8944.mask = 128'h33ffffff33ffffff0000000000100040;

	lut_sub lut_8947 ({sk[1990], i_14_, i_13_, i_12_, i_15_, n_n275, x897x}, x1241x);
	defparam lut_8947.LUT_SIZE = 7;
	defparam lut_8947.mask = 128'h33ffffff33ffffff0000003303555530;

	lut_sub lut_8954 ({sk[1991], n_n151, n_n208, x909x, n_n261, x232x, x1241x}, n_n2876);
	defparam lut_8954.LUT_SIZE = 7;
	defparam lut_8954.mask = 128'h33ffffff33ffffff00000077000f007f;

	lut_sub lut_8958 ({sk[1992], i_14_, i_13_, i_12_, i_15_, x914x, n_n247}, x1243x);
	defparam lut_8958.LUT_SIZE = 7;
	defparam lut_8958.mask = 128'h33ffffff33ffffff0537335555055550;

	lut_sub lut_8971 ({sk[1993], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x1242x);
	defparam lut_8971.LUT_SIZE = 7;
	defparam lut_8971.mask = 128'h33ffffff33ffffff3305005555055550;

	lut_sub lut_8982 ({sk[1994], n_n271, x78x, x909x, x497x, x3599x, x1242x}, x21312x);
	defparam lut_8982.LUT_SIZE = 7;
	defparam lut_8982.mask = 128'h33ffffff33ffffff3f3f3f3f3f7f3fff;

	lut_sub lut_8987 ({sk[1995], i_14_, i_13_, i_12_, i_15_, n_n253, n_n267}, x1245x);
	defparam lut_8987.LUT_SIZE = 7;
	defparam lut_8987.mask = 128'h33ffffff33ffffff0757507333003330;

	lut_sub lut_9002 ({sk[1996], i_14_, i_13_, i_12_, x900x, x906x}, x138x);
	defparam lut_9002.LUT_SIZE = 6;
	defparam lut_9002.mask = 64'h77ff77ff33050000;

	lut_sub lut_9006 ({sk[1997], n_n258, x900x, x94x, x108x, x138x}, x1244x);
	defparam lut_9006.LUT_SIZE = 6;
	defparam lut_9006.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_9011 ({sk[1998], n_n57, n_n6046, n_n49, x372x, x894x, x386x}, x21303x);
	defparam lut_9011.LUT_SIZE = 7;
	defparam lut_9011.mask = 128'h33ffffff33ffffff7f7fffff7fffffff;

	lut_sub lut_9017 ({sk[1999], n_n266, x909x, n_n222, x898x, x1090x, x1243x}, x24112x);
	defparam lut_9017.LUT_SIZE = 7;
	defparam lut_9017.mask = 128'h33ffffff33ffffffffffffffffff8880;

	lut_sub lut_9022 ({sk[2000], n_n56, n_n6035, x515x, x569x, x872x, x1091x}, x24113x);
	defparam lut_9022.LUT_SIZE = 7;
	defparam lut_9022.mask = 128'h33ffffff33ffffffc000000080000000;

	lut_sub lut_9025 ({sk[2001], i_9_, i_10_, i_11_, i_15_, n_n222}, x472x);
	defparam lut_9025.LUT_SIZE = 6;
	defparam lut_9025.mask = 64'h77ff77ff00000050;

	lut_sub lut_9028 ({sk[2002], i_7_, i_8_, i_6_, n_n110, x909x, n_n4394}, x21724x);
	defparam lut_9028.LUT_SIZE = 7;
	defparam lut_9028.mask = 128'h33ffffff33ffffff5555555555575557;

	lut_sub lut_9032 ({sk[2003], i_15_, n_n57, n_n56, n_n138, x472x, x21724x}, n_n1788);
	defparam lut_9032.LUT_SIZE = 7;
	defparam lut_9032.mask = 128'h33ffffff33ffffff55775f7f55775f7f;

	lut_sub lut_9037 ({sk[2004], n_n266, n_n271, x909x, n_n22, x212x, x426x}, n_n1791);
	defparam lut_9037.LUT_SIZE = 7;
	defparam lut_9037.mask = 128'h33ffffff33ffffff0000003f0077007f;

	lut_sub lut_9042 ({sk[2005], i_9_, i_10_, i_11_, i_15_, n_n222}, x379x);
	defparam lut_9042.LUT_SIZE = 6;
	defparam lut_9042.mask = 64'h77ff77ff00000500;

	lut_sub lut_9045 ({sk[2006], i_14_, i_13_, i_12_, i_15_, n_n242, x379x}, x1247x);
	defparam lut_9045.LUT_SIZE = 7;
	defparam lut_9045.mask = 128'h33ffffff33ffffff5757555755557755;

	lut_sub lut_9052 ({sk[2007], n_n266, n_n271, x909x, x100x, x472x, x1247x}, x21719x);
	defparam lut_9052.LUT_SIZE = 7;
	defparam lut_9052.mask = 128'h33ffffff33ffffff00000055003f007f;

	lut_sub lut_9056 ({sk[2008], i_15_, n_n57, n_n56, n_n32, n_n137, x158x}, x21736x);
	defparam lut_9056.LUT_SIZE = 7;
	defparam lut_9056.mask = 128'h33ffffff33ffffff007f557f007f557f;

	lut_sub lut_9062 ({sk[2009], n_n111, n_n57, x200x, n_n4948, n_n32, n_n4940}, x21737x);
	defparam lut_9062.LUT_SIZE = 7;
	defparam lut_9062.mask = 128'h33ffffff33ffffff5f5f7fff5f5fffff;

	lut_sub lut_9068 ({sk[2010], n_n57, n_n56, n_n76, x520x, x165x, x426x}, x24103x);
	defparam lut_9068.LUT_SIZE = 7;
	defparam lut_9068.mask = 128'h33ffffff33fffffff0f0a0a0c0008000;

	lut_sub lut_9073 ({sk[2011], n_n57, n_n56, n_n22, n_n76, n_n6190, x165x}, x21718x);
	defparam lut_9073.LUT_SIZE = 7;
	defparam lut_9073.mask = 128'h33ffffff33ffffff33337f7f33ff7fff;

	lut_sub lut_9078 ({sk[2012], n_n220, n_n57, x899x, x902x, x3096x, x3098x}, x21727x);
	defparam lut_9078.LUT_SIZE = 7;
	defparam lut_9078.mask = 128'h33ffffff33ffffff7777777777777fff;

	lut_sub lut_9083 ({sk[2013], i_14_, i_13_, i_12_, n_n3, x898x}, x5762x);
	defparam lut_9083.LUT_SIZE = 6;
	defparam lut_9083.mask = 64'h77ff77ff00000110;

	lut_sub lut_9086 ({sk[2014], i_14_, i_13_, i_12_, n_n3, x904x}, x2811x);
	defparam lut_9086.LUT_SIZE = 6;
	defparam lut_9086.mask = 64'h77ff77ff00001011;

	lut_sub lut_9090 ({sk[2015], i_14_, i_13_, i_12_, i_15_, n_n4, n_n267}, x2810x);
	defparam lut_9090.LUT_SIZE = 7;
	defparam lut_9090.mask = 128'h33ffffff33ffffff0111000000000000;

	lut_sub lut_9094 ({sk[2016], n_n208, x916x, n_n42, x5762x, x2811x, x2810x}, n_n1173);
	defparam lut_9094.LUT_SIZE = 7;
	defparam lut_9094.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_9099 ({sk[2017], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1252x);
	defparam lut_9099.LUT_SIZE = 7;
	defparam lut_9099.mask = 128'h33ffffff33ffffff0010001040004040;

	lut_sub lut_9105 ({sk[2018], n_n208, x916x, n_n197, x466x, n_n7345, x1252x}, n_n1210);
	defparam lut_9105.LUT_SIZE = 7;
	defparam lut_9105.mask = 128'h33ffffff33ffffff3f3f3f3f3f3f7fff;

	lut_sub lut_9110 ({sk[2019], i_14_, i_13_, i_12_, i_15_, n_n242, x903x}, x1254x);
	defparam lut_9110.LUT_SIZE = 7;
	defparam lut_9110.mask = 128'h33ffffff33ffffff0000007703030330;

	lut_sub lut_9118 ({sk[2020], i_7_, i_8_, i_6_, x916x, x85x, x1254x}, n_n789);
	defparam lut_9118.LUT_SIZE = 7;
	defparam lut_9118.mask = 128'h33ffffff33ffffff0000000000050003;

	lut_sub lut_9121 ({sk[2021], i_14_, i_13_, i_12_, x903x, x897x}, x320x);
	defparam lut_9121.LUT_SIZE = 6;
	defparam lut_9121.mask = 64'h77ff77ff00000503;

	lut_sub lut_9124 ({sk[2022], i_14_, i_13_, i_12_, i_15_, n_n275, x320x}, x1257x);
	defparam lut_9124.LUT_SIZE = 7;
	defparam lut_9124.mask = 128'h33ffffff33ffffff5577555575557555;

	lut_sub lut_9130 ({sk[2023], i_14_, i_13_, i_12_, i_15_, x907x, n_n259}, x22469x);
	defparam lut_9130.LUT_SIZE = 7;
	defparam lut_9130.mask = 128'h33ffffff33ffffff0000000000375050;

	lut_sub lut_9135 ({sk[2024], i_14_, i_13_, i_12_, x913x, x911x}, x292x);
	defparam lut_9135.LUT_SIZE = 6;
	defparam lut_9135.mask = 64'h77ff77ff07003000;

	lut_sub lut_9139 ({sk[2025], i_14_, i_13_, i_12_, i_15_, n_n242, x441x}, x22468x);
	defparam lut_9139.LUT_SIZE = 7;
	defparam lut_9139.mask = 128'h33ffffff33ffffff5555555555577575;

	lut_sub lut_9144 ({sk[2026], n_n271, x909x, n_n252, x22469x, x292x, x22468x}, x2309x);
	defparam lut_9144.LUT_SIZE = 7;
	defparam lut_9144.mask = 128'h33ffffff33ffffff0000000000007fff;

	lut_sub lut_9149 ({sk[2027], i_14_, i_13_, i_12_, x913x, x911x, x904x}, x22467x);
	defparam lut_9149.LUT_SIZE = 7;
	defparam lut_9149.mask = 128'h33ffffff33ffffff003f00000f550000;

	lut_sub lut_9154 ({sk[2028], n_n13, n_n57, n_n56, n_n246, x22467x, x22468x}, x22470x);
	defparam lut_9154.LUT_SIZE = 7;
	defparam lut_9154.mask = 128'h33ffffff33ffffff00007f7f00ffffff;

	lut_sub lut_9160 ({sk[2029], i_14_, i_13_, i_12_, i_15_, n_n282, n_n247}, x1736x);
	defparam lut_9160.LUT_SIZE = 7;
	defparam lut_9160.mask = 128'h33ffffff33ffffff0077000070077070;

	lut_sub lut_9173 ({sk[2030], n_n266, n_n271, x909x, n_n102, x175x, x1736x}, n_n372);
	defparam lut_9173.LUT_SIZE = 7;
	defparam lut_9173.mask = 128'h33ffffff33ffffff0000007f0055007f;

	lut_sub lut_9178 ({sk[2031], i_14_, i_13_, i_12_, x903x, x897x}, x405x);
	defparam lut_9178.LUT_SIZE = 6;
	defparam lut_9178.mask = 64'h77ff77ff07003000;

	lut_sub lut_9182 ({sk[2032], i_14_, i_13_, i_12_, i_15_, n_n270, x405x}, x1259x);
	defparam lut_9182.LUT_SIZE = 7;
	defparam lut_9182.mask = 128'h33ffffff33ffffff5577555575577575;

	lut_sub lut_9190 ({sk[2033], i_14_, i_13_, i_12_, i_15_, n_n275, n_n259}, x1258x);
	defparam lut_9190.LUT_SIZE = 7;
	defparam lut_9190.mask = 128'h33ffffff33ffffff0033000030077070;

	lut_sub lut_9200 ({sk[2034], n_n57, n_n56, x1259x, x1258x, x427x, x1609x}, x22481x);
	defparam lut_9200.LUT_SIZE = 7;
	defparam lut_9200.mask = 128'h33ffffff33ffffff000033ff5f5f7fff;

	lut_sub lut_9205 ({sk[2035], i_14_, i_13_, i_12_, x898x, x904x}, x1306x);
	defparam lut_9205.LUT_SIZE = 6;
	defparam lut_9205.mask = 64'h77ff77ff07005055;

	lut_sub lut_9211 ({sk[2036], n_n41, n_n105, n_n100, n_n94, x1306x, x229x}, x22487x);
	defparam lut_9211.LUT_SIZE = 7;
	defparam lut_9211.mask = 128'h33ffffff33ffffff03770f7f03ff0fff;

	lut_sub lut_9217 ({sk[2037], n_n151, n_n136, n_n148, x22242x, x22240x, x22241x}, x24082x);
	defparam lut_9217.LUT_SIZE = 7;
	defparam lut_9217.mask = 128'h33ffffff33ffffff8080800080800000;

	lut_sub lut_9220 ({sk[2038], i_7_, i_6_, x261x, x24082x}, x22493x);
	defparam lut_9220.LUT_SIZE = 5;
	defparam lut_9220.mask = 32'h3f3fbbbb;

	lut_sub lut_9226 ({sk[2039], i_14_, i_13_, i_12_, x907x, x915x, n_n261}, x877x);
	defparam lut_9226.LUT_SIZE = 7;
	defparam lut_9226.mask = 128'h33ffffff33ffffff0000000001000101;

	lut_sub lut_9230 ({sk[2040], i_14_, i_13_, i_12_, x915x, n_n261, x901x}, x22496x);
	defparam lut_9230.LUT_SIZE = 7;
	defparam lut_9230.mask = 128'h33ffffff33ffffff0001000000010000;

	lut_sub lut_9233 ({sk[2041], n_n94, n_n6830, n_n6829, x144x, x877x, x22496x}, n_n464);
	defparam lut_9233.LUT_SIZE = 7;
	defparam lut_9233.mask = 128'h33ffffff33ffffff77ffffff7fffffff;

	lut_sub lut_9239 ({sk[2042], x915x, x914x, n_n263, x912x, n_n256}, x688x);
	defparam lut_9239.LUT_SIZE = 6;
	defparam lut_9239.mask = 64'h77ff77ff00000105;

	lut_sub lut_9242 ({sk[2043], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x1261x);
	defparam lut_9242.LUT_SIZE = 7;
	defparam lut_9242.mask = 128'h33ffffff33ffffff0050000044004444;

	lut_sub lut_9251 ({sk[2044], n_n104, n_n94, x881x, x189x, x688x, x112x}, x22502x);
	defparam lut_9251.LUT_SIZE = 7;
	defparam lut_9251.mask = 128'h33ffffff33ffffff33ff7fff33ffffff;

	lut_sub lut_9257 ({sk[2045], x915x, n_n261, n_n263, x166x, n_n105, x229x}, n_n467);
	defparam lut_9257.LUT_SIZE = 7;
	defparam lut_9257.mask = 128'h33ffffff33ffffff00000000005f3f7f;

	lut_sub lut_9262 ({sk[2046], i_7_, i_8_, i_6_, x917x, x48x, x929x}, x22492x);
	defparam lut_9262.LUT_SIZE = 7;
	defparam lut_9262.mask = 128'h33ffffff33ffffff55575555555f555f;

	lut_sub lut_9269 ({sk[2047], n_n139, x211x, x266x, x294x, x599x, n_n3615}, x24081x);
	defparam lut_9269.LUT_SIZE = 7;
	defparam lut_9269.mask = 128'h33ffffff33ffffff8888888880000000;

	lut_sub lut_9272 ({sk[2048], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x19292x);
	defparam lut_9272.LUT_SIZE = 7;
	defparam lut_9272.mask = 128'h33ffffff33ffffff4050105010505050;

	lut_sub lut_9278 ({sk[2049], i_4_, n_n152, n_n153, x259x, x282x, x19292x}, n_n5048);
	defparam lut_9278.LUT_SIZE = 7;
	defparam lut_9278.mask = 128'h33ffffff33ffffff000f777f00007777;

	lut_sub lut_9282 ({sk[2050], i_9_, i_10_, i_11_, i_15_, n_n281, n_n279}, x19241x);
	defparam lut_9282.LUT_SIZE = 7;
	defparam lut_9282.mask = 128'h33ffffff33ffffff000000ff35ff3500;

	lut_sub lut_9289 ({sk[2051], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19233x);
	defparam lut_9289.LUT_SIZE = 7;
	defparam lut_9289.mask = 128'h33ffffff33ffffff000000800000ffff;

	lut_sub lut_9292 ({sk[2052], i_9_, i_10_, i_13_, i_12_, i_11_}, x331x);
	defparam lut_9292.LUT_SIZE = 6;
	defparam lut_9292.mask = 64'h77ff77ff00007f00;

	lut_sub lut_9296 ({sk[2053], i_14_, i_13_, i_12_, x911x, x19233x, x331x}, x19235x);
	defparam lut_9296.LUT_SIZE = 7;
	defparam lut_9296.mask = 128'h33ffffff33ffffff7f77777777777777;

	lut_sub lut_9300 ({sk[2054], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x5968x);
	defparam lut_9300.LUT_SIZE = 7;
	defparam lut_9300.mask = 128'h33ffffff33ffffff0000000000800000;

	lut_sub lut_9302 ({sk[2055], i_9_, i_10_, i_13_, i_12_, i_11_}, x454x);
	defparam lut_9302.LUT_SIZE = 6;
	defparam lut_9302.mask = 64'h77ff77ff007f0000;

	lut_sub lut_9306 ({sk[2056], i_9_, i_10_, n_n281, x912x, x5968x, x454x}, x19236x);
	defparam lut_9306.LUT_SIZE = 7;
	defparam lut_9306.mask = 128'h33ffffff33ffffffffff777f777f777f;

	lut_sub lut_9311 ({sk[2057], i_9_, i_10_, i_11_, i_15_, n_n220, x19237x}, x19240x);
	defparam lut_9311.LUT_SIZE = 7;
	defparam lut_9311.mask = 128'h33ffffff33ffffff55555555575555ff;

	lut_sub lut_9315 ({sk[2058], i_11_, i_15_, n_n281, n_n274, n_n132, n_n204}, x5960x);
	defparam lut_9315.LUT_SIZE = 7;
	defparam lut_9315.mask = 128'h33ffffff33ffffff1113111111111111;

	lut_sub lut_9318 ({sk[2059], i_9_, i_10_, n_n281, x912x, x5968x, x454x}, x19249x);
	defparam lut_9318.LUT_SIZE = 7;
	defparam lut_9318.mask = 128'h33ffffff33ffffffffff777f777f777f;

	lut_sub lut_9323 ({sk[2060], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19237x);
	defparam lut_9323.LUT_SIZE = 7;
	defparam lut_9323.mask = 128'h33ffffff33ffffff00000000222a0000;

	lut_sub lut_9326 ({sk[2061], i_9_, i_10_, i_11_, i_15_, n_n220, x19237x}, x19245x);
	defparam lut_9326.LUT_SIZE = 7;
	defparam lut_9326.mask = 128'h33ffffff33ffffff55555555575555ff;

	lut_sub lut_9330 ({sk[2062], i_14_, i_13_, i_12_, i_15_, n_n259, x284x}, x19246x);
	defparam lut_9330.LUT_SIZE = 7;
	defparam lut_9330.mask = 128'h33ffffff33ffffff5577577755777777;

	lut_sub lut_9335 ({sk[2063], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1268x);
	defparam lut_9335.LUT_SIZE = 7;
	defparam lut_9335.mask = 128'h33ffffff33ffffff4050105010505050;

	lut_sub lut_9341 ({sk[2064], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19259x);
	defparam lut_9341.LUT_SIZE = 7;
	defparam lut_9341.mask = 128'h33ffffff33ffffff000000007fff0000;

	lut_sub lut_9346 ({sk[2065], i_9_, i_10_}, x19257x);
	defparam lut_9346.LUT_SIZE = 3;
	defparam lut_9346.mask = 8'h5d;

	lut_sub lut_9349 ({sk[2066], i_8_, n_n281, n_n272, x912x, x19259x, x19257x}, x1271x);
	defparam lut_9349.LUT_SIZE = 7;
	defparam lut_9349.mask = 128'h33ffffff33ffffff00ff00ff0077007f;

	lut_sub lut_9354 ({sk[2067], i_14_, i_13_, i_12_, n_n247, x912x, x331x}, x19321x);
	defparam lut_9354.LUT_SIZE = 7;
	defparam lut_9354.mask = 128'h33ffffff33ffffff775555555f555555;

	lut_sub lut_9358 ({sk[2068], i_14_, i_13_, i_12_, x911x, x287x, x19320x}, x19322x);
	defparam lut_9358.LUT_SIZE = 7;
	defparam lut_9358.mask = 128'h33ffffff33ffffff7f77777777777777;

	lut_sub lut_9362 ({sk[2069], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1399x);
	defparam lut_9362.LUT_SIZE = 7;
	defparam lut_9362.mask = 128'h33ffffff33ffffff4050105010505050;

	lut_sub lut_9368 ({sk[2070], i_14_, i_13_, i_12_, i_15_, n_n242, x412x}, x19329x);
	defparam lut_9368.LUT_SIZE = 7;
	defparam lut_9368.mask = 128'h33ffffff33ffffff5555575557557755;

	lut_sub lut_9373 ({sk[2071], i_9_, i_10_, i_12_, i_11_, i_15_, n_n281}, x19327x);
	defparam lut_9373.LUT_SIZE = 7;
	defparam lut_9373.mask = 128'h33ffffff33ffffff0000404040400fff;

	lut_sub lut_9378 ({sk[2072], i_14_, i_13_, i_12_, x912x, n_n137, x19326x}, x19328x);
	defparam lut_9378.LUT_SIZE = 7;
	defparam lut_9378.mask = 128'h33ffffff33ffffff77777f777f777777;

	lut_sub lut_9383 ({sk[2073], i_15_, n_n281, n_n163, n_n279, n_n247, x397x}, x19324x);
	defparam lut_9383.LUT_SIZE = 7;
	defparam lut_9383.mask = 128'h33ffffff33ffffff55ff77ff57ff57ff;

	lut_sub lut_9388 ({sk[2074], n_n281, n_n165, n_n284, n_n273, x901x, x5918x}, x5855x);
	defparam lut_9388.LUT_SIZE = 7;
	defparam lut_9388.mask = 128'h33ffffff33ffffff0000000500000007;

	lut_sub lut_9391 ({sk[2075], i_14_, i_13_, i_12_, x912x, n_n137, x397x}, x19336x);
	defparam lut_9391.LUT_SIZE = 7;
	defparam lut_9391.mask = 128'h33ffffff33ffffff777777777f777777;

	lut_sub lut_9395 ({sk[2076], n_n12, x186x, x176x, n_n48, n_n53, x70x}, n_n3457);
	defparam lut_9395.LUT_SIZE = 7;
	defparam lut_9395.mask = 128'h33ffffff33ffffff05370f3f37373f3f;

	lut_sub lut_9400 ({sk[2077], i_7_, i_8_, i_6_, n_n65, x922x, x44x}, n_n3579);
	defparam lut_9400.LUT_SIZE = 7;
	defparam lut_9400.mask = 128'h33ffffff33ffffff0300110000000000;

	lut_sub lut_9403 ({sk[2078], n_n108, n_n48, n_n53, x70x, x1938x, n_n3579}, x20823x);
	defparam lut_9403.LUT_SIZE = 7;
	defparam lut_9403.mask = 128'h33ffffff33ffffff555f777f555fffff;

	lut_sub lut_9408 ({sk[2079], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1280x);
	defparam lut_9408.LUT_SIZE = 7;
	defparam lut_9408.mask = 128'h33ffffff33ffffff0105000505000404;

	lut_sub lut_9418 ({sk[2080], i_14_, i_13_, i_12_, x898x, x904x, x171x}, x1917x);
	defparam lut_9418.LUT_SIZE = 7;
	defparam lut_9418.mask = 128'h33ffffff33ffffff555f555f77555555;

	lut_sub lut_9423 ({sk[2081], i_14_, i_13_, i_12_, i_15_, n_n242, n_n138}, x194x);
	defparam lut_9423.LUT_SIZE = 7;
	defparam lut_9423.mask = 128'h33ffffff33ffffff5053505070505050;

	lut_sub lut_9427 ({sk[2082], n_n228, x902x, n_n207, x480x, x700x, n_n6824}, x20368x);
	defparam lut_9427.LUT_SIZE = 7;
	defparam lut_9427.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_9432 ({sk[2083], x913x, n_n258, n_n207, n_n59, x194x, x20368x}, n_n2875);
	defparam lut_9432.LUT_SIZE = 7;
	defparam lut_9432.mask = 128'h33ffffff33ffffff557f557f557f55ff;

	lut_sub lut_9437 ({sk[2084], i_14_, i_13_, i_12_, x900x, x906x}, x1285x);
	defparam lut_9437.LUT_SIZE = 6;
	defparam lut_9437.mask = 64'h77ff77ff30057000;

	lut_sub lut_9442 ({sk[2085], i_14_, i_13_, i_12_, x898x, x904x}, x226x);
	defparam lut_9442.LUT_SIZE = 6;
	defparam lut_9442.mask = 64'h77ff77ff30500000;

	lut_sub lut_9445 ({sk[2086], i_14_, i_13_, i_12_, i_15_, n_n253, x226x}, x1286x);
	defparam lut_9445.LUT_SIZE = 7;
	defparam lut_9445.mask = 128'h33ffffff33ffffff5557555755557755;

	lut_sub lut_9451 ({sk[2087], n_n48, n_n53, n_n80, x279x, x249x, x228x}, n_n1778);
	defparam lut_9451.LUT_SIZE = 7;
	defparam lut_9451.mask = 128'h33ffffff33ffffff00005f5f33ff7fff;

	lut_sub lut_9456 ({sk[2088], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1292x);
	defparam lut_9456.LUT_SIZE = 7;
	defparam lut_9456.mask = 128'h33ffffff33ffffff1010401000000000;

	lut_sub lut_9461 ({sk[2089], i_14_, i_13_, i_12_, x907x, x915x, n_n261}, x22231x);
	defparam lut_9461.LUT_SIZE = 7;
	defparam lut_9461.mask = 128'h33ffffff33ffffff0001000001000000;

	lut_sub lut_9464 ({sk[2090], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x1294x);
	defparam lut_9464.LUT_SIZE = 7;
	defparam lut_9464.mask = 128'h33ffffff33ffffff0555500500333300;

	lut_sub lut_9472 ({sk[2091], i_14_, i_13_, i_12_, i_15_, n_n282, n_n247}, x1293x);
	defparam lut_9472.LUT_SIZE = 7;
	defparam lut_9472.mask = 128'h33ffffff33ffffff0555500000003300;

	lut_sub lut_9479 ({sk[2092], x915x, x914x, n_n258, n_n263, x722x, x50x}, x24184x);
	defparam lut_9479.LUT_SIZE = 7;
	defparam lut_9479.mask = 128'h33ffffff33ffffffccccccccc8c8c8c0;

	lut_sub lut_9484 ({sk[2093], n_n6843, n_n6834, n_n6835, x825x, x24184x}, n_n1212);
	defparam lut_9484.LUT_SIZE = 6;
	defparam lut_9484.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_9490 ({sk[2094], i_14_, i_13_, i_12_, x907x, x915x, n_n261}, x434x);
	defparam lut_9490.LUT_SIZE = 7;
	defparam lut_9490.mask = 128'h33ffffff33ffffff0000000001000001;

	lut_sub lut_9493 ({sk[2095], i_14_, i_13_, i_12_, x908x, x902x}, x1942x);
	defparam lut_9493.LUT_SIZE = 6;
	defparam lut_9493.mask = 64'h77ff77ff55053033;

	lut_sub lut_9500 ({sk[2096], n_n4, n_n6847, n_n6829, n_n6823, n_n6824, x1942x}, x22076x);
	defparam lut_9500.LUT_SIZE = 7;
	defparam lut_9500.mask = 128'h33ffffff33ffffff3fffffff7fffffff;

	lut_sub lut_9506 ({sk[2097], i_9_, i_10_, i_11_, i_15_, x202x, n_n225}, x1298x);
	defparam lut_9506.LUT_SIZE = 7;
	defparam lut_9506.mask = 128'h33ffffff33ffffff3333333333333377;

	lut_sub lut_9510 ({sk[2098], i_14_, i_13_, i_12_, x905x, x899x}, x305x);
	defparam lut_9510.LUT_SIZE = 6;
	defparam lut_9510.mask = 64'h77ff77ff00070003;

	lut_sub lut_9514 ({sk[2099], i_7_, i_8_, i_6_, x915x, n_n65, n_n15}, x22778x);
	defparam lut_9514.LUT_SIZE = 7;
	defparam lut_9514.mask = 128'h33ffffff33ffffff0300070000000000;

	lut_sub lut_9518 ({sk[2100], x915x, n_n283, x227x, x305x, x22778x}, n_n792);
	defparam lut_9518.LUT_SIZE = 6;
	defparam lut_9518.mask = 64'h77ff77ff5555557f;

	lut_sub lut_9522 ({sk[2101], n_n31, n_n48, n_n53, x120x, x91x, x201x}, n_n830);
	defparam lut_9522.LUT_SIZE = 7;
	defparam lut_9522.mask = 128'h33ffffff33ffffff003f557f003fffff;

	lut_sub lut_9527 ({sk[2102], n_n48, n_n53, x114x, x107x, x128x, x161x}, x22700x);
	defparam lut_9527.LUT_SIZE = 7;
	defparam lut_9527.mask = 128'h33ffffff33ffffff00003f3f5fff7fff;

	lut_sub lut_9533 ({sk[2103], x915x, n_n258, x898x, n_n261, x515x, x569x}, n_n3615);
	defparam lut_9533.LUT_SIZE = 7;
	defparam lut_9533.mask = 128'h33ffffff33ffffff777777777777777f;

	lut_sub lut_9537 ({sk[2104], i_14_, i_13_, i_12_, n_n139, x913x, x911x}, x4962x);
	defparam lut_9537.LUT_SIZE = 7;
	defparam lut_9537.mask = 128'h33ffffff33ffffff0500000003000000;

	lut_sub lut_9540 ({sk[2105], i_14_, i_13_, i_12_, i_15_, n_n247, n_n267}, x1310x);
	defparam lut_9540.LUT_SIZE = 7;
	defparam lut_9540.mask = 128'h33ffffff33ffffff0077000070037070;

	lut_sub lut_9552 ({sk[2106], i_14_, i_13_, i_12_, i_15_, x901x, n_n253}, x22507x);
	defparam lut_9552.LUT_SIZE = 7;
	defparam lut_9552.mask = 128'h33ffffff33ffffff0055000000370000;

	lut_sub lut_9557 ({sk[2107], x907x, x901x, n_n256, x41x, x112x, x22507x}, x24077x);
	defparam lut_9557.LUT_SIZE = 7;
	defparam lut_9557.mask = 128'h33ffffff33ffffff8080800080008000;

	lut_sub lut_9560 ({sk[2108], n_n1, n_n2, n_n104, x112x, x1310x, x24077x}, n_n356);
	defparam lut_9560.LUT_SIZE = 7;
	defparam lut_9560.mask = 128'h33ffffff33ffffff0000aaaa3fffbfff;

	lut_sub lut_9565 ({sk[2109], i_9_, i_10_, i_11_, i_15_, n_n256}, x22516x);
	defparam lut_9565.LUT_SIZE = 6;
	defparam lut_9565.mask = 64'h77ff77ff55000000;

	lut_sub lut_9570 ({sk[2110], i_9_, i_10_, i_11_, i_15_, n_n256}, x22513x);
	defparam lut_9570.LUT_SIZE = 6;
	defparam lut_9570.mask = 64'h77ff77ff05005000;

	lut_sub lut_9575 ({sk[2111], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x22514x);
	defparam lut_9575.LUT_SIZE = 7;
	defparam lut_9575.mask = 128'h33ffffff33ffffff0000000040114040;

	lut_sub lut_9581 ({sk[2112], n_n1, n_n258, x902x, x124x, x897x, x22516x}, x2260x);
	defparam lut_9581.LUT_SIZE = 7;
	defparam lut_9581.mask = 128'h33ffffff33ffffff000000005f5f7fff;

	lut_sub lut_9586 ({sk[2113], i_14_, i_13_, i_12_, x908x, x902x}, x1734x);
	defparam lut_9586.LUT_SIZE = 6;
	defparam lut_9586.mask = 64'h77ff77ff07003033;

	lut_sub lut_9592 ({sk[2114], i_14_, i_13_, i_12_, x903x, x897x}, x1733x);
	defparam lut_9592.LUT_SIZE = 6;
	defparam lut_9592.mask = 64'h77ff77ff00003533;

	lut_sub lut_9597 ({sk[2115], n_n1, n_n2, x22513x, x22514x, x1734x, x1733x}, x22518x);
	defparam lut_9597.LUT_SIZE = 7;
	defparam lut_9597.mask = 128'h33ffffff33ffffff00005fff33337fff;

	lut_sub lut_9602 ({sk[2116], i_14_, i_13_, i_12_, i_15_, x907x, n_n282}, x1431x);
	defparam lut_9602.LUT_SIZE = 7;
	defparam lut_9602.mask = 128'h33ffffff33ffffff0037000050335000;

	lut_sub lut_9608 ({sk[2117], x915x, n_n273, n_n283, n_n54, x41x, x1431x}, n_n407);
	defparam lut_9608.LUT_SIZE = 7;
	defparam lut_9608.mask = 128'h33ffffff33ffffff0000000000553f7f;

	lut_sub lut_9612 ({sk[2118], i_7_, i_8_, i_6_, x922x, x123x}, n_n560);
	defparam lut_9612.LUT_SIZE = 6;
	defparam lut_9612.mask = 64'h77ff77ff00100000;

	lut_sub lut_9614 ({sk[2119], i_14_, i_13_, i_12_, x907x, x901x}, x233x);
	defparam lut_9614.LUT_SIZE = 6;
	defparam lut_9614.mask = 64'h77ff77ff00000503;

	lut_sub lut_9617 ({sk[2120], n_n2, n_n6872, n_n6879, x624x, n_n560, x233x}, n_n408);
	defparam lut_9617.LUT_SIZE = 7;
	defparam lut_9617.mask = 128'h33ffffff33ffffff3fffffff7fffffff;

	lut_sub lut_9623 ({sk[2121], n_n1, n_n2, x166x, n_n105, x175x, x229x}, x22524x);
	defparam lut_9623.LUT_SIZE = 7;
	defparam lut_9623.mask = 128'h33ffffff33ffffff00005fff3f3f7fff;

	lut_sub lut_9629 ({sk[2122], n_n356, x2260x, x22518x, n_n407, n_n408, x22524x}, n_n340);
	defparam lut_9629.LUT_SIZE = 7;
	defparam lut_9629.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_9636 ({sk[2123], i_9_, i_10_, i_7_, i_8_, i_6_}, x1316x);
	defparam lut_9636.LUT_SIZE = 6;
	defparam lut_9636.mask = 64'h77ff77ffb2fafafa;

	lut_sub lut_9644 ({sk[2124], i_9_, n_n273, x909x, x19302x, x24215x}, x19303x);
	defparam lut_9644.LUT_SIZE = 6;
	defparam lut_9644.mask = 64'h77ff77ffbbbbbbbf;

	lut_sub lut_9648 ({sk[2125], n_n57, n_n56, x165x, x219x, x189x, x140x}, x19703x);
	defparam lut_9648.LUT_SIZE = 7;
	defparam lut_9648.mask = 128'h33ffffff33ffffff00003f3f55ff7fff;

	lut_sub lut_9653 ({sk[2126], x268x, n_n57, n_n4940, x5325x, n_n4938, x167x}, x19704x);
	defparam lut_9653.LUT_SIZE = 7;
	defparam lut_9653.mask = 128'h33ffffff33ffffff3fff7fff3fffffff;

	lut_sub lut_9659 ({sk[2127], n_n266, n_n271, x909x, x124x, x212x, x190x}, x19709x);
	defparam lut_9659.LUT_SIZE = 7;
	defparam lut_9659.mask = 128'h33ffffff33ffffff0000005f003f007f;

	lut_sub lut_9664 ({sk[2128], n_n56, x49x, x212x, n_n30, x761x, x763x}, x19710x);
	defparam lut_9664.LUT_SIZE = 7;
	defparam lut_9664.mask = 128'h33ffffff33ffffff777777777fffffff;

	lut_sub lut_9670 ({sk[2129], i_14_, i_13_, i_12_, i_15_, x899x, n_n259}, x1319x);
	defparam lut_9670.LUT_SIZE = 7;
	defparam lut_9670.mask = 128'h33ffffff33ffffff0505005555337350;

	lut_sub lut_9681 ({sk[2130], i_14_, i_13_, i_12_, i_15_, x908x, n_n242}, x1318x);
	defparam lut_9681.LUT_SIZE = 7;
	defparam lut_9681.mask = 128'h33ffffff33ffffff0033333377057773;

	lut_sub lut_9694 ({sk[2131], n_n57, n_n56, x165x, x481x, x1319x, x1318x}, x19717x);
	defparam lut_9694.LUT_SIZE = 7;
	defparam lut_9694.mask = 128'h33ffffff33ffffff0f0f5fff3f3f7fff;

	lut_sub lut_9699 ({sk[2132], n_n266, n_n271, n_n12, x909x, x44x, x70x}, x393x);
	defparam lut_9699.LUT_SIZE = 7;
	defparam lut_9699.mask = 128'h33ffffff33ffffff00000707000f070f;

	lut_sub lut_9703 ({sk[2133], i_9_, i_10_, i_11_, i_15_, n_n225, n_n137}, x102x);
	defparam lut_9703.LUT_SIZE = 7;
	defparam lut_9703.mask = 128'h33ffffff33ffffff5050505053505050;

	lut_sub lut_9706 ({sk[2134], i_14_, i_13_, i_12_, i_15_, n_n267}, x98x);
	defparam lut_9706.LUT_SIZE = 6;
	defparam lut_9706.mask = 64'h77ff77ff14040000;

	lut_sub lut_9710 ({sk[2135], n_n283, x914x, x909x, n_n279, x904x}, x21109x);
	defparam lut_9710.LUT_SIZE = 6;
	defparam lut_9710.mask = 64'h77ff77ff00000103;

	lut_sub lut_9713 ({sk[2136], n_n255, n_n31, n_n41, n_n189, n_n54, n_n101}, x24121x);
	defparam lut_9713.LUT_SIZE = 7;
	defparam lut_9713.mask = 128'h33ffffff33fffffffafafafac8000000;

	lut_sub lut_9718 ({sk[2137], i_14_, i_13_, i_12_, x898x, x121x}, x1325x);
	defparam lut_9718.LUT_SIZE = 6;
	defparam lut_9718.mask = 64'h77ff77ff55555557;

	lut_sub lut_9721 ({sk[2138], i_14_, i_13_, i_12_, x905x, x188x}, x1324x);
	defparam lut_9721.LUT_SIZE = 6;
	defparam lut_9721.mask = 64'h77ff77ff57755555;

	lut_sub lut_9725 ({sk[2139], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1946x);
	defparam lut_9725.LUT_SIZE = 7;
	defparam lut_9725.mask = 128'h33ffffff33ffffff0000001050005040;

	lut_sub lut_9732 ({sk[2140], n_n6, n_n186, n_n48, x329x, n_n6512, n_n85}, x21568x);
	defparam lut_9732.LUT_SIZE = 7;
	defparam lut_9732.mask = 128'h33ffffff33ffffff337f337f337fffff;

	lut_sub lut_9737 ({sk[2141], i_14_, i_13_, i_12_, x914x, x912x, x102x}, x1329x);
	defparam lut_9737.LUT_SIZE = 7;
	defparam lut_9737.mask = 128'h33ffffff33ffffff77775f5555555555;

	lut_sub lut_9742 ({sk[2142], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x1328x);
	defparam lut_9742.LUT_SIZE = 7;
	defparam lut_9742.mask = 128'h33ffffff33ffffff0005000500007300;

	lut_sub lut_9747 ({sk[2143], i_14_, i_13_, i_12_, i_15_, n_n242, n_n259}, x1332x);
	defparam lut_9747.LUT_SIZE = 7;
	defparam lut_9747.mask = 128'h33ffffff33ffffff0707700700007500;

	lut_sub lut_9759 ({sk[2144], i_14_, i_13_, i_12_, i_15_, x898x, n_n242}, x1331x);
	defparam lut_9759.LUT_SIZE = 7;
	defparam lut_9759.mask = 128'h33ffffff33ffffff0505730500005500;

	lut_sub lut_9767 ({sk[2145], n_n273, n_n283, n_n220, x922x, x901x, x912x}, x21771x);
	defparam lut_9767.LUT_SIZE = 7;
	defparam lut_9767.mask = 128'h33ffffff33ffffff0000000300070007;

	lut_sub lut_9771 ({sk[2146], n_n220, x898x, n_n48, n_n53, x900x, x897x}, x24100x);
	defparam lut_9771.LUT_SIZE = 7;
	defparam lut_9771.mask = 128'h33ffffff33fffffffffffffffc88fc00;

	lut_sub lut_9776 ({sk[2147], n_n53, n_n8, n_n6521, x1331x, x21771x, x24100x}, x21779x);
	defparam lut_9776.LUT_SIZE = 7;
	defparam lut_9776.mask = 128'h33ffffff33ffffffbbffbbffbfffffff;

	lut_sub lut_9782 ({sk[2148], i_7_, i_8_, i_6_, x60x, x922x}, x4033x);
	defparam lut_9782.LUT_SIZE = 6;
	defparam lut_9782.mask = 64'h77ff77ff10000000;

	lut_sub lut_9784 ({sk[2149], i_14_, i_13_, i_12_, x903x, x897x}, x1333x);
	defparam lut_9784.LUT_SIZE = 6;
	defparam lut_9784.mask = 64'h77ff77ff00000053;

	lut_sub lut_9787 ({sk[2150], i_11_, i_15_, n_n163, n_n94, n_n225, n_n6812}, x22187x);
	defparam lut_9787.LUT_SIZE = 7;
	defparam lut_9787.mask = 128'h33ffffff33ffffff5555555555555557;

	lut_sub lut_9790 ({sk[2151], n_n197, n_n9, n_n227, n_n207, n_n21, n_n59}, x22799x);
	defparam lut_9790.LUT_SIZE = 7;
	defparam lut_9790.mask = 128'h33ffffff33ffffff057705ff05ff05ff;

	lut_sub lut_9796 ({sk[2152], n_n228, x902x, n_n207, n_n6818, x232x, x22799x}, n_n809);
	defparam lut_9796.LUT_SIZE = 7;
	defparam lut_9796.mask = 128'h33ffffff33ffffff5f7f5f7f5f7f5fff;

	lut_sub lut_9801 ({sk[2153], i_14_, i_13_, i_12_, x907x, x901x, x177x}, x1341x);
	defparam lut_9801.LUT_SIZE = 7;
	defparam lut_9801.mask = 128'h33ffffff33ffffff5555557f55775555;

	lut_sub lut_9806 ({sk[2154], i_9_, i_10_, i_11_, i_15_, n_n225}, x145x);
	defparam lut_9806.LUT_SIZE = 6;
	defparam lut_9806.mask = 64'h77ff77ff00005000;

	lut_sub lut_9809 ({sk[2155], i_9_, i_10_, i_11_, i_15_, n_n225}, x1340x);
	defparam lut_9809.LUT_SIZE = 6;
	defparam lut_9809.mask = 64'h77ff77ff50005000;

	lut_sub lut_9814 ({sk[2156], n_n88, n_n94, x368x, n_n6830, n_n6826, x1341x}, x22662x);
	defparam lut_9814.LUT_SIZE = 7;
	defparam lut_9814.mask = 128'h33ffffff33ffffff3f3f7fff3f3fffff;

	lut_sub lut_9820 ({sk[2157], i_14_, i_13_, i_12_, x915x, n_n261, x901x}, x22659x);
	defparam lut_9820.LUT_SIZE = 7;
	defparam lut_9820.mask = 128'h33ffffff33ffffff0000000001010100;

	lut_sub lut_9824 ({sk[2158], n_n100, n_n94, x1929x, x1298x, x1340x, x22659x}, x22663x);
	defparam lut_9824.LUT_SIZE = 7;
	defparam lut_9824.mask = 128'h33ffffff33ffffff55555f5f77ff7fff;

	lut_sub lut_9829 ({sk[2159], n_n103, n_n48, n_n53, x114x, x120x, x91x}, n_n831);
	defparam lut_9829.LUT_SIZE = 7;
	defparam lut_9829.mask = 128'h33ffffff33ffffff000f777f00ffffff;

	lut_sub lut_9835 ({sk[2160], n_n104, x126x, n_n53, n_n4094, n_n6504, n_n4090}, x22708x);
	defparam lut_9835.LUT_SIZE = 7;
	defparam lut_9835.mask = 128'h33ffffff33ffffff7f7f7fff7fff7fff;

	lut_sub lut_9841 ({sk[2161], i_14_, i_13_, i_12_, i_15_, x900x, n_n267}, x408x);
	defparam lut_9841.LUT_SIZE = 7;
	defparam lut_9841.mask = 128'h33ffffff33ffffff0000000000330050;

	lut_sub lut_9844 ({sk[2162], i_7_, i_8_, i_6_, x913x, x916x, n_n258}, x933x);
	defparam lut_9844.LUT_SIZE = 7;
	defparam lut_9844.mask = 128'h33ffffff33ffffff0000000000010000;

	lut_sub lut_9846 ({sk[2163], i_14_, i_13_, i_12_, i_15_, x914x, n_n247}, x22531x);
	defparam lut_9846.LUT_SIZE = 7;
	defparam lut_9846.mask = 128'h33ffffff33ffffff0037000050055050;

	lut_sub lut_9853 ({sk[2164], i_14_, i_13_, i_12_, x907x, x901x}, x414x);
	defparam lut_9853.LUT_SIZE = 6;
	defparam lut_9853.mask = 64'h77ff77ff07003000;

	lut_sub lut_9857 ({sk[2165], i_14_, i_13_, i_12_, i_15_, n_n282, x414x}, x1349x);
	defparam lut_9857.LUT_SIZE = 7;
	defparam lut_9857.mask = 128'h33ffffff33ffffff5555555555777575;

	lut_sub lut_9863 ({sk[2166], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1348x);
	defparam lut_9863.LUT_SIZE = 7;
	defparam lut_9863.mask = 128'h33ffffff33ffffff0005000004010404;

	lut_sub lut_9870 ({sk[2167], n_n208, x916x, n_n3, x408x, x933x, x1348x}, x22533x);
	defparam lut_9870.LUT_SIZE = 7;
	defparam lut_9870.mask = 128'h33ffffff33ffffff333f333f333f777f;

	lut_sub lut_9874 ({sk[2168], i_9_, i_10_, i_11_, i_15_, n_n258}, x403x);
	defparam lut_9874.LUT_SIZE = 6;
	defparam lut_9874.mask = 64'h77ff77ff04004000;

	lut_sub lut_9877 ({sk[2169], n_n265, n_n268, x22531x, x1349x, x403x, x292x}, x22534x);
	defparam lut_9877.LUT_SIZE = 7;
	defparam lut_9877.mask = 128'h33ffffff33ffffff000077ff0f0f7fff;

	lut_sub lut_9882 ({sk[2170], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1351x);
	defparam lut_9882.LUT_SIZE = 7;
	defparam lut_9882.mask = 128'h33ffffff33ffffff0000000040104040;

	lut_sub lut_9887 ({sk[2171], i_14_, i_13_, i_12_, x905x, x899x}, x187x);
	defparam lut_9887.LUT_SIZE = 6;
	defparam lut_9887.mask = 64'h77ff77ff07000000;

	lut_sub lut_9890 ({sk[2172], n_n1, n_n2, n_n216, x142x, x110x, x187x}, x22537x);
	defparam lut_9890.LUT_SIZE = 7;
	defparam lut_9890.mask = 128'h33ffffff33ffffff00003fff7fff7fff;

	lut_sub lut_9898 ({sk[2173], n_n1, n_n2, x140x, x182x, x1351x, x22537x}, n_n354);
	defparam lut_9898.LUT_SIZE = 7;
	defparam lut_9898.mask = 128'h33ffffff33ffffff55557fff77777fff;

	lut_sub lut_9904 ({sk[2174], i_7_, i_8_, i_6_, x915x, n_n240, x403x}, x22539x);
	defparam lut_9904.LUT_SIZE = 7;
	defparam lut_9904.mask = 128'h33ffffff33ffffff0700030000000000;

	lut_sub lut_9908 ({sk[2175], n_n1, n_n2, n_n257, n_n61, n_n236, x22539x}, n_n395);
	defparam lut_9908.LUT_SIZE = 7;
	defparam lut_9908.mask = 128'h33ffffff33ffffff55555fff7fff7fff;

	lut_sub lut_9915 ({sk[2176], i_14_, i_13_, i_12_, i_15_, n_n275, n_n242}, x1358x);
	defparam lut_9915.LUT_SIZE = 7;
	defparam lut_9915.mask = 128'h33ffffff33ffffff0033000030077070;

	lut_sub lut_9925 ({sk[2177], x915x, n_n283, n_n258, x904x, x187x, x22541x}, x22542x);
	defparam lut_9925.LUT_SIZE = 7;
	defparam lut_9925.mask = 128'h33ffffff33ffffff555555555555777f;

	lut_sub lut_9929 ({sk[2178], n_n268, x22533x, x22534x, n_n395, x1358x, x22542x}, x22545x);
	defparam lut_9929.LUT_SIZE = 7;
	defparam lut_9929.mask = 128'h33ffffff33ffffff5fffffff7fffffff;

	lut_sub lut_9935 ({sk[2179], i_14_, i_13_, i_12_, n_n122, x914x}, x757x);
	defparam lut_9935.LUT_SIZE = 6;
	defparam lut_9935.mask = 64'h77ff77ff00100000;

	lut_sub lut_9937 ({sk[2180], n_n41, n_n48, n_n6511, x462x, x464x, x376x}, x20253x);
	defparam lut_9937.LUT_SIZE = 7;
	defparam lut_9937.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_9943 ({sk[2181], n_n48, n_n53, n_n4094, x213x, x470x, x1913x}, x24189x);
	defparam lut_9943.LUT_SIZE = 7;
	defparam lut_9943.mask = 128'h33ffffff33ffffffcc008800c0008000;

	lut_sub lut_9948 ({sk[2182], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1360x);
	defparam lut_9948.LUT_SIZE = 7;
	defparam lut_9948.mask = 128'h33ffffff33ffffff0105000505000404;

	lut_sub lut_9958 ({sk[2183], n_n6878, x475x, x438x, x20386x, n_n6879, x680x}, x21250x);
	defparam lut_9958.LUT_SIZE = 7;
	defparam lut_9958.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_9965 ({sk[2184], x916x, n_n271, n_n3964, x1360x, x21250x}, n_n3914);
	defparam lut_9965.LUT_SIZE = 6;
	defparam lut_9965.mask = 64'h77ff77ff5f5f5f7f;

	lut_sub lut_9969 ({sk[2185], n_n281, n_n208, x916x, x908x, n_n8, x133x}, x21189x);
	defparam lut_9969.LUT_SIZE = 7;
	defparam lut_9969.mask = 128'h33ffffff33ffffff000000770000007f;

	lut_sub lut_9973 ({sk[2186], n_n9, n_n3, n_n7441, n_n61, x208x, n_n7440}, x21192x);
	defparam lut_9973.LUT_SIZE = 7;
	defparam lut_9973.mask = 128'h33ffffff33ffffff55ff7fff55ffffff;

	lut_sub lut_9979 ({sk[2187], n_n281, n_n208, x916x, x903x, x446x, x21192x}, n_n3929);
	defparam lut_9979.LUT_SIZE = 7;
	defparam lut_9979.mask = 128'h33ffffff33ffffff777777777777777f;

	lut_sub lut_9983 ({sk[2188], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1403x);
	defparam lut_9983.LUT_SIZE = 7;
	defparam lut_9983.mask = 128'h33ffffff33ffffff0101000505000504;

	lut_sub lut_9993 ({sk[2189], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x162x);
	defparam lut_9993.LUT_SIZE = 7;
	defparam lut_9993.mask = 128'h33ffffff33ffffff0101000400000000;

	lut_sub lut_9997 ({sk[2190], i_14_, i_13_, i_12_, n_n283, x922x, x908x}, x621x);
	defparam lut_9997.LUT_SIZE = 7;
	defparam lut_9997.mask = 128'h33ffffff33ffffff0001010000000000;

	lut_sub lut_10000 ({sk[2191], i_14_, i_13_, i_12_, i_15_, n_n270}, x1459x);
	defparam lut_10000.LUT_SIZE = 6;
	defparam lut_10000.mask = 64'h77ff77ff11055054;

	lut_sub lut_10010 ({sk[2192], n_n48, n_n53, n_n6860, x162x, x621x, x1459x}, x20263x);
	defparam lut_10010.LUT_SIZE = 7;
	defparam lut_10010.mask = 128'h33ffffff33ffffff33ff3fff77ff7fff;

	lut_sub lut_10015 ({sk[2193], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x203x);
	defparam lut_10015.LUT_SIZE = 7;
	defparam lut_10015.mask = 128'h33ffffff33ffffff0000000104000400;

	lut_sub lut_10019 ({sk[2194], n_n281, x907x, n_n273, n_n220, x922x, x901x}, x882x);
	defparam lut_10019.LUT_SIZE = 7;
	defparam lut_10019.mask = 128'h33ffffff33ffffff0001000100010033;

	lut_sub lut_10022 ({sk[2195], n_n281, x914x, n_n48, n_n6517, n_n6521, x463x}, x20281x);
	defparam lut_10022.LUT_SIZE = 7;
	defparam lut_10022.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_10027 ({sk[2196], n_n258, n_n53, x908x, n_n6878, x882x, x20281x}, x20282x);
	defparam lut_10027.LUT_SIZE = 7;
	defparam lut_10027.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_10032 ({sk[2197], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1536x);
	defparam lut_10032.LUT_SIZE = 7;
	defparam lut_10032.mask = 128'h33ffffff33ffffff1010005050005040;

	lut_sub lut_10042 ({sk[2198], i_7_, i_8_, i_6_, x922x, x62x, x1536x}, x4557x);
	defparam lut_10042.LUT_SIZE = 7;
	defparam lut_10042.mask = 128'h33ffffff33ffffff0000070000000000;

	lut_sub lut_10045 ({sk[2199], i_7_, i_8_, i_6_, n_n216, x922x, x62x}, x24195x);
	defparam lut_10045.LUT_SIZE = 7;
	defparam lut_10045.mask = 128'h33ffffff33ffffffecfffcffffffffff;

	lut_sub lut_10051 ({sk[2200], n_n283, n_n197, x922x, x456x, x1536x, x24195x}, x20288x);
	defparam lut_10051.LUT_SIZE = 7;
	defparam lut_10051.mask = 128'h33ffffff33ffffffafafafafafbfafff;

	lut_sub lut_10056 ({sk[2201], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x20290x);
	defparam lut_10056.LUT_SIZE = 7;
	defparam lut_10056.mask = 128'h33ffffff33ffffff0400010010041040;

	lut_sub lut_10063 ({sk[2202], i_14_, i_13_, i_12_, x906x, x188x}, x20289x);
	defparam lut_10063.LUT_SIZE = 6;
	defparam lut_10063.mask = 64'h77ff77ff75555555;

	lut_sub lut_10066 ({sk[2203], i_14_, i_13_, i_12_, i_15_, n_n259, x20289x}, x20291x);
	defparam lut_10066.LUT_SIZE = 7;
	defparam lut_10066.mask = 128'h33ffffff33ffffff5555555775557555;

	lut_sub lut_10071 ({sk[2204], i_14_, i_13_, i_12_, x900x, x906x}, x1364x);
	defparam lut_10071.LUT_SIZE = 6;
	defparam lut_10071.mask = 64'h77ff77ff50300503;

	lut_sub lut_10076 ({sk[2205], x101x, n_n48, x495x, x561x, x113x, n_n4160}, n_n3980);
	defparam lut_10076.LUT_SIZE = 7;
	defparam lut_10076.mask = 128'h33ffffff33ffffff5fff7fff5fffffff;

	lut_sub lut_10082 ({sk[2206], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x1433x);
	defparam lut_10082.LUT_SIZE = 7;
	defparam lut_10082.mask = 128'h33ffffff33ffffff1010005050005040;

	lut_sub lut_10092 ({sk[2207], i_14_, i_13_, i_12_, i_15_, n_n267, x138x}, x1367x);
	defparam lut_10092.LUT_SIZE = 7;
	defparam lut_10092.mask = 128'h33ffffff33ffffff5575755777557775;

	lut_sub lut_10102 ({sk[2208], i_14_, i_13_, i_12_, i_15_, n_n253, x138x}, x1366x);
	defparam lut_10102.LUT_SIZE = 7;
	defparam lut_10102.mask = 128'h33ffffff33ffffff5757557777557775;

	lut_sub lut_10113 ({sk[2209], i_14_, i_13_, i_12_, i_15_, n_n253, n_n267}, x1369x);
	defparam lut_10113.LUT_SIZE = 7;
	defparam lut_10113.mask = 128'h33ffffff33ffffff0757507000000000;

	lut_sub lut_10122 ({sk[2210], x915x, n_n197, n_n261, x109x, x768x, x117x}, n_n3486);
	defparam lut_10122.LUT_SIZE = 7;
	defparam lut_10122.mask = 128'h33ffffff33ffffff33333333337f33ff;

	lut_sub lut_10127 ({sk[2211], n_n216, n_n100, n_n94, n_n17, n_n6820, x514x}, x20762x);
	defparam lut_10127.LUT_SIZE = 7;
	defparam lut_10127.mask = 128'h33ffffff33ffffff337f337f337fffff;

	lut_sub lut_10132 ({sk[2212], i_7_, i_8_, i_6_, x915x, x188x, n_n1058}, x20763x);
	defparam lut_10132.LUT_SIZE = 7;
	defparam lut_10132.mask = 128'h33ffffff33ffffff5555555555555755;

	lut_sub lut_10135 ({sk[2213], n_n67, n_n216, n_n94, n_n6823, x388x, x701x}, x20764x);
	defparam lut_10135.LUT_SIZE = 7;
	defparam lut_10135.mask = 128'h33ffffff33ffffff7f7f7fff7fff7fff;

	lut_sub lut_10141 ({sk[2214], x392x, x490x, n_n241, n_n216, x386x, n_n3615}, x20770x);
	defparam lut_10141.LUT_SIZE = 7;
	defparam lut_10141.mask = 128'h33ffffff33ffffff777fffffffffffff;

	lut_sub lut_10147 ({sk[2215], n_n3486, x20762x, x20763x, x20764x, x20770x}, x20771x);
	defparam lut_10147.LUT_SIZE = 6;
	defparam lut_10147.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_10153 ({sk[2216], i_7_, i_8_, i_6_, x915x, n_n145, x225x}, n_n2713);
	defparam lut_10153.LUT_SIZE = 7;
	defparam lut_10153.mask = 128'h33ffffff33ffffff0000000005000300;

	lut_sub lut_10156 ({sk[2217], n_n57, n_n258, n_n222, x898x, x45x, x171x}, x370x);
	defparam lut_10156.LUT_SIZE = 7;
	defparam lut_10156.mask = 128'h33ffffff33ffffff00000000777f7f7f;

	lut_sub lut_10161 ({sk[2218], x218x, x911x, n_n228, n_n100, n_n94, x130x}, x493x);
	defparam lut_10161.LUT_SIZE = 7;
	defparam lut_10161.mask = 128'h33ffffff33ffffff1111111f1f1f1f1f;

	lut_sub lut_10165 ({sk[2219], x314x, n_n100, n_n3481, n_n2713, x370x, x493x}, x20782x);
	defparam lut_10165.LUT_SIZE = 7;
	defparam lut_10165.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_10171 ({sk[2220], x915x, n_n197, n_n261, n_n263, x62x, x107x}, x20773x);
	defparam lut_10171.LUT_SIZE = 7;
	defparam lut_10171.mask = 128'h33ffffff33ffffff0000000000770f7f;

	lut_sub lut_10175 ({sk[2221], n_n281, x915x, x905x, n_n263, x314x, x121x}, x20778x);
	defparam lut_10175.LUT_SIZE = 7;
	defparam lut_10175.mask = 128'h33ffffff33ffffff000007070000070f;

	lut_sub lut_10179 ({sk[2222], n_n3212, x20774x, x19564x, x19565x, x20773x, x20778x}, x20783x);
	defparam lut_10179.LUT_SIZE = 7;
	defparam lut_10179.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_10186 ({sk[2223], n_n110, n_n57, n_n56, x60x, x155x, x122x}, x19937x);
	defparam lut_10186.LUT_SIZE = 7;
	defparam lut_10186.mask = 128'h33ffffff33ffffff00777f7f00ff7fff;

	lut_sub lut_10193 ({sk[2224], i_7_, i_8_, i_6_, x909x, n_n42, x68x}, n_n4677);
	defparam lut_10193.LUT_SIZE = 7;
	defparam lut_10193.mask = 128'h33ffffff33ffffff0000000000050003;

	lut_sub lut_10196 ({sk[2225], n_n57, x82x, x111x, x19533x, x19534x, x788x}, x20786x);
	defparam lut_10196.LUT_SIZE = 7;
	defparam lut_10196.mask = 128'h33ffffff33ffffff7f7f7f7f7fffffff;

	lut_sub lut_10202 ({sk[2226], x19937x, n_n4781, x19913x, x19914x, x19932x, x19933x}, x20787x);
	defparam lut_10202.LUT_SIZE = 7;
	defparam lut_10202.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_10209 ({sk[2227], n_n266, n_n271, x909x, x68x, x55x, x788x}, x21080x);
	defparam lut_10209.LUT_SIZE = 7;
	defparam lut_10209.mask = 128'h33ffffff33ffffff5555555f5577557f;

	lut_sub lut_10213 ({sk[2228], n_n56, n_n145, n_n6046, n_n94, x45x, x171x}, x24161x);
	defparam lut_10213.LUT_SIZE = 7;
	defparam lut_10213.mask = 128'h33ffffff33ffffffff00f00088008000;

	lut_sub lut_10218 ({sk[2229], x915x, n_n258, n_n261, x91x, x897x, x1896x}, n_n2928);
	defparam lut_10218.LUT_SIZE = 7;
	defparam lut_10218.mask = 128'h33ffffff33ffffff00000000005f007f;

	lut_sub lut_10222 ({sk[2230], i_14_, i_13_, i_12_, i_15_, n_n253, n_n242}, x1370x);
	defparam lut_10222.LUT_SIZE = 7;
	defparam lut_10222.mask = 128'h33ffffff33ffffff3555535550305003;

	lut_sub lut_10235 ({sk[2231], n_n6, x188x, x411x, x1901x, x1946x, x1370x}, n_n2820);
	defparam lut_10235.LUT_SIZE = 7;
	defparam lut_10235.mask = 128'h33ffffff33ffffff00ff00ff7fffffff;

	lut_sub lut_10241 ({sk[2232], n_n208, x916x, n_n258, x902x, x601x, x382x}, x24201x);
	defparam lut_10241.LUT_SIZE = 7;
	defparam lut_10241.mask = 128'h33ffffff33ffffff8888888888888880;

	lut_sub lut_10246 ({sk[2233], n_n106, n_n100, n_n6843, x391x, x434x, x24201x}, x20374x);
	defparam lut_10246.LUT_SIZE = 7;
	defparam lut_10246.mask = 128'h33ffffff33ffffffbfffbfffbfffffff;

	lut_sub lut_10252 ({sk[2234], x183x, x909x, n_n226, n_n261, x132x, x24133x}, x20381x);
	defparam lut_10252.LUT_SIZE = 7;
	defparam lut_10252.mask = 128'h33ffffff33ffffff00000b0f00000f0f;

	lut_sub lut_10257 ({sk[2235], n_n6, x146x, x159x, x176x, x522x, x1147x}, x20382x);
	defparam lut_10257.LUT_SIZE = 7;
	defparam lut_10257.mask = 128'h33ffffff33ffffff333333337fffffff;

	lut_sub lut_10263 ({sk[2236], n_n93, n_n48, n_n53, x77x, x149x, x253x}, n_n2159);
	defparam lut_10263.LUT_SIZE = 7;
	defparam lut_10263.mask = 128'h33ffffff33ffffff005f337f005fffff;

	lut_sub lut_10268 ({sk[2237], i_14_, i_13_, i_12_, i_15_, x906x, n_n267}, x1376x);
	defparam lut_10268.LUT_SIZE = 7;
	defparam lut_10268.mask = 128'h33ffffff33ffffff0533335055000000;

	lut_sub lut_10275 ({sk[2238], n_n273, n_n283, n_n186, x51x, x922x, x1376x}, n_n2158);
	defparam lut_10275.LUT_SIZE = 7;
	defparam lut_10275.mask = 128'h33ffffff33ffffff0000033311111333;

	lut_sub lut_10279 ({sk[2239], x915x, n_n57, n_n145, n_n261, n_n263, x204x}, x21447x);
	defparam lut_10279.LUT_SIZE = 7;
	defparam lut_10279.mask = 128'h33ffffff33ffffff00005555003f557f;

	lut_sub lut_10283 ({sk[2240], i_9_, i_10_, i_11_, i_15_, n_n279}, x482x);
	defparam lut_10283.LUT_SIZE = 6;
	defparam lut_10283.mask = 64'h77ff77ff00000005;

	lut_sub lut_10286 ({sk[2241], n_n281, x913x, n_n57, x168x, x21447x, x482x}, n_n2172);
	defparam lut_10286.LUT_SIZE = 7;
	defparam lut_10286.mask = 128'h33ffffff33ffffff3377337733773f7f;

	lut_sub lut_10290 ({sk[2242], n_n56, n_n42, n_n6046, x204x, x98x, x482x}, x21453x);
	defparam lut_10290.LUT_SIZE = 7;
	defparam lut_10290.mask = 128'h33ffffff33ffffff00ff00ff7fffffff;

	lut_sub lut_10296 ({sk[2243], n_n281, x915x, n_n261, n_n263, x904x, x906x}, x21455x);
	defparam lut_10296.LUT_SIZE = 7;
	defparam lut_10296.mask = 128'h33ffffff33ffffff0000000000000577;

	lut_sub lut_10300 ({sk[2244], i_9_, i_10_, i_11_, i_15_, n_n281}, x1382x);
	defparam lut_10300.LUT_SIZE = 6;
	defparam lut_10300.mask = 64'h77ff77ff40004404;

	lut_sub lut_10305 ({sk[2245], i_14_, i_13_, i_12_, x913x, x914x}, x21456x);
	defparam lut_10305.LUT_SIZE = 6;
	defparam lut_10305.mask = 64'h77ff77ff53330000;

	lut_sub lut_10310 ({sk[2246], i_14_, i_13_, i_12_, i_15_, n_n242, x21456x}, x1381x);
	defparam lut_10310.LUT_SIZE = 7;
	defparam lut_10310.mask = 128'h33ffffff33ffffff5755555577555555;

	lut_sub lut_10315 ({sk[2247], n_n281, x915x, n_n261, n_n263, x908x, x903x}, x24164x);
	defparam lut_10315.LUT_SIZE = 7;
	defparam lut_10315.mask = 128'h33ffffff33fffffffffffffffffffa88;

	lut_sub lut_10321 ({sk[2248], x915x, n_n263, x528x, n_n2398, x1382x, x24164x}, x21462x);
	defparam lut_10321.LUT_SIZE = 7;
	defparam lut_10321.mask = 128'h33ffffff33ffffffafffafffafffbfff;

	lut_sub lut_10326 ({sk[2249], n_n100, n_n94, x21455x, x1381x, x281x, x338x}, x21463x);
	defparam lut_10326.LUT_SIZE = 7;
	defparam lut_10326.mask = 128'h33ffffff33ffffff00ff77ff0fff7fff;

	lut_sub lut_10331 ({sk[2250], i_14_, i_13_, i_12_, i_15_, n_n247, x329x}, x21464x);
	defparam lut_10331.LUT_SIZE = 7;
	defparam lut_10331.mask = 128'h33ffffff33ffffff5775557555555555;

	lut_sub lut_10336 ({sk[2251], n_n57, n_n56, x252x, n_n32, x205x, x369x}, x24186x);
	defparam lut_10336.LUT_SIZE = 7;
	defparam lut_10336.mask = 128'h33ffffff33ffffff00000f0f7fff7fff;

	lut_sub lut_10346 ({sk[2252], n_n57, n_n56, n_n45, n_n93, n_n42, x98x}, x21452x);
	defparam lut_10346.LUT_SIZE = 7;
	defparam lut_10346.mask = 128'h33ffffff33ffffff00000fff7fff7fff;

	lut_sub lut_10353 ({sk[2253], i_14_, i_13_, i_12_, x908x, x902x}, x360x);
	defparam lut_10353.LUT_SIZE = 6;
	defparam lut_10353.mask = 64'h77ff77ff55300000;

	lut_sub lut_10357 ({sk[2254], i_7_, i_8_, i_6_, x915x, x228x}, x3143x);
	defparam lut_10357.LUT_SIZE = 6;
	defparam lut_10357.mask = 64'h77ff77ff00001000;

	lut_sub lut_10359 ({sk[2255], i_14_, i_13_, i_12_, n_n94, x903x, x897x}, x21857x);
	defparam lut_10359.LUT_SIZE = 7;
	defparam lut_10359.mask = 128'h33ffffff33ffffff0000000500000700;

	lut_sub lut_10363 ({sk[2256], i_14_, i_13_, i_12_, i_15_, x900x, n_n267}, x1386x);
	defparam lut_10363.LUT_SIZE = 7;
	defparam lut_10363.mask = 128'h33ffffff33ffffff3373000550055550;

	lut_sub lut_10373 ({sk[2257], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1385x);
	defparam lut_10373.LUT_SIZE = 7;
	defparam lut_10373.mask = 128'h33ffffff33ffffff0105040104000504;

	lut_sub lut_10383 ({sk[2258], i_14_, i_13_, i_12_, i_15_, n_n253, n_n267}, x1388x);
	defparam lut_10383.LUT_SIZE = 7;
	defparam lut_10383.mask = 128'h33ffffff33ffffff0777300750055550;

	lut_sub lut_10398 ({sk[2259], i_14_, i_13_, i_12_, i_15_, n_n267}, x1387x);
	defparam lut_10398.LUT_SIZE = 6;
	defparam lut_10398.mask = 64'h77ff77ff14400154;

	lut_sub lut_10406 ({sk[2260], x915x, n_n283, n_n62, x456x, x626x, x591x}, x22040x);
	defparam lut_10406.LUT_SIZE = 7;
	defparam lut_10406.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_10411 ({sk[2261], n_n273, x922x, x409x, x42x, x479x, x869x}, x22053x);
	defparam lut_10411.LUT_SIZE = 7;
	defparam lut_10411.mask = 128'h33ffffff33ffffff77ff77ff77ff7fff;

	lut_sub lut_10416 ({sk[2262], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1389x);
	defparam lut_10416.LUT_SIZE = 7;
	defparam lut_10416.mask = 128'h33ffffff33ffffff0000000053000003;

	lut_sub lut_10420 ({sk[2263], n_n3, x993x, x21911x, n_n1159, n_n1160}, x21928x);
	defparam lut_10420.LUT_SIZE = 6;
	defparam lut_10420.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_10425 ({sk[2264], i_14_, i_13_, i_12_, n_n3, x903x}, x3678x);
	defparam lut_10425.LUT_SIZE = 6;
	defparam lut_10425.mask = 64'h77ff77ff01100000;

	lut_sub lut_10428 ({sk[2265], i_14_, i_13_, i_12_, i_15_, n_n275, n_n270}, x1391x);
	defparam lut_10428.LUT_SIZE = 7;
	defparam lut_10428.mask = 128'h33ffffff33ffffff0303000770057570;

	lut_sub lut_10441 ({sk[2266], i_14_, i_13_, i_12_, i_15_, n_n275, x257x}, x1390x);
	defparam lut_10441.LUT_SIZE = 7;
	defparam lut_10441.mask = 128'h33ffffff33ffffff5555555555557775;

	lut_sub lut_10446 ({sk[2267], i_9_, i_10_, i_14_, i_11_, i_15_, n_n254}, x1393x);
	defparam lut_10446.LUT_SIZE = 7;
	defparam lut_10446.mask = 128'h33ffffff33ffffff5040050450400000;

	lut_sub lut_10456 ({sk[2268], n_n57, n_n56, x301x, x254x, x219x, x356x}, x22625x);
	defparam lut_10456.LUT_SIZE = 7;
	defparam lut_10456.mask = 128'h33ffffff33ffffff00005fff33337fff;

	lut_sub lut_10461 ({sk[2269], n_n266, x909x, x277x, n_n4950, x1393x}, x22626x);
	defparam lut_10461.LUT_SIZE = 6;
	defparam lut_10461.mask = 64'h77ff77ff3333337f;

	lut_sub lut_10465 ({sk[2270], i_14_, i_13_, i_12_, x898x, x904x, x202x}, x1697x);
	defparam lut_10465.LUT_SIZE = 7;
	defparam lut_10465.mask = 128'h33ffffff33ffffff5555557f555f5555;

	lut_sub lut_10470 ({sk[2271], n_n9, n_n57, n_n56, n_n11, n_n63, n_n15}, x22638x);
	defparam lut_10470.LUT_SIZE = 7;
	defparam lut_10470.mask = 128'h33ffffff33ffffff007f777f007fffff;

	lut_sub lut_10477 ({sk[2272], n_n53, x571x, x665x, x737x, x1697x, x22638x}, x22640x);
	defparam lut_10477.LUT_SIZE = 7;
	defparam lut_10477.mask = 128'h33ffffff33ffffff5fffffff7fffffff;

	lut_sub lut_10483 ({sk[2273], i_14_, i_13_, i_12_, x902x, x903x, x897x}, x22641x);
	defparam lut_10483.LUT_SIZE = 7;
	defparam lut_10483.mask = 128'h33ffffff33ffffff000000770f0f0f33;

	lut_sub lut_10490 ({sk[2274], i_14_, i_13_, i_12_, x908x, x902x}, x275x);
	defparam lut_10490.LUT_SIZE = 6;
	defparam lut_10490.mask = 64'h77ff77ff00070003;

	lut_sub lut_10494 ({sk[2275], i_14_, i_13_, i_12_, x903x, x897x}, x262x);
	defparam lut_10494.LUT_SIZE = 6;
	defparam lut_10494.mask = 64'h77ff77ff00070003;

	lut_sub lut_10498 ({sk[2276], n_n56, x899x, n_n228, x902x, x309x, x24207x}, n_n838);
	defparam lut_10498.LUT_SIZE = 7;
	defparam lut_10498.mask = 128'h33ffffff33ffffffbbbbbbbbbbbfbbff;

	lut_sub lut_10503 ({sk[2277], n_n57, n_n56, x219x, x190x, x275x, x262x}, x22644x);
	defparam lut_10503.LUT_SIZE = 7;
	defparam lut_10503.mask = 128'h33ffffff33ffffff00000fff77777fff;

	lut_sub lut_10508 ({sk[2278], n_n271, x909x, x304x, n_n4930, n_n4938, x22641x}, x22645x);
	defparam lut_10508.LUT_SIZE = 7;
	defparam lut_10508.mask = 128'h33ffffff33ffffff3f3f3f3f3f3f7fff;

	lut_sub lut_10513 ({sk[2279], n_n57, n_n56, n_n65, n_n11, x275x, x1751x}, x24213x);
	defparam lut_10513.LUT_SIZE = 7;
	defparam lut_10513.mask = 128'h33ffffff33ffffffffff8800a0008000;

	lut_sub lut_10518 ({sk[2280], i_9_, i_10_, i_11_, i_15_, x202x, n_n225}, x1396x);
	defparam lut_10518.LUT_SIZE = 7;
	defparam lut_10518.mask = 128'h33ffffff33ffffff3333337733333377;

	lut_sub lut_10524 ({sk[2281], n_n54, n_n105, n_n100, n_n94, x108x, x139x}, x22667x);
	defparam lut_10524.LUT_SIZE = 7;
	defparam lut_10524.mask = 128'h33ffffff33ffffff053705ff0f3f0fff;

	lut_sub lut_10529 ({sk[2282], n_n103, n_n100, n_n94, x91x, n_n6834, x881x}, x22654x);
	defparam lut_10529.LUT_SIZE = 7;
	defparam lut_10529.mask = 128'h33ffffff33ffffff77777f7f77ffffff;

	lut_sub lut_10535 ({sk[2283], i_14_, i_13_, i_12_, i_11_, x899x, n_n269}, x412x);
	defparam lut_10535.LUT_SIZE = 7;
	defparam lut_10535.mask = 128'h33ffffff33ffffff0000330033005000;

	lut_sub lut_10539 ({sk[2284], i_9_, i_10_, i_12_, i_11_, i_15_, n_n281}, x19252x);
	defparam lut_10539.LUT_SIZE = 7;
	defparam lut_10539.mask = 128'h33ffffff33ffffff000000000fff4fff;

	lut_sub lut_10545 ({sk[2285], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19244x);
	defparam lut_10545.LUT_SIZE = 7;
	defparam lut_10545.mask = 128'h33ffffff33ffffff0000222a00000000;

	lut_sub lut_10548 ({sk[2286], n_n148, n_n163, n_n220, x911x, n_n267, x19244x}, x19256x);
	defparam lut_10548.LUT_SIZE = 7;
	defparam lut_10548.mask = 128'h33ffffff33ffffff777fffffffffffff;

	lut_sub lut_10554 ({sk[2287], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19320x);
	defparam lut_10554.LUT_SIZE = 7;
	defparam lut_10554.mask = 128'h33ffffff33ffffff00007fff0000ffff;

	lut_sub lut_10560 ({sk[2288], n_n208, x916x, n_n258, x900x, n_n228, x906x}, x546x);
	defparam lut_10560.LUT_SIZE = 7;
	defparam lut_10560.mask = 128'h33ffffff33ffffff0000000000000357;

	lut_sub lut_10563 ({sk[2289], n_n208, x916x, n_n220, x900x, n_n7407}, x634x);
	defparam lut_10563.LUT_SIZE = 6;
	defparam lut_10563.mask = 64'h77ff77ff55555557;

	lut_sub lut_10566 ({sk[2290], n_n281, n_n4, n_n9, x905x, n_n258, n_n7406}, x21255x);
	defparam lut_10566.LUT_SIZE = 7;
	defparam lut_10566.mask = 128'h33ffffff33ffffff555557ff55555fff;

	lut_sub lut_10571 ({sk[2291], n_n4, n_n12, n_n7405, x349x, x546x, x634x}, x21257x);
	defparam lut_10571.LUT_SIZE = 7;
	defparam lut_10571.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_10577 ({sk[2292], n_n53, x141x, x736x, x483x, x21255x, x21257x}, n_n3915);
	defparam lut_10577.LUT_SIZE = 7;
	defparam lut_10577.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_10583 ({sk[2293], n_n208, x916x, n_n3, n_n226, x225x, x130x}, x20790x);
	defparam lut_10583.LUT_SIZE = 7;
	defparam lut_10583.mask = 128'h33ffffff33ffffff000f000f000f777f;

	lut_sub lut_10587 ({sk[2294], n_n281, x913x, x183x, n_n3, x20790x}, n_n3406);
	defparam lut_10587.LUT_SIZE = 6;
	defparam lut_10587.mask = 64'h77ff77ff57575777;

	lut_sub lut_10591 ({sk[2295], n_n281, n_n208, x916x, x206x, x914x, n_n63}, x24205x);
	defparam lut_10591.LUT_SIZE = 7;
	defparam lut_10591.mask = 128'h33ffffff33ffffffffffffa0ffffff80;

	lut_sub lut_10596 ({sk[2296], x101x, n_n3, x113x, x24205x}, n_n3932);
	defparam lut_10596.LUT_SIZE = 5;
	defparam lut_10596.mask = 32'h3f3fabaf;

	lut_sub lut_10600 ({sk[2297], n_n281, n_n3, x904x, x409x, x83x, n_n15}, x21199x);
	defparam lut_10600.LUT_SIZE = 7;
	defparam lut_10600.mask = 128'h33ffffff33ffffff0f0f7f7f0f0f7fff;

	lut_sub lut_10605 ({sk[2298], n_n208, x916x, x898x, n_n228, x121x, x21199x}, x21201x);
	defparam lut_10605.LUT_SIZE = 7;
	defparam lut_10605.mask = 128'h33ffffff33ffffff555555555555777f;

	lut_sub lut_10609 ({sk[2299], n_n7402, n_n3, n_n65, x186x, x742x, x546x}, n_n3408);
	defparam lut_10609.LUT_SIZE = 7;
	defparam lut_10609.mask = 128'h33ffffff33ffffff77777fffffffffff;

	lut_sub lut_10615 ({sk[2300], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1408x);
	defparam lut_10615.LUT_SIZE = 7;
	defparam lut_10615.mask = 128'h33ffffff33ffffff1050005050004040;

	lut_sub lut_10625 ({sk[2301], n_n110, n_n4, n_n3, x90x, x82x, n_n3229}, x20793x);
	defparam lut_10625.LUT_SIZE = 7;
	defparam lut_10625.mask = 128'h33ffffff33ffffff55775f7f5577ffff;

	lut_sub lut_10630 ({sk[2302], i_7_, i_8_, i_6_, x916x, n_n3408, x1408x}, x20794x);
	defparam lut_10630.LUT_SIZE = 7;
	defparam lut_10630.mask = 128'h33ffffff33ffffff3337333333333333;

	lut_sub lut_10633 ({sk[2303], i_14_, i_13_, i_12_, i_15_, x60x, n_n242}, x1409x);
	defparam lut_10633.LUT_SIZE = 7;
	defparam lut_10633.mask = 128'h33ffffff33ffffff3777737777337373;

	lut_sub lut_10645 ({sk[2304], n_n4, n_n3, n_n7355, x378x, x1883x, x1409x}, n_n3375);
	defparam lut_10645.LUT_SIZE = 7;
	defparam lut_10645.mask = 128'h33ffffff33ffffff0fff5fff3fff7fff;

	lut_sub lut_10650 ({sk[2305], n_n4, n_n12, n_n7407, n_n7406, n_n7405, x349x}, x633x);
	defparam lut_10650.LUT_SIZE = 7;
	defparam lut_10650.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_10656 ({sk[2306], n_n3, x159x, n_n7441, n_n7440, n_n7442, n_n7443}, x20802x);
	defparam lut_10656.LUT_SIZE = 7;
	defparam lut_10656.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_10662 ({sk[2307], n_n3406, x20793x, x20794x, x633x, x20802x}, x20805x);
	defparam lut_10662.LUT_SIZE = 6;
	defparam lut_10662.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_10668 ({sk[2308], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1950x);
	defparam lut_10668.LUT_SIZE = 7;
	defparam lut_10668.mask = 128'h33ffffff33ffffff0010001050004040;

	lut_sub lut_10675 ({sk[2309], i_14_, i_13_, i_12_, i_15_, n_n247, n_n137}, x1902x);
	defparam lut_10675.LUT_SIZE = 7;
	defparam lut_10675.mask = 128'h33ffffff33ffffff5053505373505070;

	lut_sub lut_10682 ({sk[2310], n_n111, n_n57, x106x, x1861x, x85x, x1902x}, x20489x);
	defparam lut_10682.LUT_SIZE = 7;
	defparam lut_10682.mask = 128'h33ffffff33ffffff00007fff0000ffff;

	lut_sub lut_10688 ({sk[2311], n_n281, x911x, n_n228, x902x, x903x, x118x}, x24124x);
	defparam lut_10688.LUT_SIZE = 7;
	defparam lut_10688.mask = 128'h33ffffff33ffffffaaa0aa0088808800;

	lut_sub lut_10693 ({sk[2312], n_n208, x916x, n_n105, n_n896, x333x, x188x}, x20403x);
	defparam lut_10693.LUT_SIZE = 7;
	defparam lut_10693.mask = 128'h33ffffff33ffffff3f3f3f3f3f3f7fff;

	lut_sub lut_10698 ({sk[2313], n_n208, x916x, x51x, x94x, x138x}, x533x);
	defparam lut_10698.LUT_SIZE = 6;
	defparam lut_10698.mask = 64'h77ff77ff0000007f;

	lut_sub lut_10702 ({sk[2314], x909x, n_n261, x174x, x1905x, x20449x, x20450x}, x20452x);
	defparam lut_10702.LUT_SIZE = 7;
	defparam lut_10702.mask = 128'h33ffffff33ffffff7777777777777fff;

	lut_sub lut_10707 ({sk[2315], x20435x, x20436x, x20442x, x20443x}, x20453x);
	defparam lut_10707.LUT_SIZE = 5;
	defparam lut_10707.mask = 32'h3f3f7fff;

	lut_sub lut_10712 ({sk[2316], n_n57, x20475x, x20457x, x20458x, x1504x, x20469x}, n_n2801);
	defparam lut_10712.LUT_SIZE = 7;
	defparam lut_10712.mask = 128'h33ffffff33ffffff5fffffff7fffffff;

	lut_sub lut_10718 ({sk[2317], n_n53, x695x, x865x, x1948x, x1445x, x20478x}, x20482x);
	defparam lut_10718.LUT_SIZE = 7;
	defparam lut_10718.mask = 128'h33ffffff33ffffff55ffffff7fffffff;

	lut_sub lut_10724 ({sk[2318], x4463x, x20422x, x20430x, x20431x}, x20483x);
	defparam lut_10724.LUT_SIZE = 5;
	defparam lut_10724.mask = 32'h3f3f7fff;

	lut_sub lut_10729 ({sk[2319], n_n266, x206x, x909x, x90x, x258x, n_n6190}, x20495x);
	defparam lut_10729.LUT_SIZE = 7;
	defparam lut_10729.mask = 128'h33ffffff33ffffff55555555557f55ff;

	lut_sub lut_10734 ({sk[2320], n_n57, x155x, x122x, x20490x, x354x, x440x}, x20496x);
	defparam lut_10734.LUT_SIZE = 7;
	defparam lut_10734.mask = 128'h33ffffff33ffffff000000007fffffff;

	lut_sub lut_10740 ({sk[2321], n_n266, x909x, n_n76, x163x, x207x, x1446x}, x20550x);
	defparam lut_10740.LUT_SIZE = 7;
	defparam lut_10740.mask = 128'h33ffffff33ffffff0000000000007fff;

	lut_sub lut_10745 ({sk[2322], n_n57, n_n32, x682x, x46x, x205x, x1950x}, x24127x);
	defparam lut_10745.LUT_SIZE = 7;
	defparam lut_10745.mask = 128'h33ffffff33ffffffff00ff0080000000;

	lut_sub lut_10748 ({sk[2323], x20489x, x20495x, x20496x, x20550x, x24127x}, x20553x);
	defparam lut_10748.LUT_SIZE = 6;
	defparam lut_10748.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_10754 ({sk[2324], x20502x, x20503x, x20508x, x20509x, x4360x, x20516x}, n_n2803);
	defparam lut_10754.LUT_SIZE = 7;
	defparam lut_10754.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_10761 ({sk[2325], x915x, n_n261, x383x, x1321x, n_n2928, n_n2934}, x20544x);
	defparam lut_10761.LUT_SIZE = 7;
	defparam lut_10761.mask = 128'h33ffffff33ffffff77ff77ff77ff7fff;

	lut_sub lut_10766 ({sk[2326], x4344x, x20535x, n_n2927, x20540x}, x20545x);
	defparam lut_10766.LUT_SIZE = 5;
	defparam lut_10766.mask = 32'h3f3f7fff;

	lut_sub lut_10771 ({sk[2327], n_n1, x81x, n_n95, x136x, x98x, x20557x}, x4319x);
	defparam lut_10771.LUT_SIZE = 7;
	defparam lut_10771.mask = 128'h33ffffff33ffffff000000007fffffff;

	lut_sub lut_10777 ({sk[2328], n_n1, n_n111, x106x, x93x, n_n32, x85x}, x20562x);
	defparam lut_10777.LUT_SIZE = 7;
	defparam lut_10777.mask = 128'h33ffffff33ffffff000000007fffffff;

	lut_sub lut_10783 ({sk[2329], n_n1, x163x, n_n3162, x179x, x1623x, x1858x}, x24130x);
	defparam lut_10783.LUT_SIZE = 7;
	defparam lut_10783.mask = 128'h33ffffff33ffffffff00ff0080000000;

	lut_sub lut_10786 ({sk[2330], n_n1, n_n2860, x1949x, x92x, x1953x, x1483x}, x24131x);
	defparam lut_10786.LUT_SIZE = 7;
	defparam lut_10786.mask = 128'h33ffffff33ffffffffff000080000000;

	lut_sub lut_10789 ({sk[2331], x909x, n_n279, n_n263, x67x, x593x, x897x}, x21575x);
	defparam lut_10789.LUT_SIZE = 7;
	defparam lut_10789.mask = 128'h33ffffff33ffffff33333333333f337f;

	lut_sub lut_10793 ({sk[2332], n_n281, n_n208, x916x, n_n3, x904x, x307x}, x21518x);
	defparam lut_10793.LUT_SIZE = 7;
	defparam lut_10793.mask = 128'h33ffffff33ffffff0505050507070737;

	lut_sub lut_10797 ({sk[2333], n_n208, x916x, n_n12, n_n3, x83x, x21518x}, n_n2099);
	defparam lut_10797.LUT_SIZE = 7;
	defparam lut_10797.mask = 128'h33ffffff33ffffff575f575f575f57ff;

	lut_sub lut_10802 ({sk[2334], i_9_, i_10_, i_11_, i_15_, n_n281, n_n279}, x21477x);
	defparam lut_10802.LUT_SIZE = 7;
	defparam lut_10802.mask = 128'h33ffffff33ffffff0007550000570000;

	lut_sub lut_10810 ({sk[2335], i_14_, i_13_, i_12_, i_15_, n_n275, n_n259}, x1413x);
	defparam lut_10810.LUT_SIZE = 7;
	defparam lut_10810.mask = 128'h33ffffff33ffffff0770707077000000;

	lut_sub lut_10823 ({sk[2336], n_n281, x911x, n_n100, n_n94, n_n6813, x1413x}, x21479x);
	defparam lut_10823.LUT_SIZE = 7;
	defparam lut_10823.mask = 128'h33ffffff33ffffff3377337733773f7f;

	lut_sub lut_10827 ({sk[2337], i_14_, i_13_, i_12_, i_15_, n_n253, n_n267}, x1416x);
	defparam lut_10827.LUT_SIZE = 7;
	defparam lut_10827.mask = 128'h33ffffff33ffffff0770707077000000;

	lut_sub lut_10840 ({sk[2338], n_n57, n_n56, n_n22, x264x, x413x, x369x}, x21504x);
	defparam lut_10840.LUT_SIZE = 7;
	defparam lut_10840.mask = 128'h33ffffff33ffffff000055ff3f3f7fff;

	lut_sub lut_10845 ({sk[2339], n_n57, x258x, n_n22, x562x, n_n4924, x46x}, x21505x);
	defparam lut_10845.LUT_SIZE = 7;
	defparam lut_10845.mask = 128'h33ffffff33ffffff3f3f3f3f7fffffff;

	lut_sub lut_10851 ({sk[2340], n_n148, n_n266, n_n271, n_n108, x909x, x1096x}, x21492x);
	defparam lut_10851.LUT_SIZE = 7;
	defparam lut_10851.mask = 128'h33ffffff33ffffff0013001300333333;

	lut_sub lut_10856 ({sk[2341], n_n151, n_n57, n_n56, n_n145, n_n60, x21497x}, x21498x);
	defparam lut_10856.LUT_SIZE = 7;
	defparam lut_10856.mask = 128'h33ffffff33ffffff557f7f7f55ffffff;

	lut_sub lut_10864 ({sk[2342], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x1417x);
	defparam lut_10864.LUT_SIZE = 7;
	defparam lut_10864.mask = 128'h33ffffff33ffffff0144444405000000;

	lut_sub lut_10874 ({sk[2343], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1421x);
	defparam lut_10874.LUT_SIZE = 7;
	defparam lut_10874.mask = 128'h33ffffff33ffffff0053000000535000;

	lut_sub lut_10880 ({sk[2344], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1420x);
	defparam lut_10880.LUT_SIZE = 7;
	defparam lut_10880.mask = 128'h33ffffff33ffffff0053000000530000;

	lut_sub lut_10885 ({sk[2345], i_14_, i_13_, i_12_, i_15_, x902x, n_n270}, x350x);
	defparam lut_10885.LUT_SIZE = 7;
	defparam lut_10885.mask = 128'h33ffffff33ffffff0000000000333350;

	lut_sub lut_10889 ({sk[2346], i_14_, i_13_, i_12_, i_15_, n_n275, x350x}, x1424x);
	defparam lut_10889.LUT_SIZE = 7;
	defparam lut_10889.mask = 128'h33ffffff33ffffff5777755775557575;

	lut_sub lut_10899 ({sk[2347], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x21979x);
	defparam lut_10899.LUT_SIZE = 7;
	defparam lut_10899.mask = 128'h33ffffff33ffffff1050001040004000;

	lut_sub lut_10906 ({sk[2348], n_n1, n_n14, x337x, n_n252, x73x, x21979x}, x2825x);
	defparam lut_10906.LUT_SIZE = 7;
	defparam lut_10906.mask = 128'h33ffffff33ffffff000000007fffffff;

	lut_sub lut_10912 ({sk[2349], i_14_, i_13_, i_12_, x913x, x915x, n_n273}, x5202x);
	defparam lut_10912.LUT_SIZE = 7;
	defparam lut_10912.mask = 128'h33ffffff33ffffff0000010000000000;

	lut_sub lut_10914 ({sk[2350], i_14_, i_13_, i_12_, i_15_, x905x, n_n259}, x21975x);
	defparam lut_10914.LUT_SIZE = 7;
	defparam lut_10914.mask = 128'h33ffffff33ffffff0033330033005050;

	lut_sub lut_10920 ({sk[2351], i_14_, i_13_, i_12_, i_15_, x904x, n_n267}, x21974x);
	defparam lut_10920.LUT_SIZE = 7;
	defparam lut_10920.mask = 128'h33ffffff33ffffff0000050000730000;

	lut_sub lut_10924 ({sk[2352], n_n2, x82x, x100x, x5202x, x21975x, x21974x}, x21981x);
	defparam lut_10924.LUT_SIZE = 7;
	defparam lut_10924.mask = 128'h33ffffff33ffffff0f0f0f0f7fffffff;

	lut_sub lut_10930 ({sk[2353], i_14_, i_13_, i_12_, i_15_, n_n242, n_n270}, x1532x);
	defparam lut_10930.LUT_SIZE = 7;
	defparam lut_10930.mask = 128'h33ffffff33ffffff0777300770037330;

	lut_sub lut_10947 ({sk[2354], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1531x);
	defparam lut_10947.LUT_SIZE = 7;
	defparam lut_10947.mask = 128'h33ffffff33ffffff1050401040004040;

	lut_sub lut_10956 ({sk[2355], n_n1, n_n2, n_n76, x82x, x1532x, x1531x}, n_n1115);
	defparam lut_10956.LUT_SIZE = 7;
	defparam lut_10956.mask = 128'h33ffffff33ffffff000033ff5f5f7fff;

	lut_sub lut_10961 ({sk[2356], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1427x);
	defparam lut_10961.LUT_SIZE = 7;
	defparam lut_10961.mask = 128'h33ffffff33ffffff0300000053000000;

	lut_sub lut_10965 ({sk[2357], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1426x);
	defparam lut_10965.LUT_SIZE = 7;
	defparam lut_10965.mask = 128'h33ffffff33ffffff0000000053000003;

	lut_sub lut_10969 ({sk[2358], i_14_, i_13_, i_12_, i_15_, n_n242, x903x}, x1454x);
	defparam lut_10969.LUT_SIZE = 7;
	defparam lut_10969.mask = 128'h33ffffff33ffffff0377750330033330;

	lut_sub lut_10982 ({sk[2359], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x1453x);
	defparam lut_10982.LUT_SIZE = 7;
	defparam lut_10982.mask = 128'h33ffffff33ffffff0555000550337350;

	lut_sub lut_10992 ({sk[2360], x913x, x907x, n_n265, n_n268, n_n258, x55x}, x24211x);
	defparam lut_10992.LUT_SIZE = 7;
	defparam lut_10992.mask = 128'h33ffffff33fffffffafafac8f8f8f8c8;

	lut_sub lut_10999 ({sk[2361], i_14_, i_13_, i_12_, i_15_, n_n267}, x1428x);
	defparam lut_10999.LUT_SIZE = 6;
	defparam lut_10999.mask = 64'h77ff77ff15414054;

	lut_sub lut_11009 ({sk[2362], i_14_, i_13_, i_12_, i_15_, n_n242, x903x}, x1429x);
	defparam lut_11009.LUT_SIZE = 7;
	defparam lut_11009.mask = 128'h33ffffff33ffffff0000000000033075;

	lut_sub lut_11014 ({sk[2363], n_n6, n_n103, n_n240, n_n227, n_n207, x276x}, x24079x);
	defparam lut_11014.LUT_SIZE = 7;
	defparam lut_11014.mask = 128'h33ffffff33fffffffafac8c8fa00c800;

	lut_sub lut_11023 ({sk[2364], n_n208, x909x, n_n257, n_n263, x1429x, x24079x}, n_n416);
	defparam lut_11023.LUT_SIZE = 7;
	defparam lut_11023.mask = 128'h33ffffff33ffffffaaaaaaafaaaabbbf;

	lut_sub lut_11027 ({sk[2365], i_14_, i_13_, i_12_, i_15_, n_n282, x904x}, x1434x);
	defparam lut_11027.LUT_SIZE = 7;
	defparam lut_11027.mask = 128'h33ffffff33ffffff0377753333003330;

	lut_sub lut_11041 ({sk[2366], i_14_, i_13_, i_12_, i_15_, n_n275, n_n270}, x1436x);
	defparam lut_11041.LUT_SIZE = 7;
	defparam lut_11041.mask = 128'h33ffffff33ffffff0303003337053770;

	lut_sub lut_11055 ({sk[2367], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1435x);
	defparam lut_11055.LUT_SIZE = 7;
	defparam lut_11055.mask = 128'h33ffffff33ffffff0105040505000504;

	lut_sub lut_11067 ({sk[2368], i_14_, i_13_, i_12_, i_15_, n_n247, x1539x}, x1538x);
	defparam lut_11067.LUT_SIZE = 7;
	defparam lut_11067.mask = 128'h33ffffff33ffffff5777757555555555;

	lut_sub lut_11074 ({sk[2369], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x1537x);
	defparam lut_11074.LUT_SIZE = 7;
	defparam lut_11074.mask = 128'h33ffffff33ffffff3355505555055550;

	lut_sub lut_11087 ({sk[2370], i_7_, i_8_, i_6_, x916x, x1538x, x1537x}, n_n3909);
	defparam lut_11087.LUT_SIZE = 7;
	defparam lut_11087.mask = 128'h33ffffff33ffffff0005000300000000;

	lut_sub lut_11090 ({sk[2371], n_n208, x916x, n_n41, n_n3, x476x, x1914x}, x21233x);
	defparam lut_11090.LUT_SIZE = 7;
	defparam lut_11090.mask = 128'h33ffffff33ffffff37373737373737ff;

	lut_sub lut_11094 ({sk[2372], n_n4, n_n3, x115x, n_n54, x213x, x202x}, x21234x);
	defparam lut_11094.LUT_SIZE = 7;
	defparam lut_11094.mask = 128'h33ffffff33ffffff00005f5f33ff7fff;

	lut_sub lut_11099 ({sk[2373], i_14_, i_13_, i_12_, i_15_, n_n275, x897x}, x1441x);
	defparam lut_11099.LUT_SIZE = 7;
	defparam lut_11099.mask = 128'h33ffffff33ffffff0003000333557530;

	lut_sub lut_11108 ({sk[2374], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x20417x);
	defparam lut_11108.LUT_SIZE = 7;
	defparam lut_11108.mask = 128'h33ffffff33ffffff1440014010145040;

	lut_sub lut_11120 ({sk[2375], i_14_, i_13_, i_12_, x898x, x900x, x904x}, x440x);
	defparam lut_11120.LUT_SIZE = 7;
	defparam lut_11120.mask = 128'h33ffffff33ffffff55000f0000000033;

	lut_sub lut_11124 ({sk[2376], n_n110, n_n273, x922x, x70x, x20417x, x440x}, x4463x);
	defparam lut_11124.LUT_SIZE = 7;
	defparam lut_11124.mask = 128'h33ffffff33ffffff0000007f000000ff;

	lut_sub lut_11129 ({sk[2377], n_n281, n_n273, x914x, x922x, x901x, n_n228}, x20418x);
	defparam lut_11129.LUT_SIZE = 7;
	defparam lut_11129.mask = 128'h33ffffff33ffffff000001010000010f;

	lut_sub lut_11132 ({sk[2378], n_n108, x206x, n_n53, x155x, n_n6517, x20418x}, x20422x);
	defparam lut_11132.LUT_SIZE = 7;
	defparam lut_11132.mask = 128'h33ffffff33ffffff777f77ff77ff77ff;

	lut_sub lut_11138 ({sk[2379], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1900x);
	defparam lut_11138.LUT_SIZE = 7;
	defparam lut_11138.mask = 128'h33ffffff33ffffff0010001050004040;

	lut_sub lut_11145 ({sk[2380], i_14_, i_13_, i_12_, i_15_, n_n242, x75x}, x20423x);
	defparam lut_11145.LUT_SIZE = 7;
	defparam lut_11145.mask = 128'h33ffffff33ffffff7555555555555557;

	lut_sub lut_11149 ({sk[2381], i_14_, i_13_, i_12_, x903x, x897x, x20423x}, x1444x);
	defparam lut_11149.LUT_SIZE = 7;
	defparam lut_11149.mask = 128'h33ffffff33ffffff55557755555f5577;

	lut_sub lut_11154 ({sk[2382], n_n7, n_n53, n_n60, x475x, x626x, x1900x}, x20430x);
	defparam lut_11154.LUT_SIZE = 7;
	defparam lut_11154.mask = 128'h33ffffff33ffffff3f3f7fff3f3fffff;

	lut_sub lut_11160 ({sk[2383], i_9_, i_10_, i_11_, n_n261, x922x, n_n6878}, x20424x);
	defparam lut_11160.LUT_SIZE = 7;
	defparam lut_11160.mask = 128'h33ffffff33ffffff5755555555555555;

	lut_sub lut_11163 ({sk[2384], n_n53, x516x, x676x, x882x, x1444x, x20424x}, x20431x);
	defparam lut_11163.LUT_SIZE = 7;
	defparam lut_11163.mask = 128'h33ffffff33ffffff5fffffff7fffffff;

	lut_sub lut_11169 ({sk[2385], x389x, n_n6503, n_n6524, x495x, n_n6517, x882x}, x20449x);
	defparam lut_11169.LUT_SIZE = 7;
	defparam lut_11169.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_11176 ({sk[2386], n_n6, n_n53, x94x, x670x, n_n81, x470x}, x20450x);
	defparam lut_11176.LUT_SIZE = 7;
	defparam lut_11176.mask = 128'h33ffffff33ffffff5f5f7f7f5fff7fff;

	lut_sub lut_11181 ({sk[2387], x909x, n_n258, x115x, n_n261, x901x, x1927x}, x20435x);
	defparam lut_11181.LUT_SIZE = 7;
	defparam lut_11181.mask = 128'h33ffffff33ffffff00000000050f070f;

	lut_sub lut_11185 ({sk[2388], n_n6, n_n41, x51x, x317x, x138x, x221x}, x20436x);
	defparam lut_11185.LUT_SIZE = 7;
	defparam lut_11185.mask = 128'h33ffffff33ffffff0f0f0f0f7fffffff;

	lut_sub lut_11191 ({sk[2389], x78x, x909x, n_n261, x91x, x141x, x181x}, x20442x);
	defparam lut_11191.LUT_SIZE = 7;
	defparam lut_11191.mask = 128'h33ffffff33ffffff0000007f000000ff;

	lut_sub lut_11196 ({sk[2390], n_n6, n_n103, x593x, x1868x, x1904x, x1465x}, x20443x);
	defparam lut_11196.LUT_SIZE = 7;
	defparam lut_11196.mask = 128'h33ffffff33ffffff00ff00ff7fffffff;

	lut_sub lut_11202 ({sk[2391], n_n220, x81x, x904x, x906x, x55x, x20471x}, x24203x);
	defparam lut_11202.LUT_SIZE = 7;
	defparam lut_11202.mask = 128'h33ffffff33ffffff8888000080000000;

	lut_sub lut_11205 ({sk[2392], n_n273, x922x, x136x, x43x, x1280x, x24203x}, x20475x);
	defparam lut_11205.LUT_SIZE = 7;
	defparam lut_11205.mask = 128'h33ffffff33ffffff000000000000bfff;

	lut_sub lut_11210 ({sk[2393], i_14_, i_13_, i_12_, i_15_, n_n53, n_n282}, x20457x);
	defparam lut_11210.LUT_SIZE = 7;
	defparam lut_11210.mask = 128'h33ffffff33ffffff0111101111011110;

	lut_sub lut_11223 ({sk[2394], n_n273, x922x, x869x, x1881x, x1852x}, x20458x);
	defparam lut_11223.LUT_SIZE = 6;
	defparam lut_11223.mask = 64'h77ff77ff0f0f0f7f;

	lut_sub lut_11227 ({sk[2395], n_n148, x101x, x72x, x133x, x113x, x24129x}, x1504x);
	defparam lut_11227.LUT_SIZE = 7;
	defparam lut_11227.mask = 128'h33ffffff33ffffffbfffffffffffffff;

	lut_sub lut_11234 ({sk[2396], x218x, n_n57, n_n53, x68x, x209x, x24128x}, x20469x);
	defparam lut_11234.LUT_SIZE = 7;
	defparam lut_11234.mask = 128'h33ffffff33ffffffaaafbbbfaaafffff;

	lut_sub lut_11239 ({sk[2397], i_14_, i_13_, i_12_, x903x, x897x}, x1948x);
	defparam lut_11239.LUT_SIZE = 6;
	defparam lut_11239.mask = 64'h77ff77ff57073000;

	lut_sub lut_11246 ({sk[2398], i_14_, i_13_, i_12_, i_15_, n_n275, x897x}, x1445x);
	defparam lut_11246.LUT_SIZE = 7;
	defparam lut_11246.mask = 128'h33ffffff33ffffff0000300003557530;

	lut_sub lut_11253 ({sk[2399], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x20490x);
	defparam lut_11253.LUT_SIZE = 7;
	defparam lut_11253.mask = 128'h33ffffff33ffffff0400010000141000;

	lut_sub lut_11259 ({sk[2400], i_14_, i_13_, i_12_, x913x, x898x, x904x}, x354x);
	defparam lut_11259.LUT_SIZE = 7;
	defparam lut_11259.mask = 128'h33ffffff33ffffff00000f0000550033;

	lut_sub lut_11263 ({sk[2401], n_n266, x909x, x81x, n_n42, x55x, x20500x}, x20502x);
	defparam lut_11263.LUT_SIZE = 7;
	defparam lut_11263.mask = 128'h33ffffff33ffffff5555555555557fff;

	lut_sub lut_11268 ({sk[2402], n_n266, x909x, x179x, x43x, x98x, x370x}, x20503x);
	defparam lut_11268.LUT_SIZE = 7;
	defparam lut_11268.mask = 128'h33ffffff33ffffff5555555555557fff;

	lut_sub lut_11273 ({sk[2403], x911x, n_n258, n_n100, x83x, x121x, x107x}, x20508x);
	defparam lut_11273.LUT_SIZE = 7;
	defparam lut_11273.mask = 128'h33ffffff33ffffff007f007f007f00ff;

	lut_sub lut_11278 ({sk[2404], i_7_, i_8_, i_6_, x915x, n_n2926, x1660x}, x20509x);
	defparam lut_11278.LUT_SIZE = 7;
	defparam lut_11278.mask = 128'h33ffffff33ffffff3333333333333733;

	lut_sub lut_11281 ({sk[2405], x915x, n_n261, x176x, x132x, x20511x, x24126x}, x4360x);
	defparam lut_11281.LUT_SIZE = 7;
	defparam lut_11281.mask = 128'h33ffffff33ffffff000000000000bfff;

	lut_sub lut_11286 ({sk[2406], x146x, n_n226, n_n60, n_n100, n_n6843, x1146x}, x20516x);
	defparam lut_11286.LUT_SIZE = 7;
	defparam lut_11286.mask = 128'h33ffffff33ffffff373f3f3f3f3f3f3f;

	lut_sub lut_11292 ({sk[2407], n_n241, n_n103, n_n104, x515x, x872x, x20525x}, n_n2934);
	defparam lut_11292.LUT_SIZE = 7;
	defparam lut_11292.mask = 128'h33ffffff33ffffff7f7f7f7f7fffffff;

	lut_sub lut_11298 ({sk[2408], x915x, x51x, n_n261, x138x, x221x, x24168x}, x4344x);
	defparam lut_11298.LUT_SIZE = 7;
	defparam lut_11298.mask = 128'h33ffffff33ffffff0000000000bf00ff;

	lut_sub lut_11303 ({sk[2409], x907x, n_n279, n_n228, n_n100, x1886x, x20533x}, x20535x);
	defparam lut_11303.LUT_SIZE = 7;
	defparam lut_11303.mask = 128'h33ffffff33ffffff57575757575f5f5f;

	lut_sub lut_11308 ({sk[2410], x915x, n_n258, n_n261, x40x, x899x, x1903x}, n_n2927);
	defparam lut_11308.LUT_SIZE = 7;
	defparam lut_11308.mask = 128'h33ffffff33ffffff00000000005f007f;

	lut_sub lut_11312 ({sk[2411], x907x, n_n220, n_n100, x108x, n_n256, x20539x}, x20540x);
	defparam lut_11312.LUT_SIZE = 7;
	defparam lut_11312.mask = 128'h33ffffff33ffffff555f555f557f55ff;

	lut_sub lut_11317 ({sk[2412], i_14_, i_13_, i_12_, i_15_, x899x, n_n275}, x1446x);
	defparam lut_11317.LUT_SIZE = 7;
	defparam lut_11317.mask = 128'h33ffffff33ffffff0005500555377750;

	lut_sub lut_11329 ({sk[2413], n_n273, n_n279, x922x, x908x, x902x}, x3277x);
	defparam lut_11329.LUT_SIZE = 6;
	defparam lut_11329.mask = 64'h77ff77ff00000007;

	lut_sub lut_11332 ({sk[2414], n_n48, n_n171, x462x, x479x, x478x, x3277x}, n_n2154);
	defparam lut_11332.LUT_SIZE = 7;
	defparam lut_11332.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_11338 ({sk[2415], i_14_, i_13_, i_12_, i_15_, x913x, n_n242}, x1449x);
	defparam lut_11338.LUT_SIZE = 7;
	defparam lut_11338.mask = 128'h33ffffff33ffffff0533335055000000;

	lut_sub lut_11345 ({sk[2416], n_n208, x916x, n_n3, x62x, n_n223, x1449x}, n_n2100);
	defparam lut_11345.LUT_SIZE = 7;
	defparam lut_11345.mask = 128'h33ffffff33ffffff003f003f003f557f;

	lut_sub lut_11349 ({sk[2417], n_n1, n_n2, n_n220, x898x, x900x, x912x}, x21651x);
	defparam lut_11349.LUT_SIZE = 7;
	defparam lut_11349.mask = 128'h33ffffff33ffffff00000033007f007f;

	lut_sub lut_11354 ({sk[2418], i_14_, i_13_, i_12_, i_15_, n_n242, n_n138}, x1473x);
	defparam lut_11354.LUT_SIZE = 7;
	defparam lut_11354.mask = 128'h33ffffff33ffffff5053505070705050;

	lut_sub lut_11359 ({sk[2419], n_n257, n_n227, n_n207, x232x, x350x, x1473x}, x22088x);
	defparam lut_11359.LUT_SIZE = 7;
	defparam lut_11359.mask = 128'h33ffffff33ffffff005f337f005fffff;

	lut_sub lut_11364 ({sk[2420], x374x, x696x, x548x, x434x}, x22075x);
	defparam lut_11364.LUT_SIZE = 5;
	defparam lut_11364.mask = 32'h3f3f7fff;

	lut_sub lut_11369 ({sk[2421], x40x, n_n94, x655x, n_n6818, x380x, x22082x}, x22087x);
	defparam lut_11369.LUT_SIZE = 7;
	defparam lut_11369.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_11375 ({sk[2422], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x1456x);
	defparam lut_11375.LUT_SIZE = 7;
	defparam lut_11375.mask = 128'h33ffffff33ffffff5300000003530000;

	lut_sub lut_11381 ({sk[2423], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1458x);
	defparam lut_11381.LUT_SIZE = 7;
	defparam lut_11381.mask = 128'h33ffffff33ffffff4555155515555555;

	lut_sub lut_11388 ({sk[2424], i_14_, i_13_, i_12_, x900x, x906x}, x1924x);
	defparam lut_11388.LUT_SIZE = 6;
	defparam lut_11388.mask = 64'h77ff77ff03037055;

	lut_sub lut_11395 ({sk[2425], i_14_, i_13_, i_12_, x911x, x903x}, x377x);
	defparam lut_11395.LUT_SIZE = 6;
	defparam lut_11395.mask = 64'h77ff77ff50300003;

	lut_sub lut_11399 ({sk[2426], n_n281, x913x, n_n220, x914x, x106x, x93x}, x24115x);
	defparam lut_11399.LUT_SIZE = 7;
	defparam lut_11399.mask = 128'h33ffffff33ffffff8880888088800000;

	lut_sub lut_11404 ({sk[2427], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1480x);
	defparam lut_11404.LUT_SIZE = 7;
	defparam lut_11404.mask = 128'h33ffffff33ffffff1050005050105040;

	lut_sub lut_11416 ({sk[2428], i_14_, i_13_, i_12_, i_15_, x199x, n_n253}, x1462x);
	defparam lut_11416.LUT_SIZE = 7;
	defparam lut_11416.mask = 128'h33ffffff33ffffff3333373333733337;

	lut_sub lut_11421 ({sk[2429], x146x, x160x, n_n100, n_n94, x4847x, x1462x}, x21090x);
	defparam lut_11421.LUT_SIZE = 7;
	defparam lut_11421.mask = 128'h33ffffff33ffffff373737ff37ff37ff;

	lut_sub lut_11426 ({sk[2430], n_n228, x912x, n_n60, n_n100, n_n94, x500x}, x24165x);
	defparam lut_11426.LUT_SIZE = 7;
	defparam lut_11426.mask = 128'h33ffffff33ffffffaaa0aaa0aaa08880;

	lut_sub lut_11433 ({sk[2431], n_n42, x106x, x131x, x205x, x55x, x178x}, x24204x);
	defparam lut_11433.LUT_SIZE = 7;
	defparam lut_11433.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_11448 ({sk[2432], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1927x);
	defparam lut_11448.LUT_SIZE = 7;
	defparam lut_11448.mask = 128'h33ffffff33ffffff0000001050005040;

	lut_sub lut_11455 ({sk[2433], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x221x);
	defparam lut_11455.LUT_SIZE = 7;
	defparam lut_11455.mask = 128'h33ffffff33ffffff3305005000000000;

	lut_sub lut_11459 ({sk[2434], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1904x);
	defparam lut_11459.LUT_SIZE = 7;
	defparam lut_11459.mask = 128'h33ffffff33ffffff0101000504000400;

	lut_sub lut_11466 ({sk[2435], i_14_, i_13_, i_12_, x899x, x903x}, x1465x);
	defparam lut_11466.LUT_SIZE = 6;
	defparam lut_11466.mask = 64'h77ff77ff05500300;

	lut_sub lut_11470 ({sk[2436], i_14_, i_13_, i_12_, x913x, x90x, x70x}, x1693x);
	defparam lut_11470.LUT_SIZE = 7;
	defparam lut_11470.mask = 128'h33ffffff33ffffff77777f7777777777;

	lut_sub lut_11474 ({sk[2437], i_14_, i_13_, i_12_, i_15_, n_n275, x897x}, x1941x);
	defparam lut_11474.LUT_SIZE = 7;
	defparam lut_11474.mask = 128'h33ffffff33ffffff0000000003557530;

	lut_sub lut_11480 ({sk[2438], i_15_, x911x, n_n258, n_n138, x122x}, x1864x);
	defparam lut_11480.LUT_SIZE = 6;
	defparam lut_11480.mask = 64'h77ff77ff555f777f;

	lut_sub lut_11484 ({sk[2439], i_7_, i_8_, i_6_, x916x, n_n220, x901x}, x605x);
	defparam lut_11484.LUT_SIZE = 7;
	defparam lut_11484.mask = 128'h33ffffff33ffffff0000000000000001;

	lut_sub lut_11486 ({sk[2440], n_n48, n_n53, n_n35, n_n179, n_n113, x470x}, x21595x);
	defparam lut_11486.LUT_SIZE = 7;
	defparam lut_11486.mask = 128'h33ffffff33ffffff555555ff7f7f7fff;

	lut_sub lut_11491 ({sk[2441], i_14_, i_13_, i_12_, i_15_, n_n282, n_n253}, x1470x);
	defparam lut_11491.LUT_SIZE = 7;
	defparam lut_11491.mask = 128'h33ffffff33ffffff0770707073000000;

	lut_sub lut_11503 ({sk[2442], i_14_, i_13_, i_12_, i_15_, x904x, n_n253}, x1471x);
	defparam lut_11503.LUT_SIZE = 7;
	defparam lut_11503.mask = 128'h33ffffff33ffffff0505000533003333;

	lut_sub lut_11510 ({sk[2443], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x22003x);
	defparam lut_11510.LUT_SIZE = 7;
	defparam lut_11510.mask = 128'h33ffffff33ffffff0050030053000000;

	lut_sub lut_11515 ({sk[2444], i_14_, i_13_, i_12_, i_15_, n_n247, x897x}, x22004x);
	defparam lut_11515.LUT_SIZE = 7;
	defparam lut_11515.mask = 128'h33ffffff33ffffff0030750030003030;

	lut_sub lut_11522 ({sk[2445], i_14_, i_13_, i_12_, x915x, n_n263, x897x}, x380x);
	defparam lut_11522.LUT_SIZE = 7;
	defparam lut_11522.mask = 128'h33ffffff33ffffff0101000000000000;

	lut_sub lut_11525 ({sk[2446], i_14_, i_13_, i_12_, x905x, x900x, x73x}, x1476x);
	defparam lut_11525.LUT_SIZE = 7;
	defparam lut_11525.mask = 128'h33ffffff33ffffff555f5f5555555577;

	lut_sub lut_11530 ({sk[2447], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1481x);
	defparam lut_11530.LUT_SIZE = 7;
	defparam lut_11530.mask = 128'h33ffffff33ffffff1050005050105040;

	lut_sub lut_11542 ({sk[2448], i_14_, i_13_, i_12_, x898x, x904x, x171x}, x1877x);
	defparam lut_11542.LUT_SIZE = 7;
	defparam lut_11542.mask = 128'h33ffffff33ffffff555f555f77555555;

	lut_sub lut_11547 ({sk[2449], x559x, n_n241, n_n105, n_n177, n_n200, x524x}, x20525x);
	defparam lut_11547.LUT_SIZE = 7;
	defparam lut_11547.mask = 128'h33ffffff33ffffff575757ffffffffff;

	lut_sub lut_11552 ({sk[2450], i_14_, i_13_, i_12_, x900x, x906x, x55x}, x20557x);
	defparam lut_11552.LUT_SIZE = 7;
	defparam lut_11552.mask = 128'h33ffffff33ffffff555f775f77555555;

	lut_sub lut_11558 ({sk[2451], i_14_, i_13_, i_12_, i_15_, n_n275, x897x}, x1953x);
	defparam lut_11558.LUT_SIZE = 7;
	defparam lut_11558.mask = 128'h33ffffff33ffffff0000000003557530;

	lut_sub lut_11564 ({sk[2452], i_14_, i_13_, i_12_, i_15_, x899x, n_n275}, x1483x);
	defparam lut_11564.LUT_SIZE = 7;
	defparam lut_11564.mask = 128'h33ffffff33ffffff0550505000333300;

	lut_sub lut_11571 ({sk[2453], n_n33, n_n145, n_n280, n_n48, n_n53, x252x}, x21571x);
	defparam lut_11571.LUT_SIZE = 7;
	defparam lut_11571.mask = 128'h33ffffff33ffffff11331f3f33333f3f;

	lut_sub lut_11576 ({sk[2454], i_14_, i_13_, i_12_, i_15_, x902x, n_n275}, x21555x);
	defparam lut_11576.LUT_SIZE = 7;
	defparam lut_11576.mask = 128'h33ffffff33ffffff0550505073000000;

	lut_sub lut_11583 ({sk[2455], i_14_, i_13_, i_12_, i_15_, n_n270, x21555x}, x1487x);
	defparam lut_11583.LUT_SIZE = 7;
	defparam lut_11583.mask = 128'h33ffffff33ffffff5775757575555555;

	lut_sub lut_11590 ({sk[2456], i_14_, i_13_, i_12_, i_15_, x899x, n_n275}, x1486x);
	defparam lut_11590.LUT_SIZE = 7;
	defparam lut_11590.mask = 128'h33ffffff33ffffff0550505077000000;

	lut_sub lut_11598 ({sk[2457], i_14_, i_13_, i_12_, i_15_, n_n282, n_n270}, x1491x);
	defparam lut_11598.LUT_SIZE = 7;
	defparam lut_11598.mask = 128'h33ffffff33ffffff0707000330003070;

	lut_sub lut_11608 ({sk[2458], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x1490x);
	defparam lut_11608.LUT_SIZE = 7;
	defparam lut_11608.mask = 128'h33ffffff33ffffff1050401040005040;

	lut_sub lut_11618 ({sk[2459], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x1493x);
	defparam lut_11618.LUT_SIZE = 7;
	defparam lut_11618.mask = 128'h33ffffff33ffffff0555500550337350;

	lut_sub lut_11629 ({sk[2460], i_14_, i_13_, i_12_, i_15_, x901x, n_n247}, x1492x);
	defparam lut_11629.LUT_SIZE = 7;
	defparam lut_11629.mask = 128'h33ffffff33ffffff0550500000337750;

	lut_sub lut_11638 ({sk[2461], i_14_, i_13_, i_12_, x914x, x115x, x912x}, x1494x);
	defparam lut_11638.LUT_SIZE = 7;
	defparam lut_11638.mask = 128'h33ffffff33ffffff3333337f33333333;

	lut_sub lut_11642 ({sk[2462], i_9_, i_10_, i_14_, i_13_, i_12_, i_11_}, x19347x);
	defparam lut_11642.LUT_SIZE = 7;
	defparam lut_11642.mask = 128'h33ffffff33ffffff00007fff08880000;

	lut_sub lut_11649 ({sk[2463], i_9_, i_10_, i_12_, i_11_}, x19345x);
	defparam lut_11649.LUT_SIZE = 5;
	defparam lut_11649.mask = 32'h3f3f007f;

	lut_sub lut_11653 ({sk[2464], n_n281, x911x, x912x, x19347x, x19345x}, x1500x);
	defparam lut_11653.LUT_SIZE = 6;
	defparam lut_11653.mask = 64'h77ff77ff77777fff;

	lut_sub lut_11658 ({sk[2465], i_9_, i_10_, i_12_, i_11_, i_15_, n_n281}, x19344x);
	defparam lut_11658.LUT_SIZE = 7;
	defparam lut_11658.mask = 128'h33ffffff33ffffff0000000040404fff;

	lut_sub lut_11663 ({sk[2466], i_14_, i_13_, i_12_, i_15_, n_n242, n_n270}, x1502x);
	defparam lut_11663.LUT_SIZE = 7;
	defparam lut_11663.mask = 128'h33ffffff33ffffff0555505773007330;

	lut_sub lut_11678 ({sk[2467], x907x, n_n41, x115x, n_n222, x901x, n_n225}, x24168x);
	defparam lut_11678.LUT_SIZE = 7;
	defparam lut_11678.mask = 128'h33ffffff33ffffffee000000e0000000;

	lut_sub lut_11683 ({sk[2468], i_14_, i_13_, i_12_, x915x, n_n261, x901x}, x20533x);
	defparam lut_11683.LUT_SIZE = 7;
	defparam lut_11683.mask = 128'h33ffffff33ffffff0000000001010100;

	lut_sub lut_11687 ({sk[2469], n_n281, x911x, n_n228, x902x, x903x, x118x}, x24129x);
	defparam lut_11687.LUT_SIZE = 7;
	defparam lut_11687.mask = 128'h33ffffff33ffffffaaa0aa0088808800;

	lut_sub lut_11692 ({sk[2470], i_9_, n_n261, x922x}, x24128x);
	defparam lut_11692.LUT_SIZE = 4;
	defparam lut_11692.mask = 16'h77ef;

	lut_sub lut_11696 ({sk[2471], i_14_, i_13_, i_12_, i_15_, x911x, n_n242}, x1508x);
	defparam lut_11696.LUT_SIZE = 7;
	defparam lut_11696.mask = 128'h33ffffff33ffffff0550505073000000;

	lut_sub lut_11703 ({sk[2472], i_14_, i_13_, i_12_, i_15_, n_n282, n_n247}, x1510x);
	defparam lut_11703.LUT_SIZE = 7;
	defparam lut_11703.mask = 128'h33ffffff33ffffff0730307077000000;

	lut_sub lut_11714 ({sk[2473], i_14_, i_13_, i_12_, i_15_, x906x, n_n253}, x1511x);
	defparam lut_11714.LUT_SIZE = 7;
	defparam lut_11714.mask = 128'h33ffffff33ffffff0573735055000000;

	lut_sub lut_11723 ({sk[2474], i_14_, i_13_, i_12_, i_15_, n_n282, n_n247}, x1513x);
	defparam lut_11723.LUT_SIZE = 7;
	defparam lut_11723.mask = 128'h33ffffff33ffffff0777300770007330;

	lut_sub lut_11739 ({sk[2475], i_14_, i_13_, i_12_, i_15_, n_n247, n_n275}, x1516x);
	defparam lut_11739.LUT_SIZE = 7;
	defparam lut_11739.mask = 128'h33ffffff33ffffff0337000770037770;

	lut_sub lut_11755 ({sk[2476], i_9_, i_10_, i_11_, i_15_, n_n225, x87x}, x1859x);
	defparam lut_11755.LUT_SIZE = 7;
	defparam lut_11755.mask = 128'h33ffffff33ffffff5555555577555555;

	lut_sub lut_11759 ({sk[2477], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x1876x);
	defparam lut_11759.LUT_SIZE = 7;
	defparam lut_11759.mask = 128'h33ffffff33ffffff0000000005337350;

	lut_sub lut_11765 ({sk[2478], i_14_, i_13_, i_12_, i_15_, n_n242, n_n259}, x1524x);
	defparam lut_11765.LUT_SIZE = 7;
	defparam lut_11765.mask = 128'h33ffffff33ffffff0737307555055550;

	lut_sub lut_11781 ({sk[2479], i_14_, i_13_, i_12_, i_15_, x913x, n_n242}, x1523x);
	defparam lut_11781.LUT_SIZE = 7;
	defparam lut_11781.mask = 128'h33ffffff33ffffff0537335555055550;

	lut_sub lut_11794 ({sk[2480], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1529x);
	defparam lut_11794.LUT_SIZE = 7;
	defparam lut_11794.mask = 128'h33ffffff33ffffff0104040404000000;

	lut_sub lut_11800 ({sk[2481], i_14_, i_13_, i_12_, i_15_, n_n275, n_n270}, x1527x);
	defparam lut_11800.LUT_SIZE = 7;
	defparam lut_11800.mask = 128'h33ffffff33ffffff0730307075000000;

	lut_sub lut_11810 ({sk[2482], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x1539x);
	defparam lut_11810.LUT_SIZE = 7;
	defparam lut_11810.mask = 128'h33ffffff33ffffff3305005555055550;

	lut_sub lut_11821 ({sk[2483], i_7_, i_8_, i_6_, x48x, x896x}, x4972x);
	defparam lut_11821.LUT_SIZE = 6;
	defparam lut_11821.mask = 64'h77ff77ff00000100;

	lut_sub lut_11823 ({sk[2484], i_9_, i_10_, i_11_, i_15_, n_n279}, x371x);
	defparam lut_11823.LUT_SIZE = 6;
	defparam lut_11823.mask = 64'h77ff77ff00404000;

	lut_sub lut_11826 ({sk[2485], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, x20190x);
	defparam lut_11826.LUT_SIZE = 7;
	defparam lut_11826.mask = 128'h33ffffff33ffffff0000005000400010;

	lut_sub lut_11831 ({sk[2486], n_n163, n_n130, n_n121, n_n122, n_n109, x371x}, n_n4598);
	defparam lut_11831.LUT_SIZE = 7;
	defparam lut_11831.mask = 128'h33ffffff33ffffff075777770757ffff;

	lut_sub lut_11838 ({sk[2487], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x178x);
	defparam lut_11838.LUT_SIZE = 7;
	defparam lut_11838.mask = 128'h33ffffff33ffffff0000000010004040;

	lut_sub lut_11842 ({sk[2488], i_14_, i_13_, i_12_, i_15_, n_n247, x55x}, x1546x);
	defparam lut_11842.LUT_SIZE = 7;
	defparam lut_11842.mask = 128'h33ffffff33ffffff5557555777557575;

	lut_sub lut_11850 ({sk[2489], n_n56, x538x, x45x, x85x, x204x, x171x}, x20200x);
	defparam lut_11850.LUT_SIZE = 7;
	defparam lut_11850.mask = 128'h33ffffff33ffffff0000ffff7fffffff;

	lut_sub lut_11856 ({sk[2490], n_n57, n_n56, n_n95, x106x, x178x, x1546x}, x20201x);
	defparam lut_11856.LUT_SIZE = 7;
	defparam lut_11856.mask = 128'h33ffffff33ffffff000033ff5f5f7fff;

	lut_sub lut_11861 ({sk[2491], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1761x);
	defparam lut_11861.LUT_SIZE = 7;
	defparam lut_11861.mask = 128'h33ffffff33ffffff0105000505000404;

	lut_sub lut_11871 ({sk[2492], n_n266, n_n271, x909x, n_n32, x205x, x85x}, x20204x);
	defparam lut_11871.LUT_SIZE = 7;
	defparam lut_11871.mask = 128'h33ffffff33ffffff0000000f007f007f;

	lut_sub lut_11876 ({sk[2493], n_n266, n_n271, x909x, x131x, x205x, x178x}, x20205x);
	defparam lut_11876.LUT_SIZE = 7;
	defparam lut_11876.mask = 128'h33ffffff33ffffff0000003f005f007f;

	lut_sub lut_11881 ({sk[2494], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, x871x);
	defparam lut_11881.LUT_SIZE = 7;
	defparam lut_11881.mask = 128'h33ffffff33ffffff1010000000000000;

	lut_sub lut_11884 ({sk[2495], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, x886x);
	defparam lut_11884.LUT_SIZE = 7;
	defparam lut_11884.mask = 128'h33ffffff33ffffff0000000010100000;

	lut_sub lut_11887 ({sk[2496], i_14_, i_13_, i_12_, x903x, x897x}, x1551x);
	defparam lut_11887.LUT_SIZE = 6;
	defparam lut_11887.mask = 64'h77ff77ff33730300;

	lut_sub lut_11894 ({sk[2497], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1554x);
	defparam lut_11894.LUT_SIZE = 7;
	defparam lut_11894.mask = 128'h33ffffff33ffffff0105040504000404;

	lut_sub lut_11904 ({sk[2498], i_14_, i_13_, i_12_, i_15_, n_n275, n_n270}, x1553x);
	defparam lut_11904.LUT_SIZE = 7;
	defparam lut_11904.mask = 128'h33ffffff33ffffff0333303375057570;

	lut_sub lut_11920 ({sk[2499], n_n208, x916x, n_n3, n_n95, x204x, x1578x}, n_n3418);
	defparam lut_11920.LUT_SIZE = 7;
	defparam lut_11920.mask = 128'h33ffffff33ffffff0055005500553f7f;

	lut_sub lut_11924 ({sk[2500], n_n208, x916x, n_n3, n_n105, n_n7225, x1579x}, n_n3417);
	defparam lut_11924.LUT_SIZE = 7;
	defparam lut_11924.mask = 128'h33ffffff33ffffff3377337733773f7f;

	lut_sub lut_11928 ({sk[2501], n_n208, x916x, x68x, x45x, x171x}, x597x);
	defparam lut_11928.LUT_SIZE = 6;
	defparam lut_11928.mask = 64'h77ff77ff0000007f;

	lut_sub lut_11932 ({sk[2502], n_n208, x916x, x170x, x374x, x557x}, x19393x);
	defparam lut_11932.LUT_SIZE = 6;
	defparam lut_11932.mask = 64'h77ff77ff7777777f;

	lut_sub lut_11936 ({sk[2503], n_n1, n_n268, x124x, x190x, x137x, x132x}, x19396x);
	defparam lut_11936.LUT_SIZE = 7;
	defparam lut_11936.mask = 128'h33ffffff33ffffff00000fff77777fff;

	lut_sub lut_11941 ({sk[2504], n_n2, n_n268, x212x, x209x, x1551x, x19395x}, x19397x);
	defparam lut_11941.LUT_SIZE = 7;
	defparam lut_11941.mask = 128'h33ffffff33ffffff000033ff5f5f7fff;

	lut_sub lut_11946 ({sk[2505], n_n208, x916x, n_n236, n_n59, x633x, x132x}, x19405x);
	defparam lut_11946.LUT_SIZE = 7;
	defparam lut_11946.mask = 128'h33ffffff33ffffff3333333333337fff;

	lut_sub lut_11951 ({sk[2506], i_14_, i_13_, i_12_, i_15_, x902x, n_n275}, x19403x);
	defparam lut_11951.LUT_SIZE = 7;
	defparam lut_11951.mask = 128'h33ffffff33ffffff5000050000500037;

	lut_sub lut_11957 ({sk[2507], n_n7424, n_n3, x439x, x648x, x209x, x19403x}, x19406x);
	defparam lut_11957.LUT_SIZE = 7;
	defparam lut_11957.mask = 128'h33ffffff33ffffff0fff7fffffffffff;

	lut_sub lut_11963 ({sk[2508], n_n208, x916x, x92x, x80x, n_n7306, x1941x}, x19413x);
	defparam lut_11963.LUT_SIZE = 7;
	defparam lut_11963.mask = 128'h33ffffff33ffffff3333333333337fff;

	lut_sub lut_11968 ({sk[2509], i_14_, i_13_, i_12_, i_15_, n_n275, x46x}, x1742x);
	defparam lut_11968.LUT_SIZE = 7;
	defparam lut_11968.mask = 128'h33ffffff33ffffff5557755777557575;

	lut_sub lut_11977 ({sk[2510], n_n4, n_n3, n_n76, x163x, x56x, x1742x}, x19414x);
	defparam lut_11977.LUT_SIZE = 7;
	defparam lut_11977.mask = 128'h33ffffff33ffffff000077770fff7fff;

	lut_sub lut_11982 ({sk[2511], i_14_, i_13_, i_12_, i_15_, x902x, n_n270}, x1556x);
	defparam lut_11982.LUT_SIZE = 7;
	defparam lut_11982.mask = 128'h33ffffff33ffffff0555505555337350;

	lut_sub lut_11995 ({sk[2512], i_14_, i_13_, i_12_, i_15_, n_n275, x70x}, x1555x);
	defparam lut_11995.LUT_SIZE = 7;
	defparam lut_11995.mask = 128'h33ffffff33ffffff5775757555555555;

	lut_sub lut_12001 ({sk[2513], x913x, n_n208, x909x, x905x, n_n258, n_n227}, n_n3550);
	defparam lut_12001.LUT_SIZE = 7;
	defparam lut_12001.mask = 128'h33ffffff33ffffff0101010111111133;

	lut_sub lut_12005 ({sk[2514], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1951x);
	defparam lut_12005.LUT_SIZE = 7;
	defparam lut_12005.mask = 128'h33ffffff33ffffff0010001050004040;

	lut_sub lut_12012 ({sk[2515], x915x, n_n273, n_n283, x90x, x111x, x155x}, x20862x);
	defparam lut_12012.LUT_SIZE = 7;
	defparam lut_12012.mask = 128'h33ffffff33ffffff00000000003f5f7f;

	lut_sub lut_12017 ({sk[2516], n_n110, n_n1, n_n2, x82x, x1864x, x1951x}, x20863x);
	defparam lut_12017.LUT_SIZE = 7;
	defparam lut_12017.mask = 128'h33ffffff33ffffff005f337f00ffffff;

	lut_sub lut_12023 ({sk[2517], i_14_, i_13_, i_12_, i_15_, n_n267}, x1559x);
	defparam lut_12023.LUT_SIZE = 6;
	defparam lut_12023.mask = 64'h77ff77ff15455044;

	lut_sub lut_12034 ({sk[2518], n_n273, n_n283, x81x, x922x, n_n95, x179x}, x19509x);
	defparam lut_12034.LUT_SIZE = 7;
	defparam lut_12034.mask = 128'h33ffffff33ffffff0000000f070f070f;

	lut_sub lut_12039 ({sk[2519], n_n48, n_n42, n_n53, x68x, x204x, x98x}, x19512x);
	defparam lut_12039.LUT_SIZE = 7;
	defparam lut_12039.mask = 128'h33ffffff33ffffff005500ff3f7f3fff;

	lut_sub lut_12044 ({sk[2520], n_n273, n_n283, x922x, x43x, x1917x, x19512x}, x19513x);
	defparam lut_12044.LUT_SIZE = 7;
	defparam lut_12044.mask = 128'h33ffffff33ffffff55555577555f557f;

	lut_sub lut_12048 ({sk[2521], n_n6867, x4509x, x393x, x781x, x24197x}, x20835x);
	defparam lut_12048.LUT_SIZE = 6;
	defparam lut_12048.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_12054 ({sk[2522], n_n57, n_n2440, x159x, x741x, x406x, x20835x}, x20836x);
	defparam lut_12054.LUT_SIZE = 7;
	defparam lut_12054.mask = 128'h33ffffff33ffffff7f7fffff7fffffff;

	lut_sub lut_12060 ({sk[2523], i_14_, i_13_, i_12_, x900x, x906x}, x1578x);
	defparam lut_12060.LUT_SIZE = 6;
	defparam lut_12060.mask = 64'h77ff77ff00003375;

	lut_sub lut_12066 ({sk[2524], i_14_, i_13_, i_12_, i_15_, n_n267}, x1579x);
	defparam lut_12066.LUT_SIZE = 6;
	defparam lut_12066.mask = 64'h77ff77ff15454000;

	lut_sub lut_12074 ({sk[2525], x915x, n_n273, x739x, x225x, x130x, n_n3513}, x20810x);
	defparam lut_12074.LUT_SIZE = 7;
	defparam lut_12074.mask = 128'h33ffffff33ffffff55ff55ff55ff7fff;

	lut_sub lut_12079 ({sk[2526], i_14_, i_13_, i_12_, i_15_, x913x, n_n242}, x1616x);
	defparam lut_12079.LUT_SIZE = 7;
	defparam lut_12079.mask = 128'h33ffffff33ffffff5033373355055555;

	lut_sub lut_12092 ({sk[2527], i_14_, i_13_, i_12_, i_15_, x159x, n_n242}, x1615x);
	defparam lut_12092.LUT_SIZE = 7;
	defparam lut_12092.mask = 128'h33ffffff33ffffff7333373333733337;

	lut_sub lut_12098 ({sk[2528], x915x, n_n283, x916x, n_n271, x1616x, x1615x}, x20811x);
	defparam lut_12098.LUT_SIZE = 7;
	defparam lut_12098.mask = 128'h33ffffff33ffffff0003000300035557;

	lut_sub lut_12101 ({sk[2529], x248x, n_n222, n_n53, x901x, n_n6503, n_n6505}, x24191x);
	defparam lut_12101.LUT_SIZE = 7;
	defparam lut_12101.mask = 128'h33ffffff33ffffff8888888088008800;

	lut_sub lut_12105 ({sk[2530], n_n273, n_n283, n_n280, x922x, n_n32, x24191x}, n_n1781);
	defparam lut_12105.LUT_SIZE = 7;
	defparam lut_12105.mask = 128'h33ffffff33ffffffaaaaabafaaafabaf;

	lut_sub lut_12110 ({sk[2531], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x1562x);
	defparam lut_12110.LUT_SIZE = 7;
	defparam lut_12110.mask = 128'h33ffffff33ffffff0005000500007300;

	lut_sub lut_12115 ({sk[2532], n_n273, n_n283, x922x, x263x, x313x, x1562x}, n_n1782);
	defparam lut_12115.LUT_SIZE = 7;
	defparam lut_12115.mask = 128'h33ffffff33ffffff00000055003f007f;

	lut_sub lut_12119 ({sk[2533], n_n208, x916x, n_n3, n_n896, x1915x, x139x}, n_n785);
	defparam lut_12119.LUT_SIZE = 7;
	defparam lut_12119.mask = 128'h33ffffff33ffffff0f3f0f3f0f3f5f7f;

	lut_sub lut_12123 ({sk[2534], i_14_, i_13_, i_12_, i_15_, n_n242, x227x}, x22752x);
	defparam lut_12123.LUT_SIZE = 7;
	defparam lut_12123.mask = 128'h33ffffff33ffffff5555557757575775;

	lut_sub lut_12131 ({sk[2535], i_14_, i_13_, i_12_, i_15_, n_n242, n_n270}, x1566x);
	defparam lut_12131.LUT_SIZE = 7;
	defparam lut_12131.mask = 128'h33ffffff33ffffff0000007707070770;

	lut_sub lut_12144 ({sk[2536], n_n1, n_n2, x305x, x262x, x22752x, x1566x}, n_n751);
	defparam lut_12144.LUT_SIZE = 7;
	defparam lut_12144.mask = 128'h33ffffff33ffffff000055553fff7fff;

	lut_sub lut_12149 ({sk[2537], i_14_, i_13_, i_12_, x898x, x901x, x904x}, x22756x);
	defparam lut_12149.LUT_SIZE = 7;
	defparam lut_12149.mask = 128'h33ffffff33ffffff0000005f33333355;

	lut_sub lut_12156 ({sk[2538], i_14_, i_13_, i_12_, i_15_, n_n247, x219x}, x22754x);
	defparam lut_12156.LUT_SIZE = 7;
	defparam lut_12156.mask = 128'h33ffffff33ffffff5555557755555575;

	lut_sub lut_12161 ({sk[2539], i_14_, i_13_, i_12_, i_15_, n_n267, x22754x}, x1568x);
	defparam lut_12161.LUT_SIZE = 7;
	defparam lut_12161.mask = 128'h33ffffff33ffffff5555557757575775;

	lut_sub lut_12169 ({sk[2540], i_14_, i_13_, i_12_, x907x, x898x, x901x}, x22755x);
	defparam lut_12169.LUT_SIZE = 7;
	defparam lut_12169.mask = 128'h33ffffff33ffffff0000005f3333330f;

	lut_sub lut_12176 ({sk[2541], n_n1, n_n2, x335x, x22756x, x1568x, x22755x}, n_n753);
	defparam lut_12176.LUT_SIZE = 7;
	defparam lut_12176.mask = 128'h33ffffff33ffffff00005fff33337fff;

	lut_sub lut_12181 ({sk[2542], i_14_, i_13_, i_12_, x902x, x897x}, x22761x);
	defparam lut_12181.LUT_SIZE = 6;
	defparam lut_12181.mask = 64'h77ff77ff00007770;

	lut_sub lut_12188 ({sk[2543], i_14_, i_13_, i_12_, i_15_, n_n282, x275x}, x22762x);
	defparam lut_12188.LUT_SIZE = 7;
	defparam lut_12188.mask = 128'h33ffffff33ffffff5555557757575775;

	lut_sub lut_12196 ({sk[2544], i_14_, i_13_, i_12_, i_15_, n_n247, n_n275}, x1570x);
	defparam lut_12196.LUT_SIZE = 7;
	defparam lut_12196.mask = 128'h33ffffff33ffffff0000007707070770;

	lut_sub lut_12209 ({sk[2545], x915x, n_n273, n_n283, x22761x, x22762x, x1570x}, x22763x);
	defparam lut_12209.LUT_SIZE = 7;
	defparam lut_12209.mask = 128'h33ffffff33ffffff0000000000553f7f;

	lut_sub lut_12213 ({sk[2546], x915x, n_n263, n_n236, n_n6835, x825x, n_n6829}, x22550x);
	defparam lut_12213.LUT_SIZE = 7;
	defparam lut_12213.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_12218 ({sk[2547], i_14_, i_13_, i_12_, x915x, n_n263, x903x}, x471x);
	defparam lut_12218.LUT_SIZE = 7;
	defparam lut_12218.mask = 128'h33ffffff33ffffff0000000001000100;

	lut_sub lut_12221 ({sk[2548], x915x, n_n263, x903x, n_n256, x897x}, x658x);
	defparam lut_12221.LUT_SIZE = 6;
	defparam lut_12221.mask = 64'h77ff77ff00000013;

	lut_sub lut_12224 ({sk[2549], n_n208, x916x, n_n257, n_n227, x312x, x743x}, x22557x);
	defparam lut_12224.LUT_SIZE = 7;
	defparam lut_12224.mask = 128'h33ffffff33ffffff555f555f555f777f;

	lut_sub lut_12228 ({sk[2550], x913x, n_n258, x278x, x642x, x471x, x658x}, x22558x);
	defparam lut_12228.LUT_SIZE = 7;
	defparam lut_12228.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_12233 ({sk[2551], n_n6843, x500x, n_n6830, n_n7306, x480x, n_n6824}, x24080x);
	defparam lut_12233.LUT_SIZE = 7;
	defparam lut_12233.mask = 128'h33ffffff33ffffff8000000000000000;

	lut_sub lut_12235 ({sk[2552], x434x, x22550x, x22557x, x22558x, x24080x}, n_n359);
	defparam lut_12235.LUT_SIZE = 6;
	defparam lut_12235.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_12241 ({sk[2553], i_14_, i_13_, i_12_, i_15_, x163x, n_n270}, x1937x);
	defparam lut_12241.LUT_SIZE = 7;
	defparam lut_12241.mask = 128'h33ffffff33ffffff3333333337337373;

	lut_sub lut_12246 ({sk[2554], i_14_, i_13_, i_12_, i_11_, i_15_, x923x}, x1945x);
	defparam lut_12246.LUT_SIZE = 7;
	defparam lut_12246.mask = 128'h33ffffff33ffffff1050005040000000;

	lut_sub lut_12253 ({sk[2555], i_14_, i_13_, i_12_, x907x, x901x}, x1944x);
	defparam lut_12253.LUT_SIZE = 6;
	defparam lut_12253.mask = 64'h77ff77ff53330000;

	lut_sub lut_12258 ({sk[2556], i_9_, i_10_, i_11_, i_15_, n_n279}, x1797x);
	defparam lut_12258.LUT_SIZE = 6;
	defparam lut_12258.mask = 64'h77ff77ff00404040;

	lut_sub lut_12262 ({sk[2557], n_n139, n_n152, n_n163, n_n6036, n_n6035, x1797x}, n_n4596);
	defparam lut_12262.LUT_SIZE = 7;
	defparam lut_12262.mask = 128'h33ffffff33ffffff3f3f7f7f7fff7fff;

	lut_sub lut_12268 ({sk[2558], i_7_, i_8_, i_6_, n_n165, n_n284, x896x}, x1576x);
	defparam lut_12268.LUT_SIZE = 7;
	defparam lut_12268.mask = 128'h33ffffff33ffffff5703000000000000;

	lut_sub lut_12272 ({sk[2559], n_n266, x909x, n_n109, x171x, x371x, x1576x}, x20215x);
	defparam lut_12272.LUT_SIZE = 7;
	defparam lut_12272.mask = 128'h33ffffff33ffffff1155115511551f5f;

	lut_sub lut_12276 ({sk[2560], n_n271, x909x, x179x, n_n4681, x43x, x98x}, x20220x);
	defparam lut_12276.LUT_SIZE = 7;
	defparam lut_12276.mask = 128'h33ffffff33ffffff0f0f0f0f0f0f7fff;

	lut_sub lut_12281 ({sk[2561], n_n57, n_n56, x81x, n_n6046, x43x, x98x}, x20219x);
	defparam lut_12281.LUT_SIZE = 7;
	defparam lut_12281.mask = 128'h33ffffff33ffffff0f0f0fff7f7f7fff;

	lut_sub lut_12286 ({sk[2562], n_n283, x170x, x922x, x163x, x49x, n_n3579}, x19489x);
	defparam lut_12286.LUT_SIZE = 7;
	defparam lut_12286.mask = 128'h33ffffff33ffffff55555555557f55ff;

	lut_sub lut_12291 ({sk[2563], n_n48, n_n53, n_n22, x70x, x1930x, n_n3457}, x19490x);
	defparam lut_12291.LUT_SIZE = 7;
	defparam lut_12291.mask = 128'h33ffffff33ffffff55555fff77777fff;

	lut_sub lut_12296 ({sk[2564], i_14_, i_13_, i_12_, i_15_, n_n275, x46x}, x1583x);
	defparam lut_12296.LUT_SIZE = 7;
	defparam lut_12296.mask = 128'h33ffffff33ffffff5557555777577775;

	lut_sub lut_12306 ({sk[2565], n_n48, n_n53, n_n22, x147x, x56x, x1583x}, x19503x);
	defparam lut_12306.LUT_SIZE = 7;
	defparam lut_12306.mask = 128'h33ffffff33ffffff00003f3f55ff7fff;

	lut_sub lut_12311 ({sk[2566], n_n9, n_n7, n_n48, x44x, x209x, x133x}, x5607x);
	defparam lut_12311.LUT_SIZE = 7;
	defparam lut_12311.mask = 128'h33ffffff33ffffff007f00ff00ff00ff;

	lut_sub lut_12317 ({sk[2567], n_n53, n_n60, n_n6878, x626x, x137x, x132x}, x19495x);
	defparam lut_12317.LUT_SIZE = 7;
	defparam lut_12317.mask = 128'h33ffffff33ffffff0fff0fff7fffffff;

	lut_sub lut_12323 ({sk[2568], i_7_, i_8_, i_6_, x915x, x44x}, x5721x);
	defparam lut_12323.LUT_SIZE = 6;
	defparam lut_12323.mask = 64'h77ff77ff00100000;

	lut_sub lut_12325 ({sk[2569], i_14_, i_13_, i_12_, i_15_, x900x, n_n267}, x1867x);
	defparam lut_12325.LUT_SIZE = 7;
	defparam lut_12325.mask = 128'h33ffffff33ffffff5000050000500033;

	lut_sub lut_12330 ({sk[2570], i_7_, i_8_, i_6_, n_n281, x915x, x906x}, x5710x);
	defparam lut_12330.LUT_SIZE = 7;
	defparam lut_12330.mask = 128'h33ffffff33ffffff0000010000000000;

	lut_sub lut_12332 ({sk[2571], x909x, n_n261, n_n263, x1619x, x1618x, x217x}, n_n3388);
	defparam lut_12332.LUT_SIZE = 7;
	defparam lut_12332.mask = 128'h33ffffff33ffffff0000000000335f7f;

	lut_sub lut_12336 ({sk[2572], n_n5, x904x, n_n225, x77x, x411x, x217x}, x20842x);
	defparam lut_12336.LUT_SIZE = 7;
	defparam lut_12336.mask = 128'h33ffffff33ffffff333333337f7f7fff;

	lut_sub lut_12341 ({sk[2573], x909x, n_n261, n_n263, x99x, x1907x, x1620x}, x20843x);
	defparam lut_12341.LUT_SIZE = 7;
	defparam lut_12341.mask = 128'h33ffffff33ffffff00000000003f557f;

	lut_sub lut_12345 ({sk[2574], n_n4773, n_n4772, x19485x, n_n3388, x20842x, x20843x}, n_n3367);
	defparam lut_12345.LUT_SIZE = 7;
	defparam lut_12345.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_12352 ({sk[2575], n_n108, n_n53, n_n6870, x155x, x4033x, x286x}, x20849x);
	defparam lut_12352.LUT_SIZE = 7;
	defparam lut_12352.mask = 128'h33ffffff33ffffff77ff7fff77ffffff;

	lut_sub lut_12358 ({sk[2576], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1656x);
	defparam lut_12358.LUT_SIZE = 7;
	defparam lut_12358.mask = 128'h33ffffff33ffffff1040004010004040;

	lut_sub lut_12365 ({sk[2577], i_14_, i_13_, i_12_, i_15_, x913x, n_n242}, x20846x);
	defparam lut_12365.LUT_SIZE = 7;
	defparam lut_12365.mask = 128'h33ffffff33ffffff0005330550000000;

	lut_sub lut_12370 ({sk[2578], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1654x);
	defparam lut_12370.LUT_SIZE = 7;
	defparam lut_12370.mask = 128'h33ffffff33ffffff1040004010105040;

	lut_sub lut_12379 ({sk[2579], n_n273, n_n283, x922x, x1656x, x20846x, x1654x}, x20850x);
	defparam lut_12379.LUT_SIZE = 7;
	defparam lut_12379.mask = 128'h33ffffff33ffffff0000003f0055007f;

	lut_sub lut_12383 ({sk[2580], x183x, n_n48, x44x, x474x, n_n4774, x20853x}, x20856x);
	defparam lut_12383.LUT_SIZE = 7;
	defparam lut_12383.mask = 128'h33ffffff33ffffff7f7f7fff7f7fffff;

	lut_sub lut_12389 ({sk[2581], n_n3457, x20823x, x20849x, x20850x, x20822x}, x20857x);
	defparam lut_12389.LUT_SIZE = 6;
	defparam lut_12389.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_12395 ({sk[2582], n_n151, n_n266, x909x, n_n95, n_n100, x204x}, x20500x);
	defparam lut_12395.LUT_SIZE = 7;
	defparam lut_12395.mask = 128'h33ffffff33ffffff0000005f3333337f;

	lut_sub lut_12399 ({sk[2583], n_n106, n_n1, n_n2, x101x, x265x, x293x}, n_n2589);
	defparam lut_12399.LUT_SIZE = 7;
	defparam lut_12399.mask = 128'h33ffffff33ffffff00553f7f00ff3fff;

	lut_sub lut_12404 ({sk[2584], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1591x);
	defparam lut_12404.LUT_SIZE = 7;
	defparam lut_12404.mask = 128'h33ffffff33ffffff0105000505000404;

	lut_sub lut_12414 ({sk[2585], x915x, n_n273, n_n283, n_n111, x106x, x1858x}, x19770x);
	defparam lut_12414.LUT_SIZE = 7;
	defparam lut_12414.mask = 128'h33ffffff33ffffff00000000003f557f;

	lut_sub lut_12418 ({sk[2586], i_14_, i_13_, i_12_, i_15_, n_n253, x363x}, x1592x);
	defparam lut_12418.LUT_SIZE = 7;
	defparam lut_12418.mask = 128'h33ffffff33ffffff5555555755557755;

	lut_sub lut_12423 ({sk[2587], x917x, x266x, x294x, n_n283, n_n100, x1592x}, x21864x);
	defparam lut_12423.LUT_SIZE = 7;
	defparam lut_12423.mask = 128'h33ffffff33ffffff11111111111f1f1f;

	lut_sub lut_12427 ({sk[2588], i_14_, i_13_, i_12_, i_15_, n_n253, n_n267}, x1595x);
	defparam lut_12427.LUT_SIZE = 7;
	defparam lut_12427.mask = 128'h33ffffff33ffffff0707700700007300;

	lut_sub lut_12439 ({sk[2589], i_14_, i_13_, i_12_, i_15_, n_n267, n_n137}, x1594x);
	defparam lut_12439.LUT_SIZE = 7;
	defparam lut_12439.mask = 128'h33ffffff33ffffff0707350705053705;

	lut_sub lut_12447 ({sk[2590], n_n266, x909x, n_n222, n_n48, x900x, n_n150}, x24095x);
	defparam lut_12447.LUT_SIZE = 7;
	defparam lut_12447.mask = 128'h33ffffff33fffffffffcfffcfffcaaa8;

	lut_sub lut_12457 ({sk[2591], n_n56, n_n53, n_n144, x1286x, x1594x, x24095x}, x21839x);
	defparam lut_12457.LUT_SIZE = 7;
	defparam lut_12457.mask = 128'h33ffffff33ffffffaaaabfbfaaffbfff;

	lut_sub lut_12462 ({sk[2592], i_14_, i_13_, i_12_, x913x, x911x}, x195x);
	defparam lut_12462.LUT_SIZE = 6;
	defparam lut_12462.mask = 64'h77ff77ff50300000;

	lut_sub lut_12465 ({sk[2593], n_n62, n_n14, n_n147, n_n17, n_n8, x195x}, x1597x);
	defparam lut_12465.LUT_SIZE = 7;
	defparam lut_12465.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_12472 ({sk[2594], i_14_, i_13_, i_12_, x905x, x899x}, x240x);
	defparam lut_12472.LUT_SIZE = 6;
	defparam lut_12472.mask = 64'h77ff77ff00050070;

	lut_sub lut_12476 ({sk[2595], n_n220, x900x, x912x, n_n94, x168x, n_n1798}, x21752x);
	defparam lut_12476.LUT_SIZE = 7;
	defparam lut_12476.mask = 128'h33ffffff33ffffff55555555555f777f;

	lut_sub lut_12480 ({sk[2596], i_14_, i_13_, i_12_, i_15_, n_n259, x857x}, x1599x);
	defparam lut_12480.LUT_SIZE = 7;
	defparam lut_12480.mask = 128'h33ffffff33ffffff5757755755557755;

	lut_sub lut_12488 ({sk[2597], n_n281, x911x, n_n94, n_n256, n_n6818, n_n6823}, x24206x);
	defparam lut_12488.LUT_SIZE = 7;
	defparam lut_12488.mask = 128'h33ffffff33ffffff7777777f777777ff;

	lut_sub lut_12500 ({sk[2598], i_15_, n_n94, n_n138, n_n6820, x360x, x24206x}, x21759x);
	defparam lut_12500.LUT_SIZE = 7;
	defparam lut_12500.mask = 128'h33ffffff33ffffff5f5f7fff5f5f7f7f;

	lut_sub lut_12505 ({sk[2599], i_14_, i_13_, i_12_, i_15_, n_n270, x379x}, x236x);
	defparam lut_12505.LUT_SIZE = 7;
	defparam lut_12505.mask = 128'h33ffffff33ffffff5555555755555555;

	lut_sub lut_12508 ({sk[2600], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1730x);
	defparam lut_12508.LUT_SIZE = 7;
	defparam lut_12508.mask = 128'h33ffffff33ffffff0101040100000500;

	lut_sub lut_12515 ({sk[2601], x915x, n_n261, n_n263, x1599x, x236x, x1730x}, x21760x);
	defparam lut_12515.LUT_SIZE = 7;
	defparam lut_12515.mask = 128'h33ffffff33ffffff0000000000335f7f;

	lut_sub lut_12519 ({sk[2602], i_9_, i_10_, i_11_, i_15_, n_n222}, x494x);
	defparam lut_12519.LUT_SIZE = 6;
	defparam lut_12519.mask = 64'h77ff77ff00050000;

	lut_sub lut_12522 ({sk[2603], i_9_, i_10_, i_11_, i_15_, n_n222}, x172x);
	defparam lut_12522.LUT_SIZE = 6;
	defparam lut_12522.mask = 64'h77ff77ff00000005;

	lut_sub lut_12525 ({sk[2604], n_n56, x99x, n_n42, n_n4952, x24102x, x24159x}, x24166x);
	defparam lut_12525.LUT_SIZE = 7;
	defparam lut_12525.mask = 128'h33ffffff33ffffff1010101010000000;

	lut_sub lut_12528 ({sk[2605], n_n220, x898x, x901x, n_n94, x237x, x240x}, x3066x);
	defparam lut_12528.LUT_SIZE = 7;
	defparam lut_12528.mask = 128'h33ffffff33ffffff07070707070f0f0f;

	lut_sub lut_12533 ({sk[2606], i_9_, i_10_, i_14_, i_11_, i_15_, n_n254}, x1602x);
	defparam lut_12533.LUT_SIZE = 7;
	defparam lut_12533.mask = 128'h33ffffff33ffffff0001001040100000;

	lut_sub lut_12538 ({sk[2607], n_n208, x916x, n_n258, x898x, x202x}, x862x);
	defparam lut_12538.LUT_SIZE = 6;
	defparam lut_12538.mask = 64'h77ff77ff00000057;

	lut_sub lut_12541 ({sk[2608], n_n266, x916x, n_n271, n_n63, x1602x, x862x}, n_n787);
	defparam lut_12541.LUT_SIZE = 7;
	defparam lut_12541.mask = 128'h33ffffff33ffffff5555557755555f7f;

	lut_sub lut_12545 ({sk[2609], x907x, n_n266, x916x, x901x, x89x, n_n225}, x856x);
	defparam lut_12545.LUT_SIZE = 7;
	defparam lut_12545.mask = 128'h33ffffff33ffffff0000003700000077;

	lut_sub lut_12549 ({sk[2610], n_n268, x912x, x368x, n_n225, x55x, x856x}, x22773x);
	defparam lut_12549.LUT_SIZE = 7;
	defparam lut_12549.mask = 128'h33ffffff33ffffff5555555577ff7fff;

	lut_sub lut_12554 ({sk[2611], i_9_, i_10_, i_11_, i_15_, n_n228}, x1606x);
	defparam lut_12554.LUT_SIZE = 6;
	defparam lut_12554.mask = 64'h77ff77ff10001100;

	lut_sub lut_12558 ({sk[2612], x915x, n_n273, n_n283, n_n15, n_n59, x1606x}, x22781x);
	defparam lut_12558.LUT_SIZE = 7;
	defparam lut_12558.mask = 128'h33ffffff33ffffff00000000007f777f;

	lut_sub lut_12564 ({sk[2613], i_14_, i_13_, i_12_, x903x, x897x}, x427x);
	defparam lut_12564.LUT_SIZE = 6;
	defparam lut_12564.mask = 64'h77ff77ff00000533;

	lut_sub lut_12568 ({sk[2614], i_14_, i_13_, i_12_, i_15_, n_n270, x276x}, x1609x);
	defparam lut_12568.LUT_SIZE = 7;
	defparam lut_12568.mask = 128'h33ffffff33ffffff5577555575557555;

	lut_sub lut_12574 ({sk[2615], i_14_, i_13_, i_12_, n_n53, x908x, x902x}, x22565x);
	defparam lut_12574.LUT_SIZE = 7;
	defparam lut_12574.mask = 128'h33ffffff33ffffff0005000003050303;

	lut_sub lut_12580 ({sk[2616], n_n7441, n_n6860, n_n7405, n_n6858, x22565x}, n_n409);
	defparam lut_12580.LUT_SIZE = 6;
	defparam lut_12580.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_12586 ({sk[2617], i_14_, i_13_, i_12_, i_15_, x900x, n_n267}, x1613x);
	defparam lut_12586.LUT_SIZE = 7;
	defparam lut_12586.mask = 128'h33ffffff33ffffff0555505555335550;

	lut_sub lut_12599 ({sk[2618], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1619x);
	defparam lut_12599.LUT_SIZE = 7;
	defparam lut_12599.mask = 128'h33ffffff33ffffff1050405040004040;

	lut_sub lut_12609 ({sk[2619], i_14_, i_13_, i_12_, i_15_, n_n242, n_n259}, x1618x);
	defparam lut_12609.LUT_SIZE = 7;
	defparam lut_12609.mask = 128'h33ffffff33ffffff0333303375057570;

	lut_sub lut_12625 ({sk[2620], i_14_, i_13_, i_12_, i_15_, x899x, n_n259}, x1620x);
	defparam lut_12625.LUT_SIZE = 7;
	defparam lut_12625.mask = 128'h33ffffff33ffffff0505005555337350;

	lut_sub lut_12636 ({sk[2621], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x1622x);
	defparam lut_12636.LUT_SIZE = 7;
	defparam lut_12636.mask = 128'h33ffffff33ffffff3355505505050500;

	lut_sub lut_12646 ({sk[2622], i_14_, i_13_, i_12_, i_15_, x901x, n_n247}, x1621x);
	defparam lut_12646.LUT_SIZE = 7;
	defparam lut_12646.mask = 128'h33ffffff33ffffff3777507700000000;

	lut_sub lut_12656 ({sk[2623], i_14_, i_13_, i_12_, i_15_, n_n282, x205x}, x1623x);
	defparam lut_12656.LUT_SIZE = 7;
	defparam lut_12656.mask = 128'h33ffffff33ffffff5557555777557575;

	lut_sub lut_12664 ({sk[2624], n_n2, x82x, x1932x, x5202x, x5721x, x1867x}, x19785x);
	defparam lut_12664.LUT_SIZE = 7;
	defparam lut_12664.mask = 128'h33ffffff33ffffff3f3f3f3f7fffffff;

	lut_sub lut_12670 ({sk[2625], i_14_, i_13_, i_12_, i_15_, n_n282, n_n247}, x1624x);
	defparam lut_12670.LUT_SIZE = 7;
	defparam lut_12670.mask = 128'h33ffffff33ffffff0333003335055550;

	lut_sub lut_12682 ({sk[2626], x915x, n_n273, n_n283, x93x, n_n32, x85x}, x19776x);
	defparam lut_12682.LUT_SIZE = 7;
	defparam lut_12682.mask = 128'h33ffffff33ffffff00000000003f777f;

	lut_sub lut_12687 ({sk[2627], n_n1, n_n2, n_n76, x82x, x1899x, x1591x}, x24157x);
	defparam lut_12687.LUT_SIZE = 7;
	defparam lut_12687.mask = 128'h33ffffff33ffffffffff8800f0f08000;

	lut_sub lut_12692 ({sk[2628], n_n1, n_n2, n_n108, x90x, x60x, x1951x}, x19787x);
	defparam lut_12692.LUT_SIZE = 7;
	defparam lut_12692.mask = 128'h33ffffff33ffffff00007f7f00ff7fff;

	lut_sub lut_12697 ({sk[2629], n_n110, x915x, n_n273, n_n283, n_n2860, x1864x}, x19788x);
	defparam lut_12697.LUT_SIZE = 7;
	defparam lut_12697.mask = 128'h33ffffff33ffffff3333337733333f7f;

	lut_sub lut_12701 ({sk[2630], x915x, n_n273, x146x, x176x, n_n11, x113x}, x5185x);
	defparam lut_12701.LUT_SIZE = 7;
	defparam lut_12701.mask = 128'h33ffffff33ffffff0000000000007fff;

	lut_sub lut_12706 ({sk[2631], n_n2, x265x, n_n228, x912x, x5710x, x1879x}, x19791x);
	defparam lut_12706.LUT_SIZE = 7;
	defparam lut_12706.mask = 128'h33ffffff33ffffff33333333777fffff;

	lut_sub lut_12711 ({sk[2632], n_n1, x90x, x155x, x5204x, n_n3520, x70x}, x24142x);
	defparam lut_12711.LUT_SIZE = 7;
	defparam lut_12711.mask = 128'h33ffffff33ffffffc0c0c0c080000000;

	lut_sub lut_12714 ({sk[2633], n_n1, n_n2, n_n42, x68x, x179x, x98x}, x19798x);
	defparam lut_12714.LUT_SIZE = 7;
	defparam lut_12714.mask = 128'h33ffffff33ffffff00007f7f33ff7fff;

	lut_sub lut_12720 ({sk[2634], x915x, n_n273, n_n220, x914x, x106x, x1947x}, x19804x);
	defparam lut_12720.LUT_SIZE = 7;
	defparam lut_12720.mask = 128'h33ffffff33ffffff000000000000777f;

	lut_sub lut_12724 ({sk[2635], i_14_, i_13_, i_12_, i_15_, n_n282, n_n253}, x1846x);
	defparam lut_12724.LUT_SIZE = 7;
	defparam lut_12724.mask = 128'h33ffffff33ffffff0550505003033330;

	lut_sub lut_12734 ({sk[2636], n_n1, n_n2, x93x, x45x, x171x, x1846x}, x19805x);
	defparam lut_12734.LUT_SIZE = 7;
	defparam lut_12734.mask = 128'h33ffffff33ffffff00007f7f00ff7fff;

	lut_sub lut_12739 ({sk[2637], i_14_, i_13_, i_12_, i_15_, x101x, n_n282}, x1627x);
	defparam lut_12739.LUT_SIZE = 7;
	defparam lut_12739.mask = 128'h33ffffff33ffffff3373777337373733;

	lut_sub lut_12748 ({sk[2638], n_n6, n_n5, n_n222, x900x, n_n95, x631x}, x21791x);
	defparam lut_12748.LUT_SIZE = 7;
	defparam lut_12748.mask = 128'h33ffffff33ffffff5555555f7777777f;

	lut_sub lut_12752 ({sk[2639], n_n281, n_n6, n_n222, x898x, x129x, x21791x}, x21792x);
	defparam lut_12752.LUT_SIZE = 7;
	defparam lut_12752.mask = 128'h33ffffff33ffffff5555777f55557f7f;

	lut_sub lut_12757 ({sk[2640], i_14_, i_13_, i_12_, i_15_, n_n253, n_n267}, x1631x);
	defparam lut_12757.LUT_SIZE = 7;
	defparam lut_12757.mask = 128'h33ffffff33ffffff0707700700007300;

	lut_sub lut_12769 ({sk[2641], i_14_, i_13_, i_12_, i_15_, n_n267, n_n137}, x1630x);
	defparam lut_12769.LUT_SIZE = 7;
	defparam lut_12769.mask = 128'h33ffffff33ffffff0707350705053705;

	lut_sub lut_12777 ({sk[2642], n_n6, n_n5, x1329x, x1328x, x1631x, x1630x}, x21800x);
	defparam lut_12777.LUT_SIZE = 7;
	defparam lut_12777.mask = 128'h33ffffff33ffffff00003f3f55ff7fff;

	lut_sub lut_12782 ({sk[2643], n_n48, n_n53, n_n150, x679x, x1769x, x21786x}, n_n1773);
	defparam lut_12782.LUT_SIZE = 7;
	defparam lut_12782.mask = 128'h33ffffff33ffffff5f5f7fff5fff7fff;

	lut_sub lut_12788 ({sk[2644], n_n48, n_n6500, n_n6503, x102x, x1332x, x21784x}, x24099x);
	defparam lut_12788.LUT_SIZE = 7;
	defparam lut_12788.mask = 128'h33ffffff33ffffffaa00000080000000;

	lut_sub lut_12791 ({sk[2645], i_14_, i_13_, i_12_, x903x, x897x, x279x}, x1810x);
	defparam lut_12791.LUT_SIZE = 7;
	defparam lut_12791.mask = 128'h33ffffff33ffffff77555f5555555555;

	lut_sub lut_12795 ({sk[2646], n_n6, n_n5, n_n108, n_n80, x249x, x1810x}, x21808x);
	defparam lut_12795.LUT_SIZE = 7;
	defparam lut_12795.mask = 128'h33ffffff33ffffff00003f3f55ff7fff;

	lut_sub lut_12800 ({sk[2647], i_14_, i_13_, i_12_, i_15_, n_n242, n_n259}, x1775x);
	defparam lut_12800.LUT_SIZE = 7;
	defparam lut_12800.mask = 128'h33ffffff33ffffff0507000700007700;

	lut_sub lut_12810 ({sk[2648], i_14_, i_13_, i_12_, i_15_, n_n242, x230x}, x1774x);
	defparam lut_12810.LUT_SIZE = 7;
	defparam lut_12810.mask = 128'h33ffffff33ffffff5757755755557755;

	lut_sub lut_12818 ({sk[2649], i_7_, i_8_, i_6_, x909x, x1775x, x1774x}, x21809x);
	defparam lut_12818.LUT_SIZE = 7;
	defparam lut_12818.mask = 128'h33ffffff33ffffff0000000005000300;

	lut_sub lut_12821 ({sk[2650], n_n222, x164x, n_n207, n_n225, x897x, n_n150}, x21815x);
	defparam lut_12821.LUT_SIZE = 7;
	defparam lut_12821.mask = 128'h33ffffff33ffffff0003555700335577;

	lut_sub lut_12825 ({sk[2651], n_n6, n_n5, n_n14, n_n147, n_n8, n_n58}, x24098x);
	defparam lut_12825.LUT_SIZE = 7;
	defparam lut_12825.mask = 128'h33ffffff33ffffffffffa000c0c08000;

	lut_sub lut_12830 ({sk[2652], n_n220, x901x, x900x, x164x, x21815x, x24098x}, x21817x);
	defparam lut_12830.LUT_SIZE = 7;
	defparam lut_12830.mask = 128'h33ffffff33ffffffbbbbbbbbbbbfbfbf;

	lut_sub lut_12835 ({sk[2653], i_14_, i_13_, i_12_, i_15_, n_n282, n_n270}, x1633x);
	defparam lut_12835.LUT_SIZE = 7;
	defparam lut_12835.mask = 128'h33ffffff33ffffff0307300700007700;

	lut_sub lut_12846 ({sk[2654], i_14_, i_13_, i_12_, i_15_, x154x, n_n247}, x1632x);
	defparam lut_12846.LUT_SIZE = 7;
	defparam lut_12846.mask = 128'h33ffffff33ffffff3737733733337733;

	lut_sub lut_12854 ({sk[2655], n_n6, n_n5, x1201x, x1200x, x1633x, x1632x}, x21825x);
	defparam lut_12854.LUT_SIZE = 7;
	defparam lut_12854.mask = 128'h33ffffff33ffffff000055ff3f3f7fff;

	lut_sub lut_12859 ({sk[2656], x909x, n_n261, n_n263, n_n14, x1768x, x195x}, n_n1761);
	defparam lut_12859.LUT_SIZE = 7;
	defparam lut_12859.mask = 128'h33ffffff33ffffff0000000000335f7f;

	lut_sub lut_12863 ({sk[2657], x909x, n_n261, n_n263, n_n8, n_n58, x21814x}, x21816x);
	defparam lut_12863.LUT_SIZE = 7;
	defparam lut_12863.mask = 128'h33ffffff33ffffff55555555555f777f;

	lut_sub lut_12867 ({sk[2658], i_15_, n_n48, n_n6871, n_n138, n_n6861, x230x}, x21846x);
	defparam lut_12867.LUT_SIZE = 7;
	defparam lut_12867.mask = 128'h33ffffff33ffffff33ff77ff33ff7fff;

	lut_sub lut_12872 ({sk[2659], n_n53, n_n6868, n_n6867, n_n71, n_n72, x21846x}, x21847x);
	defparam lut_12872.LUT_SIZE = 7;
	defparam lut_12872.mask = 128'h33ffffff33ffffff55ffffff7fffffff;

	lut_sub lut_12878 ({sk[2660], n_n48, n_n1779, n_n1778, x1595x, x21839x, x21847x}, x21856x);
	defparam lut_12878.LUT_SIZE = 7;
	defparam lut_12878.mask = 128'h33ffffff33ffffff77ffffff7fffffff;

	lut_sub lut_12884 ({sk[2661], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x22677x);
	defparam lut_12884.LUT_SIZE = 7;
	defparam lut_12884.mask = 128'h33ffffff33ffffff0000000010101041;

	lut_sub lut_12890 ({sk[2662], n_n6, n_n5, n_n197, n_n216, x107x, x161x}, x22678x);
	defparam lut_12890.LUT_SIZE = 7;
	defparam lut_12890.mask = 128'h33ffffff33ffffff000077ff3f3f7fff;

	lut_sub lut_12896 ({sk[2663], x909x, n_n261, x128x, x161x, x22677x}, x2064x);
	defparam lut_12896.LUT_SIZE = 6;
	defparam lut_12896.mask = 64'h77ff77ff0000007f;

	lut_sub lut_12900 ({sk[2664], n_n5, n_n216, x114x, x109x, x128x, x2064x}, x22679x);
	defparam lut_12900.LUT_SIZE = 7;
	defparam lut_12900.mask = 128'h33ffffff33ffffff555555557fffffff;

	lut_sub lut_12906 ({sk[2665], x901x, x900x, n_n228, x164x, n_n207, x262x}, x24175x);
	defparam lut_12906.LUT_SIZE = 7;
	defparam lut_12906.mask = 128'h33ffffff33ffffffeeeeeee0eee0eee0;

	lut_sub lut_12913 ({sk[2666], n_n6, n_n228, x912x, x902x, x5130x, x24175x}, x22685x);
	defparam lut_12913.LUT_SIZE = 7;
	defparam lut_12913.mask = 128'h33ffffff33ffffffbbbbbbbbbbbbbfff;

	lut_sub lut_12918 ({sk[2667], x909x, n_n261, x899x, n_n228, x897x}, x22680x);
	defparam lut_12918.LUT_SIZE = 6;
	defparam lut_12918.mask = 64'h77ff77ff00000013;

	lut_sub lut_12921 ({sk[2668], n_n5, n_n11, n_n227, n_n15, n_n59, x275x}, x24072x);
	defparam lut_12921.LUT_SIZE = 7;
	defparam lut_12921.mask = 128'h33ffffff33ffffffffaaffaac0800000;

	lut_sub lut_12926 ({sk[2669], i_7_, i_8_, i_6_, x909x, n_n206, x190x}, x24073x);
	defparam lut_12926.LUT_SIZE = 7;
	defparam lut_12926.mask = 128'h33ffffff33fffffffffffffafcfffcff;

	lut_sub lut_12938 ({sk[2670], n_n5, n_n9, n_n226, x22680x, x24072x, x24073x}, x22686x);
	defparam lut_12938.LUT_SIZE = 7;
	defparam lut_12938.mask = 128'h33ffffff33ffffffefefefefefffffff;

	lut_sub lut_12944 ({sk[2671], i_14_, i_13_, i_12_, i_15_, n_n275, x145x}, x22688x);
	defparam lut_12944.LUT_SIZE = 7;
	defparam lut_12944.mask = 128'h33ffffff33ffffff5555555557555775;

	lut_sub lut_12949 ({sk[2672], n_n6, n_n5, n_n103, x115x, x114x, x1868x}, x22691x);
	defparam lut_12949.LUT_SIZE = 7;
	defparam lut_12949.mask = 128'h33ffffff33ffffff00000f0f77ff7fff;

	lut_sub lut_12954 ({sk[2673], n_n103, x909x, n_n263, x120x, n_n816, x22688x}, x22692x);
	defparam lut_12954.LUT_SIZE = 7;
	defparam lut_12954.mask = 128'h33ffffff33ffffff3333337f333333ff;

	lut_sub lut_12959 ({sk[2674], i_9_, i_10_, i_11_, i_15_, n_n258}, x1649x);
	defparam lut_12959.LUT_SIZE = 6;
	defparam lut_12959.mask = 64'h77ff77ff00040004;

	lut_sub lut_12962 ({sk[2675], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1652x);
	defparam lut_12962.LUT_SIZE = 7;
	defparam lut_12962.mask = 128'h33ffffff33ffffff0050000040104040;

	lut_sub lut_12969 ({sk[2676], i_14_, i_13_, i_12_, i_15_, n_n242, n_n259}, x1651x);
	defparam lut_12969.LUT_SIZE = 7;
	defparam lut_12969.mask = 128'h33ffffff33ffffff0037000070037030;

	lut_sub lut_12979 ({sk[2677], n_n5796, n_n56, x170x, n_n76, x49x, x4998x}, x19943x);
	defparam lut_12979.LUT_SIZE = 7;
	defparam lut_12979.mask = 128'h33ffffff33ffffff55557fffffffffff;

	lut_sub lut_12985 ({sk[2678], n_n266, x909x, x111x, x124x, x212x, n_n4924}, x19944x);
	defparam lut_12985.LUT_SIZE = 7;
	defparam lut_12985.mask = 128'h33ffffff33ffffff5555555555557fff;

	lut_sub lut_12990 ({sk[2679], i_7_, i_8_, i_6_, x909x, x125x, x258x}, x19932x);
	defparam lut_12990.LUT_SIZE = 7;
	defparam lut_12990.mask = 128'h33ffffff33ffffff0000000000000007;

	lut_sub lut_12993 ({sk[2680], n_n271, x909x, x90x, x60x, n_n6190}, x19933x);
	defparam lut_12993.LUT_SIZE = 6;
	defparam lut_12993.mask = 64'h77ff77ff5555557f;

	lut_sub lut_12997 ({sk[2681], x917x, n_n272, n_n5796, n_n4970, n_n4966, n_n4967}, x19953x);
	defparam lut_12997.LUT_SIZE = 7;
	defparam lut_12997.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_13003 ({sk[2682], x913x, n_n133, n_n220, x905x, n_n279, n_n107}, x19948x);
	defparam lut_13003.LUT_SIZE = 7;
	defparam lut_13003.mask = 128'h33ffffff33ffffff575fffff77ffffff;

	lut_sub lut_13010 ({sk[2683], n_n152, x299x, n_n57, x99x, x41x, x19948x}, x19954x);
	defparam lut_13010.LUT_SIZE = 7;
	defparam lut_13010.mask = 128'h33ffffff33ffffff003f003f557fffff;

	lut_sub lut_13015 ({sk[2684], n_n139, n_n110, x294x, n_n108, n_n132, x54x}, x4958x);
	defparam lut_13015.LUT_SIZE = 7;
	defparam lut_13015.mask = 128'h33ffffff33ffffff133333335fffffff;

	lut_sub lut_13024 ({sk[2685], x211x, x48x, n_n130, n_n108, n_n132, x103x}, x24180x);
	defparam lut_13024.LUT_SIZE = 7;
	defparam lut_13024.mask = 128'h33ffffff33ffffffffa0cc00ff00cc00;

	lut_sub lut_13028 ({sk[2686], n_n155, x927x, x211x, n_n128, n_n5693, x609x}, x19965x);
	defparam lut_13028.LUT_SIZE = 7;
	defparam lut_13028.mask = 128'h33ffffff33ffffff777f777f777fffff;

	lut_sub lut_13033 ({sk[2687], n_n312, x507x, n_n130, n_n111, x4972x, x19961x}, x19966x);
	defparam lut_13033.LUT_SIZE = 7;
	defparam lut_13033.mask = 128'h33ffffff33ffffff777fffffffffffff;

	lut_sub lut_13039 ({sk[2688], i_14_, i_13_, i_12_, x904x, x906x}, x1683x);
	defparam lut_13039.LUT_SIZE = 6;
	defparam lut_13039.mask = 64'h77ff77ff05553033;

	lut_sub lut_13046 ({sk[2689], i_7_, i_8_, i_6_, x909x, n_n7, x199x}, n_n3803);
	defparam lut_13046.LUT_SIZE = 7;
	defparam lut_13046.mask = 128'h33ffffff33ffffff0000000005000300;

	lut_sub lut_13049 ({sk[2690], i_14_, i_13_, i_12_, i_15_, x902x, n_n270}, x20136x);
	defparam lut_13049.LUT_SIZE = 7;
	defparam lut_13049.mask = 128'h33ffffff33ffffff0000000005053350;

	lut_sub lut_13054 ({sk[2691], n_n266, n_n271, x909x, n_n76, x82x, x1898x}, x20227x);
	defparam lut_13054.LUT_SIZE = 7;
	defparam lut_13054.mask = 128'h33ffffff33ffffff0000005f0033007f;

	lut_sub lut_13058 ({sk[2692], n_n57, x258x, x720x, x636x, x555x, x70x}, x24178x);
	defparam lut_13058.LUT_SIZE = 7;
	defparam lut_13058.mask = 128'h33ffffff33ffffffc000c00080000000;

	lut_sub lut_13061 ({sk[2693], n_n1, n_n2, n_n108, x60x, n_n42, x68x}, x20868x);
	defparam lut_13061.LUT_SIZE = 7;
	defparam lut_13061.mask = 128'h33ffffff33ffffff00005f5f33ff7fff;

	lut_sub lut_13066 ({sk[2694], x915x, n_n273, x82x, x111x, x1923x}, x20870x);
	defparam lut_13066.LUT_SIZE = 6;
	defparam lut_13066.mask = 64'h77ff77ff0000007f;

	lut_sub lut_13070 ({sk[2695], n_n2, x1873x, x45x, x171x, x20868x, x20870x}, x20872x);
	defparam lut_13070.LUT_SIZE = 7;
	defparam lut_13070.mask = 128'h33ffffff33ffffff777777777fffffff;

	lut_sub lut_13076 ({sk[2696], x915x, n_n273, n_n283, n_n12, x125x, x1879x}, x20865x);
	defparam lut_13076.LUT_SIZE = 7;
	defparam lut_13076.mask = 128'h33ffffff33ffffff0000000000770f7f;

	lut_sub lut_13080 ({sk[2697], n_n1, n_n226, x159x, x5204x, n_n3520, x70x}, x20866x);
	defparam lut_13080.LUT_SIZE = 7;
	defparam lut_13080.mask = 128'h33ffffff33ffffff3f3f3f3f7fffffff;

	lut_sub lut_13086 ({sk[2698], x20862x, x20863x, n_n3424, x20865x, x20866x}, x20873x);
	defparam lut_13086.LUT_SIZE = 6;
	defparam lut_13086.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_13092 ({sk[2699], i_14_, i_13_, i_12_, i_15_, n_n259, x187x}, x1714x);
	defparam lut_13092.LUT_SIZE = 7;
	defparam lut_13092.mask = 128'h33ffffff33ffffff5555555575577575;

	lut_sub lut_13098 ({sk[2700], n_n6, x183x, n_n5, x218x, n_n227, x1714x}, x20880x);
	defparam lut_13098.LUT_SIZE = 7;
	defparam lut_13098.mask = 128'h33ffffff33ffffff111f111f111fffff;

	lut_sub lut_13102 ({sk[2701], x915x, x400x, x911x, n_n263, x333x, n_n225}, x20887x);
	defparam lut_13102.LUT_SIZE = 7;
	defparam lut_13102.mask = 128'h33ffffff33ffffff3333333333373f3f;

	lut_sub lut_13106 ({sk[2702], n_n208, x916x, x905x, x166x, n_n225, x20887x}, x20889x);
	defparam lut_13106.LUT_SIZE = 7;
	defparam lut_13106.mask = 128'h33ffffff33ffffff5555555555555f7f;

	lut_sub lut_13110 ({sk[2703], i_14_, i_13_, i_12_, i_15_, n_n267, x19469x}, x1799x);
	defparam lut_13110.LUT_SIZE = 7;
	defparam lut_13110.mask = 128'h33ffffff33ffffff7555575555755555;

	lut_sub lut_13115 ({sk[2704], i_14_, i_13_, i_12_, i_15_, n_n267, x246x}, x1798x);
	defparam lut_13115.LUT_SIZE = 7;
	defparam lut_13115.mask = 128'h33ffffff33ffffff7555575555555555;

	lut_sub lut_13119 ({sk[2705], i_14_, i_13_, i_12_, i_11_, i_15_, n_n269}, x1659x);
	defparam lut_13119.LUT_SIZE = 7;
	defparam lut_13119.mask = 128'h33ffffff33ffffff0000010000440011;

	lut_sub lut_13125 ({sk[2706], x909x, x173x, n_n263, x100x, x281x, n_n3448}, x20894x);
	defparam lut_13125.LUT_SIZE = 7;
	defparam lut_13125.mask = 128'h33ffffff33ffffff55555555557f55ff;

	lut_sub lut_13130 ({sk[2707], n_n4809, x909x, n_n261, x539x, x1659x, x20894x}, x20895x);
	defparam lut_13130.LUT_SIZE = 7;
	defparam lut_13130.mask = 128'h33ffffff33ffffff5f5f5f7fffffffff;

	lut_sub lut_13135 ({sk[2708], n_n208, x916x, x485x, n_n223, x123x, x100x}, n_n3442);
	defparam lut_13135.LUT_SIZE = 7;
	defparam lut_13135.mask = 128'h33ffffff33ffffff00ff00ff00ff7fff;

	lut_sub lut_13140 ({sk[2709], n_n151, x909x, n_n261, n_n263, x118x, n_n3550}, x20878x);
	defparam lut_13140.LUT_SIZE = 7;
	defparam lut_13140.mask = 128'h33ffffff33ffffff55555757555557ff;

	lut_sub lut_13144 ({sk[2710], n_n208, x909x, n_n263, x72x, x480x, x1713x}, x20879x);
	defparam lut_13144.LUT_SIZE = 7;
	defparam lut_13144.mask = 128'h33ffffff33ffffff3333333f3333777f;

	lut_sub lut_13148 ({sk[2711], n_n4, n_n93, n_n6823, x381x, x455x, x388x}, x20888x);
	defparam lut_13148.LUT_SIZE = 7;
	defparam lut_13148.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_13154 ({sk[2712], x20880x, x20889x, n_n3442, x20878x, x20879x, x20888x}, x20896x);
	defparam lut_13154.LUT_SIZE = 7;
	defparam lut_13154.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_13161 ({sk[2713], i_14_, i_13_, i_12_, x913x, x898x}, x20504x);
	defparam lut_13161.LUT_SIZE = 6;
	defparam lut_13161.mask = 64'h77ff77ff03300005;

	lut_sub lut_13165 ({sk[2714], i_14_, i_13_, i_12_, i_15_, n_n242, x20504x}, x1660x);
	defparam lut_13165.LUT_SIZE = 7;
	defparam lut_13165.mask = 128'h33ffffff33ffffff5757557775557555;

	lut_sub lut_13173 ({sk[2715], i_14_, i_13_, i_12_, i_15_, x905x, n_n259}, x1662x);
	defparam lut_13173.LUT_SIZE = 7;
	defparam lut_13173.mask = 128'h33ffffff33ffffff0537333755055550;

	lut_sub lut_13186 ({sk[2716], i_14_, i_13_, i_12_, i_15_, n_n242, n_n270}, x1661x);
	defparam lut_13186.LUT_SIZE = 7;
	defparam lut_13186.mask = 128'h33ffffff33ffffff0555505530003030;

	lut_sub lut_13196 ({sk[2717], x911x, n_n258, n_n94, x381x, x140x, x1661x}, x20068x);
	defparam lut_13196.LUT_SIZE = 7;
	defparam lut_13196.mask = 128'h33ffffff33ffffff0f7f0f7f0f7f0fff;

	lut_sub lut_13201 ({sk[2718], i_14_, i_13_, i_12_, x915x, n_n263, x903x}, n_n707);
	defparam lut_13201.LUT_SIZE = 7;
	defparam lut_13201.mask = 128'h33ffffff33ffffff0000000001000101;

	lut_sub lut_13205 ({sk[2719], i_14_, i_13_, i_12_, i_15_, n_n275, x903x}, x1665x);
	defparam lut_13205.LUT_SIZE = 7;
	defparam lut_13205.mask = 128'h33ffffff33ffffff0055555503030300;

	lut_sub lut_13212 ({sk[2720], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1664x);
	defparam lut_13212.LUT_SIZE = 7;
	defparam lut_13212.mask = 128'h33ffffff33ffffff0105040505010504;

	lut_sub lut_13225 ({sk[2721], i_14_, i_13_, i_12_, x902x, x1665x}, x1663x);
	defparam lut_13225.LUT_SIZE = 6;
	defparam lut_13225.mask = 64'h77ff77ff55557775;

	lut_sub lut_13230 ({sk[2722], i_14_, i_13_, i_12_, x915x, n_n263, x897x}, x20070x);
	defparam lut_13230.LUT_SIZE = 7;
	defparam lut_13230.mask = 128'h33ffffff33ffffff0101000100000000;

	lut_sub lut_13234 ({sk[2723], n_n100, n_n94, n_n707, x1664x, x1663x, x20070x}, x20073x);
	defparam lut_13234.LUT_SIZE = 7;
	defparam lut_13234.mask = 128'h33ffffff33ffffff55ff77ff5fff7fff;

	lut_sub lut_13239 ({sk[2724], n_n4, n_n64, n_n3, n_n7406, n_n147, n_n58}, x21891x);
	defparam lut_13239.LUT_SIZE = 7;
	defparam lut_13239.mask = 128'h33ffffff33ffffff0f7f0fff3f7f3fff;

	lut_sub lut_13245 ({sk[2725], n_n4, n_n7402, n_n3, n_n62, n_n8, x21891x}, n_n1724);
	defparam lut_13245.LUT_SIZE = 7;
	defparam lut_13245.mask = 128'h33ffffff33ffffff555fffff7f7fffff;

	lut_sub lut_13251 ({sk[2726], i_14_, i_13_, i_12_, n_n273, x922x, x902x}, x544x);
	defparam lut_13251.LUT_SIZE = 7;
	defparam lut_13251.mask = 128'h33ffffff33ffffff0000000001010100;

	lut_sub lut_13255 ({sk[2727], n_n7400, n_n7440, n_n7344, x349x, n_n876, x544x}, x22793x);
	defparam lut_13255.LUT_SIZE = 7;
	defparam lut_13255.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_13262 ({sk[2728], x911x, n_n279, n_n94, x697x, x382x, x892x}, x22804x);
	defparam lut_13262.LUT_SIZE = 7;
	defparam lut_13262.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_13267 ({sk[2729], x907x, n_n228, n_n100, n_n6824, x548x, x22804x}, n_n808);
	defparam lut_13267.LUT_SIZE = 7;
	defparam lut_13267.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_13272 ({sk[2730], n_n4, n_n31, n_n11, n_n94, n_n884, x601x}, x24200x);
	defparam lut_13272.LUT_SIZE = 7;
	defparam lut_13272.mask = 128'h33ffffff33ffffff8880888088800000;

	lut_sub lut_13277 ({sk[2731], x914x, x911x, n_n228, n_n94, n_n6834, x24200x}, x22809x);
	defparam lut_13277.LUT_SIZE = 7;
	defparam lut_13277.mask = 128'h33ffffff33ffffffbbbbbbbfbbbfbbbf;

	lut_sub lut_13282 ({sk[2732], n_n4, n_n9, n_n3, n_n7224, x134x, x607x}, x22792x);
	defparam lut_13282.LUT_SIZE = 7;
	defparam lut_13282.mask = 128'h33ffffff33ffffff5f7f5f7f5f7fffff;

	lut_sub lut_13287 ({sk[2733], n_n809, n_n785, x22793x, n_n808, x22809x, x22792x}, x22815x);
	defparam lut_13287.LUT_SIZE = 7;
	defparam lut_13287.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_13294 ({sk[2734], i_7_, i_8_, i_6_, x922x, x41x}, x2328x);
	defparam lut_13294.LUT_SIZE = 6;
	defparam lut_13294.mask = 64'h77ff77ff00100000;

	lut_sub lut_13296 ({sk[2735], i_14_, i_13_, i_12_, x905x, x899x}, x441x);
	defparam lut_13296.LUT_SIZE = 6;
	defparam lut_13296.mask = 64'h77ff77ff07003000;

	lut_sub lut_13300 ({sk[2736], i_14_, i_13_, i_12_, i_15_, n_n259, x441x}, x1681x);
	defparam lut_13300.LUT_SIZE = 7;
	defparam lut_13300.mask = 128'h33ffffff33ffffff5555555555577575;

	lut_sub lut_13305 ({sk[2737], x907x, x909x, n_n258, n_n261, n_n263, x903x}, x2194x);
	defparam lut_13305.LUT_SIZE = 7;
	defparam lut_13305.mask = 128'h33ffffff33ffffff000000150000003f;

	lut_sub lut_13310 ({sk[2738], n_n6, n_n257, n_n61, n_n227, x1681x, x2194x}, x22572x);
	defparam lut_13310.LUT_SIZE = 7;
	defparam lut_13310.mask = 128'h33ffffff33ffffff5757575757ffffff;

	lut_sub lut_13315 ({sk[2739], n_n5, n_n240, n_n61, n_n246, n_n207, x292x}, x22571x);
	defparam lut_13315.LUT_SIZE = 7;
	defparam lut_13315.mask = 128'h33ffffff33ffffff111111111fffffff;

	lut_sub lut_13320 ({sk[2740], n_n416, x22572x, x22571x}, n_n360);
	defparam lut_13320.LUT_SIZE = 4;
	defparam lut_13320.mask = 16'h777f;

	lut_sub lut_13324 ({sk[2741], i_14_, i_13_, i_12_, i_15_, x902x, n_n275}, x19395x);
	defparam lut_13324.LUT_SIZE = 7;
	defparam lut_13324.mask = 128'h33ffffff33ffffff5000050000500037;

	lut_sub lut_13330 ({sk[2742], x915x, n_n273, x68x, x45x, n_n6879, x171x}, n_n3435);
	defparam lut_13330.LUT_SIZE = 7;
	defparam lut_13330.mask = 128'h33ffffff33ffffff3333333333337fff;

	lut_sub lut_13335 ({sk[2743], n_n226, n_n53, n_n6867, n_n2272, x123x, n_n952}, x20905x);
	defparam lut_13335.LUT_SIZE = 7;
	defparam lut_13335.mask = 128'h33ffffff33ffffff5fff7fff5fffffff;

	lut_sub lut_13341 ({sk[2744], i_9_, i_10_, i_11_, i_15_, x108x, n_n225}, x1699x);
	defparam lut_13341.LUT_SIZE = 7;
	defparam lut_13341.mask = 128'h33ffffff33ffffff3333337733333333;

	lut_sub lut_13345 ({sk[2745], i_14_, i_13_, i_12_, i_15_, n_n253, x1699x}, x1698x);
	defparam lut_13345.LUT_SIZE = 7;
	defparam lut_13345.mask = 128'h33ffffff33ffffff5555557757555775;

	lut_sub lut_13352 ({sk[2746], x911x, n_n258, n_n48, n_n53, x899x, n_n4073}, x22699x);
	defparam lut_13352.LUT_SIZE = 7;
	defparam lut_13352.mask = 128'h33ffffff33ffffff5555575755555fff;

	lut_sub lut_13357 ({sk[2747], n_n283, x126x, x922x, x483x, x145x}, x22707x);
	defparam lut_13357.LUT_SIZE = 6;
	defparam lut_13357.mask = 64'h77ff77ff3333373f;

	lut_sub lut_13361 ({sk[2748], n_n830, x22700x, n_n831, x22708x, x22699x, x22707x}, x22717x);
	defparam lut_13361.LUT_SIZE = 7;
	defparam lut_13361.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_13368 ({sk[2749], i_14_, i_13_, i_12_, i_15_, n_n282, n_n253}, x1719x);
	defparam lut_13368.LUT_SIZE = 7;
	defparam lut_13368.mask = 128'h33ffffff33ffffff0000005507030770;

	lut_sub lut_13378 ({sk[2750], n_n6, n_n41, x115x, x748x, x139x, x145x}, x22742x);
	defparam lut_13378.LUT_SIZE = 7;
	defparam lut_13378.mask = 128'h33ffffff33ffffff0f0f0f0f7fffffff;

	lut_sub lut_13384 ({sk[2751], x909x, n_n263, n_n819, x1719x, x22742x}, x22744x);
	defparam lut_13384.LUT_SIZE = 6;
	defparam lut_13384.mask = 64'h77ff77ff5f5f5f7f;

	lut_sub lut_13388 ({sk[2752], n_n283, x922x, n_n11, n_n6524, x495x, x670x}, x22722x);
	defparam lut_13388.LUT_SIZE = 7;
	defparam lut_13388.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_13393 ({sk[2753], n_n273, n_n283, x922x, n_n6878, n_n15, x1065x}, x22733x);
	defparam lut_13393.LUT_SIZE = 7;
	defparam lut_13393.mask = 128'h33ffffff33ffffff0f0f0f3f0f5f0f7f;

	lut_sub lut_13397 ({sk[2754], n_n824, x22723x, n_n825, x22734x, x22722x, x22733x}, x22745x);
	defparam lut_13397.LUT_SIZE = 7;
	defparam lut_13397.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_13404 ({sk[2755], n_n1, n_n53, x254x, x356x, x305x, x275x}, x22812x);
	defparam lut_13404.LUT_SIZE = 7;
	defparam lut_13404.mask = 128'h33ffffff33ffffff000077770fff7fff;

	lut_sub lut_13409 ({sk[2756], n_n2, x224x, n_n6878, n_n6875, x1119x, n_n952}, x22813x);
	defparam lut_13409.LUT_SIZE = 7;
	defparam lut_13409.mask = 128'h33ffffff33ffffff5fff5fff7fffffff;

	lut_sub lut_13415 ({sk[2757], n_n790, n_n789, n_n792, n_n787, x22773x, x22781x}, x22821x);
	defparam lut_13415.LUT_SIZE = 7;
	defparam lut_13415.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_13422 ({sk[2758], n_n784, n_n785, n_n751, n_n753, x22763x, x22818x}, x24071x);
	defparam lut_13422.LUT_SIZE = 7;
	defparam lut_13422.mask = 128'h33ffffff33ffffff8000000000000000;

	lut_sub lut_13424 ({sk[2759], n_n5, n_n103, n_n31, x208x, n_n227, n_n207}, x24162x);
	defparam lut_13424.LUT_SIZE = 7;
	defparam lut_13424.mask = 128'h33ffffff33ffffffffccaa88f0c0a080;

	lut_sub lut_13433 ({sk[2760], n_n208, x909x, x120x, x91x, x24162x}, n_n3686);
	defparam lut_13433.LUT_SIZE = 6;
	defparam lut_13433.mask = 64'h77ff77ffaaaaaabf;

	lut_sub lut_13437 ({sk[2761], i_14_, i_13_, i_12_, x913x, x911x, x142x}, x1713x);
	defparam lut_13437.LUT_SIZE = 7;
	defparam lut_13437.mask = 128'h33ffffff33ffffff557f555555775555;

	lut_sub lut_13442 ({sk[2762], x911x, n_n57, n_n56, x899x, n_n228, x897x}, x24207x);
	defparam lut_13442.LUT_SIZE = 7;
	defparam lut_13442.mask = 128'h33ffffff33ffffffffeeececffcccccc;

	lut_sub lut_13447 ({sk[2763], i_14_, i_13_, i_12_, x900x, x906x, x108x}, x1720x);
	defparam lut_13447.LUT_SIZE = 7;
	defparam lut_13447.mask = 128'h33ffffff33ffffff5555557f555f5555;

	lut_sub lut_13452 ({sk[2764], i_14_, i_13_, i_12_, n_n3, x904x}, x5683x);
	defparam lut_13452.LUT_SIZE = 6;
	defparam lut_13452.mask = 64'h77ff77ff00011011;

	lut_sub lut_13457 ({sk[2765], i_14_, i_13_, i_12_, n_n3, x898x}, x5682x);
	defparam lut_13457.LUT_SIZE = 6;
	defparam lut_13457.mask = 64'h77ff77ff00001110;

	lut_sub lut_13461 ({sk[2766], n_n4, n_n13, n_n12, n_n65, x409x, x349x}, x866x);
	defparam lut_13461.LUT_SIZE = 7;
	defparam lut_13461.mask = 128'h33ffffff33ffffff777777777fffffff;

	lut_sub lut_13467 ({sk[2767], i_14_, i_13_, i_12_, x900x, x906x}, x1787x);
	defparam lut_13467.LUT_SIZE = 6;
	defparam lut_13467.mask = 64'h77ff77ff37570000;

	lut_sub lut_13474 ({sk[2768], i_14_, i_13_, i_12_, x903x, x897x}, x19851x);
	defparam lut_13474.LUT_SIZE = 6;
	defparam lut_13474.mask = 64'h77ff77ff03335550;

	lut_sub lut_13481 ({sk[2769], i_9_, i_10_, i_14_, i_11_, i_15_, n_n278}, x1731x);
	defparam lut_13481.LUT_SIZE = 7;
	defparam lut_13481.mask = 128'h33ffffff33ffffff0100100040500000;

	lut_sub lut_13487 ({sk[2770], x905x, n_n258, n_n48, n_n53, x908x, x903x}, x22406x);
	defparam lut_13487.LUT_SIZE = 7;
	defparam lut_13487.mask = 128'h33ffffff33ffffff0000057700000fff;

	lut_sub lut_13493 ({sk[2771], i_9_, i_10_, i_11_, i_15_, n_n258, x187x}, x1738x);
	defparam lut_13493.LUT_SIZE = 7;
	defparam lut_13493.mask = 128'h33ffffff33ffffff7555555555555575;

	lut_sub lut_13497 ({sk[2772], n_n9, n_n57, n_n56, x209x, x309x, x132x}, x19520x);
	defparam lut_13497.LUT_SIZE = 7;
	defparam lut_13497.mask = 128'h33ffffff33ffffff333f7f7f33ffffff;

	lut_sub lut_13504 ({sk[2773], n_n273, x922x, x68x, x571x, x737x, x393x}, x19519x);
	defparam lut_13504.LUT_SIZE = 7;
	defparam lut_13504.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_13509 ({sk[2774], i_14_, i_13_, i_12_, i_15_, x908x, n_n270}, x1747x);
	defparam lut_13509.LUT_SIZE = 7;
	defparam lut_13509.mask = 128'h33ffffff33ffffff0537333755055550;

	lut_sub lut_13522 ({sk[2775], i_14_, i_13_, i_12_, i_15_, n_n242, n_n259}, x1751x);
	defparam lut_13522.LUT_SIZE = 7;
	defparam lut_13522.mask = 128'h33ffffff33ffffff0000007707070770;

	lut_sub lut_13535 ({sk[2776], i_14_, i_13_, i_12_, x900x, x906x}, x22377x);
	defparam lut_13535.LUT_SIZE = 6;
	defparam lut_13535.mask = 64'h77ff77ff07000055;

	lut_sub lut_13540 ({sk[2777], n_n6834, x825x, n_n6829, x892x, x548x, x434x}, n_n2671);
	defparam lut_13540.LUT_SIZE = 7;
	defparam lut_13540.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_13547 ({sk[2778], x915x, n_n261, n_n263, x1936x, x1816x, x1815x}, n_n2667);
	defparam lut_13547.LUT_SIZE = 7;
	defparam lut_13547.mask = 128'h33ffffff33ffffff0000000000335f7f;

	lut_sub lut_13551 ({sk[2779], i_14_, i_13_, i_12_, x915x, n_n261, x901x}, x20081x);
	defparam lut_13551.LUT_SIZE = 7;
	defparam lut_13551.mask = 128'h33ffffff33ffffff0000000001010100;

	lut_sub lut_13555 ({sk[2780], n_n100, n_n94, x1622x, x1621x, x1818x, x1817x}, x24138x);
	defparam lut_13555.LUT_SIZE = 7;
	defparam lut_13555.mask = 128'h33ffffff33ffffffffffaa00c0c08000;

	lut_sub lut_13560 ({sk[2781], n_n145, n_n73, x314x, n_n94, x380x, x471x}, n_n2673);
	defparam lut_13560.LUT_SIZE = 7;
	defparam lut_13560.mask = 128'h33ffffff33ffffff777f7f7f7f7f7f7f;

	lut_sub lut_13566 ({sk[2782], n_n22, n_n94, n_n6823, x381x, n_n6824, x388x}, x20104x);
	defparam lut_13566.LUT_SIZE = 7;
	defparam lut_13566.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_13572 ({sk[2783], i_14_, i_13_, i_12_, i_15_, x173x, n_n267}, x1763x);
	defparam lut_13572.LUT_SIZE = 7;
	defparam lut_13572.mask = 128'h33ffffff33ffffff7333373333333333;

	lut_sub lut_13576 ({sk[2784], i_14_, i_13_, i_12_, i_15_, x900x, n_n267}, x1762x);
	defparam lut_13576.LUT_SIZE = 7;
	defparam lut_13576.mask = 128'h33ffffff33ffffff5000050000500033;

	lut_sub lut_13581 ({sk[2785], i_14_, i_13_, i_12_, i_15_, n_n267, x246x}, x1764x);
	defparam lut_13581.LUT_SIZE = 7;
	defparam lut_13581.mask = 128'h33ffffff33ffffff7555575555555555;

	lut_sub lut_13585 ({sk[2786], i_14_, i_13_, i_12_, i_15_, n_n275, n_n259}, x1766x);
	defparam lut_13585.LUT_SIZE = 7;
	defparam lut_13585.mask = 128'h33ffffff33ffffff0737307555005550;

	lut_sub lut_13600 ({sk[2787], i_14_, i_13_, i_12_, i_15_, n_n270}, x1765x);
	defparam lut_13600.LUT_SIZE = 6;
	defparam lut_13600.mask = 64'h77ff77ff11055154;

	lut_sub lut_13611 ({sk[2788], n_n197, n_n57, n_n56, x3567x, x1766x, x1765x}, n_n2434);
	defparam lut_13611.LUT_SIZE = 7;
	defparam lut_13611.mask = 128'h33ffffff33ffffff0f5f3f7f0f5fffff;

	lut_sub lut_13616 ({sk[2789], n_n111, n_n48, n_n53, n_n6505, n_n34, x629x}, x21784x);
	defparam lut_13616.LUT_SIZE = 7;
	defparam lut_13616.mask = 128'h33ffffff33ffffff5f7f5f7f5f7fffff;

	lut_sub lut_13621 ({sk[2790], i_14_, i_13_, i_12_, x905x, x899x}, x375x);
	defparam lut_13621.LUT_SIZE = 6;
	defparam lut_13621.mask = 64'h77ff77ff50300000;

	lut_sub lut_13624 ({sk[2791], i_14_, i_13_, i_12_, i_15_, n_n259, x375x}, x1768x);
	defparam lut_13624.LUT_SIZE = 7;
	defparam lut_13624.mask = 128'h33ffffff33ffffff5557555755557755;

	lut_sub lut_13630 ({sk[2792], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1769x);
	defparam lut_13630.LUT_SIZE = 7;
	defparam lut_13630.mask = 128'h33ffffff33ffffff0000011000004000;

	lut_sub lut_13634 ({sk[2793], n_n273, n_n283, n_n222, x922x, x901x, n_n144}, x21786x);
	defparam lut_13634.LUT_SIZE = 7;
	defparam lut_13634.mask = 128'h33ffffff33ffffff0000050500030507;

	lut_sub lut_13637 ({sk[2794], n_n4, n_n9, n_n3, n_n226, n_n11, n_n59}, x22832x);
	defparam lut_13637.LUT_SIZE = 7;
	defparam lut_13637.mask = 128'h33ffffff33ffffff007f00ff557f55ff;

	lut_sub lut_13643 ({sk[2795], n_n4, n_n9, n_n3, n_n7440, n_n206, x22832x}, n_n775);
	defparam lut_13643.LUT_SIZE = 7;
	defparam lut_13643.mask = 128'h33ffffff33ffffff5f7f5f7f7f7fffff;

	lut_sub lut_13649 ({sk[2796], i_14_, i_13_, i_12_, i_15_, x201x, n_n242}, x1778x);
	defparam lut_13649.LUT_SIZE = 7;
	defparam lut_13649.mask = 128'h33ffffff33ffffff3333333337373773;

	lut_sub lut_13655 ({sk[2797], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1781x);
	defparam lut_13655.LUT_SIZE = 7;
	defparam lut_13655.mask = 128'h33ffffff33ffffff1010005040004000;

	lut_sub lut_13662 ({sk[2798], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1780x);
	defparam lut_13662.LUT_SIZE = 7;
	defparam lut_13662.mask = 128'h33ffffff33ffffff1010005050105040;

	lut_sub lut_13673 ({sk[2799], i_14_, i_13_, i_12_, i_15_, x902x, n_n275}, x1782x);
	defparam lut_13673.LUT_SIZE = 7;
	defparam lut_13673.mask = 128'h33ffffff33ffffff0555505555335550;

	lut_sub lut_13686 ({sk[2800], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1789x);
	defparam lut_13686.LUT_SIZE = 7;
	defparam lut_13686.mask = 128'h33ffffff33ffffff1010005050105040;

	lut_sub lut_13697 ({sk[2801], i_14_, i_13_, i_12_, i_15_, n_n259, n_n267}, x1795x);
	defparam lut_13697.LUT_SIZE = 7;
	defparam lut_13697.mask = 128'h33ffffff33ffffff0007000070007000;

	lut_sub lut_13704 ({sk[2802], n_n208, x916x, n_n61, x518x, x1795x, x24078x}, x22579x);
	defparam lut_13704.LUT_SIZE = 7;
	defparam lut_13704.mask = 128'h33ffffff33ffffffafafafafafafbfff;

	lut_sub lut_13709 ({sk[2803], i_14_, i_13_, i_12_, x900x, x904x}, x19469x);
	defparam lut_13709.LUT_SIZE = 6;
	defparam lut_13709.mask = 64'h77ff77ff50000003;

	lut_sub lut_13712 ({sk[2804], i_14_, i_13_, i_12_, i_15_, x908x, n_n270}, x1801x);
	defparam lut_13712.LUT_SIZE = 7;
	defparam lut_13712.mask = 128'h33ffffff33ffffff0537335550005000;

	lut_sub lut_13721 ({sk[2805], x915x, n_n261, n_n263, x21869x, x21870x, x1850x}, n_n1721);
	defparam lut_13721.LUT_SIZE = 7;
	defparam lut_13721.mask = 128'h33ffffff33ffffff00000000003f557f;

	lut_sub lut_13725 ({sk[2806], i_7_, i_8_, i_6_, x917x, x927x, x48x}, x21862x);
	defparam lut_13725.LUT_SIZE = 7;
	defparam lut_13725.mask = 128'h33ffffff33ffffff373333333f333f33;

	lut_sub lut_13732 ({sk[2807], i_7_, i_6_, x918x, x24148x}, x21863x);
	defparam lut_13732.LUT_SIZE = 5;
	defparam lut_13732.mask = 32'h3f3fbbbb;

	lut_sub lut_13738 ({sk[2808], i_15_, n_n94, n_n6834, n_n137, n_n6835, x1834x}, x21874x);
	defparam lut_13738.LUT_SIZE = 7;
	defparam lut_13738.mask = 128'h33ffffff33ffffff33ff7fff33ff7fff;

	lut_sub lut_13744 ({sk[2809], n_n100, n_n6814, x360x, x3143x, x21857x, x1835x}, x21875x);
	defparam lut_13744.LUT_SIZE = 7;
	defparam lut_13744.mask = 128'h33ffffff33ffffff3f3fffff7fffffff;

	lut_sub lut_13750 ({sk[2810], x21864x, n_n1721, x21862x, x21863x, x21874x, x21875x}, n_n1692);
	defparam lut_13750.LUT_SIZE = 7;
	defparam lut_13750.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_13757 ({sk[2811], n_n57, n_n56, x208x, n_n59, x50x, x156x}, n_n2442);
	defparam lut_13757.LUT_SIZE = 7;
	defparam lut_13757.mask = 128'h33ffffff33ffffff00005f5f3fff7fff;

	lut_sub lut_13763 ({sk[2812], i_14_, i_13_, i_12_, i_15_, n_n282, n_n247}, x1808x);
	defparam lut_13763.LUT_SIZE = 7;
	defparam lut_13763.mask = 128'h33ffffff33ffffff7000070000700007;

	lut_sub lut_13772 ({sk[2813], i_14_, i_13_, i_12_, i_15_, n_n282, x199x}, x1807x);
	defparam lut_13772.LUT_SIZE = 7;
	defparam lut_13772.mask = 128'h33ffffff33ffffff7555575555755557;

	lut_sub lut_13778 ({sk[2814], i_14_, i_13_, i_12_, i_15_, n_n242, x897x}, x1813x);
	defparam lut_13778.LUT_SIZE = 7;
	defparam lut_13778.mask = 128'h33ffffff33ffffff0033000075577530;

	lut_sub lut_13788 ({sk[2815], i_14_, i_13_, i_12_, i_15_, x904x, n_n253}, x1816x);
	defparam lut_13788.LUT_SIZE = 7;
	defparam lut_13788.mask = 128'h33ffffff33ffffff0555505537053733;

	lut_sub lut_13801 ({sk[2816], i_14_, i_13_, i_12_, i_15_, n_n247, x906x}, x1815x);
	defparam lut_13801.LUT_SIZE = 7;
	defparam lut_13801.mask = 128'h33ffffff33ffffff0055555533033330;

	lut_sub lut_13811 ({sk[2817], i_14_, i_13_, i_12_, i_15_, x900x, n_n253}, x1818x);
	defparam lut_13811.LUT_SIZE = 7;
	defparam lut_13811.mask = 128'h33ffffff33ffffff0555505577377750;

	lut_sub lut_13827 ({sk[2818], i_14_, i_13_, i_12_, i_15_, x900x, n_n267}, x1817x);
	defparam lut_13827.LUT_SIZE = 7;
	defparam lut_13827.mask = 128'h33ffffff33ffffff0555505573337350;

	lut_sub lut_13840 ({sk[2819], i_14_, i_13_, i_12_, x905x, x899x, x902x}, x21894x);
	defparam lut_13840.LUT_SIZE = 7;
	defparam lut_13840.mask = 128'h33ffffff33ffffff33005f0000000000;

	lut_sub lut_13844 ({sk[2820], i_14_, i_13_, i_12_, i_15_, n_n259, x21894x}, x1824x);
	defparam lut_13844.LUT_SIZE = 7;
	defparam lut_13844.mask = 128'h33ffffff33ffffff5557575755557755;

	lut_sub lut_13851 ({sk[2821], i_9_, i_10_, i_11_, i_15_, n_n281, n_n220}, x1823x);
	defparam lut_13851.LUT_SIZE = 7;
	defparam lut_13851.mask = 128'h33ffffff33ffffff0005530000000005;

	lut_sub lut_13856 ({sk[2822], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x20173x);
	defparam lut_13856.LUT_SIZE = 7;
	defparam lut_13856.mask = 128'h33ffffff33ffffff4000110000440001;

	lut_sub lut_13863 ({sk[2823], n_n281, x206x, x914x, x156x, x113x}, x24136x);
	defparam lut_13863.LUT_SIZE = 6;
	defparam lut_13863.mask = 64'h77ff77ff88008000;

	lut_sub lut_13866 ({sk[2824], i_14_, i_13_, i_12_, i_15_, n_n247, n_n267}, x1827x);
	defparam lut_13866.LUT_SIZE = 7;
	defparam lut_13866.mask = 128'h33ffffff33ffffff7000070000700007;

	lut_sub lut_13875 ({sk[2825], i_14_, i_13_, i_12_, x913x, x914x, x912x}, x1844x);
	defparam lut_13875.LUT_SIZE = 7;
	defparam lut_13875.mask = 128'h33ffffff33ffffff55003f003f000000;

	lut_sub lut_13881 ({sk[2826], i_14_, i_13_, i_12_, i_15_, x901x, n_n282}, x21343x);
	defparam lut_13881.LUT_SIZE = 7;
	defparam lut_13881.mask = 128'h33ffffff33ffffff3305005550005000;

	lut_sub lut_13888 ({sk[2827], i_14_, i_13_, i_12_, i_15_, n_n282, n_n270}, x21344x);
	defparam lut_13888.LUT_SIZE = 7;
	defparam lut_13888.mask = 128'h33ffffff33ffffff0030300007050770;

	lut_sub lut_13898 ({sk[2828], i_14_, i_13_, i_12_, i_15_, x914x, n_n247}, x1830x);
	defparam lut_13898.LUT_SIZE = 7;
	defparam lut_13898.mask = 128'h33ffffff33ffffff0537335555055550;

	lut_sub lut_13911 ({sk[2829], n_n266, n_n271, x909x, x21343x, x21344x, x1830x}, n_n2436);
	defparam lut_13911.LUT_SIZE = 7;
	defparam lut_13911.mask = 128'h33ffffff33ffffff00000055003f007f;

	lut_sub lut_13915 ({sk[2830], i_14_, i_13_, i_12_, i_15_, n_n275, n_n270}, x1833x);
	defparam lut_13915.LUT_SIZE = 7;
	defparam lut_13915.mask = 128'h33ffffff33ffffff0505005773037330;

	lut_sub lut_13929 ({sk[2831], i_14_, i_13_, i_12_, i_11_, i_15_, n_n163}, x1832x);
	defparam lut_13929.LUT_SIZE = 7;
	defparam lut_13929.mask = 128'h33ffffff33ffffff0105040505000504;

	lut_sub lut_13941 ({sk[2832], n_n103, n_n57, n_n56, x3569x, x1833x, x1832x}, x21351x);
	defparam lut_13941.LUT_SIZE = 7;
	defparam lut_13941.mask = 128'h33ffffff33ffffff0f5f3f7f0fff3fff;

	lut_sub lut_13946 ({sk[2833], n_n222, x898x, x901x, x904x, n_n225, x158x}, x21869x);
	defparam lut_13946.LUT_SIZE = 7;
	defparam lut_13946.mask = 128'h33ffffff33ffffff557777775f7fffff;

	lut_sub lut_13952 ({sk[2834], i_14_, i_13_, i_12_, i_15_, n_n267, x363x}, x21870x);
	defparam lut_13952.LUT_SIZE = 7;
	defparam lut_13952.mask = 128'h33ffffff33ffffff5757755755557755;

	lut_sub lut_13960 ({sk[2835], i_14_, i_13_, i_12_, i_15_, n_n267, x21867x}, x1850x);
	defparam lut_13960.LUT_SIZE = 7;
	defparam lut_13960.mask = 128'h33ffffff33ffffff5757755755557755;

	lut_sub lut_13968 ({sk[2836], i_14_, i_13_, i_12_, i_15_, n_n282, x236x}, x1835x);
	defparam lut_13968.LUT_SIZE = 7;
	defparam lut_13968.mask = 128'h33ffffff33ffffff5757755755557755;

	lut_sub lut_13976 ({sk[2837], i_9_, i_10_, i_11_, i_15_, x154x, n_n256}, x339x);
	defparam lut_13976.LUT_SIZE = 7;
	defparam lut_13976.mask = 128'h33ffffff33ffffff3733333333333333;

	lut_sub lut_13979 ({sk[2838], i_14_, i_13_, i_12_, i_15_, n_n247, x339x}, x1834x);
	defparam lut_13979.LUT_SIZE = 7;
	defparam lut_13979.mask = 128'h33ffffff33ffffff5755755555555555;

	lut_sub lut_13983 ({sk[2839], i_9_, i_10_, i_14_, i_11_, i_15_, n_n254}, x22836x);
	defparam lut_13983.LUT_SIZE = 7;
	defparam lut_13983.mask = 128'h33ffffff33ffffff0000500000100001;

	lut_sub lut_13988 ({sk[2840], i_14_, i_13_, i_12_, i_15_, n_n247, x428x}, x21867x);
	defparam lut_13988.LUT_SIZE = 7;
	defparam lut_13988.mask = 128'h33ffffff33ffffff5757755555555555;

	lut_sub lut_13993 ({sk[2841], i_14_, i_13_, i_12_, x907x, x901x}, x291x);
	defparam lut_13993.LUT_SIZE = 6;
	defparam lut_13993.mask = 64'h77ff77ff00500300;

	lut_sub lut_13996 ({sk[2842], i_14_, i_13_, i_12_, x898x, x904x}, x1879x);
	defparam lut_13996.LUT_SIZE = 6;
	defparam lut_13996.mask = 64'h77ff77ff50300503;

	lut_sub lut_14001 ({sk[2843], i_14_, i_13_, i_12_, i_11_, i_15_, n_n274}, x1880x);
	defparam lut_14001.LUT_SIZE = 7;
	defparam lut_14001.mask = 128'h33ffffff33ffffff1050005050004040;

	lut_sub lut_14011 ({sk[2844], i_14_, i_13_, i_12_, i_15_, n_n247, x205x}, x1884x);
	defparam lut_14011.LUT_SIZE = 7;
	defparam lut_14011.mask = 128'h33ffffff33ffffff5555555557557575;

	lut_sub lut_14016 ({sk[2845], i_7_, i_5_, i_6_, i_3_, i_4_}, x1887x);
	defparam lut_14016.LUT_SIZE = 6;
	defparam lut_14016.mask = 64'h77ff77ffc08c0cc4;

	lut_sub lut_14025 ({sk[2846], i_14_, i_13_, i_12_, x903x, x897x}, x1919x);
	defparam lut_14025.LUT_SIZE = 6;
	defparam lut_14025.mask = 64'h77ff77ff53330000;

	lut_sub lut_14030 ({sk[2847], i_14_, i_13_, i_12_, i_15_, n_n275, x897x}, x1921x);
	defparam lut_14030.LUT_SIZE = 7;
	defparam lut_14030.mask = 128'h33ffffff33ffffff0000000003557530;

	lut_sub lut_14036 ({sk[2848], i_7_, i_8_, i_6_, x916x, x107x, x22836x}, x458x);
	defparam lut_14036.LUT_SIZE = 7;
	defparam lut_14036.mask = 128'h33ffffff33ffffff0000000700000000;

	lut_sub lut_14039 ({sk[2849], i_7_, i_8_, i_6_, x916x, x114x, x128x}, x607x);
	defparam lut_14039.LUT_SIZE = 7;
	defparam lut_14039.mask = 128'h33ffffff33ffffff0000000700000000;

	lut_sub lut_14042 ({sk[2850], i_7_, i_8_, i_6_, x909x, n_n240, n_n236}, x2319x);
	defparam lut_14042.LUT_SIZE = 7;
	defparam lut_14042.mask = 128'h33ffffff33ffffff0000000000070007;

	lut_sub lut_14047 ({sk[2851], i_9_, i_10_, i_11_, i_15_, n_n57, n_n258}, x2321x);
	defparam lut_14047.LUT_SIZE = 7;
	defparam lut_14047.mask = 128'h33ffffff33ffffff1000000000101000;

	lut_sub lut_14051 ({sk[2852], i_14_, i_13_, i_12_, x900x, x906x, x220x}, x22274x);
	defparam lut_14051.LUT_SIZE = 7;
	defparam lut_14051.mask = 128'h33ffffff33ffffff55555f5555775555;

	lut_sub lut_14055 ({sk[2853], i_7_, i_8_, i_6_, x909x, n_n62, n_n58}, x3096x);
	defparam lut_14055.LUT_SIZE = 7;
	defparam lut_14055.mask = 128'h33ffffff33ffffff0000000000070007;

	lut_sub lut_14060 ({sk[2854], i_9_, i_10_, i_11_, i_15_, n_n220, n_n56}, x3098x);
	defparam lut_14060.LUT_SIZE = 7;
	defparam lut_14060.mask = 128'h33ffffff33ffffff0000010001010000;

	lut_sub lut_14064 ({sk[2855], i_14_, i_13_, i_12_, n_n3, x900x}, x3192x);
	defparam lut_14064.LUT_SIZE = 6;
	defparam lut_14064.mask = 64'h77ff77ff00000010;

	lut_sub lut_14066 ({sk[2856], x915x, n_n273, n_n283, n_n220, x911x, x897x}, x3201x);
	defparam lut_14066.LUT_SIZE = 7;
	defparam lut_14066.mask = 128'h33ffffff33ffffff0000000000070707;

	lut_sub lut_14071 ({sk[2857], i_9_, i_10_, i_11_, i_15_, n_n1, n_n220}, x3203x);
	defparam lut_14071.LUT_SIZE = 7;
	defparam lut_14071.mask = 128'h33ffffff33ffffff0100000000010100;

	lut_sub lut_14075 ({sk[2858], i_9_, i_10_, i_11_, n_n263, x922x}, x3821x);
	defparam lut_14075.LUT_SIZE = 6;
	defparam lut_14075.mask = 64'h77ff77ff00001101;

	lut_sub lut_14079 ({sk[2859], i_14_, i_13_, i_12_, i_15_, n_n247, x160x}, x20511x);
	defparam lut_14079.LUT_SIZE = 7;
	defparam lut_14079.mask = 128'h33ffffff33ffffff7555575555555555;

	lut_sub lut_14083 ({sk[2860], n_n281, x183x, x159x, x901x, n_n228, x906x}, x24126x);
	defparam lut_14083.LUT_SIZE = 7;
	defparam lut_14083.mask = 128'h33ffffff33fffffffc000000a8000000;

	lut_sub lut_14088 ({sk[2861], i_7_, i_8_, i_6_, x909x, x72x}, x4763x);
	defparam lut_14088.LUT_SIZE = 6;
	defparam lut_14088.mask = 64'h77ff77ff00000100;

	lut_sub lut_14090 ({sk[2862], n_n2, x218x, x146x, x72x, n_n206, x118x}, x5153x);
	defparam lut_14090.LUT_SIZE = 7;
	defparam lut_14090.mask = 128'h33ffffff33ffffff000000007fffffff;

	lut_sub lut_14096 ({sk[2863], i_7_, i_8_, i_6_, n_n165, n_n106, n_n284}, x5444x);
	defparam lut_14096.LUT_SIZE = 7;
	defparam lut_14096.mask = 128'h33ffffff33ffffff0000010100000000;

	lut_sub lut_14099 ({sk[2864], n_n271, x896x, n_n220, x912x, x328x, x19237x}, x5848x);
	defparam lut_14099.LUT_SIZE = 7;
	defparam lut_14099.mask = 128'h33ffffff33ffffff000000000000777f;

	lut_sub lut_14103 ({sk[2865], i_7_, i_6_, i_4_, x910x, x259x, x1316x}, x19302x);
	defparam lut_14103.LUT_SIZE = 7;
	defparam lut_14103.mask = 128'h33ffffff33ffffff11001f0f1f0f1f0f;

	lut_sub lut_14107 ({sk[2866], i_9_, i_10_, x260x, n_n273, n_n283, x910x}, x24215x);
	defparam lut_14107.LUT_SIZE = 7;
	defparam lut_14107.mask = 128'h33ffffff33ffffffeeccfaf0faf0eac0;

	lut_sub lut_14113 ({sk[2867], i_9_, i_10_, i_12_, i_11_}, x19326x);
	defparam lut_14113.LUT_SIZE = 5;
	defparam lut_14113.mask = 32'h3f3f0770;

	lut_sub lut_14118 ({sk[2868], i_7_, i_8_, i_6_, x917x, n_n151, x927x}, x19369x);
	defparam lut_14118.LUT_SIZE = 7;
	defparam lut_14118.mask = 128'h33ffffff33ffffff55005703000f000f;

	lut_sub lut_14123 ({sk[2869], x917x, n_n312, n_n4476, x266x, x294x, n_n283}, x19373x);
	defparam lut_14123.LUT_SIZE = 7;
	defparam lut_14123.mask = 128'h33ffffff33ffffff00ffffff15ffffff;

	lut_sub lut_14128 ({sk[2870], i_14_, i_13_, i_12_, n_n273, x922x, x902x}, x19451x);
	defparam lut_14128.LUT_SIZE = 7;
	defparam lut_14128.mask = 128'h33ffffff33ffffff0101000101010100;

	lut_sub lut_14135 ({sk[2871], n_n7424, n_n6878, x438x, x626x, n_n2274, n_n639}, x19453x);
	defparam lut_14135.LUT_SIZE = 7;
	defparam lut_14135.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_14142 ({sk[2872], n_n1, n_n7402, n_n7407, x68x, x1877x, x19451x}, x19454x);
	defparam lut_14142.LUT_SIZE = 7;
	defparam lut_14142.mask = 128'h33ffffff33ffffff55ffffff7fffffff;

	lut_sub lut_14148 ({sk[2873], i_7_, i_8_, i_6_, n_n9, x909x, n_n59}, x19475x);
	defparam lut_14148.LUT_SIZE = 7;
	defparam lut_14148.mask = 128'h33ffffff33ffffff0013001300000000;

	lut_sub lut_14153 ({sk[2874], x909x, n_n261, n_n228, x897x, x50x, x19475x}, x19477x);
	defparam lut_14153.LUT_SIZE = 7;
	defparam lut_14153.mask = 128'h33ffffff33ffffff555555555555777f;

	lut_sub lut_14157 ({sk[2875], n_n5, x114x, x201x, n_n227, x156x, n_n3803}, x19478x);
	defparam lut_14157.LUT_SIZE = 7;
	defparam lut_14157.mask = 128'h33ffffff33ffffff555f5f5f777f7f7f;

	lut_sub lut_14162 ({sk[2876], n_n258, n_n100, n_n94, n_n225, x897x, x471x}, x19551x);
	defparam lut_14162.LUT_SIZE = 7;
	defparam lut_14162.mask = 128'h33ffffff33ffffff5557555755577777;

	lut_sub lut_14166 ({sk[2877], n_n863, x19554x, x768x, x383x, x380x, x19551x}, x19587x);
	defparam lut_14166.LUT_SIZE = 7;
	defparam lut_14166.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_14173 ({sk[2878], i_7_, i_6_, n_n118, n_n264, n_n284, n_n116}, x19642x);
	defparam lut_14173.LUT_SIZE = 7;
	defparam lut_14173.mask = 128'h33ffffff33ffffff0000000000330537;

	lut_sub lut_14177 ({sk[2879], i_5_, i_3_, i_4_, n_n118, x116x, x19642x}, x19643x);
	defparam lut_14177.LUT_SIZE = 7;
	defparam lut_14177.mask = 128'h33ffffff33ffffff5557555557575555;

	lut_sub lut_14182 ({sk[2880], i_7_, i_6_, x927x, n_n5672, x924x, x880x}, x24167x);
	defparam lut_14182.LUT_SIZE = 7;
	defparam lut_14182.mask = 128'h33ffffff33ffffffa0a080808000a0a0;

	lut_sub lut_14188 ({sk[2881], x146x, x909x, n_n261, n_n263, n_n11, x44x}, x19651x);
	defparam lut_14188.LUT_SIZE = 7;
	defparam lut_14188.mask = 128'h33ffffff33ffffff00000537000005ff;

	lut_sub lut_14192 ({sk[2882], x909x, n_n261, n_n263, x265x, n_n60, x137x}, x19652x);
	defparam lut_14192.LUT_SIZE = 7;
	defparam lut_14192.mask = 128'h33ffffff33ffffff00000000005f337f;

	lut_sub lut_14196 ({sk[2883], n_n12, x909x, n_n261, n_n263, x293x, x70x}, x19653x);
	defparam lut_14196.LUT_SIZE = 7;
	defparam lut_14196.mask = 128'h33ffffff33ffffff00000707000007ff;

	lut_sub lut_14200 ({sk[2884], i_7_, i_8_, i_6_, x909x, x265x, x498x}, x19654x);
	defparam lut_14200.LUT_SIZE = 7;
	defparam lut_14200.mask = 128'h33ffffff33ffffff5555555555555755;

	lut_sub lut_14203 ({sk[2885], x909x, n_n261, n_n263, x81x, n_n95, n_n49}, x19670x);
	defparam lut_14203.LUT_SIZE = 7;
	defparam lut_14203.mask = 128'h33ffffff33ffffff00000000000f777f;

	lut_sub lut_14207 ({sk[2886], x183x, n_n4223, n_n4224, x390x, x909x, n_n261}, x19761x);
	defparam lut_14207.LUT_SIZE = 7;
	defparam lut_14207.mask = 128'h33ffffff33ffffff0fffffff1fffffff;

	lut_sub lut_14212 ({sk[2887], x19659x, x19660x, x19651x, x19652x, x19653x, x19654x}, x19762x);
	defparam lut_14212.LUT_SIZE = 7;
	defparam lut_14212.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_14219 ({sk[2888], x915x, n_n273, n_n283, x81x, n_n42, n_n95}, x19796x);
	defparam lut_14219.LUT_SIZE = 7;
	defparam lut_14219.mask = 128'h33ffffff33ffffff00000000003f5f7f;

	lut_sub lut_14224 ({sk[2889], i_7_, i_8_, i_6_, x915x, x43x, x98x}, x19797x);
	defparam lut_14224.LUT_SIZE = 7;
	defparam lut_14224.mask = 128'h33ffffff33ffffff0300070000000000;

	lut_sub lut_14228 ({sk[2890], n_n151, x183x, n_n1, x5159x, x72x, x118x}, x19819x);
	defparam lut_14228.LUT_SIZE = 7;
	defparam lut_14228.mask = 128'h33ffffff33ffffff0f7f0fff0fff0fff;

	lut_sub lut_14234 ({sk[2891], n_n266, x916x, x268x, n_n280, x64x, x112x}, x19857x);
	defparam lut_14234.LUT_SIZE = 7;
	defparam lut_14234.mask = 128'h33ffffff33ffffff0000000000007fff;

	lut_sub lut_14239 ({sk[2892], i_9_, i_10_, n_n155, x924x, x260x, n_n283}, x19961x);
	defparam lut_14239.LUT_SIZE = 7;
	defparam lut_14239.mask = 128'h33ffffff33ffffff000f111f000f000f;

	lut_sub lut_14242 ({sk[2893], n_n4807, x390x, n_n5796, n_n5, x218x, n_n4809}, x19987x);
	defparam lut_14242.LUT_SIZE = 7;
	defparam lut_14242.mask = 128'h33ffffff33ffffff57ffffffffffffff;

	lut_sub lut_14248 ({sk[2894], x913x, n_n130, n_n220, n_n121, x914x, x905x}, x20011x);
	defparam lut_14248.LUT_SIZE = 7;
	defparam lut_14248.mask = 128'h33ffffff33ffffff00030077000300ff;

	lut_sub lut_14253 ({sk[2895], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, x20030x);
	defparam lut_14253.LUT_SIZE = 7;
	defparam lut_14253.mask = 128'h33ffffff33ffffff4040101000000000;

	lut_sub lut_14258 ({sk[2896], i_7_, i_6_, x927x, n_n5674, x260x, x20030x}, x20032x);
	defparam lut_14258.LUT_SIZE = 7;
	defparam lut_14258.mask = 128'h33ffffff33ffffff5fff7fff7f7f5f5f;

	lut_sub lut_14265 ({sk[2897], n_n151, n_n6843, n_n94, n_n6847, x601x, x377x}, x20111x);
	defparam lut_14265.LUT_SIZE = 7;
	defparam lut_14265.mask = 128'h33ffffff33ffffff3f7fffff3fffffff;

	lut_sub lut_14271 ({sk[2898], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, x20189x);
	defparam lut_14271.LUT_SIZE = 7;
	defparam lut_14271.mask = 128'h33ffffff33ffffff0050000000100000;

	lut_sub lut_14275 ({sk[2899], i_7_, i_8_, i_6_, x909x, x45x, x204x}, x20214x);
	defparam lut_14275.LUT_SIZE = 7;
	defparam lut_14275.mask = 128'h33ffffff33ffffff0000000000000007;

	lut_sub lut_14278 ({sk[2900], i_7_, i_6_, n_n118, n_n264, n_n284, n_n116}, x20236x);
	defparam lut_14278.LUT_SIZE = 7;
	defparam lut_14278.mask = 128'h33ffffff33ffffff0000003300000537;

	lut_sub lut_14282 ({sk[2901], i_7_, i_6_, x919x, x918x, x261x, x20236x}, x20237x);
	defparam lut_14282.LUT_SIZE = 7;
	defparam lut_14282.mask = 128'h33ffffff33ffffff55557fff55557fff;

	lut_sub lut_14290 ({sk[2902], n_n271, x896x, x371x, x20190x, x20189x, x20237x}, x20238x);
	defparam lut_14290.LUT_SIZE = 7;
	defparam lut_14290.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_14295 ({sk[2903], n_n103, n_n48, n_n53, x91x, x141x, x203x}, x20269x);
	defparam lut_14295.LUT_SIZE = 7;
	defparam lut_14295.mask = 128'h33ffffff33ffffff007f007f00ffffff;

	lut_sub lut_14301 ({sk[2904], n_n48, x40x, x479x, x478x, x1403x, x578x}, x20270x);
	defparam lut_14301.LUT_SIZE = 7;
	defparam lut_14301.mask = 128'h33ffffff33ffffff5fff5fff7fffffff;

	lut_sub lut_14307 ({sk[2905], n_n48, n_n53, x121x, n_n15, x1364x, x1476x}, x20293x);
	defparam lut_14307.LUT_SIZE = 7;
	defparam lut_14307.mask = 128'h33ffffff33ffffff00003fff5f5f7fff;

	lut_sub lut_14313 ({sk[2906], n_n281, x184x, x901x, x160x, n_n228, x906x}, x24133x);
	defparam lut_14313.LUT_SIZE = 7;
	defparam lut_14313.mask = 128'h33ffffff33fffffff0c00000a0800000;

	lut_sub lut_14318 ({sk[2907], n_n4, n_n7402, n_n13, n_n12, n_n7440, x20394x}, x24153x);
	defparam lut_14318.LUT_SIZE = 7;
	defparam lut_14318.mask = 128'h33ffffff33ffffff7777ffff7fffffff;

	lut_sub lut_14331 ({sk[2908], n_n4, n_n9, n_n65, n_n7425, x446x, x24153x}, x20410x);
	defparam lut_14331.LUT_SIZE = 7;
	defparam lut_14331.mask = 128'h33ffffff33ffffff7f7f7f7f7fffffff;

	lut_sub lut_14337 ({sk[2909], i_14_, i_13_, i_12_, i_15_, n_n267}, x20471x);
	defparam lut_14337.LUT_SIZE = 6;
	defparam lut_14337.mask = 64'h77ff77ff14041044;

	lut_sub lut_14344 ({sk[2910], i_7_, i_8_, i_6_, x922x, x111x, x406x}, x20478x);
	defparam lut_14344.LUT_SIZE = 7;
	defparam lut_14344.mask = 128'h33ffffff33ffffff5555575555555555;

	lut_sub lut_14347 ({sk[2911], x915x, n_n258, n_n261, x900x, x94x, x77x}, x20539x);
	defparam lut_14347.LUT_SIZE = 7;
	defparam lut_14347.mask = 128'h33ffffff33ffffff000000000077007f;

	lut_sub lut_14351 ({sk[2912], n_n4, x206x, n_n7402, n_n13, x410x, n_n12}, x20622x);
	defparam lut_14351.LUT_SIZE = 7;
	defparam lut_14351.mask = 128'h33ffffff33ffffff00ff00ff7fffffff;

	lut_sub lut_14357 ({sk[2913], i_7_, i_5_, i_6_, i_3_, i_4_, n_n116}, x24151x);
	defparam lut_14357.LUT_SIZE = 7;
	defparam lut_14357.mask = 128'h33ffffff33ffffffefffafffefffefff;

	lut_sub lut_14363 ({sk[2914], i_7_, i_8_, i_6_, x909x, x119x}, x20696x);
	defparam lut_14363.LUT_SIZE = 6;
	defparam lut_14363.mask = 64'h77ff77ff00000101;

	lut_sub lut_14366 ({sk[2915], n_n5796, n_n57, n_n56, x170x, x49x, x124x}, x20697x);
	defparam lut_14366.LUT_SIZE = 7;
	defparam lut_14366.mask = 128'h33ffffff33ffffff003f557fffffffff;

	lut_sub lut_14371 ({sk[2916], i_7_, i_8_, i_6_, x909x, x157x, x190x}, x24171x);
	defparam lut_14371.LUT_SIZE = 7;
	defparam lut_14371.mask = 128'h33ffffff33fffffffffffffffff8ffff;

	lut_sub lut_14377 ({sk[2917], n_n266, x909x, x140x, n_n4940, x167x, x24171x}, x20740x);
	defparam lut_14377.LUT_SIZE = 7;
	defparam lut_14377.mask = 128'h33ffffff33ffffffafafafafafafbfff;

	lut_sub lut_14382 ({sk[2918], n_n6, x183x, n_n4223, n_n4224, x390x, n_n5796}, x20748x);
	defparam lut_14382.LUT_SIZE = 7;
	defparam lut_14382.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_14388 ({sk[2919], x19659x, x19660x, x19651x, x19652x, x19653x, x19654x}, x20749x);
	defparam lut_14388.LUT_SIZE = 7;
	defparam lut_14388.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_14395 ({sk[2920], n_n4, x111x, x557x, n_n7345, n_n7344, x933x}, x20814x);
	defparam lut_14395.LUT_SIZE = 7;
	defparam lut_14395.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_14401 ({sk[2921], n_n3, n_n7224, n_n7225, n_n3418, x597x, x1579x}, x20817x);
	defparam lut_14401.LUT_SIZE = 7;
	defparam lut_14401.mask = 128'h33ffffff33ffffff3fffffff7fffffff;

	lut_sub lut_14407 ({sk[2922], x19390x, x19391x, x20810x, x20811x, x20814x}, x20818x);
	defparam lut_14407.LUT_SIZE = 6;
	defparam lut_14407.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_14413 ({sk[2923], n_n110, n_n273, n_n283, x258x, x922x, x82x}, x20822x);
	defparam lut_14413.LUT_SIZE = 7;
	defparam lut_14413.mask = 128'h33ffffff33ffffff0013001300133333;

	lut_sub lut_14417 ({sk[2924], n_n57, n_n226, n_n53, x111x, x579x, x309x}, x24197x);
	defparam lut_14417.LUT_SIZE = 7;
	defparam lut_14417.mask = 128'h33ffffff33ffffff8880888088800000;

	lut_sub lut_14422 ({sk[2925], n_n283, x159x, x922x, n_n6875, x475x, n_n6879}, x20853x);
	defparam lut_14422.LUT_SIZE = 7;
	defparam lut_14422.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_14427 ({sk[2926], n_n7441, n_n53, n_n6868, n_n71, x475x, x634x}, x20904x);
	defparam lut_14427.LUT_SIZE = 7;
	defparam lut_14427.mask = 128'h33ffffff33ffffff77ff7fffffffffff;

	lut_sub lut_14433 ({sk[2927], n_n4, x476x, n_n1356, x5683x, x5682x, x1787x}, x20909x);
	defparam lut_14433.LUT_SIZE = 7;
	defparam lut_14433.mask = 128'h33ffffff33ffffff3fffffff7fffffff;

	lut_sub lut_14439 ({sk[2928], n_n7440, n_n7442, n_n7443, x866x, x20909x}, x20910x);
	defparam lut_14439.LUT_SIZE = 6;
	defparam lut_14439.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_14445 ({sk[2929], x19440x, n_n3435, x20905x, x19438x, x19439x, x20904x}, x20911x);
	defparam lut_14445.LUT_SIZE = 7;
	defparam lut_14445.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_14452 ({sk[2930], n_n6, n_n5, x159x, x522x, x523x, x208x}, x20955x);
	defparam lut_14452.LUT_SIZE = 7;
	defparam lut_14452.mask = 128'h33ffffff33ffffff3f3f7f7f3fff7fff;

	lut_sub lut_14457 ({sk[2931], n_n281, x909x, x905x, n_n263, x685x}, x20982x);
	defparam lut_14457.LUT_SIZE = 6;
	defparam lut_14457.mask = 64'h77ff77ff55555557;

	lut_sub lut_14460 ({sk[2932], n_n9, n_n257, n_n6830, x278x, x655x, x20982x}, x20984x);
	defparam lut_14460.LUT_SIZE = 7;
	defparam lut_14460.mask = 128'h33ffffff33ffffff77ff7fff7fff7fff;

	lut_sub lut_14466 ({sk[2933], n_n4, n_n9, n_n7407, x409x, x476x, x446x}, x20993x);
	defparam lut_14466.LUT_SIZE = 7;
	defparam lut_14466.mask = 128'h33ffffff33ffffff7fff7fff7fffffff;

	lut_sub lut_14472 ({sk[2934], n_n3, n_n7425, n_n7440, n_n15, x20394x, x1914x}, x20994x);
	defparam lut_14472.LUT_SIZE = 7;
	defparam lut_14472.mask = 128'h33ffffff33ffffff33ffffff7fffffff;

	lut_sub lut_14478 ({sk[2935], n_n283, x170x, x922x, n_n76, x49x, x207x}, x21058x);
	defparam lut_14478.LUT_SIZE = 7;
	defparam lut_14478.mask = 128'h33ffffff33ffffff00000000007f00ff;

	lut_sub lut_14483 ({sk[2936], n_n48, n_n53, x111x, x163x, x478x, x20344x}, x24156x);
	defparam lut_14483.LUT_SIZE = 7;
	defparam lut_14483.mask = 128'h33ffffff33ffffff8888880080808000;

	lut_sub lut_14488 ({sk[2937], n_n6, n_n5, x188x, x1325x, x1324x, x1946x}, x21126x);
	defparam lut_14488.LUT_SIZE = 7;
	defparam lut_14488.mask = 128'h33ffffff33ffffff000033335fff7fff;

	lut_sub lut_14493 ({sk[2938], n_n3172, x20956x, n_n3167, x3870x, x20955x, x20984x}, x21128x);
	defparam lut_14493.LUT_SIZE = 7;
	defparam lut_14493.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_14500 ({sk[2939], n_n3964, x736x, x20392x, x876x, x20993x, x20994x}, x24198x);
	defparam lut_14500.LUT_SIZE = 7;
	defparam lut_14500.mask = 128'h33ffffff33ffffff8000000000000000;

	lut_sub lut_14502 ({sk[2940], n_n4, n_n9, n_n3, x439x, x648x, x953x}, x21151x);
	defparam lut_14502.LUT_SIZE = 7;
	defparam lut_14502.mask = 128'h33ffffff33ffffff3f7f3f7f3f7fffff;

	lut_sub lut_14507 ({sk[2941], i_7_, i_6_, n_n264, x918x, x879x, n_n116}, x21171x);
	defparam lut_14507.LUT_SIZE = 7;
	defparam lut_14507.mask = 128'h33ffffff33ffffff3f3f333333773377;

	lut_sub lut_14512 ({sk[2942], i_7_, i_8_, i_6_, x917x, x211x, n_n133}, x24149x);
	defparam lut_14512.LUT_SIZE = 7;
	defparam lut_14512.mask = 128'h33ffffff33fffffffcfafffffff0fff0;

	lut_sub lut_14520 ({sk[2943], n_n4, n_n7402, n_n12, n_n3, x176x, x546x}, x21200x);
	defparam lut_14520.LUT_SIZE = 7;
	defparam lut_14520.mask = 128'h33ffffff33ffffff575fffff57ffffff;

	lut_sub lut_14526 ({sk[2944], n_n208, x916x, n_n9, n_n3, x159x, n_n61}, x21239x);
	defparam lut_14526.LUT_SIZE = 7;
	defparam lut_14526.mask = 128'h33ffffff33ffffff03030303030357ff;

	lut_sub lut_14530 ({sk[2945], n_n281, n_n4, x206x, n_n3, x914x, x290x}, x21240x);
	defparam lut_14530.LUT_SIZE = 7;
	defparam lut_14530.mask = 128'h33ffffff33ffffff000f555f030f575f;

	lut_sub lut_14534 ({sk[2946], n_n266, x909x, x159x, n_n7, x899x, n_n228}, x21362x);
	defparam lut_14534.LUT_SIZE = 7;
	defparam lut_14534.mask = 128'h33ffffff33ffffff0000000000001fff;

	lut_sub lut_14538 ({sk[2947], n_n208, x916x, n_n3, n_n60, n_n223, x253x}, x21430x);
	defparam lut_14538.LUT_SIZE = 7;
	defparam lut_14538.mask = 128'h33ffffff33ffffff0055005500553f7f;

	lut_sub lut_14542 ({sk[2948], n_n281, x905x, n_n53, x908x, x413x, x369x}, x24108x);
	defparam lut_14542.LUT_SIZE = 7;
	defparam lut_14542.mask = 128'h33ffffff33ffffffff88ff88ff80ff00;

	lut_sub lut_14546 ({sk[2949], n_n266, n_n271, x909x, n_n7, n_n186, n_n53}, x21497x);
	defparam lut_14546.LUT_SIZE = 7;
	defparam lut_14546.mask = 128'h33ffffff33ffffff1111111f111f111f;

	lut_sub lut_14550 ({sk[2950], x915x, n_n261, n_n263, n_n35, x382x, x330x}, x24111x);
	defparam lut_14550.LUT_SIZE = 7;
	defparam lut_14550.mask = 128'h33ffffff33ffffffcccccccccc88c080;

	lut_sub lut_14556 ({sk[2951], n_n106, x909x, n_n145, n_n261, n_n263, n_n60}, x21532x);
	defparam lut_14556.LUT_SIZE = 7;
	defparam lut_14556.mask = 128'h33ffffff33ffffff0000050f00003f3f;

	lut_sub lut_14561 ({sk[2952], n_n6, n_n5, x307x, x411x, x1034x, x1486x}, x21556x);
	defparam lut_14561.LUT_SIZE = 7;
	defparam lut_14561.mask = 128'h33ffffff33ffffff0f0f3f3f5fff7fff;

	lut_sub lut_14566 ({sk[2953], n_n48, n_n53, n_n223, n_n171, x1529x, x1527x}, x21611x);
	defparam lut_14566.LUT_SIZE = 7;
	defparam lut_14566.mask = 128'h33ffffff33ffffff00003fff55557fff;

	lut_sub lut_14571 ({sk[2954], n_n281, x913x, n_n208, x916x, n_n3, x905x}, x21614x);
	defparam lut_14571.LUT_SIZE = 7;
	defparam lut_14571.mask = 128'h33ffffff33ffffff000000001111333f;

	lut_sub lut_14575 ({sk[2955], x21372x, x21373x, x21525x, n_n2099, n_n2100, x21614x}, x21616x);
	defparam lut_14575.LUT_SIZE = 7;
	defparam lut_14575.mask = 128'h33ffffff33ffffff7fffffffffffffff;

	lut_sub lut_14582 ({sk[2956], n_n151, x295x, n_n126, n_n5769, n_n127, n_n5660}, x21630x);
	defparam lut_14582.LUT_SIZE = 7;
	defparam lut_14582.mask = 128'h33ffffff33ffffff5f5f7f7f5fff7fff;

	lut_sub lut_14587 ({sk[2957], i_7_, i_8_, i_6_, x909x, n_n80, n_n144}, x21814x);
	defparam lut_14587.LUT_SIZE = 7;
	defparam lut_14587.mask = 128'h33ffffff33ffffff0003000005000500;

	lut_sub lut_14591 ({sk[2958], n_n111, n_n48, n_n53, n_n6511, n_n6512, x249x}, x24194x);
	defparam lut_14591.LUT_SIZE = 7;
	defparam lut_14591.mask = 128'h33ffffff33ffffffc080c080c0800000;

	lut_sub lut_14596 ({sk[2959], n_n273, n_n283, x922x, n_n80, x102x, x24194x}, x21853x);
	defparam lut_14596.LUT_SIZE = 7;
	defparam lut_14596.mask = 128'h33ffffff33ffffffaaaaaabbaaafaabf;

	lut_sub lut_14600 ({sk[2960], n_n281, x913x, n_n152, x211x, n_n142, x914x}, x24148x);
	defparam lut_14600.LUT_SIZE = 7;
	defparam lut_14600.mask = 128'h33ffffff33fffffffff0fff0eee0ccc0;

	lut_sub lut_14607 ({sk[2961], n_n220, n_n4, n_n3, x911x, x899x, x1823x}, x21897x);
	defparam lut_14607.LUT_SIZE = 7;
	defparam lut_14607.mask = 128'h33ffffff33ffffff00005555000f7f7f;

	lut_sub lut_14612 ({sk[2962], i_15_, n_n4, n_n3, x957x, x154x, n_n137}, x21900x);
	defparam lut_14612.LUT_SIZE = 7;
	defparam lut_14612.mask = 128'h33ffffff33ffffff00330f3f00770f7f;

	lut_sub lut_14616 ({sk[2963], n_n3, x21885x, x21886x, n_n1724, x1824x, x21897x}, x21903x);
	defparam lut_14616.LUT_SIZE = 7;
	defparam lut_14616.mask = 128'h33ffffff33ffffff5fffffff7fffffff;

	lut_sub lut_14622 ({sk[2964], n_n4, n_n7402, n_n3, n_n258, x906x, x73x}, x24083x);
	defparam lut_14622.LUT_SIZE = 7;
	defparam lut_14622.mask = 128'h33ffffff33ffffffffaa0000fca80000;

	lut_sub lut_14629 ({sk[2965], n_n208, x916x, n_n7406, n_n7405, x1389x, x24083x}, x21925x);
	defparam lut_14629.LUT_SIZE = 7;
	defparam lut_14629.mask = 128'h33ffffff33ffffffafffafffafffbfff;

	lut_sub lut_14634 ({sk[2966], n_n1, n_n2, n_n220, n_n257, x899x, x75x}, x24087x);
	defparam lut_14634.LUT_SIZE = 7;
	defparam lut_14634.mask = 128'h33ffffff33ffffff00005f7f55775f7f;

	lut_sub lut_14645 ({sk[2967], n_n1, n_n2, n_n62, n_n10, x680x, x24087x}, x21990x);
	defparam lut_14645.LUT_SIZE = 7;
	defparam lut_14645.mask = 128'h33ffffff33ffffff77777fff7f7f7fff;

	lut_sub lut_14651 ({sk[2968], n_n1, n_n2, x1421x, x1420x, x1427x, x1426x}, x21991x);
	defparam lut_14651.LUT_SIZE = 7;
	defparam lut_14651.mask = 128'h33ffffff33ffffff00005f5f33ff7fff;

	lut_sub lut_14656 ({sk[2969], n_n1, n_n2, n_n42, x68x, x43x, x1387x}, x22061x);
	defparam lut_14656.LUT_SIZE = 7;
	defparam lut_14656.mask = 128'h33ffffff33ffffff00007f7f00ff7fff;

	lut_sub lut_14661 ({sk[2970], i_14_, i_13_, i_12_, x915x, n_n263, x903x}, x22082x);
	defparam lut_14661.LUT_SIZE = 7;
	defparam lut_14661.mask = 128'h33ffffff33ffffff0000000001000100;

	lut_sub lut_14664 ({sk[2971], n_n281, n_n208, x916x, x899x, n_n228, x906x}, x22090x);
	defparam lut_14664.LUT_SIZE = 7;
	defparam lut_14664.mask = 128'h33ffffff33ffffff000000110000001f;

	lut_sub lut_14667 ({sk[2972], n_n208, x916x, x94x, x333x, x455x, x22090x}, x22093x);
	defparam lut_14667.LUT_SIZE = 7;
	defparam lut_14667.mask = 128'h33ffffff33ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_14672 ({sk[2973], n_n6, n_n5, n_n246, n_n147, x1456x, x291x}, x22097x);
	defparam lut_14672.LUT_SIZE = 7;
	defparam lut_14672.mask = 128'h33ffffff33ffffff00005fff33337fff;

	lut_sub lut_14677 ({sk[2974], i_7_, i_8_, i_6_, x922x, x163x, x1002x}, x22174x);
	defparam lut_14677.LUT_SIZE = 7;
	defparam lut_14677.mask = 128'h33ffffff33ffffff0300050000000000;

	lut_sub lut_14680 ({sk[2975], n_n31, n_n48, n_n22, x4600x, x5627x, x1003x}, x22175x);
	defparam lut_14680.LUT_SIZE = 7;
	defparam lut_14680.mask = 128'h33ffffff33ffffff3f3f7fff3f3fffff;

	lut_sub lut_14686 ({sk[2976], i_9_, i_10_, i_11_, i_15_, n_n220, n_n258}, x24090x);
	defparam lut_14686.LUT_SIZE = 7;
	defparam lut_14686.mask = 128'h33ffffff33ffffffacffffacacacffac;

	lut_sub lut_14692 ({sk[2977], n_n222, x76x, n_n53, x900x, x43x, x416x}, x22300x);
	defparam lut_14692.LUT_SIZE = 7;
	defparam lut_14692.mask = 128'h33ffffff33ffffff007700ff007f00ff;

	lut_sub lut_14697 ({sk[2978], x51x, x81x, n_n48, x619x, x5574x, x1177x}, x22301x);
	defparam lut_14697.LUT_SIZE = 7;
	defparam lut_14697.mask = 128'h33ffffff33ffffff3f7f3fff3fff3fff;

	lut_sub lut_14703 ({sk[2979], i_7_, i_8_, i_6_, x915x, n_n258, x897x}, x22384x);
	defparam lut_14703.LUT_SIZE = 7;
	defparam lut_14703.mask = 128'h33ffffff33ffffff0000000001000100;

	lut_sub lut_14706 ({sk[2980], n_n31, n_n216, n_n94, x552x, x140x, x182x}, x22391x);
	defparam lut_14706.LUT_SIZE = 7;
	defparam lut_14706.mask = 128'h33ffffff33ffffff0f7f0fff0fff0fff;

	lut_sub lut_14712 ({sk[2981], n_n100, x1070x, x182x, x658x, n_n707, x22384x}, x22392x);
	defparam lut_14712.LUT_SIZE = 7;
	defparam lut_14712.mask = 128'h33ffffff33ffffff7f7f7f7f7fffffff;

	lut_sub lut_14718 ({sk[2982], n_n1, n_n2, n_n13, n_n246, n_n10, n_n252}, x22541x);
	defparam lut_14718.LUT_SIZE = 7;
	defparam lut_14718.mask = 128'h33ffffff33ffffff000033ff7fff7fff;

	lut_sub lut_14725 ({sk[2983], n_n4, n_n13, n_n3, n_n7224, n_n70, n_n49}, x24078x);
	defparam lut_14725.LUT_SIZE = 7;
	defparam lut_14725.mask = 128'h33ffffff33fffffff0a0f0a0c0800000;

	lut_sub lut_14730 ({sk[2984], x913x, n_n4, n_n3, x905x, n_n258, x908x}, x22591x);
	defparam lut_14730.LUT_SIZE = 7;
	defparam lut_14730.mask = 128'h33ffffff33ffffff0013031300333333;

	lut_sub lut_14736 ({sk[2985], x907x, n_n4, n_n3, x914x, n_n258, x903x}, x24075x);
	defparam lut_14736.LUT_SIZE = 7;
	defparam lut_14736.mask = 128'h33ffffff33ffffffffecececffcccccc;

	lut_sub lut_14740 ({sk[2986], n_n4, n_n13, n_n7405, n_n7425, x22591x, x24075x}, x22592x);
	defparam lut_14740.LUT_SIZE = 7;
	defparam lut_14740.mask = 128'h33ffffff33ffffffbfffbfffbfffffff;

	lut_sub lut_14746 ({sk[2987], n_n41, n_n54, n_n48, n_n53, n_n105, x1699x}, x22714x);
	defparam lut_14746.LUT_SIZE = 7;
	defparam lut_14746.mask = 128'h33ffffff33ffffff070707ff0f0f0fff;

	lut_sub lut_14751 ({sk[2988], n_n104, n_n48, n_n53, x177x, x1494x, x1698x}, x22715x);
	defparam lut_14751.LUT_SIZE = 7;
	defparam lut_14751.mask = 128'h33ffffff33ffffff00335f7f0033ffff;

	lut_sub lut_14756 ({sk[2989], n_n208, x916x, n_n3, n_n105, x134x, x1720x}, x22818x);
	defparam lut_14756.LUT_SIZE = 7;
	defparam lut_14756.mask = 128'h33ffffff33ffffff0055005500553f7f;

	lut_sub lut_14760 ({sk[2990], n_n208, x916x, n_n31, n_n3, x126x, x960x}, x22843x);
	defparam lut_14760.LUT_SIZE = 7;
	defparam lut_14760.mask = 128'h33ffffff33ffffff05050505050537ff;

	lut_sub lut_14764 ({sk[2991], x22602x, x22603x, x22839x, n_n775, x458x}, x22846x);
	defparam lut_14764.LUT_SIZE = 6;
	defparam lut_14764.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_14770 ({sk[2992], n_n266, n_n271, x909x, n_n137, x494x, x172x}, x24102x);
	defparam lut_14770.LUT_SIZE = 7;
	defparam lut_14770.mask = 128'h33ffffff33ffffffffffff88fff0ff80;

	lut_sub lut_14776 ({sk[2993], n_n266, n_n271, x909x, n_n42, n_n95, x494x}, x24159x);
	defparam lut_14776.LUT_SIZE = 7;
	defparam lut_14776.mask = 128'h33ffffff33ffffffffffffccffa0ff80;


endmodule