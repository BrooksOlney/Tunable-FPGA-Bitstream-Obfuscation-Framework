module s298x6xv (s298_in_0_, s298_in_2_, s298_in_1_, clock, s298_out_0_, s298_out_1_, s298_out_2_, s298_out_3_, s298_out_4_, s298_out_5_);

	input s298_in_0_;
	input s298_in_2_;
	input s298_in_1_;
	input clock;
	output s298_out_0_;
	output s298_out_1_;
	output s298_out_2_;
	output s298_out_3_;
	output s298_out_4_;
	output s298_out_5_;

	wire [978 : 0] sk /* synthesis noprune */;

	lut_sub lut_11 ({sk[0], n_n854, n_n855, n_n856, n_n857, n_n858, n_n859}, s298_out_0_);
	defparam lut_11.LUT_SIZE = 7;
	defparam lut_11.mask = 128'h37373737373737374445444444674444;

	lut_sub lut_15 ({sk[1], n_n854, n_n855, n_n856, n_n857, n_n858, n_n859}, s298_out_1_);
	defparam lut_15.LUT_SIZE = 7;
	defparam lut_15.mask = 128'h1155ffffffffffff2020202220002022;

	lut_sub lut_20 ({sk[2], n_n855, n_n856, n_n857, n_n858, n_n859}, s298_out_2_);
	defparam lut_20.LUT_SIZE = 6;
	defparam lut_20.mask = 64'h5f5f5f5f131a131b;

	lut_sub lut_27 ({sk[3], n_n856, n_n857, n_n858, n_n859}, s298_out_3_);
	defparam lut_27.LUT_SIZE = 5;
	defparam lut_27.mask = 32'h37ff0200;

	lut_sub lut_29 ({sk[4], n_n855, n_n856, n_n857, n_n858, n_n859}, s298_out_4_);
	defparam lut_29.LUT_SIZE = 6;
	defparam lut_29.mask = 64'h5f5f5f5f111a111b;

	lut_sub lut_35 ({sk[5], n_n855, n_n856, n_n857, n_n858, n_n859}, s298_out_5_);
	defparam lut_35.LUT_SIZE = 6;
	defparam lut_35.mask = 64'h5f5f5f5f64656464;

	lut_sub lut_39 ({sk[6], x7228x, x7229x, x7230x, x7231x, x7232x}, n_n45);
	defparam lut_39.LUT_SIZE = 6;
	defparam lut_39.mask = 64'h5f5f5f5f7fffffff;

	lut_sub lut_45 ({sk[7], x8000x, x8001x, x8002x, x8003x, x8004x}, n_n46);
	defparam lut_45.LUT_SIZE = 6;
	defparam lut_45.mask = 64'h0f0fffff7fffffff;

	lut_sub lut_51 ({sk[8], x8741x, x8742x, x8743x, x8744x, x8745x, x8746x}, n_n47);
	defparam lut_51.LUT_SIZE = 7;
	defparam lut_51.mask = 128'h33333333ffffffff7fffffffffffffff;

	lut_sub lut_58 ({sk[9], x9156x, x9157x, x9158x, x9159x}, n_n48);
	defparam lut_58.LUT_SIZE = 5;
	defparam lut_58.mask = 32'h01ff7fff;

	lut_sub lut_63 ({sk[10], x6375x, x6355x, x6356x, x6357x, x6358x, x6374x}, n_n49);
	defparam lut_63.LUT_SIZE = 7;
	defparam lut_63.mask = 128'h33333333ffffffff7fffffffffffffff;

	lut_sub lut_70 ({sk[11], x6018x, x510x, x511x, x513x, x518x, x6017x}, n_n50);
	defparam lut_70.LUT_SIZE = 7;
	defparam lut_70.mask = 128'h33333333ffffffff7fffffffffffffff;

	lut_sub lut_77 ({sk[12], x5705x, x5676x, x5677x, x5693x, x5701x}, n_n51);
	defparam lut_77.LUT_SIZE = 6;
	defparam lut_77.mask = 64'h0f0fffff7fffffff;

	lut_sub lut_83 ({sk[13], x5785x, x5786x, x5787x, x5788x, x5789x}, n_n52);
	defparam lut_83.LUT_SIZE = 6;
	defparam lut_83.mask = 64'h33ff33ff7fffffff;

	lut_sub lut_89 ({sk[14], n_n49, x6384x, x7092x, x7096x, x441x, x7200x}, x7228x);
	defparam lut_89.LUT_SIZE = 7;
	defparam lut_89.mask = 128'h0f0fffff0f0fffff7777ffff7fff7fff;

	lut_sub lut_95 ({sk[15], n_n49, x6421x, x6428x, x7202x, x7204x, x7205x}, x7229x);
	defparam lut_95.LUT_SIZE = 7;
	defparam lut_95.mask = 128'h0f0fffff0f0fffff7fffffff7f7f7f7f;

	lut_sub lut_101 ({sk[16], x7206x, x7207x, x7208x, x7209x}, x7230x);
	defparam lut_101.LUT_SIZE = 5;
	defparam lut_101.mask = 32'h57ff7fff;

	lut_sub lut_106 ({sk[17], n_n49, x6974x, x6979x, x7210x, x7211x, x7212x}, x7231x);
	defparam lut_106.LUT_SIZE = 7;
	defparam lut_106.mask = 128'h555555ffffffffff7f7fffff7fff7fff;

	lut_sub lut_112 ({sk[18], n_n49, x7004x, x7009x, x7014x, x7088x, x12832x}, x7232x);
	defparam lut_112.LUT_SIZE = 7;
	defparam lut_112.mask = 128'h555555ffffffffffbbbbbbbbafffffff;

	lut_sub lut_118 ({sk[19], n_n49, x7970x, x7971x, x7972x, x12831x}, x8000x);
	defparam lut_118.LUT_SIZE = 6;
	defparam lut_118.mask = 64'h33ffffffbfff3fff;

	lut_sub lut_123 ({sk[20], n_n49, x7744x, x7749x, x7974x, x7975x, x7976x}, x8001x);
	defparam lut_123.LUT_SIZE = 7;
	defparam lut_123.mask = 128'h555555ffffffffff7fffffff7f7f7f7f;

	lut_sub lut_129 ({sk[21], n_n49, x7774x, x7779x, x7784x, x7789x, x12830x}, x8002x);
	defparam lut_129.LUT_SIZE = 7;
	defparam lut_129.mask = 128'h555555ffffffffffaaaaaaaabfffffff;

	lut_sub lut_135 ({sk[22], n_n49, x7853x, x7857x, x7861x, x7865x, x12829x}, x8003x);
	defparam lut_135.LUT_SIZE = 7;
	defparam lut_135.mask = 128'h555555ffffffffffaaaaaaaabfffffff;

	lut_sub lut_141 ({sk[23], x7967x, x7968x, x7969x, x7987x, x12824x}, x8004x);
	defparam lut_141.LUT_SIZE = 6;
	defparam lut_141.mask = 64'h33ffffffbfffffff;

	lut_sub lut_147 ({sk[24], x8705x, x8706x, x8707x, x8708x}, x8741x);
	defparam lut_147.LUT_SIZE = 5;
	defparam lut_147.mask = 32'h57ff7fff;

	lut_sub lut_152 ({sk[25], x8709x, x8710x, x8711x, x8712x}, x8742x);
	defparam lut_152.LUT_SIZE = 5;
	defparam lut_152.mask = 32'h57ff7fff;

	lut_sub lut_157 ({sk[26], n_n49, x8444x, x8449x, x8713x, x8714x, x8715x}, x8743x);
	defparam lut_157.LUT_SIZE = 7;
	defparam lut_157.mask = 128'h555555ffffffffff7fffffff7f7f7f7f;

	lut_sub lut_163 ({sk[27], n_n49, x8474x, x8479x, x8484x, x8489x, x12820x}, x8744x);
	defparam lut_163.LUT_SIZE = 7;
	defparam lut_163.mask = 128'h555555ffffffffffaaaaaaaabfffffff;

	lut_sub lut_169 ({sk[28], n_n49, x8514x, x8519x, x8573x, x8577x, x12819x}, x8745x);
	defparam lut_169.LUT_SIZE = 7;
	defparam lut_169.mask = 128'h0f0f0fff3f3f3fffbfbfbfbfaaffffff;

	lut_sub lut_175 ({sk[29], n_n49, x8597x, x8601x, x8605x, x8609x, x12818x}, x8746x);
	defparam lut_175.LUT_SIZE = 7;
	defparam lut_175.mask = 128'h0f0f0fff3f3f3fffaaaaaaaabfffffff;

	lut_sub lut_181 ({sk[30], x9132x, x9133x, x9134x, x9135x}, x9156x);
	defparam lut_181.LUT_SIZE = 5;
	defparam lut_181.mask = 32'h5f7f7fff;

	lut_sub lut_186 ({sk[31], n_n49, x8920x, x8925x, x8930x, x8935x, x12817x}, x9157x);
	defparam lut_186.LUT_SIZE = 7;
	defparam lut_186.mask = 128'h0f3fffff0f3fffffaaaaffffbfffbfff;

	lut_sub lut_192 ({sk[32], n_n49, x9022x, x9026x, x9030x, x9034x, x12816x}, x9158x);
	defparam lut_192.LUT_SIZE = 7;
	defparam lut_192.mask = 128'h0f3fffff0f3fffffaaaaffffbfffbfff;

	lut_sub lut_198 ({sk[33], x9130x, x9131x, x9144x, x9145x, x9146x}, x9159x);
	defparam lut_198.LUT_SIZE = 6;
	defparam lut_198.mask = 64'h333333337fffffff;

	lut_sub lut_204 ({sk[34], x6365x, x6366x, x12843x}, x6375x);
	defparam lut_204.LUT_SIZE = 4;
	defparam lut_204.mask = 16'h5fbf;

	lut_sub lut_208 ({sk[35], x6018x, x6025x, x6016x, x6017x, x6352x, x6353x}, x6355x);
	defparam lut_208.LUT_SIZE = 7;
	defparam lut_208.mask = 128'h0f3fffff0f3fffff7777f77777777777;

	lut_sub lut_212 ({sk[36], n_n52, x6018x, x6031x, x6016x, x6017x, x6036x}, x6356x);
	defparam lut_212.LUT_SIZE = 7;
	defparam lut_212.mask = 128'h00ff00ffffffffff40c0000000c00000;

	lut_sub lut_215 ({sk[37], s298_out_4_, x6018x, x6016x, x6017x, x6042x, x6048x}, x6357x);
	defparam lut_215.LUT_SIZE = 7;
	defparam lut_215.mask = 128'h00ff00ffffffffff0000000070000000;

	lut_sub lut_218 ({sk[38], s298_out_0_, x6018x, x6055x, x6016x, x6017x, x6060x}, x6358x);
	defparam lut_218.LUT_SIZE = 7;
	defparam lut_218.mask = 128'h00ff00ffffffffff00c0000015d55555;

	lut_sub lut_223 ({sk[39], x6359x, x6360x, x6361x, x6362x}, x6374x);
	defparam lut_223.LUT_SIZE = 5;
	defparam lut_223.mask = 32'h33ff7fff;

	lut_sub lut_228 ({sk[40], x536x, x542x, x544x, x6007x, x6008x}, x6018x);
	defparam lut_228.LUT_SIZE = 6;
	defparam lut_228.mask = 64'h5f5f5f5f7fffffff;

	lut_sub lut_234 ({sk[41], x5824x, x5785x, x5786x, x5787x, x5788x, x5789x}, x510x);
	defparam lut_234.LUT_SIZE = 7;
	defparam lut_234.mask = 128'h00ff00ffffffffff0000000080000000;

	lut_sub lut_236 ({sk[42], x5830x, x5785x, x5786x, x5787x, x5788x, x5789x}, x511x);
	defparam lut_236.LUT_SIZE = 7;
	defparam lut_236.mask = 128'h00ff00ffffffffff0000000080000000;

	lut_sub lut_238 ({sk[43], x5842x, x5785x, x5786x, x5787x, x5788x, x5789x}, x513x);
	defparam lut_238.LUT_SIZE = 7;
	defparam lut_238.mask = 128'h00ff00ffffffffff0000000080000000;

	lut_sub lut_240 ({sk[44], x5868x, x5785x, x5786x, x5787x, x5788x, x5789x}, x518x);
	defparam lut_240.LUT_SIZE = 7;
	defparam lut_240.mask = 128'h77ff77ff77ff77ff000000007fffffff;

	lut_sub lut_246 ({sk[45], x519x, x526x, x531x, x535x}, x6017x);
	defparam lut_246.LUT_SIZE = 5;
	defparam lut_246.mask = 32'h5fff7fff;

	lut_sub lut_251 ({sk[46], x603x, x604x, x5687x, x5696x, x5703x}, x5705x);
	defparam lut_251.LUT_SIZE = 6;
	defparam lut_251.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_257 ({sk[47], x5548x, x5549x, x5554x, x5555x}, x5676x);
	defparam lut_257.LUT_SIZE = 5;
	defparam lut_257.mask = 32'h5fff111f;

	lut_sub lut_260 ({sk[48], n_n854, n_n855, n_n856, n_n857, x5560x, x5566x}, x5677x);
	defparam lut_260.LUT_SIZE = 7;
	defparam lut_260.mask = 128'h77ff77ff77ff77ff0003000000050000;

	lut_sub lut_263 ({sk[49], x5572x, x5573x, x5578x, x5579x, x589x, x590x}, x5693x);
	defparam lut_263.LUT_SIZE = 7;
	defparam lut_263.mask = 128'h77ff77ff77ff77ff777f777f777fffff;

	lut_sub lut_268 ({sk[50], x591x, x592x, x595x, x596x, x5681x, x5683x}, x5701x);
	defparam lut_268.LUT_SIZE = 7;
	defparam lut_268.mask = 128'h77ff77ff77ff77ff7fffffffffffffff;

	lut_sub lut_275 ({sk[51], s298_out_0_, n_n854, n_n855, n_n51}, x5785x);
	defparam lut_275.LUT_SIZE = 5;
	defparam lut_275.mask = 32'h5fff00a2;

	lut_sub lut_278 ({sk[52], n_n51, x548x, x5772x, x5775x, x12837x}, x5786x);
	defparam lut_278.LUT_SIZE = 6;
	defparam lut_278.mask = 64'h3f3f3f3fbfff3fff;

	lut_sub lut_283 ({sk[53], x550x, x556x, x558x, x5767x, x5768x, x5780x}, x5787x);
	defparam lut_283.LUT_SIZE = 7;
	defparam lut_283.mask = 128'h77ff77ff77ff77ff7fffffffffffffff;

	lut_sub lut_290 ({sk[54], s298_out_0_, n_n852, n_n853, n_n51, x5740x, x5781x}, x5788x);
	defparam lut_290.LUT_SIZE = 7;
	defparam lut_290.mask = 128'h5555ffffffffffff55555555f7777777;

	lut_sub lut_294 ({sk[55], s298_in_2_, s298_out_0_, s298_out_4_, n_n51, n_n859, x5783x}, x5789x);
	defparam lut_294.LUT_SIZE = 7;
	defparam lut_294.mask = 128'h5555ffffffffffff5555d5d55555d5ff;

	lut_sub lut_298 ({sk[56], n_n854, n_n855, n_n856, n_n857, n_n858, n_n859}, x5527x);
	defparam lut_298.LUT_SIZE = 7;
	defparam lut_298.mask = 128'h5555ffffffffffff2020202200002022;

	lut_sub lut_302 ({sk[57], x6018x, x6294x, x6298x, x6016x, x6017x}, x6365x);
	defparam lut_302.LUT_SIZE = 6;
	defparam lut_302.mask = 64'h77ff77ff078f0f0f;

	lut_sub lut_307 ({sk[58], x6018x, x6313x, x6315x, x6016x, x6017x}, x6366x);
	defparam lut_307.LUT_SIZE = 6;
	defparam lut_307.mask = 64'h77ff77ff087f00ff;

	lut_sub lut_312 ({sk[59], x6018x, x6274x, x6282x, x6016x, x6017x, x12835x}, x12843x);
	defparam lut_312.LUT_SIZE = 7;
	defparam lut_312.mask = 128'h5555ffffffffffff7f3f3f3fffffffff;

	lut_sub lut_317 ({sk[60], x5947x, x5785x, x5786x, x5787x, x5788x, x5789x}, x536x);
	defparam lut_317.LUT_SIZE = 7;
	defparam lut_317.mask = 128'h5555ffffffffffff000000007fffffff;

	lut_sub lut_323 ({sk[61], x5967x, x5785x, x5786x, x5787x, x5788x, x5789x}, x542x);
	defparam lut_323.LUT_SIZE = 7;
	defparam lut_323.mask = 128'h5555ffffffffffff0000000080000000;

	lut_sub lut_325 ({sk[62], x5973x, x5785x, x5786x, x5787x, x5788x, x5789x}, x544x);
	defparam lut_325.LUT_SIZE = 7;
	defparam lut_325.mask = 128'h5555ffffffffffff0000000080000000;

	lut_sub lut_327 ({sk[63], x5997x, x5998x, x6003x}, x6007x);
	defparam lut_327.LUT_SIZE = 4;
	defparam lut_327.mask = 16'h3f7f;

	lut_sub lut_331 ({sk[64], x5999x, x6000x, x6001x, x6002x}, x6008x);
	defparam lut_331.LUT_SIZE = 5;
	defparam lut_331.mask = 32'h3fff7fff;

	lut_sub lut_336 ({sk[65], n_n854, n_n855, n_n856, n_n858, n_n859}, x603x);
	defparam lut_336.LUT_SIZE = 6;
	defparam lut_336.mask = 64'h00ff00ff20000000;

	lut_sub lut_338 ({sk[66], s298_in_2_, n_n852, n_n853, n_n855, n_n859}, x604x);
	defparam lut_338.LUT_SIZE = 6;
	defparam lut_338.mask = 64'h00ff00ff00080000;

	lut_sub lut_340 ({sk[67], s298_in_2_, n_n852, n_n855, n_n856, n_n857, n_n859}, x5687x);
	defparam lut_340.LUT_SIZE = 7;
	defparam lut_340.mask = 128'h33ffffffffffffff0000a00000008000;

	lut_sub lut_343 ({sk[68], x600x, x602x, x12839x}, x5696x);
	defparam lut_343.LUT_SIZE = 4;
	defparam lut_343.mask = 16'h3fbf;

	lut_sub lut_347 ({sk[69], x5672x, x5673x, x5674x, x5689x, x12838x}, x5703x);
	defparam lut_347.LUT_SIZE = 6;
	defparam lut_347.mask = 64'h00ff00ffbfffffff;

	lut_sub lut_353 ({sk[70], s298_in_0_, s298_in_2_, n_n855, n_n856, n_n857}, x8757x);
	defparam lut_353.LUT_SIZE = 6;
	defparam lut_353.mask = 64'h33ff33ff20000000;

	lut_sub lut_355 ({sk[71], s298_in_1_, n_n852, n_n853, n_n854, x8757x}, x8758x);
	defparam lut_355.LUT_SIZE = 6;
	defparam lut_355.mask = 64'h33ff33ff00040000;

	lut_sub lut_357 ({sk[72], s298_in_1_, n_n852, n_n854, n_n855}, x8763x);
	defparam lut_357.LUT_SIZE = 5;
	defparam lut_357.mask = 32'h0f0f4000;

	lut_sub lut_359 ({sk[73], s298_in_0_, s298_in_2_, n_n50, n_n857, x8763x}, x8765x);
	defparam lut_359.LUT_SIZE = 6;
	defparam lut_359.mask = 64'h33ff33ff40000000;

	lut_sub lut_361 ({sk[74], s298_in_1_, n_n852, n_n853, n_n854}, x8777x);
	defparam lut_361.LUT_SIZE = 5;
	defparam lut_361.mask = 32'h0f0f8000;

	lut_sub lut_363 ({sk[75], s298_in_0_, s298_in_2_, s298_out_5_, n_n857, n_n52, x8777x}, x27x);
	defparam lut_363.LUT_SIZE = 7;
	defparam lut_363.mask = 128'h7777ffff7777ffff0001000000000000;

	lut_sub lut_365 ({sk[76], s298_in_1_, n_n852, n_n855, n_n856}, x8784x);
	defparam lut_365.LUT_SIZE = 5;
	defparam lut_365.mask = 32'h33ff0800;

	lut_sub lut_367 ({sk[77], s298_in_0_, s298_in_2_, s298_out_3_, n_n858, x8784x}, x8786x);
	defparam lut_367.LUT_SIZE = 6;
	defparam lut_367.mask = 64'h55ffffff10000000;

	lut_sub lut_369 ({sk[78], s298_in_0_, s298_in_2_, s298_in_1_, n_n853}, x8791x);
	defparam lut_369.LUT_SIZE = 5;
	defparam lut_369.mask = 32'h33ff2000;

	lut_sub lut_371 ({sk[79], n_n855, n_n856, n_n858, n_n52, n_n859, x8791x}, x29x);
	defparam lut_371.LUT_SIZE = 7;
	defparam lut_371.mask = 128'h0fff5fffffffffff0000001000000000;

	lut_sub lut_373 ({sk[80], s298_in_0_, s298_in_2_, n_n856, n_n858, n_n859}, x8800x);
	defparam lut_373.LUT_SIZE = 6;
	defparam lut_373.mask = 64'h55ffffff00000100;

	lut_sub lut_375 ({sk[81], s298_in_1_, n_n853, n_n854, n_n855}, x8883x);
	defparam lut_375.LUT_SIZE = 5;
	defparam lut_375.mask = 32'h33ff0010;

	lut_sub lut_377 ({sk[82], s298_in_0_, s298_in_2_, s298_out_4_, n_n856, x8883x}, x44x);
	defparam lut_377.LUT_SIZE = 6;
	defparam lut_377.mask = 64'h3fff3fff04000000;

	lut_sub lut_379 ({sk[83], s298_in_2_, s298_in_1_, s298_out_1_, n_n854, n_n855, n_n50}, x8895x);
	defparam lut_379.LUT_SIZE = 7;
	defparam lut_379.mask = 128'h0fff3fff0fff3fff0000002000000000;

	lut_sub lut_381 ({sk[84], s298_in_2_, s298_out_5_, n_n853, n_n854, n_n857, n_n51}, x8900x);
	defparam lut_381.LUT_SIZE = 7;
	defparam lut_381.mask = 128'h0fff3fff0fff3fff0040000000000000;

	lut_sub lut_383 ({sk[85], s298_in_2_, s298_out_3_, s298_out_5_, n_n854, n_n855, n_n52}, x8905x);
	defparam lut_383.LUT_SIZE = 7;
	defparam lut_383.mask = 128'h0fff3fff0fff3fff1000000000000000;

	lut_sub lut_385 ({sk[86], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n51, n_n52}, x8910x);
	defparam lut_385.LUT_SIZE = 7;
	defparam lut_385.mask = 128'h0fff3fff0fff3fff0400000000000000;

	lut_sub lut_387 ({sk[87], s298_in_2_, n_n853, n_n855, n_n856, n_n52, n_n859}, x8915x);
	defparam lut_387.LUT_SIZE = 7;
	defparam lut_387.mask = 128'h0fff3fff0fff3fff0010000000000000;

	lut_sub lut_389 ({sk[88], s298_in_2_, n_n853, n_n855, n_n856, n_n52, n_n859}, x8920x);
	defparam lut_389.LUT_SIZE = 7;
	defparam lut_389.mask = 128'h0fff3fff0fff3fff0000100000000000;

	lut_sub lut_391 ({sk[89], s298_in_0_, s298_in_1_, n_n852, n_n855, n_n50, n_n857}, x8925x);
	defparam lut_391.LUT_SIZE = 7;
	defparam lut_391.mask = 128'h0fff3fff0fff3fff0000004000000000;

	lut_sub lut_393 ({sk[90], s298_in_0_, s298_in_1_, s298_out_0_, n_n852, n_n854, n_n857}, x8930x);
	defparam lut_393.LUT_SIZE = 7;
	defparam lut_393.mask = 128'h0f0fffffffffffff1000000000000000;

	lut_sub lut_395 ({sk[91], s298_in_0_, s298_in_1_, s298_out_0_, n_n852, n_n855, n_n856}, x8935x);
	defparam lut_395.LUT_SIZE = 7;
	defparam lut_395.mask = 128'h0f0fffffffffffff0000000000000080;

	lut_sub lut_397 ({sk[92], s298_in_0_, s298_in_1_, n_n853, n_n854, n_n857, n_n51}, x8940x);
	defparam lut_397.LUT_SIZE = 7;
	defparam lut_397.mask = 128'h0f0fffffffffffff0000000080000000;

	lut_sub lut_399 ({sk[93], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n857, n_n52}, x8945x);
	defparam lut_399.LUT_SIZE = 7;
	defparam lut_399.mask = 128'h0f0fffffffffffff0000000000020000;

	lut_sub lut_401 ({sk[94], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_1_, n_n853, n_n52}, x8950x);
	defparam lut_401.LUT_SIZE = 7;
	defparam lut_401.mask = 128'h0f0fffffffffffff0000000008000000;

	lut_sub lut_403 ({sk[95], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n854, n_n856}, x8955x);
	defparam lut_403.LUT_SIZE = 7;
	defparam lut_403.mask = 128'h0f0fffffffffffff0004000000000000;

	lut_sub lut_405 ({sk[96], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n855, n_n856}, x8960x);
	defparam lut_405.LUT_SIZE = 7;
	defparam lut_405.mask = 128'h0f0fffffffffffff0000000000010000;

	lut_sub lut_407 ({sk[97], s298_in_2_, n_n853, n_n854, n_n855, n_n856, n_n857}, x8965x);
	defparam lut_407.LUT_SIZE = 7;
	defparam lut_407.mask = 128'h0f0fffffffffffff0200000000000000;

	lut_sub lut_409 ({sk[98], s298_in_0_, s298_in_1_, n_n852, n_n854, n_n855, n_n859}, x8970x);
	defparam lut_409.LUT_SIZE = 7;
	defparam lut_409.mask = 128'h0f0fffffffffffff0000000000000800;

	lut_sub lut_411 ({sk[99], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n854, n_n857}, x8975x);
	defparam lut_411.LUT_SIZE = 7;
	defparam lut_411.mask = 128'h0f0fffffffffffff0000000000002000;

	lut_sub lut_413 ({sk[100], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n855, n_n858}, x8980x);
	defparam lut_413.LUT_SIZE = 7;
	defparam lut_413.mask = 128'h0f0fffffffffffff0000000004000000;

	lut_sub lut_415 ({sk[101], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n856, n_n858}, x8990x);
	defparam lut_415.LUT_SIZE = 7;
	defparam lut_415.mask = 128'h0f0fffffffffffff0000000000020000;

	lut_sub lut_417 ({sk[102], s298_in_0_, s298_in_1_, s298_out_2_, n_n852, n_n853, n_n51}, x8995x);
	defparam lut_417.LUT_SIZE = 7;
	defparam lut_417.mask = 128'h0f0fffffffffffff0004000000000000;

	lut_sub lut_419 ({sk[103], s298_in_2_, n_n853, n_n854, n_n855, n_n856, n_n857}, x9000x);
	defparam lut_419.LUT_SIZE = 7;
	defparam lut_419.mask = 128'h0f0fffffffffffff0000008000000000;

	lut_sub lut_421 ({sk[104], s298_in_2_, n_n852, n_n853, n_n854, n_n855, n_n857}, x9005x);
	defparam lut_421.LUT_SIZE = 7;
	defparam lut_421.mask = 128'h0f0fffffffffffff0000020000000000;

	lut_sub lut_423 ({sk[105], s298_in_0_, s298_in_2_, n_n859}, x9009x);
	defparam lut_423.LUT_SIZE = 4;
	defparam lut_423.mask = 16'h3f80;

	lut_sub lut_425 ({sk[106], s298_in_2_, s298_out_4_, n_n852, n_n856, n_n50}, x9014x);
	defparam lut_425.LUT_SIZE = 6;
	defparam lut_425.mask = 64'h5f5fffff00200000;

	lut_sub lut_427 ({sk[107], s298_in_2_, s298_out_4_, n_n853, n_n855, n_n857}, x9018x);
	defparam lut_427.LUT_SIZE = 6;
	defparam lut_427.mask = 64'h5f5fffff00020000;

	lut_sub lut_429 ({sk[108], s298_in_2_, n_n852, n_n854, n_n856, n_n52}, x9022x);
	defparam lut_429.LUT_SIZE = 6;
	defparam lut_429.mask = 64'h5f5fffff00040000;

	lut_sub lut_431 ({sk[109], s298_in_0_, n_n854, n_n856, n_n50, n_n858}, x9026x);
	defparam lut_431.LUT_SIZE = 6;
	defparam lut_431.mask = 64'h33ff33ff00002000;

	lut_sub lut_433 ({sk[110], s298_in_0_, s298_in_1_, n_n853, n_n856, n_n50}, x9030x);
	defparam lut_433.LUT_SIZE = 6;
	defparam lut_433.mask = 64'h33ff33ff00100000;

	lut_sub lut_435 ({sk[111], s298_out_4_, n_n853, n_n854, n_n856, n_n52}, x9034x);
	defparam lut_435.LUT_SIZE = 6;
	defparam lut_435.mask = 64'h33ff33ff01000000;

	lut_sub lut_437 ({sk[112], s298_in_0_, s298_out_1_, s298_out_5_, n_n853, n_n52}, x9038x);
	defparam lut_437.LUT_SIZE = 6;
	defparam lut_437.mask = 64'h33ff33ff00020000;

	lut_sub lut_439 ({sk[113], s298_in_1_, s298_out_5_, n_n855, n_n52, n_n859}, x9042x);
	defparam lut_439.LUT_SIZE = 6;
	defparam lut_439.mask = 64'h33ff33ff02000000;

	lut_sub lut_441 ({sk[114], n_n855, n_n856, n_n858, n_n52, n_n859}, x9046x);
	defparam lut_441.LUT_SIZE = 6;
	defparam lut_441.mask = 64'h33ff33ff00000020;

	lut_sub lut_443 ({sk[115], n_n852, n_n854, n_n856, n_n858, n_n52}, x9050x);
	defparam lut_443.LUT_SIZE = 6;
	defparam lut_443.mask = 64'h33ff33ff00000100;

	lut_sub lut_445 ({sk[116], s298_in_2_, s298_out_2_, n_n853, n_n855, n_n856, n_n857}, x81x);
	defparam lut_445.LUT_SIZE = 7;
	defparam lut_445.mask = 128'h1fff1fffffffffff0004000000000000;

	lut_sub lut_447 ({sk[117], x510x, x511x, x513x, x518x}, x6016x);
	defparam lut_447.LUT_SIZE = 5;
	defparam lut_447.mask = 32'h33337fff;

	lut_sub lut_452 ({sk[118], s298_out_1_, n_n852, n_n854, x6018x, x6016x, x6017x}, x9061x);
	defparam lut_452.LUT_SIZE = 7;
	defparam lut_452.mask = 128'h1fff1fffffffffff000000000000007f;

	lut_sub lut_456 ({sk[119], s298_out_0_, n_n852, n_n856, n_n858}, x9067x);
	defparam lut_456.LUT_SIZE = 5;
	defparam lut_456.mask = 32'h33330100;

	lut_sub lut_458 ({sk[120], s298_in_1_, s298_out_0_, n_n854, n_n858}, x9076x);
	defparam lut_458.LUT_SIZE = 5;
	defparam lut_458.mask = 32'h33332000;

	lut_sub lut_460 ({sk[121], s298_out_0_, n_n853, n_n854, n_n856}, x9082x);
	defparam lut_460.LUT_SIZE = 5;
	defparam lut_460.mask = 32'h5f5f0008;

	lut_sub lut_462 ({sk[122], n_n51, n_n859, x6018x, x6016x, x6017x}, x9090x);
	defparam lut_462.LUT_SIZE = 6;
	defparam lut_462.mask = 64'h000077ff7f000000;

	lut_sub lut_466 ({sk[123], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x8012x);
	defparam lut_466.LUT_SIZE = 5;
	defparam lut_466.mask = 32'h5f5f8000;

	lut_sub lut_468 ({sk[124], s298_out_4_, n_n853, n_n854, n_n855, n_n857, x8012x}, x8015x);
	defparam lut_468.LUT_SIZE = 7;
	defparam lut_468.mask = 128'h0fffffff0fffffff4000000000000000;

	lut_sub lut_470 ({sk[125], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n854}, x8020x);
	defparam lut_470.LUT_SIZE = 7;
	defparam lut_470.mask = 128'h0fffffff0fffffff0000000008000000;

	lut_sub lut_472 ({sk[126], s298_out_5_, x6018x, x6016x, x6017x, x8020x}, x8022x);
	defparam lut_472.LUT_SIZE = 6;
	defparam lut_472.mask = 64'h000077ff00004000;

	lut_sub lut_474 ({sk[127], s298_in_1_, n_n852, n_n853, n_n854}, x8041x);
	defparam lut_474.LUT_SIZE = 5;
	defparam lut_474.mask = 32'h5f5f0100;

	lut_sub lut_476 ({sk[128], s298_in_0_, s298_in_2_, n_n51, n_n858, x8041x}, x8043x);
	defparam lut_476.LUT_SIZE = 6;
	defparam lut_476.mask = 64'h0f0f3f3f00004000;

	lut_sub lut_478 ({sk[129], s298_in_2_, s298_in_1_, n_n852, n_n853}, x8054x);
	defparam lut_478.LUT_SIZE = 5;
	defparam lut_478.mask = 32'h55ff8000;

	lut_sub lut_480 ({sk[130], s298_out_1_, s298_out_3_, n_n854, n_n855, n_n50, x8054x}, x101x);
	defparam lut_480.LUT_SIZE = 7;
	defparam lut_480.mask = 128'h3333ffffffffffff0004000000000000;

	lut_sub lut_482 ({sk[131], s298_in_1_, n_n852, n_n853, n_n855}, x8076x);
	defparam lut_482.LUT_SIZE = 5;
	defparam lut_482.mask = 32'h55ff8000;

	lut_sub lut_484 ({sk[132], s298_in_0_, s298_in_2_, s298_out_0_, n_n858, n_n52, x8076x}, x104x);
	defparam lut_484.LUT_SIZE = 7;
	defparam lut_484.mask = 128'h3333ffffffffffff0100000000000000;

	lut_sub lut_486 ({sk[133], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x8090x);
	defparam lut_486.LUT_SIZE = 5;
	defparam lut_486.mask = 32'h5f5f2000;

	lut_sub lut_488 ({sk[134], s298_out_0_, n_n853, n_n854, n_n856, n_n858, x8090x}, x106x);
	defparam lut_488.LUT_SIZE = 7;
	defparam lut_488.mask = 128'h5555ffffffffffff0000000000040000;

	lut_sub lut_490 ({sk[135], s298_in_0_, s298_in_2_, s298_in_1_, n_n853}, x8097x);
	defparam lut_490.LUT_SIZE = 5;
	defparam lut_490.mask = 32'h5f5f0020;

	lut_sub lut_492 ({sk[136], n_n854, n_n855, n_n858, n_n52, n_n859, x8097x}, x107x);
	defparam lut_492.LUT_SIZE = 7;
	defparam lut_492.mask = 128'h5555ffffffffffff0000000000100000;

	lut_sub lut_494 ({sk[137], s298_in_2_, s298_in_1_, n_n852, n_n853}, x8104x);
	defparam lut_494.LUT_SIZE = 5;
	defparam lut_494.mask = 32'h5f5f8000;

	lut_sub lut_496 ({sk[138], n_n854, n_n855, n_n857, n_n858, n_n52, x8104x}, x108x);
	defparam lut_496.LUT_SIZE = 7;
	defparam lut_496.mask = 128'h5555ffffffffffff0000000400000000;

	lut_sub lut_498 ({sk[139], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x8111x);
	defparam lut_498.LUT_SIZE = 5;
	defparam lut_498.mask = 32'h5f5f4000;

	lut_sub lut_500 ({sk[140], n_n853, n_n854, n_n856, n_n857, x8111x}, x8113x);
	defparam lut_500.LUT_SIZE = 6;
	defparam lut_500.mask = 64'h5fff5fff40000000;

	lut_sub lut_502 ({sk[141], n_n852, n_n853, n_n854, n_n856}, x8118x);
	defparam lut_502.LUT_SIZE = 5;
	defparam lut_502.mask = 32'h5f5f0020;

	lut_sub lut_504 ({sk[142], s298_in_2_, s298_in_1_, s298_out_2_, n_n857, n_n52, x8118x}, x110x);
	defparam lut_504.LUT_SIZE = 7;
	defparam lut_504.mask = 128'h5555ffffffffffff0000010000000000;

	lut_sub lut_506 ({sk[143], s298_in_0_, s298_in_2_, n_n856, n_n857, n_n859}, x8127x);
	defparam lut_506.LUT_SIZE = 6;
	defparam lut_506.mask = 64'h5fff5fff00001000;

	lut_sub lut_508 ({sk[144], s298_in_0_, s298_in_2_, n_n855, n_n856, n_n859}, x8134x);
	defparam lut_508.LUT_SIZE = 6;
	defparam lut_508.mask = 64'h5fff5fff00004000;

	lut_sub lut_510 ({sk[145], s298_in_0_, s298_in_2_, n_n855, n_n857, n_n859}, x8141x);
	defparam lut_510.LUT_SIZE = 6;
	defparam lut_510.mask = 64'h5fff5fff04000000;

	lut_sub lut_512 ({sk[146], s298_in_0_, s298_in_2_, n_n855, n_n858, n_n859}, x8148x);
	defparam lut_512.LUT_SIZE = 6;
	defparam lut_512.mask = 64'h5fff5fff10000000;

	lut_sub lut_514 ({sk[147], s298_in_0_, s298_in_2_, n_n855, n_n856, n_n858}, x8155x);
	defparam lut_514.LUT_SIZE = 6;
	defparam lut_514.mask = 64'h5fff5fff10000000;

	lut_sub lut_516 ({sk[148], s298_in_0_, s298_in_2_, n_n855, n_n856, n_n858}, x8162x);
	defparam lut_516.LUT_SIZE = 6;
	defparam lut_516.mask = 64'h5fff5fff08000000;

	lut_sub lut_518 ({sk[149], s298_in_0_, s298_in_2_, n_n855, n_n856, n_n857}, x8169x);
	defparam lut_518.LUT_SIZE = 6;
	defparam lut_518.mask = 64'h5fff5fff00000100;

	lut_sub lut_520 ({sk[150], s298_in_1_, n_n853, n_n854, n_n855}, x8175x);
	defparam lut_520.LUT_SIZE = 5;
	defparam lut_520.mask = 32'h5f5f0020;

	lut_sub lut_522 ({sk[151], s298_in_0_, s298_in_2_, n_n856, n_n857, n_n858}, x8176x);
	defparam lut_522.LUT_SIZE = 6;
	defparam lut_522.mask = 64'h5555777702000000;

	lut_sub lut_524 ({sk[152], s298_in_1_, n_n853, n_n854, n_n858}, x8265x);
	defparam lut_524.LUT_SIZE = 5;
	defparam lut_524.mask = 32'h0f5f0400;

	lut_sub lut_526 ({sk[153], s298_in_0_, s298_in_2_, s298_out_1_, n_n859, x8265x}, x133x);
	defparam lut_526.LUT_SIZE = 6;
	defparam lut_526.mask = 64'h5555777740000000;

	lut_sub lut_528 ({sk[154], s298_in_1_, s298_out_3_, n_n853, n_n854, n_n857, n_n859}, x8301x);
	defparam lut_528.LUT_SIZE = 7;
	defparam lut_528.mask = 128'h77ff7fff77ff7fff0200000000000000;

	lut_sub lut_530 ({sk[155], s298_out_0_, n_n52, x8301x}, x139x);
	defparam lut_530.LUT_SIZE = 4;
	defparam lut_530.mask = 16'h3310;

	lut_sub lut_532 ({sk[156], s298_in_1_, n_n852, n_n853, n_n854}, x8313x);
	defparam lut_532.LUT_SIZE = 5;
	defparam lut_532.mask = 32'h0f5f0080;

	lut_sub lut_534 ({sk[157], s298_in_0_, s298_in_2_, s298_out_4_, n_n856, x8313x}, x141x);
	defparam lut_534.LUT_SIZE = 6;
	defparam lut_534.mask = 64'h5555777704000000;

	lut_sub lut_536 ({sk[158], n_n852, n_n853, n_n854, n_n855}, x8367x);
	defparam lut_536.LUT_SIZE = 5;
	defparam lut_536.mask = 32'h0f5f0001;

	lut_sub lut_538 ({sk[159], s298_in_0_, s298_in_1_, s298_out_5_, n_n858, x8367x}, x150x);
	defparam lut_538.LUT_SIZE = 6;
	defparam lut_538.mask = 64'h5555777700004000;

	lut_sub lut_540 ({sk[160], n_n852, n_n853, n_n855, n_n856}, x8397x);
	defparam lut_540.LUT_SIZE = 5;
	defparam lut_540.mask = 32'h0f5f4000;

	lut_sub lut_542 ({sk[161], s298_in_2_, s298_in_1_, n_n857, n_n52, x8397x}, x155x);
	defparam lut_542.LUT_SIZE = 6;
	defparam lut_542.mask = 64'h5555777700010000;

	lut_sub lut_544 ({sk[162], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x8409x);
	defparam lut_544.LUT_SIZE = 5;
	defparam lut_544.mask = 32'h0f5f0040;

	lut_sub lut_546 ({sk[163], n_n853, n_n855, n_n856, n_n859}, x8410x);
	defparam lut_546.LUT_SIZE = 5;
	defparam lut_546.mask = 32'h0f5f0400;

	lut_sub lut_548 ({sk[164], s298_in_0_, s298_in_2_, n_n852, n_n853}, x8415x);
	defparam lut_548.LUT_SIZE = 5;
	defparam lut_548.mask = 32'h0f5f4000;

	lut_sub lut_550 ({sk[165], n_n854, n_n855, n_n857, n_n858}, x8416x);
	defparam lut_550.LUT_SIZE = 5;
	defparam lut_550.mask = 32'h0f5f2000;

	lut_sub lut_552 ({sk[166], n_n853, n_n854, n_n855, n_n858}, x8422x);
	defparam lut_552.LUT_SIZE = 5;
	defparam lut_552.mask = 32'h0f5f0080;

	lut_sub lut_554 ({sk[167], n_n854, n_n855, n_n856, n_n857}, x8428x);
	defparam lut_554.LUT_SIZE = 5;
	defparam lut_554.mask = 32'h0f5f0010;

	lut_sub lut_556 ({sk[168], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x8433x);
	defparam lut_556.LUT_SIZE = 5;
	defparam lut_556.mask = 32'h0f5f0040;

	lut_sub lut_558 ({sk[169], n_n853, n_n854, n_n856, n_n858, x8433x}, x161x);
	defparam lut_558.LUT_SIZE = 6;
	defparam lut_558.mask = 64'h5555777700010000;

	lut_sub lut_560 ({sk[170], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_1_, n_n853, n_n854}, x8439x);
	defparam lut_560.LUT_SIZE = 7;
	defparam lut_560.mask = 128'h77ff7fff77ff7fff0000000002000000;

	lut_sub lut_562 ({sk[171], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_1_, n_n852, n_n856}, x8444x);
	defparam lut_562.LUT_SIZE = 7;
	defparam lut_562.mask = 128'h77ff7fff77ff7fff0002000000000000;

	lut_sub lut_564 ({sk[172], s298_in_2_, s298_in_1_, s298_out_4_, n_n854, n_n856, n_n50}, x8449x);
	defparam lut_564.LUT_SIZE = 7;
	defparam lut_564.mask = 128'h77ff7fff77ff7fff0000000200000000;

	lut_sub lut_566 ({sk[173], s298_in_1_, s298_out_3_, n_n853, n_n856, n_n50, n_n52}, x8454x);
	defparam lut_566.LUT_SIZE = 7;
	defparam lut_566.mask = 128'h77ff7fff77ff7fff0000000010000000;

	lut_sub lut_568 ({sk[174], s298_in_0_, s298_out_0_, n_n853, n_n854, n_n855, n_n858}, x8459x);
	defparam lut_568.LUT_SIZE = 7;
	defparam lut_568.mask = 128'h77ff7fff77ff7fff0000000008000000;

	lut_sub lut_570 ({sk[175], s298_in_0_, n_n852, n_n854, n_n856, n_n52, n_n859}, x8464x);
	defparam lut_570.LUT_SIZE = 7;
	defparam lut_570.mask = 128'h77ff7fff77ff7fff0000000000000200;

	lut_sub lut_572 ({sk[176], s298_out_1_, n_n852, n_n853, n_n854, n_n855, n_n856}, x8469x);
	defparam lut_572.LUT_SIZE = 7;
	defparam lut_572.mask = 128'h77ff7fff77ff7fff0000010000000000;

	lut_sub lut_574 ({sk[177], s298_in_0_, s298_in_1_, s298_out_0_, n_n852, n_n854, n_n50}, x8474x);
	defparam lut_574.LUT_SIZE = 7;
	defparam lut_574.mask = 128'h77ff7fff77ff7fff0000008000000000;

	lut_sub lut_576 ({sk[178], s298_in_0_, s298_out_0_, n_n852, n_n854, n_n50, n_n858}, x8479x);
	defparam lut_576.LUT_SIZE = 7;
	defparam lut_576.mask = 128'h77ff7fff77ff7fff0000000000000800;

	lut_sub lut_578 ({sk[179], s298_in_0_, n_n852, n_n855, n_n856, n_n50, n_n857}, x8484x);
	defparam lut_578.LUT_SIZE = 7;
	defparam lut_578.mask = 128'h77ff7fff77ff7fff0000000800000000;

	lut_sub lut_580 ({sk[180], s298_in_0_, s298_in_1_, n_n852, n_n50, n_n857, n_n51}, x8489x);
	defparam lut_580.LUT_SIZE = 7;
	defparam lut_580.mask = 128'h77ff7fff77ff7fff0000000000020000;

	lut_sub lut_582 ({sk[181], s298_in_0_, s298_in_1_, n_n853, n_n854, n_n856, n_n50}, x8494x);
	defparam lut_582.LUT_SIZE = 7;
	defparam lut_582.mask = 128'h77ff7fff77ff7fff0000000010000000;

	lut_sub lut_584 ({sk[182], s298_in_0_, s298_in_1_, s298_out_0_, n_n852, n_n855, n_n857}, x8499x);
	defparam lut_584.LUT_SIZE = 7;
	defparam lut_584.mask = 128'h77ff7fff77ff7fff0010000000000000;

	lut_sub lut_586 ({sk[183], s298_in_0_, s298_in_1_, s298_out_0_, n_n853, n_n855, n_n858}, x8504x);
	defparam lut_586.LUT_SIZE = 7;
	defparam lut_586.mask = 128'h77ff7fff77ff7fff0000000000000080;

	lut_sub lut_588 ({sk[184], s298_in_0_, s298_in_1_, s298_out_4_, n_n852, n_n853, n_n854}, x8509x);
	defparam lut_588.LUT_SIZE = 7;
	defparam lut_588.mask = 128'h77ff7fff77ff7fff0000000000200000;

	lut_sub lut_590 ({sk[185], s298_in_0_, s298_in_1_, s298_out_5_, n_n853, n_n854, n_n858}, x8514x);
	defparam lut_590.LUT_SIZE = 7;
	defparam lut_590.mask = 128'h77ff7fff77ff7fff2000000000000000;

	lut_sub lut_592 ({sk[186], s298_in_0_, s298_in_1_, n_n853, n_n854, n_n856, n_n857}, x8519x);
	defparam lut_592.LUT_SIZE = 7;
	defparam lut_592.mask = 128'h77ff7fff77ff7fff0000001000000000;

	lut_sub lut_594 ({sk[187], s298_in_2_, s298_in_1_, s298_out_4_, n_n854, n_n855, n_n52}, x8524x);
	defparam lut_594.LUT_SIZE = 7;
	defparam lut_594.mask = 128'h77ff7fff77ff7fff0000004000000000;

	lut_sub lut_596 ({sk[188], s298_in_2_, s298_in_1_, s298_out_4_, n_n853, n_n854, n_n855}, x8529x);
	defparam lut_596.LUT_SIZE = 7;
	defparam lut_596.mask = 128'h77ff7fff77ff7fff0000000100000000;

	lut_sub lut_598 ({sk[189], s298_in_0_, s298_in_1_, s298_out_4_, n_n852, n_n853, n_n859}, x8534x);
	defparam lut_598.LUT_SIZE = 7;
	defparam lut_598.mask = 128'h77ff7fff77ff7fff0000000000000040;

	lut_sub lut_600 ({sk[190], s298_in_0_, s298_in_1_, s298_out_5_, n_n852, n_n853, n_n858}, x8539x);
	defparam lut_600.LUT_SIZE = 7;
	defparam lut_600.mask = 128'h77ff7fff77ff7fff0000000000000200;

	lut_sub lut_602 ({sk[191], s298_in_0_, s298_in_1_, n_n853, n_n854, n_n856, n_n858}, x8544x);
	defparam lut_602.LUT_SIZE = 7;
	defparam lut_602.mask = 128'h77ff7fff77ff7fff0000000200000000;

	lut_sub lut_604 ({sk[192], s298_in_0_, n_n852, n_n854, n_n855, n_n856, n_n858}, x8549x);
	defparam lut_604.LUT_SIZE = 7;
	defparam lut_604.mask = 128'h77ff7fff77ff7fff0000000008000000;

	lut_sub lut_606 ({sk[193], s298_in_0_, n_n852, n_n853, n_n854, n_n855, n_n858}, x8554x);
	defparam lut_606.LUT_SIZE = 7;
	defparam lut_606.mask = 128'h77ff7fff77ff7fff0002000000000000;

	lut_sub lut_608 ({sk[194], s298_in_0_, s298_in_2_, n_n852, n_n853, n_n854, n_n855}, x8559x);
	defparam lut_608.LUT_SIZE = 7;
	defparam lut_608.mask = 128'h77ff7fff77ff7fff0000000004000000;

	lut_sub lut_610 ({sk[195], s298_in_2_, s298_in_1_, n_n852, n_n854, n_n855, n_n857}, x8564x);
	defparam lut_610.LUT_SIZE = 7;
	defparam lut_610.mask = 128'h77ff7fff77ff7fff0000001000000000;

	lut_sub lut_612 ({sk[196], s298_in_0_, s298_in_1_, n_n853, n_n854, n_n855, n_n857}, x8569x);
	defparam lut_612.LUT_SIZE = 7;
	defparam lut_612.mask = 128'h77ff7fff77ff7fff0000800000000000;

	lut_sub lut_614 ({sk[197], s298_in_1_, s298_out_1_, n_n853, n_n856, n_n50}, x8573x);
	defparam lut_614.LUT_SIZE = 6;
	defparam lut_614.mask = 64'h5555777700020000;

	lut_sub lut_616 ({sk[198], s298_in_0_, s298_in_1_, s298_out_1_, n_n855, n_n51}, x8577x);
	defparam lut_616.LUT_SIZE = 6;
	defparam lut_616.mask = 64'h5555777700000004;

	lut_sub lut_618 ({sk[199], s298_in_2_, n_n854, n_n50, n_n857, n_n51}, x8581x);
	defparam lut_618.LUT_SIZE = 6;
	defparam lut_618.mask = 64'h5555777700040000;

	lut_sub lut_620 ({sk[200], s298_in_1_, n_n854, n_n855, n_n50, n_n857}, x8585x);
	defparam lut_620.LUT_SIZE = 6;
	defparam lut_620.mask = 64'h5555777700200000;

	lut_sub lut_622 ({sk[201], s298_out_1_, n_n852, n_n51, n_n858, n_n859}, x8589x);
	defparam lut_622.LUT_SIZE = 6;
	defparam lut_622.mask = 64'h5555777702000000;

	lut_sub lut_624 ({sk[202], s298_out_4_, n_n852, n_n855, n_n856, n_n52}, x8593x);
	defparam lut_624.LUT_SIZE = 6;
	defparam lut_624.mask = 64'h5555777700000002;

	lut_sub lut_626 ({sk[203], s298_in_1_, n_n853, n_n854, n_n855, n_n52}, x8597x);
	defparam lut_626.LUT_SIZE = 6;
	defparam lut_626.mask = 64'h5555777702000000;

	lut_sub lut_628 ({sk[204], s298_in_0_, n_n853, n_n856, n_n857, n_n52}, x8601x);
	defparam lut_628.LUT_SIZE = 6;
	defparam lut_628.mask = 64'h5555777700020000;

	lut_sub lut_630 ({sk[205], s298_in_0_, s298_in_1_, n_n852, n_n854, n_n859}, x8605x);
	defparam lut_630.LUT_SIZE = 6;
	defparam lut_630.mask = 64'h5555777700008000;

	lut_sub lut_632 ({sk[206], s298_in_1_, n_n852, n_n854, n_n855, n_n857}, x8609x);
	defparam lut_632.LUT_SIZE = 6;
	defparam lut_632.mask = 64'h5555777700400000;

	lut_sub lut_634 ({sk[207], s298_in_1_, s298_out_0_, n_n852, n_n855, n_n856, n_n858}, x199x);
	defparam lut_634.LUT_SIZE = 7;
	defparam lut_634.mask = 128'h77ff7fff77ff7fff0020000000000000;

	lut_sub lut_636 ({sk[208], s298_in_0_, s298_in_2_, n_n852, n_n853, n_n858}, x8617x);
	defparam lut_636.LUT_SIZE = 6;
	defparam lut_636.mask = 64'h5555777700004000;

	lut_sub lut_638 ({sk[209], s298_in_1_, n_n853, n_n855, n_n856, n_n858}, x8621x);
	defparam lut_638.LUT_SIZE = 6;
	defparam lut_638.mask = 64'h5555777700000002;

	lut_sub lut_640 ({sk[210], s298_in_0_, s298_in_2_, n_n855}, x8624x);
	defparam lut_640.LUT_SIZE = 4;
	defparam lut_640.mask = 16'h3308;

	lut_sub lut_642 ({sk[211], s298_in_2_, s298_out_0_, n_n853, n_n859}, x8631x);
	defparam lut_642.LUT_SIZE = 5;
	defparam lut_642.mask = 32'h0f5f0800;

	lut_sub lut_644 ({sk[212], s298_in_2_, s298_out_1_, s298_out_4_, n_n854}, x205x);
	defparam lut_644.LUT_SIZE = 5;
	defparam lut_644.mask = 32'h0f5f0001;

	lut_sub lut_646 ({sk[213], n_n855, n_n857, n_n859}, x8637x);
	defparam lut_646.LUT_SIZE = 4;
	defparam lut_646.mask = 16'h3340;

	lut_sub lut_648 ({sk[214], s298_in_0_, s298_in_2_, n_n855, n_n857, n_n858}, x7242x);
	defparam lut_648.LUT_SIZE = 6;
	defparam lut_648.mask = 64'h5555777700008000;

	lut_sub lut_650 ({sk[215], s298_in_1_, s298_out_5_, n_n852, n_n853, n_n854, x7242x}, x209x);
	defparam lut_650.LUT_SIZE = 7;
	defparam lut_650.mask = 128'h77ff7fff77ff7fff0100000000000000;

	lut_sub lut_652 ({sk[216], s298_in_1_, n_n852, n_n855, n_n857}, x7255x);
	defparam lut_652.LUT_SIZE = 5;
	defparam lut_652.mask = 32'h0f5f0001;

	lut_sub lut_654 ({sk[217], s298_in_0_, s298_in_2_, s298_out_4_, n_n859, x7255x}, x7257x);
	defparam lut_654.LUT_SIZE = 6;
	defparam lut_654.mask = 64'h5555777700000100;

	lut_sub lut_656 ({sk[218], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7276x);
	defparam lut_656.LUT_SIZE = 5;
	defparam lut_656.mask = 32'h0f5f2000;

	lut_sub lut_658 ({sk[219], s298_out_1_, n_n853, n_n854, n_n856, n_n858, x7276x}, x214x);
	defparam lut_658.LUT_SIZE = 7;
	defparam lut_658.mask = 128'h77ff7fff77ff7fff0100000000000000;

	lut_sub lut_660 ({sk[220], s298_in_1_, n_n852, n_n853, n_n854}, x7283x);
	defparam lut_660.LUT_SIZE = 5;
	defparam lut_660.mask = 32'h0f5f2000;

	lut_sub lut_662 ({sk[221], s298_in_0_, s298_in_2_, n_n50, n_n857, n_n51, x7283x}, x215x);
	defparam lut_662.LUT_SIZE = 7;
	defparam lut_662.mask = 128'h77ff7fff77ff7fff0001000000000000;

	lut_sub lut_664 ({sk[222], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7304x);
	defparam lut_664.LUT_SIZE = 5;
	defparam lut_664.mask = 32'h0f5f2000;

	lut_sub lut_666 ({sk[223], s298_out_0_, n_n854, n_n855, n_n856, n_n857, x7304x}, x218x);
	defparam lut_666.LUT_SIZE = 7;
	defparam lut_666.mask = 128'h77ff7fff77ff7fff0000400000000000;

	lut_sub lut_668 ({sk[224], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7311x);
	defparam lut_668.LUT_SIZE = 5;
	defparam lut_668.mask = 32'h0f5f2000;

	lut_sub lut_670 ({sk[225], s298_out_0_, n_n853, n_n854, n_n855, n_n858, x7311x}, x219x);
	defparam lut_670.LUT_SIZE = 7;
	defparam lut_670.mask = 128'h77ff7fff77ff7fff0000000000000040;

	lut_sub lut_672 ({sk[226], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7318x);
	defparam lut_672.LUT_SIZE = 5;
	defparam lut_672.mask = 32'h0f5f1000;

	lut_sub lut_674 ({sk[227], s298_out_0_, n_n853, n_n854, n_n855, n_n857, x7318x}, x220x);
	defparam lut_674.LUT_SIZE = 7;
	defparam lut_674.mask = 128'h77ff7fff77ff7fff0000000000000004;

	lut_sub lut_676 ({sk[228], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7325x);
	defparam lut_676.LUT_SIZE = 5;
	defparam lut_676.mask = 32'h0f5f8000;

	lut_sub lut_678 ({sk[229], n_n853, n_n855, n_n857, n_n858, x7325x}, x7327x);
	defparam lut_678.LUT_SIZE = 6;
	defparam lut_678.mask = 64'h5555777704000000;

	lut_sub lut_680 ({sk[230], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7332x);
	defparam lut_680.LUT_SIZE = 5;
	defparam lut_680.mask = 32'h0f5f0020;

	lut_sub lut_682 ({sk[231], s298_out_4_, n_n853, n_n854, n_n855, n_n857, x7332x}, x222x);
	defparam lut_682.LUT_SIZE = 7;
	defparam lut_682.mask = 128'h77ff7fff77ff7fff0000001000000000;

	lut_sub lut_684 ({sk[232], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7339x);
	defparam lut_684.LUT_SIZE = 5;
	defparam lut_684.mask = 32'h0f5f8000;

	lut_sub lut_686 ({sk[233], s298_out_4_, n_n853, n_n855, n_n856, n_n857, x7339x}, x223x);
	defparam lut_686.LUT_SIZE = 7;
	defparam lut_686.mask = 128'h77ff7fff77ff7fff0000040000000000;

	lut_sub lut_688 ({sk[234], s298_in_1_, n_n852, n_n854, n_n855}, x7346x);
	defparam lut_688.LUT_SIZE = 5;
	defparam lut_688.mask = 32'h0f5f0400;

	lut_sub lut_690 ({sk[235], s298_in_0_, s298_in_2_, s298_out_4_, n_n856, n_n52, x7346x}, x224x);
	defparam lut_690.LUT_SIZE = 7;
	defparam lut_690.mask = 128'h77ff7fff77ff7fff0000000000400000;

	lut_sub lut_692 ({sk[236], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7353x);
	defparam lut_692.LUT_SIZE = 5;
	defparam lut_692.mask = 32'h0f5f2000;

	lut_sub lut_694 ({sk[237], n_n853, n_n854, n_n855, n_n856, x7353x}, x7355x);
	defparam lut_694.LUT_SIZE = 6;
	defparam lut_694.mask = 64'h5555777700000004;

	lut_sub lut_696 ({sk[238], s298_in_2_, s298_in_1_, n_n852, n_n853}, x7360x);
	defparam lut_696.LUT_SIZE = 5;
	defparam lut_696.mask = 32'h0f5f8000;

	lut_sub lut_698 ({sk[239], n_n854, n_n855, n_n858, n_n52, n_n859, x7360x}, x226x);
	defparam lut_698.LUT_SIZE = 7;
	defparam lut_698.mask = 128'h77ff7fff77ff7fff0000000000100000;

	lut_sub lut_700 ({sk[240], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7367x);
	defparam lut_700.LUT_SIZE = 5;
	defparam lut_700.mask = 32'h0f5f0020;

	lut_sub lut_702 ({sk[241], n_n853, n_n855, n_n856, n_n859, x7367x}, x7369x);
	defparam lut_702.LUT_SIZE = 6;
	defparam lut_702.mask = 64'h5555777710000000;

	lut_sub lut_704 ({sk[242], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7374x);
	defparam lut_704.LUT_SIZE = 5;
	defparam lut_704.mask = 32'h0f5f2000;

	lut_sub lut_706 ({sk[243], n_n853, n_n854, n_n855, n_n857, n_n52, x7374x}, x228x);
	defparam lut_706.LUT_SIZE = 7;
	defparam lut_706.mask = 128'h77ff7fff77ff7fff1000000000000000;

	lut_sub lut_708 ({sk[244], s298_in_0_, s298_in_2_, s298_in_1_, n_n853}, x7381x);
	defparam lut_708.LUT_SIZE = 5;
	defparam lut_708.mask = 32'h0f5f8000;

	lut_sub lut_710 ({sk[245], n_n854, n_n855, n_n856, n_n857, n_n52, x7381x}, x229x);
	defparam lut_710.LUT_SIZE = 7;
	defparam lut_710.mask = 128'h77ff7fff77ff7fff0000001000000000;

	lut_sub lut_712 ({sk[246], n_n853, n_n854, n_n856, n_n858}, x7389x);
	defparam lut_712.LUT_SIZE = 5;
	defparam lut_712.mask = 32'h0f5f0040;

	lut_sub lut_714 ({sk[247], s298_in_1_, n_n852, n_n853, n_n854}, x7396x);
	defparam lut_714.LUT_SIZE = 5;
	defparam lut_714.mask = 32'h0f5f0002;

	lut_sub lut_716 ({sk[248], s298_in_0_, s298_in_2_, n_n857, n_n858, n_n859}, x7397x);
	defparam lut_716.LUT_SIZE = 6;
	defparam lut_716.mask = 64'h5555777701000000;

	lut_sub lut_718 ({sk[249], s298_in_0_, s298_in_2_, n_n856, n_n857, n_n859}, x7404x);
	defparam lut_718.LUT_SIZE = 6;
	defparam lut_718.mask = 64'h5555777740000000;

	lut_sub lut_720 ({sk[250], s298_in_0_, s298_in_2_, n_n856, n_n857, n_n858}, x7411x);
	defparam lut_720.LUT_SIZE = 6;
	defparam lut_720.mask = 64'h5555777700000100;

	lut_sub lut_722 ({sk[251], s298_in_1_, n_n852, n_n853, n_n854, x7411x}, x233x);
	defparam lut_722.LUT_SIZE = 6;
	defparam lut_722.mask = 64'h5555777700000040;

	lut_sub lut_724 ({sk[252], s298_in_0_, s298_in_2_, n_n856, n_n857, n_n858}, x7418x);
	defparam lut_724.LUT_SIZE = 6;
	defparam lut_724.mask = 64'h5555777708000000;

	lut_sub lut_726 ({sk[253], s298_in_1_, n_n852, n_n853, n_n854}, x7549x);
	defparam lut_726.LUT_SIZE = 5;
	defparam lut_726.mask = 32'h0f5f0008;

	lut_sub lut_728 ({sk[254], s298_in_0_, s298_in_2_, n_n857, x7549x}, x7550x);
	defparam lut_728.LUT_SIZE = 5;
	defparam lut_728.mask = 32'h0f5f1000;

	lut_sub lut_730 ({sk[255], s298_in_1_, n_n853, n_n855, n_n856}, x7555x);
	defparam lut_730.LUT_SIZE = 5;
	defparam lut_730.mask = 32'h0f5f4000;

	lut_sub lut_732 ({sk[256], s298_in_0_, s298_in_2_, s298_out_0_, n_n858, x7555x}, x257x);
	defparam lut_732.LUT_SIZE = 6;
	defparam lut_732.mask = 64'h5555777700004000;

	lut_sub lut_734 ({sk[257], s298_in_1_, n_n852, n_n853, n_n854}, x7567x);
	defparam lut_734.LUT_SIZE = 5;
	defparam lut_734.mask = 32'h0f5f0800;

	lut_sub lut_736 ({sk[258], s298_in_0_, s298_in_2_, s298_out_0_, n_n856, x7567x}, x259x);
	defparam lut_736.LUT_SIZE = 6;
	defparam lut_736.mask = 64'h5555777700000400;

	lut_sub lut_738 ({sk[259], s298_in_1_, n_n852, n_n853, n_n855}, x7591x);
	defparam lut_738.LUT_SIZE = 5;
	defparam lut_738.mask = 32'h0f5f0100;

	lut_sub lut_740 ({sk[260], s298_in_0_, s298_in_2_, s298_out_0_, n_n856, x7591x}, x263x);
	defparam lut_740.LUT_SIZE = 6;
	defparam lut_740.mask = 64'h5555777701000000;

	lut_sub lut_742 ({sk[261], s298_in_1_, n_n852, n_n854, n_n855}, x7597x);
	defparam lut_742.LUT_SIZE = 5;
	defparam lut_742.mask = 32'h0f5f0100;

	lut_sub lut_744 ({sk[262], s298_in_0_, s298_in_2_, s298_out_4_, n_n858, x7597x}, x264x);
	defparam lut_744.LUT_SIZE = 6;
	defparam lut_744.mask = 64'h5555777700001000;

	lut_sub lut_746 ({sk[263], s298_in_1_, n_n852, n_n855, n_n856}, x7621x);
	defparam lut_746.LUT_SIZE = 5;
	defparam lut_746.mask = 32'h0f5f8000;

	lut_sub lut_748 ({sk[264], s298_in_0_, s298_in_2_, s298_out_4_, n_n857, x7621x}, x268x);
	defparam lut_748.LUT_SIZE = 6;
	defparam lut_748.mask = 64'h5555777701000000;

	lut_sub lut_750 ({sk[265], s298_in_1_, n_n852, n_n853, n_n856}, x7627x);
	defparam lut_750.LUT_SIZE = 5;
	defparam lut_750.mask = 32'h0f5f0400;

	lut_sub lut_752 ({sk[266], s298_in_0_, s298_in_2_, s298_out_4_, n_n857, x7627x}, x269x);
	defparam lut_752.LUT_SIZE = 6;
	defparam lut_752.mask = 64'h5555777700000400;

	lut_sub lut_754 ({sk[267], n_n852, n_n854, n_n855, n_n856}, x7639x);
	defparam lut_754.LUT_SIZE = 5;
	defparam lut_754.mask = 32'h0f5f0002;

	lut_sub lut_756 ({sk[268], s298_in_2_, s298_in_1_, s298_out_5_, n_n858, x7639x}, x271x);
	defparam lut_756.LUT_SIZE = 6;
	defparam lut_756.mask = 64'h5555777700400000;

	lut_sub lut_758 ({sk[269], s298_in_1_, n_n853, n_n854, n_n855}, x7645x);
	defparam lut_758.LUT_SIZE = 5;
	defparam lut_758.mask = 32'h0f5f0010;

	lut_sub lut_760 ({sk[270], s298_in_0_, s298_in_2_, s298_out_5_, n_n858, x7645x}, x272x);
	defparam lut_760.LUT_SIZE = 6;
	defparam lut_760.mask = 64'h5555777740000000;

	lut_sub lut_762 ({sk[271], n_n852, n_n853, n_n854, n_n856}, x7681x);
	defparam lut_762.LUT_SIZE = 5;
	defparam lut_762.mask = 32'h0f5f0100;

	lut_sub lut_764 ({sk[272], s298_in_2_, s298_in_1_, n_n857, n_n52, x7681x}, x278x);
	defparam lut_764.LUT_SIZE = 6;
	defparam lut_764.mask = 64'h5555777700010000;

	lut_sub lut_766 ({sk[273], s298_in_1_, n_n852, n_n853, n_n855}, x7687x);
	defparam lut_766.LUT_SIZE = 5;
	defparam lut_766.mask = 32'h0f5f0200;

	lut_sub lut_768 ({sk[274], s298_in_0_, s298_in_2_, s298_out_3_, n_n857, x7687x}, x279x);
	defparam lut_768.LUT_SIZE = 6;
	defparam lut_768.mask = 64'h5555777700001000;

	lut_sub lut_770 ({sk[275], s298_in_0_, s298_in_2_, n_n852, n_n853}, x7693x);
	defparam lut_770.LUT_SIZE = 5;
	defparam lut_770.mask = 32'h0f5f2000;

	lut_sub lut_772 ({sk[276], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7699x);
	defparam lut_772.LUT_SIZE = 5;
	defparam lut_772.mask = 32'h0f5f0010;

	lut_sub lut_774 ({sk[277], n_n853, n_n854, n_n857, n_n859, x7699x}, x281x);
	defparam lut_774.LUT_SIZE = 6;
	defparam lut_774.mask = 64'h5555777700000400;

	lut_sub lut_776 ({sk[278], s298_in_2_, s298_in_1_, n_n852, n_n853}, x7705x);
	defparam lut_776.LUT_SIZE = 5;
	defparam lut_776.mask = 32'h0f5f2000;

	lut_sub lut_778 ({sk[279], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7711x);
	defparam lut_778.LUT_SIZE = 5;
	defparam lut_778.mask = 32'h0f5f0080;

	lut_sub lut_780 ({sk[280], n_n853, n_n854, n_n857, n_n858, x7711x}, x283x);
	defparam lut_780.LUT_SIZE = 6;
	defparam lut_780.mask = 64'h5555777700000400;

	lut_sub lut_782 ({sk[281], s298_in_0_, s298_in_2_, s298_out_1_, n_n854, n_n855, n_n51}, x7729x);
	defparam lut_782.LUT_SIZE = 7;
	defparam lut_782.mask = 128'h77ff7fff77ff7fff0004000000000000;

	lut_sub lut_784 ({sk[282], s298_in_2_, s298_in_1_, s298_out_4_, n_n852, n_n855, n_n50}, x7734x);
	defparam lut_784.LUT_SIZE = 7;
	defparam lut_784.mask = 128'h77ff7fff77ff7fff0000000800000000;

	lut_sub lut_786 ({sk[283], s298_in_1_, n_n852, n_n855, n_n50, n_n858, n_n859}, x7739x);
	defparam lut_786.LUT_SIZE = 7;
	defparam lut_786.mask = 128'h77ff7fff77ff7fff0000000000000200;

	lut_sub lut_788 ({sk[284], s298_in_2_, s298_in_1_, s298_out_0_, n_n853, n_n856, n_n857}, x7744x);
	defparam lut_788.LUT_SIZE = 7;
	defparam lut_788.mask = 128'h77ff7fff77ff7fff0000000800000000;

	lut_sub lut_790 ({sk[285], s298_in_2_, s298_in_1_, s298_out_5_, n_n856, n_n857, n_n51}, x7749x);
	defparam lut_790.LUT_SIZE = 7;
	defparam lut_790.mask = 128'h77ff7fff77ff7fff0000400000000000;

	lut_sub lut_792 ({sk[286], s298_in_0_, s298_in_1_, s298_out_0_, n_n852, n_n50, n_n857}, x7754x);
	defparam lut_792.LUT_SIZE = 7;
	defparam lut_792.mask = 128'h77ff7fff77ff7fff0000000040000000;

	lut_sub lut_794 ({sk[287], s298_in_0_, s298_in_1_, s298_out_0_, n_n853, n_n854, n_n50}, x7759x);
	defparam lut_794.LUT_SIZE = 7;
	defparam lut_794.mask = 128'h77ff7fff77ff7fff0000000000020000;

	lut_sub lut_796 ({sk[288], s298_in_1_, s298_out_4_, n_n853, n_n855, n_n856, n_n50}, x7764x);
	defparam lut_796.LUT_SIZE = 7;
	defparam lut_796.mask = 128'h77ff7fff77ff7fff0000000000000020;

	lut_sub lut_798 ({sk[289], s298_in_1_, s298_out_5_, n_n852, n_n854, n_n50, n_n51}, x7769x);
	defparam lut_798.LUT_SIZE = 7;
	defparam lut_798.mask = 128'h77ff7fff77ff7fff0040000000000000;

	lut_sub lut_800 ({sk[290], s298_in_0_, s298_in_1_, s298_out_5_, n_n852, n_n855, n_n50}, x7774x);
	defparam lut_800.LUT_SIZE = 7;
	defparam lut_800.mask = 128'h77ff7fff77ff7fff0800000000000000;

	lut_sub lut_802 ({sk[291], s298_in_0_, s298_in_1_, s298_out_0_, n_n852, n_n856, n_n50}, x7779x);
	defparam lut_802.LUT_SIZE = 7;
	defparam lut_802.mask = 128'h77ff7fff77ff7fff0000000000000004;

	lut_sub lut_804 ({sk[292], s298_in_0_, s298_in_1_, n_n852, n_n50, n_n857, n_n51}, x7784x);
	defparam lut_804.LUT_SIZE = 7;
	defparam lut_804.mask = 128'h77ff7fff77ff7fff0000080000000000;

	lut_sub lut_806 ({sk[293], s298_in_0_, s298_in_1_, s298_out_4_, n_n852, n_n854, n_n857}, x7789x);
	defparam lut_806.LUT_SIZE = 7;
	defparam lut_806.mask = 128'h77ff7fff77ff7fff0000000000000080;

	lut_sub lut_808 ({sk[294], s298_in_0_, s298_in_1_, s298_out_5_, n_n853, n_n856, n_n857}, x7794x);
	defparam lut_808.LUT_SIZE = 7;
	defparam lut_808.mask = 128'h77ff7fff77ff7fff0000000000000200;

	lut_sub lut_810 ({sk[295], s298_in_0_, s298_in_1_, n_n852, n_n856, n_n857, n_n51}, x7799x);
	defparam lut_810.LUT_SIZE = 7;
	defparam lut_810.mask = 128'h77ff7fff77ff7fff1000000000000000;

	lut_sub lut_812 ({sk[296], s298_in_0_, s298_in_1_, n_n852, n_n854, n_n856, n_n52}, x7804x);
	defparam lut_812.LUT_SIZE = 7;
	defparam lut_812.mask = 128'h77ff7fff77ff7fff8000000000000000;

	lut_sub lut_814 ({sk[297], s298_in_0_, s298_in_1_, n_n852, n_n855, n_n856, n_n857}, x7809x);
	defparam lut_814.LUT_SIZE = 7;
	defparam lut_814.mask = 128'h77ff7fff77ff7fff0000000000000002;

	lut_sub lut_816 ({sk[298], s298_in_2_, s298_in_1_, s298_out_0_, n_n853, n_n854, n_n856}, x7814x);
	defparam lut_816.LUT_SIZE = 7;
	defparam lut_816.mask = 128'h77ff7fff77ff7fff0008000000000000;

	lut_sub lut_818 ({sk[299], s298_in_2_, s298_in_1_, s298_out_4_, n_n852, n_n855, n_n52}, x7819x);
	defparam lut_818.LUT_SIZE = 7;
	defparam lut_818.mask = 128'h77ff7fff77ff7fff0010000000000000;

	lut_sub lut_820 ({sk[300], s298_in_0_, s298_in_1_, s298_out_0_, n_n852, n_n855, n_n856}, x7824x);
	defparam lut_820.LUT_SIZE = 7;
	defparam lut_820.mask = 128'h77ff7fff77ff7fff0002000000000000;

	lut_sub lut_822 ({sk[301], s298_in_1_, n_n853, n_n854, n_n856, n_n857, n_n858}, x7829x);
	defparam lut_822.LUT_SIZE = 7;
	defparam lut_822.mask = 128'h77ff7fff77ff7fff0002000000000000;

	lut_sub lut_824 ({sk[302], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n855, n_n856}, x7834x);
	defparam lut_824.LUT_SIZE = 7;
	defparam lut_824.mask = 128'h77ff7fff77ff7fff0040000000000000;

	lut_sub lut_826 ({sk[303], s298_in_2_, s298_in_1_, s298_out_0_, n_n853, n_n855, n_n856}, x7839x);
	defparam lut_826.LUT_SIZE = 7;
	defparam lut_826.mask = 128'h77ff7fff77ff7fff0000010000000000;

	lut_sub lut_828 ({sk[304], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n855, n_n857}, x7844x);
	defparam lut_828.LUT_SIZE = 7;
	defparam lut_828.mask = 128'h77ff7fff77ff7fff0000000010000000;

	lut_sub lut_830 ({sk[305], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n855, n_n857}, x7849x);
	defparam lut_830.LUT_SIZE = 7;
	defparam lut_830.mask = 128'h77ff7fff77ff7fff0000000010000000;

	lut_sub lut_832 ({sk[306], s298_in_0_, s298_out_1_, s298_out_4_, n_n853, n_n858}, x7853x);
	defparam lut_832.LUT_SIZE = 6;
	defparam lut_832.mask = 64'h5555777740000000;

	lut_sub lut_834 ({sk[307], s298_in_0_, s298_out_1_, n_n852, n_n854, n_n855}, x7857x);
	defparam lut_834.LUT_SIZE = 6;
	defparam lut_834.mask = 64'h5555777700000008;

	lut_sub lut_836 ({sk[308], s298_in_1_, n_n854, n_n855, n_n50, n_n51}, x7861x);
	defparam lut_836.LUT_SIZE = 6;
	defparam lut_836.mask = 64'h5555777720000000;

	lut_sub lut_838 ({sk[309], s298_in_1_, s298_out_0_, n_n854, n_n855, n_n857}, x7865x);
	defparam lut_838.LUT_SIZE = 6;
	defparam lut_838.mask = 64'h5555777700000080;

	lut_sub lut_840 ({sk[310], s298_in_0_, s298_in_1_, s298_out_0_, n_n852, n_n855}, x7869x);
	defparam lut_840.LUT_SIZE = 6;
	defparam lut_840.mask = 64'h5555777700000400;

	lut_sub lut_842 ({sk[311], s298_in_1_, s298_out_4_, n_n854, n_n855, n_n856}, x7873x);
	defparam lut_842.LUT_SIZE = 6;
	defparam lut_842.mask = 64'h5555777700010000;

	lut_sub lut_844 ({sk[312], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n859}, x7877x);
	defparam lut_844.LUT_SIZE = 6;
	defparam lut_844.mask = 64'h5555777700008000;

	lut_sub lut_846 ({sk[313], s298_in_2_, s298_in_1_, s298_out_4_, n_n852, n_n859}, x7881x);
	defparam lut_846.LUT_SIZE = 6;
	defparam lut_846.mask = 64'h5555777700800000;

	lut_sub lut_848 ({sk[314], s298_in_1_, n_n855, n_n856, n_n858, n_n859}, x7890x);
	defparam lut_848.LUT_SIZE = 6;
	defparam lut_848.mask = 64'h5555777700000010;

	lut_sub lut_850 ({sk[315], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6381x);
	defparam lut_850.LUT_SIZE = 5;
	defparam lut_850.mask = 32'h0f5f0040;

	lut_sub lut_852 ({sk[316], s298_out_4_, n_n853, n_n854, n_n856, n_n857, x6381x}, x6384x);
	defparam lut_852.LUT_SIZE = 7;
	defparam lut_852.mask = 128'h77ff7fff77ff7fff0000400000000000;

	lut_sub lut_854 ({sk[317], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6397x);
	defparam lut_854.LUT_SIZE = 5;
	defparam lut_854.mask = 32'h0f5f4000;

	lut_sub lut_856 ({sk[318], s298_out_5_, n_n853, n_n855, n_n856, n_n857, x6397x}, x6400x);
	defparam lut_856.LUT_SIZE = 7;
	defparam lut_856.mask = 128'h77ff7fff77ff7fff4000000000000000;

	lut_sub lut_858 ({sk[319], s298_in_1_, n_n852, n_n853, n_n854}, x6419x);
	defparam lut_858.LUT_SIZE = 5;
	defparam lut_858.mask = 32'h0f5f0004;

	lut_sub lut_860 ({sk[320], s298_in_0_, s298_in_2_, s298_out_0_, n_n858, x6419x}, x6421x);
	defparam lut_860.LUT_SIZE = 6;
	defparam lut_860.mask = 64'h5555777700001000;

	lut_sub lut_862 ({sk[321], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n855}, x6426x);
	defparam lut_862.LUT_SIZE = 7;
	defparam lut_862.mask = 128'h77ff7fff77ff7fff0000000000080000;

	lut_sub lut_864 ({sk[322], n_n856, n_n857, n_n858, n_n859, x6426x}, x6428x);
	defparam lut_864.LUT_SIZE = 6;
	defparam lut_864.mask = 64'h5555777740444000;

	lut_sub lut_868 ({sk[323], s298_in_1_, n_n852, n_n853, n_n854}, x6482x);
	defparam lut_868.LUT_SIZE = 5;
	defparam lut_868.mask = 32'h0f5f4000;

	lut_sub lut_870 ({sk[324], s298_in_0_, s298_in_2_, s298_out_4_, n_n855, x6482x}, x6484x);
	defparam lut_870.LUT_SIZE = 6;
	defparam lut_870.mask = 64'h5555777700000400;

	lut_sub lut_872 ({sk[325], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6503x);
	defparam lut_872.LUT_SIZE = 5;
	defparam lut_872.mask = 32'h0f5f2000;

	lut_sub lut_874 ({sk[326], n_n853, n_n854, n_n855, n_n857, x6503x}, x6505x);
	defparam lut_874.LUT_SIZE = 6;
	defparam lut_874.mask = 64'h5555777700400000;

	lut_sub lut_876 ({sk[327], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6510x);
	defparam lut_876.LUT_SIZE = 5;
	defparam lut_876.mask = 32'h0f5f1000;

	lut_sub lut_878 ({sk[328], n_n853, n_n854, n_n857, n_n859, x6510x}, x6512x);
	defparam lut_878.LUT_SIZE = 6;
	defparam lut_878.mask = 64'h5555777700000010;

	lut_sub lut_880 ({sk[329], s298_in_1_, n_n852, n_n853, n_n854}, x6524x);
	defparam lut_880.LUT_SIZE = 5;
	defparam lut_880.mask = 32'h0f5f0400;

	lut_sub lut_882 ({sk[330], s298_in_0_, s298_in_2_, s298_out_0_, n_n855, x6524x}, x6526x);
	defparam lut_882.LUT_SIZE = 6;
	defparam lut_882.mask = 64'h5555777700000400;

	lut_sub lut_884 ({sk[331], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6531x);
	defparam lut_884.LUT_SIZE = 5;
	defparam lut_884.mask = 32'h0f5f8000;

	lut_sub lut_886 ({sk[332], s298_out_0_, n_n853, n_n854, n_n855, n_n856, x6531x}, x345x);
	defparam lut_886.LUT_SIZE = 7;
	defparam lut_886.mask = 128'h77ff7fff77ff7fff0000000001000000;

	lut_sub lut_888 ({sk[333], s298_in_1_, n_n852, n_n853, n_n854}, x6538x);
	defparam lut_888.LUT_SIZE = 5;
	defparam lut_888.mask = 32'h0f5f0020;

	lut_sub lut_890 ({sk[334], s298_in_0_, s298_in_2_, s298_out_4_, n_n857, n_n52, x6538x}, x346x);
	defparam lut_890.LUT_SIZE = 7;
	defparam lut_890.mask = 128'h77ff7fff77ff7fff0100000000000000;

	lut_sub lut_892 ({sk[335], s298_in_0_, s298_in_2_, s298_in_1_, n_n853}, x6545x);
	defparam lut_892.LUT_SIZE = 5;
	defparam lut_892.mask = 32'h0f5f8000;

	lut_sub lut_894 ({sk[336], s298_out_4_, n_n854, n_n855, n_n858, n_n859, x6545x}, x347x);
	defparam lut_894.LUT_SIZE = 7;
	defparam lut_894.mask = 128'h77ff7fff77ff7fff0400000000000000;

	lut_sub lut_896 ({sk[337], s298_in_0_, s298_in_2_, s298_in_1_, n_n853}, x6566x);
	defparam lut_896.LUT_SIZE = 5;
	defparam lut_896.mask = 32'h0f5f0080;

	lut_sub lut_898 ({sk[338], s298_out_4_, n_n854, n_n855, n_n856, n_n858, x6566x}, x350x);
	defparam lut_898.LUT_SIZE = 7;
	defparam lut_898.mask = 128'h77ff7fff77ff7fff0000100000000000;

	lut_sub lut_900 ({sk[339], s298_in_1_, n_n852, n_n853, n_n855}, x6573x);
	defparam lut_900.LUT_SIZE = 5;
	defparam lut_900.mask = 32'h0f5f8000;

	lut_sub lut_902 ({sk[340], s298_in_0_, s298_in_2_, s298_out_4_, n_n856, n_n52, x6573x}, x351x);
	defparam lut_902.LUT_SIZE = 7;
	defparam lut_902.mask = 128'h77ff7fff77ff7fff0040000000000000;

	lut_sub lut_904 ({sk[341], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6580x);
	defparam lut_904.LUT_SIZE = 5;
	defparam lut_904.mask = 32'h0f5f2000;

	lut_sub lut_906 ({sk[342], s298_out_4_, n_n853, n_n854, n_n855, n_n857, x6580x}, x352x);
	defparam lut_906.LUT_SIZE = 7;
	defparam lut_906.mask = 128'h77ff7fff77ff7fff0000000004000000;

	lut_sub lut_908 ({sk[343], s298_in_1_, n_n852, n_n853, n_n854}, x6587x);
	defparam lut_908.LUT_SIZE = 5;
	defparam lut_908.mask = 32'h0f5f0200;

	lut_sub lut_910 ({sk[344], s298_in_0_, s298_in_2_, s298_out_5_, n_n856, n_n52, x6587x}, x353x);
	defparam lut_910.LUT_SIZE = 7;
	defparam lut_910.mask = 128'h77ff7fff77ff7fff0100000000000000;

	lut_sub lut_912 ({sk[345], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6594x);
	defparam lut_912.LUT_SIZE = 5;
	defparam lut_912.mask = 32'h0f5f0040;

	lut_sub lut_914 ({sk[346], n_n853, n_n854, n_n855, n_n858, x6594x}, x6596x);
	defparam lut_914.LUT_SIZE = 6;
	defparam lut_914.mask = 64'h5555777700040000;

	lut_sub lut_916 ({sk[347], s298_in_1_, n_n852, n_n855, n_n856}, x6601x);
	defparam lut_916.LUT_SIZE = 5;
	defparam lut_916.mask = 32'h0f5f0010;

	lut_sub lut_918 ({sk[348], s298_in_0_, s298_in_2_, n_n857, n_n51, n_n52, x6601x}, x355x);
	defparam lut_918.LUT_SIZE = 7;
	defparam lut_918.mask = 128'h77ff7fff77ff7fff0000000010000000;

	lut_sub lut_920 ({sk[349], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6622x);
	defparam lut_920.LUT_SIZE = 5;
	defparam lut_920.mask = 32'h0f5f0040;

	lut_sub lut_922 ({sk[350], n_n853, n_n854, n_n856, n_n857, x6622x}, x6624x);
	defparam lut_922.LUT_SIZE = 6;
	defparam lut_922.mask = 64'h5555777700100000;

	lut_sub lut_924 ({sk[351], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6629x);
	defparam lut_924.LUT_SIZE = 5;
	defparam lut_924.mask = 32'h0f5f0040;

	lut_sub lut_926 ({sk[352], n_n853, n_n854, n_n855, n_n856, x6629x}, x6631x);
	defparam lut_926.LUT_SIZE = 6;
	defparam lut_926.mask = 64'h5555777740000000;

	lut_sub lut_928 ({sk[353], s298_in_0_, s298_in_2_, n_n856, n_n857, n_n859}, x6645x);
	defparam lut_928.LUT_SIZE = 6;
	defparam lut_928.mask = 64'h5555777780000000;

	lut_sub lut_930 ({sk[354], s298_in_0_, s298_in_2_, n_n855, n_n856, n_n859}, x6652x);
	defparam lut_930.LUT_SIZE = 6;
	defparam lut_930.mask = 64'h5555777740000000;

	lut_sub lut_932 ({sk[355], s298_in_1_, n_n852, n_n853, n_n854, x6652x}, x362x);
	defparam lut_932.LUT_SIZE = 6;
	defparam lut_932.mask = 64'h5555777700000040;

	lut_sub lut_934 ({sk[356], s298_in_0_, s298_in_2_, n_n856, n_n857, n_n859}, x6659x);
	defparam lut_934.LUT_SIZE = 6;
	defparam lut_934.mask = 64'h5555777704000000;

	lut_sub lut_936 ({sk[357], s298_in_0_, s298_in_2_, n_n855, n_n856, n_n858}, x6666x);
	defparam lut_936.LUT_SIZE = 6;
	defparam lut_936.mask = 64'h5555777700004000;

	lut_sub lut_938 ({sk[358], s298_in_1_, n_n852, n_n853, n_n854, x6666x}, x364x);
	defparam lut_938.LUT_SIZE = 6;
	defparam lut_938.mask = 64'h5555777700004000;

	lut_sub lut_940 ({sk[359], s298_in_0_, s298_in_2_, n_n855, n_n857, n_n858}, x6687x);
	defparam lut_940.LUT_SIZE = 6;
	defparam lut_940.mask = 64'h5555777700002000;

	lut_sub lut_942 ({sk[360], s298_in_0_, s298_in_2_, n_n856, n_n857, n_n858}, x6694x);
	defparam lut_942.LUT_SIZE = 6;
	defparam lut_942.mask = 64'h5555777700000200;

	lut_sub lut_944 ({sk[361], s298_in_1_, n_n852, n_n854, n_n855, x6694x}, x368x);
	defparam lut_944.LUT_SIZE = 6;
	defparam lut_944.mask = 64'h5555777700000004;

	lut_sub lut_946 ({sk[362], s298_in_0_, s298_in_2_, n_n856, n_n857, n_n858}, x6701x);
	defparam lut_946.LUT_SIZE = 6;
	defparam lut_946.mask = 64'h5555777701000000;

	lut_sub lut_948 ({sk[363], s298_in_1_, n_n852, n_n853, n_n855}, x6820x);
	defparam lut_948.LUT_SIZE = 5;
	defparam lut_948.mask = 32'h0f5f0020;

	lut_sub lut_950 ({sk[364], s298_in_0_, s298_in_2_, n_n856, x6820x}, x6821x);
	defparam lut_950.LUT_SIZE = 5;
	defparam lut_950.mask = 32'h0f5f0010;

	lut_sub lut_952 ({sk[365], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n854, n_n855}, x6832x);
	defparam lut_952.LUT_SIZE = 7;
	defparam lut_952.mask = 128'h77ff7fff77ff7fff0000000040000000;

	lut_sub lut_954 ({sk[366], s298_out_4_, n_n52, x6832x}, x391x);
	defparam lut_954.LUT_SIZE = 4;
	defparam lut_954.mask = 16'h3304;

	lut_sub lut_956 ({sk[367], s298_in_1_, n_n852, n_n853, n_n854}, x6850x);
	defparam lut_956.LUT_SIZE = 5;
	defparam lut_956.mask = 32'h0f5f0400;

	lut_sub lut_958 ({sk[368], s298_in_0_, s298_in_2_, s298_out_4_, n_n855, x6850x}, x394x);
	defparam lut_958.LUT_SIZE = 6;
	defparam lut_958.mask = 64'h5555777704000000;

	lut_sub lut_960 ({sk[369], s298_in_1_, n_n852, n_n853, n_n856}, x6856x);
	defparam lut_960.LUT_SIZE = 5;
	defparam lut_960.mask = 32'h0f5f0100;

	lut_sub lut_962 ({sk[370], s298_in_0_, s298_in_2_, s298_out_4_, n_n857, x6856x}, x395x);
	defparam lut_962.LUT_SIZE = 6;
	defparam lut_962.mask = 64'h5555777700000400;

	lut_sub lut_964 ({sk[371], s298_in_1_, n_n852, n_n853, n_n855}, x6874x);
	defparam lut_964.LUT_SIZE = 5;
	defparam lut_964.mask = 32'h0f5f1000;

	lut_sub lut_966 ({sk[372], s298_in_0_, s298_in_2_, n_n856, n_n52, x6874x}, x398x);
	defparam lut_966.LUT_SIZE = 6;
	defparam lut_966.mask = 64'h5555777700000400;

	lut_sub lut_968 ({sk[373], n_n852, n_n853, n_n855, n_n856}, x6880x);
	defparam lut_968.LUT_SIZE = 5;
	defparam lut_968.mask = 32'h0f5f0010;

	lut_sub lut_970 ({sk[374], s298_in_2_, s298_in_1_, n_n857, x6880x}, x6881x);
	defparam lut_970.LUT_SIZE = 5;
	defparam lut_970.mask = 32'h0f5f4000;

	lut_sub lut_972 ({sk[375], s298_in_1_, n_n854, n_n855, n_n856}, x6892x);
	defparam lut_972.LUT_SIZE = 5;
	defparam lut_972.mask = 32'h0f5f0100;

	lut_sub lut_974 ({sk[376], s298_in_0_, s298_in_2_, n_n857, n_n52, x6892x}, x401x);
	defparam lut_974.LUT_SIZE = 6;
	defparam lut_974.mask = 64'h5555777701000000;

	lut_sub lut_976 ({sk[377], s298_in_1_, n_n852, n_n854, n_n856}, x6898x);
	defparam lut_976.LUT_SIZE = 5;
	defparam lut_976.mask = 32'h0f5f0008;

	lut_sub lut_978 ({sk[378], s298_in_0_, s298_in_2_, s298_out_2_, n_n857, x6898x}, x402x);
	defparam lut_978.LUT_SIZE = 6;
	defparam lut_978.mask = 64'h5555777700001000;

	lut_sub lut_980 ({sk[379], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6910x);
	defparam lut_980.LUT_SIZE = 5;
	defparam lut_980.mask = 32'h0f5f0010;

	lut_sub lut_982 ({sk[380], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6916x);
	defparam lut_982.LUT_SIZE = 5;
	defparam lut_982.mask = 32'h0f5f4000;

	lut_sub lut_984 ({sk[381], n_n853, n_n856, n_n858, n_n859}, x6923x);
	defparam lut_984.LUT_SIZE = 5;
	defparam lut_984.mask = 32'h0f5f0002;

	lut_sub lut_986 ({sk[382], n_n855, n_n856, n_n858, n_n859}, x6929x);
	defparam lut_986.LUT_SIZE = 5;
	defparam lut_986.mask = 32'h0f5f0200;

	lut_sub lut_988 ({sk[383], s298_in_0_, s298_in_2_, s298_in_1_, n_n853}, x6934x);
	defparam lut_988.LUT_SIZE = 5;
	defparam lut_988.mask = 32'h0f5f0020;

	lut_sub lut_990 ({sk[384], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6940x);
	defparam lut_990.LUT_SIZE = 5;
	defparam lut_990.mask = 32'h0f5f0080;

	lut_sub lut_992 ({sk[385], n_n853, n_n854, n_n856, n_n857, x6940x}, x409x);
	defparam lut_992.LUT_SIZE = 6;
	defparam lut_992.mask = 64'h5555777700001000;

	lut_sub lut_994 ({sk[386], n_n853, n_n856, n_n857, n_n858}, x6947x);
	defparam lut_994.LUT_SIZE = 5;
	defparam lut_994.mask = 32'h0f5f0200;

	lut_sub lut_996 ({sk[387], n_n853, n_n855, n_n857, n_n858}, x6953x);
	defparam lut_996.LUT_SIZE = 5;
	defparam lut_996.mask = 32'h0f5f0010;

	lut_sub lut_998 ({sk[388], s298_in_0_, s298_in_2_, s298_in_1_, n_n853}, x6958x);
	defparam lut_998.LUT_SIZE = 5;
	defparam lut_998.mask = 32'h0f5f1000;

	lut_sub lut_1000 ({sk[389], n_n855, n_n856, n_n857, n_n858}, x6959x);
	defparam lut_1000.LUT_SIZE = 5;
	defparam lut_1000.mask = 32'h0f5f0200;

	lut_sub lut_1002 ({sk[390], s298_in_2_, s298_in_1_, s298_out_4_, n_n855, n_n856, n_n50}, x6964x);
	defparam lut_1002.LUT_SIZE = 7;
	defparam lut_1002.mask = 128'h77ff7fff77ff7fff0000002000000000;

	lut_sub lut_1004 ({sk[391], s298_in_1_, s298_out_5_, n_n854, n_n855, n_n50, n_n857}, x6969x);
	defparam lut_1004.LUT_SIZE = 7;
	defparam lut_1004.mask = 128'h77ff7fff77ff7fff0000002000000000;

	lut_sub lut_1006 ({sk[392], s298_in_2_, s298_in_1_, n_n852, n_n854, n_n856, n_n858}, x6974x);
	defparam lut_1006.LUT_SIZE = 7;
	defparam lut_1006.mask = 128'h77ff7fff77ff7fff0000002000000000;

	lut_sub lut_1008 ({sk[393], s298_in_1_, s298_out_0_, n_n854, n_n855, n_n856, n_n50}, x6979x);
	defparam lut_1008.LUT_SIZE = 7;
	defparam lut_1008.mask = 128'h77ff7fff77ff7fff0000000000000100;

	lut_sub lut_1010 ({sk[394], s298_in_1_, s298_out_5_, n_n853, n_n854, n_n855, n_n856}, x6984x);
	defparam lut_1010.LUT_SIZE = 7;
	defparam lut_1010.mask = 128'h77ff7fff77ff7fff0008000000000000;

	lut_sub lut_1012 ({sk[395], s298_in_0_, s298_in_1_, s298_out_5_, n_n852, n_n853, n_n855}, x6989x);
	defparam lut_1012.LUT_SIZE = 7;
	defparam lut_1012.mask = 128'h77ff7fff77ff7fff0000000000000100;

	lut_sub lut_1014 ({sk[396], s298_in_1_, s298_out_5_, n_n853, n_n854, n_n856, n_n857}, x6994x);
	defparam lut_1014.LUT_SIZE = 7;
	defparam lut_1014.mask = 128'h77ff7fff77ff7fff0000008000000000;

	lut_sub lut_1016 ({sk[397], s298_in_1_, n_n852, n_n853, n_n854, n_n856, n_n52}, x6999x);
	defparam lut_1016.LUT_SIZE = 7;
	defparam lut_1016.mask = 128'h77ff7fff77ff7fff0000000001000000;

	lut_sub lut_1018 ({sk[398], s298_in_0_, s298_in_1_, n_n853, n_n854, n_n855, n_n859}, x7004x);
	defparam lut_1018.LUT_SIZE = 7;
	defparam lut_1018.mask = 128'h77ff7fff77ff7fff4000000000000000;

	lut_sub lut_1020 ({sk[399], s298_in_0_, s298_in_1_, n_n853, n_n854, n_n855, n_n856}, x7009x);
	defparam lut_1020.LUT_SIZE = 7;
	defparam lut_1020.mask = 128'h77ff7fff77ff7fff0000000000000002;

	lut_sub lut_1022 ({sk[400], s298_in_1_, n_n852, n_n855, n_n856, n_n857, n_n858}, x7014x);
	defparam lut_1022.LUT_SIZE = 7;
	defparam lut_1022.mask = 128'h77ff7fff77ff7fff0000000200000000;

	lut_sub lut_1024 ({sk[401], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_1_, n_n853, n_n855}, x7019x);
	defparam lut_1024.LUT_SIZE = 7;
	defparam lut_1024.mask = 128'h77ff7fff77ff7fff0000000000040000;

	lut_sub lut_1026 ({sk[402], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_1_, n_n852, n_n51}, x7024x);
	defparam lut_1026.LUT_SIZE = 7;
	defparam lut_1026.mask = 128'h77ff7fff77ff7fff0000000008000000;

	lut_sub lut_1028 ({sk[403], s298_in_2_, s298_in_1_, n_n852, n_n853, n_n855, n_n856}, x7029x);
	defparam lut_1028.LUT_SIZE = 7;
	defparam lut_1028.mask = 128'h77ff7fff77ff7fff0000100000000000;

	lut_sub lut_1030 ({sk[404], s298_in_2_, s298_in_1_, n_n852, n_n853, n_n855, n_n856}, x7034x);
	defparam lut_1030.LUT_SIZE = 7;
	defparam lut_1030.mask = 128'h77ff7fff77ff7fff0000000100000000;

	lut_sub lut_1032 ({sk[405], s298_in_2_, s298_in_1_, n_n853, n_n856, n_n52, n_n859}, x7039x);
	defparam lut_1032.LUT_SIZE = 7;
	defparam lut_1032.mask = 128'h77ff7fff77ff7fff0800000000000000;

	lut_sub lut_1034 ({sk[406], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_3_, n_n852, n_n855}, x7044x);
	defparam lut_1034.LUT_SIZE = 7;
	defparam lut_1034.mask = 128'h77ff7fff77ff7fff0004000000000000;

	lut_sub lut_1036 ({sk[407], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n855, n_n51}, x7049x);
	defparam lut_1036.LUT_SIZE = 7;
	defparam lut_1036.mask = 128'h77ff7fff77ff7fff0000000800000000;

	lut_sub lut_1038 ({sk[408], s298_in_0_, s298_in_1_, n_n852, n_n854, n_n857, n_n51}, x7054x);
	defparam lut_1038.LUT_SIZE = 7;
	defparam lut_1038.mask = 128'h77ff7fff77ff7fff0000000000000400;

	lut_sub lut_1040 ({sk[409], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_4_, n_n853, n_n856}, x7059x);
	defparam lut_1040.LUT_SIZE = 7;
	defparam lut_1040.mask = 128'h77ff7fff77ff7fff0000000002000000;

	lut_sub lut_1042 ({sk[410], s298_in_2_, s298_in_1_, n_n852, n_n853, n_n855, n_n857}, x7064x);
	defparam lut_1042.LUT_SIZE = 7;
	defparam lut_1042.mask = 128'h77ff7fff77ff7fff0000400000000000;

	lut_sub lut_1044 ({sk[411], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n855, n_n856}, x7069x);
	defparam lut_1044.LUT_SIZE = 7;
	defparam lut_1044.mask = 128'h77ff7fff77ff7fff0002000000000000;

	lut_sub lut_1046 ({sk[412], s298_in_2_, s298_in_1_, n_n852, n_n853, n_n855, n_n857}, x7074x);
	defparam lut_1046.LUT_SIZE = 7;
	defparam lut_1046.mask = 128'h77ff7fff77ff7fff0100000000000000;

	lut_sub lut_1048 ({sk[413], s298_in_2_, s298_in_1_, n_n852, n_n855, n_n856, n_n857}, x7079x);
	defparam lut_1048.LUT_SIZE = 7;
	defparam lut_1048.mask = 128'h77ff7fff77ff7fff0000100000000000;

	lut_sub lut_1050 ({sk[414], s298_in_1_, n_n855, n_n857, n_n858}, x7084x);
	defparam lut_1050.LUT_SIZE = 5;
	defparam lut_1050.mask = 32'h0f5f0002;

	lut_sub lut_1052 ({sk[415], s298_in_1_, s298_out_4_, n_n855, n_n856, n_n50}, x7088x);
	defparam lut_1052.LUT_SIZE = 6;
	defparam lut_1052.mask = 64'h5555777700040000;

	lut_sub lut_1054 ({sk[416], s298_in_1_, s298_out_0_, n_n853, n_n857, n_n858}, x7092x);
	defparam lut_1054.LUT_SIZE = 6;
	defparam lut_1054.mask = 64'h5555777700000010;

	lut_sub lut_1056 ({sk[417], s298_in_0_, s298_in_1_, s298_out_4_, n_n852, n_n856}, x7096x);
	defparam lut_1056.LUT_SIZE = 6;
	defparam lut_1056.mask = 64'h5555777701000000;

	lut_sub lut_1058 ({sk[418], s298_in_1_, n_n852, n_n853, n_n49, n_n856, n_n858}, x441x);
	defparam lut_1058.LUT_SIZE = 7;
	defparam lut_1058.mask = 128'h77ff7fff77ff7fff0000040000000000;

	lut_sub lut_1060 ({sk[419], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_1_, n_n854, n_n855}, x442x);
	defparam lut_1060.LUT_SIZE = 7;
	defparam lut_1060.mask = 128'h77ff7fff77ff7fff0002000000000000;

	lut_sub lut_1062 ({sk[420], s298_in_1_, s298_out_4_, n_n853, n_n51, n_n859}, x7108x);
	defparam lut_1062.LUT_SIZE = 6;
	defparam lut_1062.mask = 64'h5555777700010000;

	lut_sub lut_1064 ({sk[421], s298_in_2_, s298_in_1_, s298_out_2_, n_n852, n_n51, n_n52}, x444x);
	defparam lut_1064.LUT_SIZE = 7;
	defparam lut_1064.mask = 128'h77ff7fff77ff7fff0000000200000000;

	lut_sub lut_1066 ({sk[422], s298_in_0_, s298_in_2_, n_n855, n_n856, n_n858}, x5520x);
	defparam lut_1066.LUT_SIZE = 6;
	defparam lut_1066.mask = 64'h5555777708000000;

	lut_sub lut_1068 ({sk[423], s298_in_2_, s298_in_1_, n_n852, n_n853, n_n855, n_n856}, x5797x);
	defparam lut_1068.LUT_SIZE = 7;
	defparam lut_1068.mask = 128'h77ff7fff77ff7fff0000200000000000;

	lut_sub lut_1070 ({sk[424], s298_out_5_, n_n856, n_n859, x5527x, x5797x}, x5798x);
	defparam lut_1070.LUT_SIZE = 6;
	defparam lut_1070.mask = 64'h5555777711115111;

	lut_sub lut_1073 ({sk[425], x5798x, x5785x, x5786x, x5787x, x5788x, x5789x}, x447x);
	defparam lut_1073.LUT_SIZE = 7;
	defparam lut_1073.mask = 128'h77ff7fff77ff7fff0000000080000000;

	lut_sub lut_1075 ({sk[426], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n855}, x6024x);
	defparam lut_1075.LUT_SIZE = 7;
	defparam lut_1075.mask = 128'h77ff7fff77ff7fff0040000000000000;

	lut_sub lut_1077 ({sk[427], s298_out_0_, x6024x}, x6025x);
	defparam lut_1077.LUT_SIZE = 3;
	defparam lut_1077.mask = 8'h51;

	lut_sub lut_1079 ({sk[428], s298_in_2_, n_n852, n_n853, n_n854, n_n855, n_n858}, x6030x);
	defparam lut_1079.LUT_SIZE = 7;
	defparam lut_1079.mask = 128'h77ff7fff77ff7fff0040000000000000;

	lut_sub lut_1081 ({sk[429], n_n855, n_n856, n_n857, n_n858, n_n859, x6030x}, x6031x);
	defparam lut_1081.LUT_SIZE = 7;
	defparam lut_1081.mask = 128'h77ff7fff77ff7fff5454541154545410;

	lut_sub lut_1086 ({sk[430], s298_in_2_, n_n852, n_n853, n_n854}, x6053x);
	defparam lut_1086.LUT_SIZE = 5;
	defparam lut_1086.mask = 32'h05ff0400;

	lut_sub lut_1088 ({sk[431], n_n856, n_n857, n_n858, n_n859, x6053x}, x6055x);
	defparam lut_1088.LUT_SIZE = 6;
	defparam lut_1088.mask = 64'h337f337f00010005;

	lut_sub lut_1091 ({sk[432], s298_in_1_, n_n852, n_n854, n_n855}, x6072x);
	defparam lut_1091.LUT_SIZE = 5;
	defparam lut_1091.mask = 32'h05ff0004;

	lut_sub lut_1093 ({sk[433], s298_in_0_, s298_in_2_, n_n857, x6072x}, x6073x);
	defparam lut_1093.LUT_SIZE = 5;
	defparam lut_1093.mask = 32'h05ff0040;

	lut_sub lut_1095 ({sk[434], s298_in_0_, s298_in_2_, n_n852, n_n853, n_n854, n_n857}, x6078x);
	defparam lut_1095.LUT_SIZE = 7;
	defparam lut_1095.mask = 128'h77ff7fff77ff7fff0000000000400000;

	lut_sub lut_1097 ({sk[435], n_n855, n_n856, n_n857, n_n858, n_n859, x6078x}, x6079x);
	defparam lut_1097.LUT_SIZE = 7;
	defparam lut_1097.mask = 128'h77ff7fff77ff7fff0101014401010145;

	lut_sub lut_1103 ({sk[436], x6079x, x5785x, x5786x, x5787x, x5788x, x5789x}, x457x);
	defparam lut_1103.LUT_SIZE = 7;
	defparam lut_1103.mask = 128'h77ff7fff77ff7fff0000000080000000;

	lut_sub lut_1105 ({sk[437], s298_in_1_, n_n852, n_n853, n_n854}, x6084x);
	defparam lut_1105.LUT_SIZE = 5;
	defparam lut_1105.mask = 32'h05ff0001;

	lut_sub lut_1107 ({sk[438], s298_in_0_, s298_in_2_, s298_out_4_, n_n857, x6084x}, x458x);
	defparam lut_1107.LUT_SIZE = 6;
	defparam lut_1107.mask = 64'h337f337f00000100;

	lut_sub lut_1109 ({sk[439], s298_in_1_, n_n852, n_n853, n_n857}, x6102x);
	defparam lut_1109.LUT_SIZE = 5;
	defparam lut_1109.mask = 32'h05ff0010;

	lut_sub lut_1111 ({sk[440], s298_in_0_, s298_in_2_, n_n858, x6102x}, x6103x);
	defparam lut_1111.LUT_SIZE = 5;
	defparam lut_1111.mask = 32'h05ff0040;

	lut_sub lut_1113 ({sk[441], n_n852, n_n853, n_n854, n_n856}, x6108x);
	defparam lut_1113.LUT_SIZE = 5;
	defparam lut_1113.mask = 32'h05ff0004;

	lut_sub lut_1115 ({sk[442], s298_in_0_, s298_in_2_, n_n857, x6108x}, x6109x);
	defparam lut_1115.LUT_SIZE = 5;
	defparam lut_1115.mask = 32'h05ff1000;

	lut_sub lut_1117 ({sk[443], x6109x, x5785x, x5786x, x5787x, x5788x, x5789x}, x462x);
	defparam lut_1117.LUT_SIZE = 7;
	defparam lut_1117.mask = 128'h77ff7fff77ff7fff0000000080000000;

	lut_sub lut_1119 ({sk[444], s298_in_1_, n_n852, n_n854, n_n856}, x6114x);
	defparam lut_1119.LUT_SIZE = 5;
	defparam lut_1119.mask = 32'h05ff0200;

	lut_sub lut_1121 ({sk[445], s298_in_0_, s298_in_2_, n_n859, x6114x}, x6115x);
	defparam lut_1121.LUT_SIZE = 5;
	defparam lut_1121.mask = 32'h05ff0040;

	lut_sub lut_1123 ({sk[446], x6115x, x5785x, x5786x, x5787x, x5788x, x5789x}, x463x);
	defparam lut_1123.LUT_SIZE = 7;
	defparam lut_1123.mask = 128'h77ff7fff77ff7fff000000007fffffff;

	lut_sub lut_1129 ({sk[447], s298_in_1_, n_n852, n_n854, n_n855}, x6120x);
	defparam lut_1129.LUT_SIZE = 5;
	defparam lut_1129.mask = 32'h05ff0100;

	lut_sub lut_1131 ({sk[448], s298_in_0_, s298_in_2_, s298_out_2_, n_n857, x6120x}, x464x);
	defparam lut_1131.LUT_SIZE = 6;
	defparam lut_1131.mask = 64'h337f337f10000000;

	lut_sub lut_1133 ({sk[449], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6126x);
	defparam lut_1133.LUT_SIZE = 5;
	defparam lut_1133.mask = 32'h05ff0010;

	lut_sub lut_1135 ({sk[450], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6132x);
	defparam lut_1135.LUT_SIZE = 5;
	defparam lut_1135.mask = 32'h05ff1000;

	lut_sub lut_1137 ({sk[451], s298_in_0_, s298_in_2_, s298_out_1_, n_n852, n_n853, n_n854}, x6150x);
	defparam lut_1137.LUT_SIZE = 7;
	defparam lut_1137.mask = 128'h77ff7fff77ff7fff0001000000000000;

	lut_sub lut_1139 ({sk[452], s298_in_2_, n_n852, n_n853, n_n854, n_n855, n_n856}, x6155x);
	defparam lut_1139.LUT_SIZE = 7;
	defparam lut_1139.mask = 128'h77ff7fff77ff7fff0000800000000000;

	lut_sub lut_1141 ({sk[453], s298_in_2_, s298_in_1_, n_n852, n_n853, n_n854, n_n855}, x6160x);
	defparam lut_1141.LUT_SIZE = 7;
	defparam lut_1141.mask = 128'h77ff7fff77ff7fff0000002000000000;

	lut_sub lut_1143 ({sk[454], s298_in_0_, s298_in_1_, s298_out_0_, n_n857, n_n51, n_n52}, x6165x);
	defparam lut_1143.LUT_SIZE = 7;
	defparam lut_1143.mask = 128'h77ff7fff77ff7fff0000001000000000;

	lut_sub lut_1145 ({sk[455], s298_in_0_, s298_in_1_, s298_out_0_, n_n852, n_n854, n_n855}, x6170x);
	defparam lut_1145.LUT_SIZE = 7;
	defparam lut_1145.mask = 128'h77ff7fff77ff7fff0000000400000000;

	lut_sub lut_1147 ({sk[456], s298_in_0_, s298_in_1_, s298_out_4_, n_n854, n_n855, n_n856}, x6175x);
	defparam lut_1147.LUT_SIZE = 7;
	defparam lut_1147.mask = 128'h77ff7fff77ff7fff0000000000020000;

	lut_sub lut_1149 ({sk[457], s298_in_0_, s298_in_1_, s298_out_5_, n_n852, n_n857, n_n859}, x6180x);
	defparam lut_1149.LUT_SIZE = 7;
	defparam lut_1149.mask = 128'h77ff7fff77ff7fff0800000000000000;

	lut_sub lut_1151 ({sk[458], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n854, n_n52}, x6185x);
	defparam lut_1151.LUT_SIZE = 7;
	defparam lut_1151.mask = 128'h77ff7fff77ff7fff0000001000000000;

	lut_sub lut_1153 ({sk[459], s298_in_0_, s298_in_1_, n_n854, n_n855, n_n856, n_n857}, x6190x);
	defparam lut_1153.LUT_SIZE = 7;
	defparam lut_1153.mask = 128'h77ff7fff77ff7fff0000000000800000;

	lut_sub lut_1155 ({sk[460], s298_in_2_, n_n852, n_n855, n_n856, n_n857, n_n858}, x6195x);
	defparam lut_1155.LUT_SIZE = 7;
	defparam lut_1155.mask = 128'h77ff7fff77ff7fff0000000200000000;

	lut_sub lut_1157 ({sk[461], s298_in_2_, s298_out_0_, n_n852, n_n855, n_n856, n_n857}, x6200x);
	defparam lut_1157.LUT_SIZE = 7;
	defparam lut_1157.mask = 128'h77ff7fff77ff7fff0008000000000000;

	lut_sub lut_1159 ({sk[462], x6200x, x5785x, x5786x, x5787x, x5788x, x5789x}, x479x);
	defparam lut_1159.LUT_SIZE = 7;
	defparam lut_1159.mask = 128'h77ff7fff77ff7fff000000007fffffff;

	lut_sub lut_1165 ({sk[463], s298_in_2_, n_n853, n_n854, n_n855, n_n857, n_n858}, x6210x);
	defparam lut_1165.LUT_SIZE = 7;
	defparam lut_1165.mask = 128'h77ff7fff77ff7fff0000200000000000;

	lut_sub lut_1167 ({sk[464], s298_in_2_, n_n852, n_n854, n_n855, n_n856, n_n857}, x6215x);
	defparam lut_1167.LUT_SIZE = 7;
	defparam lut_1167.mask = 128'h77ff7fff77ff7fff0000000800000000;

	lut_sub lut_1169 ({sk[465], s298_in_2_, s298_in_1_, s298_out_4_, n_n852, n_n854, n_n857}, x6220x);
	defparam lut_1169.LUT_SIZE = 7;
	defparam lut_1169.mask = 128'h77ff7fff77ff7fff0000000400000000;

	lut_sub lut_1171 ({sk[466], x6220x, x5785x, x5786x, x5787x, x5788x, x5789x}, x483x);
	defparam lut_1171.LUT_SIZE = 7;
	defparam lut_1171.mask = 128'h77ff7fff77ff7fff0000000080000000;

	lut_sub lut_1173 ({sk[467], s298_in_2_, s298_in_1_, s298_out_4_, n_n853, n_n854, n_n857}, x6225x);
	defparam lut_1173.LUT_SIZE = 7;
	defparam lut_1173.mask = 128'h77ff7fff77ff7fff0001000000000000;

	lut_sub lut_1175 ({sk[468], x6225x, x5785x, x5786x, x5787x, x5788x, x5789x}, x484x);
	defparam lut_1175.LUT_SIZE = 7;
	defparam lut_1175.mask = 128'h77ff7fff77ff7fff0000000080000000;

	lut_sub lut_1177 ({sk[469], s298_in_2_, s298_out_4_, n_n853, n_n854, n_n855, n_n856}, x6230x);
	defparam lut_1177.LUT_SIZE = 7;
	defparam lut_1177.mask = 128'h77ff7fff77ff7fff0000000800000000;

	lut_sub lut_1179 ({sk[470], x6230x, x5785x, x5786x, x5787x, x5788x, x5789x}, x485x);
	defparam lut_1179.LUT_SIZE = 7;
	defparam lut_1179.mask = 128'h77ff7fff77ff7fff0000000080000000;

	lut_sub lut_1181 ({sk[471], s298_in_2_, n_n853, n_n854, n_n855, n_n856, n_n857}, x6235x);
	defparam lut_1181.LUT_SIZE = 7;
	defparam lut_1181.mask = 128'h77ff7fff77ff7fff0000080000000000;

	lut_sub lut_1183 ({sk[472], s298_in_2_, s298_out_5_, n_n852, n_n854, n_n855, n_n856}, x6240x);
	defparam lut_1183.LUT_SIZE = 7;
	defparam lut_1183.mask = 128'h77ff7fff77ff7fff4000000000000000;

	lut_sub lut_1185 ({sk[473], s298_in_2_, n_n852, n_n853, n_n854, n_n855, n_n858}, x6245x);
	defparam lut_1185.LUT_SIZE = 7;
	defparam lut_1185.mask = 128'h77ff7fff77ff7fff0200000000000000;

	lut_sub lut_1187 ({sk[474], s298_in_2_, n_n852, n_n853, n_n855, n_n856, n_n858}, x6250x);
	defparam lut_1187.LUT_SIZE = 7;
	defparam lut_1187.mask = 128'h77ff7fff77ff7fff2000000000000000;

	lut_sub lut_1189 ({sk[475], s298_in_2_, n_n852, n_n853, n_n854, n_n855, n_n856}, x6255x);
	defparam lut_1189.LUT_SIZE = 7;
	defparam lut_1189.mask = 128'h77ff7fff77ff7fff1000000000000000;

	lut_sub lut_1191 ({sk[476], s298_in_2_, n_n853, n_n854, n_n855, n_n856, n_n857}, x6260x);
	defparam lut_1191.LUT_SIZE = 7;
	defparam lut_1191.mask = 128'h77ff7fff77ff7fff0000000400000000;

	lut_sub lut_1193 ({sk[477], s298_in_2_, n_n852, n_n853, n_n855, n_n856, n_n857}, x6265x);
	defparam lut_1193.LUT_SIZE = 7;
	defparam lut_1193.mask = 128'h77ff7fff77ff7fff0400000000000000;

	lut_sub lut_1195 ({sk[478], s298_in_1_, n_n854, n_n857, n_n858}, x6270x);
	defparam lut_1195.LUT_SIZE = 5;
	defparam lut_1195.mask = 32'h05ff0002;

	lut_sub lut_1197 ({sk[479], s298_in_2_, s298_out_1_, n_n852, n_n854, n_n856}, x6274x);
	defparam lut_1197.LUT_SIZE = 6;
	defparam lut_1197.mask = 64'h337f337f00010000;

	lut_sub lut_1199 ({sk[480], s298_in_0_, s298_in_2_, n_n852, n_n853, n_n855}, x6278x);
	defparam lut_1199.LUT_SIZE = 6;
	defparam lut_1199.mask = 64'h337f337f00002000;

	lut_sub lut_1201 ({sk[481], s298_in_2_, s298_out_0_, n_n852, n_n853, n_n51}, x6282x);
	defparam lut_1201.LUT_SIZE = 6;
	defparam lut_1201.mask = 64'h337f337f00100000;

	lut_sub lut_1203 ({sk[482], s298_in_2_, n_n856, n_n857, n_n51, n_n858}, x6294x);
	defparam lut_1203.LUT_SIZE = 6;
	defparam lut_1203.mask = 64'h337f337f00800000;

	lut_sub lut_1205 ({sk[483], s298_in_2_, n_n852, n_n854, n_n855, n_n859}, x6298x);
	defparam lut_1205.LUT_SIZE = 6;
	defparam lut_1205.mask = 64'h337f337f00080000;

	lut_sub lut_1207 ({sk[484], s298_in_2_, n_n853, n_n854, n_n856, n_n858}, x6306x);
	defparam lut_1207.LUT_SIZE = 6;
	defparam lut_1207.mask = 64'h337f337f00080000;

	lut_sub lut_1209 ({sk[485], s298_in_2_, n_n853, n_n854, n_n855, n_n857, n_n858}, x503x);
	defparam lut_1209.LUT_SIZE = 7;
	defparam lut_1209.mask = 128'h77ff7fff77ff7fff0000080000000000;

	lut_sub lut_1211 ({sk[486], s298_in_0_, s298_in_2_, s298_out_0_, n_n859}, x6313x);
	defparam lut_1211.LUT_SIZE = 5;
	defparam lut_1211.mask = 32'h05ff0020;

	lut_sub lut_1213 ({sk[487], s298_in_2_, n_n856, n_n857, n_n51, n_n858, n_n859}, x6315x);
	defparam lut_1213.LUT_SIZE = 7;
	defparam lut_1213.mask = 128'h77ff7fff77ff7fff0002000000000000;

	lut_sub lut_1215 ({sk[488], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x5803x);
	defparam lut_1215.LUT_SIZE = 5;
	defparam lut_1215.mask = 32'h05ff0040;

	lut_sub lut_1217 ({sk[489], s298_out_0_, n_n854, n_n855, n_n856, n_n857, x5803x}, x507x);
	defparam lut_1217.LUT_SIZE = 7;
	defparam lut_1217.mask = 128'h77ff7fff77ff7fff0000000000040000;

	lut_sub lut_1219 ({sk[490], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x5810x);
	defparam lut_1219.LUT_SIZE = 5;
	defparam lut_1219.mask = 32'h05ff8000;

	lut_sub lut_1221 ({sk[491], n_n854, n_n856, n_n857, n_n858, x5810x}, x5812x);
	defparam lut_1221.LUT_SIZE = 6;
	defparam lut_1221.mask = 64'h337f337f00000040;

	lut_sub lut_1223 ({sk[492], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n854, n_n857}, x5823x);
	defparam lut_1223.LUT_SIZE = 7;
	defparam lut_1223.mask = 128'h77ff7fff77ff7fff0000000004000000;

	lut_sub lut_1225 ({sk[493], n_n855, n_n856, n_n857, n_n858, n_n859, x5823x}, x5824x);
	defparam lut_1225.LUT_SIZE = 7;
	defparam lut_1225.mask = 128'h77ff7fff77ff7fff0101014401010145;

	lut_sub lut_1231 ({sk[494], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n854, n_n856}, x5829x);
	defparam lut_1231.LUT_SIZE = 7;
	defparam lut_1231.mask = 128'h77ff7fff77ff7fff0001000000000000;

	lut_sub lut_1233 ({sk[495], n_n855, n_n856, n_n857, n_n858, n_n859, x5829x}, x5830x);
	defparam lut_1233.LUT_SIZE = 7;
	defparam lut_1233.mask = 128'h77ff7fff77ff7fff0101014401010145;

	lut_sub lut_1239 ({sk[496], s298_in_1_, n_n852, n_n853, n_n854}, x5841x);
	defparam lut_1239.LUT_SIZE = 5;
	defparam lut_1239.mask = 32'h05ff0800;

	lut_sub lut_1241 ({sk[497], s298_in_0_, s298_in_2_, n_n857, x5841x}, x5842x);
	defparam lut_1241.LUT_SIZE = 5;
	defparam lut_1241.mask = 32'h05ff1000;

	lut_sub lut_1243 ({sk[498], s298_in_0_, s298_in_2_, n_n852, n_n854}, x5847x);
	defparam lut_1243.LUT_SIZE = 5;
	defparam lut_1243.mask = 32'h05ff1000;

	lut_sub lut_1245 ({sk[499], n_n855, n_n856, n_n857, n_n858}, x5848x);
	defparam lut_1245.LUT_SIZE = 5;
	defparam lut_1245.mask = 32'h05ff0400;

	lut_sub lut_1247 ({sk[500], s298_in_2_, s298_out_3_, n_n852, n_n853, n_n854, n_n857}, x5858x);
	defparam lut_1247.LUT_SIZE = 7;
	defparam lut_1247.mask = 128'h77ff7fff77ff7fff0400000000000000;

	lut_sub lut_1249 ({sk[501], s298_in_2_, s298_out_0_, n_n852, n_n853, n_n854, n_n856}, x5868x);
	defparam lut_1249.LUT_SIZE = 7;
	defparam lut_1249.mask = 128'h77ff7fff77ff7fff0000040000000000;

	lut_sub lut_1251 ({sk[502], s298_in_2_, s298_out_0_, n_n853, n_n854, n_n856, n_n857}, x5873x);
	defparam lut_1251.LUT_SIZE = 7;
	defparam lut_1251.mask = 128'h77ff7fff77ff7fff0000000400000000;

	lut_sub lut_1253 ({sk[503], x5873x, x5785x, x5786x, x5787x, x5788x, x5789x}, x519x);
	defparam lut_1253.LUT_SIZE = 7;
	defparam lut_1253.mask = 128'h77ff7fff77ff7fff000000007fffffff;

	lut_sub lut_1259 ({sk[504], s298_in_2_, n_n852, n_n854, n_n855, n_n856, n_n857}, x5878x);
	defparam lut_1259.LUT_SIZE = 7;
	defparam lut_1259.mask = 128'h77ff7fff77ff7fff0800000000000000;

	lut_sub lut_1261 ({sk[505], s298_in_2_, n_n852, n_n855, n_n856, n_n857, n_n858}, x5883x);
	defparam lut_1261.LUT_SIZE = 7;
	defparam lut_1261.mask = 128'h77ff7fff77ff7fff0800000000000000;

	lut_sub lut_1263 ({sk[506], s298_in_2_, s298_out_5_, n_n852, n_n854, n_n855, n_n856}, x5888x);
	defparam lut_1263.LUT_SIZE = 7;
	defparam lut_1263.mask = 128'h77ff7fff77ff7fff0100000000000000;

	lut_sub lut_1265 ({sk[507], n_n852, n_n853, n_n854, n_n855, n_n858, n_n859}, x5893x);
	defparam lut_1265.LUT_SIZE = 7;
	defparam lut_1265.mask = 128'h77ff7fff77ff7fff0020000000000000;

	lut_sub lut_1267 ({sk[508], n_n852, n_n853, n_n854, n_n856, n_n857, n_n858}, x5898x);
	defparam lut_1267.LUT_SIZE = 7;
	defparam lut_1267.mask = 128'h77ff7fff77ff7fff0000000000000002;

	lut_sub lut_1269 ({sk[509], s298_in_0_, s298_in_2_, n_n857}, x5902x);
	defparam lut_1269.LUT_SIZE = 4;
	defparam lut_1269.mask = 16'h3f04;

	lut_sub lut_1271 ({sk[510], n_n853, n_n854, n_n855, n_n856}, x5903x);
	defparam lut_1271.LUT_SIZE = 5;
	defparam lut_1271.mask = 32'h05ff0100;

	lut_sub lut_1273 ({sk[511], s298_in_2_, s298_out_0_, s298_out_2_, n_n852, n_n855}, x5907x);
	defparam lut_1273.LUT_SIZE = 6;
	defparam lut_1273.mask = 64'h337f337f02000000;

	lut_sub lut_1275 ({sk[512], x5907x, x5785x, x5786x, x5787x, x5788x, x5789x}, x526x);
	defparam lut_1275.LUT_SIZE = 7;
	defparam lut_1275.mask = 128'h77ff7fff77ff7fff000000007fffffff;

	lut_sub lut_1281 ({sk[513], s298_in_2_, n_n853, n_n854, n_n856, n_n857}, x5911x);
	defparam lut_1281.LUT_SIZE = 6;
	defparam lut_1281.mask = 64'h337f337f01000000;

	lut_sub lut_1283 ({sk[514], s298_in_0_, s298_in_2_, s298_out_0_, n_n852, n_n853, n_n859}, x528x);
	defparam lut_1283.LUT_SIZE = 7;
	defparam lut_1283.mask = 128'h77ff7fff77ff7fff0000000000800000;

	lut_sub lut_1285 ({sk[515], s298_in_2_, n_n853, n_n854, n_n856, n_n857}, x5919x);
	defparam lut_1285.LUT_SIZE = 6;
	defparam lut_1285.mask = 64'h337f337f00800000;

	lut_sub lut_1287 ({sk[516], s298_in_2_, s298_out_0_, n_n852, n_n853, n_n857, n_n858}, x530x);
	defparam lut_1287.LUT_SIZE = 7;
	defparam lut_1287.mask = 128'h77ff7fff77ff7fff0000080000000000;

	lut_sub lut_1289 ({sk[517], s298_in_2_, s298_out_4_, n_n852, n_n51, n_n858}, x5927x);
	defparam lut_1289.LUT_SIZE = 6;
	defparam lut_1289.mask = 64'h337f337f01000000;

	lut_sub lut_1291 ({sk[518], x5927x, x5785x, x5786x, x5787x, x5788x, x5789x}, x531x);
	defparam lut_1291.LUT_SIZE = 7;
	defparam lut_1291.mask = 128'h77ff7fff77ff7fff000000007fffffff;

	lut_sub lut_1297 ({sk[519], s298_in_2_, s298_out_4_, n_n853, n_n854, n_n855, n_n856}, x532x);
	defparam lut_1297.LUT_SIZE = 7;
	defparam lut_1297.mask = 128'h77ff7fff77ff7fff0000004000000000;

	lut_sub lut_1299 ({sk[520], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_3_, n_n853}, x5935x);
	defparam lut_1299.LUT_SIZE = 6;
	defparam lut_1299.mask = 64'h337f337f00000100;

	lut_sub lut_1301 ({sk[521], s298_in_2_, n_n852, n_n853, n_n854, n_n857}, x5943x);
	defparam lut_1301.LUT_SIZE = 6;
	defparam lut_1301.mask = 64'h337f337f10000000;

	lut_sub lut_1303 ({sk[522], x5943x, x5785x, x5786x, x5787x, x5788x, x5789x}, x535x);
	defparam lut_1303.LUT_SIZE = 7;
	defparam lut_1303.mask = 128'h77ff7fff77ff7fff000000007fffffff;

	lut_sub lut_1309 ({sk[523], s298_in_2_, n_n853, n_n855, n_n856, n_n857}, x5947x);
	defparam lut_1309.LUT_SIZE = 6;
	defparam lut_1309.mask = 64'h337f337f00020000;

	lut_sub lut_1311 ({sk[524], s298_in_2_, n_n852, n_n854, n_n855, n_n856, n_n857}, x537x);
	defparam lut_1311.LUT_SIZE = 7;
	defparam lut_1311.mask = 128'h77ff7fff77ff7fff0000100000000000;

	lut_sub lut_1313 ({sk[525], s298_in_2_, n_n854, n_n855, n_n856, n_n857, n_n858}, x538x);
	defparam lut_1313.LUT_SIZE = 7;
	defparam lut_1313.mask = 128'h77ff7fff77ff7fff0100000000000000;

	lut_sub lut_1315 ({sk[526], s298_in_2_, n_n854, n_n857, n_n858}, x5961x);
	defparam lut_1315.LUT_SIZE = 5;
	defparam lut_1315.mask = 32'h05ff0200;

	lut_sub lut_1317 ({sk[527], n_n854, n_n855, n_n856, n_n858, n_n859}, x5967x);
	defparam lut_1317.LUT_SIZE = 6;
	defparam lut_1317.mask = 64'h337f337f40000000;

	lut_sub lut_1319 ({sk[528], s298_in_0_, s298_in_2_, n_n853, n_n859}, x5970x);
	defparam lut_1319.LUT_SIZE = 5;
	defparam lut_1319.mask = 32'h05ff2000;

	lut_sub lut_1321 ({sk[529], n_n854, n_n855, n_n856, n_n857, n_n858, n_n859}, x5973x);
	defparam lut_1321.LUT_SIZE = 7;
	defparam lut_1321.mask = 128'h77ff7fff77ff7fff000000e400000000;

	lut_sub lut_1324 ({sk[530], s298_in_0_, s298_out_1_, s298_out_4_, n_n852, n_n853, n_n854}, x548x);
	defparam lut_1324.LUT_SIZE = 7;
	defparam lut_1324.mask = 128'h77ff7fff77ff7fff0000000400000000;

	lut_sub lut_1326 ({sk[531], n_n852, n_n853, n_n854, n_n855, n_n856}, x5535x);
	defparam lut_1326.LUT_SIZE = 6;
	defparam lut_1326.mask = 64'h337f337f00000020;

	lut_sub lut_1328 ({sk[532], s298_in_0_, s298_in_1_, s298_out_4_, n_n853, n_n854, n_n859}, x550x);
	defparam lut_1328.LUT_SIZE = 7;
	defparam lut_1328.mask = 128'h77ff7fff77ff7fff0000000000000020;

	lut_sub lut_1330 ({sk[533], n_n853, n_n854, n_n855, n_n856, n_n857}, x5543x);
	defparam lut_1330.LUT_SIZE = 6;
	defparam lut_1330.mask = 64'h337f337f00000002;

	lut_sub lut_1332 ({sk[534], s298_out_3_, n_n852, n_n853, n_n854, n_n856, n_n857}, x553x);
	defparam lut_1332.LUT_SIZE = 7;
	defparam lut_1332.mask = 128'h77ff7fff77ff7fff0400000000000000;

	lut_sub lut_1334 ({sk[535], n_n852, n_n853, n_n854, n_n855, n_n856, n_n857}, x554x);
	defparam lut_1334.LUT_SIZE = 7;
	defparam lut_1334.mask = 128'h77ff7fff77ff7fff0000000000020000;

	lut_sub lut_1336 ({sk[536], s298_out_0_, s298_out_2_, n_n852, n_n855, n_n857}, x556x);
	defparam lut_1336.LUT_SIZE = 6;
	defparam lut_1336.mask = 64'h337f337f00040000;

	lut_sub lut_1338 ({sk[537], n_n853, n_n855, n_n856, n_n857}, x5729x);
	defparam lut_1338.LUT_SIZE = 5;
	defparam lut_1338.mask = 32'h05ff0040;

	lut_sub lut_1340 ({sk[538], s298_out_2_, n_n853, n_n854, n_n855, n_n859}, x558x);
	defparam lut_1340.LUT_SIZE = 6;
	defparam lut_1340.mask = 64'h337f337f02000000;

	lut_sub lut_1342 ({sk[539], s298_in_1_, s298_out_4_, n_n852}, x5740x);
	defparam lut_1342.LUT_SIZE = 4;
	defparam lut_1342.mask = 16'h3f20;

	lut_sub lut_1344 ({sk[540], s298_in_1_, n_n857, n_n859}, x5748x);
	defparam lut_1344.LUT_SIZE = 4;
	defparam lut_1344.mask = 16'h3f08;

	lut_sub lut_1346 ({sk[541], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x5548x);
	defparam lut_1346.LUT_SIZE = 5;
	defparam lut_1346.mask = 32'h05ff2000;

	lut_sub lut_1348 ({sk[542], n_n853, n_n854, n_n856, n_n859}, x5549x);
	defparam lut_1348.LUT_SIZE = 5;
	defparam lut_1348.mask = 32'h05ff0200;

	lut_sub lut_1350 ({sk[543], s298_in_2_, s298_in_1_, n_n852, n_n853}, x5554x);
	defparam lut_1350.LUT_SIZE = 5;
	defparam lut_1350.mask = 32'h05ff4000;

	lut_sub lut_1352 ({sk[544], n_n854, n_n855, n_n856, n_n857}, x5555x);
	defparam lut_1352.LUT_SIZE = 5;
	defparam lut_1352.mask = 32'h05ff1000;

	lut_sub lut_1354 ({sk[545], s298_in_0_, s298_in_2_, n_n852, n_n853}, x5560x);
	defparam lut_1354.LUT_SIZE = 5;
	defparam lut_1354.mask = 32'h05ff0040;

	lut_sub lut_1356 ({sk[546], s298_in_2_, s298_in_1_, n_n852, n_n853}, x5566x);
	defparam lut_1356.LUT_SIZE = 5;
	defparam lut_1356.mask = 32'h05ff8000;

	lut_sub lut_1358 ({sk[547], s298_in_0_, s298_in_2_, n_n852, n_n853}, x5572x);
	defparam lut_1358.LUT_SIZE = 5;
	defparam lut_1358.mask = 32'h05ff8000;

	lut_sub lut_1360 ({sk[548], n_n854, n_n855, n_n856, n_n857}, x5573x);
	defparam lut_1360.LUT_SIZE = 5;
	defparam lut_1360.mask = 32'h05ff0010;

	lut_sub lut_1362 ({sk[549], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x5578x);
	defparam lut_1362.LUT_SIZE = 5;
	defparam lut_1362.mask = 32'h05ff4000;

	lut_sub lut_1364 ({sk[550], n_n854, n_n855, n_n856, n_n858}, x5579x);
	defparam lut_1364.LUT_SIZE = 5;
	defparam lut_1364.mask = 32'h05ff0002;

	lut_sub lut_1366 ({sk[551], s298_in_2_, n_n852, n_n853, n_n855, n_n857, n_n859}, x589x);
	defparam lut_1366.LUT_SIZE = 7;
	defparam lut_1366.mask = 128'h77ff7fff77ff7fff0000080000000000;

	lut_sub lut_1368 ({sk[552], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n855, n_n859}, x590x);
	defparam lut_1368.LUT_SIZE = 7;
	defparam lut_1368.mask = 128'h77ff7fff77ff7fff0000000008000000;

	lut_sub lut_1370 ({sk[553], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n856, n_n859}, x591x);
	defparam lut_1370.LUT_SIZE = 7;
	defparam lut_1370.mask = 128'h77ff7fff77ff7fff0000000000020000;

	lut_sub lut_1372 ({sk[554], n_n852, n_n853, n_n854, n_n856, n_n857, n_n858}, x592x);
	defparam lut_1372.LUT_SIZE = 7;
	defparam lut_1372.mask = 128'h77ff7fff77ff7fff2000000000000000;

	lut_sub lut_1374 ({sk[555], n_n852, n_n853, n_n854, n_n855, n_n856, n_n857}, x595x);
	defparam lut_1374.LUT_SIZE = 7;
	defparam lut_1374.mask = 128'h77ff7fff77ff7fff0000000000000010;

	lut_sub lut_1376 ({sk[556], s298_in_2_, n_n852, n_n853, n_n854, n_n856, n_n858}, x596x);
	defparam lut_1376.LUT_SIZE = 7;
	defparam lut_1376.mask = 128'h77ff7fff77ff7fff0000000200000000;

	lut_sub lut_1378 ({sk[557], s298_in_2_, n_n853, n_n854, n_n856, n_n857, n_n858}, x600x);
	defparam lut_1378.LUT_SIZE = 7;
	defparam lut_1378.mask = 128'h77ff7fff77ff7fff0000000800000000;

	lut_sub lut_1380 ({sk[558], n_n853, n_n854, n_n855, n_n857, n_n859}, x602x);
	defparam lut_1380.LUT_SIZE = 6;
	defparam lut_1380.mask = 64'h337f337f08000000;

	lut_sub lut_1382 ({sk[559], n_n852, n_n853, n_n854, n_n857, n_n859}, x5672x);
	defparam lut_1382.LUT_SIZE = 6;
	defparam lut_1382.mask = 64'h337f337f00a02020;

	lut_sub lut_1385 ({sk[560], s298_in_2_, n_n852, n_n854, n_n856, n_n857, n_n859}, x5673x);
	defparam lut_1385.LUT_SIZE = 7;
	defparam lut_1385.mask = 128'h77ff7fff77ff7fff0800aa0008000800;

	lut_sub lut_1388 ({sk[561], n_n853, n_n854, n_n855, n_n857, n_n858, n_n859}, x5674x);
	defparam lut_1388.LUT_SIZE = 7;
	defparam lut_1388.mask = 128'h77ff7fff77ff7fff00008888000a888a;

	lut_sub lut_1391 ({sk[562], n_n852, n_n853, n_n854, n_n855, n_n857, n_n858}, x5681x);
	defparam lut_1391.LUT_SIZE = 7;
	defparam lut_1391.mask = 128'h77ff7fff77ff7fff0210000000000000;

	lut_sub lut_1394 ({sk[563], n_n852, n_n854, n_n855, n_n856, n_n857, n_n858}, x5683x);
	defparam lut_1394.LUT_SIZE = 7;
	defparam lut_1394.mask = 128'h77ff7fff77ff7fff0000000000002008;

	lut_sub lut_1397 ({sk[564], n_n852, n_n853, n_n854, n_n855, n_n857, n_n858}, x5689x);
	defparam lut_1397.LUT_SIZE = 7;
	defparam lut_1397.mask = 128'h77ff7fff77ff7fff0000100010001000;

	lut_sub lut_1400 ({sk[565], n_n853, n_n854, n_n855, n_n856, n_n857, n_n858}, x12839x);
	defparam lut_1400.LUT_SIZE = 7;
	defparam lut_1400.mask = 128'h77ff7fff77ff7fffffffffffffffdff7;

	lut_sub lut_1410 ({sk[566], n_n853, n_n855, n_n856, n_n857, n_n858, n_n859}, x12838x);
	defparam lut_1410.LUT_SIZE = 7;
	defparam lut_1410.mask = 128'h77ff7fff77ff7ffffffe77555ffe7755;

	lut_sub lut_1423 ({sk[567], n_n852, n_n853, n_n854, n_n855, n_n857, n_n858}, x5765x);
	defparam lut_1423.LUT_SIZE = 7;
	defparam lut_1423.mask = 128'h77ff7fff77ff7fff00000202aa000202;

	lut_sub lut_1426 ({sk[568], x553x, x5765x}, x5767x);
	defparam lut_1426.LUT_SIZE = 3;
	defparam lut_1426.mask = 8'h57;

	lut_sub lut_1429 ({sk[569], s298_out_5_, n_n855, n_n857, n_n858, x5543x, x554x}, x5768x);
	defparam lut_1429.LUT_SIZE = 7;
	defparam lut_1429.mask = 128'h77ff7fff77ff7ffff7777777f5555555;

	lut_sub lut_1433 ({sk[570], s298_in_2_, s298_in_1_, s298_out_5_, n_n856, n_n858}, x5770x);
	defparam lut_1433.LUT_SIZE = 6;
	defparam lut_1433.mask = 64'h337f337f8000a0a0;

	lut_sub lut_1436 ({sk[571], s298_in_0_, s298_out_5_, n_n852, n_n858, x5748x, x5770x}, x5772x);
	defparam lut_1436.LUT_SIZE = 7;
	defparam lut_1436.mask = 128'h77ff7fff77ff7fff77f7555577775555;

	lut_sub lut_1440 ({sk[572], s298_out_1_, s298_out_4_, n_n854, n_n855, n_n858, x5535x}, x5775x);
	defparam lut_1440.LUT_SIZE = 7;
	defparam lut_1440.mask = 128'h77ff7fff77ff7fff3000000055555555;

	lut_sub lut_1443 ({sk[573], s298_out_0_, n_n852, n_n855, n_n858, x5729x}, x5780x);
	defparam lut_1443.LUT_SIZE = 6;
	defparam lut_1443.mask = 64'h337f337fd5550000;

	lut_sub lut_1446 ({sk[574], s298_in_0_, s298_out_0_, n_n852, n_n853, n_n856, n_n858}, x5781x);
	defparam lut_1446.LUT_SIZE = 7;
	defparam lut_1446.mask = 128'h77ff7fff77ff7fff20200000aa200000;

	lut_sub lut_1449 ({sk[575], s298_out_0_, n_n852, n_n853, n_n857, n_n859}, x5783x);
	defparam lut_1449.LUT_SIZE = 6;
	defparam lut_1449.mask = 64'h337f337f0000440a;

	lut_sub lut_1452 ({sk[576], n_n852, n_n853, n_n854, n_n855, n_n856, n_n857}, x12837x);
	defparam lut_1452.LUT_SIZE = 7;
	defparam lut_1452.mask = 128'h77ff7fff77ff7fffbb3fbbffbbffbbff;

	lut_sub lut_1461 ({sk[577], s298_in_0_, s298_in_2_, n_n857}, x5816x);
	defparam lut_1461.LUT_SIZE = 4;
	defparam lut_1461.mask = 16'h3f04;

	lut_sub lut_1463 ({sk[578], s298_in_1_, n_n852, n_n854, n_n856}, x5817x);
	defparam lut_1463.LUT_SIZE = 5;
	defparam lut_1463.mask = 32'h05ff0010;

	lut_sub lut_1465 ({sk[579], s298_in_1_, n_n853, n_n855, n_n858}, x5835x);
	defparam lut_1465.LUT_SIZE = 5;
	defparam lut_1465.mask = 32'h05ff0040;

	lut_sub lut_1467 ({sk[580], s298_in_2_, n_n852, n_n854, n_n855, n_n856}, x5852x);
	defparam lut_1467.LUT_SIZE = 6;
	defparam lut_1467.mask = 64'h337f337f00040000;

	lut_sub lut_1469 ({sk[581], s298_in_2_, n_n853, n_n854, n_n856, n_n857}, x5862x);
	defparam lut_1469.LUT_SIZE = 6;
	defparam lut_1469.mask = 64'h337f337f40000000;

	lut_sub lut_1471 ({sk[582], x5847x, x5848x, x5902x, x5903x, x537x, x538x}, x5983x);
	defparam lut_1471.LUT_SIZE = 7;
	defparam lut_1471.mask = 128'h77ff7fff77ff7fff777f777f777fffff;

	lut_sub lut_1476 ({sk[583], s298_in_0_, s298_in_2_, s298_out_5_, n_n859, x5893x, x5835x}, x5984x);
	defparam lut_1476.LUT_SIZE = 7;
	defparam lut_1476.mask = 128'h77ff7fff77ff7fff7300330033003300;

	lut_sub lut_1479 ({sk[584], x532x, x5983x, x5984x}, x5986x);
	defparam lut_1479.LUT_SIZE = 4;
	defparam lut_1479.mask = 16'h3f7f;

	lut_sub lut_1483 ({sk[585], s298_out_0_, s298_out_4_, x5816x, x5817x, x5852x}, x5992x);
	defparam lut_1483.LUT_SIZE = 6;
	defparam lut_1483.mask = 64'h337f337f03570000;

	lut_sub lut_1486 ({sk[586], s298_in_2_, s298_out_0_, n_n855, n_n857, n_n51, x5961x}, x5997x);
	defparam lut_1486.LUT_SIZE = 7;
	defparam lut_1486.mask = 128'h77ff7fff77ff7fff5557000055550000;

	lut_sub lut_1489 ({sk[587], s298_out_0_, n_n852, n_n853, n_n857, n_n51, x5970x}, x5998x);
	defparam lut_1489.LUT_SIZE = 7;
	defparam lut_1489.mask = 128'h77ff7fff77ff7fff0000000055555575;

	lut_sub lut_1492 ({sk[588], n_n51, x5812x, x5888x, x5898x, x5986x}, x5999x);
	defparam lut_1492.LUT_SIZE = 6;
	defparam lut_1492.mask = 64'h337f337f55ff7f7f;

	lut_sub lut_1497 ({sk[589], s298_in_2_, n_n852, n_n854, n_n855, n_n856, n_n857}, x12836x);
	defparam lut_1497.LUT_SIZE = 7;
	defparam lut_1497.mask = 128'h77ff7fff77ff7ffffffff8fffffffaff;

	lut_sub lut_1503 ({sk[590], s298_out_4_, n_n854, n_n855, n_n51, x5935x, x12836x}, x6000x);
	defparam lut_1503.LUT_SIZE = 7;
	defparam lut_1503.mask = 128'h77ff7fff77ff7fff0b0b0b0b0b0f0b0b;

	lut_sub lut_1507 ({sk[591], n_n853, n_n855, n_n857, n_n51, x507x, x5992x}, x6001x);
	defparam lut_1507.LUT_SIZE = 7;
	defparam lut_1507.mask = 128'h77ff7fff77ff7fff777777777777777f;

	lut_sub lut_1511 ({sk[592], s298_out_0_, n_n51, x5858x, x5878x, x5883x, x5862x}, x6002x);
	defparam lut_1511.LUT_SIZE = 7;
	defparam lut_1511.mask = 128'h77ff7fff77ff7fff00ff00ff7f7f3f3f;

	lut_sub lut_1516 ({sk[593], s298_out_0_, x5911x, x528x, x5919x, x530x}, x6003x);
	defparam lut_1516.LUT_SIZE = 6;
	defparam lut_1516.mask = 64'h337f337f5fff7f7f;

	lut_sub lut_1521 ({sk[594], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_4_, n_n854, n_n856}, x6036x);
	defparam lut_1521.LUT_SIZE = 7;
	defparam lut_1521.mask = 128'h77ff7fff77ff7fff0000000000010000;

	lut_sub lut_1523 ({sk[595], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n854}, x6042x);
	defparam lut_1523.LUT_SIZE = 7;
	defparam lut_1523.mask = 128'h77ff7fff77ff7fff0000000001000000;

	lut_sub lut_1525 ({sk[596], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n856}, x6048x);
	defparam lut_1525.LUT_SIZE = 7;
	defparam lut_1525.mask = 128'h77ff7fff77ff7fff0010000000000000;

	lut_sub lut_1527 ({sk[597], s298_in_0_, s298_in_1_, n_n854, n_n855, n_n856, n_n857}, x6060x);
	defparam lut_1527.LUT_SIZE = 7;
	defparam lut_1527.mask = 128'h77ff7fff77ff7fff0000000000000004;

	lut_sub lut_1529 ({sk[598], s298_in_0_, s298_in_2_, n_n853, n_n854}, x6065x);
	defparam lut_1529.LUT_SIZE = 5;
	defparam lut_1529.mask = 32'h05ff1000;

	lut_sub lut_1531 ({sk[599], n_n856, n_n857, n_n858, n_n859}, x6066x);
	defparam lut_1531.LUT_SIZE = 5;
	defparam lut_1531.mask = 32'h05ff2022;

	lut_sub lut_1534 ({sk[600], s298_in_1_, n_n852, n_n853, n_n855}, x6090x);
	defparam lut_1534.LUT_SIZE = 5;
	defparam lut_1534.mask = 32'h05ff1000;

	lut_sub lut_1536 ({sk[601], s298_in_0_, s298_in_2_, n_n858}, x6095x);
	defparam lut_1536.LUT_SIZE = 4;
	defparam lut_1536.mask = 16'h3f08;

	lut_sub lut_1538 ({sk[602], s298_in_1_, n_n852, n_n853, n_n855}, x6096x);
	defparam lut_1538.LUT_SIZE = 5;
	defparam lut_1538.mask = 32'h05ff1000;

	lut_sub lut_1540 ({sk[603], s298_in_2_, n_n852, n_n854, n_n856, n_n857}, x6204x);
	defparam lut_1540.LUT_SIZE = 6;
	defparam lut_1540.mask = 64'h337f337f00100000;

	lut_sub lut_1542 ({sk[604], s298_in_2_, n_n852, n_n854, n_n855}, x6301x);
	defparam lut_1542.LUT_SIZE = 5;
	defparam lut_1542.mask = 32'h05ff0400;

	lut_sub lut_1544 ({sk[605], n_n853, n_n854, n_n856, n_n858, x6126x, x6132x}, x6318x);
	defparam lut_1544.LUT_SIZE = 7;
	defparam lut_1544.mask = 128'h77ff7fff77ff7fff0030000000500000;

	lut_sub lut_1547 ({sk[606], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n854}, x12834x);
	defparam lut_1547.LUT_SIZE = 7;
	defparam lut_1547.mask = 128'h77ff7fff77ff7fffbfbfffff15bfffff;

	lut_sub lut_1557 ({sk[607], n_n855, n_n856, n_n857, n_n858, x12834x}, x6319x);
	defparam lut_1557.LUT_SIZE = 6;
	defparam lut_1557.mask = 64'h337f337f00080000;

	lut_sub lut_1559 ({sk[608], s298_in_0_, s298_in_2_, n_n859, x6270x, x503x}, x6320x);
	defparam lut_1559.LUT_SIZE = 6;
	defparam lut_1559.mask = 64'h337f337f75555555;

	lut_sub lut_1562 ({sk[609], s298_in_1_, n_n852, n_n853, n_n854, x5520x, x6318x}, x6321x);
	defparam lut_1562.LUT_SIZE = 7;
	defparam lut_1562.mask = 128'h77ff7fff77ff7fff7555555555555555;

	lut_sub lut_1565 ({sk[610], s298_out_5_, x6245x, x6250x, x6306x, x6095x, x6096x}, x6326x);
	defparam lut_1565.LUT_SIZE = 7;
	defparam lut_1565.mask = 128'h77ff7fff77ff7fff1fffffff00000000;

	lut_sub lut_1570 ({sk[611], s298_in_0_, s298_in_2_, s298_out_4_, n_n856, x6235x, x6090x}, x6328x);
	defparam lut_1570.LUT_SIZE = 7;
	defparam lut_1570.mask = 128'h77ff7fff77ff7fff0073003300330033;

	lut_sub lut_1573 ({sk[612], s298_out_1_, s298_out_4_, s298_out_5_, n_n858, x6278x, x6301x}, x6331x);
	defparam lut_1573.LUT_SIZE = 7;
	defparam lut_1573.mask = 128'h77ff7fff77ff7fff5000000073333333;

	lut_sub lut_1576 ({sk[613], s298_out_1_, x464x, x6155x, x6160x, x6326x}, x6336x);
	defparam lut_1576.LUT_SIZE = 6;
	defparam lut_1576.mask = 64'h337f337f55ff7fff;

	lut_sub lut_1581 ({sk[614], x458x, x6319x, x6320x, x6321x, x6328x, x6331x}, x6337x);
	defparam lut_1581.LUT_SIZE = 7;
	defparam lut_1581.mask = 128'h77ff7fff77ff7fff7fffffffffffffff;

	lut_sub lut_1588 ({sk[615], s298_out_0_, n_n855, n_n857, n_n51, x6103x, x6150x}, x6340x);
	defparam lut_1588.LUT_SIZE = 7;
	defparam lut_1588.mask = 128'h77ff7fff77ff7fff070707070f070707;

	lut_sub lut_1592 ({sk[616], n_n51, x6240x, x6255x, x6260x, x6265x}, x6341x);
	defparam lut_1592.LUT_SIZE = 6;
	defparam lut_1592.mask = 64'h337f337f3f3f55ff;

	lut_sub lut_1597 ({sk[617], s298_out_0_, n_n51, x6073x, x6210x, x6215x, x6204x}, x6343x);
	defparam lut_1597.LUT_SIZE = 7;
	defparam lut_1597.mask = 128'h77ff7fff77ff7fff000000007fff3fff;

	lut_sub lut_1602 ({sk[618], x6336x, x6337x, x6340x, x6341x, x6343x}, x6346x);
	defparam lut_1602.LUT_SIZE = 6;
	defparam lut_1602.mask = 64'h337f337f7fffffff;

	lut_sub lut_1608 ({sk[619], x457x, x462x, x463x, x479x}, x6352x);
	defparam lut_1608.LUT_SIZE = 5;
	defparam lut_1608.mask = 32'h05ff7fff;

	lut_sub lut_1613 ({sk[620], x447x, x483x, x484x, x485x, x6346x}, x6353x);
	defparam lut_1613.LUT_SIZE = 6;
	defparam lut_1613.mask = 64'h337f337f7fffffff;

	lut_sub lut_1619 ({sk[621], x6018x, x6165x, x6016x, x6017x, x6065x, x6066x}, x6359x);
	defparam lut_1619.LUT_SIZE = 7;
	defparam lut_1619.mask = 128'h77ff7fff77ff7fff01110fff1111ffff;

	lut_sub lut_1626 ({sk[622], x6018x, x6170x, x6175x, x6016x, x6017x}, x6360x);
	defparam lut_1626.LUT_SIZE = 6;
	defparam lut_1626.mask = 64'h337f337f07770fff;

	lut_sub lut_1633 ({sk[623], x6018x, x6180x, x6185x, x6016x, x6017x}, x6361x);
	defparam lut_1633.LUT_SIZE = 6;
	defparam lut_1633.mask = 64'h337f337f07770fff;

	lut_sub lut_1640 ({sk[624], x6018x, x6190x, x6195x, x6016x, x6017x}, x6362x);
	defparam lut_1640.LUT_SIZE = 6;
	defparam lut_1640.mask = 64'h337f337f07770fff;

	lut_sub lut_1647 ({sk[625], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6389x);
	defparam lut_1647.LUT_SIZE = 5;
	defparam lut_1647.mask = 32'h05ff1000;

	lut_sub lut_1649 ({sk[626], n_n853, n_n855, n_n856, n_n857}, x6390x);
	defparam lut_1649.LUT_SIZE = 5;
	defparam lut_1649.mask = 32'h05ff0800;

	lut_sub lut_1651 ({sk[627], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n859}, x6405x);
	defparam lut_1651.LUT_SIZE = 7;
	defparam lut_1651.mask = 128'h77ff7fff77ff7fff0000000080000000;

	lut_sub lut_1653 ({sk[628], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_5_, n_n852, n_n853}, x6412x);
	defparam lut_1653.LUT_SIZE = 7;
	defparam lut_1653.mask = 128'h77ff7fff77ff7fff0800000000000000;

	lut_sub lut_1655 ({sk[629], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n856}, x6433x);
	defparam lut_1655.LUT_SIZE = 7;
	defparam lut_1655.mask = 128'h77ff7fff77ff7fff0000000000020000;

	lut_sub lut_1657 ({sk[630], s298_in_0_, s298_in_2_, n_n857}, x6439x);
	defparam lut_1657.LUT_SIZE = 4;
	defparam lut_1657.mask = 16'h3f80;

	lut_sub lut_1659 ({sk[631], s298_in_1_, n_n852, n_n853, n_n854}, x6440x);
	defparam lut_1659.LUT_SIZE = 5;
	defparam lut_1659.mask = 32'h05ff0080;

	lut_sub lut_1661 ({sk[632], s298_in_0_, s298_in_2_, n_n857}, x6446x);
	defparam lut_1661.LUT_SIZE = 4;
	defparam lut_1661.mask = 16'h3f08;

	lut_sub lut_1663 ({sk[633], s298_in_1_, n_n852, n_n853, n_n856}, x6447x);
	defparam lut_1663.LUT_SIZE = 5;
	defparam lut_1663.mask = 32'h05ff0020;

	lut_sub lut_1665 ({sk[634], s298_in_0_, s298_in_2_, s298_in_1_, n_n853}, x6454x);
	defparam lut_1665.LUT_SIZE = 5;
	defparam lut_1665.mask = 32'h05ff0080;

	lut_sub lut_1667 ({sk[635], n_n854, n_n855, n_n856, n_n857}, x6455x);
	defparam lut_1667.LUT_SIZE = 5;
	defparam lut_1667.mask = 32'h05ff0800;

	lut_sub lut_1669 ({sk[636], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6461x);
	defparam lut_1669.LUT_SIZE = 5;
	defparam lut_1669.mask = 32'h05ff0040;

	lut_sub lut_1671 ({sk[637], n_n853, n_n854, n_n856, n_n857}, x6462x);
	defparam lut_1671.LUT_SIZE = 5;
	defparam lut_1671.mask = 32'h05ff0002;

	lut_sub lut_1673 ({sk[638], s298_in_0_, s298_in_2_, n_n855}, x6467x);
	defparam lut_1673.LUT_SIZE = 4;
	defparam lut_1673.mask = 16'h3f40;

	lut_sub lut_1675 ({sk[639], s298_in_1_, n_n852, n_n853, n_n854}, x6468x);
	defparam lut_1675.LUT_SIZE = 5;
	defparam lut_1675.mask = 32'h05ff0010;

	lut_sub lut_1677 ({sk[640], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n854, n_n855}, x6475x);
	defparam lut_1677.LUT_SIZE = 7;
	defparam lut_1677.mask = 128'h77ff7fff77ff7fff0020000000000000;

	lut_sub lut_1679 ({sk[641], s298_in_1_, n_n853, n_n854, n_n855}, x6489x);
	defparam lut_1679.LUT_SIZE = 5;
	defparam lut_1679.mask = 32'h05ff4000;

	lut_sub lut_1681 ({sk[642], s298_in_0_, s298_in_2_, n_n856, n_n857, n_n858, n_n859}, x6490x);
	defparam lut_1681.LUT_SIZE = 7;
	defparam lut_1681.mask = 128'h77ff7fff77ff7fff0d0f000000000000;

	lut_sub lut_1685 ({sk[643], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6496x);
	defparam lut_1685.LUT_SIZE = 5;
	defparam lut_1685.mask = 32'h05ff4000;

	lut_sub lut_1687 ({sk[644], n_n853, n_n855, n_n856, n_n859}, x6497x);
	defparam lut_1687.LUT_SIZE = 5;
	defparam lut_1687.mask = 32'h05ff0040;

	lut_sub lut_1689 ({sk[645], s298_in_1_, n_n852, n_n853, n_n854}, x6517x);
	defparam lut_1689.LUT_SIZE = 5;
	defparam lut_1689.mask = 32'h05ff0008;

	lut_sub lut_1691 ({sk[646], s298_in_0_, s298_in_2_, n_n855, x6517x}, x6518x);
	defparam lut_1691.LUT_SIZE = 5;
	defparam lut_1691.mask = 32'h05ff0040;

	lut_sub lut_1693 ({sk[647], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6552x);
	defparam lut_1693.LUT_SIZE = 5;
	defparam lut_1693.mask = 32'h05ff8000;

	lut_sub lut_1695 ({sk[648], n_n853, n_n855, n_n857, n_n859}, x6553x);
	defparam lut_1695.LUT_SIZE = 5;
	defparam lut_1695.mask = 32'h05ff2000;

	lut_sub lut_1697 ({sk[649], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6559x);
	defparam lut_1697.LUT_SIZE = 5;
	defparam lut_1697.mask = 32'h05ff0020;

	lut_sub lut_1699 ({sk[650], n_n853, n_n854, n_n855, n_n858}, x6560x);
	defparam lut_1699.LUT_SIZE = 5;
	defparam lut_1699.mask = 32'h05ff0004;

	lut_sub lut_1701 ({sk[651], s298_in_0_, s298_in_2_, n_n857}, x6607x);
	defparam lut_1701.LUT_SIZE = 4;
	defparam lut_1701.mask = 16'h3f40;

	lut_sub lut_1703 ({sk[652], s298_in_1_, n_n852, n_n853, n_n856}, x6608x);
	defparam lut_1703.LUT_SIZE = 5;
	defparam lut_1703.mask = 32'h05ff0008;

	lut_sub lut_1705 ({sk[653], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6615x);
	defparam lut_1705.LUT_SIZE = 5;
	defparam lut_1705.mask = 32'h05ff0040;

	lut_sub lut_1707 ({sk[654], n_n853, n_n854, n_n855, n_n856}, x6616x);
	defparam lut_1707.LUT_SIZE = 5;
	defparam lut_1707.mask = 32'h05ff4000;

	lut_sub lut_1709 ({sk[655], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x6636x);
	defparam lut_1709.LUT_SIZE = 5;
	defparam lut_1709.mask = 32'h05ff0080;

	lut_sub lut_1711 ({sk[656], n_n853, n_n854, n_n855, n_n856}, x6637x);
	defparam lut_1711.LUT_SIZE = 5;
	defparam lut_1711.mask = 32'h05ff0080;

	lut_sub lut_1713 ({sk[657], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n859}, x6706x);
	defparam lut_1713.LUT_SIZE = 7;
	defparam lut_1713.mask = 128'h77ff7fff77ff7fff0002000000000000;

	lut_sub lut_1715 ({sk[658], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n855, n_n856}, x6712x);
	defparam lut_1715.LUT_SIZE = 7;
	defparam lut_1715.mask = 128'h77ff7fff77ff7fff0008000000000000;

	lut_sub lut_1717 ({sk[659], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_0_, n_n852, n_n854}, x6718x);
	defparam lut_1717.LUT_SIZE = 7;
	defparam lut_1717.mask = 128'h77ff7fff77ff7fff0000000008000000;

	lut_sub lut_1719 ({sk[660], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_4_, n_n852, n_n853}, x6724x);
	defparam lut_1719.LUT_SIZE = 7;
	defparam lut_1719.mask = 128'h77ff7fff77ff7fff0004000000000000;

	lut_sub lut_1721 ({sk[661], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_4_, n_n852, n_n855}, x6730x);
	defparam lut_1721.LUT_SIZE = 7;
	defparam lut_1721.mask = 128'h77ff7fff77ff7fff1000000000000000;

	lut_sub lut_1723 ({sk[662], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_4_, n_n854, n_n857}, x6736x);
	defparam lut_1723.LUT_SIZE = 7;
	defparam lut_1723.mask = 128'h77ff7fff77ff7fff0000000000100000;

	lut_sub lut_1725 ({sk[663], s298_in_2_, s298_in_1_, n_n852, n_n853, n_n854, n_n856}, x6742x);
	defparam lut_1725.LUT_SIZE = 7;
	defparam lut_1725.mask = 128'h77ff7fff77ff7fff1000000000000000;

	lut_sub lut_1727 ({sk[664], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n857}, x6748x);
	defparam lut_1727.LUT_SIZE = 7;
	defparam lut_1727.mask = 128'h77ff7fff77ff7fff2000000000000000;

	lut_sub lut_1729 ({sk[665], s298_in_0_, s298_in_2_, n_n858}, x6753x);
	defparam lut_1729.LUT_SIZE = 4;
	defparam lut_1729.mask = 16'h3f08;

	lut_sub lut_1731 ({sk[666], s298_in_1_, n_n852, n_n854, n_n856}, x6754x);
	defparam lut_1731.LUT_SIZE = 5;
	defparam lut_1731.mask = 32'h05ff4000;

	lut_sub lut_1733 ({sk[667], s298_in_0_, s298_in_2_, n_n856}, x6759x);
	defparam lut_1733.LUT_SIZE = 4;
	defparam lut_1733.mask = 16'h3f08;

	lut_sub lut_1735 ({sk[668], s298_in_1_, n_n852, n_n853, n_n854}, x6760x);
	defparam lut_1735.LUT_SIZE = 5;
	defparam lut_1735.mask = 32'h05ff0001;

	lut_sub lut_1737 ({sk[669], s298_in_0_, s298_in_1_, s298_out_5_, n_n853, n_n855, n_n856}, x6766x);
	defparam lut_1737.LUT_SIZE = 7;
	defparam lut_1737.mask = 128'h77ff7fff77ff7fff0000000000040000;

	lut_sub lut_1739 ({sk[670], s298_in_1_, n_n852, n_n853, n_n854, n_n855, n_n51}, x6772x);
	defparam lut_1739.LUT_SIZE = 7;
	defparam lut_1739.mask = 128'h77ff7fff77ff7fff0010000000000000;

	lut_sub lut_1741 ({sk[671], s298_in_1_, n_n852, n_n857}, x6777x);
	defparam lut_1741.LUT_SIZE = 4;
	defparam lut_1741.mask = 16'h3f02;

	lut_sub lut_1743 ({sk[672], n_n853, n_n854, n_n855, n_n856}, x6778x);
	defparam lut_1743.LUT_SIZE = 5;
	defparam lut_1743.mask = 32'h05ff1000;

	lut_sub lut_1745 ({sk[673], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n855, n_n856}, x6784x);
	defparam lut_1745.LUT_SIZE = 7;
	defparam lut_1745.mask = 128'h77ff7fff77ff7fff0000000000400000;

	lut_sub lut_1747 ({sk[674], s298_in_2_, s298_in_1_, s298_out_0_, n_n852, n_n854, n_n855}, x6790x);
	defparam lut_1747.LUT_SIZE = 7;
	defparam lut_1747.mask = 128'h77ff7fff77ff7fff0000002000000000;

	lut_sub lut_1749 ({sk[675], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n855, n_n856}, x6796x);
	defparam lut_1749.LUT_SIZE = 7;
	defparam lut_1749.mask = 128'h77ff7fff77ff7fff0004000000000000;

	lut_sub lut_1751 ({sk[676], s298_in_0_, s298_in_2_, s298_in_1_, n_n854, n_n855, n_n856}, x6802x);
	defparam lut_1751.LUT_SIZE = 7;
	defparam lut_1751.mask = 128'h77ff7fff77ff7fff0000000000400000;

	lut_sub lut_1753 ({sk[677], s298_in_2_, s298_in_1_, n_n853, n_n854, n_n855, n_n856}, x6808x);
	defparam lut_1753.LUT_SIZE = 7;
	defparam lut_1753.mask = 128'h77ff7fff77ff7fff0000002000000000;

	lut_sub lut_1755 ({sk[678], n_n852, n_n854, n_n855, n_n857}, x6814x);
	defparam lut_1755.LUT_SIZE = 5;
	defparam lut_1755.mask = 32'h05ff0002;

	lut_sub lut_1757 ({sk[679], s298_in_1_, n_n852, n_n855, n_n857}, x6826x);
	defparam lut_1757.LUT_SIZE = 5;
	defparam lut_1757.mask = 32'h05ff0040;

	lut_sub lut_1759 ({sk[680], s298_in_1_, n_n853, n_n854, n_n855}, x6838x);
	defparam lut_1759.LUT_SIZE = 5;
	defparam lut_1759.mask = 32'h05ff0400;

	lut_sub lut_1761 ({sk[681], s298_in_1_, n_n852, n_n854, n_n855}, x6844x);
	defparam lut_1761.LUT_SIZE = 5;
	defparam lut_1761.mask = 32'h05ff0010;

	lut_sub lut_1763 ({sk[682], s298_in_1_, n_n852, n_n854, n_n856}, x6862x);
	defparam lut_1763.LUT_SIZE = 5;
	defparam lut_1763.mask = 32'h05ff0040;

	lut_sub lut_1765 ({sk[683], s298_in_0_, s298_in_2_, n_n853, n_n854, n_n855, n_n857}, x6868x);
	defparam lut_1765.LUT_SIZE = 7;
	defparam lut_1765.mask = 128'h77ff7fff77ff7fff1000000000000000;

	lut_sub lut_1767 ({sk[684], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n854, n_n859}, x6886x);
	defparam lut_1767.LUT_SIZE = 7;
	defparam lut_1767.mask = 128'h77ff7fff77ff7fff0200000000000000;

	lut_sub lut_1769 ({sk[685], s298_in_0_, s298_in_2_, n_n857}, x6903x);
	defparam lut_1769.LUT_SIZE = 4;
	defparam lut_1769.mask = 16'h3f40;

	lut_sub lut_1771 ({sk[686], s298_in_1_, n_n854, n_n855, n_n856}, x6904x);
	defparam lut_1771.LUT_SIZE = 5;
	defparam lut_1771.mask = 32'h05ff0002;

	lut_sub lut_1773 ({sk[687], n_n853, n_n854, n_n856, n_n859, x6910x, x6916x}, x7116x);
	defparam lut_1773.LUT_SIZE = 7;
	defparam lut_1773.mask = 128'h77ff7fff77ff7fff0000005000300000;

	lut_sub lut_1776 ({sk[688], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, x6923x, x6929x}, x7117x);
	defparam lut_1776.LUT_SIZE = 7;
	defparam lut_1776.mask = 128'h77ff7fff77ff7fff0530000000000000;

	lut_sub lut_1779 ({sk[689], n_n854, n_n856, n_n857, n_n859, x6934x, x409x}, x7118x);
	defparam lut_1779.LUT_SIZE = 7;
	defparam lut_1779.mask = 128'h77ff7fff77ff7fff5557555555555555;

	lut_sub lut_1782 ({sk[690], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, x6947x, x6953x}, x7119x);
	defparam lut_1782.LUT_SIZE = 7;
	defparam lut_1782.mask = 128'h77ff7fff77ff7fff0300000005000000;

	lut_sub lut_1785 ({sk[691], s298_in_0_, s298_in_2_, n_n859, x6958x, x6959x, x7084x}, x7120x);
	defparam lut_1785.LUT_SIZE = 7;
	defparam lut_1785.mask = 128'h77ff7fff77ff7fff0303030357030303;

	lut_sub lut_1788 ({sk[692], s298_in_1_, n_n852, n_n853, n_n855, x6645x, x362x}, x7121x);
	defparam lut_1788.LUT_SIZE = 7;
	defparam lut_1788.mask = 128'h77ff7fff77ff7fff5555555755555555;

	lut_sub lut_1791 ({sk[693], s298_in_1_, n_n852, n_n853, n_n855, x6659x, x364x}, x7122x);
	defparam lut_1791.LUT_SIZE = 7;
	defparam lut_1791.mask = 128'h77ff7fff77ff7fff5575555555555555;

	lut_sub lut_1794 ({sk[694], s298_in_0_, s298_in_2_, n_n855, n_n856, n_n857, n_n858}, x12833x);
	defparam lut_1794.LUT_SIZE = 7;
	defparam lut_1794.mask = 128'h77ff7fff77ff7fffff3fffffff5fffff;

	lut_sub lut_1801 ({sk[695], s298_in_1_, n_n852, n_n853, n_n854, x12833x}, x7123x);
	defparam lut_1801.LUT_SIZE = 6;
	defparam lut_1801.mask = 64'h337f337f20000000;

	lut_sub lut_1803 ({sk[696], s298_in_1_, n_n852, n_n853, n_n854, x6687x, x368x}, x7124x);
	defparam lut_1803.LUT_SIZE = 7;
	defparam lut_1803.mask = 128'h77ff7fff77ff7fff5557555555555555;

	lut_sub lut_1806 ({sk[697], s298_in_1_, n_n852, n_n853, n_n855, x6701x, x7116x}, x7125x);
	defparam lut_1806.LUT_SIZE = 7;
	defparam lut_1806.mask = 128'h77ff7fff77ff7fff5555555555555755;

	lut_sub lut_1809 ({sk[698], s298_in_0_, s298_in_2_, s298_out_5_, n_n859, x6596x, x6862x}, x7128x);
	defparam lut_1809.LUT_SIZE = 7;
	defparam lut_1809.mask = 128'h77ff7fff77ff7fff7300330033003300;

	lut_sub lut_1812 ({sk[699], x7121x, x7122x, x7123x, x7124x}, x7133x);
	defparam lut_1812.LUT_SIZE = 5;
	defparam lut_1812.mask = 32'h05ff7fff;

	lut_sub lut_1817 ({sk[700], s298_out_4_, x6552x, x6553x, x6559x, x6560x}, x7135x);
	defparam lut_1817.LUT_SIZE = 6;
	defparam lut_1817.mask = 64'h337f337f111f0000;

	lut_sub lut_1820 ({sk[701], s298_in_0_, s298_in_2_, s298_out_4_, n_n856, x6838x, x6844x}, x7137x);
	defparam lut_1820.LUT_SIZE = 7;
	defparam lut_1820.mask = 128'h77ff7fff77ff7fff0003000000500000;

	lut_sub lut_1823 ({sk[702], s298_out_4_, x7064x, x7069x}, x7139x);
	defparam lut_1823.LUT_SIZE = 4;
	defparam lut_1823.mask = 16'h3f07;

	lut_sub lut_1826 ({sk[703], s298_out_1_, x6454x, x6455x, x6461x, x6462x}, x7141x);
	defparam lut_1826.LUT_SIZE = 6;
	defparam lut_1826.mask = 64'h337f337f111f0000;

	lut_sub lut_1829 ({sk[704], s298_out_1_, s298_out_2_, x7029x, x6903x, x6904x}, x7143x);
	defparam lut_1829.LUT_SIZE = 6;
	defparam lut_1829.mask = 64'h337f337f11001f0f;

	lut_sub lut_1832 ({sk[705], x347x, x7117x, x7118x, x7125x, x7135x}, x7145x);
	defparam lut_1832.LUT_SIZE = 6;
	defparam lut_1832.mask = 64'h337f337f7fffffff;

	lut_sub lut_1838 ({sk[706], n_n51, x6400x, x7119x, x7120x, x7128x, x7133x}, x7148x);
	defparam lut_1838.LUT_SIZE = 7;
	defparam lut_1838.mask = 128'h77ff7fff77ff7fff7fff7fff7fffffff;

	lut_sub lut_1844 ({sk[707], s298_out_2_, n_n51, x6607x, x6608x, x6615x, x6616x}, x7149x);
	defparam lut_1844.LUT_SIZE = 7;
	defparam lut_1844.mask = 128'h77ff7fff77ff7fff0000111f00001111;

	lut_sub lut_1847 ({sk[708], s298_out_2_, x402x, x6636x, x6637x, x7143x}, x7152x);
	defparam lut_1847.LUT_SIZE = 6;
	defparam lut_1847.mask = 64'h337f337f55ff57ff;

	lut_sub lut_1851 ({sk[709], x350x, x352x, x394x, x395x, x7137x, x7139x}, x7154x);
	defparam lut_1851.LUT_SIZE = 7;
	defparam lut_1851.mask = 128'h77ff7fff77ff7fff7fffffffffffffff;

	lut_sub lut_1858 ({sk[710], s298_in_0_, s298_in_2_, s298_out_0_, n_n858, x6821x, x6826x}, x7156x);
	defparam lut_1858.LUT_SIZE = 7;
	defparam lut_1858.mask = 128'h77ff7fff77ff7fff3350330033003300;

	lut_sub lut_1861 ({sk[711], s298_out_1_, n_n51, x6624x, x7074x, x6784x, x7141x}, x7158x);
	defparam lut_1861.LUT_SIZE = 7;
	defparam lut_1861.mask = 128'h77ff7fff77ff7fff55557fff55555fff;

	lut_sub lut_1866 ({sk[712], s298_out_1_, x7034x, x442x, x7145x, x7152x}, x7159x);
	defparam lut_1866.LUT_SIZE = 6;
	defparam lut_1866.mask = 64'h337f337f7f7f7fff;

	lut_sub lut_1871 ({sk[713], s298_out_0_, n_n51, x345x, x6518x, x7154x}, x7160x);
	defparam lut_1871.LUT_SIZE = 6;
	defparam lut_1871.mask = 64'h337f337f5f5f7f5f;

	lut_sub lut_1875 ({sk[714], x7148x, x7149x, x7156x, x7158x, x7159x, x7160x}, x7164x);
	defparam lut_1875.LUT_SIZE = 7;
	defparam lut_1875.mask = 128'h77ff7fff77ff7fff7fffffffffffffff;

	lut_sub lut_1882 ({sk[715], x346x, x351x, x353x, x355x}, x7174x);
	defparam lut_1882.LUT_SIZE = 5;
	defparam lut_1882.mask = 32'h05ff7fff;

	lut_sub lut_1887 ({sk[716], n_n51, n_n52, x6631x, x391x, x398x, x6868x}, x7175x);
	defparam lut_1887.LUT_SIZE = 7;
	defparam lut_1887.mask = 128'h77ff7fff77ff7fff3fff3f3f3fff7f7f;

	lut_sub lut_1892 ({sk[717], s298_out_2_, n_n52, x6881x, x401x, x7024x, x6886x}, x7176x);
	defparam lut_1892.LUT_SIZE = 7;
	defparam lut_1892.mask = 128'h77ff7fff77ff7fff3fff0f0f3fff5f5f;

	lut_sub lut_1897 ({sk[718], n_n52, x6526x, x7059x, x7079x, x444x, x7164x}, x7177x);
	defparam lut_1897.LUT_SIZE = 7;
	defparam lut_1897.mask = 128'h77ff7fff77ff7fff777777777fffffff;

	lut_sub lut_1903 ({sk[719], s298_out_0_, n_n50, x6389x, x6390x, x6467x, x6468x}, x7181x);
	defparam lut_1903.LUT_SIZE = 7;
	defparam lut_1903.mask = 128'h77ff7fff77ff7fff111f000000000000;

	lut_sub lut_1906 ({sk[720], s298_out_0_, n_n50, n_n52, x6484x, x6475x}, x7182x);
	defparam lut_1906.LUT_SIZE = 6;
	defparam lut_1906.mask = 64'h337f337f33003700;

	lut_sub lut_1909 ({sk[721], n_n50, x6489x, x6490x, x6496x, x6497x}, x7183x);
	defparam lut_1909.LUT_SIZE = 6;
	defparam lut_1909.mask = 64'h337f337f111f0000;

	lut_sub lut_1912 ({sk[722], s298_out_0_, n_n50, n_n52, x6790x, x6796x}, x7185x);
	defparam lut_1912.LUT_SIZE = 6;
	defparam lut_1912.mask = 64'h337f337f03005700;

	lut_sub lut_1915 ({sk[723], s298_out_4_, n_n50, n_n52, x6802x, x6808x}, x7186x);
	defparam lut_1915.LUT_SIZE = 6;
	defparam lut_1915.mask = 64'h337f337f50007300;

	lut_sub lut_1918 ({sk[724], s298_in_2_, s298_in_1_, n_n50, n_n859, x7019x, x6814x}, x7187x);
	defparam lut_1918.LUT_SIZE = 7;
	defparam lut_1918.mask = 128'h77ff7fff77ff7fff3300370033003300;

	lut_sub lut_1921 ({sk[725], x6018x, x7039x, x7044x, x6016x, x6017x}, x7188x);
	defparam lut_1921.LUT_SIZE = 6;
	defparam lut_1921.mask = 64'h337f337f08880000;

	lut_sub lut_1924 ({sk[726], s298_in_1_, s298_out_0_, n_n852, n_n50, n_n858, x7108x}, x7190x);
	defparam lut_1924.LUT_SIZE = 7;
	defparam lut_1924.mask = 128'h77ff7fff77ff7fff0505050705050505;

	lut_sub lut_1927 ({sk[727], x7174x, x7175x, x7176x, x7177x, x7181x, x7190x}, x7196x);
	defparam lut_1927.LUT_SIZE = 7;
	defparam lut_1927.mask = 128'h77ff7fff77ff7fff7fffffffffffffff;

	lut_sub lut_1934 ({sk[728], n_n50, x6505x, x6512x, x7182x, x7183x, x7185x}, x7197x);
	defparam lut_1934.LUT_SIZE = 7;
	defparam lut_1934.mask = 128'h77ff7fff77ff7fff7f7fffff7fff7fff;

	lut_sub lut_1940 ({sk[729], n_n50, x7049x, x7054x, x7186x, x7187x, x7188x}, x7198x);
	defparam lut_1940.LUT_SIZE = 7;
	defparam lut_1940.mask = 128'h77ff7fff77ff7fff7f7f7f7f7fffffff;

	lut_sub lut_1946 ({sk[730], x7196x, x7197x, x7198x}, x7200x);
	defparam lut_1946.LUT_SIZE = 4;
	defparam lut_1946.mask = 16'h3f7f;

	lut_sub lut_1950 ({sk[731], s298_out_5_, n_n49, n_n50, n_n52, x6405x, x6412x}, x7202x);
	defparam lut_1950.LUT_SIZE = 7;
	defparam lut_1950.mask = 128'h77ff7fff77ff7fff7300000050000000;

	lut_sub lut_1953 ({sk[732], s298_out_4_, n_n49, n_n52, x6433x, x6439x, x6440x}, x7204x);
	defparam lut_1953.LUT_SIZE = 7;
	defparam lut_1953.mask = 128'h77ff7fff77ff7fff001100000f110000;

	lut_sub lut_1956 ({sk[733], s298_out_1_, n_n49, n_n52, x6446x, x6447x, x6706x}, x7205x);
	defparam lut_1956.LUT_SIZE = 7;
	defparam lut_1956.mask = 128'h77ff7fff77ff7fff5557000000030000;

	lut_sub lut_1959 ({sk[734], s298_out_1_, n_n49, n_n50, x6712x, x6718x}, x7206x);
	defparam lut_1959.LUT_SIZE = 6;
	defparam lut_1959.mask = 64'h337f337f50007300;

	lut_sub lut_1962 ({sk[735], n_n49, n_n50, n_n51, x6724x, x6730x}, x7207x);
	defparam lut_1962.LUT_SIZE = 6;
	defparam lut_1962.mask = 64'h337f337f73500000;

	lut_sub lut_1965 ({sk[736], s298_out_4_, n_n49, n_n52, x6736x, x6742x}, x7208x);
	defparam lut_1965.LUT_SIZE = 6;
	defparam lut_1965.mask = 64'h337f337f03005700;

	lut_sub lut_1968 ({sk[737], n_n49, n_n52, x6748x, x6753x, x6754x}, x7209x);
	defparam lut_1968.LUT_SIZE = 6;
	defparam lut_1968.mask = 64'h337f337f111f0000;

	lut_sub lut_1971 ({sk[738], n_n49, n_n51, x6759x, x6760x, x6766x}, x7210x);
	defparam lut_1971.LUT_SIZE = 6;
	defparam lut_1971.mask = 64'h337f337f03035500;

	lut_sub lut_1974 ({sk[739], n_n49, n_n52, x6772x, x6777x, x6778x}, x7211x);
	defparam lut_1974.LUT_SIZE = 6;
	defparam lut_1974.mask = 64'h337f337f0000111f;

	lut_sub lut_1977 ({sk[740], n_n49, x6964x, x6969x}, x7212x);
	defparam lut_1977.LUT_SIZE = 4;
	defparam lut_1977.mask = 16'h3f70;

	lut_sub lut_1980 ({sk[741], n_n49, x6984x, x6989x, x6994x, x6999x}, x12832x);
	defparam lut_1980.LUT_SIZE = 6;
	defparam lut_1980.mask = 64'h337f337fffff8000;

	lut_sub lut_1983 ({sk[742], s298_in_0_, s298_in_2_, s298_out_3_, n_n853, n_n854, n_n855}, x7248x);
	defparam lut_1983.LUT_SIZE = 7;
	defparam lut_1983.mask = 128'h77ff7fff77ff7fff0000000040000000;

	lut_sub lut_1985 ({sk[743], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n855, n_n856}, x7262x);
	defparam lut_1985.LUT_SIZE = 7;
	defparam lut_1985.mask = 128'h77ff7fff77ff7fff0200000000000000;

	lut_sub lut_1987 ({sk[744], s298_in_0_, s298_in_1_, n_n858}, x7268x);
	defparam lut_1987.LUT_SIZE = 4;
	defparam lut_1987.mask = 16'h3f20;

	lut_sub lut_1989 ({sk[745], n_n852, n_n853, n_n854, n_n857}, x7269x);
	defparam lut_1989.LUT_SIZE = 5;
	defparam lut_1989.mask = 32'h05ff0001;

	lut_sub lut_1991 ({sk[746], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7290x);
	defparam lut_1991.LUT_SIZE = 5;
	defparam lut_1991.mask = 32'h05ff4000;

	lut_sub lut_1993 ({sk[747], n_n853, n_n854, n_n855, n_n856}, x7291x);
	defparam lut_1993.LUT_SIZE = 5;
	defparam lut_1993.mask = 32'h05ff0020;

	lut_sub lut_1995 ({sk[748], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7297x);
	defparam lut_1995.LUT_SIZE = 5;
	defparam lut_1995.mask = 32'h05ff0080;

	lut_sub lut_1997 ({sk[749], n_n853, n_n854, n_n855, n_n857}, x7298x);
	defparam lut_1997.LUT_SIZE = 5;
	defparam lut_1997.mask = 32'h05ff0001;

	lut_sub lut_1999 ({sk[750], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x7388x);
	defparam lut_1999.LUT_SIZE = 5;
	defparam lut_1999.mask = 32'h05ff1000;

	lut_sub lut_2001 ({sk[751], s298_in_0_, s298_in_2_, s298_out_1_, n_n852, n_n853, n_n855}, x7423x);
	defparam lut_2001.LUT_SIZE = 7;
	defparam lut_2001.mask = 128'h77ff7fff77ff7fff0000000000400000;

	lut_sub lut_2003 ({sk[752], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n856, n_n859}, x7429x);
	defparam lut_2003.LUT_SIZE = 7;
	defparam lut_2003.mask = 128'h77ff7fff77ff7fff0200000000000000;

	lut_sub lut_2005 ({sk[753], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n856}, x7435x);
	defparam lut_2005.LUT_SIZE = 7;
	defparam lut_2005.mask = 128'h77ff7fff77ff7fff0008000000000000;

	lut_sub lut_2007 ({sk[754], s298_in_2_, s298_in_1_, n_n852, n_n854, n_n855, n_n857}, x7441x);
	defparam lut_2007.LUT_SIZE = 7;
	defparam lut_2007.mask = 128'h77ff7fff77ff7fff0000200000000000;

	lut_sub lut_2009 ({sk[755], s298_in_2_, s298_in_1_, n_n852, n_n853, n_n856, n_n857}, x7447x);
	defparam lut_2009.LUT_SIZE = 7;
	defparam lut_2009.mask = 128'h77ff7fff77ff7fff0000800000000000;

	lut_sub lut_2011 ({sk[756], n_n853, n_n854, n_n855, n_n856}, x7453x);
	defparam lut_2011.LUT_SIZE = 5;
	defparam lut_2011.mask = 32'h05ff0040;

	lut_sub lut_2013 ({sk[757], n_n853, n_n854, n_n855, n_n858}, x7459x);
	defparam lut_2013.LUT_SIZE = 5;
	defparam lut_2013.mask = 32'h05ff0004;

	lut_sub lut_2015 ({sk[758], s298_in_1_, n_n852, n_n854, n_n855}, x7465x);
	defparam lut_2015.LUT_SIZE = 5;
	defparam lut_2015.mask = 32'h05ff0080;

	lut_sub lut_2017 ({sk[759], s298_in_1_, n_n853, n_n854, n_n855}, x7471x);
	defparam lut_2017.LUT_SIZE = 5;
	defparam lut_2017.mask = 32'h05ff0400;

	lut_sub lut_2019 ({sk[760], s298_in_0_, s298_in_2_, n_n858}, x7476x);
	defparam lut_2019.LUT_SIZE = 4;
	defparam lut_2019.mask = 16'h3f04;

	lut_sub lut_2021 ({sk[761], s298_in_1_, n_n852, n_n853, n_n856}, x7477x);
	defparam lut_2021.LUT_SIZE = 5;
	defparam lut_2021.mask = 32'h05ff4000;

	lut_sub lut_2023 ({sk[762], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n855, n_n52}, x7483x);
	defparam lut_2023.LUT_SIZE = 7;
	defparam lut_2023.mask = 128'h77ff7fff77ff7fff0100000000000000;

	lut_sub lut_2025 ({sk[763], n_n853, n_n854, n_n855, n_n856}, x7489x);
	defparam lut_2025.LUT_SIZE = 5;
	defparam lut_2025.mask = 32'h05ff1000;

	lut_sub lut_2027 ({sk[764], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n854}, x7495x);
	defparam lut_2027.LUT_SIZE = 7;
	defparam lut_2027.mask = 128'h77ff7fff77ff7fff0020000000000000;

	lut_sub lut_2029 ({sk[765], s298_in_0_, s298_in_2_, n_n856}, x7500x);
	defparam lut_2029.LUT_SIZE = 4;
	defparam lut_2029.mask = 16'h3f08;

	lut_sub lut_2031 ({sk[766], s298_in_1_, n_n852, n_n853, n_n855}, x7501x);
	defparam lut_2031.LUT_SIZE = 5;
	defparam lut_2031.mask = 32'h05ff0004;

	lut_sub lut_2033 ({sk[767], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n855, n_n856}, x7507x);
	defparam lut_2033.LUT_SIZE = 7;
	defparam lut_2033.mask = 128'h77ff7fff77ff7fff0010000000000000;

	lut_sub lut_2035 ({sk[768], s298_in_2_, s298_in_1_, n_n858}, x7512x);
	defparam lut_2035.LUT_SIZE = 4;
	defparam lut_2035.mask = 16'h3f80;

	lut_sub lut_2037 ({sk[769], n_n852, n_n854, n_n855, n_n856}, x7513x);
	defparam lut_2037.LUT_SIZE = 5;
	defparam lut_2037.mask = 32'h05ff1000;

	lut_sub lut_2039 ({sk[770], s298_in_2_, s298_in_1_, n_n858}, x7518x);
	defparam lut_2039.LUT_SIZE = 4;
	defparam lut_2039.mask = 16'h3f80;

	lut_sub lut_2041 ({sk[771], n_n852, n_n854, n_n855, n_n856}, x7519x);
	defparam lut_2041.LUT_SIZE = 5;
	defparam lut_2041.mask = 32'h05ff0004;

	lut_sub lut_2043 ({sk[772], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_3_, n_n852, n_n856}, x7525x);
	defparam lut_2043.LUT_SIZE = 7;
	defparam lut_2043.mask = 128'h77ff7fff77ff7fff0000000020000000;

	lut_sub lut_2045 ({sk[773], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_2_, n_n852, n_n853}, x7531x);
	defparam lut_2045.LUT_SIZE = 7;
	defparam lut_2045.mask = 128'h77ff7fff77ff7fff0008000000000000;

	lut_sub lut_2047 ({sk[774], s298_in_0_, s298_in_1_, n_n859}, x7536x);
	defparam lut_2047.LUT_SIZE = 4;
	defparam lut_2047.mask = 16'h3f01;

	lut_sub lut_2049 ({sk[775], n_n852, n_n853, n_n854, n_n858}, x7537x);
	defparam lut_2049.LUT_SIZE = 5;
	defparam lut_2049.mask = 32'h05ff0400;

	lut_sub lut_2051 ({sk[776], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n854, n_n857}, x7543x);
	defparam lut_2051.LUT_SIZE = 7;
	defparam lut_2051.mask = 128'h77ff7fff77ff7fff0100000000000000;

	lut_sub lut_2053 ({sk[777], s298_in_0_, s298_in_2_, n_n852, n_n853, n_n855, n_n858}, x7561x);
	defparam lut_2053.LUT_SIZE = 7;
	defparam lut_2053.mask = 128'h77ff7fff77ff7fff0000000000080000;

	lut_sub lut_2055 ({sk[778], s298_in_1_, n_n852, n_n853, n_n854}, x7573x);
	defparam lut_2055.LUT_SIZE = 5;
	defparam lut_2055.mask = 32'h05ff4000;

	lut_sub lut_2057 ({sk[779], n_n852, n_n853, n_n854, n_n855}, x7579x);
	defparam lut_2057.LUT_SIZE = 5;
	defparam lut_2057.mask = 32'h05ff0010;

	lut_sub lut_2059 ({sk[780], s298_in_1_, n_n853, n_n854, n_n856}, x7585x);
	defparam lut_2059.LUT_SIZE = 5;
	defparam lut_2059.mask = 32'h05ff0020;

	lut_sub lut_2061 ({sk[781], s298_in_2_, s298_in_1_, n_n852, n_n854, n_n855, n_n856}, x7603x);
	defparam lut_2061.LUT_SIZE = 7;
	defparam lut_2061.mask = 128'h77ff7fff77ff7fff8000000000000000;

	lut_sub lut_2063 ({sk[782], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n853, n_n855}, x7633x);
	defparam lut_2063.LUT_SIZE = 7;
	defparam lut_2063.mask = 128'h77ff7fff77ff7fff0000000000100000;

	lut_sub lut_2065 ({sk[783], s298_in_2_, s298_in_1_, n_n852, n_n853, n_n854, n_n855}, x7651x);
	defparam lut_2065.LUT_SIZE = 7;
	defparam lut_2065.mask = 128'h77ff7fff77ff7fff0100000000000000;

	lut_sub lut_2067 ({sk[784], s298_in_0_, s298_in_2_, n_n856}, x7656x);
	defparam lut_2067.LUT_SIZE = 4;
	defparam lut_2067.mask = 16'h3f04;

	lut_sub lut_2069 ({sk[785], s298_in_1_, n_n852, n_n853, n_n854}, x7657x);
	defparam lut_2069.LUT_SIZE = 5;
	defparam lut_2069.mask = 32'h05ff4000;

	lut_sub lut_2071 ({sk[786], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n854, n_n857}, x7663x);
	defparam lut_2071.LUT_SIZE = 7;
	defparam lut_2071.mask = 128'h77ff7fff77ff7fff1000000000000000;

	lut_sub lut_2073 ({sk[787], n_n854, n_n857, n_n858, n_n859, x7693x, x281x}, x7895x);
	defparam lut_2073.LUT_SIZE = 7;
	defparam lut_2073.mask = 128'h77ff7fff77ff7fff5555755555555555;

	lut_sub lut_2076 ({sk[788], n_n854, n_n856, n_n858, n_n859, x7705x, x283x}, x7896x);
	defparam lut_2076.LUT_SIZE = 7;
	defparam lut_2076.mask = 128'h77ff7fff77ff7fff5555555555555575;

	lut_sub lut_2079 ({sk[789], n_n853, n_n854, n_n855, n_n856, n_n857}, x12828x);
	defparam lut_2079.LUT_SIZE = 6;
	defparam lut_2079.mask = 64'h337f337fffff7c7f;

	lut_sub lut_2088 ({sk[790], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, x12828x}, x7897x);
	defparam lut_2088.LUT_SIZE = 6;
	defparam lut_2088.mask = 64'h337f337f00000200;

	lut_sub lut_2090 ({sk[791], s298_out_3_, x7389x, x7396x, x7397x, x7388x}, x7898x);
	defparam lut_2090.LUT_SIZE = 6;
	defparam lut_2090.mask = 64'h337f337f03570303;

	lut_sub lut_2093 ({sk[792], s298_in_1_, n_n853, n_n854, n_n855, x7404x, x233x}, x7899x);
	defparam lut_2093.LUT_SIZE = 7;
	defparam lut_2093.mask = 128'h77ff7fff77ff7fff5557555555555555;

	lut_sub lut_2096 ({sk[793], s298_in_1_, n_n852, n_n853, n_n854, x7418x, x279x}, x7900x);
	defparam lut_2096.LUT_SIZE = 7;
	defparam lut_2096.mask = 128'h77ff7fff77ff7fff5555555557555555;

	lut_sub lut_2099 ({sk[794], x209x, x269x, x271x, x272x, x7897x}, x7910x);
	defparam lut_2099.LUT_SIZE = 6;
	defparam lut_2099.mask = 64'h337f337f7fffffff;

	lut_sub lut_2105 ({sk[795], x214x, x7895x, x7896x, x7898x, x7899x, x7900x}, x7911x);
	defparam lut_2105.LUT_SIZE = 7;
	defparam lut_2105.mask = 128'h77ff7fff77ff7fff7fffffffffffffff;

	lut_sub lut_2112 ({sk[796], s298_out_1_, s298_out_5_, x7495x, x7500x, x7501x}, x7912x);
	defparam lut_2112.LUT_SIZE = 6;
	defparam lut_2112.mask = 64'h337f337f0000111f;

	lut_sub lut_2115 ({sk[797], s298_out_2_, n_n51, x7656x, x7657x, x7663x}, x7916x);
	defparam lut_2115.LUT_SIZE = 6;
	defparam lut_2115.mask = 64'h337f337f03550300;

	lut_sub lut_2118 ({sk[798], x218x, x222x, x223x, x264x, x268x}, x7920x);
	defparam lut_2118.LUT_SIZE = 6;
	defparam lut_2118.mask = 64'h337f337f7fffffff;

	lut_sub lut_2124 ({sk[799], s298_in_0_, s298_in_2_, s298_out_0_, n_n856, x7573x, x7579x}, x7925x);
	defparam lut_2124.LUT_SIZE = 7;
	defparam lut_2124.mask = 128'h77ff7fff77ff7fff0030000000050000;

	lut_sub lut_2127 ({sk[800], s298_in_0_, s298_in_2_, s298_out_0_, n_n857, x263x, x7585x}, x7926x);
	defparam lut_2127.LUT_SIZE = 7;
	defparam lut_2127.mask = 128'h77ff7fff77ff7fff3333333333733333;

	lut_sub lut_2130 ({sk[801], s298_out_0_, n_n51, x7355x, x7844x, x7910x}, x7927x);
	defparam lut_2130.LUT_SIZE = 6;
	defparam lut_2130.mask = 64'h337f337f5f557f77;

	lut_sub lut_2134 ({sk[802], s298_out_5_, n_n51, x7633x, x7651x, x7916x}, x7928x);
	defparam lut_2134.LUT_SIZE = 6;
	defparam lut_2134.mask = 64'h337f337f555f5577;

	lut_sub lut_2138 ({sk[803], s298_in_0_, s298_in_2_, n_n859, x12842x}, x12827x);
	defparam lut_2138.LUT_SIZE = 5;
	defparam lut_2138.mask = 32'h05ffff7f;

	lut_sub lut_2143 ({sk[804], n_n51, x7849x, x7881x, x12827x}, x7929x);
	defparam lut_2143.LUT_SIZE = 5;
	defparam lut_2143.mask = 32'h05ff33af;

	lut_sub lut_2147 ({sk[805], s298_out_0_, n_n51, x219x, x220x, x7327x, x7543x}, x7931x);
	defparam lut_2147.LUT_SIZE = 7;
	defparam lut_2147.mask = 128'h77ff7fff77ff7fff5fff0fff3fff3fff;

	lut_sub lut_2152 ({sk[806], s298_out_0_, n_n51, x7550x, x257x, x259x, x7561x}, x7932x);
	defparam lut_2152.LUT_SIZE = 7;
	defparam lut_2152.mask = 128'h77ff7fff77ff7fff3fff3fff3f3f7f7f;

	lut_sub lut_2157 ({sk[807], x7925x, x7926x, x7927x, x7928x}, x7937x);
	defparam lut_2157.LUT_SIZE = 5;
	defparam lut_2157.mask = 32'h05ff7fff;

	lut_sub lut_2162 ({sk[808], x7911x, x7912x, x7920x, x7929x, x7931x, x7932x}, x7938x);
	defparam lut_2162.LUT_SIZE = 7;
	defparam lut_2162.mask = 128'h77ff7fff77ff7fff7fffffffffffffff;

	lut_sub lut_2169 ({sk[809], x224x, x226x, x7937x, x7938x}, x7945x);
	defparam lut_2169.LUT_SIZE = 5;
	defparam lut_2169.mask = 32'h05ff7fff;

	lut_sub lut_2174 ({sk[810], s298_out_4_, n_n52, x7369x, x228x, x229x, x7603x}, x7946x);
	defparam lut_2174.LUT_SIZE = 7;
	defparam lut_2174.mask = 128'h77ff7fff77ff7fff3f3f3fff7f7f3fff;

	lut_sub lut_2179 ({sk[811], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n854, n_n856}, x12826x);
	defparam lut_2179.LUT_SIZE = 7;
	defparam lut_2179.mask = 128'h77ff7fff77ff7fffffffffffdffdffff;

	lut_sub lut_2186 ({sk[812], s298_out_4_, n_n52, x278x, x7839x, x12826x}, x7947x);
	defparam lut_2186.LUT_SIZE = 6;
	defparam lut_2186.mask = 64'h337f337f0f3faf3f;

	lut_sub lut_2190 ({sk[813], n_n50, x7290x, x7291x, x7297x, x7298x}, x7951x);
	defparam lut_2190.LUT_SIZE = 6;
	defparam lut_2190.mask = 64'h337f337f0000111f;

	lut_sub lut_2193 ({sk[814], s298_out_4_, n_n50, x7507x, x7512x, x7513x}, x7952x);
	defparam lut_2193.LUT_SIZE = 6;
	defparam lut_2193.mask = 64'h337f337f11001f00;

	lut_sub lut_2196 ({sk[815], s298_out_5_, n_n50, x7518x, x7519x, x7525x}, x7953x);
	defparam lut_2196.LUT_SIZE = 6;
	defparam lut_2196.mask = 64'h337f337f03550300;

	lut_sub lut_2199 ({sk[816], n_n50, n_n52, x7531x, x7536x, x7537x}, x7954x);
	defparam lut_2199.LUT_SIZE = 6;
	defparam lut_2199.mask = 64'h337f337f00001f11;

	lut_sub lut_2202 ({sk[817], s298_in_1_, s298_out_4_, n_n854, n_n50, n_n857, x7834x}, x7957x);
	defparam lut_2202.LUT_SIZE = 7;
	defparam lut_2202.mask = 128'h77ff7fff77ff7fff0505050505050d05;

	lut_sub lut_2205 ({sk[818], n_n852, n_n50, n_n51, n_n859, x7890x}, x7958x);
	defparam lut_2205.LUT_SIZE = 6;
	defparam lut_2205.mask = 64'h337f337f005500d5;

	lut_sub lut_2208 ({sk[819], n_n50, x7814x, x7819x, x7952x, x7953x, x7954x}, x7964x);
	defparam lut_2208.LUT_SIZE = 7;
	defparam lut_2208.mask = 128'h77ff7fff77ff7fff7fffffff7f7f7f7f;

	lut_sub lut_2214 ({sk[820], n_n50, x7824x, x7829x, x7945x, x7946x, x7947x}, x12825x);
	defparam lut_2214.LUT_SIZE = 7;
	defparam lut_2214.mask = 128'h77ff7fff77ff7fff8080808080000000;

	lut_sub lut_2217 ({sk[821], x215x, x7951x, x7957x, x7958x, x12825x}, x7965x);
	defparam lut_2217.LUT_SIZE = 6;
	defparam lut_2217.mask = 64'h337f337fbfffffff;

	lut_sub lut_2223 ({sk[822], n_n49, n_n50, n_n51, x7248x, x7964x, x7965x}, x7967x);
	defparam lut_2223.LUT_SIZE = 7;
	defparam lut_2223.mask = 128'h77ff7fff77ff7fff7777777f77777777;

	lut_sub lut_2227 ({sk[823], n_n49, n_n51, n_n52, x7257x, x7262x}, x7968x);
	defparam lut_2227.LUT_SIZE = 6;
	defparam lut_2227.mask = 64'h337f337f73330000;

	lut_sub lut_2230 ({sk[824], n_n49, n_n51, x7268x, x7269x, x7423x}, x7969x);
	defparam lut_2230.LUT_SIZE = 6;
	defparam lut_2230.mask = 64'h337f337f00550003;

	lut_sub lut_2233 ({sk[825], s298_out_0_, n_n49, n_n50, x7429x, x7435x}, x7970x);
	defparam lut_2233.LUT_SIZE = 6;
	defparam lut_2233.mask = 64'h337f337f30007500;

	lut_sub lut_2236 ({sk[826], n_n49, n_n51, x7441x, x7447x}, x7971x);
	defparam lut_2236.LUT_SIZE = 5;
	defparam lut_2236.mask = 32'h05ff3500;

	lut_sub lut_2239 ({sk[827], s298_in_2_, s298_in_1_, n_n49, n_n859, x7453x, x7459x}, x7972x);
	defparam lut_2239.LUT_SIZE = 7;
	defparam lut_2239.mask = 128'h77ff7fff77ff7fff3500000000000000;

	lut_sub lut_2242 ({sk[828], n_n49, n_n50, x7476x, x7477x, x7483x}, x7974x);
	defparam lut_2242.LUT_SIZE = 6;
	defparam lut_2242.mask = 64'h337f337f03035500;

	lut_sub lut_2245 ({sk[829], s298_in_0_, s298_in_1_, n_n49, n_n857, x7729x, x7489x}, x7975x);
	defparam lut_2245.LUT_SIZE = 7;
	defparam lut_2245.mask = 128'h77ff7fff77ff7fff3300330533003300;

	lut_sub lut_2248 ({sk[830], n_n49, x7734x, x7739x}, x7976x);
	defparam lut_2248.LUT_SIZE = 4;
	defparam lut_2248.mask = 16'h3f70;

	lut_sub lut_2251 ({sk[831], s298_out_0_, n_n852, n_n49, n_n51, n_n859, x7877x}, x7987x);
	defparam lut_2251.LUT_SIZE = 7;
	defparam lut_2251.mask = 128'h77ff7fff77ff7fff00550055005d0055;

	lut_sub lut_2254 ({sk[832], s298_in_0_, s298_in_2_, n_n856, n_n858, x7465x, x7471x}, x12831x);
	defparam lut_2254.LUT_SIZE = 7;
	defparam lut_2254.mask = 128'h77ff7fff77ff7fffffaaffffcfcfffff;

	lut_sub lut_2264 ({sk[833], n_n49, x7754x, x7759x, x7764x, x7769x}, x12830x);
	defparam lut_2264.LUT_SIZE = 6;
	defparam lut_2264.mask = 64'h337f337fffff8000;

	lut_sub lut_2267 ({sk[834], n_n49, x7794x, x7799x, x7804x, x7809x}, x12829x);
	defparam lut_2267.LUT_SIZE = 6;
	defparam lut_2267.mask = 64'h337f337fffff8000;

	lut_sub lut_2270 ({sk[835], s298_out_0_, n_n49, n_n856, n_n51, x7869x, x7873x}, x12824x);
	defparam lut_2270.LUT_SIZE = 7;
	defparam lut_2270.mask = 128'h77ff7fff77ff7fffffff8888ffff8088;

	lut_sub lut_2275 ({sk[836], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n854, n_n855}, x8027x);
	defparam lut_2275.LUT_SIZE = 7;
	defparam lut_2275.mask = 128'h77ff7fff77ff7fff0000000000400000;

	lut_sub lut_2277 ({sk[837], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n854, n_n856}, x8034x);
	defparam lut_2277.LUT_SIZE = 7;
	defparam lut_2277.mask = 128'h77ff7fff77ff7fff0004000000000000;

	lut_sub lut_2279 ({sk[838], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x8048x);
	defparam lut_2279.LUT_SIZE = 5;
	defparam lut_2279.mask = 32'h05ff4000;

	lut_sub lut_2281 ({sk[839], n_n853, n_n854, n_n857, n_n858}, x8049x);
	defparam lut_2281.LUT_SIZE = 5;
	defparam lut_2281.mask = 32'h05ff0080;

	lut_sub lut_2283 ({sk[840], s298_in_0_, s298_in_2_, s298_in_1_, n_n852}, x8062x);
	defparam lut_2283.LUT_SIZE = 5;
	defparam lut_2283.mask = 32'h05ff0010;

	lut_sub lut_2285 ({sk[841], n_n853, n_n854, n_n855, n_n856}, x8063x);
	defparam lut_2285.LUT_SIZE = 5;
	defparam lut_2285.mask = 32'h05ff1000;

	lut_sub lut_2287 ({sk[842], s298_in_1_, n_n852, n_n853, n_n854}, x8069x);
	defparam lut_2287.LUT_SIZE = 5;
	defparam lut_2287.mask = 32'h05ff1000;

	lut_sub lut_2289 ({sk[843], s298_in_0_, s298_in_2_, n_n856, x8069x}, x8070x);
	defparam lut_2289.LUT_SIZE = 5;
	defparam lut_2289.mask = 32'h05ff0010;

	lut_sub lut_2291 ({sk[844], s298_in_1_, n_n853, n_n854, n_n855}, x8083x);
	defparam lut_2291.LUT_SIZE = 5;
	defparam lut_2291.mask = 32'h05ff8000;

	lut_sub lut_2293 ({sk[845], s298_in_0_, s298_in_2_, n_n856, x8083x}, x8084x);
	defparam lut_2293.LUT_SIZE = 5;
	defparam lut_2293.mask = 32'h05ff1000;

	lut_sub lut_2295 ({sk[846], s298_in_0_, s298_in_2_, n_n852, n_n855, n_n857, n_n859}, x8181x);
	defparam lut_2295.LUT_SIZE = 7;
	defparam lut_2295.mask = 128'h77ff7fff77ff7fff0000000004000000;

	lut_sub lut_2297 ({sk[847], s298_in_2_, s298_in_1_, n_n852, n_n854, n_n856, n_n858}, x8187x);
	defparam lut_2297.LUT_SIZE = 7;
	defparam lut_2297.mask = 128'h77ff7fff77ff7fff0000080000000000;

	lut_sub lut_2299 ({sk[848], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n854, n_n856}, x8193x);
	defparam lut_2299.LUT_SIZE = 7;
	defparam lut_2299.mask = 128'h77ff7fff77ff7fff0000000080000000;

	lut_sub lut_2301 ({sk[849], s298_in_0_, s298_in_1_, n_n853, n_n854, n_n855, n_n856}, x8199x);
	defparam lut_2301.LUT_SIZE = 7;
	defparam lut_2301.mask = 128'h77ff7fff77ff7fff0000000000000040;

	lut_sub lut_2303 ({sk[850], s298_in_0_, s298_out_5_, n_n852, n_n853, n_n856, n_n857}, x8205x);
	defparam lut_2303.LUT_SIZE = 7;
	defparam lut_2303.mask = 128'h77ff7fff77ff7fff0080000000000000;

	lut_sub lut_2305 ({sk[851], s298_in_0_, s298_in_2_, s298_out_5_, n_n854, n_n855, n_n856}, x8211x);
	defparam lut_2305.LUT_SIZE = 7;
	defparam lut_2305.mask = 128'h77ff7fff77ff7fff0800000000000000;

	lut_sub lut_2307 ({sk[852], s298_in_0_, s298_in_2_, n_n852, n_n853, n_n856, n_n858}, x8217x);
	defparam lut_2307.LUT_SIZE = 7;
	defparam lut_2307.mask = 128'h77ff7fff77ff7fff0100000000000000;

	lut_sub lut_2309 ({sk[853], s298_in_0_, s298_in_2_, s298_in_1_, n_n854, n_n855, n_n856}, x8223x);
	defparam lut_2309.LUT_SIZE = 7;
	defparam lut_2309.mask = 128'h77ff7fff77ff7fff0000000002000000;

	lut_sub lut_2311 ({sk[854], s298_in_0_, s298_in_2_, n_n857}, x8228x);
	defparam lut_2311.LUT_SIZE = 4;
	defparam lut_2311.mask = 16'h3f80;

	lut_sub lut_2313 ({sk[855], n_n852, n_n854, n_n855, n_n856}, x8229x);
	defparam lut_2313.LUT_SIZE = 5;
	defparam lut_2313.mask = 32'h05ff0020;

	lut_sub lut_2315 ({sk[856], s298_in_2_, s298_in_1_, n_n858}, x8234x);
	defparam lut_2315.LUT_SIZE = 4;
	defparam lut_2315.mask = 16'h3f40;

	lut_sub lut_2317 ({sk[857], n_n852, n_n853, n_n854, n_n855}, x8235x);
	defparam lut_2317.LUT_SIZE = 5;
	defparam lut_2317.mask = 32'h05ff0002;

	lut_sub lut_2319 ({sk[858], s298_in_0_, n_n852, n_n853, n_n854, n_n855, n_n856}, x8241x);
	defparam lut_2319.LUT_SIZE = 7;
	defparam lut_2319.mask = 128'h77ff7fff77ff7fff0000001000000000;

	lut_sub lut_2321 ({sk[859], s298_in_0_, s298_in_1_, n_n852, n_n854, n_n855, n_n857}, x8247x);
	defparam lut_2321.LUT_SIZE = 7;
	defparam lut_2321.mask = 128'h77ff7fff77ff7fff0000000800000000;

	lut_sub lut_2323 ({sk[860], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n856, n_n857}, x8253x);
	defparam lut_2323.LUT_SIZE = 7;
	defparam lut_2323.mask = 128'h77ff7fff77ff7fff0000000000020000;

	lut_sub lut_2325 ({sk[861], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n856, n_n857}, x8259x);
	defparam lut_2325.LUT_SIZE = 7;
	defparam lut_2325.mask = 128'h77ff7fff77ff7fff0000000000000800;

	lut_sub lut_2327 ({sk[862], s298_in_2_, s298_in_1_, n_n852, n_n854, n_n855, n_n857}, x8271x);
	defparam lut_2327.LUT_SIZE = 7;
	defparam lut_2327.mask = 128'h77ff7fff77ff7fff0000008000000000;

	lut_sub lut_2329 ({sk[863], s298_in_0_, s298_in_2_, n_n859}, x8276x);
	defparam lut_2329.LUT_SIZE = 4;
	defparam lut_2329.mask = 16'h3f80;

	lut_sub lut_2331 ({sk[864], s298_in_1_, n_n852, n_n853, n_n855}, x8277x);
	defparam lut_2331.LUT_SIZE = 5;
	defparam lut_2331.mask = 32'h05ff1000;

	lut_sub lut_2333 ({sk[865], s298_in_0_, s298_in_1_, n_n852, n_n854, n_n856, n_n857}, x8283x);
	defparam lut_2333.LUT_SIZE = 7;
	defparam lut_2333.mask = 128'h77ff7fff77ff7fff2000000000000000;

	lut_sub lut_2335 ({sk[866], s298_in_0_, s298_in_1_, s298_out_5_, n_n852, n_n853, n_n857}, x8289x);
	defparam lut_2335.LUT_SIZE = 7;
	defparam lut_2335.mask = 128'h77ff7fff77ff7fff0000100000000000;

	lut_sub lut_2337 ({sk[867], s298_in_0_, s298_in_1_, n_n853, n_n855, n_n856, n_n857}, x8295x);
	defparam lut_2337.LUT_SIZE = 7;
	defparam lut_2337.mask = 128'h77ff7fff77ff7fff0400000000000000;

	lut_sub lut_2339 ({sk[868], s298_in_0_, s298_in_2_, s298_in_1_, n_n854, n_n855, n_n857}, x8307x);
	defparam lut_2339.LUT_SIZE = 7;
	defparam lut_2339.mask = 128'h77ff7fff77ff7fff0010000000000000;

	lut_sub lut_2341 ({sk[869], s298_in_1_, n_n852, n_n854, n_n856}, x8319x);
	defparam lut_2341.LUT_SIZE = 5;
	defparam lut_2341.mask = 32'h05ff4000;

	lut_sub lut_2343 ({sk[870], s298_in_1_, n_n852, n_n853, n_n855}, x8337x);
	defparam lut_2343.LUT_SIZE = 5;
	defparam lut_2343.mask = 32'h05ff0100;

	lut_sub lut_2345 ({sk[871], s298_in_0_, s298_in_1_, n_n853, n_n854, n_n856, n_n857}, x8343x);
	defparam lut_2345.LUT_SIZE = 7;
	defparam lut_2345.mask = 128'h77ff7fff77ff7fff0000000000008000;

	lut_sub lut_2347 ({sk[872], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n856, n_n857}, x8349x);
	defparam lut_2347.LUT_SIZE = 7;
	defparam lut_2347.mask = 128'h77ff7fff77ff7fff0000800000000000;

	lut_sub lut_2349 ({sk[873], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n854, n_n856}, x8355x);
	defparam lut_2349.LUT_SIZE = 7;
	defparam lut_2349.mask = 128'h77ff7fff77ff7fff0000000000004000;

	lut_sub lut_2351 ({sk[874], s298_in_1_, n_n852, n_n853, n_n858}, x8361x);
	defparam lut_2351.LUT_SIZE = 5;
	defparam lut_2351.mask = 32'h05ff4000;

	lut_sub lut_2353 ({sk[875], n_n852, n_n853, n_n854, n_n855}, x8373x);
	defparam lut_2353.LUT_SIZE = 5;
	defparam lut_2353.mask = 32'h05ff0200;

	lut_sub lut_2355 ({sk[876], s298_in_1_, n_n853, n_n854, n_n855}, x8379x);
	defparam lut_2355.LUT_SIZE = 5;
	defparam lut_2355.mask = 32'h05ff2000;

	lut_sub lut_2357 ({sk[877], s298_in_1_, n_n852, n_n853, n_n855}, x8403x);
	defparam lut_2357.LUT_SIZE = 5;
	defparam lut_2357.mask = 32'h05ff0004;

	lut_sub lut_2359 ({sk[878], x8409x, x8410x, x8415x, x8416x}, x8639x);
	defparam lut_2359.LUT_SIZE = 5;
	defparam lut_2359.mask = 32'h05ff111f;

	lut_sub lut_2362 ({sk[879], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, x8422x, x8428x}, x8640x);
	defparam lut_2362.LUT_SIZE = 7;
	defparam lut_2362.mask = 128'h77ff7fff77ff7fff5000000030000000;

	lut_sub lut_2365 ({sk[880], s298_in_1_, n_n852, n_n854, n_n855, x8127x, x161x}, x8641x);
	defparam lut_2365.LUT_SIZE = 7;
	defparam lut_2365.mask = 128'h77ff7fff77ff7fff5555555555557555;

	lut_sub lut_2368 ({sk[881], s298_in_1_, n_n852, n_n853, n_n854, x8134x, x8141x}, x8642x);
	defparam lut_2368.LUT_SIZE = 7;
	defparam lut_2368.mask = 128'h77ff7fff77ff7fff0000000500030000;

	lut_sub lut_2371 ({sk[882], s298_in_1_, n_n852, n_n853, n_n854, x8148x, x8155x}, x8643x);
	defparam lut_2371.LUT_SIZE = 7;
	defparam lut_2371.mask = 128'h77ff7fff77ff7fff0000000000005003;

	lut_sub lut_2374 ({sk[883], s298_in_1_, n_n852, n_n853, n_n854, x8162x, x8169x}, x8644x);
	defparam lut_2374.LUT_SIZE = 7;
	defparam lut_2374.mask = 128'h77ff7fff77ff7fff0005000000000030;

	lut_sub lut_2377 ({sk[884], s298_in_1_, s298_out_3_, n_n852, x8175x, x8176x, x8624x}, x8645x);
	defparam lut_2377.LUT_SIZE = 7;
	defparam lut_2377.mask = 128'h77ff7fff77ff7fff0303570303030303;

	lut_sub lut_2380 ({sk[885], s298_in_0_, s298_in_2_, s298_out_5_, n_n859, x150x, x8361x}, x8647x);
	defparam lut_2380.LUT_SIZE = 7;
	defparam lut_2380.mask = 128'h77ff7fff77ff7fff7333333333333333;

	lut_sub lut_2383 ({sk[886], s298_in_0_, s298_in_2_, s298_out_5_, n_n857, x8549x, x8373x}, x8648x);
	defparam lut_2383.LUT_SIZE = 7;
	defparam lut_2383.mask = 128'h77ff7fff77ff7fff3350330033003300;

	lut_sub lut_2386 ({sk[887], s298_out_5_, x8554x, x8621x}, x8649x);
	defparam lut_2386.LUT_SIZE = 4;
	defparam lut_2386.mask = 16'h3f70;

	lut_sub lut_2389 ({sk[888], s298_in_0_, s298_in_2_, s298_out_4_, n_n856, n_n858, x8337x}, x8658x);
	defparam lut_2389.LUT_SIZE = 7;
	defparam lut_2389.mask = 128'h77ff7fff77ff7fff005000cc000000cc;

	lut_sub lut_2392 ({sk[889], x133x, x8639x, x8640x, x8643x, x8644x, x8645x}, x8660x);
	defparam lut_2392.LUT_SIZE = 7;
	defparam lut_2392.mask = 128'h77ff7fff77ff7fff7fffffffffffffff;

	lut_sub lut_2399 ({sk[890], s298_in_0_, s298_in_2_, s298_out_2_, n_n859, x205x, x8403x}, x8661x);
	defparam lut_2399.LUT_SIZE = 7;
	defparam lut_2399.mask = 128'h77ff7fff77ff7fff3373333333333333;

	lut_sub lut_2402 ({sk[891], x8641x, x8642x, x8647x, x8648x, x8649x, x8658x}, x8663x);
	defparam lut_2402.LUT_SIZE = 7;
	defparam lut_2402.mask = 128'h77ff7fff77ff7fff7fffffffffffffff;

	lut_sub lut_2409 ({sk[892], s298_in_0_, s298_in_2_, n_n856, n_n51, x8559x, x8379x}, x8665x);
	defparam lut_2409.LUT_SIZE = 7;
	defparam lut_2409.mask = 128'h77ff7fff77ff7fff5303030303030303;

	lut_sub lut_2412 ({sk[893], s298_in_0_, s298_in_2_, s298_out_4_, n_n857, x8319x, x12823x}, x12841x);
	defparam lut_2412.LUT_SIZE = 7;
	defparam lut_2412.mask = 128'h77ff7fff77ff7fffffcffffffff5ffff;

	lut_sub lut_2422 ({sk[894], x141x, x8661x, x12841x}, x8668x);
	defparam lut_2422.LUT_SIZE = 4;
	defparam lut_2422.mask = 16'h3fbf;

	lut_sub lut_2426 ({sk[895], s298_in_2_, s298_out_0_, s298_out_1_, s298_out_3_, n_n51, x8617x}, x8672x);
	defparam lut_2426.LUT_SIZE = 7;
	defparam lut_2426.mask = 128'h77ff7fff77ff7fff0000555530005555;

	lut_sub lut_2429 ({sk[896], s298_out_5_, n_n51, x8343x, x8349x, x8665x}, x8673x);
	defparam lut_2429.LUT_SIZE = 6;
	defparam lut_2429.mask = 64'h337f337f557f5555;

	lut_sub lut_2433 ({sk[897], n_n51, x8564x, x8569x, x8637x, x8660x}, x8674x);
	defparam lut_2433.LUT_SIZE = 6;
	defparam lut_2433.mask = 64'h337f337f55557fff;

	lut_sub lut_2438 ({sk[898], s298_out_0_, n_n51, x8070x, x8663x, x8668x}, x8675x);
	defparam lut_2438.LUT_SIZE = 6;
	defparam lut_2438.mask = 64'h337f337f7f777777;

	lut_sub lut_2442 ({sk[899], s298_out_0_, n_n51, x106x, x8544x, x199x, x8084x}, x8676x);
	defparam lut_2442.LUT_SIZE = 7;
	defparam lut_2442.mask = 128'h77ff7fff77ff7fff3fff3fff77ff33ff;

	lut_sub lut_2447 ({sk[900], x8672x, x8673x, x8674x, x8675x, x8676x}, x8680x);
	defparam lut_2447.LUT_SIZE = 6;
	defparam lut_2447.mask = 64'h337f337f7fffffff;

	lut_sub lut_2453 ({sk[901], x104x, x107x, x108x, x8680x}, x8687x);
	defparam lut_2453.LUT_SIZE = 5;
	defparam lut_2453.mask = 32'h05ff7fff;

	lut_sub lut_2458 ({sk[902], s298_out_4_, n_n52, x8113x, x110x, x139x, x8307x}, x8688x);
	defparam lut_2458.LUT_SIZE = 7;
	defparam lut_2458.mask = 128'h77ff7fff77ff7fff3fff3f3f7fff3f3f;

	lut_sub lut_2463 ({sk[903], s298_in_0_, s298_in_2_, n_n855, n_n52, x12840x}, x12822x);
	defparam lut_2463.LUT_SIZE = 6;
	defparam lut_2463.mask = 64'h337f337fffff7fff;

	lut_sub lut_2469 ({sk[904], s298_out_5_, n_n52, x155x, x8355x, x12822x}, x8689x);
	defparam lut_2469.LUT_SIZE = 6;
	defparam lut_2469.mask = 64'h337f337fafbfafaf;

	lut_sub lut_2473 ({sk[905], s298_out_0_, n_n50, x8062x, x8063x, x8271x}, x8693x);
	defparam lut_2473.LUT_SIZE = 6;
	defparam lut_2473.mask = 64'h337f337f03005700;

	lut_sub lut_2476 ({sk[906], s298_out_0_, n_n50, x8276x, x8277x, x8283x}, x8694x);
	defparam lut_2476.LUT_SIZE = 6;
	defparam lut_2476.mask = 64'h337f337f03000355;

	lut_sub lut_2479 ({sk[907], s298_in_2_, s298_out_4_, n_n50, n_n51, x8631x}, x8698x);
	defparam lut_2479.LUT_SIZE = 6;
	defparam lut_2479.mask = 64'h337f337f05053505;

	lut_sub lut_2482 ({sk[908], x101x, x8687x, x8688x, x8689x, x8693x, x8698x}, x8702x);
	defparam lut_2482.LUT_SIZE = 7;
	defparam lut_2482.mask = 128'h77ff7fff77ff7fff7fffffffffffffff;

	lut_sub lut_2489 ({sk[909], n_n50, n_n52, x8524x, x8529x, x8289x, x8295x}, x12821x);
	defparam lut_2489.LUT_SIZE = 7;
	defparam lut_2489.mask = 128'h77ff7fff77ff7ffff000f000ffff8888;

	lut_sub lut_2495 ({sk[910], n_n50, x8534x, x8539x, x8694x, x12821x}, x8703x);
	defparam lut_2495.LUT_SIZE = 6;
	defparam lut_2495.mask = 64'h337f337fbbbbbfff;

	lut_sub lut_2500 ({sk[911], n_n49, x8015x, x8702x, x8703x}, x8705x);
	defparam lut_2500.LUT_SIZE = 5;
	defparam lut_2500.mask = 32'h05ff7f77;

	lut_sub lut_2504 ({sk[912], s298_out_0_, n_n49, n_n51, x8022x, x8027x}, x8706x);
	defparam lut_2504.LUT_SIZE = 6;
	defparam lut_2504.mask = 64'h337f337f33007300;

	lut_sub lut_2507 ({sk[913], s298_out_4_, n_n49, n_n52, x8043x, x8034x}, x8707x);
	defparam lut_2507.LUT_SIZE = 6;
	defparam lut_2507.mask = 64'h337f337f33007300;

	lut_sub lut_2510 ({sk[914], n_n49, n_n50, x8048x, x8049x, x8181x}, x8708x);
	defparam lut_2510.LUT_SIZE = 6;
	defparam lut_2510.mask = 64'h337f337f57030000;

	lut_sub lut_2513 ({sk[915], n_n49, x6018x, x6016x, x6017x, x8187x, x8193x}, x8709x);
	defparam lut_2513.LUT_SIZE = 7;
	defparam lut_2513.mask = 128'h77ff7fff77ff7fff3555555500000000;

	lut_sub lut_2518 ({sk[916], n_n49, n_n50, n_n51, x8199x, x8205x}, x8710x);
	defparam lut_2518.LUT_SIZE = 6;
	defparam lut_2518.mask = 64'h337f337f05370000;

	lut_sub lut_2521 ({sk[917], n_n49, n_n51, n_n52, x8211x, x8217x}, x8711x);
	defparam lut_2521.LUT_SIZE = 6;
	defparam lut_2521.mask = 64'h337f337f30750000;

	lut_sub lut_2524 ({sk[918], n_n49, n_n52, x8223x, x8228x, x8229x}, x8712x);
	defparam lut_2524.LUT_SIZE = 6;
	defparam lut_2524.mask = 64'h337f337f111f0000;

	lut_sub lut_2527 ({sk[919], s298_out_5_, n_n49, x8234x, x8235x, x8241x}, x8713x);
	defparam lut_2527.LUT_SIZE = 6;
	defparam lut_2527.mask = 64'h337f337f03550300;

	lut_sub lut_2530 ({sk[920], s298_out_5_, n_n49, n_n51, x8247x, x8253x}, x8714x);
	defparam lut_2530.LUT_SIZE = 6;
	defparam lut_2530.mask = 64'h337f337f00730050;

	lut_sub lut_2533 ({sk[921], n_n49, n_n52, x8439x, x8259x}, x8715x);
	defparam lut_2533.LUT_SIZE = 5;
	defparam lut_2533.mask = 32'h05ff3305;

	lut_sub lut_2536 ({sk[922], n_n49, x8454x, x8459x, x8464x, x8469x}, x12820x);
	defparam lut_2536.LUT_SIZE = 6;
	defparam lut_2536.mask = 64'h337f337fc000aaaa;

	lut_sub lut_2539 ({sk[923], n_n49, x8494x, x8499x, x8504x, x8509x}, x12819x);
	defparam lut_2539.LUT_SIZE = 6;
	defparam lut_2539.mask = 64'h337f337fffff8000;

	lut_sub lut_2542 ({sk[924], n_n49, x8581x, x8585x, x8589x, x8593x}, x12818x);
	defparam lut_2542.LUT_SIZE = 6;
	defparam lut_2542.mask = 64'h337f337ff0008888;

	lut_sub lut_2546 ({sk[925], s298_in_2_, s298_in_1_, n_n858}, x8769x);
	defparam lut_2546.LUT_SIZE = 4;
	defparam lut_2546.mask = 16'h3f20;

	lut_sub lut_2548 ({sk[926], n_n852, n_n854, n_n855, n_n857}, x8770x);
	defparam lut_2548.LUT_SIZE = 5;
	defparam lut_2548.mask = 32'h05ff4000;

	lut_sub lut_2550 ({sk[927], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_4_, n_n852, n_n857}, x8805x);
	defparam lut_2550.LUT_SIZE = 7;
	defparam lut_2550.mask = 128'h77ff7fff77ff7fff0000000004000000;

	lut_sub lut_2552 ({sk[928], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n854, n_n855}, x8811x);
	defparam lut_2552.LUT_SIZE = 7;
	defparam lut_2552.mask = 128'h77ff7fff77ff7fff0000000000040000;

	lut_sub lut_2554 ({sk[929], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n854, n_n856}, x8817x);
	defparam lut_2554.LUT_SIZE = 7;
	defparam lut_2554.mask = 128'h77ff7fff77ff7fff0000000002000000;

	lut_sub lut_2556 ({sk[930], s298_in_0_, s298_in_2_, s298_in_1_, s298_out_5_, n_n854, n_n857}, x8823x);
	defparam lut_2556.LUT_SIZE = 7;
	defparam lut_2556.mask = 128'h77ff7fff77ff7fff0000000080000000;

	lut_sub lut_2558 ({sk[931], s298_in_0_, s298_in_2_, s298_in_1_, n_n852, n_n854, n_n858}, x8829x);
	defparam lut_2558.LUT_SIZE = 7;
	defparam lut_2558.mask = 128'h77ff7fff77ff7fff2000000000000000;

	lut_sub lut_2560 ({sk[932], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n854, n_n51}, x8835x);
	defparam lut_2560.LUT_SIZE = 7;
	defparam lut_2560.mask = 128'h77ff7fff77ff7fff0000000001000000;

	lut_sub lut_2562 ({sk[933], s298_in_0_, s298_in_1_, n_n853, n_n855, n_n857, n_n858}, x8841x);
	defparam lut_2562.LUT_SIZE = 7;
	defparam lut_2562.mask = 128'h77ff7fff77ff7fff0000000000000020;

	lut_sub lut_2564 ({sk[934], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n856, n_n857}, x8847x);
	defparam lut_2564.LUT_SIZE = 7;
	defparam lut_2564.mask = 128'h77ff7fff77ff7fff0000000000008000;

	lut_sub lut_2566 ({sk[935], s298_in_0_, s298_in_2_, s298_in_1_, n_n853, n_n854, n_n856}, x8853x);
	defparam lut_2566.LUT_SIZE = 7;
	defparam lut_2566.mask = 128'h77ff7fff77ff7fff4000000000000000;

	lut_sub lut_2568 ({sk[936], s298_in_0_, s298_in_2_, n_n858}, x8858x);
	defparam lut_2568.LUT_SIZE = 4;
	defparam lut_2568.mask = 16'h3f04;

	lut_sub lut_2570 ({sk[937], s298_in_1_, n_n852, n_n854, n_n856}, x8859x);
	defparam lut_2570.LUT_SIZE = 5;
	defparam lut_2570.mask = 32'h05ff0040;

	lut_sub lut_2572 ({sk[938], s298_in_0_, s298_in_1_, n_n852, n_n853, n_n855, n_n858}, x8865x);
	defparam lut_2572.LUT_SIZE = 7;
	defparam lut_2572.mask = 128'h77ff7fff77ff7fff0000080000000000;

	lut_sub lut_2574 ({sk[939], s298_in_0_, s298_in_2_, n_n856}, x8870x);
	defparam lut_2574.LUT_SIZE = 4;
	defparam lut_2574.mask = 16'h3f40;

	lut_sub lut_2576 ({sk[940], s298_in_1_, n_n852, n_n853, n_n855}, x8871x);
	defparam lut_2576.LUT_SIZE = 5;
	defparam lut_2576.mask = 32'h05ff0008;

	lut_sub lut_2578 ({sk[941], s298_in_0_, s298_in_2_, n_n856}, x8876x);
	defparam lut_2578.LUT_SIZE = 4;
	defparam lut_2578.mask = 16'h3f08;

	lut_sub lut_2580 ({sk[942], s298_in_1_, n_n852, n_n853, n_n854}, x8877x);
	defparam lut_2580.LUT_SIZE = 5;
	defparam lut_2580.mask = 32'h05ff4000;

	lut_sub lut_2582 ({sk[943], s298_in_0_, s298_in_1_, s298_out_2_, n_n852, n_n853, n_n854}, x8889x);
	defparam lut_2582.LUT_SIZE = 7;
	defparam lut_2582.mask = 128'h77ff7fff77ff7fff0000000000020000;

	lut_sub lut_2584 ({sk[944], s298_in_2_, s298_out_3_, n_n852, n_n853, n_n855}, x8984x);
	defparam lut_2584.LUT_SIZE = 6;
	defparam lut_2584.mask = 64'h337f337f20000000;

	lut_sub lut_2586 ({sk[945], s298_in_0_, s298_in_2_, n_n854, n_n856}, x9053x);
	defparam lut_2586.LUT_SIZE = 5;
	defparam lut_2586.mask = 32'h05ff8000;

	lut_sub lut_2588 ({sk[946], s298_in_1_, n_n852, n_n853, n_n854, x8800x, x9009x}, x9093x);
	defparam lut_2588.LUT_SIZE = 7;
	defparam lut_2588.mask = 128'h77ff7fff77ff7fff0000000000500003;

	lut_sub lut_2591 ({sk[947], s298_out_5_, n_n51, x8786x, x44x, x8990x, x9093x}, x9098x);
	defparam lut_2591.LUT_SIZE = 7;
	defparam lut_2591.mask = 128'h77ff7fff77ff7fff7f7f7fff5f5f5fff;

	lut_sub lut_2596 ({sk[948], s298_out_0_, s298_out_1_, x8960x, x81x, x8870x, x8871x}, x9100x);
	defparam lut_2596.LUT_SIZE = 7;
	defparam lut_2596.mask = 128'h77ff7fff77ff7fff1f1f1fff0f0f0fff;

	lut_sub lut_2600 ({sk[949], s298_out_0_, n_n51, x8876x, x8877x, x8984x}, x9101x);
	defparam lut_2600.LUT_SIZE = 6;
	defparam lut_2600.mask = 64'h337f337f00550303;

	lut_sub lut_2603 ({sk[950], s298_out_1_, n_n51, x8758x, x8955x, x9000x, x9100x}, x9103x);
	defparam lut_2603.LUT_SIZE = 7;
	defparam lut_2603.mask = 128'h77ff7fff77ff7fff55ff77ff5f5f7f7f;

	lut_sub lut_2608 ({sk[951], s298_out_0_, n_n51, x9053x, x9098x, x9101x, x9103x}, x9105x);
	defparam lut_2608.LUT_SIZE = 7;
	defparam lut_2608.mask = 128'h77ff7fff77ff7fff7f7f7f7f7f7f7fff;

	lut_sub lut_2613 ({sk[952], n_n51, n_n52, x8995x, x8889x}, x12815x);
	defparam lut_2613.LUT_SIZE = 5;
	defparam lut_2613.mask = 32'h05ffcf8f;

	lut_sub lut_2617 ({sk[953], n_n52, x27x, x29x, x9005x, x9105x, x12815x}, x9110x);
	defparam lut_2617.LUT_SIZE = 7;
	defparam lut_2617.mask = 128'h77ff7fff77ff7fffbfffffffbbffffff;

	lut_sub lut_2623 ({sk[954], n_n50, n_n51, x8858x, x8859x, x8865x}, x9112x);
	defparam lut_2623.LUT_SIZE = 6;
	defparam lut_2623.mask = 64'h337f337f03035500;

	lut_sub lut_2626 ({sk[955], x6018x, x8970x, x8975x, x6016x, x6017x}, x9114x);
	defparam lut_2626.LUT_SIZE = 6;
	defparam lut_2626.mask = 64'h337f337f07770fff;

	lut_sub lut_2633 ({sk[956], x6018x, x8980x, x9038x, x6016x, x6017x}, x9115x);
	defparam lut_2633.LUT_SIZE = 6;
	defparam lut_2633.mask = 64'h337f337f07770fff;

	lut_sub lut_2640 ({sk[957], s298_in_0_, s298_out_1_, n_n852, n_n853, n_n50, x9050x}, x9117x);
	defparam lut_2640.LUT_SIZE = 7;
	defparam lut_2640.mask = 128'h77ff7fff77ff7fff1111111111111311;

	lut_sub lut_2643 ({sk[958], s298_out_0_, n_n855, n_n50, n_n857, n_n51, x9076x}, x9118x);
	defparam lut_2643.LUT_SIZE = 7;
	defparam lut_2643.mask = 128'h77ff7fff77ff7fff0055005500550075;

	lut_sub lut_2646 ({sk[959], s298_in_1_, s298_out_4_, n_n853, n_n50, n_n858, x9082x}, x9119x);
	defparam lut_2646.LUT_SIZE = 7;
	defparam lut_2646.mask = 128'h77ff7fff77ff7fff0505050d05050505;

	lut_sub lut_2649 ({sk[960], s298_in_0_, s298_in_2_, s298_out_5_, n_n854, n_n50, n_n858}, x9120x);
	defparam lut_2649.LUT_SIZE = 7;
	defparam lut_2649.mask = 128'h77ff7fff77ff7fff0200333300003333;

	lut_sub lut_2652 ({sk[961], n_n50, x9042x, x9046x, x9115x, x9117x, x9118x}, x9127x);
	defparam lut_2652.LUT_SIZE = 7;
	defparam lut_2652.mask = 128'h77ff7fff77ff7fff7f7f7f7f7fffffff;

	lut_sub lut_2658 ({sk[962], n_n50, n_n51, x8950x, x8965x, x8853x, x9110x}, x12814x);
	defparam lut_2658.LUT_SIZE = 7;
	defparam lut_2658.mask = 128'h77ff7fff77ff7fffa0008000aaaaaaaa;

	lut_sub lut_2662 ({sk[963], x9112x, x9114x, x9119x, x9120x, x12814x}, x9128x);
	defparam lut_2662.LUT_SIZE = 6;
	defparam lut_2662.mask = 64'h337f337fbfffffff;

	lut_sub lut_2668 ({sk[964], n_n49, x8765x, x9127x, x9128x}, x9130x);
	defparam lut_2668.LUT_SIZE = 5;
	defparam lut_2668.mask = 32'h05ff7f77;

	lut_sub lut_2672 ({sk[965], s298_out_0_, n_n49, n_n52, x8769x, x8770x, x8805x}, x9131x);
	defparam lut_2672.LUT_SIZE = 7;
	defparam lut_2672.mask = 128'h77ff7fff77ff7fff0055000003570000;

	lut_sub lut_2675 ({sk[966], s298_out_4_, n_n49, x8811x, x8817x}, x9132x);
	defparam lut_2675.LUT_SIZE = 5;
	defparam lut_2675.mask = 32'h05ff0070;

	lut_sub lut_2678 ({sk[967], n_n49, n_n51, x8823x, x8829x}, x9133x);
	defparam lut_2678.LUT_SIZE = 5;
	defparam lut_2678.mask = 32'h05ff0700;

	lut_sub lut_2681 ({sk[968], n_n49, x6018x, x6016x, x6017x, x8835x, x8841x}, x9134x);
	defparam lut_2681.LUT_SIZE = 7;
	defparam lut_2681.mask = 128'h77ff7fff77ff7fff0000000035555555;

	lut_sub lut_2686 ({sk[969], n_n49, n_n52, x8895x, x8847x}, x9135x);
	defparam lut_2686.LUT_SIZE = 5;
	defparam lut_2686.mask = 32'h05ff3305;

	lut_sub lut_2689 ({sk[970], s298_out_0_, n_n853, n_n854, n_n49, n_n856, x9061x}, x9144x);
	defparam lut_2689.LUT_SIZE = 7;
	defparam lut_2689.mask = 128'h77ff7fff77ff7fff5050505350505050;

	lut_sub lut_2692 ({sk[971], n_n855, n_n49, n_n856, n_n858, n_n859, x9067x}, x9145x);
	defparam lut_2692.LUT_SIZE = 7;
	defparam lut_2692.mask = 128'h77ff7fff77ff7fff0000555700005555;

	lut_sub lut_2695 ({sk[972], n_n854, n_n855, n_n49, n_n858, x9090x}, x9146x);
	defparam lut_2695.LUT_SIZE = 6;
	defparam lut_2695.mask = 64'h337f337f07050505;

	lut_sub lut_2698 ({sk[973], n_n49, x8900x, x8905x, x8910x, x8915x}, x12817x);
	defparam lut_2698.LUT_SIZE = 6;
	defparam lut_2698.mask = 64'h337f337f8000ffff;

	lut_sub lut_2701 ({sk[974], n_n49, x8940x, x8945x, x9014x, x9018x}, x12816x);
	defparam lut_2701.LUT_SIZE = 6;
	defparam lut_2701.mask = 64'h337f337f8888f000;

	lut_sub lut_2705 ({sk[975], s298_in_1_, n_n852, n_n853, n_n854}, x12840x);
	defparam lut_2705.LUT_SIZE = 5;
	defparam lut_2705.mask = 32'h05fffddf;

	lut_sub lut_2710 ({sk[976], n_n852, n_n853, n_n854, n_n855, n_n856}, x12823x);
	defparam lut_2710.LUT_SIZE = 6;
	defparam lut_2710.mask = 64'h337f337fffddf5ff;

	lut_sub lut_2719 ({sk[977], s298_in_1_, n_n852, n_n853, n_n854, n_n857, n_n858}, x12842x);
	defparam lut_2719.LUT_SIZE = 7;
	defparam lut_2719.mask = 128'h77ff7fff77ff7fffccfffffafffffffa;

	lut_sub lut_2734 ({sk[978], s298_in_2_, s298_out_4_, n_n852, n_n854, n_n855, n_n856}, x12835x);
	defparam lut_2734.LUT_SIZE = 7;
	defparam lut_2734.mask = 128'h77ff7fff77ff7ffffffffbbbffffffff;


endmodule