module apex2x5xv (i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_28_, i_13_, i_4_, i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_, i_16_, i_22_, i_15_, i_32_, i_31_, i_34_, i_33_, i_19_, i_36_, i_35_, i_38_, i_29_, i_37_, o_1_, o_2_, o_0_);

	input i_30_;
	input i_20_;
	input i_9_;
	input i_10_;
	input i_7_;
	input i_8_;
	input i_5_;
	input i_6_;
	input i_27_;
	input i_14_;
	input i_3_;
	input i_28_;
	input i_13_;
	input i_4_;
	input i_25_;
	input i_12_;
	input i_1_;
	input i_26_;
	input i_11_;
	input i_2_;
	input i_23_;
	input i_18_;
	input i_24_;
	input i_17_;
	input i_0_;
	input i_21_;
	input i_16_;
	input i_22_;
	input i_15_;
	input i_32_;
	input i_31_;
	input i_34_;
	input i_33_;
	input i_19_;
	input i_36_;
	input i_35_;
	input i_38_;
	input i_29_;
	input i_37_;
	output o_1_;
	output o_2_;
	output o_0_;

	wire [1337 : 0] sk /* synthesis noprune */;

	lut_sub lut_3 ({sk[0], x7257x, x7252x, x7044x, x7045x, x7250x}, o_1_);
	defparam lut_3.LUT_SIZE = 6;
	defparam lut_3.mask = 64'h55ffffff7fffffff;

	lut_sub lut_9 ({sk[1], x7747x, n_n1811, x7746x}, o_2_);
	defparam lut_9.LUT_SIZE = 4;
	defparam lut_9.mask = 16'h557f;

	lut_sub lut_13 ({sk[2], x8098x, x8080x, x8054x, x8055x}, o_0_);
	defparam lut_13.LUT_SIZE = 5;
	defparam lut_13.mask = 32'h37377fff;

	lut_sub lut_18 ({sk[3], n_n1696, n_n1695, x1465x}, x7257x);
	defparam lut_18.LUT_SIZE = 4;
	defparam lut_18.mask = 16'h557f;

	lut_sub lut_22 ({sk[4], n_n1710, x7094x, x7240x, x7241x}, x7252x);
	defparam lut_22.LUT_SIZE = 5;
	defparam lut_22.mask = 32'h0f0f7fff;

	lut_sub lut_27 ({sk[5], n_n1720, x6992x, n_n1722, x7040x, x7041x}, x7044x);
	defparam lut_27.LUT_SIZE = 6;
	defparam lut_27.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_33 ({sk[6], x7023x, n_n1723, x7020x, x7021x}, x7045x);
	defparam lut_33.LUT_SIZE = 5;
	defparam lut_33.mask = 32'h0f0f7fff;

	lut_sub lut_38 ({sk[7], n_n1707, n_n1706, n_n1708, n_n1713, x7246x}, x7250x);
	defparam lut_38.LUT_SIZE = 6;
	defparam lut_38.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_44 ({sk[8], x7349x, x7350x, n_n1829, n_n1812}, x7747x);
	defparam lut_44.LUT_SIZE = 5;
	defparam lut_44.mask = 32'h0f0f7fff;

	lut_sub lut_49 ({sk[9], n_n1831, x7599x, n_n1818, n_n1835, x7713x}, n_n1811);
	defparam lut_49.LUT_SIZE = 6;
	defparam lut_49.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_55 ({sk[10], x7486x, n_n1822, n_n1821, x7744x}, x7746x);
	defparam lut_55.LUT_SIZE = 5;
	defparam lut_55.mask = 32'h0f0f7fff;

	lut_sub lut_60 ({sk[11], n_n1558, n_n1559, n_n1560, x8095x}, x8098x);
	defparam lut_60.LUT_SIZE = 5;
	defparam lut_60.mask = 32'h0f0f7fff;

	lut_sub lut_65 ({sk[12], n_n1549, n_n1548, x7922x, x8079x}, x8080x);
	defparam lut_65.LUT_SIZE = 5;
	defparam lut_65.mask = 32'h0f0f7fff;

	lut_sub lut_70 ({sk[13], x7955x, x7956x, x8037x, x8038x, x8051x}, x8054x);
	defparam lut_70.LUT_SIZE = 6;
	defparam lut_70.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_76 ({sk[14], n_n1571, n_n1570, n_n1572, x8049x}, x8055x);
	defparam lut_76.LUT_SIZE = 5;
	defparam lut_76.mask = 32'h0f0f7fff;

	lut_sub lut_81 ({sk[15], x6898x, x10x, n_n1318, x1759x, x603x}, n_n1696);
	defparam lut_81.LUT_SIZE = 6;
	defparam lut_81.mask = 64'h37ff37ff0307ffff;

	lut_sub lut_85 ({sk[16], n_n26, x1748x, x6916x, x6917x, x6918x}, n_n1695);
	defparam lut_85.LUT_SIZE = 6;
	defparam lut_85.mask = 64'h37ff37ff77777fff;

	lut_sub lut_90 ({sk[17], i_33_, i_37_, x1469x, n_n178, x357x}, x1465x);
	defparam lut_90.LUT_SIZE = 6;
	defparam lut_90.mask = 64'h37ff37ff001f0000;

	lut_sub lut_93 ({sk[18], x1457x, x7267x, x7291x, n_n1860}, x7349x);
	defparam lut_93.LUT_SIZE = 5;
	defparam lut_93.mask = 32'h0f0f7fff;

	lut_sub lut_98 ({sk[19], x7315x, x7316x, n_n1859, n_n1861}, x7350x);
	defparam lut_98.LUT_SIZE = 5;
	defparam lut_98.mask = 32'h0f0f7fff;

	lut_sub lut_103 ({sk[20], x7408x, x1347x, x7396x, x7406x}, n_n1829);
	defparam lut_103.LUT_SIZE = 5;
	defparam lut_103.mask = 32'h0f0f7fff;

	lut_sub lut_108 ({sk[21], n_n1842, n_n1843, x7434x, x1296x, x7440x}, n_n1812);
	defparam lut_108.LUT_SIZE = 6;
	defparam lut_108.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_114 ({sk[22], i_36_, x7760x, x25x, x7759x, x273x}, n_n1558);
	defparam lut_114.LUT_SIZE = 6;
	defparam lut_114.mask = 64'h37ff37ff00ff37ff;

	lut_sub lut_118 ({sk[23], i_36_, x7771x, x7767x, x7768x}, n_n1559);
	defparam lut_118.LUT_SIZE = 5;
	defparam lut_118.mask = 32'h0f0f0f7f;

	lut_sub lut_122 ({sk[24], x945x, x944x, x7780x}, n_n1560);
	defparam lut_122.LUT_SIZE = 4;
	defparam lut_122.mask = 16'h777f;

	lut_sub lut_126 ({sk[25], x19x, x493x, x6x, x22x, x32x}, x8095x);
	defparam lut_126.LUT_SIZE = 6;
	defparam lut_126.mask = 64'h37ff37ff7f7f7fff;

	lut_sub lut_131 ({sk[26], n_n1307, n_n1278, n_n1100, x219x, x326x}, x19x);
	defparam lut_131.LUT_SIZE = 6;
	defparam lut_131.mask = 64'h37ff37ff00330537;

	lut_sub lut_134 ({sk[27], i_9_, n_n1406, n_n1303, n_n1213, n_n629}, x233x);
	defparam lut_134.LUT_SIZE = 6;
	defparam lut_134.mask = 64'h37ff37ff00010000;

	lut_sub lut_136 ({sk[28], i_27_, i_35_, i_37_, x42x, n_n1311}, x492x);
	defparam lut_136.LUT_SIZE = 6;
	defparam lut_136.mask = 64'h37ff37ff00010000;

	lut_sub lut_138 ({sk[29], i_10_, i_13_, i_33_, i_37_, n_n245}, x6880x);
	defparam lut_138.LUT_SIZE = 6;
	defparam lut_138.mask = 64'h37ff37ff10000000;

	lut_sub lut_140 ({sk[30], x1766x, n_n129, x267x, n_n130, x246x}, x1756x);
	defparam lut_140.LUT_SIZE = 6;
	defparam lut_140.mask = 64'h37ff37ff00010505;

	lut_sub lut_143 ({sk[31], x19x, x233x, x492x, x6880x, x1756x}, x6898x);
	defparam lut_143.LUT_SIZE = 6;
	defparam lut_143.mask = 64'h37ff37ff55775f7f;

	lut_sub lut_147 ({sk[32], i_14_, i_16_}, x10x);
	defparam lut_147.LUT_SIZE = 3;
	defparam lut_147.mask = 8'h58;

	lut_sub lut_149 ({sk[33], i_35_, i_37_}, n_n1318);
	defparam lut_149.LUT_SIZE = 3;
	defparam lut_149.mask = 8'h54;

	lut_sub lut_151 ({sk[34], i_14_, i_17_, i_16_, x63x, x604x}, x1759x);
	defparam lut_151.LUT_SIZE = 6;
	defparam lut_151.mask = 64'h37ff37ff10000000;

	lut_sub lut_153 ({sk[35], i_9_, n_n1118, n_n26, n_n21, x1762x}, x603x);
	defparam lut_153.LUT_SIZE = 6;
	defparam lut_153.mask = 64'h37ff37ff55575555;

	lut_sub lut_156 ({sk[36], i_3_, i_4_, i_0_}, n_n26);
	defparam lut_156.LUT_SIZE = 4;
	defparam lut_156.mask = 16'h7708;

	lut_sub lut_158 ({sk[37], i_9_, i_37_, n_n1278, x1753x, x1754x}, x1748x);
	defparam lut_158.LUT_SIZE = 6;
	defparam lut_158.mask = 64'h37ff37ff00070000;

	lut_sub lut_161 ({sk[38], i_9_, x43x, n_n21, x606x, x1750x}, x6916x);
	defparam lut_161.LUT_SIZE = 6;
	defparam lut_161.mask = 64'h37ff37ff55575555;

	lut_sub lut_164 ({sk[39], n_n504, n_n178, n_n18, x487x, x1745x}, x6917x);
	defparam lut_164.LUT_SIZE = 6;
	defparam lut_164.mask = 64'h37ff37ff55555557;

	lut_sub lut_167 ({sk[40], i_11_, x268x, x357x, x508x, x6901x}, x6918x);
	defparam lut_167.LUT_SIZE = 6;
	defparam lut_167.mask = 64'h37ff37ff111f1111;

	lut_sub lut_170 ({sk[41], i_0_, i_37_, x7062x, x1634x, x769x}, n_n1710);
	defparam lut_170.LUT_SIZE = 6;
	defparam lut_170.mask = 64'h37ff37ff0f7f0f3f;

	lut_sub lut_174 ({sk[42], x1619x, x7077x, x1608x, x7090x, x7091x}, x7094x);
	defparam lut_174.LUT_SIZE = 6;
	defparam lut_174.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_180 ({sk[43], n_n1697, n_n1701, n_n1702, x7235x}, x7240x);
	defparam lut_180.LUT_SIZE = 5;
	defparam lut_180.mask = 32'h0f0f7fff;

	lut_sub lut_185 ({sk[44], n_n1698, n_n1699, n_n1703, n_n1704, n_n1705}, x7241x);
	defparam lut_185.LUT_SIZE = 6;
	defparam lut_185.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_191 ({sk[45], i_33_, i_37_}, x59x);
	defparam lut_191.LUT_SIZE = 3;
	defparam lut_191.mask = 8'h54;

	lut_sub lut_193 ({sk[46], i_11_, i_17_, i_16_, i_19_}, x431x);
	defparam lut_193.LUT_SIZE = 5;
	defparam lut_193.mask = 32'h0f0f8000;

	lut_sub lut_195 ({sk[47], i_7_, i_8_, i_6_, x88x}, x508x);
	defparam lut_195.LUT_SIZE = 5;
	defparam lut_195.mask = 32'h0f0f4000;

	lut_sub lut_197 ({sk[48], i_8_, n_n1278, n_n132, n_n26, x274x}, x1471x);
	defparam lut_197.LUT_SIZE = 6;
	defparam lut_197.mask = 64'h37ff37ff00010000;

	lut_sub lut_199 ({sk[49], i_9_, i_13_, x431x, x508x, x1471x}, x1469x);
	defparam lut_199.LUT_SIZE = 6;
	defparam lut_199.mask = 64'h37ff37ff57000000;

	lut_sub lut_202 ({sk[50], i_38_, x52x, x1462x, x9219x}, x1457x);
	defparam lut_202.LUT_SIZE = 5;
	defparam lut_202.mask = 32'h0f0f003b;

	lut_sub lut_205 ({sk[51], n_n762, n_n416, x70x, n_n706, x579x}, x7267x);
	defparam lut_205.LUT_SIZE = 6;
	defparam lut_205.mask = 64'h37ff37ff030f575f;

	lut_sub lut_209 ({sk[52], x1449x, x1437x, x1450x, x7282x, x7289x}, x7291x);
	defparam lut_209.LUT_SIZE = 6;
	defparam lut_209.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_215 ({sk[53], i_34_, n_n1300, x715x, x7337x, x7338x}, n_n1860);
	defparam lut_215.LUT_SIZE = 6;
	defparam lut_215.mask = 64'h37ff37ff7777777f;

	lut_sub lut_219 ({sk[54], i_25_, n_n1486, x1431x, x7304x, x354x}, x7315x);
	defparam lut_219.LUT_SIZE = 6;
	defparam lut_219.mask = 64'h37ff37ff3f7f3f3f;

	lut_sub lut_223 ({sk[55], n_n1128, x623x, x1408x, x1419x, x7312x}, x7316x);
	defparam lut_223.LUT_SIZE = 6;
	defparam lut_223.mask = 64'h37ff37ff7f7f7fff;

	lut_sub lut_228 ({sk[56], i_32_, x1399x, x7326x, x9218x}, n_n1859);
	defparam lut_228.LUT_SIZE = 5;
	defparam lut_228.mask = 32'h0f0fbf3f;

	lut_sub lut_232 ({sk[57], x223x, x7346x, x346x, x379x, x1383x}, n_n1861);
	defparam lut_232.LUT_SIZE = 6;
	defparam lut_232.mask = 64'h37ff37ff57ff77ff;

	lut_sub lut_237 ({sk[58], i_9_, i_8_, i_18_, n_n1278, n_n787}, n_n416);
	defparam lut_237.LUT_SIZE = 6;
	defparam lut_237.mask = 64'h37ff37ff10000000;

	lut_sub lut_239 ({sk[59], i_28_, i_25_, i_38_, i_29_, x73x}, x456x);
	defparam lut_239.LUT_SIZE = 6;
	defparam lut_239.mask = 64'h37ff37ff04000000;

	lut_sub lut_241 ({sk[60], i_32_, i_38_, i_29_, n_n1478, x26x}, x1367x);
	defparam lut_241.LUT_SIZE = 6;
	defparam lut_241.mask = 64'h37ff37ff00100000;

	lut_sub lut_243 ({sk[61], i_31_, x261x, n_n316, x218x, x387x}, x7368x);
	defparam lut_243.LUT_SIZE = 6;
	defparam lut_243.mask = 64'h37ff37ff03570055;

	lut_sub lut_246 ({sk[62], x1364x, x1365x, x1366x, x1369x}, x7369x);
	defparam lut_246.LUT_SIZE = 5;
	defparam lut_246.mask = 32'h0f0f7fff;

	lut_sub lut_251 ({sk[63], n_n416, x456x, x1367x, x7368x, x7369x}, n_n1863);
	defparam lut_251.LUT_SIZE = 6;
	defparam lut_251.mask = 64'h37ff37ff7f7f7fff;

	lut_sub lut_256 ({sk[64], i_31_, x53x, x421x, x1374x, x9233x}, x7359x);
	defparam lut_256.LUT_SIZE = 6;
	defparam lut_256.mask = 64'h37ff37ffbbbfbbbb;

	lut_sub lut_260 ({sk[65], n_n706, x456x, x714x, x7352x, x1375x}, x7360x);
	defparam lut_260.LUT_SIZE = 6;
	defparam lut_260.mask = 64'h37ff37ff575757ff;

	lut_sub lut_264 ({sk[66], i_13_, x377x, x7375x, x37x}, x1356x);
	defparam lut_264.LUT_SIZE = 5;
	defparam lut_264.mask = 32'h0f0f0703;

	lut_sub lut_267 ({sk[67], i_13_, i_31_, n_n316, x207x, x310x}, x7380x);
	defparam lut_267.LUT_SIZE = 6;
	defparam lut_267.mask = 64'h37ff37ff03005755;

	lut_sub lut_270 ({sk[68], i_10_, x15x, x387x, x1353x, x1354x}, x7381x);
	defparam lut_270.LUT_SIZE = 6;
	defparam lut_270.mask = 64'h37ff37ff777f7777;

	lut_sub lut_274 ({sk[69], x7359x, x7360x, x1356x, x7380x, x7381x}, x7384x);
	defparam lut_274.LUT_SIZE = 6;
	defparam lut_274.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_280 ({sk[70], i_30_, i_28_, i_29_}, n_n1489);
	defparam lut_280.LUT_SIZE = 4;
	defparam lut_280.mask = 16'h7780;

	lut_sub lut_282 ({sk[71], x261x, x388x, x70x, x346x, x1334x}, x7401x);
	defparam lut_282.LUT_SIZE = 6;
	defparam lut_282.mask = 64'h37ff37ff575757ff;

	lut_sub lut_286 ({sk[72], i_13_, x239x, n_n1422, n_n1058, x436x}, x1338x);
	defparam lut_286.LUT_SIZE = 6;
	defparam lut_286.mask = 64'h37ff37ff00070005;

	lut_sub lut_289 ({sk[73], i_24_, i_38_, n_n1437, x425x, x454x}, x1339x);
	defparam lut_289.LUT_SIZE = 6;
	defparam lut_289.mask = 64'h37ff37ff00070000;

	lut_sub lut_292 ({sk[74], i_38_, x261x, x52x, x223x, x1330x}, x1327x);
	defparam lut_292.LUT_SIZE = 6;
	defparam lut_292.mask = 64'h37ff37ff0000575f;

	lut_sub lut_296 ({sk[75], n_n1489, x7401x, x1338x, x1339x, x1327x}, x7408x);
	defparam lut_296.LUT_SIZE = 6;
	defparam lut_296.mask = 64'h37ff37ff55ff7fff;

	lut_sub lut_301 ({sk[76], i_33_, n_n1361, x1349x, x1351x, x9217x}, x1347x);
	defparam lut_301.LUT_SIZE = 6;
	defparam lut_301.mask = 64'h37ff37ff00bf0000;

	lut_sub lut_305 ({sk[77], x1344x, x1345x, x1346x, x1348x}, x7396x);
	defparam lut_305.LUT_SIZE = 5;
	defparam lut_305.mask = 32'h0f0f7fff;

	lut_sub lut_310 ({sk[78], i_24_, i_38_, x78x, x346x, x9216x}, x7406x);
	defparam lut_310.LUT_SIZE = 6;
	defparam lut_310.mask = 64'h37ff37ffaaabaaaa;

	lut_sub lut_313 ({sk[79], i_19_, x520x, x28x, x1318x, x1317x}, n_n1842);
	defparam lut_313.LUT_SIZE = 6;
	defparam lut_313.mask = 64'h37ff37ff7777777f;

	lut_sub lut_317 ({sk[80], x288x, x12x, x20x, x1315x, x1314x}, n_n1843);
	defparam lut_317.LUT_SIZE = 6;
	defparam lut_317.mask = 64'h37ff37ff7777777f;

	lut_sub lut_321 ({sk[81], n_n300, x100x, x98x, x1309x, x7432x}, x7434x);
	defparam lut_321.LUT_SIZE = 6;
	defparam lut_321.mask = 64'h37ff37ff77777fff;

	lut_sub lut_326 ({sk[82], i_19_, x21x, x28x, x276x, x7438x}, x1296x);
	defparam lut_326.LUT_SIZE = 6;
	defparam lut_326.mask = 64'h37ff37ff00331333;

	lut_sub lut_330 ({sk[83], x20x, x276x, x1297x, x1304x, x9215x}, x7440x);
	defparam lut_330.LUT_SIZE = 6;
	defparam lut_330.mask = 64'h37ff37ffbfbfbfff;

	lut_sub lut_335 ({sk[84], n_n805, n_n1466, x4x, x30x, x7450x}, x651x);
	defparam lut_335.LUT_SIZE = 6;
	defparam lut_335.mask = 64'h37ff37ff05050537;

	lut_sub lut_338 ({sk[85], i_8_, i_18_, x60x, n_n706, x387x}, x1286x);
	defparam lut_338.LUT_SIZE = 6;
	defparam lut_338.mask = 64'h37ff37ff15111111;

	lut_sub lut_341 ({sk[86], x61x, x226x, x231x, x521x, x1285x}, x7451x);
	defparam lut_341.LUT_SIZE = 6;
	defparam lut_341.mask = 64'h37ff37ff5555557f;

	lut_sub lut_345 ({sk[87], x1290x, x7445x, x1240x, x7481x, x7482x}, x7485x);
	defparam lut_345.LUT_SIZE = 6;
	defparam lut_345.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_351 ({sk[88], i_31_, x651x, x1286x, x7451x, x7485x}, x7486x);
	defparam lut_351.LUT_SIZE = 6;
	defparam lut_351.mask = 64'h37ff37ff7fff7f7f;

	lut_sub lut_356 ({sk[89], x7550x, x7551x, n_n1876, x7568x, x7569x}, n_n1831);
	defparam lut_356.LUT_SIZE = 6;
	defparam lut_356.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_362 ({sk[90], n_n1872, n_n1877, x7596x, x7597x}, x7599x);
	defparam lut_362.LUT_SIZE = 5;
	defparam lut_362.mask = 32'h0f0f7fff;

	lut_sub lut_367 ({sk[91], n_n1891, n_n1889, n_n1837, x7621x, x7642x}, n_n1818);
	defparam lut_367.LUT_SIZE = 6;
	defparam lut_367.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_373 ({sk[92], x1013x, x7699x, x7707x, x7708x}, n_n1835);
	defparam lut_373.LUT_SIZE = 5;
	defparam lut_373.mask = 32'h0f0f7fff;

	lut_sub lut_378 ({sk[93], n_n1880, n_n1883, x7681x, x7710x}, x7713x);
	defparam lut_378.LUT_SIZE = 5;
	defparam lut_378.mask = 32'h0f0f7fff;

	lut_sub lut_383 ({sk[94], i_29_, n_n416, n_n1300, n_n1497, n_n706}, x990x);
	defparam lut_383.LUT_SIZE = 6;
	defparam lut_383.mask = 64'h37ff37ff01030000;

	lut_sub lut_386 ({sk[95], i_32_, i_33_, i_38_, n_n1486, x26x}, x991x);
	defparam lut_386.LUT_SIZE = 6;
	defparam lut_386.mask = 64'h37ff37ff01000000;

	lut_sub lut_388 ({sk[96], i_34_, n_n1361, n_n1302, n_n849, x994x}, x992x);
	defparam lut_388.LUT_SIZE = 6;
	defparam lut_388.mask = 64'h37ff37ff00000057;

	lut_sub lut_391 ({sk[97], i_32_, x218x, x408x, x421x, x66x}, x993x);
	defparam lut_391.LUT_SIZE = 6;
	defparam lut_391.mask = 64'h37ff37ff15551515;

	lut_sub lut_395 ({sk[98], x990x, x991x, x992x, x993x}, n_n1866);
	defparam lut_395.LUT_SIZE = 5;
	defparam lut_395.mask = 32'h0f0f7fff;

	lut_sub lut_400 ({sk[99], i_34_, i_35_, i_38_}, n_n805);
	defparam lut_400.LUT_SIZE = 4;
	defparam lut_400.mask = 16'h7704;

	lut_sub lut_402 ({sk[100], i_28_, i_25_, i_29_}, n_n1466);
	defparam lut_402.LUT_SIZE = 4;
	defparam lut_402.mask = 16'h7780;

	lut_sub lut_404 ({sk[101], i_9_, i_10_, i_8_, i_24_, x11x}, n_n849);
	defparam lut_404.LUT_SIZE = 6;
	defparam lut_404.mask = 64'h37ff37ff00004000;

	lut_sub lut_406 ({sk[102], i_24_, i_34_, n_n1361, x344x, x335x}, x982x);
	defparam lut_406.LUT_SIZE = 6;
	defparam lut_406.mask = 64'h37ff37ff00010000;

	lut_sub lut_408 ({sk[103], i_32_, i_31_, i_29_, x207x, x315x}, x984x);
	defparam lut_408.LUT_SIZE = 6;
	defparam lut_408.mask = 64'h37ff37ff10000000;

	lut_sub lut_410 ({sk[104], n_n805, n_n1466, n_n849, x982x, x984x}, x7729x);
	defparam lut_410.LUT_SIZE = 6;
	defparam lut_410.mask = 64'h37ff37ff7777777f;

	lut_sub lut_414 ({sk[105], i_28_, i_32_, i_33_, n_n1361, n_n1523}, n_n316);
	defparam lut_414.LUT_SIZE = 6;
	defparam lut_414.mask = 64'h37ff37ff10000000;

	lut_sub lut_416 ({sk[106], i_9_, n_n1497, x5x, x349x, x989x}, x763x);
	defparam lut_416.LUT_SIZE = 6;
	defparam lut_416.mask = 64'h37ff37ff5555557f;

	lut_sub lut_420 ({sk[107], i_2_, i_33_, i_35_, i_38_, x3x}, x7724x);
	defparam lut_420.LUT_SIZE = 6;
	defparam lut_420.mask = 64'h37ff37ff20000000;

	lut_sub lut_422 ({sk[108], i_9_, i_10_, i_6_, i_12_, n_n1307}, x7726x);
	defparam lut_422.LUT_SIZE = 6;
	defparam lut_422.mask = 64'h37ff37ff00004000;

	lut_sub lut_424 ({sk[109], i_10_, x310x}, x986x);
	defparam lut_424.LUT_SIZE = 3;
	defparam lut_424.mask = 8'h54;

	lut_sub lut_426 ({sk[110], n_n316, x763x, x7724x, x7726x, x986x}, x7730x);
	defparam lut_426.LUT_SIZE = 6;
	defparam lut_426.mask = 64'h37ff37ff555f777f;

	lut_sub lut_430 ({sk[111], i_35_, i_38_}, n_n1361);
	defparam lut_430.LUT_SIZE = 3;
	defparam lut_430.mask = 8'h54;

	lut_sub lut_432 ({sk[112], i_28_, i_25_, i_26_, i_29_, x12x}, x330x);
	defparam lut_432.LUT_SIZE = 6;
	defparam lut_432.mask = 64'h37ff37ff40000000;

	lut_sub lut_434 ({sk[113], i_10_, i_13_, i_31_, n_n1307, n_n841}, x790x);
	defparam lut_434.LUT_SIZE = 6;
	defparam lut_434.mask = 64'h37ff37ff10100010;

	lut_sub lut_437 ({sk[114], x73x, n_n1486, n_n1288, x335x, x394x}, x9212x);
	defparam lut_437.LUT_SIZE = 6;
	defparam lut_437.mask = 64'h37ff37ffffaafca8;

	lut_sub lut_444 ({sk[115], i_33_, n_n1361, x330x, x790x, x9212x}, x7740x);
	defparam lut_444.LUT_SIZE = 6;
	defparam lut_444.mask = 64'h37ff37ff03ab0303;

	lut_sub lut_447 ({sk[116], i_36_, i_35_}, n_n880);
	defparam lut_447.LUT_SIZE = 3;
	defparam lut_447.mask = 8'h52;

	lut_sub lut_449 ({sk[117], i_9_, i_4_, x224x, x44x, x7749x}, x64x);
	defparam lut_449.LUT_SIZE = 6;
	defparam lut_449.mask = 64'h37ff37ff01000000;

	lut_sub lut_451 ({sk[118], i_23_, i_17_, i_21_, x43x, x45x}, x463x);
	defparam lut_451.LUT_SIZE = 6;
	defparam lut_451.mask = 64'h37ff37ff10000000;

	lut_sub lut_453 ({sk[119], i_8_, x204x, x232x, n_n841, x338x}, x547x);
	defparam lut_453.LUT_SIZE = 6;
	defparam lut_453.mask = 64'h37ff37ff111f1111;

	lut_sub lut_456 ({sk[120], i_3_, i_13_, n_n132, n_n576, x431x}, x7751x);
	defparam lut_456.LUT_SIZE = 6;
	defparam lut_456.mask = 64'h37ff37ff11001300;

	lut_sub lut_459 ({sk[121], n_n880, x64x, x463x, x547x, x7751x}, x7760x);
	defparam lut_459.LUT_SIZE = 6;
	defparam lut_459.mask = 64'h37ff37ff00550357;

	lut_sub lut_462 ({sk[122], i_18_, i_19_, x263x, n_n29, n_n129}, x25x);
	defparam lut_462.LUT_SIZE = 6;
	defparam lut_462.mask = 64'h37ff37ff07030500;

	lut_sub lut_465 ({sk[123], i_14_, i_13_, x15x, x373x, x7758x}, x7759x);
	defparam lut_465.LUT_SIZE = 6;
	defparam lut_465.mask = 64'h37ff37ff55575555;

	lut_sub lut_468 ({sk[124], i_27_, i_23_, i_24_, i_34_, x42x}, x273x);
	defparam lut_468.LUT_SIZE = 6;
	defparam lut_468.mask = 64'h37ff37ff10000000;

	lut_sub lut_470 ({sk[125], i_34_, i_36_, i_35_, i_29_, n_n1216}, x396x);
	defparam lut_470.LUT_SIZE = 6;
	defparam lut_470.mask = 64'h37ff37ff00000040;

	lut_sub lut_472 ({sk[126], i_8_, i_5_, i_6_, x219x}, x498x);
	defparam lut_472.LUT_SIZE = 5;
	defparam lut_472.mask = 32'h0f0f4000;

	lut_sub lut_474 ({sk[127], i_5_, i_4_, i_2_, n_n841, x326x}, x522x);
	defparam lut_474.LUT_SIZE = 6;
	defparam lut_474.mask = 64'h37ff37ff10000000;

	lut_sub lut_476 ({sk[128], i_9_, i_4_, x224x, n_n916, x363x}, x952x);
	defparam lut_476.LUT_SIZE = 6;
	defparam lut_476.mask = 64'h37ff37ff01000000;

	lut_sub lut_478 ({sk[129], i_13_, i_17_, x10x, x64x, x7769x}, x955x);
	defparam lut_478.LUT_SIZE = 6;
	defparam lut_478.mask = 64'h37ff37ff00000100;

	lut_sub lut_480 ({sk[130], x396x, x498x, x522x, x952x, x955x}, x7771x);
	defparam lut_480.LUT_SIZE = 6;
	defparam lut_480.mask = 64'h37ff37ff77777fff;

	lut_sub lut_485 ({sk[131], i_7_, x224x, x256x, x219x, x956x}, x7767x);
	defparam lut_485.LUT_SIZE = 6;
	defparam lut_485.mask = 64'h37ff37ff55575555;

	lut_sub lut_488 ({sk[132], i_10_, x43x, n_n82, x87x, x373x}, x7768x);
	defparam lut_488.LUT_SIZE = 6;
	defparam lut_488.mask = 64'h37ff37ff05370505;

	lut_sub lut_491 ({sk[133], i_13_, i_16_}, x43x);
	defparam lut_491.LUT_SIZE = 3;
	defparam lut_491.mask = 8'h58;

	lut_sub lut_493 ({sk[134], i_10_, i_7_, i_32_, i_36_, x64x}, x949x);
	defparam lut_493.LUT_SIZE = 6;
	defparam lut_493.mask = 64'h37ff37ff10000000;

	lut_sub lut_495 ({sk[135], x484x, x489x}, x7x);
	defparam lut_495.LUT_SIZE = 3;
	defparam lut_495.mask = 8'h57;

	lut_sub lut_498 ({sk[136], i_32_, i_36_, i_35_, i_29_, n_n1441}, x7779x);
	defparam lut_498.LUT_SIZE = 6;
	defparam lut_498.mask = 64'h37ff37ff00400000;

	lut_sub lut_500 ({sk[137], i_17_, x43x, x949x, x7x, x7779x}, x945x);
	defparam lut_500.LUT_SIZE = 6;
	defparam lut_500.mask = 64'h37ff37ff001f0000;

	lut_sub lut_503 ({sk[138], i_9_, n_n461, n_n301, x363x, x946x}, x944x);
	defparam lut_503.LUT_SIZE = 6;
	defparam lut_503.mask = 64'h37ff37ff00570000;

	lut_sub lut_506 ({sk[139], x42x, x498x, x522x, x368x, x942x}, x7780x);
	defparam lut_506.LUT_SIZE = 6;
	defparam lut_506.mask = 64'h37ff37ff55555777;

	lut_sub lut_510 ({sk[140], x7825x, n_n1566, x7852x, x906x, x7824x}, n_n1549);
	defparam lut_510.LUT_SIZE = 6;
	defparam lut_510.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_516 ({sk[141], n_n1561, n_n1563, x850x, x851x, x7880x}, n_n1548);
	defparam lut_516.LUT_SIZE = 6;
	defparam lut_516.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_522 ({sk[142], n_n1567, n_n1569, n_n1568}, x7922x);
	defparam lut_522.LUT_SIZE = 4;
	defparam lut_522.mask = 16'h777f;

	lut_sub lut_526 ({sk[143], n_n1556, x8074x, x8075x, x8076x}, x8079x);
	defparam lut_526.LUT_SIZE = 5;
	defparam lut_526.mask = 32'h0f0f7fff;

	lut_sub lut_531 ({sk[144], i_5_, i_4_, i_2_}, n_n1307);
	defparam lut_531.LUT_SIZE = 4;
	defparam lut_531.mask = 16'h7780;

	lut_sub lut_533 ({sk[145], i_7_, i_5_, i_6_}, n_n1278);
	defparam lut_533.LUT_SIZE = 4;
	defparam lut_533.mask = 16'h7780;

	lut_sub lut_535 ({sk[146], i_9_, i_7_, i_6_}, n_n1100);
	defparam lut_535.LUT_SIZE = 4;
	defparam lut_535.mask = 16'h7780;

	lut_sub lut_537 ({sk[147], i_9_, i_18_, x43x, x242x, n_n787}, x219x);
	defparam lut_537.LUT_SIZE = 6;
	defparam lut_537.mask = 64'h37ff37ff01000000;

	lut_sub lut_539 ({sk[148], i_11_, i_23_, i_17_, i_19_, x43x}, x326x);
	defparam lut_539.LUT_SIZE = 6;
	defparam lut_539.mask = 64'h37ff37ff40000000;

	lut_sub lut_541 ({sk[149], i_9_, i_8_, i_13_, n_n1278, n_n787}, n_n29);
	defparam lut_541.LUT_SIZE = 6;
	defparam lut_541.mask = 64'h37ff37ff10000000;

	lut_sub lut_543 ({sk[150], i_18_, i_17_, i_16_, n_n29}, x1766x);
	defparam lut_543.LUT_SIZE = 5;
	defparam lut_543.mask = 32'h0f0f4000;

	lut_sub lut_545 ({sk[151], i_17_, i_16_}, x263x);
	defparam lut_545.LUT_SIZE = 3;
	defparam lut_545.mask = 8'h58;

	lut_sub lut_547 ({sk[152], i_9_, i_13_, i_11_, n_n1307, n_n1303}, n_n129);
	defparam lut_547.LUT_SIZE = 6;
	defparam lut_547.mask = 64'h37ff37ff10000000;

	lut_sub lut_549 ({sk[153], i_11_, i_19_}, x204x);
	defparam lut_549.LUT_SIZE = 3;
	defparam lut_549.mask = 8'h58;

	lut_sub lut_551 ({sk[154], i_5_, i_6_, i_4_}, n_n461);
	defparam lut_551.LUT_SIZE = 4;
	defparam lut_551.mask = 16'h7780;

	lut_sub lut_553 ({sk[155], i_9_, i_5_, i_6_, i_4_}, x232x);
	defparam lut_553.LUT_SIZE = 5;
	defparam lut_553.mask = 32'h0f0f8000;

	lut_sub lut_555 ({sk[156], i_23_, i_21_}, x296x);
	defparam lut_555.LUT_SIZE = 3;
	defparam lut_555.mask = 8'h58;

	lut_sub lut_557 ({sk[157], i_27_, i_28_, i_23_}, n_n793);
	defparam lut_557.LUT_SIZE = 4;
	defparam lut_557.mask = 16'h7780;

	lut_sub lut_559 ({sk[158], i_34_, i_35_, i_29_, n_n793}, x378x);
	defparam lut_559.LUT_SIZE = 5;
	defparam lut_559.mask = 32'h0f0f0400;

	lut_sub lut_561 ({sk[159], i_27_, i_26_, i_24_, i_36_}, x79x);
	defparam lut_561.LUT_SIZE = 5;
	defparam lut_561.mask = 32'h0f0f4000;

	lut_sub lut_563 ({sk[160], i_13_, i_17_, i_16_}, n_n1443);
	defparam lut_563.LUT_SIZE = 4;
	defparam lut_563.mask = 16'h7780;

	lut_sub lut_565 ({sk[161], i_26_, i_24_}, x73x);
	defparam lut_565.LUT_SIZE = 3;
	defparam lut_565.mask = 8'h58;

	lut_sub lut_567 ({sk[162], i_28_, i_32_, i_29_}, n_n460);
	defparam lut_567.LUT_SIZE = 4;
	defparam lut_567.mask = 16'h7740;

	lut_sub lut_569 ({sk[163], i_27_, i_36_, n_n1443, x73x, n_n460}, x462x);
	defparam lut_569.LUT_SIZE = 6;
	defparam lut_569.mask = 64'h37ff37ff00010000;

	lut_sub lut_571 ({sk[164], i_27_, i_28_, i_29_}, n_n1375);
	defparam lut_571.LUT_SIZE = 4;
	defparam lut_571.mask = 16'h7780;

	lut_sub lut_573 ({sk[165], i_32_, i_34_, i_36_, i_35_}, x227x);
	defparam lut_573.LUT_SIZE = 5;
	defparam lut_573.mask = 32'h0f0f1000;

	lut_sub lut_575 ({sk[166], i_32_, i_34_, i_35_}, n_n1202);
	defparam lut_575.LUT_SIZE = 4;
	defparam lut_575.mask = 16'h7740;

	lut_sub lut_577 ({sk[167], i_27_, i_28_, i_36_, i_29_, n_n1202}, x493x);
	defparam lut_577.LUT_SIZE = 6;
	defparam lut_577.mask = 64'h37ff37ff04000000;

	lut_sub lut_579 ({sk[168], i_9_, i_6_}, x280x);
	defparam lut_579.LUT_SIZE = 3;
	defparam lut_579.mask = 8'h58;

	lut_sub lut_581 ({sk[169], i_5_, i_3_, i_4_, i_18_}, x338x);
	defparam lut_581.LUT_SIZE = 5;
	defparam lut_581.mask = 32'h0f0f0800;

	lut_sub lut_583 ({sk[170], i_7_, i_23_, x462x, x280x, x338x}, x102x);
	defparam lut_583.LUT_SIZE = 6;
	defparam lut_583.mask = 64'h37ff37ff01000000;

	lut_sub lut_585 ({sk[171], i_27_, i_28_, i_26_}, n_n1441);
	defparam lut_585.LUT_SIZE = 4;
	defparam lut_585.mask = 16'h7780;

	lut_sub lut_587 ({sk[172], i_32_, i_31_}, x302x);
	defparam lut_587.LUT_SIZE = 3;
	defparam lut_587.mask = 8'h58;

	lut_sub lut_589 ({sk[173], i_32_, i_31_, i_34_}, n_n1433);
	defparam lut_589.LUT_SIZE = 4;
	defparam lut_589.mask = 16'h7740;

	lut_sub lut_591 ({sk[174], i_30_, i_28_, i_26_}, n_n1425);
	defparam lut_591.LUT_SIZE = 4;
	defparam lut_591.mask = 16'h7780;

	lut_sub lut_593 ({sk[175], i_23_, i_24_}, x54x);
	defparam lut_593.LUT_SIZE = 3;
	defparam lut_593.mask = 8'h58;

	lut_sub lut_595 ({sk[176], i_25_, i_23_, i_24_}, n_n1396);
	defparam lut_595.LUT_SIZE = 4;
	defparam lut_595.mask = 16'h7708;

	lut_sub lut_597 ({sk[177], i_14_, i_12_, i_16_}, n_n1404);
	defparam lut_597.LUT_SIZE = 4;
	defparam lut_597.mask = 16'h7780;

	lut_sub lut_599 ({sk[178], i_23_, i_24_, i_16_}, n_n1390);
	defparam lut_599.LUT_SIZE = 4;
	defparam lut_599.mask = 16'h7780;

	lut_sub lut_601 ({sk[179], i_7_, i_14_, i_12_}, n_n1372);
	defparam lut_601.LUT_SIZE = 4;
	defparam lut_601.mask = 16'h7708;

	lut_sub lut_603 ({sk[180], i_27_, i_26_, i_24_}, n_n1369);
	defparam lut_603.LUT_SIZE = 4;
	defparam lut_603.mask = 16'h7780;

	lut_sub lut_605 ({sk[181], i_13_, i_12_, i_16_}, n_n1429);
	defparam lut_605.LUT_SIZE = 4;
	defparam lut_605.mask = 16'h7780;

	lut_sub lut_607 ({sk[182], i_25_, i_26_, i_24_}, n_n1454);
	defparam lut_607.LUT_SIZE = 4;
	defparam lut_607.mask = 16'h7780;

	lut_sub lut_609 ({sk[183], i_28_, i_29_}, x42x);
	defparam lut_609.LUT_SIZE = 3;
	defparam lut_609.mask = 8'h58;

	lut_sub lut_611 ({sk[184], i_9_, i_10_, i_8_}, n_n1353);
	defparam lut_611.LUT_SIZE = 4;
	defparam lut_611.mask = 16'h7708;

	lut_sub lut_613 ({sk[185], i_28_, i_25_, i_24_}, n_n1423);
	defparam lut_613.LUT_SIZE = 4;
	defparam lut_613.mask = 16'h7780;

	lut_sub lut_615 ({sk[186], i_34_, i_37_}, n_n1295);
	defparam lut_615.LUT_SIZE = 3;
	defparam lut_615.mask = 8'h51;

	lut_sub lut_617 ({sk[187], i_30_, i_32_}, x3x);
	defparam lut_617.LUT_SIZE = 3;
	defparam lut_617.mask = 8'h57;

	lut_sub lut_620 ({sk[188], i_30_, i_32_, i_31_}, n_n1438);
	defparam lut_620.LUT_SIZE = 4;
	defparam lut_620.mask = 16'h7780;

	lut_sub lut_622 ({sk[189], i_34_, i_35_}, n_n1397);
	defparam lut_622.LUT_SIZE = 3;
	defparam lut_622.mask = 8'h54;

	lut_sub lut_624 ({sk[190], i_23_, i_17_}, x242x);
	defparam lut_624.LUT_SIZE = 3;
	defparam lut_624.mask = 8'h58;

	lut_sub lut_626 ({sk[191], i_20_, i_23_, i_17_}, n_n1274);
	defparam lut_626.LUT_SIZE = 4;
	defparam lut_626.mask = 16'h7780;

	lut_sub lut_628 ({sk[192], i_31_, i_34_}, n_n1334);
	defparam lut_628.LUT_SIZE = 3;
	defparam lut_628.mask = 8'h51;

	lut_sub lut_630 ({sk[193], i_27_, i_28_, i_24_}, n_n1216);
	defparam lut_630.LUT_SIZE = 4;
	defparam lut_630.mask = 16'h7780;

	lut_sub lut_632 ({sk[194], i_13_, i_12_}, x290x);
	defparam lut_632.LUT_SIZE = 3;
	defparam lut_632.mask = 8'h58;

	lut_sub lut_634 ({sk[195], i_7_, i_13_, i_12_}, n_n1391);
	defparam lut_634.LUT_SIZE = 4;
	defparam lut_634.mask = 16'h7708;

	lut_sub lut_636 ({sk[196], i_28_, i_25_, i_26_}, n_n1478);
	defparam lut_636.LUT_SIZE = 4;
	defparam lut_636.mask = 16'h7780;

	lut_sub lut_638 ({sk[197], i_4_, i_2_}, x292x);
	defparam lut_638.LUT_SIZE = 3;
	defparam lut_638.mask = 8'h58;

	lut_sub lut_640 ({sk[198], i_34_, i_33_}, n_n1374);
	defparam lut_640.LUT_SIZE = 3;
	defparam lut_640.mask = 8'h51;

	lut_sub lut_642 ({sk[199], i_31_, i_34_, i_35_}, n_n1504);
	defparam lut_642.LUT_SIZE = 4;
	defparam lut_642.mask = 16'h7704;

	lut_sub lut_644 ({sk[200], i_9_, i_8_, i_6_}, n_n841);
	defparam lut_644.LUT_SIZE = 4;
	defparam lut_644.mask = 16'h7780;

	lut_sub lut_646 ({sk[201], i_9_, i_10_, i_6_}, n_n853);
	defparam lut_646.LUT_SIZE = 4;
	defparam lut_646.mask = 16'h7780;

	lut_sub lut_648 ({sk[202], i_9_, i_7_, i_12_}, n_n1315);
	defparam lut_648.LUT_SIZE = 4;
	defparam lut_648.mask = 16'h7720;

	lut_sub lut_650 ({sk[203], i_20_, i_23_, i_21_}, n_n1092);
	defparam lut_650.LUT_SIZE = 4;
	defparam lut_650.mask = 16'h7708;

	lut_sub lut_652 ({sk[204], i_27_, i_28_, i_29_}, n_n1406);
	defparam lut_652.LUT_SIZE = 4;
	defparam lut_652.mask = 16'h7740;

	lut_sub lut_654 ({sk[205], i_5_, i_6_}, x224x);
	defparam lut_654.LUT_SIZE = 3;
	defparam lut_654.mask = 8'h58;

	lut_sub lut_656 ({sk[206], i_3_, i_4_, i_2_}, n_n787);
	defparam lut_656.LUT_SIZE = 4;
	defparam lut_656.mask = 16'h7708;

	lut_sub lut_658 ({sk[207], i_30_, i_32_, i_33_, i_35_, i_38_}, n_n762);
	defparam lut_658.LUT_SIZE = 6;
	defparam lut_658.mask = 64'h37ff37ff40000000;

	lut_sub lut_660 ({sk[208], i_13_, i_12_, i_19_}, n_n582);
	defparam lut_660.LUT_SIZE = 4;
	defparam lut_660.mask = 16'h7710;

	lut_sub lut_662 ({sk[209], i_9_, i_8_, i_3_}, n_n1038);
	defparam lut_662.LUT_SIZE = 4;
	defparam lut_662.mask = 16'h7708;

	lut_sub lut_664 ({sk[210], i_13_, i_23_, i_16_}, n_n1314);
	defparam lut_664.LUT_SIZE = 4;
	defparam lut_664.mask = 16'h7780;

	lut_sub lut_666 ({sk[211], i_7_, i_8_}, x13x);
	defparam lut_666.LUT_SIZE = 3;
	defparam lut_666.mask = 8'h58;

	lut_sub lut_668 ({sk[212], i_7_, i_8_, i_12_}, n_n1141);
	defparam lut_668.LUT_SIZE = 4;
	defparam lut_668.mask = 16'h7780;

	lut_sub lut_670 ({sk[213], i_5_, i_6_, i_4_, i_12_, i_2_}, x11x);
	defparam lut_670.LUT_SIZE = 6;
	defparam lut_670.mask = 64'h37ff37ff80000000;

	lut_sub lut_672 ({sk[214], i_13_, i_23_, i_24_, i_16_, x11x}, n_n544);
	defparam lut_672.LUT_SIZE = 6;
	defparam lut_672.mask = 64'h37ff37ff40000000;

	lut_sub lut_674 ({sk[215], i_28_, i_26_, i_29_}, n_n1486);
	defparam lut_674.LUT_SIZE = 4;
	defparam lut_674.mask = 16'h7780;

	lut_sub lut_676 ({sk[216], i_14_, i_17_, i_16_}, n_n1408);
	defparam lut_676.LUT_SIZE = 4;
	defparam lut_676.mask = 16'h7780;

	lut_sub lut_678 ({sk[217], i_33_, i_35_, i_37_}, n_n504);
	defparam lut_678.LUT_SIZE = 4;
	defparam lut_678.mask = 16'h7740;

	lut_sub lut_680 ({sk[218], i_9_, i_7_, i_5_, i_6_, n_n787}, x60x);
	defparam lut_680.LUT_SIZE = 6;
	defparam lut_680.mask = 64'h37ff37ff40000000;

	lut_sub lut_682 ({sk[219], i_9_, i_7_, i_18_, x224x, n_n787}, x297x);
	defparam lut_682.LUT_SIZE = 6;
	defparam lut_682.mask = 64'h37ff37ff10000000;

	lut_sub lut_684 ({sk[220], i_32_, i_29_}, x243x);
	defparam lut_684.LUT_SIZE = 3;
	defparam lut_684.mask = 8'h58;

	lut_sub lut_686 ({sk[221], i_32_, i_33_, i_29_}, n_n1305);
	defparam lut_686.LUT_SIZE = 4;
	defparam lut_686.mask = 16'h7780;

	lut_sub lut_688 ({sk[222], i_8_, i_5_, i_6_}, n_n1118);
	defparam lut_688.LUT_SIZE = 4;
	defparam lut_688.mask = 16'h7780;

	lut_sub lut_690 ({sk[223], i_4_, i_1_, i_2_}, n_n1279);
	defparam lut_690.LUT_SIZE = 4;
	defparam lut_690.mask = 16'h7780;

	lut_sub lut_692 ({sk[224], i_7_, i_5_, i_6_, n_n1408, n_n1279}, n_n358);
	defparam lut_692.LUT_SIZE = 6;
	defparam lut_692.mask = 64'h37ff37ff10000000;

	lut_sub lut_694 ({sk[225], i_9_, i_13_, i_18_}, n_n1048);
	defparam lut_694.LUT_SIZE = 4;
	defparam lut_694.mask = 16'h7704;

	lut_sub lut_696 ({sk[226], i_8_, i_6_, i_12_, n_n1307}, x76x);
	defparam lut_696.LUT_SIZE = 5;
	defparam lut_696.mask = 32'h0f0f4000;

	lut_sub lut_698 ({sk[227], i_9_, i_13_, i_18_, x76x}, n_n307);
	defparam lut_698.LUT_SIZE = 5;
	defparam lut_698.mask = 32'h0f0f0010;

	lut_sub lut_700 ({sk[228], i_14_, i_23_, i_16_}, n_n1263);
	defparam lut_700.LUT_SIZE = 4;
	defparam lut_700.mask = 16'h7780;

	lut_sub lut_702 ({sk[229], i_7_, i_6_, i_12_}, n_n1306);
	defparam lut_702.LUT_SIZE = 4;
	defparam lut_702.mask = 16'h7780;

	lut_sub lut_704 ({sk[230], i_5_, i_4_, i_2_, n_n1306}, x321x);
	defparam lut_704.LUT_SIZE = 5;
	defparam lut_704.mask = 32'h0f0f4000;

	lut_sub lut_706 ({sk[231], i_14_, i_23_, i_16_, n_n1307, n_n1306}, n_n620);
	defparam lut_706.LUT_SIZE = 6;
	defparam lut_706.mask = 64'h37ff37ff10000000;

	lut_sub lut_708 ({sk[232], i_28_, i_32_, i_29_}, n_n1288);
	defparam lut_708.LUT_SIZE = 4;
	defparam lut_708.mask = 16'h7780;

	lut_sub lut_710 ({sk[233], i_27_, i_23_, i_24_}, n_n1018);
	defparam lut_710.LUT_SIZE = 4;
	defparam lut_710.mask = 16'h7780;

	lut_sub lut_712 ({sk[234], i_3_, i_13_, i_4_, i_12_, i_2_}, x213x);
	defparam lut_712.LUT_SIZE = 6;
	defparam lut_712.mask = 64'h37ff37ff80000000;

	lut_sub lut_714 ({sk[235], i_9_, i_5_, i_6_, i_11_}, x7425x);
	defparam lut_714.LUT_SIZE = 5;
	defparam lut_714.mask = 32'h0f0f0040;

	lut_sub lut_716 ({sk[236], i_13_, i_17_, i_16_, n_n1278, n_n1279}, n_n458);
	defparam lut_716.LUT_SIZE = 6;
	defparam lut_716.mask = 64'h37ff37ff10000000;

	lut_sub lut_718 ({sk[237], i_3_, i_4_, i_1_, i_2_, x224x}, x208x);
	defparam lut_718.LUT_SIZE = 6;
	defparam lut_718.mask = 64'h37ff37ff40000000;

	lut_sub lut_720 ({sk[238], i_9_, i_13_, i_11_, x208x}, n_n372);
	defparam lut_720.LUT_SIZE = 5;
	defparam lut_720.mask = 32'h0f0f0010;

	lut_sub lut_722 ({sk[239], i_32_, i_35_, i_38_}, n_n1179);
	defparam lut_722.LUT_SIZE = 4;
	defparam lut_722.mask = 16'h7740;

	lut_sub lut_724 ({sk[240], i_28_, i_25_, i_26_, i_24_, i_22_}, x257x);
	defparam lut_724.LUT_SIZE = 6;
	defparam lut_724.mask = 64'h37ff37ff80000000;

	lut_sub lut_726 ({sk[241], i_32_, i_35_, i_38_, x257x}, n_n300);
	defparam lut_726.LUT_SIZE = 5;
	defparam lut_726.mask = 32'h0f0f1000;

	lut_sub lut_728 ({sk[242], i_28_, i_34_, i_29_}, n_n1225);
	defparam lut_728.LUT_SIZE = 4;
	defparam lut_728.mask = 16'h7720;

	lut_sub lut_730 ({sk[243], i_9_, i_13_, i_19_, x208x}, n_n294);
	defparam lut_730.LUT_SIZE = 5;
	defparam lut_730.mask = 32'h0f0f0010;

	lut_sub lut_732 ({sk[244], i_10_, i_13_, i_16_}, n_n301);
	defparam lut_732.LUT_SIZE = 4;
	defparam lut_732.mask = 16'h7780;

	lut_sub lut_734 ({sk[245], i_5_, i_6_, i_4_, i_1_, i_2_}, x51x);
	defparam lut_734.LUT_SIZE = 6;
	defparam lut_734.mask = 64'h37ff37ff80000000;

	lut_sub lut_736 ({sk[246], i_23_, i_17_, i_16_}, n_n1322);
	defparam lut_736.LUT_SIZE = 4;
	defparam lut_736.mask = 16'h7780;

	lut_sub lut_738 ({sk[247], i_14_, i_23_, i_17_, i_16_}, x260x);
	defparam lut_738.LUT_SIZE = 5;
	defparam lut_738.mask = 32'h0f0f8000;

	lut_sub lut_740 ({sk[248], i_14_, i_23_, i_17_, i_16_, x51x}, n_n437);
	defparam lut_740.LUT_SIZE = 6;
	defparam lut_740.mask = 64'h37ff37ff40000000;

	lut_sub lut_742 ({sk[249], i_17_, i_21_, i_16_}, n_n825);
	defparam lut_742.LUT_SIZE = 4;
	defparam lut_742.mask = 16'h7780;

	lut_sub lut_744 ({sk[250], i_34_, i_33_, i_35_}, n_n1437);
	defparam lut_744.LUT_SIZE = 4;
	defparam lut_744.mask = 16'h7708;

	lut_sub lut_746 ({sk[251], i_32_, i_34_, i_33_}, n_n1340);
	defparam lut_746.LUT_SIZE = 4;
	defparam lut_746.mask = 16'h7720;

	lut_sub lut_748 ({sk[252], i_18_, i_17_, i_16_}, n_n132);
	defparam lut_748.LUT_SIZE = 4;
	defparam lut_748.mask = 16'h7780;

	lut_sub lut_750 ({sk[253], i_4_, i_1_, i_0_}, n_n152);
	defparam lut_750.LUT_SIZE = 4;
	defparam lut_750.mask = 16'h7780;

	lut_sub lut_752 ({sk[254], i_33_, i_38_}, n_n1300);
	defparam lut_752.LUT_SIZE = 3;
	defparam lut_752.mask = 8'h54;

	lut_sub lut_754 ({sk[255], i_30_, i_32_, i_29_}, n_n1472);
	defparam lut_754.LUT_SIZE = 4;
	defparam lut_754.mask = 16'h7780;

	lut_sub lut_756 ({sk[256], i_9_, i_6_, i_13_, n_n1307, x13x}, x261x);
	defparam lut_756.LUT_SIZE = 6;
	defparam lut_756.mask = 64'h37ff37ff01000000;

	lut_sub lut_758 ({sk[257], i_7_, i_8_, i_6_}, n_n1303);
	defparam lut_758.LUT_SIZE = 4;
	defparam lut_758.mask = 16'h7780;

	lut_sub lut_760 ({sk[258], i_9_, i_13_, i_24_, n_n1307, n_n1303}, n_n928);
	defparam lut_760.LUT_SIZE = 6;
	defparam lut_760.mask = 64'h37ff37ff00100000;

	lut_sub lut_762 ({sk[259], i_8_, i_5_, i_6_, i_1_, x292x}, x50x);
	defparam lut_762.LUT_SIZE = 6;
	defparam lut_762.mask = 64'h37ff37ff40000000;

	lut_sub lut_764 ({sk[260], i_28_, i_25_, i_26_, i_24_, i_22_}, x52x);
	defparam lut_764.LUT_SIZE = 6;
	defparam lut_764.mask = 64'h37ff37ff80000000;

	lut_sub lut_766 ({sk[261], i_9_, i_7_, i_6_, n_n1307}, x14x);
	defparam lut_766.LUT_SIZE = 5;
	defparam lut_766.mask = 32'h0f0f4000;

	lut_sub lut_768 ({sk[262], i_9_, i_7_, i_8_, i_6_, n_n1307}, x15x);
	defparam lut_768.LUT_SIZE = 6;
	defparam lut_768.mask = 64'h37ff37ff40000000;

	lut_sub lut_770 ({sk[263], i_9_, i_10_, i_6_, n_n1307, x13x}, x223x);
	defparam lut_770.LUT_SIZE = 6;
	defparam lut_770.mask = 64'h37ff37ff10000000;

	lut_sub lut_772 ({sk[264], i_28_, i_24_, i_38_, n_n1437}, x237x);
	defparam lut_772.LUT_SIZE = 5;
	defparam lut_772.mask = 32'h0f0f1000;

	lut_sub lut_774 ({sk[265], i_31_, i_35_, i_38_}, x264x);
	defparam lut_774.LUT_SIZE = 4;
	defparam lut_774.mask = 16'h7740;

	lut_sub lut_776 ({sk[266], i_34_, i_38_}, x266x);
	defparam lut_776.LUT_SIZE = 3;
	defparam lut_776.mask = 8'h51;

	lut_sub lut_778 ({sk[267], i_28_, i_26_, i_24_, i_22_}, x61x);
	defparam lut_778.LUT_SIZE = 5;
	defparam lut_778.mask = 32'h0f0f8000;

	lut_sub lut_780 ({sk[268], i_28_, i_26_, i_24_}, n_n1497);
	defparam lut_780.LUT_SIZE = 4;
	defparam lut_780.mask = 16'h7780;

	lut_sub lut_782 ({sk[269], i_22_, i_33_, i_38_, n_n1497}, x388x);
	defparam lut_782.LUT_SIZE = 5;
	defparam lut_782.mask = 32'h0f0f1000;

	lut_sub lut_784 ({sk[270], i_10_, i_24_, i_22_}, n_n1191);
	defparam lut_784.LUT_SIZE = 4;
	defparam lut_784.mask = 16'h7780;

	lut_sub lut_786 ({sk[271], i_10_, i_28_, i_26_, i_24_, i_22_}, x518x);
	defparam lut_786.LUT_SIZE = 6;
	defparam lut_786.mask = 64'h37ff37ff80000000;

	lut_sub lut_788 ({sk[272], i_9_, i_3_, i_13_, i_11_}, x262x);
	defparam lut_788.LUT_SIZE = 5;
	defparam lut_788.mask = 32'h0f0f0040;

	lut_sub lut_790 ({sk[273], i_9_, i_3_, i_11_}, n_n1058);
	defparam lut_790.LUT_SIZE = 4;
	defparam lut_790.mask = 16'h7704;

	lut_sub lut_792 ({sk[274], i_9_, i_3_, i_13_, i_18_}, x18x);
	defparam lut_792.LUT_SIZE = 5;
	defparam lut_792.mask = 32'h0f0f00c4;

	lut_sub lut_795 ({sk[275], i_9_, i_13_, i_11_, i_18_}, x436x);
	defparam lut_795.LUT_SIZE = 5;
	defparam lut_795.mask = 32'h0f0f0010;

	lut_sub lut_797 ({sk[276], i_13_, i_19_, n_n1058, x18x, x436x}, x529x);
	defparam lut_797.LUT_SIZE = 6;
	defparam lut_797.mask = 64'h37ff37ff5f7f5577;

	lut_sub lut_801 ({sk[277], i_32_, i_33_, i_38_, x14x, x518x}, x1216x);
	defparam lut_801.LUT_SIZE = 6;
	defparam lut_801.mask = 64'h37ff37ff01000000;

	lut_sub lut_803 ({sk[278], i_32_, i_31_, n_n1361, x51x, x52x}, x1217x);
	defparam lut_803.LUT_SIZE = 6;
	defparam lut_803.mask = 64'h37ff37ff01000000;

	lut_sub lut_805 ({sk[279], n_n1472, x237x, x529x, x1216x, x1217x}, x7513x);
	defparam lut_805.LUT_SIZE = 6;
	defparam lut_805.mask = 64'h37ff37ff7777777f;

	lut_sub lut_809 ({sk[280], i_28_, i_25_, i_34_, i_38_, i_29_}, x7509x);
	defparam lut_809.LUT_SIZE = 6;
	defparam lut_809.mask = 64'h37ff37ff02000000;

	lut_sub lut_811 ({sk[281], i_31_, i_35_, i_38_, x257x, x50x}, x1219x);
	defparam lut_811.LUT_SIZE = 6;
	defparam lut_811.mask = 64'h37ff37ff01000000;

	lut_sub lut_813 ({sk[282], n_n928, x223x, x388x, x7509x, x1219x}, x7514x);
	defparam lut_813.LUT_SIZE = 6;
	defparam lut_813.mask = 64'h37ff37ff555f777f;

	lut_sub lut_817 ({sk[283], i_7_, i_13_, i_12_}, n_n1147);
	defparam lut_817.LUT_SIZE = 4;
	defparam lut_817.mask = 16'h7780;

	lut_sub lut_819 ({sk[284], i_7_, i_14_, i_12_}, n_n1089);
	defparam lut_819.LUT_SIZE = 4;
	defparam lut_819.mask = 16'h7780;

	lut_sub lut_821 ({sk[285], i_24_, i_34_}, x298x);
	defparam lut_821.LUT_SIZE = 3;
	defparam lut_821.mask = 8'h54;

	lut_sub lut_823 ({sk[286], i_16_, i_36_, n_n1441, x54x, n_n1472}, x362x);
	defparam lut_823.LUT_SIZE = 6;
	defparam lut_823.mask = 64'h37ff37ff00010000;

	lut_sub lut_825 ({sk[287], i_30_, i_34_, i_36_, i_29_, n_n1216}, x374x);
	defparam lut_825.LUT_SIZE = 6;
	defparam lut_825.mask = 64'h37ff37ff00040000;

	lut_sub lut_827 ({sk[288], i_27_, i_23_, i_24_, i_17_, x42x}, x48x);
	defparam lut_827.LUT_SIZE = 6;
	defparam lut_827.mask = 64'h37ff37ff40000000;

	lut_sub lut_829 ({sk[289], i_34_, i_36_}, x244x);
	defparam lut_829.LUT_SIZE = 3;
	defparam lut_829.mask = 8'h51;

	lut_sub lut_831 ({sk[290], i_30_, i_7_, i_32_, x48x, x244x}, x410x);
	defparam lut_831.LUT_SIZE = 6;
	defparam lut_831.mask = 64'h37ff37ff10000000;

	lut_sub lut_833 ({sk[291], i_30_, i_32_, n_n1375, n_n1390, x244x}, x467x);
	defparam lut_833.LUT_SIZE = 6;
	defparam lut_833.mask = 64'h37ff37ff01000000;

	lut_sub lut_835 ({sk[292], i_23_, i_24_, i_17_, n_n1441}, x74x);
	defparam lut_835.LUT_SIZE = 5;
	defparam lut_835.mask = 32'h0f0f4000;

	lut_sub lut_837 ({sk[293], i_7_, i_36_, i_29_, x3x, x74x}, x516x);
	defparam lut_837.LUT_SIZE = 6;
	defparam lut_837.mask = 64'h37ff37ff00400000;

	lut_sub lut_839 ({sk[294], i_12_, n_n1489, x13x, n_n1263, x260x}, x531x);
	defparam lut_839.LUT_SIZE = 6;
	defparam lut_839.mask = 64'h37ff37ff00070005;

	lut_sub lut_842 ({sk[295], i_13_, i_12_, i_23_, i_16_, x13x}, x323x);
	defparam lut_842.LUT_SIZE = 6;
	defparam lut_842.mask = 64'h37ff37ff40000000;

	lut_sub lut_844 ({sk[296], i_7_, i_8_, i_13_, i_16_, x242x}, x291x);
	defparam lut_844.LUT_SIZE = 6;
	defparam lut_844.mask = 64'h37ff37ff40000000;

	lut_sub lut_846 ({sk[297], i_13_, i_23_, i_16_, n_n1141, x291x}, x530x);
	defparam lut_846.LUT_SIZE = 6;
	defparam lut_846.mask = 64'h37ff37ff75555555;

	lut_sub lut_849 ({sk[298], i_28_, i_29_, n_n1438, n_n1092, x298x}, x933x);
	defparam lut_849.LUT_SIZE = 6;
	defparam lut_849.mask = 64'h37ff37ff00010000;

	lut_sub lut_851 ({sk[299], x79x, x374x, x531x, x530x, x933x}, x7796x);
	defparam lut_851.LUT_SIZE = 6;
	defparam lut_851.mask = 64'h37ff37ff55775f7f;

	lut_sub lut_855 ({sk[300], i_14_, i_16_, n_n1147, x467x, x516x}, x9206x);
	defparam lut_855.LUT_SIZE = 6;
	defparam lut_855.mask = 64'h37ff37ffa8fcfcfc;

	lut_sub lut_862 ({sk[301], x43x, n_n1089, x362x, x410x, x9206x}, x7797x);
	defparam lut_862.LUT_SIZE = 6;
	defparam lut_862.mask = 64'h37ff37ffaaafbbbf;

	lut_sub lut_866 ({sk[302], i_28_, i_34_, i_29_}, n_n1326);
	defparam lut_866.LUT_SIZE = 4;
	defparam lut_866.mask = 16'h7740;

	lut_sub lut_868 ({sk[303], i_20_, i_34_, i_29_, x296x, n_n1216}, x209x);
	defparam lut_868.LUT_SIZE = 6;
	defparam lut_868.mask = 64'h37ff37ff00000001;

	lut_sub lut_870 ({sk[304], i_23_, i_24_, i_21_}, n_n1312);
	defparam lut_870.LUT_SIZE = 4;
	defparam lut_870.mask = 16'h7740;

	lut_sub lut_872 ({sk[305], i_23_, i_24_, i_21_, i_34_}, x245x);
	defparam lut_872.LUT_SIZE = 5;
	defparam lut_872.mask = 32'h0f0f1000;

	lut_sub lut_874 ({sk[306], i_30_, i_28_}, x277x);
	defparam lut_874.LUT_SIZE = 3;
	defparam lut_874.mask = 8'h58;

	lut_sub lut_876 ({sk[307], i_28_, i_31_, i_34_}, n_n1511);
	defparam lut_876.LUT_SIZE = 4;
	defparam lut_876.mask = 16'h7710;

	lut_sub lut_878 ({sk[308], i_27_, i_23_, i_24_, i_21_, n_n1511}, x300x);
	defparam lut_878.LUT_SIZE = 6;
	defparam lut_878.mask = 64'h37ff37ff10000000;

	lut_sub lut_880 ({sk[309], i_32_, i_31_, i_33_}, n_n1393);
	defparam lut_880.LUT_SIZE = 4;
	defparam lut_880.mask = 16'h7740;

	lut_sub lut_882 ({sk[310], i_14_, i_32_, i_31_, i_33_}, x340x);
	defparam lut_882.LUT_SIZE = 5;
	defparam lut_882.mask = 32'h0f0f0040;

	lut_sub lut_884 ({sk[311], i_20_, i_26_, i_23_, i_24_, n_n1406}, x222x);
	defparam lut_884.LUT_SIZE = 6;
	defparam lut_884.mask = 64'h37ff37ff40000000;

	lut_sub lut_886 ({sk[312], i_26_, i_23_, i_24_}, n_n1213);
	defparam lut_886.LUT_SIZE = 4;
	defparam lut_886.mask = 16'h7780;

	lut_sub lut_888 ({sk[313], i_20_, i_2_, i_21_, n_n1406, n_n1213}, x432x);
	defparam lut_888.LUT_SIZE = 6;
	defparam lut_888.mask = 64'h37ff37ff00100000;

	lut_sub lut_890 ({sk[314], i_20_, i_21_, x73x, n_n1438, n_n1326}, x924x);
	defparam lut_890.LUT_SIZE = 6;
	defparam lut_890.mask = 64'h37ff37ff00000100;

	lut_sub lut_892 ({sk[315], i_7_, i_8_, i_14_, n_n1322, x374x}, x925x);
	defparam lut_892.LUT_SIZE = 6;
	defparam lut_892.mask = 64'h37ff37ff10000000;

	lut_sub lut_894 ({sk[316], i_12_, x10x, x432x, x924x, x925x}, x7808x);
	defparam lut_894.LUT_SIZE = 6;
	defparam lut_894.mask = 64'h37ff37ff777f7777;

	lut_sub lut_898 ({sk[317], i_30_, i_28_, i_34_, n_n1312, x340x}, x926x);
	defparam lut_898.LUT_SIZE = 6;
	defparam lut_898.mask = 64'h37ff37ff01000000;

	lut_sub lut_900 ({sk[318], x43x, n_n1315, x263x, x300x, n_n1323}, x927x);
	defparam lut_900.LUT_SIZE = 6;
	defparam lut_900.mask = 64'h37ff37ff01010133;

	lut_sub lut_903 ({sk[319], i_13_, i_12_, i_17_, i_16_, x209x}, x928x);
	defparam lut_903.LUT_SIZE = 6;
	defparam lut_903.mask = 64'h37ff37ff44400000;

	lut_sub lut_906 ({sk[320], x10x, x410x, x926x, x927x, x928x}, x7809x);
	defparam lut_906.LUT_SIZE = 6;
	defparam lut_906.mask = 64'h37ff37ff7f7f7fff;

	lut_sub lut_911 ({sk[321], i_27_, i_28_, i_24_, i_29_}, x80x);
	defparam lut_911.LUT_SIZE = 5;
	defparam lut_911.mask = 32'h0f0f8000;

	lut_sub lut_913 ({sk[322], i_9_, i_7_, i_14_}, n_n1285);
	defparam lut_913.LUT_SIZE = 4;
	defparam lut_913.mask = 16'h7720;

	lut_sub lut_915 ({sk[323], i_23_, x10x, n_n1315, n_n1322, n_n1285}, x535x);
	defparam lut_915.LUT_SIZE = 6;
	defparam lut_915.mask = 64'h37ff37ff111f1111;

	lut_sub lut_918 ({sk[324], i_28_, i_33_, i_29_}, n_n1257);
	defparam lut_918.LUT_SIZE = 4;
	defparam lut_918.mask = 16'h7720;

	lut_sub lut_920 ({sk[325], i_27_, i_25_, i_23_, n_n1397, n_n1257}, x82x);
	defparam lut_920.LUT_SIZE = 6;
	defparam lut_920.mask = 64'h37ff37ff00100000;

	lut_sub lut_922 ({sk[326], i_12_, x10x, n_n1312, x82x, x485x}, x916x);
	defparam lut_922.LUT_SIZE = 6;
	defparam lut_922.mask = 64'h37ff37ff00370000;

	lut_sub lut_925 ({sk[327], i_13_, i_12_, i_16_, x432x, x916x}, x7814x);
	defparam lut_925.LUT_SIZE = 6;
	defparam lut_925.mask = 64'h37ff37ff75555555;

	lut_sub lut_928 ({sk[328], i_12_, i_17_}, x240x);
	defparam lut_928.LUT_SIZE = 3;
	defparam lut_928.mask = 8'h51;

	lut_sub lut_930 ({sk[329], i_12_, i_24_, i_17_}, n_n1519);
	defparam lut_930.LUT_SIZE = 4;
	defparam lut_930.mask = 16'h7704;

	lut_sub lut_932 ({sk[330], i_28_, i_33_, i_29_}, n_n1302);
	defparam lut_932.LUT_SIZE = 4;
	defparam lut_932.mask = 16'h7780;

	lut_sub lut_934 ({sk[331], i_7_, i_13_, i_16_}, n_n1401);
	defparam lut_934.LUT_SIZE = 4;
	defparam lut_934.mask = 16'h7708;

	lut_sub lut_936 ({sk[332], i_9_, i_8_, i_2_}, n_n1192);
	defparam lut_936.LUT_SIZE = 4;
	defparam lut_936.mask = 16'h7708;

	lut_sub lut_938 ({sk[333], i_9_, i_7_, i_13_}, n_n1323);
	defparam lut_938.LUT_SIZE = 4;
	defparam lut_938.mask = 16'h7720;

	lut_sub lut_940 ({sk[334], i_32_, i_31_, i_29_}, n_n1133);
	defparam lut_940.LUT_SIZE = 4;
	defparam lut_940.mask = 16'h7780;

	lut_sub lut_942 ({sk[335], i_28_, i_31_, i_29_}, n_n1128);
	defparam lut_942.LUT_SIZE = 4;
	defparam lut_942.mask = 16'h7780;

	lut_sub lut_944 ({sk[336], i_13_, i_12_, i_11_}, n_n586);
	defparam lut_944.LUT_SIZE = 4;
	defparam lut_944.mask = 16'h7710;

	lut_sub lut_946 ({sk[337], i_26_, i_24_, i_22_}, n_n1523);
	defparam lut_946.LUT_SIZE = 4;
	defparam lut_946.mask = 16'h7780;

	lut_sub lut_948 ({sk[338], i_13_, i_23_, i_16_, n_n1307, n_n1306}, n_n269);
	defparam lut_948.LUT_SIZE = 6;
	defparam lut_948.mask = 64'h37ff37ff10000000;

	lut_sub lut_950 ({sk[339], i_8_, i_13_, i_16_}, x259x);
	defparam lut_950.LUT_SIZE = 4;
	defparam lut_950.mask = 16'h7780;

	lut_sub lut_952 ({sk[340], i_7_, i_5_, i_6_, n_n1279, x259x}, n_n242);
	defparam lut_952.LUT_SIZE = 6;
	defparam lut_952.mask = 64'h37ff37ff10000000;

	lut_sub lut_954 ({sk[341], i_8_, i_14_, i_16_, n_n1278, n_n1279}, n_n355);
	defparam lut_954.LUT_SIZE = 6;
	defparam lut_954.mask = 64'h37ff37ff10000000;

	lut_sub lut_956 ({sk[342], i_30_, i_28_, i_31_}, n_n1345);
	defparam lut_956.LUT_SIZE = 4;
	defparam lut_956.mask = 16'h7780;

	lut_sub lut_958 ({sk[343], i_9_, i_5_, i_6_, i_1_, x292x}, x229x);
	defparam lut_958.LUT_SIZE = 6;
	defparam lut_958.mask = 64'h37ff37ff00004000;

	lut_sub lut_960 ({sk[344], i_13_, i_11_, i_18_, x229x}, n_n371);
	defparam lut_960.LUT_SIZE = 5;
	defparam lut_960.mask = 32'h0f0f0100;

	lut_sub lut_962 ({sk[345], i_22_, i_33_, i_35_, i_38_, x73x}, x389x);
	defparam lut_962.LUT_SIZE = 6;
	defparam lut_962.mask = 64'h37ff37ff10000000;

	lut_sub lut_964 ({sk[346], i_28_, i_33_, i_35_, i_38_, n_n1523}, x53x);
	defparam lut_964.LUT_SIZE = 6;
	defparam lut_964.mask = 64'h37ff37ff10000000;

	lut_sub lut_966 ({sk[347], i_13_, i_18_, i_19_}, n_n735);
	defparam lut_966.LUT_SIZE = 4;
	defparam lut_966.mask = 16'h7710;

	lut_sub lut_968 ({sk[348], i_9_, i_13_, i_18_, i_19_, x11x}, n_n315);
	defparam lut_968.LUT_SIZE = 6;
	defparam lut_968.mask = 64'h37ff37ff00000100;

	lut_sub lut_970 ({sk[349], i_27_, i_28_, i_31_}, n_n984);
	defparam lut_970.LUT_SIZE = 4;
	defparam lut_970.mask = 16'h7740;

	lut_sub lut_972 ({sk[350], i_32_, i_33_, i_35_}, n_n1458);
	defparam lut_972.LUT_SIZE = 4;
	defparam lut_972.mask = 16'h7780;

	lut_sub lut_974 ({sk[351], i_34_, i_33_, i_29_}, n_n1241);
	defparam lut_974.LUT_SIZE = 4;
	defparam lut_974.mask = 16'h7708;

	lut_sub lut_976 ({sk[352], i_5_, i_4_, i_0_}, n_n245);
	defparam lut_976.LUT_SIZE = 4;
	defparam lut_976.mask = 16'h7780;

	lut_sub lut_978 ({sk[353], i_30_, i_28_, i_32_}, n_n1431);
	defparam lut_978.LUT_SIZE = 4;
	defparam lut_978.mask = 16'h7780;

	lut_sub lut_980 ({sk[354], i_26_, i_23_, i_24_, n_n1406}, x46x);
	defparam lut_980.LUT_SIZE = 5;
	defparam lut_980.mask = 32'h0f0f4000;

	lut_sub lut_982 ({sk[355], i_20_, i_21_, i_22_}, x7491x);
	defparam lut_982.LUT_SIZE = 4;
	defparam lut_982.mask = 16'h7708;

	lut_sub lut_984 ({sk[356], i_26_, i_23_, i_24_, n_n1406, x7491x}, x62x);
	defparam lut_984.LUT_SIZE = 6;
	defparam lut_984.mask = 64'h37ff37ff10000000;

	lut_sub lut_986 ({sk[357], i_28_, i_22_, i_33_, i_38_, x73x}, x70x);
	defparam lut_986.LUT_SIZE = 6;
	defparam lut_986.mask = 64'h37ff37ff10000000;

	lut_sub lut_988 ({sk[358], i_7_, i_8_, i_6_, i_12_, n_n1307}, x72x);
	defparam lut_988.LUT_SIZE = 6;
	defparam lut_988.mask = 64'h37ff37ff40000000;

	lut_sub lut_990 ({sk[359], i_8_, i_24_, i_38_}, x7492x);
	defparam lut_990.LUT_SIZE = 4;
	defparam lut_990.mask = 16'h7740;

	lut_sub lut_992 ({sk[360], i_7_, i_5_, i_6_, n_n1279, x7492x}, x212x);
	defparam lut_992.LUT_SIZE = 6;
	defparam lut_992.mask = 64'h37ff37ff10000000;

	lut_sub lut_994 ({sk[361], i_24_, i_38_}, x9x);
	defparam lut_994.LUT_SIZE = 3;
	defparam lut_994.mask = 8'h54;

	lut_sub lut_996 ({sk[362], i_25_, i_24_, i_38_}, x239x);
	defparam lut_996.LUT_SIZE = 4;
	defparam lut_996.mask = 16'h7740;

	lut_sub lut_998 ({sk[363], i_7_, i_5_, i_6_, i_38_, n_n1279}, x250x);
	defparam lut_998.LUT_SIZE = 6;
	defparam lut_998.mask = 64'h37ff37ff10000000;

	lut_sub lut_1000 ({sk[364], i_28_, i_34_, i_33_, i_29_}, x288x);
	defparam lut_1000.LUT_SIZE = 5;
	defparam lut_1000.mask = 32'h0f0f0800;

	lut_sub lut_1002 ({sk[365], i_12_, i_32_, n_n1307, n_n1306, n_n1303}, x538x);
	defparam lut_1002.LUT_SIZE = 6;
	defparam lut_1002.mask = 64'h37ff37ff07050300;

	lut_sub lut_1005 ({sk[366], i_32_, i_34_, i_29_, n_n1423}, x476x);
	defparam lut_1005.LUT_SIZE = 5;
	defparam lut_1005.mask = 32'h0f0f0400;

	lut_sub lut_1007 ({sk[367], i_28_, i_24_, i_29_, n_n1340}, x477x);
	defparam lut_1007.LUT_SIZE = 5;
	defparam lut_1007.mask = 32'h0f0f4000;

	lut_sub lut_1009 ({sk[368], i_28_, n_n1241, x70x, x212x, x538x}, x7495x);
	defparam lut_1009.LUT_SIZE = 6;
	defparam lut_1009.mask = 64'h37ff37ff05370505;

	lut_sub lut_1012 ({sk[369], i_9_, i_10_, i_2_, x389x, n_n1431}, x1230x);
	defparam lut_1012.LUT_SIZE = 6;
	defparam lut_1012.mask = 64'h37ff37ff00001000;

	lut_sub lut_1014 ({sk[370], n_n1423, x250x, x477x, x7409x, x1234x}, x7494x);
	defparam lut_1014.LUT_SIZE = 6;
	defparam lut_1014.mask = 64'h37ff37ff555f557f;

	lut_sub lut_1018 ({sk[371], n_n1225, x72x, x239x, x1230x, x7494x}, x7496x);
	defparam lut_1018.LUT_SIZE = 6;
	defparam lut_1018.mask = 64'h37ff37ff7777777f;

	lut_sub lut_1022 ({sk[372], i_32_, i_36_, i_35_}, n_n576);
	defparam lut_1022.LUT_SIZE = 4;
	defparam lut_1022.mask = 16'h7720;

	lut_sub lut_1024 ({sk[373], i_28_, i_31_, i_29_}, n_n1499);
	defparam lut_1024.LUT_SIZE = 4;
	defparam lut_1024.mask = 16'h7720;

	lut_sub lut_1026 ({sk[374], i_9_, i_2_, x463x, x578x}, x902x);
	defparam lut_1026.LUT_SIZE = 5;
	defparam lut_1026.mask = 32'h0f0f0100;

	lut_sub lut_1028 ({sk[375], i_28_, i_36_, n_n1369, n_n355, n_n1282}, x907x);
	defparam lut_1028.LUT_SIZE = 6;
	defparam lut_1028.mask = 64'h37ff37ff00010000;

	lut_sub lut_1030 ({sk[376], n_n1307, n_n841, x221x, x367x, x384x}, x9211x);
	defparam lut_1030.LUT_SIZE = 6;
	defparam lut_1030.mask = 64'h37ff37fffcfcfca8;

	lut_sub lut_1037 ({sk[377], i_34_, n_n880, x902x, x907x, x9211x}, x7825x);
	defparam lut_1037.LUT_SIZE = 6;
	defparam lut_1037.mask = 64'h37ff37ff3f3f3fbf;

	lut_sub lut_1041 ({sk[378], i_23_, x493x, x10x, n_n1307, n_n1306}, x898x);
	defparam lut_1041.LUT_SIZE = 6;
	defparam lut_1041.mask = 64'h37ff37ff00010000;

	lut_sub lut_1043 ({sk[379], i_28_, i_36_, n_n1369, n_n242, n_n1282}, x899x);
	defparam lut_1043.LUT_SIZE = 6;
	defparam lut_1043.mask = 64'h37ff37ff00010000;

	lut_sub lut_1045 ({sk[380], n_n358, n_n1288, n_n1018, x48x, n_n355}, x9210x);
	defparam lut_1045.LUT_SIZE = 6;
	defparam lut_1045.mask = 64'h37ff37ffeeeeeee0;

	lut_sub lut_1052 ({sk[381], i_34_, i_36_, x898x, x899x, x9210x}, x7840x);
	defparam lut_1052.LUT_SIZE = 6;
	defparam lut_1052.mask = 64'h37ff37ff3f3f3fbf;

	lut_sub lut_1056 ({sk[382], x325x, x328x, x7830x, x894x}, x7836x);
	defparam lut_1056.LUT_SIZE = 5;
	defparam lut_1056.mask = 32'h0f0f5777;

	lut_sub lut_1060 ({sk[383], i_36_, x378x, n_n363, x895x}, x7837x);
	defparam lut_1060.LUT_SIZE = 5;
	defparam lut_1060.mask = 32'h0f0f5557;

	lut_sub lut_1063 ({sk[384], x7840x, x7836x, x7837x}, n_n1566);
	defparam lut_1063.LUT_SIZE = 4;
	defparam lut_1063.mask = 16'h777f;

	lut_sub lut_1067 ({sk[385], i_10_, i_7_, i_3_, i_18_}, x437x);
	defparam lut_1067.LUT_SIZE = 5;
	defparam lut_1067.mask = 32'h0f0f0002;

	lut_sub lut_1069 ({sk[386], i_10_, i_7_, i_11_, i_19_, x437x}, x16x);
	defparam lut_1069.LUT_SIZE = 6;
	defparam lut_1069.mask = 64'h37ff37ff555555d5;

	lut_sub lut_1072 ({sk[387], i_5_, i_4_, i_2_, n_n841}, x41x);
	defparam lut_1072.LUT_SIZE = 5;
	defparam lut_1072.mask = 32'h0f0f4000;

	lut_sub lut_1074 ({sk[388], i_23_, i_24_, i_17_, i_29_, n_n1441}, x458x);
	defparam lut_1074.LUT_SIZE = 6;
	defparam lut_1074.mask = 64'h37ff37ff40000000;

	lut_sub lut_1076 ({sk[389], i_29_, n_n1307, n_n841, x74x}, x217x);
	defparam lut_1076.LUT_SIZE = 5;
	defparam lut_1076.mask = 32'h0f0f0100;

	lut_sub lut_1078 ({sk[390], i_23_, i_24_, i_21_, n_n1441}, x228x);
	defparam lut_1078.LUT_SIZE = 5;
	defparam lut_1078.mask = 32'h0f0f4000;

	lut_sub lut_1080 ({sk[391], i_27_, i_28_, i_26_, i_29_}, x44x);
	defparam lut_1080.LUT_SIZE = 5;
	defparam lut_1080.mask = 32'h0f0f4000;

	lut_sub lut_1082 ({sk[392], i_23_, i_24_, i_21_}, x7749x);
	defparam lut_1082.LUT_SIZE = 4;
	defparam lut_1082.mask = 16'h7780;

	lut_sub lut_1084 ({sk[393], i_31_, n_n461, n_n576, x44x, x7749x}, x307x);
	defparam lut_1084.LUT_SIZE = 6;
	defparam lut_1084.mask = 64'h37ff37ff00010000;

	lut_sub lut_1086 ({sk[394], i_13_, i_12_, i_17_, i_16_, x9230x}, x882x);
	defparam lut_1086.LUT_SIZE = 6;
	defparam lut_1086.mask = 64'h37ff37ff88800000;

	lut_sub lut_1089 ({sk[395], i_21_, i_32_, i_36_, n_n1441, x54x}, x7845x);
	defparam lut_1089.LUT_SIZE = 6;
	defparam lut_1089.mask = 64'h37ff37ff01000000;

	lut_sub lut_1091 ({sk[396], n_n576, n_n329, x468x, x67x, x367x}, x885x);
	defparam lut_1091.LUT_SIZE = 6;
	defparam lut_1091.mask = 64'h37ff37ff0000111f;

	lut_sub lut_1094 ({sk[397], n_n1429, n_n301, n_n880, x217x, x307x}, x7850x);
	defparam lut_1094.LUT_SIZE = 6;
	defparam lut_1094.mask = 64'h37ff37ff00035557;

	lut_sub lut_1097 ({sk[398], n_n358, x882x, x7845x, x885x, x7850x}, x7852x);
	defparam lut_1097.LUT_SIZE = 6;
	defparam lut_1097.mask = 64'h37ff37ff77ff7fff;

	lut_sub lut_1102 ({sk[399], n_n576, x265x, x312x, x67x, x495x}, x906x);
	defparam lut_1102.LUT_SIZE = 6;
	defparam lut_1102.mask = 64'h37ff37ff00031113;

	lut_sub lut_1105 ({sk[400], i_36_, i_35_, x217x, n_n916, x903x}, x7824x);
	defparam lut_1105.LUT_SIZE = 6;
	defparam lut_1105.mask = 64'h37ff37ff55555755;

	lut_sub lut_1108 ({sk[401], i_9_, i_10_, i_13_, n_n1307, n_n1303}, n_n82);
	defparam lut_1108.LUT_SIZE = 6;
	defparam lut_1108.mask = 64'h37ff37ff10000000;

	lut_sub lut_1110 ({sk[402], i_14_, i_17_, i_16_, n_n1118, n_n1279}, n_n195);
	defparam lut_1110.LUT_SIZE = 6;
	defparam lut_1110.mask = 64'h37ff37ff10000000;

	lut_sub lut_1112 ({sk[403], i_23_, i_17_, i_16_, i_29_, n_n1216}, x391x);
	defparam lut_1112.LUT_SIZE = 6;
	defparam lut_1112.mask = 64'h37ff37ff40000000;

	lut_sub lut_1114 ({sk[404], i_13_, i_32_, x10x, x14x, x48x}, x147x);
	defparam lut_1114.LUT_SIZE = 6;
	defparam lut_1114.mask = 64'h37ff37ff00000100;

	lut_sub lut_1116 ({sk[405], i_14_, x261x, x244x, x391x, x147x}, x877x);
	defparam lut_1116.LUT_SIZE = 6;
	defparam lut_1116.mask = 64'h37ff37ff05070505;

	lut_sub lut_1119 ({sk[406], n_n825, n_n576, x881x, x7858x, x7859x}, x875x);
	defparam lut_1119.LUT_SIZE = 6;
	defparam lut_1119.mask = 64'h37ff37ff0000001f;

	lut_sub lut_1122 ({sk[407], x228x, x265x, x559x, x873x, x876x}, x7865x);
	defparam lut_1122.LUT_SIZE = 6;
	defparam lut_1122.mask = 64'h37ff37ff7777777f;

	lut_sub lut_1126 ({sk[408], x877x, x875x, x7865x}, n_n1561);
	defparam lut_1126.LUT_SIZE = 4;
	defparam lut_1126.mask = 16'h777f;

	lut_sub lut_1130 ({sk[409], i_34_, i_36_, i_35_, n_n1018, n_n1128}, x500x);
	defparam lut_1130.LUT_SIZE = 6;
	defparam lut_1130.mask = 64'h37ff37ff00000010;

	lut_sub lut_1132 ({sk[410], i_13_, i_17_, i_16_, n_n1118, n_n1279}, x312x);
	defparam lut_1132.LUT_SIZE = 6;
	defparam lut_1132.mask = 64'h37ff37ff10000000;

	lut_sub lut_1134 ({sk[411], n_n437, n_n576, x483x, n_n329, x468x}, x9209x);
	defparam lut_1134.LUT_SIZE = 6;
	defparam lut_1134.mask = 64'h37ff37fffcfcfca8;

	lut_sub lut_1141 ({sk[412], n_n1404, x307x, x500x, x312x, x9209x}, x7876x);
	defparam lut_1141.LUT_SIZE = 6;
	defparam lut_1141.mask = 64'h37ff37ffabababff;

	lut_sub lut_1145 ({sk[413], i_14_, n_n195, x265x, x67x, x501x}, x863x);
	defparam lut_1145.LUT_SIZE = 6;
	defparam lut_1145.mask = 64'h37ff37ff05070003;

	lut_sub lut_1148 ({sk[414], i_36_, x384x, x7868x, x871x, x872x}, x864x);
	defparam lut_1148.LUT_SIZE = 6;
	defparam lut_1148.mask = 64'h37ff37ff0000777f;

	lut_sub lut_1152 ({sk[415], x7876x, x863x, x864x}, n_n1563);
	defparam lut_1152.LUT_SIZE = 4;
	defparam lut_1152.mask = 16'h777f;

	lut_sub lut_1156 ({sk[416], i_23_, i_34_, i_35_, n_n984}, x275x);
	defparam lut_1156.LUT_SIZE = 5;
	defparam lut_1156.mask = 32'h0f0f1000;

	lut_sub lut_1158 ({sk[417], i_34_, i_36_, i_35_, n_n1216, n_n1133}, x483x);
	defparam lut_1158.LUT_SIZE = 6;
	defparam lut_1158.mask = 64'h37ff37ff00000010;

	lut_sub lut_1160 ({sk[418], i_14_, i_13_, i_16_, x48x, x41x}, x144x);
	defparam lut_1160.LUT_SIZE = 6;
	defparam lut_1160.mask = 64'h37ff37ff00100000;

	lut_sub lut_1162 ({sk[419], i_21_, n_n1443, n_n1429, x437x, x16x}, x856x);
	defparam lut_1162.LUT_SIZE = 6;
	defparam lut_1162.mask = 64'h37ff37ff00000537;

	lut_sub lut_1165 ({sk[420], i_17_, x43x, x275x, x856x, x440x}, x850x);
	defparam lut_1165.LUT_SIZE = 6;
	defparam lut_1165.mask = 64'h37ff37ff03070303;

	lut_sub lut_1168 ({sk[421], i_34_, n_n880, x144x, x221x, x495x}, x851x);
	defparam lut_1168.LUT_SIZE = 6;
	defparam lut_1168.mask = 64'h37ff37ff0000001f;

	lut_sub lut_1171 ({sk[422], n_n82, n_n195, x500x, x7878x, x853x}, x7880x);
	defparam lut_1171.LUT_SIZE = 6;
	defparam lut_1171.mask = 64'h37ff37ff555f777f;

	lut_sub lut_1175 ({sk[423], n_n458, n_n355, x458x, x846x, x7889x}, x609x);
	defparam lut_1175.LUT_SIZE = 6;
	defparam lut_1175.mask = 64'h37ff37ff333f777f;

	lut_sub lut_1179 ({sk[424], i_23_, i_21_, n_n1334, n_n1216, x610x}, x840x);
	defparam lut_1179.LUT_SIZE = 6;
	defparam lut_1179.mask = 64'h37ff37ff00010000;

	lut_sub lut_1181 ({sk[425], n_n242, x360x, x839x, x7887x, x7888x}, x7894x);
	defparam lut_1181.LUT_SIZE = 6;
	defparam lut_1181.mask = 64'h37ff37ff0f3f5f7f;

	lut_sub lut_1185 ({sk[426], i_36_, x609x, x840x, x7894x}, n_n1567);
	defparam lut_1185.LUT_SIZE = 5;
	defparam lut_1185.mask = 32'h0f0f777f;

	lut_sub lut_1189 ({sk[427], n_n458, n_n242, x458x, x838x, x7902x}, x670x);
	defparam lut_1189.LUT_SIZE = 6;
	defparam lut_1189.mask = 64'h37ff37ff333f777f;

	lut_sub lut_1193 ({sk[428], i_10_, i_17_, x43x, x332x, x832x}, x7907x);
	defparam lut_1193.LUT_SIZE = 6;
	defparam lut_1193.mask = 64'h37ff37ff57555555;

	lut_sub lut_1196 ({sk[429], i_7_, x290x, x383x, x831x, x9208x}, x7908x);
	defparam lut_1196.LUT_SIZE = 6;
	defparam lut_1196.mask = 64'h37ff37ffbbbfbbbb;

	lut_sub lut_1200 ({sk[430], i_36_, x670x, x7907x, x7908x}, n_n1569);
	defparam lut_1200.LUT_SIZE = 5;
	defparam lut_1200.mask = 32'h0f0f777f;

	lut_sub lut_1204 ({sk[431], n_n880, x468x, x515x, x827x, x828x}, x823x);
	defparam lut_1204.LUT_SIZE = 6;
	defparam lut_1204.mask = 64'h37ff37ff0000777f;

	lut_sub lut_1208 ({sk[432], i_32_, i_36_, n_n358, x67x, x822x}, x7916x);
	defparam lut_1208.LUT_SIZE = 6;
	defparam lut_1208.mask = 64'h37ff37ff55575555;

	lut_sub lut_1211 ({sk[433], i_23_, x43x, x396x, x360x, x824x}, x7917x);
	defparam lut_1211.LUT_SIZE = 6;
	defparam lut_1211.mask = 64'h37ff37ff55575555;

	lut_sub lut_1214 ({sk[434], i_13_, n_n1408, n_n1089, x332x, x383x}, x7918x);
	defparam lut_1214.LUT_SIZE = 6;
	defparam lut_1214.mask = 64'h37ff37ff05050537;

	lut_sub lut_1217 ({sk[435], x823x, x7916x, x7917x, x7918x}, n_n1568);
	defparam lut_1217.LUT_SIZE = 5;
	defparam lut_1217.mask = 32'h0f0f7fff;

	lut_sub lut_1222 ({sk[436], i_14_, i_13_, i_12_}, n_n1384);
	defparam lut_1222.LUT_SIZE = 4;
	defparam lut_1222.mask = 16'h7708;

	lut_sub lut_1224 ({sk[437], i_23_, i_17_, i_21_}, n_n1282);
	defparam lut_1224.LUT_SIZE = 4;
	defparam lut_1224.mask = 16'h7780;

	lut_sub lut_1226 ({sk[438], i_9_, i_6_, i_13_}, n_n839);
	defparam lut_1226.LUT_SIZE = 4;
	defparam lut_1226.mask = 16'h7740;

	lut_sub lut_1228 ({sk[439], i_32_, i_34_, i_33_}, n_n1311);
	defparam lut_1228.LUT_SIZE = 4;
	defparam lut_1228.mask = 16'h7780;

	lut_sub lut_1230 ({sk[440], i_13_, i_12_, i_16_, n_n1307, n_n1303}, n_n263);
	defparam lut_1230.LUT_SIZE = 6;
	defparam lut_1230.mask = 64'h37ff37ff10000000;

	lut_sub lut_1232 ({sk[441], i_14_, i_12_, i_16_, n_n1307, n_n1303}, n_n363);
	defparam lut_1232.LUT_SIZE = 6;
	defparam lut_1232.mask = 64'h37ff37ff10000000;

	lut_sub lut_1234 ({sk[442], i_13_, i_12_, i_18_}, n_n584);
	defparam lut_1234.LUT_SIZE = 4;
	defparam lut_1234.mask = 16'h7710;

	lut_sub lut_1236 ({sk[443], i_9_, i_8_, i_11_}, n_n1033);
	defparam lut_1236.LUT_SIZE = 4;
	defparam lut_1236.mask = 16'h7704;

	lut_sub lut_1238 ({sk[444], i_9_, i_8_, i_5_, i_6_}, x7420x);
	defparam lut_1238.LUT_SIZE = 5;
	defparam lut_1238.mask = 32'h0f0f0080;

	lut_sub lut_1240 ({sk[445], i_13_, i_18_, i_19_, x229x}, n_n284);
	defparam lut_1240.LUT_SIZE = 5;
	defparam lut_1240.mask = 32'h0f0f0100;

	lut_sub lut_1242 ({sk[446], i_9_, i_8_, i_13_}, n_n1028);
	defparam lut_1242.LUT_SIZE = 4;
	defparam lut_1242.mask = 16'h7708;

	lut_sub lut_1244 ({sk[447], i_13_, i_11_, i_16_}, n_n178);
	defparam lut_1244.LUT_SIZE = 4;
	defparam lut_1244.mask = 16'h7780;

	lut_sub lut_1246 ({sk[448], i_30_, i_29_}, x57x);
	defparam lut_1246.LUT_SIZE = 3;
	defparam lut_1246.mask = 8'h58;

	lut_sub lut_1248 ({sk[449], i_30_, i_7_, i_8_}, x77x);
	defparam lut_1248.LUT_SIZE = 4;
	defparam lut_1248.mask = 16'h7780;

	lut_sub lut_1250 ({sk[450], i_28_, i_22_}, x83x);
	defparam lut_1250.LUT_SIZE = 3;
	defparam lut_1250.mask = 8'h54;

	lut_sub lut_1252 ({sk[451], i_28_, i_34_, i_35_, i_29_}, x372x);
	defparam lut_1252.LUT_SIZE = 5;
	defparam lut_1252.mask = 32'h0f0f1000;

	lut_sub lut_1254 ({sk[452], i_28_, i_26_, i_33_, i_38_, i_29_}, x380x);
	defparam lut_1254.LUT_SIZE = 6;
	defparam lut_1254.mask = 64'h37ff37ff20000000;

	lut_sub lut_1256 ({sk[453], i_28_, i_25_, i_26_, i_29_}, x71x);
	defparam lut_1256.LUT_SIZE = 5;
	defparam lut_1256.mask = 32'h0f0f8000;

	lut_sub lut_1258 ({sk[454], i_25_, i_26_, i_24_, i_38_, x42x}, x395x);
	defparam lut_1258.LUT_SIZE = 6;
	defparam lut_1258.mask = 64'h37ff37ff10000000;

	lut_sub lut_1260 ({sk[455], i_30_, i_7_, i_28_, i_32_, i_29_}, x474x);
	defparam lut_1260.LUT_SIZE = 6;
	defparam lut_1260.mask = 64'h37ff37ff80000000;

	lut_sub lut_1262 ({sk[456], i_26_, i_24_, i_33_, i_38_}, x503x);
	defparam lut_1262.LUT_SIZE = 5;
	defparam lut_1262.mask = 32'h0f0f4000;

	lut_sub lut_1264 ({sk[457], i_27_, i_23_, i_16_}, n_n1251);
	defparam lut_1264.LUT_SIZE = 4;
	defparam lut_1264.mask = 16'h7780;

	lut_sub lut_1266 ({sk[458], i_14_, i_31_, i_33_, n_n1397, n_n1251}, x545x);
	defparam lut_1266.LUT_SIZE = 6;
	defparam lut_1266.mask = 64'h37ff37ff00220323;

	lut_sub lut_1269 ({sk[459], i_30_, i_7_, i_32_, x9x, x71x}, x1132x);
	defparam lut_1269.LUT_SIZE = 6;
	defparam lut_1269.mask = 64'h37ff37ff10000000;

	lut_sub lut_1271 ({sk[460], i_20_, i_22_, x372x, x1131x}, x7606x);
	defparam lut_1271.LUT_SIZE = 5;
	defparam lut_1271.mask = 32'h0f0f5575;

	lut_sub lut_1274 ({sk[461], i_24_, x77x, x380x, x474x, x503x}, x7607x);
	defparam lut_1274.LUT_SIZE = 6;
	defparam lut_1274.mask = 64'h37ff37ff111f1111;

	lut_sub lut_1277 ({sk[462], x83x, x545x, x1132x, x7606x, x7607x}, n_n1891);
	defparam lut_1277.LUT_SIZE = 6;
	defparam lut_1277.mask = 64'h37ff37ff7f7f7fff;

	lut_sub lut_1282 ({sk[463], i_14_, i_13_, i_16_}, n_n1387);
	defparam lut_1282.LUT_SIZE = 4;
	defparam lut_1282.mask = 16'h7708;

	lut_sub lut_1284 ({sk[464], i_9_, i_10_, i_24_}, n_n1359);
	defparam lut_1284.LUT_SIZE = 4;
	defparam lut_1284.mask = 16'h7708;

	lut_sub lut_1286 ({sk[465], i_23_, i_21_, i_16_}, n_n1254);
	defparam lut_1286.LUT_SIZE = 4;
	defparam lut_1286.mask = 16'h7780;

	lut_sub lut_1288 ({sk[466], i_27_, i_34_, i_33_, x42x, x38x}, x145x);
	defparam lut_1288.LUT_SIZE = 6;
	defparam lut_1288.mask = 64'h37ff37ff00010000;

	lut_sub lut_1290 ({sk[467], i_26_, i_24_, i_34_}, x452x);
	defparam lut_1290.LUT_SIZE = 4;
	defparam lut_1290.mask = 16'h7780;

	lut_sub lut_1292 ({sk[468], i_7_, i_36_, n_n1438, x214x, x464x}, x812x);
	defparam lut_1292.LUT_SIZE = 6;
	defparam lut_1292.mask = 64'h37ff37ff00570000;

	lut_sub lut_1295 ({sk[469], n_n1489, x340x, x145x, x452x, x812x}, x7929x);
	defparam lut_1295.LUT_SIZE = 6;
	defparam lut_1295.mask = 64'h37ff37ff5f5f5f7f;

	lut_sub lut_1299 ({sk[470], i_25_, i_33_, x42x, n_n1438, n_n1397}, x126x);
	defparam lut_1299.LUT_SIZE = 6;
	defparam lut_1299.mask = 64'h37ff37ff00000001;

	lut_sub lut_1301 ({sk[471], i_14_, i_33_, x42x, n_n1438, n_n1397}, x128x);
	defparam lut_1301.LUT_SIZE = 6;
	defparam lut_1301.mask = 64'h37ff37ff00000001;

	lut_sub lut_1303 ({sk[472], i_30_, i_28_, i_29_, n_n1393, x806x}, x196x);
	defparam lut_1303.LUT_SIZE = 6;
	defparam lut_1303.mask = 64'h37ff37ff10000000;

	lut_sub lut_1305 ({sk[473], x7929x, x126x, x128x, x196x}, n_n1585);
	defparam lut_1305.LUT_SIZE = 5;
	defparam lut_1305.mask = 32'h0f0f7fff;

	lut_sub lut_1310 ({sk[474], i_32_, i_34_, i_35_}, n_n1422);
	defparam lut_1310.LUT_SIZE = 4;
	defparam lut_1310.mask = 16'h7720;

	lut_sub lut_1312 ({sk[475], i_14_, i_12_, i_17_, i_16_}, x8x);
	defparam lut_1312.LUT_SIZE = 5;
	defparam lut_1312.mask = 32'h0f0fa800;

	lut_sub lut_1315 ({sk[476], i_17_, i_16_, x54x, n_n1384, n_n1387}, x38x);
	defparam lut_1315.LUT_SIZE = 6;
	defparam lut_1315.mask = 64'h37ff37ff07050300;

	lut_sub lut_1318 ({sk[477], i_23_, i_24_, i_22_, i_34_, n_n1406}, x308x);
	defparam lut_1318.LUT_SIZE = 6;
	defparam lut_1318.mask = 64'h37ff37ff01000000;

	lut_sub lut_1320 ({sk[478], i_13_, i_12_, i_17_, i_16_, x308x}, x1661x);
	defparam lut_1320.LUT_SIZE = 6;
	defparam lut_1320.mask = 64'h37ff37ff44400000;

	lut_sub lut_1323 ({sk[479], i_24_, i_34_, i_29_, x302x, n_n1425}, x1663x);
	defparam lut_1323.LUT_SIZE = 6;
	defparam lut_1323.mask = 64'h37ff37ff01000000;

	lut_sub lut_1325 ({sk[480], n_n1433, x54x, x6984x, x44x, x805x}, x1664x);
	defparam lut_1325.LUT_SIZE = 6;
	defparam lut_1325.mask = 64'h37ff37ff0011001f;

	lut_sub lut_1328 ({sk[481], i_22_, x1661x, x1663x, x1664x}, x90x);
	defparam lut_1328.LUT_SIZE = 5;
	defparam lut_1328.mask = 32'h0f0f0f7f;

	lut_sub lut_1332 ({sk[482], i_23_, i_24_, i_34_, n_n1489, x340x}, x112x);
	defparam lut_1332.LUT_SIZE = 6;
	defparam lut_1332.mask = 64'h37ff37ff01000000;

	lut_sub lut_1334 ({sk[483], i_30_, i_22_, i_32_, i_31_, x372x}, x127x);
	defparam lut_1334.LUT_SIZE = 6;
	defparam lut_1334.mask = 64'h37ff37ff00400000;

	lut_sub lut_1336 ({sk[484], i_27_, i_28_, i_26_, i_33_}, x6958x);
	defparam lut_1336.LUT_SIZE = 5;
	defparam lut_1336.mask = 32'h0f0f4000;

	lut_sub lut_1338 ({sk[485], i_25_, i_23_, i_24_, i_33_, n_n1441}, x309x);
	defparam lut_1338.LUT_SIZE = 6;
	defparam lut_1338.mask = 64'h37ff37ff00001000;

	lut_sub lut_1340 ({sk[486], i_30_, i_31_, i_29_}, n_n1459);
	defparam lut_1340.LUT_SIZE = 4;
	defparam lut_1340.mask = 16'h7780;

	lut_sub lut_1342 ({sk[487], i_28_, i_23_, i_24_, i_31_, x57x}, x419x);
	defparam lut_1342.LUT_SIZE = 6;
	defparam lut_1342.mask = 64'h37ff37ff40000000;

	lut_sub lut_1344 ({sk[488], i_30_, i_31_, i_29_, n_n1497}, x513x);
	defparam lut_1344.LUT_SIZE = 5;
	defparam lut_1344.mask = 32'h0f0f4000;

	lut_sub lut_1346 ({sk[489], x112x, x127x, x507x, x7934x, x9207x}, x7938x);
	defparam lut_1346.LUT_SIZE = 6;
	defparam lut_1346.mask = 64'h37ff37ffbfffffff;

	lut_sub lut_1352 ({sk[490], n_n1585, x90x, x7938x}, n_n1556);
	defparam lut_1352.LUT_SIZE = 4;
	defparam lut_1352.mask = 16'h777f;

	lut_sub lut_1356 ({sk[491], i_7_, i_14_, i_16_}, n_n1377);
	defparam lut_1356.LUT_SIZE = 4;
	defparam lut_1356.mask = 16'h7708;

	lut_sub lut_1358 ({sk[492], i_30_, i_34_, i_36_, i_35_}, n_n820);
	defparam lut_1358.LUT_SIZE = 5;
	defparam lut_1358.mask = 32'h0f0f1000;

	lut_sub lut_1360 ({sk[493], i_9_, i_11_, i_19_, n_n1307, n_n1303}, n_n706);
	defparam lut_1360.LUT_SIZE = 6;
	defparam lut_1360.mask = 64'h37ff37ff10000000;

	lut_sub lut_1362 ({sk[494], i_14_, i_23_, i_24_, i_16_, x11x}, n_n608);
	defparam lut_1362.LUT_SIZE = 6;
	defparam lut_1362.mask = 64'h37ff37ff40000000;

	lut_sub lut_1364 ({sk[495], i_14_, i_13_, i_16_}, n_n916);
	defparam lut_1364.LUT_SIZE = 4;
	defparam lut_1364.mask = 16'h7720;

	lut_sub lut_1366 ({sk[496], i_20_, i_17_, i_16_}, n_n629);
	defparam lut_1366.LUT_SIZE = 4;
	defparam lut_1366.mask = 16'h7780;

	lut_sub lut_1368 ({sk[497], i_24_, i_35_, i_38_}, x12x);
	defparam lut_1368.LUT_SIZE = 4;
	defparam lut_1368.mask = 16'h7740;

	lut_sub lut_1370 ({sk[498], i_28_, i_24_, i_35_, i_38_, n_n1241}, x520x);
	defparam lut_1370.LUT_SIZE = 6;
	defparam lut_1370.mask = 64'h37ff37ff10000000;

	lut_sub lut_1372 ({sk[499], i_28_, i_24_, i_19_, n_n1361, n_n1241}, n_n338);
	defparam lut_1372.LUT_SIZE = 6;
	defparam lut_1372.mask = 64'h37ff37ff01000000;

	lut_sub lut_1374 ({sk[500], i_27_, i_28_, i_26_, i_24_, i_29_}, x45x);
	defparam lut_1374.LUT_SIZE = 6;
	defparam lut_1374.mask = 64'h37ff37ff40000000;

	lut_sub lut_1376 ({sk[501], i_27_, i_34_, i_35_, x42x, n_n1322}, x373x);
	defparam lut_1376.LUT_SIZE = 6;
	defparam lut_1376.mask = 64'h37ff37ff01000000;

	lut_sub lut_1378 ({sk[502], x14x, n_n916, x256x, x87x, x326x}, x7758x);
	defparam lut_1378.LUT_SIZE = 6;
	defparam lut_1378.mask = 64'h37ff37ff00330537;

	lut_sub lut_1381 ({sk[503], i_20_, i_34_, i_35_, x296x, n_n1406}, x255x);
	defparam lut_1381.LUT_SIZE = 6;
	defparam lut_1381.mask = 64'h37ff37ff00000100;

	lut_sub lut_1383 ({sk[504], x43x, n_n1315, x263x, n_n1323, x299x}, x450x);
	defparam lut_1383.LUT_SIZE = 6;
	defparam lut_1383.mask = 64'h37ff37ff01010155;

	lut_sub lut_1386 ({sk[505], n_n1375, n_n1429, n_n846, x342x, x478x}, x9205x);
	defparam lut_1386.LUT_SIZE = 6;
	defparam lut_1386.mask = 64'h37ff37ffffaafca8;

	lut_sub lut_1393 ({sk[506], i_17_, x43x, x255x, x450x, x9205x}, x7955x);
	defparam lut_1393.LUT_SIZE = 6;
	defparam lut_1393.mask = 64'h37ff37ffbbbfbbbb;

	lut_sub lut_1397 ({sk[507], i_7_, i_8_, n_n1375, n_n1322, n_n820}, x517x);
	defparam lut_1397.LUT_SIZE = 6;
	defparam lut_1397.mask = 64'h37ff37ff01000000;

	lut_sub lut_1399 ({sk[508], i_2_, i_21_, i_36_, x263x, x65x}, x481x);
	defparam lut_1399.LUT_SIZE = 6;
	defparam lut_1399.mask = 64'h37ff37ff01000000;

	lut_sub lut_1401 ({sk[509], i_14_, i_13_, i_16_, x337x, x511x}, x9204x);
	defparam lut_1401.LUT_SIZE = 6;
	defparam lut_1401.mask = 64'h37ff37ff8acfaaff;

	lut_sub lut_1408 ({sk[510], i_14_, x517x, x481x, x9204x}, x7956x);
	defparam lut_1408.LUT_SIZE = 5;
	defparam lut_1408.mask = 32'h0f0fbfaa;

	lut_sub lut_1412 ({sk[511], i_32_, i_36_, n_n1489, n_n1397, n_n1251}, x472x);
	defparam lut_1412.LUT_SIZE = 6;
	defparam lut_1412.mask = 64'h37ff37ff00010000;

	lut_sub lut_1414 ({sk[512], i_2_, i_36_, n_n1443, x228x, x77x}, x364x);
	defparam lut_1414.LUT_SIZE = 6;
	defparam lut_1414.mask = 64'h37ff37ff00010000;

	lut_sub lut_1416 ({sk[513], i_36_, i_35_, n_n1441, n_n1459, x342x}, x392x);
	defparam lut_1416.LUT_SIZE = 6;
	defparam lut_1416.mask = 64'h37ff37ff00000100;

	lut_sub lut_1418 ({sk[514], i_8_, i_14_, i_16_, x48x, n_n846}, x397x);
	defparam lut_1418.LUT_SIZE = 6;
	defparam lut_1418.mask = 64'h37ff37ff10000000;

	lut_sub lut_1420 ({sk[515], n_n1147, x472x, x364x, x392x, x397x}, x7966x);
	defparam lut_1420.LUT_SIZE = 6;
	defparam lut_1420.mask = 64'h37ff37ff7f7f7fff;

	lut_sub lut_1425 ({sk[516], i_20_, i_21_, x234x, x9229x}, x7978x);
	defparam lut_1425.LUT_SIZE = 5;
	defparam lut_1425.mask = 32'h0f0f33b3;

	lut_sub lut_1428 ({sk[517], i_26_, x54x, n_n984, x325x, x328x}, x9195x);
	defparam lut_1428.LUT_SIZE = 6;
	defparam lut_1428.mask = 64'h37ff37fffff8ffff;

	lut_sub lut_1439 ({sk[518], n_n1141, n_n1263, x374x, x7978x, x9195x}, x7982x);
	defparam lut_1439.LUT_SIZE = 6;
	defparam lut_1439.mask = 64'h37ff37ffbbbbbbbf;

	lut_sub lut_1443 ({sk[519], i_24_, i_21_, i_34_, n_n1425}, x441x);
	defparam lut_1443.LUT_SIZE = 5;
	defparam lut_1443.mask = 32'h0f0f0400;

	lut_sub lut_1445 ({sk[520], i_21_, i_36_, n_n1141, n_n1213, x7053x}, x301x);
	defparam lut_1445.LUT_SIZE = 6;
	defparam lut_1445.mask = 64'h37ff37ff00010000;

	lut_sub lut_1447 ({sk[521], i_7_, x290x, n_n1089, x467x, x514x}, x9194x);
	defparam lut_1447.LUT_SIZE = 6;
	defparam lut_1447.mask = 64'h37ff37fffca8fcfc;

	lut_sub lut_1454 ({sk[522], x43x, x340x, x441x, x301x, x9194x}, x7983x);
	defparam lut_1454.LUT_SIZE = 6;
	defparam lut_1454.mask = 64'h37ff37ffaaafbbbf;

	lut_sub lut_1458 ({sk[523], i_8_, n_n1441, x10x, x74x, x348x}, x667x);
	defparam lut_1458.LUT_SIZE = 6;
	defparam lut_1458.mask = 64'h37ff37ff03570055;

	lut_sub lut_1461 ({sk[524], i_25_, i_21_, n_n1404, n_n1408, x505x}, x192x);
	defparam lut_1461.LUT_SIZE = 6;
	defparam lut_1461.mask = 64'h37ff37ff00000015;

	lut_sub lut_1464 ({sk[525], i_27_, x42x, n_n1504, n_n1322, n_n1285}, x194x);
	defparam lut_1464.LUT_SIZE = 6;
	defparam lut_1464.mask = 64'h37ff37ff00010000;

	lut_sub lut_1466 ({sk[526], n_n880, n_n1459, x667x, x192x, x194x}, x7992x);
	defparam lut_1466.LUT_SIZE = 6;
	defparam lut_1466.mask = 64'h37ff37ff7777777f;

	lut_sub lut_1470 ({sk[527], i_27_, i_28_, i_29_, n_n1504, n_n1315}, x486x);
	defparam lut_1470.LUT_SIZE = 6;
	defparam lut_1470.mask = 64'h37ff37ff10000000;

	lut_sub lut_1472 ({sk[528], n_n1089, x48x, x259x, n_n846, x514x}, x9193x);
	defparam lut_1472.LUT_SIZE = 6;
	defparam lut_1472.mask = 64'h37ff37fffffcaaa8;

	lut_sub lut_1479 ({sk[529], i_23_, x10x, x301x, x486x, x9193x}, x7993x);
	defparam lut_1479.LUT_SIZE = 6;
	defparam lut_1479.mask = 64'h37ff37ffaabfaaaf;

	lut_sub lut_1483 ({sk[530], i_14_, i_28_, i_33_, n_n1438, n_n1397}, x189x);
	defparam lut_1483.LUT_SIZE = 6;
	defparam lut_1483.mask = 64'h37ff37ff00000100;

	lut_sub lut_1485 ({sk[531], i_27_, i_17_, x54x, n_n1511, n_n1285}, x190x);
	defparam lut_1485.LUT_SIZE = 6;
	defparam lut_1485.mask = 64'h37ff37ff01000000;

	lut_sub lut_1487 ({sk[532], i_23_, i_34_, i_33_, n_n1216, n_n1384}, x191x);
	defparam lut_1487.LUT_SIZE = 6;
	defparam lut_1487.mask = 64'h37ff37ff00010000;

	lut_sub lut_1489 ({sk[533], i_21_, i_16_, x189x, x190x, x191x}, x186x);
	defparam lut_1489.LUT_SIZE = 6;
	defparam lut_1489.mask = 64'h37ff37ff00007f0f;

	lut_sub lut_1493 ({sk[534], i_14_, i_16_, n_n1315, x300x}, x183x);
	defparam lut_1493.LUT_SIZE = 5;
	defparam lut_1493.mask = 32'h0f0f1000;

	lut_sub lut_1495 ({sk[535], i_23_, x43x, x486x, x182x, x184x}, x8003x);
	defparam lut_1495.LUT_SIZE = 6;
	defparam lut_1495.mask = 64'h37ff37ff777f7777;

	lut_sub lut_1499 ({sk[536], n_n1404, n_n1408, x209x, x183x, x8003x}, x8004x);
	defparam lut_1499.LUT_SIZE = 6;
	defparam lut_1499.mask = 64'h37ff37ff777f7f7f;

	lut_sub lut_1504 ({sk[537], i_27_, i_36_, x73x, n_n620, n_n1288}, x173x);
	defparam lut_1504.LUT_SIZE = 6;
	defparam lut_1504.mask = 64'h37ff37ff00010000;

	lut_sub lut_1506 ({sk[538], i_14_, x245x, n_n984, x511x, x325x}, x9199x);
	defparam lut_1506.LUT_SIZE = 6;
	defparam lut_1506.mask = 64'h37ff37ffccc8fffa;

	lut_sub lut_1513 ({sk[539], i_12_, x10x, x255x, x173x, x9199x}, x8016x);
	defparam lut_1513.LUT_SIZE = 6;
	defparam lut_1513.mask = 64'h37ff37ffbbbfbbbb;

	lut_sub lut_1517 ({sk[540], i_36_, n_n269, x256x, x9198x}, x174x);
	defparam lut_1517.LUT_SIZE = 5;
	defparam lut_1517.mask = 32'h0f0f00ab;

	lut_sub lut_1520 ({sk[541], i_13_, i_16_, x295x, x352x}, x8015x);
	defparam lut_1520.LUT_SIZE = 5;
	defparam lut_1520.mask = 32'h0f0f7500;

	lut_sub lut_1523 ({sk[542], x8016x, x174x, x8015x}, n_n1571);
	defparam lut_1523.LUT_SIZE = 4;
	defparam lut_1523.mask = 16'h777f;

	lut_sub lut_1527 ({sk[543], i_36_, i_35_, n_n1441, n_n544, n_n1133}, x162x);
	defparam lut_1527.LUT_SIZE = 6;
	defparam lut_1527.mask = 64'h37ff37ff00000100;

	lut_sub lut_1529 ({sk[544], i_21_, i_34_, x54x, n_n984, x328x}, x163x);
	defparam lut_1529.LUT_SIZE = 6;
	defparam lut_1529.mask = 64'h37ff37ff00000001;

	lut_sub lut_1531 ({sk[545], i_12_, i_17_, x43x, x393x, x382x}, x9197x);
	defparam lut_1531.LUT_SIZE = 6;
	defparam lut_1531.mask = 64'h37ff37fff8faf8ff;

	lut_sub lut_1536 ({sk[546], n_n1375, n_n1334, x162x, x163x, x9197x}, x8025x);
	defparam lut_1536.LUT_SIZE = 6;
	defparam lut_1536.mask = 64'h37ff37ff3f3f3fbf;

	lut_sub lut_1540 ({sk[547], i_36_, n_n620, n_n363, x273x, x256x}, x165x);
	defparam lut_1540.LUT_SIZE = 6;
	defparam lut_1540.mask = 64'h37ff37ff00000357;

	lut_sub lut_1543 ({sk[548], i_14_, i_16_, x295x, x352x}, x8024x);
	defparam lut_1543.LUT_SIZE = 5;
	defparam lut_1543.mask = 32'h0f0f7500;

	lut_sub lut_1546 ({sk[549], x8025x, x165x, x8024x}, n_n1570);
	defparam lut_1546.LUT_SIZE = 4;
	defparam lut_1546.mask = 16'h777f;

	lut_sub lut_1550 ({sk[550], i_27_, x42x, n_n1141, n_n1263, n_n820}, x158x);
	defparam lut_1550.LUT_SIZE = 6;
	defparam lut_1550.mask = 64'h37ff37ff00010000;

	lut_sub lut_1552 ({sk[551], i_34_, n_n1018, n_n1499, x325x, x328x}, x9203x);
	defparam lut_1552.LUT_SIZE = 6;
	defparam lut_1552.mask = 64'h37ff37fffffffff8;

	lut_sub lut_1563 ({sk[552], i_12_, x43x, x255x, x158x, x9203x}, x8037x);
	defparam lut_1563.LUT_SIZE = 6;
	defparam lut_1563.mask = 64'h37ff37ffbbbfbbbb;

	lut_sub lut_1567 ({sk[553], i_2_, i_36_, n_n1408, x228x, x77x}, x156x);
	defparam lut_1567.LUT_SIZE = 6;
	defparam lut_1567.mask = 64'h37ff37ff00010000;

	lut_sub lut_1569 ({sk[554], i_31_, n_n1441, n_n1443, x393x, x382x}, x9201x);
	defparam lut_1569.LUT_SIZE = 6;
	defparam lut_1569.mask = 64'h37ff37fffffffff8;

	lut_sub lut_1580 ({sk[555], x79x, n_n1288, n_n1089, n_n269, x472x}, x9202x);
	defparam lut_1580.LUT_SIZE = 6;
	defparam lut_1580.mask = 64'h37ff37fffafafac8;

	lut_sub lut_1587 ({sk[556], x156x, x9201x, x9202x}, x8038x);
	defparam lut_1587.LUT_SIZE = 4;
	defparam lut_1587.mask = 16'h77ef;

	lut_sub lut_1591 ({sk[557], i_17_, n_n1387, x505x, x151x, x153x}, x730x);
	defparam lut_1591.LUT_SIZE = 6;
	defparam lut_1591.mask = 64'h37ff37ff777f3333;

	lut_sub lut_1595 ({sk[558], i_36_, n_n1404, n_n263, x478x, x67x}, x8046x);
	defparam lut_1595.LUT_SIZE = 6;
	defparam lut_1595.mask = 64'h37ff37ff00330537;

	lut_sub lut_1598 ({sk[559], i_17_, x10x, x255x, x142x, x9196x}, x8047x);
	defparam lut_1598.LUT_SIZE = 6;
	defparam lut_1598.mask = 64'h37ff37ffbbbfbbbb;

	lut_sub lut_1602 ({sk[560], i_21_, x730x, x8046x, x8047x}, n_n1572);
	defparam lut_1602.LUT_SIZE = 5;
	defparam lut_1602.mask = 32'h0f0f777f;

	lut_sub lut_1606 ({sk[561], x7966x, x186x, x8004x, x412x, x7965x}, x8051x);
	defparam lut_1606.LUT_SIZE = 6;
	defparam lut_1606.mask = 64'h37ff37ff7fffffff;

	lut_sub lut_1612 ({sk[562], x7982x, x7983x, x7992x, x7993x}, x8049x);
	defparam lut_1612.LUT_SIZE = 5;
	defparam lut_1612.mask = 32'h0f0f7fff;

	lut_sub lut_1617 ({sk[563], i_27_, i_16_}, x103x);
	defparam lut_1617.LUT_SIZE = 3;
	defparam lut_1617.mask = 8'h57;

	lut_sub lut_1620 ({sk[564], i_25_, i_24_, i_19_}, n_n998);
	defparam lut_1620.LUT_SIZE = 4;
	defparam lut_1620.mask = 16'h7740;

	lut_sub lut_1622 ({sk[565], i_27_, i_23_, i_22_, i_35_, n_n1326}, x40x);
	defparam lut_1622.LUT_SIZE = 6;
	defparam lut_1622.mask = 64'h37ff37ff01000000;

	lut_sub lut_1624 ({sk[566], i_27_, i_23_, i_17_, i_34_, i_35_}, x318x);
	defparam lut_1624.LUT_SIZE = 6;
	defparam lut_1624.mask = 64'h37ff37ff40000000;

	lut_sub lut_1626 ({sk[567], i_28_, i_33_, i_29_, n_n1387, x318x}, x124x);
	defparam lut_1626.LUT_SIZE = 6;
	defparam lut_1626.mask = 64'h37ff37ff00100000;

	lut_sub lut_1628 ({sk[568], i_34_, i_35_, n_n1257, n_n1384, n_n1251}, x132x);
	defparam lut_1628.LUT_SIZE = 6;
	defparam lut_1628.mask = 64'h37ff37ff00010000;

	lut_sub lut_1630 ({sk[569], i_27_, i_28_, i_26_, i_24_, i_31_}, x236x);
	defparam lut_1630.LUT_SIZE = 6;
	defparam lut_1630.mask = 64'h37ff37ff40000000;

	lut_sub lut_1632 ({sk[570], i_27_, i_28_, i_0_, i_29_, x73x}, x355x);
	defparam lut_1632.LUT_SIZE = 6;
	defparam lut_1632.mask = 64'h37ff37ff01000000;

	lut_sub lut_1634 ({sk[571], n_n1404, n_n1315, n_n1263, x40x, x236x}, x8060x);
	defparam lut_1634.LUT_SIZE = 6;
	defparam lut_1634.mask = 64'h37ff37ff00053337;

	lut_sub lut_1637 ({sk[572], n_n1257, n_n1387, x318x, x132x, x8060x}, x8062x);
	defparam lut_1637.LUT_SIZE = 6;
	defparam lut_1637.mask = 64'h37ff37ff7777777f;

	lut_sub lut_1641 ({sk[573], i_25_, x245x, x277x, n_n1393, x441x}, x129x);
	defparam lut_1641.LUT_SIZE = 6;
	defparam lut_1641.mask = 64'h37ff37ff00001113;

	lut_sub lut_1644 ({sk[574], x10x, x290x, n_n1282, n_n1254, x355x}, x131x);
	defparam lut_1644.LUT_SIZE = 6;
	defparam lut_1644.mask = 64'h37ff37ff00110515;

	lut_sub lut_1647 ({sk[575], i_17_, x43x, x62x, x129x, x131x}, x8063x);
	defparam lut_1647.LUT_SIZE = 6;
	defparam lut_1647.mask = 64'h37ff37ff777f7777;

	lut_sub lut_1651 ({sk[576], i_28_, i_34_, i_33_, i_35_, n_n1438}, x287x);
	defparam lut_1651.LUT_SIZE = 6;
	defparam lut_1651.mask = 64'h37ff37ff01000000;

	lut_sub lut_1653 ({sk[577], n_n1315, n_n1314, n_n1322, x80x, n_n1323}, x554x);
	defparam lut_1653.LUT_SIZE = 6;
	defparam lut_1653.mask = 64'h37ff37ff01010133;

	lut_sub lut_1656 ({sk[578], i_27_, i_28_, i_25_, i_34_, i_33_}, x485x);
	defparam lut_1656.LUT_SIZE = 6;
	defparam lut_1656.mask = 64'h37ff37ff01000000;

	lut_sub lut_1658 ({sk[579], n_n1429, n_n1406, n_n1213, x7491x, x8x}, x118x);
	defparam lut_1658.LUT_SIZE = 6;
	defparam lut_1658.mask = 64'h37ff37ff00010003;

	lut_sub lut_1661 ({sk[580], n_n1408, n_n1312, x82x, x485x, x118x}, x8068x);
	defparam lut_1661.LUT_SIZE = 6;
	defparam lut_1661.mask = 64'h37ff37ff55555f7f;

	lut_sub lut_1665 ({sk[581], i_14_, i_12_, i_16_, x296x, x355x}, x116x);
	defparam lut_1665.LUT_SIZE = 6;
	defparam lut_1665.mask = 64'h37ff37ff10000000;

	lut_sub lut_1667 ({sk[582], i_25_, i_21_, x287x}, x117x);
	defparam lut_1667.LUT_SIZE = 4;
	defparam lut_1667.mask = 16'h7701;

	lut_sub lut_1669 ({sk[583], i_31_, i_34_, x554x, x116x, x117x}, x8069x);
	defparam lut_1669.LUT_SIZE = 6;
	defparam lut_1669.mask = 64'h37ff37ff7777777f;

	lut_sub lut_1673 ({sk[584], i_25_, i_23_, i_24_, i_34_, i_33_}, x6944x);
	defparam lut_1673.LUT_SIZE = 6;
	defparam lut_1673.mask = 64'h37ff37ff00001000;

	lut_sub lut_1675 ({sk[585], n_n1375, n_n1443, n_n1408, x40x, x6944x}, x104x);
	defparam lut_1675.LUT_SIZE = 6;
	defparam lut_1675.mask = 64'h37ff37ff00330537;

	lut_sub lut_1678 ({sk[586], i_27_, i_28_, i_29_, n_n1396, n_n1374}, x252x);
	defparam lut_1678.LUT_SIZE = 6;
	defparam lut_1678.mask = 64'h37ff37ff10000000;

	lut_sub lut_1680 ({sk[587], n_n1315, n_n1314, n_n1322, n_n1323, n_n1285}, x555x);
	defparam lut_1680.LUT_SIZE = 6;
	defparam lut_1680.mask = 64'h37ff37ff070707ff;

	lut_sub lut_1684 ({sk[588], i_14_, i_12_, i_16_, x104x, x252x}, x8072x);
	defparam lut_1684.LUT_SIZE = 6;
	defparam lut_1684.mask = 64'h37ff37ff73333333;

	lut_sub lut_1687 ({sk[589], i_13_, i_21_, i_16_, x242x, x355x}, x108x);
	defparam lut_1687.LUT_SIZE = 6;
	defparam lut_1687.mask = 64'h37ff37ff10000000;

	lut_sub lut_1689 ({sk[590], i_13_, i_12_, i_16_, n_n1408, x40x}, x110x);
	defparam lut_1689.LUT_SIZE = 6;
	defparam lut_1689.mask = 64'h37ff37ff51111111;

	lut_sub lut_1692 ({sk[591], x236x, x555x, x108x, x110x}, x8073x);
	defparam lut_1692.LUT_SIZE = 5;
	defparam lut_1692.mask = 32'h0f0f777f;

	lut_sub lut_1696 ({sk[592], i_28_, i_34_, i_35_, i_29_}, x214x);
	defparam lut_1696.LUT_SIZE = 5;
	defparam lut_1696.mask = 32'h0f0f2000;

	lut_sub lut_1698 ({sk[593], i_31_, i_36_, i_35_}, x265x);
	defparam lut_1698.LUT_SIZE = 4;
	defparam lut_1698.mask = 16'h7720;

	lut_sub lut_1700 ({sk[594], i_27_, i_28_, i_23_, i_29_}, x267x);
	defparam lut_1700.LUT_SIZE = 5;
	defparam lut_1700.mask = 32'h0f0f8000;

	lut_sub lut_1702 ({sk[595], i_9_, i_10_, i_13_, n_n461, x46x}, x881x);
	defparam lut_1702.LUT_SIZE = 6;
	defparam lut_1702.mask = 64'h37ff37ff10000000;

	lut_sub lut_1704 ({sk[596], i_14_, i_13_, i_17_, i_16_, x50x}, x559x);
	defparam lut_1704.LUT_SIZE = 6;
	defparam lut_1704.mask = 64'h37ff37ff40404000;

	lut_sub lut_1707 ({sk[597], i_13_, i_23_, i_17_, i_16_, x51x}, n_n329);
	defparam lut_1707.LUT_SIZE = 6;
	defparam lut_1707.mask = 64'h37ff37ff40000000;

	lut_sub lut_1709 ({sk[598], i_27_, i_26_, i_24_, i_31_, x42x}, x468x);
	defparam lut_1709.LUT_SIZE = 6;
	defparam lut_1709.mask = 64'h37ff37ff40000000;

	lut_sub lut_1711 ({sk[599], i_25_, i_26_, i_23_, i_24_, i_34_}, x806x);
	defparam lut_1711.LUT_SIZE = 6;
	defparam lut_1711.mask = 64'h37ff37ff0000c840;

	lut_sub lut_1714 ({sk[600], i_30_, i_23_, i_24_, n_n1433, x42x}, x464x);
	defparam lut_1714.LUT_SIZE = 6;
	defparam lut_1714.mask = 64'h37ff37ff10000000;

	lut_sub lut_1716 ({sk[601], i_7_, i_8_, i_36_, n_n1282, x45x}, x363x);
	defparam lut_1716.LUT_SIZE = 6;
	defparam lut_1716.mask = 64'h37ff37ff01000000;

	lut_sub lut_1718 ({sk[602], i_7_, i_32_, i_36_}, x7769x);
	defparam lut_1718.LUT_SIZE = 4;
	defparam lut_1718.mask = 16'h7740;

	lut_sub lut_1720 ({sk[603], i_32_, i_34_, i_29_, n_n1216}, x256x);
	defparam lut_1720.LUT_SIZE = 5;
	defparam lut_1720.mask = 32'h0f0f0400;

	lut_sub lut_1722 ({sk[604], n_n1375, n_n1443, n_n1422, x484x, x489x}, x956x);
	defparam lut_1722.LUT_SIZE = 6;
	defparam lut_1722.mask = 64'h37ff37ff00000007;

	lut_sub lut_1725 ({sk[605], i_27_, i_34_, i_35_, x242x, x272x}, x87x);
	defparam lut_1725.LUT_SIZE = 6;
	defparam lut_1725.mask = 64'h37ff37ff01000000;

	lut_sub lut_1727 ({sk[606], i_27_, i_26_, i_24_, i_36_, i_35_}, x368x);
	defparam lut_1727.LUT_SIZE = 6;
	defparam lut_1727.mask = 64'h37ff37ff20000000;

	lut_sub lut_1729 ({sk[607], i_10_, i_14_, i_13_, i_17_, i_16_}, x571x);
	defparam lut_1729.LUT_SIZE = 6;
	defparam lut_1729.mask = 64'h37ff37ff88800800;

	lut_sub lut_1732 ({sk[608], i_14_, i_13_, n_n825, x46x, n_n576}, x946x);
	defparam lut_1732.LUT_SIZE = 6;
	defparam lut_1732.mask = 64'h37ff37ff00010000;

	lut_sub lut_1734 ({sk[609], i_17_, i_16_, i_19_}, n_n130);
	defparam lut_1734.LUT_SIZE = 4;
	defparam lut_1734.mask = 16'h7780;

	lut_sub lut_1736 ({sk[610], i_34_, i_33_, i_35_, i_38_}, n_n1059);
	defparam lut_1736.LUT_SIZE = 5;
	defparam lut_1736.mask = 32'h0f0f1000;

	lut_sub lut_1738 ({sk[611], i_20_, i_17_, i_19_, n_n1406, n_n1213}, n_n18);
	defparam lut_1738.LUT_SIZE = 6;
	defparam lut_1738.mask = 64'h37ff37ff10000000;

	lut_sub lut_1740 ({sk[612], i_30_, i_31_, i_34_, i_36_, i_35_}, n_n846);
	defparam lut_1740.LUT_SIZE = 6;
	defparam lut_1740.mask = 64'h37ff37ff02000000;

	lut_sub lut_1742 ({sk[613], i_20_, i_18_, i_17_, n_n1406, n_n1213}, n_n21);
	defparam lut_1742.LUT_SIZE = 6;
	defparam lut_1742.mask = 64'h37ff37ff10000000;

	lut_sub lut_1744 ({sk[614], i_21_, i_31_, i_34_, i_35_, n_n793}, x299x);
	defparam lut_1744.LUT_SIZE = 6;
	defparam lut_1744.mask = 64'h37ff37ff00000010;

	lut_sub lut_1746 ({sk[615], i_7_, i_27_, x227x, n_n1489, x242x}, x337x);
	defparam lut_1746.LUT_SIZE = 6;
	defparam lut_1746.mask = 64'h37ff37ff01000000;

	lut_sub lut_1748 ({sk[616], i_8_, i_14_, i_12_, i_16_, x54x}, x342x);
	defparam lut_1748.LUT_SIZE = 6;
	defparam lut_1748.mask = 64'h37ff37ff40000000;

	lut_sub lut_1750 ({sk[617], i_21_, n_n1441, x54x, n_n1438, n_n880}, x478x);
	defparam lut_1750.LUT_SIZE = 6;
	defparam lut_1750.mask = 64'h37ff37ff00010000;

	lut_sub lut_1752 ({sk[618], i_8_, i_12_, n_n1345, n_n1254, x368x}, x511x);
	defparam lut_1752.LUT_SIZE = 6;
	defparam lut_1752.mask = 64'h37ff37ff01000000;

	lut_sub lut_1754 ({sk[619], i_7_, i_26_, i_32_, x54x, x7053x}, x65x);
	defparam lut_1754.LUT_SIZE = 6;
	defparam lut_1754.mask = 64'h37ff37ff10000000;

	lut_sub lut_1756 ({sk[620], i_2_, i_36_}, x433x);
	defparam lut_1756.LUT_SIZE = 3;
	defparam lut_1756.mask = 8'h54;

	lut_sub lut_1758 ({sk[621], i_27_, i_28_, i_26_, i_29_, x54x}, x67x);
	defparam lut_1758.LUT_SIZE = 6;
	defparam lut_1758.mask = 64'h37ff37ff40000000;

	lut_sub lut_1760 ({sk[622], i_8_, i_12_, n_n461, n_n1254, x45x}, x501x);
	defparam lut_1760.LUT_SIZE = 6;
	defparam lut_1760.mask = 64'h37ff37ff01000000;

	lut_sub lut_1762 ({sk[623], i_3_, i_11_, i_18_, i_19_}, x578x);
	defparam lut_1762.LUT_SIZE = 5;
	defparam lut_1762.mask = 32'h0f0fa0ec;

	lut_sub lut_1765 ({sk[624], i_8_, i_18_, x60x, x257x}, x1462x);
	defparam lut_1765.LUT_SIZE = 5;
	defparam lut_1765.mask = 32'h0f0f1000;

	lut_sub lut_1767 ({sk[625], i_3_, i_13_, i_18_, i_22_, i_19_}, x5x);
	defparam lut_1767.LUT_SIZE = 6;
	defparam lut_1767.mask = 64'h37ff37ff44000400;

	lut_sub lut_1770 ({sk[626], i_13_, i_11_, i_18_, i_22_}, x349x);
	defparam lut_1770.LUT_SIZE = 5;
	defparam lut_1770.mask = 32'h0f0f0200;

	lut_sub lut_1772 ({sk[627], i_9_, i_28_, i_12_, i_26_, i_24_}, x7261x);
	defparam lut_1772.LUT_SIZE = 6;
	defparam lut_1772.mask = 64'h37ff37ff00000800;

	lut_sub lut_1774 ({sk[628], i_28_, i_12_, i_26_, i_24_, i_22_}, x7263x);
	defparam lut_1774.LUT_SIZE = 6;
	defparam lut_1774.mask = 64'h37ff37ff00800000;

	lut_sub lut_1776 ({sk[629], x262x, x5x, x349x, x7261x, x7263x}, x579x);
	defparam lut_1776.LUT_SIZE = 6;
	defparam lut_1776.mask = 64'h37ff37ff03335777;

	lut_sub lut_1780 ({sk[630], i_11_, i_32_, i_19_, x297x, x14x}, x9219x);
	defparam lut_1780.LUT_SIZE = 6;
	defparam lut_1780.mask = 64'h37ff37ff8cffccff;

	lut_sub lut_1785 ({sk[631], i_9_, i_8_, i_13_, i_11_, x208x}, x423x);
	defparam lut_1785.LUT_SIZE = 6;
	defparam lut_1785.mask = 64'h37ff37ff00001000;

	lut_sub lut_1787 ({sk[632], i_9_, i_13_, i_11_, i_18_, x50x}, x435x);
	defparam lut_1787.LUT_SIZE = 6;
	defparam lut_1787.mask = 64'h37ff37ff00000100;

	lut_sub lut_1789 ({sk[633], i_13_, x208x, n_n1033, x435x}, x20x);
	defparam lut_1789.LUT_SIZE = 5;
	defparam lut_1789.mask = 32'h0f0f5755;

	lut_sub lut_1792 ({sk[634], i_13_, i_11_, i_18_, i_22_, x5x}, x23x);
	defparam lut_1792.LUT_SIZE = 6;
	defparam lut_1792.mask = 64'h37ff37ff555d5555;

	lut_sub lut_1795 ({sk[635], i_24_, i_35_, i_38_, x42x, n_n1340}, x253x);
	defparam lut_1795.LUT_SIZE = 6;
	defparam lut_1795.mask = 64'h37ff37ff01000000;

	lut_sub lut_1797 ({sk[636], i_10_, i_12_}, x405x);
	defparam lut_1797.LUT_SIZE = 3;
	defparam lut_1797.mask = 8'h51;

	lut_sub lut_1799 ({sk[637], i_33_, i_35_, i_38_, n_n1497}, x509x);
	defparam lut_1799.LUT_SIZE = 5;
	defparam lut_1799.mask = 32'h0f0f1000;

	lut_sub lut_1801 ({sk[638], i_11_, x11x, n_n1048, x213x, x7425x}, x100x);
	defparam lut_1801.LUT_SIZE = 6;
	defparam lut_1801.mask = 64'h37ff37ff1111111f;

	lut_sub lut_1804 ({sk[639], i_9_, i_19_, x224x, x213x, x100x}, x24x);
	defparam lut_1804.LUT_SIZE = 6;
	defparam lut_1804.mask = 64'h37ff37ff55555557;

	lut_sub lut_1807 ({sk[640], i_35_, i_38_, n_n315, x477x, x24x}, x1282x);
	defparam lut_1807.LUT_SIZE = 6;
	defparam lut_1807.mask = 64'h37ff37ff00130000;

	lut_sub lut_1810 ({sk[641], i_10_, i_12_, n_n1438, x23x, x509x}, x1281x);
	defparam lut_1810.LUT_SIZE = 6;
	defparam lut_1810.mask = 64'h37ff37ff00000001;

	lut_sub lut_1812 ({sk[642], x423x, x435x, x330x, x1282x, x1281x}, n_n1847);
	defparam lut_1812.LUT_SIZE = 6;
	defparam lut_1812.mask = 64'h37ff37ff777f7f7f;

	lut_sub lut_1817 ({sk[643], i_25_, i_24_, i_38_, x474x}, x1130x);
	defparam lut_1817.LUT_SIZE = 5;
	defparam lut_1817.mask = 32'h0f0f1000;

	lut_sub lut_1819 ({sk[644], i_25_, i_24_, i_38_, x42x, x77x}, x1129x);
	defparam lut_1819.LUT_SIZE = 6;
	defparam lut_1819.mask = 64'h37ff37ff01000000;

	lut_sub lut_1821 ({sk[645], i_30_, i_32_, n_n1519, x83x, x1129x}, x7614x);
	defparam lut_1821.LUT_SIZE = 6;
	defparam lut_1821.mask = 64'h37ff37ff55575757;

	lut_sub lut_1825 ({sk[646], i_14_, i_13_}, x285x);
	defparam lut_1825.LUT_SIZE = 3;
	defparam lut_1825.mask = 8'h51;

	lut_sub lut_1827 ({sk[647], i_28_, i_29_, n_n1504, x240x, x285x}, x1123x);
	defparam lut_1827.LUT_SIZE = 6;
	defparam lut_1827.mask = 64'h37ff37ff07000000;

	lut_sub lut_1830 ({sk[648], x3x, n_n1300, x298x, x369x, x345x}, x1124x);
	defparam lut_1830.LUT_SIZE = 6;
	defparam lut_1830.mask = 64'h37ff37ff00030507;

	lut_sub lut_1833 ({sk[649], i_34_, x1130x, x7614x, x1123x, x1124x}, n_n1889);
	defparam lut_1833.LUT_SIZE = 6;
	defparam lut_1833.mask = 64'h37ff37ff77777fff;

	lut_sub lut_1838 ({sk[650], i_7_, i_28_}, x409x);
	defparam lut_1838.LUT_SIZE = 3;
	defparam lut_1838.mask = 8'h58;

	lut_sub lut_1840 ({sk[651], i_30_, i_27_, i_23_, i_32_}, x95x);
	defparam lut_1840.LUT_SIZE = 5;
	defparam lut_1840.mask = 32'h0f0f1537;

	lut_sub lut_1844 ({sk[652], i_30_, i_27_, i_16_, i_32_}, x96x);
	defparam lut_1844.LUT_SIZE = 5;
	defparam lut_1844.mask = 32'h0f0f113f;

	lut_sub lut_1848 ({sk[653], i_9_, i_6_, i_11_, i_19_}, x361x);
	defparam lut_1848.LUT_SIZE = 5;
	defparam lut_1848.mask = 32'h0f0f8000;

	lut_sub lut_1850 ({sk[654], i_9_, i_5_, i_6_, i_18_}, x353x);
	defparam lut_1850.LUT_SIZE = 5;
	defparam lut_1850.mask = 32'h0f0f8000;

	lut_sub lut_1852 ({sk[655], n_n1307, n_n787, x361x, x353x}, x4x);
	defparam lut_1852.LUT_SIZE = 5;
	defparam lut_1852.mask = 32'h0f0f0537;

	lut_sub lut_1855 ({sk[656], i_11_, i_19_, n_n1307, n_n841}, x521x);
	defparam lut_1855.LUT_SIZE = 5;
	defparam lut_1855.mask = 32'h0f0f1000;

	lut_sub lut_1857 ({sk[657], i_9_, i_18_, n_n787, n_n1118, x521x}, x801x);
	defparam lut_1857.LUT_SIZE = 6;
	defparam lut_1857.mask = 64'h37ff37ff57555555;

	lut_sub lut_1860 ({sk[658], i_24_, x801x}, x30x);
	defparam lut_1860.LUT_SIZE = 3;
	defparam lut_1860.mask = 8'h54;

	lut_sub lut_1862 ({sk[659], i_25_, i_24_, i_22_, n_n1425}, x313x);
	defparam lut_1862.LUT_SIZE = 5;
	defparam lut_1862.mask = 32'h0f0f4000;

	lut_sub lut_1864 ({sk[660], i_35_, i_38_, x313x}, x56x);
	defparam lut_1864.LUT_SIZE = 4;
	defparam lut_1864.mask = 16'h7710;

	lut_sub lut_1866 ({sk[661], i_10_, i_3_, i_13_, i_12_, i_11_}, x210x);
	defparam lut_1866.LUT_SIZE = 6;
	defparam lut_1866.mask = 64'h37ff37ff00001000;

	lut_sub lut_1868 ({sk[662], i_31_, i_33_, i_35_, i_38_}, x226x);
	defparam lut_1868.LUT_SIZE = 5;
	defparam lut_1868.mask = 32'h0f0f4000;

	lut_sub lut_1870 ({sk[663], i_7_, i_26_, i_24_, i_22_, n_n1431}, x282x);
	defparam lut_1870.LUT_SIZE = 6;
	defparam lut_1870.mask = 64'h37ff37ff40000000;

	lut_sub lut_1872 ({sk[664], i_26_, i_24_, i_38_, n_n1458}, x294x);
	defparam lut_1872.LUT_SIZE = 5;
	defparam lut_1872.mask = 32'h0f0f1000;

	lut_sub lut_1874 ({sk[665], i_13_, i_12_, i_11_, i_19_, n_n1038}, x1451x);
	defparam lut_1874.LUT_SIZE = 6;
	defparam lut_1874.mask = 64'h37ff37ff00150000;

	lut_sub lut_1877 ({sk[666], i_28_, i_26_, i_29_, x30x, x226x}, x1449x);
	defparam lut_1877.LUT_SIZE = 6;
	defparam lut_1877.mask = 64'h37ff37ff10000000;

	lut_sub lut_1879 ({sk[667], i_25_, i_26_, i_24_, i_35_, i_38_}, x81x);
	defparam lut_1879.LUT_SIZE = 6;
	defparam lut_1879.mask = 64'h37ff37ff40000000;

	lut_sub lut_1881 ({sk[668], i_33_, i_35_, i_38_, x277x, n_n1523}, x377x);
	defparam lut_1881.LUT_SIZE = 6;
	defparam lut_1881.mask = 64'h37ff37ff01000000;

	lut_sub lut_1883 ({sk[669], i_13_, i_12_, i_11_, i_19_, n_n1038}, x1444x);
	defparam lut_1883.LUT_SIZE = 6;
	defparam lut_1883.mask = 64'h37ff37ff00150000;

	lut_sub lut_1886 ({sk[670], i_9_, i_12_, i_22_, x262x, x23x}, x591x);
	defparam lut_1886.LUT_SIZE = 6;
	defparam lut_1886.mask = 64'h37ff37ff00300075;

	lut_sub lut_1889 ({sk[671], i_30_, i_28_, i_32_, x81x, x591x}, x1437x);
	defparam lut_1889.LUT_SIZE = 6;
	defparam lut_1889.mask = 64'h37ff37ff10000000;

	lut_sub lut_1891 ({sk[672], n_n584, n_n1033, x56x, x1451x, x414x}, x1450x);
	defparam lut_1891.LUT_SIZE = 6;
	defparam lut_1891.mask = 64'h37ff37ff0707070f;

	lut_sub lut_1895 ({sk[673], i_31_, x42x, x4x, x294x, x1448x}, x7282x);
	defparam lut_1895.LUT_SIZE = 6;
	defparam lut_1895.mask = 64'h37ff37ff55575555;

	lut_sub lut_1898 ({sk[674], i_38_, x204x, x257x, x15x, x1439x}, x7289x);
	defparam lut_1898.LUT_SIZE = 6;
	defparam lut_1898.mask = 64'h37ff37ff55555557;

	lut_sub lut_1901 ({sk[675], i_10_, i_3_, n_n582, x7302x}, x406x);
	defparam lut_1901.LUT_SIZE = 5;
	defparam lut_1901.mask = 32'h0f0f0075;

	lut_sub lut_1904 ({sk[676], i_7_, i_32_, i_38_, x313x}, x249x);
	defparam lut_1904.LUT_SIZE = 5;
	defparam lut_1904.mask = 32'h0f0f1000;

	lut_sub lut_1906 ({sk[677], i_10_, i_3_, n_n586, x406x, x249x}, x1431x);
	defparam lut_1906.LUT_SIZE = 6;
	defparam lut_1906.mask = 64'h37ff37ff11111511;

	lut_sub lut_1909 ({sk[678], i_10_, i_18_, n_n586, x329x}, x1428x);
	defparam lut_1909.LUT_SIZE = 5;
	defparam lut_1909.mask = 32'h0f0f0001;

	lut_sub lut_1911 ({sk[679], i_31_, i_35_, i_38_, i_29_, n_n1478}, x7296x);
	defparam lut_1911.LUT_SIZE = 6;
	defparam lut_1911.mask = 64'h37ff37ff04000000;

	lut_sub lut_1913 ({sk[680], x210x, x281x, x7300x, x7298x, x7299x}, x1430x);
	defparam lut_1913.LUT_SIZE = 6;
	defparam lut_1913.mask = 64'h37ff37ff00030507;

	lut_sub lut_1916 ({sk[681], i_24_, x801x, x1428x, x7296x, x1430x}, x7304x);
	defparam lut_1916.LUT_SIZE = 6;
	defparam lut_1916.mask = 64'h37ff37ff5f7f5f5f;

	lut_sub lut_1920 ({sk[682], i_24_, i_32_, i_31_, n_n1361, x4x}, x354x);
	defparam lut_1920.LUT_SIZE = 6;
	defparam lut_1920.mask = 64'h37ff37ff10000000;

	lut_sub lut_1922 ({sk[683], i_38_, n_n1437, x30x, x624x, x7310x}, x623x);
	defparam lut_1922.LUT_SIZE = 6;
	defparam lut_1922.mask = 64'h37ff37ff1111111f;

	lut_sub lut_1925 ({sk[684], n_n1425, n_n1300, x282x, x406x, x595x}, x1408x);
	defparam lut_1925.LUT_SIZE = 6;
	defparam lut_1925.mask = 64'h37ff37ff00030057;

	lut_sub lut_1928 ({sk[685], i_34_, i_35_, i_38_, x36x, x344x}, x1419x);
	defparam lut_1928.LUT_SIZE = 6;
	defparam lut_1928.mask = 64'h37ff37ff00010000;

	lut_sub lut_1930 ({sk[686], i_31_, x243x, x237x, x4x, x1418x}, x7312x);
	defparam lut_1930.LUT_SIZE = 6;
	defparam lut_1930.mask = 64'h37ff37ff55575555;

	lut_sub lut_1933 ({sk[687], i_29_, n_n1423, n_n416, x266x, n_n706}, x1399x);
	defparam lut_1933.LUT_SIZE = 6;
	defparam lut_1933.mask = 64'h37ff37ff00130000;

	lut_sub lut_1936 ({sk[688], n_n1300, n_n706, x447x, x1400x, x1401x}, x7326x);
	defparam lut_1936.LUT_SIZE = 6;
	defparam lut_1936.mask = 64'h37ff37ff7777777f;

	lut_sub lut_1940 ({sk[689], n_n1466, x266x, x388x, x36x, x26x}, x9218x);
	defparam lut_1940.LUT_SIZE = 6;
	defparam lut_1940.mask = 64'h37ff37fffcfcfca8;

	lut_sub lut_1947 ({sk[690], i_24_, x297x, n_n1288, x1398x, x1406x}, x715x);
	defparam lut_1947.LUT_SIZE = 6;
	defparam lut_1947.mask = 64'h37ff37ff373f3333;

	lut_sub lut_1951 ({sk[691], i_31_, x261x, x276x, x379x, x421x}, x7337x);
	defparam lut_1951.LUT_SIZE = 6;
	defparam lut_1951.mask = 64'h37ff37ff05370033;

	lut_sub lut_1954 ({sk[692], x1390x, x1391x, x1393x, x1394x}, x7338x);
	defparam lut_1954.LUT_SIZE = 5;
	defparam lut_1954.mask = 32'h0f0f7fff;

	lut_sub lut_1959 ({sk[693], i_8_, i_5_, i_6_, n_n1279, n_n1359}, x394x);
	defparam lut_1959.LUT_SIZE = 6;
	defparam lut_1959.mask = 64'h37ff37ff10000000;

	lut_sub lut_1961 ({sk[694], i_35_, i_38_, n_n1353, x11x, x52x}, x1380x);
	defparam lut_1961.LUT_SIZE = 6;
	defparam lut_1961.mask = 64'h37ff37ff00010000;

	lut_sub lut_1963 ({sk[695], i_32_, i_31_, n_n1361, x257x, x207x}, x1381x);
	defparam lut_1963.LUT_SIZE = 6;
	defparam lut_1963.mask = 64'h37ff37ff01000000;

	lut_sub lut_1965 ({sk[696], n_n805, n_n1466, x394x, x1380x, x1381x}, x7346x);
	defparam lut_1965.LUT_SIZE = 6;
	defparam lut_1965.mask = 64'h37ff37ff7777777f;

	lut_sub lut_1969 ({sk[697], i_7_, i_13_, i_32_, n_n1307, x280x}, x346x);
	defparam lut_1969.LUT_SIZE = 6;
	defparam lut_1969.mask = 64'h37ff37ff00100000;

	lut_sub lut_1971 ({sk[698], i_25_, i_34_, i_35_, i_38_, x42x}, x379x);
	defparam lut_1971.LUT_SIZE = 6;
	defparam lut_1971.mask = 64'h37ff37ff01000000;

	lut_sub lut_1973 ({sk[699], i_13_, n_n1361, x313x, x7344x, x37x}, x1383x);
	defparam lut_1973.LUT_SIZE = 6;
	defparam lut_1973.mask = 64'h37ff37ff00070003;

	lut_sub lut_1976 ({sk[700], i_23_, i_31_, i_34_, n_n1216}, x84x);
	defparam lut_1976.LUT_SIZE = 5;
	defparam lut_1976.mask = 32'h0f0f0100;

	lut_sub lut_1978 ({sk[701], i_20_, i_23_, i_17_, x45x}, x319x);
	defparam lut_1978.LUT_SIZE = 5;
	defparam lut_1978.mask = 32'h0f0f4000;

	lut_sub lut_1980 ({sk[702], i_20_, i_7_, i_13_, i_17_, i_16_}, x399x);
	defparam lut_1980.LUT_SIZE = 6;
	defparam lut_1980.mask = 64'h37ff37ff00000080;

	lut_sub lut_1982 ({sk[703], i_23_, i_24_, i_21_, i_34_, n_n1406}, x488x);
	defparam lut_1982.LUT_SIZE = 6;
	defparam lut_1982.mask = 64'h37ff37ff01000000;

	lut_sub lut_1984 ({sk[704], i_23_, i_24_, i_34_, n_n1425, x277x}, x599x);
	defparam lut_1984.LUT_SIZE = 6;
	defparam lut_1984.mask = 64'h37ff37ff35003000;

	lut_sub lut_1987 ({sk[705], n_n1396, n_n1429, n_n1408, x6958x, x488x}, x6963x);
	defparam lut_1987.LUT_SIZE = 6;
	defparam lut_1987.mask = 64'h37ff37ff05550577;

	lut_sub lut_1991 ({sk[706], i_20_, i_25_, i_33_, x302x, x599x}, x1705x);
	defparam lut_1991.LUT_SIZE = 6;
	defparam lut_1991.mask = 64'h37ff37ff00000001;

	lut_sub lut_1993 ({sk[707], i_14_, i_2_, i_16_, n_n1274, x45x}, x1706x);
	defparam lut_1993.LUT_SIZE = 6;
	defparam lut_1993.mask = 64'h37ff37ff00100000;

	lut_sub lut_1995 ({sk[708], i_21_, n_n1438, n_n1302, x372x, x6957x}, x1707x);
	defparam lut_1995.LUT_SIZE = 6;
	defparam lut_1995.mask = 64'h37ff37ff00050037;

	lut_sub lut_1998 ({sk[709], x84x, x399x, x1705x, x1706x, x1707x}, x6964x);
	defparam lut_1998.LUT_SIZE = 6;
	defparam lut_1998.mask = 64'h37ff37ff7f7f7fff;

	lut_sub lut_2003 ({sk[710], i_27_, i_34_, i_37_, x54x, n_n1302}, x317x);
	defparam lut_2003.LUT_SIZE = 6;
	defparam lut_2003.mask = 64'h37ff37ff00010000;

	lut_sub lut_2005 ({sk[711], i_27_, i_28_, i_29_, i_37_}, x365x);
	defparam lut_2005.LUT_SIZE = 5;
	defparam lut_2005.mask = 32'h0f0f4000;

	lut_sub lut_2007 ({sk[712], i_14_, i_17_, i_16_, x50x, x273x}, x1739x);
	defparam lut_2007.LUT_SIZE = 6;
	defparam lut_2007.mask = 64'h37ff37ff10000000;

	lut_sub lut_2009 ({sk[713], n_n1295, n_n1216, n_n1305, n_n269, x1734x}, x6931x);
	defparam lut_2009.LUT_SIZE = 6;
	defparam lut_2009.mask = 64'h37ff37ff55555557;

	lut_sub lut_2012 ({sk[714], n_n1318, n_n437, x1739x, x256x, x6931x}, x6933x);
	defparam lut_2012.LUT_SIZE = 6;
	defparam lut_2012.mask = 64'h37ff37ff55555f7f;

	lut_sub lut_2016 ({sk[715], n_n1295, n_n358, x48x, n_n355, x221x}, x1737x);
	defparam lut_2016.LUT_SIZE = 6;
	defparam lut_2016.mask = 64'h37ff37ff00000357;

	lut_sub lut_2019 ({sk[716], n_n263, n_n363, x317x, x1732x, x6924x}, x6932x);
	defparam lut_2019.LUT_SIZE = 6;
	defparam lut_2019.mask = 64'h37ff37ff33773f7f;

	lut_sub lut_2023 ({sk[717], x6933x, x1737x, x6932x}, n_n1707);
	defparam lut_2023.LUT_SIZE = 4;
	defparam lut_2023.mask = 16'h777f;

	lut_sub lut_2027 ({sk[718], i_34_, i_33_, i_35_, i_37_}, x246x);
	defparam lut_2027.LUT_SIZE = 5;
	defparam lut_2027.mask = 32'h0f0f1000;

	lut_sub lut_2029 ({sk[719], i_20_, i_27_, i_23_, x73x, n_n460}, x63x);
	defparam lut_2029.LUT_SIZE = 6;
	defparam lut_2029.mask = 64'h37ff37ff10000000;

	lut_sub lut_2031 ({sk[720], n_n245, n_n26, x361x, x353x}, x604x);
	defparam lut_2031.LUT_SIZE = 5;
	defparam lut_2031.mask = 32'h0f0f0537;

	lut_sub lut_2034 ({sk[721], i_14_, i_16_, i_37_}, x268x);
	defparam lut_2034.LUT_SIZE = 4;
	defparam lut_2034.mask = 16'h7740;

	lut_sub lut_2036 ({sk[722], i_7_, i_32_, x280x, n_n245, n_n18}, x357x);
	defparam lut_2036.LUT_SIZE = 6;
	defparam lut_2036.mask = 64'h37ff37ff01000000;

	lut_sub lut_2038 ({sk[723], i_13_, i_17_, i_16_, i_33_, n_n1318}, x461x);
	defparam lut_2038.LUT_SIZE = 6;
	defparam lut_2038.mask = 64'h37ff37ff40000000;

	lut_sub lut_2040 ({sk[724], i_9_, i_8_, i_6_, n_n245}, x487x);
	defparam lut_2040.LUT_SIZE = 5;
	defparam lut_2040.mask = 32'h0f0f4000;

	lut_sub lut_2042 ({sk[725], i_20_, i_23_, i_24_, n_n245, x44x}, x88x);
	defparam lut_2042.LUT_SIZE = 6;
	defparam lut_2042.mask = 64'h37ff37ff10000000;

	lut_sub lut_2044 ({sk[726], i_8_, i_14_, i_18_, x263x, x274x}, x1753x);
	defparam lut_2044.LUT_SIZE = 6;
	defparam lut_2044.mask = 64'h37ff37ff10000000;

	lut_sub lut_2046 ({sk[727], i_14_, i_16_, i_32_, n_n21}, x1754x);
	defparam lut_2046.LUT_SIZE = 5;
	defparam lut_2046.mask = 32'h0f0f4000;

	lut_sub lut_2048 ({sk[728], i_32_, x59x, n_n1278, n_n504, n_n1118}, x606x);
	defparam lut_2048.LUT_SIZE = 6;
	defparam lut_2048.mask = 64'h37ff37ff111f1111;

	lut_sub lut_2051 ({sk[729], i_17_, x43x, n_n504, x63x, x353x}, x1750x);
	defparam lut_2051.LUT_SIZE = 6;
	defparam lut_2051.mask = 64'h37ff37ff00010000;

	lut_sub lut_2053 ({sk[730], i_30_, i_27_, i_28_}, x7053x);
	defparam lut_2053.LUT_SIZE = 4;
	defparam lut_2053.mask = 16'h7780;

	lut_sub lut_2055 ({sk[731], i_27_, i_36_, x73x, n_n1431, n_n1254}, x514x);
	defparam lut_2055.LUT_SIZE = 6;
	defparam lut_2055.mask = 64'h37ff37ff00010000;

	lut_sub lut_2057 ({sk[732], i_10_, i_7_, i_13_, i_17_, x10x}, x325x);
	defparam lut_2057.LUT_SIZE = 6;
	defparam lut_2057.mask = 64'h37ff37ff00000004;

	lut_sub lut_2059 ({sk[733], i_10_, i_7_, i_13_, i_12_, x10x}, x328x);
	defparam lut_2059.LUT_SIZE = 6;
	defparam lut_2059.mask = 64'h37ff37ff00000004;

	lut_sub lut_2061 ({sk[734], i_8_, i_6_, i_12_, i_31_, n_n1307}, x360x);
	defparam lut_2061.LUT_SIZE = 6;
	defparam lut_2061.mask = 64'h37ff37ff40000000;

	lut_sub lut_2063 ({sk[735], i_12_, i_17_, x43x, x437x, x16x}, x610x);
	defparam lut_2063.LUT_SIZE = 6;
	defparam lut_2063.mask = 64'h37ff37ff07030500;

	lut_sub lut_2066 ({sk[736], i_21_, n_n461, n_n1406, n_n1141, n_n1213}, x356x);
	defparam lut_2066.LUT_SIZE = 6;
	defparam lut_2066.mask = 64'h37ff37ff00010000;

	lut_sub lut_2068 ({sk[737], i_14_, i_16_, x356x}, x846x);
	defparam lut_2068.LUT_SIZE = 4;
	defparam lut_2068.mask = 16'h7740;

	lut_sub lut_2070 ({sk[738], i_28_, i_32_, i_34_, i_29_, n_n1018}, x7889x);
	defparam lut_2070.LUT_SIZE = 6;
	defparam lut_2070.mask = 64'h37ff37ff04000000;

	lut_sub lut_2072 ({sk[739], i_32_, i_31_, i_33_, i_35_, i_38_}, n_n1149);
	defparam lut_2072.LUT_SIZE = 6;
	defparam lut_2072.mask = 64'h37ff37ff40000000;

	lut_sub lut_2074 ({sk[740], i_28_, i_24_, i_34_, i_29_}, x447x);
	defparam lut_2074.LUT_SIZE = 5;
	defparam lut_2074.mask = 32'h0f0f2000;

	lut_sub lut_2076 ({sk[741], i_13_, i_12_, x292x, n_n1118, n_n1058}, x422x);
	defparam lut_2076.LUT_SIZE = 6;
	defparam lut_2076.mask = 64'h37ff37ff01000000;

	lut_sub lut_2078 ({sk[742], i_13_, i_18_, x11x, n_n1033}, x434x);
	defparam lut_2078.LUT_SIZE = 5;
	defparam lut_2078.mask = 32'h0f0f0100;

	lut_sub lut_2080 ({sk[743], i_13_, i_18_, x11x, n_n1033, x422x}, x21x);
	defparam lut_2080.LUT_SIZE = 6;
	defparam lut_2080.mask = 64'h37ff37ff55575555;

	lut_sub lut_2083 ({sk[744], n_n1118, n_n1279, n_n1048, x208x, n_n1028}, x28x);
	defparam lut_2083.LUT_SIZE = 6;
	defparam lut_2083.mask = 64'h37ff37ff1111111f;

	lut_sub lut_2086 ({sk[745], i_8_, i_33_, n_n1361, n_n1523, n_n1345}, x235x);
	defparam lut_2086.LUT_SIZE = 6;
	defparam lut_2086.mask = 64'h37ff37ff01000000;

	lut_sub lut_2088 ({sk[746], i_25_, i_24_, i_19_, i_35_, i_38_}, x371x);
	defparam lut_2088.LUT_SIZE = 6;
	defparam lut_2088.mask = 64'h37ff37ff04000000;

	lut_sub lut_2090 ({sk[747], i_13_, i_12_, i_11_, i_18_, i_19_}, x7302x);
	defparam lut_2090.LUT_SIZE = 6;
	defparam lut_2090.mask = 64'h37ff37ff00130000;

	lut_sub lut_2093 ({sk[748], i_10_, i_3_, n_n586, x235x, x406x}, x1265x);
	defparam lut_2093.LUT_SIZE = 6;
	defparam lut_2093.mask = 64'h37ff37ff11111311;

	lut_sub lut_2096 ({sk[749], n_n1486, x520x, x21x, x28x, x371x}, x7467x);
	defparam lut_2096.LUT_SIZE = 6;
	defparam lut_2096.mask = 64'h37ff37ff000f111f;

	lut_sub lut_2099 ({sk[750], x213x, x7420x, n_n338, x1265x, x7467x}, n_n1846);
	defparam lut_2099.LUT_SIZE = 6;
	defparam lut_2099.mask = 64'h37ff37ff7777777f;

	lut_sub lut_2103 ({sk[751], i_30_, i_32_, i_31_, i_34_, x42x}, x616x);
	defparam lut_2103.LUT_SIZE = 6;
	defparam lut_2103.mask = 64'h37ff37ff01111111;

	lut_sub lut_2107 ({sk[752], i_12_, i_24_, i_17_, x285x, x616x}, x1107x);
	defparam lut_2107.LUT_SIZE = 6;
	defparam lut_2107.mask = 64'h37ff37ff11001500;

	lut_sub lut_2110 ({sk[753], i_12_, i_17_, i_29_, x61x, x285x}, x1105x);
	defparam lut_2110.LUT_SIZE = 6;
	defparam lut_2110.mask = 64'h37ff37ff01010103;

	lut_sub lut_2113 ({sk[754], i_21_, i_22_, x372x, x1105x}, x7625x);
	defparam lut_2113.LUT_SIZE = 5;
	defparam lut_2113.mask = 32'h0f0f5575;

	lut_sub lut_2116 ({sk[755], i_30_, i_27_, i_16_, i_32_}, x35x);
	defparam lut_2116.LUT_SIZE = 5;
	defparam lut_2116.mask = 32'h0f0f151f;

	lut_sub lut_2120 ({sk[756], i_30_, i_27_, i_23_, i_16_, i_32_}, x618x);
	defparam lut_2120.LUT_SIZE = 6;
	defparam lut_2120.mask = 64'h0fff0fff15553fff;

	lut_sub lut_2127 ({sk[757], i_24_, n_n1511, x83x, x620x, x7629x}, x1097x);
	defparam lut_2127.LUT_SIZE = 6;
	defparam lut_2127.mask = 64'h0fff0fff03570000;

	lut_sub lut_2130 ({sk[758], i_28_, i_26_, x3x, n_n1519, x1093x}, x7631x);
	defparam lut_2130.LUT_SIZE = 6;
	defparam lut_2130.mask = 64'h0fff0fff57555555;

	lut_sub lut_2133 ({sk[759], x42x, n_n1504, n_n1251, x214x, x618x}, x7632x);
	defparam lut_2133.LUT_SIZE = 6;
	defparam lut_2133.mask = 64'h0fff0fff111111f1;

	lut_sub lut_2136 ({sk[760], x1107x, x7625x, x1097x, x7631x, x7632x}, n_n1837);
	defparam lut_2136.LUT_SIZE = 6;
	defparam lut_2136.mask = 64'h0fff0fff7fffffff;

	lut_sub lut_2142 ({sk[761], i_28_, i_25_, i_26_, i_38_}, x311x);
	defparam lut_2142.LUT_SIZE = 5;
	defparam lut_2142.mask = 32'h55574000;

	lut_sub lut_2144 ({sk[762], i_28_, i_25_, i_26_, i_22_}, x78x);
	defparam lut_2144.LUT_SIZE = 5;
	defparam lut_2144.mask = 32'h55578000;

	lut_sub lut_2146 ({sk[763], i_30_, i_24_, i_38_, x13x, x78x}, x329x);
	defparam lut_2146.LUT_SIZE = 6;
	defparam lut_2146.mask = 64'h0fff0fff01000000;

	lut_sub lut_2148 ({sk[764], i_11_, i_18_, i_19_, x60x, x14x}, x36x);
	defparam lut_2148.LUT_SIZE = 6;
	defparam lut_2148.mask = 64'h0fff0fff73503300;

	lut_sub lut_2151 ({sk[765], i_28_, i_32_, i_33_, i_29_}, x344x);
	defparam lut_2151.LUT_SIZE = 5;
	defparam lut_2151.mask = 32'h55578000;

	lut_sub lut_2153 ({sk[766], n_n1307, n_n787, x361x, x353x}, x624x);
	defparam lut_2153.LUT_SIZE = 5;
	defparam lut_2153.mask = 32'h55570537;

	lut_sub lut_2156 ({sk[767], i_25_, i_24_, i_38_, n_n1422}, x7310x);
	defparam lut_2156.LUT_SIZE = 5;
	defparam lut_2156.mask = 32'h55571000;

	lut_sub lut_2158 ({sk[768], i_5_, i_13_, i_4_, i_2_, n_n841}, x421x);
	defparam lut_2158.LUT_SIZE = 6;
	defparam lut_2158.mask = 64'h0fff0fff00400000;

	lut_sub lut_2160 ({sk[769], i_28_, i_32_, i_29_, x238x, x335x}, x1374x);
	defparam lut_2160.LUT_SIZE = 6;
	defparam lut_2160.mask = 64'h0fff0fff10000000;

	lut_sub lut_2162 ({sk[770], i_10_, i_32_, n_n1307, n_n1100, x379x}, x9233x);
	defparam lut_2162.LUT_SIZE = 6;
	defparam lut_2162.mask = 64'h0fff0ffffeffffff;

	lut_sub lut_2174 ({sk[771], i_9_, i_22_, x5x, x349x, x343x}, x714x);
	defparam lut_2174.LUT_SIZE = 6;
	defparam lut_2174.mask = 64'h0fff0fff55007f3f;

	lut_sub lut_2178 ({sk[772], i_30_, i_28_, i_2_, i_32_, x81x}, x7352x);
	defparam lut_2178.LUT_SIZE = 6;
	defparam lut_2178.mask = 64'h0fff0fff40000000;

	lut_sub lut_2180 ({sk[773], i_32_, i_35_, i_38_, x78x, x327x}, x1375x);
	defparam lut_2180.LUT_SIZE = 6;
	defparam lut_2180.mask = 64'h0fff0fff01000000;

	lut_sub lut_2182 ({sk[774], i_9_, i_10_, i_6_, n_n1307}, x207x);
	defparam lut_2182.LUT_SIZE = 5;
	defparam lut_2182.mask = 32'h55574000;

	lut_sub lut_2184 ({sk[775], i_5_, i_4_, i_2_, n_n839}, x218x);
	defparam lut_2184.LUT_SIZE = 5;
	defparam lut_2184.mask = 32'h55574000;

	lut_sub lut_2186 ({sk[776], i_25_, i_24_, i_34_, i_35_, i_38_}, x238x);
	defparam lut_2186.LUT_SIZE = 6;
	defparam lut_2186.mask = 64'h0fff0fff04000000;

	lut_sub lut_2188 ({sk[777], i_35_, i_38_, x42x, x14x, n_n1311}, x310x);
	defparam lut_2188.LUT_SIZE = 6;
	defparam lut_2188.mask = 64'h0fff0fff00000001;

	lut_sub lut_2190 ({sk[778], i_34_, i_35_, i_38_, n_n1423}, x315x);
	defparam lut_2190.LUT_SIZE = 5;
	defparam lut_2190.mask = 32'h55570010;

	lut_sub lut_2192 ({sk[779], i_34_, i_33_, i_35_, i_38_, x42x}, x387x);
	defparam lut_2192.LUT_SIZE = 6;
	defparam lut_2192.mask = 64'h0fff0fff01000000;

	lut_sub lut_2194 ({sk[780], i_10_, i_5_, i_4_, i_2_, n_n841}, x408x);
	defparam lut_2194.LUT_SIZE = 6;
	defparam lut_2194.mask = 64'h0fff0fff40000000;

	lut_sub lut_2196 ({sk[781], i_9_, i_3_, i_13_, i_11_}, x343x);
	defparam lut_2196.LUT_SIZE = 5;
	defparam lut_2196.mask = 32'h55570040;

	lut_sub lut_2198 ({sk[782], i_9_, i_8_, i_2_, n_n735, x343x}, x7375x);
	defparam lut_2198.LUT_SIZE = 6;
	defparam lut_2198.mask = 64'h0fff0fff50007000;

	lut_sub lut_2201 ({sk[783], i_10_, i_13_, x73x, n_n1128, x41x}, x1349x);
	defparam lut_2201.LUT_SIZE = 6;
	defparam lut_2201.mask = 64'h0fff0fff01010001;

	lut_sub lut_2204 ({sk[784], i_32_, i_31_, i_29_, n_n1497, x207x}, x1351x);
	defparam lut_2204.LUT_SIZE = 6;
	defparam lut_2204.mask = 64'h0fff0fff10000000;

	lut_sub lut_2206 ({sk[785], i_26_, i_32_, x42x, n_n849, x327x}, x9217x);
	defparam lut_2206.LUT_SIZE = 6;
	defparam lut_2206.mask = 64'h0fff0ffff8fcffff;

	lut_sub lut_2211 ({sk[786], i_32_, i_31_, i_29_, x509x, x218x}, x1344x);
	defparam lut_2211.LUT_SIZE = 6;
	defparam lut_2211.mask = 64'h0fff0fff10000000;

	lut_sub lut_2213 ({sk[787], i_35_, i_38_, i_29_, n_n1478, n_n849}, x1345x);
	defparam lut_2213.LUT_SIZE = 6;
	defparam lut_2213.mask = 64'h0fff0fff00100000;

	lut_sub lut_2215 ({sk[788], i_28_, i_31_, i_29_, x207x, x270x}, x1346x);
	defparam lut_2215.LUT_SIZE = 6;
	defparam lut_2215.mask = 64'h0fff0fff10000000;

	lut_sub lut_2217 ({sk[789], i_32_, n_n1361, x11x, x71x, n_n1359}, x1348x);
	defparam lut_2217.LUT_SIZE = 6;
	defparam lut_2217.mask = 64'h0fff0fff00010000;

	lut_sub lut_2219 ({sk[790], i_32_, i_38_, n_n1478, x14x, n_n1191}, x1334x);
	defparam lut_2219.LUT_SIZE = 6;
	defparam lut_2219.mask = 64'h0fff0fff00010000;

	lut_sub lut_2221 ({sk[791], i_30_, i_24_}, x278x);
	defparam lut_2221.LUT_SIZE = 3;
	defparam lut_2221.mask = 8'h58;

	lut_sub lut_2223 ({sk[792], i_30_, x42x, n_n1422, n_n998, x18x}, x1330x);
	defparam lut_2223.LUT_SIZE = 6;
	defparam lut_2223.mask = 64'h0fff0fff00010000;

	lut_sub lut_2225 ({sk[793], i_13_, i_11_, i_18_, n_n1038, n_n1033}, x425x);
	defparam lut_2225.LUT_SIZE = 6;
	defparam lut_2225.mask = 64'h0fff0fff05370000;

	lut_sub lut_2228 ({sk[794], i_13_, i_18_, i_19_, n_n1038, n_n1028}, x454x);
	defparam lut_2228.LUT_SIZE = 6;
	defparam lut_2228.mask = 64'h0fff0fff03070005;

	lut_sub lut_2231 ({sk[795], i_27_, i_28_, i_31_, i_34_, i_29_}, x320x);
	defparam lut_2231.LUT_SIZE = 6;
	defparam lut_2231.mask = 64'h0fff0fff02000000;

	lut_sub lut_2233 ({sk[796], i_14_, i_35_, i_37_}, x416x);
	defparam lut_2233.LUT_SIZE = 4;
	defparam lut_2233.mask = 16'h5740;

	lut_sub lut_2235 ({sk[797], i_32_, i_31_, i_33_}, x6967x);
	defparam lut_2235.LUT_SIZE = 4;
	defparam lut_2235.mask = 16'h5780;

	lut_sub lut_2237 ({sk[798], i_14_, i_28_, i_23_, i_24_, i_29_}, x6970x);
	defparam lut_2237.LUT_SIZE = 6;
	defparam lut_2237.mask = 64'h0fff0fff80000000;

	lut_sub lut_2239 ({sk[799], x54x, n_n1489, n_n1438, x6967x, x6970x}, x631x);
	defparam lut_2239.LUT_SIZE = 6;
	defparam lut_2239.mask = 64'h0fff0fff05050537;

	lut_sub lut_2242 ({sk[800], i_32_, i_31_, n_n1489, x452x, x416x}, x1715x);
	defparam lut_2242.LUT_SIZE = 6;
	defparam lut_2242.mask = 64'h0fff0fff01000000;

	lut_sub lut_2244 ({sk[801], i_23_, i_24_, i_16_, n_n1372, x320x}, x1717x);
	defparam lut_2244.LUT_SIZE = 6;
	defparam lut_2244.mask = 64'h0fff0fff10000000;

	lut_sub lut_2246 ({sk[802], i_7_, n_n1295, x631x, x1715x, x1717x}, x6976x);
	defparam lut_2246.LUT_SIZE = 6;
	defparam lut_2246.mask = 64'h0fff0fff777f7777;

	lut_sub lut_2250 ({sk[803], i_13_, i_2_, i_16_, n_n1274, x45x}, x1718x);
	defparam lut_2250.LUT_SIZE = 6;
	defparam lut_2250.mask = 64'h0fff0fff00100000;

	lut_sub lut_2252 ({sk[804], i_17_, x43x, n_n1396, x6958x, x488x}, x1720x);
	defparam lut_2252.LUT_SIZE = 6;
	defparam lut_2252.mask = 64'h0fff0fff00570000;

	lut_sub lut_2255 ({sk[805], n_n1404, n_n1408, x40x, x1718x, x1720x}, x6977x);
	defparam lut_2255.LUT_SIZE = 6;
	defparam lut_2255.mask = 64'h0fff0fff777f7f7f;

	lut_sub lut_2260 ({sk[806], i_34_, i_35_, i_37_}, x248x);
	defparam lut_2260.LUT_SIZE = 4;
	defparam lut_2260.mask = 16'h5704;

	lut_sub lut_2262 ({sk[807], i_10_, i_14_, i_16_}, x334x);
	defparam lut_2262.LUT_SIZE = 4;
	defparam lut_2262.mask = 16'h5780;

	lut_sub lut_2264 ({sk[808], i_17_, i_32_, i_35_, i_37_, x10x}, x303x);
	defparam lut_2264.LUT_SIZE = 6;
	defparam lut_2264.mask = 64'h0fff0fff10000000;

	lut_sub lut_2266 ({sk[809], i_10_, n_n1307, x280x, n_n839, x303x}, x1730x);
	defparam lut_2266.LUT_SIZE = 6;
	defparam lut_2266.mask = 64'h0fff0fff00150011;

	lut_sub lut_2269 ({sk[810], i_27_, i_23_, i_24_, n_n1302, x312x}, x1728x);
	defparam lut_2269.LUT_SIZE = 6;
	defparam lut_2269.mask = 64'h0fff0fff10000000;

	lut_sub lut_2271 ({sk[811], i_10_, i_13_, i_35_, i_37_, x10x}, x6935x);
	defparam lut_2271.LUT_SIZE = 6;
	defparam lut_2271.mask = 64'h0fff0fff10100010;

	lut_sub lut_2274 ({sk[812], i_29_, n_n793, n_n263, x246x}, x1724x);
	defparam lut_2274.LUT_SIZE = 5;
	defparam lut_2274.mask = 32'h55570100;

	lut_sub lut_2276 ({sk[813], i_23_, x43x, n_n1307, n_n1306, x492x}, x1727x);
	defparam lut_2276.LUT_SIZE = 6;
	defparam lut_2276.mask = 64'h0fff0fff00010000;

	lut_sub lut_2278 ({sk[814], x217x, x6935x, x1724x, x1727x}, x6942x);
	defparam lut_2278.LUT_SIZE = 5;
	defparam lut_2278.mask = 32'h5557777f;

	lut_sub lut_2282 ({sk[815], n_n1216, n_n1305, n_n329, x248x, x1728x}, x1725x);
	defparam lut_2282.LUT_SIZE = 6;
	defparam lut_2282.mask = 64'h0fff0fff11111113;

	lut_sub lut_2285 ({sk[816], i_33_, n_n1318, x312x, x67x, x1730x}, x1726x);
	defparam lut_2285.LUT_SIZE = 6;
	defparam lut_2285.mask = 64'h0fff0fff11131111;

	lut_sub lut_2288 ({sk[817], x6942x, x1725x, x1726x}, n_n1706);
	defparam lut_2288.LUT_SIZE = 4;
	defparam lut_2288.mask = 16'h577f;

	lut_sub lut_2292 ({sk[818], i_8_, x60x, n_n132, x15x, x431x}, x31x);
	defparam lut_2292.LUT_SIZE = 6;
	defparam lut_2292.mask = 64'h0fff0fff111f1111;

	lut_sub lut_2295 ({sk[819], i_20_, i_23_, i_24_, i_29_, n_n1441}, x274x);
	defparam lut_2295.LUT_SIZE = 6;
	defparam lut_2295.mask = 64'h0fff0fff10000000;

	lut_sub lut_2297 ({sk[820], i_11_, i_19_, x242x, x14x, x268x}, x351x);
	defparam lut_2297.LUT_SIZE = 6;
	defparam lut_2297.mask = 64'h0fff0fff01000000;

	lut_sub lut_2299 ({sk[821], i_18_, i_37_, x10x, x242x, x60x}, x1574x);
	defparam lut_2299.LUT_SIZE = 6;
	defparam lut_2299.mask = 64'h0fff0fff00010000;

	lut_sub lut_2301 ({sk[822], i_14_, i_13_, i_37_, x233x}, x1568x);
	defparam lut_2301.LUT_SIZE = 5;
	defparam lut_2301.mask = 32'h55570100;

	lut_sub lut_2303 ({sk[823], i_14_, i_13_, i_16_, i_37_, x314x}, x1570x);
	defparam lut_2303.LUT_SIZE = 6;
	defparam lut_2303.mask = 64'h0fff0fff00100000;

	lut_sub lut_2305 ({sk[824], x59x, n_n841, n_n504, x45x, x314x}, x9228x);
	defparam lut_2305.LUT_SIZE = 6;
	defparam lut_2305.mask = 64'h0fff0ffffffcaaa8;

	lut_sub lut_2312 ({sk[825], i_20_, x242x, n_n301, x1570x, x9228x}, x1569x);
	defparam lut_2312.LUT_SIZE = 6;
	defparam lut_2312.mask = 64'h0fff0fff003b0000;

	lut_sub lut_2315 ({sk[826], i_14_, i_37_, x378x, x31x}, x1566x);
	defparam lut_2315.LUT_SIZE = 5;
	defparam lut_2315.mask = 32'h55570100;

	lut_sub lut_2317 ({sk[827], i_32_, n_n853, x461x, x88x, x1565x}, x7132x);
	defparam lut_2317.LUT_SIZE = 6;
	defparam lut_2317.mask = 64'h0fff0fff55575555;

	lut_sub lut_2320 ({sk[828], n_n245, x1568x, x1569x, x1566x, x7132x}, n_n1697);
	defparam lut_2320.LUT_SIZE = 6;
	defparam lut_2320.mask = 64'h0fff0fff77777fff;

	lut_sub lut_2325 ({sk[829], i_14_, n_n1318, n_n1311, x513x, x464x}, x9224x);
	defparam lut_2325.LUT_SIZE = 6;
	defparam lut_2325.mask = 64'h0fff0fffffa8fffc;

	lut_sub lut_2331 ({sk[830], n_n1404, n_n1390, n_n1391, x252x, x320x}, x9225x);
	defparam lut_2331.LUT_SIZE = 6;
	defparam lut_2331.mask = 64'h0fff0ffffffaccc8;

	lut_sub lut_2338 ({sk[831], i_29_, x302x, x441x, x9224x, x9225x}, x6991x);
	defparam lut_2338.LUT_SIZE = 6;
	defparam lut_2338.mask = 64'h0fff0fffeeeeeeef;

	lut_sub lut_2342 ({sk[832], i_32_, i_34_, i_33_, i_35_, i_37_}, x499x);
	defparam lut_2342.LUT_SIZE = 6;
	defparam lut_2342.mask = 64'h0fff0fff00400000;

	lut_sub lut_2344 ({sk[833], i_7_, i_31_, i_34_, x10x, x48x}, x1699x);
	defparam lut_2344.LUT_SIZE = 6;
	defparam lut_2344.mask = 64'h0fff0fff00000001;

	lut_sub lut_2346 ({sk[834], n_n1433, n_n1429, n_n1312, x40x, x6984x}, x6987x);
	defparam lut_2346.LUT_SIZE = 6;
	defparam lut_2346.mask = 64'h0fff0fff00330537;

	lut_sub lut_2349 ({sk[835], x419x, x6991x, x499x, x1699x, x6987x}, n_n1720);
	defparam lut_2349.LUT_SIZE = 6;
	defparam lut_2349.mask = 64'h0fff0fff77ff7fff;

	lut_sub lut_2354 ({sk[836], x6963x, x6964x, x6976x, x6977x}, x6992x);
	defparam lut_2354.LUT_SIZE = 5;
	defparam lut_2354.mask = 32'h55577fff;

	lut_sub lut_2359 ({sk[837], i_20_, i_23_, i_24_, x485x}, x322x);
	defparam lut_2359.LUT_SIZE = 5;
	defparam lut_2359.mask = 32'h55570040;

	lut_sub lut_2361 ({sk[838], n_n1397, n_n1377, n_n1251, x318x, x661x}, x658x);
	defparam lut_2361.LUT_SIZE = 6;
	defparam lut_2361.mask = 64'h0fff0fff00330537;

	lut_sub lut_2364 ({sk[839], n_n1404, x82x, n_n1499, x322x, x658x}, x7002x);
	defparam lut_2364.LUT_SIZE = 6;
	defparam lut_2364.mask = 64'h0fff0fff050537ff;

	lut_sub lut_2368 ({sk[840], i_8_, n_n1441, x10x, x74x, x342x}, x660x);
	defparam lut_2368.LUT_SIZE = 6;
	defparam lut_2368.mask = 64'h0fff0fff03570055;

	lut_sub lut_2371 ({sk[841], i_30_, i_35_, i_29_, i_37_}, x6994x);
	defparam lut_2371.LUT_SIZE = 5;
	defparam lut_2371.mask = 32'h55574000;

	lut_sub lut_2373 ({sk[842], i_13_, i_12_, i_16_, x432x}, x1690x);
	defparam lut_2373.LUT_SIZE = 5;
	defparam lut_2373.mask = 32'h55574000;

	lut_sub lut_2375 ({sk[843], n_n1443, x252x, x660x, x6994x, x1690x}, x7003x);
	defparam lut_2375.LUT_SIZE = 6;
	defparam lut_2375.mask = 64'h0fff0fff575757ff;

	lut_sub lut_2379 ({sk[844], i_27_, n_n1429, x42x, x6944x, x247x}, x1682x);
	defparam lut_2379.LUT_SIZE = 6;
	defparam lut_2379.mask = 64'h0fff0fff00570055;

	lut_sub lut_2382 ({sk[845], i_14_, i_12_, i_16_, x432x, x1682x}, x7012x);
	defparam lut_2382.LUT_SIZE = 6;
	defparam lut_2382.mask = 64'h0fff0fff75555555;

	lut_sub lut_2385 ({sk[846], i_8_, n_n1375, x10x, x48x, x342x}, x703x);
	defparam lut_2385.LUT_SIZE = 6;
	defparam lut_2385.mask = 64'h0fff0fff03570055;

	lut_sub lut_2388 ({sk[847], i_31_, i_37_, x3x, x8x, x67x}, x1681x);
	defparam lut_2388.LUT_SIZE = 6;
	defparam lut_2388.mask = 64'h0fff0fff00000010;

	lut_sub lut_2390 ({sk[848], n_n1443, x13x, x260x, x247x, x524x}, x9222x);
	defparam lut_2390.LUT_SIZE = 6;
	defparam lut_2390.mask = 64'h0fff0ffffffaccc8;

	lut_sub lut_2397 ({sk[849], i_30_, x248x, x703x, x1681x, x9222x}, x7013x);
	defparam lut_2397.LUT_SIZE = 6;
	defparam lut_2397.mask = 64'h0fff0fffbbbfbbbb;

	lut_sub lut_2401 ({sk[850], x7002x, x7003x, x7012x, x7013x}, x7023x);
	defparam lut_2401.LUT_SIZE = 5;
	defparam lut_2401.mask = 32'h55577fff;

	lut_sub lut_2406 ({sk[851], i_7_, i_31_, x43x, x74x, x90x}, n_n1723);
	defparam lut_2406.LUT_SIZE = 6;
	defparam lut_2406.mask = 64'h0fff0fff55555557;

	lut_sub lut_2409 ({sk[852], i_23_, i_21_, i_22_, x45x}, x55x);
	defparam lut_2409.LUT_SIZE = 5;
	defparam lut_2409.mask = 32'h55570400;

	lut_sub lut_2411 ({sk[853], i_31_, n_n1441, n_n1390, n_n1372, n_n1391}, x1653x);
	defparam lut_2411.LUT_SIZE = 6;
	defparam lut_2411.mask = 64'h0fff0fff00000007;

	lut_sub lut_2414 ({sk[854], i_7_, i_31_, x10x, x74x, x127x}, x7034x);
	defparam lut_2414.LUT_SIZE = 6;
	defparam lut_2414.mask = 64'h0fff0fff55555557;

	lut_sub lut_2417 ({sk[855], i_12_, i_17_, x10x, x308x, x309x}, x9223x);
	defparam lut_2417.LUT_SIZE = 6;
	defparam lut_2417.mask = 64'h0fff0ffff8f8f8ff;

	lut_sub lut_2421 ({sk[856], n_n1443, x55x, x1653x, x7034x, x9223x}, n_n1722);
	defparam lut_2421.LUT_SIZE = 6;
	defparam lut_2421.mask = 64'h0fff0fffbfbfbfff;

	lut_sub lut_2426 ({sk[857], i_23_, i_21_, i_22_}, x7033x);
	defparam lut_2426.LUT_SIZE = 4;
	defparam lut_2426.mask = 16'h5720;

	lut_sub lut_2428 ({sk[858], n_n1429, x8x, x45x, x196x, x7033x}, x7040x);
	defparam lut_2428.LUT_SIZE = 6;
	defparam lut_2428.mask = 64'h0fff0fff33373737;

	lut_sub lut_2432 ({sk[859], n_n1334, x48x, n_n1401, x104x, x126x}, x7041x);
	defparam lut_2432.LUT_SIZE = 6;
	defparam lut_2432.mask = 64'h0fff0fff7777777f;

	lut_sub lut_2436 ({sk[860], n_n1408, x82x, x322x, x1667x, x1668x}, x7020x);
	defparam lut_2436.LUT_SIZE = 6;
	defparam lut_2436.mask = 64'h0fff0fff77777fff;

	lut_sub lut_2441 ({sk[861], i_20_, n_n1404, x488x, x1672x, x9221x}, x7021x);
	defparam lut_2441.LUT_SIZE = 6;
	defparam lut_2441.mask = 64'h0fff0fff333fbbbf;

	lut_sub lut_2445 ({sk[862], i_10_, i_7_, i_11_, i_21_, i_19_}, x440x);
	defparam lut_2445.LUT_SIZE = 6;
	defparam lut_2445.mask = 64'h0fff0fff00000020;

	lut_sub lut_2447 ({sk[863], i_9_, i_10_, i_24_, n_n1307, n_n1303}, n_n1086);
	defparam lut_2447.LUT_SIZE = 6;
	defparam lut_2447.mask = 64'h0fff0fff10000000;

	lut_sub lut_2449 ({sk[864], i_30_, i_16_, i_34_}, x143x);
	defparam lut_2449.LUT_SIZE = 4;
	defparam lut_2449.mask = 16'h5701;

	lut_sub lut_2451 ({sk[865], i_23_, x3x, x298x, n_n1497, x83x}, x1087x);
	defparam lut_2451.LUT_SIZE = 6;
	defparam lut_2451.mask = 64'h0fff0fff00000537;

	lut_sub lut_2454 ({sk[866], i_24_, x42x, n_n1334, x103x, x143x}, x9235x);
	defparam lut_2454.LUT_SIZE = 6;
	defparam lut_2454.mask = 64'h0fff0fffffa8ffff;

	lut_sub lut_2465 ({sk[867], i_24_, i_34_, x42x, x35x, x9235x}, x7635x);
	defparam lut_2465.LUT_SIZE = 6;
	defparam lut_2465.mask = 64'h0fff0fffaaabaaaa;

	lut_sub lut_2468 ({sk[868], i_27_, i_23_, i_16_, i_31_}, x1082x);
	defparam lut_2468.LUT_SIZE = 5;
	defparam lut_2468.mask = 32'h55571555;

	lut_sub lut_2472 ({sk[869], i_28_, i_23_, i_24_, i_34_, i_29_}, x1081x);
	defparam lut_2472.LUT_SIZE = 6;
	defparam lut_2472.mask = 64'h0fff0fff00200000;

	lut_sub lut_2474 ({sk[870], i_30_, i_14_, i_16_, i_33_}, x7636x);
	defparam lut_2474.LUT_SIZE = 5;
	defparam lut_2474.mask = 32'h55570537;

	lut_sub lut_2477 ({sk[871], n_n1497, x35x, x1082x, x1081x, x7636x}, n_n1897);
	defparam lut_2477.LUT_SIZE = 6;
	defparam lut_2477.mask = 64'h0fff0fff33337fff;

	lut_sub lut_2482 ({sk[872], i_9_, i_19_, x224x, x213x, n_n315}, x98x);
	defparam lut_2482.LUT_SIZE = 6;
	defparam lut_2482.mask = 64'h0fff0fff55555557;

	lut_sub lut_2485 ({sk[873], i_33_, i_35_, i_38_, x243x, n_n1497}, x254x);
	defparam lut_2485.LUT_SIZE = 6;
	defparam lut_2485.mask = 64'h0fff0fff01000000;

	lut_sub lut_2487 ({sk[874], i_28_, i_32_, i_29_, n_n1454, n_n1361}, x381x);
	defparam lut_2487.LUT_SIZE = 6;
	defparam lut_2487.mask = 64'h0fff0fff10000000;

	lut_sub lut_2489 ({sk[875], i_28_, i_26_, i_33_, i_29_}, x430x);
	defparam lut_2489.LUT_SIZE = 5;
	defparam lut_2489.mask = 32'h55578000;

	lut_sub lut_2491 ({sk[876], i_13_, i_18_, x11x, n_n1033, x422x}, x7442x);
	defparam lut_2491.LUT_SIZE = 6;
	defparam lut_2491.mask = 64'h0fff0fff55575555;

	lut_sub lut_2494 ({sk[877], i_9_, i_8_, x224x, n_n307, x213x}, x33x);
	defparam lut_2494.LUT_SIZE = 6;
	defparam lut_2494.mask = 64'h0fff0fff33333733;

	lut_sub lut_2497 ({sk[878], i_19_, x12x, x430x, x7442x, x33x}, x1290x);
	defparam lut_2497.LUT_SIZE = 6;
	defparam lut_2497.mask = 64'h0fff0fff00030007;

	lut_sub lut_2500 ({sk[879], n_n1288, x24x, x81x, x98x, x254x}, x7445x);
	defparam lut_2500.LUT_SIZE = 6;
	defparam lut_2500.mask = 64'h0fff0fff1111111f;

	lut_sub lut_2503 ({sk[880], i_25_, i_34_, i_35_, i_38_}, x429x);
	defparam lut_2503.LUT_SIZE = 5;
	defparam lut_2503.mask = 32'h55571000;

	lut_sub lut_2505 ({sk[881], i_9_, i_8_, i_18_, x224x, n_n787}, x231x);
	defparam lut_2505.LUT_SIZE = 6;
	defparam lut_2505.mask = 64'h0fff0fff10000000;

	lut_sub lut_2507 ({sk[882], i_28_, i_22_, i_38_, x73x, n_n1458}, x7450x);
	defparam lut_2507.LUT_SIZE = 6;
	defparam lut_2507.mask = 64'h0fff0fff01000000;

	lut_sub lut_2509 ({sk[883], i_19_, x53x, x422x, x434x, x33x}, x1318x);
	defparam lut_2509.LUT_SIZE = 6;
	defparam lut_2509.mask = 64'h0fff0fff003f007f;

	lut_sub lut_2513 ({sk[884], n_n1361, n_n372, n_n294, n_n371, x476x}, x1317x);
	defparam lut_2513.LUT_SIZE = 6;
	defparam lut_2513.mask = 64'h0fff0fff00001555;

	lut_sub lut_2517 ({sk[885], i_28_, i_32_, x389x, n_n315, x24x}, x1315x);
	defparam lut_2517.LUT_SIZE = 6;
	defparam lut_2517.mask = 64'h0fff0fff07000000;

	lut_sub lut_2520 ({sk[886], n_n294, x229x, n_n371, n_n735, x253x}, x1314x);
	defparam lut_2520.LUT_SIZE = 6;
	defparam lut_2520.mask = 64'h0fff0fff05155555;

	lut_sub lut_2524 ({sk[887], i_34_, i_35_, i_38_, n_n1423, x243x}, x75x);
	defparam lut_2524.LUT_SIZE = 6;
	defparam lut_2524.mask = 64'h0fff0fff00000100;

	lut_sub lut_2526 ({sk[888], i_28_, i_25_, i_34_, i_29_, x12x}, x293x);
	defparam lut_2526.LUT_SIZE = 6;
	defparam lut_2526.mask = 64'h0fff0fff04000000;

	lut_sub lut_2528 ({sk[889], i_13_, x208x, n_n1033, x435x, x293x}, x1309x);
	defparam lut_2528.LUT_SIZE = 6;
	defparam lut_2528.mask = 64'h0fff0fff11151111;

	lut_sub lut_2531 ({sk[890], n_n1225, n_n284, x28x, x371x, x75x}, x7432x);
	defparam lut_2531.LUT_SIZE = 6;
	defparam lut_2531.mask = 64'h0fff0fff00550357;

	lut_sub lut_2534 ({sk[891], i_24_, i_22_, i_35_, i_38_, n_n1478}, x276x);
	defparam lut_2534.LUT_SIZE = 6;
	defparam lut_2534.mask = 64'h0fff0fff10000000;

	lut_sub lut_2536 ({sk[892], i_7_, i_14_, i_13_, i_12_}, x661x);
	defparam lut_2536.LUT_SIZE = 5;
	defparam lut_2536.mask = 32'h555700a8;

	lut_sub lut_2539 ({sk[893], i_27_, i_26_, i_24_, n_n1100, n_n460}, x314x);
	defparam lut_2539.LUT_SIZE = 6;
	defparam lut_2539.mask = 64'h0fff0fff10000000;

	lut_sub lut_2541 ({sk[894], i_20_, i_14_, i_16_, x242x, x314x}, x1562x);
	defparam lut_2541.LUT_SIZE = 6;
	defparam lut_2541.mask = 64'h0fff0fff10000000;

	lut_sub lut_2543 ({sk[895], i_14_, x233x, x1562x, x7138x}, x1556x);
	defparam lut_2543.LUT_SIZE = 5;
	defparam lut_2543.mask = 32'h55571511;

	lut_sub lut_2546 ({sk[896], i_34_, i_37_, x19x, n_n1216, n_n1305}, x1557x);
	defparam lut_2546.LUT_SIZE = 6;
	defparam lut_2546.mask = 64'h0fff0fff00000001;

	lut_sub lut_2548 ({sk[897], n_n132, n_n29, n_n129, n_n130, x317x}, x1559x);
	defparam lut_2548.LUT_SIZE = 6;
	defparam lut_2548.mask = 64'h0fff0fff01010155;

	lut_sub lut_2551 ({sk[898], n_n839, x88x, x303x, x9227x}, x7141x);
	defparam lut_2551.LUT_SIZE = 5;
	defparam lut_2551.mask = 32'h5557aaab;

	lut_sub lut_2554 ({sk[899], x1556x, x1557x, x1559x, x7141x}, n_n1698);
	defparam lut_2554.LUT_SIZE = 5;
	defparam lut_2554.mask = 32'h55577fff;

	lut_sub lut_2559 ({sk[900], i_20_, i_25_, i_23_, n_n1397, x7058x}, x331x);
	defparam lut_2559.LUT_SIZE = 6;
	defparam lut_2559.mask = 64'h0fff0fff00000010;

	lut_sub lut_2561 ({sk[901], i_13_, n_n1375, n_n1322, x77x, x246x}, x1628x);
	defparam lut_2561.LUT_SIZE = 6;
	defparam lut_2561.mask = 64'h0fff0fff00010000;

	lut_sub lut_2563 ({sk[902], i_35_, i_29_, n_n1295, n_n1216, x515x}, x1629x);
	defparam lut_2563.LUT_SIZE = 6;
	defparam lut_2563.mask = 64'h0fff0fff01000000;

	lut_sub lut_2565 ({sk[903], i_27_, i_37_, x42x, n_n1422, n_n608}, x1630x);
	defparam lut_2565.LUT_SIZE = 6;
	defparam lut_2565.mask = 64'h0fff0fff00010000;

	lut_sub lut_2567 ({sk[904], n_n1429, x331x, x1628x, x1629x, x1630x}, x7062x);
	defparam lut_2567.LUT_SIZE = 6;
	defparam lut_2567.mask = 64'h0fff0fff7f7f7fff;

	lut_sub lut_2572 ({sk[905], i_32_, i_34_, i_29_, n_n1216, n_n620}, x1634x);
	defparam lut_2572.LUT_SIZE = 6;
	defparam lut_2572.mask = 64'h0fff0fff00100000;

	lut_sub lut_2574 ({sk[906], i_20_, n_n1404, x65x, x251x, x7057x}, x769x);
	defparam lut_2574.LUT_SIZE = 6;
	defparam lut_2574.mask = 64'h0fff0fff557f5577;

	lut_sub lut_2578 ({sk[907], i_20_, n_n1404, x773x, x1623x, x1625x}, x772x);
	defparam lut_2578.LUT_SIZE = 6;
	defparam lut_2578.mask = 64'h0fff0fff777f7777;

	lut_sub lut_2582 ({sk[908], i_0_, i_35_, i_37_, x772x}, x1619x);
	defparam lut_2582.LUT_SIZE = 5;
	defparam lut_2582.mask = 32'h55571000;

	lut_sub lut_2584 ({sk[909], i_37_, n_n1404, n_n1408, n_n1202, x445x}, x1618x);
	defparam lut_2584.LUT_SIZE = 6;
	defparam lut_2584.mask = 64'h0fff0fff00000111;

	lut_sub lut_2587 ({sk[910], i_28_, i_29_, n_n1369, n_n1318, x515x}, x1620x);
	defparam lut_2587.LUT_SIZE = 6;
	defparam lut_2587.mask = 64'h0fff0fff01000000;

	lut_sub lut_2589 ({sk[911], i_32_, i_29_, n_n1441, n_n1318, n_n608}, x1621x);
	defparam lut_2589.LUT_SIZE = 6;
	defparam lut_2589.mask = 64'h0fff0fff01000000;

	lut_sub lut_2591 ({sk[912], n_n1443, x331x, x1618x, x1620x, x1621x}, x7077x);
	defparam lut_2591.LUT_SIZE = 6;
	defparam lut_2591.mask = 64'h0fff0fff7f7f7fff;

	lut_sub lut_2596 ({sk[913], i_13_, i_12_, i_17_, i_16_}, x29x);
	defparam lut_2596.LUT_SIZE = 5;
	defparam lut_2596.mask = 32'h5557a800;

	lut_sub lut_2599 ({sk[914], i_27_, i_28_, i_26_, i_35_, i_37_}, x366x);
	defparam lut_2599.LUT_SIZE = 6;
	defparam lut_2599.mask = 64'h0fff0fff40000000;

	lut_sub lut_2601 ({sk[915], i_30_, i_31_, i_29_, n_n793}, x445x);
	defparam lut_2601.LUT_SIZE = 5;
	defparam lut_2601.mask = 32'h55570400;

	lut_sub lut_2603 ({sk[916], i_20_, i_13_, i_12_, i_23_, i_16_}, x1616x);
	defparam lut_2603.LUT_SIZE = 6;
	defparam lut_2603.mask = 64'h0fff0fff80000000;

	lut_sub lut_2605 ({sk[917], x43x, n_n1369, n_n1274, n_n1431, x1616x}, x1614x);
	defparam lut_2605.LUT_SIZE = 6;
	defparam lut_2605.mask = 64'h0fff0fff00110013;

	lut_sub lut_2608 ({sk[918], i_8_, i_26_, i_23_, i_24_, x7053x}, x202x);
	defparam lut_2608.LUT_SIZE = 6;
	defparam lut_2608.mask = 64'h0fff0fff40000000;

	lut_sub lut_2610 ({sk[919], i_20_, i_13_, i_17_, i_16_, x202x}, x1615x);
	defparam lut_2610.LUT_SIZE = 6;
	defparam lut_2610.mask = 64'h0fff0fff40000000;

	lut_sub lut_2612 ({sk[920], i_0_, i_33_, n_n1318, x1614x, x1615x}, x1608x);
	defparam lut_2612.LUT_SIZE = 6;
	defparam lut_2612.mask = 64'h0fff0fff07000000;

	lut_sub lut_2615 ({sk[921], i_33_, n_n544, x243x, x366x, x1609x}, x7090x);
	defparam lut_2615.LUT_SIZE = 6;
	defparam lut_2615.mask = 64'h0fff0fff55575555;

	lut_sub lut_2618 ({sk[922], i_37_, n_n363, x273x, x1606x, x1607x}, x7091x);
	defparam lut_2618.LUT_SIZE = 6;
	defparam lut_2618.mask = 64'h0fff0fff7777777f;

	lut_sub lut_2622 ({sk[923], i_27_, i_28_, i_33_}, x7058x);
	defparam lut_2622.LUT_SIZE = 4;
	defparam lut_2622.mask = 16'h5740;

	lut_sub lut_2624 ({sk[924], i_23_, i_34_, i_35_, x7058x}, x505x);
	defparam lut_2624.LUT_SIZE = 5;
	defparam lut_2624.mask = 32'h55571000;

	lut_sub lut_2626 ({sk[925], i_8_, i_13_, i_12_, i_16_, x54x}, x348x);
	defparam lut_2626.LUT_SIZE = 6;
	defparam lut_2626.mask = 64'h0fff0fff40000000;

	lut_sub lut_2628 ({sk[926], i_9_, i_2_, i_29_, n_n1441, x7749x}, x332x);
	defparam lut_2628.LUT_SIZE = 6;
	defparam lut_2628.mask = 64'h0fff0fff00010000;

	lut_sub lut_2630 ({sk[927], i_4_, x79x, x224x, n_n460, n_n1254}, x383x);
	defparam lut_2630.LUT_SIZE = 6;
	defparam lut_2630.mask = 64'h0fff0fff00010000;

	lut_sub lut_2632 ({sk[928], i_10_, i_7_, i_11_, i_19_, x54x}, x393x);
	defparam lut_2632.LUT_SIZE = 6;
	defparam lut_2632.mask = 64'h0fff0fff00000040;

	lut_sub lut_2634 ({sk[929], i_13_, i_16_, x356x}, x838x);
	defparam lut_2634.LUT_SIZE = 4;
	defparam lut_2634.mask = 16'h5740;

	lut_sub lut_2636 ({sk[930], i_27_, i_28_, i_32_, i_29_, n_n1213}, x7902x);
	defparam lut_2636.LUT_SIZE = 6;
	defparam lut_2636.mask = 64'h0fff0fff40000000;

	lut_sub lut_2638 ({sk[931], i_22_, i_33_, i_35_, i_38_, n_n1497}, x390x);
	defparam lut_2638.LUT_SIZE = 6;
	defparam lut_2638.mask = 64'h0fff0fff10000000;

	lut_sub lut_2640 ({sk[932], i_9_, i_8_, i_13_, x208x}, x1279x);
	defparam lut_2640.LUT_SIZE = 5;
	defparam lut_2640.mask = 32'h55570040;

	lut_sub lut_2642 ({sk[933], i_19_, n_n1048, x50x, x20x, x1279x}, x672x);
	defparam lut_2642.LUT_SIZE = 6;
	defparam lut_2642.mask = 64'h0fff0fff3333777f;

	lut_sub lut_2646 ({sk[934], i_30_, i_32_, i_31_, x210x, x390x}, x1275x);
	defparam lut_2646.LUT_SIZE = 6;
	defparam lut_2646.mask = 64'h0fff0fff10000000;

	lut_sub lut_2648 ({sk[935], n_n372, n_n294, n_n371, n_n284, x381x}, x1276x);
	defparam lut_2648.LUT_SIZE = 6;
	defparam lut_2648.mask = 64'h0fff0fff15555555;

	lut_sub lut_2653 ({sk[936], x12x, x430x, x672x, x1275x, x1276x}, n_n1848);
	defparam lut_2653.LUT_SIZE = 6;
	defparam lut_2653.mask = 64'h0fff0fff7777777f;

	lut_sub lut_2657 ({sk[937], n_n372, n_n294, n_n371, n_n284, x254x}, x1269x);
	defparam lut_2657.LUT_SIZE = 6;
	defparam lut_2657.mask = 64'h0fff0fff15555555;

	lut_sub lut_2662 ({sk[938], n_n1486, n_n315, x371x, x381x, x33x}, x7461x);
	defparam lut_2662.LUT_SIZE = 6;
	defparam lut_2662.mask = 64'h0fff0fff00330537;

	lut_sub lut_2665 ({sk[939], x71x, x12x, x21x, x1269x, x7461x}, x7463x);
	defparam lut_2665.LUT_SIZE = 6;
	defparam lut_2665.mask = 64'h0fff0fff7777777f;

	lut_sub lut_2669 ({sk[940], n_n1847, n_n1848, x7463x}, n_n1822);
	defparam lut_2669.LUT_SIZE = 4;
	defparam lut_2669.mask = 16'h577f;

	lut_sub lut_2673 ({sk[941], i_8_, i_31_}, x284x);
	defparam lut_2673.LUT_SIZE = 3;
	defparam lut_2673.mask = 8'h58;

	lut_sub lut_2675 ({sk[942], i_10_, i_11_, n_n584, x1262x}, x1260x);
	defparam lut_2675.LUT_SIZE = 5;
	defparam lut_2675.mask = 32'h55570057;

	lut_sub lut_2678 ({sk[943], n_n735, x405x, x56x, x284x, x1260x}, x1256x);
	defparam lut_2678.LUT_SIZE = 6;
	defparam lut_2678.mask = 64'h0fff0fff01010103;

	lut_sub lut_2681 ({sk[944], n_n372, n_n1225, x253x, x371x, x33x}, x7471x);
	defparam lut_2681.LUT_SIZE = 6;
	defparam lut_2681.mask = 64'h0fff0fff00110f1f;

	lut_sub lut_2684 ({sk[945], x422x, x434x, x293x, x1256x, x7471x}, n_n1844);
	defparam lut_2684.LUT_SIZE = 6;
	defparam lut_2684.mask = 64'h0fff0fff777f7f7f;

	lut_sub lut_2689 ({sk[946], i_25_, i_26_, i_24_, i_32_, n_n1361}, x270x);
	defparam lut_2689.LUT_SIZE = 6;
	defparam lut_2689.mask = 64'h0fff0fff40000000;

	lut_sub lut_2691 ({sk[947], i_3_, i_12_, i_22_, n_n586, x349x}, x679x);
	defparam lut_2691.LUT_SIZE = 6;
	defparam lut_2691.mask = 64'h0fff0fff30750055;

	lut_sub lut_2694 ({sk[948], i_10_, i_12_, x5x, x679x}, x678x);
	defparam lut_2694.LUT_SIZE = 5;
	defparam lut_2694.mask = 32'h55570057;

	lut_sub lut_2697 ({sk[949], i_11_, x11x, n_n1048, x213x, x7425x}, x7475x);
	defparam lut_2697.LUT_SIZE = 6;
	defparam lut_2697.mask = 64'h0fff0fff1111111f;

	lut_sub lut_2700 ({sk[950], n_n307, n_n1345, n_n338, x270x, x678x}, x7476x);
	defparam lut_2700.LUT_SIZE = 6;
	defparam lut_2700.mask = 64'h0fff0fff00110f1f;

	lut_sub lut_2703 ({sk[951], n_n1361, x476x, x98x, x7475x, x7476x}, x7477x);
	defparam lut_2703.LUT_SIZE = 6;
	defparam lut_2703.mask = 64'h0fff0fff5555557f;

	lut_sub lut_2707 ({sk[952], n_n1846, n_n1844, x7477x}, n_n1821);
	defparam lut_2707.LUT_SIZE = 4;
	defparam lut_2707.mask = 16'h577f;

	lut_sub lut_2711 ({sk[953], i_28_, i_32_, i_29_, n_n1307, n_n1100}, x272x);
	defparam lut_2711.LUT_SIZE = 6;
	defparam lut_2711.mask = 64'h0fff0fff10000000;

	lut_sub lut_2713 ({sk[954], i_20_, i_23_, i_24_, n_n1441, x77x}, x251x);
	defparam lut_2713.LUT_SIZE = 6;
	defparam lut_2713.mask = 64'h0fff0fff10000000;

	lut_sub lut_2715 ({sk[955], i_26_, i_23_, i_24_, x7053x, x9231x}, x1602x);
	defparam lut_2715.LUT_SIZE = 6;
	defparam lut_2715.mask = 64'h0fff0fff20000000;

	lut_sub lut_2717 ({sk[956], n_n504, x470x, x202x, x251x, x402x}, x9220x);
	defparam lut_2717.LUT_SIZE = 6;
	defparam lut_2717.mask = 64'h0fff0fffffccfac8;

	lut_sub lut_2724 ({sk[957], x59x, n_n1443, x251x, x1602x, x9220x}, x681x);
	defparam lut_2724.LUT_SIZE = 6;
	defparam lut_2724.mask = 64'h0fff0fffaaaabbbf;

	lut_sub lut_2728 ({sk[958], i_27_, i_28_, i_29_, n_n544, x499x}, x1594x);
	defparam lut_2728.LUT_SIZE = 6;
	defparam lut_2728.mask = 64'h0fff0fff10000000;

	lut_sub lut_2730 ({sk[959], i_35_, i_37_, n_n1369, n_n1288, n_n437}, x1595x);
	defparam lut_2730.LUT_SIZE = 6;
	defparam lut_2730.mask = 64'h0fff0fff00010000;

	lut_sub lut_2732 ({sk[960], i_27_, i_35_, i_37_, x42x, n_n1213}, x7097x);
	defparam lut_2732.LUT_SIZE = 6;
	defparam lut_2732.mask = 64'h0fff0fff01000000;

	lut_sub lut_2734 ({sk[961], n_n1216, n_n1314, n_n1318, x76x, n_n1241}, x1598x);
	defparam lut_2734.LUT_SIZE = 6;
	defparam lut_2734.mask = 64'h0fff0fff00000001;

	lut_sub lut_2736 ({sk[962], n_n195, x1594x, x1595x, x7097x, x1598x}, x7104x);
	defparam lut_2736.LUT_SIZE = 6;
	defparam lut_2736.mask = 64'h0fff0fff5fff7fff;

	lut_sub lut_2741 ({sk[963], i_0_, x681x, x7104x}, n_n1708);
	defparam lut_2741.LUT_SIZE = 4;
	defparam lut_2741.mask = 16'h5775;

	lut_sub lut_2744 ({sk[964], i_11_, i_19_, x54x, n_n1307, x280x}, x484x);
	defparam lut_2744.LUT_SIZE = 6;
	defparam lut_2744.mask = 64'h0fff0fff01000000;

	lut_sub lut_2746 ({sk[965], i_9_, i_18_, x54x, x224x, n_n787}, x489x);
	defparam lut_2746.LUT_SIZE = 6;
	defparam lut_2746.mask = 64'h0fff0fff01000000;

	lut_sub lut_2748 ({sk[966], i_10_, i_13_, x15x, x373x}, x1551x);
	defparam lut_2748.LUT_SIZE = 5;
	defparam lut_2748.mask = 32'h55571000;

	lut_sub lut_2750 ({sk[967], i_32_, n_n1443, x259x, x319x, x274x}, x9226x);
	defparam lut_2750.LUT_SIZE = 6;
	defparam lut_2750.mask = 64'h0fff0ffffca8fcfc;

	lut_sub lut_2757 ({sk[968], n_n1278, n_n301, n_n152, x87x, x9226x}, x7155x);
	defparam lut_2757.LUT_SIZE = 6;
	defparam lut_2757.mask = 64'h0fff0fff00330a3b;

	lut_sub lut_2760 ({sk[969], n_n1216, n_n1318, n_n1241, x498x, x522x}, x1548x);
	defparam lut_2760.LUT_SIZE = 6;
	defparam lut_2760.mask = 64'h0fff0fff00000007;

	lut_sub lut_2763 ({sk[970], n_n853, x88x, x303x, x7x, x7151x}, x7156x);
	defparam lut_2763.LUT_SIZE = 6;
	defparam lut_2763.mask = 64'h0fff0fff1111111f;

	lut_sub lut_2766 ({sk[971], x59x, x1551x, x7155x, x1548x, x7156x}, n_n1699);
	defparam lut_2766.LUT_SIZE = 6;
	defparam lut_2766.mask = 64'h0fff0fff77777fff;

	lut_sub lut_2771 ({sk[972], i_9_, i_12_}, x68x);
	defparam lut_2771.LUT_SIZE = 3;
	defparam lut_2771.mask = 8'h51;

	lut_sub lut_2773 ({sk[973], i_5_, i_4_, i_2_, i_38_, n_n1306}, x206x);
	defparam lut_2773.LUT_SIZE = 6;
	defparam lut_2773.mask = 64'h0fff0fff10000000;

	lut_sub lut_2775 ({sk[974], x72x, x9x, x288x, x124x, x132x}, x7504x);
	defparam lut_2775.LUT_SIZE = 6;
	defparam lut_2775.mask = 64'h0fff0fff7777777f;

	lut_sub lut_2779 ({sk[975], n_n1278, n_n1279, x7492x, x71x, x430x}, x1224x);
	defparam lut_2779.LUT_SIZE = 6;
	defparam lut_2779.mask = 64'h0fff0fff00000007;

	lut_sub lut_2782 ({sk[976], n_n1454, n_n1288, x250x, x329x, x68x}, x9213x);
	defparam lut_2782.LUT_SIZE = 6;
	defparam lut_2782.mask = 64'h0fff0fffeeeeeee0;

	lut_sub lut_2789 ({sk[977], x476x, x477x, x206x, x1224x, x9213x}, x7505x);
	defparam lut_2789.LUT_SIZE = 6;
	defparam lut_2789.mask = 64'h0fff0fffbbbfbfbf;

	lut_sub lut_2794 ({sk[978], i_32_, i_31_, n_n1489, n_n1295, n_n1018}, x216x);
	defparam lut_2794.LUT_SIZE = 6;
	defparam lut_2794.mask = 64'h0fff0fff00010000;

	lut_sub lut_2796 ({sk[979], i_27_, i_23_, i_21_, i_35_, n_n1326}, x247x);
	defparam lut_2796.LUT_SIZE = 6;
	defparam lut_2796.mask = 64'h0fff0fff01000000;

	lut_sub lut_2798 ({sk[980], i_30_, i_34_, i_29_, i_37_, n_n1216}, x524x);
	defparam lut_2798.LUT_SIZE = 6;
	defparam lut_2798.mask = 64'h0fff0fff00100000;

	lut_sub lut_2800 ({sk[981], i_17_, n_n1441, x54x, x259x, x348x}, x695x);
	defparam lut_2800.LUT_SIZE = 6;
	defparam lut_2800.mask = 64'h0fff0fff00570055;

	lut_sub lut_2803 ({sk[982], n_n1141, n_n1263, x8x, x216x, x524x}, x7111x);
	defparam lut_2803.LUT_SIZE = 6;
	defparam lut_2803.mask = 64'h0fff0fff03030357;

	lut_sub lut_2806 ({sk[983], i_20_, i_16_, n_n1391, x275x, x399x}, x1588x);
	defparam lut_2806.LUT_SIZE = 6;
	defparam lut_2806.mask = 64'h0fff0fff11111311;

	lut_sub lut_2809 ({sk[984], i_14_, i_12_, i_17_, i_16_, x247x}, x1589x);
	defparam lut_2809.LUT_SIZE = 6;
	defparam lut_2809.mask = 64'h0fff0fff44400000;

	lut_sub lut_2812 ({sk[985], n_n504, x57x, x695x, x1588x, x1589x}, x7112x);
	defparam lut_2812.LUT_SIZE = 6;
	defparam lut_2812.mask = 64'h0fff0fff7777777f;

	lut_sub lut_2816 ({sk[986], i_32_, n_n1306, x222x, n_n245}, x358x);
	defparam lut_2816.LUT_SIZE = 5;
	defparam lut_2816.mask = 32'h55570100;

	lut_sub lut_2818 ({sk[987], i_13_, i_12_, i_16_, i_33_, i_37_}, x470x);
	defparam lut_2818.LUT_SIZE = 6;
	defparam lut_2818.mask = 64'h0fff0fff40000000;

	lut_sub lut_2820 ({sk[988], i_13_, i_17_, i_16_, n_n1307, n_n853}, x367x);
	defparam lut_2820.LUT_SIZE = 6;
	defparam lut_2820.mask = 64'h0fff0fff10000000;

	lut_sub lut_2822 ({sk[989], i_10_, x43x, n_n1307, n_n841, x48x}, x1544x);
	defparam lut_2822.LUT_SIZE = 6;
	defparam lut_2822.mask = 64'h0fff0fff00010000;

	lut_sub lut_2824 ({sk[990], n_n1288, n_n1018, n_n1437, x367x, x1544x}, x1543x);
	defparam lut_2824.LUT_SIZE = 6;
	defparam lut_2824.mask = 64'h0fff0fff05050507;

	lut_sub lut_2827 ({sk[991], i_10_, i_13_, i_16_, x48x}, x384x);
	defparam lut_2827.LUT_SIZE = 5;
	defparam lut_2827.mask = 32'h55574000;

	lut_sub lut_2829 ({sk[992], i_34_, i_35_, n_n793, n_n1305, n_n458}, x1540x);
	defparam lut_2829.LUT_SIZE = 6;
	defparam lut_2829.mask = 64'h0fff0fff00010000;

	lut_sub lut_2831 ({sk[993], i_28_, i_33_, i_29_, n_n242, x318x}, x1542x);
	defparam lut_2831.LUT_SIZE = 6;
	defparam lut_2831.mask = 64'h0fff0fff10000000;

	lut_sub lut_2833 ({sk[994], n_n1340, x14x, x384x, x1540x, x1542x}, x7170x);
	defparam lut_2833.LUT_SIZE = 6;
	defparam lut_2833.mask = 64'h0fff0fff7777777f;

	lut_sub lut_2837 ({sk[995], i_8_, i_6_, i_12_, x43x, x222x}, x1538x);
	defparam lut_2837.LUT_SIZE = 6;
	defparam lut_2837.mask = 64'h0fff0fff10000000;

	lut_sub lut_2839 ({sk[996], i_6_, i_13_, i_12_, i_16_, x63x}, x1539x);
	defparam lut_2839.LUT_SIZE = 6;
	defparam lut_2839.mask = 64'h0fff0fff40000000;

	lut_sub lut_2841 ({sk[997], i_7_, i_8_, i_6_, x88x, x470x}, x1537x);
	defparam lut_2841.LUT_SIZE = 6;
	defparam lut_2841.mask = 64'h0fff0fff10000000;

	lut_sub lut_2843 ({sk[998], n_n504, n_n245, x1538x, x1539x, x1535x}, x7171x);
	defparam lut_2843.LUT_SIZE = 6;
	defparam lut_2843.mask = 64'h0fff0fff5555557f;

	lut_sub lut_2847 ({sk[999], i_37_, x1543x, x7170x, x1537x, x7171x}, n_n1703);
	defparam lut_2847.LUT_SIZE = 6;
	defparam lut_2847.mask = 64'h0fff0fff77777fff;

	lut_sub lut_2852 ({sk[1000], i_2_, n_n1369, n_n1345, n_n576, n_n1282}, x295x);
	defparam lut_2852.LUT_SIZE = 6;
	defparam lut_2852.mask = 64'h0fff0fff00010000;

	lut_sub lut_2854 ({sk[1001], i_2_, i_21_, x263x, x265x, x202x}, x352x);
	defparam lut_2854.LUT_SIZE = 6;
	defparam lut_2854.mask = 64'h0fff0fff01000000;

	lut_sub lut_2856 ({sk[1002], i_34_, n_n1307, n_n1100, x9x, x344x}, x286x);
	defparam lut_2856.LUT_SIZE = 6;
	defparam lut_2856.mask = 64'h0fff0fff00000001;

	lut_sub lut_2858 ({sk[1003], n_n1466, x266x, n_n1202, x250x, n_n1086}, x1211x);
	defparam lut_2858.LUT_SIZE = 6;
	defparam lut_2858.mask = 64'h0fff0fff00000357;

	lut_sub lut_2861 ({sk[1004], i_13_, x286x, x1206x, x1207x}, x7527x);
	defparam lut_2861.LUT_SIZE = 5;
	defparam lut_2861.mask = 32'h5557777f;

	lut_sub lut_2865 ({sk[1005], n_n928, x53x, x7520x, x1209x, x7522x}, x7528x);
	defparam lut_2865.LUT_SIZE = 6;
	defparam lut_2865.mask = 64'h0fff0fff33773f7f;

	lut_sub lut_2869 ({sk[1006], x1211x, x7527x, x7528x}, n_n1872);
	defparam lut_2869.LUT_SIZE = 4;
	defparam lut_2869.mask = 16'h577f;

	lut_sub lut_2873 ({sk[1007], i_30_, i_32_, i_31_, n_n1375, n_n1213}, x306x);
	defparam lut_2873.LUT_SIZE = 6;
	defparam lut_2873.mask = 64'h0fff0fff01000000;

	lut_sub lut_2875 ({sk[1008], i_30_, i_28_, i_29_}, x6984x);
	defparam lut_2875.LUT_SIZE = 4;
	defparam lut_2875.mask = 16'h5740;

	lut_sub lut_2877 ({sk[1009], i_14_, i_13_, n_n1322, x15x, x80x}, x1532x);
	defparam lut_2877.LUT_SIZE = 6;
	defparam lut_2877.mask = 64'h0fff0fff00010000;

	lut_sub lut_2879 ({sk[1010], i_10_, i_32_, x10x, x14x, x48x}, x9234x);
	defparam lut_2879.LUT_SIZE = 6;
	defparam lut_2879.mask = 64'h0fff0ffffeffffff;

	lut_sub lut_2891 ({sk[1011], x260x, x223x, x80x, x147x, x9234x}, x7182x);
	defparam lut_2891.LUT_SIZE = 6;
	defparam lut_2891.mask = 64'h0fff0fffbbbbbbbf;

	lut_sub lut_2895 ({sk[1012], i_32_, i_29_, n_n793, n_n358}, x1528x);
	defparam lut_2895.LUT_SIZE = 5;
	defparam lut_2895.mask = 32'h55571000;

	lut_sub lut_2897 ({sk[1013], i_27_, i_28_, i_29_, x242x, n_n355}, x1529x);
	defparam lut_2897.LUT_SIZE = 6;
	defparam lut_2897.mask = 64'h0fff0fff10000000;

	lut_sub lut_2899 ({sk[1014], i_14_, i_12_, i_16_, n_n1303, x88x}, x1527x);
	defparam lut_2899.LUT_SIZE = 6;
	defparam lut_2899.mask = 64'h0fff0fff10000000;

	lut_sub lut_2901 ({sk[1015], i_37_, n_n1458, x67x, x1527x, x367x}, x1524x);
	defparam lut_2901.LUT_SIZE = 6;
	defparam lut_2901.mask = 64'h0fff0fff00003337;

	lut_sub lut_2904 ({sk[1016], x217x, x1528x, x1529x, x7175x, x7176x}, x7183x);
	defparam lut_2904.LUT_SIZE = 6;
	defparam lut_2904.mask = 64'h0fff0fff03335777;

	lut_sub lut_2908 ({sk[1017], n_n1295, x1532x, x7182x, x1524x, x7183x}, n_n1704);
	defparam lut_2908.LUT_SIZE = 6;
	defparam lut_2908.mask = 64'h0fff0fff77777fff;

	lut_sub lut_2913 ({sk[1018], i_28_, i_32_, i_29_, n_n1018, n_n458}, x1515x);
	defparam lut_2913.LUT_SIZE = 6;
	defparam lut_2913.mask = 64'h0fff0fff10000000;

	lut_sub lut_2915 ({sk[1019], i_8_, i_6_, i_12_, x10x, x222x}, x1513x);
	defparam lut_2915.LUT_SIZE = 6;
	defparam lut_2915.mask = 64'h0fff0fff10000000;

	lut_sub lut_2917 ({sk[1020], i_6_, i_14_, i_12_, i_16_, x63x}, x1514x);
	defparam lut_2917.LUT_SIZE = 6;
	defparam lut_2917.mask = 64'h0fff0fff40000000;

	lut_sub lut_2919 ({sk[1021], i_5_, i_4_, i_0_, i_35_, i_37_}, x7187x);
	defparam lut_2919.LUT_SIZE = 6;
	defparam lut_2919.mask = 64'h0fff0fff40000000;

	lut_sub lut_2921 ({sk[1022], x268x, x358x, x1513x, x1514x, x7187x}, x7192x);
	defparam lut_2921.LUT_SIZE = 6;
	defparam lut_2921.mask = 64'h0fff0fff151515ff;

	lut_sub lut_2925 ({sk[1023], i_33_, n_n1295, x48x, n_n242, x1515x}, x1510x);
	defparam lut_2925.LUT_SIZE = 6;
	defparam lut_2925.mask = 64'h0fff0fff00570000;

	lut_sub lut_2928 ({sk[1024], x144x, x248x, x221x, x710x, x1517x}, x1511x);
	defparam lut_2928.LUT_SIZE = 6;
	defparam lut_2928.mask = 64'h0fff0fff005700ff;

	lut_sub lut_2932 ({sk[1025], x7192x, x1510x, x1511x}, n_n1705);
	defparam lut_2932.LUT_SIZE = 4;
	defparam lut_2932.mask = 16'h577f;

	lut_sub lut_2936 ({sk[1026], i_9_, i_10_, i_24_, x11x}, x327x);
	defparam lut_2936.LUT_SIZE = 5;
	defparam lut_2936.mask = 32'h55570040;

	lut_sub lut_2938 ({sk[1027], i_9_, i_10_, i_5_, i_6_, n_n1279}, x335x);
	defparam lut_2938.LUT_SIZE = 6;
	defparam lut_2938.mask = 64'h0fff0fff00004000;

	lut_sub lut_2940 ({sk[1028], i_8_, i_28_, i_24_, i_29_, x297x}, x1398x);
	defparam lut_2940.LUT_SIZE = 6;
	defparam lut_2940.mask = 64'h0fff0fff40000000;

	lut_sub lut_2942 ({sk[1029], i_7_, i_11_, i_19_, n_n1307, x280x}, x1406x);
	defparam lut_2942.LUT_SIZE = 6;
	defparam lut_2942.mask = 64'h0fff0fff10000000;

	lut_sub lut_2944 ({sk[1030], i_9_, i_18_, x242x, n_n787, n_n1118}, x1507x);
	defparam lut_2944.LUT_SIZE = 6;
	defparam lut_2944.mask = 64'h0fff0fff01000000;

	lut_sub lut_2946 ({sk[1031], i_11_, i_19_, x242x, x41x, x1507x}, x27x);
	defparam lut_2946.LUT_SIZE = 6;
	defparam lut_2946.mask = 64'h0fff0fff57555555;

	lut_sub lut_2949 ({sk[1032], i_14_, i_13_, i_16_, x318x, x272x}, x1506x);
	defparam lut_2949.LUT_SIZE = 6;
	defparam lut_2949.mask = 64'h0fff0fff00100000;

	lut_sub lut_2951 ({sk[1033], i_8_, x10x, n_n1278, n_n152, x319x}, x1504x);
	defparam lut_2951.LUT_SIZE = 6;
	defparam lut_2951.mask = 64'h0fff0fff00010000;

	lut_sub lut_2953 ({sk[1034], i_14_, i_34_, i_35_, n_n1375, n_n1322}, x7204x);
	defparam lut_2953.LUT_SIZE = 6;
	defparam lut_2953.mask = 64'h0fff0fff01000000;

	lut_sub lut_2955 ({sk[1035], i_37_, x223x, x1506x, x1504x, x7204x}, x1501x);
	defparam lut_2955.LUT_SIZE = 6;
	defparam lut_2955.mask = 64'h0fff0fff00003f7f;

	lut_sub lut_2959 ({sk[1036], n_n1408, n_n1422, x365x, x7x, x9232x}, x1500x);
	defparam lut_2959.LUT_SIZE = 6;
	defparam lut_2959.mask = 64'h0fff0fff0a0a0a0b;

	lut_sub lut_2962 ({sk[1037], x60x, x27x, x7195x, x7199x}, x7206x);
	defparam lut_2962.LUT_SIZE = 5;
	defparam lut_2962.mask = 32'h55570537;

	lut_sub lut_2965 ({sk[1038], x1501x, x1500x, x7206x}, n_n1701);
	defparam lut_2965.LUT_SIZE = 4;
	defparam lut_2965.mask = 16'h577f;

	lut_sub lut_2969 ({sk[1039], i_5_, i_6_, n_n152, x46x, n_n629}, x386x);
	defparam lut_2969.LUT_SIZE = 6;
	defparam lut_2969.mask = 64'h0fff0fff01000000;

	lut_sub lut_2971 ({sk[1040], i_7_, i_5_, i_6_, i_32_, i_37_}, x1496x);
	defparam lut_2971.LUT_SIZE = 6;
	defparam lut_2971.mask = 64'h0fff0fff40000000;

	lut_sub lut_2973 ({sk[1041], n_n1318, n_n1118, n_n152, x274x, x1496x}, x1494x);
	defparam lut_2973.LUT_SIZE = 6;
	defparam lut_2973.mask = 64'h0fff0fff01010103;

	lut_sub lut_2976 ({sk[1042], i_16_, i_37_, x242x, n_n1216, n_n1241}, x7210x);
	defparam lut_2976.LUT_SIZE = 6;
	defparam lut_2976.mask = 64'h0fff0fff00010000;

	lut_sub lut_2978 ({sk[1043], i_10_, n_n82, x268x, x87x, x7210x}, x7221x);
	defparam lut_2978.LUT_SIZE = 6;
	defparam lut_2978.mask = 64'h0fff0fff03570055;

	lut_sub lut_2981 ({sk[1044], n_n1408, x243x, x366x, x7x, x1494x}, x1493x);
	defparam lut_2981.LUT_SIZE = 6;
	defparam lut_2981.mask = 64'h0fff0fff00005557;

	lut_sub lut_2984 ({sk[1045], i_32_, x416x, x27x, x386x, x7212x}, x7220x);
	defparam lut_2984.LUT_SIZE = 6;
	defparam lut_2984.mask = 64'h0fff0fff05370505;

	lut_sub lut_2987 ({sk[1046], x7221x, x1493x, x7220x}, n_n1702);
	defparam lut_2987.LUT_SIZE = 4;
	defparam lut_2987.mask = 16'h577f;

	lut_sub lut_2991 ({sk[1047], i_10_, i_7_, i_3_, i_18_, x54x}, x382x);
	defparam lut_2991.LUT_SIZE = 6;
	defparam lut_2991.mask = 64'h0fff0fff00000004;

	lut_sub lut_2993 ({sk[1048], i_9_, i_8_, i_2_, n_n735, x343x}, x7344x);
	defparam lut_2993.LUT_SIZE = 6;
	defparam lut_2993.mask = 64'h0fff0fff50007000;

	lut_sub lut_2996 ({sk[1049], i_7_, i_14_, i_12_, i_17_, i_16_}, x94x);
	defparam lut_2996.LUT_SIZE = 6;
	defparam lut_2996.mask = 64'h0fff0fff0000a800;

	lut_sub lut_2999 ({sk[1050], i_27_, x42x, x48x, x259x, x348x}, x729x);
	defparam lut_2999.LUT_SIZE = 6;
	defparam lut_2999.mask = 64'h0fff0fff03570303;

	lut_sub lut_3002 ({sk[1051], i_12_, i_17_, x10x, x331x, x1579x}, x7116x);
	defparam lut_3002.LUT_SIZE = 6;
	defparam lut_3002.mask = 64'h0fff0fff57575755;

	lut_sub lut_3006 ({sk[1052], x59x, n_n1443, x322x, x306x, x7116x}, x7118x);
	defparam lut_3006.LUT_SIZE = 6;
	defparam lut_3006.mask = 64'h0fff0fff555f557f;

	lut_sub lut_3010 ({sk[1053], i_30_, i_34_, i_33_, i_35_, i_37_}, x7114x);
	defparam lut_3010.LUT_SIZE = 6;
	defparam lut_3010.mask = 64'h0fff0fff00400000;

	lut_sub lut_3012 ({sk[1054], n_n1429, x322x, x729x, x7118x, x7114x}, n_n1713);
	defparam lut_3012.LUT_SIZE = 6;
	defparam lut_3012.mask = 64'h0fff0fff373737ff;

	lut_sub lut_3016 ({sk[1055], i_23_, i_16_, n_n1397, n_n1384, x7058x}, x151x);
	defparam lut_3016.LUT_SIZE = 6;
	defparam lut_3016.mask = 64'h0fff0fff01000000;

	lut_sub lut_3018 ({sk[1056], i_16_, i_31_, n_n793, n_n1397, n_n1285}, x153x);
	defparam lut_3018.LUT_SIZE = 6;
	defparam lut_3018.mask = 64'h0fff0fff00010000;

	lut_sub lut_3020 ({sk[1057], i_30_, i_7_, i_8_, i_28_, i_29_}, x369x);
	defparam lut_3020.LUT_SIZE = 6;
	defparam lut_3020.mask = 64'h0fff0fff80000000;

	lut_sub lut_3022 ({sk[1058], i_30_, i_28_, i_22_, i_32_, x285x}, x1028x);
	defparam lut_3022.LUT_SIZE = 6;
	defparam lut_3022.mask = 64'h0fff0fff01000500;

	lut_sub lut_3025 ({sk[1059], i_25_, i_34_, i_33_, i_35_, i_38_}, x733x);
	defparam lut_3025.LUT_SIZE = 6;
	defparam lut_3025.mask = 64'h0fff0fff11001000;

	lut_sub lut_3028 ({sk[1060], n_n1489, x13x, x238x, x284x, x733x}, x7688x);
	defparam lut_3028.LUT_SIZE = 6;
	defparam lut_3028.mask = 64'h0fff0fff00000357;

	lut_sub lut_3031 ({sk[1061], i_28_, i_24_, i_33_, i_29_}, x7547x);
	defparam lut_3031.LUT_SIZE = 5;
	defparam lut_3031.mask = 32'h55578000;

	lut_sub lut_3033 ({sk[1062], i_31_, i_34_, i_35_, i_38_, x7547x}, x66x);
	defparam lut_3033.LUT_SIZE = 6;
	defparam lut_3033.mask = 64'h0fff0fff00100000;

	lut_sub lut_3035 ({sk[1063], i_28_, i_31_, i_29_, n_n1340, x12x}, x502x);
	defparam lut_3035.LUT_SIZE = 6;
	defparam lut_3035.mask = 64'h0fff0fff10000000;

	lut_sub lut_3037 ({sk[1064], i_9_, i_8_, i_3_, i_11_, i_18_}, x17x);
	defparam lut_3037.LUT_SIZE = 6;
	defparam lut_3037.mask = 64'h0fff0fff00003100;

	lut_sub lut_3040 ({sk[1065], i_13_, i_19_, n_n1038, x17x}, x1197x);
	defparam lut_3040.LUT_SIZE = 5;
	defparam lut_3040.mask = 32'h55575700;

	lut_sub lut_3043 ({sk[1066], i_18_, i_19_, n_n1028, x1197x}, x736x);
	defparam lut_3043.LUT_SIZE = 5;
	defparam lut_3043.mask = 32'h55575557;

	lut_sub lut_3046 ({sk[1067], i_28_, i_25_, i_26_, i_38_, i_29_}, x7544x);
	defparam lut_3046.LUT_SIZE = 6;
	defparam lut_3046.mask = 64'h0fff0fff20000000;

	lut_sub lut_3048 ({sk[1068], i_22_, i_32_, x11x, n_n1497, x226x}, x1192x);
	defparam lut_3048.LUT_SIZE = 6;
	defparam lut_3048.mask = 64'h0fff0fff01000000;

	lut_sub lut_3050 ({sk[1069], x51x, n_n928, x502x, x7544x, x1192x}, x7550x);
	defparam lut_3050.LUT_SIZE = 6;
	defparam lut_3050.mask = 64'h0fff0fff55775f7f;

	lut_sub lut_3054 ({sk[1070], i_33_, i_35_, i_38_, n_n1486, x278x}, x7543x);
	defparam lut_3054.LUT_SIZE = 6;
	defparam lut_3054.mask = 64'h0fff0fff01000000;

	lut_sub lut_3056 ({sk[1071], i_8_, i_5_, i_6_, n_n1279, x66x}, x1195x);
	defparam lut_3056.LUT_SIZE = 6;
	defparam lut_3056.mask = 64'h0fff0fff10000000;

	lut_sub lut_3058 ({sk[1072], x53x, x360x, x736x, x7543x, x1195x}, x7551x);
	defparam lut_3058.LUT_SIZE = 6;
	defparam lut_3058.mask = 64'h0fff0fff575757ff;

	lut_sub lut_3062 ({sk[1073], i_31_, i_29_, n_n1118, n_n1279, x315x}, x1200x);
	defparam lut_3062.LUT_SIZE = 6;
	defparam lut_3062.mask = 64'h0fff0fff01000000;

	lut_sub lut_3064 ({sk[1074], i_8_, x42x, n_n1278, n_n1279, n_n1059}, x1201x);
	defparam lut_3064.LUT_SIZE = 6;
	defparam lut_3064.mask = 64'h0fff0fff00010000;

	lut_sub lut_3066 ({sk[1075], i_30_, i_24_, i_29_, n_n1361, n_n1478}, x7534x);
	defparam lut_3066.LUT_SIZE = 6;
	defparam lut_3066.mask = 64'h0fff0fff10000000;

	lut_sub lut_3068 ({sk[1076], x425x, x454x, x1200x, x1201x, x7534x}, x7539x);
	defparam lut_3068.LUT_SIZE = 6;
	defparam lut_3068.mask = 64'h0fff0fff3f7f7f7f;

	lut_sub lut_3073 ({sk[1077], i_28_, i_34_, i_33_, i_38_, i_29_}, x7535x);
	defparam lut_3073.LUT_SIZE = 6;
	defparam lut_3073.mask = 64'h0fff0fff00200000;

	lut_sub lut_3075 ({sk[1078], i_31_, i_35_, i_38_, x76x, x257x}, x1204x);
	defparam lut_3075.LUT_SIZE = 6;
	defparam lut_3075.mask = 64'h0fff0fff01000000;

	lut_sub lut_3077 ({sk[1079], i_10_, n_n1086, x286x, x7535x, x1204x}, x7540x);
	defparam lut_3077.LUT_SIZE = 6;
	defparam lut_3077.mask = 64'h0fff0fff5f7f5577;

	lut_sub lut_3081 ({sk[1080], i_29_, x360x, x311x, x315x, n_n1086}, x1184x);
	defparam lut_3081.LUT_SIZE = 6;
	defparam lut_3081.mask = 64'h0fff0fff05370000;

	lut_sub lut_3084 ({sk[1081], i_32_, x42x, x321x, x72x, n_n1059}, x1183x);
	defparam lut_3084.LUT_SIZE = 6;
	defparam lut_3084.mask = 64'h0fff0fff00150011;

	lut_sub lut_3087 ({sk[1082], n_n1489, x395x, x294x, x346x, x744x}, x7553x);
	defparam lut_3087.LUT_SIZE = 6;
	defparam lut_3087.mask = 64'h0fff0fff00330537;

	lut_sub lut_3090 ({sk[1083], x1184x, x1183x, x7553x}, n_n1876);
	defparam lut_3090.LUT_SIZE = 4;
	defparam lut_3090.mask = 16'h577f;

	lut_sub lut_3094 ({sk[1084], x1171x, x1173x, x1174x, x1175x}, x7568x);
	defparam lut_3094.LUT_SIZE = 5;
	defparam lut_3094.mask = 32'h55577fff;

	lut_sub lut_3099 ({sk[1085], x51x, x465x, x751x, x7559x, x1176x}, x7569x);
	defparam lut_3099.LUT_SIZE = 6;
	defparam lut_3099.mask = 64'h0fff0fff575757ff;

	lut_sub lut_3103 ({sk[1086], x395x, x1152x, x1153x, x7585x, x1155x}, x7590x);
	defparam lut_3103.LUT_SIZE = 6;
	defparam lut_3103.mask = 64'h0fff0fff5fff7fff;

	lut_sub lut_3108 ({sk[1087], x11x, x76x, x66x, x502x, x465x}, x7589x);
	defparam lut_3108.LUT_SIZE = 6;
	defparam lut_3108.mask = 64'h0fff0fff000f777f;

	lut_sub lut_3112 ({sk[1088], n_n928, x380x, n_n1086, x7590x, x7589x}, n_n1877);
	defparam lut_3112.LUT_SIZE = 6;
	defparam lut_3112.mask = 64'h0fff0fff777f77ff;

	lut_sub lut_3117 ({sk[1089], i_10_, x56x, x284x, x1166x, x9214x}, x777x);
	defparam lut_3117.LUT_SIZE = 6;
	defparam lut_3117.mask = 64'h0fff0fffbbbf333f;

	lut_sub lut_3121 ({sk[1090], x51x, x776x, x1159x, x1160x, x1161x}, x7581x);
	defparam lut_3121.LUT_SIZE = 6;
	defparam lut_3121.mask = 64'h0fff0fff7f7f7fff;

	lut_sub lut_3126 ({sk[1091], x76x, x62x, x8x, x781x, x1142x}, x7593x);
	defparam lut_3126.LUT_SIZE = 6;
	defparam lut_3126.mask = 64'h0fff0fff555f777f;

	lut_sub lut_3130 ({sk[1092], i_9_, i_12_, x11x, x783x, x782x}, x7594x);
	defparam lut_3130.LUT_SIZE = 6;
	defparam lut_3130.mask = 64'h0fff0fff03030357;

	lut_sub lut_3133 ({sk[1093], x68x, x777x, x7581x, x7593x, x7594x}, x7596x);
	defparam lut_3133.LUT_SIZE = 6;
	defparam lut_3133.mask = 64'h0fff0fff7f7f7fff;

	lut_sub lut_3138 ({sk[1094], x7513x, x7514x, x7539x, x7540x}, x7597x);
	defparam lut_3138.LUT_SIZE = 5;
	defparam lut_3138.mask = 32'h55577fff;

	lut_sub lut_3143 ({sk[1095], i_20_, i_24_, i_21_, i_22_, i_34_}, x1078x);
	defparam lut_3143.LUT_SIZE = 6;
	defparam lut_3143.mask = 64'h0fff0fff04004400;

	lut_sub lut_3146 ({sk[1096], i_24_, i_31_, x3x, x240x, x285x}, x738x);
	defparam lut_3146.LUT_SIZE = 6;
	defparam lut_3146.mask = 64'h0fff0fff05770000;

	lut_sub lut_3150 ({sk[1097], n_n1397, x83x, x95x, x96x, x7620x}, x7621x);
	defparam lut_3150.LUT_SIZE = 6;
	defparam lut_3150.mask = 64'h0fff0fff5555557f;

	lut_sub lut_3154 ({sk[1098], x1087x, x7635x, n_n1897, x1070x, x1071x}, x7642x);
	defparam lut_3154.LUT_SIZE = 6;
	defparam lut_3154.mask = 64'h0fff0fff7fffffff;

	lut_sub lut_3160 ({sk[1099], i_7_, i_5_, i_6_, n_n1279, x70x}, x1069x);
	defparam lut_3160.LUT_SIZE = 6;
	defparam lut_3160.mask = 64'h0fff0fff10000000;

	lut_sub lut_3162 ({sk[1100], i_32_, x257x, x250x, x206x, x1069x}, x1064x);
	defparam lut_3162.LUT_SIZE = 6;
	defparam lut_3162.mask = 64'h0fff0fff557f0000;

	lut_sub lut_3166 ({sk[1101], n_n1191, n_n1192, x787x, x1063x}, x7650x);
	defparam lut_3166.LUT_SIZE = 5;
	defparam lut_3166.mask = 32'h55575557;

	lut_sub lut_3169 ({sk[1102], x72x, x9x, x78x, x1060x, x1062x}, x7651x);
	defparam lut_3169.LUT_SIZE = 6;
	defparam lut_3169.mask = 64'h0fff0fff7777777f;

	lut_sub lut_3173 ({sk[1103], x1064x, x7650x, x7651x}, n_n1880);
	defparam lut_3173.LUT_SIZE = 4;
	defparam lut_3173.mask = 16'h577f;

	lut_sub lut_3177 ({sk[1104], i_7_, i_8_, n_n1300, x282x, x466x}, x1046x);
	defparam lut_3177.LUT_SIZE = 6;
	defparam lut_3177.mask = 64'h0fff0fff07030303;

	lut_sub lut_3180 ({sk[1105], n_n1305, x250x, n_n1497, x206x, x1045x}, x7667x);
	defparam lut_3180.LUT_SIZE = 6;
	defparam lut_3180.mask = 64'h0fff0fff5555575f;

	lut_sub lut_3184 ({sk[1106], x72x, x9x, x430x, x1041x, x1042x}, x7668x);
	defparam lut_3184.LUT_SIZE = 6;
	defparam lut_3184.mask = 64'h0fff0fff7777777f;

	lut_sub lut_3188 ({sk[1107], x249x, x68x, x1046x, x7667x, x7668x}, n_n1883);
	defparam lut_3188.LUT_SIZE = 6;
	defparam lut_3188.mask = 64'h0fff0fff777f77ff;

	lut_sub lut_3193 ({sk[1108], n_n1404, n_n1408, x55x, x1050x, x1051x}, x7661x);
	defparam lut_3193.LUT_SIZE = 6;
	defparam lut_3193.mask = 64'h0fff0fff777f7f7f;

	lut_sub lut_3198 ({sk[1109], n_n1353, n_n1359, x1059x, x7659x, x746x}, x7662x);
	defparam lut_3198.LUT_SIZE = 6;
	defparam lut_3198.mask = 64'h0fff0fff003f557f;

	lut_sub lut_3202 ({sk[1110], n_n1443, n_n1429, x128x, x55x, x1030x}, x7678x);
	defparam lut_3202.LUT_SIZE = 6;
	defparam lut_3202.mask = 64'h0fff0fff5f7f7f7f;

	lut_sub lut_3207 ({sk[1111], x145x, x1029x, x1031x, x1032x}, x7679x);
	defparam lut_3207.LUT_SIZE = 5;
	defparam lut_3207.mask = 32'h55577fff;

	lut_sub lut_3212 ({sk[1112], x7661x, x7662x, x7678x, x7679x}, x7681x);
	defparam lut_3212.LUT_SIZE = 5;
	defparam lut_3212.mask = 32'h55577fff;

	lut_sub lut_3217 ({sk[1113], i_2_, i_38_, x795x, x1017x, x1018x}, x1013x);
	defparam lut_3217.LUT_SIZE = 6;
	defparam lut_3217.mask = 64'h0fff0fff007f0077;

	lut_sub lut_3221 ({sk[1114], i_2_, x70x, x77x, x1010x, x7698x}, x7699x);
	defparam lut_3221.LUT_SIZE = 6;
	defparam lut_3221.mask = 64'h0fff0fff777f7777;

	lut_sub lut_3225 ({sk[1115], n_n1489, x214x, x797x, x796x, x1000x}, x7707x);
	defparam lut_3225.LUT_SIZE = 6;
	defparam lut_3225.mask = 64'h0fff0fff555f777f;

	lut_sub lut_3229 ({sk[1116], x7688x, x999x, x1001x, x1025x, x7687x}, x7708x);
	defparam lut_3229.LUT_SIZE = 6;
	defparam lut_3229.mask = 64'h0fff0fff7fffffff;

	lut_sub lut_3235 ({sk[1117], x1484x, x1485x, x7231x, x7232x}, x7235x);
	defparam lut_3235.LUT_SIZE = 5;
	defparam lut_3235.mask = 32'h55577fff;

	lut_sub lut_3240 ({sk[1118], i_13_, i_19_, n_n1058, x18x, x436x}, x744x);
	defparam lut_3240.LUT_SIZE = 6;
	defparam lut_3240.mask = 64'h0fff0fff5f7f5577;

	lut_sub lut_3244 ({sk[1119], i_18_, i_24_, x204x, x60x, x14x}, x26x);
	defparam lut_3244.LUT_SIZE = 6;
	defparam lut_3244.mask = 64'h0fff0fff37000500;

	lut_sub lut_3247 ({sk[1120], i_30_, i_32_, i_34_, n_n1361, n_n1466}, x1059x);
	defparam lut_3247.LUT_SIZE = 6;
	defparam lut_3247.mask = 64'h0fff0fff01000000;

	lut_sub lut_3249 ({sk[1121], n_n1489, n_n1361, n_n1478, n_n1340, n_n1472}, x7659x);
	defparam lut_3249.LUT_SIZE = 6;
	defparam lut_3249.mask = 64'h0fff0fff00050037;

	lut_sub lut_3252 ({sk[1122], i_30_, x42x, n_n805, x81x, x7547x}, x746x);
	defparam lut_3252.LUT_SIZE = 6;
	defparam lut_3252.mask = 64'h0fff0fff05370000;

	lut_sub lut_3255 ({sk[1123], i_8_, i_2_, i_22_, n_n1345, x81x}, x1050x);
	defparam lut_3255.LUT_SIZE = 6;
	defparam lut_3255.mask = 64'h0fff0fff10000000;

	lut_sub lut_3257 ({sk[1124], i_30_, i_2_, i_32_, i_31_, x276x}, x1051x);
	defparam lut_3257.LUT_SIZE = 6;
	defparam lut_3257.mask = 64'h0fff0fff40000000;

	lut_sub lut_3259 ({sk[1125], i_28_, i_25_, i_32_, i_29_, x327x}, x994x);
	defparam lut_3259.LUT_SIZE = 6;
	defparam lut_3259.mask = 64'h0fff0fff40000000;

	lut_sub lut_3261 ({sk[1126], i_28_, i_25_, i_29_, n_n1433, x12x}, x465x);
	defparam lut_3261.LUT_SIZE = 6;
	defparam lut_3261.mask = 64'h0fff0fff10000000;

	lut_sub lut_3263 ({sk[1127], i_28_, i_25_, i_26_, i_24_, i_29_}, x7557x);
	defparam lut_3263.LUT_SIZE = 6;
	defparam lut_3263.mask = 64'h0fff0fff80000000;

	lut_sub lut_3265 ({sk[1128], n_n1486, n_n998, x18x, x436x, x7557x}, x751x);
	defparam lut_3265.LUT_SIZE = 6;
	defparam lut_3265.mask = 64'h0fff0fff1111111f;

	lut_sub lut_3268 ({sk[1129], i_13_, i_12_, i_17_, i_16_, x216x}, x1480x);
	defparam lut_3268.LUT_SIZE = 6;
	defparam lut_3268.mask = 64'h0fff0fff44400000;

	lut_sub lut_3271 ({sk[1130], i_30_, i_12_, x13x, n_n1263, x260x}, x756x);
	defparam lut_3271.LUT_SIZE = 6;
	defparam lut_3271.mask = 64'h0fff0fff07050000;

	lut_sub lut_3274 ({sk[1131], i_33_, x323x, x291x, x524x, x1480x}, x1474x);
	defparam lut_3274.LUT_SIZE = 6;
	defparam lut_3274.mask = 64'h0fff0fff57770000;

	lut_sub lut_3278 ({sk[1132], i_27_, i_34_, i_35_, i_37_, x42x}, x7242x);
	defparam lut_3278.LUT_SIZE = 6;
	defparam lut_3278.mask = 64'h0fff0fff01000000;

	lut_sub lut_3280 ({sk[1133], i_12_, i_33_, i_37_, x43x, x306x}, x1475x);
	defparam lut_3280.LUT_SIZE = 6;
	defparam lut_3280.mask = 64'h0fff0fff01000000;

	lut_sub lut_3282 ({sk[1134], x82x, x29x, x756x, x7242x, x1475x}, x7245x);
	defparam lut_3282.LUT_SIZE = 6;
	defparam lut_3282.mask = 64'h0fff0fff575757ff;

	lut_sub lut_3286 ({sk[1135], i_30_, i_28_, i_26_, i_24_, i_22_}, x466x);
	defparam lut_3286.LUT_SIZE = 6;
	defparam lut_3286.mask = 64'h0fff0fff80000000;

	lut_sub lut_3288 ({sk[1136], i_28_, i_26_, i_24_, i_22_, x343x}, x989x);
	defparam lut_3288.LUT_SIZE = 6;
	defparam lut_3288.mask = 64'h0fff0fff40000000;

	lut_sub lut_3290 ({sk[1137], i_3_, i_13_, i_12_, i_11_, i_19_}, x1262x);
	defparam lut_3290.LUT_SIZE = 6;
	defparam lut_3290.mask = 64'h0fff0fff07000000;

	lut_sub lut_3293 ({sk[1138], i_14_, i_23_, i_16_, x76x}, x515x);
	defparam lut_3293.LUT_SIZE = 5;
	defparam lut_3293.mask = 32'h55574000;

	lut_sub lut_3295 ({sk[1139], i_27_, i_23_, x73x, n_n1431, x202x}, x773x);
	defparam lut_3295.LUT_SIZE = 6;
	defparam lut_3295.mask = 64'h0fff0fff57555555;

	lut_sub lut_3298 ({sk[1140], i_14_, i_16_, n_n1369, n_n1274, n_n1431}, x1623x);
	defparam lut_3298.LUT_SIZE = 6;
	defparam lut_3298.mask = 64'h0fff0fff01000000;

	lut_sub lut_3300 ({sk[1141], i_20_, i_14_, i_17_, i_16_, x202x}, x1625x);
	defparam lut_3300.LUT_SIZE = 6;
	defparam lut_3300.mask = 64'h0fff0fff40000000;

	lut_sub lut_3302 ({sk[1142], i_30_, i_28_, i_22_, i_31_, x270x}, x1166x);
	defparam lut_3302.LUT_SIZE = 6;
	defparam lut_3302.mask = 64'h0fff0fff40000000;

	lut_sub lut_3304 ({sk[1143], i_32_, n_n1361, x389x, n_n1431, x313x}, x9214x);
	defparam lut_3304.LUT_SIZE = 6;
	defparam lut_3304.mask = 64'h0fff0ffffca8fcfc;

	lut_sub lut_3311 ({sk[1144], i_28_, i_26_, i_24_, i_29_}, x7576x);
	defparam lut_3311.LUT_SIZE = 5;
	defparam lut_3311.mask = 32'h55578000;

	lut_sub lut_3313 ({sk[1145], n_n1478, n_n1133, x12x, n_n1149, x7576x}, x776x);
	defparam lut_3313.LUT_SIZE = 6;
	defparam lut_3313.mask = 64'h0fff0fff1111111f;

	lut_sub lut_3316 ({sk[1146], i_12_, i_33_, n_n1353, n_n1361, x466x}, x1159x);
	defparam lut_3316.LUT_SIZE = 6;
	defparam lut_3316.mask = 64'h0fff0fff00000100;

	lut_sub lut_3318 ({sk[1147], i_10_, i_26_, i_24_, n_n1300, x272x}, x1160x);
	defparam lut_3318.LUT_SIZE = 6;
	defparam lut_3318.mask = 64'h0fff0fff10000000;

	lut_sub lut_3320 ({sk[1148], i_29_, n_n1118, n_n1279, n_n1497, x226x}, x1161x);
	defparam lut_3320.LUT_SIZE = 6;
	defparam lut_3320.mask = 64'h0fff0fff00010000;

	lut_sub lut_3322 ({sk[1149], i_30_, i_12_, n_n1353, x12x, x78x}, x1152x);
	defparam lut_3322.LUT_SIZE = 6;
	defparam lut_3322.mask = 64'h0fff0fff00010000;

	lut_sub lut_3324 ({sk[1150], i_13_, i_26_, i_24_, n_n1300, x272x}, x1153x);
	defparam lut_3324.LUT_SIZE = 6;
	defparam lut_3324.mask = 64'h0fff0fff00001000;

	lut_sub lut_3326 ({sk[1151], i_10_, i_7_, i_32_, n_n1307, x280x}, x7585x);
	defparam lut_3326.LUT_SIZE = 6;
	defparam lut_3326.mask = 64'h0fff0fff10000000;

	lut_sub lut_3328 ({sk[1152], i_28_, i_31_, i_29_, x50x, x81x}, x1155x);
	defparam lut_3328.LUT_SIZE = 6;
	defparam lut_3328.mask = 64'h0fff0fff10000000;

	lut_sub lut_3330 ({sk[1153], n_n1478, n_n1133, x12x, n_n1149, x7576x}, x783x);
	defparam lut_3330.LUT_SIZE = 6;
	defparam lut_3330.mask = 64'h0fff0fff1111111f;

	lut_sub lut_3333 ({sk[1154], i_33_, n_n1361, n_n1438, x61x, x235x}, x782x);
	defparam lut_3333.LUT_SIZE = 6;
	defparam lut_3333.mask = 64'h0fff0fff55575555;

	lut_sub lut_3336 ({sk[1155], i_29_, n_n1128, n_n1497, x226x, x81x}, x781x);
	defparam lut_3336.LUT_SIZE = 6;
	defparam lut_3336.mask = 64'h0fff0fff03570055;

	lut_sub lut_3339 ({sk[1156], i_30_, i_33_, n_n1425, n_n1361, n_n1478}, x787x);
	defparam lut_3339.LUT_SIZE = 6;
	defparam lut_3339.mask = 64'h0fff0fff13110300;

	lut_sub lut_3342 ({sk[1157], i_14_, i_28_, i_13_, i_22_}, x345x);
	defparam lut_3342.LUT_SIZE = 5;
	defparam lut_3342.mask = 32'h55570010;

	lut_sub lut_3344 ({sk[1158], i_28_, i_12_, i_17_, i_22_}, x1015x);
	defparam lut_3344.LUT_SIZE = 5;
	defparam lut_3344.mask = 32'h55570100;

	lut_sub lut_3346 ({sk[1159], i_7_, i_8_, n_n1431, x313x, x7695x}, x795x);
	defparam lut_3346.LUT_SIZE = 6;
	defparam lut_3346.mask = 64'h0fff0fff37050505;

	lut_sub lut_3349 ({sk[1160], i_30_, i_31_, i_29_, n_n1423, n_n1422}, x1017x);
	defparam lut_3349.LUT_SIZE = 6;
	defparam lut_3349.mask = 64'h0fff0fff10000000;

	lut_sub lut_3351 ({sk[1161], i_28_, i_24_, i_29_, n_n1438, n_n1437}, x1018x);
	defparam lut_3351.LUT_SIZE = 6;
	defparam lut_3351.mask = 64'h0fff0fff10000000;

	lut_sub lut_3353 ({sk[1162], i_30_, i_8_, i_31_, i_29_, x237x}, x1010x);
	defparam lut_3353.LUT_SIZE = 6;
	defparam lut_3353.mask = 64'h0fff0fff40000000;

	lut_sub lut_3355 ({sk[1163], n_n1504, x474x, n_n1059, x345x, x1015x}, x7698x);
	defparam lut_3355.LUT_SIZE = 6;
	defparam lut_3355.mask = 64'h0fff0fff000f777f;

	lut_sub lut_3359 ({sk[1164], i_30_, i_12_, i_17_, i_32_, x285x}, x797x);
	defparam lut_3359.LUT_SIZE = 6;
	defparam lut_3359.mask = 64'h0fff0fff1113555f;

	lut_sub lut_3364 ({sk[1165], i_8_, i_31_, x73x, x226x, x270x}, x796x);
	defparam lut_3364.LUT_SIZE = 6;
	defparam lut_3364.mask = 64'h0fff0fff57035500;

	lut_sub lut_3367 ({sk[1166], i_9_, i_8_, i_11_, i_2_, i_18_}, x1388x);
	defparam lut_3367.LUT_SIZE = 6;
	defparam lut_3367.mask = 64'h0fff0fff00000400;

	lut_sub lut_3369 ({sk[1167], i_2_, i_19_, n_n1038, x1388x}, x37x);
	defparam lut_3369.LUT_SIZE = 5;
	defparam lut_3369.mask = 32'h55575755;

	lut_sub lut_3372 ({sk[1168], i_32_, i_34_, i_29_}, x7409x);
	defparam lut_3372.LUT_SIZE = 4;
	defparam lut_3372.mask = 16'h5720;

	lut_sub lut_3374 ({sk[1169], i_14_, i_13_, i_12_, i_17_, i_16_}, x805x);
	defparam lut_3374.LUT_SIZE = 6;
	defparam lut_3374.mask = 64'h0fff0fffa8a8a800;

	lut_sub lut_3379 ({sk[1170], i_10_, i_7_, i_8_, i_24_, i_22_}, x281x);
	defparam lut_3379.LUT_SIZE = 6;
	defparam lut_3379.mask = 64'h0fff0fff00008000;

	lut_sub lut_3381 ({sk[1171], i_27_, i_28_, i_32_, i_29_, x54x}, x221x);
	defparam lut_3381.LUT_SIZE = 6;
	defparam lut_3381.mask = 64'h0fff0fff40000000;

	lut_sub lut_3383 ({sk[1172], i_20_, i_13_, i_12_, i_16_}, x402x);
	defparam lut_3383.LUT_SIZE = 5;
	defparam lut_3383.mask = 32'h55578000;

	lut_sub lut_3385 ({sk[1173], i_9_, i_8_, i_12_, n_n735}, x414x);
	defparam lut_3385.LUT_SIZE = 5;
	defparam lut_3385.mask = 32'h55570010;

	lut_sub lut_3387 ({sk[1174], i_14_, i_17_, i_16_, n_n1307, n_n839}, x495x);
	defparam lut_3387.LUT_SIZE = 6;
	defparam lut_3387.mask = 64'h0fff0fff10000000;

	lut_sub lut_3389 ({sk[1175], i_7_, i_8_, i_19_, x232x, n_n178}, x105x);
	defparam lut_3389.LUT_SIZE = 6;
	defparam lut_3389.mask = 64'h0fff0fff10000000;

	lut_sub lut_3391 ({sk[1176], i_9_, i_13_, i_16_, n_n1303, x338x}, x107x);
	defparam lut_3391.LUT_SIZE = 6;
	defparam lut_3391.mask = 64'h0fff0fff10000000;

	lut_sub lut_3393 ({sk[1177], i_13_, i_12_, i_11_, i_18_, i_19_}, x596x);
	defparam lut_3393.LUT_SIZE = 6;
	defparam lut_3393.mask = 64'h0fff0fff00130000;

	lut_sub lut_3396 ({sk[1178], i_3_, i_13_, i_12_, i_19_}, x7298x);
	defparam lut_3396.LUT_SIZE = 5;
	defparam lut_3396.mask = 32'h55571000;

	lut_sub lut_3398 ({sk[1179], i_7_, i_8_, i_24_, i_22_}, x7299x);
	defparam lut_3398.LUT_SIZE = 5;
	defparam lut_3398.mask = 32'h55578000;

	lut_sub lut_3400 ({sk[1180], x210x, x281x, x596x, x7298x, x7299x}, x595x);
	defparam lut_3400.LUT_SIZE = 6;
	defparam lut_3400.mask = 64'h0fff0fff003f557f;

	lut_sub lut_3404 ({sk[1181], i_11_, n_n841, n_n245, n_n18}, x1762x);
	defparam lut_3404.LUT_SIZE = 5;
	defparam lut_3404.mask = 32'h55570100;

	lut_sub lut_3406 ({sk[1182], i_30_, i_14_, i_16_, i_34_, i_33_}, x620x);
	defparam lut_3406.LUT_SIZE = 6;
	defparam lut_3406.mask = 64'h0fff0fff00110313;

	lut_sub lut_3409 ({sk[1183], i_9_, i_8_, x224x, n_n307, x213x}, x7438x);
	defparam lut_3409.LUT_SIZE = 6;
	defparam lut_3409.mask = 64'h0fff0fff33333733;

	lut_sub lut_3412 ({sk[1184], i_7_, i_13_, i_32_, n_n629, x402x}, x9231x);
	defparam lut_3412.LUT_SIZE = 6;
	defparam lut_3412.mask = 64'h0fff0fff8fafffff;

	lut_sub lut_3423 ({sk[1185], i_17_, x10x, n_n1307, n_n853, n_n839}, x710x);
	defparam lut_3423.LUT_SIZE = 6;
	defparam lut_3423.mask = 64'h0fff0fff00070000;

	lut_sub lut_3426 ({sk[1186], i_14_, n_n1408, n_n629, x65x, x251x}, x7057x);
	defparam lut_3426.LUT_SIZE = 6;
	defparam lut_3426.mask = 64'h0fff0fff03570055;

	lut_sub lut_3429 ({sk[1187], i_7_, i_25_, i_26_, i_24_, i_22_}, x7695x);
	defparam lut_3429.LUT_SIZE = 6;
	defparam lut_3429.mask = 64'h0fff0fff80000000;

	lut_sub lut_3431 ({sk[1188], i_7_, x204x, x232x, x296x, x462x}, x6x);
	defparam lut_3431.LUT_SIZE = 6;
	defparam lut_3431.mask = 64'h0fff0fff00010000;

	lut_sub lut_3433 ({sk[1189], i_36_, i_29_, x25x, n_n793, n_n1397}, x22x);
	defparam lut_3433.LUT_SIZE = 6;
	defparam lut_3433.mask = 64'h0fff0fff00000100;

	lut_sub lut_3435 ({sk[1190], i_26_, i_17_, i_36_, x54x, n_n1406}, x8090x);
	defparam lut_3435.LUT_SIZE = 6;
	defparam lut_3435.mask = 64'h0fff0fff01000000;

	lut_sub lut_3437 ({sk[1191], i_21_, x102x, x105x, x107x, x8090x}, x32x);
	defparam lut_3437.LUT_SIZE = 6;
	defparam lut_3437.mask = 64'h0fff0fff15ff0000;

	lut_sub lut_3441 ({sk[1192], i_14_, i_16_, n_n1315, x299x}, x142x);
	defparam lut_3441.LUT_SIZE = 5;
	defparam lut_3441.mask = 32'h55571000;

	lut_sub lut_3443 ({sk[1193], n_n1375, n_n1213, n_n263, n_n363, x273x}, x9198x);
	defparam lut_3443.LUT_SIZE = 6;
	defparam lut_3443.mask = 64'h0fff0ffffafafac8;

	lut_sub lut_3450 ({sk[1194], i_36_, i_35_, x74x, x259x, n_n1459}, x182x);
	defparam lut_3450.LUT_SIZE = 6;
	defparam lut_3450.mask = 64'h0fff0fff00000100;

	lut_sub lut_3452 ({sk[1195], i_27_, x42x, n_n1504, n_n1322, n_n1323}, x184x);
	defparam lut_3452.LUT_SIZE = 6;
	defparam lut_3452.mask = 64'h0fff0fff00010000;

	lut_sub lut_3454 ({sk[1196], i_21_, x242x, n_n1216, n_n1374, n_n1387}, x234x);
	defparam lut_3454.LUT_SIZE = 6;
	defparam lut_3454.mask = 64'h0fff0fff00000001;

	lut_sub lut_3456 ({sk[1197], i_13_, n_n825, x517x, x433x, x65x}, x412x);
	defparam lut_3456.LUT_SIZE = 6;
	defparam lut_3456.mask = 64'h0fff0fff0f1f0000;

	lut_sub lut_3459 ({sk[1198], i_32_, i_34_, i_36_, i_35_, x419x}, x497x);
	defparam lut_3459.LUT_SIZE = 6;
	defparam lut_3459.mask = 64'h0fff0fff00040000;

	lut_sub lut_3461 ({sk[1199], i_14_, i_12_, i_17_, i_16_, x309x}, x507x);
	defparam lut_3461.LUT_SIZE = 6;
	defparam lut_3461.mask = 64'h0fff0fff44400000;

	lut_sub lut_3464 ({sk[1200], i_36_, i_29_, n_n793, n_n1397, n_n263}, x822x);
	defparam lut_3464.LUT_SIZE = 6;
	defparam lut_3464.mask = 64'h0fff0fff00000100;

	lut_sub lut_3466 ({sk[1201], i_32_, i_31_, i_29_, n_n1441, n_n608}, x827x);
	defparam lut_3466.LUT_SIZE = 6;
	defparam lut_3466.mask = 64'h0fff0fff10000000;

	lut_sub lut_3468 ({sk[1202], i_27_, i_28_, i_29_, n_n1433, n_n544}, x828x);
	defparam lut_3468.LUT_SIZE = 6;
	defparam lut_3468.mask = 64'h0fff0fff10000000;

	lut_sub lut_3470 ({sk[1203], i_23_, x493x, x43x, n_n1307, n_n1306}, x824x);
	defparam lut_3470.LUT_SIZE = 6;
	defparam lut_3470.mask = 64'h0fff0fff00010000;

	lut_sub lut_3472 ({sk[1204], i_23_, x43x, x76x, n_n1128, x368x}, x831x);
	defparam lut_3472.LUT_SIZE = 6;
	defparam lut_3472.mask = 64'h0fff0fff00010000;

	lut_sub lut_3474 ({sk[1205], i_13_, i_12_, i_16_, x320x, x393x}, x832x);
	defparam lut_3474.LUT_SIZE = 6;
	defparam lut_3474.mask = 64'h0fff0fff10000000;

	lut_sub lut_3476 ({sk[1206], i_36_, i_35_, n_n1375, n_n1433, n_n608}, x839x);
	defparam lut_3476.LUT_SIZE = 6;
	defparam lut_3476.mask = 64'h0fff0fff00000100;

	lut_sub lut_3478 ({sk[1207], i_14_, i_23_, i_16_, x396x}, x7887x);
	defparam lut_3478.LUT_SIZE = 5;
	defparam lut_3478.mask = 32'h55574000;

	lut_sub lut_3480 ({sk[1208], i_17_, i_34_, i_36_, n_n1375, x54x}, x7888x);
	defparam lut_3480.LUT_SIZE = 6;
	defparam lut_3480.mask = 64'h0fff0fff00010000;

	lut_sub lut_3482 ({sk[1209], i_16_, i_34_, i_36_, x242x, x80x}, x7878x);
	defparam lut_3482.LUT_SIZE = 6;
	defparam lut_3482.mask = 64'h0fff0fff00010000;

	lut_sub lut_3484 ({sk[1210], i_14_, i_16_, x242x, x51x, x483x}, x853x);
	defparam lut_3484.LUT_SIZE = 6;
	defparam lut_3484.mask = 64'h0fff0fff01000000;

	lut_sub lut_3486 ({sk[1211], i_7_, i_32_, i_34_, n_n1307, x280x}, x7868x);
	defparam lut_3486.LUT_SIZE = 6;
	defparam lut_3486.mask = 64'h0fff0fff01000000;

	lut_sub lut_3488 ({sk[1212], i_32_, i_34_, i_35_, n_n458, x267x}, x871x);
	defparam lut_3488.LUT_SIZE = 6;
	defparam lut_3488.mask = 64'h0fff0fff01000000;

	lut_sub lut_3490 ({sk[1213], i_27_, i_23_, i_17_, n_n242, x214x}, x872x);
	defparam lut_3490.LUT_SIZE = 6;
	defparam lut_3490.mask = 64'h0fff0fff10000000;

	lut_sub lut_3492 ({sk[1214], i_27_, i_36_, x242x, n_n355, x214x}, x873x);
	defparam lut_3492.LUT_SIZE = 6;
	defparam lut_3492.mask = 64'h0fff0fff00010000;

	lut_sub lut_3494 ({sk[1215], i_14_, i_13_, i_26_, i_23_, i_24_}, x7858x);
	defparam lut_3494.LUT_SIZE = 6;
	defparam lut_3494.mask = 64'h0fff0fff80808000;

	lut_sub lut_3497 ({sk[1216], i_27_, i_28_, i_31_, x224x, n_n1279}, x7859x);
	defparam lut_3497.LUT_SIZE = 6;
	defparam lut_3497.mask = 64'h0fff0fff10000000;

	lut_sub lut_3499 ({sk[1217], i_32_, i_36_, n_n1397, n_n358, x267x}, x876x);
	defparam lut_3499.LUT_SIZE = 6;
	defparam lut_3499.mask = 64'h0fff0fff00010000;

	lut_sub lut_3501 ({sk[1218], i_27_, i_23_, n_n1397, n_n1499, x16x}, x9230x);
	defparam lut_3501.LUT_SIZE = 6;
	defparam lut_3501.mask = 64'h0fff0ffffeffffff;

	lut_sub lut_3513 ({sk[1219], i_27_, i_28_, i_23_, i_21_, n_n1504}, x7830x);
	defparam lut_3513.LUT_SIZE = 6;
	defparam lut_3513.mask = 64'h0fff0fff10000000;

	lut_sub lut_3515 ({sk[1220], i_32_, i_36_, n_n458, x228x}, x894x);
	defparam lut_3515.LUT_SIZE = 5;
	defparam lut_3515.mask = 32'h55570100;

	lut_sub lut_3517 ({sk[1221], i_13_, i_12_, i_16_, x84x, x440x}, x895x);
	defparam lut_3517.LUT_SIZE = 6;
	defparam lut_3517.mask = 64'h0fff0fff10000000;

	lut_sub lut_3519 ({sk[1222], i_13_, i_31_, i_36_, i_35_, x501x}, x903x);
	defparam lut_3519.LUT_SIZE = 6;
	defparam lut_3519.mask = 64'h0fff0fff04000000;

	lut_sub lut_3521 ({sk[1223], i_36_, n_n1369, n_n1489, x323x, x291x}, x915x);
	defparam lut_3521.LUT_SIZE = 6;
	defparam lut_3521.mask = 64'h0fff0fff00000007;

	lut_sub lut_3524 ({sk[1224], i_8_, i_36_, i_35_, x64x, x571x}, x942x);
	defparam lut_3524.LUT_SIZE = 6;
	defparam lut_3524.mask = 64'h0fff0fff00100000;

	lut_sub lut_3526 ({sk[1225], i_35_, i_38_, i_29_, n_n1478, x394x}, x972x);
	defparam lut_3526.LUT_SIZE = 6;
	defparam lut_3526.mask = 64'h0fff0fff00100000;

	lut_sub lut_3528 ({sk[1226], i_34_, i_35_, i_38_, x344x, x327x}, x973x);
	defparam lut_3528.LUT_SIZE = 6;
	defparam lut_3528.mask = 64'h0fff0fff00000100;

	lut_sub lut_3530 ({sk[1227], i_28_, i_31_, i_29_, x218x, x270x}, x974x);
	defparam lut_3530.LUT_SIZE = 6;
	defparam lut_3530.mask = 64'h0fff0fff10000000;

	lut_sub lut_3532 ({sk[1228], i_30_, i_7_, i_2_, i_32_, x388x}, x999x);
	defparam lut_3532.LUT_SIZE = 6;
	defparam lut_3532.mask = 64'h0fff0fff40000000;

	lut_sub lut_3534 ({sk[1229], i_31_, i_38_, n_n1458, n_n1497, x57x}, x1000x);
	defparam lut_3534.LUT_SIZE = 6;
	defparam lut_3534.mask = 64'h0fff0fff00010000;

	lut_sub lut_3536 ({sk[1230], i_30_, i_8_, i_31_, x71x, x12x}, x1001x);
	defparam lut_3536.LUT_SIZE = 6;
	defparam lut_3536.mask = 64'h0fff0fff10000000;

	lut_sub lut_3538 ({sk[1231], x3x, n_n1397, x240x, x83x, x1028x}, x1025x);
	defparam lut_3538.LUT_SIZE = 6;
	defparam lut_3538.mask = 64'h0fff0fff00550057;

	lut_sub lut_3541 ({sk[1232], i_30_, i_8_, i_2_, x61x, x226x}, x1029x);
	defparam lut_3541.LUT_SIZE = 6;
	defparam lut_3541.mask = 64'h0fff0fff10000000;

	lut_sub lut_3543 ({sk[1233], i_30_, i_29_, n_n1353, x509x}, x1030x);
	defparam lut_3543.LUT_SIZE = 5;
	defparam lut_3543.mask = 32'h55571000;

	lut_sub lut_3545 ({sk[1234], i_2_, i_32_, x226x, x466x}, x1031x);
	defparam lut_3545.LUT_SIZE = 5;
	defparam lut_3545.mask = 32'h55571000;

	lut_sub lut_3547 ({sk[1235], i_28_, i_26_, i_29_, n_n762, n_n1359}, x1032x);
	defparam lut_3547.LUT_SIZE = 6;
	defparam lut_3547.mask = 64'h0fff0fff10000000;

	lut_sub lut_3549 ({sk[1236], i_30_, i_29_, n_n1353, n_n1423, n_n805}, x1041x);
	defparam lut_3549.LUT_SIZE = 6;
	defparam lut_3549.mask = 64'h0fff0fff01000000;

	lut_sub lut_3551 ({sk[1237], i_25_, i_26_, i_24_, n_n1288, x206x}, x1042x);
	defparam lut_3551.LUT_SIZE = 6;
	defparam lut_3551.mask = 64'h0fff0fff10000000;

	lut_sub lut_3553 ({sk[1238], i_6_, i_12_, n_n1307, x13x, x395x}, x1045x);
	defparam lut_3553.LUT_SIZE = 6;
	defparam lut_3553.mask = 64'h0fff0fff01000000;

	lut_sub lut_3555 ({sk[1239], i_9_, i_10_, i_2_, n_n1179, x313x}, x1060x);
	defparam lut_3555.LUT_SIZE = 6;
	defparam lut_3555.mask = 64'h0fff0fff00001000;

	lut_sub lut_3557 ({sk[1240], i_28_, i_25_, i_34_, i_29_, x212x}, x1062x);
	defparam lut_3557.LUT_SIZE = 6;
	defparam lut_3557.mask = 64'h0fff0fff04000000;

	lut_sub lut_3559 ({sk[1241], i_7_, i_8_, x224x, n_n1279, x70x}, x1063x);
	defparam lut_3559.LUT_SIZE = 6;
	defparam lut_3559.mask = 64'h0fff0fff01000000;

	lut_sub lut_3561 ({sk[1242], i_28_, i_26_, x738x}, x1070x);
	defparam lut_3561.LUT_SIZE = 4;
	defparam lut_3561.mask = 16'h5740;

	lut_sub lut_3563 ({sk[1243], i_28_, i_29_, n_n1523, n_n1251, x1078x}, x1071x);
	defparam lut_3563.LUT_SIZE = 6;
	defparam lut_3563.mask = 64'h0fff0fff005d0000;

	lut_sub lut_3566 ({sk[1244], i_28_, i_24_, i_22_, i_34_, x35x}, x1093x);
	defparam lut_3566.LUT_SIZE = 6;
	defparam lut_3566.mask = 64'h0fff0fff01000000;

	lut_sub lut_3568 ({sk[1245], i_27_, i_16_, i_22_}, x7629x);
	defparam lut_3568.LUT_SIZE = 4;
	defparam lut_3568.mask = 16'h5715;

	lut_sub lut_3571 ({sk[1246], i_24_, i_22_, n_n1511, x240x, x285x}, x1114x);
	defparam lut_3571.LUT_SIZE = 6;
	defparam lut_3571.mask = 64'h0fff0fff00070000;

	lut_sub lut_3574 ({sk[1247], i_7_, i_8_, n_n1478, x9x, x57x}, x1131x);
	defparam lut_3574.LUT_SIZE = 6;
	defparam lut_3574.mask = 64'h0fff0fff01000000;

	lut_sub lut_3576 ({sk[1248], i_28_, i_25_, i_26_, i_22_, x212x}, x1142x);
	defparam lut_3576.LUT_SIZE = 6;
	defparam lut_3576.mask = 64'h0fff0fff40000000;

	lut_sub lut_3578 ({sk[1249], i_25_, i_38_, x72x, x214x}, x1171x);
	defparam lut_3578.LUT_SIZE = 5;
	defparam lut_3578.mask = 32'h55570100;

	lut_sub lut_3580 ({sk[1250], i_30_, i_32_, i_35_, i_38_}, x7559x);
	defparam lut_3580.LUT_SIZE = 5;
	defparam lut_3580.mask = 32'h55574000;

	lut_sub lut_3582 ({sk[1251], i_30_, i_24_, n_n1179, x262x, x71x}, x1173x);
	defparam lut_3582.LUT_SIZE = 6;
	defparam lut_3582.mask = 64'h0fff0fff01000000;

	lut_sub lut_3584 ({sk[1252], i_32_, i_31_, n_n1361, x11x, x52x}, x1174x);
	defparam lut_3584.LUT_SIZE = 6;
	defparam lut_3584.mask = 64'h0fff0fff01000000;

	lut_sub lut_3586 ({sk[1253], i_28_, i_25_, i_29_, n_n1202, x206x}, x1175x);
	defparam lut_3586.LUT_SIZE = 6;
	defparam lut_3586.mask = 64'h0fff0fff10000000;

	lut_sub lut_3588 ({sk[1254], i_7_, x224x, n_n1279, n_n1288, n_n1059}, x1176x);
	defparam lut_3588.LUT_SIZE = 6;
	defparam lut_3588.mask = 64'h0fff0fff00010000;

	lut_sub lut_3590 ({sk[1255], i_10_, i_13_, i_34_, x239x, x272x}, x1206x);
	defparam lut_3590.LUT_SIZE = 6;
	defparam lut_3590.mask = 64'h0fff0fff01010001;

	lut_sub lut_3593 ({sk[1256], i_8_, i_25_, x250x, x214x}, x1207x);
	defparam lut_3593.LUT_SIZE = 5;
	defparam lut_3593.mask = 32'h55571000;

	lut_sub lut_3595 ({sk[1257], i_28_, i_34_, i_33_, i_38_, i_29_}, x7520x);
	defparam lut_3595.LUT_SIZE = 6;
	defparam lut_3595.mask = 64'h0fff0fff00200000;

	lut_sub lut_3597 ({sk[1258], i_22_, i_32_, x51x, n_n1497, x226x}, x1209x);
	defparam lut_3597.LUT_SIZE = 6;
	defparam lut_3597.mask = 64'h0fff0fff01000000;

	lut_sub lut_3599 ({sk[1259], i_8_, i_5_, i_6_, i_31_, n_n1279}, x7522x);
	defparam lut_3599.LUT_SIZE = 6;
	defparam lut_3599.mask = 64'h0fff0fff40000000;

	lut_sub lut_3601 ({sk[1260], i_12_, i_17_, x43x, x46x, x7491x}, x1234x);
	defparam lut_3601.LUT_SIZE = 6;
	defparam lut_3601.mask = 64'h0fff0fff01010100;

	lut_sub lut_3604 ({sk[1261], i_11_, i_19_, x429x, x272x}, x1239x);
	defparam lut_3604.LUT_SIZE = 5;
	defparam lut_3604.mask = 32'h55571000;

	lut_sub lut_3606 ({sk[1262], i_8_, i_18_, x60x, n_n706, x379x}, x1240x);
	defparam lut_3606.LUT_SIZE = 6;
	defparam lut_3606.mask = 64'h0fff0fff15111111;

	lut_sub lut_3609 ({sk[1263], i_18_, i_32_, x42x, x60x, x429x}, x1285x);
	defparam lut_3609.LUT_SIZE = 6;
	defparam lut_3609.mask = 64'h0fff0fff01000000;

	lut_sub lut_3611 ({sk[1264], n_n372, n_n294, n_n371, n_n316, n_n284}, x1297x);
	defparam lut_3611.LUT_SIZE = 6;
	defparam lut_3611.mask = 64'h0fff0fff13333333;

	lut_sub lut_3616 ({sk[1265], n_n372, n_n300, n_n294, n_n371, n_n284}, x1304x);
	defparam lut_3616.LUT_SIZE = 6;
	defparam lut_3616.mask = 64'h0fff0fff007f00ff;

	lut_sub lut_3621 ({sk[1266], i_28_, i_31_, i_29_, x238x, x408x}, x1353x);
	defparam lut_3621.LUT_SIZE = 6;
	defparam lut_3621.mask = 64'h0fff0fff10000000;

	lut_sub lut_3623 ({sk[1267], i_32_, i_31_, i_29_, x218x, x315x}, x1354x);
	defparam lut_3623.LUT_SIZE = 6;
	defparam lut_3623.mask = 64'h0fff0fff10000000;

	lut_sub lut_3625 ({sk[1268], n_n1307, n_n841, x518x, x226x}, x1364x);
	defparam lut_3625.LUT_SIZE = 5;
	defparam lut_3625.mask = 32'h55570001;

	lut_sub lut_3627 ({sk[1269], i_28_, i_31_, i_29_, x238x, x421x}, x1365x);
	defparam lut_3627.LUT_SIZE = 6;
	defparam lut_3627.mask = 64'h0fff0fff10000000;

	lut_sub lut_3629 ({sk[1270], i_34_, i_35_, i_38_, n_n1302, x394x}, x1366x);
	defparam lut_3629.LUT_SIZE = 6;
	defparam lut_3629.mask = 64'h0fff0fff00000100;

	lut_sub lut_3631 ({sk[1271], i_9_, i_10_, i_8_, x11x, x390x}, x1369x);
	defparam lut_3631.LUT_SIZE = 6;
	defparam lut_3631.mask = 64'h0fff0fff00001000;

	lut_sub lut_3633 ({sk[1272], i_32_, i_33_, n_n1361, x518x, x229x}, x1390x);
	defparam lut_3633.LUT_SIZE = 6;
	defparam lut_3633.mask = 64'h0fff0fff01000000;

	lut_sub lut_3635 ({sk[1273], i_31_, n_n1361, n_n1478, n_n1191, x41x}, x1391x);
	defparam lut_3635.LUT_SIZE = 6;
	defparam lut_3635.mask = 64'h0fff0fff00010000;

	lut_sub lut_3637 ({sk[1274], i_9_, i_10_, n_n1118, n_n1279, x390x}, x1393x);
	defparam lut_3637.LUT_SIZE = 6;
	defparam lut_3637.mask = 64'h0fff0fff00000100;

	lut_sub lut_3639 ({sk[1275], i_32_, i_31_, n_n1361, x257x, x218x}, x1394x);
	defparam lut_3639.LUT_SIZE = 6;
	defparam lut_3639.mask = 64'h0fff0fff01000000;

	lut_sub lut_3641 ({sk[1276], i_9_, i_10_, n_n1361, x50x, x52x}, x1400x);
	defparam lut_3641.LUT_SIZE = 6;
	defparam lut_3641.mask = 64'h0fff0fff00000100;

	lut_sub lut_3643 ({sk[1277], i_32_, n_n1361, n_n1478, n_n1191, x229x}, x1401x);
	defparam lut_3643.LUT_SIZE = 6;
	defparam lut_3643.mask = 64'h0fff0fff00010000;

	lut_sub lut_3645 ({sk[1278], i_10_, i_19_, n_n584, x329x}, x1418x);
	defparam lut_3645.LUT_SIZE = 5;
	defparam lut_3645.mask = 32'h55570001;

	lut_sub lut_3647 ({sk[1279], i_30_, i_28_, i_25_, i_26_, i_38_}, x7300x);
	defparam lut_3647.LUT_SIZE = 6;
	defparam lut_3647.mask = 64'h0fff0fff40000000;

	lut_sub lut_3649 ({sk[1280], n_n584, n_n1033, x377x, x1444x, x414x}, x1439x);
	defparam lut_3649.LUT_SIZE = 6;
	defparam lut_3649.mask = 64'h0fff0fff0707070f;

	lut_sub lut_3653 ({sk[1281], i_33_, i_38_, x210x, x282x}, x1448x);
	defparam lut_3653.LUT_SIZE = 5;
	defparam lut_3653.mask = 32'h55570100;

	lut_sub lut_3655 ({sk[1282], i_13_, i_37_, n_n1458, x386x}, x1482x);
	defparam lut_3655.LUT_SIZE = 5;
	defparam lut_3655.mask = 32'h55570100;

	lut_sub lut_3657 ({sk[1283], i_13_, i_17_, i_16_, n_n1305, x366x}, x7228x);
	defparam lut_3657.LUT_SIZE = 6;
	defparam lut_3657.mask = 64'h0fff0fff10000000;

	lut_sub lut_3659 ({sk[1284], n_n1369, n_n1318, n_n1302, x498x, x522x}, x1484x);
	defparam lut_3659.LUT_SIZE = 6;
	defparam lut_3659.mask = 64'h0fff0fff00000007;

	lut_sub lut_3662 ({sk[1285], i_14_, i_37_, n_n1018, n_n1225, x31x}, x1485x);
	defparam lut_3662.LUT_SIZE = 6;
	defparam lut_3662.mask = 64'h0fff0fff00010000;

	lut_sub lut_3664 ({sk[1286], i_14_, i_16_, n_n1369, x42x, n_n1318}, x7212x);
	defparam lut_3664.LUT_SIZE = 6;
	defparam lut_3664.mask = 64'h0fff0fff01000000;

	lut_sub lut_3666 ({sk[1287], i_23_, i_18_, i_17_, x268x, x256x}, x7195x);
	defparam lut_3666.LUT_SIZE = 6;
	defparam lut_3666.mask = 64'h0fff0fff10000000;

	lut_sub lut_3668 ({sk[1288], i_14_, i_16_, i_29_, n_n1216, x248x}, x7199x);
	defparam lut_3668.LUT_SIZE = 6;
	defparam lut_3668.mask = 64'h0fff0fff10000000;

	lut_sub lut_3670 ({sk[1289], i_14_, i_34_, i_35_, n_n1322, x261x}, x9232x);
	defparam lut_3670.LUT_SIZE = 6;
	defparam lut_3670.mask = 64'h0fff0ffffeffffff;

	lut_sub lut_3682 ({sk[1290], i_10_, i_14_, i_16_, x48x, x41x}, x1517x);
	defparam lut_3682.LUT_SIZE = 6;
	defparam lut_3682.mask = 64'h0fff0fff10000000;

	lut_sub lut_3684 ({sk[1291], i_34_, i_35_, i_37_}, x7175x);
	defparam lut_3684.LUT_SIZE = 4;
	defparam lut_3684.mask = 16'h5710;

	lut_sub lut_3686 ({sk[1292], i_10_, i_33_, i_35_, i_37_, x43x}, x7176x);
	defparam lut_3686.LUT_SIZE = 6;
	defparam lut_3686.mask = 64'h0fff0fff10000000;

	lut_sub lut_3688 ({sk[1293], i_13_, i_16_, i_33_, i_37_, x358x}, x1535x);
	defparam lut_3688.LUT_SIZE = 6;
	defparam lut_3688.mask = 64'h0fff0fff10000000;

	lut_sub lut_3690 ({sk[1294], i_27_, i_28_, i_29_, n_n1443, x499x}, x7151x);
	defparam lut_3690.LUT_SIZE = 6;
	defparam lut_3690.mask = 64'h0fff0fff10000000;

	lut_sub lut_3692 ({sk[1295], i_10_, i_5_, i_4_, i_0_, i_37_}, x7138x);
	defparam lut_3692.LUT_SIZE = 6;
	defparam lut_3692.mask = 64'h0fff0fff40000000;

	lut_sub lut_3694 ({sk[1296], i_27_, x42x, n_n1202, x351x, x1574x}, x1565x);
	defparam lut_3694.LUT_SIZE = 6;
	defparam lut_3694.mask = 64'h0fff0fff00070000;

	lut_sub lut_3697 ({sk[1297], i_20_, i_23_, n_n1397, n_n984, x94x}, x1579x);
	defparam lut_3697.LUT_SIZE = 6;
	defparam lut_3697.mask = 64'h0fff0fff00000100;

	lut_sub lut_3699 ({sk[1298], i_35_, i_37_, n_n1311, x29x, x445x}, x1606x);
	defparam lut_3699.LUT_SIZE = 6;
	defparam lut_3699.mask = 64'h0fff0fff00000001;

	lut_sub lut_3701 ({sk[1299], i_30_, i_27_, x42x, x323x, x246x}, x1607x);
	defparam lut_3701.LUT_SIZE = 6;
	defparam lut_3701.mask = 64'h0fff0fff01000000;

	lut_sub lut_3703 ({sk[1300], n_n1369, n_n1314, n_n1318, x76x, n_n1302}, x1609x);
	defparam lut_3703.LUT_SIZE = 6;
	defparam lut_3703.mask = 64'h0fff0fff00000001;

	lut_sub lut_3705 ({sk[1301], i_14_, i_37_, n_n1202, n_n1459, x409x}, x1667x);
	defparam lut_3705.LUT_SIZE = 6;
	defparam lut_3705.mask = 64'h0fff0fff00010000;

	lut_sub lut_3707 ({sk[1302], i_7_, i_13_, i_16_, n_n1499, x318x}, x1668x);
	defparam lut_3707.LUT_SIZE = 6;
	defparam lut_3707.mask = 64'h0fff0fff00001000;

	lut_sub lut_3709 ({sk[1303], i_20_, i_7_, i_16_, x290x, x84x}, x1672x);
	defparam lut_3709.LUT_SIZE = 6;
	defparam lut_3709.mask = 64'h0fff0fff00000010;

	lut_sub lut_3711 ({sk[1304], i_7_, i_34_, i_35_, i_37_}, x6957x);
	defparam lut_3711.LUT_SIZE = 5;
	defparam lut_3711.mask = 32'h55571000;

	lut_sub lut_3713 ({sk[1305], i_27_, x73x, n_n504, n_n1288, n_n329}, x1732x);
	defparam lut_3713.LUT_SIZE = 6;
	defparam lut_3713.mask = 64'h0fff0fff00010000;

	lut_sub lut_3715 ({sk[1306], i_34_, i_35_, i_29_, i_37_, n_n793}, x6924x);
	defparam lut_3715.LUT_SIZE = 6;
	defparam lut_3715.mask = 64'h0fff0fff00100000;

	lut_sub lut_3717 ({sk[1307], i_32_, i_34_, i_35_, n_n620, x365x}, x1734x);
	defparam lut_3717.LUT_SIZE = 6;
	defparam lut_3717.mask = 64'h0fff0fff01000000;

	lut_sub lut_3719 ({sk[1308], i_9_, i_14_, i_11_, i_37_, n_n130}, x6901x);
	defparam lut_3719.LUT_SIZE = 6;
	defparam lut_3719.mask = 64'h0fff0fff10000000;

	lut_sub lut_3721 ({sk[1309], n_n1443, n_n504, n_n245, x63x, x361x}, x1745x);
	defparam lut_3721.LUT_SIZE = 6;
	defparam lut_3721.mask = 64'h0fff0fff00000001;

	lut_sub lut_3723 ({sk[1310], i_25_, x287x, x84x, x94x}, x9221x);
	defparam lut_3723.LUT_SIZE = 5;
	defparam lut_3723.mask = 32'h5557eee0;

	lut_sub lut_3728 ({sk[1311], n_n1318, n_n916, x319x, x487x, x334x}, x9227x);
	defparam lut_3728.LUT_SIZE = 6;
	defparam lut_3728.mask = 64'h0fff0ffffffffefc;

	lut_sub lut_3739 ({sk[1312], n_n1118, n_n152, x461x, x274x, x1482x}, x7231x);
	defparam lut_3739.LUT_SIZE = 6;
	defparam lut_3739.mask = 64'h0fff0fff55555557;

	lut_sub lut_3742 ({sk[1313], x351x, x484x, x489x, x256x, x7228x}, x7232x);
	defparam lut_3742.LUT_SIZE = 6;
	defparam lut_3742.mask = 64'h0fff0fff05553777;

	lut_sub lut_3746 ({sk[1314], x7111x, x7112x, x1474x, x7245x}, x7246x);
	defparam lut_3746.LUT_SIZE = 5;
	defparam lut_3746.mask = 32'h55577fff;

	lut_sub lut_3751 ({sk[1315], n_n805, n_n1466, x278x, x425x, x454x}, x9216x);
	defparam lut_3751.LUT_SIZE = 6;
	defparam lut_3751.mask = 64'h0fff0ffffffffff8;

	lut_sub lut_3762 ({sk[1316], i_19_, x53x, x423x, x435x, x28x}, x9215x);
	defparam lut_3762.LUT_SIZE = 6;
	defparam lut_3762.mask = 64'h0fff0fffffc0ff80;

	lut_sub lut_3766 ({sk[1317], x52x, x264x, x231x, x521x, x1239x}, x7481x);
	defparam lut_3766.LUT_SIZE = 6;
	defparam lut_3766.mask = 64'h0fff0fff5555557f;

	lut_sub lut_3770 ({sk[1318], i_22_, n_n1478, x354x, x100x, x254x}, x7482x);
	defparam lut_3770.LUT_SIZE = 6;
	defparam lut_3770.mask = 64'h0fff0fff111f1111;

	lut_sub lut_3773 ({sk[1319], n_n1300, n_n1472, x298x, x409x, x1114x}, x7620x);
	defparam lut_3773.LUT_SIZE = 6;
	defparam lut_3773.mask = 64'h0fff0fff55555557;

	lut_sub lut_3776 ({sk[1320], i_7_, i_28_, n_n1472, x112x, x429x}, x7687x);
	defparam lut_3776.LUT_SIZE = 6;
	defparam lut_3776.mask = 64'h0fff0fff37333333;

	lut_sub lut_3779 ({sk[1321], x7495x, x7496x, x7504x, x7505x}, x7710x);
	defparam lut_3779.LUT_SIZE = 5;
	defparam lut_3779.mask = 32'h55577fff;

	lut_sub lut_3784 ({sk[1322], i_24_, n_n1179, x71x, x335x, x974x}, x7738x);
	defparam lut_3784.LUT_SIZE = 6;
	defparam lut_3784.mask = 64'h0fff0fff55575555;

	lut_sub lut_3787 ({sk[1323], i_32_, x207x, x66x, x972x, x973x}, x7739x);
	defparam lut_3787.LUT_SIZE = 6;
	defparam lut_3787.mask = 64'h0fff0fff777f7777;

	lut_sub lut_3791 ({sk[1324], x7729x, x7730x, x7740x, x7738x, x7739x}, x7742x);
	defparam lut_3791.LUT_SIZE = 6;
	defparam lut_3791.mask = 64'h0fff0fff7fffffff;

	lut_sub lut_3797 ({sk[1325], n_n1863, x7384x, n_n1866, x7742x}, x7744x);
	defparam lut_3797.LUT_SIZE = 5;
	defparam lut_3797.mask = 32'h55577fff;

	lut_sub lut_3802 ({sk[1326], i_31_, i_34_, x80x, x535x, x915x}, x7812x);
	defparam lut_3802.LUT_SIZE = 6;
	defparam lut_3802.mask = 64'h0fff0fff55555557;

	lut_sub lut_3805 ({sk[1327], i_13_, i_16_, n_n1147, x362x, x516x}, x7813x);
	defparam lut_3805.LUT_SIZE = 6;
	defparam lut_3805.mask = 64'h0fff0fff57030303;

	lut_sub lut_3808 ({sk[1328], i_31_, n_n1397, x267x, x325x, x328x}, x9208x);
	defparam lut_3808.LUT_SIZE = 6;
	defparam lut_3808.mask = 64'h0fff0ffffffffff8;

	lut_sub lut_3819 ({sk[1329], i_32_, i_34_, n_n880, x513x, x497x}, x7934x);
	defparam lut_3819.LUT_SIZE = 6;
	defparam lut_3819.mask = 64'h0fff0fff57555555;

	lut_sub lut_3822 ({sk[1330], i_33_, n_n1441, x8x, x38x, x308x}, x9207x);
	defparam lut_3822.LUT_SIZE = 6;
	defparam lut_3822.mask = 64'h0fff0ffffafafac8;

	lut_sub lut_3829 ({sk[1331], n_n1314, n_n1141, n_n820, n_n846, x348x}, x9200x);
	defparam lut_3829.LUT_SIZE = 6;
	defparam lut_3829.mask = 64'h0fff0fffeeeeeee0;

	lut_sub lut_3836 ({sk[1332], i_13_, i_16_, n_n1375, x337x, x9200x}, x7965x);
	defparam lut_3836.LUT_SIZE = 6;
	defparam lut_3836.mask = 64'h0fff0fff3b0a0a0a;

	lut_sub lut_3839 ({sk[1333], i_30_, i_28_, i_31_, i_29_, n_n1202}, x9229x);
	defparam lut_3839.LUT_SIZE = 6;
	defparam lut_3839.mask = 64'h0fff0fffefffffff;

	lut_sub lut_3851 ({sk[1334], i_31_, n_n1441, n_n1429, x393x, x382x}, x9196x);
	defparam lut_3851.LUT_SIZE = 6;
	defparam lut_3851.mask = 64'h0fff0ffffffffff8;

	lut_sub lut_3862 ({sk[1335], x7796x, x7797x, x7808x, x7809x}, x8074x);
	defparam lut_3862.LUT_SIZE = 5;
	defparam lut_3862.mask = 32'h55577fff;

	lut_sub lut_3867 ({sk[1336], x7814x, x8062x, x8063x, x7812x, x7813x}, x8075x);
	defparam lut_3867.LUT_SIZE = 6;
	defparam lut_3867.mask = 64'h0fff0fff7fffffff;

	lut_sub lut_3873 ({sk[1337], x8068x, x8069x, x8072x, x8073x}, x8076x);
	defparam lut_3873.LUT_SIZE = 5;
	defparam lut_3873.mask = 32'h55577fff;


endmodule