module seq (
	i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, 
	i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, 
	i_18_, i_19_, i_20_, i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, 
	i_28_, i_29_, i_30_, i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, 
	i_38_, i_39_, i_40_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, 
	o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, 
	o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, 
	o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_);

input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, i_18_, i_19_, i_20_, i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_, i_30_, i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_, i_39_, i_40_;

output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_;

wire n1, n2, n5, n6, n7, n8, n9, n10, n14, n16, n18, n19, n20, n23, n24, n25, n26, n22, n28, n29, n27, n32, n33, n30, n35, n36, n37, n34, n41, n38, n44, n45, n46, n47, n48, n43, n50, n51, n52, n53, n54, n55, n49, n58, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70, n71, n73, n78, n79, n80, n81, n82, n76, n83, n84, n86, n87, n88, n90, n85, n94, n95, n97, n98, n99, n96, n101, n103, n100, n104, n105, n106, n107, n115, n113, n112, n118, n119, n120, n117, n125, n126, n133, n131, n135, n136, n138, n134, n141, n140, n139, n145, n143, n142, n146, n147, n152, n157, n154, n160, n158, n161, n162, n165, n163, n164, n167, n166, n170, n171, n169, n173, n174, n172, n179, n177, n178, n175, n180, n181, n182, n184, n185, n183, n188, n186, n190, n196, n197, n198, n199, n195, n202, n201, n200, n205, n204, n203, n209, n207, n206, n210, n217, n215, n214, n221, n222, n219, n220, n218, n223, n227, n228, n226, n224, n231, n232, n230, n229, n234, n235, n233, n239, n237, n238, n236, n241, n240, n244, n242, n247, n246, n250, n251, n249, n253, n256, n259, n263, n264, n265, n266, n267, n268, n269, n270, n262, n271, n274, n275, n276, n277, n273, n278, n284, n283, n290, n288, n289, n287, n292, n291, n295, n294, n293, n297, n296, n298, n304, n306, n307, n302, n309, n312, n308, n316, n317, n314, n315, n313, n320, n318, n324, n325, n322, n323, n321, n326, n331, n332, n329, n330, n328, n335, n336, n334, n333, n337, n340, n341, n339, n343, n344, n345, n342, n347, n348, n346, n350, n349, n353, n352, n351, n355, n356, n357, n358, n354, n359, n363, n362, n365, n367, n364, n369, n374, n375, n376, n380, n381, n379, n378, n384, n385, n383, n382, n387, n386, n390, n391, n389, n388, n392, n396, n395, n394, n400, n398, n397, n401, n403, n404, n402, n406, n407, n405, n408, n410, n414, n418, n419, n420, n421, n422, n423, n424, n417, n427, n426, n425, n430, n431, n429, n428, n433, n434, n435, n432, n438, n439, n440, n436, n441, n443, n444, n442, n445, n451, n450, n457, n458, n455, n456, n454, n460, n459, n462, n461, n464, n463, n470, n468, n474, n473, n472, n477, n476, n475, n479, n478, n481, n484, n482, n486, n487, n485, n490, n491, n489, n494, n492, n495, n500, n506, n507, n509, n510, n511, n504, n514, n512, n516, n515, n517, n520, n526, n528, n525, n529, n537, n535, n534, n540, n541, n539, n538, n542, n545, n544, n551, n550, n548, n549, n547, n554, n553, n552, n557, n558, n556, n555, n562, n560, n561, n559, n566, n563, n567, n570, n573, n574, n575, n576, n578, n579, n572, n580, n581, n584, n583, n582, n585, n591, n590, n594, n595, n593, n592, n599, n597, n598, n596, n602, n603, n601, n600, n604, n605, n610, n609, n614, n613, n612, n617, n615, n619, n620, n618, n623, n627, n632, n633, n634, n635, n636, n637, n631, n638, n640, n643, n646, n644, n649, n653, n651, n656, n654, n660, n658, n659, n657, n663, n661, n666, n665, n664, n668, n667, n670, n671, n669, n673, n674, n675, n676, n677, n672, n680, n678, n679, n683, n682, n681, n685, n684, n687, n689, n686, n690, n691, n696, n697, n695, n699, n702, n701, n703, n707, n709, n711, n712, n713, n715, n714, n716, n718, n719, n717, n722, n723, n721, n720, n725, n724, n726, n727, n728, n729, n730, n735, n733, n731, n736, n740, n739, n742, n746, n751, n750, n752, n756, n755, n754, n760, n758, n762, n761, n765, n770, n768, n771, n772, n773, n774, n775, n784, n783, n786, n785, n789, n787, n792, n793, n791, n794, n796, n797, n795, n799, n800, n804, n803, n807, n808, n806, n810, n809, n811, n818, n816, n815, n820, n821, n822, n823, n819, n825, n824, n827, n828, n826, n830, n829, n832, n831, n834, n833, n837, n836, n835, n838, n841, n840, n843, n844, n845, n846, n847, n842, n849, n848, n850, n853, n856, n857, n858, n855, n860, n859, n862, n863, n864, n861, n865, n871, n868, n872, n878, n877, n882, n883, n884, n885, n886, n881, n889, n890, n888, n892, n891, n895, n894, n893, n897, n896, n899, n900, n898, n902, n901, n905, n904, n903, n906, n907, n910, n909, n913, n912, n916, n915, n914, n917, n919, n923, n921, n922, n920, n926, n924, n928, n927, n932, n929, n933, n936, n937, n938, n939, n940, n935, n942, n941, n944, n943, n945, n948, n946, n949, n951, n952, n950, n953, n957, n954, n963, n964, n965, n968, n966, n969, n970, n971, n972, n973, n975, n976, n980, n977, n982, n981, n984, n985, n983, n987, n990, n989, n993, n992, n995, n994, n997, n996, n998, n1001, n1004, n1008, n1012, n1013, n1014, n1015, n1016, n1011, n1017, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1027, n1029, n1030, n1032, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1064, n1065, n1066, n1067, n1068, n1069, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1088, n1089, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1113, n1114, n1116, n1117, n1119, n1120, n1122, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1139, n1140, n1143, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1155, n1154, n1157, n1158, n1160, n1162, n1161, n1163, n1165, n1167, n1168, n1169, n1172, n1173, n1175, n1174, n1177, n1176, n1179, n1178, n1180, n1181, n1182, n1183, n1184, n1187, n1185, n1188, n1189, n1190, n1192, n1191, n1194, n1195, n1196, n1197, n1199, n1198, n1201, n1202, n1204, n1205, n1206, n1210, n1214, n1213, n1215, n1218, n1220, n1221, n1223, n1224, n1229, n1228, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1241, n1245, n1248, n1247, n1249, n1250, n1251, n1252, n1254, n1255, n1256, n1257, n1258, n1260, n1259, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1270, n1271, n1272, n1274, n1273, n1276, n1277, n1278, n1279, n1280, n1282, n1283, n1284, n1288, n1287, n1289, n1291, n1295, n1294, n1296, n1297, n1301, n1302, n1303, n1305, n1309, n1308, n1307, n1310, n1311, n1312, n1314, n1313, n1318, n1319, n1321, n1323, n1324, n1325, n1327, n1328, n1330, n1333, n1334, n1335, n1336, n1337, n1342;

assign o_0_ = ( (~ n1011) ) ;
 assign o_1_ = ( (~ n881) ) ;
 assign o_2_ = ( (~ n672) ) ;
 assign o_3_ = ( (~ n504) ) ;
 assign o_4_ = ( (~ n417) ) ;
 assign o_5_ = ( n104 ) | ( n105 ) | ( n106 ) | ( n107 ) | ( (~ n1176) ) | ( (~ n1178) ) | ( (~ n1183) ) | ( (~ n1188) ) ;
 assign o_6_ = ( (~ n262) ) ;
 assign o_7_ = ( (~ n100) ) ;
 assign o_8_ = ( (~ n1) ) ;
 assign o_9_ = ( (~ n96) ) ;
 assign o_10_ = ( (~ n86) ) | ( n94 ) | ( n95 ) | ( (~ n972) ) | ( (~ n983) ) ;
 assign o_11_ = ( (~ n85) ) ;
 assign o_12_ = ( i_8_  &  n2  &  (~ n398)  &  (~ n827) ) ;
 assign o_13_ = ( (~ n84) ) ;
 assign o_14_ = ( (~ n83) ) ;
 assign o_15_ = ( (~ n52) ) ;
 assign o_16_ = ( (~ n76) ) ;
 assign o_17_ = ( n69 ) | ( n70 ) | ( n71 ) | ( n73 ) | ( (~ n432) ) | ( (~ n953) ) | ( (~ n1310) ) | ( (~ n1312) ) ;
 assign o_18_ = ( (~ n935) ) ;
 assign o_19_ = ( (~ n67) ) ;
 assign o_20_ = ( (~ n842) ) ;
 assign o_21_ = ( (~ n66) ) ;
 assign o_22_ = ( n58 ) | ( n60 ) | ( n61 ) | ( n62 ) | ( n63 ) | ( n64 ) | ( n65 ) | ( (~ n754) ) ;
 assign o_23_ = ( (~ n49) ) ;
 assign o_24_ = ( (~ n43) ) ;
 assign o_25_ = ( (~ n34) ) ;
 assign o_26_ = ( (~ n30) ) ;
 assign o_27_ = ( (~ n27) ) ;
 assign o_28_ = ( (~ n22) ) ;
 assign o_29_ = ( (~ n686) ) ;
 assign o_30_ = ( n19 ) | ( n20 ) | ( (~ n1247) ) ;
 assign o_31_ = ( n5 ) | ( n6 ) | ( n7 ) | ( n8 ) | ( n9 ) | ( (~ n22) ) ;
 assign o_32_ = ( (~ n1254) ) ;
 assign o_33_ = ( (~ n631) ) ;
 assign o_34_ = ( (~ n572) ) ;
 assign n1 = ( n165  &  n52  &  n163 ) | ( n165  &  n52  &  n164 ) ;
 assign n2 = ( (~ i_37_)  &  (~ n1337) ) | ( (~ n244)  &  (~ n561)  &  (~ n1337) ) ;
 assign n5 = ( n125  &  (~ n834) ) | ( (~ i_39_)  &  n125  &  (~ n230) ) ;
 assign n6 = ( n484  &  n640  &  (~ n683) ) ;
 assign n7 = ( (~ n162)  &  (~ n203)  &  n643 ) ;
 assign n8 = ( n113  &  n125 ) ;
 assign n9 = ( n374  &  (~ n376) ) | ( n374  &  (~ n834) ) ;
 assign n10 = ( (~ n403)  &  (~ n1047)  &  (~ n1084) ) ;
 assign n14 = ( (~ n403)  &  (~ n1047)  &  (~ n1081) ) ;
 assign n16 = ( (~ n407)  &  (~ n1047)  &  (~ n1084) ) ;
 assign n18 = ( (~ n407)  &  (~ n1047)  &  (~ n1081) ) ;
 assign n19 = ( n649  &  (~ n1129) ) | ( (~ n820)  &  (~ n1129) ) | ( (~ n1032)  &  (~ n1129) ) ;
 assign n20 = ( n16 ) | ( n18 ) | ( n10 ) | ( n14 ) ;
 assign n23 = ( n334 ) | ( n1086 ) ;
 assign n24 = ( n238 ) | ( n580 ) | ( n638 ) ;
 assign n25 = ( n238 ) | ( n638 ) | ( n553 ) ;
 assign n26 = ( n895 ) | ( n964 ) | ( n1074 ) ;
 assign n22 = ( n23  &  n24  &  n25  &  n26 ) ;
 assign n28 = ( (~ n9)  &  n44  &  (~ n113) ) | ( (~ n9)  &  n44  &  n707 ) ;
 assign n29 = ( n273  &  n287  &  n304  &  n690  &  (~ n691)  &  (~ n695)  &  n1140  &  n1143 ) ;
 assign n27 = ( n28  &  n29 ) ;
 assign n32 = ( n490 ) | ( n339 ) | ( n712 ) ;
 assign n33 = ( n35  &  (~ n112)  &  (~ n117) ) ;
 assign n30 = ( n32  &  n33  &  (~ n131) ) ;
 assign n35 = ( (~ i_34_) ) | ( n682 ) | ( n1042 ) | ( n1065 ) ;
 assign n36 = ( n680  &  n678 ) | ( n680  &  n679 ) ;
 assign n37 = ( n29  &  (~ n126) ) ;
 assign n34 = ( n22  &  n35  &  n36  &  n28  &  n37 ) ;
 assign n41 = ( (~ i_37_)  &  i_39_  &  (~ n665) ) ;
 assign n38 = ( n41  &  (~ n1077) ) | ( (~ n271)  &  (~ n665)  &  (~ n1077) ) ;
 assign n44 = ( (~ n5)  &  (~ n20)  &  (~ n38)  &  n283  &  n689  &  (~ n701)  &  (~ n703)  &  n1139 ) ;
 assign n45 = ( (~ n9)  &  n23  &  (~ n131)  &  n713 ) ;
 assign n46 = ( n297 ) | ( i_39_ ) | ( n638 ) ;
 assign n47 = ( (~ n113) ) | ( n707 ) ;
 assign n48 = ( n25  &  n26  &  n1254 ) ;
 assign n43 = ( n36  &  n44  &  n33  &  n37  &  n45  &  n46  &  n47  &  n48 ) ;
 assign n50 = ( n238 ) | ( n474 ) | ( n398 ) | ( n726 ) ;
 assign n51 = ( n721 ) | ( n271 ) | ( i_35_ ) | ( i_34_ ) ;
 assign n52 = ( (~ i_7_) ) | ( (~ i_33_) ) ;
 assign n53 = ( (~ i_37_) ) | ( n389 ) | ( n728 ) ;
 assign n54 = ( n553 ) | ( n727 ) | ( n728 ) ;
 assign n55 = ( n556 ) | ( n729 ) | ( n730 ) ;
 assign n49 = ( n50  &  n51  &  n52  &  n53  &  n54  &  n55  &  (~ n731)  &  (~ n1267) ) ;
 assign n58 = ( (~ n173)  &  (~ n761) ) | ( (~ n334)  &  (~ n761) ) | ( (~ n729)  &  (~ n761) ) ;
 assign n60 = ( (~ i_40_)  &  n765 ) | ( (~ i_40_)  &  (~ n315)  &  n760 ) ;
 assign n61 = ( (~ n682)  &  n760 ) ;
 assign n62 = ( n772  &  n773  &  n774 ) ;
 assign n63 = ( (~ n768)  &  (~ n796) ) | ( n775  &  (~ n796)  &  (~ n1097) ) ;
 assign n64 = ( (~ i_7_)  &  i_32_  &  n772 ) ;
 assign n65 = ( i_37_  &  (~ n312)  &  n771  &  (~ n827) ) ;
 assign n66 = ( n794  &  i_33_  &  i_7_ ) | ( n794  &  i_33_  &  n787 ) ;
 assign n67 = ( n899  &  n900  &  n898 ) | ( n899  &  n900  &  n219 ) ;
 assign n69 = ( (~ i_29_)  &  n957  &  (~ n1336) ) | ( n957  &  n954  &  (~ n1336) ) ;
 assign n70 = ( n735  &  n733  &  (~ n1024) ) ;
 assign n71 = ( (~ n554)  &  (~ n1104) ) | ( (~ n784)  &  (~ n1104) ) ;
 assign n73 = ( (~ n426)  &  (~ n1307) ) | ( (~ n426)  &  n484  &  (~ n683) ) ;
 assign n78 = ( n315 ) | ( n969 ) ;
 assign n79 = ( n970 ) | ( n554 ) ;
 assign n80 = ( n963 ) | ( n964 ) | ( n712 ) | ( n490 ) ;
 assign n81 = ( n828 ) | ( n926 ) | ( n312 ) | ( n271 ) ;
 assign n82 = ( n965 ) | ( i_40_ ) | ( n455 ) ;
 assign n76 = ( n78  &  n79  &  n80  &  n81  &  n82  &  (~ n966) ) ;
 assign n83 = ( (~ i_13_)  &  n515 ) | ( n398  &  n515 ) | ( n515  &  n971 ) ;
 assign n84 = ( n515  &  n580 ) | ( n515  &  n312 ) | ( n515  &  n581 ) ;
 assign n86 = ( n965 ) | ( n597 ) ;
 assign n87 = ( n394 ) | ( n1094 ) | ( n1095 ) ;
 assign n88 = ( n451 ) | ( n975 ) | ( n976 ) ;
 assign n90 = ( n972  &  n164 ) | ( n972  &  n965 ) ;
 assign n85 = ( n86  &  n87  &  n88  &  n90  &  (~ n977) ) ;
 assign n94 = ( i_20_  &  i_21_  &  n987  &  i_15_ ) ;
 assign n95 = ( n640  &  n981 ) | ( n613  &  n640  &  (~ n656) ) ;
 assign n97 = ( n462 ) | ( n329 ) | ( n1022 ) | ( n653 ) ;
 assign n98 = ( n161 ) | ( n158 ) | ( n162 ) ;
 assign n99 = ( n52  &  n139  &  (~ n147) ) | ( n52  &  (~ n147)  &  n152 ) ;
 assign n96 = ( n97  &  n98  &  n99 ) ;
 assign n101 = ( n180  &  n97  &  n181  &  n182 ) ;
 assign n103 = ( n165  &  n1039 ) | ( n165  &  n820  &  n185 ) ;
 assign n100 = ( n99  &  n101  &  n103  &  (~ n186) ) ;
 assign n104 = ( n251  &  n359 ) | ( (~ i_23_)  &  n251  &  (~ n354) ) ;
 assign n105 = ( (~ n1061)  &  (~ n1085) ) | ( (~ i_37_)  &  (~ n271)  &  (~ n1085) ) ;
 assign n106 = ( n113  &  n374 ) | ( n374  &  (~ n1083) ) ;
 assign n107 = ( n113  &  n369 ) | ( n326  &  n369 ) | ( n113  &  (~ n1134) ) | ( n326  &  (~ n1134) ) ;
 assign n115 = ( i_2_ ) | ( i_3_ ) | ( i_1_ ) | ( i_4_ ) ;
 assign n113 = ( i_39_  &  n740 ) ;
 assign n112 = ( n115  &  n113  &  (~ n1068) ) | ( n115  &  (~ n235)  &  (~ n1068) ) ;
 assign n118 = ( (~ n309)  &  n709 ) | ( i_0_  &  i_4_  &  (~ n309) ) ;
 assign n119 = ( (~ n312)  &  n711 ) ;
 assign n120 = ( (~ n164)  &  (~ n1111) ) ;
 assign n117 = ( n118  &  n120 ) | ( n119  &  n120 ) | ( n118  &  (~ n1146) ) | ( n119  &  (~ n1146) ) ;
 assign n125 = ( (~ i_24_)  &  (~ n357)  &  (~ n407) ) ;
 assign n126 = ( (~ n666)  &  (~ n679) ) | ( (~ n514)  &  (~ n666)  &  (~ n1075) ) ;
 assign n133 = ( i_2_  &  (~ n341) ) ;
 assign n131 = ( n120  &  n133  &  (~ n312) ) | ( n133  &  (~ n312)  &  (~ n1146) ) ;
 assign n135 = ( i_11_ ) | ( (~ n1027) ) ;
 assign n136 = ( (~ i_17_) ) | ( n284 ) ;
 assign n138 = ( i_12_ ) | ( n406 ) ;
 assign n134 = ( n135  &  n138 ) | ( n136  &  n138 ) | ( n135  &  (~ n171) ) | ( n136  &  (~ n171) ) ;
 assign n141 = ( n145  &  (~ n849) ) | ( n145  &  n1152  &  n1153 ) ;
 assign n140 = ( (~ i_16_) ) | ( n284 ) ;
 assign n139 = ( n134  &  n141  &  n135 ) | ( n134  &  n141  &  n140 ) ;
 assign n145 = ( i_12_ ) | ( (~ i_15_) ) | ( (~ i_17_) ) | ( (~ n171) ) ;
 assign n143 = ( n1153  &  n1152 ) ;
 assign n142 = ( n145  &  n143 ) | ( n145  &  (~ n849) ) ;
 assign n146 = ( n134  &  n135 ) | ( n134  &  n140 ) ;
 assign n147 = ( (~ n142)  &  (~ n619)  &  (~ n1029) ) | ( (~ n146)  &  (~ n619)  &  (~ n1029) ) ;
 assign n152 = ( n619 ) | ( n289 ) ;
 assign n157 = ( (~ i_18_) ) | ( n426 ) ;
 assign n154 = ( (~ i_15_)  &  n157 ) | ( n157  &  (~ n1155) ) ;
 assign n160 = ( n395 ) | ( (~ n1155) ) ;
 assign n158 = ( (~ i_19_)  &  n160 ) | ( i_21_  &  n160 ) | ( n154  &  n160 ) ;
 assign n161 = ( (~ i_23_) ) | ( n184 ) ;
 assign n162 = ( n1032 ) | ( n312 ) ;
 assign n165 = ( n237 ) | ( n786 ) | ( n863 ) | ( (~ n1017) ) ;
 assign n163 = ( n997 ) | ( n535 ) ;
 assign n164 = ( (~ i_38_) ) | ( n904 ) ;
 assign n167 = ( i_12_  &  n1027 ) ;
 assign n166 = ( i_22_  &  (~ n157) ) | ( i_15_  &  i_22_  &  n167 ) ;
 assign n170 = ( i_15_  &  i_22_ ) ;
 assign n171 = ( i_11_  &  n1027 ) ;
 assign n169 = ( i_19_  &  n166 ) | ( i_19_  &  n170  &  n171 ) ;
 assign n173 = ( (~ i_40_) ) | ( n440 ) ;
 assign n174 = ( (~ i_38_) ) | ( i_39_ ) ;
 assign n172 = ( n173  &  n174 ) ;
 assign n179 = ( n221 ) | ( n685 ) | ( n426 ) | ( n646 ) ;
 assign n177 = ( (~ i_33_) ) | ( (~ i_34_) ) | ( i_35_ ) ;
 assign n178 = ( i_32_ ) | ( n426 ) | ( n916 ) ;
 assign n175 = ( (~ i_21_)  &  n179 ) | ( n179  &  n177 ) | ( n179  &  n178 ) ;
 assign n180 = ( n164 ) | ( n556 ) | ( n1021 ) | ( n653 ) ;
 assign n181 = ( (~ i_22_)  &  n1036 ) | ( n175  &  n1036 ) | ( (~ i_22_)  &  (~ n1154) ) | ( n175  &  (~ n1154) ) ;
 assign n182 = ( n1157  &  n1032 ) | ( n1157  &  n1039 ) ;
 assign n184 = ( (~ i_22_) ) | ( (~ i_24_) ) ;
 assign n185 = ( n1040 ) | ( n668 ) ;
 assign n183 = ( n184 ) | ( n154 ) | ( n185 ) ;
 assign n188 = ( (~ n164) ) | ( (~ n804) ) ;
 assign n186 = ( (~ n183)  &  (~ n312) ) | ( n188  &  (~ n312)  &  (~ n581) ) ;
 assign n190 = ( (~ n1042)  &  (~ n1158) ) | ( (~ n164)  &  (~ n1042)  &  (~ n1045) ) ;
 assign n196 = ( (~ n113) ) | ( (~ n640) ) | ( n751 ) | ( n1036 ) ;
 assign n197 = ( i_37_ ) | ( n329 ) | ( n898 ) ;
 assign n198 = ( (~ i_24_) ) | ( (~ n251) ) | ( n357 ) | ( n658 ) ;
 assign n199 = ( (~ n190)  &  n580 ) | ( (~ n190)  &  n910 ) | ( (~ n190)  &  n1045 ) ;
 assign n195 = ( n196  &  n197  &  n198  &  n199 ) ;
 assign n202 = ( (~ i_18_) ) | ( n201 ) ;
 assign n201 = ( n284  &  n276 ) ;
 assign n200 = ( (~ i_19_)  &  n202 ) | ( n202  &  n201 ) ;
 assign n205 = ( (~ i_15_) ) | ( (~ i_18_) ) | ( (~ i_19_) ) | ( (~ n251) ) ;
 assign n204 = ( (~ i_9_) ) | ( n294 ) ;
 assign n203 = ( n205  &  n200 ) | ( n205  &  n204 ) ;
 assign n209 = ( i_29_  &  n348 ) | ( (~ i_29_)  &  n975 ) | ( n348  &  n975 ) ;
 assign n207 = ( i_29_ ) | ( n294 ) ;
 assign n206 = ( (~ i_30_)  &  n209 ) | ( n209  &  n207 ) ;
 assign n210 = ( (~ n367)  &  (~ n479) ) | ( (~ n230)  &  (~ n237)  &  (~ n367) ) ;
 assign n217 = ( n204 ) | ( (~ n702) ) | ( n726 ) ;
 assign n215 = ( n1082  &  n1067 ) ;
 assign n214 = ( n206  &  (~ n210)  &  n217 ) | ( (~ n210)  &  n217  &  n215 ) ;
 assign n221 = ( n1024 ) | ( n389 ) ;
 assign n222 = ( n389  &  n490 ) | ( n487  &  n490 ) | ( n389  &  n1045 ) | ( n487  &  n1045 ) ;
 assign n219 = ( (~ i_40_) ) | ( n1046 ) ;
 assign n220 = ( (~ i_34_) ) | ( n1023 ) ;
 assign n218 = ( n221  &  n222  &  n219 ) | ( n221  &  n222  &  n220 ) ;
 assign n223 = ( i_10_  &  i_27_ ) ;
 assign n227 = ( n1051 ) | ( n295 ) | ( n1061 ) ;
 assign n228 = ( n965  &  n462 ) | ( n315  &  n462 ) | ( n965  &  n1058 ) | ( n315  &  n1058 ) ;
 assign n226 = ( n1061 ) | ( n841 ) | ( n862 ) ;
 assign n224 = ( (~ i_11_)  &  n227  &  n228 ) | ( n227  &  n228  &  n226 ) ;
 assign n231 = ( n237 ) | ( n292 ) ;
 assign n232 = ( i_36_ ) | ( n271 ) ;
 assign n230 = ( i_36_ ) | ( n729 ) ;
 assign n229 = ( (~ i_39_)  &  n231  &  n232 ) | ( n231  &  n232  &  n230 ) ;
 assign n234 = ( n387 ) | ( (~ n740) ) ;
 assign n235 = ( i_39_ ) | ( n462 ) ;
 assign n233 = ( n234  &  n235  &  n229 ) ;
 assign n239 = ( n580 ) | ( n535 ) ;
 assign n237 = ( (~ i_39_) ) | ( (~ i_40_) ) ;
 assign n238 = ( i_37_ ) | ( n1023 ) ;
 assign n236 = ( n239  &  n237 ) | ( n239  &  n238 ) ;
 assign n241 = ( (~ i_40_)  &  n238 ) | ( n238  &  n297 ) | ( (~ i_40_)  &  n440 ) | ( n297  &  n440 ) ;
 assign n240 = ( n241  &  n236 ) ;
 assign n244 = ( (~ i_38_) ) | ( i_40_ ) ;
 assign n242 = ( (~ i_37_)  &  (~ n188) ) | ( (~ n188)  &  n244 ) ;
 assign n247 = ( i_12_ ) | ( i_11_ ) ;
 assign n246 = ( n170  &  (~ n204)  &  n247 ) ;
 assign n250 = ( i_18_  &  n170 ) ;
 assign n251 = ( (~ n403) ) | ( (~ n407) ) ;
 assign n249 = ( n246  &  (~ n685) ) | ( n250  &  n251  &  (~ n685) ) ;
 assign n253 = ( (~ i_37_)  &  n249  &  (~ n610) ) | ( (~ i_37_)  &  (~ n610)  &  (~ n910) ) ;
 assign n256 = ( n253  &  (~ n389) ) | ( (~ n389)  &  (~ n487)  &  (~ n910) ) ;
 assign n259 = ( n113  &  (~ n1058) ) | ( (~ n682)  &  (~ n1058) ) ;
 assign n263 = ( n204 ) | ( n539 ) | ( (~ n702) ) | ( n1048 ) ;
 assign n264 = ( n1047 ) | ( n367 ) | ( i_32_ ) | ( i_13_ ) ;
 assign n265 = ( n904 ) | ( n1045 ) | ( n1050 ) ;
 assign n266 = ( n1160  &  n215 ) | ( n1160  &  n1022 ) | ( n1160  &  n347 ) ;
 assign n267 = ( n242  &  (~ n256)  &  n1163 ) | ( (~ n256)  &  n314  &  n1163 ) ;
 assign n268 = ( (~ i_40_)  &  n233 ) | ( n224  &  n233 ) | ( (~ i_40_)  &  n1060 ) | ( n224  &  n1060 ) ;
 assign n269 = ( n1165  &  n218 ) | ( n1165  &  n1059 ) ;
 assign n270 = ( n195  &  n1168  &  n1069 ) | ( n195  &  n1168  &  n821 ) ;
 assign n262 = ( n263  &  n264  &  n265  &  n266  &  n267  &  n268  &  n269  &  n270 ) ;
 assign n271 = ( i_38_ ) | ( (~ i_40_) ) ;
 assign n274 = ( n276 ) | ( n1076 ) ;
 assign n275 = ( n271 ) | ( n665 ) ;
 assign n276 = ( (~ i_11_) ) | ( (~ i_15_) ) ;
 assign n277 = ( n474 ) | ( n1051 ) | ( n1078 ) ;
 assign n273 = ( n274  &  n276 ) | ( n275  &  n276 ) | ( n274  &  n277 ) | ( n275  &  n277 ) ;
 assign n278 = ( (~ n455)  &  (~ n990)  &  (~ n1051) ) | ( (~ n804)  &  (~ n990)  &  (~ n1051) ) ;
 assign n284 = ( (~ i_12_) ) | ( (~ i_15_) ) ;
 assign n283 = ( (~ n8)  &  n277  &  (~ n278) ) | ( (~ n8)  &  (~ n278)  &  n284 ) ;
 assign n290 = ( n201 ) | ( n152 ) | ( n1078 ) ;
 assign n288 = ( n1077  &  n274 ) ;
 assign n289 = ( n665 ) | ( n1030 ) ;
 assign n287 = ( n290  &  n288 ) | ( n290  &  n289 ) ;
 assign n292 = ( i_36_ ) | ( i_37_ ) ;
 assign n291 = ( (~ i_39_)  &  n232  &  n235 ) | ( n232  &  n235  &  n292 ) ;
 assign n295 = ( i_15_ ) | ( n294 ) ;
 assign n294 = ( i_7_ ) | ( i_5_ ) ;
 assign n293 = ( n295  &  i_12_ ) | ( n295  &  n294 ) ;
 assign n297 = ( i_38_ ) | ( n1023 ) ;
 assign n296 = ( (~ i_39_)  &  (~ i_40_) ) | ( (~ i_40_)  &  n238 ) | ( (~ i_39_)  &  n297 ) | ( n238  &  n297 ) ;
 assign n298 = ( (~ n293)  &  (~ n358)  &  (~ n1051) ) | ( (~ n358)  &  (~ n404)  &  (~ n1051) ) ;
 assign n304 = ( (~ n41) ) | ( n274 ) ;
 assign n306 = ( n1169  &  n291 ) | ( n1169  &  n1060 ) ;
 assign n307 = ( (~ n113)  &  n289 ) | ( n289  &  n1172 ) | ( (~ n113)  &  (~ n1342) ) | ( n1172  &  (~ n1342) ) ;
 assign n302 = ( (~ n38)  &  (~ n112)  &  n273  &  n283  &  n287  &  n304  &  n306  &  n307 ) ;
 assign n309 = ( i_7_ ) | ( n312 ) ;
 assign n312 = ( i_34_ ) | ( n398 ) ;
 assign n308 = ( n309  &  n312 ) | ( n309  &  (~ n1091) ) | ( n312  &  (~ n1173) ) | ( (~ n1091)  &  (~ n1173) ) ;
 assign n316 = ( n226  &  n308 ) | ( (~ n247)  &  n308 ) | ( n226  &  n1093 ) | ( (~ n247)  &  n1093 ) ;
 assign n317 = ( n1174  &  n970 ) | ( n1174  &  n455  &  n597 ) ;
 assign n314 = ( n898 ) | ( n473 ) ;
 assign n315 = ( (~ i_37_) ) | ( n174 ) ;
 assign n313 = ( n316  &  n317  &  n314 ) | ( n316  &  n317  &  n315 ) ;
 assign n320 = ( (~ i_15_) ) | ( (~ n247) ) | ( n990 ) ;
 assign n318 = ( (~ i_15_)  &  n320 ) | ( i_18_  &  n320 ) | ( (~ n251)  &  n320 ) ;
 assign n324 = ( n284 ) | ( n1089 ) ;
 assign n325 = ( n276 ) | ( n1089 ) ;
 assign n322 = ( i_21_ ) | ( n398 ) ;
 assign n323 = ( i_19_ ) | ( n318 ) ;
 assign n321 = ( n324  &  n325  &  n322 ) | ( n324  &  n325  &  n323 ) ;
 assign n326 = ( (~ i_40_)  &  (~ n1083) ) ;
 assign n331 = ( i_34_ ) | ( n1073 ) | ( n928 ) ;
 assign n332 = ( n389  &  n561 ) | ( n1088  &  n561 ) | ( n389  &  n1061 ) | ( n1088  &  n1061 ) ;
 assign n329 = ( (~ i_39_) ) | ( i_40_ ) ;
 assign n330 = ( n473 ) | ( n727 ) ;
 assign n328 = ( n331  &  n332  &  n329 ) | ( n331  &  n332  &  n330 ) ;
 assign n335 = ( n619 ) | ( n173 ) | ( n295 ) ;
 assign n336 = ( i_38_ ) | ( n638 ) ;
 assign n334 = ( (~ i_38_) ) | ( n387 ) ;
 assign n333 = ( n335  &  n336  &  n288 ) | ( n335  &  n336  &  n334 ) ;
 assign n337 = ( (~ i_25_)  &  i_26_ ) ;
 assign n340 = ( i_4_  &  i_1_ ) ;
 assign n341 = ( (~ i_0_) ) | ( i_7_ ) ;
 assign n339 = ( n340  &  (~ n1091) ) | ( n341  &  (~ n1091) ) ;
 assign n343 = ( n1172 ) | ( n1083 ) ;
 assign n344 = ( n339 ) | ( n312 ) | ( n1092 ) ;
 assign n345 = ( n1049 ) | ( n597 ) | ( n556 ) | ( n1048 ) ;
 assign n342 = ( n343  &  n344  &  n345  &  n86 ) ;
 assign n347 = ( (~ i_29_) ) | ( n294 ) ;
 assign n348 = ( (~ i_28_) ) | ( n294 ) ;
 assign n346 = ( (~ i_30_)  &  n347  &  n348 ) | ( n294  &  n347  &  n348 ) ;
 assign n350 = ( n238 ) | ( n668 ) ;
 assign n349 = ( n350  &  n289 ) ;
 assign n353 = ( n284 ) | ( n403 ) | ( i_14_ ) | ( n349 ) ;
 assign n352 = ( i_34_ ) | ( n491 ) ;
 assign n351 = ( n353  &  n346 ) | ( n353  &  n329 ) | ( n353  &  n352 ) ;
 assign n355 = ( (~ i_15_) ) | ( i_21_ ) ;
 assign n356 = ( n580 ) | ( n439 ) | ( n312 ) ;
 assign n357 = ( n751 ) | ( n1044 ) ;
 assign n358 = ( i_40_ ) | ( n1024 ) ;
 assign n354 = ( n355  &  n357 ) | ( n356  &  n357 ) | ( n355  &  n358 ) | ( n356  &  n358 ) ;
 assign n359 = ( (~ n177)  &  (~ n916)  &  (~ n1081) ) | ( (~ n177)  &  (~ n916)  &  (~ n1084) ) ;
 assign n363 = ( (~ i_0_) ) | ( n751 ) | ( n841 ) ;
 assign n362 = ( i_36_ ) | ( (~ i_37_) ) | ( n329 ) | ( n363 ) ;
 assign n365 = ( n234 ) | ( n808 ) ;
 assign n367 = ( i_12_ ) | ( n404 ) ;
 assign n364 = ( (~ i_13_) ) | ( i_31_ ) | ( n365 ) | ( n367 ) ;
 assign n369 = ( (~ n403)  &  (~ n751)  &  (~ n1084) ) ;
 assign n374 = ( (~ i_24_)  &  (~ n357)  &  (~ n403) ) ;
 assign n375 = ( n206  &  i_30_ ) | ( n206  &  n347 ) ;
 assign n376 = ( i_39_  &  (~ n113) ) | ( (~ n113)  &  n230 ) ;
 assign n380 = ( n1147 ) | ( n1096 ) ;
 assign n381 = ( i_40_ ) | ( n970 ) | ( n455 ) ;
 assign n379 = ( (~ i_13_) ) | ( n1057 ) ;
 assign n378 = ( n380  &  n381  &  n376 ) | ( n380  &  n381  &  n379 ) ;
 assign n384 = ( i_13_ ) | ( n230 ) | ( n237 ) | ( (~ n1017) ) ;
 assign n385 = ( (~ i_40_) ) | ( n389 ) | ( n398 ) | ( n554 ) ;
 assign n383 = ( i_32_ ) | ( (~ i_39_) ) | ( n177 ) | ( n462 ) ;
 assign n382 = ( (~ i_13_)  &  n384  &  n385 ) | ( n384  &  n385  &  n383 ) ;
 assign n387 = ( i_39_ ) | ( i_40_ ) ;
 assign n386 = ( (~ i_37_)  &  n219 ) | ( n219  &  n387 ) ;
 assign n390 = ( i_34_ ) | ( n164 ) | ( n1041 ) ;
 assign n391 = ( n330  &  n561 ) | ( n804  &  n561 ) | ( n330  &  n358 ) | ( n804  &  n358 ) ;
 assign n389 = ( i_36_ ) | ( n1038 ) ;
 assign n388 = ( n390  &  n391  &  n386 ) | ( n390  &  n391  &  n389 ) ;
 assign n392 = ( (~ i_24_)  &  n295 ) | ( n295  &  n294 ) ;
 assign n396 = ( n204 ) | ( (~ n247) ) | ( n355 ) ;
 assign n395 = ( (~ i_18_) ) | ( n355 ) ;
 assign n394 = ( (~ n251)  &  n396 ) | ( n396  &  n395 ) ;
 assign n400 = ( (~ i_17_) ) | ( n398 ) ;
 assign n398 = ( i_32_ ) | ( (~ i_33_) ) ;
 assign n397 = ( (~ i_16_)  &  n400 ) | ( n400  &  n398 ) ;
 assign n401 = ( i_12_  &  i_11_ ) | ( n276  &  i_11_ ) | ( i_12_  &  n284 ) | ( n276  &  n284 ) ;
 assign n403 = ( (~ i_11_) ) | ( n294 ) ;
 assign n404 = ( i_11_ ) | ( n294 ) ;
 assign n402 = ( n138  &  n140 ) | ( n403  &  n140 ) | ( n138  &  n404 ) | ( n403  &  n404 ) ;
 assign n406 = ( (~ i_15_) ) | ( (~ i_16_) ) ;
 assign n407 = ( (~ i_12_) ) | ( n294 ) ;
 assign n405 = ( n402  &  i_14_ ) | ( n402  &  n406 ) | ( n402  &  n407 ) ;
 assign n408 = ( n204  &  n400 ) | ( n204  &  n405 ) | ( n400  &  (~ n1190) ) | ( n405  &  (~ n1190) ) ;
 assign n410 = ( (~ n294)  &  (~ n312)  &  (~ n1149) ) | ( (~ n294)  &  (~ n312)  &  (~ n1189) ) ;
 assign n414 = ( (~ i_39_)  &  (~ n1064) ) | ( (~ i_39_)  &  (~ n1177) ) ;
 assign n418 = ( i_40_  &  (~ n1330) ) | ( n86  &  n1148  &  (~ n1330) ) ;
 assign n419 = ( n1205  &  n1085 ) | ( n1205  &  n928 ) ;
 assign n420 = ( n388  &  n219 ) | ( n1042  &  n219 ) | ( n388  &  n970 ) | ( n1042  &  n970 ) ;
 assign n421 = ( n1204  &  n810 ) | ( n1204  &  n408 ) ;
 assign n422 = ( (~ n414)  &  n487 ) | ( (~ n414)  &  n1096  &  n1202 ) ;
 assign n423 = ( (~ i_31_)  &  n1198 ) | ( (~ n410)  &  n1198  &  n1201 ) ;
 assign n424 = ( n1194  &  n1195  &  n1196  &  n87  &  n35  &  n1197 ) ;
 assign n417 = ( n418  &  n378  &  n419  &  n420  &  n421  &  n422  &  n423  &  n424 ) ;
 assign n427 = ( n426 ) | ( n389 ) | ( n1107 ) ;
 assign n426 = ( n1019  &  i_5_ ) | ( n1019  &  n276 ) ;
 assign n425 = ( n427  &  n426 ) | ( n427  &  n389 ) | ( n427  &  n322 ) ;
 assign n430 = ( (~ i_3_) ) | ( n429 ) ;
 assign n431 = ( (~ i_2_) ) | ( n429 ) ;
 assign n429 = ( (~ i_0_) ) | ( i_32_ ) ;
 assign n428 = ( n430  &  n431  &  n340 ) | ( n430  &  n431  &  n429 ) ;
 assign n433 = ( (~ n223) ) | ( n387 ) | ( n890 ) | ( (~ n1017) ) ;
 assign n434 = ( (~ n735) ) | ( (~ n733) ) | ( n1030 ) ;
 assign n435 = ( n1024  &  n1103 ) | ( n1103  &  n1104 ) | ( n1024  &  (~ n1224) ) | ( n1104  &  (~ n1224) ) ;
 assign n432 = ( n433  &  n52  &  n434  &  n435 ) ;
 assign n438 = ( i_5_ ) | ( (~ i_31_) ) | ( n1023 ) ;
 assign n439 = ( (~ i_35_) ) | ( i_36_ ) | ( (~ i_37_) ) ;
 assign n440 = ( i_38_ ) | ( (~ i_39_) ) ;
 assign n436 = ( (~ n284)  &  n439 ) | ( n438  &  n439 ) | ( (~ n284)  &  n440 ) | ( n438  &  n440 ) ;
 assign n441 = ( (~ i_39_)  &  n271 ) ;
 assign n443 = ( (~ i_35_) ) | ( n1073 ) ;
 assign n444 = ( (~ i_36_) ) | ( n1100 ) ;
 assign n442 = ( n387  &  n237 ) | ( n443  &  n237 ) | ( n387  &  n444 ) | ( n443  &  n444 ) ;
 assign n445 = ( (~ n329)  &  (~ n1092) ) | ( (~ n329)  &  (~ n456)  &  (~ n944) ) ;
 assign n451 = ( i_29_ ) | ( i_30_ ) ;
 assign n450 = ( (~ i_5_)  &  i_28_  &  (~ n1082) ) | ( (~ i_5_)  &  n451  &  (~ n1082) ) ;
 assign n457 = ( (~ i_15_) ) | ( i_17_ ) | ( n591 ) | ( n948 ) ;
 assign n458 = ( (~ i_36_)  &  (~ n450) ) | ( n173  &  (~ n450) ) | ( (~ n450)  &  n863 ) ;
 assign n455 = ( (~ i_37_) ) | ( n474 ) ;
 assign n456 = ( i_9_ ) | ( i_5_ ) ;
 assign n454 = ( n457  &  n458  &  n455 ) | ( n457  &  n458  &  n456 ) ;
 assign n460 = ( (~ i_4_)  &  i_32_ ) | ( i_32_  &  n429 ) | ( (~ i_4_)  &  (~ n709) ) | ( n429  &  (~ n709) ) ;
 assign n459 = ( n430  &  n431  &  n460 ) ;
 assign n462 = ( i_36_ ) | ( n491 ) ;
 assign n461 = ( i_36_  &  n462 ) | ( (~ i_39_)  &  n462 ) ;
 assign n464 = ( i_11_  &  (~ n456) ) ;
 assign n463 = ( (~ n1106)  &  (~ n1218) ) | ( n464  &  (~ n1037)  &  (~ n1106) ) ;
 assign n470 = ( i_36_ ) | ( (~ n1030) ) | ( n1110 ) ;
 assign n468 = ( (~ i_40_)  &  (~ n463)  &  n470 ) | ( (~ n463)  &  n470  &  (~ n1215) ) ;
 assign n474 = ( (~ i_38_) ) | ( (~ i_39_) ) ;
 assign n473 = ( (~ i_0_) ) | ( n1054 ) ;
 assign n472 = ( n244  &  n474  &  n473 ) | ( n244  &  n474  &  n387 ) ;
 assign n477 = ( (~ i_9_) ) | ( (~ i_14_) ) | ( (~ n726) ) | ( n860 ) ;
 assign n476 = ( (~ i_14_) ) | ( (~ n726) ) ;
 assign n475 = ( n477  &  n476 ) | ( n477  &  (~ n849) ) ;
 assign n479 = ( n462 ) | ( n904 ) ;
 assign n478 = ( i_13_  &  (~ i_15_) ) | ( (~ i_15_)  &  n479 ) | ( i_13_  &  (~ n702) ) | ( n479  &  (~ n702) ) ;
 assign n481 = ( n53  &  i_5_ ) | ( n53  &  n398 ) | ( n53  &  n352 ) ;
 assign n484 = ( (~ i_23_)  &  (~ n398) ) ;
 assign n482 = ( (~ n322)  &  (~ n804)  &  (~ n1045) ) | ( n484  &  (~ n804)  &  (~ n1045) ) ;
 assign n486 = ( n1107  &  n322 ) ;
 assign n487 = ( (~ i_37_) ) | ( n271 ) ;
 assign n485 = ( n220  &  (~ n482) ) | ( (~ n482)  &  n486 ) | ( (~ n482)  &  n487 ) ;
 assign n490 = ( i_40_ ) | ( n580 ) ;
 assign n491 = ( (~ i_37_) ) | ( i_38_ ) ;
 assign n489 = ( n490  &  n491 ) ;
 assign n494 = ( n556 ) | ( n897 ) | ( n1106 ) ;
 assign n492 = ( i_18_  &  n494 ) | ( n355  &  n494 ) | ( n494  &  (~ n982) ) ;
 assign n495 = ( (~ n808)  &  (~ n1213) ) | ( (~ n475)  &  (~ n808)  &  (~ n821) ) ;
 assign n500 = ( (~ n312)  &  (~ n436) ) | ( (~ n312)  &  (~ n1221) ) | ( (~ n312)  &  (~ n1223) ) ;
 assign n506 = ( n454  &  n580 ) | ( n580  &  (~ n1017) ) | ( n454  &  n1104 ) | ( (~ n1017)  &  n1104 ) ;
 assign n507 = ( n472  &  n784 ) | ( n894  &  n784 ) | ( n472  &  n163 ) | ( n894  &  n163 ) ;
 assign n509 = ( n1024  &  n468 ) | ( n427  &  n468 ) | ( n1024  &  n539 ) | ( n427  &  n539 ) ;
 assign n510 = ( n1232  &  n1233  &  n426 ) | ( n1232  &  n1233  &  n485 ) ;
 assign n511 = ( n1105  &  n1230  &  n1231 ) | ( (~ n1210)  &  n1230  &  n1231 ) ;
 assign n504 = ( n432  &  (~ n495)  &  (~ n500)  &  n506  &  n507  &  n509  &  n510  &  n511 ) ;
 assign n514 = ( i_31_ ) | ( n312 ) ;
 assign n512 = ( n152  &  n350 ) | ( n350  &  (~ n476) ) | ( n152  &  n514 ) | ( (~ n476)  &  n514 ) ;
 assign n516 = ( n312 ) | ( n1040 ) ;
 assign n515 = ( n52  &  n516 ) | ( n52  &  n173  &  n334 ) ;
 assign n517 = ( i_9_  &  (~ n1079) ) | ( (~ n773)  &  (~ n1079) ) ;
 assign n520 = ( (~ i_31_)  &  (~ n234)  &  (~ n247) ) | ( (~ i_31_)  &  (~ n240)  &  (~ n247) ) ;
 assign n526 = ( (~ i_5_) ) | ( n517 ) | ( n1023 ) ;
 assign n528 = ( n490  &  n926 ) | ( n1111  &  n926 ) | ( n490  &  n804 ) | ( n1111  &  n804 ) ;
 assign n525 = ( (~ n520)  &  n526  &  n528 ) ;
 assign n529 = ( (~ i_34_)  &  (~ n292)  &  (~ n474) ) | ( (~ i_34_)  &  (~ n292)  &  (~ n580) ) ;
 assign n537 = ( n389  &  n665 ) | ( n665  &  n784 ) | ( n389  &  (~ n1030) ) | ( n784  &  (~ n1030) ) ;
 assign n535 = ( (~ i_37_) ) | ( n1023 ) ;
 assign n534 = ( n173  &  (~ n529)  &  n537 ) | ( (~ n529)  &  n537  &  n535 ) ;
 assign n540 = ( n897 ) | ( n836 ) ;
 assign n541 = ( n539 ) | ( n235 ) ;
 assign n539 = ( i_35_ ) | ( n1020 ) ;
 assign n538 = ( n540  &  n541  &  n229 ) | ( n540  &  n541  &  n539 ) ;
 assign n542 = ( (~ i_15_)  &  i_39_  &  (~ n238) ) ;
 assign n545 = ( (~ i_35_)  &  (~ i_37_)  &  (~ n804) ) ;
 assign n544 = ( (~ n514)  &  n542 ) | ( (~ n514)  &  n545  &  (~ n726) ) ;
 assign n551 = ( n862 ) | ( n1114 ) | ( n963 ) ;
 assign n550 = ( (~ i_0_) ) | ( i_1_ ) | ( i_2_ ) ;
 assign n548 = ( n751 ) | ( n444 ) ;
 assign n549 = ( n177 ) | ( n230 ) | ( (~ n237) ) ;
 assign n547 = ( n551  &  n550 ) | ( n551  &  n548  &  n549 ) ;
 assign n554 = ( i_37_ ) | ( n580 ) ;
 assign n553 = ( i_38_ ) | ( i_40_ ) ;
 assign n552 = ( n554  &  i_37_ ) | ( n554  &  n553 ) ;
 assign n557 = ( (~ i_40_)  &  n548 ) | ( n315  &  n548 ) | ( n548  &  n862 ) ;
 assign n558 = ( n804  &  n539 ) | ( n836  &  n539 ) | ( n804  &  n1024 ) | ( n836  &  n1024 ) ;
 assign n556 = ( (~ i_33_) ) | ( n1023 ) ;
 assign n555 = ( n557  &  n558  &  n552 ) | ( n557  &  n558  &  n556 ) ;
 assign n562 = ( (~ i_40_) ) | ( n220 ) | ( n455 ) ;
 assign n560 = ( n1025  &  n1052 ) ;
 assign n561 = ( (~ i_36_) ) | ( n1038 ) ;
 assign n559 = ( n562  &  n560 ) | ( n562  &  n561 ) ;
 assign n566 = ( (~ i_3_)  &  (~ i_4_)  &  (~ n550) ) ;
 assign n563 = ( n566  &  (~ n825) ) | ( i_39_  &  n566  &  (~ n890) ) ;
 assign n567 = ( (~ i_5_)  &  (~ n563) ) | ( i_36_  &  (~ n563) ) | ( (~ n563)  &  (~ n775) ) ;
 assign n570 = ( i_9_  &  n544 ) | ( i_9_  &  (~ n512)  &  (~ n1079) ) ;
 assign n573 = ( n525  &  n512 ) | ( n312  &  n512 ) | ( n525  &  n773 ) | ( n312  &  n773 ) ;
 assign n574 = ( n163  &  n538 ) | ( n334  &  n538 ) | ( n163  &  n1048 ) | ( n334  &  n1048 ) ;
 assign n575 = ( n534 ) | ( n1116 ) ;
 assign n576 = ( n555  &  n547 ) | ( n730  &  n547 ) | ( n555  &  n1103 ) | ( n730  &  n1103 ) ;
 assign n578 = ( n559  &  n567 ) | ( n559  &  (~ n1017) ) | ( n567  &  n1113 ) | ( (~ n1017)  &  n1113 ) ;
 assign n579 = ( (~ i_11_)  &  n882 ) | ( n598  &  n882 ) | ( n864  &  n882 ) ;
 assign n572 = ( n515  &  (~ n570)  &  n573  &  n574  &  n575  &  n576  &  n578  &  n579 ) ;
 assign n580 = ( i_38_ ) | ( i_39_ ) ;
 assign n581 = ( (~ i_35_) ) | ( n1041 ) ;
 assign n584 = ( (~ i_17_) ) | ( n583 ) ;
 assign n583 = ( i_32_ ) | ( i_31_ ) ;
 assign n582 = ( (~ i_16_)  &  n584 ) | ( n584  &  n583 ) ;
 assign n585 = ( (~ n541)  &  (~ n582) ) | ( (~ n539)  &  (~ n582)  &  (~ n591) ) ;
 assign n591 = ( i_36_ ) | ( n474 ) ;
 assign n590 = ( (~ i_40_)  &  n541 ) | ( n541  &  n539 ) | ( n541  &  n591 ) ;
 assign n594 = ( i_14_ ) | ( n582 ) | ( n590 ) ;
 assign n595 = ( i_15_  &  i_12_ ) | ( n1122  &  i_12_ ) | ( i_15_  &  n1235 ) | ( n1122  &  n1235 ) ;
 assign n593 = ( n474 ) | ( n535 ) ;
 assign n592 = ( n594  &  n595  &  n514 ) | ( n594  &  n595  &  n593 ) ;
 assign n599 = ( n904 ) | ( n312 ) | ( n890 ) ;
 assign n597 = ( i_37_ ) | ( n174 ) ;
 assign n598 = ( n398 ) | ( n1066 ) ;
 assign n596 = ( n599  &  n223 ) | ( n599  &  n597 ) | ( n599  &  n598 ) ;
 assign n602 = ( n1236  &  n154 ) | ( n1236  &  n184 ) | ( n1236  &  n1124 ) ;
 assign n603 = ( n1237  &  n329 ) | ( n1237  &  n890 ) ;
 assign n601 = ( i_15_ ) | ( i_5_ ) | ( i_31_ ) ;
 assign n600 = ( n602  &  n603  &  n240 ) | ( n602  &  n603  &  n601 ) ;
 assign n604 = ( n548  &  n177 ) | ( n548  &  n230 ) ;
 assign n605 = ( i_36_  &  (~ n490)  &  (~ n751)  &  (~ n963) ) ;
 assign n610 = ( (~ i_38_) ) | ( (~ i_40_) ) ;
 assign n609 = ( n487  &  n610 ) | ( n561  &  n610 ) | ( n487  &  (~ n1150) ) | ( n561  &  (~ n1150) ) ;
 assign n614 = ( (~ i_13_)  &  (~ n398) ) ;
 assign n613 = ( (~ n173)  &  (~ n220) ) ;
 assign n612 = ( n614  &  n613 ) | ( (~ n490)  &  n614  &  (~ n1045) ) ;
 assign n617 = ( (~ n1030) ) | ( (~ n1061) ) ;
 assign n615 = ( (~ n271)  &  (~ n1051) ) | ( n617  &  (~ n1051) ) | ( (~ n905)  &  (~ n1051) ) ;
 assign n619 = ( i_31_ ) | ( n398 ) ;
 assign n620 = ( n238 ) | ( n334 ) ;
 assign n618 = ( (~ n612)  &  (~ n615)  &  n619 ) | ( (~ n612)  &  (~ n615)  &  n620 ) ;
 assign n623 = ( (~ n1039)  &  (~ n1124) ) | ( (~ n1039)  &  (~ n1125) ) ;
 assign n627 = ( n605  &  (~ n1103) ) | ( (~ n550)  &  (~ n604)  &  (~ n1103) ) ;
 assign n632 = ( (~ i_32_)  &  n135 ) | ( i_33_  &  n135 ) | ( (~ i_32_)  &  n1235 ) | ( i_33_  &  n1235 ) ;
 assign n633 = ( n312  &  n942 ) | ( n600  &  n942 ) | ( n312  &  (~ n1126) ) | ( n600  &  (~ n1126) ) ;
 assign n634 = ( n365  &  n592 ) | ( n592  &  n601 ) | ( n365  &  (~ n1027) ) | ( n601  &  (~ n1027) ) ;
 assign n635 = ( (~ n623)  &  n1109 ) | ( n162  &  (~ n623)  &  n1117 ) ;
 assign n636 = ( (~ n247)  &  n1238 ) | ( n598  &  n1238 ) | ( n864  &  n1238 ) ;
 assign n637 = ( (~ n627)  &  n1114  &  n1241 ) | ( (~ n627)  &  n1120  &  n1241 ) ;
 assign n631 = ( n596  &  n101  &  n632  &  n633  &  n634  &  n635  &  n636  &  n637 ) ;
 assign n638 = ( n997 ) | ( n964 ) | ( n1074 ) ;
 assign n640 = ( n251  &  n1043 ) ;
 assign n643 = ( (~ i_23_)  &  n1098 ) ;
 assign n646 = ( (~ i_21_) ) | ( (~ i_23_) ) ;
 assign n644 = ( n646  &  (~ n804)  &  (~ n1040) ) ;
 assign n649 = ( (~ n474)  &  (~ n1040) ) ;
 assign n653 = ( i_5_ ) | ( i_29_ ) | ( i_28_ ) ;
 assign n651 = ( i_5_  &  n653 ) | ( n653  &  (~ n1151) ) ;
 assign n656 = ( (~ i_25_) ) | ( n398 ) ;
 assign n654 = ( (~ i_26_)  &  n656 ) | ( n398  &  n656 ) ;
 assign n660 = ( n997 ) | ( n620 ) ;
 assign n658 = ( i_37_ ) | ( n904 ) ;
 assign n659 = ( n389 ) | ( n685 ) ;
 assign n657 = ( n660  &  n426 ) | ( n660  &  n658 ) | ( n660  &  n659 ) ;
 assign n663 = ( (~ i_22_) ) | ( n355 ) ;
 assign n661 = ( n157  &  n663 ) | ( n663  &  (~ n1098) ) | ( n157  &  (~ n1155) ) | ( (~ n1098)  &  (~ n1155) ) ;
 assign n666 = ( n535 ) | ( n928 ) ;
 assign n665 = ( i_34_ ) | ( n1023 ) ;
 assign n664 = ( n666  &  n665 ) | ( n666  &  n164 ) ;
 assign n668 = ( (~ i_38_) ) | ( n237 ) ;
 assign n667 = ( n668  &  n490 ) ;
 assign n670 = ( n1249  &  n904 ) | ( n1249  &  n1040 ) | ( n1249  &  n1109 ) ;
 assign n671 = ( n1250  &  n581 ) | ( n1111  &  n581 ) | ( n1250  &  n804 ) | ( n1111  &  n804 ) ;
 assign n669 = ( n670  &  n671  &  n667 ) | ( n670  &  n671  &  n439 ) ;
 assign n673 = ( n658  &  n942 ) | ( n658  &  n1120 ) | ( n942  &  (~ n1126) ) | ( n1120  &  (~ n1126) ) ;
 assign n674 = ( n669  &  n654 ) | ( n312  &  n654 ) | ( n669  &  n971 ) | ( n312  &  n971 ) ;
 assign n675 = ( n163 ) | ( n928 ) ;
 assign n676 = ( n1251  &  n661 ) | ( n1251  &  n668 ) | ( n1251  &  n659 ) ;
 assign n677 = ( n158 ) | ( n161 ) | ( n356 ) ;
 assign n672 = ( n657  &  n596  &  n673  &  n99  &  n674  &  n675  &  n676  &  n677 ) ;
 assign n680 = ( n678 ) | ( n514 ) | ( n1075 ) ;
 assign n678 = ( n904 ) | ( n944 ) ;
 assign n679 = ( n348 ) | ( n514 ) | ( n451 ) ;
 assign n683 = ( n389 ) | ( n358 ) ;
 assign n682 = ( i_40_ ) | ( n554 ) ;
 assign n681 = ( n683  &  n389 ) | ( n683  &  n682 ) ;
 assign n685 = ( (~ i_24_) ) | ( n398 ) ;
 assign n684 = ( n163  &  n681 ) | ( n173  &  n681 ) | ( n163  &  n685 ) | ( n173  &  n685 ) ;
 assign n687 = ( (~ n251) ) | ( n663 ) | ( n684 ) ;
 assign n689 = ( n898 ) | ( n1067 ) ;
 assign n686 = ( n36  &  (~ n126)  &  n687  &  n689 ) ;
 assign n690 = ( i_23_ ) | ( n162 ) | ( (~ n251) ) | ( n355 ) ;
 assign n691 = ( (~ n221)  &  (~ n324) ) | ( (~ n221)  &  (~ n325) ) ;
 assign n696 = ( (~ n403)  &  n1080 ) ;
 assign n697 = ( (~ n407)  &  n1080 ) ;
 assign n695 = ( (~ n289)  &  n696 ) | ( (~ n289)  &  n697 ) ;
 assign n699 = ( (~ i_23_)  &  n251  &  (~ n357) ) ;
 assign n702 = ( (~ n329)  &  n740 ) ;
 assign n701 = ( n369  &  n702 ) | ( n699  &  n702 ) | ( n702  &  (~ n1134) ) ;
 assign n703 = ( n113  &  (~ n1133) ) | ( (~ n1132)  &  (~ n1133) ) ;
 assign n707 = ( n751 ) | ( n403 ) | ( n1081 ) ;
 assign n709 = ( i_0_  &  i_1_ ) ;
 assign n711 = ( i_3_  &  (~ n341) ) ;
 assign n712 = ( n312 ) | ( n443 ) ;
 assign n713 = ( n712 ) | ( n339 ) | ( n553 ) ;
 assign n715 = ( n473  &  i_37_ ) | ( n1100  &  i_37_ ) | ( n473  &  n804 ) | ( n1100  &  n804 ) ;
 assign n714 = ( n658  &  n554  &  n715 ) ;
 assign n716 = ( n247  &  i_9_ ) | ( n247  &  i_16_ ) ;
 assign n718 = ( i_9_ ) | ( i_16_ ) | ( i_36_ ) | ( (~ i_39_) ) ;
 assign n719 = ( n1037 ) | ( n247 ) ;
 assign n717 = ( n718  &  n719  &  n271 ) | ( n718  &  n719  &  n716 ) ;
 assign n722 = ( (~ i_37_)  &  n1333 ) | ( n730  &  n1333 ) | ( n1020  &  n1333 ) ;
 assign n723 = ( n1255  &  n1256  &  n1066 ) | ( n1255  &  n1256  &  n728 ) ;
 assign n721 = ( i_15_ ) | ( n398 ) ;
 assign n720 = ( n722  &  n723  &  n238 ) | ( n722  &  n723  &  n721 ) ;
 assign n725 = ( i_3_ ) | ( n1074 ) ;
 assign n724 = ( n725 ) | ( i_38_ ) ;
 assign n726 = ( i_11_  &  i_12_ ) ;
 assign n727 = ( (~ i_37_) ) | ( n1038 ) ;
 assign n728 = ( (~ i_0_) ) | ( n398 ) ;
 assign n729 = ( i_38_ ) | ( i_37_ ) ;
 assign n730 = ( i_0_ ) | ( (~ i_5_) ) | ( i_32_ ) ;
 assign n735 = ( (~ n220)  &  (~ n398) ) ;
 assign n733 = ( i_2_ ) | ( i_3_ ) | ( n1054 ) ;
 assign n731 = ( (~ n724)  &  n735 ) | ( (~ n491)  &  n735  &  n733 ) ;
 assign n736 = ( (~ n997)  &  (~ n1257) ) | ( n237  &  (~ n944)  &  (~ n997) ) ;
 assign n740 = ( i_38_  &  (~ n292) ) ;
 assign n739 = ( (~ n808)  &  (~ n1258) ) | ( i_40_  &  n740  &  (~ n808) ) ;
 assign n742 = ( (~ n665)  &  (~ n1099) ) | ( (~ n665)  &  (~ n1116) ) | ( (~ n665)  &  (~ n1259) ) ;
 assign n746 = ( (~ n312)  &  (~ n1263) ) | ( (~ n312)  &  (~ n1264) ) | ( (~ n312)  &  (~ n1265) ) ;
 assign n751 = ( (~ i_35_) ) | ( n1020 ) ;
 assign n750 = ( (~ n113)  &  n219 ) | ( (~ n113)  &  n556 ) | ( n219  &  n751 ) | ( n556  &  n751 ) ;
 assign n752 = ( (~ n827)  &  (~ n1271) ) | ( (~ n312)  &  (~ n827)  &  (~ n1146) ) ;
 assign n756 = ( (~ i_5_) ) | ( n841 ) ;
 assign n755 = ( n751  &  n554 ) | ( n834  &  n554 ) | ( n751  &  n836 ) | ( n834  &  n836 ) ;
 assign n754 = ( (~ n752)  &  n756 ) | ( n750  &  (~ n752)  &  n755 ) ;
 assign n760 = ( (~ i_7_)  &  n932 ) ;
 assign n758 = ( n760  &  (~ n1270) ) | ( i_9_  &  (~ n284)  &  n760 ) ;
 assign n762 = ( i_7_ ) | ( (~ i_9_) ) | ( (~ i_11_) ) ;
 assign n761 = ( (~ i_15_)  &  (~ n758) ) | ( (~ n758)  &  n762 ) | ( (~ n758)  &  (~ n932) ) ;
 assign n765 = ( (~ i_31_)  &  (~ i_37_)  &  (~ n284)  &  (~ n762)  &  (~ n1097) ) ;
 assign n770 = ( n174  &  n244  &  n440  &  (~ n1079)  &  n1100 ) ;
 assign n768 = ( (~ i_33_) ) | ( n665 ) | ( n770 ) ;
 assign n771 = ( (~ i_35_)  &  (~ n164) ) | ( i_35_  &  (~ n804) ) | ( (~ n164)  &  (~ n804) ) ;
 assign n772 = ( i_33_  &  (~ n665) ) ;
 assign n773 = ( (~ i_16_) ) | ( (~ i_17_) ) ;
 assign n774 = ( (~ i_9_)  &  (~ n796) ) ;
 assign n775 = ( (~ i_15_) ) | ( n476 ) ;
 assign n784 = ( i_38_ ) | ( n904 ) ;
 assign n783 = ( n668  &  n784 ) | ( n581  &  n784 ) | ( n668  &  n443 ) | ( n581  &  n443 ) ;
 assign n786 = ( (~ i_36_) ) | ( n729 ) ;
 assign n785 = ( n220  &  i_35_ ) | ( n220  &  n786 ) | ( n220  &  n387 ) ;
 assign n789 = ( i_6_ ) | ( (~ i_34_) ) | ( n535 ) | ( n668 ) ;
 assign n787 = ( (~ i_32_)  &  n789  &  (~ n1334) ) | ( n785  &  n789  &  (~ n1334) ) ;
 assign n792 = ( n1272  &  n561 ) | ( n1272  &  n1100 ) ;
 assign n793 = ( n1025  &  n727 ) | ( n1066  &  n727 ) | ( n1025  &  n804 ) | ( n1066  &  n804 ) ;
 assign n791 = ( n792  &  n793  &  n552 ) | ( n792  &  n793  &  n220 ) ;
 assign n794 = ( i_0_ ) | ( n791 ) | ( n294 ) ;
 assign n796 = ( (~ i_5_) ) | ( i_7_ ) ;
 assign n797 = ( i_17_ ) | ( n398 ) ;
 assign n795 = ( n398  &  n796 ) | ( (~ n774)  &  n796 ) | ( n398  &  n797 ) | ( (~ n774)  &  n797 ) ;
 assign n799 = ( i_16_  &  (~ n774) ) | ( i_16_  &  n797 ) | ( (~ n774)  &  n795 ) | ( n797  &  n795 ) ;
 assign n800 = ( (~ n289)  &  (~ n397) ) | ( (~ n397)  &  (~ n665)  &  (~ n1024) ) ;
 assign n804 = ( (~ i_38_) ) | ( n329 ) ;
 assign n803 = ( n238  &  (~ n800) ) | ( n312  &  (~ n800) ) | ( (~ n800)  &  n804 ) ;
 assign n807 = ( n462 ) | ( n237 ) ;
 assign n808 = ( i_35_ ) | ( n398 ) ;
 assign n806 = ( n807  &  (~ n982) ) | ( n808  &  (~ n982) ) ;
 assign n810 = ( n289  &  n1029 ) ;
 assign n809 = ( n810 ) | ( i_14_ ) | ( n397 ) ;
 assign n811 = ( i_9_  &  (~ n809) ) | ( i_9_  &  (~ i_12_)  &  (~ n803) ) ;
 assign n818 = ( (~ i_16_) ) | ( n400 ) | ( (~ n476) ) | ( n810 ) ;
 assign n816 = ( n665 ) | ( n1099 ) ;
 assign n815 = ( n517  &  (~ n811)  &  n818 ) | ( (~ n811)  &  n818  &  n816 ) ;
 assign n820 = ( n1040 ) | ( n490 ) ;
 assign n821 = ( n237 ) | ( (~ n740) ) ;
 assign n822 = ( n904  &  n440 ) | ( n297  &  n440 ) | ( n904  &  n238 ) | ( n297  &  n238 ) ;
 assign n823 = ( (~ i_13_)  &  n479 ) | ( i_36_  &  n479 ) | ( n479  &  n784 ) ;
 assign n819 = ( n620  &  n239  &  n820  &  n821  &  n822  &  n823 ) ;
 assign n825 = ( n904 ) | ( n444 ) ;
 assign n824 = ( n825  &  i_40_ ) | ( n825  &  n591 ) ;
 assign n827 = ( i_0_ ) | ( n796 ) ;
 assign n828 = ( i_7_ ) | ( n247 ) ;
 assign n826 = ( n824  &  n819 ) | ( n827  &  n819 ) | ( n824  &  n828 ) | ( n827  &  n828 ) ;
 assign n830 = ( n1037  &  n915  &  n921 ) ;
 assign n829 = ( n830  &  i_36_ ) | ( n830  &  n244 ) ;
 assign n832 = ( (~ i_31_) ) | ( n841 ) ;
 assign n831 = ( n829  &  n830 ) | ( n832  &  n830 ) | ( n829  &  n756 ) | ( n832  &  n756 ) ;
 assign n834 = ( (~ i_40_) ) | ( n1083 ) ;
 assign n833 = ( (~ i_39_)  &  n234  &  n834 ) | ( n230  &  n234  &  n834 ) ;
 assign n837 = ( n1276  &  n541  &  n833 ) | ( n1276  &  n541  &  n539 ) ;
 assign n836 = ( i_36_ ) | ( n1020 ) ;
 assign n835 = ( n750  &  n837  &  n560 ) | ( n750  &  n837  &  n836 ) ;
 assign n838 = ( (~ i_9_)  &  (~ i_13_) ) | ( (~ i_13_)  &  (~ n113) ) | ( (~ i_9_)  &  n834 ) | ( (~ n113)  &  n834 ) ;
 assign n841 = ( i_7_ ) | ( i_32_ ) ;
 assign n840 = ( n838  &  n835 ) | ( n309  &  n835 ) | ( n838  &  n841 ) | ( n309  &  n841 ) ;
 assign n843 = ( i_7_ ) | ( (~ i_9_) ) | ( i_11_ ) | ( n803 ) ;
 assign n844 = ( n826  &  i_7_ ) | ( n312  &  i_7_ ) | ( n826  &  n815 ) | ( n312  &  n815 ) ;
 assign n845 = ( n806 ) | ( n828 ) ;
 assign n846 = ( i_15_  &  n831 ) | ( n840  &  n831 ) | ( i_15_  &  n539 ) | ( n840  &  n539 ) ;
 assign n847 = ( n1277  &  n1278  &  n799 ) | ( n1277  &  n1278  &  n665 ) ;
 assign n842 = ( n754  &  n843  &  n844  &  n845  &  n846  &  n847 ) ;
 assign n849 = ( i_15_  &  (~ n773) ) ;
 assign n848 = ( (~ i_5_)  &  i_12_  &  n849 ) ;
 assign n850 = ( (~ i_14_)  &  n848 ) | ( (~ i_14_)  &  n167  &  (~ n860) ) ;
 assign n853 = ( (~ n142)  &  (~ n239) ) | ( (~ n146)  &  (~ n239) ) | ( (~ n239)  &  n850 ) ;
 assign n856 = ( n1282  &  n1109 ) | ( n1282  &  n1280  &  n236 ) ;
 assign n857 = ( n439  &  (~ n853) ) | ( n237  &  n334  &  (~ n853) ) ;
 assign n858 = ( n1249  &  n581 ) | ( n1249  &  n329  &  n440 ) ;
 assign n855 = ( n856  &  n436  &  n857  &  n858 ) ;
 assign n860 = ( (~ i_15_) ) | ( n1079 ) ;
 assign n859 = ( n426  &  n860 ) | ( n773  &  n860 ) | ( n426  &  (~ n1155) ) | ( n773  &  (~ n1155) ) ;
 assign n862 = ( (~ i_36_) ) | ( n1020 ) ;
 assign n863 = ( i_11_ ) | ( (~ i_12_) ) ;
 assign n864 = ( (~ i_40_) ) | ( n1061 ) ;
 assign n861 = ( n862 ) | ( n863 ) | ( n864 ) ;
 assign n865 = ( i_37_  &  (~ n617) ) | ( (~ i_40_)  &  (~ n617) ) | ( (~ n174)  &  (~ n617) ) ;
 assign n871 = ( n614  &  n1119 ) ;
 assign n868 = ( n871  &  (~ n1279) ) | ( (~ n665)  &  (~ n865)  &  n871 ) ;
 assign n872 = ( (~ n365)  &  (~ n1109) ) | ( (~ n806)  &  (~ n1109) ) | ( (~ n1053)  &  (~ n1109) ) ;
 assign n878 = ( (~ n539)  &  (~ n821) ) ;
 assign n877 = ( (~ i_32_)  &  (~ n861) ) | ( (~ i_32_)  &  (~ n859)  &  n878 ) ;
 assign n882 = ( n475 ) | ( n312 ) | ( n350 ) ;
 assign n883 = ( n1283  &  n654 ) | ( n1283  &  n729 ) | ( n1283  &  n561 ) ;
 assign n884 = ( (~ n1030)  &  n1284 ) | ( n1097  &  n1284 ) | ( n1110  &  n1284 ) ;
 assign n885 = ( n855  &  n1025 ) | ( n312  &  n1025 ) | ( n855  &  n1120 ) | ( n312  &  n1120 ) ;
 assign n886 = ( (~ n872)  &  (~ n1126) ) | ( n487  &  (~ n872)  &  n1147 ) ;
 assign n881 = ( n52  &  n657  &  (~ n877)  &  n882  &  n883  &  n884  &  n885  &  n886 ) ;
 assign n889 = ( (~ i_36_) ) | ( n491 ) ;
 assign n890 = ( (~ i_38_) ) | ( n1041 ) ;
 assign n888 = ( (~ i_40_)  &  n237 ) | ( n237  &  n889 ) | ( (~ i_40_)  &  n890 ) | ( n889  &  n890 ) ;
 assign n892 = ( n237 ) | ( n177 ) | ( n1101 ) ;
 assign n891 = ( n892  &  n888 ) | ( n892  &  n751 ) ;
 assign n895 = ( (~ i_38_) ) | ( n712 ) ;
 assign n894 = ( n997 ) | ( n238 ) ;
 assign n893 = ( n895  &  n894 ) | ( n895  &  n580  &  n553 ) ;
 assign n897 = ( i_40_ ) | ( n597 ) ;
 assign n896 = ( n864  &  n897 ) ;
 assign n899 = ( n896  &  n970 ) | ( n1127  &  n970 ) | ( n896  &  n1114 ) | ( n1127  &  n1114 ) ;
 assign n900 = ( n1287  &  n462 ) | ( n1287  &  n387 ) | ( n1287  &  n1069 ) ;
 assign n898 = ( n1042 ) | ( n561 ) ;
 assign n902 = ( (~ i_15_) ) | ( i_40_ ) | ( (~ n726) ) | ( n944 ) ;
 assign n901 = ( n593  &  n902 ) ;
 assign n905 = ( i_37_ ) | ( n237 ) ;
 assign n904 = ( i_39_ ) | ( (~ i_40_) ) ;
 assign n903 = ( (~ i_37_)  &  n244  &  n905 ) | ( n244  &  n905  &  n904 ) ;
 assign n906 = ( n223  &  i_11_ ) | ( n244  &  i_11_ ) | ( n223  &  n271 ) | ( n244  &  n271 ) ;
 assign n907 = ( (~ n315)  &  (~ n1042) ) | ( (~ n1042)  &  (~ n1088) ) ;
 assign n910 = ( (~ n251) ) | ( n685 ) | ( (~ n1043) ) ;
 assign n909 = ( (~ n907)  &  n910 ) | ( n491  &  n610  &  (~ n907) ) ;
 assign n913 = ( (~ i_37_) ) | ( (~ i_39_) ) ;
 assign n912 = ( n913  &  n658  &  n804  &  n784 ) ;
 assign n916 = ( (~ i_40_) ) | ( n1037 ) ;
 assign n915 = ( i_36_ ) | ( n174 ) ;
 assign n914 = ( n916  &  n230  &  i_40_ ) | ( n916  &  n230  &  n915 ) ;
 assign n917 = ( (~ i_7_)  &  (~ n476)  &  n849 ) ;
 assign n919 = ( n201  &  (~ n251) ) | ( n204  &  (~ n251) ) | ( n201  &  n406 ) | ( n204  &  n406 ) ;
 assign n923 = ( n1092 ) | ( n963 ) | ( n312 ) | ( n964 ) ;
 assign n921 = ( n1101  &  n230 ) ;
 assign n922 = ( i_31_ ) | ( n539 ) ;
 assign n920 = ( n923  &  n921 ) | ( n923  &  n294 ) | ( n923  &  n922 ) ;
 assign n926 = ( i_37_ ) | ( n1065 ) ;
 assign n924 = ( (~ i_38_)  &  n490 ) | ( n330  &  n490 ) | ( (~ i_38_)  &  n926 ) | ( n330  &  n926 ) ;
 assign n928 = ( i_38_ ) | ( n329 ) ;
 assign n927 = ( n928  &  i_39_ ) | ( n928  &  i_37_ ) ;
 assign n932 = ( (~ i_31_)  &  n772 ) ;
 assign n929 = ( (~ n164)  &  (~ n375)  &  n932 ) | ( (~ n375)  &  n932  &  (~ n1067) ) ;
 assign n933 = ( (~ n174)  &  (~ n965) ) | ( i_37_  &  (~ n329)  &  (~ n965) ) ;
 assign n936 = ( (~ i_36_)  &  n1335 ) | ( n906  &  n1335 ) | ( n1062  &  n1335 ) ;
 assign n937 = ( n1303  &  n658 ) | ( n1303  &  n1058 ) ;
 assign n938 = ( n969  &  n1020 ) | ( n1020  &  n1100 ) | ( n969  &  (~ n1291) ) | ( n1100  &  (~ n1291) ) ;
 assign n939 = ( n1301  &  n1302  &  n920 ) | ( n1301  &  n1302  &  n387 ) ;
 assign n940 = ( (~ n64)  &  (~ n929)  &  (~ n933)  &  n972  &  n1148  &  n1294  &  n1296  &  n1297 ) ;
 assign n935 = ( n936  &  n195  &  n937  &  n938  &  n939  &  n940 ) ;
 assign n942 = ( n1052  &  n1024 ) ;
 assign n941 = ( n942  &  n682 ) ;
 assign n944 = ( (~ i_38_) ) | ( n1023 ) ;
 assign n943 = ( (~ i_39_)  &  n239 ) | ( n239  &  n944 ) ;
 assign n945 = ( n296  &  n943  &  n238 ) | ( n296  &  n943  &  n244 ) ;
 assign n948 = ( (~ i_12_) ) | ( n456 ) ;
 assign n946 = ( (~ n464)  &  n948 ) ;
 assign n949 = ( n593  &  n329 ) | ( n593  &  n944 ) ;
 assign n951 = ( (~ i_15_) ) | ( i_17_ ) | ( n943 ) | ( n946 ) ;
 assign n952 = ( (~ i_15_) ) | ( i_16_ ) | ( n945 ) | ( n946 ) ;
 assign n950 = ( n951  &  n952  &  n949 ) | ( n951  &  n952  &  n456 ) ;
 assign n953 = ( n889 ) | ( n751 ) | ( n428 ) | ( i_40_ ) ;
 assign n957 = ( (~ i_5_)  &  (~ n1082) ) | ( (~ i_5_)  &  (~ n329)  &  (~ n462) ) ;
 assign n954 = ( (~ i_28_)  &  i_30_  &  (~ i_31_)  &  n1017 ) ;
 assign n963 = ( i_2_ ) | ( (~ n709) ) ;
 assign n964 = ( i_3_ ) | ( (~ i_4_) ) | ( i_7_ ) ;
 assign n965 = ( n1042 ) | ( n220 ) ;
 assign n968 = ( (~ n309)  &  n566 ) ;
 assign n966 = ( n968  &  (~ n1146) ) | ( (~ n174)  &  n968  &  (~ n1111) ) ;
 assign n969 = ( (~ i_40_)  &  n970 ) | ( i_40_  &  n1127 ) | ( n970  &  n1127 ) ;
 assign n970 = ( n1042 ) | ( n1066 ) ;
 assign n971 = ( n561 ) | ( n554 ) ;
 assign n972 = ( n965 ) | ( n864 ) ;
 assign n973 = ( (~ n204)  &  (~ n401)  &  (~ n582) ) ;
 assign n975 = ( i_28_ ) | ( n294 ) ;
 assign n976 = ( i_31_ ) | ( n808 ) | ( n1082 ) ;
 assign n980 = ( (~ n541) ) | ( n878 ) ;
 assign n977 = ( n973  &  n980 ) | ( (~ n402)  &  (~ n584)  &  n980 ) ;
 assign n982 = ( (~ n312)  &  n649 ) ;
 assign n981 = ( i_25_  &  n982  &  i_23_  &  i_24_ ) ;
 assign n984 = ( (~ n1035)  &  n1094  &  n1276 ) ;
 assign n985 = ( (~ i_24_) ) | ( i_32_ ) ;
 assign n983 = ( (~ i_25_) ) | ( (~ n251) ) | ( n984 ) | ( n985 ) | ( (~ n1043) ) ;
 assign n987 = ( n251  &  (~ n1313) ) | ( (~ n161)  &  n251  &  n982 ) ;
 assign n990 = ( i_9_ ) | ( n294 ) ;
 assign n989 = ( n202 ) | ( n985 ) | ( n990 ) | ( (~ n1035) ) ;
 assign n993 = ( n1030 ) | ( n389 ) ;
 assign n992 = ( (~ i_40_) ) | ( n200 ) | ( n204 ) | ( n685 ) | ( n993 ) ;
 assign n995 = ( i_12_ ) | ( i_17_ ) | ( n403 ) | ( n1106 ) | ( n922 ) ;
 assign n994 = ( (~ i_21_)  &  n995 ) | ( (~ n251)  &  n995 ) | ( n357  &  n995 ) ;
 assign n997 = ( (~ i_34_) ) | ( n398 ) ;
 assign n996 = ( n237 ) | ( n997 ) | ( n297 ) ;
 assign n998 = ( (~ i_18_)  &  (~ n162)  &  (~ n320) ) | ( (~ i_18_)  &  (~ n320)  &  n982 ) ;
 assign n1001 = ( n251  &  n613  &  (~ n1105) ) | ( n251  &  (~ n681)  &  (~ n1105) ) ;
 assign n1004 = ( (~ n976)  &  (~ n1075) ) | ( (~ n348)  &  (~ n451)  &  (~ n976) ) ;
 assign n1008 = ( n643  &  (~ n989) ) | ( n643  &  (~ n992) ) ;
 assign n1012 = ( n302  &  n1328  &  n329 ) | ( n302  &  n1328  &  n1148 ) ;
 assign n1013 = ( n1327  &  n1325  &  n784 ) | ( n1327  &  n1325  &  n1096 ) ;
 assign n1014 = ( n996  &  (~ n1004)  &  n1323 ) | ( (~ n1004)  &  n1049  &  n1323 ) ;
 assign n1015 = ( n1321  &  n1319  &  n162 ) | ( n1321  &  n1319  &  n323 ) ;
 assign n1016 = ( (~ n5)  &  (~ n117)  &  (~ n126)  &  n689  &  (~ n998)  &  n1140  &  n1277  &  n1318 ) ;
 assign n1011 = ( n45  &  n378  &  n90  &  n1012  &  n1013  &  n1014  &  n1015  &  n1016 ) ;
 assign n1017 = ( (~ i_32_)  &  (~ n539) ) ;
 assign n1019 = ( i_5_ ) | ( n284 ) ;
 assign n1020 = ( (~ i_33_) ) | ( i_34_ ) ;
 assign n1021 = ( i_30_ ) | ( n583 ) ;
 assign n1022 = ( n1021 ) | ( n539 ) ;
 assign n1023 = ( i_36_ ) | ( i_35_ ) ;
 assign n1024 = ( i_37_ ) | ( n474 ) ;
 assign n1025 = ( (~ i_40_) ) | ( n1024 ) ;
 assign n1027 = ( (~ i_5_)  &  i_9_ ) ;
 assign n1029 = ( n1025 ) | ( n665 ) ;
 assign n1030 = ( (~ i_37_) ) | ( n580 ) ;
 assign n1032 = ( n439 ) | ( n784 ) ;
 assign n1035 = ( (~ n479)  &  (~ n751) ) ;
 assign n1036 = ( (~ i_23_) ) | ( n985 ) ;
 assign n1037 = ( i_36_ ) | ( n440 ) ;
 assign n1038 = ( i_34_ ) | ( (~ i_35_) ) ;
 assign n1039 = ( (~ i_21_) ) | ( n184 ) | ( n312 ) | ( n426 ) ;
 assign n1040 = ( (~ i_35_) ) | ( n292 ) ;
 assign n1041 = ( (~ i_36_) ) | ( i_37_ ) ;
 assign n1042 = ( i_7_ ) | ( n398 ) ;
 assign n1043 = ( n170  &  i_21_ ) ;
 assign n1044 = ( (~ i_15_) ) | ( i_32_ ) ;
 assign n1045 = ( i_37_ ) | ( n1038 ) ;
 assign n1046 = ( (~ i_37_) ) | ( n440 ) ;
 assign n1047 = ( n177 ) | ( n807 ) ;
 assign n1048 = ( i_15_ ) | ( n583 ) ;
 assign n1049 = ( (~ i_13_) ) | ( n294 ) ;
 assign n1050 = ( n1049 ) | ( n721 ) ;
 assign n1051 = ( n665 ) | ( n619 ) ;
 assign n1052 = ( (~ i_40_) ) | ( n1030 ) ;
 assign n1053 = ( n271 ) | ( n439 ) | ( n312 ) ;
 assign n1054 = ( i_4_ ) | ( i_1_ ) ;
 assign n1056 = ( (~ i_13_) ) | ( n367 ) | ( n514 ) ;
 assign n1057 = ( i_32_ ) | ( n751 ) | ( n367 ) ;
 assign n1058 = ( i_13_ ) | ( n1057 ) ;
 assign n1059 = ( i_13_ ) | ( n294 ) | ( n721 ) ;
 assign n1060 = ( n539 ) | ( n1048 ) | ( n1049 ) ;
 assign n1061 = ( i_37_ ) | ( n440 ) ;
 assign n1062 = ( i_7_ ) | ( (~ n1017) ) ;
 assign n1064 = ( n223 ) | ( n1062 ) | ( n890 ) ;
 assign n1065 = ( i_35_ ) | ( (~ i_36_) ) ;
 assign n1066 = ( i_34_ ) | ( n1065 ) ;
 assign n1067 = ( i_40_ ) | ( n1046 ) ;
 assign n1068 = ( n177 ) | ( n841 ) ;
 assign n1069 = ( n733 ) | ( n1068 ) ;
 assign n1073 = ( (~ i_36_) ) | ( (~ i_37_) ) ;
 assign n1074 = ( (~ i_0_) ) | ( i_1_ ) | ( (~ i_2_) ) ;
 assign n1075 = ( (~ i_29_) ) | ( (~ i_30_) ) | ( n975 ) ;
 assign n1076 = ( i_16_ ) | ( n619 ) | ( n990 ) ;
 assign n1077 = ( n284 ) | ( n1076 ) ;
 assign n1078 = ( i_17_ ) | ( n990 ) ;
 assign n1079 = ( (~ i_16_)  &  (~ i_17_) ) ;
 assign n1080 = ( i_15_  &  (~ n619)  &  n1079 ) ;
 assign n1081 = ( i_22_ ) | ( n1044 ) ;
 assign n1082 = ( (~ i_40_) ) | ( n915 ) ;
 assign n1083 = ( i_36_ ) | ( n580 ) ;
 assign n1084 = ( i_32_ ) | ( n355 ) ;
 assign n1085 = ( n473 ) | ( n965 ) ;
 assign n1086 = ( (~ n223) ) | ( n309 ) | ( n926 ) ;
 assign n1088 = ( (~ i_37_) ) | ( n553 ) ;
 assign n1089 = ( i_18_ ) | ( n990 ) | ( n322 ) ;
 assign n1091 = ( n711 ) | ( n133 ) ;
 assign n1092 = ( (~ i_35_) ) | ( n491 ) ;
 assign n1093 = ( (~ i_38_) ) | ( n1065 ) ;
 assign n1094 = ( n751 ) | ( n821 ) ;
 assign n1095 = ( i_32_ ) | ( n184 ) ;
 assign n1096 = ( n389 ) | ( n1050 ) ;
 assign n1097 = ( i_36_ ) | ( n539 ) ;
 assign n1098 = ( (~ i_21_)  &  i_22_ ) ;
 assign n1099 = ( (~ i_31_) ) | ( n398 ) ;
 assign n1100 = ( (~ i_37_) ) | ( (~ i_38_) ) ;
 assign n1101 = ( i_36_ ) | ( n1100 ) ;
 assign n1103 = ( i_3_ ) | ( (~ i_4_) ) | ( i_32_ ) ;
 assign n1104 = ( n398 ) | ( n389 ) | ( i_24_ ) | ( n426 ) ;
 assign n1105 = ( (~ i_15_) ) | ( n398 ) ;
 assign n1106 = ( i_16_ ) | ( n1044 ) ;
 assign n1107 = ( i_22_ ) | ( n398 ) ;
 assign n1108 = ( n1074 ) | ( n1103 ) | ( i_40_ ) | ( n177 ) ;
 assign n1109 = ( i_15_ ) | ( i_5_ ) | ( i_13_ ) ;
 assign n1110 = ( i_5_ ) | ( (~ i_31_) ) | ( i_32_ ) ;
 assign n1111 = ( (~ i_37_) ) | ( n1065 ) ;
 assign n1113 = ( (~ i_6_) ) | ( n398 ) ;
 assign n1114 = ( i_40_ ) | ( n1030 ) ;
 assign n1116 = ( (~ i_5_) ) | ( n398 ) ;
 assign n1117 = ( (~ n982)  &  n996 ) ;
 assign n1119 = ( (~ i_5_)  &  (~ n247) ) ;
 assign n1120 = ( (~ n735) ) | ( n733 ) ;
 assign n1122 = ( i_34_ ) | ( (~ n545) ) | ( n619 ) ;
 assign n1124 = ( n237 ) | ( n1040 ) ;
 assign n1125 = ( (~ i_35_) ) | ( n387 ) | ( n729 ) ;
 assign n1126 = ( (~ n389)  &  n871 ) ;
 assign n1127 = ( n389 ) | ( n1042 ) ;
 assign n1128 = ( (~ i_15_) ) | ( (~ i_24_) ) | ( n312 ) ;
 assign n1129 = ( i_22_ ) | ( (~ n251) ) | ( n1128 ) ;
 assign n1130 = ( n230 ) | ( n387 ) ;
 assign n1131 = ( n389 ) | ( n1052 ) ;
 assign n1132 = ( n1130  &  n479 ) ;
 assign n1133 = ( n751 ) | ( n407 ) | ( n1081 ) ;
 assign n1134 = ( n751 ) | ( n407 ) | ( n1084 ) ;
 assign n1139 = ( n1130  &  n1132 ) | ( n1134  &  n1132 ) | ( n1130  &  n707 ) | ( n1134  &  n707 ) ;
 assign n1140 = ( n665 ) | ( n244 ) | ( i_37_ ) | ( n288 ) ;
 assign n1143 = ( n1252  &  n321 ) | ( n1252  &  n1131 ) ;
 assign n1146 = ( n668 ) | ( n926 ) ;
 assign n1147 = ( n554  &  n1024 ) ;
 assign n1148 = ( n363 ) | ( n1101 ) ;
 assign n1149 = ( (~ i_38_)  &  n238 ) | ( i_38_  &  n535 ) | ( n238  &  n535 ) ;
 assign n1150 = ( i_37_  &  (~ n220) ) | ( (~ i_37_)  &  (~ n561) ) | ( (~ n220)  &  (~ n561) ) ;
 assign n1151 = ( i_28_  &  i_29_ ) | ( i_28_  &  i_30_ ) | ( i_29_  &  (~ i_30_) ) ;
 assign n1152 = ( i_5_ ) | ( n863 ) ;
 assign n1153 = ( i_5_ ) | ( (~ i_11_) ) | ( i_12_ ) ;
 assign n1155 = ( n167 ) | ( n171 ) ;
 assign n1154 = ( n1035  &  n169 ) | ( n1035  &  n250  &  n1155 ) ;
 assign n1157 = ( n172  &  n997 ) | ( n894  &  n997 ) | ( n172  &  n678 ) | ( n894  &  n678 ) ;
 assign n1158 = ( n729  &  n389 ) | ( n561  &  n389 ) | ( n729  &  n1046 ) | ( n561  &  n1046 ) ;
 assign n1160 = ( n163 ) | ( n173 ) | ( (~ n640) ) ;
 assign n1162 = ( n1051 ) | ( n295 ) | ( n1052 ) ;
 assign n1161 = ( i_31_  &  n1162 ) | ( n214  &  n1162 ) | ( (~ n1017)  &  n1162 ) ;
 assign n1163 = ( n1161  &  n203 ) | ( n1161  &  n161 ) | ( n1161  &  n1053 ) ;
 assign n1165 = ( (~ n259)  &  n1056 ) | ( n240  &  (~ n259)  &  n620 ) ;
 assign n1167 = ( n387  &  n970 ) | ( n1064  &  n970 ) | ( n387  &  n1067 ) | ( n1064  &  n1067 ) ;
 assign n1168 = ( n1167  &  n658 ) | ( n1167  &  n379 ) ;
 assign n1169 = ( (~ n298)  &  n1056 ) | ( n239  &  n296  &  (~ n298) ) ;
 assign n1172 = ( n1133  &  n707 ) ;
 assign n1173 = ( n1054  &  i_0_ ) ;
 assign n1175 = ( n367 ) | ( n1061 ) | ( n583 ) | ( n556 ) ;
 assign n1174 = ( n1175  &  n389 ) | ( n1175  &  n554 ) | ( n1175  &  n1059 ) ;
 assign n1177 = ( n751 ) | ( n841 ) | ( n337 ) | ( n786 ) ;
 assign n1176 = ( n1177  &  n362  &  n364  &  n26  &  n680  &  n197 ) ;
 assign n1179 = ( n1022 ) | ( n207 ) | ( n1082 ) ;
 assign n1178 = ( n1179  &  n904 ) | ( n1179  &  n230 ) | ( n1179  &  n1058 ) ;
 assign n1180 = ( n351  &  n174 ) | ( n619  &  n174 ) | ( n351  &  n1086 ) | ( n619  &  n1086 ) ;
 assign n1181 = ( n1180  &  n965 ) | ( n1180  &  n905 ) ;
 assign n1182 = ( n333  &  n328 ) | ( n238  &  n328 ) | ( n333  &  n1042 ) | ( n238  &  n1042 ) ;
 assign n1183 = ( n350  &  n1181  &  n1182 ) | ( n1181  &  n1182  &  (~ n1342) ) ;
 assign n1184 = ( n1172  &  n321 ) | ( n235  &  n321 ) | ( n1172  &  n993 ) | ( n235  &  n993 ) ;
 assign n1187 = ( i_40_  &  n313 ) | ( (~ i_40_)  &  n342 ) | ( n313  &  n342 ) ;
 assign n1185 = ( (~ n125)  &  n302  &  n1187 ) | ( n302  &  n1083  &  n1187 ) ;
 assign n1188 = ( n1184  &  n1185  &  n1052 ) | ( n1184  &  n1185  &  n970 ) ;
 assign n1189 = ( (~ i_39_)  &  (~ n237) ) | ( (~ n237)  &  n297 ) | ( (~ i_39_)  &  n944 ) | ( n297  &  n944 ) ;
 assign n1190 = ( (~ n397)  &  (~ n401) ) | ( (~ i_14_)  &  (~ n284)  &  (~ n397) ) ;
 assign n1192 = ( n665 ) | ( n1059 ) | ( n1061 ) ;
 assign n1191 = ( n1192  &  n462 ) | ( n1192  &  n379 ) ;
 assign n1194 = ( n451 ) | ( n975 ) | ( (~ n1017) ) | ( n1082 ) ;
 assign n1195 = ( i_5_ ) | ( n832 ) | ( (~ n1079) ) | ( n1097 ) ;
 assign n1196 = ( n1046 ) | ( n1050 ) | ( n220 ) ;
 assign n1197 = ( i_38_ ) | ( n863 ) | ( n237 ) | ( n1065 ) | ( n309 ) ;
 assign n1199 = ( n392 ) | ( n784 ) | ( n516 ) ;
 assign n1198 = ( n1199  &  n375 ) | ( n1199  &  n398 ) | ( n1199  &  n666 ) ;
 assign n1201 = ( i_36_ ) | ( (~ n773) ) | ( n990 ) | ( (~ n1017) ) ;
 assign n1202 = ( (~ i_23_) ) | ( n203 ) | ( n659 ) | ( (~ n1098) ) ;
 assign n1204 = ( n293  &  n382 ) | ( n816  &  n382 ) | ( n293  &  n367 ) | ( n816  &  n367 ) ;
 assign n1205 = ( n965  &  n164 ) | ( n1067  &  n164 ) | ( n965  &  n314 ) | ( n1067  &  n314 ) ;
 assign n1206 = ( (~ i_32_)  &  (~ n541) ) | ( (~ i_32_)  &  (~ n556)  &  (~ n1025) ) ;
 assign n1210 = ( (~ n143)  &  (~ n289) ) | ( (~ n143)  &  (~ n238)  &  (~ n474) ) ;
 assign n1214 = ( i_12_ ) | ( i_5_ ) | ( n478 ) ;
 assign n1213 = ( n1109  &  n1214 ) | ( n479  &  (~ n702)  &  n1214 ) ;
 assign n1215 = ( (~ n459)  &  (~ n1073) ) | ( i_36_  &  (~ n459)  &  (~ n474) ) ;
 assign n1218 = ( n461  &  n946 ) | ( n948  &  n946 ) | ( n461  &  n232 ) | ( n948  &  n232 ) ;
 assign n1220 = ( n442  &  n441 ) | ( n473  &  n441 ) | ( n442  &  n1111 ) | ( n473  &  n1111 ) ;
 assign n1221 = ( i_14_  &  (~ n445)  &  n1220 ) | ( n438  &  (~ n445)  &  n1220 ) ;
 assign n1223 = ( (~ n188)  &  n439 ) | ( (~ n188)  &  n553 ) | ( n439  &  n581 ) | ( n553  &  n581 ) ;
 assign n1224 = ( (~ n548)  &  (~ n1074) ) | ( (~ n177)  &  (~ n1074)  &  (~ n1083) ) ;
 assign n1229 = ( n541 ) | ( n948 ) | ( i_17_ ) | ( n1044 ) ;
 assign n1228 = ( n1019  &  n1229 ) | ( (~ n1079)  &  n1229 ) | ( (~ n1206)  &  n1229 ) ;
 assign n1230 = ( n1228  &  i_25_ ) | ( n1228  &  n398 ) | ( n1228  &  n971 ) ;
 assign n1231 = ( n428 ) | ( n751 ) | ( n1088 ) ;
 assign n1232 = ( n946  &  n425 ) | ( n492  &  n425 ) | ( n946  &  n489 ) | ( n492  &  n489 ) ;
 assign n1233 = ( n481  &  n292 ) | ( n329  &  n292 ) | ( n481  &  n1108 ) | ( n329  &  n1108 ) ;
 assign n1234 = ( (~ i_5_)  &  n476  &  n980 ) ;
 assign n1235 = ( (~ n585)  &  n1122 ) ;
 assign n1236 = ( n1109 ) | ( n1125 ) ;
 assign n1237 = ( n173  &  n490 ) | ( n443  &  n490 ) | ( n173  &  n1111 ) | ( n443  &  n1111 ) ;
 assign n1238 = ( (~ i_16_)  &  n84 ) | ( n84  &  n584 ) | ( n84  &  (~ n1234) ) ;
 assign n1241 = ( n609  &  n618 ) | ( n618  &  n1113 ) | ( n609  &  (~ n1119) ) | ( n1113  &  (~ n1119) ) ;
 assign n1245 = ( n251  &  n644 ) | ( (~ i_21_)  &  n251  &  (~ n820) ) ;
 assign n1248 = ( i_21_ ) | ( i_23_ ) | ( (~ i_24_) ) | ( n162 ) | ( n203 ) ;
 assign n1247 = ( n23  &  n1128  &  n1248 ) | ( n23  &  (~ n1245)  &  n1248 ) ;
 assign n1249 = ( (~ i_35_) ) | ( i_37_ ) | ( n164 ) ;
 assign n1250 = ( n271  &  n440 ) ;
 assign n1251 = ( n651 ) | ( n664 ) | ( n619 ) ;
 assign n1252 = ( (~ n369)  &  n1029 ) | ( n1029  &  n1130 ) | ( (~ n369)  &  (~ n1342) ) | ( n1130  &  (~ n1342) ) ;
 assign n1254 = ( i_40_ ) | ( n315 ) | ( n1127 ) ;
 assign n1255 = ( i_34_ ) | ( i_35_ ) | ( n1116 ) ;
 assign n1256 = ( n398 ) | ( n727 ) | ( n725 ) ;
 assign n1257 = ( n1250  &  n238 ) | ( n535  &  n238 ) | ( n1250  &  n473 ) | ( n535  &  n473 ) ;
 assign n1258 = ( n1082  &  n786 ) | ( n1082  &  n387 ) ;
 assign n1260 = ( i_9_ ) | ( n398 ) | ( n474 ) ;
 assign n1259 = ( n1260  &  n440 ) | ( n1260  &  n721 ) ;
 assign n1261 = ( (~ i_35_)  &  n271 ) | ( n271  &  n714 ) | ( (~ i_35_)  &  n1065 ) | ( n714  &  n1065 ) ;
 assign n1262 = ( n329  &  n174 ) | ( n1092  &  n174 ) | ( n329  &  n926 ) | ( n1092  &  n926 ) ;
 assign n1263 = ( n1261  &  n1262  &  i_40_ ) | ( n1261  &  n1262  &  n1093 ) ;
 assign n1264 = ( i_38_  &  n439 ) | ( n439  &  n581 ) | ( i_38_  &  (~ n804) ) | ( n581  &  (~ n804) ) ;
 assign n1265 = ( (~ i_39_)  &  (~ n237) ) | ( (~ i_39_)  &  n462 ) | ( (~ n237)  &  n1111 ) | ( n462  &  n1111 ) ;
 assign n1266 = ( (~ i_38_)  &  n717 ) | ( n717  &  n720 ) | ( (~ i_38_)  &  (~ n1017) ) | ( n720  &  (~ n1017) ) ;
 assign n1267 = ( n736 ) | ( n739 ) | ( n742 ) | ( n746 ) | ( (~ n1117) ) | ( (~ n1266) ) ;
 assign n1270 = ( (~ i_16_)  &  n140 ) | ( n140  &  n276 ) ;
 assign n1271 = ( n230  &  n895 ) | ( (~ n237)  &  n895 ) | ( n808  &  n895 ) ;
 assign n1272 = ( i_34_ ) | ( n164 ) | ( n1073 ) ;
 assign n1274 = ( i_0_ ) | ( n490 ) | ( n443 ) ;
 assign n1273 = ( n1274  &  i_6_ ) | ( n1274  &  n783 ) ;
 assign n1276 = ( n751 ) | ( n1130 ) ;
 assign n1277 = ( (~ i_11_) ) | ( n237 ) | ( n786 ) | ( n1062 ) ;
 assign n1278 = ( n358 ) | ( n836 ) | ( n756 ) ;
 assign n1279 = ( n620  &  n535 ) | ( n620  &  n173 ) ;
 assign n1280 = ( n1250  &  n580 ) | ( n238  &  n580 ) | ( n1250  &  n1040 ) | ( n238  &  n1040 ) ;
 assign n1282 = ( n668 ) | ( n1111 ) ;
 assign n1283 = ( i_5_ ) | ( n517 ) | ( n816 ) ;
 assign n1284 = ( n490  &  (~ n868) ) | ( (~ n868)  &  n926 ) | ( (~ n868)  &  n997 ) ;
 assign n1288 = ( (~ i_6_) ) | ( n841 ) | ( n891 ) ;
 assign n1287 = ( n1288  &  n893 ) | ( n1288  &  n964 ) | ( n1288  &  n550 ) ;
 assign n1289 = ( i_14_  &  (~ n140) ) | ( i_14_  &  i_17_  &  (~ n284) ) ;
 assign n1291 = ( n917  &  (~ n1308) ) | ( (~ n762)  &  n1289  &  (~ n1308) ) ;
 assign n1295 = ( n1020 ) | ( n204 ) | ( i_31_ ) | ( n901 ) ;
 assign n1294 = ( n1295  &  n914 ) | ( n1295  &  n919 ) | ( n1295  &  n922 ) ;
 assign n1296 = ( n927  &  n924 ) | ( n1085  &  n924 ) | ( n927  &  n1042 ) | ( n1085  &  n1042 ) ;
 assign n1297 = ( (~ i_40_) ) | ( (~ n968) ) | ( n1093 ) ;
 assign n1301 = ( n904 ) | ( n1045 ) | ( n1059 ) ;
 assign n1302 = ( (~ n640) ) | ( n996 ) ;
 assign n1303 = ( n912  &  n909 ) | ( n970  &  n909 ) | ( n912  &  n389 ) | ( n970  &  n389 ) ;
 assign n1305 = ( (~ n459)  &  (~ n825) ) | ( (~ n237)  &  (~ n459)  &  (~ n890) ) ;
 assign n1309 = ( n486 ) | ( n219 ) | ( n220 ) ;
 assign n1308 = ( n239  &  n350 ) ;
 assign n1307 = ( n514  &  n1309 ) | ( (~ n1079)  &  n1309 ) | ( n1309  &  n1308 ) ;
 assign n1310 = ( n514  &  n539 ) | ( n539  &  n950 ) | ( n514  &  (~ n1305) ) | ( n950  &  (~ n1305) ) ;
 assign n1311 = ( n425  &  n230 ) | ( n941  &  n230 ) | ( n425  &  n1108 ) | ( n941  &  n1108 ) ;
 assign n1312 = ( n1311  &  n712 ) | ( n1311  &  n928 ) ;
 assign n1314 = ( (~ i_22_) ) | ( n173 ) | ( (~ n735) ) ;
 assign n1313 = ( n1314  &  n984 ) | ( n1314  &  n1095 ) ;
 assign n1318 = ( i_25_ ) | ( i_26_ ) | ( n580 ) | ( n581 ) | ( n309 ) ;
 assign n1319 = ( n604  &  (~ n1001) ) | ( n725  &  (~ n1001) ) | ( n841  &  (~ n1001) ) ;
 assign n1321 = ( n238 ) | ( n244 ) | ( n1056 ) ;
 assign n1323 = ( i_40_ ) | ( (~ n740) ) | ( n1060 ) ;
 assign n1324 = ( n314  &  n379 ) | ( n1100  &  n379 ) | ( n314  &  n834 ) | ( n1100  &  n834 ) ;
 assign n1325 = ( (~ n113)  &  (~ n1008)  &  n1324 ) | ( n994  &  (~ n1008)  &  n1324 ) ;
 assign n1327 = ( n1032  &  n910 ) | ( n1129  &  n910 ) | ( n1032  &  n1131 ) | ( n1129  &  n1131 ) ;
 assign n1328 = ( (~ n697)  &  n729 ) | ( n729  &  n1029 ) | ( (~ n697)  &  n1085 ) | ( n1029  &  n1085 ) ;
 assign n1330 = ( i_40_  &  (~ n1191) ) | ( i_40_  &  (~ n554)  &  (~ n1085) ) ;
 assign n1333 = ( i_32_ ) | ( n716 ) | ( n556 ) | ( i_37_ ) ;
 assign n1334 = ( (~ i_34_)  &  (~ n1273) ) | ( i_32_  &  (~ i_34_)  &  n1023 ) ;
 assign n1335 = ( n903 ) | ( n1069 ) | ( i_36_ ) ;
 assign n1336 = ( (~ i_28_)  &  (~ i_29_) ) | ( (~ i_29_)  &  n1022 ) ;
 assign n1337 = ( (~ i_37_)  &  n220 ) | ( (~ i_37_)  &  n553 ) ;
 assign n1342 = ( n696 ) | ( n697 ) ;


endmodule

