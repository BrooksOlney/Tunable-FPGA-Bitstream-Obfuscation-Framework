module ks_sin_qmap_map (sk, ax22x, ax5x, ax3x, ax2x, ax0x, ax1x, ax4x, ax21x, ax19x, ax17x, ax16x, ax13x, ax11x, ax9x, ax7x, ax6x, ax8x, ax10x, ax12x, ax14x, ax15x, ax18x, ax20x, ax23x, sinx0x, sinx1x, sinx2x, sinx3x, sinx4x, sinx5x, sinx6x, sinx7x, sinx8x, sinx9x, sinx10x, sinx11x, sinx12x, sinx13x, sinx14x, sinx15x, sinx16x, sinx17x, sinx18x, sinx19x, sinx20x, sinx21x, sinx22x, sinx23x, sinx24x);

	input ax22x;
	input ax5x;
	input ax3x;
	input ax2x;
	input ax0x;
	input ax1x;
	input ax4x;
	input ax21x;
	input ax19x;
	input ax17x;
	input ax16x;
	input ax13x;
	input ax11x;
	input ax9x;
	input ax7x;
	input ax6x;
	input ax8x;
	input ax10x;
	input ax12x;
	input ax14x;
	input ax15x;
	input ax18x;
	input ax20x;
	input ax23x;
	output sinx0x;
	output sinx1x;
	output sinx2x;
	output sinx3x;
	output sinx4x;
	output sinx5x;
	output sinx6x;
	output sinx7x;
	output sinx8x;
	output sinx9x;
	output sinx10x;
	output sinx11x;
	output sinx12x;
	output sinx13x;
	output sinx14x;
	output sinx15x;
	output sinx16x;
	output sinx17x;
	output sinx18x;
	output sinx19x;
	output sinx20x;
	output sinx21x;
	output sinx22x;
	output sinx23x;
	output sinx24x;

	input [127 : 0] sk /* synthesis noprune */;


	wire g1067, g1107, g1134, g1208, g1231, g1280, g1303, g1339, g1419, g1431, g1441, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10;
	wire g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31;
	wire g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g52;
	wire g53, g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73;
	wire g74, g75, g76, g77, g78, g79, g80, g81, g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93, g94;
	wire g95, g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115;
	wire g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g136;
	wire g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157;
	wire g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178;
	wire g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195, g196, g197, g198, g199;
	wire g200, g201, g202, g203, g204, g205, g206, g207, g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219, g220;
	wire g221, g222, g223, g224, g225, g226, g227, g228, g229, g230, g231, g232, g233, g234, g235, g236, g237, g238, g239, g240, g241;
	wire g242, g243, g244, g245, g246, g247, g248, g249, g250, g251, g252, g253, g254, g255, g256, g257, g258, g259, g260, g261, g262;
	wire g263, g264, g265, g266, g267, g268, g269, g270, g271, g272, g273, g274, g275, g276, g277, g278, g279, g280, g281, g282, g283;
	wire g284, g285, g286, g287, g288, g289, g290, g291, g292, g293, g294, g295, g296, g297, g298, g299, g300, g301, g302, g303, g304;
	wire g305, g306, g307, g308, g309, g310, g311, g312, g313, g314, g315, g316, g317, g318, g319, g320, g321, g322, g323, g324, g325;
	wire g326, g327, g328, g329, g330, g331, g332, g333, g334, g335, g336, g337, g338, g339, g340, g341, g342, g343, g344, g345, g346;
	wire g347, g348, g349, g350, g351, g352, g353, g354, g355, g356, g357, g358, g359, g360, g361, g362, g363, g364, g365, g366, g367;
	wire g368, g369, g370, g371, g372, g373, g374, g375, g376, g377, g378, g379, g380, g381, g382, g383, g384, g385, g386, g387, g388;
	wire g389, g390, g391, g392, g393, g394, g395, g396, g397, g398, g399, g400, g401, g402, g403, g404, g405, g406, g407, g408, g409;
	wire g410, g411, g412, g413, g414, g415, g416, g417, g418, g419, g420, g421, g422, g423, g424, g425, g426, g427, g428, g429, g430;
	wire g431, g432, g433, g434, g435, g436, g437, g438, g439, g440, g441, g442, g443, g444, g445, g446, g447, g448, g449, g450, g451;
	wire g452, g453, g454, g455, g456, g457, g458, g459, g460, g461, g462, g463, g464, g465, g466, g467, g468, g469, g470, g471, g472;
	wire g473, g474, g475, g476, g477, g478, g479, g480, g481, g482, g483, g484, g485, g486, g487, g488, g489, g490, g491, g492, g493;
	wire g494, g495, g496, g497, g498, g499, g500, g501, g502, g503, g504, g505, g506, g507, g508, g509, g510, g511, g512, g513, g514;
	wire g515, g516, g517, g518, g519, g520, g521, g522, g523, g524, g525, g526, g527, g528, g529, g530, g531, g532, g533, g534, g535;
	wire g536, g537, g538, g539, g540, g541, g542, g543, g544, g545, g546, g547, g548, g549, g550, g551, g552, g553, g554, g555, g556;
	wire g557, g558, g559, g560, g561, g562, g563, g564, g565, g566, g567, g568, g569, g570, g571, g572, g573, g574, g575, g576, g577;
	wire g578, g579, g580, g581, g582, g583, g584, g585, g586, g587, g588, g589, g590, g591, g592, g593, g594, g595, g596, g597, g598;
	wire g599, g600, g601, g602, g603, g604, g605, g606, g607, g608, g609, g610, g611, g612, g613, g614, g615, g616, g617, g618, g619;
	wire g620, g621, g622, g623, g624, g625, g626, g627, g628, g629, g630, g631, g632, g633, g634, g635, g636, g637, g638, g639, g640;
	wire g641, g642, g643, g644, g645, g646, g647, g648, g649, g650, g651, g652, g653, g654, g655, g656, g657, g658, g659, g660, g661;
	wire g662, g663, g664, g665, g666, g667, g668, g669, g670, g671, g672, g673, g674, g675, g676, g677, g678, g679, g680, g681, g682;
	wire g683, g684, g685, g686, g687, g688, g689, g690, g691, g692, g693, g694, g695, g696, g697, g698, g699, g700, g701, g702, g703;
	wire g704, g705, g706, g707, g708, g709, g710, g711, g712, g713, g714, g715, g716, g717, g718, g719, g720, g721, g722, g723, g724;
	wire g725, g726, g727, g728, g729, g730, g731, g732, g733, g734, g735, g736, g737, g738, g739, g740, g741, g742, g743, g744, g745;
	wire g746, g747, g748, g749, g750, g751, g752, g753, g754, g755, g756, g757, g758, g759, g760, g761, g762, g763, g764, g765, g766;
	wire g767, g768, g769, g770, g771, g772, g773, g774, g775, g776, g777, g778, g779, g780, g781, g782, g783, g784, g785, g786, g787;
	wire g788, g789, g790, g791, g792, g793, g794, g795, g796, g797, g798, g799, g800, g801, g802, g803, g804, g805, g806, g807, g808;
	wire g809, g810, g811, g812, g813, g814, g815, g816, g817, g818, g819, g820, g821, g822, g823, g824, g825, g826, g827, g828, g829;
	wire g830, g831, g832, g833, g834, g835, g836, g837, g838, g839, g840, g841, g842, g843, g844, g845, g846, g847, g848, g849, g850;
	wire g851, g852, g853, g854, g855, g856, g857, g858, g859, g860, g861, g862, g863, g864, g865, g866, g867, g868, g869, g870, g871;
	wire g872, g873, g874, g875, g876, g877, g878, g879, g880, g881, g882, g883, g884, g885, g886, g887, g888, g889, g890, g891, g892;
	wire g893, g894, g895, g896, g897, g898, g899, g900, g901, g902, g903, g904, g905, g906, g907, g908, g909, g910, g911, g912, g913;
	wire g914, g915, g916, g917, g918, g919, g920, g921, g922, g923, g924, g925, g926, g927, g928, g929, g930, g931, g932, g933, g934;
	wire g935, g936, g937, g938, g939, g940, g941, g942, g943, g944, g945, g946, g947, g948, g949, g950, g951, g952, g953, g954, g955;
	wire g956, g957, g958, g959, g960, g961, g962, g963, g964, g965, g966, g967, g968, g969, g970, g971, g972, g973, g974, g975, g976;
	wire g977, g978, g979, g980, g981, g982, g983, g984, g985, g986, g1447, g987, g988, g989, g990, g991, g992, g993, g994, g995, g996;
	wire g997, g998, g999, g1000, g1001, g1002, g1003, g1004, g1005, g1006, g1007, g1008, g1009, g1010, g1011, g1012, g1013, g1014, g1015, g1016, g1017;
	wire g1018, g1019, g1020, g1021, g1022, g1023, g1024, g1025, g1026, g1027, g1028, g1029, g1030, g1031, g1032, g1033, g1034, g1035, g1036, g1037, g1038;
	wire g1039, g1040, g1041, g1042, g1043, g1044, g1045, g1046, g1047, g1048, g1049, g1050, g1051, g1052, g1053, g1054, g1055, g1056, g1057, g1058, g1059;
	wire g1060, g1061, g1062, g1063, g1064, g1065, g1066, g1068, g1069, g1070, g1071, g1072, g1073, g1074, g1075, g1076, g1077, g1078, g1079, g1080, g1081;
	wire g1082, g1083, g1084, g1085, g1086, g1087, g1088, g1089, g1090, g1091, g1092, g1093, g1094, g1095, g1096, g1097, g1098, g1099, g1100, g1101, g1102;
	wire g1103, g1104, g1105, g1106, g1108, g1109, g1110, g1111, g1112, g1113, g1114, g1115, g1116, g1117, g1118, g1119, g1120, g1121, g1122, g1123, g1124;
	wire g1125, g1126, g1127, g1128, g1129, g1130, g1131, g1132, g1133, g1135, g1136, g1137, g1138, g1139, g1140, g1141, g1142, g1143, g1144, g1145, g1146;
	wire g1147, g1148, g1149, g1150, g1151, g1152, g1153, g1154, g1155, g1156, g1157, g1158, g1160, g1161, g1162, g1163, g1164, g1165, g1166, g1167, g1168;
	wire g1169, g1170, g1171, g1172, g1173, g1174, g1175, g1176, g1177, g1178, g1179, g1180, g1181, g1182, g1183, g1185, g1186, g1187, g1188, g1189, g1190;
	wire g1191, g1192, g1193, g1194, g1195, g1196, g1197, g1198, g1199, g1200, g1201, g1202, g1203, g1204, g1205, g1206, g1207, g1209, g1210, g1211, g1212;
	wire g1213, g1214, g1215, g1216, g1217, g1218, g1219, g1220, g1221, g1222, g1223, g1224, g1225, g1226, g1227, g1228, g1229, g1230, g1232, g1233, g1234;
	wire g1235, g1236, g1237, g1238, g1239, g1240, g1241, g1242, g1243, g1244, g1245, g1246, g1247, g1248, g1249, g1250, g1251, g1252, g1253, g1254, g1255;
	wire g1257, g1258, g1259, g1260, g1261, g1262, g1263, g1264, g1265, g1266, g1267, g1268, g1269, g1270, g1271, g1272, g1273, g1274, g1275, g1276, g1277;
	wire g1278, g1279, g1281, g1282, g1283, g1284, g1285, g1286, g1287, g1288, g1289, g1290, g1291, g1292, g1293, g1294, g1295, g1296, g1297, g1298, g1299;
	wire g1300, g1301, g1302, g1304, g1305, g1306, g1307, g1308, g1309, g1310, g1311, g1312, g1313, g1314, g1315, g1316, g1317, g1318, g1320, g1321, g1322;
	wire g1323, g1324, g1325, g1326, g1327, g1328, g1329, g1330, g1331, g1332, g1333, g1334, g1335, g1336, g1337, g1338, g1340, g1341, g1342, g1343, g1344;
	wire g1345, g1346, g1347, g1348, g1349, g1350, g1351, g1352, g1354, g1355, g1356, g1357, g1358, g1359, g1360, g1361, g1362, g1363, g1364, g1365, g1366;
	wire g1367, g1369, g1370, g1371, g1372, g1373, g1374, g1375, g1376, g1377, g1378, g1379, g1380, g1381, g1382, g1383, g1385, g1386, g1387, g1388, g1389;
	wire g1390, g1391, g1392, g1393, g1394, g1396, g1397, g1398, g1399, g1400, g1401, g1402, g1403, g1404, g1405, g1406, g1407, g1409, g1410, g1411, g1412;
	wire g1414, g1415, g1416, g1417, g1418, g1420, g1421, g1422, g1423, g1424, g1426, g1427, g1428, g1429, g1430, g1432, g1433, g1434, g1435, g1437, g1438;
	wire g1439, g1440, g1442, g1443, g1445, g1448, g1449, g1450, g1453, g1451, g1452, g1456, g1457, g1454, g1455, g1458, g1459;

	assign sinx0x = (((sk[0]) & (!g1067)));
	assign sinx1x = (((sk[1]) & (!g1107)));
	assign sinx2x = (((sk[2]) & (!g1134)));
	assign sinx5x = (((sk[3]) & (!g1208)));
	assign sinx6x = (((sk[4]) & (!g1231)));
	assign sinx8x = (((sk[5]) & (!g1280)));
	assign sinx9x = (((sk[6]) & (!g1303)));
	assign sinx11x = (((sk[7]) & (!g1339)));
	assign sinx18x = (((sk[8]) & (!g1419)));
	assign sinx20x = (((sk[9]) & (!g1431)));
	assign sinx22x = (((sk[10]) & (!g1441)));
	assign g1 = (((!ax3x) & (!ax2x) & (!ax0x) & (!sk[11]) & (ax1x)) + ((!ax3x) & (!ax2x) & (!ax0x) & (sk[11]) & (!ax1x)) + ((!ax3x) & (!ax2x) & (ax0x) & (!sk[11]) & (ax1x)) + ((!ax3x) & (ax2x) & (!ax0x) & (!sk[11]) & (!ax1x)) + ((!ax3x) & (ax2x) & (!ax0x) & (!sk[11]) & (ax1x)) + ((!ax3x) & (ax2x) & (ax0x) & (!sk[11]) & (!ax1x)) + ((!ax3x) & (ax2x) & (ax0x) & (!sk[11]) & (ax1x)) + ((ax3x) & (!ax2x) & (!ax0x) & (!sk[11]) & (ax1x)) + ((ax3x) & (!ax2x) & (ax0x) & (!sk[11]) & (!ax1x)) + ((ax3x) & (!ax2x) & (ax0x) & (!sk[11]) & (ax1x)) + ((ax3x) & (ax2x) & (!ax0x) & (!sk[11]) & (!ax1x)) + ((ax3x) & (ax2x) & (!ax0x) & (!sk[11]) & (ax1x)) + ((ax3x) & (ax2x) & (ax0x) & (!sk[11]) & (!ax1x)) + ((ax3x) & (ax2x) & (ax0x) & (!sk[11]) & (ax1x)));
	assign g2 = (((!ax22x) & (!ax5x) & (!g1) & (!sk[12]) & (ax4x)) + ((!ax22x) & (!ax5x) & (!g1) & (sk[12]) & (!ax4x)) + ((!ax22x) & (!ax5x) & (!g1) & (sk[12]) & (ax4x)) + ((!ax22x) & (!ax5x) & (g1) & (!sk[12]) & (ax4x)) + ((!ax22x) & (!ax5x) & (g1) & (sk[12]) & (ax4x)) + ((!ax22x) & (ax5x) & (!g1) & (!sk[12]) & (!ax4x)) + ((!ax22x) & (ax5x) & (!g1) & (!sk[12]) & (ax4x)) + ((!ax22x) & (ax5x) & (g1) & (!sk[12]) & (!ax4x)) + ((!ax22x) & (ax5x) & (g1) & (!sk[12]) & (ax4x)) + ((!ax22x) & (ax5x) & (g1) & (sk[12]) & (!ax4x)) + ((ax22x) & (!ax5x) & (!g1) & (!sk[12]) & (ax4x)) + ((ax22x) & (!ax5x) & (g1) & (!sk[12]) & (!ax4x)) + ((ax22x) & (!ax5x) & (g1) & (!sk[12]) & (ax4x)) + ((ax22x) & (ax5x) & (!g1) & (!sk[12]) & (!ax4x)) + ((ax22x) & (ax5x) & (!g1) & (!sk[12]) & (ax4x)) + ((ax22x) & (ax5x) & (!g1) & (sk[12]) & (!ax4x)) + ((ax22x) & (ax5x) & (!g1) & (sk[12]) & (ax4x)) + ((ax22x) & (ax5x) & (g1) & (!sk[12]) & (!ax4x)) + ((ax22x) & (ax5x) & (g1) & (!sk[12]) & (ax4x)) + ((ax22x) & (ax5x) & (g1) & (sk[12]) & (!ax4x)) + ((ax22x) & (ax5x) & (g1) & (sk[12]) & (ax4x)));
	assign g3 = (((!ax5x) & (!ax3x) & (!ax2x) & (!ax0x) & (!ax1x) & (!ax4x)));
	assign g4 = (((!ax9x) & (!ax7x) & (g3) & (!ax6x) & (!ax8x) & (!ax10x)));
	assign g5 = (((!ax13x) & (!ax11x) & (g4) & (!ax12x) & (!ax14x) & (!ax15x)));
	assign g6 = (((!ax19x) & (!ax17x) & (!ax16x) & (g5) & (!sk[16]) & (ax18x)) + ((!ax19x) & (!ax17x) & (!ax16x) & (g5) & (sk[16]) & (!ax18x)) + ((!ax19x) & (!ax17x) & (ax16x) & (g5) & (!sk[16]) & (ax18x)) + ((!ax19x) & (ax17x) & (!ax16x) & (!g5) & (!sk[16]) & (ax18x)) + ((!ax19x) & (ax17x) & (!ax16x) & (g5) & (!sk[16]) & (ax18x)) + ((!ax19x) & (ax17x) & (ax16x) & (!g5) & (!sk[16]) & (ax18x)) + ((!ax19x) & (ax17x) & (ax16x) & (g5) & (!sk[16]) & (ax18x)) + ((ax19x) & (!ax17x) & (!ax16x) & (!g5) & (!sk[16]) & (ax18x)) + ((ax19x) & (!ax17x) & (!ax16x) & (g5) & (!sk[16]) & (ax18x)) + ((ax19x) & (!ax17x) & (ax16x) & (!g5) & (!sk[16]) & (ax18x)) + ((ax19x) & (!ax17x) & (ax16x) & (g5) & (!sk[16]) & (ax18x)) + ((ax19x) & (ax17x) & (!ax16x) & (!g5) & (!sk[16]) & (ax18x)) + ((ax19x) & (ax17x) & (!ax16x) & (g5) & (!sk[16]) & (ax18x)) + ((ax19x) & (ax17x) & (ax16x) & (!g5) & (!sk[16]) & (ax18x)) + ((ax19x) & (ax17x) & (ax16x) & (g5) & (!sk[16]) & (ax18x)));
	assign g7 = (((!ax13x) & (!ax11x) & (!sk[17]) & (g4) & (!ax12x)) + ((!ax13x) & (!ax11x) & (!sk[17]) & (g4) & (ax12x)) + ((!ax13x) & (!ax11x) & (sk[17]) & (g4) & (!ax12x)) + ((!ax13x) & (ax11x) & (!sk[17]) & (g4) & (!ax12x)) + ((!ax13x) & (ax11x) & (!sk[17]) & (g4) & (ax12x)) + ((ax13x) & (!ax11x) & (!sk[17]) & (!g4) & (!ax12x)) + ((ax13x) & (!ax11x) & (!sk[17]) & (!g4) & (ax12x)) + ((ax13x) & (!ax11x) & (!sk[17]) & (g4) & (!ax12x)) + ((ax13x) & (!ax11x) & (!sk[17]) & (g4) & (ax12x)) + ((ax13x) & (ax11x) & (!sk[17]) & (!g4) & (!ax12x)) + ((ax13x) & (ax11x) & (!sk[17]) & (!g4) & (ax12x)) + ((ax13x) & (ax11x) & (!sk[17]) & (g4) & (!ax12x)) + ((ax13x) & (ax11x) & (!sk[17]) & (g4) & (ax12x)));
	assign g8 = (((!ax22x) & (!g7) & (!ax14x) & (sk[18]) & (!ax15x)) + ((!ax22x) & (!g7) & (ax14x) & (!sk[18]) & (!ax15x)) + ((!ax22x) & (!g7) & (ax14x) & (!sk[18]) & (ax15x)) + ((!ax22x) & (!g7) & (ax14x) & (sk[18]) & (!ax15x)) + ((!ax22x) & (g7) & (!ax14x) & (sk[18]) & (ax15x)) + ((!ax22x) & (g7) & (ax14x) & (!sk[18]) & (!ax15x)) + ((!ax22x) & (g7) & (ax14x) & (!sk[18]) & (ax15x)) + ((!ax22x) & (g7) & (ax14x) & (sk[18]) & (!ax15x)) + ((ax22x) & (!g7) & (!ax14x) & (!sk[18]) & (!ax15x)) + ((ax22x) & (!g7) & (!ax14x) & (!sk[18]) & (ax15x)) + ((ax22x) & (!g7) & (!ax14x) & (sk[18]) & (ax15x)) + ((ax22x) & (!g7) & (ax14x) & (!sk[18]) & (!ax15x)) + ((ax22x) & (!g7) & (ax14x) & (!sk[18]) & (ax15x)) + ((ax22x) & (!g7) & (ax14x) & (sk[18]) & (ax15x)) + ((ax22x) & (g7) & (!ax14x) & (!sk[18]) & (!ax15x)) + ((ax22x) & (g7) & (!ax14x) & (!sk[18]) & (ax15x)) + ((ax22x) & (g7) & (!ax14x) & (sk[18]) & (ax15x)) + ((ax22x) & (g7) & (ax14x) & (!sk[18]) & (!ax15x)) + ((ax22x) & (g7) & (ax14x) & (!sk[18]) & (ax15x)) + ((ax22x) & (g7) & (ax14x) & (sk[18]) & (ax15x)));
	assign g9 = (((!ax22x) & (!ax21x) & (!sk[19]) & (!g6) & (ax20x) & (!g8)) + ((!ax22x) & (!ax21x) & (!sk[19]) & (!g6) & (ax20x) & (g8)) + ((!ax22x) & (!ax21x) & (!sk[19]) & (g6) & (ax20x) & (!g8)) + ((!ax22x) & (!ax21x) & (!sk[19]) & (g6) & (ax20x) & (g8)) + ((!ax22x) & (!ax21x) & (sk[19]) & (!g6) & (!ax20x) & (!g8)) + ((!ax22x) & (!ax21x) & (sk[19]) & (g6) & (ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[19]) & (!g6) & (!ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[19]) & (!g6) & (!ax20x) & (g8)) + ((!ax22x) & (ax21x) & (!sk[19]) & (!g6) & (ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[19]) & (!g6) & (ax20x) & (g8)) + ((!ax22x) & (ax21x) & (!sk[19]) & (g6) & (!ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[19]) & (g6) & (!ax20x) & (g8)) + ((!ax22x) & (ax21x) & (!sk[19]) & (g6) & (ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[19]) & (g6) & (ax20x) & (g8)) + ((ax22x) & (!ax21x) & (!sk[19]) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (!sk[19]) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (!ax21x) & (!sk[19]) & (g6) & (!ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (!sk[19]) & (g6) & (!ax20x) & (g8)) + ((ax22x) & (!ax21x) & (!sk[19]) & (g6) & (ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (!sk[19]) & (g6) & (ax20x) & (g8)) + ((ax22x) & (ax21x) & (!sk[19]) & (!g6) & (!ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!sk[19]) & (!g6) & (!ax20x) & (g8)) + ((ax22x) & (ax21x) & (!sk[19]) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!sk[19]) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (ax21x) & (!sk[19]) & (g6) & (!ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!sk[19]) & (g6) & (!ax20x) & (g8)) + ((ax22x) & (ax21x) & (!sk[19]) & (g6) & (ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!sk[19]) & (g6) & (ax20x) & (g8)) + ((ax22x) & (ax21x) & (sk[19]) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (ax21x) & (sk[19]) & (g6) & (ax20x) & (!g8)));
	assign g10 = (((!ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)));
	assign g11 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g10)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g10)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g10)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g10)));
	assign g12 = (((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)));
	assign g13 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g12)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g12)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g12)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g12)));
	assign g14 = (((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)));
	assign g15 = (((!g9) & (!g11) & (!g13) & (sk[25]) & (!g14)) + ((!g9) & (!g11) & (!g13) & (sk[25]) & (g14)) + ((!g9) & (!g11) & (g13) & (!sk[25]) & (!g14)) + ((!g9) & (!g11) & (g13) & (!sk[25]) & (g14)) + ((!g9) & (g11) & (g13) & (!sk[25]) & (!g14)) + ((!g9) & (g11) & (g13) & (!sk[25]) & (g14)) + ((g9) & (!g11) & (!g13) & (!sk[25]) & (!g14)) + ((g9) & (!g11) & (!g13) & (!sk[25]) & (g14)) + ((g9) & (!g11) & (!g13) & (sk[25]) & (!g14)) + ((g9) & (!g11) & (g13) & (!sk[25]) & (!g14)) + ((g9) & (!g11) & (g13) & (!sk[25]) & (g14)) + ((g9) & (g11) & (!g13) & (!sk[25]) & (!g14)) + ((g9) & (g11) & (!g13) & (!sk[25]) & (g14)) + ((g9) & (g11) & (g13) & (!sk[25]) & (!g14)) + ((g9) & (g11) & (g13) & (!sk[25]) & (g14)));
	assign g16 = (((!ax22x) & (!ax21x) & (!g6) & (!sk[26]) & (ax20x) & (!g8)) + ((!ax22x) & (!ax21x) & (!g6) & (!sk[26]) & (ax20x) & (g8)) + ((!ax22x) & (!ax21x) & (!g6) & (sk[26]) & (!ax20x) & (g8)) + ((!ax22x) & (!ax21x) & (g6) & (!sk[26]) & (ax20x) & (!g8)) + ((!ax22x) & (!ax21x) & (g6) & (!sk[26]) & (ax20x) & (g8)) + ((!ax22x) & (!ax21x) & (g6) & (sk[26]) & (ax20x) & (g8)) + ((!ax22x) & (ax21x) & (!g6) & (!sk[26]) & (!ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!g6) & (!sk[26]) & (!ax20x) & (g8)) + ((!ax22x) & (ax21x) & (!g6) & (!sk[26]) & (ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!g6) & (!sk[26]) & (ax20x) & (g8)) + ((!ax22x) & (ax21x) & (g6) & (!sk[26]) & (!ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (g6) & (!sk[26]) & (!ax20x) & (g8)) + ((!ax22x) & (ax21x) & (g6) & (!sk[26]) & (ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (g6) & (!sk[26]) & (ax20x) & (g8)) + ((ax22x) & (!ax21x) & (!g6) & (!sk[26]) & (ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (!g6) & (!sk[26]) & (ax20x) & (g8)) + ((ax22x) & (!ax21x) & (g6) & (!sk[26]) & (!ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (g6) & (!sk[26]) & (!ax20x) & (g8)) + ((ax22x) & (!ax21x) & (g6) & (!sk[26]) & (ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (g6) & (!sk[26]) & (ax20x) & (g8)) + ((ax22x) & (ax21x) & (!g6) & (!sk[26]) & (!ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!g6) & (!sk[26]) & (!ax20x) & (g8)) + ((ax22x) & (ax21x) & (!g6) & (!sk[26]) & (ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!g6) & (!sk[26]) & (ax20x) & (g8)) + ((ax22x) & (ax21x) & (!g6) & (sk[26]) & (ax20x) & (g8)) + ((ax22x) & (ax21x) & (g6) & (!sk[26]) & (!ax20x) & (!g8)) + ((ax22x) & (ax21x) & (g6) & (!sk[26]) & (!ax20x) & (g8)) + ((ax22x) & (ax21x) & (g6) & (!sk[26]) & (ax20x) & (!g8)) + ((ax22x) & (ax21x) & (g6) & (!sk[26]) & (ax20x) & (g8)) + ((ax22x) & (ax21x) & (g6) & (sk[26]) & (ax20x) & (g8)));
	assign g17 = (((!ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)));
	assign g18 = (((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)));
	assign g19 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g12)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g12)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g12)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g12)));
	assign g20 = (((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)));
	assign g21 = (((!ax22x) & (!ax21x) & (!sk[31]) & (!g6) & (ax20x) & (!g20)) + ((!ax22x) & (!ax21x) & (!sk[31]) & (!g6) & (ax20x) & (g20)) + ((!ax22x) & (!ax21x) & (!sk[31]) & (g6) & (ax20x) & (!g20)) + ((!ax22x) & (!ax21x) & (!sk[31]) & (g6) & (ax20x) & (g20)) + ((!ax22x) & (!ax21x) & (sk[31]) & (!g6) & (ax20x) & (g20)) + ((!ax22x) & (ax21x) & (!sk[31]) & (!g6) & (!ax20x) & (!g20)) + ((!ax22x) & (ax21x) & (!sk[31]) & (!g6) & (!ax20x) & (g20)) + ((!ax22x) & (ax21x) & (!sk[31]) & (!g6) & (ax20x) & (!g20)) + ((!ax22x) & (ax21x) & (!sk[31]) & (!g6) & (ax20x) & (g20)) + ((!ax22x) & (ax21x) & (!sk[31]) & (g6) & (!ax20x) & (!g20)) + ((!ax22x) & (ax21x) & (!sk[31]) & (g6) & (!ax20x) & (g20)) + ((!ax22x) & (ax21x) & (!sk[31]) & (g6) & (ax20x) & (!g20)) + ((!ax22x) & (ax21x) & (!sk[31]) & (g6) & (ax20x) & (g20)) + ((!ax22x) & (ax21x) & (sk[31]) & (g6) & (!ax20x) & (g20)) + ((ax22x) & (!ax21x) & (!sk[31]) & (!g6) & (ax20x) & (!g20)) + ((ax22x) & (!ax21x) & (!sk[31]) & (!g6) & (ax20x) & (g20)) + ((ax22x) & (!ax21x) & (!sk[31]) & (g6) & (!ax20x) & (!g20)) + ((ax22x) & (!ax21x) & (!sk[31]) & (g6) & (!ax20x) & (g20)) + ((ax22x) & (!ax21x) & (!sk[31]) & (g6) & (ax20x) & (!g20)) + ((ax22x) & (!ax21x) & (!sk[31]) & (g6) & (ax20x) & (g20)) + ((ax22x) & (ax21x) & (!sk[31]) & (!g6) & (!ax20x) & (!g20)) + ((ax22x) & (ax21x) & (!sk[31]) & (!g6) & (!ax20x) & (g20)) + ((ax22x) & (ax21x) & (!sk[31]) & (!g6) & (ax20x) & (!g20)) + ((ax22x) & (ax21x) & (!sk[31]) & (!g6) & (ax20x) & (g20)) + ((ax22x) & (ax21x) & (!sk[31]) & (g6) & (!ax20x) & (!g20)) + ((ax22x) & (ax21x) & (!sk[31]) & (g6) & (!ax20x) & (g20)) + ((ax22x) & (ax21x) & (!sk[31]) & (g6) & (ax20x) & (!g20)) + ((ax22x) & (ax21x) & (!sk[31]) & (g6) & (ax20x) & (g20)) + ((ax22x) & (ax21x) & (sk[31]) & (!g6) & (!ax20x) & (g20)) + ((ax22x) & (ax21x) & (sk[31]) & (g6) & (!ax20x) & (g20)));
	assign g22 = (((!sk[32]) & (!g16) & (!g17) & (!g18) & (g19) & (!g21)) + ((!sk[32]) & (!g16) & (!g17) & (!g18) & (g19) & (g21)) + ((!sk[32]) & (!g16) & (!g17) & (g18) & (g19) & (!g21)) + ((!sk[32]) & (!g16) & (!g17) & (g18) & (g19) & (g21)) + ((!sk[32]) & (!g16) & (g17) & (!g18) & (!g19) & (!g21)) + ((!sk[32]) & (!g16) & (g17) & (!g18) & (!g19) & (g21)) + ((!sk[32]) & (!g16) & (g17) & (!g18) & (g19) & (!g21)) + ((!sk[32]) & (!g16) & (g17) & (!g18) & (g19) & (g21)) + ((!sk[32]) & (!g16) & (g17) & (g18) & (!g19) & (!g21)) + ((!sk[32]) & (!g16) & (g17) & (g18) & (!g19) & (g21)) + ((!sk[32]) & (!g16) & (g17) & (g18) & (g19) & (!g21)) + ((!sk[32]) & (!g16) & (g17) & (g18) & (g19) & (g21)) + ((!sk[32]) & (g16) & (!g17) & (!g18) & (g19) & (!g21)) + ((!sk[32]) & (g16) & (!g17) & (!g18) & (g19) & (g21)) + ((!sk[32]) & (g16) & (!g17) & (g18) & (!g19) & (!g21)) + ((!sk[32]) & (g16) & (!g17) & (g18) & (!g19) & (g21)) + ((!sk[32]) & (g16) & (!g17) & (g18) & (g19) & (!g21)) + ((!sk[32]) & (g16) & (!g17) & (g18) & (g19) & (g21)) + ((!sk[32]) & (g16) & (g17) & (!g18) & (!g19) & (!g21)) + ((!sk[32]) & (g16) & (g17) & (!g18) & (!g19) & (g21)) + ((!sk[32]) & (g16) & (g17) & (!g18) & (g19) & (!g21)) + ((!sk[32]) & (g16) & (g17) & (!g18) & (g19) & (g21)) + ((!sk[32]) & (g16) & (g17) & (g18) & (!g19) & (!g21)) + ((!sk[32]) & (g16) & (g17) & (g18) & (!g19) & (g21)) + ((!sk[32]) & (g16) & (g17) & (g18) & (g19) & (!g21)) + ((!sk[32]) & (g16) & (g17) & (g18) & (g19) & (g21)) + ((sk[32]) & (!g16) & (!g17) & (!g18) & (!g19) & (!g21)) + ((sk[32]) & (!g16) & (!g17) & (g18) & (!g19) & (!g21)) + ((sk[32]) & (!g16) & (g17) & (!g18) & (!g19) & (!g21)) + ((sk[32]) & (!g16) & (g17) & (g18) & (!g19) & (!g21)) + ((sk[32]) & (g16) & (!g17) & (!g18) & (!g19) & (!g21)));
	assign g23 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)));
	assign g24 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g23)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g23)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g23)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g23)));
	assign g25 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)));
	assign g26 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g25)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g25)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g25)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g25)));
	assign g27 = (((!ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)));
	assign g28 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g27)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g27)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g27)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g27)));
	assign g29 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g27)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g27)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g27)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g27)));
	assign g30 = (((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)));
	assign g31 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g30)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g30)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g30)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g30)));
	assign g32 = (((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)));
	assign g33 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g32)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g32)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g32)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g32)));
	assign g34 = (((!g24) & (!g26) & (!g28) & (!g29) & (!g31) & (!g33)));
	assign g35 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g25)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g25)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g25)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g25)));
	assign g36 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g30)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g30)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g30)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g30)));
	assign g37 = (((!g35) & (!sk[47]) & (g36)) + ((!g35) & (sk[47]) & (!g36)) + ((g35) & (!sk[47]) & (g36)));
	assign g38 = (((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)));
	assign g39 = (((!g38) & (!g9) & (!sk[49]) & (g16) & (!g30)) + ((!g38) & (!g9) & (!sk[49]) & (g16) & (g30)) + ((!g38) & (!g9) & (sk[49]) & (!g16) & (!g30)) + ((!g38) & (!g9) & (sk[49]) & (!g16) & (g30)) + ((!g38) & (!g9) & (sk[49]) & (g16) & (!g30)) + ((!g38) & (g9) & (!sk[49]) & (g16) & (!g30)) + ((!g38) & (g9) & (!sk[49]) & (g16) & (g30)) + ((!g38) & (g9) & (sk[49]) & (!g16) & (!g30)) + ((!g38) & (g9) & (sk[49]) & (g16) & (!g30)) + ((g38) & (!g9) & (!sk[49]) & (!g16) & (!g30)) + ((g38) & (!g9) & (!sk[49]) & (!g16) & (g30)) + ((g38) & (!g9) & (!sk[49]) & (g16) & (!g30)) + ((g38) & (!g9) & (!sk[49]) & (g16) & (g30)) + ((g38) & (!g9) & (sk[49]) & (!g16) & (!g30)) + ((g38) & (!g9) & (sk[49]) & (!g16) & (g30)) + ((g38) & (!g9) & (sk[49]) & (g16) & (!g30)) + ((g38) & (g9) & (!sk[49]) & (!g16) & (!g30)) + ((g38) & (g9) & (!sk[49]) & (!g16) & (g30)) + ((g38) & (g9) & (!sk[49]) & (g16) & (!g30)) + ((g38) & (g9) & (!sk[49]) & (g16) & (g30)));
	assign g40 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)));
	assign g41 = (((!ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)));
	assign g42 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)));
	assign g43 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g42)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g42)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g42)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g42)));
	assign g44 = (((!g9) & (!g16) & (!g12) & (!g40) & (!g41) & (!g43)) + ((!g9) & (!g16) & (!g12) & (!g40) & (g41) & (!g43)) + ((!g9) & (!g16) & (!g12) & (g40) & (!g41) & (!g43)) + ((!g9) & (!g16) & (!g12) & (g40) & (g41) & (!g43)) + ((!g9) & (!g16) & (g12) & (!g40) & (!g41) & (!g43)) + ((!g9) & (!g16) & (g12) & (!g40) & (g41) & (!g43)) + ((!g9) & (!g16) & (g12) & (g40) & (!g41) & (!g43)) + ((!g9) & (!g16) & (g12) & (g40) & (g41) & (!g43)) + ((!g9) & (g16) & (!g12) & (!g40) & (!g41) & (!g43)) + ((!g9) & (g16) & (!g12) & (!g40) & (g41) & (!g43)) + ((g9) & (!g16) & (!g12) & (!g40) & (!g41) & (!g43)) + ((g9) & (!g16) & (g12) & (!g40) & (!g41) & (!g43)) + ((g9) & (g16) & (!g12) & (!g40) & (!g41) & (!g43)));
	assign g45 = (((g15) & (g22) & (g34) & (g37) & (g39) & (g44)));
	assign g46 = (((!ax22x) & (!ax21x) & (!sk[56]) & (!g6) & (ax20x) & (!g8)) + ((!ax22x) & (!ax21x) & (!sk[56]) & (!g6) & (ax20x) & (g8)) + ((!ax22x) & (!ax21x) & (!sk[56]) & (g6) & (ax20x) & (!g8)) + ((!ax22x) & (!ax21x) & (!sk[56]) & (g6) & (ax20x) & (g8)) + ((!ax22x) & (!ax21x) & (sk[56]) & (!g6) & (ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[56]) & (!g6) & (!ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[56]) & (!g6) & (!ax20x) & (g8)) + ((!ax22x) & (ax21x) & (!sk[56]) & (!g6) & (ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[56]) & (!g6) & (ax20x) & (g8)) + ((!ax22x) & (ax21x) & (!sk[56]) & (g6) & (!ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[56]) & (g6) & (!ax20x) & (g8)) + ((!ax22x) & (ax21x) & (!sk[56]) & (g6) & (ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[56]) & (g6) & (ax20x) & (g8)) + ((!ax22x) & (ax21x) & (sk[56]) & (g6) & (!ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (!sk[56]) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (!sk[56]) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (!ax21x) & (!sk[56]) & (g6) & (!ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (!sk[56]) & (g6) & (!ax20x) & (g8)) + ((ax22x) & (!ax21x) & (!sk[56]) & (g6) & (ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (!sk[56]) & (g6) & (ax20x) & (g8)) + ((ax22x) & (ax21x) & (!sk[56]) & (!g6) & (!ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!sk[56]) & (!g6) & (!ax20x) & (g8)) + ((ax22x) & (ax21x) & (!sk[56]) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!sk[56]) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (ax21x) & (!sk[56]) & (g6) & (!ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!sk[56]) & (g6) & (!ax20x) & (g8)) + ((ax22x) & (ax21x) & (!sk[56]) & (g6) & (ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!sk[56]) & (g6) & (ax20x) & (g8)) + ((ax22x) & (ax21x) & (sk[56]) & (!g6) & (!ax20x) & (!g8)) + ((ax22x) & (ax21x) & (sk[56]) & (g6) & (!ax20x) & (!g8)));
	assign g47 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g10)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g10)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g10)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g10)));
	assign g48 = (((!sk[58]) & (!g17) & (!g46) & (g47)) + ((!sk[58]) & (!g17) & (g46) & (g47)) + ((!sk[58]) & (g17) & (!g46) & (!g47)) + ((!sk[58]) & (g17) & (!g46) & (g47)) + ((!sk[58]) & (g17) & (g46) & (!g47)) + ((!sk[58]) & (g17) & (g46) & (g47)) + ((sk[58]) & (!g17) & (!g46) & (!g47)) + ((sk[58]) & (!g17) & (g46) & (!g47)) + ((sk[58]) & (g17) & (!g46) & (!g47)));
	assign g49 = (((!ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)));
	assign g50 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g49)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g49)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g49)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g49)));
	assign g51 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g17)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g17)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g17)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g17)));
	assign g52 = (((!sk[62]) & (!g50) & (g51)) + ((!sk[62]) & (g50) & (g51)) + ((sk[62]) & (!g50) & (!g51)));
	assign g53 = (((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)));
	assign g54 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g53)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g53)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g53)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g53)));
	assign g55 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g20)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g20)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g20)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g20)));
	assign g56 = (((!sk[66]) & (!g54) & (g55)) + ((!sk[66]) & (g54) & (g55)) + ((sk[66]) & (!g54) & (!g55)));
	assign g57 = (((!ax22x) & (!ax21x) & (!g6) & (sk[67]) & (ax20x)) + ((!ax22x) & (!ax21x) & (g6) & (!sk[67]) & (!ax20x)) + ((!ax22x) & (!ax21x) & (g6) & (!sk[67]) & (ax20x)) + ((!ax22x) & (ax21x) & (g6) & (!sk[67]) & (!ax20x)) + ((!ax22x) & (ax21x) & (g6) & (!sk[67]) & (ax20x)) + ((!ax22x) & (ax21x) & (g6) & (sk[67]) & (!ax20x)) + ((ax22x) & (!ax21x) & (!g6) & (!sk[67]) & (!ax20x)) + ((ax22x) & (!ax21x) & (!g6) & (!sk[67]) & (ax20x)) + ((ax22x) & (!ax21x) & (g6) & (!sk[67]) & (!ax20x)) + ((ax22x) & (!ax21x) & (g6) & (!sk[67]) & (ax20x)) + ((ax22x) & (ax21x) & (!g6) & (!sk[67]) & (!ax20x)) + ((ax22x) & (ax21x) & (!g6) & (!sk[67]) & (ax20x)) + ((ax22x) & (ax21x) & (!g6) & (sk[67]) & (!ax20x)) + ((ax22x) & (ax21x) & (g6) & (!sk[67]) & (!ax20x)) + ((ax22x) & (ax21x) & (g6) & (!sk[67]) & (ax20x)) + ((ax22x) & (ax21x) & (g6) & (sk[67]) & (!ax20x)));
	assign g58 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)));
	assign g59 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g49)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g49)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g49)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g49)));
	assign g60 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g20)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g20)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g20)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g20)));
	assign g61 = (((!g57) & (!g58) & (!g32) & (!g59) & (sk[71]) & (!g60)) + ((!g57) & (!g58) & (!g32) & (g59) & (!sk[71]) & (!g60)) + ((!g57) & (!g58) & (!g32) & (g59) & (!sk[71]) & (g60)) + ((!g57) & (!g58) & (g32) & (!g59) & (sk[71]) & (!g60)) + ((!g57) & (!g58) & (g32) & (g59) & (!sk[71]) & (!g60)) + ((!g57) & (!g58) & (g32) & (g59) & (!sk[71]) & (g60)) + ((!g57) & (g58) & (!g32) & (!g59) & (!sk[71]) & (!g60)) + ((!g57) & (g58) & (!g32) & (!g59) & (!sk[71]) & (g60)) + ((!g57) & (g58) & (!g32) & (!g59) & (sk[71]) & (!g60)) + ((!g57) & (g58) & (!g32) & (g59) & (!sk[71]) & (!g60)) + ((!g57) & (g58) & (!g32) & (g59) & (!sk[71]) & (g60)) + ((!g57) & (g58) & (g32) & (!g59) & (!sk[71]) & (!g60)) + ((!g57) & (g58) & (g32) & (!g59) & (!sk[71]) & (g60)) + ((!g57) & (g58) & (g32) & (!g59) & (sk[71]) & (!g60)) + ((!g57) & (g58) & (g32) & (g59) & (!sk[71]) & (!g60)) + ((!g57) & (g58) & (g32) & (g59) & (!sk[71]) & (g60)) + ((g57) & (!g58) & (!g32) & (!g59) & (sk[71]) & (!g60)) + ((g57) & (!g58) & (!g32) & (g59) & (!sk[71]) & (!g60)) + ((g57) & (!g58) & (!g32) & (g59) & (!sk[71]) & (g60)) + ((g57) & (!g58) & (g32) & (!g59) & (!sk[71]) & (!g60)) + ((g57) & (!g58) & (g32) & (!g59) & (!sk[71]) & (g60)) + ((g57) & (!g58) & (g32) & (g59) & (!sk[71]) & (!g60)) + ((g57) & (!g58) & (g32) & (g59) & (!sk[71]) & (g60)) + ((g57) & (g58) & (!g32) & (!g59) & (!sk[71]) & (!g60)) + ((g57) & (g58) & (!g32) & (!g59) & (!sk[71]) & (g60)) + ((g57) & (g58) & (!g32) & (g59) & (!sk[71]) & (!g60)) + ((g57) & (g58) & (!g32) & (g59) & (!sk[71]) & (g60)) + ((g57) & (g58) & (g32) & (!g59) & (!sk[71]) & (!g60)) + ((g57) & (g58) & (g32) & (!g59) & (!sk[71]) & (g60)) + ((g57) & (g58) & (g32) & (g59) & (!sk[71]) & (!g60)) + ((g57) & (g58) & (g32) & (g59) & (!sk[71]) & (g60)));
	assign g62 = (((!sk[72]) & (!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8)) + ((!sk[72]) & (!ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8)) + ((!sk[72]) & (!ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8)) + ((!sk[72]) & (!ax22x) & (!ax21x) & (g6) & (ax20x) & (g8)) + ((!sk[72]) & (!ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8)) + ((!sk[72]) & (!ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8)) + ((!sk[72]) & (!ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8)) + ((!sk[72]) & (!ax22x) & (ax21x) & (!g6) & (ax20x) & (g8)) + ((!sk[72]) & (!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8)) + ((!sk[72]) & (!ax22x) & (ax21x) & (g6) & (!ax20x) & (g8)) + ((!sk[72]) & (!ax22x) & (ax21x) & (g6) & (ax20x) & (!g8)) + ((!sk[72]) & (!ax22x) & (ax21x) & (g6) & (ax20x) & (g8)) + ((!sk[72]) & (ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8)) + ((!sk[72]) & (ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8)) + ((!sk[72]) & (ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8)) + ((!sk[72]) & (ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8)) + ((!sk[72]) & (ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8)) + ((!sk[72]) & (ax22x) & (!ax21x) & (g6) & (ax20x) & (g8)) + ((!sk[72]) & (ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8)) + ((!sk[72]) & (ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8)) + ((!sk[72]) & (ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8)) + ((!sk[72]) & (ax22x) & (ax21x) & (!g6) & (ax20x) & (g8)) + ((!sk[72]) & (ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8)) + ((!sk[72]) & (ax22x) & (ax21x) & (g6) & (!ax20x) & (g8)) + ((!sk[72]) & (ax22x) & (ax21x) & (g6) & (ax20x) & (!g8)) + ((!sk[72]) & (ax22x) & (ax21x) & (g6) & (ax20x) & (g8)) + ((sk[72]) & (!ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8)) + ((sk[72]) & (!ax22x) & (ax21x) & (g6) & (!ax20x) & (g8)) + ((sk[72]) & (ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8)) + ((sk[72]) & (ax22x) & (ax21x) & (g6) & (!ax20x) & (g8)));
	assign g63 = (((!ax22x) & (!sk[73]) & (!ax21x) & (!g6) & (ax20x) & (!g25)) + ((!ax22x) & (!sk[73]) & (!ax21x) & (!g6) & (ax20x) & (g25)) + ((!ax22x) & (!sk[73]) & (!ax21x) & (g6) & (ax20x) & (!g25)) + ((!ax22x) & (!sk[73]) & (!ax21x) & (g6) & (ax20x) & (g25)) + ((!ax22x) & (!sk[73]) & (ax21x) & (!g6) & (!ax20x) & (!g25)) + ((!ax22x) & (!sk[73]) & (ax21x) & (!g6) & (!ax20x) & (g25)) + ((!ax22x) & (!sk[73]) & (ax21x) & (!g6) & (ax20x) & (!g25)) + ((!ax22x) & (!sk[73]) & (ax21x) & (!g6) & (ax20x) & (g25)) + ((!ax22x) & (!sk[73]) & (ax21x) & (g6) & (!ax20x) & (!g25)) + ((!ax22x) & (!sk[73]) & (ax21x) & (g6) & (!ax20x) & (g25)) + ((!ax22x) & (!sk[73]) & (ax21x) & (g6) & (ax20x) & (!g25)) + ((!ax22x) & (!sk[73]) & (ax21x) & (g6) & (ax20x) & (g25)) + ((!ax22x) & (sk[73]) & (!ax21x) & (!g6) & (!ax20x) & (g25)) + ((!ax22x) & (sk[73]) & (!ax21x) & (g6) & (ax20x) & (g25)) + ((ax22x) & (!sk[73]) & (!ax21x) & (!g6) & (ax20x) & (!g25)) + ((ax22x) & (!sk[73]) & (!ax21x) & (!g6) & (ax20x) & (g25)) + ((ax22x) & (!sk[73]) & (!ax21x) & (g6) & (!ax20x) & (!g25)) + ((ax22x) & (!sk[73]) & (!ax21x) & (g6) & (!ax20x) & (g25)) + ((ax22x) & (!sk[73]) & (!ax21x) & (g6) & (ax20x) & (!g25)) + ((ax22x) & (!sk[73]) & (!ax21x) & (g6) & (ax20x) & (g25)) + ((ax22x) & (!sk[73]) & (ax21x) & (!g6) & (!ax20x) & (!g25)) + ((ax22x) & (!sk[73]) & (ax21x) & (!g6) & (!ax20x) & (g25)) + ((ax22x) & (!sk[73]) & (ax21x) & (!g6) & (ax20x) & (!g25)) + ((ax22x) & (!sk[73]) & (ax21x) & (!g6) & (ax20x) & (g25)) + ((ax22x) & (!sk[73]) & (ax21x) & (g6) & (!ax20x) & (!g25)) + ((ax22x) & (!sk[73]) & (ax21x) & (g6) & (!ax20x) & (g25)) + ((ax22x) & (!sk[73]) & (ax21x) & (g6) & (ax20x) & (!g25)) + ((ax22x) & (!sk[73]) & (ax21x) & (g6) & (ax20x) & (g25)) + ((ax22x) & (sk[73]) & (ax21x) & (!g6) & (ax20x) & (g25)) + ((ax22x) & (sk[73]) & (ax21x) & (g6) & (ax20x) & (g25)));
	assign g64 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g58)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g58)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g58)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g58)));
	assign g65 = (((!g38) & (!g62) & (!g46) & (!g63) & (!g42) & (!g64)) + ((!g38) & (!g62) & (!g46) & (!g63) & (g42) & (!g64)) + ((!g38) & (!g62) & (g46) & (!g63) & (!g42) & (!g64)) + ((!g38) & (g62) & (!g46) & (!g63) & (!g42) & (!g64)) + ((!g38) & (g62) & (!g46) & (!g63) & (g42) & (!g64)) + ((!g38) & (g62) & (g46) & (!g63) & (!g42) & (!g64)) + ((g38) & (!g62) & (!g46) & (!g63) & (!g42) & (!g64)) + ((g38) & (!g62) & (!g46) & (!g63) & (g42) & (!g64)));
	assign g66 = (((!ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)));
	assign g67 = (((!g38) & (!g9) & (!g16) & (!g41) & (!g42) & (!g66)) + ((!g38) & (!g9) & (!g16) & (!g41) & (!g42) & (g66)) + ((!g38) & (!g9) & (!g16) & (!g41) & (g42) & (!g66)) + ((!g38) & (!g9) & (!g16) & (!g41) & (g42) & (g66)) + ((!g38) & (!g9) & (!g16) & (g41) & (!g42) & (!g66)) + ((!g38) & (!g9) & (!g16) & (g41) & (!g42) & (g66)) + ((!g38) & (!g9) & (!g16) & (g41) & (g42) & (!g66)) + ((!g38) & (!g9) & (!g16) & (g41) & (g42) & (g66)) + ((!g38) & (!g9) & (g16) & (!g41) & (!g42) & (!g66)) + ((!g38) & (g9) & (!g16) & (!g41) & (!g42) & (!g66)) + ((!g38) & (g9) & (!g16) & (g41) & (!g42) & (!g66)) + ((!g38) & (g9) & (g16) & (!g41) & (!g42) & (!g66)) + ((g38) & (!g9) & (!g16) & (!g41) & (!g42) & (!g66)) + ((g38) & (!g9) & (!g16) & (!g41) & (!g42) & (g66)) + ((g38) & (!g9) & (!g16) & (!g41) & (g42) & (!g66)) + ((g38) & (!g9) & (!g16) & (!g41) & (g42) & (g66)) + ((g38) & (!g9) & (!g16) & (g41) & (!g42) & (!g66)) + ((g38) & (!g9) & (!g16) & (g41) & (!g42) & (g66)) + ((g38) & (!g9) & (!g16) & (g41) & (g42) & (!g66)) + ((g38) & (!g9) & (!g16) & (g41) & (g42) & (g66)) + ((g38) & (g9) & (!g16) & (!g41) & (!g42) & (!g66)) + ((g38) & (g9) & (!g16) & (g41) & (!g42) & (!g66)));
	assign g68 = (((g48) & (g52) & (g56) & (g61) & (g65) & (g67)));
	assign g69 = (((!g45) & (!sk[79]) & (g68)) + ((g45) & (!sk[79]) & (g68)) + ((g45) & (sk[79]) & (g68)));
	assign g70 = (((!sk[80]) & (!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8)) + ((!sk[80]) & (!ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8)) + ((!sk[80]) & (!ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8)) + ((!sk[80]) & (!ax22x) & (!ax21x) & (g6) & (ax20x) & (g8)) + ((!sk[80]) & (!ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8)) + ((!sk[80]) & (!ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8)) + ((!sk[80]) & (!ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8)) + ((!sk[80]) & (!ax22x) & (ax21x) & (!g6) & (ax20x) & (g8)) + ((!sk[80]) & (!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8)) + ((!sk[80]) & (!ax22x) & (ax21x) & (g6) & (!ax20x) & (g8)) + ((!sk[80]) & (!ax22x) & (ax21x) & (g6) & (ax20x) & (!g8)) + ((!sk[80]) & (!ax22x) & (ax21x) & (g6) & (ax20x) & (g8)) + ((!sk[80]) & (ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8)) + ((!sk[80]) & (ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8)) + ((!sk[80]) & (ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8)) + ((!sk[80]) & (ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8)) + ((!sk[80]) & (ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8)) + ((!sk[80]) & (ax22x) & (!ax21x) & (g6) & (ax20x) & (g8)) + ((!sk[80]) & (ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8)) + ((!sk[80]) & (ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8)) + ((!sk[80]) & (ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8)) + ((!sk[80]) & (ax22x) & (ax21x) & (!g6) & (ax20x) & (g8)) + ((!sk[80]) & (ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8)) + ((!sk[80]) & (ax22x) & (ax21x) & (g6) & (!ax20x) & (g8)) + ((!sk[80]) & (ax22x) & (ax21x) & (g6) & (ax20x) & (!g8)) + ((!sk[80]) & (ax22x) & (ax21x) & (g6) & (ax20x) & (g8)) + ((sk[80]) & (!ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8)) + ((sk[80]) & (!ax22x) & (ax21x) & (!g6) & (ax20x) & (g8)) + ((sk[80]) & (ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8)) + ((sk[80]) & (ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8)));
	assign g71 = (((!ax22x) & (!ax21x) & (!sk[81]) & (!g6) & (ax20x) & (!g8)) + ((!ax22x) & (!ax21x) & (!sk[81]) & (!g6) & (ax20x) & (g8)) + ((!ax22x) & (!ax21x) & (!sk[81]) & (g6) & (ax20x) & (!g8)) + ((!ax22x) & (!ax21x) & (!sk[81]) & (g6) & (ax20x) & (g8)) + ((!ax22x) & (ax21x) & (!sk[81]) & (!g6) & (!ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[81]) & (!g6) & (!ax20x) & (g8)) + ((!ax22x) & (ax21x) & (!sk[81]) & (!g6) & (ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[81]) & (!g6) & (ax20x) & (g8)) + ((!ax22x) & (ax21x) & (!sk[81]) & (g6) & (!ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[81]) & (g6) & (!ax20x) & (g8)) + ((!ax22x) & (ax21x) & (!sk[81]) & (g6) & (ax20x) & (!g8)) + ((!ax22x) & (ax21x) & (!sk[81]) & (g6) & (ax20x) & (g8)) + ((!ax22x) & (ax21x) & (sk[81]) & (!g6) & (!ax20x) & (g8)) + ((!ax22x) & (ax21x) & (sk[81]) & (g6) & (ax20x) & (g8)) + ((ax22x) & (!ax21x) & (!sk[81]) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (!sk[81]) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (!ax21x) & (!sk[81]) & (g6) & (!ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (!sk[81]) & (g6) & (!ax20x) & (g8)) + ((ax22x) & (!ax21x) & (!sk[81]) & (g6) & (ax20x) & (!g8)) + ((ax22x) & (!ax21x) & (!sk[81]) & (g6) & (ax20x) & (g8)) + ((ax22x) & (!ax21x) & (sk[81]) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (!ax21x) & (sk[81]) & (g6) & (ax20x) & (g8)) + ((ax22x) & (ax21x) & (!sk[81]) & (!g6) & (!ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!sk[81]) & (!g6) & (!ax20x) & (g8)) + ((ax22x) & (ax21x) & (!sk[81]) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!sk[81]) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (ax21x) & (!sk[81]) & (g6) & (!ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!sk[81]) & (g6) & (!ax20x) & (g8)) + ((ax22x) & (ax21x) & (!sk[81]) & (g6) & (ax20x) & (!g8)) + ((ax22x) & (ax21x) & (!sk[81]) & (g6) & (ax20x) & (g8)));
	assign g72 = (((!g70) & (!sk[82]) & (!g10) & (g71) & (!g20)) + ((!g70) & (!sk[82]) & (!g10) & (g71) & (g20)) + ((!g70) & (!sk[82]) & (g10) & (g71) & (!g20)) + ((!g70) & (!sk[82]) & (g10) & (g71) & (g20)) + ((!g70) & (sk[82]) & (!g10) & (g71) & (g20)) + ((!g70) & (sk[82]) & (g10) & (g71) & (g20)) + ((g70) & (!sk[82]) & (!g10) & (!g71) & (!g20)) + ((g70) & (!sk[82]) & (!g10) & (!g71) & (g20)) + ((g70) & (!sk[82]) & (!g10) & (g71) & (!g20)) + ((g70) & (!sk[82]) & (!g10) & (g71) & (g20)) + ((g70) & (!sk[82]) & (g10) & (!g71) & (!g20)) + ((g70) & (!sk[82]) & (g10) & (!g71) & (g20)) + ((g70) & (!sk[82]) & (g10) & (g71) & (!g20)) + ((g70) & (!sk[82]) & (g10) & (g71) & (g20)) + ((g70) & (sk[82]) & (!g10) & (g71) & (g20)) + ((g70) & (sk[82]) & (g10) & (!g71) & (!g20)) + ((g70) & (sk[82]) & (g10) & (!g71) & (g20)) + ((g70) & (sk[82]) & (g10) & (g71) & (!g20)) + ((g70) & (sk[82]) & (g10) & (g71) & (g20)));
	assign g73 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g12)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g12)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g12)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g12)));
	assign g74 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g20)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g20)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g20)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g20)));
	assign g75 = (((!g70) & (!sk[85]) & (!g18) & (g74)) + ((!g70) & (!sk[85]) & (g18) & (g74)) + ((!g70) & (sk[85]) & (!g18) & (!g74)) + ((!g70) & (sk[85]) & (g18) & (!g74)) + ((g70) & (!sk[85]) & (!g18) & (!g74)) + ((g70) & (!sk[85]) & (!g18) & (g74)) + ((g70) & (!sk[85]) & (g18) & (!g74)) + ((g70) & (!sk[85]) & (g18) & (g74)) + ((g70) & (sk[85]) & (!g18) & (!g74)));
	assign g76 = (((!ax22x) & (g38) & (ax21x) & (!g6) & (!ax20x) & (!g8)) + ((!ax22x) & (g38) & (ax21x) & (g6) & (ax20x) & (!g8)) + ((ax22x) & (g38) & (!ax21x) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (g38) & (!ax21x) & (g6) & (ax20x) & (!g8)));
	assign g77 = (((!g76) & (!sk[87]) & (g28)) + ((!g76) & (sk[87]) & (!g28)) + ((g76) & (!sk[87]) & (g28)));
	assign g78 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g49)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g49)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g49)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g49)));
	assign g79 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g17)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g17)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g17)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g17)));
	assign g80 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g10)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g10)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g10)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g10)));
	assign g81 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g32)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g32)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g32)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g32)));
	assign g82 = (((!g78) & (!g79) & (!g35) & (!g60) & (!g80) & (!g81)));
	assign g83 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g18)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g18)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g18)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g18)));
	assign g84 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8) & (g49)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g49)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g49)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8) & (g49)));
	assign g85 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g42)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g42)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g42)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g42)));
	assign g86 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g30)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g30)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g30)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g30)));
	assign g87 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g17)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g17)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g17)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g17)));
	assign g88 = (((!g83) & (!g84) & (!g85) & (!g86) & (sk[98]) & (!g87)) + ((!g83) & (!g84) & (!g85) & (g86) & (!sk[98]) & (!g87)) + ((!g83) & (!g84) & (!g85) & (g86) & (!sk[98]) & (g87)) + ((!g83) & (!g84) & (g85) & (g86) & (!sk[98]) & (!g87)) + ((!g83) & (!g84) & (g85) & (g86) & (!sk[98]) & (g87)) + ((!g83) & (g84) & (!g85) & (!g86) & (!sk[98]) & (!g87)) + ((!g83) & (g84) & (!g85) & (!g86) & (!sk[98]) & (g87)) + ((!g83) & (g84) & (!g85) & (g86) & (!sk[98]) & (!g87)) + ((!g83) & (g84) & (!g85) & (g86) & (!sk[98]) & (g87)) + ((!g83) & (g84) & (g85) & (!g86) & (!sk[98]) & (!g87)) + ((!g83) & (g84) & (g85) & (!g86) & (!sk[98]) & (g87)) + ((!g83) & (g84) & (g85) & (g86) & (!sk[98]) & (!g87)) + ((!g83) & (g84) & (g85) & (g86) & (!sk[98]) & (g87)) + ((g83) & (!g84) & (!g85) & (g86) & (!sk[98]) & (!g87)) + ((g83) & (!g84) & (!g85) & (g86) & (!sk[98]) & (g87)) + ((g83) & (!g84) & (g85) & (!g86) & (!sk[98]) & (!g87)) + ((g83) & (!g84) & (g85) & (!g86) & (!sk[98]) & (g87)) + ((g83) & (!g84) & (g85) & (g86) & (!sk[98]) & (!g87)) + ((g83) & (!g84) & (g85) & (g86) & (!sk[98]) & (g87)) + ((g83) & (g84) & (!g85) & (!g86) & (!sk[98]) & (!g87)) + ((g83) & (g84) & (!g85) & (!g86) & (!sk[98]) & (g87)) + ((g83) & (g84) & (!g85) & (g86) & (!sk[98]) & (!g87)) + ((g83) & (g84) & (!g85) & (g86) & (!sk[98]) & (g87)) + ((g83) & (g84) & (g85) & (!g86) & (!sk[98]) & (!g87)) + ((g83) & (g84) & (g85) & (!g86) & (!sk[98]) & (g87)) + ((g83) & (g84) & (g85) & (g86) & (!sk[98]) & (!g87)) + ((g83) & (g84) & (g85) & (g86) & (!sk[98]) & (g87)));
	assign g89 = (((!g72) & (!g73) & (g75) & (g77) & (g82) & (g88)));
	assign g90 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g40)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g40)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g40)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g40)));
	assign g91 = (((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)));
	assign g92 = (((!g62) & (!sk[102]) & (!g90) & (g91)) + ((!g62) & (!sk[102]) & (g90) & (g91)) + ((!g62) & (sk[102]) & (!g90) & (!g91)) + ((!g62) & (sk[102]) & (!g90) & (g91)) + ((g62) & (!sk[102]) & (!g90) & (!g91)) + ((g62) & (!sk[102]) & (!g90) & (g91)) + ((g62) & (!sk[102]) & (g90) & (!g91)) + ((g62) & (!sk[102]) & (g90) & (g91)) + ((g62) & (sk[102]) & (!g90) & (!g91)));
	assign g93 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8) & (g66)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g66)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g66)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8) & (g66)));
	assign g94 = (((!g71) & (!g25) & (!sk[104]) & (g41) & (!g93)) + ((!g71) & (!g25) & (!sk[104]) & (g41) & (g93)) + ((!g71) & (!g25) & (sk[104]) & (!g41) & (!g93)) + ((!g71) & (!g25) & (sk[104]) & (g41) & (!g93)) + ((!g71) & (g25) & (!sk[104]) & (g41) & (!g93)) + ((!g71) & (g25) & (!sk[104]) & (g41) & (g93)) + ((!g71) & (g25) & (sk[104]) & (!g41) & (!g93)) + ((!g71) & (g25) & (sk[104]) & (g41) & (!g93)) + ((g71) & (!g25) & (!sk[104]) & (!g41) & (!g93)) + ((g71) & (!g25) & (!sk[104]) & (!g41) & (g93)) + ((g71) & (!g25) & (!sk[104]) & (g41) & (!g93)) + ((g71) & (!g25) & (!sk[104]) & (g41) & (g93)) + ((g71) & (!g25) & (sk[104]) & (!g41) & (!g93)) + ((g71) & (g25) & (!sk[104]) & (!g41) & (!g93)) + ((g71) & (g25) & (!sk[104]) & (!g41) & (g93)) + ((g71) & (g25) & (!sk[104]) & (g41) & (!g93)) + ((g71) & (g25) & (!sk[104]) & (g41) & (g93)));
	assign g95 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g20)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g20)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g20)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g20)));
	assign g96 = (((!sk[106]) & (!g17) & (!g71) & (g95)) + ((!sk[106]) & (!g17) & (g71) & (g95)) + ((!sk[106]) & (g17) & (!g71) & (!g95)) + ((!sk[106]) & (g17) & (!g71) & (g95)) + ((!sk[106]) & (g17) & (g71) & (!g95)) + ((!sk[106]) & (g17) & (g71) & (g95)) + ((sk[106]) & (!g17) & (!g71) & (!g95)) + ((sk[106]) & (!g17) & (g71) & (!g95)) + ((sk[106]) & (g17) & (!g71) & (!g95)));
	assign g97 = (((!sk[107]) & (!ax22x) & (!ax17x) & (ax16x) & (!g5)) + ((!sk[107]) & (!ax22x) & (!ax17x) & (ax16x) & (g5)) + ((!sk[107]) & (!ax22x) & (ax17x) & (ax16x) & (!g5)) + ((!sk[107]) & (!ax22x) & (ax17x) & (ax16x) & (g5)) + ((!sk[107]) & (ax22x) & (!ax17x) & (!ax16x) & (!g5)) + ((!sk[107]) & (ax22x) & (!ax17x) & (!ax16x) & (g5)) + ((!sk[107]) & (ax22x) & (!ax17x) & (ax16x) & (!g5)) + ((!sk[107]) & (ax22x) & (!ax17x) & (ax16x) & (g5)) + ((!sk[107]) & (ax22x) & (ax17x) & (!ax16x) & (!g5)) + ((!sk[107]) & (ax22x) & (ax17x) & (!ax16x) & (g5)) + ((!sk[107]) & (ax22x) & (ax17x) & (ax16x) & (!g5)) + ((!sk[107]) & (ax22x) & (ax17x) & (ax16x) & (g5)) + ((sk[107]) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5)) + ((sk[107]) & (!ax22x) & (!ax17x) & (ax16x) & (!g5)) + ((sk[107]) & (!ax22x) & (!ax17x) & (ax16x) & (g5)) + ((sk[107]) & (!ax22x) & (ax17x) & (!ax16x) & (g5)) + ((sk[107]) & (ax22x) & (ax17x) & (!ax16x) & (!g5)) + ((sk[107]) & (ax22x) & (ax17x) & (!ax16x) & (g5)) + ((sk[107]) & (ax22x) & (ax17x) & (ax16x) & (!g5)) + ((sk[107]) & (ax22x) & (ax17x) & (ax16x) & (g5)));
	assign g98 = (((!ax22x) & (!sk[108]) & (!ax16x) & (g5)) + ((!ax22x) & (!sk[108]) & (ax16x) & (g5)) + ((!ax22x) & (sk[108]) & (!ax16x) & (!g5)) + ((!ax22x) & (sk[108]) & (ax16x) & (g5)) + ((ax22x) & (!sk[108]) & (!ax16x) & (!g5)) + ((ax22x) & (!sk[108]) & (!ax16x) & (g5)) + ((ax22x) & (!sk[108]) & (ax16x) & (!g5)) + ((ax22x) & (!sk[108]) & (ax16x) & (g5)) + ((ax22x) & (sk[108]) & (ax16x) & (!g5)) + ((ax22x) & (sk[108]) & (ax16x) & (g5)));
	assign g99 = (((!ax22x) & (!sk[109]) & (!ax21x) & (!g6) & (ax20x) & (!g8)) + ((!ax22x) & (!sk[109]) & (!ax21x) & (!g6) & (ax20x) & (g8)) + ((!ax22x) & (!sk[109]) & (!ax21x) & (g6) & (ax20x) & (!g8)) + ((!ax22x) & (!sk[109]) & (!ax21x) & (g6) & (ax20x) & (g8)) + ((!ax22x) & (!sk[109]) & (ax21x) & (!g6) & (!ax20x) & (!g8)) + ((!ax22x) & (!sk[109]) & (ax21x) & (!g6) & (!ax20x) & (g8)) + ((!ax22x) & (!sk[109]) & (ax21x) & (!g6) & (ax20x) & (!g8)) + ((!ax22x) & (!sk[109]) & (ax21x) & (!g6) & (ax20x) & (g8)) + ((!ax22x) & (!sk[109]) & (ax21x) & (g6) & (!ax20x) & (!g8)) + ((!ax22x) & (!sk[109]) & (ax21x) & (g6) & (!ax20x) & (g8)) + ((!ax22x) & (!sk[109]) & (ax21x) & (g6) & (ax20x) & (!g8)) + ((!ax22x) & (!sk[109]) & (ax21x) & (g6) & (ax20x) & (g8)) + ((!ax22x) & (sk[109]) & (ax21x) & (!g6) & (!ax20x) & (!g8)) + ((!ax22x) & (sk[109]) & (ax21x) & (g6) & (ax20x) & (!g8)) + ((ax22x) & (!sk[109]) & (!ax21x) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (!sk[109]) & (!ax21x) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (!sk[109]) & (!ax21x) & (g6) & (!ax20x) & (!g8)) + ((ax22x) & (!sk[109]) & (!ax21x) & (g6) & (!ax20x) & (g8)) + ((ax22x) & (!sk[109]) & (!ax21x) & (g6) & (ax20x) & (!g8)) + ((ax22x) & (!sk[109]) & (!ax21x) & (g6) & (ax20x) & (g8)) + ((ax22x) & (!sk[109]) & (ax21x) & (!g6) & (!ax20x) & (!g8)) + ((ax22x) & (!sk[109]) & (ax21x) & (!g6) & (!ax20x) & (g8)) + ((ax22x) & (!sk[109]) & (ax21x) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (!sk[109]) & (ax21x) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (!sk[109]) & (ax21x) & (g6) & (!ax20x) & (!g8)) + ((ax22x) & (!sk[109]) & (ax21x) & (g6) & (!ax20x) & (g8)) + ((ax22x) & (!sk[109]) & (ax21x) & (g6) & (ax20x) & (!g8)) + ((ax22x) & (!sk[109]) & (ax21x) & (g6) & (ax20x) & (g8)) + ((ax22x) & (sk[109]) & (!ax21x) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (sk[109]) & (!ax21x) & (g6) & (ax20x) & (!g8)));
	assign g100 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)));
	assign g101 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8) & (g41)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g41)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g41)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8) & (g41)));
	assign g102 = (((!g97) & (!g98) & (!g99) & (!g100) & (!g62) & (!g101)) + ((!g97) & (!g98) & (!g99) & (!g100) & (g62) & (!g101)) + ((!g97) & (!g98) & (!g99) & (g100) & (!g62) & (!g101)) + ((!g97) & (!g98) & (!g99) & (g100) & (g62) & (!g101)) + ((!g97) & (!g98) & (g99) & (!g100) & (!g62) & (!g101)) + ((!g97) & (!g98) & (g99) & (!g100) & (g62) & (!g101)) + ((!g97) & (!g98) & (g99) & (g100) & (!g62) & (!g101)) + ((!g97) & (!g98) & (g99) & (g100) & (g62) & (!g101)) + ((!g97) & (g98) & (!g99) & (!g100) & (!g62) & (!g101)) + ((!g97) & (g98) & (!g99) & (!g100) & (g62) & (!g101)) + ((!g97) & (g98) & (!g99) & (g100) & (!g62) & (!g101)) + ((!g97) & (g98) & (g99) & (!g100) & (!g62) & (!g101)) + ((!g97) & (g98) & (g99) & (!g100) & (g62) & (!g101)) + ((g97) & (!g98) & (!g99) & (!g100) & (!g62) & (!g101)) + ((g97) & (!g98) & (!g99) & (!g100) & (g62) & (!g101)) + ((g97) & (!g98) & (!g99) & (g100) & (!g62) & (!g101)) + ((g97) & (!g98) & (!g99) & (g100) & (g62) & (!g101)) + ((g97) & (!g98) & (g99) & (!g100) & (!g62) & (!g101)) + ((g97) & (!g98) & (g99) & (!g100) & (g62) & (!g101)) + ((g97) & (g98) & (!g99) & (!g100) & (!g62) & (!g101)) + ((g97) & (g98) & (!g99) & (!g100) & (g62) & (!g101)) + ((g97) & (g98) & (!g99) & (g100) & (!g62) & (!g101)) + ((g97) & (g98) & (g99) & (!g100) & (!g62) & (!g101)) + ((g97) & (g98) & (g99) & (!g100) & (g62) & (!g101)) + ((g97) & (g98) & (g99) & (g100) & (!g62) & (!g101)));
	assign g103 = (((!g9) & (!g10) & (!g99) & (!sk[113]) & (g12) & (!g20)) + ((!g9) & (!g10) & (!g99) & (!sk[113]) & (g12) & (g20)) + ((!g9) & (!g10) & (!g99) & (sk[113]) & (!g12) & (!g20)) + ((!g9) & (!g10) & (!g99) & (sk[113]) & (!g12) & (g20)) + ((!g9) & (!g10) & (!g99) & (sk[113]) & (g12) & (!g20)) + ((!g9) & (!g10) & (!g99) & (sk[113]) & (g12) & (g20)) + ((!g9) & (!g10) & (g99) & (!sk[113]) & (g12) & (!g20)) + ((!g9) & (!g10) & (g99) & (!sk[113]) & (g12) & (g20)) + ((!g9) & (!g10) & (g99) & (sk[113]) & (!g12) & (!g20)) + ((!g9) & (!g10) & (g99) & (sk[113]) & (!g12) & (g20)) + ((!g9) & (!g10) & (g99) & (sk[113]) & (g12) & (!g20)) + ((!g9) & (!g10) & (g99) & (sk[113]) & (g12) & (g20)) + ((!g9) & (g10) & (!g99) & (!sk[113]) & (!g12) & (!g20)) + ((!g9) & (g10) & (!g99) & (!sk[113]) & (!g12) & (g20)) + ((!g9) & (g10) & (!g99) & (!sk[113]) & (g12) & (!g20)) + ((!g9) & (g10) & (!g99) & (!sk[113]) & (g12) & (g20)) + ((!g9) & (g10) & (!g99) & (sk[113]) & (!g12) & (!g20)) + ((!g9) & (g10) & (!g99) & (sk[113]) & (!g12) & (g20)) + ((!g9) & (g10) & (!g99) & (sk[113]) & (g12) & (!g20)) + ((!g9) & (g10) & (!g99) & (sk[113]) & (g12) & (g20)) + ((!g9) & (g10) & (g99) & (!sk[113]) & (!g12) & (!g20)) + ((!g9) & (g10) & (g99) & (!sk[113]) & (!g12) & (g20)) + ((!g9) & (g10) & (g99) & (!sk[113]) & (g12) & (!g20)) + ((!g9) & (g10) & (g99) & (!sk[113]) & (g12) & (g20)) + ((g9) & (!g10) & (!g99) & (!sk[113]) & (g12) & (!g20)) + ((g9) & (!g10) & (!g99) & (!sk[113]) & (g12) & (g20)) + ((g9) & (!g10) & (!g99) & (sk[113]) & (!g12) & (!g20)) + ((g9) & (!g10) & (g99) & (!sk[113]) & (!g12) & (!g20)) + ((g9) & (!g10) & (g99) & (!sk[113]) & (!g12) & (g20)) + ((g9) & (!g10) & (g99) & (!sk[113]) & (g12) & (!g20)) + ((g9) & (!g10) & (g99) & (!sk[113]) & (g12) & (g20)) + ((g9) & (!g10) & (g99) & (sk[113]) & (!g12) & (!g20)) + ((g9) & (g10) & (!g99) & (!sk[113]) & (!g12) & (!g20)) + ((g9) & (g10) & (!g99) & (!sk[113]) & (!g12) & (g20)) + ((g9) & (g10) & (!g99) & (!sk[113]) & (g12) & (!g20)) + ((g9) & (g10) & (!g99) & (!sk[113]) & (g12) & (g20)) + ((g9) & (g10) & (!g99) & (sk[113]) & (!g12) & (!g20)) + ((g9) & (g10) & (g99) & (!sk[113]) & (!g12) & (!g20)) + ((g9) & (g10) & (g99) & (!sk[113]) & (!g12) & (g20)) + ((g9) & (g10) & (g99) & (!sk[113]) & (g12) & (!g20)) + ((g9) & (g10) & (g99) & (!sk[113]) & (g12) & (g20)));
	assign g104 = (((!ax22x) & (!sk[114]) & (!ax21x) & (!g6) & (ax20x) & (!g8)) + ((!ax22x) & (!sk[114]) & (!ax21x) & (!g6) & (ax20x) & (g8)) + ((!ax22x) & (!sk[114]) & (!ax21x) & (g6) & (ax20x) & (!g8)) + ((!ax22x) & (!sk[114]) & (!ax21x) & (g6) & (ax20x) & (g8)) + ((!ax22x) & (!sk[114]) & (ax21x) & (!g6) & (!ax20x) & (!g8)) + ((!ax22x) & (!sk[114]) & (ax21x) & (!g6) & (!ax20x) & (g8)) + ((!ax22x) & (!sk[114]) & (ax21x) & (!g6) & (ax20x) & (!g8)) + ((!ax22x) & (!sk[114]) & (ax21x) & (!g6) & (ax20x) & (g8)) + ((!ax22x) & (!sk[114]) & (ax21x) & (g6) & (!ax20x) & (!g8)) + ((!ax22x) & (!sk[114]) & (ax21x) & (g6) & (!ax20x) & (g8)) + ((!ax22x) & (!sk[114]) & (ax21x) & (g6) & (ax20x) & (!g8)) + ((!ax22x) & (!sk[114]) & (ax21x) & (g6) & (ax20x) & (g8)) + ((!ax22x) & (sk[114]) & (!ax21x) & (g6) & (!ax20x) & (!g8)) + ((!ax22x) & (sk[114]) & (ax21x) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (!sk[114]) & (!ax21x) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (!sk[114]) & (!ax21x) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (!sk[114]) & (!ax21x) & (g6) & (!ax20x) & (!g8)) + ((ax22x) & (!sk[114]) & (!ax21x) & (g6) & (!ax20x) & (g8)) + ((ax22x) & (!sk[114]) & (!ax21x) & (g6) & (ax20x) & (!g8)) + ((ax22x) & (!sk[114]) & (!ax21x) & (g6) & (ax20x) & (g8)) + ((ax22x) & (!sk[114]) & (ax21x) & (!g6) & (!ax20x) & (!g8)) + ((ax22x) & (!sk[114]) & (ax21x) & (!g6) & (!ax20x) & (g8)) + ((ax22x) & (!sk[114]) & (ax21x) & (!g6) & (ax20x) & (!g8)) + ((ax22x) & (!sk[114]) & (ax21x) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (!sk[114]) & (ax21x) & (g6) & (!ax20x) & (!g8)) + ((ax22x) & (!sk[114]) & (ax21x) & (g6) & (!ax20x) & (g8)) + ((ax22x) & (!sk[114]) & (ax21x) & (g6) & (ax20x) & (!g8)) + ((ax22x) & (!sk[114]) & (ax21x) & (g6) & (ax20x) & (g8)) + ((ax22x) & (sk[114]) & (!ax21x) & (!g6) & (!ax20x) & (!g8)) + ((ax22x) & (sk[114]) & (!ax21x) & (g6) & (!ax20x) & (!g8)));
	assign g105 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g66)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g66)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g66)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g66)));
	assign g106 = (((!g38) & (!g70) & (!g104) & (sk[116]) & (!g105)) + ((!g38) & (!g70) & (g104) & (!sk[116]) & (!g105)) + ((!g38) & (!g70) & (g104) & (!sk[116]) & (g105)) + ((!g38) & (!g70) & (g104) & (sk[116]) & (!g105)) + ((!g38) & (g70) & (!g104) & (sk[116]) & (!g105)) + ((!g38) & (g70) & (g104) & (!sk[116]) & (!g105)) + ((!g38) & (g70) & (g104) & (!sk[116]) & (g105)) + ((!g38) & (g70) & (g104) & (sk[116]) & (!g105)) + ((g38) & (!g70) & (!g104) & (!sk[116]) & (!g105)) + ((g38) & (!g70) & (!g104) & (!sk[116]) & (g105)) + ((g38) & (!g70) & (!g104) & (sk[116]) & (!g105)) + ((g38) & (!g70) & (g104) & (!sk[116]) & (!g105)) + ((g38) & (!g70) & (g104) & (!sk[116]) & (g105)) + ((g38) & (g70) & (!g104) & (!sk[116]) & (!g105)) + ((g38) & (g70) & (!g104) & (!sk[116]) & (g105)) + ((g38) & (g70) & (g104) & (!sk[116]) & (!g105)) + ((g38) & (g70) & (g104) & (!sk[116]) & (g105)));
	assign g107 = (((g92) & (g94) & (g96) & (g102) & (g103) & (g106)));
	assign g108 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8) & (g40)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g40)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g40)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8) & (g40)));
	assign g109 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)));
	assign g110 = (((!g99) & (!g30) & (!g18) & (!g104) & (!g25) & (!g32)) + ((!g99) & (!g30) & (!g18) & (!g104) & (!g25) & (g32)) + ((!g99) & (!g30) & (!g18) & (!g104) & (g25) & (!g32)) + ((!g99) & (!g30) & (!g18) & (!g104) & (g25) & (g32)) + ((!g99) & (!g30) & (!g18) & (g104) & (!g25) & (!g32)) + ((!g99) & (!g30) & (g18) & (!g104) & (!g25) & (!g32)) + ((!g99) & (!g30) & (g18) & (!g104) & (!g25) & (g32)) + ((!g99) & (!g30) & (g18) & (!g104) & (g25) & (!g32)) + ((!g99) & (!g30) & (g18) & (!g104) & (g25) & (g32)) + ((!g99) & (!g30) & (g18) & (g104) & (!g25) & (!g32)) + ((!g99) & (g30) & (!g18) & (!g104) & (!g25) & (!g32)) + ((!g99) & (g30) & (!g18) & (!g104) & (!g25) & (g32)) + ((!g99) & (g30) & (!g18) & (!g104) & (g25) & (!g32)) + ((!g99) & (g30) & (!g18) & (!g104) & (g25) & (g32)) + ((!g99) & (g30) & (!g18) & (g104) & (!g25) & (!g32)) + ((!g99) & (g30) & (g18) & (!g104) & (!g25) & (!g32)) + ((!g99) & (g30) & (g18) & (!g104) & (!g25) & (g32)) + ((!g99) & (g30) & (g18) & (!g104) & (g25) & (!g32)) + ((!g99) & (g30) & (g18) & (!g104) & (g25) & (g32)) + ((!g99) & (g30) & (g18) & (g104) & (!g25) & (!g32)) + ((g99) & (!g30) & (!g18) & (!g104) & (!g25) & (!g32)) + ((g99) & (!g30) & (!g18) & (!g104) & (!g25) & (g32)) + ((g99) & (!g30) & (!g18) & (!g104) & (g25) & (!g32)) + ((g99) & (!g30) & (!g18) & (!g104) & (g25) & (g32)) + ((g99) & (!g30) & (!g18) & (g104) & (!g25) & (!g32)));
	assign g111 = (((!g9) & (!g29) & (!sk[121]) & (!g108) & (g109) & (!g110)) + ((!g9) & (!g29) & (!sk[121]) & (!g108) & (g109) & (g110)) + ((!g9) & (!g29) & (!sk[121]) & (g108) & (g109) & (!g110)) + ((!g9) & (!g29) & (!sk[121]) & (g108) & (g109) & (g110)) + ((!g9) & (!g29) & (sk[121]) & (!g108) & (!g109) & (g110)) + ((!g9) & (!g29) & (sk[121]) & (!g108) & (g109) & (g110)) + ((!g9) & (g29) & (!sk[121]) & (!g108) & (!g109) & (!g110)) + ((!g9) & (g29) & (!sk[121]) & (!g108) & (!g109) & (g110)) + ((!g9) & (g29) & (!sk[121]) & (!g108) & (g109) & (!g110)) + ((!g9) & (g29) & (!sk[121]) & (!g108) & (g109) & (g110)) + ((!g9) & (g29) & (!sk[121]) & (g108) & (!g109) & (!g110)) + ((!g9) & (g29) & (!sk[121]) & (g108) & (!g109) & (g110)) + ((!g9) & (g29) & (!sk[121]) & (g108) & (g109) & (!g110)) + ((!g9) & (g29) & (!sk[121]) & (g108) & (g109) & (g110)) + ((g9) & (!g29) & (!sk[121]) & (!g108) & (g109) & (!g110)) + ((g9) & (!g29) & (!sk[121]) & (!g108) & (g109) & (g110)) + ((g9) & (!g29) & (!sk[121]) & (g108) & (!g109) & (!g110)) + ((g9) & (!g29) & (!sk[121]) & (g108) & (!g109) & (g110)) + ((g9) & (!g29) & (!sk[121]) & (g108) & (g109) & (!g110)) + ((g9) & (!g29) & (!sk[121]) & (g108) & (g109) & (g110)) + ((g9) & (!g29) & (sk[121]) & (!g108) & (!g109) & (g110)) + ((g9) & (g29) & (!sk[121]) & (!g108) & (!g109) & (!g110)) + ((g9) & (g29) & (!sk[121]) & (!g108) & (!g109) & (g110)) + ((g9) & (g29) & (!sk[121]) & (!g108) & (g109) & (!g110)) + ((g9) & (g29) & (!sk[121]) & (!g108) & (g109) & (g110)) + ((g9) & (g29) & (!sk[121]) & (g108) & (!g109) & (!g110)) + ((g9) & (g29) & (!sk[121]) & (g108) & (!g109) & (g110)) + ((g9) & (g29) & (!sk[121]) & (g108) & (g109) & (!g110)) + ((g9) & (g29) & (!sk[121]) & (g108) & (g109) & (g110)));
	assign g112 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)));
	assign g113 = (((!ax22x) & (!ax17x) & (!sk[123]) & (!ax16x) & (g5) & (!ax18x)) + ((!ax22x) & (!ax17x) & (!sk[123]) & (!ax16x) & (g5) & (ax18x)) + ((!ax22x) & (!ax17x) & (!sk[123]) & (ax16x) & (g5) & (!ax18x)) + ((!ax22x) & (!ax17x) & (!sk[123]) & (ax16x) & (g5) & (ax18x)) + ((!ax22x) & (!ax17x) & (sk[123]) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax22x) & (!ax17x) & (sk[123]) & (!ax16x) & (g5) & (ax18x)) + ((!ax22x) & (!ax17x) & (sk[123]) & (ax16x) & (!g5) & (!ax18x)) + ((!ax22x) & (!ax17x) & (sk[123]) & (ax16x) & (g5) & (!ax18x)) + ((!ax22x) & (ax17x) & (!sk[123]) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax22x) & (ax17x) & (!sk[123]) & (!ax16x) & (!g5) & (ax18x)) + ((!ax22x) & (ax17x) & (!sk[123]) & (!ax16x) & (g5) & (!ax18x)) + ((!ax22x) & (ax17x) & (!sk[123]) & (!ax16x) & (g5) & (ax18x)) + ((!ax22x) & (ax17x) & (!sk[123]) & (ax16x) & (!g5) & (!ax18x)) + ((!ax22x) & (ax17x) & (!sk[123]) & (ax16x) & (!g5) & (ax18x)) + ((!ax22x) & (ax17x) & (!sk[123]) & (ax16x) & (g5) & (!ax18x)) + ((!ax22x) & (ax17x) & (!sk[123]) & (ax16x) & (g5) & (ax18x)) + ((!ax22x) & (ax17x) & (sk[123]) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax22x) & (ax17x) & (sk[123]) & (!ax16x) & (g5) & (!ax18x)) + ((!ax22x) & (ax17x) & (sk[123]) & (ax16x) & (!g5) & (!ax18x)) + ((!ax22x) & (ax17x) & (sk[123]) & (ax16x) & (g5) & (!ax18x)) + ((ax22x) & (!ax17x) & (!sk[123]) & (!ax16x) & (g5) & (!ax18x)) + ((ax22x) & (!ax17x) & (!sk[123]) & (!ax16x) & (g5) & (ax18x)) + ((ax22x) & (!ax17x) & (!sk[123]) & (ax16x) & (!g5) & (!ax18x)) + ((ax22x) & (!ax17x) & (!sk[123]) & (ax16x) & (!g5) & (ax18x)) + ((ax22x) & (!ax17x) & (!sk[123]) & (ax16x) & (g5) & (!ax18x)) + ((ax22x) & (!ax17x) & (!sk[123]) & (ax16x) & (g5) & (ax18x)) + ((ax22x) & (!ax17x) & (sk[123]) & (!ax16x) & (!g5) & (ax18x)) + ((ax22x) & (!ax17x) & (sk[123]) & (!ax16x) & (g5) & (ax18x)) + ((ax22x) & (!ax17x) & (sk[123]) & (ax16x) & (!g5) & (ax18x)) + ((ax22x) & (!ax17x) & (sk[123]) & (ax16x) & (g5) & (ax18x)) + ((ax22x) & (ax17x) & (!sk[123]) & (!ax16x) & (!g5) & (!ax18x)) + ((ax22x) & (ax17x) & (!sk[123]) & (!ax16x) & (!g5) & (ax18x)) + ((ax22x) & (ax17x) & (!sk[123]) & (!ax16x) & (g5) & (!ax18x)) + ((ax22x) & (ax17x) & (!sk[123]) & (!ax16x) & (g5) & (ax18x)) + ((ax22x) & (ax17x) & (!sk[123]) & (ax16x) & (!g5) & (!ax18x)) + ((ax22x) & (ax17x) & (!sk[123]) & (ax16x) & (!g5) & (ax18x)) + ((ax22x) & (ax17x) & (!sk[123]) & (ax16x) & (g5) & (!ax18x)) + ((ax22x) & (ax17x) & (!sk[123]) & (ax16x) & (g5) & (ax18x)) + ((ax22x) & (ax17x) & (sk[123]) & (!ax16x) & (!g5) & (ax18x)) + ((ax22x) & (ax17x) & (sk[123]) & (!ax16x) & (g5) & (ax18x)) + ((ax22x) & (ax17x) & (sk[123]) & (ax16x) & (!g5) & (ax18x)) + ((ax22x) & (ax17x) & (sk[123]) & (ax16x) & (g5) & (ax18x)));
	assign g114 = (((!ax22x) & (!sk[124]) & (!ax21x) & (g6) & (!ax20x)) + ((!ax22x) & (!sk[124]) & (!ax21x) & (g6) & (ax20x)) + ((!ax22x) & (!sk[124]) & (ax21x) & (g6) & (!ax20x)) + ((!ax22x) & (!sk[124]) & (ax21x) & (g6) & (ax20x)) + ((!ax22x) & (sk[124]) & (!ax21x) & (!g6) & (!ax20x)) + ((!ax22x) & (sk[124]) & (!ax21x) & (!g6) & (ax20x)) + ((!ax22x) & (sk[124]) & (!ax21x) & (g6) & (ax20x)) + ((!ax22x) & (sk[124]) & (ax21x) & (g6) & (!ax20x)) + ((ax22x) & (!sk[124]) & (!ax21x) & (!g6) & (!ax20x)) + ((ax22x) & (!sk[124]) & (!ax21x) & (!g6) & (ax20x)) + ((ax22x) & (!sk[124]) & (!ax21x) & (g6) & (!ax20x)) + ((ax22x) & (!sk[124]) & (!ax21x) & (g6) & (ax20x)) + ((ax22x) & (!sk[124]) & (ax21x) & (!g6) & (!ax20x)) + ((ax22x) & (!sk[124]) & (ax21x) & (!g6) & (ax20x)) + ((ax22x) & (!sk[124]) & (ax21x) & (g6) & (!ax20x)) + ((ax22x) & (!sk[124]) & (ax21x) & (g6) & (ax20x)) + ((ax22x) & (sk[124]) & (ax21x) & (!g6) & (!ax20x)) + ((ax22x) & (sk[124]) & (ax21x) & (!g6) & (ax20x)) + ((ax22x) & (sk[124]) & (ax21x) & (g6) & (!ax20x)) + ((ax22x) & (sk[124]) & (ax21x) & (g6) & (ax20x)));
	assign g115 = (((!ax22x) & (!sk[125]) & (!g6) & (ax20x)) + ((!ax22x) & (!sk[125]) & (g6) & (ax20x)) + ((!ax22x) & (sk[125]) & (!g6) & (!ax20x)) + ((!ax22x) & (sk[125]) & (g6) & (ax20x)) + ((ax22x) & (!sk[125]) & (!g6) & (!ax20x)) + ((ax22x) & (!sk[125]) & (!g6) & (ax20x)) + ((ax22x) & (!sk[125]) & (g6) & (!ax20x)) + ((ax22x) & (!sk[125]) & (g6) & (ax20x)) + ((ax22x) & (sk[125]) & (!g6) & (ax20x)) + ((ax22x) & (sk[125]) & (g6) & (ax20x)));
	assign g116 = (((!ax22x) & (!ax17x) & (!ax16x) & (sk[126]) & (!g5)) + ((!ax22x) & (!ax17x) & (ax16x) & (!sk[126]) & (!g5)) + ((!ax22x) & (!ax17x) & (ax16x) & (!sk[126]) & (g5)) + ((!ax22x) & (!ax17x) & (ax16x) & (sk[126]) & (g5)) + ((!ax22x) & (ax17x) & (ax16x) & (!sk[126]) & (!g5)) + ((!ax22x) & (ax17x) & (ax16x) & (!sk[126]) & (g5)) + ((ax22x) & (!ax17x) & (!ax16x) & (!sk[126]) & (!g5)) + ((ax22x) & (!ax17x) & (!ax16x) & (!sk[126]) & (g5)) + ((ax22x) & (!ax17x) & (ax16x) & (!sk[126]) & (!g5)) + ((ax22x) & (!ax17x) & (ax16x) & (!sk[126]) & (g5)) + ((ax22x) & (ax17x) & (!ax16x) & (!sk[126]) & (!g5)) + ((ax22x) & (ax17x) & (!ax16x) & (!sk[126]) & (g5)) + ((ax22x) & (ax17x) & (ax16x) & (!sk[126]) & (!g5)) + ((ax22x) & (ax17x) & (ax16x) & (!sk[126]) & (g5)) + ((ax22x) & (ax17x) & (ax16x) & (sk[126]) & (!g5)) + ((ax22x) & (ax17x) & (ax16x) & (sk[126]) & (g5)));
	assign g117 = (((!g112) & (!g113) & (!g114) & (g115) & (!g8) & (g116)) + ((!g112) & (g113) & (g114) & (!g115) & (g8) & (g116)) + ((!g112) & (g113) & (g114) & (g115) & (g8) & (g116)) + ((g112) & (!g113) & (!g114) & (!g115) & (!g8) & (g116)) + ((g112) & (!g113) & (!g114) & (g115) & (g8) & (g116)) + ((g112) & (g113) & (!g114) & (!g115) & (g8) & (g116)));
	assign g118 = (((!sk[0]) & (!g30) & (!g62) & (!g46) & (g41) & (!g66)) + ((!sk[0]) & (!g30) & (!g62) & (!g46) & (g41) & (g66)) + ((!sk[0]) & (!g30) & (!g62) & (g46) & (g41) & (!g66)) + ((!sk[0]) & (!g30) & (!g62) & (g46) & (g41) & (g66)) + ((!sk[0]) & (!g30) & (g62) & (!g46) & (!g41) & (!g66)) + ((!sk[0]) & (!g30) & (g62) & (!g46) & (!g41) & (g66)) + ((!sk[0]) & (!g30) & (g62) & (!g46) & (g41) & (!g66)) + ((!sk[0]) & (!g30) & (g62) & (!g46) & (g41) & (g66)) + ((!sk[0]) & (!g30) & (g62) & (g46) & (!g41) & (!g66)) + ((!sk[0]) & (!g30) & (g62) & (g46) & (!g41) & (g66)) + ((!sk[0]) & (!g30) & (g62) & (g46) & (g41) & (!g66)) + ((!sk[0]) & (!g30) & (g62) & (g46) & (g41) & (g66)) + ((!sk[0]) & (g30) & (!g62) & (!g46) & (g41) & (!g66)) + ((!sk[0]) & (g30) & (!g62) & (!g46) & (g41) & (g66)) + ((!sk[0]) & (g30) & (!g62) & (g46) & (!g41) & (!g66)) + ((!sk[0]) & (g30) & (!g62) & (g46) & (!g41) & (g66)) + ((!sk[0]) & (g30) & (!g62) & (g46) & (g41) & (!g66)) + ((!sk[0]) & (g30) & (!g62) & (g46) & (g41) & (g66)) + ((!sk[0]) & (g30) & (g62) & (!g46) & (!g41) & (!g66)) + ((!sk[0]) & (g30) & (g62) & (!g46) & (!g41) & (g66)) + ((!sk[0]) & (g30) & (g62) & (!g46) & (g41) & (!g66)) + ((!sk[0]) & (g30) & (g62) & (!g46) & (g41) & (g66)) + ((!sk[0]) & (g30) & (g62) & (g46) & (!g41) & (!g66)) + ((!sk[0]) & (g30) & (g62) & (g46) & (!g41) & (g66)) + ((!sk[0]) & (g30) & (g62) & (g46) & (g41) & (!g66)) + ((!sk[0]) & (g30) & (g62) & (g46) & (g41) & (g66)) + ((sk[0]) & (!g30) & (!g62) & (!g46) & (!g41) & (!g66)) + ((sk[0]) & (!g30) & (!g62) & (!g46) & (!g41) & (g66)) + ((sk[0]) & (!g30) & (!g62) & (!g46) & (g41) & (!g66)) + ((sk[0]) & (!g30) & (!g62) & (!g46) & (g41) & (g66)) + ((sk[0]) & (!g30) & (!g62) & (g46) & (!g41) & (!g66)) + ((sk[0]) & (!g30) & (!g62) & (g46) & (!g41) & (g66)) + ((sk[0]) & (!g30) & (g62) & (!g46) & (!g41) & (!g66)) + ((sk[0]) & (!g30) & (g62) & (!g46) & (g41) & (!g66)) + ((sk[0]) & (!g30) & (g62) & (g46) & (!g41) & (!g66)) + ((sk[0]) & (g30) & (!g62) & (!g46) & (!g41) & (!g66)) + ((sk[0]) & (g30) & (!g62) & (!g46) & (!g41) & (g66)) + ((sk[0]) & (g30) & (!g62) & (!g46) & (g41) & (!g66)) + ((sk[0]) & (g30) & (!g62) & (!g46) & (g41) & (g66)) + ((sk[0]) & (g30) & (!g62) & (g46) & (!g41) & (!g66)) + ((sk[0]) & (g30) & (!g62) & (g46) & (!g41) & (g66)));
	assign g119 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)));
	assign g120 = (((!g38) & (!g114) & (!g115) & (g8) & (!g10) & (g27)) + ((!g38) & (!g114) & (!g115) & (g8) & (g10) & (g27)) + ((!g38) & (!g114) & (g115) & (g8) & (g10) & (!g27)) + ((!g38) & (!g114) & (g115) & (g8) & (g10) & (g27)) + ((g38) & (!g114) & (!g115) & (g8) & (!g10) & (g27)) + ((g38) & (!g114) & (!g115) & (g8) & (g10) & (g27)) + ((g38) & (!g114) & (g115) & (g8) & (g10) & (!g27)) + ((g38) & (!g114) & (g115) & (g8) & (g10) & (g27)) + ((g38) & (g114) & (!g115) & (!g8) & (!g10) & (!g27)) + ((g38) & (g114) & (!g115) & (!g8) & (!g10) & (g27)) + ((g38) & (g114) & (!g115) & (!g8) & (g10) & (!g27)) + ((g38) & (g114) & (!g115) & (!g8) & (g10) & (g27)) + ((g38) & (g114) & (!g115) & (g8) & (!g10) & (!g27)) + ((g38) & (g114) & (!g115) & (g8) & (!g10) & (g27)) + ((g38) & (g114) & (!g115) & (g8) & (g10) & (!g27)) + ((g38) & (g114) & (!g115) & (g8) & (g10) & (g27)));
	assign g121 = (((!g9) & (!g16) & (!g18) & (g118) & (!g119) & (!g120)) + ((!g9) & (!g16) & (!g18) & (g118) & (g119) & (!g120)) + ((!g9) & (!g16) & (g18) & (g118) & (!g119) & (!g120)) + ((!g9) & (!g16) & (g18) & (g118) & (g119) & (!g120)) + ((!g9) & (g16) & (!g18) & (g118) & (!g119) & (!g120)) + ((!g9) & (g16) & (g18) & (g118) & (!g119) & (!g120)) + ((g9) & (!g16) & (!g18) & (g118) & (!g119) & (!g120)) + ((g9) & (!g16) & (!g18) & (g118) & (g119) & (!g120)) + ((g9) & (g16) & (!g18) & (g118) & (!g119) & (!g120)));
	assign g122 = (((!g89) & (!sk[4]) & (!g107) & (!g111) & (g117) & (!g121)) + ((!g89) & (!sk[4]) & (!g107) & (!g111) & (g117) & (g121)) + ((!g89) & (!sk[4]) & (!g107) & (g111) & (g117) & (!g121)) + ((!g89) & (!sk[4]) & (!g107) & (g111) & (g117) & (g121)) + ((!g89) & (!sk[4]) & (g107) & (!g111) & (!g117) & (!g121)) + ((!g89) & (!sk[4]) & (g107) & (!g111) & (!g117) & (g121)) + ((!g89) & (!sk[4]) & (g107) & (!g111) & (g117) & (!g121)) + ((!g89) & (!sk[4]) & (g107) & (!g111) & (g117) & (g121)) + ((!g89) & (!sk[4]) & (g107) & (g111) & (!g117) & (!g121)) + ((!g89) & (!sk[4]) & (g107) & (g111) & (!g117) & (g121)) + ((!g89) & (!sk[4]) & (g107) & (g111) & (g117) & (!g121)) + ((!g89) & (!sk[4]) & (g107) & (g111) & (g117) & (g121)) + ((g89) & (!sk[4]) & (!g107) & (!g111) & (g117) & (!g121)) + ((g89) & (!sk[4]) & (!g107) & (!g111) & (g117) & (g121)) + ((g89) & (!sk[4]) & (!g107) & (g111) & (!g117) & (!g121)) + ((g89) & (!sk[4]) & (!g107) & (g111) & (!g117) & (g121)) + ((g89) & (!sk[4]) & (!g107) & (g111) & (g117) & (!g121)) + ((g89) & (!sk[4]) & (!g107) & (g111) & (g117) & (g121)) + ((g89) & (!sk[4]) & (g107) & (!g111) & (!g117) & (!g121)) + ((g89) & (!sk[4]) & (g107) & (!g111) & (!g117) & (g121)) + ((g89) & (!sk[4]) & (g107) & (!g111) & (g117) & (!g121)) + ((g89) & (!sk[4]) & (g107) & (!g111) & (g117) & (g121)) + ((g89) & (!sk[4]) & (g107) & (g111) & (!g117) & (!g121)) + ((g89) & (!sk[4]) & (g107) & (g111) & (!g117) & (g121)) + ((g89) & (!sk[4]) & (g107) & (g111) & (g117) & (!g121)) + ((g89) & (!sk[4]) & (g107) & (g111) & (g117) & (g121)) + ((g89) & (sk[4]) & (g107) & (g111) & (!g117) & (g121)));
	assign g123 = (((!sk[5]) & (!g9) & (!g46) & (!g41) & (g66) & (!g43)) + ((!sk[5]) & (!g9) & (!g46) & (!g41) & (g66) & (g43)) + ((!sk[5]) & (!g9) & (!g46) & (g41) & (g66) & (!g43)) + ((!sk[5]) & (!g9) & (!g46) & (g41) & (g66) & (g43)) + ((!sk[5]) & (!g9) & (g46) & (!g41) & (!g66) & (!g43)) + ((!sk[5]) & (!g9) & (g46) & (!g41) & (!g66) & (g43)) + ((!sk[5]) & (!g9) & (g46) & (!g41) & (g66) & (!g43)) + ((!sk[5]) & (!g9) & (g46) & (!g41) & (g66) & (g43)) + ((!sk[5]) & (!g9) & (g46) & (g41) & (!g66) & (!g43)) + ((!sk[5]) & (!g9) & (g46) & (g41) & (!g66) & (g43)) + ((!sk[5]) & (!g9) & (g46) & (g41) & (g66) & (!g43)) + ((!sk[5]) & (!g9) & (g46) & (g41) & (g66) & (g43)) + ((!sk[5]) & (g9) & (!g46) & (!g41) & (g66) & (!g43)) + ((!sk[5]) & (g9) & (!g46) & (!g41) & (g66) & (g43)) + ((!sk[5]) & (g9) & (!g46) & (g41) & (!g66) & (!g43)) + ((!sk[5]) & (g9) & (!g46) & (g41) & (!g66) & (g43)) + ((!sk[5]) & (g9) & (!g46) & (g41) & (g66) & (!g43)) + ((!sk[5]) & (g9) & (!g46) & (g41) & (g66) & (g43)) + ((!sk[5]) & (g9) & (g46) & (!g41) & (!g66) & (!g43)) + ((!sk[5]) & (g9) & (g46) & (!g41) & (!g66) & (g43)) + ((!sk[5]) & (g9) & (g46) & (!g41) & (g66) & (!g43)) + ((!sk[5]) & (g9) & (g46) & (!g41) & (g66) & (g43)) + ((!sk[5]) & (g9) & (g46) & (g41) & (!g66) & (!g43)) + ((!sk[5]) & (g9) & (g46) & (g41) & (!g66) & (g43)) + ((!sk[5]) & (g9) & (g46) & (g41) & (g66) & (!g43)) + ((!sk[5]) & (g9) & (g46) & (g41) & (g66) & (g43)) + ((sk[5]) & (!g9) & (!g46) & (!g41) & (!g66) & (!g43)) + ((sk[5]) & (!g9) & (!g46) & (!g41) & (g66) & (!g43)) + ((sk[5]) & (!g9) & (!g46) & (g41) & (!g66) & (!g43)) + ((sk[5]) & (!g9) & (!g46) & (g41) & (g66) & (!g43)) + ((sk[5]) & (!g9) & (g46) & (!g41) & (!g66) & (!g43)) + ((sk[5]) & (!g9) & (g46) & (!g41) & (g66) & (!g43)) + ((sk[5]) & (g9) & (!g46) & (!g41) & (!g66) & (!g43)) + ((sk[5]) & (g9) & (!g46) & (g41) & (!g66) & (!g43)) + ((sk[5]) & (g9) & (g46) & (!g41) & (!g66) & (!g43)));
	assign g124 = (((!ax22x) & (g38) & (!ax21x) & (!g6) & (ax20x) & (!g8)) + ((!ax22x) & (g38) & (ax21x) & (g6) & (!ax20x) & (!g8)) + ((ax22x) & (g38) & (ax21x) & (!g6) & (!ax20x) & (!g8)) + ((ax22x) & (g38) & (ax21x) & (g6) & (!ax20x) & (!g8)));
	assign g125 = (((!g70) & (!sk[7]) & (!g16) & (!g12) & (g30) & (!g124)) + ((!g70) & (!sk[7]) & (!g16) & (!g12) & (g30) & (g124)) + ((!g70) & (!sk[7]) & (!g16) & (g12) & (g30) & (!g124)) + ((!g70) & (!sk[7]) & (!g16) & (g12) & (g30) & (g124)) + ((!g70) & (!sk[7]) & (g16) & (!g12) & (!g30) & (!g124)) + ((!g70) & (!sk[7]) & (g16) & (!g12) & (!g30) & (g124)) + ((!g70) & (!sk[7]) & (g16) & (!g12) & (g30) & (!g124)) + ((!g70) & (!sk[7]) & (g16) & (!g12) & (g30) & (g124)) + ((!g70) & (!sk[7]) & (g16) & (g12) & (!g30) & (!g124)) + ((!g70) & (!sk[7]) & (g16) & (g12) & (!g30) & (g124)) + ((!g70) & (!sk[7]) & (g16) & (g12) & (g30) & (!g124)) + ((!g70) & (!sk[7]) & (g16) & (g12) & (g30) & (g124)) + ((!g70) & (sk[7]) & (!g16) & (!g12) & (!g30) & (!g124)) + ((!g70) & (sk[7]) & (!g16) & (!g12) & (g30) & (!g124)) + ((!g70) & (sk[7]) & (!g16) & (g12) & (!g30) & (!g124)) + ((!g70) & (sk[7]) & (!g16) & (g12) & (g30) & (!g124)) + ((!g70) & (sk[7]) & (g16) & (!g12) & (!g30) & (!g124)) + ((!g70) & (sk[7]) & (g16) & (g12) & (!g30) & (!g124)) + ((g70) & (!sk[7]) & (!g16) & (!g12) & (g30) & (!g124)) + ((g70) & (!sk[7]) & (!g16) & (!g12) & (g30) & (g124)) + ((g70) & (!sk[7]) & (!g16) & (g12) & (!g30) & (!g124)) + ((g70) & (!sk[7]) & (!g16) & (g12) & (!g30) & (g124)) + ((g70) & (!sk[7]) & (!g16) & (g12) & (g30) & (!g124)) + ((g70) & (!sk[7]) & (!g16) & (g12) & (g30) & (g124)) + ((g70) & (!sk[7]) & (g16) & (!g12) & (!g30) & (!g124)) + ((g70) & (!sk[7]) & (g16) & (!g12) & (!g30) & (g124)) + ((g70) & (!sk[7]) & (g16) & (!g12) & (g30) & (!g124)) + ((g70) & (!sk[7]) & (g16) & (!g12) & (g30) & (g124)) + ((g70) & (!sk[7]) & (g16) & (g12) & (!g30) & (!g124)) + ((g70) & (!sk[7]) & (g16) & (g12) & (!g30) & (g124)) + ((g70) & (!sk[7]) & (g16) & (g12) & (g30) & (!g124)) + ((g70) & (!sk[7]) & (g16) & (g12) & (g30) & (g124)) + ((g70) & (sk[7]) & (!g16) & (!g12) & (!g30) & (!g124)) + ((g70) & (sk[7]) & (!g16) & (!g12) & (g30) & (!g124)) + ((g70) & (sk[7]) & (g16) & (!g12) & (!g30) & (!g124)));
	assign g126 = (((!sk[8]) & (!g123) & (g125)) + ((!sk[8]) & (g123) & (g125)) + ((sk[8]) & (g123) & (g125)));
	assign g127 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g30)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g30)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g30)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g30)));
	assign g128 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)));
	assign g129 = (((!g128) & (!g97) & (!g98) & (g9) & (!sk[11]) & (!g71)) + ((!g128) & (!g97) & (!g98) & (g9) & (!sk[11]) & (g71)) + ((!g128) & (!g97) & (g98) & (g9) & (!sk[11]) & (!g71)) + ((!g128) & (!g97) & (g98) & (g9) & (!sk[11]) & (g71)) + ((!g128) & (g97) & (!g98) & (!g9) & (!sk[11]) & (!g71)) + ((!g128) & (g97) & (!g98) & (!g9) & (!sk[11]) & (g71)) + ((!g128) & (g97) & (!g98) & (g9) & (!sk[11]) & (!g71)) + ((!g128) & (g97) & (!g98) & (g9) & (!sk[11]) & (g71)) + ((!g128) & (g97) & (g98) & (!g9) & (!sk[11]) & (!g71)) + ((!g128) & (g97) & (g98) & (!g9) & (!sk[11]) & (g71)) + ((!g128) & (g97) & (g98) & (g9) & (!sk[11]) & (!g71)) + ((!g128) & (g97) & (g98) & (g9) & (!sk[11]) & (g71)) + ((g128) & (!g97) & (!g98) & (g9) & (!sk[11]) & (!g71)) + ((g128) & (!g97) & (!g98) & (g9) & (!sk[11]) & (g71)) + ((g128) & (!g97) & (!g98) & (g9) & (sk[11]) & (!g71)) + ((g128) & (!g97) & (!g98) & (g9) & (sk[11]) & (g71)) + ((g128) & (!g97) & (g98) & (!g9) & (!sk[11]) & (!g71)) + ((g128) & (!g97) & (g98) & (!g9) & (!sk[11]) & (g71)) + ((g128) & (!g97) & (g98) & (!g9) & (sk[11]) & (g71)) + ((g128) & (!g97) & (g98) & (g9) & (!sk[11]) & (!g71)) + ((g128) & (!g97) & (g98) & (g9) & (!sk[11]) & (g71)) + ((g128) & (!g97) & (g98) & (g9) & (sk[11]) & (g71)) + ((g128) & (g97) & (!g98) & (!g9) & (!sk[11]) & (!g71)) + ((g128) & (g97) & (!g98) & (!g9) & (!sk[11]) & (g71)) + ((g128) & (g97) & (!g98) & (g9) & (!sk[11]) & (!g71)) + ((g128) & (g97) & (!g98) & (g9) & (!sk[11]) & (g71)) + ((g128) & (g97) & (!g98) & (g9) & (sk[11]) & (!g71)) + ((g128) & (g97) & (!g98) & (g9) & (sk[11]) & (g71)) + ((g128) & (g97) & (g98) & (!g9) & (!sk[11]) & (!g71)) + ((g128) & (g97) & (g98) & (!g9) & (!sk[11]) & (g71)) + ((g128) & (g97) & (g98) & (g9) & (!sk[11]) & (!g71)) + ((g128) & (g97) & (g98) & (g9) & (!sk[11]) & (g71)) + ((g128) & (g97) & (g98) & (g9) & (sk[11]) & (!g71)) + ((g128) & (g97) & (g98) & (g9) & (sk[11]) & (g71)));
	assign g130 = (((!sk[12]) & (!g90) & (g11)) + ((!sk[12]) & (g90) & (g11)) + ((sk[12]) & (!g90) & (!g11)));
	assign g131 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g66)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g66)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g66)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g66)));
	assign g132 = (((!g70) & (!g99) & (!g42) & (!g20) & (!g131) & (!g73)) + ((!g70) & (!g99) & (!g42) & (g20) & (!g131) & (!g73)) + ((!g70) & (!g99) & (g42) & (!g20) & (!g131) & (!g73)) + ((!g70) & (!g99) & (g42) & (g20) & (!g131) & (!g73)) + ((!g70) & (g99) & (!g42) & (!g20) & (!g131) & (!g73)) + ((!g70) & (g99) & (!g42) & (g20) & (!g131) & (!g73)) + ((g70) & (!g99) & (!g42) & (!g20) & (!g131) & (!g73)) + ((g70) & (!g99) & (g42) & (!g20) & (!g131) & (!g73)) + ((g70) & (g99) & (!g42) & (!g20) & (!g131) & (!g73)));
	assign g133 = (((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)));
	assign g134 = (((!g9) & (!g16) & (!g42) & (!g20) & (!g36) & (!g133)) + ((!g9) & (!g16) & (!g42) & (!g20) & (!g36) & (g133)) + ((!g9) & (!g16) & (!g42) & (g20) & (!g36) & (!g133)) + ((!g9) & (!g16) & (!g42) & (g20) & (!g36) & (g133)) + ((!g9) & (!g16) & (g42) & (!g20) & (!g36) & (!g133)) + ((!g9) & (!g16) & (g42) & (!g20) & (!g36) & (g133)) + ((!g9) & (!g16) & (g42) & (g20) & (!g36) & (!g133)) + ((!g9) & (!g16) & (g42) & (g20) & (!g36) & (g133)) + ((!g9) & (g16) & (!g42) & (!g20) & (!g36) & (!g133)) + ((!g9) & (g16) & (!g42) & (!g20) & (!g36) & (g133)) + ((g9) & (!g16) & (!g42) & (!g20) & (!g36) & (!g133)) + ((g9) & (!g16) & (!g42) & (g20) & (!g36) & (!g133)) + ((g9) & (!g16) & (g42) & (!g20) & (!g36) & (!g133)) + ((g9) & (!g16) & (g42) & (g20) & (!g36) & (!g133)) + ((g9) & (g16) & (!g42) & (!g20) & (!g36) & (!g133)));
	assign g135 = (((!g127) & (!g129) & (!g130) & (g132) & (!sk[17]) & (!g134)) + ((!g127) & (!g129) & (!g130) & (g132) & (!sk[17]) & (g134)) + ((!g127) & (!g129) & (g130) & (g132) & (!sk[17]) & (!g134)) + ((!g127) & (!g129) & (g130) & (g132) & (!sk[17]) & (g134)) + ((!g127) & (!g129) & (g130) & (g132) & (sk[17]) & (g134)) + ((!g127) & (g129) & (!g130) & (!g132) & (!sk[17]) & (!g134)) + ((!g127) & (g129) & (!g130) & (!g132) & (!sk[17]) & (g134)) + ((!g127) & (g129) & (!g130) & (g132) & (!sk[17]) & (!g134)) + ((!g127) & (g129) & (!g130) & (g132) & (!sk[17]) & (g134)) + ((!g127) & (g129) & (g130) & (!g132) & (!sk[17]) & (!g134)) + ((!g127) & (g129) & (g130) & (!g132) & (!sk[17]) & (g134)) + ((!g127) & (g129) & (g130) & (g132) & (!sk[17]) & (!g134)) + ((!g127) & (g129) & (g130) & (g132) & (!sk[17]) & (g134)) + ((g127) & (!g129) & (!g130) & (g132) & (!sk[17]) & (!g134)) + ((g127) & (!g129) & (!g130) & (g132) & (!sk[17]) & (g134)) + ((g127) & (!g129) & (g130) & (!g132) & (!sk[17]) & (!g134)) + ((g127) & (!g129) & (g130) & (!g132) & (!sk[17]) & (g134)) + ((g127) & (!g129) & (g130) & (g132) & (!sk[17]) & (!g134)) + ((g127) & (!g129) & (g130) & (g132) & (!sk[17]) & (g134)) + ((g127) & (g129) & (!g130) & (!g132) & (!sk[17]) & (!g134)) + ((g127) & (g129) & (!g130) & (!g132) & (!sk[17]) & (g134)) + ((g127) & (g129) & (!g130) & (g132) & (!sk[17]) & (!g134)) + ((g127) & (g129) & (!g130) & (g132) & (!sk[17]) & (g134)) + ((g127) & (g129) & (g130) & (!g132) & (!sk[17]) & (!g134)) + ((g127) & (g129) & (g130) & (!g132) & (!sk[17]) & (g134)) + ((g127) & (g129) & (g130) & (g132) & (!sk[17]) & (!g134)) + ((g127) & (g129) & (g130) & (g132) & (!sk[17]) & (g134)));
	assign g136 = (((!g16) & (!g58) & (!g25) & (!sk[18]) & (g55) & (!g95)) + ((!g16) & (!g58) & (!g25) & (!sk[18]) & (g55) & (g95)) + ((!g16) & (!g58) & (!g25) & (sk[18]) & (!g55) & (!g95)) + ((!g16) & (!g58) & (g25) & (!sk[18]) & (g55) & (!g95)) + ((!g16) & (!g58) & (g25) & (!sk[18]) & (g55) & (g95)) + ((!g16) & (!g58) & (g25) & (sk[18]) & (!g55) & (!g95)) + ((!g16) & (g58) & (!g25) & (!sk[18]) & (!g55) & (!g95)) + ((!g16) & (g58) & (!g25) & (!sk[18]) & (!g55) & (g95)) + ((!g16) & (g58) & (!g25) & (!sk[18]) & (g55) & (!g95)) + ((!g16) & (g58) & (!g25) & (!sk[18]) & (g55) & (g95)) + ((!g16) & (g58) & (!g25) & (sk[18]) & (!g55) & (!g95)) + ((!g16) & (g58) & (g25) & (!sk[18]) & (!g55) & (!g95)) + ((!g16) & (g58) & (g25) & (!sk[18]) & (!g55) & (g95)) + ((!g16) & (g58) & (g25) & (!sk[18]) & (g55) & (!g95)) + ((!g16) & (g58) & (g25) & (!sk[18]) & (g55) & (g95)) + ((!g16) & (g58) & (g25) & (sk[18]) & (!g55) & (!g95)) + ((g16) & (!g58) & (!g25) & (!sk[18]) & (g55) & (!g95)) + ((g16) & (!g58) & (!g25) & (!sk[18]) & (g55) & (g95)) + ((g16) & (!g58) & (!g25) & (sk[18]) & (!g55) & (!g95)) + ((g16) & (!g58) & (g25) & (!sk[18]) & (!g55) & (!g95)) + ((g16) & (!g58) & (g25) & (!sk[18]) & (!g55) & (g95)) + ((g16) & (!g58) & (g25) & (!sk[18]) & (g55) & (!g95)) + ((g16) & (!g58) & (g25) & (!sk[18]) & (g55) & (g95)) + ((g16) & (g58) & (!g25) & (!sk[18]) & (!g55) & (!g95)) + ((g16) & (g58) & (!g25) & (!sk[18]) & (!g55) & (g95)) + ((g16) & (g58) & (!g25) & (!sk[18]) & (g55) & (!g95)) + ((g16) & (g58) & (!g25) & (!sk[18]) & (g55) & (g95)) + ((g16) & (g58) & (g25) & (!sk[18]) & (!g55) & (!g95)) + ((g16) & (g58) & (g25) & (!sk[18]) & (!g55) & (g95)) + ((g16) & (g58) & (g25) & (!sk[18]) & (g55) & (!g95)) + ((g16) & (g58) & (g25) & (!sk[18]) & (g55) & (g95)));
	assign g137 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g40)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g40)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g40)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g40)));
	assign g138 = (((!g10) & (!g17) & (!g99) & (!g12) & (!g46) & (!g137)) + ((!g10) & (!g17) & (!g99) & (!g12) & (g46) & (!g137)) + ((!g10) & (!g17) & (!g99) & (g12) & (!g46) & (!g137)) + ((!g10) & (!g17) & (!g99) & (g12) & (g46) & (!g137)) + ((!g10) & (!g17) & (g99) & (!g12) & (!g46) & (!g137)) + ((!g10) & (!g17) & (g99) & (!g12) & (g46) & (!g137)) + ((!g10) & (g17) & (!g99) & (!g12) & (!g46) & (!g137)) + ((!g10) & (g17) & (!g99) & (g12) & (!g46) & (!g137)) + ((!g10) & (g17) & (g99) & (!g12) & (!g46) & (!g137)) + ((g10) & (!g17) & (!g99) & (!g12) & (!g46) & (!g137)) + ((g10) & (!g17) & (!g99) & (g12) & (!g46) & (!g137)) + ((g10) & (!g17) & (g99) & (!g12) & (!g46) & (!g137)) + ((g10) & (g17) & (!g99) & (!g12) & (!g46) & (!g137)) + ((g10) & (g17) & (!g99) & (g12) & (!g46) & (!g137)) + ((g10) & (g17) & (g99) & (!g12) & (!g46) & (!g137)));
	assign g139 = (((!sk[21]) & (!g49) & (!g62) & (g46) & (!g18)) + ((!sk[21]) & (!g49) & (!g62) & (g46) & (g18)) + ((!sk[21]) & (!g49) & (g62) & (g46) & (!g18)) + ((!sk[21]) & (!g49) & (g62) & (g46) & (g18)) + ((!sk[21]) & (g49) & (!g62) & (!g46) & (!g18)) + ((!sk[21]) & (g49) & (!g62) & (!g46) & (g18)) + ((!sk[21]) & (g49) & (!g62) & (g46) & (!g18)) + ((!sk[21]) & (g49) & (!g62) & (g46) & (g18)) + ((!sk[21]) & (g49) & (g62) & (!g46) & (!g18)) + ((!sk[21]) & (g49) & (g62) & (!g46) & (g18)) + ((!sk[21]) & (g49) & (g62) & (g46) & (!g18)) + ((!sk[21]) & (g49) & (g62) & (g46) & (g18)) + ((sk[21]) & (!g49) & (g62) & (!g46) & (g18)) + ((sk[21]) & (!g49) & (g62) & (g46) & (g18)) + ((sk[21]) & (g49) & (!g62) & (g46) & (!g18)) + ((sk[21]) & (g49) & (!g62) & (g46) & (g18)) + ((sk[21]) & (g49) & (g62) & (!g46) & (g18)) + ((sk[21]) & (g49) & (g62) & (g46) & (!g18)) + ((sk[21]) & (g49) & (g62) & (g46) & (g18)));
	assign g140 = (((!g9) & (!sk[22]) & (!g30) & (!g87) & (g138) & (!g139)) + ((!g9) & (!sk[22]) & (!g30) & (!g87) & (g138) & (g139)) + ((!g9) & (!sk[22]) & (!g30) & (g87) & (g138) & (!g139)) + ((!g9) & (!sk[22]) & (!g30) & (g87) & (g138) & (g139)) + ((!g9) & (!sk[22]) & (g30) & (!g87) & (!g138) & (!g139)) + ((!g9) & (!sk[22]) & (g30) & (!g87) & (!g138) & (g139)) + ((!g9) & (!sk[22]) & (g30) & (!g87) & (g138) & (!g139)) + ((!g9) & (!sk[22]) & (g30) & (!g87) & (g138) & (g139)) + ((!g9) & (!sk[22]) & (g30) & (g87) & (!g138) & (!g139)) + ((!g9) & (!sk[22]) & (g30) & (g87) & (!g138) & (g139)) + ((!g9) & (!sk[22]) & (g30) & (g87) & (g138) & (!g139)) + ((!g9) & (!sk[22]) & (g30) & (g87) & (g138) & (g139)) + ((!g9) & (sk[22]) & (!g30) & (!g87) & (g138) & (!g139)) + ((!g9) & (sk[22]) & (g30) & (!g87) & (g138) & (!g139)) + ((g9) & (!sk[22]) & (!g30) & (!g87) & (g138) & (!g139)) + ((g9) & (!sk[22]) & (!g30) & (!g87) & (g138) & (g139)) + ((g9) & (!sk[22]) & (!g30) & (g87) & (!g138) & (!g139)) + ((g9) & (!sk[22]) & (!g30) & (g87) & (!g138) & (g139)) + ((g9) & (!sk[22]) & (!g30) & (g87) & (g138) & (!g139)) + ((g9) & (!sk[22]) & (!g30) & (g87) & (g138) & (g139)) + ((g9) & (!sk[22]) & (g30) & (!g87) & (!g138) & (!g139)) + ((g9) & (!sk[22]) & (g30) & (!g87) & (!g138) & (g139)) + ((g9) & (!sk[22]) & (g30) & (!g87) & (g138) & (!g139)) + ((g9) & (!sk[22]) & (g30) & (!g87) & (g138) & (g139)) + ((g9) & (!sk[22]) & (g30) & (g87) & (!g138) & (!g139)) + ((g9) & (!sk[22]) & (g30) & (g87) & (!g138) & (g139)) + ((g9) & (!sk[22]) & (g30) & (g87) & (g138) & (!g139)) + ((g9) & (!sk[22]) & (g30) & (g87) & (g138) & (g139)) + ((g9) & (sk[22]) & (!g30) & (!g87) & (g138) & (!g139)));
	assign g141 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g27)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g27)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g27)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g27)));
	assign g142 = (((!g12) & (!sk[24]) & (!g71) & (g58)) + ((!g12) & (!sk[24]) & (g71) & (g58)) + ((!g12) & (sk[24]) & (g71) & (g58)) + ((g12) & (!sk[24]) & (!g71) & (!g58)) + ((g12) & (!sk[24]) & (!g71) & (g58)) + ((g12) & (!sk[24]) & (g71) & (!g58)) + ((g12) & (!sk[24]) & (g71) & (g58)) + ((g12) & (sk[24]) & (g71) & (!g58)) + ((g12) & (sk[24]) & (g71) & (g58)));
	assign g143 = (((!g62) & (!g27) & (!sk[25]) & (g35)) + ((!g62) & (!g27) & (sk[25]) & (!g35)) + ((!g62) & (g27) & (!sk[25]) & (g35)) + ((!g62) & (g27) & (sk[25]) & (!g35)) + ((g62) & (!g27) & (!sk[25]) & (!g35)) + ((g62) & (!g27) & (!sk[25]) & (g35)) + ((g62) & (!g27) & (sk[25]) & (!g35)) + ((g62) & (g27) & (!sk[25]) & (!g35)) + ((g62) & (g27) & (!sk[25]) & (g35)));
	assign g144 = (((!g38) & (!g16) & (!g17) & (!g99) & (sk[26]) & (!g81)) + ((!g38) & (!g16) & (!g17) & (g99) & (!sk[26]) & (!g81)) + ((!g38) & (!g16) & (!g17) & (g99) & (!sk[26]) & (g81)) + ((!g38) & (!g16) & (!g17) & (g99) & (sk[26]) & (!g81)) + ((!g38) & (!g16) & (g17) & (!g99) & (sk[26]) & (!g81)) + ((!g38) & (!g16) & (g17) & (g99) & (!sk[26]) & (!g81)) + ((!g38) & (!g16) & (g17) & (g99) & (!sk[26]) & (g81)) + ((!g38) & (g16) & (!g17) & (!g99) & (!sk[26]) & (!g81)) + ((!g38) & (g16) & (!g17) & (!g99) & (!sk[26]) & (g81)) + ((!g38) & (g16) & (!g17) & (!g99) & (sk[26]) & (!g81)) + ((!g38) & (g16) & (!g17) & (g99) & (!sk[26]) & (!g81)) + ((!g38) & (g16) & (!g17) & (g99) & (!sk[26]) & (g81)) + ((!g38) & (g16) & (!g17) & (g99) & (sk[26]) & (!g81)) + ((!g38) & (g16) & (g17) & (!g99) & (!sk[26]) & (!g81)) + ((!g38) & (g16) & (g17) & (!g99) & (!sk[26]) & (g81)) + ((!g38) & (g16) & (g17) & (!g99) & (sk[26]) & (!g81)) + ((!g38) & (g16) & (g17) & (g99) & (!sk[26]) & (!g81)) + ((!g38) & (g16) & (g17) & (g99) & (!sk[26]) & (g81)) + ((g38) & (!g16) & (!g17) & (!g99) & (sk[26]) & (!g81)) + ((g38) & (!g16) & (!g17) & (g99) & (!sk[26]) & (!g81)) + ((g38) & (!g16) & (!g17) & (g99) & (!sk[26]) & (g81)) + ((g38) & (!g16) & (!g17) & (g99) & (sk[26]) & (!g81)) + ((g38) & (!g16) & (g17) & (!g99) & (!sk[26]) & (!g81)) + ((g38) & (!g16) & (g17) & (!g99) & (!sk[26]) & (g81)) + ((g38) & (!g16) & (g17) & (!g99) & (sk[26]) & (!g81)) + ((g38) & (!g16) & (g17) & (g99) & (!sk[26]) & (!g81)) + ((g38) & (!g16) & (g17) & (g99) & (!sk[26]) & (g81)) + ((g38) & (g16) & (!g17) & (!g99) & (!sk[26]) & (!g81)) + ((g38) & (g16) & (!g17) & (!g99) & (!sk[26]) & (g81)) + ((g38) & (g16) & (!g17) & (g99) & (!sk[26]) & (!g81)) + ((g38) & (g16) & (!g17) & (g99) & (!sk[26]) & (g81)) + ((g38) & (g16) & (g17) & (!g99) & (!sk[26]) & (!g81)) + ((g38) & (g16) & (g17) & (!g99) & (!sk[26]) & (g81)) + ((g38) & (g16) & (g17) & (g99) & (!sk[26]) & (!g81)) + ((g38) & (g16) & (g17) & (g99) & (!sk[26]) & (g81)));
	assign g145 = (((!g99) & (!g18) & (!g141) & (!g142) & (g143) & (g144)) + ((!g99) & (g18) & (!g141) & (!g142) & (g143) & (g144)) + ((g99) & (!g18) & (!g141) & (!g142) & (g143) & (g144)));
	assign g146 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g58)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g58)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g58)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g58)));
	assign g147 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g27)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g27)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g27)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g27)));
	assign g148 = (((!g58) & (!g104) & (!sk[30]) & (g147)) + ((!g58) & (!g104) & (sk[30]) & (!g147)) + ((!g58) & (g104) & (!sk[30]) & (g147)) + ((!g58) & (g104) & (sk[30]) & (!g147)) + ((g58) & (!g104) & (!sk[30]) & (!g147)) + ((g58) & (!g104) & (!sk[30]) & (g147)) + ((g58) & (!g104) & (sk[30]) & (!g147)) + ((g58) & (g104) & (!sk[30]) & (!g147)) + ((g58) & (g104) & (!sk[30]) & (g147)));
	assign g149 = (((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)));
	assign g150 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g149)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g149)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g149)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g149)));
	assign g151 = (((!g38) & (!g70) & (!g17) & (!g99) & (!g40) & (!g150)) + ((!g38) & (!g70) & (!g17) & (!g99) & (g40) & (!g150)) + ((!g38) & (!g70) & (!g17) & (g99) & (!g40) & (!g150)) + ((!g38) & (!g70) & (g17) & (!g99) & (!g40) & (!g150)) + ((!g38) & (!g70) & (g17) & (!g99) & (g40) & (!g150)) + ((!g38) & (!g70) & (g17) & (g99) & (!g40) & (!g150)) + ((!g38) & (g70) & (!g17) & (!g99) & (!g40) & (!g150)) + ((!g38) & (g70) & (!g17) & (!g99) & (g40) & (!g150)) + ((!g38) & (g70) & (!g17) & (g99) & (!g40) & (!g150)) + ((g38) & (!g70) & (!g17) & (!g99) & (!g40) & (!g150)) + ((g38) & (!g70) & (!g17) & (!g99) & (g40) & (!g150)) + ((g38) & (!g70) & (!g17) & (g99) & (!g40) & (!g150)) + ((g38) & (!g70) & (g17) & (!g99) & (!g40) & (!g150)) + ((g38) & (!g70) & (g17) & (!g99) & (g40) & (!g150)) + ((g38) & (!g70) & (g17) & (g99) & (!g40) & (!g150)));
	assign g152 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g10)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g10)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g10)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g10)));
	assign g153 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g58)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g58)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g58)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g58)));
	assign g154 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g42)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g42)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g42)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g42)));
	assign g155 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)));
	assign g156 = (((!g70) & (!g54) & (!g153) & (!g13) & (!g154) & (!g155)) + ((!g70) & (!g54) & (!g153) & (!g13) & (!g154) & (g155)) + ((g70) & (!g54) & (!g153) & (!g13) & (!g154) & (!g155)));
	assign g157 = (((!g38) & (!sk[39]) & (!g62) & (!g104) & (g32) & (!g74)) + ((!g38) & (!sk[39]) & (!g62) & (!g104) & (g32) & (g74)) + ((!g38) & (!sk[39]) & (!g62) & (g104) & (g32) & (!g74)) + ((!g38) & (!sk[39]) & (!g62) & (g104) & (g32) & (g74)) + ((!g38) & (!sk[39]) & (g62) & (!g104) & (!g32) & (!g74)) + ((!g38) & (!sk[39]) & (g62) & (!g104) & (!g32) & (g74)) + ((!g38) & (!sk[39]) & (g62) & (!g104) & (g32) & (!g74)) + ((!g38) & (!sk[39]) & (g62) & (!g104) & (g32) & (g74)) + ((!g38) & (!sk[39]) & (g62) & (g104) & (!g32) & (!g74)) + ((!g38) & (!sk[39]) & (g62) & (g104) & (!g32) & (g74)) + ((!g38) & (!sk[39]) & (g62) & (g104) & (g32) & (!g74)) + ((!g38) & (!sk[39]) & (g62) & (g104) & (g32) & (g74)) + ((!g38) & (sk[39]) & (!g62) & (!g104) & (!g32) & (!g74)) + ((!g38) & (sk[39]) & (!g62) & (!g104) & (g32) & (!g74)) + ((!g38) & (sk[39]) & (!g62) & (g104) & (!g32) & (!g74)) + ((!g38) & (sk[39]) & (g62) & (!g104) & (!g32) & (!g74)) + ((!g38) & (sk[39]) & (g62) & (!g104) & (g32) & (!g74)) + ((!g38) & (sk[39]) & (g62) & (g104) & (!g32) & (!g74)) + ((g38) & (!sk[39]) & (!g62) & (!g104) & (g32) & (!g74)) + ((g38) & (!sk[39]) & (!g62) & (!g104) & (g32) & (g74)) + ((g38) & (!sk[39]) & (!g62) & (g104) & (!g32) & (!g74)) + ((g38) & (!sk[39]) & (!g62) & (g104) & (!g32) & (g74)) + ((g38) & (!sk[39]) & (!g62) & (g104) & (g32) & (!g74)) + ((g38) & (!sk[39]) & (!g62) & (g104) & (g32) & (g74)) + ((g38) & (!sk[39]) & (g62) & (!g104) & (!g32) & (!g74)) + ((g38) & (!sk[39]) & (g62) & (!g104) & (!g32) & (g74)) + ((g38) & (!sk[39]) & (g62) & (!g104) & (g32) & (!g74)) + ((g38) & (!sk[39]) & (g62) & (!g104) & (g32) & (g74)) + ((g38) & (!sk[39]) & (g62) & (g104) & (!g32) & (!g74)) + ((g38) & (!sk[39]) & (g62) & (g104) & (!g32) & (g74)) + ((g38) & (!sk[39]) & (g62) & (g104) & (g32) & (!g74)) + ((g38) & (!sk[39]) & (g62) & (g104) & (g32) & (g74)) + ((g38) & (sk[39]) & (!g62) & (!g104) & (!g32) & (!g74)) + ((g38) & (sk[39]) & (!g62) & (!g104) & (g32) & (!g74)) + ((g38) & (sk[39]) & (!g62) & (g104) & (!g32) & (!g74)));
	assign g158 = (((!g146) & (g148) & (g151) & (!g152) & (g156) & (g157)));
	assign g159 = (((g126) & (g135) & (g136) & (g140) & (g145) & (g158)));
	assign g160 = (((!sk[42]) & (!g78) & (g13)) + ((!sk[42]) & (g78) & (g13)) + ((sk[42]) & (!g78) & (!g13)));
	assign g161 = (((!sk[43]) & (!g16) & (!g99) & (g12) & (!g30)) + ((!sk[43]) & (!g16) & (!g99) & (g12) & (g30)) + ((!sk[43]) & (!g16) & (g99) & (g12) & (!g30)) + ((!sk[43]) & (!g16) & (g99) & (g12) & (g30)) + ((!sk[43]) & (g16) & (!g99) & (!g12) & (!g30)) + ((!sk[43]) & (g16) & (!g99) & (!g12) & (g30)) + ((!sk[43]) & (g16) & (!g99) & (g12) & (!g30)) + ((!sk[43]) & (g16) & (!g99) & (g12) & (g30)) + ((!sk[43]) & (g16) & (g99) & (!g12) & (!g30)) + ((!sk[43]) & (g16) & (g99) & (!g12) & (g30)) + ((!sk[43]) & (g16) & (g99) & (g12) & (!g30)) + ((!sk[43]) & (g16) & (g99) & (g12) & (g30)) + ((sk[43]) & (!g16) & (g99) & (g12) & (!g30)) + ((sk[43]) & (!g16) & (g99) & (g12) & (g30)) + ((sk[43]) & (g16) & (!g99) & (!g12) & (g30)) + ((sk[43]) & (g16) & (!g99) & (g12) & (g30)) + ((sk[43]) & (g16) & (g99) & (!g12) & (g30)) + ((sk[43]) & (g16) & (g99) & (g12) & (!g30)) + ((sk[43]) & (g16) & (g99) & (g12) & (g30)));
	assign g162 = (((!sk[44]) & (!g9) & (!g17) & (g12) & (!g46)) + ((!sk[44]) & (!g9) & (!g17) & (g12) & (g46)) + ((!sk[44]) & (!g9) & (g17) & (g12) & (!g46)) + ((!sk[44]) & (!g9) & (g17) & (g12) & (g46)) + ((!sk[44]) & (g9) & (!g17) & (!g12) & (!g46)) + ((!sk[44]) & (g9) & (!g17) & (!g12) & (g46)) + ((!sk[44]) & (g9) & (!g17) & (g12) & (!g46)) + ((!sk[44]) & (g9) & (!g17) & (g12) & (g46)) + ((!sk[44]) & (g9) & (g17) & (!g12) & (!g46)) + ((!sk[44]) & (g9) & (g17) & (!g12) & (g46)) + ((!sk[44]) & (g9) & (g17) & (g12) & (!g46)) + ((!sk[44]) & (g9) & (g17) & (g12) & (g46)) + ((sk[44]) & (!g9) & (g17) & (!g12) & (g46)) + ((sk[44]) & (!g9) & (g17) & (g12) & (g46)) + ((sk[44]) & (g9) & (!g17) & (g12) & (!g46)) + ((sk[44]) & (g9) & (!g17) & (g12) & (g46)) + ((sk[44]) & (g9) & (g17) & (!g12) & (g46)) + ((sk[44]) & (g9) & (g17) & (g12) & (!g46)) + ((sk[44]) & (g9) & (g17) & (g12) & (g46)));
	assign g163 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g17)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g17)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g17)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g17)));
	assign g164 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g32)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g32)) + ((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g32)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g32)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g32)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g32)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g32)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g32)));
	assign g165 = (((!g163) & (!g104) & (!g42) & (!g27) & (!g21) & (!g164)) + ((!g163) & (!g104) & (!g42) & (g27) & (!g21) & (!g164)) + ((!g163) & (!g104) & (g42) & (!g27) & (!g21) & (!g164)) + ((!g163) & (!g104) & (g42) & (g27) & (!g21) & (!g164)) + ((!g163) & (g104) & (!g42) & (!g27) & (!g21) & (!g164)));
	assign g166 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8) & (g27)) + ((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g27)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g27)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g27)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g27)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g27)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (g8) & (g27)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g27)));
	assign g167 = (((!g70) & (!g42) & (!sk[49]) & (g29) & (!g166)) + ((!g70) & (!g42) & (!sk[49]) & (g29) & (g166)) + ((!g70) & (!g42) & (sk[49]) & (!g29) & (!g166)) + ((!g70) & (g42) & (!sk[49]) & (g29) & (!g166)) + ((!g70) & (g42) & (!sk[49]) & (g29) & (g166)) + ((!g70) & (g42) & (sk[49]) & (!g29) & (!g166)) + ((g70) & (!g42) & (!sk[49]) & (!g29) & (!g166)) + ((g70) & (!g42) & (!sk[49]) & (!g29) & (g166)) + ((g70) & (!g42) & (!sk[49]) & (g29) & (!g166)) + ((g70) & (!g42) & (!sk[49]) & (g29) & (g166)) + ((g70) & (!g42) & (sk[49]) & (!g29) & (!g166)) + ((g70) & (g42) & (!sk[49]) & (!g29) & (!g166)) + ((g70) & (g42) & (!sk[49]) & (!g29) & (g166)) + ((g70) & (g42) & (!sk[49]) & (g29) & (!g166)) + ((g70) & (g42) & (!sk[49]) & (g29) & (g166)));
	assign g168 = (((g160) & (!g161) & (!g162) & (g132) & (g165) & (g167)));
	assign g169 = (((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (!ax18x)));
	assign g170 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g169)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g169)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g169)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g169)));
	assign g171 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g42)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g42)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g42)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g42)));
	assign g172 = (((!sk[54]) & (!g38) & (!g9) & (g85) & (!g171)) + ((!sk[54]) & (!g38) & (!g9) & (g85) & (g171)) + ((!sk[54]) & (!g38) & (g9) & (g85) & (!g171)) + ((!sk[54]) & (!g38) & (g9) & (g85) & (g171)) + ((!sk[54]) & (g38) & (!g9) & (!g85) & (!g171)) + ((!sk[54]) & (g38) & (!g9) & (!g85) & (g171)) + ((!sk[54]) & (g38) & (!g9) & (g85) & (!g171)) + ((!sk[54]) & (g38) & (!g9) & (g85) & (g171)) + ((!sk[54]) & (g38) & (g9) & (!g85) & (!g171)) + ((!sk[54]) & (g38) & (g9) & (!g85) & (g171)) + ((!sk[54]) & (g38) & (g9) & (g85) & (!g171)) + ((!sk[54]) & (g38) & (g9) & (g85) & (g171)) + ((sk[54]) & (!g38) & (!g9) & (!g85) & (!g171)) + ((sk[54]) & (!g38) & (g9) & (!g85) & (!g171)) + ((sk[54]) & (g38) & (!g9) & (!g85) & (!g171)));
	assign g173 = (((!g16) & (!g47) & (!g66) & (g52) & (!g170) & (g172)) + ((!g16) & (!g47) & (g66) & (g52) & (!g170) & (g172)) + ((g16) & (!g47) & (!g66) & (g52) & (!g170) & (g172)));
	assign g174 = (((!sk[56]) & (!g70) & (!g17) & (g58)) + ((!sk[56]) & (!g70) & (g17) & (g58)) + ((!sk[56]) & (g70) & (!g17) & (!g58)) + ((!sk[56]) & (g70) & (!g17) & (g58)) + ((!sk[56]) & (g70) & (g17) & (!g58)) + ((!sk[56]) & (g70) & (g17) & (g58)) + ((sk[56]) & (g70) & (!g17) & (g58)) + ((sk[56]) & (g70) & (g17) & (!g58)) + ((sk[56]) & (g70) & (g17) & (g58)));
	assign g175 = (((!g9) & (!g30) & (!g42) & (!g26) & (!g152) & (!g87)) + ((!g9) & (!g30) & (g42) & (!g26) & (!g152) & (!g87)) + ((!g9) & (g30) & (!g42) & (!g26) & (!g152) & (!g87)) + ((!g9) & (g30) & (g42) & (!g26) & (!g152) & (!g87)) + ((g9) & (!g30) & (!g42) & (!g26) & (!g152) & (!g87)));
	assign g176 = (((!g99) & (!sk[58]) & (!g30) & (!g25) & (g93) & (!g137)) + ((!g99) & (!sk[58]) & (!g30) & (!g25) & (g93) & (g137)) + ((!g99) & (!sk[58]) & (!g30) & (g25) & (g93) & (!g137)) + ((!g99) & (!sk[58]) & (!g30) & (g25) & (g93) & (g137)) + ((!g99) & (!sk[58]) & (g30) & (!g25) & (!g93) & (!g137)) + ((!g99) & (!sk[58]) & (g30) & (!g25) & (!g93) & (g137)) + ((!g99) & (!sk[58]) & (g30) & (!g25) & (g93) & (!g137)) + ((!g99) & (!sk[58]) & (g30) & (!g25) & (g93) & (g137)) + ((!g99) & (!sk[58]) & (g30) & (g25) & (!g93) & (!g137)) + ((!g99) & (!sk[58]) & (g30) & (g25) & (!g93) & (g137)) + ((!g99) & (!sk[58]) & (g30) & (g25) & (g93) & (!g137)) + ((!g99) & (!sk[58]) & (g30) & (g25) & (g93) & (g137)) + ((!g99) & (sk[58]) & (!g30) & (!g25) & (!g93) & (!g137)) + ((!g99) & (sk[58]) & (!g30) & (g25) & (!g93) & (!g137)) + ((!g99) & (sk[58]) & (g30) & (!g25) & (!g93) & (!g137)) + ((!g99) & (sk[58]) & (g30) & (g25) & (!g93) & (!g137)) + ((g99) & (!sk[58]) & (!g30) & (!g25) & (g93) & (!g137)) + ((g99) & (!sk[58]) & (!g30) & (!g25) & (g93) & (g137)) + ((g99) & (!sk[58]) & (!g30) & (g25) & (!g93) & (!g137)) + ((g99) & (!sk[58]) & (!g30) & (g25) & (!g93) & (g137)) + ((g99) & (!sk[58]) & (!g30) & (g25) & (g93) & (!g137)) + ((g99) & (!sk[58]) & (!g30) & (g25) & (g93) & (g137)) + ((g99) & (!sk[58]) & (g30) & (!g25) & (!g93) & (!g137)) + ((g99) & (!sk[58]) & (g30) & (!g25) & (!g93) & (g137)) + ((g99) & (!sk[58]) & (g30) & (!g25) & (g93) & (!g137)) + ((g99) & (!sk[58]) & (g30) & (!g25) & (g93) & (g137)) + ((g99) & (!sk[58]) & (g30) & (g25) & (!g93) & (!g137)) + ((g99) & (!sk[58]) & (g30) & (g25) & (!g93) & (g137)) + ((g99) & (!sk[58]) & (g30) & (g25) & (g93) & (!g137)) + ((g99) & (!sk[58]) & (g30) & (g25) & (g93) & (g137)) + ((g99) & (sk[58]) & (!g30) & (!g25) & (!g93) & (!g137)));
	assign g177 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g25)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g25)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g25)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g25)));
	assign g178 = (((!g9) & (!g153) & (!g41) & (!g177) & (!g108) & (!g81)) + ((!g9) & (!g153) & (g41) & (!g177) & (!g108) & (!g81)) + ((g9) & (!g153) & (!g41) & (!g177) & (!g108) & (!g81)));
	assign g179 = (((!g9) & (!g17) & (!g76) & (!g71) & (!g58) & (!g41)) + ((!g9) & (!g17) & (!g76) & (!g71) & (!g58) & (g41)) + ((!g9) & (!g17) & (!g76) & (!g71) & (g58) & (!g41)) + ((!g9) & (!g17) & (!g76) & (!g71) & (g58) & (g41)) + ((!g9) & (!g17) & (!g76) & (g71) & (!g58) & (!g41)) + ((!g9) & (!g17) & (!g76) & (g71) & (g58) & (!g41)) + ((!g9) & (g17) & (!g76) & (!g71) & (!g58) & (!g41)) + ((!g9) & (g17) & (!g76) & (!g71) & (!g58) & (g41)) + ((!g9) & (g17) & (!g76) & (!g71) & (g58) & (!g41)) + ((!g9) & (g17) & (!g76) & (!g71) & (g58) & (g41)) + ((g9) & (!g17) & (!g76) & (!g71) & (!g58) & (!g41)) + ((g9) & (!g17) & (!g76) & (!g71) & (!g58) & (g41)) + ((g9) & (!g17) & (!g76) & (g71) & (!g58) & (!g41)) + ((g9) & (g17) & (!g76) & (!g71) & (!g58) & (!g41)) + ((g9) & (g17) & (!g76) & (!g71) & (!g58) & (g41)));
	assign g180 = (((!sk[62]) & (!g174) & (!g175) & (!g176) & (g178) & (!g179)) + ((!sk[62]) & (!g174) & (!g175) & (!g176) & (g178) & (g179)) + ((!sk[62]) & (!g174) & (!g175) & (g176) & (g178) & (!g179)) + ((!sk[62]) & (!g174) & (!g175) & (g176) & (g178) & (g179)) + ((!sk[62]) & (!g174) & (g175) & (!g176) & (!g178) & (!g179)) + ((!sk[62]) & (!g174) & (g175) & (!g176) & (!g178) & (g179)) + ((!sk[62]) & (!g174) & (g175) & (!g176) & (g178) & (!g179)) + ((!sk[62]) & (!g174) & (g175) & (!g176) & (g178) & (g179)) + ((!sk[62]) & (!g174) & (g175) & (g176) & (!g178) & (!g179)) + ((!sk[62]) & (!g174) & (g175) & (g176) & (!g178) & (g179)) + ((!sk[62]) & (!g174) & (g175) & (g176) & (g178) & (!g179)) + ((!sk[62]) & (!g174) & (g175) & (g176) & (g178) & (g179)) + ((!sk[62]) & (g174) & (!g175) & (!g176) & (g178) & (!g179)) + ((!sk[62]) & (g174) & (!g175) & (!g176) & (g178) & (g179)) + ((!sk[62]) & (g174) & (!g175) & (g176) & (!g178) & (!g179)) + ((!sk[62]) & (g174) & (!g175) & (g176) & (!g178) & (g179)) + ((!sk[62]) & (g174) & (!g175) & (g176) & (g178) & (!g179)) + ((!sk[62]) & (g174) & (!g175) & (g176) & (g178) & (g179)) + ((!sk[62]) & (g174) & (g175) & (!g176) & (!g178) & (!g179)) + ((!sk[62]) & (g174) & (g175) & (!g176) & (!g178) & (g179)) + ((!sk[62]) & (g174) & (g175) & (!g176) & (g178) & (!g179)) + ((!sk[62]) & (g174) & (g175) & (!g176) & (g178) & (g179)) + ((!sk[62]) & (g174) & (g175) & (g176) & (!g178) & (!g179)) + ((!sk[62]) & (g174) & (g175) & (g176) & (!g178) & (g179)) + ((!sk[62]) & (g174) & (g175) & (g176) & (g178) & (!g179)) + ((!sk[62]) & (g174) & (g175) & (g176) & (g178) & (g179)) + ((sk[62]) & (!g174) & (g175) & (g176) & (g178) & (g179)));
	assign g181 = (((!sk[63]) & (!g35) & (g101)) + ((!sk[63]) & (g35) & (g101)) + ((sk[63]) & (!g35) & (!g101)));
	assign g182 = (((!g38) & (!sk[64]) & (!g62) & (g83) & (!g32)) + ((!g38) & (!sk[64]) & (!g62) & (g83) & (g32)) + ((!g38) & (!sk[64]) & (g62) & (g83) & (!g32)) + ((!g38) & (!sk[64]) & (g62) & (g83) & (g32)) + ((!g38) & (sk[64]) & (!g62) & (!g83) & (!g32)) + ((!g38) & (sk[64]) & (!g62) & (!g83) & (g32)) + ((!g38) & (sk[64]) & (g62) & (!g83) & (!g32)) + ((g38) & (!sk[64]) & (!g62) & (!g83) & (!g32)) + ((g38) & (!sk[64]) & (!g62) & (!g83) & (g32)) + ((g38) & (!sk[64]) & (!g62) & (g83) & (!g32)) + ((g38) & (!sk[64]) & (!g62) & (g83) & (g32)) + ((g38) & (!sk[64]) & (g62) & (!g83) & (!g32)) + ((g38) & (!sk[64]) & (g62) & (!g83) & (g32)) + ((g38) & (!sk[64]) & (g62) & (g83) & (!g32)) + ((g38) & (!sk[64]) & (g62) & (g83) & (g32)) + ((g38) & (sk[64]) & (!g62) & (!g83) & (!g32)) + ((g38) & (sk[64]) & (!g62) & (!g83) & (g32)));
	assign g183 = (((!g70) & (!g16) & (!g40) & (!g25) & (g181) & (g182)) + ((!g70) & (!g16) & (!g40) & (g25) & (g181) & (g182)) + ((!g70) & (!g16) & (g40) & (!g25) & (g181) & (g182)) + ((!g70) & (!g16) & (g40) & (g25) & (g181) & (g182)) + ((!g70) & (g16) & (!g40) & (!g25) & (g181) & (g182)) + ((!g70) & (g16) & (!g40) & (g25) & (g181) & (g182)) + ((g70) & (!g16) & (!g40) & (!g25) & (g181) & (g182)) + ((g70) & (!g16) & (g40) & (!g25) & (g181) & (g182)) + ((g70) & (g16) & (!g40) & (!g25) & (g181) & (g182)));
	assign g184 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g58)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g58)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g58)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g58)));
	assign g185 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g41)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g41)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g41)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g41)));
	assign g186 = (((!g16) & (!g42) & (!sk[68]) & (g146)) + ((!g16) & (!g42) & (sk[68]) & (!g146)) + ((!g16) & (g42) & (!sk[68]) & (g146)) + ((!g16) & (g42) & (sk[68]) & (!g146)) + ((g16) & (!g42) & (!sk[68]) & (!g146)) + ((g16) & (!g42) & (!sk[68]) & (g146)) + ((g16) & (!g42) & (sk[68]) & (!g146)) + ((g16) & (g42) & (!sk[68]) & (!g146)) + ((g16) & (g42) & (!sk[68]) & (g146)));
	assign g187 = (((!ax22x) & (g38) & (!ax21x) & (g6) & (!ax20x) & (g8)) + ((!ax22x) & (g38) & (ax21x) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (g38) & (!ax21x) & (!g6) & (!ax20x) & (g8)) + ((ax22x) & (g38) & (!ax21x) & (g6) & (!ax20x) & (g8)));
	assign g188 = (((!g62) & (!g18) & (!g42) & (!sk[70]) & (g11) & (!g187)) + ((!g62) & (!g18) & (!g42) & (!sk[70]) & (g11) & (g187)) + ((!g62) & (!g18) & (!g42) & (sk[70]) & (!g11) & (!g187)) + ((!g62) & (!g18) & (g42) & (!sk[70]) & (g11) & (!g187)) + ((!g62) & (!g18) & (g42) & (!sk[70]) & (g11) & (g187)) + ((!g62) & (!g18) & (g42) & (sk[70]) & (!g11) & (!g187)) + ((!g62) & (g18) & (!g42) & (!sk[70]) & (!g11) & (!g187)) + ((!g62) & (g18) & (!g42) & (!sk[70]) & (!g11) & (g187)) + ((!g62) & (g18) & (!g42) & (!sk[70]) & (g11) & (!g187)) + ((!g62) & (g18) & (!g42) & (!sk[70]) & (g11) & (g187)) + ((!g62) & (g18) & (!g42) & (sk[70]) & (!g11) & (!g187)) + ((!g62) & (g18) & (g42) & (!sk[70]) & (!g11) & (!g187)) + ((!g62) & (g18) & (g42) & (!sk[70]) & (!g11) & (g187)) + ((!g62) & (g18) & (g42) & (!sk[70]) & (g11) & (!g187)) + ((!g62) & (g18) & (g42) & (!sk[70]) & (g11) & (g187)) + ((!g62) & (g18) & (g42) & (sk[70]) & (!g11) & (!g187)) + ((g62) & (!g18) & (!g42) & (!sk[70]) & (g11) & (!g187)) + ((g62) & (!g18) & (!g42) & (!sk[70]) & (g11) & (g187)) + ((g62) & (!g18) & (!g42) & (sk[70]) & (!g11) & (!g187)) + ((g62) & (!g18) & (g42) & (!sk[70]) & (!g11) & (!g187)) + ((g62) & (!g18) & (g42) & (!sk[70]) & (!g11) & (g187)) + ((g62) & (!g18) & (g42) & (!sk[70]) & (g11) & (!g187)) + ((g62) & (!g18) & (g42) & (!sk[70]) & (g11) & (g187)) + ((g62) & (g18) & (!g42) & (!sk[70]) & (!g11) & (!g187)) + ((g62) & (g18) & (!g42) & (!sk[70]) & (!g11) & (g187)) + ((g62) & (g18) & (!g42) & (!sk[70]) & (g11) & (!g187)) + ((g62) & (g18) & (!g42) & (!sk[70]) & (g11) & (g187)) + ((g62) & (g18) & (g42) & (!sk[70]) & (!g11) & (!g187)) + ((g62) & (g18) & (g42) & (!sk[70]) & (!g11) & (g187)) + ((g62) & (g18) & (g42) & (!sk[70]) & (g11) & (!g187)) + ((g62) & (g18) & (g42) & (!sk[70]) & (g11) & (g187)));
	assign g189 = (((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)));
	assign g190 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (g8) & (g189)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g189)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (g8) & (g189)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g189)));
	assign g191 = (((!g104) & (!sk[73]) & (!g40) & (!g20) & (g19) & (!g190)) + ((!g104) & (!sk[73]) & (!g40) & (!g20) & (g19) & (g190)) + ((!g104) & (!sk[73]) & (!g40) & (g20) & (g19) & (!g190)) + ((!g104) & (!sk[73]) & (!g40) & (g20) & (g19) & (g190)) + ((!g104) & (!sk[73]) & (g40) & (!g20) & (!g19) & (!g190)) + ((!g104) & (!sk[73]) & (g40) & (!g20) & (!g19) & (g190)) + ((!g104) & (!sk[73]) & (g40) & (!g20) & (g19) & (!g190)) + ((!g104) & (!sk[73]) & (g40) & (!g20) & (g19) & (g190)) + ((!g104) & (!sk[73]) & (g40) & (g20) & (!g19) & (!g190)) + ((!g104) & (!sk[73]) & (g40) & (g20) & (!g19) & (g190)) + ((!g104) & (!sk[73]) & (g40) & (g20) & (g19) & (!g190)) + ((!g104) & (!sk[73]) & (g40) & (g20) & (g19) & (g190)) + ((!g104) & (sk[73]) & (!g40) & (!g20) & (!g19) & (!g190)) + ((!g104) & (sk[73]) & (!g40) & (g20) & (!g19) & (!g190)) + ((!g104) & (sk[73]) & (g40) & (!g20) & (!g19) & (!g190)) + ((!g104) & (sk[73]) & (g40) & (g20) & (!g19) & (!g190)) + ((g104) & (!sk[73]) & (!g40) & (!g20) & (g19) & (!g190)) + ((g104) & (!sk[73]) & (!g40) & (!g20) & (g19) & (g190)) + ((g104) & (!sk[73]) & (!g40) & (g20) & (!g19) & (!g190)) + ((g104) & (!sk[73]) & (!g40) & (g20) & (!g19) & (g190)) + ((g104) & (!sk[73]) & (!g40) & (g20) & (g19) & (!g190)) + ((g104) & (!sk[73]) & (!g40) & (g20) & (g19) & (g190)) + ((g104) & (!sk[73]) & (g40) & (!g20) & (!g19) & (!g190)) + ((g104) & (!sk[73]) & (g40) & (!g20) & (!g19) & (g190)) + ((g104) & (!sk[73]) & (g40) & (!g20) & (g19) & (!g190)) + ((g104) & (!sk[73]) & (g40) & (!g20) & (g19) & (g190)) + ((g104) & (!sk[73]) & (g40) & (g20) & (!g19) & (!g190)) + ((g104) & (!sk[73]) & (g40) & (g20) & (!g19) & (g190)) + ((g104) & (!sk[73]) & (g40) & (g20) & (g19) & (!g190)) + ((g104) & (!sk[73]) & (g40) & (g20) & (g19) & (g190)) + ((g104) & (sk[73]) & (!g40) & (!g20) & (!g19) & (!g190)));
	assign g192 = (((!g184) & (!g185) & (!g186) & (g188) & (!sk[74]) & (!g191)) + ((!g184) & (!g185) & (!g186) & (g188) & (!sk[74]) & (g191)) + ((!g184) & (!g185) & (g186) & (g188) & (!sk[74]) & (!g191)) + ((!g184) & (!g185) & (g186) & (g188) & (!sk[74]) & (g191)) + ((!g184) & (!g185) & (g186) & (g188) & (sk[74]) & (g191)) + ((!g184) & (g185) & (!g186) & (!g188) & (!sk[74]) & (!g191)) + ((!g184) & (g185) & (!g186) & (!g188) & (!sk[74]) & (g191)) + ((!g184) & (g185) & (!g186) & (g188) & (!sk[74]) & (!g191)) + ((!g184) & (g185) & (!g186) & (g188) & (!sk[74]) & (g191)) + ((!g184) & (g185) & (g186) & (!g188) & (!sk[74]) & (!g191)) + ((!g184) & (g185) & (g186) & (!g188) & (!sk[74]) & (g191)) + ((!g184) & (g185) & (g186) & (g188) & (!sk[74]) & (!g191)) + ((!g184) & (g185) & (g186) & (g188) & (!sk[74]) & (g191)) + ((g184) & (!g185) & (!g186) & (g188) & (!sk[74]) & (!g191)) + ((g184) & (!g185) & (!g186) & (g188) & (!sk[74]) & (g191)) + ((g184) & (!g185) & (g186) & (!g188) & (!sk[74]) & (!g191)) + ((g184) & (!g185) & (g186) & (!g188) & (!sk[74]) & (g191)) + ((g184) & (!g185) & (g186) & (g188) & (!sk[74]) & (!g191)) + ((g184) & (!g185) & (g186) & (g188) & (!sk[74]) & (g191)) + ((g184) & (g185) & (!g186) & (!g188) & (!sk[74]) & (!g191)) + ((g184) & (g185) & (!g186) & (!g188) & (!sk[74]) & (g191)) + ((g184) & (g185) & (!g186) & (g188) & (!sk[74]) & (!g191)) + ((g184) & (g185) & (!g186) & (g188) & (!sk[74]) & (g191)) + ((g184) & (g185) & (g186) & (!g188) & (!sk[74]) & (!g191)) + ((g184) & (g185) & (g186) & (!g188) & (!sk[74]) & (g191)) + ((g184) & (g185) & (g186) & (g188) & (!sk[74]) & (!g191)) + ((g184) & (g185) & (g186) & (g188) & (!sk[74]) & (g191)));
	assign g193 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g18)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g18)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g18)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g18)));
	assign g194 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g41)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g41)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g41)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g41)));
	assign g195 = (((!g62) & (!g104) & (!sk[77]) & (!g66) & (g193) & (!g194)) + ((!g62) & (!g104) & (!sk[77]) & (!g66) & (g193) & (g194)) + ((!g62) & (!g104) & (!sk[77]) & (g66) & (g193) & (!g194)) + ((!g62) & (!g104) & (!sk[77]) & (g66) & (g193) & (g194)) + ((!g62) & (!g104) & (sk[77]) & (!g66) & (!g193) & (!g194)) + ((!g62) & (!g104) & (sk[77]) & (g66) & (!g193) & (!g194)) + ((!g62) & (g104) & (!sk[77]) & (!g66) & (!g193) & (!g194)) + ((!g62) & (g104) & (!sk[77]) & (!g66) & (!g193) & (g194)) + ((!g62) & (g104) & (!sk[77]) & (!g66) & (g193) & (!g194)) + ((!g62) & (g104) & (!sk[77]) & (!g66) & (g193) & (g194)) + ((!g62) & (g104) & (!sk[77]) & (g66) & (!g193) & (!g194)) + ((!g62) & (g104) & (!sk[77]) & (g66) & (!g193) & (g194)) + ((!g62) & (g104) & (!sk[77]) & (g66) & (g193) & (!g194)) + ((!g62) & (g104) & (!sk[77]) & (g66) & (g193) & (g194)) + ((!g62) & (g104) & (sk[77]) & (!g66) & (!g193) & (!g194)) + ((g62) & (!g104) & (!sk[77]) & (!g66) & (g193) & (!g194)) + ((g62) & (!g104) & (!sk[77]) & (!g66) & (g193) & (g194)) + ((g62) & (!g104) & (!sk[77]) & (g66) & (!g193) & (!g194)) + ((g62) & (!g104) & (!sk[77]) & (g66) & (!g193) & (g194)) + ((g62) & (!g104) & (!sk[77]) & (g66) & (g193) & (!g194)) + ((g62) & (!g104) & (!sk[77]) & (g66) & (g193) & (g194)) + ((g62) & (!g104) & (sk[77]) & (!g66) & (!g193) & (!g194)) + ((g62) & (g104) & (!sk[77]) & (!g66) & (!g193) & (!g194)) + ((g62) & (g104) & (!sk[77]) & (!g66) & (!g193) & (g194)) + ((g62) & (g104) & (!sk[77]) & (!g66) & (g193) & (!g194)) + ((g62) & (g104) & (!sk[77]) & (!g66) & (g193) & (g194)) + ((g62) & (g104) & (!sk[77]) & (g66) & (!g193) & (!g194)) + ((g62) & (g104) & (!sk[77]) & (g66) & (!g193) & (g194)) + ((g62) & (g104) & (!sk[77]) & (g66) & (g193) & (!g194)) + ((g62) & (g104) & (!sk[77]) & (g66) & (g193) & (g194)) + ((g62) & (g104) & (sk[77]) & (!g66) & (!g193) & (!g194)));
	assign g196 = (((g168) & (g173) & (g180) & (g183) & (g192) & (g195)));
	assign g197 = (((!g122) & (!sk[79]) & (!g159) & (g196)) + ((!g122) & (!sk[79]) & (g159) & (g196)) + ((!g122) & (sk[79]) & (!g159) & (g196)) + ((!g122) & (sk[79]) & (g159) & (!g196)) + ((!g122) & (sk[79]) & (g159) & (g196)) + ((g122) & (!sk[79]) & (!g159) & (!g196)) + ((g122) & (!sk[79]) & (!g159) & (g196)) + ((g122) & (!sk[79]) & (g159) & (!g196)) + ((g122) & (!sk[79]) & (g159) & (g196)));
	assign g198 = (((!ax22x) & (!ax7x) & (!sk[80]) & (g3) & (!ax6x)) + ((!ax22x) & (!ax7x) & (!sk[80]) & (g3) & (ax6x)) + ((!ax22x) & (!ax7x) & (sk[80]) & (!g3) & (!ax6x)) + ((!ax22x) & (!ax7x) & (sk[80]) & (!g3) & (ax6x)) + ((!ax22x) & (!ax7x) & (sk[80]) & (g3) & (ax6x)) + ((!ax22x) & (ax7x) & (!sk[80]) & (g3) & (!ax6x)) + ((!ax22x) & (ax7x) & (!sk[80]) & (g3) & (ax6x)) + ((!ax22x) & (ax7x) & (sk[80]) & (g3) & (!ax6x)) + ((ax22x) & (!ax7x) & (!sk[80]) & (!g3) & (!ax6x)) + ((ax22x) & (!ax7x) & (!sk[80]) & (!g3) & (ax6x)) + ((ax22x) & (!ax7x) & (!sk[80]) & (g3) & (!ax6x)) + ((ax22x) & (!ax7x) & (!sk[80]) & (g3) & (ax6x)) + ((ax22x) & (ax7x) & (!sk[80]) & (!g3) & (!ax6x)) + ((ax22x) & (ax7x) & (!sk[80]) & (!g3) & (ax6x)) + ((ax22x) & (ax7x) & (!sk[80]) & (g3) & (!ax6x)) + ((ax22x) & (ax7x) & (!sk[80]) & (g3) & (ax6x)) + ((ax22x) & (ax7x) & (sk[80]) & (!g3) & (!ax6x)) + ((ax22x) & (ax7x) & (sk[80]) & (!g3) & (ax6x)) + ((ax22x) & (ax7x) & (sk[80]) & (g3) & (!ax6x)) + ((ax22x) & (ax7x) & (sk[80]) & (g3) & (ax6x)));
	assign g199 = (((!ax7x) & (!sk[81]) & (!g3) & (ax6x)) + ((!ax7x) & (!sk[81]) & (g3) & (ax6x)) + ((!ax7x) & (sk[81]) & (g3) & (!ax6x)) + ((ax7x) & (!sk[81]) & (!g3) & (!ax6x)) + ((ax7x) & (!sk[81]) & (!g3) & (ax6x)) + ((ax7x) & (!sk[81]) & (g3) & (!ax6x)) + ((ax7x) & (!sk[81]) & (g3) & (ax6x)));
	assign g200 = (((!ax22x) & (!sk[82]) & (!g199) & (ax8x)) + ((!ax22x) & (!sk[82]) & (g199) & (ax8x)) + ((!ax22x) & (sk[82]) & (!g199) & (!ax8x)) + ((!ax22x) & (sk[82]) & (g199) & (ax8x)) + ((ax22x) & (!sk[82]) & (!g199) & (!ax8x)) + ((ax22x) & (!sk[82]) & (!g199) & (ax8x)) + ((ax22x) & (!sk[82]) & (g199) & (!ax8x)) + ((ax22x) & (!sk[82]) & (g199) & (ax8x)) + ((ax22x) & (sk[82]) & (!g199) & (ax8x)) + ((ax22x) & (sk[82]) & (g199) & (ax8x)));
	assign g201 = (((!g69) & (!g197) & (!g198) & (sk[83]) & (g200)) + ((!g69) & (!g197) & (g198) & (!sk[83]) & (!g200)) + ((!g69) & (!g197) & (g198) & (!sk[83]) & (g200)) + ((!g69) & (!g197) & (g198) & (sk[83]) & (!g200)) + ((!g69) & (!g197) & (g198) & (sk[83]) & (g200)) + ((!g69) & (g197) & (g198) & (!sk[83]) & (!g200)) + ((!g69) & (g197) & (g198) & (!sk[83]) & (g200)) + ((!g69) & (g197) & (g198) & (sk[83]) & (g200)) + ((g69) & (!g197) & (!g198) & (!sk[83]) & (!g200)) + ((g69) & (!g197) & (!g198) & (!sk[83]) & (g200)) + ((g69) & (!g197) & (g198) & (!sk[83]) & (!g200)) + ((g69) & (!g197) & (g198) & (!sk[83]) & (g200)) + ((g69) & (g197) & (!g198) & (!sk[83]) & (!g200)) + ((g69) & (g197) & (!g198) & (!sk[83]) & (g200)) + ((g69) & (g197) & (g198) & (!sk[83]) & (!g200)) + ((g69) & (g197) & (g198) & (!sk[83]) & (g200)));
	assign g202 = (((!sk[84]) & (!ax22x) & (!ax11x) & (g4)) + ((!sk[84]) & (!ax22x) & (ax11x) & (g4)) + ((!sk[84]) & (ax22x) & (!ax11x) & (!g4)) + ((!sk[84]) & (ax22x) & (!ax11x) & (g4)) + ((!sk[84]) & (ax22x) & (ax11x) & (!g4)) + ((!sk[84]) & (ax22x) & (ax11x) & (g4)) + ((sk[84]) & (!ax22x) & (!ax11x) & (!g4)) + ((sk[84]) & (!ax22x) & (ax11x) & (g4)) + ((sk[84]) & (ax22x) & (ax11x) & (!g4)) + ((sk[84]) & (ax22x) & (ax11x) & (g4)));
	assign g203 = (((!sk[85]) & (!g38) & (!g99) & (g25)) + ((!sk[85]) & (!g38) & (g99) & (g25)) + ((!sk[85]) & (g38) & (!g99) & (!g25)) + ((!sk[85]) & (g38) & (!g99) & (g25)) + ((!sk[85]) & (g38) & (g99) & (!g25)) + ((!sk[85]) & (g38) & (g99) & (g25)) + ((sk[85]) & (!g38) & (g99) & (g25)) + ((sk[85]) & (g38) & (g99) & (!g25)) + ((sk[85]) & (g38) & (g99) & (g25)));
	assign g204 = (((!g99) & (!g46) & (!sk[86]) & (g40) & (!g42)) + ((!g99) & (!g46) & (!sk[86]) & (g40) & (g42)) + ((!g99) & (g46) & (!sk[86]) & (g40) & (!g42)) + ((!g99) & (g46) & (!sk[86]) & (g40) & (g42)) + ((!g99) & (g46) & (sk[86]) & (g40) & (!g42)) + ((!g99) & (g46) & (sk[86]) & (g40) & (g42)) + ((g99) & (!g46) & (!sk[86]) & (!g40) & (!g42)) + ((g99) & (!g46) & (!sk[86]) & (!g40) & (g42)) + ((g99) & (!g46) & (!sk[86]) & (g40) & (!g42)) + ((g99) & (!g46) & (!sk[86]) & (g40) & (g42)) + ((g99) & (!g46) & (sk[86]) & (!g40) & (g42)) + ((g99) & (!g46) & (sk[86]) & (g40) & (g42)) + ((g99) & (g46) & (!sk[86]) & (!g40) & (!g42)) + ((g99) & (g46) & (!sk[86]) & (!g40) & (g42)) + ((g99) & (g46) & (!sk[86]) & (g40) & (!g42)) + ((g99) & (g46) & (!sk[86]) & (g40) & (g42)) + ((g99) & (g46) & (sk[86]) & (!g40) & (g42)) + ((g99) & (g46) & (sk[86]) & (g40) & (!g42)) + ((g99) & (g46) & (sk[86]) & (g40) & (g42)));
	assign g205 = (((!g112) & (!g113) & (!g97) & (g98) & (!g71) & (g46)) + ((!g112) & (!g113) & (!g97) & (g98) & (g71) & (g46)) + ((!g112) & (!g113) & (g97) & (g98) & (!g71) & (g46)) + ((!g112) & (!g113) & (g97) & (g98) & (g71) & (g46)) + ((g112) & (!g113) & (g97) & (!g98) & (g71) & (!g46)) + ((g112) & (!g113) & (g97) & (!g98) & (g71) & (g46)) + ((g112) & (g113) & (g97) & (g98) & (g71) & (!g46)) + ((g112) & (g113) & (g97) & (g98) & (g71) & (g46)));
	assign g206 = (((!g112) & (!g113) & (!g97) & (!g98) & (g62) & (!g46)) + ((!g112) & (!g113) & (!g97) & (!g98) & (g62) & (g46)) + ((!g112) & (!g113) & (!g97) & (g98) & (g62) & (!g46)) + ((!g112) & (!g113) & (!g97) & (g98) & (g62) & (g46)) + ((!g112) & (!g113) & (g97) & (!g98) & (!g62) & (g46)) + ((!g112) & (!g113) & (g97) & (!g98) & (g62) & (!g46)) + ((!g112) & (!g113) & (g97) & (!g98) & (g62) & (g46)) + ((!g112) & (!g113) & (g97) & (g98) & (g62) & (!g46)) + ((!g112) & (!g113) & (g97) & (g98) & (g62) & (g46)) + ((!g112) & (g113) & (g97) & (!g98) & (!g62) & (g46)) + ((!g112) & (g113) & (g97) & (!g98) & (g62) & (g46)));
	assign g207 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!sk[89]) & (!g58)) + ((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!sk[89]) & (g58)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (!sk[89]) & (!g58)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (!sk[89]) & (g58)) + ((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (!sk[89]) & (!g58)) + ((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (!sk[89]) & (g58)) + ((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (sk[89]) & (g58)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (!sk[89]) & (!g58)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (!sk[89]) & (g58)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!sk[89]) & (!g58)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!sk[89]) & (g58)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (!sk[89]) & (!g58)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (!sk[89]) & (g58)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (sk[89]) & (g58)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (!sk[89]) & (!g58)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (!sk[89]) & (g58)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (sk[89]) & (g58)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (!sk[89]) & (!g58)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (!sk[89]) & (g58)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (!sk[89]) & (!g58)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (!sk[89]) & (g58)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (sk[89]) & (g58)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!sk[89]) & (!g58)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!sk[89]) & (g58)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (!sk[89]) & (!g58)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (!sk[89]) & (g58)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!sk[89]) & (!g58)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!sk[89]) & (g58)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (!sk[89]) & (!g58)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (!sk[89]) & (g58)));
	assign g208 = (((!g128) & (!g97) & (!g98) & (!g99) & (!g71) & (!g207)) + ((!g128) & (!g97) & (!g98) & (!g99) & (g71) & (!g207)) + ((!g128) & (!g97) & (!g98) & (g99) & (!g71) & (!g207)) + ((!g128) & (!g97) & (!g98) & (g99) & (g71) & (!g207)) + ((!g128) & (!g97) & (g98) & (!g99) & (!g71) & (!g207)) + ((!g128) & (!g97) & (g98) & (!g99) & (g71) & (!g207)) + ((!g128) & (!g97) & (g98) & (g99) & (!g71) & (!g207)) + ((!g128) & (!g97) & (g98) & (g99) & (g71) & (!g207)) + ((!g128) & (g97) & (!g98) & (!g99) & (!g71) & (!g207)) + ((!g128) & (g97) & (!g98) & (!g99) & (g71) & (!g207)) + ((!g128) & (g97) & (!g98) & (g99) & (!g71) & (!g207)) + ((!g128) & (g97) & (!g98) & (g99) & (g71) & (!g207)) + ((!g128) & (g97) & (g98) & (!g99) & (!g71) & (!g207)) + ((!g128) & (g97) & (g98) & (!g99) & (g71) & (!g207)) + ((!g128) & (g97) & (g98) & (g99) & (!g71) & (!g207)) + ((!g128) & (g97) & (g98) & (g99) & (g71) & (!g207)) + ((g128) & (!g97) & (!g98) & (!g99) & (!g71) & (!g207)) + ((g128) & (!g97) & (!g98) & (g99) & (!g71) & (!g207)) + ((g128) & (!g97) & (g98) & (!g99) & (!g71) & (!g207)) + ((g128) & (g97) & (!g98) & (!g99) & (!g71) & (!g207)) + ((g128) & (g97) & (!g98) & (g99) & (!g71) & (!g207)) + ((g128) & (g97) & (g98) & (!g99) & (!g71) & (!g207)) + ((g128) & (g97) & (g98) & (!g99) & (g71) & (!g207)) + ((g128) & (g97) & (g98) & (g99) & (!g71) & (!g207)) + ((g128) & (g97) & (g98) & (g99) & (g71) & (!g207)));
	assign g209 = (((!g203) & (!g204) & (!g205) & (!sk[91]) & (g206) & (!g208)) + ((!g203) & (!g204) & (!g205) & (!sk[91]) & (g206) & (g208)) + ((!g203) & (!g204) & (!g205) & (sk[91]) & (!g206) & (g208)) + ((!g203) & (!g204) & (g205) & (!sk[91]) & (g206) & (!g208)) + ((!g203) & (!g204) & (g205) & (!sk[91]) & (g206) & (g208)) + ((!g203) & (g204) & (!g205) & (!sk[91]) & (!g206) & (!g208)) + ((!g203) & (g204) & (!g205) & (!sk[91]) & (!g206) & (g208)) + ((!g203) & (g204) & (!g205) & (!sk[91]) & (g206) & (!g208)) + ((!g203) & (g204) & (!g205) & (!sk[91]) & (g206) & (g208)) + ((!g203) & (g204) & (g205) & (!sk[91]) & (!g206) & (!g208)) + ((!g203) & (g204) & (g205) & (!sk[91]) & (!g206) & (g208)) + ((!g203) & (g204) & (g205) & (!sk[91]) & (g206) & (!g208)) + ((!g203) & (g204) & (g205) & (!sk[91]) & (g206) & (g208)) + ((g203) & (!g204) & (!g205) & (!sk[91]) & (g206) & (!g208)) + ((g203) & (!g204) & (!g205) & (!sk[91]) & (g206) & (g208)) + ((g203) & (!g204) & (g205) & (!sk[91]) & (!g206) & (!g208)) + ((g203) & (!g204) & (g205) & (!sk[91]) & (!g206) & (g208)) + ((g203) & (!g204) & (g205) & (!sk[91]) & (g206) & (!g208)) + ((g203) & (!g204) & (g205) & (!sk[91]) & (g206) & (g208)) + ((g203) & (g204) & (!g205) & (!sk[91]) & (!g206) & (!g208)) + ((g203) & (g204) & (!g205) & (!sk[91]) & (!g206) & (g208)) + ((g203) & (g204) & (!g205) & (!sk[91]) & (g206) & (!g208)) + ((g203) & (g204) & (!g205) & (!sk[91]) & (g206) & (g208)) + ((g203) & (g204) & (g205) & (!sk[91]) & (!g206) & (!g208)) + ((g203) & (g204) & (g205) & (!sk[91]) & (!g206) & (g208)) + ((g203) & (g204) & (g205) & (!sk[91]) & (g206) & (!g208)) + ((g203) & (g204) & (g205) & (!sk[91]) & (g206) & (g208)));
	assign g210 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g91)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g91)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g91)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g91)));
	assign g211 = (((!g128) & (!g97) & (!g98) & (!sk[93]) & (g70) & (!g104)) + ((!g128) & (!g97) & (!g98) & (!sk[93]) & (g70) & (g104)) + ((!g128) & (!g97) & (g98) & (!sk[93]) & (g70) & (!g104)) + ((!g128) & (!g97) & (g98) & (!sk[93]) & (g70) & (g104)) + ((!g128) & (g97) & (!g98) & (!sk[93]) & (!g70) & (!g104)) + ((!g128) & (g97) & (!g98) & (!sk[93]) & (!g70) & (g104)) + ((!g128) & (g97) & (!g98) & (!sk[93]) & (g70) & (!g104)) + ((!g128) & (g97) & (!g98) & (!sk[93]) & (g70) & (g104)) + ((!g128) & (g97) & (g98) & (!sk[93]) & (!g70) & (!g104)) + ((!g128) & (g97) & (g98) & (!sk[93]) & (!g70) & (g104)) + ((!g128) & (g97) & (g98) & (!sk[93]) & (g70) & (!g104)) + ((!g128) & (g97) & (g98) & (!sk[93]) & (g70) & (g104)) + ((g128) & (!g97) & (!g98) & (!sk[93]) & (g70) & (!g104)) + ((g128) & (!g97) & (!g98) & (!sk[93]) & (g70) & (g104)) + ((g128) & (!g97) & (!g98) & (sk[93]) & (g70) & (!g104)) + ((g128) & (!g97) & (!g98) & (sk[93]) & (g70) & (g104)) + ((g128) & (!g97) & (g98) & (!sk[93]) & (!g70) & (!g104)) + ((g128) & (!g97) & (g98) & (!sk[93]) & (!g70) & (g104)) + ((g128) & (!g97) & (g98) & (!sk[93]) & (g70) & (!g104)) + ((g128) & (!g97) & (g98) & (!sk[93]) & (g70) & (g104)) + ((g128) & (!g97) & (g98) & (sk[93]) & (!g70) & (g104)) + ((g128) & (!g97) & (g98) & (sk[93]) & (g70) & (!g104)) + ((g128) & (!g97) & (g98) & (sk[93]) & (g70) & (g104)) + ((g128) & (g97) & (!g98) & (!sk[93]) & (!g70) & (!g104)) + ((g128) & (g97) & (!g98) & (!sk[93]) & (!g70) & (g104)) + ((g128) & (g97) & (!g98) & (!sk[93]) & (g70) & (!g104)) + ((g128) & (g97) & (!g98) & (!sk[93]) & (g70) & (g104)) + ((g128) & (g97) & (g98) & (!sk[93]) & (!g70) & (!g104)) + ((g128) & (g97) & (g98) & (!sk[93]) & (!g70) & (g104)) + ((g128) & (g97) & (g98) & (!sk[93]) & (g70) & (!g104)) + ((g128) & (g97) & (g98) & (!sk[93]) & (g70) & (g104)) + ((g128) & (g97) & (g98) & (sk[93]) & (g70) & (!g104)) + ((g128) & (g97) & (g98) & (sk[93]) & (g70) & (g104)));
	assign g212 = (((!g38) & (!g70) & (!g99) & (!g104) & (!g40) & (!g42)) + ((!g38) & (!g70) & (!g99) & (!g104) & (!g40) & (g42)) + ((!g38) & (!g70) & (!g99) & (!g104) & (g40) & (!g42)) + ((!g38) & (!g70) & (!g99) & (!g104) & (g40) & (g42)) + ((!g38) & (!g70) & (!g99) & (g104) & (!g40) & (!g42)) + ((!g38) & (!g70) & (!g99) & (g104) & (g40) & (!g42)) + ((!g38) & (!g70) & (g99) & (!g104) & (!g40) & (!g42)) + ((!g38) & (!g70) & (g99) & (!g104) & (!g40) & (g42)) + ((!g38) & (!g70) & (g99) & (g104) & (!g40) & (!g42)) + ((!g38) & (g70) & (!g99) & (!g104) & (!g40) & (!g42)) + ((!g38) & (g70) & (!g99) & (!g104) & (!g40) & (g42)) + ((!g38) & (g70) & (!g99) & (!g104) & (g40) & (!g42)) + ((!g38) & (g70) & (!g99) & (!g104) & (g40) & (g42)) + ((!g38) & (g70) & (!g99) & (g104) & (!g40) & (!g42)) + ((!g38) & (g70) & (!g99) & (g104) & (g40) & (!g42)) + ((!g38) & (g70) & (g99) & (!g104) & (!g40) & (!g42)) + ((!g38) & (g70) & (g99) & (!g104) & (!g40) & (g42)) + ((!g38) & (g70) & (g99) & (g104) & (!g40) & (!g42)) + ((g38) & (!g70) & (!g99) & (!g104) & (!g40) & (!g42)) + ((g38) & (!g70) & (!g99) & (!g104) & (!g40) & (g42)) + ((g38) & (!g70) & (!g99) & (!g104) & (g40) & (!g42)) + ((g38) & (!g70) & (!g99) & (!g104) & (g40) & (g42)) + ((g38) & (!g70) & (g99) & (!g104) & (!g40) & (!g42)) + ((g38) & (!g70) & (g99) & (!g104) & (!g40) & (g42)));
	assign g213 = (((!sk[95]) & (!g70) & (!g58) & (!g104) & (g25) & (!g32)) + ((!sk[95]) & (!g70) & (!g58) & (!g104) & (g25) & (g32)) + ((!sk[95]) & (!g70) & (!g58) & (g104) & (g25) & (!g32)) + ((!sk[95]) & (!g70) & (!g58) & (g104) & (g25) & (g32)) + ((!sk[95]) & (!g70) & (g58) & (!g104) & (!g25) & (!g32)) + ((!sk[95]) & (!g70) & (g58) & (!g104) & (!g25) & (g32)) + ((!sk[95]) & (!g70) & (g58) & (!g104) & (g25) & (!g32)) + ((!sk[95]) & (!g70) & (g58) & (!g104) & (g25) & (g32)) + ((!sk[95]) & (!g70) & (g58) & (g104) & (!g25) & (!g32)) + ((!sk[95]) & (!g70) & (g58) & (g104) & (!g25) & (g32)) + ((!sk[95]) & (!g70) & (g58) & (g104) & (g25) & (!g32)) + ((!sk[95]) & (!g70) & (g58) & (g104) & (g25) & (g32)) + ((!sk[95]) & (g70) & (!g58) & (!g104) & (g25) & (!g32)) + ((!sk[95]) & (g70) & (!g58) & (!g104) & (g25) & (g32)) + ((!sk[95]) & (g70) & (!g58) & (g104) & (!g25) & (!g32)) + ((!sk[95]) & (g70) & (!g58) & (g104) & (!g25) & (g32)) + ((!sk[95]) & (g70) & (!g58) & (g104) & (g25) & (!g32)) + ((!sk[95]) & (g70) & (!g58) & (g104) & (g25) & (g32)) + ((!sk[95]) & (g70) & (g58) & (!g104) & (!g25) & (!g32)) + ((!sk[95]) & (g70) & (g58) & (!g104) & (!g25) & (g32)) + ((!sk[95]) & (g70) & (g58) & (!g104) & (g25) & (!g32)) + ((!sk[95]) & (g70) & (g58) & (!g104) & (g25) & (g32)) + ((!sk[95]) & (g70) & (g58) & (g104) & (!g25) & (!g32)) + ((!sk[95]) & (g70) & (g58) & (g104) & (!g25) & (g32)) + ((!sk[95]) & (g70) & (g58) & (g104) & (g25) & (!g32)) + ((!sk[95]) & (g70) & (g58) & (g104) & (g25) & (g32)) + ((sk[95]) & (!g70) & (!g58) & (!g104) & (!g25) & (!g32)) + ((sk[95]) & (!g70) & (!g58) & (!g104) & (!g25) & (g32)) + ((sk[95]) & (!g70) & (!g58) & (!g104) & (g25) & (!g32)) + ((sk[95]) & (!g70) & (!g58) & (!g104) & (g25) & (g32)) + ((sk[95]) & (!g70) & (!g58) & (g104) & (!g25) & (!g32)) + ((sk[95]) & (!g70) & (!g58) & (g104) & (!g25) & (g32)) + ((sk[95]) & (!g70) & (g58) & (!g104) & (!g25) & (!g32)) + ((sk[95]) & (!g70) & (g58) & (!g104) & (!g25) & (g32)) + ((sk[95]) & (!g70) & (g58) & (!g104) & (g25) & (!g32)) + ((sk[95]) & (!g70) & (g58) & (!g104) & (g25) & (g32)) + ((sk[95]) & (g70) & (!g58) & (!g104) & (!g25) & (!g32)) + ((sk[95]) & (g70) & (!g58) & (!g104) & (g25) & (!g32)) + ((sk[95]) & (g70) & (!g58) & (g104) & (!g25) & (!g32)));
	assign g214 = (((!sk[96]) & (!g70) & (!g12) & (!g104) & (g32) & (!g20)) + ((!sk[96]) & (!g70) & (!g12) & (!g104) & (g32) & (g20)) + ((!sk[96]) & (!g70) & (!g12) & (g104) & (g32) & (!g20)) + ((!sk[96]) & (!g70) & (!g12) & (g104) & (g32) & (g20)) + ((!sk[96]) & (!g70) & (g12) & (!g104) & (!g32) & (!g20)) + ((!sk[96]) & (!g70) & (g12) & (!g104) & (!g32) & (g20)) + ((!sk[96]) & (!g70) & (g12) & (!g104) & (g32) & (!g20)) + ((!sk[96]) & (!g70) & (g12) & (!g104) & (g32) & (g20)) + ((!sk[96]) & (!g70) & (g12) & (g104) & (!g32) & (!g20)) + ((!sk[96]) & (!g70) & (g12) & (g104) & (!g32) & (g20)) + ((!sk[96]) & (!g70) & (g12) & (g104) & (g32) & (!g20)) + ((!sk[96]) & (!g70) & (g12) & (g104) & (g32) & (g20)) + ((!sk[96]) & (g70) & (!g12) & (!g104) & (g32) & (!g20)) + ((!sk[96]) & (g70) & (!g12) & (!g104) & (g32) & (g20)) + ((!sk[96]) & (g70) & (!g12) & (g104) & (!g32) & (!g20)) + ((!sk[96]) & (g70) & (!g12) & (g104) & (!g32) & (g20)) + ((!sk[96]) & (g70) & (!g12) & (g104) & (g32) & (!g20)) + ((!sk[96]) & (g70) & (!g12) & (g104) & (g32) & (g20)) + ((!sk[96]) & (g70) & (g12) & (!g104) & (!g32) & (!g20)) + ((!sk[96]) & (g70) & (g12) & (!g104) & (!g32) & (g20)) + ((!sk[96]) & (g70) & (g12) & (!g104) & (g32) & (!g20)) + ((!sk[96]) & (g70) & (g12) & (!g104) & (g32) & (g20)) + ((!sk[96]) & (g70) & (g12) & (g104) & (!g32) & (!g20)) + ((!sk[96]) & (g70) & (g12) & (g104) & (!g32) & (g20)) + ((!sk[96]) & (g70) & (g12) & (g104) & (g32) & (!g20)) + ((!sk[96]) & (g70) & (g12) & (g104) & (g32) & (g20)) + ((sk[96]) & (!g70) & (!g12) & (!g104) & (!g32) & (!g20)) + ((sk[96]) & (!g70) & (!g12) & (!g104) & (!g32) & (g20)) + ((sk[96]) & (!g70) & (!g12) & (!g104) & (g32) & (!g20)) + ((sk[96]) & (!g70) & (!g12) & (!g104) & (g32) & (g20)) + ((sk[96]) & (!g70) & (!g12) & (g104) & (!g32) & (!g20)) + ((sk[96]) & (!g70) & (!g12) & (g104) & (!g32) & (g20)) + ((sk[96]) & (!g70) & (g12) & (!g104) & (!g32) & (!g20)) + ((sk[96]) & (!g70) & (g12) & (!g104) & (!g32) & (g20)) + ((sk[96]) & (!g70) & (g12) & (!g104) & (g32) & (!g20)) + ((sk[96]) & (!g70) & (g12) & (!g104) & (g32) & (g20)) + ((sk[96]) & (g70) & (!g12) & (!g104) & (!g32) & (!g20)) + ((sk[96]) & (g70) & (!g12) & (!g104) & (g32) & (!g20)) + ((sk[96]) & (g70) & (!g12) & (g104) & (!g32) & (!g20)));
	assign g215 = (((g92) & (!g210) & (!g211) & (g212) & (g213) & (g214)));
	assign g216 = (((!g112) & (!g113) & (!g97) & (g98) & (!g99) & (g71)) + ((!g112) & (!g113) & (!g97) & (g98) & (g99) & (!g71)) + ((!g112) & (!g113) & (!g97) & (g98) & (g99) & (g71)) + ((!g112) & (!g113) & (g97) & (!g98) & (!g99) & (g71)) + ((!g112) & (!g113) & (g97) & (!g98) & (g99) & (!g71)) + ((!g112) & (!g113) & (g97) & (!g98) & (g99) & (g71)) + ((!g112) & (!g113) & (g97) & (g98) & (!g99) & (g71)) + ((!g112) & (!g113) & (g97) & (g98) & (g99) & (!g71)) + ((!g112) & (!g113) & (g97) & (g98) & (g99) & (g71)) + ((!g112) & (g113) & (!g97) & (!g98) & (!g99) & (g71)) + ((!g112) & (g113) & (!g97) & (!g98) & (g99) & (!g71)) + ((!g112) & (g113) & (!g97) & (!g98) & (g99) & (g71)) + ((!g112) & (g113) & (!g97) & (g98) & (g99) & (!g71)) + ((!g112) & (g113) & (!g97) & (g98) & (g99) & (g71)));
	assign g217 = (((!g112) & (g113) & (!g97) & (g98) & (!g99) & (g71)) + ((!g112) & (g113) & (!g97) & (g98) & (g99) & (g71)) + ((!g112) & (g113) & (g97) & (!g98) & (!g99) & (g71)) + ((!g112) & (g113) & (g97) & (!g98) & (g99) & (!g71)) + ((!g112) & (g113) & (g97) & (!g98) & (g99) & (g71)) + ((!g112) & (g113) & (g97) & (g98) & (!g99) & (g71)) + ((!g112) & (g113) & (g97) & (g98) & (g99) & (!g71)) + ((!g112) & (g113) & (g97) & (g98) & (g99) & (g71)) + ((g112) & (!g113) & (!g97) & (!g98) & (!g99) & (g71)) + ((g112) & (!g113) & (!g97) & (!g98) & (g99) & (!g71)) + ((g112) & (!g113) & (!g97) & (!g98) & (g99) & (g71)) + ((g112) & (!g113) & (!g97) & (g98) & (!g99) & (g71)) + ((g112) & (!g113) & (!g97) & (g98) & (g99) & (!g71)) + ((g112) & (!g113) & (!g97) & (g98) & (g99) & (g71)) + ((g112) & (!g113) & (g97) & (!g98) & (g99) & (!g71)) + ((g112) & (!g113) & (g97) & (!g98) & (g99) & (g71)));
	assign g218 = (((g45) & (g68) & (!g209) & (!g215) & (!g216) & (!g217)) + ((g45) & (g68) & (!g209) & (!g215) & (!g216) & (g217)) + ((g45) & (g68) & (!g209) & (!g215) & (g216) & (!g217)) + ((g45) & (g68) & (!g209) & (!g215) & (g216) & (g217)) + ((g45) & (g68) & (!g209) & (g215) & (!g216) & (!g217)) + ((g45) & (g68) & (!g209) & (g215) & (!g216) & (g217)) + ((g45) & (g68) & (!g209) & (g215) & (g216) & (!g217)) + ((g45) & (g68) & (!g209) & (g215) & (g216) & (g217)) + ((g45) & (g68) & (g209) & (!g215) & (!g216) & (!g217)) + ((g45) & (g68) & (g209) & (!g215) & (!g216) & (g217)) + ((g45) & (g68) & (g209) & (!g215) & (g216) & (!g217)) + ((g45) & (g68) & (g209) & (!g215) & (g216) & (g217)) + ((g45) & (g68) & (g209) & (g215) & (!g216) & (g217)) + ((g45) & (g68) & (g209) & (g215) & (g216) & (!g217)) + ((g45) & (g68) & (g209) & (g215) & (g216) & (g217)));
	assign g219 = (((!g62) & (!g46) & (!sk[101]) & (g91) & (!g217)) + ((!g62) & (!g46) & (!sk[101]) & (g91) & (g217)) + ((!g62) & (!g46) & (sk[101]) & (!g91) & (!g217)) + ((!g62) & (!g46) & (sk[101]) & (g91) & (!g217)) + ((!g62) & (g46) & (!sk[101]) & (g91) & (!g217)) + ((!g62) & (g46) & (!sk[101]) & (g91) & (g217)) + ((!g62) & (g46) & (sk[101]) & (!g91) & (!g217)) + ((g62) & (!g46) & (!sk[101]) & (!g91) & (!g217)) + ((g62) & (!g46) & (!sk[101]) & (!g91) & (g217)) + ((g62) & (!g46) & (!sk[101]) & (g91) & (!g217)) + ((g62) & (!g46) & (!sk[101]) & (g91) & (g217)) + ((g62) & (!g46) & (sk[101]) & (!g91) & (!g217)) + ((g62) & (g46) & (!sk[101]) & (!g91) & (!g217)) + ((g62) & (g46) & (!sk[101]) & (!g91) & (g217)) + ((g62) & (g46) & (!sk[101]) & (g91) & (!g217)) + ((g62) & (g46) & (!sk[101]) & (g91) & (g217)) + ((g62) & (g46) & (sk[101]) & (!g91) & (!g217)));
	assign g220 = (((!g209) & (!g215) & (g216) & (!sk[102]) & (!g219)) + ((!g209) & (!g215) & (g216) & (!sk[102]) & (g219)) + ((!g209) & (g215) & (g216) & (!sk[102]) & (!g219)) + ((!g209) & (g215) & (g216) & (!sk[102]) & (g219)) + ((g209) & (!g215) & (!g216) & (!sk[102]) & (!g219)) + ((g209) & (!g215) & (!g216) & (!sk[102]) & (g219)) + ((g209) & (!g215) & (!g216) & (sk[102]) & (g219)) + ((g209) & (!g215) & (g216) & (!sk[102]) & (!g219)) + ((g209) & (!g215) & (g216) & (!sk[102]) & (g219)) + ((g209) & (g215) & (!g216) & (!sk[102]) & (!g219)) + ((g209) & (g215) & (!g216) & (!sk[102]) & (g219)) + ((g209) & (g215) & (!g216) & (sk[102]) & (!g219)) + ((g209) & (g215) & (g216) & (!sk[102]) & (!g219)) + ((g209) & (g215) & (g216) & (!sk[102]) & (g219)) + ((g209) & (g215) & (g216) & (sk[102]) & (!g219)) + ((g209) & (g215) & (g216) & (sk[102]) & (g219)));
	assign g221 = (((!g45) & (!g68) & (g209) & (!g215) & (!g216) & (g219)) + ((!g45) & (!g68) & (g209) & (g215) & (!g216) & (!g219)) + ((!g45) & (!g68) & (g209) & (g215) & (!g216) & (g219)) + ((!g45) & (!g68) & (g209) & (g215) & (g216) & (!g219)) + ((!g45) & (!g68) & (g209) & (g215) & (g216) & (g219)) + ((!g45) & (g68) & (g209) & (!g215) & (!g216) & (g219)) + ((!g45) & (g68) & (g209) & (g215) & (!g216) & (!g219)) + ((!g45) & (g68) & (g209) & (g215) & (!g216) & (g219)) + ((!g45) & (g68) & (g209) & (g215) & (g216) & (!g219)) + ((!g45) & (g68) & (g209) & (g215) & (g216) & (g219)) + ((g45) & (!g68) & (g209) & (!g215) & (!g216) & (g219)) + ((g45) & (!g68) & (g209) & (g215) & (!g216) & (!g219)) + ((g45) & (!g68) & (g209) & (g215) & (!g216) & (g219)) + ((g45) & (!g68) & (g209) & (g215) & (g216) & (!g219)) + ((g45) & (!g68) & (g209) & (g215) & (g216) & (g219)));
	assign g222 = (((!ax22x) & (!ax9x) & (!sk[104]) & (!g199) & (ax8x) & (!ax10x)) + ((!ax22x) & (!ax9x) & (!sk[104]) & (!g199) & (ax8x) & (ax10x)) + ((!ax22x) & (!ax9x) & (!sk[104]) & (g199) & (ax8x) & (!ax10x)) + ((!ax22x) & (!ax9x) & (!sk[104]) & (g199) & (ax8x) & (ax10x)) + ((!ax22x) & (!ax9x) & (sk[104]) & (!g199) & (!ax8x) & (!ax10x)) + ((!ax22x) & (!ax9x) & (sk[104]) & (!g199) & (ax8x) & (!ax10x)) + ((!ax22x) & (!ax9x) & (sk[104]) & (g199) & (!ax8x) & (ax10x)) + ((!ax22x) & (!ax9x) & (sk[104]) & (g199) & (ax8x) & (!ax10x)) + ((!ax22x) & (ax9x) & (!sk[104]) & (!g199) & (!ax8x) & (!ax10x)) + ((!ax22x) & (ax9x) & (!sk[104]) & (!g199) & (!ax8x) & (ax10x)) + ((!ax22x) & (ax9x) & (!sk[104]) & (!g199) & (ax8x) & (!ax10x)) + ((!ax22x) & (ax9x) & (!sk[104]) & (!g199) & (ax8x) & (ax10x)) + ((!ax22x) & (ax9x) & (!sk[104]) & (g199) & (!ax8x) & (!ax10x)) + ((!ax22x) & (ax9x) & (!sk[104]) & (g199) & (!ax8x) & (ax10x)) + ((!ax22x) & (ax9x) & (!sk[104]) & (g199) & (ax8x) & (!ax10x)) + ((!ax22x) & (ax9x) & (!sk[104]) & (g199) & (ax8x) & (ax10x)) + ((!ax22x) & (ax9x) & (sk[104]) & (!g199) & (!ax8x) & (!ax10x)) + ((!ax22x) & (ax9x) & (sk[104]) & (!g199) & (ax8x) & (!ax10x)) + ((!ax22x) & (ax9x) & (sk[104]) & (g199) & (!ax8x) & (!ax10x)) + ((!ax22x) & (ax9x) & (sk[104]) & (g199) & (ax8x) & (!ax10x)) + ((ax22x) & (!ax9x) & (!sk[104]) & (!g199) & (ax8x) & (!ax10x)) + ((ax22x) & (!ax9x) & (!sk[104]) & (!g199) & (ax8x) & (ax10x)) + ((ax22x) & (!ax9x) & (!sk[104]) & (g199) & (!ax8x) & (!ax10x)) + ((ax22x) & (!ax9x) & (!sk[104]) & (g199) & (!ax8x) & (ax10x)) + ((ax22x) & (!ax9x) & (!sk[104]) & (g199) & (ax8x) & (!ax10x)) + ((ax22x) & (!ax9x) & (!sk[104]) & (g199) & (ax8x) & (ax10x)) + ((ax22x) & (!ax9x) & (sk[104]) & (!g199) & (!ax8x) & (ax10x)) + ((ax22x) & (!ax9x) & (sk[104]) & (!g199) & (ax8x) & (ax10x)) + ((ax22x) & (!ax9x) & (sk[104]) & (g199) & (!ax8x) & (ax10x)) + ((ax22x) & (!ax9x) & (sk[104]) & (g199) & (ax8x) & (ax10x)) + ((ax22x) & (ax9x) & (!sk[104]) & (!g199) & (!ax8x) & (!ax10x)) + ((ax22x) & (ax9x) & (!sk[104]) & (!g199) & (!ax8x) & (ax10x)) + ((ax22x) & (ax9x) & (!sk[104]) & (!g199) & (ax8x) & (!ax10x)) + ((ax22x) & (ax9x) & (!sk[104]) & (!g199) & (ax8x) & (ax10x)) + ((ax22x) & (ax9x) & (!sk[104]) & (g199) & (!ax8x) & (!ax10x)) + ((ax22x) & (ax9x) & (!sk[104]) & (g199) & (!ax8x) & (ax10x)) + ((ax22x) & (ax9x) & (!sk[104]) & (g199) & (ax8x) & (!ax10x)) + ((ax22x) & (ax9x) & (!sk[104]) & (g199) & (ax8x) & (ax10x)) + ((ax22x) & (ax9x) & (sk[104]) & (!g199) & (!ax8x) & (ax10x)) + ((ax22x) & (ax9x) & (sk[104]) & (!g199) & (ax8x) & (ax10x)) + ((ax22x) & (ax9x) & (sk[104]) & (g199) & (!ax8x) & (ax10x)) + ((ax22x) & (ax9x) & (sk[104]) & (g199) & (ax8x) & (ax10x)));
	assign g223 = (((!g202) & (!g218) & (!g220) & (!sk[105]) & (g221) & (!g222)) + ((!g202) & (!g218) & (!g220) & (!sk[105]) & (g221) & (g222)) + ((!g202) & (!g218) & (!g220) & (sk[105]) & (g221) & (!g222)) + ((!g202) & (!g218) & (g220) & (!sk[105]) & (g221) & (!g222)) + ((!g202) & (!g218) & (g220) & (!sk[105]) & (g221) & (g222)) + ((!g202) & (!g218) & (g220) & (sk[105]) & (g221) & (!g222)) + ((!g202) & (!g218) & (g220) & (sk[105]) & (g221) & (g222)) + ((!g202) & (g218) & (!g220) & (!sk[105]) & (!g221) & (!g222)) + ((!g202) & (g218) & (!g220) & (!sk[105]) & (!g221) & (g222)) + ((!g202) & (g218) & (!g220) & (!sk[105]) & (g221) & (!g222)) + ((!g202) & (g218) & (!g220) & (!sk[105]) & (g221) & (g222)) + ((!g202) & (g218) & (!g220) & (sk[105]) & (!g221) & (g222)) + ((!g202) & (g218) & (!g220) & (sk[105]) & (g221) & (!g222)) + ((!g202) & (g218) & (!g220) & (sk[105]) & (g221) & (g222)) + ((!g202) & (g218) & (g220) & (!sk[105]) & (!g221) & (!g222)) + ((!g202) & (g218) & (g220) & (!sk[105]) & (!g221) & (g222)) + ((!g202) & (g218) & (g220) & (!sk[105]) & (g221) & (!g222)) + ((!g202) & (g218) & (g220) & (!sk[105]) & (g221) & (g222)) + ((!g202) & (g218) & (g220) & (sk[105]) & (g221) & (!g222)) + ((!g202) & (g218) & (g220) & (sk[105]) & (g221) & (g222)) + ((g202) & (!g218) & (!g220) & (!sk[105]) & (g221) & (!g222)) + ((g202) & (!g218) & (!g220) & (!sk[105]) & (g221) & (g222)) + ((g202) & (!g218) & (!g220) & (sk[105]) & (g221) & (!g222)) + ((g202) & (!g218) & (g220) & (!sk[105]) & (!g221) & (!g222)) + ((g202) & (!g218) & (g220) & (!sk[105]) & (!g221) & (g222)) + ((g202) & (!g218) & (g220) & (!sk[105]) & (g221) & (!g222)) + ((g202) & (!g218) & (g220) & (!sk[105]) & (g221) & (g222)) + ((g202) & (g218) & (!g220) & (!sk[105]) & (!g221) & (!g222)) + ((g202) & (g218) & (!g220) & (!sk[105]) & (!g221) & (g222)) + ((g202) & (g218) & (!g220) & (!sk[105]) & (g221) & (!g222)) + ((g202) & (g218) & (!g220) & (!sk[105]) & (g221) & (g222)) + ((g202) & (g218) & (!g220) & (sk[105]) & (!g221) & (g222)) + ((g202) & (g218) & (!g220) & (sk[105]) & (g221) & (!g222)) + ((g202) & (g218) & (!g220) & (sk[105]) & (g221) & (g222)) + ((g202) & (g218) & (g220) & (!sk[105]) & (!g221) & (!g222)) + ((g202) & (g218) & (g220) & (!sk[105]) & (!g221) & (g222)) + ((g202) & (g218) & (g220) & (!sk[105]) & (g221) & (!g222)) + ((g202) & (g218) & (g220) & (!sk[105]) & (g221) & (g222)) + ((g202) & (g218) & (g220) & (sk[105]) & (!g221) & (!g222)) + ((g202) & (g218) & (g220) & (sk[105]) & (!g221) & (g222)) + ((g202) & (g218) & (g220) & (sk[105]) & (g221) & (!g222)) + ((g202) & (g218) & (g220) & (sk[105]) & (g221) & (g222)));
	assign g224 = (((!g99) & (!sk[106]) & (!g18) & (g60)) + ((!g99) & (!sk[106]) & (g18) & (g60)) + ((!g99) & (sk[106]) & (!g18) & (!g60)) + ((!g99) & (sk[106]) & (g18) & (!g60)) + ((g99) & (!sk[106]) & (!g18) & (!g60)) + ((g99) & (!sk[106]) & (!g18) & (g60)) + ((g99) & (!sk[106]) & (g18) & (!g60)) + ((g99) & (!sk[106]) & (g18) & (g60)) + ((g99) & (sk[106]) & (!g18) & (!g60)));
	assign g225 = (((!g9) & (!g16) & (!sk[107]) & (!g12) & (g30) & (!g23)) + ((!g9) & (!g16) & (!sk[107]) & (!g12) & (g30) & (g23)) + ((!g9) & (!g16) & (!sk[107]) & (g12) & (g30) & (!g23)) + ((!g9) & (!g16) & (!sk[107]) & (g12) & (g30) & (g23)) + ((!g9) & (!g16) & (sk[107]) & (!g12) & (!g30) & (!g23)) + ((!g9) & (!g16) & (sk[107]) & (!g12) & (!g30) & (g23)) + ((!g9) & (!g16) & (sk[107]) & (!g12) & (g30) & (!g23)) + ((!g9) & (!g16) & (sk[107]) & (!g12) & (g30) & (g23)) + ((!g9) & (!g16) & (sk[107]) & (g12) & (!g30) & (!g23)) + ((!g9) & (!g16) & (sk[107]) & (g12) & (!g30) & (g23)) + ((!g9) & (!g16) & (sk[107]) & (g12) & (g30) & (!g23)) + ((!g9) & (!g16) & (sk[107]) & (g12) & (g30) & (g23)) + ((!g9) & (g16) & (!sk[107]) & (!g12) & (!g30) & (!g23)) + ((!g9) & (g16) & (!sk[107]) & (!g12) & (!g30) & (g23)) + ((!g9) & (g16) & (!sk[107]) & (!g12) & (g30) & (!g23)) + ((!g9) & (g16) & (!sk[107]) & (!g12) & (g30) & (g23)) + ((!g9) & (g16) & (!sk[107]) & (g12) & (!g30) & (!g23)) + ((!g9) & (g16) & (!sk[107]) & (g12) & (!g30) & (g23)) + ((!g9) & (g16) & (!sk[107]) & (g12) & (g30) & (!g23)) + ((!g9) & (g16) & (!sk[107]) & (g12) & (g30) & (g23)) + ((!g9) & (g16) & (sk[107]) & (!g12) & (!g30) & (!g23)) + ((!g9) & (g16) & (sk[107]) & (!g12) & (!g30) & (g23)) + ((!g9) & (g16) & (sk[107]) & (!g12) & (g30) & (!g23)) + ((!g9) & (g16) & (sk[107]) & (!g12) & (g30) & (g23)) + ((g9) & (!g16) & (!sk[107]) & (!g12) & (g30) & (!g23)) + ((g9) & (!g16) & (!sk[107]) & (!g12) & (g30) & (g23)) + ((g9) & (!g16) & (!sk[107]) & (g12) & (!g30) & (!g23)) + ((g9) & (!g16) & (!sk[107]) & (g12) & (!g30) & (g23)) + ((g9) & (!g16) & (!sk[107]) & (g12) & (g30) & (!g23)) + ((g9) & (!g16) & (!sk[107]) & (g12) & (g30) & (g23)) + ((g9) & (!g16) & (sk[107]) & (!g12) & (!g30) & (!g23)) + ((g9) & (!g16) & (sk[107]) & (g12) & (!g30) & (!g23)) + ((g9) & (g16) & (!sk[107]) & (!g12) & (!g30) & (!g23)) + ((g9) & (g16) & (!sk[107]) & (!g12) & (!g30) & (g23)) + ((g9) & (g16) & (!sk[107]) & (!g12) & (g30) & (!g23)) + ((g9) & (g16) & (!sk[107]) & (!g12) & (g30) & (g23)) + ((g9) & (g16) & (!sk[107]) & (g12) & (!g30) & (!g23)) + ((g9) & (g16) & (!sk[107]) & (g12) & (!g30) & (g23)) + ((g9) & (g16) & (!sk[107]) & (g12) & (g30) & (!g23)) + ((g9) & (g16) & (!sk[107]) & (g12) & (g30) & (g23)) + ((g9) & (g16) & (sk[107]) & (!g12) & (!g30) & (!g23)));
	assign g226 = (((!g38) & (!g70) & (!g10) & (!g49) & (!g99) & (!g62)) + ((!g38) & (!g70) & (!g10) & (!g49) & (!g99) & (g62)) + ((!g38) & (!g70) & (!g10) & (!g49) & (g99) & (!g62)) + ((!g38) & (!g70) & (!g10) & (!g49) & (g99) & (g62)) + ((!g38) & (!g70) & (!g10) & (g49) & (!g99) & (!g62)) + ((!g38) & (!g70) & (!g10) & (g49) & (!g99) & (g62)) + ((!g38) & (!g70) & (g10) & (!g49) & (!g99) & (!g62)) + ((!g38) & (!g70) & (g10) & (!g49) & (!g99) & (g62)) + ((!g38) & (!g70) & (g10) & (!g49) & (g99) & (!g62)) + ((!g38) & (!g70) & (g10) & (!g49) & (g99) & (g62)) + ((!g38) & (!g70) & (g10) & (g49) & (!g99) & (!g62)) + ((!g38) & (!g70) & (g10) & (g49) & (!g99) & (g62)) + ((!g38) & (g70) & (!g10) & (!g49) & (!g99) & (!g62)) + ((!g38) & (g70) & (!g10) & (!g49) & (!g99) & (g62)) + ((!g38) & (g70) & (!g10) & (!g49) & (g99) & (!g62)) + ((!g38) & (g70) & (!g10) & (!g49) & (g99) & (g62)) + ((!g38) & (g70) & (!g10) & (g49) & (!g99) & (!g62)) + ((!g38) & (g70) & (!g10) & (g49) & (!g99) & (g62)) + ((g38) & (!g70) & (!g10) & (!g49) & (!g99) & (!g62)) + ((g38) & (!g70) & (!g10) & (g49) & (!g99) & (!g62)) + ((g38) & (!g70) & (g10) & (!g49) & (!g99) & (!g62)) + ((g38) & (!g70) & (g10) & (g49) & (!g99) & (!g62)) + ((g38) & (g70) & (!g10) & (!g49) & (!g99) & (!g62)) + ((g38) & (g70) & (!g10) & (g49) & (!g99) & (!g62)));
	assign g227 = (((!sk[109]) & (!g38) & (!g114) & (!g115) & (g8) & (!g17)) + ((!sk[109]) & (!g38) & (!g114) & (!g115) & (g8) & (g17)) + ((!sk[109]) & (!g38) & (!g114) & (g115) & (g8) & (!g17)) + ((!sk[109]) & (!g38) & (!g114) & (g115) & (g8) & (g17)) + ((!sk[109]) & (!g38) & (g114) & (!g115) & (!g8) & (!g17)) + ((!sk[109]) & (!g38) & (g114) & (!g115) & (!g8) & (g17)) + ((!sk[109]) & (!g38) & (g114) & (!g115) & (g8) & (!g17)) + ((!sk[109]) & (!g38) & (g114) & (!g115) & (g8) & (g17)) + ((!sk[109]) & (!g38) & (g114) & (g115) & (!g8) & (!g17)) + ((!sk[109]) & (!g38) & (g114) & (g115) & (!g8) & (g17)) + ((!sk[109]) & (!g38) & (g114) & (g115) & (g8) & (!g17)) + ((!sk[109]) & (!g38) & (g114) & (g115) & (g8) & (g17)) + ((!sk[109]) & (g38) & (!g114) & (!g115) & (g8) & (!g17)) + ((!sk[109]) & (g38) & (!g114) & (!g115) & (g8) & (g17)) + ((!sk[109]) & (g38) & (!g114) & (g115) & (!g8) & (!g17)) + ((!sk[109]) & (g38) & (!g114) & (g115) & (!g8) & (g17)) + ((!sk[109]) & (g38) & (!g114) & (g115) & (g8) & (!g17)) + ((!sk[109]) & (g38) & (!g114) & (g115) & (g8) & (g17)) + ((!sk[109]) & (g38) & (g114) & (!g115) & (!g8) & (!g17)) + ((!sk[109]) & (g38) & (g114) & (!g115) & (!g8) & (g17)) + ((!sk[109]) & (g38) & (g114) & (!g115) & (g8) & (!g17)) + ((!sk[109]) & (g38) & (g114) & (!g115) & (g8) & (g17)) + ((!sk[109]) & (g38) & (g114) & (g115) & (!g8) & (!g17)) + ((!sk[109]) & (g38) & (g114) & (g115) & (!g8) & (g17)) + ((!sk[109]) & (g38) & (g114) & (g115) & (g8) & (!g17)) + ((!sk[109]) & (g38) & (g114) & (g115) & (g8) & (g17)) + ((sk[109]) & (!g38) & (!g114) & (!g115) & (g8) & (g17)) + ((sk[109]) & (!g38) & (g114) & (g115) & (!g8) & (g17)) + ((sk[109]) & (g38) & (!g114) & (!g115) & (g8) & (g17)) + ((sk[109]) & (g38) & (!g114) & (g115) & (g8) & (!g17)) + ((sk[109]) & (g38) & (!g114) & (g115) & (g8) & (g17)) + ((sk[109]) & (g38) & (g114) & (g115) & (!g8) & (g17)) + ((sk[109]) & (g38) & (g114) & (g115) & (g8) & (!g17)) + ((sk[109]) & (g38) & (g114) & (g115) & (g8) & (g17)));
	assign g228 = (((!g163) & (!g54) & (!sk[110]) & (!g225) & (g226) & (!g227)) + ((!g163) & (!g54) & (!sk[110]) & (!g225) & (g226) & (g227)) + ((!g163) & (!g54) & (!sk[110]) & (g225) & (g226) & (!g227)) + ((!g163) & (!g54) & (!sk[110]) & (g225) & (g226) & (g227)) + ((!g163) & (!g54) & (sk[110]) & (g225) & (g226) & (!g227)) + ((!g163) & (g54) & (!sk[110]) & (!g225) & (!g226) & (!g227)) + ((!g163) & (g54) & (!sk[110]) & (!g225) & (!g226) & (g227)) + ((!g163) & (g54) & (!sk[110]) & (!g225) & (g226) & (!g227)) + ((!g163) & (g54) & (!sk[110]) & (!g225) & (g226) & (g227)) + ((!g163) & (g54) & (!sk[110]) & (g225) & (!g226) & (!g227)) + ((!g163) & (g54) & (!sk[110]) & (g225) & (!g226) & (g227)) + ((!g163) & (g54) & (!sk[110]) & (g225) & (g226) & (!g227)) + ((!g163) & (g54) & (!sk[110]) & (g225) & (g226) & (g227)) + ((g163) & (!g54) & (!sk[110]) & (!g225) & (g226) & (!g227)) + ((g163) & (!g54) & (!sk[110]) & (!g225) & (g226) & (g227)) + ((g163) & (!g54) & (!sk[110]) & (g225) & (!g226) & (!g227)) + ((g163) & (!g54) & (!sk[110]) & (g225) & (!g226) & (g227)) + ((g163) & (!g54) & (!sk[110]) & (g225) & (g226) & (!g227)) + ((g163) & (!g54) & (!sk[110]) & (g225) & (g226) & (g227)) + ((g163) & (g54) & (!sk[110]) & (!g225) & (!g226) & (!g227)) + ((g163) & (g54) & (!sk[110]) & (!g225) & (!g226) & (g227)) + ((g163) & (g54) & (!sk[110]) & (!g225) & (g226) & (!g227)) + ((g163) & (g54) & (!sk[110]) & (!g225) & (g226) & (g227)) + ((g163) & (g54) & (!sk[110]) & (g225) & (!g226) & (!g227)) + ((g163) & (g54) & (!sk[110]) & (g225) & (!g226) & (g227)) + ((g163) & (g54) & (!sk[110]) & (g225) & (g226) & (!g227)) + ((g163) & (g54) & (!sk[110]) & (g225) & (g226) & (g227)));
	assign g229 = (((!sk[111]) & (!g99) & (!g184) & (g40)) + ((!sk[111]) & (!g99) & (g184) & (g40)) + ((!sk[111]) & (g99) & (!g184) & (!g40)) + ((!sk[111]) & (g99) & (!g184) & (g40)) + ((!sk[111]) & (g99) & (g184) & (!g40)) + ((!sk[111]) & (g99) & (g184) & (g40)) + ((sk[111]) & (!g99) & (!g184) & (!g40)) + ((sk[111]) & (!g99) & (!g184) & (g40)) + ((sk[111]) & (g99) & (!g184) & (!g40)));
	assign g230 = (((!g58) & (!g104) & (!sk[112]) & (g90)) + ((!g58) & (!g104) & (sk[112]) & (!g90)) + ((!g58) & (g104) & (!sk[112]) & (g90)) + ((!g58) & (g104) & (sk[112]) & (!g90)) + ((g58) & (!g104) & (!sk[112]) & (!g90)) + ((g58) & (!g104) & (!sk[112]) & (g90)) + ((g58) & (!g104) & (sk[112]) & (!g90)) + ((g58) & (g104) & (!sk[112]) & (!g90)) + ((g58) & (g104) & (!sk[112]) & (g90)));
	assign g231 = (((!g38) & (!sk[113]) & (!g9) & (g80)) + ((!g38) & (!sk[113]) & (g9) & (g80)) + ((!g38) & (sk[113]) & (!g9) & (!g80)) + ((!g38) & (sk[113]) & (g9) & (!g80)) + ((g38) & (!sk[113]) & (!g9) & (!g80)) + ((g38) & (!sk[113]) & (!g9) & (g80)) + ((g38) & (!sk[113]) & (g9) & (!g80)) + ((g38) & (!sk[113]) & (g9) & (g80)) + ((g38) & (sk[113]) & (!g9) & (!g80)));
	assign g232 = (((!sk[114]) & (!g70) & (!g30) & (g57) & (!g58)) + ((!sk[114]) & (!g70) & (!g30) & (g57) & (g58)) + ((!sk[114]) & (!g70) & (g30) & (g57) & (!g58)) + ((!sk[114]) & (!g70) & (g30) & (g57) & (g58)) + ((!sk[114]) & (g70) & (!g30) & (!g57) & (!g58)) + ((!sk[114]) & (g70) & (!g30) & (!g57) & (g58)) + ((!sk[114]) & (g70) & (!g30) & (g57) & (!g58)) + ((!sk[114]) & (g70) & (!g30) & (g57) & (g58)) + ((!sk[114]) & (g70) & (g30) & (!g57) & (!g58)) + ((!sk[114]) & (g70) & (g30) & (!g57) & (g58)) + ((!sk[114]) & (g70) & (g30) & (g57) & (!g58)) + ((!sk[114]) & (g70) & (g30) & (g57) & (g58)) + ((sk[114]) & (!g70) & (g30) & (g57) & (!g58)) + ((sk[114]) & (!g70) & (g30) & (g57) & (g58)) + ((sk[114]) & (g70) & (!g30) & (!g57) & (g58)) + ((sk[114]) & (g70) & (!g30) & (g57) & (g58)) + ((sk[114]) & (g70) & (g30) & (!g57) & (g58)) + ((sk[114]) & (g70) & (g30) & (g57) & (!g58)) + ((sk[114]) & (g70) & (g30) & (g57) & (g58)));
	assign g233 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g66)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g66)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g66)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g66)));
	assign g234 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (!ax18x)) + ((!ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (!ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (ax18x)));
	assign g235 = (((!g70) & (!g16) & (!g42) & (!g233) & (!g234) & (!g166)) + ((!g70) & (!g16) & (!g42) & (!g233) & (g234) & (!g166)) + ((!g70) & (!g16) & (g42) & (!g233) & (!g234) & (!g166)) + ((!g70) & (!g16) & (g42) & (!g233) & (g234) & (!g166)) + ((!g70) & (g16) & (!g42) & (!g233) & (!g234) & (!g166)) + ((!g70) & (g16) & (g42) & (!g233) & (!g234) & (!g166)) + ((g70) & (!g16) & (!g42) & (!g233) & (!g234) & (!g166)) + ((g70) & (!g16) & (!g42) & (!g233) & (g234) & (!g166)) + ((g70) & (g16) & (!g42) & (!g233) & (!g234) & (!g166)));
	assign g236 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g10)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g10)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g10)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g10)));
	assign g237 = (((!g59) & (!g50) & (!g154) & (!g93) & (sk[119]) & (!g236)) + ((!g59) & (!g50) & (!g154) & (g93) & (!sk[119]) & (!g236)) + ((!g59) & (!g50) & (!g154) & (g93) & (!sk[119]) & (g236)) + ((!g59) & (!g50) & (g154) & (g93) & (!sk[119]) & (!g236)) + ((!g59) & (!g50) & (g154) & (g93) & (!sk[119]) & (g236)) + ((!g59) & (g50) & (!g154) & (!g93) & (!sk[119]) & (!g236)) + ((!g59) & (g50) & (!g154) & (!g93) & (!sk[119]) & (g236)) + ((!g59) & (g50) & (!g154) & (g93) & (!sk[119]) & (!g236)) + ((!g59) & (g50) & (!g154) & (g93) & (!sk[119]) & (g236)) + ((!g59) & (g50) & (g154) & (!g93) & (!sk[119]) & (!g236)) + ((!g59) & (g50) & (g154) & (!g93) & (!sk[119]) & (g236)) + ((!g59) & (g50) & (g154) & (g93) & (!sk[119]) & (!g236)) + ((!g59) & (g50) & (g154) & (g93) & (!sk[119]) & (g236)) + ((g59) & (!g50) & (!g154) & (g93) & (!sk[119]) & (!g236)) + ((g59) & (!g50) & (!g154) & (g93) & (!sk[119]) & (g236)) + ((g59) & (!g50) & (g154) & (!g93) & (!sk[119]) & (!g236)) + ((g59) & (!g50) & (g154) & (!g93) & (!sk[119]) & (g236)) + ((g59) & (!g50) & (g154) & (g93) & (!sk[119]) & (!g236)) + ((g59) & (!g50) & (g154) & (g93) & (!sk[119]) & (g236)) + ((g59) & (g50) & (!g154) & (!g93) & (!sk[119]) & (!g236)) + ((g59) & (g50) & (!g154) & (!g93) & (!sk[119]) & (g236)) + ((g59) & (g50) & (!g154) & (g93) & (!sk[119]) & (!g236)) + ((g59) & (g50) & (!g154) & (g93) & (!sk[119]) & (g236)) + ((g59) & (g50) & (g154) & (!g93) & (!sk[119]) & (!g236)) + ((g59) & (g50) & (g154) & (!g93) & (!sk[119]) & (g236)) + ((g59) & (g50) & (g154) & (g93) & (!sk[119]) & (!g236)) + ((g59) & (g50) & (g154) & (g93) & (!sk[119]) & (g236)));
	assign g238 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g12)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g12)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g12)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g12)));
	assign g239 = (((!g16) & (!g30) & (!g238) & (!g153) & (!g83) & (!g63)) + ((!g16) & (g30) & (!g238) & (!g153) & (!g83) & (!g63)) + ((g16) & (!g30) & (!g238) & (!g153) & (!g83) & (!g63)));
	assign g240 = (((g230) & (g231) & (!g232) & (g235) & (g237) & (g239)));
	assign g241 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g42)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g42)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g42)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g42)));
	assign g242 = (((!g70) & (!g99) & (!g241) & (!g32) & (!g20) & (!g193)) + ((!g70) & (!g99) & (!g241) & (!g32) & (g20) & (!g193)) + ((!g70) & (!g99) & (!g241) & (g32) & (!g20) & (!g193)) + ((!g70) & (!g99) & (!g241) & (g32) & (g20) & (!g193)) + ((!g70) & (g99) & (!g241) & (!g32) & (!g20) & (!g193)) + ((!g70) & (g99) & (!g241) & (g32) & (!g20) & (!g193)) + ((g70) & (!g99) & (!g241) & (!g32) & (!g20) & (!g193)) + ((g70) & (!g99) & (!g241) & (!g32) & (g20) & (!g193)) + ((g70) & (g99) & (!g241) & (!g32) & (!g20) & (!g193)));
	assign g243 = (((!sk[125]) & (!g99) & (!g71) & (g42) & (!g87)) + ((!sk[125]) & (!g99) & (!g71) & (g42) & (g87)) + ((!sk[125]) & (!g99) & (g71) & (g42) & (!g87)) + ((!sk[125]) & (!g99) & (g71) & (g42) & (g87)) + ((!sk[125]) & (g99) & (!g71) & (!g42) & (!g87)) + ((!sk[125]) & (g99) & (!g71) & (!g42) & (g87)) + ((!sk[125]) & (g99) & (!g71) & (g42) & (!g87)) + ((!sk[125]) & (g99) & (!g71) & (g42) & (g87)) + ((!sk[125]) & (g99) & (g71) & (!g42) & (!g87)) + ((!sk[125]) & (g99) & (g71) & (!g42) & (g87)) + ((!sk[125]) & (g99) & (g71) & (g42) & (!g87)) + ((!sk[125]) & (g99) & (g71) & (g42) & (g87)) + ((sk[125]) & (!g99) & (!g71) & (!g42) & (!g87)) + ((sk[125]) & (!g99) & (!g71) & (g42) & (!g87)) + ((sk[125]) & (!g99) & (g71) & (!g42) & (!g87)) + ((sk[125]) & (g99) & (!g71) & (!g42) & (!g87)) + ((sk[125]) & (g99) & (g71) & (!g42) & (!g87)));
	assign g244 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g30)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (g8) & (g30)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g30)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (g8) & (g30)));
	assign g245 = (((!g99) & (!g12) & (!g26) & (!g11) & (!g244) & (!g55)) + ((!g99) & (g12) & (!g26) & (!g11) & (!g244) & (!g55)) + ((g99) & (!g12) & (!g26) & (!g11) & (!g244) & (!g55)));
	assign g246 = (((!g49) & (!g99) & (!g62) & (!g32) & (!g124) & (!g95)) + ((!g49) & (!g99) & (!g62) & (g32) & (!g124) & (!g95)) + ((!g49) & (!g99) & (g62) & (!g32) & (!g124) & (!g95)) + ((!g49) & (g99) & (!g62) & (!g32) & (!g124) & (!g95)) + ((!g49) & (g99) & (g62) & (!g32) & (!g124) & (!g95)) + ((g49) & (!g99) & (!g62) & (!g32) & (!g124) & (!g95)) + ((g49) & (!g99) & (!g62) & (g32) & (!g124) & (!g95)) + ((g49) & (g99) & (!g62) & (!g32) & (!g124) & (!g95)));
	assign g247 = (((!ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)) + ((!ax19x) & (!ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (ax16x) & (!g5) & (ax18x)) + ((!ax19x) & (ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (ax16x) & (!g5) & (!ax18x)) + ((!ax19x) & (ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (!ax22x) & (!ax17x) & (ax16x) & (g5) & (ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (!ax16x) & (!g5) & (!ax18x)) + ((ax19x) & (!ax22x) & (ax17x) & (ax16x) & (g5) & (!ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (!g5) & (ax18x)) + ((ax19x) & (ax22x) & (!ax17x) & (!ax16x) & (g5) & (ax18x)));
	assign g248 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g247)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g247)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g247)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g247)));
	assign g249 = (((!g62) & (!g18) & (!g104) & (!g25) & (!g27) & (!g248)) + ((!g62) & (!g18) & (!g104) & (!g25) & (g27) & (!g248)) + ((!g62) & (!g18) & (!g104) & (g25) & (!g27) & (!g248)) + ((!g62) & (!g18) & (!g104) & (g25) & (g27) & (!g248)) + ((!g62) & (!g18) & (g104) & (!g25) & (!g27) & (!g248)) + ((!g62) & (g18) & (!g104) & (!g25) & (!g27) & (!g248)) + ((!g62) & (g18) & (!g104) & (!g25) & (g27) & (!g248)) + ((!g62) & (g18) & (!g104) & (g25) & (!g27) & (!g248)) + ((!g62) & (g18) & (!g104) & (g25) & (g27) & (!g248)) + ((!g62) & (g18) & (g104) & (!g25) & (!g27) & (!g248)) + ((g62) & (!g18) & (!g104) & (!g25) & (!g27) & (!g248)) + ((g62) & (!g18) & (!g104) & (g25) & (!g27) & (!g248)) + ((g62) & (!g18) & (g104) & (!g25) & (!g27) & (!g248)));
	assign g250 = (((!g71) & (!g20) & (g243) & (g245) & (g246) & (g249)) + ((!g71) & (g20) & (g243) & (g245) & (g246) & (g249)) + ((g71) & (!g20) & (g243) & (g245) & (g246) & (g249)));
	assign g251 = (((g224) & (g228) & (g229) & (g240) & (g242) & (g250)));
	assign g252 = (((!sk[6]) & (!ax22x) & (!g7) & (ax14x)) + ((!sk[6]) & (!ax22x) & (g7) & (ax14x)) + ((!sk[6]) & (ax22x) & (!g7) & (!ax14x)) + ((!sk[6]) & (ax22x) & (!g7) & (ax14x)) + ((!sk[6]) & (ax22x) & (g7) & (!ax14x)) + ((!sk[6]) & (ax22x) & (g7) & (ax14x)) + ((sk[6]) & (!ax22x) & (!g7) & (!ax14x)) + ((sk[6]) & (!ax22x) & (g7) & (ax14x)) + ((sk[6]) & (ax22x) & (!g7) & (ax14x)) + ((sk[6]) & (ax22x) & (g7) & (ax14x)));
	assign g253 = (((!ax22x) & (!ax13x) & (!ax11x) & (!sk[7]) & (g4) & (!ax12x)) + ((!ax22x) & (!ax13x) & (!ax11x) & (!sk[7]) & (g4) & (ax12x)) + ((!ax22x) & (!ax13x) & (!ax11x) & (sk[7]) & (!g4) & (!ax12x)) + ((!ax22x) & (!ax13x) & (!ax11x) & (sk[7]) & (!g4) & (ax12x)) + ((!ax22x) & (!ax13x) & (!ax11x) & (sk[7]) & (g4) & (ax12x)) + ((!ax22x) & (!ax13x) & (ax11x) & (!sk[7]) & (g4) & (!ax12x)) + ((!ax22x) & (!ax13x) & (ax11x) & (!sk[7]) & (g4) & (ax12x)) + ((!ax22x) & (!ax13x) & (ax11x) & (sk[7]) & (!g4) & (!ax12x)) + ((!ax22x) & (!ax13x) & (ax11x) & (sk[7]) & (!g4) & (ax12x)) + ((!ax22x) & (!ax13x) & (ax11x) & (sk[7]) & (g4) & (!ax12x)) + ((!ax22x) & (!ax13x) & (ax11x) & (sk[7]) & (g4) & (ax12x)) + ((!ax22x) & (ax13x) & (!ax11x) & (!sk[7]) & (!g4) & (!ax12x)) + ((!ax22x) & (ax13x) & (!ax11x) & (!sk[7]) & (!g4) & (ax12x)) + ((!ax22x) & (ax13x) & (!ax11x) & (!sk[7]) & (g4) & (!ax12x)) + ((!ax22x) & (ax13x) & (!ax11x) & (!sk[7]) & (g4) & (ax12x)) + ((!ax22x) & (ax13x) & (!ax11x) & (sk[7]) & (g4) & (!ax12x)) + ((!ax22x) & (ax13x) & (ax11x) & (!sk[7]) & (!g4) & (!ax12x)) + ((!ax22x) & (ax13x) & (ax11x) & (!sk[7]) & (!g4) & (ax12x)) + ((!ax22x) & (ax13x) & (ax11x) & (!sk[7]) & (g4) & (!ax12x)) + ((!ax22x) & (ax13x) & (ax11x) & (!sk[7]) & (g4) & (ax12x)) + ((ax22x) & (!ax13x) & (!ax11x) & (!sk[7]) & (g4) & (!ax12x)) + ((ax22x) & (!ax13x) & (!ax11x) & (!sk[7]) & (g4) & (ax12x)) + ((ax22x) & (!ax13x) & (ax11x) & (!sk[7]) & (!g4) & (!ax12x)) + ((ax22x) & (!ax13x) & (ax11x) & (!sk[7]) & (!g4) & (ax12x)) + ((ax22x) & (!ax13x) & (ax11x) & (!sk[7]) & (g4) & (!ax12x)) + ((ax22x) & (!ax13x) & (ax11x) & (!sk[7]) & (g4) & (ax12x)) + ((ax22x) & (ax13x) & (!ax11x) & (!sk[7]) & (!g4) & (!ax12x)) + ((ax22x) & (ax13x) & (!ax11x) & (!sk[7]) & (!g4) & (ax12x)) + ((ax22x) & (ax13x) & (!ax11x) & (!sk[7]) & (g4) & (!ax12x)) + ((ax22x) & (ax13x) & (!ax11x) & (!sk[7]) & (g4) & (ax12x)) + ((ax22x) & (ax13x) & (!ax11x) & (sk[7]) & (!g4) & (!ax12x)) + ((ax22x) & (ax13x) & (!ax11x) & (sk[7]) & (!g4) & (ax12x)) + ((ax22x) & (ax13x) & (!ax11x) & (sk[7]) & (g4) & (!ax12x)) + ((ax22x) & (ax13x) & (!ax11x) & (sk[7]) & (g4) & (ax12x)) + ((ax22x) & (ax13x) & (ax11x) & (!sk[7]) & (!g4) & (!ax12x)) + ((ax22x) & (ax13x) & (ax11x) & (!sk[7]) & (!g4) & (ax12x)) + ((ax22x) & (ax13x) & (ax11x) & (!sk[7]) & (g4) & (!ax12x)) + ((ax22x) & (ax13x) & (ax11x) & (!sk[7]) & (g4) & (ax12x)) + ((ax22x) & (ax13x) & (ax11x) & (sk[7]) & (!g4) & (!ax12x)) + ((ax22x) & (ax13x) & (ax11x) & (sk[7]) & (!g4) & (ax12x)) + ((ax22x) & (ax13x) & (ax11x) & (sk[7]) & (g4) & (!ax12x)) + ((ax22x) & (ax13x) & (ax11x) & (sk[7]) & (g4) & (ax12x)));
	assign g254 = (((!g17) & (!g99) & (g71) & (!sk[8]) & (!g32)) + ((!g17) & (!g99) & (g71) & (!sk[8]) & (g32)) + ((!g17) & (g99) & (!g71) & (sk[8]) & (g32)) + ((!g17) & (g99) & (g71) & (!sk[8]) & (!g32)) + ((!g17) & (g99) & (g71) & (!sk[8]) & (g32)) + ((!g17) & (g99) & (g71) & (sk[8]) & (g32)) + ((g17) & (!g99) & (!g71) & (!sk[8]) & (!g32)) + ((g17) & (!g99) & (!g71) & (!sk[8]) & (g32)) + ((g17) & (!g99) & (g71) & (!sk[8]) & (!g32)) + ((g17) & (!g99) & (g71) & (!sk[8]) & (g32)) + ((g17) & (!g99) & (g71) & (sk[8]) & (!g32)) + ((g17) & (!g99) & (g71) & (sk[8]) & (g32)) + ((g17) & (g99) & (!g71) & (!sk[8]) & (!g32)) + ((g17) & (g99) & (!g71) & (!sk[8]) & (g32)) + ((g17) & (g99) & (!g71) & (sk[8]) & (g32)) + ((g17) & (g99) & (g71) & (!sk[8]) & (!g32)) + ((g17) & (g99) & (g71) & (!sk[8]) & (g32)) + ((g17) & (g99) & (g71) & (sk[8]) & (!g32)) + ((g17) & (g99) & (g71) & (sk[8]) & (g32)));
	assign g255 = (((!g38) & (!sk[9]) & (!g16) & (!g49) & (g62) & (!g41)) + ((!g38) & (!sk[9]) & (!g16) & (!g49) & (g62) & (g41)) + ((!g38) & (!sk[9]) & (!g16) & (g49) & (g62) & (!g41)) + ((!g38) & (!sk[9]) & (!g16) & (g49) & (g62) & (g41)) + ((!g38) & (!sk[9]) & (g16) & (!g49) & (!g62) & (!g41)) + ((!g38) & (!sk[9]) & (g16) & (!g49) & (!g62) & (g41)) + ((!g38) & (!sk[9]) & (g16) & (!g49) & (g62) & (!g41)) + ((!g38) & (!sk[9]) & (g16) & (!g49) & (g62) & (g41)) + ((!g38) & (!sk[9]) & (g16) & (g49) & (!g62) & (!g41)) + ((!g38) & (!sk[9]) & (g16) & (g49) & (!g62) & (g41)) + ((!g38) & (!sk[9]) & (g16) & (g49) & (g62) & (!g41)) + ((!g38) & (!sk[9]) & (g16) & (g49) & (g62) & (g41)) + ((!g38) & (sk[9]) & (!g16) & (!g49) & (!g62) & (!g41)) + ((!g38) & (sk[9]) & (!g16) & (!g49) & (!g62) & (g41)) + ((!g38) & (sk[9]) & (!g16) & (!g49) & (g62) & (!g41)) + ((!g38) & (sk[9]) & (!g16) & (!g49) & (g62) & (g41)) + ((!g38) & (sk[9]) & (!g16) & (g49) & (!g62) & (!g41)) + ((!g38) & (sk[9]) & (!g16) & (g49) & (!g62) & (g41)) + ((!g38) & (sk[9]) & (g16) & (!g49) & (!g62) & (!g41)) + ((!g38) & (sk[9]) & (g16) & (!g49) & (g62) & (!g41)) + ((!g38) & (sk[9]) & (g16) & (g49) & (!g62) & (!g41)) + ((g38) & (!sk[9]) & (!g16) & (!g49) & (g62) & (!g41)) + ((g38) & (!sk[9]) & (!g16) & (!g49) & (g62) & (g41)) + ((g38) & (!sk[9]) & (!g16) & (g49) & (!g62) & (!g41)) + ((g38) & (!sk[9]) & (!g16) & (g49) & (!g62) & (g41)) + ((g38) & (!sk[9]) & (!g16) & (g49) & (g62) & (!g41)) + ((g38) & (!sk[9]) & (!g16) & (g49) & (g62) & (g41)) + ((g38) & (!sk[9]) & (g16) & (!g49) & (!g62) & (!g41)) + ((g38) & (!sk[9]) & (g16) & (!g49) & (!g62) & (g41)) + ((g38) & (!sk[9]) & (g16) & (!g49) & (g62) & (!g41)) + ((g38) & (!sk[9]) & (g16) & (!g49) & (g62) & (g41)) + ((g38) & (!sk[9]) & (g16) & (g49) & (!g62) & (!g41)) + ((g38) & (!sk[9]) & (g16) & (g49) & (!g62) & (g41)) + ((g38) & (!sk[9]) & (g16) & (g49) & (g62) & (!g41)) + ((g38) & (!sk[9]) & (g16) & (g49) & (g62) & (g41)) + ((g38) & (sk[9]) & (!g16) & (!g49) & (!g62) & (!g41)) + ((g38) & (sk[9]) & (!g16) & (!g49) & (!g62) & (g41)) + ((g38) & (sk[9]) & (!g16) & (!g49) & (g62) & (!g41)) + ((g38) & (sk[9]) & (!g16) & (!g49) & (g62) & (g41)) + ((g38) & (sk[9]) & (!g16) & (g49) & (!g62) & (!g41)) + ((g38) & (sk[9]) & (!g16) & (g49) & (!g62) & (g41)));
	assign g256 = (((!g38) & (!g9) & (!g17) & (!g99) & (!g80) & (!g64)) + ((!g38) & (!g9) & (!g17) & (g99) & (!g80) & (!g64)) + ((!g38) & (!g9) & (g17) & (!g99) & (!g80) & (!g64)) + ((!g38) & (g9) & (!g17) & (!g99) & (!g80) & (!g64)) + ((!g38) & (g9) & (!g17) & (g99) & (!g80) & (!g64)) + ((!g38) & (g9) & (g17) & (!g99) & (!g80) & (!g64)) + ((g38) & (!g9) & (!g17) & (!g99) & (!g80) & (!g64)) + ((g38) & (!g9) & (!g17) & (g99) & (!g80) & (!g64)) + ((g38) & (!g9) & (g17) & (!g99) & (!g80) & (!g64)));
	assign g257 = (((!ax22x) & (!g6) & (!sk[11]) & (!ax20x) & (g8) & (!g49)) + ((!ax22x) & (!g6) & (!sk[11]) & (!ax20x) & (g8) & (g49)) + ((!ax22x) & (!g6) & (!sk[11]) & (ax20x) & (g8) & (!g49)) + ((!ax22x) & (!g6) & (!sk[11]) & (ax20x) & (g8) & (g49)) + ((!ax22x) & (!g6) & (sk[11]) & (ax20x) & (!g8) & (g49)) + ((!ax22x) & (g6) & (!sk[11]) & (!ax20x) & (!g8) & (!g49)) + ((!ax22x) & (g6) & (!sk[11]) & (!ax20x) & (!g8) & (g49)) + ((!ax22x) & (g6) & (!sk[11]) & (!ax20x) & (g8) & (!g49)) + ((!ax22x) & (g6) & (!sk[11]) & (!ax20x) & (g8) & (g49)) + ((!ax22x) & (g6) & (!sk[11]) & (ax20x) & (!g8) & (!g49)) + ((!ax22x) & (g6) & (!sk[11]) & (ax20x) & (!g8) & (g49)) + ((!ax22x) & (g6) & (!sk[11]) & (ax20x) & (g8) & (!g49)) + ((!ax22x) & (g6) & (!sk[11]) & (ax20x) & (g8) & (g49)) + ((!ax22x) & (g6) & (sk[11]) & (!ax20x) & (!g8) & (g49)) + ((ax22x) & (!g6) & (!sk[11]) & (!ax20x) & (g8) & (!g49)) + ((ax22x) & (!g6) & (!sk[11]) & (!ax20x) & (g8) & (g49)) + ((ax22x) & (!g6) & (!sk[11]) & (ax20x) & (!g8) & (!g49)) + ((ax22x) & (!g6) & (!sk[11]) & (ax20x) & (!g8) & (g49)) + ((ax22x) & (!g6) & (!sk[11]) & (ax20x) & (g8) & (!g49)) + ((ax22x) & (!g6) & (!sk[11]) & (ax20x) & (g8) & (g49)) + ((ax22x) & (!g6) & (sk[11]) & (!ax20x) & (!g8) & (g49)) + ((ax22x) & (g6) & (!sk[11]) & (!ax20x) & (!g8) & (!g49)) + ((ax22x) & (g6) & (!sk[11]) & (!ax20x) & (!g8) & (g49)) + ((ax22x) & (g6) & (!sk[11]) & (!ax20x) & (g8) & (!g49)) + ((ax22x) & (g6) & (!sk[11]) & (!ax20x) & (g8) & (g49)) + ((ax22x) & (g6) & (!sk[11]) & (ax20x) & (!g8) & (!g49)) + ((ax22x) & (g6) & (!sk[11]) & (ax20x) & (!g8) & (g49)) + ((ax22x) & (g6) & (!sk[11]) & (ax20x) & (g8) & (!g49)) + ((ax22x) & (g6) & (!sk[11]) & (ax20x) & (g8) & (g49)) + ((ax22x) & (g6) & (sk[11]) & (!ax20x) & (!g8) & (g49)));
	assign g258 = (((!g9) & (!g23) & (!g18) & (!sk[12]) & (g27) & (!g257)) + ((!g9) & (!g23) & (!g18) & (!sk[12]) & (g27) & (g257)) + ((!g9) & (!g23) & (!g18) & (sk[12]) & (!g27) & (!g257)) + ((!g9) & (!g23) & (!g18) & (sk[12]) & (g27) & (!g257)) + ((!g9) & (!g23) & (g18) & (!sk[12]) & (g27) & (!g257)) + ((!g9) & (!g23) & (g18) & (!sk[12]) & (g27) & (g257)) + ((!g9) & (!g23) & (g18) & (sk[12]) & (!g27) & (!g257)) + ((!g9) & (!g23) & (g18) & (sk[12]) & (g27) & (!g257)) + ((!g9) & (g23) & (!g18) & (!sk[12]) & (!g27) & (!g257)) + ((!g9) & (g23) & (!g18) & (!sk[12]) & (!g27) & (g257)) + ((!g9) & (g23) & (!g18) & (!sk[12]) & (g27) & (!g257)) + ((!g9) & (g23) & (!g18) & (!sk[12]) & (g27) & (g257)) + ((!g9) & (g23) & (!g18) & (sk[12]) & (!g27) & (!g257)) + ((!g9) & (g23) & (!g18) & (sk[12]) & (g27) & (!g257)) + ((!g9) & (g23) & (g18) & (!sk[12]) & (!g27) & (!g257)) + ((!g9) & (g23) & (g18) & (!sk[12]) & (!g27) & (g257)) + ((!g9) & (g23) & (g18) & (!sk[12]) & (g27) & (!g257)) + ((!g9) & (g23) & (g18) & (!sk[12]) & (g27) & (g257)) + ((!g9) & (g23) & (g18) & (sk[12]) & (!g27) & (!g257)) + ((!g9) & (g23) & (g18) & (sk[12]) & (g27) & (!g257)) + ((g9) & (!g23) & (!g18) & (!sk[12]) & (g27) & (!g257)) + ((g9) & (!g23) & (!g18) & (!sk[12]) & (g27) & (g257)) + ((g9) & (!g23) & (!g18) & (sk[12]) & (!g27) & (!g257)) + ((g9) & (!g23) & (g18) & (!sk[12]) & (!g27) & (!g257)) + ((g9) & (!g23) & (g18) & (!sk[12]) & (!g27) & (g257)) + ((g9) & (!g23) & (g18) & (!sk[12]) & (g27) & (!g257)) + ((g9) & (!g23) & (g18) & (!sk[12]) & (g27) & (g257)) + ((g9) & (g23) & (!g18) & (!sk[12]) & (!g27) & (!g257)) + ((g9) & (g23) & (!g18) & (!sk[12]) & (!g27) & (g257)) + ((g9) & (g23) & (!g18) & (!sk[12]) & (g27) & (!g257)) + ((g9) & (g23) & (!g18) & (!sk[12]) & (g27) & (g257)) + ((g9) & (g23) & (g18) & (!sk[12]) & (!g27) & (!g257)) + ((g9) & (g23) & (g18) & (!sk[12]) & (!g27) & (g257)) + ((g9) & (g23) & (g18) & (!sk[12]) & (g27) & (!g257)) + ((g9) & (g23) & (g18) & (!sk[12]) & (g27) & (g257)));
	assign g259 = (((!g95) & (!g254) & (g255) & (g256) & (g258) & (g151)));
	assign g260 = (((!g16) & (!g30) & (!sk[14]) & (g131)) + ((!g16) & (!g30) & (sk[14]) & (!g131)) + ((!g16) & (g30) & (!sk[14]) & (g131)) + ((!g16) & (g30) & (sk[14]) & (!g131)) + ((g16) & (!g30) & (!sk[14]) & (!g131)) + ((g16) & (!g30) & (!sk[14]) & (g131)) + ((g16) & (!g30) & (sk[14]) & (!g131)) + ((g16) & (g30) & (!sk[14]) & (!g131)) + ((g16) & (g30) & (!sk[14]) & (g131)));
	assign g261 = (((!g9) & (!g66) & (!sk[15]) & (g29)) + ((!g9) & (!g66) & (sk[15]) & (!g29)) + ((!g9) & (g66) & (!sk[15]) & (g29)) + ((!g9) & (g66) & (sk[15]) & (!g29)) + ((g9) & (!g66) & (!sk[15]) & (!g29)) + ((g9) & (!g66) & (!sk[15]) & (g29)) + ((g9) & (!g66) & (sk[15]) & (!g29)) + ((g9) & (g66) & (!sk[15]) & (!g29)) + ((g9) & (g66) & (!sk[15]) & (g29)));
	assign g262 = (((!sk[16]) & (!g9) & (!g16) & (!g12) & (g25) & (!g85)) + ((!sk[16]) & (!g9) & (!g16) & (!g12) & (g25) & (g85)) + ((!sk[16]) & (!g9) & (!g16) & (g12) & (g25) & (!g85)) + ((!sk[16]) & (!g9) & (!g16) & (g12) & (g25) & (g85)) + ((!sk[16]) & (!g9) & (g16) & (!g12) & (!g25) & (!g85)) + ((!sk[16]) & (!g9) & (g16) & (!g12) & (!g25) & (g85)) + ((!sk[16]) & (!g9) & (g16) & (!g12) & (g25) & (!g85)) + ((!sk[16]) & (!g9) & (g16) & (!g12) & (g25) & (g85)) + ((!sk[16]) & (!g9) & (g16) & (g12) & (!g25) & (!g85)) + ((!sk[16]) & (!g9) & (g16) & (g12) & (!g25) & (g85)) + ((!sk[16]) & (!g9) & (g16) & (g12) & (g25) & (!g85)) + ((!sk[16]) & (!g9) & (g16) & (g12) & (g25) & (g85)) + ((!sk[16]) & (g9) & (!g16) & (!g12) & (g25) & (!g85)) + ((!sk[16]) & (g9) & (!g16) & (!g12) & (g25) & (g85)) + ((!sk[16]) & (g9) & (!g16) & (g12) & (!g25) & (!g85)) + ((!sk[16]) & (g9) & (!g16) & (g12) & (!g25) & (g85)) + ((!sk[16]) & (g9) & (!g16) & (g12) & (g25) & (!g85)) + ((!sk[16]) & (g9) & (!g16) & (g12) & (g25) & (g85)) + ((!sk[16]) & (g9) & (g16) & (!g12) & (!g25) & (!g85)) + ((!sk[16]) & (g9) & (g16) & (!g12) & (!g25) & (g85)) + ((!sk[16]) & (g9) & (g16) & (!g12) & (g25) & (!g85)) + ((!sk[16]) & (g9) & (g16) & (!g12) & (g25) & (g85)) + ((!sk[16]) & (g9) & (g16) & (g12) & (!g25) & (!g85)) + ((!sk[16]) & (g9) & (g16) & (g12) & (!g25) & (g85)) + ((!sk[16]) & (g9) & (g16) & (g12) & (g25) & (!g85)) + ((!sk[16]) & (g9) & (g16) & (g12) & (g25) & (g85)) + ((sk[16]) & (!g9) & (!g16) & (!g12) & (!g25) & (!g85)) + ((sk[16]) & (!g9) & (!g16) & (!g12) & (g25) & (!g85)) + ((sk[16]) & (!g9) & (!g16) & (g12) & (!g25) & (!g85)) + ((sk[16]) & (!g9) & (!g16) & (g12) & (g25) & (!g85)) + ((sk[16]) & (!g9) & (g16) & (!g12) & (!g25) & (!g85)) + ((sk[16]) & (!g9) & (g16) & (!g12) & (g25) & (!g85)) + ((sk[16]) & (g9) & (!g16) & (!g12) & (!g25) & (!g85)) + ((sk[16]) & (g9) & (!g16) & (g12) & (!g25) & (!g85)) + ((sk[16]) & (g9) & (g16) & (!g12) & (!g25) & (!g85)));
	assign g263 = (((!g114) & (!g115) & (g8) & (g12) & (!g25) & (!g42)) + ((!g114) & (!g115) & (g8) & (g12) & (!g25) & (g42)) + ((!g114) & (!g115) & (g8) & (g12) & (g25) & (!g42)) + ((!g114) & (!g115) & (g8) & (g12) & (g25) & (g42)) + ((!g114) & (g115) & (!g8) & (!g12) & (!g25) & (g42)) + ((!g114) & (g115) & (!g8) & (!g12) & (g25) & (g42)) + ((!g114) & (g115) & (!g8) & (g12) & (!g25) & (g42)) + ((!g114) & (g115) & (!g8) & (g12) & (g25) & (g42)) + ((!g114) & (g115) & (g8) & (g12) & (!g25) & (!g42)) + ((!g114) & (g115) & (g8) & (g12) & (!g25) & (g42)) + ((!g114) & (g115) & (g8) & (g12) & (g25) & (!g42)) + ((!g114) & (g115) & (g8) & (g12) & (g25) & (g42)) + ((g114) & (!g115) & (g8) & (!g12) & (g25) & (!g42)) + ((g114) & (!g115) & (g8) & (!g12) & (g25) & (g42)) + ((g114) & (!g115) & (g8) & (g12) & (g25) & (!g42)) + ((g114) & (!g115) & (g8) & (g12) & (g25) & (g42)));
	assign g264 = (((!g38) & (!sk[18]) & (!g62) & (!g147) & (g36) & (!g81)) + ((!g38) & (!sk[18]) & (!g62) & (!g147) & (g36) & (g81)) + ((!g38) & (!sk[18]) & (!g62) & (g147) & (g36) & (!g81)) + ((!g38) & (!sk[18]) & (!g62) & (g147) & (g36) & (g81)) + ((!g38) & (!sk[18]) & (g62) & (!g147) & (!g36) & (!g81)) + ((!g38) & (!sk[18]) & (g62) & (!g147) & (!g36) & (g81)) + ((!g38) & (!sk[18]) & (g62) & (!g147) & (g36) & (!g81)) + ((!g38) & (!sk[18]) & (g62) & (!g147) & (g36) & (g81)) + ((!g38) & (!sk[18]) & (g62) & (g147) & (!g36) & (!g81)) + ((!g38) & (!sk[18]) & (g62) & (g147) & (!g36) & (g81)) + ((!g38) & (!sk[18]) & (g62) & (g147) & (g36) & (!g81)) + ((!g38) & (!sk[18]) & (g62) & (g147) & (g36) & (g81)) + ((!g38) & (sk[18]) & (!g62) & (!g147) & (!g36) & (!g81)) + ((!g38) & (sk[18]) & (g62) & (!g147) & (!g36) & (!g81)) + ((g38) & (!sk[18]) & (!g62) & (!g147) & (g36) & (!g81)) + ((g38) & (!sk[18]) & (!g62) & (!g147) & (g36) & (g81)) + ((g38) & (!sk[18]) & (!g62) & (g147) & (!g36) & (!g81)) + ((g38) & (!sk[18]) & (!g62) & (g147) & (!g36) & (g81)) + ((g38) & (!sk[18]) & (!g62) & (g147) & (g36) & (!g81)) + ((g38) & (!sk[18]) & (!g62) & (g147) & (g36) & (g81)) + ((g38) & (!sk[18]) & (g62) & (!g147) & (!g36) & (!g81)) + ((g38) & (!sk[18]) & (g62) & (!g147) & (!g36) & (g81)) + ((g38) & (!sk[18]) & (g62) & (!g147) & (g36) & (!g81)) + ((g38) & (!sk[18]) & (g62) & (!g147) & (g36) & (g81)) + ((g38) & (!sk[18]) & (g62) & (g147) & (!g36) & (!g81)) + ((g38) & (!sk[18]) & (g62) & (g147) & (!g36) & (g81)) + ((g38) & (!sk[18]) & (g62) & (g147) & (g36) & (!g81)) + ((g38) & (!sk[18]) & (g62) & (g147) & (g36) & (g81)) + ((g38) & (sk[18]) & (!g62) & (!g147) & (!g36) & (!g81)));
	assign g265 = (((!g38) & (!g99) & (!sk[19]) & (!g104) & (g25) & (!g33)) + ((!g38) & (!g99) & (!sk[19]) & (!g104) & (g25) & (g33)) + ((!g38) & (!g99) & (!sk[19]) & (g104) & (g25) & (!g33)) + ((!g38) & (!g99) & (!sk[19]) & (g104) & (g25) & (g33)) + ((!g38) & (!g99) & (sk[19]) & (!g104) & (!g25) & (!g33)) + ((!g38) & (!g99) & (sk[19]) & (!g104) & (g25) & (!g33)) + ((!g38) & (!g99) & (sk[19]) & (g104) & (!g25) & (!g33)) + ((!g38) & (g99) & (!sk[19]) & (!g104) & (!g25) & (!g33)) + ((!g38) & (g99) & (!sk[19]) & (!g104) & (!g25) & (g33)) + ((!g38) & (g99) & (!sk[19]) & (!g104) & (g25) & (!g33)) + ((!g38) & (g99) & (!sk[19]) & (!g104) & (g25) & (g33)) + ((!g38) & (g99) & (!sk[19]) & (g104) & (!g25) & (!g33)) + ((!g38) & (g99) & (!sk[19]) & (g104) & (!g25) & (g33)) + ((!g38) & (g99) & (!sk[19]) & (g104) & (g25) & (!g33)) + ((!g38) & (g99) & (!sk[19]) & (g104) & (g25) & (g33)) + ((!g38) & (g99) & (sk[19]) & (!g104) & (!g25) & (!g33)) + ((!g38) & (g99) & (sk[19]) & (g104) & (!g25) & (!g33)) + ((g38) & (!g99) & (!sk[19]) & (!g104) & (g25) & (!g33)) + ((g38) & (!g99) & (!sk[19]) & (!g104) & (g25) & (g33)) + ((g38) & (!g99) & (!sk[19]) & (g104) & (!g25) & (!g33)) + ((g38) & (!g99) & (!sk[19]) & (g104) & (!g25) & (g33)) + ((g38) & (!g99) & (!sk[19]) & (g104) & (g25) & (!g33)) + ((g38) & (!g99) & (!sk[19]) & (g104) & (g25) & (g33)) + ((g38) & (!g99) & (sk[19]) & (!g104) & (!g25) & (!g33)) + ((g38) & (!g99) & (sk[19]) & (!g104) & (g25) & (!g33)) + ((g38) & (g99) & (!sk[19]) & (!g104) & (!g25) & (!g33)) + ((g38) & (g99) & (!sk[19]) & (!g104) & (!g25) & (g33)) + ((g38) & (g99) & (!sk[19]) & (!g104) & (g25) & (!g33)) + ((g38) & (g99) & (!sk[19]) & (!g104) & (g25) & (g33)) + ((g38) & (g99) & (!sk[19]) & (g104) & (!g25) & (!g33)) + ((g38) & (g99) & (!sk[19]) & (g104) & (!g25) & (g33)) + ((g38) & (g99) & (!sk[19]) & (g104) & (g25) & (!g33)) + ((g38) & (g99) & (!sk[19]) & (g104) & (g25) & (g33)) + ((g38) & (g99) & (sk[19]) & (!g104) & (!g25) & (!g33)));
	assign g266 = (((g260) & (g261) & (g262) & (!g263) & (g264) & (g265)));
	assign g267 = (((!ax22x) & (g38) & (ax21x) & (!g6) & (!ax20x) & (g8)) + ((!ax22x) & (g38) & (ax21x) & (g6) & (ax20x) & (g8)) + ((ax22x) & (g38) & (!ax21x) & (!g6) & (ax20x) & (g8)) + ((ax22x) & (g38) & (!ax21x) & (g6) & (ax20x) & (g8)));
	assign g268 = (((!sk[22]) & (!g62) & (!g104) & (g41) & (!g27)) + ((!sk[22]) & (!g62) & (!g104) & (g41) & (g27)) + ((!sk[22]) & (!g62) & (g104) & (g41) & (!g27)) + ((!sk[22]) & (!g62) & (g104) & (g41) & (g27)) + ((!sk[22]) & (g62) & (!g104) & (!g41) & (!g27)) + ((!sk[22]) & (g62) & (!g104) & (!g41) & (g27)) + ((!sk[22]) & (g62) & (!g104) & (g41) & (!g27)) + ((!sk[22]) & (g62) & (!g104) & (g41) & (g27)) + ((!sk[22]) & (g62) & (g104) & (!g41) & (!g27)) + ((!sk[22]) & (g62) & (g104) & (!g41) & (g27)) + ((!sk[22]) & (g62) & (g104) & (g41) & (!g27)) + ((!sk[22]) & (g62) & (g104) & (g41) & (g27)) + ((sk[22]) & (!g62) & (g104) & (!g41) & (g27)) + ((sk[22]) & (!g62) & (g104) & (g41) & (g27)) + ((sk[22]) & (g62) & (!g104) & (g41) & (!g27)) + ((sk[22]) & (g62) & (!g104) & (g41) & (g27)) + ((sk[22]) & (g62) & (g104) & (!g41) & (g27)) + ((sk[22]) & (g62) & (g104) & (g41) & (!g27)) + ((sk[22]) & (g62) & (g104) & (g41) & (g27)));
	assign g269 = (((!sk[23]) & (!g78) & (!g104) & (g41) & (!g32)) + ((!sk[23]) & (!g78) & (!g104) & (g41) & (g32)) + ((!sk[23]) & (!g78) & (g104) & (g41) & (!g32)) + ((!sk[23]) & (!g78) & (g104) & (g41) & (g32)) + ((!sk[23]) & (g78) & (!g104) & (!g41) & (!g32)) + ((!sk[23]) & (g78) & (!g104) & (!g41) & (g32)) + ((!sk[23]) & (g78) & (!g104) & (g41) & (!g32)) + ((!sk[23]) & (g78) & (!g104) & (g41) & (g32)) + ((!sk[23]) & (g78) & (g104) & (!g41) & (!g32)) + ((!sk[23]) & (g78) & (g104) & (!g41) & (g32)) + ((!sk[23]) & (g78) & (g104) & (g41) & (!g32)) + ((!sk[23]) & (g78) & (g104) & (g41) & (g32)) + ((sk[23]) & (!g78) & (!g104) & (!g41) & (!g32)) + ((sk[23]) & (!g78) & (!g104) & (!g41) & (g32)) + ((sk[23]) & (!g78) & (!g104) & (g41) & (!g32)) + ((sk[23]) & (!g78) & (!g104) & (g41) & (g32)) + ((sk[23]) & (!g78) & (g104) & (!g41) & (!g32)));
	assign g270 = (((!g62) & (!g267) & (!g66) & (!g84) & (!g268) & (g269)) + ((!g62) & (!g267) & (g66) & (!g84) & (!g268) & (g269)) + ((g62) & (!g267) & (!g66) & (!g84) & (!g268) & (g269)));
	assign g271 = (((!sk[25]) & (!g71) & (!g25) & (g66)) + ((!sk[25]) & (!g71) & (g25) & (g66)) + ((!sk[25]) & (g71) & (!g25) & (!g66)) + ((!sk[25]) & (g71) & (!g25) & (g66)) + ((!sk[25]) & (g71) & (g25) & (!g66)) + ((!sk[25]) & (g71) & (g25) & (g66)) + ((sk[25]) & (g71) & (!g25) & (g66)) + ((sk[25]) & (g71) & (g25) & (!g66)) + ((sk[25]) & (g71) & (g25) & (g66)));
	assign g272 = (((!ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g66)) + ((!ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g66)) + ((ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g66)) + ((ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g66)));
	assign g273 = (((!g16) & (!sk[27]) & (!g25) & (g19)) + ((!g16) & (!sk[27]) & (g25) & (g19)) + ((!g16) & (sk[27]) & (!g25) & (!g19)) + ((!g16) & (sk[27]) & (g25) & (!g19)) + ((g16) & (!sk[27]) & (!g25) & (!g19)) + ((g16) & (!sk[27]) & (!g25) & (g19)) + ((g16) & (!sk[27]) & (g25) & (!g19)) + ((g16) & (!sk[27]) & (g25) & (g19)) + ((g16) & (sk[27]) & (!g25) & (!g19)));
	assign g274 = (((!sk[28]) & (!g31) & (g13)) + ((!sk[28]) & (g31) & (g13)) + ((sk[28]) & (!g31) & (!g13)));
	assign g275 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (g8) & (g20)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g20)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (g8) & (g20)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (g8) & (g20)));
	assign g276 = (((!g70) & (!g58) & (!g193) & (sk[30]) & (!g275)) + ((!g70) & (!g58) & (g193) & (!sk[30]) & (!g275)) + ((!g70) & (!g58) & (g193) & (!sk[30]) & (g275)) + ((!g70) & (g58) & (!g193) & (sk[30]) & (!g275)) + ((!g70) & (g58) & (g193) & (!sk[30]) & (!g275)) + ((!g70) & (g58) & (g193) & (!sk[30]) & (g275)) + ((g70) & (!g58) & (!g193) & (!sk[30]) & (!g275)) + ((g70) & (!g58) & (!g193) & (!sk[30]) & (g275)) + ((g70) & (!g58) & (!g193) & (sk[30]) & (!g275)) + ((g70) & (!g58) & (g193) & (!sk[30]) & (!g275)) + ((g70) & (!g58) & (g193) & (!sk[30]) & (g275)) + ((g70) & (g58) & (!g193) & (!sk[30]) & (!g275)) + ((g70) & (g58) & (!g193) & (!sk[30]) & (g275)) + ((g70) & (g58) & (g193) & (!sk[30]) & (!g275)) + ((g70) & (g58) & (g193) & (!sk[30]) & (g275)));
	assign g277 = (((!g9) & (!g16) & (!g30) & (!g90) & (!g42) & (!g101)) + ((!g9) & (!g16) & (!g30) & (!g90) & (g42) & (!g101)) + ((!g9) & (!g16) & (g30) & (!g90) & (!g42) & (!g101)) + ((!g9) & (!g16) & (g30) & (!g90) & (g42) & (!g101)) + ((!g9) & (g16) & (!g30) & (!g90) & (!g42) & (!g101)) + ((!g9) & (g16) & (g30) & (!g90) & (!g42) & (!g101)) + ((g9) & (!g16) & (!g30) & (!g90) & (!g42) & (!g101)) + ((g9) & (g16) & (!g30) & (!g90) & (!g42) & (!g101)));
	assign g278 = (((!g70) & (!g99) & (!sk[32]) & (!g30) & (g27) & (!g124)) + ((!g70) & (!g99) & (!sk[32]) & (!g30) & (g27) & (g124)) + ((!g70) & (!g99) & (!sk[32]) & (g30) & (g27) & (!g124)) + ((!g70) & (!g99) & (!sk[32]) & (g30) & (g27) & (g124)) + ((!g70) & (!g99) & (sk[32]) & (!g30) & (!g27) & (!g124)) + ((!g70) & (!g99) & (sk[32]) & (!g30) & (g27) & (!g124)) + ((!g70) & (!g99) & (sk[32]) & (g30) & (!g27) & (!g124)) + ((!g70) & (!g99) & (sk[32]) & (g30) & (g27) & (!g124)) + ((!g70) & (g99) & (!sk[32]) & (!g30) & (!g27) & (!g124)) + ((!g70) & (g99) & (!sk[32]) & (!g30) & (!g27) & (g124)) + ((!g70) & (g99) & (!sk[32]) & (!g30) & (g27) & (!g124)) + ((!g70) & (g99) & (!sk[32]) & (!g30) & (g27) & (g124)) + ((!g70) & (g99) & (!sk[32]) & (g30) & (!g27) & (!g124)) + ((!g70) & (g99) & (!sk[32]) & (g30) & (!g27) & (g124)) + ((!g70) & (g99) & (!sk[32]) & (g30) & (g27) & (!g124)) + ((!g70) & (g99) & (!sk[32]) & (g30) & (g27) & (g124)) + ((!g70) & (g99) & (sk[32]) & (!g30) & (!g27) & (!g124)) + ((!g70) & (g99) & (sk[32]) & (!g30) & (g27) & (!g124)) + ((g70) & (!g99) & (!sk[32]) & (!g30) & (g27) & (!g124)) + ((g70) & (!g99) & (!sk[32]) & (!g30) & (g27) & (g124)) + ((g70) & (!g99) & (!sk[32]) & (g30) & (!g27) & (!g124)) + ((g70) & (!g99) & (!sk[32]) & (g30) & (!g27) & (g124)) + ((g70) & (!g99) & (!sk[32]) & (g30) & (g27) & (!g124)) + ((g70) & (!g99) & (!sk[32]) & (g30) & (g27) & (g124)) + ((g70) & (!g99) & (sk[32]) & (!g30) & (!g27) & (!g124)) + ((g70) & (g99) & (!sk[32]) & (!g30) & (!g27) & (!g124)) + ((g70) & (g99) & (!sk[32]) & (!g30) & (!g27) & (g124)) + ((g70) & (g99) & (!sk[32]) & (!g30) & (g27) & (!g124)) + ((g70) & (g99) & (!sk[32]) & (!g30) & (g27) & (g124)) + ((g70) & (g99) & (!sk[32]) & (g30) & (!g27) & (!g124)) + ((g70) & (g99) & (!sk[32]) & (g30) & (!g27) & (g124)) + ((g70) & (g99) & (!sk[32]) & (g30) & (g27) & (!g124)) + ((g70) & (g99) & (!sk[32]) & (g30) & (g27) & (g124)) + ((g70) & (g99) & (sk[32]) & (!g30) & (!g27) & (!g124)));
	assign g279 = (((!g272) & (g273) & (g274) & (g276) & (g277) & (g278)));
	assign g280 = (((!g259) & (!g266) & (!g270) & (g271) & (!sk[34]) & (!g279)) + ((!g259) & (!g266) & (!g270) & (g271) & (!sk[34]) & (g279)) + ((!g259) & (!g266) & (g270) & (g271) & (!sk[34]) & (!g279)) + ((!g259) & (!g266) & (g270) & (g271) & (!sk[34]) & (g279)) + ((!g259) & (g266) & (!g270) & (!g271) & (!sk[34]) & (!g279)) + ((!g259) & (g266) & (!g270) & (!g271) & (!sk[34]) & (g279)) + ((!g259) & (g266) & (!g270) & (g271) & (!sk[34]) & (!g279)) + ((!g259) & (g266) & (!g270) & (g271) & (!sk[34]) & (g279)) + ((!g259) & (g266) & (g270) & (!g271) & (!sk[34]) & (!g279)) + ((!g259) & (g266) & (g270) & (!g271) & (!sk[34]) & (g279)) + ((!g259) & (g266) & (g270) & (g271) & (!sk[34]) & (!g279)) + ((!g259) & (g266) & (g270) & (g271) & (!sk[34]) & (g279)) + ((g259) & (!g266) & (!g270) & (g271) & (!sk[34]) & (!g279)) + ((g259) & (!g266) & (!g270) & (g271) & (!sk[34]) & (g279)) + ((g259) & (!g266) & (g270) & (!g271) & (!sk[34]) & (!g279)) + ((g259) & (!g266) & (g270) & (!g271) & (!sk[34]) & (g279)) + ((g259) & (!g266) & (g270) & (g271) & (!sk[34]) & (!g279)) + ((g259) & (!g266) & (g270) & (g271) & (!sk[34]) & (g279)) + ((g259) & (g266) & (!g270) & (!g271) & (!sk[34]) & (!g279)) + ((g259) & (g266) & (!g270) & (!g271) & (!sk[34]) & (g279)) + ((g259) & (g266) & (!g270) & (g271) & (!sk[34]) & (!g279)) + ((g259) & (g266) & (!g270) & (g271) & (!sk[34]) & (g279)) + ((g259) & (g266) & (g270) & (!g271) & (!sk[34]) & (!g279)) + ((g259) & (g266) & (g270) & (!g271) & (!sk[34]) & (g279)) + ((g259) & (g266) & (g270) & (!g271) & (sk[34]) & (g279)) + ((g259) & (g266) & (g270) & (g271) & (!sk[34]) & (!g279)) + ((g259) & (g266) & (g270) & (g271) & (!sk[34]) & (g279)));
	assign g281 = (((!g251) & (!sk[35]) & (!g252) & (!g253) & (g122) & (!g280)) + ((!g251) & (!sk[35]) & (!g252) & (!g253) & (g122) & (g280)) + ((!g251) & (!sk[35]) & (!g252) & (g253) & (g122) & (!g280)) + ((!g251) & (!sk[35]) & (!g252) & (g253) & (g122) & (g280)) + ((!g251) & (!sk[35]) & (g252) & (!g253) & (!g122) & (!g280)) + ((!g251) & (!sk[35]) & (g252) & (!g253) & (!g122) & (g280)) + ((!g251) & (!sk[35]) & (g252) & (!g253) & (g122) & (!g280)) + ((!g251) & (!sk[35]) & (g252) & (!g253) & (g122) & (g280)) + ((!g251) & (!sk[35]) & (g252) & (g253) & (!g122) & (!g280)) + ((!g251) & (!sk[35]) & (g252) & (g253) & (!g122) & (g280)) + ((!g251) & (!sk[35]) & (g252) & (g253) & (g122) & (!g280)) + ((!g251) & (!sk[35]) & (g252) & (g253) & (g122) & (g280)) + ((!g251) & (sk[35]) & (!g252) & (!g253) & (!g122) & (g280)) + ((!g251) & (sk[35]) & (!g252) & (!g253) & (g122) & (!g280)) + ((!g251) & (sk[35]) & (!g252) & (!g253) & (g122) & (g280)) + ((!g251) & (sk[35]) & (!g252) & (g253) & (!g122) & (g280)) + ((!g251) & (sk[35]) & (!g252) & (g253) & (g122) & (!g280)) + ((!g251) & (sk[35]) & (g252) & (!g253) & (g122) & (g280)) + ((g251) & (!sk[35]) & (!g252) & (!g253) & (g122) & (!g280)) + ((g251) & (!sk[35]) & (!g252) & (!g253) & (g122) & (g280)) + ((g251) & (!sk[35]) & (!g252) & (g253) & (!g122) & (!g280)) + ((g251) & (!sk[35]) & (!g252) & (g253) & (!g122) & (g280)) + ((g251) & (!sk[35]) & (!g252) & (g253) & (g122) & (!g280)) + ((g251) & (!sk[35]) & (!g252) & (g253) & (g122) & (g280)) + ((g251) & (!sk[35]) & (g252) & (!g253) & (!g122) & (!g280)) + ((g251) & (!sk[35]) & (g252) & (!g253) & (!g122) & (g280)) + ((g251) & (!sk[35]) & (g252) & (!g253) & (g122) & (!g280)) + ((g251) & (!sk[35]) & (g252) & (!g253) & (g122) & (g280)) + ((g251) & (!sk[35]) & (g252) & (g253) & (!g122) & (!g280)) + ((g251) & (!sk[35]) & (g252) & (g253) & (!g122) & (g280)) + ((g251) & (!sk[35]) & (g252) & (g253) & (g122) & (!g280)) + ((g251) & (!sk[35]) & (g252) & (g253) & (g122) & (g280)) + ((g251) & (sk[35]) & (!g252) & (g253) & (!g122) & (!g280)) + ((g251) & (sk[35]) & (g252) & (!g253) & (!g122) & (g280)) + ((g251) & (sk[35]) & (g252) & (!g253) & (g122) & (!g280)) + ((g251) & (sk[35]) & (g252) & (g253) & (!g122) & (!g280)) + ((g251) & (sk[35]) & (g252) & (g253) & (!g122) & (g280)) + ((g251) & (sk[35]) & (g252) & (g253) & (g122) & (!g280)));
	assign g282 = (((!g70) & (!g10) & (!sk[36]) & (!g42) & (g50) & (!g33)) + ((!g70) & (!g10) & (!sk[36]) & (!g42) & (g50) & (g33)) + ((!g70) & (!g10) & (!sk[36]) & (g42) & (g50) & (!g33)) + ((!g70) & (!g10) & (!sk[36]) & (g42) & (g50) & (g33)) + ((!g70) & (!g10) & (sk[36]) & (!g42) & (!g50) & (!g33)) + ((!g70) & (!g10) & (sk[36]) & (g42) & (!g50) & (!g33)) + ((!g70) & (g10) & (!sk[36]) & (!g42) & (!g50) & (!g33)) + ((!g70) & (g10) & (!sk[36]) & (!g42) & (!g50) & (g33)) + ((!g70) & (g10) & (!sk[36]) & (!g42) & (g50) & (!g33)) + ((!g70) & (g10) & (!sk[36]) & (!g42) & (g50) & (g33)) + ((!g70) & (g10) & (!sk[36]) & (g42) & (!g50) & (!g33)) + ((!g70) & (g10) & (!sk[36]) & (g42) & (!g50) & (g33)) + ((!g70) & (g10) & (!sk[36]) & (g42) & (g50) & (!g33)) + ((!g70) & (g10) & (!sk[36]) & (g42) & (g50) & (g33)) + ((!g70) & (g10) & (sk[36]) & (!g42) & (!g50) & (!g33)) + ((!g70) & (g10) & (sk[36]) & (g42) & (!g50) & (!g33)) + ((g70) & (!g10) & (!sk[36]) & (!g42) & (g50) & (!g33)) + ((g70) & (!g10) & (!sk[36]) & (!g42) & (g50) & (g33)) + ((g70) & (!g10) & (!sk[36]) & (g42) & (!g50) & (!g33)) + ((g70) & (!g10) & (!sk[36]) & (g42) & (!g50) & (g33)) + ((g70) & (!g10) & (!sk[36]) & (g42) & (g50) & (!g33)) + ((g70) & (!g10) & (!sk[36]) & (g42) & (g50) & (g33)) + ((g70) & (!g10) & (sk[36]) & (!g42) & (!g50) & (!g33)) + ((g70) & (g10) & (!sk[36]) & (!g42) & (!g50) & (!g33)) + ((g70) & (g10) & (!sk[36]) & (!g42) & (!g50) & (g33)) + ((g70) & (g10) & (!sk[36]) & (!g42) & (g50) & (!g33)) + ((g70) & (g10) & (!sk[36]) & (!g42) & (g50) & (g33)) + ((g70) & (g10) & (!sk[36]) & (g42) & (!g50) & (!g33)) + ((g70) & (g10) & (!sk[36]) & (g42) & (!g50) & (g33)) + ((g70) & (g10) & (!sk[36]) & (g42) & (g50) & (!g33)) + ((g70) & (g10) & (!sk[36]) & (g42) & (g50) & (g33)));
	assign g283 = (((!g9) & (!g30) & (!g87) & (!g131) & (g123) & (g282)) + ((!g9) & (g30) & (!g87) & (!g131) & (g123) & (g282)) + ((g9) & (!g30) & (!g87) & (!g131) & (g123) & (g282)));
	assign g284 = (((!g38) & (!sk[38]) & (!g16) & (g12) & (!g104)) + ((!g38) & (!sk[38]) & (!g16) & (g12) & (g104)) + ((!g38) & (!sk[38]) & (g16) & (g12) & (!g104)) + ((!g38) & (!sk[38]) & (g16) & (g12) & (g104)) + ((!g38) & (sk[38]) & (g16) & (g12) & (!g104)) + ((!g38) & (sk[38]) & (g16) & (g12) & (g104)) + ((g38) & (!sk[38]) & (!g16) & (!g12) & (!g104)) + ((g38) & (!sk[38]) & (!g16) & (!g12) & (g104)) + ((g38) & (!sk[38]) & (!g16) & (g12) & (!g104)) + ((g38) & (!sk[38]) & (!g16) & (g12) & (g104)) + ((g38) & (!sk[38]) & (g16) & (!g12) & (!g104)) + ((g38) & (!sk[38]) & (g16) & (!g12) & (g104)) + ((g38) & (!sk[38]) & (g16) & (g12) & (!g104)) + ((g38) & (!sk[38]) & (g16) & (g12) & (g104)) + ((g38) & (sk[38]) & (!g16) & (!g12) & (g104)) + ((g38) & (sk[38]) & (!g16) & (g12) & (g104)) + ((g38) & (sk[38]) & (g16) & (!g12) & (g104)) + ((g38) & (sk[38]) & (g16) & (g12) & (!g104)) + ((g38) & (sk[38]) & (g16) & (g12) & (g104)));
	assign g285 = (((!g114) & (!g115) & (!g8) & (g10) & (!g12) & (!g18)) + ((!g114) & (!g115) & (!g8) & (g10) & (!g12) & (g18)) + ((!g114) & (!g115) & (!g8) & (g10) & (g12) & (!g18)) + ((!g114) & (!g115) & (!g8) & (g10) & (g12) & (g18)) + ((!g114) & (!g115) & (g8) & (!g10) & (!g12) & (g18)) + ((!g114) & (!g115) & (g8) & (!g10) & (g12) & (g18)) + ((!g114) & (!g115) & (g8) & (g10) & (!g12) & (g18)) + ((!g114) & (!g115) & (g8) & (g10) & (g12) & (g18)) + ((!g114) & (g115) & (!g8) & (g10) & (!g12) & (!g18)) + ((!g114) & (g115) & (!g8) & (g10) & (!g12) & (g18)) + ((!g114) & (g115) & (!g8) & (g10) & (g12) & (!g18)) + ((!g114) & (g115) & (!g8) & (g10) & (g12) & (g18)) + ((g114) & (g115) & (!g8) & (!g10) & (g12) & (!g18)) + ((g114) & (g115) & (!g8) & (!g10) & (g12) & (g18)) + ((g114) & (g115) & (!g8) & (g10) & (!g12) & (!g18)) + ((g114) & (g115) & (!g8) & (g10) & (!g12) & (g18)) + ((g114) & (g115) & (!g8) & (g10) & (g12) & (!g18)) + ((g114) & (g115) & (!g8) & (g10) & (g12) & (g18)));
	assign g286 = (((!g71) & (!g20) & (!g284) & (g130) & (!sk[40]) & (!g285)) + ((!g71) & (!g20) & (!g284) & (g130) & (!sk[40]) & (g285)) + ((!g71) & (!g20) & (!g284) & (g130) & (sk[40]) & (!g285)) + ((!g71) & (!g20) & (g284) & (g130) & (!sk[40]) & (!g285)) + ((!g71) & (!g20) & (g284) & (g130) & (!sk[40]) & (g285)) + ((!g71) & (g20) & (!g284) & (!g130) & (!sk[40]) & (!g285)) + ((!g71) & (g20) & (!g284) & (!g130) & (!sk[40]) & (g285)) + ((!g71) & (g20) & (!g284) & (g130) & (!sk[40]) & (!g285)) + ((!g71) & (g20) & (!g284) & (g130) & (!sk[40]) & (g285)) + ((!g71) & (g20) & (!g284) & (g130) & (sk[40]) & (!g285)) + ((!g71) & (g20) & (g284) & (!g130) & (!sk[40]) & (!g285)) + ((!g71) & (g20) & (g284) & (!g130) & (!sk[40]) & (g285)) + ((!g71) & (g20) & (g284) & (g130) & (!sk[40]) & (!g285)) + ((!g71) & (g20) & (g284) & (g130) & (!sk[40]) & (g285)) + ((g71) & (!g20) & (!g284) & (g130) & (!sk[40]) & (!g285)) + ((g71) & (!g20) & (!g284) & (g130) & (!sk[40]) & (g285)) + ((g71) & (!g20) & (!g284) & (g130) & (sk[40]) & (!g285)) + ((g71) & (!g20) & (g284) & (!g130) & (!sk[40]) & (!g285)) + ((g71) & (!g20) & (g284) & (!g130) & (!sk[40]) & (g285)) + ((g71) & (!g20) & (g284) & (g130) & (!sk[40]) & (!g285)) + ((g71) & (!g20) & (g284) & (g130) & (!sk[40]) & (g285)) + ((g71) & (g20) & (!g284) & (!g130) & (!sk[40]) & (!g285)) + ((g71) & (g20) & (!g284) & (!g130) & (!sk[40]) & (g285)) + ((g71) & (g20) & (!g284) & (g130) & (!sk[40]) & (!g285)) + ((g71) & (g20) & (!g284) & (g130) & (!sk[40]) & (g285)) + ((g71) & (g20) & (g284) & (!g130) & (!sk[40]) & (!g285)) + ((g71) & (g20) & (g284) & (!g130) & (!sk[40]) & (g285)) + ((g71) & (g20) & (g284) & (g130) & (!sk[40]) & (!g285)) + ((g71) & (g20) & (g284) & (g130) & (!sk[40]) & (g285)));
	assign g287 = (((!g9) & (!sk[41]) & (!g99) & (g41) & (!g20)) + ((!g9) & (!sk[41]) & (!g99) & (g41) & (g20)) + ((!g9) & (!sk[41]) & (g99) & (g41) & (!g20)) + ((!g9) & (!sk[41]) & (g99) & (g41) & (g20)) + ((!g9) & (sk[41]) & (g99) & (!g41) & (g20)) + ((!g9) & (sk[41]) & (g99) & (g41) & (g20)) + ((g9) & (!sk[41]) & (!g99) & (!g41) & (!g20)) + ((g9) & (!sk[41]) & (!g99) & (!g41) & (g20)) + ((g9) & (!sk[41]) & (!g99) & (g41) & (!g20)) + ((g9) & (!sk[41]) & (!g99) & (g41) & (g20)) + ((g9) & (!sk[41]) & (g99) & (!g41) & (!g20)) + ((g9) & (!sk[41]) & (g99) & (!g41) & (g20)) + ((g9) & (!sk[41]) & (g99) & (g41) & (!g20)) + ((g9) & (!sk[41]) & (g99) & (g41) & (g20)) + ((g9) & (sk[41]) & (!g99) & (!g41) & (g20)) + ((g9) & (sk[41]) & (!g99) & (g41) & (!g20)) + ((g9) & (sk[41]) & (!g99) & (g41) & (g20)) + ((g9) & (sk[41]) & (g99) & (!g41) & (g20)) + ((g9) & (sk[41]) & (g99) & (g41) & (!g20)) + ((g9) & (sk[41]) & (g99) & (g41) & (g20)));
	assign g288 = (((!ax22x) & (!ax21x) & (!g6) & (ax20x) & (!g8) & (g27)) + ((!ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g27)) + ((ax22x) & (ax21x) & (!g6) & (!ax20x) & (!g8) & (g27)) + ((ax22x) & (ax21x) & (g6) & (!ax20x) & (!g8) & (g27)));
	assign g289 = (((!g70) & (!sk[43]) & (!g163) & (g25) & (!g288)) + ((!g70) & (!sk[43]) & (!g163) & (g25) & (g288)) + ((!g70) & (!sk[43]) & (g163) & (g25) & (!g288)) + ((!g70) & (!sk[43]) & (g163) & (g25) & (g288)) + ((!g70) & (sk[43]) & (!g163) & (!g25) & (!g288)) + ((!g70) & (sk[43]) & (!g163) & (g25) & (!g288)) + ((g70) & (!sk[43]) & (!g163) & (!g25) & (!g288)) + ((g70) & (!sk[43]) & (!g163) & (!g25) & (g288)) + ((g70) & (!sk[43]) & (!g163) & (g25) & (!g288)) + ((g70) & (!sk[43]) & (!g163) & (g25) & (g288)) + ((g70) & (!sk[43]) & (g163) & (!g25) & (!g288)) + ((g70) & (!sk[43]) & (g163) & (!g25) & (g288)) + ((g70) & (!sk[43]) & (g163) & (g25) & (!g288)) + ((g70) & (!sk[43]) & (g163) & (g25) & (g288)) + ((g70) & (sk[43]) & (!g163) & (!g25) & (!g288)));
	assign g290 = (((!g16) & (!g238) & (!sk[44]) & (g40)) + ((!g16) & (!g238) & (sk[44]) & (!g40)) + ((!g16) & (!g238) & (sk[44]) & (g40)) + ((!g16) & (g238) & (!sk[44]) & (g40)) + ((g16) & (!g238) & (!sk[44]) & (!g40)) + ((g16) & (!g238) & (!sk[44]) & (g40)) + ((g16) & (!g238) & (sk[44]) & (!g40)) + ((g16) & (g238) & (!sk[44]) & (!g40)) + ((g16) & (g238) & (!sk[44]) & (g40)));
	assign g291 = (((!g59) & (!g84) & (!sk[45]) & (g137)) + ((!g59) & (!g84) & (sk[45]) & (!g137)) + ((!g59) & (g84) & (!sk[45]) & (g137)) + ((g59) & (!g84) & (!sk[45]) & (!g137)) + ((g59) & (!g84) & (!sk[45]) & (g137)) + ((g59) & (g84) & (!sk[45]) & (!g137)) + ((g59) & (g84) & (!sk[45]) & (g137)));
	assign g292 = (((!sk[46]) & (!g114) & (!g115) & (!g8) & (g18) & (!g42)) + ((!sk[46]) & (!g114) & (!g115) & (!g8) & (g18) & (g42)) + ((!sk[46]) & (!g114) & (!g115) & (g8) & (g18) & (!g42)) + ((!sk[46]) & (!g114) & (!g115) & (g8) & (g18) & (g42)) + ((!sk[46]) & (!g114) & (g115) & (!g8) & (!g18) & (!g42)) + ((!sk[46]) & (!g114) & (g115) & (!g8) & (!g18) & (g42)) + ((!sk[46]) & (!g114) & (g115) & (!g8) & (g18) & (!g42)) + ((!sk[46]) & (!g114) & (g115) & (!g8) & (g18) & (g42)) + ((!sk[46]) & (!g114) & (g115) & (g8) & (!g18) & (!g42)) + ((!sk[46]) & (!g114) & (g115) & (g8) & (!g18) & (g42)) + ((!sk[46]) & (!g114) & (g115) & (g8) & (g18) & (!g42)) + ((!sk[46]) & (!g114) & (g115) & (g8) & (g18) & (g42)) + ((!sk[46]) & (g114) & (!g115) & (!g8) & (g18) & (!g42)) + ((!sk[46]) & (g114) & (!g115) & (!g8) & (g18) & (g42)) + ((!sk[46]) & (g114) & (!g115) & (g8) & (!g18) & (!g42)) + ((!sk[46]) & (g114) & (!g115) & (g8) & (!g18) & (g42)) + ((!sk[46]) & (g114) & (!g115) & (g8) & (g18) & (!g42)) + ((!sk[46]) & (g114) & (!g115) & (g8) & (g18) & (g42)) + ((!sk[46]) & (g114) & (g115) & (!g8) & (!g18) & (!g42)) + ((!sk[46]) & (g114) & (g115) & (!g8) & (!g18) & (g42)) + ((!sk[46]) & (g114) & (g115) & (!g8) & (g18) & (!g42)) + ((!sk[46]) & (g114) & (g115) & (!g8) & (g18) & (g42)) + ((!sk[46]) & (g114) & (g115) & (g8) & (!g18) & (!g42)) + ((!sk[46]) & (g114) & (g115) & (g8) & (!g18) & (g42)) + ((!sk[46]) & (g114) & (g115) & (g8) & (g18) & (!g42)) + ((!sk[46]) & (g114) & (g115) & (g8) & (g18) & (g42)) + ((sk[46]) & (!g114) & (!g115) & (!g8) & (g18) & (!g42)) + ((sk[46]) & (!g114) & (!g115) & (!g8) & (g18) & (g42)) + ((sk[46]) & (g114) & (!g115) & (g8) & (g18) & (!g42)) + ((sk[46]) & (g114) & (!g115) & (g8) & (g18) & (g42)) + ((sk[46]) & (g114) & (g115) & (g8) & (!g18) & (g42)) + ((sk[46]) & (g114) & (g115) & (g8) & (g18) & (g42)));
	assign g293 = (((!g287) & (!sk[47]) & (!g289) & (!g290) & (g291) & (!g292)) + ((!g287) & (!sk[47]) & (!g289) & (!g290) & (g291) & (g292)) + ((!g287) & (!sk[47]) & (!g289) & (g290) & (g291) & (!g292)) + ((!g287) & (!sk[47]) & (!g289) & (g290) & (g291) & (g292)) + ((!g287) & (!sk[47]) & (g289) & (!g290) & (!g291) & (!g292)) + ((!g287) & (!sk[47]) & (g289) & (!g290) & (!g291) & (g292)) + ((!g287) & (!sk[47]) & (g289) & (!g290) & (g291) & (!g292)) + ((!g287) & (!sk[47]) & (g289) & (!g290) & (g291) & (g292)) + ((!g287) & (!sk[47]) & (g289) & (g290) & (!g291) & (!g292)) + ((!g287) & (!sk[47]) & (g289) & (g290) & (!g291) & (g292)) + ((!g287) & (!sk[47]) & (g289) & (g290) & (g291) & (!g292)) + ((!g287) & (!sk[47]) & (g289) & (g290) & (g291) & (g292)) + ((!g287) & (sk[47]) & (g289) & (g290) & (g291) & (!g292)) + ((g287) & (!sk[47]) & (!g289) & (!g290) & (g291) & (!g292)) + ((g287) & (!sk[47]) & (!g289) & (!g290) & (g291) & (g292)) + ((g287) & (!sk[47]) & (!g289) & (g290) & (!g291) & (!g292)) + ((g287) & (!sk[47]) & (!g289) & (g290) & (!g291) & (g292)) + ((g287) & (!sk[47]) & (!g289) & (g290) & (g291) & (!g292)) + ((g287) & (!sk[47]) & (!g289) & (g290) & (g291) & (g292)) + ((g287) & (!sk[47]) & (g289) & (!g290) & (!g291) & (!g292)) + ((g287) & (!sk[47]) & (g289) & (!g290) & (!g291) & (g292)) + ((g287) & (!sk[47]) & (g289) & (!g290) & (g291) & (!g292)) + ((g287) & (!sk[47]) & (g289) & (!g290) & (g291) & (g292)) + ((g287) & (!sk[47]) & (g289) & (g290) & (!g291) & (!g292)) + ((g287) & (!sk[47]) & (g289) & (g290) & (!g291) & (g292)) + ((g287) & (!sk[47]) & (g289) & (g290) & (g291) & (!g292)) + ((g287) & (!sk[47]) & (g289) & (g290) & (g291) & (g292)));
	assign g294 = (((!g9) & (!g62) & (!g40) & (!g66) & (sk[48]) & (!g171)) + ((!g9) & (!g62) & (!g40) & (g66) & (!sk[48]) & (!g171)) + ((!g9) & (!g62) & (!g40) & (g66) & (!sk[48]) & (g171)) + ((!g9) & (!g62) & (!g40) & (g66) & (sk[48]) & (!g171)) + ((!g9) & (!g62) & (g40) & (!g66) & (sk[48]) & (!g171)) + ((!g9) & (!g62) & (g40) & (g66) & (!sk[48]) & (!g171)) + ((!g9) & (!g62) & (g40) & (g66) & (!sk[48]) & (g171)) + ((!g9) & (!g62) & (g40) & (g66) & (sk[48]) & (!g171)) + ((!g9) & (g62) & (!g40) & (!g66) & (!sk[48]) & (!g171)) + ((!g9) & (g62) & (!g40) & (!g66) & (!sk[48]) & (g171)) + ((!g9) & (g62) & (!g40) & (!g66) & (sk[48]) & (!g171)) + ((!g9) & (g62) & (!g40) & (g66) & (!sk[48]) & (!g171)) + ((!g9) & (g62) & (!g40) & (g66) & (!sk[48]) & (g171)) + ((!g9) & (g62) & (g40) & (!g66) & (!sk[48]) & (!g171)) + ((!g9) & (g62) & (g40) & (!g66) & (!sk[48]) & (g171)) + ((!g9) & (g62) & (g40) & (!g66) & (sk[48]) & (!g171)) + ((!g9) & (g62) & (g40) & (g66) & (!sk[48]) & (!g171)) + ((!g9) & (g62) & (g40) & (g66) & (!sk[48]) & (g171)) + ((g9) & (!g62) & (!g40) & (!g66) & (sk[48]) & (!g171)) + ((g9) & (!g62) & (!g40) & (g66) & (!sk[48]) & (!g171)) + ((g9) & (!g62) & (!g40) & (g66) & (!sk[48]) & (g171)) + ((g9) & (!g62) & (!g40) & (g66) & (sk[48]) & (!g171)) + ((g9) & (!g62) & (g40) & (!g66) & (!sk[48]) & (!g171)) + ((g9) & (!g62) & (g40) & (!g66) & (!sk[48]) & (g171)) + ((g9) & (!g62) & (g40) & (g66) & (!sk[48]) & (!g171)) + ((g9) & (!g62) & (g40) & (g66) & (!sk[48]) & (g171)) + ((g9) & (g62) & (!g40) & (!g66) & (!sk[48]) & (!g171)) + ((g9) & (g62) & (!g40) & (!g66) & (!sk[48]) & (g171)) + ((g9) & (g62) & (!g40) & (!g66) & (sk[48]) & (!g171)) + ((g9) & (g62) & (!g40) & (g66) & (!sk[48]) & (!g171)) + ((g9) & (g62) & (!g40) & (g66) & (!sk[48]) & (g171)) + ((g9) & (g62) & (g40) & (!g66) & (!sk[48]) & (!g171)) + ((g9) & (g62) & (g40) & (!g66) & (!sk[48]) & (g171)) + ((g9) & (g62) & (g40) & (g66) & (!sk[48]) & (!g171)) + ((g9) & (g62) & (g40) & (g66) & (!sk[48]) & (g171)));
	assign g295 = (((!g16) & (!g25) & (!g241) & (!g152) & (!g161) & (g294)) + ((!g16) & (g25) & (!g241) & (!g152) & (!g161) & (g294)) + ((g16) & (!g25) & (!g241) & (!g152) & (!g161) & (g294)));
	assign g296 = (((!g83) & (!g29) & (!g60) & (sk[50]) & (!g154)) + ((!g83) & (!g29) & (g60) & (!sk[50]) & (!g154)) + ((!g83) & (!g29) & (g60) & (!sk[50]) & (g154)) + ((!g83) & (g29) & (g60) & (!sk[50]) & (!g154)) + ((!g83) & (g29) & (g60) & (!sk[50]) & (g154)) + ((g83) & (!g29) & (!g60) & (!sk[50]) & (!g154)) + ((g83) & (!g29) & (!g60) & (!sk[50]) & (g154)) + ((g83) & (!g29) & (g60) & (!sk[50]) & (!g154)) + ((g83) & (!g29) & (g60) & (!sk[50]) & (g154)) + ((g83) & (g29) & (!g60) & (!sk[50]) & (!g154)) + ((g83) & (g29) & (!g60) & (!sk[50]) & (g154)) + ((g83) & (g29) & (g60) & (!sk[50]) & (!g154)) + ((g83) & (g29) & (g60) & (!sk[50]) & (g154)));
	assign g297 = (((!g49) & (!sk[51]) & (!g62) & (g71) & (!g27)) + ((!g49) & (!sk[51]) & (!g62) & (g71) & (g27)) + ((!g49) & (!sk[51]) & (g62) & (g71) & (!g27)) + ((!g49) & (!sk[51]) & (g62) & (g71) & (g27)) + ((!g49) & (sk[51]) & (g62) & (!g71) & (g27)) + ((!g49) & (sk[51]) & (g62) & (g71) & (g27)) + ((g49) & (!sk[51]) & (!g62) & (!g71) & (!g27)) + ((g49) & (!sk[51]) & (!g62) & (!g71) & (g27)) + ((g49) & (!sk[51]) & (!g62) & (g71) & (!g27)) + ((g49) & (!sk[51]) & (!g62) & (g71) & (g27)) + ((g49) & (!sk[51]) & (g62) & (!g71) & (!g27)) + ((g49) & (!sk[51]) & (g62) & (!g71) & (g27)) + ((g49) & (!sk[51]) & (g62) & (g71) & (!g27)) + ((g49) & (!sk[51]) & (g62) & (g71) & (g27)) + ((g49) & (sk[51]) & (!g62) & (g71) & (!g27)) + ((g49) & (sk[51]) & (!g62) & (g71) & (g27)) + ((g49) & (sk[51]) & (g62) & (!g71) & (g27)) + ((g49) & (sk[51]) & (g62) & (g71) & (!g27)) + ((g49) & (sk[51]) & (g62) & (g71) & (g27)));
	assign g298 = (((!g70) & (!g30) & (!g79) & (!g46) & (sk[52]) & (!g40)) + ((!g70) & (!g30) & (!g79) & (!g46) & (sk[52]) & (g40)) + ((!g70) & (!g30) & (!g79) & (g46) & (!sk[52]) & (!g40)) + ((!g70) & (!g30) & (!g79) & (g46) & (!sk[52]) & (g40)) + ((!g70) & (!g30) & (!g79) & (g46) & (sk[52]) & (!g40)) + ((!g70) & (!g30) & (g79) & (g46) & (!sk[52]) & (!g40)) + ((!g70) & (!g30) & (g79) & (g46) & (!sk[52]) & (g40)) + ((!g70) & (g30) & (!g79) & (!g46) & (!sk[52]) & (!g40)) + ((!g70) & (g30) & (!g79) & (!g46) & (!sk[52]) & (g40)) + ((!g70) & (g30) & (!g79) & (!g46) & (sk[52]) & (!g40)) + ((!g70) & (g30) & (!g79) & (!g46) & (sk[52]) & (g40)) + ((!g70) & (g30) & (!g79) & (g46) & (!sk[52]) & (!g40)) + ((!g70) & (g30) & (!g79) & (g46) & (!sk[52]) & (g40)) + ((!g70) & (g30) & (!g79) & (g46) & (sk[52]) & (!g40)) + ((!g70) & (g30) & (g79) & (!g46) & (!sk[52]) & (!g40)) + ((!g70) & (g30) & (g79) & (!g46) & (!sk[52]) & (g40)) + ((!g70) & (g30) & (g79) & (g46) & (!sk[52]) & (!g40)) + ((!g70) & (g30) & (g79) & (g46) & (!sk[52]) & (g40)) + ((g70) & (!g30) & (!g79) & (!g46) & (sk[52]) & (!g40)) + ((g70) & (!g30) & (!g79) & (!g46) & (sk[52]) & (g40)) + ((g70) & (!g30) & (!g79) & (g46) & (!sk[52]) & (!g40)) + ((g70) & (!g30) & (!g79) & (g46) & (!sk[52]) & (g40)) + ((g70) & (!g30) & (!g79) & (g46) & (sk[52]) & (!g40)) + ((g70) & (!g30) & (g79) & (!g46) & (!sk[52]) & (!g40)) + ((g70) & (!g30) & (g79) & (!g46) & (!sk[52]) & (g40)) + ((g70) & (!g30) & (g79) & (g46) & (!sk[52]) & (!g40)) + ((g70) & (!g30) & (g79) & (g46) & (!sk[52]) & (g40)) + ((g70) & (g30) & (!g79) & (!g46) & (!sk[52]) & (!g40)) + ((g70) & (g30) & (!g79) & (!g46) & (!sk[52]) & (g40)) + ((g70) & (g30) & (!g79) & (g46) & (!sk[52]) & (!g40)) + ((g70) & (g30) & (!g79) & (g46) & (!sk[52]) & (g40)) + ((g70) & (g30) & (g79) & (!g46) & (!sk[52]) & (!g40)) + ((g70) & (g30) & (g79) & (!g46) & (!sk[52]) & (g40)) + ((g70) & (g30) & (g79) & (g46) & (!sk[52]) & (!g40)) + ((g70) & (g30) & (g79) & (g46) & (!sk[52]) & (g40)));
	assign g299 = (((!g9) & (!sk[53]) & (!g62) & (!g25) & (g41) & (!g86)) + ((!g9) & (!sk[53]) & (!g62) & (!g25) & (g41) & (g86)) + ((!g9) & (!sk[53]) & (!g62) & (g25) & (g41) & (!g86)) + ((!g9) & (!sk[53]) & (!g62) & (g25) & (g41) & (g86)) + ((!g9) & (!sk[53]) & (g62) & (!g25) & (!g41) & (!g86)) + ((!g9) & (!sk[53]) & (g62) & (!g25) & (!g41) & (g86)) + ((!g9) & (!sk[53]) & (g62) & (!g25) & (g41) & (!g86)) + ((!g9) & (!sk[53]) & (g62) & (!g25) & (g41) & (g86)) + ((!g9) & (!sk[53]) & (g62) & (g25) & (!g41) & (!g86)) + ((!g9) & (!sk[53]) & (g62) & (g25) & (!g41) & (g86)) + ((!g9) & (!sk[53]) & (g62) & (g25) & (g41) & (!g86)) + ((!g9) & (!sk[53]) & (g62) & (g25) & (g41) & (g86)) + ((!g9) & (sk[53]) & (!g62) & (!g25) & (!g41) & (!g86)) + ((!g9) & (sk[53]) & (!g62) & (!g25) & (g41) & (!g86)) + ((!g9) & (sk[53]) & (!g62) & (g25) & (!g41) & (!g86)) + ((!g9) & (sk[53]) & (!g62) & (g25) & (g41) & (!g86)) + ((!g9) & (sk[53]) & (g62) & (!g25) & (!g41) & (!g86)) + ((!g9) & (sk[53]) & (g62) & (g25) & (!g41) & (!g86)) + ((g9) & (!sk[53]) & (!g62) & (!g25) & (g41) & (!g86)) + ((g9) & (!sk[53]) & (!g62) & (!g25) & (g41) & (g86)) + ((g9) & (!sk[53]) & (!g62) & (g25) & (!g41) & (!g86)) + ((g9) & (!sk[53]) & (!g62) & (g25) & (!g41) & (g86)) + ((g9) & (!sk[53]) & (!g62) & (g25) & (g41) & (!g86)) + ((g9) & (!sk[53]) & (!g62) & (g25) & (g41) & (g86)) + ((g9) & (!sk[53]) & (g62) & (!g25) & (!g41) & (!g86)) + ((g9) & (!sk[53]) & (g62) & (!g25) & (!g41) & (g86)) + ((g9) & (!sk[53]) & (g62) & (!g25) & (g41) & (!g86)) + ((g9) & (!sk[53]) & (g62) & (!g25) & (g41) & (g86)) + ((g9) & (!sk[53]) & (g62) & (g25) & (!g41) & (!g86)) + ((g9) & (!sk[53]) & (g62) & (g25) & (!g41) & (g86)) + ((g9) & (!sk[53]) & (g62) & (g25) & (g41) & (!g86)) + ((g9) & (!sk[53]) & (g62) & (g25) & (g41) & (g86)) + ((g9) & (sk[53]) & (!g62) & (!g25) & (!g41) & (!g86)) + ((g9) & (sk[53]) & (!g62) & (!g25) & (g41) & (!g86)) + ((g9) & (sk[53]) & (g62) & (!g25) & (!g41) & (!g86)));
	assign g300 = (((!g296) & (!g297) & (g298) & (!sk[54]) & (!g299)) + ((!g296) & (!g297) & (g298) & (!sk[54]) & (g299)) + ((!g296) & (g297) & (g298) & (!sk[54]) & (!g299)) + ((!g296) & (g297) & (g298) & (!sk[54]) & (g299)) + ((g296) & (!g297) & (!g298) & (!sk[54]) & (!g299)) + ((g296) & (!g297) & (!g298) & (!sk[54]) & (g299)) + ((g296) & (!g297) & (g298) & (!sk[54]) & (!g299)) + ((g296) & (!g297) & (g298) & (!sk[54]) & (g299)) + ((g296) & (!g297) & (g298) & (sk[54]) & (g299)) + ((g296) & (g297) & (!g298) & (!sk[54]) & (!g299)) + ((g296) & (g297) & (!g298) & (!sk[54]) & (g299)) + ((g296) & (g297) & (g298) & (!sk[54]) & (!g299)) + ((g296) & (g297) & (g298) & (!sk[54]) & (g299)));
	assign g301 = (((g259) & (g283) & (g286) & (g293) & (g295) & (g300)));
	assign g302 = (((!g209) & (!sk[56]) & (g215)) + ((g209) & (!sk[56]) & (g215)) + ((g209) & (sk[56]) & (g215)));
	assign g303 = (((!ax22x) & (!ax11x) & (!g4) & (sk[57]) & (!ax12x)) + ((!ax22x) & (!ax11x) & (g4) & (!sk[57]) & (!ax12x)) + ((!ax22x) & (!ax11x) & (g4) & (!sk[57]) & (ax12x)) + ((!ax22x) & (!ax11x) & (g4) & (sk[57]) & (ax12x)) + ((!ax22x) & (ax11x) & (!g4) & (sk[57]) & (!ax12x)) + ((!ax22x) & (ax11x) & (g4) & (!sk[57]) & (!ax12x)) + ((!ax22x) & (ax11x) & (g4) & (!sk[57]) & (ax12x)) + ((!ax22x) & (ax11x) & (g4) & (sk[57]) & (!ax12x)) + ((ax22x) & (!ax11x) & (!g4) & (!sk[57]) & (!ax12x)) + ((ax22x) & (!ax11x) & (!g4) & (!sk[57]) & (ax12x)) + ((ax22x) & (!ax11x) & (!g4) & (sk[57]) & (ax12x)) + ((ax22x) & (!ax11x) & (g4) & (!sk[57]) & (!ax12x)) + ((ax22x) & (!ax11x) & (g4) & (!sk[57]) & (ax12x)) + ((ax22x) & (!ax11x) & (g4) & (sk[57]) & (ax12x)) + ((ax22x) & (ax11x) & (!g4) & (!sk[57]) & (!ax12x)) + ((ax22x) & (ax11x) & (!g4) & (!sk[57]) & (ax12x)) + ((ax22x) & (ax11x) & (!g4) & (sk[57]) & (ax12x)) + ((ax22x) & (ax11x) & (g4) & (!sk[57]) & (!ax12x)) + ((ax22x) & (ax11x) & (g4) & (!sk[57]) & (ax12x)) + ((ax22x) & (ax11x) & (g4) & (sk[57]) & (ax12x)));
	assign g304 = (((!g202) & (!g301) & (!sk[58]) & (!g251) & (g302) & (!g303)) + ((!g202) & (!g301) & (!sk[58]) & (!g251) & (g302) & (g303)) + ((!g202) & (!g301) & (!sk[58]) & (g251) & (g302) & (!g303)) + ((!g202) & (!g301) & (!sk[58]) & (g251) & (g302) & (g303)) + ((!g202) & (!g301) & (sk[58]) & (g251) & (!g302) & (!g303)) + ((!g202) & (!g301) & (sk[58]) & (g251) & (g302) & (g303)) + ((!g202) & (g301) & (!sk[58]) & (!g251) & (!g302) & (!g303)) + ((!g202) & (g301) & (!sk[58]) & (!g251) & (!g302) & (g303)) + ((!g202) & (g301) & (!sk[58]) & (!g251) & (g302) & (!g303)) + ((!g202) & (g301) & (!sk[58]) & (!g251) & (g302) & (g303)) + ((!g202) & (g301) & (!sk[58]) & (g251) & (!g302) & (!g303)) + ((!g202) & (g301) & (!sk[58]) & (g251) & (!g302) & (g303)) + ((!g202) & (g301) & (!sk[58]) & (g251) & (g302) & (!g303)) + ((!g202) & (g301) & (!sk[58]) & (g251) & (g302) & (g303)) + ((!g202) & (g301) & (sk[58]) & (!g251) & (!g302) & (!g303)) + ((!g202) & (g301) & (sk[58]) & (!g251) & (g302) & (g303)) + ((!g202) & (g301) & (sk[58]) & (g251) & (!g302) & (!g303)) + ((!g202) & (g301) & (sk[58]) & (g251) & (!g302) & (g303)) + ((g202) & (!g301) & (!sk[58]) & (!g251) & (g302) & (!g303)) + ((g202) & (!g301) & (!sk[58]) & (!g251) & (g302) & (g303)) + ((g202) & (!g301) & (!sk[58]) & (g251) & (!g302) & (!g303)) + ((g202) & (!g301) & (!sk[58]) & (g251) & (!g302) & (g303)) + ((g202) & (!g301) & (!sk[58]) & (g251) & (g302) & (!g303)) + ((g202) & (!g301) & (!sk[58]) & (g251) & (g302) & (g303)) + ((g202) & (!g301) & (sk[58]) & (!g251) & (g302) & (!g303)) + ((g202) & (!g301) & (sk[58]) & (!g251) & (g302) & (g303)) + ((g202) & (!g301) & (sk[58]) & (g251) & (!g302) & (!g303)) + ((g202) & (!g301) & (sk[58]) & (g251) & (g302) & (g303)) + ((g202) & (g301) & (!sk[58]) & (!g251) & (!g302) & (!g303)) + ((g202) & (g301) & (!sk[58]) & (!g251) & (!g302) & (g303)) + ((g202) & (g301) & (!sk[58]) & (!g251) & (g302) & (!g303)) + ((g202) & (g301) & (!sk[58]) & (!g251) & (g302) & (g303)) + ((g202) & (g301) & (!sk[58]) & (g251) & (!g302) & (!g303)) + ((g202) & (g301) & (!sk[58]) & (g251) & (!g302) & (g303)) + ((g202) & (g301) & (!sk[58]) & (g251) & (g302) & (!g303)) + ((g202) & (g301) & (!sk[58]) & (g251) & (g302) & (g303)) + ((g202) & (g301) & (sk[58]) & (!g251) & (!g302) & (!g303)) + ((g202) & (g301) & (sk[58]) & (!g251) & (g302) & (g303)));
	assign g305 = (((!sk[59]) & (!ax22x) & (!ax9x) & (g199) & (!ax8x)) + ((!sk[59]) & (!ax22x) & (!ax9x) & (g199) & (ax8x)) + ((!sk[59]) & (!ax22x) & (ax9x) & (g199) & (!ax8x)) + ((!sk[59]) & (!ax22x) & (ax9x) & (g199) & (ax8x)) + ((!sk[59]) & (ax22x) & (!ax9x) & (!g199) & (!ax8x)) + ((!sk[59]) & (ax22x) & (!ax9x) & (!g199) & (ax8x)) + ((!sk[59]) & (ax22x) & (!ax9x) & (g199) & (!ax8x)) + ((!sk[59]) & (ax22x) & (!ax9x) & (g199) & (ax8x)) + ((!sk[59]) & (ax22x) & (ax9x) & (!g199) & (!ax8x)) + ((!sk[59]) & (ax22x) & (ax9x) & (!g199) & (ax8x)) + ((!sk[59]) & (ax22x) & (ax9x) & (g199) & (!ax8x)) + ((!sk[59]) & (ax22x) & (ax9x) & (g199) & (ax8x)) + ((sk[59]) & (!ax22x) & (!ax9x) & (!g199) & (!ax8x)) + ((sk[59]) & (!ax22x) & (!ax9x) & (!g199) & (ax8x)) + ((sk[59]) & (!ax22x) & (!ax9x) & (g199) & (ax8x)) + ((sk[59]) & (!ax22x) & (ax9x) & (g199) & (!ax8x)) + ((sk[59]) & (ax22x) & (ax9x) & (!g199) & (!ax8x)) + ((sk[59]) & (ax22x) & (ax9x) & (!g199) & (ax8x)) + ((sk[59]) & (ax22x) & (ax9x) & (g199) & (!ax8x)) + ((sk[59]) & (ax22x) & (ax9x) & (g199) & (ax8x)));
	assign g306 = (((!g218) & (!sk[60]) & (!g220) & (!g221) & (g305) & (!g222)) + ((!g218) & (!sk[60]) & (!g220) & (!g221) & (g305) & (g222)) + ((!g218) & (!sk[60]) & (!g220) & (g221) & (g305) & (!g222)) + ((!g218) & (!sk[60]) & (!g220) & (g221) & (g305) & (g222)) + ((!g218) & (!sk[60]) & (g220) & (!g221) & (!g305) & (!g222)) + ((!g218) & (!sk[60]) & (g220) & (!g221) & (!g305) & (g222)) + ((!g218) & (!sk[60]) & (g220) & (!g221) & (g305) & (!g222)) + ((!g218) & (!sk[60]) & (g220) & (!g221) & (g305) & (g222)) + ((!g218) & (!sk[60]) & (g220) & (g221) & (!g305) & (!g222)) + ((!g218) & (!sk[60]) & (g220) & (g221) & (!g305) & (g222)) + ((!g218) & (!sk[60]) & (g220) & (g221) & (g305) & (!g222)) + ((!g218) & (!sk[60]) & (g220) & (g221) & (g305) & (g222)) + ((!g218) & (sk[60]) & (!g220) & (g221) & (!g305) & (!g222)) + ((!g218) & (sk[60]) & (!g220) & (g221) & (!g305) & (g222)) + ((!g218) & (sk[60]) & (g220) & (g221) & (!g305) & (!g222)) + ((!g218) & (sk[60]) & (g220) & (g221) & (g305) & (!g222)) + ((g218) & (!sk[60]) & (!g220) & (!g221) & (g305) & (!g222)) + ((g218) & (!sk[60]) & (!g220) & (!g221) & (g305) & (g222)) + ((g218) & (!sk[60]) & (!g220) & (g221) & (!g305) & (!g222)) + ((g218) & (!sk[60]) & (!g220) & (g221) & (!g305) & (g222)) + ((g218) & (!sk[60]) & (!g220) & (g221) & (g305) & (!g222)) + ((g218) & (!sk[60]) & (!g220) & (g221) & (g305) & (g222)) + ((g218) & (!sk[60]) & (g220) & (!g221) & (!g305) & (!g222)) + ((g218) & (!sk[60]) & (g220) & (!g221) & (!g305) & (g222)) + ((g218) & (!sk[60]) & (g220) & (!g221) & (g305) & (!g222)) + ((g218) & (!sk[60]) & (g220) & (!g221) & (g305) & (g222)) + ((g218) & (!sk[60]) & (g220) & (g221) & (!g305) & (!g222)) + ((g218) & (!sk[60]) & (g220) & (g221) & (!g305) & (g222)) + ((g218) & (!sk[60]) & (g220) & (g221) & (g305) & (!g222)) + ((g218) & (!sk[60]) & (g220) & (g221) & (g305) & (g222)) + ((g218) & (sk[60]) & (!g220) & (!g221) & (g305) & (!g222)) + ((g218) & (sk[60]) & (!g220) & (!g221) & (g305) & (g222)) + ((g218) & (sk[60]) & (!g220) & (g221) & (!g305) & (!g222)) + ((g218) & (sk[60]) & (!g220) & (g221) & (!g305) & (g222)) + ((g218) & (sk[60]) & (!g220) & (g221) & (g305) & (!g222)) + ((g218) & (sk[60]) & (!g220) & (g221) & (g305) & (g222)) + ((g218) & (sk[60]) & (g220) & (!g221) & (!g305) & (g222)) + ((g218) & (sk[60]) & (g220) & (!g221) & (g305) & (g222)) + ((g218) & (sk[60]) & (g220) & (g221) & (!g305) & (!g222)) + ((g218) & (sk[60]) & (g220) & (g221) & (!g305) & (g222)) + ((g218) & (sk[60]) & (g220) & (g221) & (g305) & (!g222)) + ((g218) & (sk[60]) & (g220) & (g221) & (g305) & (g222)));
	assign g307 = (((!g201) & (!sk[61]) & (!g223) & (!g281) & (g304) & (!g306)) + ((!g201) & (!sk[61]) & (!g223) & (!g281) & (g304) & (g306)) + ((!g201) & (!sk[61]) & (!g223) & (g281) & (g304) & (!g306)) + ((!g201) & (!sk[61]) & (!g223) & (g281) & (g304) & (g306)) + ((!g201) & (!sk[61]) & (g223) & (!g281) & (!g304) & (!g306)) + ((!g201) & (!sk[61]) & (g223) & (!g281) & (!g304) & (g306)) + ((!g201) & (!sk[61]) & (g223) & (!g281) & (g304) & (!g306)) + ((!g201) & (!sk[61]) & (g223) & (!g281) & (g304) & (g306)) + ((!g201) & (!sk[61]) & (g223) & (g281) & (!g304) & (!g306)) + ((!g201) & (!sk[61]) & (g223) & (g281) & (!g304) & (g306)) + ((!g201) & (!sk[61]) & (g223) & (g281) & (g304) & (!g306)) + ((!g201) & (!sk[61]) & (g223) & (g281) & (g304) & (g306)) + ((!g201) & (sk[61]) & (g223) & (!g281) & (g304) & (g306)) + ((!g201) & (sk[61]) & (g223) & (g281) & (!g304) & (g306)) + ((!g201) & (sk[61]) & (g223) & (g281) & (g304) & (!g306)) + ((!g201) & (sk[61]) & (g223) & (g281) & (g304) & (g306)) + ((g201) & (!sk[61]) & (!g223) & (!g281) & (g304) & (!g306)) + ((g201) & (!sk[61]) & (!g223) & (!g281) & (g304) & (g306)) + ((g201) & (!sk[61]) & (!g223) & (g281) & (!g304) & (!g306)) + ((g201) & (!sk[61]) & (!g223) & (g281) & (!g304) & (g306)) + ((g201) & (!sk[61]) & (!g223) & (g281) & (g304) & (!g306)) + ((g201) & (!sk[61]) & (!g223) & (g281) & (g304) & (g306)) + ((g201) & (!sk[61]) & (g223) & (!g281) & (!g304) & (!g306)) + ((g201) & (!sk[61]) & (g223) & (!g281) & (!g304) & (g306)) + ((g201) & (!sk[61]) & (g223) & (!g281) & (g304) & (!g306)) + ((g201) & (!sk[61]) & (g223) & (!g281) & (g304) & (g306)) + ((g201) & (!sk[61]) & (g223) & (g281) & (!g304) & (!g306)) + ((g201) & (!sk[61]) & (g223) & (g281) & (!g304) & (g306)) + ((g201) & (!sk[61]) & (g223) & (g281) & (g304) & (!g306)) + ((g201) & (!sk[61]) & (g223) & (g281) & (g304) & (g306)) + ((g201) & (sk[61]) & (!g223) & (!g281) & (g304) & (g306)) + ((g201) & (sk[61]) & (!g223) & (g281) & (!g304) & (g306)) + ((g201) & (sk[61]) & (!g223) & (g281) & (g304) & (!g306)) + ((g201) & (sk[61]) & (!g223) & (g281) & (g304) & (g306)) + ((g201) & (sk[61]) & (g223) & (!g281) & (!g304) & (!g306)) + ((g201) & (sk[61]) & (g223) & (!g281) & (!g304) & (g306)) + ((g201) & (sk[61]) & (g223) & (!g281) & (g304) & (!g306)) + ((g201) & (sk[61]) & (g223) & (!g281) & (g304) & (g306)) + ((g201) & (sk[61]) & (g223) & (g281) & (!g304) & (!g306)) + ((g201) & (sk[61]) & (g223) & (g281) & (!g304) & (g306)) + ((g201) & (sk[61]) & (g223) & (g281) & (g304) & (!g306)) + ((g201) & (sk[61]) & (g223) & (g281) & (g304) & (g306)));
	assign g308 = (((!g251) & (!g122) & (!sk[62]) & (g280)) + ((!g251) & (!g122) & (sk[62]) & (g280)) + ((!g251) & (g122) & (!sk[62]) & (g280)) + ((!g251) & (g122) & (sk[62]) & (!g280)) + ((!g251) & (g122) & (sk[62]) & (g280)) + ((g251) & (!g122) & (!sk[62]) & (!g280)) + ((g251) & (!g122) & (!sk[62]) & (g280)) + ((g251) & (g122) & (!sk[62]) & (!g280)) + ((g251) & (g122) & (!sk[62]) & (g280)));
	assign g309 = (((!g69) & (!g305) & (!g308) & (sk[63]) & (g222)) + ((!g69) & (!g305) & (g308) & (!sk[63]) & (!g222)) + ((!g69) & (!g305) & (g308) & (!sk[63]) & (g222)) + ((!g69) & (!g305) & (g308) & (sk[63]) & (!g222)) + ((!g69) & (g305) & (!g308) & (sk[63]) & (!g222)) + ((!g69) & (g305) & (g308) & (!sk[63]) & (!g222)) + ((!g69) & (g305) & (g308) & (!sk[63]) & (g222)) + ((!g69) & (g305) & (g308) & (sk[63]) & (g222)) + ((g69) & (!g305) & (!g308) & (!sk[63]) & (!g222)) + ((g69) & (!g305) & (!g308) & (!sk[63]) & (g222)) + ((g69) & (!g305) & (g308) & (!sk[63]) & (!g222)) + ((g69) & (!g305) & (g308) & (!sk[63]) & (g222)) + ((g69) & (!g305) & (g308) & (sk[63]) & (!g222)) + ((g69) & (!g305) & (g308) & (sk[63]) & (g222)) + ((g69) & (g305) & (!g308) & (!sk[63]) & (!g222)) + ((g69) & (g305) & (!g308) & (!sk[63]) & (g222)) + ((g69) & (g305) & (g308) & (!sk[63]) & (!g222)) + ((g69) & (g305) & (g308) & (!sk[63]) & (g222)) + ((g69) & (g305) & (g308) & (sk[63]) & (!g222)) + ((g69) & (g305) & (g308) & (sk[63]) & (g222)));
	assign g310 = (((!sk[64]) & (!g202) & (!g218) & (!g220) & (g303) & (!g221)) + ((!sk[64]) & (!g202) & (!g218) & (!g220) & (g303) & (g221)) + ((!sk[64]) & (!g202) & (!g218) & (g220) & (g303) & (!g221)) + ((!sk[64]) & (!g202) & (!g218) & (g220) & (g303) & (g221)) + ((!sk[64]) & (!g202) & (g218) & (!g220) & (!g303) & (!g221)) + ((!sk[64]) & (!g202) & (g218) & (!g220) & (!g303) & (g221)) + ((!sk[64]) & (!g202) & (g218) & (!g220) & (g303) & (!g221)) + ((!sk[64]) & (!g202) & (g218) & (!g220) & (g303) & (g221)) + ((!sk[64]) & (!g202) & (g218) & (g220) & (!g303) & (!g221)) + ((!sk[64]) & (!g202) & (g218) & (g220) & (!g303) & (g221)) + ((!sk[64]) & (!g202) & (g218) & (g220) & (g303) & (!g221)) + ((!sk[64]) & (!g202) & (g218) & (g220) & (g303) & (g221)) + ((!sk[64]) & (g202) & (!g218) & (!g220) & (g303) & (!g221)) + ((!sk[64]) & (g202) & (!g218) & (!g220) & (g303) & (g221)) + ((!sk[64]) & (g202) & (!g218) & (g220) & (!g303) & (!g221)) + ((!sk[64]) & (g202) & (!g218) & (g220) & (!g303) & (g221)) + ((!sk[64]) & (g202) & (!g218) & (g220) & (g303) & (!g221)) + ((!sk[64]) & (g202) & (!g218) & (g220) & (g303) & (g221)) + ((!sk[64]) & (g202) & (g218) & (!g220) & (!g303) & (!g221)) + ((!sk[64]) & (g202) & (g218) & (!g220) & (!g303) & (g221)) + ((!sk[64]) & (g202) & (g218) & (!g220) & (g303) & (!g221)) + ((!sk[64]) & (g202) & (g218) & (!g220) & (g303) & (g221)) + ((!sk[64]) & (g202) & (g218) & (g220) & (!g303) & (!g221)) + ((!sk[64]) & (g202) & (g218) & (g220) & (!g303) & (g221)) + ((!sk[64]) & (g202) & (g218) & (g220) & (g303) & (!g221)) + ((!sk[64]) & (g202) & (g218) & (g220) & (g303) & (g221)) + ((sk[64]) & (!g202) & (!g218) & (!g220) & (!g303) & (g221)) + ((sk[64]) & (!g202) & (!g218) & (!g220) & (g303) & (g221)) + ((sk[64]) & (!g202) & (!g218) & (g220) & (!g303) & (g221)) + ((sk[64]) & (!g202) & (g218) & (!g220) & (!g303) & (g221)) + ((sk[64]) & (!g202) & (g218) & (!g220) & (g303) & (g221)) + ((sk[64]) & (!g202) & (g218) & (g220) & (!g303) & (g221)) + ((sk[64]) & (!g202) & (g218) & (g220) & (g303) & (!g221)) + ((sk[64]) & (!g202) & (g218) & (g220) & (g303) & (g221)) + ((sk[64]) & (g202) & (!g218) & (g220) & (!g303) & (g221)) + ((sk[64]) & (g202) & (g218) & (!g220) & (!g303) & (!g221)) + ((sk[64]) & (g202) & (g218) & (!g220) & (!g303) & (g221)) + ((sk[64]) & (g202) & (g218) & (!g220) & (g303) & (!g221)) + ((sk[64]) & (g202) & (g218) & (!g220) & (g303) & (g221)) + ((sk[64]) & (g202) & (g218) & (g220) & (!g303) & (g221)) + ((sk[64]) & (g202) & (g218) & (g220) & (g303) & (!g221)) + ((sk[64]) & (g202) & (g218) & (g220) & (g303) & (g221)));
	assign g311 = (((!g301) & (!sk[65]) & (!g251) & (!g302) & (g252) & (!g253)) + ((!g301) & (!sk[65]) & (!g251) & (!g302) & (g252) & (g253)) + ((!g301) & (!sk[65]) & (!g251) & (g302) & (g252) & (!g253)) + ((!g301) & (!sk[65]) & (!g251) & (g302) & (g252) & (g253)) + ((!g301) & (!sk[65]) & (g251) & (!g302) & (!g252) & (!g253)) + ((!g301) & (!sk[65]) & (g251) & (!g302) & (!g252) & (g253)) + ((!g301) & (!sk[65]) & (g251) & (!g302) & (g252) & (!g253)) + ((!g301) & (!sk[65]) & (g251) & (!g302) & (g252) & (g253)) + ((!g301) & (!sk[65]) & (g251) & (g302) & (!g252) & (!g253)) + ((!g301) & (!sk[65]) & (g251) & (g302) & (!g252) & (g253)) + ((!g301) & (!sk[65]) & (g251) & (g302) & (g252) & (!g253)) + ((!g301) & (!sk[65]) & (g251) & (g302) & (g252) & (g253)) + ((!g301) & (sk[65]) & (!g251) & (g302) & (!g252) & (g253)) + ((!g301) & (sk[65]) & (!g251) & (g302) & (g252) & (g253)) + ((!g301) & (sk[65]) & (g251) & (!g302) & (!g252) & (!g253)) + ((!g301) & (sk[65]) & (g251) & (!g302) & (!g252) & (g253)) + ((!g301) & (sk[65]) & (g251) & (g302) & (g252) & (!g253)) + ((!g301) & (sk[65]) & (g251) & (g302) & (g252) & (g253)) + ((g301) & (!sk[65]) & (!g251) & (!g302) & (g252) & (!g253)) + ((g301) & (!sk[65]) & (!g251) & (!g302) & (g252) & (g253)) + ((g301) & (!sk[65]) & (!g251) & (g302) & (!g252) & (!g253)) + ((g301) & (!sk[65]) & (!g251) & (g302) & (!g252) & (g253)) + ((g301) & (!sk[65]) & (!g251) & (g302) & (g252) & (!g253)) + ((g301) & (!sk[65]) & (!g251) & (g302) & (g252) & (g253)) + ((g301) & (!sk[65]) & (g251) & (!g302) & (!g252) & (!g253)) + ((g301) & (!sk[65]) & (g251) & (!g302) & (!g252) & (g253)) + ((g301) & (!sk[65]) & (g251) & (!g302) & (g252) & (!g253)) + ((g301) & (!sk[65]) & (g251) & (!g302) & (g252) & (g253)) + ((g301) & (!sk[65]) & (g251) & (g302) & (!g252) & (!g253)) + ((g301) & (!sk[65]) & (g251) & (g302) & (!g252) & (g253)) + ((g301) & (!sk[65]) & (g251) & (g302) & (g252) & (!g253)) + ((g301) & (!sk[65]) & (g251) & (g302) & (g252) & (g253)) + ((g301) & (sk[65]) & (!g251) & (!g302) & (!g252) & (!g253)) + ((g301) & (sk[65]) & (!g251) & (!g302) & (!g252) & (g253)) + ((g301) & (sk[65]) & (!g251) & (g302) & (g252) & (!g253)) + ((g301) & (sk[65]) & (!g251) & (g302) & (g252) & (g253)) + ((g301) & (sk[65]) & (g251) & (!g302) & (!g252) & (!g253)) + ((g301) & (sk[65]) & (g251) & (!g302) & (g252) & (!g253)));
	assign g312 = (((!g251) & (!sk[66]) & (!g252) & (g122) & (!g280)) + ((!g251) & (!sk[66]) & (!g252) & (g122) & (g280)) + ((!g251) & (!sk[66]) & (g252) & (g122) & (!g280)) + ((!g251) & (!sk[66]) & (g252) & (g122) & (g280)) + ((!g251) & (sk[66]) & (!g252) & (!g122) & (g280)) + ((!g251) & (sk[66]) & (!g252) & (g122) & (!g280)) + ((!g251) & (sk[66]) & (!g252) & (g122) & (g280)) + ((!g251) & (sk[66]) & (g252) & (!g122) & (g280)) + ((!g251) & (sk[66]) & (g252) & (g122) & (!g280)) + ((g251) & (!sk[66]) & (!g252) & (!g122) & (!g280)) + ((g251) & (!sk[66]) & (!g252) & (!g122) & (g280)) + ((g251) & (!sk[66]) & (!g252) & (g122) & (!g280)) + ((g251) & (!sk[66]) & (!g252) & (g122) & (g280)) + ((g251) & (!sk[66]) & (g252) & (!g122) & (!g280)) + ((g251) & (!sk[66]) & (g252) & (!g122) & (g280)) + ((g251) & (!sk[66]) & (g252) & (g122) & (!g280)) + ((g251) & (!sk[66]) & (g252) & (g122) & (g280)) + ((g251) & (sk[66]) & (g252) & (!g122) & (!g280)));
	assign g313 = (((!g301) & (!sk[67]) & (!g251) & (!g302) & (g253) & (!g303)) + ((!g301) & (!sk[67]) & (!g251) & (!g302) & (g253) & (g303)) + ((!g301) & (!sk[67]) & (!g251) & (g302) & (g253) & (!g303)) + ((!g301) & (!sk[67]) & (!g251) & (g302) & (g253) & (g303)) + ((!g301) & (!sk[67]) & (g251) & (!g302) & (!g253) & (!g303)) + ((!g301) & (!sk[67]) & (g251) & (!g302) & (!g253) & (g303)) + ((!g301) & (!sk[67]) & (g251) & (!g302) & (g253) & (!g303)) + ((!g301) & (!sk[67]) & (g251) & (!g302) & (g253) & (g303)) + ((!g301) & (!sk[67]) & (g251) & (g302) & (!g253) & (!g303)) + ((!g301) & (!sk[67]) & (g251) & (g302) & (!g253) & (g303)) + ((!g301) & (!sk[67]) & (g251) & (g302) & (g253) & (!g303)) + ((!g301) & (!sk[67]) & (g251) & (g302) & (g253) & (g303)) + ((!g301) & (sk[67]) & (!g251) & (g302) & (!g253) & (g303)) + ((!g301) & (sk[67]) & (!g251) & (g302) & (g253) & (g303)) + ((!g301) & (sk[67]) & (g251) & (!g302) & (!g253) & (!g303)) + ((!g301) & (sk[67]) & (g251) & (!g302) & (!g253) & (g303)) + ((!g301) & (sk[67]) & (g251) & (g302) & (g253) & (!g303)) + ((!g301) & (sk[67]) & (g251) & (g302) & (g253) & (g303)) + ((g301) & (!sk[67]) & (!g251) & (!g302) & (g253) & (!g303)) + ((g301) & (!sk[67]) & (!g251) & (!g302) & (g253) & (g303)) + ((g301) & (!sk[67]) & (!g251) & (g302) & (!g253) & (!g303)) + ((g301) & (!sk[67]) & (!g251) & (g302) & (!g253) & (g303)) + ((g301) & (!sk[67]) & (!g251) & (g302) & (g253) & (!g303)) + ((g301) & (!sk[67]) & (!g251) & (g302) & (g253) & (g303)) + ((g301) & (!sk[67]) & (g251) & (!g302) & (!g253) & (!g303)) + ((g301) & (!sk[67]) & (g251) & (!g302) & (!g253) & (g303)) + ((g301) & (!sk[67]) & (g251) & (!g302) & (g253) & (!g303)) + ((g301) & (!sk[67]) & (g251) & (!g302) & (g253) & (g303)) + ((g301) & (!sk[67]) & (g251) & (g302) & (!g253) & (!g303)) + ((g301) & (!sk[67]) & (g251) & (g302) & (!g253) & (g303)) + ((g301) & (!sk[67]) & (g251) & (g302) & (g253) & (!g303)) + ((g301) & (!sk[67]) & (g251) & (g302) & (g253) & (g303)) + ((g301) & (sk[67]) & (!g251) & (!g302) & (!g253) & (!g303)) + ((g301) & (sk[67]) & (!g251) & (!g302) & (!g253) & (g303)) + ((g301) & (sk[67]) & (!g251) & (g302) & (g253) & (!g303)) + ((g301) & (sk[67]) & (!g251) & (g302) & (g253) & (g303)) + ((g301) & (sk[67]) & (g251) & (!g302) & (!g253) & (!g303)) + ((g301) & (sk[67]) & (g251) & (!g302) & (g253) & (!g303)));
	assign g314 = (((!g69) & (!g305) & (!g312) & (sk[68]) & (!g313)) + ((!g69) & (!g305) & (g312) & (!sk[68]) & (!g313)) + ((!g69) & (!g305) & (g312) & (!sk[68]) & (g313)) + ((!g69) & (g305) & (!g312) & (sk[68]) & (!g313)) + ((!g69) & (g305) & (!g312) & (sk[68]) & (g313)) + ((!g69) & (g305) & (g312) & (!sk[68]) & (!g313)) + ((!g69) & (g305) & (g312) & (!sk[68]) & (g313)) + ((!g69) & (g305) & (g312) & (sk[68]) & (!g313)) + ((g69) & (!g305) & (!g312) & (!sk[68]) & (!g313)) + ((g69) & (!g305) & (!g312) & (!sk[68]) & (g313)) + ((g69) & (!g305) & (!g312) & (sk[68]) & (!g313)) + ((g69) & (!g305) & (g312) & (!sk[68]) & (!g313)) + ((g69) & (!g305) & (g312) & (!sk[68]) & (g313)) + ((g69) & (g305) & (!g312) & (!sk[68]) & (!g313)) + ((g69) & (g305) & (!g312) & (!sk[68]) & (g313)) + ((g69) & (g305) & (!g312) & (sk[68]) & (!g313)) + ((g69) & (g305) & (g312) & (!sk[68]) & (!g313)) + ((g69) & (g305) & (g312) & (!sk[68]) & (g313)));
	assign g315 = (((!g310) & (!g311) & (!sk[69]) & (g314)) + ((!g310) & (!g311) & (sk[69]) & (!g314)) + ((!g310) & (g311) & (!sk[69]) & (g314)) + ((!g310) & (g311) & (sk[69]) & (g314)) + ((g310) & (!g311) & (!sk[69]) & (!g314)) + ((g310) & (!g311) & (!sk[69]) & (g314)) + ((g310) & (!g311) & (sk[69]) & (g314)) + ((g310) & (g311) & (!sk[69]) & (!g314)) + ((g310) & (g311) & (!sk[69]) & (g314)) + ((g310) & (g311) & (sk[69]) & (!g314)));
	assign g316 = (((!g307) & (!g309) & (!sk[70]) & (g315)) + ((!g307) & (!g309) & (sk[70]) & (g315)) + ((!g307) & (g309) & (!sk[70]) & (g315)) + ((g307) & (!g309) & (!sk[70]) & (!g315)) + ((g307) & (!g309) & (!sk[70]) & (g315)) + ((g307) & (!g309) & (sk[70]) & (!g315)) + ((g307) & (!g309) & (sk[70]) & (g315)) + ((g307) & (g309) & (!sk[70]) & (!g315)) + ((g307) & (g309) & (!sk[70]) & (g315)) + ((g307) & (g309) & (sk[70]) & (g315)));
	assign g317 = (((!g69) & (!g305) & (!sk[71]) & (g308) & (!g222)) + ((!g69) & (!g305) & (!sk[71]) & (g308) & (g222)) + ((!g69) & (!g305) & (sk[71]) & (!g308) & (g222)) + ((!g69) & (g305) & (!sk[71]) & (g308) & (!g222)) + ((!g69) & (g305) & (!sk[71]) & (g308) & (g222)) + ((!g69) & (g305) & (sk[71]) & (!g308) & (!g222)) + ((!g69) & (g305) & (sk[71]) & (!g308) & (g222)) + ((!g69) & (g305) & (sk[71]) & (g308) & (g222)) + ((g69) & (!g305) & (!sk[71]) & (!g308) & (!g222)) + ((g69) & (!g305) & (!sk[71]) & (!g308) & (g222)) + ((g69) & (!g305) & (!sk[71]) & (g308) & (!g222)) + ((g69) & (!g305) & (!sk[71]) & (g308) & (g222)) + ((g69) & (g305) & (!sk[71]) & (!g308) & (!g222)) + ((g69) & (g305) & (!sk[71]) & (!g308) & (g222)) + ((g69) & (g305) & (!sk[71]) & (g308) & (!g222)) + ((g69) & (g305) & (!sk[71]) & (g308) & (g222)));
	assign g318 = (((!sk[72]) & (!g310) & (!g311) & (g314)) + ((!sk[72]) & (!g310) & (g311) & (g314)) + ((!sk[72]) & (g310) & (!g311) & (!g314)) + ((!sk[72]) & (g310) & (!g311) & (g314)) + ((!sk[72]) & (g310) & (g311) & (!g314)) + ((!sk[72]) & (g310) & (g311) & (g314)) + ((sk[72]) & (!g310) & (g311) & (!g314)) + ((sk[72]) & (g310) & (!g311) & (!g314)) + ((sk[72]) & (g310) & (g311) & (!g314)) + ((sk[72]) & (g310) & (g311) & (g314)));
	assign g319 = (((!sk[73]) & (!g301) & (!g251) & (g302) & (!g252)) + ((!sk[73]) & (!g301) & (!g251) & (g302) & (g252)) + ((!sk[73]) & (!g301) & (g251) & (g302) & (!g252)) + ((!sk[73]) & (!g301) & (g251) & (g302) & (g252)) + ((!sk[73]) & (g301) & (!g251) & (!g302) & (!g252)) + ((!sk[73]) & (g301) & (!g251) & (!g302) & (g252)) + ((!sk[73]) & (g301) & (!g251) & (g302) & (!g252)) + ((!sk[73]) & (g301) & (!g251) & (g302) & (g252)) + ((!sk[73]) & (g301) & (g251) & (!g302) & (!g252)) + ((!sk[73]) & (g301) & (g251) & (!g302) & (g252)) + ((!sk[73]) & (g301) & (g251) & (g302) & (!g252)) + ((!sk[73]) & (g301) & (g251) & (g302) & (g252)) + ((sk[73]) & (!g301) & (!g251) & (g302) & (g252)) + ((sk[73]) & (!g301) & (g251) & (!g302) & (!g252)) + ((sk[73]) & (!g301) & (g251) & (!g302) & (g252)) + ((sk[73]) & (g301) & (!g251) & (!g302) & (!g252)) + ((sk[73]) & (g301) & (!g251) & (!g302) & (g252)) + ((sk[73]) & (g301) & (g251) & (!g302) & (!g252)));
	assign g320 = (((!g218) & (!g253) & (!g220) & (!sk[74]) & (g303) & (!g221)) + ((!g218) & (!g253) & (!g220) & (!sk[74]) & (g303) & (g221)) + ((!g218) & (!g253) & (!g220) & (sk[74]) & (!g303) & (g221)) + ((!g218) & (!g253) & (g220) & (!sk[74]) & (g303) & (!g221)) + ((!g218) & (!g253) & (g220) & (!sk[74]) & (g303) & (g221)) + ((!g218) & (!g253) & (g220) & (sk[74]) & (!g303) & (g221)) + ((!g218) & (!g253) & (g220) & (sk[74]) & (g303) & (g221)) + ((!g218) & (g253) & (!g220) & (!sk[74]) & (!g303) & (!g221)) + ((!g218) & (g253) & (!g220) & (!sk[74]) & (!g303) & (g221)) + ((!g218) & (g253) & (!g220) & (!sk[74]) & (g303) & (!g221)) + ((!g218) & (g253) & (!g220) & (!sk[74]) & (g303) & (g221)) + ((!g218) & (g253) & (!g220) & (sk[74]) & (!g303) & (g221)) + ((!g218) & (g253) & (g220) & (!sk[74]) & (!g303) & (!g221)) + ((!g218) & (g253) & (g220) & (!sk[74]) & (!g303) & (g221)) + ((!g218) & (g253) & (g220) & (!sk[74]) & (g303) & (!g221)) + ((!g218) & (g253) & (g220) & (!sk[74]) & (g303) & (g221)) + ((g218) & (!g253) & (!g220) & (!sk[74]) & (g303) & (!g221)) + ((g218) & (!g253) & (!g220) & (!sk[74]) & (g303) & (g221)) + ((g218) & (!g253) & (!g220) & (sk[74]) & (!g303) & (g221)) + ((g218) & (!g253) & (!g220) & (sk[74]) & (g303) & (!g221)) + ((g218) & (!g253) & (!g220) & (sk[74]) & (g303) & (g221)) + ((g218) & (!g253) & (g220) & (!sk[74]) & (!g303) & (!g221)) + ((g218) & (!g253) & (g220) & (!sk[74]) & (!g303) & (g221)) + ((g218) & (!g253) & (g220) & (!sk[74]) & (g303) & (!g221)) + ((g218) & (!g253) & (g220) & (!sk[74]) & (g303) & (g221)) + ((g218) & (!g253) & (g220) & (sk[74]) & (!g303) & (g221)) + ((g218) & (!g253) & (g220) & (sk[74]) & (g303) & (g221)) + ((g218) & (g253) & (!g220) & (!sk[74]) & (!g303) & (!g221)) + ((g218) & (g253) & (!g220) & (!sk[74]) & (!g303) & (g221)) + ((g218) & (g253) & (!g220) & (!sk[74]) & (g303) & (!g221)) + ((g218) & (g253) & (!g220) & (!sk[74]) & (g303) & (g221)) + ((g218) & (g253) & (!g220) & (sk[74]) & (!g303) & (g221)) + ((g218) & (g253) & (!g220) & (sk[74]) & (g303) & (!g221)) + ((g218) & (g253) & (!g220) & (sk[74]) & (g303) & (g221)) + ((g218) & (g253) & (g220) & (!sk[74]) & (!g303) & (!g221)) + ((g218) & (g253) & (g220) & (!sk[74]) & (!g303) & (g221)) + ((g218) & (g253) & (g220) & (!sk[74]) & (g303) & (!g221)) + ((g218) & (g253) & (g220) & (!sk[74]) & (g303) & (g221)) + ((g218) & (g253) & (g220) & (sk[74]) & (!g303) & (!g221)) + ((g218) & (g253) & (g220) & (sk[74]) & (!g303) & (g221)) + ((g218) & (g253) & (g220) & (sk[74]) & (g303) & (!g221)) + ((g218) & (g253) & (g220) & (sk[74]) & (g303) & (g221)));
	assign g321 = (((!g202) & (!g69) & (!sk[75]) & (g319) & (!g320)) + ((!g202) & (!g69) & (!sk[75]) & (g319) & (g320)) + ((!g202) & (!g69) & (sk[75]) & (!g319) & (g320)) + ((!g202) & (!g69) & (sk[75]) & (g319) & (!g320)) + ((!g202) & (g69) & (!sk[75]) & (g319) & (!g320)) + ((!g202) & (g69) & (!sk[75]) & (g319) & (g320)) + ((!g202) & (g69) & (sk[75]) & (!g319) & (g320)) + ((!g202) & (g69) & (sk[75]) & (g319) & (!g320)) + ((g202) & (!g69) & (!sk[75]) & (!g319) & (!g320)) + ((g202) & (!g69) & (!sk[75]) & (!g319) & (g320)) + ((g202) & (!g69) & (!sk[75]) & (g319) & (!g320)) + ((g202) & (!g69) & (!sk[75]) & (g319) & (g320)) + ((g202) & (!g69) & (sk[75]) & (!g319) & (!g320)) + ((g202) & (!g69) & (sk[75]) & (g319) & (g320)) + ((g202) & (g69) & (!sk[75]) & (!g319) & (!g320)) + ((g202) & (g69) & (!sk[75]) & (!g319) & (g320)) + ((g202) & (g69) & (!sk[75]) & (g319) & (!g320)) + ((g202) & (g69) & (!sk[75]) & (g319) & (g320)) + ((g202) & (g69) & (sk[75]) & (!g319) & (g320)) + ((g202) & (g69) & (sk[75]) & (g319) & (!g320)));
	assign g322 = (((!g317) & (!g318) & (!sk[76]) & (g321)) + ((!g317) & (!g318) & (sk[76]) & (!g321)) + ((!g317) & (g318) & (!sk[76]) & (g321)) + ((!g317) & (g318) & (sk[76]) & (g321)) + ((g317) & (!g318) & (!sk[76]) & (!g321)) + ((g317) & (!g318) & (!sk[76]) & (g321)) + ((g317) & (!g318) & (sk[76]) & (g321)) + ((g317) & (g318) & (!sk[76]) & (!g321)) + ((g317) & (g318) & (!sk[76]) & (g321)) + ((g317) & (g318) & (sk[76]) & (!g321)));
	assign g323 = (((!g218) & (!g220) & (!g221) & (g305) & (!sk[77]) & (!g200)) + ((!g218) & (!g220) & (!g221) & (g305) & (!sk[77]) & (g200)) + ((!g218) & (!g220) & (g221) & (!g305) & (sk[77]) & (!g200)) + ((!g218) & (!g220) & (g221) & (g305) & (!sk[77]) & (!g200)) + ((!g218) & (!g220) & (g221) & (g305) & (!sk[77]) & (g200)) + ((!g218) & (!g220) & (g221) & (g305) & (sk[77]) & (!g200)) + ((!g218) & (g220) & (!g221) & (!g305) & (!sk[77]) & (!g200)) + ((!g218) & (g220) & (!g221) & (!g305) & (!sk[77]) & (g200)) + ((!g218) & (g220) & (!g221) & (g305) & (!sk[77]) & (!g200)) + ((!g218) & (g220) & (!g221) & (g305) & (!sk[77]) & (g200)) + ((!g218) & (g220) & (g221) & (!g305) & (!sk[77]) & (!g200)) + ((!g218) & (g220) & (g221) & (!g305) & (!sk[77]) & (g200)) + ((!g218) & (g220) & (g221) & (!g305) & (sk[77]) & (!g200)) + ((!g218) & (g220) & (g221) & (!g305) & (sk[77]) & (g200)) + ((!g218) & (g220) & (g221) & (g305) & (!sk[77]) & (!g200)) + ((!g218) & (g220) & (g221) & (g305) & (!sk[77]) & (g200)) + ((g218) & (!g220) & (!g221) & (!g305) & (sk[77]) & (g200)) + ((g218) & (!g220) & (!g221) & (g305) & (!sk[77]) & (!g200)) + ((g218) & (!g220) & (!g221) & (g305) & (!sk[77]) & (g200)) + ((g218) & (!g220) & (!g221) & (g305) & (sk[77]) & (g200)) + ((g218) & (!g220) & (g221) & (!g305) & (!sk[77]) & (!g200)) + ((g218) & (!g220) & (g221) & (!g305) & (!sk[77]) & (g200)) + ((g218) & (!g220) & (g221) & (!g305) & (sk[77]) & (!g200)) + ((g218) & (!g220) & (g221) & (!g305) & (sk[77]) & (g200)) + ((g218) & (!g220) & (g221) & (g305) & (!sk[77]) & (!g200)) + ((g218) & (!g220) & (g221) & (g305) & (!sk[77]) & (g200)) + ((g218) & (!g220) & (g221) & (g305) & (sk[77]) & (!g200)) + ((g218) & (!g220) & (g221) & (g305) & (sk[77]) & (g200)) + ((g218) & (g220) & (!g221) & (!g305) & (!sk[77]) & (!g200)) + ((g218) & (g220) & (!g221) & (!g305) & (!sk[77]) & (g200)) + ((g218) & (g220) & (!g221) & (g305) & (!sk[77]) & (!g200)) + ((g218) & (g220) & (!g221) & (g305) & (!sk[77]) & (g200)) + ((g218) & (g220) & (!g221) & (g305) & (sk[77]) & (!g200)) + ((g218) & (g220) & (!g221) & (g305) & (sk[77]) & (g200)) + ((g218) & (g220) & (g221) & (!g305) & (!sk[77]) & (!g200)) + ((g218) & (g220) & (g221) & (!g305) & (!sk[77]) & (g200)) + ((g218) & (g220) & (g221) & (!g305) & (sk[77]) & (!g200)) + ((g218) & (g220) & (g221) & (!g305) & (sk[77]) & (g200)) + ((g218) & (g220) & (g221) & (g305) & (!sk[77]) & (!g200)) + ((g218) & (g220) & (g221) & (g305) & (!sk[77]) & (g200)) + ((g218) & (g220) & (g221) & (g305) & (sk[77]) & (!g200)) + ((g218) & (g220) & (g221) & (g305) & (sk[77]) & (g200)));
	assign g324 = (((!g202) & (!g301) & (!sk[78]) & (!g251) & (g302) & (!g222)) + ((!g202) & (!g301) & (!sk[78]) & (!g251) & (g302) & (g222)) + ((!g202) & (!g301) & (!sk[78]) & (g251) & (g302) & (!g222)) + ((!g202) & (!g301) & (!sk[78]) & (g251) & (g302) & (g222)) + ((!g202) & (!g301) & (sk[78]) & (!g251) & (g302) & (g222)) + ((!g202) & (!g301) & (sk[78]) & (g251) & (!g302) & (!g222)) + ((!g202) & (!g301) & (sk[78]) & (g251) & (!g302) & (g222)) + ((!g202) & (g301) & (!sk[78]) & (!g251) & (!g302) & (!g222)) + ((!g202) & (g301) & (!sk[78]) & (!g251) & (!g302) & (g222)) + ((!g202) & (g301) & (!sk[78]) & (!g251) & (g302) & (!g222)) + ((!g202) & (g301) & (!sk[78]) & (!g251) & (g302) & (g222)) + ((!g202) & (g301) & (!sk[78]) & (g251) & (!g302) & (!g222)) + ((!g202) & (g301) & (!sk[78]) & (g251) & (!g302) & (g222)) + ((!g202) & (g301) & (!sk[78]) & (g251) & (g302) & (!g222)) + ((!g202) & (g301) & (!sk[78]) & (g251) & (g302) & (g222)) + ((!g202) & (g301) & (sk[78]) & (!g251) & (!g302) & (!g222)) + ((!g202) & (g301) & (sk[78]) & (!g251) & (!g302) & (g222)) + ((!g202) & (g301) & (sk[78]) & (g251) & (!g302) & (!g222)) + ((g202) & (!g301) & (!sk[78]) & (!g251) & (g302) & (!g222)) + ((g202) & (!g301) & (!sk[78]) & (!g251) & (g302) & (g222)) + ((g202) & (!g301) & (!sk[78]) & (g251) & (!g302) & (!g222)) + ((g202) & (!g301) & (!sk[78]) & (g251) & (!g302) & (g222)) + ((g202) & (!g301) & (!sk[78]) & (g251) & (g302) & (!g222)) + ((g202) & (!g301) & (!sk[78]) & (g251) & (g302) & (g222)) + ((g202) & (!g301) & (sk[78]) & (!g251) & (g302) & (g222)) + ((g202) & (!g301) & (sk[78]) & (g251) & (g302) & (!g222)) + ((g202) & (!g301) & (sk[78]) & (g251) & (g302) & (g222)) + ((g202) & (g301) & (!sk[78]) & (!g251) & (!g302) & (!g222)) + ((g202) & (g301) & (!sk[78]) & (!g251) & (!g302) & (g222)) + ((g202) & (g301) & (!sk[78]) & (!g251) & (g302) & (!g222)) + ((g202) & (g301) & (!sk[78]) & (!g251) & (g302) & (g222)) + ((g202) & (g301) & (!sk[78]) & (g251) & (!g302) & (!g222)) + ((g202) & (g301) & (!sk[78]) & (g251) & (!g302) & (g222)) + ((g202) & (g301) & (!sk[78]) & (g251) & (g302) & (!g222)) + ((g202) & (g301) & (!sk[78]) & (g251) & (g302) & (g222)) + ((g202) & (g301) & (sk[78]) & (!g251) & (g302) & (!g222)) + ((g202) & (g301) & (sk[78]) & (!g251) & (g302) & (g222)) + ((g202) & (g301) & (sk[78]) & (g251) & (!g302) & (!g222)));
	assign g325 = (((!sk[79]) & (!g168) & (!g173) & (!g180) & (g183) & (!g192)) + ((!sk[79]) & (!g168) & (!g173) & (!g180) & (g183) & (g192)) + ((!sk[79]) & (!g168) & (!g173) & (g180) & (g183) & (!g192)) + ((!sk[79]) & (!g168) & (!g173) & (g180) & (g183) & (g192)) + ((!sk[79]) & (!g168) & (g173) & (!g180) & (!g183) & (!g192)) + ((!sk[79]) & (!g168) & (g173) & (!g180) & (!g183) & (g192)) + ((!sk[79]) & (!g168) & (g173) & (!g180) & (g183) & (!g192)) + ((!sk[79]) & (!g168) & (g173) & (!g180) & (g183) & (g192)) + ((!sk[79]) & (!g168) & (g173) & (g180) & (!g183) & (!g192)) + ((!sk[79]) & (!g168) & (g173) & (g180) & (!g183) & (g192)) + ((!sk[79]) & (!g168) & (g173) & (g180) & (g183) & (!g192)) + ((!sk[79]) & (!g168) & (g173) & (g180) & (g183) & (g192)) + ((!sk[79]) & (g168) & (!g173) & (!g180) & (g183) & (!g192)) + ((!sk[79]) & (g168) & (!g173) & (!g180) & (g183) & (g192)) + ((!sk[79]) & (g168) & (!g173) & (g180) & (!g183) & (!g192)) + ((!sk[79]) & (g168) & (!g173) & (g180) & (!g183) & (g192)) + ((!sk[79]) & (g168) & (!g173) & (g180) & (g183) & (!g192)) + ((!sk[79]) & (g168) & (!g173) & (g180) & (g183) & (g192)) + ((!sk[79]) & (g168) & (g173) & (!g180) & (!g183) & (!g192)) + ((!sk[79]) & (g168) & (g173) & (!g180) & (!g183) & (g192)) + ((!sk[79]) & (g168) & (g173) & (!g180) & (g183) & (!g192)) + ((!sk[79]) & (g168) & (g173) & (!g180) & (g183) & (g192)) + ((!sk[79]) & (g168) & (g173) & (g180) & (!g183) & (!g192)) + ((!sk[79]) & (g168) & (g173) & (g180) & (!g183) & (g192)) + ((!sk[79]) & (g168) & (g173) & (g180) & (g183) & (!g192)) + ((!sk[79]) & (g168) & (g173) & (g180) & (g183) & (g192)) + ((sk[79]) & (g168) & (g173) & (g180) & (g183) & (g192)));
	assign g326 = (((!g85) & (!sk[80]) & (!g124) & (g86)) + ((!g85) & (!sk[80]) & (g124) & (g86)) + ((!g85) & (sk[80]) & (!g124) & (!g86)) + ((g85) & (!sk[80]) & (!g124) & (!g86)) + ((g85) & (!sk[80]) & (!g124) & (g86)) + ((g85) & (!sk[80]) & (g124) & (!g86)) + ((g85) & (!sk[80]) & (g124) & (g86)));
	assign g327 = (((!g70) & (!g241) & (!sk[81]) & (g32)) + ((!g70) & (!g241) & (sk[81]) & (!g32)) + ((!g70) & (!g241) & (sk[81]) & (g32)) + ((!g70) & (g241) & (!sk[81]) & (g32)) + ((g70) & (!g241) & (!sk[81]) & (!g32)) + ((g70) & (!g241) & (!sk[81]) & (g32)) + ((g70) & (!g241) & (sk[81]) & (!g32)) + ((g70) & (g241) & (!sk[81]) & (!g32)) + ((g70) & (g241) & (!sk[81]) & (g32)));
	assign g328 = (((!g16) & (!sk[82]) & (!g25) & (g288)) + ((!g16) & (!sk[82]) & (g25) & (g288)) + ((!g16) & (sk[82]) & (!g25) & (!g288)) + ((!g16) & (sk[82]) & (g25) & (!g288)) + ((g16) & (!sk[82]) & (!g25) & (!g288)) + ((g16) & (!sk[82]) & (!g25) & (g288)) + ((g16) & (!sk[82]) & (g25) & (!g288)) + ((g16) & (!sk[82]) & (g25) & (g288)) + ((g16) & (sk[82]) & (!g25) & (!g288)));
	assign g329 = (((!g38) & (!g49) & (!g99) & (!g71) & (!g41) & (!g233)) + ((!g38) & (!g49) & (!g99) & (!g71) & (g41) & (!g233)) + ((!g38) & (!g49) & (!g99) & (g71) & (!g41) & (!g233)) + ((!g38) & (!g49) & (g99) & (!g71) & (!g41) & (!g233)) + ((!g38) & (!g49) & (g99) & (g71) & (!g41) & (!g233)) + ((!g38) & (g49) & (!g99) & (!g71) & (!g41) & (!g233)) + ((!g38) & (g49) & (!g99) & (!g71) & (g41) & (!g233)) + ((!g38) & (g49) & (!g99) & (g71) & (!g41) & (!g233)) + ((g38) & (!g49) & (!g99) & (!g71) & (!g41) & (!g233)) + ((g38) & (!g49) & (!g99) & (!g71) & (g41) & (!g233)) + ((g38) & (!g49) & (g99) & (!g71) & (!g41) & (!g233)) + ((g38) & (g49) & (!g99) & (!g71) & (!g41) & (!g233)) + ((g38) & (g49) & (!g99) & (!g71) & (g41) & (!g233)));
	assign g330 = (((g326) & (g327) & (g134) & (g138) & (g328) & (g329)));
	assign g331 = (((!g70) & (!g17) & (!sk[85]) & (g71) & (!g20)) + ((!g70) & (!g17) & (!sk[85]) & (g71) & (g20)) + ((!g70) & (g17) & (!sk[85]) & (g71) & (!g20)) + ((!g70) & (g17) & (!sk[85]) & (g71) & (g20)) + ((!g70) & (g17) & (sk[85]) & (g71) & (!g20)) + ((!g70) & (g17) & (sk[85]) & (g71) & (g20)) + ((g70) & (!g17) & (!sk[85]) & (!g71) & (!g20)) + ((g70) & (!g17) & (!sk[85]) & (!g71) & (g20)) + ((g70) & (!g17) & (!sk[85]) & (g71) & (!g20)) + ((g70) & (!g17) & (!sk[85]) & (g71) & (g20)) + ((g70) & (!g17) & (sk[85]) & (!g71) & (g20)) + ((g70) & (!g17) & (sk[85]) & (g71) & (g20)) + ((g70) & (g17) & (!sk[85]) & (!g71) & (!g20)) + ((g70) & (g17) & (!sk[85]) & (!g71) & (g20)) + ((g70) & (g17) & (!sk[85]) & (g71) & (!g20)) + ((g70) & (g17) & (!sk[85]) & (g71) & (g20)) + ((g70) & (g17) & (sk[85]) & (!g71) & (g20)) + ((g70) & (g17) & (sk[85]) & (g71) & (!g20)) + ((g70) & (g17) & (sk[85]) & (g71) & (g20)));
	assign g332 = (((!sk[86]) & (!g70) & (!g16) & (g40) & (!g272)) + ((!sk[86]) & (!g70) & (!g16) & (g40) & (g272)) + ((!sk[86]) & (!g70) & (g16) & (g40) & (!g272)) + ((!sk[86]) & (!g70) & (g16) & (g40) & (g272)) + ((!sk[86]) & (g70) & (!g16) & (!g40) & (!g272)) + ((!sk[86]) & (g70) & (!g16) & (!g40) & (g272)) + ((!sk[86]) & (g70) & (!g16) & (g40) & (!g272)) + ((!sk[86]) & (g70) & (!g16) & (g40) & (g272)) + ((!sk[86]) & (g70) & (g16) & (!g40) & (!g272)) + ((!sk[86]) & (g70) & (g16) & (!g40) & (g272)) + ((!sk[86]) & (g70) & (g16) & (g40) & (!g272)) + ((!sk[86]) & (g70) & (g16) & (g40) & (g272)) + ((sk[86]) & (!g70) & (!g16) & (!g40) & (!g272)) + ((sk[86]) & (!g70) & (!g16) & (g40) & (!g272)) + ((sk[86]) & (!g70) & (g16) & (!g40) & (!g272)) + ((sk[86]) & (g70) & (!g16) & (!g40) & (!g272)) + ((sk[86]) & (g70) & (g16) & (!g40) & (!g272)));
	assign g333 = (((!g331) & (!g260) & (!sk[87]) & (g143) & (!g332)) + ((!g331) & (!g260) & (!sk[87]) & (g143) & (g332)) + ((!g331) & (g260) & (!sk[87]) & (g143) & (!g332)) + ((!g331) & (g260) & (!sk[87]) & (g143) & (g332)) + ((!g331) & (g260) & (sk[87]) & (g143) & (g332)) + ((g331) & (!g260) & (!sk[87]) & (!g143) & (!g332)) + ((g331) & (!g260) & (!sk[87]) & (!g143) & (g332)) + ((g331) & (!g260) & (!sk[87]) & (g143) & (!g332)) + ((g331) & (!g260) & (!sk[87]) & (g143) & (g332)) + ((g331) & (g260) & (!sk[87]) & (!g143) & (!g332)) + ((g331) & (g260) & (!sk[87]) & (!g143) & (g332)) + ((g331) & (g260) & (!sk[87]) & (g143) & (!g332)) + ((g331) & (g260) & (!sk[87]) & (g143) & (g332)));
	assign g334 = (((!sk[88]) & (!g70) & (!g163) & (g58)) + ((!sk[88]) & (!g70) & (g163) & (g58)) + ((!sk[88]) & (g70) & (!g163) & (!g58)) + ((!sk[88]) & (g70) & (!g163) & (g58)) + ((!sk[88]) & (g70) & (g163) & (!g58)) + ((!sk[88]) & (g70) & (g163) & (g58)) + ((sk[88]) & (!g70) & (!g163) & (!g58)) + ((sk[88]) & (!g70) & (!g163) & (g58)) + ((sk[88]) & (g70) & (!g163) & (!g58)));
	assign g335 = (((!sk[89]) & (!g71) & (!g20) & (g13)) + ((!sk[89]) & (!g71) & (g20) & (g13)) + ((!sk[89]) & (g71) & (!g20) & (!g13)) + ((!sk[89]) & (g71) & (!g20) & (g13)) + ((!sk[89]) & (g71) & (g20) & (!g13)) + ((!sk[89]) & (g71) & (g20) & (g13)) + ((sk[89]) & (!g71) & (!g20) & (!g13)) + ((sk[89]) & (!g71) & (g20) & (!g13)) + ((sk[89]) & (g71) & (!g20) & (!g13)));
	assign g336 = (((!g9) & (!g62) & (!g71) & (!g18) & (!g25) & (!g66)) + ((!g9) & (!g62) & (!g71) & (!g18) & (!g25) & (g66)) + ((!g9) & (!g62) & (!g71) & (!g18) & (g25) & (!g66)) + ((!g9) & (!g62) & (!g71) & (!g18) & (g25) & (g66)) + ((!g9) & (!g62) & (!g71) & (g18) & (!g25) & (!g66)) + ((!g9) & (!g62) & (!g71) & (g18) & (!g25) & (g66)) + ((!g9) & (!g62) & (!g71) & (g18) & (g25) & (!g66)) + ((!g9) & (!g62) & (!g71) & (g18) & (g25) & (g66)) + ((!g9) & (!g62) & (g71) & (!g18) & (!g25) & (!g66)) + ((!g9) & (!g62) & (g71) & (!g18) & (!g25) & (g66)) + ((!g9) & (!g62) & (g71) & (g18) & (!g25) & (!g66)) + ((!g9) & (!g62) & (g71) & (g18) & (!g25) & (g66)) + ((!g9) & (g62) & (!g71) & (!g18) & (!g25) & (!g66)) + ((!g9) & (g62) & (!g71) & (!g18) & (g25) & (!g66)) + ((!g9) & (g62) & (g71) & (!g18) & (!g25) & (!g66)) + ((g9) & (!g62) & (!g71) & (!g18) & (!g25) & (!g66)) + ((g9) & (!g62) & (!g71) & (!g18) & (!g25) & (g66)) + ((g9) & (!g62) & (!g71) & (g18) & (!g25) & (!g66)) + ((g9) & (!g62) & (!g71) & (g18) & (!g25) & (g66)) + ((g9) & (!g62) & (g71) & (!g18) & (!g25) & (!g66)) + ((g9) & (!g62) & (g71) & (!g18) & (!g25) & (g66)) + ((g9) & (!g62) & (g71) & (g18) & (!g25) & (!g66)) + ((g9) & (!g62) & (g71) & (g18) & (!g25) & (g66)) + ((g9) & (g62) & (!g71) & (!g18) & (!g25) & (!g66)) + ((g9) & (g62) & (g71) & (!g18) & (!g25) & (!g66)));
	assign g337 = (((!g99) & (!g83) & (!g25) & (!g84) & (sk[91]) & (!g152)) + ((!g99) & (!g83) & (!g25) & (g84) & (!sk[91]) & (!g152)) + ((!g99) & (!g83) & (!g25) & (g84) & (!sk[91]) & (g152)) + ((!g99) & (!g83) & (g25) & (!g84) & (sk[91]) & (!g152)) + ((!g99) & (!g83) & (g25) & (g84) & (!sk[91]) & (!g152)) + ((!g99) & (!g83) & (g25) & (g84) & (!sk[91]) & (g152)) + ((!g99) & (g83) & (!g25) & (!g84) & (!sk[91]) & (!g152)) + ((!g99) & (g83) & (!g25) & (!g84) & (!sk[91]) & (g152)) + ((!g99) & (g83) & (!g25) & (g84) & (!sk[91]) & (!g152)) + ((!g99) & (g83) & (!g25) & (g84) & (!sk[91]) & (g152)) + ((!g99) & (g83) & (g25) & (!g84) & (!sk[91]) & (!g152)) + ((!g99) & (g83) & (g25) & (!g84) & (!sk[91]) & (g152)) + ((!g99) & (g83) & (g25) & (g84) & (!sk[91]) & (!g152)) + ((!g99) & (g83) & (g25) & (g84) & (!sk[91]) & (g152)) + ((g99) & (!g83) & (!g25) & (!g84) & (sk[91]) & (!g152)) + ((g99) & (!g83) & (!g25) & (g84) & (!sk[91]) & (!g152)) + ((g99) & (!g83) & (!g25) & (g84) & (!sk[91]) & (g152)) + ((g99) & (!g83) & (g25) & (!g84) & (!sk[91]) & (!g152)) + ((g99) & (!g83) & (g25) & (!g84) & (!sk[91]) & (g152)) + ((g99) & (!g83) & (g25) & (g84) & (!sk[91]) & (!g152)) + ((g99) & (!g83) & (g25) & (g84) & (!sk[91]) & (g152)) + ((g99) & (g83) & (!g25) & (!g84) & (!sk[91]) & (!g152)) + ((g99) & (g83) & (!g25) & (!g84) & (!sk[91]) & (g152)) + ((g99) & (g83) & (!g25) & (g84) & (!sk[91]) & (!g152)) + ((g99) & (g83) & (!g25) & (g84) & (!sk[91]) & (g152)) + ((g99) & (g83) & (g25) & (!g84) & (!sk[91]) & (!g152)) + ((g99) & (g83) & (g25) & (!g84) & (!sk[91]) & (g152)) + ((g99) & (g83) & (g25) & (g84) & (!sk[91]) & (!g152)) + ((g99) & (g83) & (g25) & (g84) & (!sk[91]) & (g152)));
	assign g338 = (((!g9) & (!g10) & (!g27) & (!g105) & (!g275) & (!g150)) + ((!g9) & (!g10) & (g27) & (!g105) & (!g275) & (!g150)) + ((!g9) & (g10) & (!g27) & (!g105) & (!g275) & (!g150)) + ((!g9) & (g10) & (g27) & (!g105) & (!g275) & (!g150)) + ((g9) & (!g10) & (!g27) & (!g105) & (!g275) & (!g150)));
	assign g339 = (((g237) & (g334) & (g335) & (g336) & (g337) & (g338)));
	assign g340 = (((!g70) & (!sk[94]) & (!g12) & (g18) & (!g104)) + ((!g70) & (!sk[94]) & (!g12) & (g18) & (g104)) + ((!g70) & (!sk[94]) & (g12) & (g18) & (!g104)) + ((!g70) & (!sk[94]) & (g12) & (g18) & (g104)) + ((!g70) & (sk[94]) & (!g12) & (g18) & (g104)) + ((!g70) & (sk[94]) & (g12) & (g18) & (g104)) + ((g70) & (!sk[94]) & (!g12) & (!g18) & (!g104)) + ((g70) & (!sk[94]) & (!g12) & (!g18) & (g104)) + ((g70) & (!sk[94]) & (!g12) & (g18) & (!g104)) + ((g70) & (!sk[94]) & (!g12) & (g18) & (g104)) + ((g70) & (!sk[94]) & (g12) & (!g18) & (!g104)) + ((g70) & (!sk[94]) & (g12) & (!g18) & (g104)) + ((g70) & (!sk[94]) & (g12) & (g18) & (!g104)) + ((g70) & (!sk[94]) & (g12) & (g18) & (g104)) + ((g70) & (sk[94]) & (!g12) & (g18) & (g104)) + ((g70) & (sk[94]) & (g12) & (!g18) & (!g104)) + ((g70) & (sk[94]) & (g12) & (!g18) & (g104)) + ((g70) & (sk[94]) & (g12) & (g18) & (!g104)) + ((g70) & (sk[94]) & (g12) & (g18) & (g104)));
	assign g341 = (((!g57) & (!g71) & (!g18) & (!g32) & (!g187) & (!g207)) + ((!g57) & (!g71) & (!g18) & (g32) & (!g187) & (!g207)) + ((!g57) & (!g71) & (g18) & (!g32) & (!g187) & (!g207)) + ((!g57) & (!g71) & (g18) & (g32) & (!g187) & (!g207)) + ((!g57) & (g71) & (!g18) & (!g32) & (!g187) & (!g207)) + ((g57) & (!g71) & (!g18) & (!g32) & (!g187) & (!g207)) + ((g57) & (!g71) & (g18) & (!g32) & (!g187) & (!g207)) + ((g57) & (g71) & (!g18) & (!g32) & (!g187) & (!g207)));
	assign g342 = (((!g340) & (!sk[96]) & (g341)) + ((!g340) & (sk[96]) & (g341)) + ((g340) & (!sk[96]) & (g341)));
	assign g343 = (((!g330) & (!sk[97]) & (!g333) & (g339) & (!g342)) + ((!g330) & (!sk[97]) & (!g333) & (g339) & (g342)) + ((!g330) & (!sk[97]) & (g333) & (g339) & (!g342)) + ((!g330) & (!sk[97]) & (g333) & (g339) & (g342)) + ((g330) & (!sk[97]) & (!g333) & (!g339) & (!g342)) + ((g330) & (!sk[97]) & (!g333) & (!g339) & (g342)) + ((g330) & (!sk[97]) & (!g333) & (g339) & (!g342)) + ((g330) & (!sk[97]) & (!g333) & (g339) & (g342)) + ((g330) & (!sk[97]) & (g333) & (!g339) & (!g342)) + ((g330) & (!sk[97]) & (g333) & (!g339) & (g342)) + ((g330) & (!sk[97]) & (g333) & (g339) & (!g342)) + ((g330) & (!sk[97]) & (g333) & (g339) & (g342)) + ((g330) & (sk[97]) & (g333) & (g339) & (g342)));
	assign g344 = (((!g325) & (!sk[98]) & (g343)) + ((g325) & (!sk[98]) & (g343)) + ((g325) & (sk[98]) & (g343)));
	assign g345 = (((!g104) & (!sk[99]) & (!g40) & (g19)) + ((!g104) & (!sk[99]) & (g40) & (g19)) + ((!g104) & (sk[99]) & (!g40) & (!g19)) + ((!g104) & (sk[99]) & (g40) & (!g19)) + ((g104) & (!sk[99]) & (!g40) & (!g19)) + ((g104) & (!sk[99]) & (!g40) & (g19)) + ((g104) & (!sk[99]) & (g40) & (!g19)) + ((g104) & (!sk[99]) & (g40) & (g19)) + ((g104) & (sk[99]) & (!g40) & (!g19)));
	assign g346 = (((!g38) & (!g62) & (!sk[100]) & (g127) & (!g87)) + ((!g38) & (!g62) & (!sk[100]) & (g127) & (g87)) + ((!g38) & (!g62) & (sk[100]) & (!g127) & (!g87)) + ((!g38) & (g62) & (!sk[100]) & (g127) & (!g87)) + ((!g38) & (g62) & (!sk[100]) & (g127) & (g87)) + ((!g38) & (g62) & (sk[100]) & (!g127) & (!g87)) + ((g38) & (!g62) & (!sk[100]) & (!g127) & (!g87)) + ((g38) & (!g62) & (!sk[100]) & (!g127) & (g87)) + ((g38) & (!g62) & (!sk[100]) & (g127) & (!g87)) + ((g38) & (!g62) & (!sk[100]) & (g127) & (g87)) + ((g38) & (!g62) & (sk[100]) & (!g127) & (!g87)) + ((g38) & (g62) & (!sk[100]) & (!g127) & (!g87)) + ((g38) & (g62) & (!sk[100]) & (!g127) & (g87)) + ((g38) & (g62) & (!sk[100]) & (g127) & (!g87)) + ((g38) & (g62) & (!sk[100]) & (g127) & (g87)));
	assign g347 = (((g345) & (g330) & (g333) & (g339) & (g342) & (g346)));
	assign g348 = (((!g9) & (!g16) & (!g40) & (sk[102]) & (!g80)) + ((!g9) & (!g16) & (g40) & (!sk[102]) & (!g80)) + ((!g9) & (!g16) & (g40) & (!sk[102]) & (g80)) + ((!g9) & (!g16) & (g40) & (sk[102]) & (!g80)) + ((!g9) & (g16) & (!g40) & (sk[102]) & (!g80)) + ((!g9) & (g16) & (g40) & (!sk[102]) & (!g80)) + ((!g9) & (g16) & (g40) & (!sk[102]) & (g80)) + ((g9) & (!g16) & (!g40) & (!sk[102]) & (!g80)) + ((g9) & (!g16) & (!g40) & (!sk[102]) & (g80)) + ((g9) & (!g16) & (!g40) & (sk[102]) & (!g80)) + ((g9) & (!g16) & (g40) & (!sk[102]) & (!g80)) + ((g9) & (!g16) & (g40) & (!sk[102]) & (g80)) + ((g9) & (g16) & (!g40) & (!sk[102]) & (!g80)) + ((g9) & (g16) & (!g40) & (!sk[102]) & (g80)) + ((g9) & (g16) & (!g40) & (sk[102]) & (!g80)) + ((g9) & (g16) & (g40) & (!sk[102]) & (!g80)) + ((g9) & (g16) & (g40) & (!sk[102]) & (g80)));
	assign g349 = (((!g153) & (!sk[103]) & (g177)) + ((!g153) & (sk[103]) & (!g177)) + ((g153) & (!sk[103]) & (g177)));
	assign g350 = (((!g70) & (!g16) & (!g41) & (!g13) & (!g171) & (!g87)) + ((!g70) & (!g16) & (g41) & (!g13) & (!g171) & (!g87)) + ((!g70) & (g16) & (!g41) & (!g13) & (!g171) & (!g87)) + ((g70) & (!g16) & (!g41) & (!g13) & (!g171) & (!g87)) + ((g70) & (g16) & (!g41) & (!g13) & (!g171) & (!g87)));
	assign g351 = (((!g70) & (!g62) & (!sk[105]) & (g18) & (!g91)) + ((!g70) & (!g62) & (!sk[105]) & (g18) & (g91)) + ((!g70) & (g62) & (!sk[105]) & (g18) & (!g91)) + ((!g70) & (g62) & (!sk[105]) & (g18) & (g91)) + ((!g70) & (g62) & (sk[105]) & (!g18) & (g91)) + ((!g70) & (g62) & (sk[105]) & (g18) & (g91)) + ((g70) & (!g62) & (!sk[105]) & (!g18) & (!g91)) + ((g70) & (!g62) & (!sk[105]) & (!g18) & (g91)) + ((g70) & (!g62) & (!sk[105]) & (g18) & (!g91)) + ((g70) & (!g62) & (!sk[105]) & (g18) & (g91)) + ((g70) & (!g62) & (sk[105]) & (g18) & (!g91)) + ((g70) & (!g62) & (sk[105]) & (g18) & (g91)) + ((g70) & (g62) & (!sk[105]) & (!g18) & (!g91)) + ((g70) & (g62) & (!sk[105]) & (!g18) & (g91)) + ((g70) & (g62) & (!sk[105]) & (g18) & (!g91)) + ((g70) & (g62) & (!sk[105]) & (g18) & (g91)) + ((g70) & (g62) & (sk[105]) & (!g18) & (g91)) + ((g70) & (g62) & (sk[105]) & (g18) & (!g91)) + ((g70) & (g62) & (sk[105]) & (g18) & (g91)));
	assign g352 = (((g348) & (!g232) & (g349) & (g157) & (g350) & (!g351)));
	assign g353 = (((!g112) & (!g113) & (!g97) & (g98) & (!g16) & (g62)) + ((!g112) & (!g113) & (!g97) & (g98) & (g16) & (g62)) + ((!g112) & (!g113) & (g97) & (!g98) & (!g16) & (g62)) + ((!g112) & (!g113) & (g97) & (!g98) & (g16) & (g62)) + ((!g112) & (g113) & (g97) & (!g98) & (g16) & (!g62)) + ((!g112) & (g113) & (g97) & (!g98) & (g16) & (g62)) + ((g112) & (!g113) & (!g97) & (g98) & (!g16) & (g62)) + ((g112) & (!g113) & (!g97) & (g98) & (g16) & (g62)) + ((g112) & (g113) & (!g97) & (!g98) & (g16) & (!g62)) + ((g112) & (g113) & (!g97) & (!g98) & (g16) & (g62)) + ((g112) & (g113) & (g97) & (g98) & (g16) & (!g62)) + ((g112) & (g113) & (g97) & (g98) & (g16) & (g62)));
	assign g354 = (((!ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g49)) + ((!ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g49)) + ((ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g49)) + ((ax22x) & (!ax21x) & (g6) & (!ax20x) & (!g8) & (g49)));
	assign g355 = (((!g238) & (!g241) & (!g50) & (!g354) & (!g147) & (!g51)));
	assign g356 = (((!g38) & (!g9) & (!g32) & (!g60) & (!g95) & (!g190)) + ((!g38) & (!g9) & (g32) & (!g60) & (!g95) & (!g190)) + ((!g38) & (g9) & (!g32) & (!g60) & (!g95) & (!g190)) + ((g38) & (!g9) & (!g32) & (!g60) & (!g95) & (!g190)) + ((g38) & (!g9) & (g32) & (!g60) & (!g95) & (!g190)));
	assign g357 = (((g298) & (!g340) & (g341) & (!g353) & (g355) & (g356)));
	assign g358 = (((!g128) & (!g97) & (!sk[112]) & (g71) & (!g127)) + ((!g128) & (!g97) & (!sk[112]) & (g71) & (g127)) + ((!g128) & (!g97) & (sk[112]) & (!g71) & (!g127)) + ((!g128) & (!g97) & (sk[112]) & (g71) & (!g127)) + ((!g128) & (g97) & (!sk[112]) & (g71) & (!g127)) + ((!g128) & (g97) & (!sk[112]) & (g71) & (g127)) + ((!g128) & (g97) & (sk[112]) & (!g71) & (!g127)) + ((!g128) & (g97) & (sk[112]) & (g71) & (!g127)) + ((g128) & (!g97) & (!sk[112]) & (!g71) & (!g127)) + ((g128) & (!g97) & (!sk[112]) & (!g71) & (g127)) + ((g128) & (!g97) & (!sk[112]) & (g71) & (!g127)) + ((g128) & (!g97) & (!sk[112]) & (g71) & (g127)) + ((g128) & (!g97) & (sk[112]) & (!g71) & (!g127)) + ((g128) & (g97) & (!sk[112]) & (!g71) & (!g127)) + ((g128) & (g97) & (!sk[112]) & (!g71) & (g127)) + ((g128) & (g97) & (!sk[112]) & (g71) & (!g127)) + ((g128) & (g97) & (!sk[112]) & (g71) & (g127)) + ((g128) & (g97) & (sk[112]) & (!g71) & (!g127)) + ((g128) & (g97) & (sk[112]) & (g71) & (!g127)));
	assign g359 = (((!ax22x) & (!ax21x) & (!g6) & (!ax20x) & (!g8) & (g91)) + ((!ax22x) & (!ax21x) & (g6) & (ax20x) & (!g8) & (g91)) + ((ax22x) & (ax21x) & (!g6) & (ax20x) & (!g8) & (g91)) + ((ax22x) & (ax21x) & (g6) & (ax20x) & (!g8) & (g91)));
	assign g360 = (((!sk[114]) & (!g17) & (!g99) & (!g18) & (g40) & (!g66)) + ((!sk[114]) & (!g17) & (!g99) & (!g18) & (g40) & (g66)) + ((!sk[114]) & (!g17) & (!g99) & (g18) & (g40) & (!g66)) + ((!sk[114]) & (!g17) & (!g99) & (g18) & (g40) & (g66)) + ((!sk[114]) & (!g17) & (g99) & (!g18) & (!g40) & (!g66)) + ((!sk[114]) & (!g17) & (g99) & (!g18) & (!g40) & (g66)) + ((!sk[114]) & (!g17) & (g99) & (!g18) & (g40) & (!g66)) + ((!sk[114]) & (!g17) & (g99) & (!g18) & (g40) & (g66)) + ((!sk[114]) & (!g17) & (g99) & (g18) & (!g40) & (!g66)) + ((!sk[114]) & (!g17) & (g99) & (g18) & (!g40) & (g66)) + ((!sk[114]) & (!g17) & (g99) & (g18) & (g40) & (!g66)) + ((!sk[114]) & (!g17) & (g99) & (g18) & (g40) & (g66)) + ((!sk[114]) & (g17) & (!g99) & (!g18) & (g40) & (!g66)) + ((!sk[114]) & (g17) & (!g99) & (!g18) & (g40) & (g66)) + ((!sk[114]) & (g17) & (!g99) & (g18) & (!g40) & (!g66)) + ((!sk[114]) & (g17) & (!g99) & (g18) & (!g40) & (g66)) + ((!sk[114]) & (g17) & (!g99) & (g18) & (g40) & (!g66)) + ((!sk[114]) & (g17) & (!g99) & (g18) & (g40) & (g66)) + ((!sk[114]) & (g17) & (g99) & (!g18) & (!g40) & (!g66)) + ((!sk[114]) & (g17) & (g99) & (!g18) & (!g40) & (g66)) + ((!sk[114]) & (g17) & (g99) & (!g18) & (g40) & (!g66)) + ((!sk[114]) & (g17) & (g99) & (!g18) & (g40) & (g66)) + ((!sk[114]) & (g17) & (g99) & (g18) & (!g40) & (!g66)) + ((!sk[114]) & (g17) & (g99) & (g18) & (!g40) & (g66)) + ((!sk[114]) & (g17) & (g99) & (g18) & (g40) & (!g66)) + ((!sk[114]) & (g17) & (g99) & (g18) & (g40) & (g66)) + ((sk[114]) & (!g17) & (g99) & (!g18) & (!g40) & (g66)) + ((sk[114]) & (!g17) & (g99) & (!g18) & (g40) & (!g66)) + ((sk[114]) & (!g17) & (g99) & (!g18) & (g40) & (g66)) + ((sk[114]) & (!g17) & (g99) & (g18) & (!g40) & (!g66)) + ((sk[114]) & (!g17) & (g99) & (g18) & (!g40) & (g66)) + ((sk[114]) & (!g17) & (g99) & (g18) & (g40) & (!g66)) + ((sk[114]) & (!g17) & (g99) & (g18) & (g40) & (g66)) + ((sk[114]) & (g17) & (g99) & (!g18) & (!g40) & (!g66)) + ((sk[114]) & (g17) & (g99) & (!g18) & (!g40) & (g66)) + ((sk[114]) & (g17) & (g99) & (!g18) & (g40) & (!g66)) + ((sk[114]) & (g17) & (g99) & (!g18) & (g40) & (g66)) + ((sk[114]) & (g17) & (g99) & (g18) & (!g40) & (!g66)) + ((sk[114]) & (g17) & (g99) & (g18) & (!g40) & (g66)) + ((sk[114]) & (g17) & (g99) & (g18) & (g40) & (!g66)) + ((sk[114]) & (g17) & (g99) & (g18) & (g40) & (g66)));
	assign g361 = (((!g54) & (!g297) & (g358) & (!g203) & (!g359) & (!g360)));
	assign g362 = (((!g70) & (!g17) & (!g184) & (!g104) & (!g40) & (!g41)) + ((!g70) & (!g17) & (!g184) & (!g104) & (!g40) & (g41)) + ((!g70) & (!g17) & (!g184) & (!g104) & (g40) & (!g41)) + ((!g70) & (!g17) & (!g184) & (!g104) & (g40) & (g41)) + ((!g70) & (!g17) & (!g184) & (g104) & (!g40) & (!g41)) + ((!g70) & (g17) & (!g184) & (!g104) & (!g40) & (!g41)) + ((!g70) & (g17) & (!g184) & (!g104) & (!g40) & (g41)) + ((!g70) & (g17) & (!g184) & (!g104) & (g40) & (!g41)) + ((!g70) & (g17) & (!g184) & (!g104) & (g40) & (g41)) + ((!g70) & (g17) & (!g184) & (g104) & (!g40) & (!g41)) + ((g70) & (!g17) & (!g184) & (!g104) & (!g40) & (!g41)) + ((g70) & (!g17) & (!g184) & (!g104) & (!g40) & (g41)) + ((g70) & (!g17) & (!g184) & (g104) & (!g40) & (!g41)));
	assign g363 = (((!sk[117]) & (!g9) & (!g58) & (g194)) + ((!sk[117]) & (!g9) & (g58) & (g194)) + ((!sk[117]) & (g9) & (!g58) & (!g194)) + ((!sk[117]) & (g9) & (!g58) & (g194)) + ((!sk[117]) & (g9) & (g58) & (!g194)) + ((!sk[117]) & (g9) & (g58) & (g194)) + ((sk[117]) & (!g9) & (!g58) & (!g194)) + ((sk[117]) & (!g9) & (g58) & (!g194)) + ((sk[117]) & (g9) & (!g58) & (!g194)));
	assign g364 = (((!g85) & (!g29) & (!sk[118]) & (!g86) & (g254) & (!g363)) + ((!g85) & (!g29) & (!sk[118]) & (!g86) & (g254) & (g363)) + ((!g85) & (!g29) & (!sk[118]) & (g86) & (g254) & (!g363)) + ((!g85) & (!g29) & (!sk[118]) & (g86) & (g254) & (g363)) + ((!g85) & (!g29) & (sk[118]) & (!g86) & (!g254) & (g363)) + ((!g85) & (g29) & (!sk[118]) & (!g86) & (!g254) & (!g363)) + ((!g85) & (g29) & (!sk[118]) & (!g86) & (!g254) & (g363)) + ((!g85) & (g29) & (!sk[118]) & (!g86) & (g254) & (!g363)) + ((!g85) & (g29) & (!sk[118]) & (!g86) & (g254) & (g363)) + ((!g85) & (g29) & (!sk[118]) & (g86) & (!g254) & (!g363)) + ((!g85) & (g29) & (!sk[118]) & (g86) & (!g254) & (g363)) + ((!g85) & (g29) & (!sk[118]) & (g86) & (g254) & (!g363)) + ((!g85) & (g29) & (!sk[118]) & (g86) & (g254) & (g363)) + ((g85) & (!g29) & (!sk[118]) & (!g86) & (g254) & (!g363)) + ((g85) & (!g29) & (!sk[118]) & (!g86) & (g254) & (g363)) + ((g85) & (!g29) & (!sk[118]) & (g86) & (!g254) & (!g363)) + ((g85) & (!g29) & (!sk[118]) & (g86) & (!g254) & (g363)) + ((g85) & (!g29) & (!sk[118]) & (g86) & (g254) & (!g363)) + ((g85) & (!g29) & (!sk[118]) & (g86) & (g254) & (g363)) + ((g85) & (g29) & (!sk[118]) & (!g86) & (!g254) & (!g363)) + ((g85) & (g29) & (!sk[118]) & (!g86) & (!g254) & (g363)) + ((g85) & (g29) & (!sk[118]) & (!g86) & (g254) & (!g363)) + ((g85) & (g29) & (!sk[118]) & (!g86) & (g254) & (g363)) + ((g85) & (g29) & (!sk[118]) & (g86) & (!g254) & (!g363)) + ((g85) & (g29) & (!sk[118]) & (g86) & (!g254) & (g363)) + ((g85) & (g29) & (!sk[118]) & (g86) & (g254) & (!g363)) + ((g85) & (g29) & (!sk[118]) & (g86) & (g254) & (g363)));
	assign g365 = (((!g275) & (g352) & (g357) & (g361) & (g362) & (g364)));
	assign g366 = (((!sk[120]) & (!g196) & (!g347) & (g365)) + ((!sk[120]) & (!g196) & (g347) & (g365)) + ((!sk[120]) & (g196) & (!g347) & (!g365)) + ((!sk[120]) & (g196) & (!g347) & (g365)) + ((!sk[120]) & (g196) & (g347) & (!g365)) + ((!sk[120]) & (g196) & (g347) & (g365)) + ((sk[120]) & (!g196) & (!g347) & (g365)));
	assign g367 = (((!sk[121]) & (!ax22x) & (!g3) & (ax6x)) + ((!sk[121]) & (!ax22x) & (g3) & (ax6x)) + ((!sk[121]) & (ax22x) & (!g3) & (!ax6x)) + ((!sk[121]) & (ax22x) & (!g3) & (ax6x)) + ((!sk[121]) & (ax22x) & (g3) & (!ax6x)) + ((!sk[121]) & (ax22x) & (g3) & (ax6x)) + ((sk[121]) & (!ax22x) & (!g3) & (!ax6x)) + ((sk[121]) & (!ax22x) & (g3) & (ax6x)) + ((sk[121]) & (ax22x) & (!g3) & (ax6x)) + ((sk[121]) & (ax22x) & (g3) & (ax6x)));
	assign g368 = (((!g45) & (!sk[122]) & (!g68) & (g367)) + ((!g45) & (!sk[122]) & (g68) & (g367)) + ((!g45) & (sk[122]) & (!g68) & (g367)) + ((!g45) & (sk[122]) & (g68) & (g367)) + ((g45) & (!sk[122]) & (!g68) & (!g367)) + ((g45) & (!sk[122]) & (!g68) & (g367)) + ((g45) & (!sk[122]) & (g68) & (!g367)) + ((g45) & (!sk[122]) & (g68) & (g367)) + ((g45) & (sk[122]) & (!g68) & (g367)));
	assign g369 = (((!sk[123]) & (!g323) & (!g324) & (!g344) & (g366) & (!g368)) + ((!sk[123]) & (!g323) & (!g324) & (!g344) & (g366) & (g368)) + ((!sk[123]) & (!g323) & (!g324) & (g344) & (g366) & (!g368)) + ((!sk[123]) & (!g323) & (!g324) & (g344) & (g366) & (g368)) + ((!sk[123]) & (!g323) & (g324) & (!g344) & (!g366) & (!g368)) + ((!sk[123]) & (!g323) & (g324) & (!g344) & (!g366) & (g368)) + ((!sk[123]) & (!g323) & (g324) & (!g344) & (g366) & (!g368)) + ((!sk[123]) & (!g323) & (g324) & (!g344) & (g366) & (g368)) + ((!sk[123]) & (!g323) & (g324) & (g344) & (!g366) & (!g368)) + ((!sk[123]) & (!g323) & (g324) & (g344) & (!g366) & (g368)) + ((!sk[123]) & (!g323) & (g324) & (g344) & (g366) & (!g368)) + ((!sk[123]) & (!g323) & (g324) & (g344) & (g366) & (g368)) + ((!sk[123]) & (g323) & (!g324) & (!g344) & (g366) & (!g368)) + ((!sk[123]) & (g323) & (!g324) & (!g344) & (g366) & (g368)) + ((!sk[123]) & (g323) & (!g324) & (g344) & (!g366) & (!g368)) + ((!sk[123]) & (g323) & (!g324) & (g344) & (!g366) & (g368)) + ((!sk[123]) & (g323) & (!g324) & (g344) & (g366) & (!g368)) + ((!sk[123]) & (g323) & (!g324) & (g344) & (g366) & (g368)) + ((!sk[123]) & (g323) & (g324) & (!g344) & (!g366) & (!g368)) + ((!sk[123]) & (g323) & (g324) & (!g344) & (!g366) & (g368)) + ((!sk[123]) & (g323) & (g324) & (!g344) & (g366) & (!g368)) + ((!sk[123]) & (g323) & (g324) & (!g344) & (g366) & (g368)) + ((!sk[123]) & (g323) & (g324) & (g344) & (!g366) & (!g368)) + ((!sk[123]) & (g323) & (g324) & (g344) & (!g366) & (g368)) + ((!sk[123]) & (g323) & (g324) & (g344) & (g366) & (!g368)) + ((!sk[123]) & (g323) & (g324) & (g344) & (g366) & (g368)) + ((sk[123]) & (!g323) & (!g324) & (!g344) & (!g366) & (!g368)) + ((sk[123]) & (!g323) & (!g324) & (!g344) & (!g366) & (g368)) + ((sk[123]) & (!g323) & (!g324) & (!g344) & (g366) & (!g368)) + ((sk[123]) & (!g323) & (!g324) & (!g344) & (g366) & (g368)) + ((sk[123]) & (!g323) & (!g324) & (g344) & (!g366) & (!g368)) + ((sk[123]) & (!g323) & (!g324) & (g344) & (!g366) & (g368)) + ((sk[123]) & (!g323) & (!g324) & (g344) & (g366) & (!g368)) + ((sk[123]) & (!g323) & (!g324) & (g344) & (g366) & (g368)) + ((sk[123]) & (!g323) & (g324) & (!g344) & (!g366) & (!g368)) + ((sk[123]) & (!g323) & (g324) & (!g344) & (g366) & (!g368)) + ((sk[123]) & (!g323) & (g324) & (!g344) & (g366) & (g368)) + ((sk[123]) & (g323) & (!g324) & (!g344) & (!g366) & (!g368)) + ((sk[123]) & (g323) & (!g324) & (!g344) & (g366) & (!g368)) + ((sk[123]) & (g323) & (!g324) & (!g344) & (g366) & (g368)));
	assign g370 = (((!g252) & (!g122) & (!g159) & (sk[124]) & (g196)) + ((!g252) & (!g122) & (g159) & (!sk[124]) & (!g196)) + ((!g252) & (!g122) & (g159) & (!sk[124]) & (g196)) + ((!g252) & (!g122) & (g159) & (sk[124]) & (!g196)) + ((!g252) & (!g122) & (g159) & (sk[124]) & (g196)) + ((!g252) & (g122) & (g159) & (!sk[124]) & (!g196)) + ((!g252) & (g122) & (g159) & (!sk[124]) & (g196)) + ((g252) & (!g122) & (!g159) & (!sk[124]) & (!g196)) + ((g252) & (!g122) & (!g159) & (!sk[124]) & (g196)) + ((g252) & (!g122) & (!g159) & (sk[124]) & (g196)) + ((g252) & (!g122) & (g159) & (!sk[124]) & (!g196)) + ((g252) & (!g122) & (g159) & (!sk[124]) & (g196)) + ((g252) & (!g122) & (g159) & (sk[124]) & (!g196)) + ((g252) & (g122) & (!g159) & (!sk[124]) & (!g196)) + ((g252) & (g122) & (!g159) & (!sk[124]) & (g196)) + ((g252) & (g122) & (!g159) & (sk[124]) & (!g196)) + ((g252) & (g122) & (g159) & (!sk[124]) & (!g196)) + ((g252) & (g122) & (g159) & (!sk[124]) & (g196)));
	assign g371 = (((!sk[125]) & (!g251) & (!g253) & (!g303) & (g122) & (!g280)) + ((!sk[125]) & (!g251) & (!g253) & (!g303) & (g122) & (g280)) + ((!sk[125]) & (!g251) & (!g253) & (g303) & (g122) & (!g280)) + ((!sk[125]) & (!g251) & (!g253) & (g303) & (g122) & (g280)) + ((!sk[125]) & (!g251) & (g253) & (!g303) & (!g122) & (!g280)) + ((!sk[125]) & (!g251) & (g253) & (!g303) & (!g122) & (g280)) + ((!sk[125]) & (!g251) & (g253) & (!g303) & (g122) & (!g280)) + ((!sk[125]) & (!g251) & (g253) & (!g303) & (g122) & (g280)) + ((!sk[125]) & (!g251) & (g253) & (g303) & (!g122) & (!g280)) + ((!sk[125]) & (!g251) & (g253) & (g303) & (!g122) & (g280)) + ((!sk[125]) & (!g251) & (g253) & (g303) & (g122) & (!g280)) + ((!sk[125]) & (!g251) & (g253) & (g303) & (g122) & (g280)) + ((!sk[125]) & (g251) & (!g253) & (!g303) & (g122) & (!g280)) + ((!sk[125]) & (g251) & (!g253) & (!g303) & (g122) & (g280)) + ((!sk[125]) & (g251) & (!g253) & (g303) & (!g122) & (!g280)) + ((!sk[125]) & (g251) & (!g253) & (g303) & (!g122) & (g280)) + ((!sk[125]) & (g251) & (!g253) & (g303) & (g122) & (!g280)) + ((!sk[125]) & (g251) & (!g253) & (g303) & (g122) & (g280)) + ((!sk[125]) & (g251) & (g253) & (!g303) & (!g122) & (!g280)) + ((!sk[125]) & (g251) & (g253) & (!g303) & (!g122) & (g280)) + ((!sk[125]) & (g251) & (g253) & (!g303) & (g122) & (!g280)) + ((!sk[125]) & (g251) & (g253) & (!g303) & (g122) & (g280)) + ((!sk[125]) & (g251) & (g253) & (g303) & (!g122) & (!g280)) + ((!sk[125]) & (g251) & (g253) & (g303) & (!g122) & (g280)) + ((!sk[125]) & (g251) & (g253) & (g303) & (g122) & (!g280)) + ((!sk[125]) & (g251) & (g253) & (g303) & (g122) & (g280)) + ((sk[125]) & (!g251) & (!g253) & (!g303) & (!g122) & (g280)) + ((sk[125]) & (!g251) & (!g253) & (!g303) & (g122) & (!g280)) + ((sk[125]) & (!g251) & (!g253) & (!g303) & (g122) & (g280)) + ((sk[125]) & (!g251) & (!g253) & (g303) & (!g122) & (g280)) + ((sk[125]) & (!g251) & (!g253) & (g303) & (g122) & (!g280)) + ((sk[125]) & (!g251) & (g253) & (!g303) & (g122) & (g280)) + ((sk[125]) & (g251) & (!g253) & (g303) & (!g122) & (!g280)) + ((sk[125]) & (g251) & (g253) & (!g303) & (!g122) & (g280)) + ((sk[125]) & (g251) & (g253) & (!g303) & (g122) & (!g280)) + ((sk[125]) & (g251) & (g253) & (g303) & (!g122) & (!g280)) + ((sk[125]) & (g251) & (g253) & (g303) & (!g122) & (g280)) + ((sk[125]) & (g251) & (g253) & (g303) & (g122) & (!g280)));
	assign g372 = (((!sk[126]) & (!g69) & (!g198) & (g370) & (!g371)) + ((!sk[126]) & (!g69) & (!g198) & (g370) & (g371)) + ((!sk[126]) & (!g69) & (g198) & (g370) & (!g371)) + ((!sk[126]) & (!g69) & (g198) & (g370) & (g371)) + ((!sk[126]) & (g69) & (!g198) & (!g370) & (!g371)) + ((!sk[126]) & (g69) & (!g198) & (!g370) & (g371)) + ((!sk[126]) & (g69) & (!g198) & (g370) & (!g371)) + ((!sk[126]) & (g69) & (!g198) & (g370) & (g371)) + ((!sk[126]) & (g69) & (g198) & (!g370) & (!g371)) + ((!sk[126]) & (g69) & (g198) & (!g370) & (g371)) + ((!sk[126]) & (g69) & (g198) & (g370) & (!g371)) + ((!sk[126]) & (g69) & (g198) & (g370) & (g371)) + ((sk[126]) & (!g69) & (!g198) & (!g370) & (!g371)) + ((sk[126]) & (!g69) & (g198) & (!g370) & (!g371)) + ((sk[126]) & (!g69) & (g198) & (!g370) & (g371)) + ((sk[126]) & (!g69) & (g198) & (g370) & (!g371)) + ((sk[126]) & (g69) & (!g198) & (!g370) & (!g371)) + ((sk[126]) & (g69) & (g198) & (!g370) & (!g371)));
	assign g373 = (((!g69) & (!g197) & (!g198) & (!g200) & (!g369) & (!g372)) + ((!g69) & (!g197) & (!g198) & (!g200) & (!g369) & (g372)) + ((!g69) & (!g197) & (!g198) & (!g200) & (g369) & (!g372)) + ((!g69) & (!g197) & (!g198) & (g200) & (!g369) & (!g372)) + ((!g69) & (!g197) & (g198) & (!g200) & (!g369) & (!g372)) + ((!g69) & (!g197) & (g198) & (g200) & (!g369) & (!g372)) + ((!g69) & (!g197) & (g198) & (g200) & (!g369) & (g372)) + ((!g69) & (!g197) & (g198) & (g200) & (g369) & (!g372)) + ((!g69) & (g197) & (!g198) & (!g200) & (!g369) & (!g372)) + ((!g69) & (g197) & (!g198) & (g200) & (!g369) & (!g372)) + ((!g69) & (g197) & (!g198) & (g200) & (!g369) & (g372)) + ((!g69) & (g197) & (!g198) & (g200) & (g369) & (!g372)) + ((!g69) & (g197) & (g198) & (!g200) & (!g369) & (!g372)) + ((!g69) & (g197) & (g198) & (!g200) & (!g369) & (g372)) + ((!g69) & (g197) & (g198) & (!g200) & (g369) & (!g372)) + ((!g69) & (g197) & (g198) & (g200) & (!g369) & (!g372)) + ((g69) & (!g197) & (!g198) & (!g200) & (!g369) & (!g372)) + ((g69) & (!g197) & (!g198) & (!g200) & (!g369) & (g372)) + ((g69) & (!g197) & (!g198) & (!g200) & (g369) & (!g372)) + ((g69) & (!g197) & (!g198) & (g200) & (!g369) & (!g372)) + ((g69) & (!g197) & (!g198) & (g200) & (!g369) & (g372)) + ((g69) & (!g197) & (!g198) & (g200) & (g369) & (!g372)) + ((g69) & (!g197) & (g198) & (!g200) & (!g369) & (!g372)) + ((g69) & (!g197) & (g198) & (!g200) & (!g369) & (g372)) + ((g69) & (!g197) & (g198) & (!g200) & (g369) & (!g372)) + ((g69) & (!g197) & (g198) & (g200) & (!g369) & (!g372)) + ((g69) & (!g197) & (g198) & (g200) & (!g369) & (g372)) + ((g69) & (!g197) & (g198) & (g200) & (g369) & (!g372)) + ((g69) & (g197) & (!g198) & (!g200) & (!g369) & (!g372)) + ((g69) & (g197) & (!g198) & (g200) & (!g369) & (!g372)) + ((g69) & (g197) & (g198) & (!g200) & (!g369) & (!g372)) + ((g69) & (g197) & (g198) & (g200) & (!g369) & (!g372)));
	assign g374 = (((!g69) & (!g305) & (!sk[0]) & (g312) & (!g313)) + ((!g69) & (!g305) & (!sk[0]) & (g312) & (g313)) + ((!g69) & (!g305) & (sk[0]) & (!g312) & (g313)) + ((!g69) & (!g305) & (sk[0]) & (g312) & (!g313)) + ((!g69) & (g305) & (!sk[0]) & (g312) & (!g313)) + ((!g69) & (g305) & (!sk[0]) & (g312) & (g313)) + ((!g69) & (g305) & (sk[0]) & (!g312) & (!g313)) + ((!g69) & (g305) & (sk[0]) & (g312) & (g313)) + ((g69) & (!g305) & (!sk[0]) & (!g312) & (!g313)) + ((g69) & (!g305) & (!sk[0]) & (!g312) & (g313)) + ((g69) & (!g305) & (!sk[0]) & (g312) & (!g313)) + ((g69) & (!g305) & (!sk[0]) & (g312) & (g313)) + ((g69) & (!g305) & (sk[0]) & (!g312) & (g313)) + ((g69) & (!g305) & (sk[0]) & (g312) & (!g313)) + ((g69) & (g305) & (!sk[0]) & (!g312) & (!g313)) + ((g69) & (g305) & (!sk[0]) & (!g312) & (g313)) + ((g69) & (g305) & (!sk[0]) & (g312) & (!g313)) + ((g69) & (g305) & (!sk[0]) & (g312) & (g313)) + ((g69) & (g305) & (sk[0]) & (!g312) & (g313)) + ((g69) & (g305) & (sk[0]) & (g312) & (!g313)));
	assign g375 = (((!sk[1]) & (!g201) & (!g223) & (!g281) & (g304) & (!g306)) + ((!sk[1]) & (!g201) & (!g223) & (!g281) & (g304) & (g306)) + ((!sk[1]) & (!g201) & (!g223) & (g281) & (g304) & (!g306)) + ((!sk[1]) & (!g201) & (!g223) & (g281) & (g304) & (g306)) + ((!sk[1]) & (!g201) & (g223) & (!g281) & (!g304) & (!g306)) + ((!sk[1]) & (!g201) & (g223) & (!g281) & (!g304) & (g306)) + ((!sk[1]) & (!g201) & (g223) & (!g281) & (g304) & (!g306)) + ((!sk[1]) & (!g201) & (g223) & (!g281) & (g304) & (g306)) + ((!sk[1]) & (!g201) & (g223) & (g281) & (!g304) & (!g306)) + ((!sk[1]) & (!g201) & (g223) & (g281) & (!g304) & (g306)) + ((!sk[1]) & (!g201) & (g223) & (g281) & (g304) & (!g306)) + ((!sk[1]) & (!g201) & (g223) & (g281) & (g304) & (g306)) + ((!sk[1]) & (g201) & (!g223) & (!g281) & (g304) & (!g306)) + ((!sk[1]) & (g201) & (!g223) & (!g281) & (g304) & (g306)) + ((!sk[1]) & (g201) & (!g223) & (g281) & (!g304) & (!g306)) + ((!sk[1]) & (g201) & (!g223) & (g281) & (!g304) & (g306)) + ((!sk[1]) & (g201) & (!g223) & (g281) & (g304) & (!g306)) + ((!sk[1]) & (g201) & (!g223) & (g281) & (g304) & (g306)) + ((!sk[1]) & (g201) & (g223) & (!g281) & (!g304) & (!g306)) + ((!sk[1]) & (g201) & (g223) & (!g281) & (!g304) & (g306)) + ((!sk[1]) & (g201) & (g223) & (!g281) & (g304) & (!g306)) + ((!sk[1]) & (g201) & (g223) & (!g281) & (g304) & (g306)) + ((!sk[1]) & (g201) & (g223) & (g281) & (!g304) & (!g306)) + ((!sk[1]) & (g201) & (g223) & (g281) & (!g304) & (g306)) + ((!sk[1]) & (g201) & (g223) & (g281) & (g304) & (!g306)) + ((!sk[1]) & (g201) & (g223) & (g281) & (g304) & (g306)) + ((sk[1]) & (!g201) & (!g223) & (!g281) & (g304) & (g306)) + ((sk[1]) & (!g201) & (!g223) & (g281) & (!g304) & (g306)) + ((sk[1]) & (!g201) & (!g223) & (g281) & (g304) & (!g306)) + ((sk[1]) & (!g201) & (!g223) & (g281) & (g304) & (g306)) + ((sk[1]) & (!g201) & (g223) & (!g281) & (!g304) & (!g306)) + ((sk[1]) & (!g201) & (g223) & (!g281) & (!g304) & (g306)) + ((sk[1]) & (!g201) & (g223) & (!g281) & (g304) & (!g306)) + ((sk[1]) & (!g201) & (g223) & (g281) & (!g304) & (!g306)) + ((sk[1]) & (g201) & (!g223) & (!g281) & (!g304) & (!g306)) + ((sk[1]) & (g201) & (!g223) & (!g281) & (!g304) & (g306)) + ((sk[1]) & (g201) & (!g223) & (!g281) & (g304) & (!g306)) + ((sk[1]) & (g201) & (!g223) & (g281) & (!g304) & (!g306)) + ((sk[1]) & (g201) & (g223) & (!g281) & (g304) & (g306)) + ((sk[1]) & (g201) & (g223) & (g281) & (!g304) & (g306)) + ((sk[1]) & (g201) & (g223) & (g281) & (g304) & (!g306)) + ((sk[1]) & (g201) & (g223) & (g281) & (g304) & (g306)));
	assign g376 = (((!sk[2]) & (!g373) & (!g374) & (g375)) + ((!sk[2]) & (!g373) & (g374) & (g375)) + ((!sk[2]) & (g373) & (!g374) & (!g375)) + ((!sk[2]) & (g373) & (!g374) & (g375)) + ((!sk[2]) & (g373) & (g374) & (!g375)) + ((!sk[2]) & (g373) & (g374) & (g375)) + ((sk[2]) & (!g373) & (!g374) & (g375)) + ((sk[2]) & (g373) & (!g374) & (!g375)) + ((sk[2]) & (g373) & (!g374) & (g375)) + ((sk[2]) & (g373) & (g374) & (g375)));
	assign g377 = (((!g307) & (!sk[3]) & (!g309) & (g315)) + ((!g307) & (!sk[3]) & (g309) & (g315)) + ((!g307) & (sk[3]) & (!g309) & (g315)) + ((!g307) & (sk[3]) & (g309) & (!g315)) + ((g307) & (!sk[3]) & (!g309) & (!g315)) + ((g307) & (!sk[3]) & (!g309) & (g315)) + ((g307) & (!sk[3]) & (g309) & (!g315)) + ((g307) & (!sk[3]) & (g309) & (g315)) + ((g307) & (sk[3]) & (!g309) & (!g315)) + ((g307) & (sk[3]) & (g309) & (g315)));
	assign g378 = (((!g301) & (!g251) & (!sk[4]) & (!g302) & (g305) & (!g222)) + ((!g301) & (!g251) & (!sk[4]) & (!g302) & (g305) & (g222)) + ((!g301) & (!g251) & (!sk[4]) & (g302) & (g305) & (!g222)) + ((!g301) & (!g251) & (!sk[4]) & (g302) & (g305) & (g222)) + ((!g301) & (!g251) & (sk[4]) & (g302) & (g305) & (!g222)) + ((!g301) & (!g251) & (sk[4]) & (g302) & (g305) & (g222)) + ((!g301) & (g251) & (!sk[4]) & (!g302) & (!g305) & (!g222)) + ((!g301) & (g251) & (!sk[4]) & (!g302) & (!g305) & (g222)) + ((!g301) & (g251) & (!sk[4]) & (!g302) & (g305) & (!g222)) + ((!g301) & (g251) & (!sk[4]) & (!g302) & (g305) & (g222)) + ((!g301) & (g251) & (!sk[4]) & (g302) & (!g305) & (!g222)) + ((!g301) & (g251) & (!sk[4]) & (g302) & (!g305) & (g222)) + ((!g301) & (g251) & (!sk[4]) & (g302) & (g305) & (!g222)) + ((!g301) & (g251) & (!sk[4]) & (g302) & (g305) & (g222)) + ((!g301) & (g251) & (sk[4]) & (!g302) & (!g305) & (!g222)) + ((!g301) & (g251) & (sk[4]) & (!g302) & (g305) & (!g222)) + ((!g301) & (g251) & (sk[4]) & (g302) & (!g305) & (g222)) + ((!g301) & (g251) & (sk[4]) & (g302) & (g305) & (g222)) + ((g301) & (!g251) & (!sk[4]) & (!g302) & (g305) & (!g222)) + ((g301) & (!g251) & (!sk[4]) & (!g302) & (g305) & (g222)) + ((g301) & (!g251) & (!sk[4]) & (g302) & (!g305) & (!g222)) + ((g301) & (!g251) & (!sk[4]) & (g302) & (!g305) & (g222)) + ((g301) & (!g251) & (!sk[4]) & (g302) & (g305) & (!g222)) + ((g301) & (!g251) & (!sk[4]) & (g302) & (g305) & (g222)) + ((g301) & (!g251) & (sk[4]) & (!g302) & (!g305) & (!g222)) + ((g301) & (!g251) & (sk[4]) & (!g302) & (g305) & (!g222)) + ((g301) & (!g251) & (sk[4]) & (g302) & (!g305) & (g222)) + ((g301) & (!g251) & (sk[4]) & (g302) & (g305) & (g222)) + ((g301) & (g251) & (!sk[4]) & (!g302) & (!g305) & (!g222)) + ((g301) & (g251) & (!sk[4]) & (!g302) & (!g305) & (g222)) + ((g301) & (g251) & (!sk[4]) & (!g302) & (g305) & (!g222)) + ((g301) & (g251) & (!sk[4]) & (!g302) & (g305) & (g222)) + ((g301) & (g251) & (!sk[4]) & (g302) & (!g305) & (!g222)) + ((g301) & (g251) & (!sk[4]) & (g302) & (!g305) & (g222)) + ((g301) & (g251) & (!sk[4]) & (g302) & (g305) & (!g222)) + ((g301) & (g251) & (!sk[4]) & (g302) & (g305) & (g222)) + ((g301) & (g251) & (sk[4]) & (!g302) & (!g305) & (!g222)) + ((g301) & (g251) & (sk[4]) & (!g302) & (!g305) & (g222)));
	assign g379 = (((!g218) & (!g220) & (sk[5]) & (g221) & (!g198) & (!g200)) + ((!g218) & (!g220) & (sk[5]) & (g221) & (!g198) & (g200)) + ((!g218) & (g220) & (!sk[5]) & (!g221) & (!g198) & (!g200)) + ((!g218) & (g220) & (!sk[5]) & (!g221) & (!g198) & (g200)) + ((!g218) & (g220) & (!sk[5]) & (!g221) & (g198) & (!g200)) + ((!g218) & (g220) & (!sk[5]) & (!g221) & (g198) & (g200)) + ((!g218) & (g220) & (!sk[5]) & (g221) & (!g198) & (!g200)) + ((!g218) & (g220) & (!sk[5]) & (g221) & (!g198) & (g200)) + ((!g218) & (g220) & (!sk[5]) & (g221) & (g198) & (!g200)) + ((!g218) & (g220) & (!sk[5]) & (g221) & (g198) & (g200)) + ((!g218) & (g220) & (sk[5]) & (g221) & (!g198) & (!g200)) + ((!g218) & (g220) & (sk[5]) & (g221) & (g198) & (!g200)) + ((g218) & (!g220) & (sk[5]) & (!g221) & (g198) & (!g200)) + ((g218) & (!g220) & (sk[5]) & (!g221) & (g198) & (g200)) + ((g218) & (!g220) & (sk[5]) & (g221) & (!g198) & (!g200)) + ((g218) & (!g220) & (sk[5]) & (g221) & (!g198) & (g200)) + ((g218) & (!g220) & (sk[5]) & (g221) & (g198) & (!g200)) + ((g218) & (!g220) & (sk[5]) & (g221) & (g198) & (g200)) + ((g218) & (g220) & (!sk[5]) & (!g221) & (!g198) & (!g200)) + ((g218) & (g220) & (!sk[5]) & (!g221) & (!g198) & (g200)) + ((g218) & (g220) & (!sk[5]) & (!g221) & (g198) & (!g200)) + ((g218) & (g220) & (!sk[5]) & (!g221) & (g198) & (g200)) + ((g218) & (g220) & (!sk[5]) & (g221) & (!g198) & (!g200)) + ((g218) & (g220) & (!sk[5]) & (g221) & (!g198) & (g200)) + ((g218) & (g220) & (!sk[5]) & (g221) & (g198) & (!g200)) + ((g218) & (g220) & (!sk[5]) & (g221) & (g198) & (g200)) + ((g218) & (g220) & (sk[5]) & (!g221) & (!g198) & (g200)) + ((g218) & (g220) & (sk[5]) & (!g221) & (g198) & (g200)) + ((g218) & (g220) & (sk[5]) & (g221) & (!g198) & (!g200)) + ((g218) & (g220) & (sk[5]) & (g221) & (!g198) & (g200)) + ((g218) & (g220) & (sk[5]) & (g221) & (g198) & (!g200)) + ((g218) & (g220) & (sk[5]) & (g221) & (g198) & (g200)));
	assign g380 = (((!g252) & (!g253) & (!sk[6]) & (g122) & (!g159) & (!g196)) + ((!g252) & (!g253) & (!sk[6]) & (g122) & (!g159) & (g196)) + ((!g252) & (!g253) & (!sk[6]) & (g122) & (g159) & (!g196)) + ((!g252) & (!g253) & (!sk[6]) & (g122) & (g159) & (g196)) + ((!g252) & (!g253) & (sk[6]) & (!g122) & (!g159) & (g196)) + ((!g252) & (!g253) & (sk[6]) & (!g122) & (g159) & (!g196)) + ((!g252) & (!g253) & (sk[6]) & (!g122) & (g159) & (g196)) + ((!g252) & (g253) & (!sk[6]) & (g122) & (!g159) & (!g196)) + ((!g252) & (g253) & (!sk[6]) & (g122) & (!g159) & (g196)) + ((!g252) & (g253) & (!sk[6]) & (g122) & (g159) & (!g196)) + ((!g252) & (g253) & (!sk[6]) & (g122) & (g159) & (g196)) + ((!g252) & (g253) & (sk[6]) & (!g122) & (!g159) & (g196)) + ((!g252) & (g253) & (sk[6]) & (!g122) & (g159) & (!g196)) + ((!g252) & (g253) & (sk[6]) & (g122) & (!g159) & (!g196)) + ((g252) & (!g253) & (!sk[6]) & (!g122) & (!g159) & (!g196)) + ((g252) & (!g253) & (!sk[6]) & (!g122) & (!g159) & (g196)) + ((g252) & (!g253) & (!sk[6]) & (!g122) & (g159) & (!g196)) + ((g252) & (!g253) & (!sk[6]) & (!g122) & (g159) & (g196)) + ((g252) & (!g253) & (!sk[6]) & (g122) & (!g159) & (!g196)) + ((g252) & (!g253) & (!sk[6]) & (g122) & (!g159) & (g196)) + ((g252) & (!g253) & (!sk[6]) & (g122) & (g159) & (!g196)) + ((g252) & (!g253) & (!sk[6]) & (g122) & (g159) & (g196)) + ((g252) & (!g253) & (sk[6]) & (!g122) & (g159) & (g196)) + ((g252) & (!g253) & (sk[6]) & (g122) & (!g159) & (g196)) + ((g252) & (!g253) & (sk[6]) & (g122) & (g159) & (!g196)) + ((g252) & (g253) & (!sk[6]) & (!g122) & (!g159) & (!g196)) + ((g252) & (g253) & (!sk[6]) & (!g122) & (!g159) & (g196)) + ((g252) & (g253) & (!sk[6]) & (!g122) & (g159) & (!g196)) + ((g252) & (g253) & (!sk[6]) & (!g122) & (g159) & (g196)) + ((g252) & (g253) & (!sk[6]) & (g122) & (!g159) & (!g196)) + ((g252) & (g253) & (!sk[6]) & (g122) & (!g159) & (g196)) + ((g252) & (g253) & (!sk[6]) & (g122) & (g159) & (!g196)) + ((g252) & (g253) & (!sk[6]) & (g122) & (g159) & (g196)) + ((g252) & (g253) & (sk[6]) & (g122) & (!g159) & (!g196)) + ((g252) & (g253) & (sk[6]) & (g122) & (!g159) & (g196)) + ((g252) & (g253) & (sk[6]) & (g122) & (g159) & (!g196)));
	assign g381 = (((!g378) & (!g379) & (!sk[7]) & (g380)) + ((!g378) & (g379) & (!sk[7]) & (g380)) + ((!g378) & (g379) & (sk[7]) & (g380)) + ((g378) & (!g379) & (!sk[7]) & (g380)) + ((g378) & (!g379) & (sk[7]) & (g380)) + ((g378) & (g379) & (!sk[7]) & (g380)) + ((g378) & (g379) & (sk[7]) & (!g380)) + ((g378) & (g379) & (sk[7]) & (g380)));
	assign g382 = (((!sk[8]) & (!g69) & (g198) & (g370) & (!g371)) + ((!sk[8]) & (!g69) & (g198) & (g370) & (g371)) + ((!sk[8]) & (g69) & (!g198) & (g370) & (!g371)) + ((!sk[8]) & (g69) & (!g198) & (g370) & (g371)) + ((!sk[8]) & (g69) & (g198) & (!g370) & (!g371)) + ((!sk[8]) & (g69) & (g198) & (!g370) & (g371)) + ((!sk[8]) & (g69) & (g198) & (g370) & (!g371)) + ((!sk[8]) & (g69) & (g198) & (g370) & (g371)) + ((sk[8]) & (!g69) & (!g198) & (!g370) & (!g371)) + ((sk[8]) & (!g69) & (!g198) & (g370) & (g371)) + ((sk[8]) & (!g69) & (g198) & (!g370) & (g371)) + ((sk[8]) & (!g69) & (g198) & (g370) & (!g371)) + ((sk[8]) & (g69) & (!g198) & (!g370) & (!g371)) + ((sk[8]) & (g69) & (!g198) & (g370) & (g371)) + ((sk[8]) & (g69) & (g198) & (!g370) & (!g371)) + ((sk[8]) & (g69) & (g198) & (g370) & (g371)));
	assign g383 = (((!g323) & (!g324) & (sk[9]) & (!g344) & (!g366) & (g368)) + ((!g323) & (!g324) & (sk[9]) & (g344) & (!g366) & (!g368)) + ((!g323) & (!g324) & (sk[9]) & (g344) & (!g366) & (g368)) + ((!g323) & (!g324) & (sk[9]) & (g344) & (g366) & (!g368)) + ((!g323) & (!g324) & (sk[9]) & (g344) & (g366) & (g368)) + ((!g323) & (g324) & (!sk[9]) & (g344) & (!g366) & (!g368)) + ((!g323) & (g324) & (!sk[9]) & (g344) & (!g366) & (g368)) + ((!g323) & (g324) & (!sk[9]) & (g344) & (g366) & (!g368)) + ((!g323) & (g324) & (!sk[9]) & (g344) & (g366) & (g368)) + ((!g323) & (g324) & (sk[9]) & (!g344) & (!g366) & (!g368)) + ((!g323) & (g324) & (sk[9]) & (!g344) & (g366) & (!g368)) + ((!g323) & (g324) & (sk[9]) & (!g344) & (g366) & (g368)) + ((g323) & (!g324) & (!sk[9]) & (g344) & (!g366) & (!g368)) + ((g323) & (!g324) & (!sk[9]) & (g344) & (!g366) & (g368)) + ((g323) & (!g324) & (!sk[9]) & (g344) & (g366) & (!g368)) + ((g323) & (!g324) & (!sk[9]) & (g344) & (g366) & (g368)) + ((g323) & (!g324) & (sk[9]) & (!g344) & (!g366) & (!g368)) + ((g323) & (!g324) & (sk[9]) & (!g344) & (g366) & (!g368)) + ((g323) & (!g324) & (sk[9]) & (!g344) & (g366) & (g368)) + ((g323) & (g324) & (!sk[9]) & (!g344) & (!g366) & (!g368)) + ((g323) & (g324) & (!sk[9]) & (!g344) & (!g366) & (g368)) + ((g323) & (g324) & (!sk[9]) & (!g344) & (g366) & (!g368)) + ((g323) & (g324) & (!sk[9]) & (!g344) & (g366) & (g368)) + ((g323) & (g324) & (!sk[9]) & (g344) & (!g366) & (!g368)) + ((g323) & (g324) & (!sk[9]) & (g344) & (!g366) & (g368)) + ((g323) & (g324) & (!sk[9]) & (g344) & (g366) & (!g368)) + ((g323) & (g324) & (!sk[9]) & (g344) & (g366) & (g368)) + ((g323) & (g324) & (sk[9]) & (!g344) & (!g366) & (g368)) + ((g323) & (g324) & (sk[9]) & (g344) & (!g366) & (!g368)) + ((g323) & (g324) & (sk[9]) & (g344) & (!g366) & (g368)) + ((g323) & (g324) & (sk[9]) & (g344) & (g366) & (!g368)) + ((g323) & (g324) & (sk[9]) & (g344) & (g366) & (g368)));
	assign g384 = (((!g381) & (!sk[10]) & (!g382) & (g383)) + ((!g381) & (!sk[10]) & (g382) & (g383)) + ((!g381) & (sk[10]) & (g382) & (g383)) + ((g381) & (!sk[10]) & (!g382) & (g383)) + ((g381) & (!sk[10]) & (g382) & (g383)) + ((g381) & (sk[10]) & (!g382) & (g383)) + ((g381) & (sk[10]) & (g382) & (!g383)) + ((g381) & (sk[10]) & (g382) & (g383)));
	assign g385 = (((!sk[11]) & (!g281) & (!g304) & (g306)) + ((!sk[11]) & (!g281) & (g304) & (g306)) + ((!sk[11]) & (g281) & (!g304) & (g306)) + ((!sk[11]) & (g281) & (g304) & (g306)) + ((sk[11]) & (!g281) & (!g304) & (g306)) + ((sk[11]) & (!g281) & (g304) & (!g306)) + ((sk[11]) & (g281) & (!g304) & (!g306)) + ((sk[11]) & (g281) & (g304) & (g306)));
	assign g386 = (((!g69) & (!g197) & (!g198) & (!g200) & (!g369) & (!g372)) + ((!g69) & (!g197) & (!g198) & (!g200) & (g369) & (g372)) + ((!g69) & (!g197) & (!g198) & (g200) & (!g369) & (g372)) + ((!g69) & (!g197) & (!g198) & (g200) & (g369) & (!g372)) + ((!g69) & (!g197) & (g198) & (!g200) & (!g369) & (g372)) + ((!g69) & (!g197) & (g198) & (!g200) & (g369) & (!g372)) + ((!g69) & (!g197) & (g198) & (g200) & (!g369) & (!g372)) + ((!g69) & (!g197) & (g198) & (g200) & (g369) & (g372)) + ((!g69) & (g197) & (!g198) & (!g200) & (!g369) & (g372)) + ((!g69) & (g197) & (!g198) & (!g200) & (g369) & (!g372)) + ((!g69) & (g197) & (!g198) & (g200) & (!g369) & (!g372)) + ((!g69) & (g197) & (!g198) & (g200) & (g369) & (g372)) + ((!g69) & (g197) & (g198) & (!g200) & (!g369) & (!g372)) + ((!g69) & (g197) & (g198) & (!g200) & (g369) & (g372)) + ((!g69) & (g197) & (g198) & (g200) & (!g369) & (g372)) + ((!g69) & (g197) & (g198) & (g200) & (g369) & (!g372)) + ((g69) & (!g197) & (!g198) & (!g200) & (!g369) & (!g372)) + ((g69) & (!g197) & (!g198) & (!g200) & (g369) & (g372)) + ((g69) & (!g197) & (!g198) & (g200) & (!g369) & (!g372)) + ((g69) & (!g197) & (!g198) & (g200) & (g369) & (g372)) + ((g69) & (!g197) & (g198) & (!g200) & (!g369) & (!g372)) + ((g69) & (!g197) & (g198) & (!g200) & (g369) & (g372)) + ((g69) & (!g197) & (g198) & (g200) & (!g369) & (!g372)) + ((g69) & (!g197) & (g198) & (g200) & (g369) & (g372)) + ((g69) & (g197) & (!g198) & (!g200) & (!g369) & (g372)) + ((g69) & (g197) & (!g198) & (!g200) & (g369) & (!g372)) + ((g69) & (g197) & (!g198) & (g200) & (!g369) & (g372)) + ((g69) & (g197) & (!g198) & (g200) & (g369) & (!g372)) + ((g69) & (g197) & (g198) & (!g200) & (!g369) & (g372)) + ((g69) & (g197) & (g198) & (!g200) & (g369) & (!g372)) + ((g69) & (g197) & (g198) & (g200) & (!g369) & (g372)) + ((g69) & (g197) & (g198) & (g200) & (g369) & (!g372)));
	assign g387 = (((!g384) & (!g385) & (!sk[13]) & (g386)) + ((!g384) & (g385) & (!sk[13]) & (g386)) + ((!g384) & (g385) & (sk[13]) & (g386)) + ((g384) & (!g385) & (!sk[13]) & (g386)) + ((g384) & (!g385) & (sk[13]) & (g386)) + ((g384) & (g385) & (!sk[13]) & (g386)) + ((g384) & (g385) & (sk[13]) & (!g386)) + ((g384) & (g385) & (sk[13]) & (g386)));
	assign g388 = (((!g373) & (!sk[14]) & (!g374) & (g375)) + ((!g373) & (!sk[14]) & (g374) & (g375)) + ((!g373) & (sk[14]) & (!g374) & (!g375)) + ((!g373) & (sk[14]) & (g374) & (g375)) + ((g373) & (!sk[14]) & (!g374) & (g375)) + ((g373) & (!sk[14]) & (g374) & (g375)) + ((g373) & (sk[14]) & (!g374) & (g375)) + ((g373) & (sk[14]) & (g374) & (!g375)));
	assign g389 = (((!g202) & (!g251) & (!sk[15]) & (!g303) & (!g122) & (g280)) + ((!g202) & (!g251) & (!sk[15]) & (!g303) & (g122) & (g280)) + ((!g202) & (!g251) & (!sk[15]) & (g303) & (!g122) & (g280)) + ((!g202) & (!g251) & (!sk[15]) & (g303) & (g122) & (g280)) + ((!g202) & (!g251) & (sk[15]) & (!g303) & (!g122) & (g280)) + ((!g202) & (!g251) & (sk[15]) & (!g303) & (g122) & (!g280)) + ((!g202) & (!g251) & (sk[15]) & (!g303) & (g122) & (g280)) + ((!g202) & (!g251) & (sk[15]) & (g303) & (g122) & (g280)) + ((!g202) & (g251) & (!sk[15]) & (!g303) & (!g122) & (g280)) + ((!g202) & (g251) & (!sk[15]) & (!g303) & (g122) & (!g280)) + ((!g202) & (g251) & (!sk[15]) & (!g303) & (g122) & (g280)) + ((!g202) & (g251) & (!sk[15]) & (g303) & (!g122) & (g280)) + ((!g202) & (g251) & (!sk[15]) & (g303) & (g122) & (!g280)) + ((!g202) & (g251) & (!sk[15]) & (g303) & (g122) & (g280)) + ((!g202) & (g251) & (sk[15]) & (g303) & (!g122) & (g280)) + ((!g202) & (g251) & (sk[15]) & (g303) & (g122) & (!g280)) + ((g202) & (!g251) & (!sk[15]) & (!g303) & (!g122) & (g280)) + ((g202) & (!g251) & (!sk[15]) & (!g303) & (g122) & (g280)) + ((g202) & (!g251) & (!sk[15]) & (g303) & (!g122) & (g280)) + ((g202) & (!g251) & (!sk[15]) & (g303) & (g122) & (g280)) + ((g202) & (!g251) & (sk[15]) & (!g303) & (!g122) & (g280)) + ((g202) & (!g251) & (sk[15]) & (!g303) & (g122) & (!g280)) + ((g202) & (g251) & (!sk[15]) & (!g303) & (!g122) & (g280)) + ((g202) & (g251) & (!sk[15]) & (!g303) & (g122) & (!g280)) + ((g202) & (g251) & (!sk[15]) & (!g303) & (g122) & (g280)) + ((g202) & (g251) & (!sk[15]) & (g303) & (!g122) & (g280)) + ((g202) & (g251) & (!sk[15]) & (g303) & (g122) & (!g280)) + ((g202) & (g251) & (!sk[15]) & (g303) & (g122) & (g280)) + ((g202) & (g251) & (sk[15]) & (!g303) & (!g122) & (!g280)) + ((g202) & (g251) & (sk[15]) & (g303) & (!g122) & (!g280)) + ((g202) & (g251) & (sk[15]) & (g303) & (!g122) & (g280)) + ((g202) & (g251) & (sk[15]) & (g303) & (g122) & (!g280)));
	assign g390 = (((!g325) & (!g196) & (!g343) & (!g347) & (!g365) & (g368)) + ((!g325) & (!g196) & (!g343) & (!g347) & (g365) & (!g368)) + ((!g325) & (!g196) & (!g343) & (g347) & (!g365) & (g368)) + ((!g325) & (!g196) & (!g343) & (g347) & (g365) & (g368)) + ((!g325) & (!g196) & (g343) & (!g347) & (!g365) & (g368)) + ((!g325) & (!g196) & (g343) & (!g347) & (g365) & (!g368)) + ((!g325) & (!g196) & (g343) & (g347) & (!g365) & (g368)) + ((!g325) & (!g196) & (g343) & (g347) & (g365) & (g368)) + ((!g325) & (g196) & (!g343) & (!g347) & (!g365) & (g368)) + ((!g325) & (g196) & (!g343) & (!g347) & (g365) & (g368)) + ((!g325) & (g196) & (!g343) & (g347) & (!g365) & (g368)) + ((!g325) & (g196) & (!g343) & (g347) & (g365) & (g368)) + ((!g325) & (g196) & (g343) & (!g347) & (!g365) & (g368)) + ((!g325) & (g196) & (g343) & (!g347) & (g365) & (g368)) + ((!g325) & (g196) & (g343) & (g347) & (!g365) & (g368)) + ((!g325) & (g196) & (g343) & (g347) & (g365) & (g368)) + ((g325) & (!g196) & (!g343) & (!g347) & (!g365) & (g368)) + ((g325) & (!g196) & (!g343) & (!g347) & (g365) & (!g368)) + ((g325) & (!g196) & (!g343) & (g347) & (!g365) & (g368)) + ((g325) & (!g196) & (!g343) & (g347) & (g365) & (g368)) + ((g325) & (!g196) & (g343) & (!g347) & (!g365) & (!g368)) + ((g325) & (!g196) & (g343) & (!g347) & (g365) & (!g368)) + ((g325) & (!g196) & (g343) & (g347) & (!g365) & (!g368)) + ((g325) & (!g196) & (g343) & (g347) & (g365) & (!g368)) + ((g325) & (g196) & (!g343) & (!g347) & (!g365) & (g368)) + ((g325) & (g196) & (!g343) & (!g347) & (g365) & (g368)) + ((g325) & (g196) & (!g343) & (g347) & (!g365) & (g368)) + ((g325) & (g196) & (!g343) & (g347) & (g365) & (g368)) + ((g325) & (g196) & (g343) & (!g347) & (!g365) & (!g368)) + ((g325) & (g196) & (g343) & (!g347) & (g365) & (!g368)) + ((g325) & (g196) & (g343) & (g347) & (!g365) & (!g368)) + ((g325) & (g196) & (g343) & (g347) & (g365) & (!g368)));
	assign g391 = (((!g2) & (!sk[17]) & (!g69) & (g347)) + ((!g2) & (!sk[17]) & (g69) & (g347)) + ((g2) & (!sk[17]) & (!g69) & (g347)) + ((g2) & (!sk[17]) & (g69) & (g347)) + ((g2) & (sk[17]) & (!g69) & (!g347)));
	assign g392 = (((!g2) & (!sk[18]) & (!g69) & (g347)) + ((!g2) & (!sk[18]) & (g69) & (g347)) + ((!g2) & (sk[18]) & (!g69) & (g347)) + ((!g2) & (sk[18]) & (g69) & (g347)) + ((g2) & (!sk[18]) & (!g69) & (g347)) + ((g2) & (!sk[18]) & (g69) & (g347)) + ((g2) & (sk[18]) & (g69) & (g347)));
	assign g393 = (((g330) & (g333) & (g339) & (g352) & (g357) & (g361)));
	assign g394 = (((!sk[20]) & (!g252) & (!g196) & (!g347) & (!g365) & (g393)) + ((!sk[20]) & (!g252) & (!g196) & (!g347) & (g365) & (g393)) + ((!sk[20]) & (!g252) & (!g196) & (g347) & (!g365) & (g393)) + ((!sk[20]) & (!g252) & (!g196) & (g347) & (g365) & (g393)) + ((!sk[20]) & (!g252) & (g196) & (!g347) & (!g365) & (g393)) + ((!sk[20]) & (!g252) & (g196) & (!g347) & (g365) & (!g393)) + ((!sk[20]) & (!g252) & (g196) & (!g347) & (g365) & (g393)) + ((!sk[20]) & (!g252) & (g196) & (g347) & (!g365) & (g393)) + ((!sk[20]) & (!g252) & (g196) & (g347) & (g365) & (!g393)) + ((!sk[20]) & (!g252) & (g196) & (g347) & (g365) & (g393)) + ((!sk[20]) & (g252) & (!g196) & (!g347) & (!g365) & (g393)) + ((!sk[20]) & (g252) & (!g196) & (!g347) & (g365) & (g393)) + ((!sk[20]) & (g252) & (!g196) & (g347) & (!g365) & (g393)) + ((!sk[20]) & (g252) & (!g196) & (g347) & (g365) & (g393)) + ((!sk[20]) & (g252) & (g196) & (!g347) & (!g365) & (g393)) + ((!sk[20]) & (g252) & (g196) & (!g347) & (g365) & (!g393)) + ((!sk[20]) & (g252) & (g196) & (!g347) & (g365) & (g393)) + ((!sk[20]) & (g252) & (g196) & (g347) & (!g365) & (g393)) + ((!sk[20]) & (g252) & (g196) & (g347) & (g365) & (!g393)) + ((!sk[20]) & (g252) & (g196) & (g347) & (g365) & (g393)) + ((sk[20]) & (!g252) & (!g196) & (!g347) & (g365) & (!g393)) + ((sk[20]) & (!g252) & (!g196) & (!g347) & (g365) & (g393)) + ((sk[20]) & (!g252) & (!g196) & (g347) & (!g365) & (!g393)) + ((sk[20]) & (!g252) & (!g196) & (g347) & (!g365) & (g393)) + ((sk[20]) & (!g252) & (!g196) & (g347) & (g365) & (!g393)) + ((sk[20]) & (!g252) & (!g196) & (g347) & (g365) & (g393)) + ((sk[20]) & (g252) & (!g196) & (!g347) & (g365) & (!g393)) + ((sk[20]) & (g252) & (!g196) & (!g347) & (g365) & (g393)) + ((sk[20]) & (g252) & (!g196) & (g347) & (!g365) & (!g393)) + ((sk[20]) & (g252) & (!g196) & (g347) & (!g365) & (g393)) + ((sk[20]) & (g252) & (g196) & (!g347) & (!g365) & (!g393)) + ((sk[20]) & (g252) & (g196) & (g347) & (g365) & (!g393)));
	assign g395 = (((!g389) & (!g390) & (!sk[21]) & (!g391) & (!g392) & (g394)) + ((!g389) & (!g390) & (!sk[21]) & (!g391) & (g392) & (g394)) + ((!g389) & (!g390) & (!sk[21]) & (g391) & (!g392) & (g394)) + ((!g389) & (!g390) & (!sk[21]) & (g391) & (g392) & (g394)) + ((!g389) & (!g390) & (sk[21]) & (!g391) & (!g392) & (!g394)) + ((!g389) & (!g390) & (sk[21]) & (!g391) & (g392) & (!g394)) + ((!g389) & (!g390) & (sk[21]) & (!g391) & (g392) & (g394)) + ((!g389) & (g390) & (!sk[21]) & (!g391) & (!g392) & (g394)) + ((!g389) & (g390) & (!sk[21]) & (!g391) & (g392) & (!g394)) + ((!g389) & (g390) & (!sk[21]) & (!g391) & (g392) & (g394)) + ((!g389) & (g390) & (!sk[21]) & (g391) & (!g392) & (g394)) + ((!g389) & (g390) & (!sk[21]) & (g391) & (g392) & (!g394)) + ((!g389) & (g390) & (!sk[21]) & (g391) & (g392) & (g394)) + ((!g389) & (g390) & (sk[21]) & (!g391) & (!g392) & (!g394)) + ((!g389) & (g390) & (sk[21]) & (!g391) & (!g392) & (g394)) + ((!g389) & (g390) & (sk[21]) & (!g391) & (g392) & (!g394)) + ((!g389) & (g390) & (sk[21]) & (!g391) & (g392) & (g394)) + ((!g389) & (g390) & (sk[21]) & (g391) & (!g392) & (!g394)) + ((!g389) & (g390) & (sk[21]) & (g391) & (!g392) & (g394)) + ((!g389) & (g390) & (sk[21]) & (g391) & (g392) & (!g394)) + ((!g389) & (g390) & (sk[21]) & (g391) & (g392) & (g394)) + ((g389) & (!g390) & (!sk[21]) & (!g391) & (!g392) & (g394)) + ((g389) & (!g390) & (!sk[21]) & (!g391) & (g392) & (g394)) + ((g389) & (!g390) & (!sk[21]) & (g391) & (!g392) & (g394)) + ((g389) & (!g390) & (!sk[21]) & (g391) & (g392) & (g394)) + ((g389) & (g390) & (!sk[21]) & (!g391) & (!g392) & (g394)) + ((g389) & (g390) & (!sk[21]) & (!g391) & (g392) & (!g394)) + ((g389) & (g390) & (!sk[21]) & (!g391) & (g392) & (g394)) + ((g389) & (g390) & (!sk[21]) & (g391) & (!g392) & (g394)) + ((g389) & (g390) & (!sk[21]) & (g391) & (g392) & (!g394)) + ((g389) & (g390) & (!sk[21]) & (g391) & (g392) & (g394)) + ((g389) & (g390) & (sk[21]) & (!g391) & (!g392) & (!g394)) + ((g389) & (g390) & (sk[21]) & (!g391) & (g392) & (!g394)) + ((g389) & (g390) & (sk[21]) & (!g391) & (g392) & (g394)));
	assign g396 = (((!g253) & (!g303) & (!g122) & (!sk[22]) & (!g159) & (g196)) + ((!g253) & (!g303) & (!g122) & (!sk[22]) & (g159) & (g196)) + ((!g253) & (!g303) & (!g122) & (sk[22]) & (!g159) & (g196)) + ((!g253) & (!g303) & (!g122) & (sk[22]) & (g159) & (!g196)) + ((!g253) & (!g303) & (!g122) & (sk[22]) & (g159) & (g196)) + ((!g253) & (!g303) & (g122) & (!sk[22]) & (!g159) & (g196)) + ((!g253) & (!g303) & (g122) & (!sk[22]) & (g159) & (g196)) + ((!g253) & (g303) & (!g122) & (!sk[22]) & (!g159) & (!g196)) + ((!g253) & (g303) & (!g122) & (!sk[22]) & (!g159) & (g196)) + ((!g253) & (g303) & (!g122) & (!sk[22]) & (g159) & (!g196)) + ((!g253) & (g303) & (!g122) & (!sk[22]) & (g159) & (g196)) + ((!g253) & (g303) & (!g122) & (sk[22]) & (!g159) & (g196)) + ((!g253) & (g303) & (!g122) & (sk[22]) & (g159) & (!g196)) + ((!g253) & (g303) & (g122) & (!sk[22]) & (!g159) & (!g196)) + ((!g253) & (g303) & (g122) & (!sk[22]) & (!g159) & (g196)) + ((!g253) & (g303) & (g122) & (!sk[22]) & (g159) & (!g196)) + ((!g253) & (g303) & (g122) & (!sk[22]) & (g159) & (g196)) + ((!g253) & (g303) & (g122) & (sk[22]) & (!g159) & (!g196)) + ((g253) & (!g303) & (!g122) & (!sk[22]) & (!g159) & (g196)) + ((g253) & (!g303) & (!g122) & (!sk[22]) & (g159) & (g196)) + ((g253) & (!g303) & (!g122) & (sk[22]) & (g159) & (g196)) + ((g253) & (!g303) & (g122) & (!sk[22]) & (!g159) & (g196)) + ((g253) & (!g303) & (g122) & (!sk[22]) & (g159) & (g196)) + ((g253) & (!g303) & (g122) & (sk[22]) & (!g159) & (g196)) + ((g253) & (!g303) & (g122) & (sk[22]) & (g159) & (!g196)) + ((g253) & (g303) & (!g122) & (!sk[22]) & (!g159) & (!g196)) + ((g253) & (g303) & (!g122) & (!sk[22]) & (!g159) & (g196)) + ((g253) & (g303) & (!g122) & (!sk[22]) & (g159) & (!g196)) + ((g253) & (g303) & (!g122) & (!sk[22]) & (g159) & (g196)) + ((g253) & (g303) & (g122) & (!sk[22]) & (!g159) & (!g196)) + ((g253) & (g303) & (g122) & (!sk[22]) & (!g159) & (g196)) + ((g253) & (g303) & (g122) & (!sk[22]) & (g159) & (!g196)) + ((g253) & (g303) & (g122) & (!sk[22]) & (g159) & (g196)) + ((g253) & (g303) & (g122) & (sk[22]) & (!g159) & (!g196)) + ((g253) & (g303) & (g122) & (sk[22]) & (!g159) & (g196)) + ((g253) & (g303) & (g122) & (sk[22]) & (g159) & (!g196)));
	assign g397 = (((!g202) & (!g251) & (!g122) & (!g280) & (!sk[23]) & (g222)) + ((!g202) & (!g251) & (!g122) & (g280) & (!sk[23]) & (g222)) + ((!g202) & (!g251) & (!g122) & (g280) & (sk[23]) & (!g222)) + ((!g202) & (!g251) & (!g122) & (g280) & (sk[23]) & (g222)) + ((!g202) & (!g251) & (g122) & (!g280) & (!sk[23]) & (g222)) + ((!g202) & (!g251) & (g122) & (!g280) & (sk[23]) & (!g222)) + ((!g202) & (!g251) & (g122) & (!g280) & (sk[23]) & (g222)) + ((!g202) & (!g251) & (g122) & (g280) & (!sk[23]) & (g222)) + ((!g202) & (!g251) & (g122) & (g280) & (sk[23]) & (!g222)) + ((!g202) & (g251) & (!g122) & (!g280) & (!sk[23]) & (!g222)) + ((!g202) & (g251) & (!g122) & (!g280) & (!sk[23]) & (g222)) + ((!g202) & (g251) & (!g122) & (!g280) & (sk[23]) & (g222)) + ((!g202) & (g251) & (!g122) & (g280) & (!sk[23]) & (!g222)) + ((!g202) & (g251) & (!g122) & (g280) & (!sk[23]) & (g222)) + ((!g202) & (g251) & (g122) & (!g280) & (!sk[23]) & (!g222)) + ((!g202) & (g251) & (g122) & (!g280) & (!sk[23]) & (g222)) + ((!g202) & (g251) & (g122) & (g280) & (!sk[23]) & (!g222)) + ((!g202) & (g251) & (g122) & (g280) & (!sk[23]) & (g222)) + ((g202) & (!g251) & (!g122) & (!g280) & (!sk[23]) & (g222)) + ((g202) & (!g251) & (!g122) & (g280) & (!sk[23]) & (g222)) + ((g202) & (!g251) & (g122) & (!g280) & (!sk[23]) & (g222)) + ((g202) & (!g251) & (g122) & (g280) & (!sk[23]) & (g222)) + ((g202) & (!g251) & (g122) & (g280) & (sk[23]) & (!g222)) + ((g202) & (g251) & (!g122) & (!g280) & (!sk[23]) & (!g222)) + ((g202) & (g251) & (!g122) & (!g280) & (!sk[23]) & (g222)) + ((g202) & (g251) & (!g122) & (!g280) & (sk[23]) & (g222)) + ((g202) & (g251) & (!g122) & (g280) & (!sk[23]) & (!g222)) + ((g202) & (g251) & (!g122) & (g280) & (!sk[23]) & (g222)) + ((g202) & (g251) & (!g122) & (g280) & (sk[23]) & (!g222)) + ((g202) & (g251) & (!g122) & (g280) & (sk[23]) & (g222)) + ((g202) & (g251) & (g122) & (!g280) & (!sk[23]) & (!g222)) + ((g202) & (g251) & (g122) & (!g280) & (!sk[23]) & (g222)) + ((g202) & (g251) & (g122) & (!g280) & (sk[23]) & (!g222)) + ((g202) & (g251) & (g122) & (!g280) & (sk[23]) & (g222)) + ((g202) & (g251) & (g122) & (g280) & (!sk[23]) & (!g222)) + ((g202) & (g251) & (g122) & (g280) & (!sk[23]) & (g222)));
	assign g398 = (((!g301) & (!g251) & (!g302) & (!g305) & (!sk[24]) & (g200)) + ((!g301) & (!g251) & (!g302) & (g305) & (!sk[24]) & (g200)) + ((!g301) & (!g251) & (g302) & (!g305) & (!sk[24]) & (g200)) + ((!g301) & (!g251) & (g302) & (!g305) & (sk[24]) & (g200)) + ((!g301) & (!g251) & (g302) & (g305) & (!sk[24]) & (g200)) + ((!g301) & (!g251) & (g302) & (g305) & (sk[24]) & (g200)) + ((!g301) & (g251) & (!g302) & (!g305) & (!sk[24]) & (!g200)) + ((!g301) & (g251) & (!g302) & (!g305) & (!sk[24]) & (g200)) + ((!g301) & (g251) & (!g302) & (!g305) & (sk[24]) & (!g200)) + ((!g301) & (g251) & (!g302) & (!g305) & (sk[24]) & (g200)) + ((!g301) & (g251) & (!g302) & (g305) & (!sk[24]) & (!g200)) + ((!g301) & (g251) & (!g302) & (g305) & (!sk[24]) & (g200)) + ((!g301) & (g251) & (g302) & (!g305) & (!sk[24]) & (!g200)) + ((!g301) & (g251) & (g302) & (!g305) & (!sk[24]) & (g200)) + ((!g301) & (g251) & (g302) & (g305) & (!sk[24]) & (!g200)) + ((!g301) & (g251) & (g302) & (g305) & (!sk[24]) & (g200)) + ((!g301) & (g251) & (g302) & (g305) & (sk[24]) & (!g200)) + ((!g301) & (g251) & (g302) & (g305) & (sk[24]) & (g200)) + ((g301) & (!g251) & (!g302) & (!g305) & (!sk[24]) & (g200)) + ((g301) & (!g251) & (!g302) & (!g305) & (sk[24]) & (!g200)) + ((g301) & (!g251) & (!g302) & (!g305) & (sk[24]) & (g200)) + ((g301) & (!g251) & (!g302) & (g305) & (!sk[24]) & (g200)) + ((g301) & (!g251) & (g302) & (!g305) & (!sk[24]) & (g200)) + ((g301) & (!g251) & (g302) & (g305) & (!sk[24]) & (g200)) + ((g301) & (!g251) & (g302) & (g305) & (sk[24]) & (!g200)) + ((g301) & (!g251) & (g302) & (g305) & (sk[24]) & (g200)) + ((g301) & (g251) & (!g302) & (!g305) & (!sk[24]) & (!g200)) + ((g301) & (g251) & (!g302) & (!g305) & (!sk[24]) & (g200)) + ((g301) & (g251) & (!g302) & (!g305) & (sk[24]) & (!g200)) + ((g301) & (g251) & (!g302) & (g305) & (!sk[24]) & (!g200)) + ((g301) & (g251) & (!g302) & (g305) & (!sk[24]) & (g200)) + ((g301) & (g251) & (!g302) & (g305) & (sk[24]) & (!g200)) + ((g301) & (g251) & (g302) & (!g305) & (!sk[24]) & (!g200)) + ((g301) & (g251) & (g302) & (!g305) & (!sk[24]) & (g200)) + ((g301) & (g251) & (g302) & (g305) & (!sk[24]) & (!g200)) + ((g301) & (g251) & (g302) & (g305) & (!sk[24]) & (g200)));
	assign g399 = (((!g396) & (!sk[25]) & (!g397) & (g398)) + ((!g396) & (!sk[25]) & (g397) & (!g398)) + ((!g396) & (!sk[25]) & (g397) & (g398)) + ((!g396) & (sk[25]) & (g397) & (g398)) + ((g396) & (!sk[25]) & (!g397) & (g398)) + ((g396) & (!sk[25]) & (g397) & (!g398)) + ((g396) & (!sk[25]) & (g397) & (g398)) + ((g396) & (sk[25]) & (!g397) & (g398)) + ((g396) & (sk[25]) & (g397) & (!g398)) + ((g396) & (sk[25]) & (g397) & (g398)));
	assign g400 = (((!sk[26]) & (!g378) & (!g379) & (g380)) + ((!sk[26]) & (!g378) & (g379) & (!g380)) + ((!sk[26]) & (!g378) & (g379) & (g380)) + ((!sk[26]) & (g378) & (!g379) & (g380)) + ((!sk[26]) & (g378) & (g379) & (!g380)) + ((!sk[26]) & (g378) & (g379) & (g380)) + ((sk[26]) & (!g378) & (!g379) & (!g380)) + ((sk[26]) & (!g378) & (g379) & (g380)) + ((sk[26]) & (g378) & (!g379) & (g380)) + ((sk[26]) & (g378) & (g379) & (!g380)));
	assign g401 = (((!ax22x) & (!sk[27]) & (!g1) & (ax4x)) + ((!ax22x) & (!sk[27]) & (g1) & (!ax4x)) + ((!ax22x) & (!sk[27]) & (g1) & (ax4x)) + ((!ax22x) & (sk[27]) & (!g1) & (!ax4x)) + ((!ax22x) & (sk[27]) & (g1) & (ax4x)) + ((ax22x) & (!sk[27]) & (!g1) & (ax4x)) + ((ax22x) & (!sk[27]) & (g1) & (!ax4x)) + ((ax22x) & (!sk[27]) & (g1) & (ax4x)) + ((ax22x) & (sk[27]) & (!g1) & (ax4x)) + ((ax22x) & (sk[27]) & (g1) & (ax4x)));
	assign g402 = (((!g69) & (!g347) & (!sk[28]) & (g401)) + ((!g69) & (!g347) & (sk[28]) & (g401)) + ((!g69) & (g347) & (!sk[28]) & (!g401)) + ((!g69) & (g347) & (!sk[28]) & (g401)) + ((g69) & (!g347) & (!sk[28]) & (g401)) + ((g69) & (g347) & (!sk[28]) & (!g401)) + ((g69) & (g347) & (!sk[28]) & (g401)));
	assign g403 = (((!g252) & (!g253) & (!g196) & (!g347) & (g365) & (!g393)) + ((!g252) & (!g253) & (!g196) & (!g347) & (g365) & (g393)) + ((!g252) & (!g253) & (!g196) & (g347) & (!g365) & (!g393)) + ((!g252) & (!g253) & (!g196) & (g347) & (!g365) & (g393)) + ((!g252) & (!g253) & (!g196) & (g347) & (g365) & (!g393)) + ((!g252) & (!g253) & (!g196) & (g347) & (g365) & (g393)) + ((!g252) & (g253) & (!g196) & (!g347) & (g365) & (!g393)) + ((!g252) & (g253) & (!g196) & (!g347) & (g365) & (g393)) + ((!g252) & (g253) & (!g196) & (g347) & (!g365) & (!g393)) + ((!g252) & (g253) & (!g196) & (g347) & (!g365) & (g393)) + ((!g252) & (g253) & (g196) & (!g347) & (!g365) & (!g393)) + ((!g252) & (g253) & (g196) & (g347) & (g365) & (!g393)) + ((g252) & (!g253) & (!g196) & (g347) & (g365) & (!g393)) + ((g252) & (!g253) & (!g196) & (g347) & (g365) & (g393)) + ((g252) & (!g253) & (g196) & (!g347) & (g365) & (!g393)) + ((g252) & (!g253) & (g196) & (g347) & (!g365) & (!g393)) + ((g252) & (g253) & (g196) & (!g347) & (!g365) & (!g393)) + ((g252) & (g253) & (g196) & (!g347) & (g365) & (!g393)) + ((g252) & (g253) & (g196) & (g347) & (!g365) & (!g393)) + ((g252) & (g253) & (g196) & (g347) & (g365) & (!g393)));
	assign g404 = (((!sk[30]) & (!g69) & (g347) & (!g401) & (!g403)) + ((!sk[30]) & (!g69) & (g347) & (!g401) & (g403)) + ((!sk[30]) & (!g69) & (g347) & (g401) & (!g403)) + ((!sk[30]) & (!g69) & (g347) & (g401) & (g403)) + ((!sk[30]) & (g69) & (g347) & (!g401) & (!g403)) + ((!sk[30]) & (g69) & (g347) & (!g401) & (g403)) + ((!sk[30]) & (g69) & (g347) & (g401) & (!g403)) + ((!sk[30]) & (g69) & (g347) & (g401) & (g403)) + ((sk[30]) & (!g69) & (!g347) & (!g401) & (g403)) + ((sk[30]) & (!g69) & (g347) & (g401) & (g403)) + ((sk[30]) & (g69) & (!g347) & (!g401) & (g403)) + ((sk[30]) & (g69) & (!g347) & (g401) & (g403)));
	assign g405 = (((!g218) & (!g220) & (!g221) & (!g198) & (!sk[31]) & (g367)) + ((!g218) & (!g220) & (!g221) & (g198) & (!sk[31]) & (g367)) + ((!g218) & (!g220) & (g221) & (!g198) & (!sk[31]) & (g367)) + ((!g218) & (!g220) & (g221) & (!g198) & (sk[31]) & (!g367)) + ((!g218) & (!g220) & (g221) & (g198) & (!sk[31]) & (g367)) + ((!g218) & (!g220) & (g221) & (g198) & (sk[31]) & (!g367)) + ((!g218) & (g220) & (!g221) & (!g198) & (!sk[31]) & (!g367)) + ((!g218) & (g220) & (!g221) & (!g198) & (!sk[31]) & (g367)) + ((!g218) & (g220) & (!g221) & (g198) & (!sk[31]) & (!g367)) + ((!g218) & (g220) & (!g221) & (g198) & (!sk[31]) & (g367)) + ((!g218) & (g220) & (g221) & (!g198) & (!sk[31]) & (!g367)) + ((!g218) & (g220) & (g221) & (!g198) & (!sk[31]) & (g367)) + ((!g218) & (g220) & (g221) & (!g198) & (sk[31]) & (!g367)) + ((!g218) & (g220) & (g221) & (!g198) & (sk[31]) & (g367)) + ((!g218) & (g220) & (g221) & (g198) & (!sk[31]) & (!g367)) + ((!g218) & (g220) & (g221) & (g198) & (!sk[31]) & (g367)) + ((g218) & (!g220) & (!g221) & (!g198) & (!sk[31]) & (g367)) + ((g218) & (!g220) & (!g221) & (!g198) & (sk[31]) & (g367)) + ((g218) & (!g220) & (!g221) & (g198) & (!sk[31]) & (g367)) + ((g218) & (!g220) & (!g221) & (g198) & (sk[31]) & (g367)) + ((g218) & (!g220) & (g221) & (!g198) & (!sk[31]) & (g367)) + ((g218) & (!g220) & (g221) & (!g198) & (sk[31]) & (!g367)) + ((g218) & (!g220) & (g221) & (!g198) & (sk[31]) & (g367)) + ((g218) & (!g220) & (g221) & (g198) & (!sk[31]) & (g367)) + ((g218) & (!g220) & (g221) & (g198) & (sk[31]) & (!g367)) + ((g218) & (!g220) & (g221) & (g198) & (sk[31]) & (g367)) + ((g218) & (g220) & (!g221) & (!g198) & (!sk[31]) & (!g367)) + ((g218) & (g220) & (!g221) & (!g198) & (!sk[31]) & (g367)) + ((g218) & (g220) & (!g221) & (g198) & (!sk[31]) & (!g367)) + ((g218) & (g220) & (!g221) & (g198) & (!sk[31]) & (g367)) + ((g218) & (g220) & (!g221) & (g198) & (sk[31]) & (!g367)) + ((g218) & (g220) & (!g221) & (g198) & (sk[31]) & (g367)) + ((g218) & (g220) & (g221) & (!g198) & (!sk[31]) & (!g367)) + ((g218) & (g220) & (g221) & (!g198) & (!sk[31]) & (g367)) + ((g218) & (g220) & (g221) & (!g198) & (sk[31]) & (!g367)) + ((g218) & (g220) & (g221) & (!g198) & (sk[31]) & (g367)) + ((g218) & (g220) & (g221) & (g198) & (!sk[31]) & (!g367)) + ((g218) & (g220) & (g221) & (g198) & (!sk[31]) & (g367)) + ((g218) & (g220) & (g221) & (g198) & (sk[31]) & (!g367)) + ((g218) & (g220) & (g221) & (g198) & (sk[31]) & (g367)));
	assign g406 = (((!g251) & (!g305) & (!g122) & (!sk[32]) & (g280) & (!g222)) + ((!g251) & (!g305) & (!g122) & (!sk[32]) & (g280) & (g222)) + ((!g251) & (!g305) & (!g122) & (sk[32]) & (g280) & (!g222)) + ((!g251) & (!g305) & (g122) & (!sk[32]) & (!g280) & (!g222)) + ((!g251) & (!g305) & (g122) & (!sk[32]) & (!g280) & (g222)) + ((!g251) & (!g305) & (g122) & (!sk[32]) & (g280) & (!g222)) + ((!g251) & (!g305) & (g122) & (!sk[32]) & (g280) & (g222)) + ((!g251) & (!g305) & (g122) & (sk[32]) & (!g280) & (!g222)) + ((!g251) & (!g305) & (g122) & (sk[32]) & (g280) & (!g222)) + ((!g251) & (!g305) & (g122) & (sk[32]) & (g280) & (g222)) + ((!g251) & (g305) & (!g122) & (!sk[32]) & (!g280) & (!g222)) + ((!g251) & (g305) & (!g122) & (!sk[32]) & (!g280) & (g222)) + ((!g251) & (g305) & (!g122) & (!sk[32]) & (g280) & (!g222)) + ((!g251) & (g305) & (!g122) & (!sk[32]) & (g280) & (g222)) + ((!g251) & (g305) & (!g122) & (sk[32]) & (g280) & (!g222)) + ((!g251) & (g305) & (g122) & (!sk[32]) & (!g280) & (!g222)) + ((!g251) & (g305) & (g122) & (!sk[32]) & (!g280) & (g222)) + ((!g251) & (g305) & (g122) & (!sk[32]) & (g280) & (!g222)) + ((!g251) & (g305) & (g122) & (!sk[32]) & (g280) & (g222)) + ((!g251) & (g305) & (g122) & (sk[32]) & (!g280) & (!g222)) + ((g251) & (!g305) & (!g122) & (!sk[32]) & (g280) & (!g222)) + ((g251) & (!g305) & (!g122) & (!sk[32]) & (g280) & (g222)) + ((g251) & (!g305) & (!g122) & (sk[32]) & (g280) & (g222)) + ((g251) & (!g305) & (g122) & (!sk[32]) & (!g280) & (!g222)) + ((g251) & (!g305) & (g122) & (!sk[32]) & (!g280) & (g222)) + ((g251) & (!g305) & (g122) & (!sk[32]) & (g280) & (!g222)) + ((g251) & (!g305) & (g122) & (!sk[32]) & (g280) & (g222)) + ((g251) & (!g305) & (g122) & (sk[32]) & (!g280) & (g222)) + ((g251) & (g305) & (!g122) & (!sk[32]) & (!g280) & (!g222)) + ((g251) & (g305) & (!g122) & (!sk[32]) & (!g280) & (g222)) + ((g251) & (g305) & (!g122) & (!sk[32]) & (g280) & (!g222)) + ((g251) & (g305) & (!g122) & (!sk[32]) & (g280) & (g222)) + ((g251) & (g305) & (!g122) & (sk[32]) & (!g280) & (!g222)) + ((g251) & (g305) & (!g122) & (sk[32]) & (!g280) & (g222)) + ((g251) & (g305) & (!g122) & (sk[32]) & (g280) & (g222)) + ((g251) & (g305) & (g122) & (!sk[32]) & (!g280) & (!g222)) + ((g251) & (g305) & (g122) & (!sk[32]) & (!g280) & (g222)) + ((g251) & (g305) & (g122) & (!sk[32]) & (g280) & (!g222)) + ((g251) & (g305) & (g122) & (!sk[32]) & (g280) & (g222)) + ((g251) & (g305) & (g122) & (sk[32]) & (!g280) & (g222)));
	assign g407 = (((!sk[33]) & (!g202) & (!g303) & (!g122) & (g159) & (!g196)) + ((!sk[33]) & (!g202) & (!g303) & (!g122) & (g159) & (g196)) + ((!sk[33]) & (!g202) & (!g303) & (g122) & (!g159) & (!g196)) + ((!sk[33]) & (!g202) & (!g303) & (g122) & (!g159) & (g196)) + ((!sk[33]) & (!g202) & (!g303) & (g122) & (g159) & (!g196)) + ((!sk[33]) & (!g202) & (!g303) & (g122) & (g159) & (g196)) + ((!sk[33]) & (!g202) & (g303) & (!g122) & (!g159) & (!g196)) + ((!sk[33]) & (!g202) & (g303) & (!g122) & (!g159) & (g196)) + ((!sk[33]) & (!g202) & (g303) & (!g122) & (g159) & (!g196)) + ((!sk[33]) & (!g202) & (g303) & (!g122) & (g159) & (g196)) + ((!sk[33]) & (!g202) & (g303) & (g122) & (!g159) & (!g196)) + ((!sk[33]) & (!g202) & (g303) & (g122) & (!g159) & (g196)) + ((!sk[33]) & (!g202) & (g303) & (g122) & (g159) & (!g196)) + ((!sk[33]) & (!g202) & (g303) & (g122) & (g159) & (g196)) + ((!sk[33]) & (g202) & (!g303) & (!g122) & (g159) & (!g196)) + ((!sk[33]) & (g202) & (!g303) & (!g122) & (g159) & (g196)) + ((!sk[33]) & (g202) & (!g303) & (g122) & (!g159) & (!g196)) + ((!sk[33]) & (g202) & (!g303) & (g122) & (!g159) & (g196)) + ((!sk[33]) & (g202) & (!g303) & (g122) & (g159) & (!g196)) + ((!sk[33]) & (g202) & (!g303) & (g122) & (g159) & (g196)) + ((!sk[33]) & (g202) & (g303) & (!g122) & (!g159) & (!g196)) + ((!sk[33]) & (g202) & (g303) & (!g122) & (!g159) & (g196)) + ((!sk[33]) & (g202) & (g303) & (!g122) & (g159) & (!g196)) + ((!sk[33]) & (g202) & (g303) & (!g122) & (g159) & (g196)) + ((!sk[33]) & (g202) & (g303) & (g122) & (!g159) & (!g196)) + ((!sk[33]) & (g202) & (g303) & (g122) & (!g159) & (g196)) + ((!sk[33]) & (g202) & (g303) & (g122) & (g159) & (!g196)) + ((!sk[33]) & (g202) & (g303) & (g122) & (g159) & (g196)) + ((sk[33]) & (!g202) & (!g303) & (!g122) & (!g159) & (g196)) + ((sk[33]) & (!g202) & (!g303) & (!g122) & (g159) & (!g196)) + ((sk[33]) & (!g202) & (!g303) & (!g122) & (g159) & (g196)) + ((sk[33]) & (!g202) & (g303) & (!g122) & (g159) & (g196)) + ((sk[33]) & (!g202) & (g303) & (g122) & (!g159) & (g196)) + ((sk[33]) & (!g202) & (g303) & (g122) & (g159) & (!g196)) + ((sk[33]) & (g202) & (!g303) & (!g122) & (!g159) & (g196)) + ((sk[33]) & (g202) & (!g303) & (!g122) & (g159) & (!g196)) + ((sk[33]) & (g202) & (!g303) & (g122) & (!g159) & (!g196)) + ((sk[33]) & (g202) & (g303) & (g122) & (!g159) & (!g196)) + ((sk[33]) & (g202) & (g303) & (g122) & (!g159) & (g196)) + ((sk[33]) & (g202) & (g303) & (g122) & (g159) & (!g196)));
	assign g408 = (((!sk[34]) & (!g301) & (!g251) & (!g302) & (g198) & (!g200)) + ((!sk[34]) & (!g301) & (!g251) & (!g302) & (g198) & (g200)) + ((!sk[34]) & (!g301) & (!g251) & (g302) & (!g198) & (!g200)) + ((!sk[34]) & (!g301) & (!g251) & (g302) & (!g198) & (g200)) + ((!sk[34]) & (!g301) & (!g251) & (g302) & (g198) & (!g200)) + ((!sk[34]) & (!g301) & (!g251) & (g302) & (g198) & (g200)) + ((!sk[34]) & (!g301) & (g251) & (!g302) & (!g198) & (!g200)) + ((!sk[34]) & (!g301) & (g251) & (!g302) & (!g198) & (g200)) + ((!sk[34]) & (!g301) & (g251) & (!g302) & (g198) & (!g200)) + ((!sk[34]) & (!g301) & (g251) & (!g302) & (g198) & (g200)) + ((!sk[34]) & (!g301) & (g251) & (g302) & (!g198) & (!g200)) + ((!sk[34]) & (!g301) & (g251) & (g302) & (!g198) & (g200)) + ((!sk[34]) & (!g301) & (g251) & (g302) & (g198) & (!g200)) + ((!sk[34]) & (!g301) & (g251) & (g302) & (g198) & (g200)) + ((!sk[34]) & (g301) & (!g251) & (!g302) & (g198) & (!g200)) + ((!sk[34]) & (g301) & (!g251) & (!g302) & (g198) & (g200)) + ((!sk[34]) & (g301) & (!g251) & (g302) & (!g198) & (!g200)) + ((!sk[34]) & (g301) & (!g251) & (g302) & (!g198) & (g200)) + ((!sk[34]) & (g301) & (!g251) & (g302) & (g198) & (!g200)) + ((!sk[34]) & (g301) & (!g251) & (g302) & (g198) & (g200)) + ((!sk[34]) & (g301) & (g251) & (!g302) & (!g198) & (!g200)) + ((!sk[34]) & (g301) & (g251) & (!g302) & (!g198) & (g200)) + ((!sk[34]) & (g301) & (g251) & (!g302) & (g198) & (!g200)) + ((!sk[34]) & (g301) & (g251) & (!g302) & (g198) & (g200)) + ((!sk[34]) & (g301) & (g251) & (g302) & (!g198) & (!g200)) + ((!sk[34]) & (g301) & (g251) & (g302) & (!g198) & (g200)) + ((!sk[34]) & (g301) & (g251) & (g302) & (g198) & (!g200)) + ((!sk[34]) & (g301) & (g251) & (g302) & (g198) & (g200)) + ((sk[34]) & (!g301) & (!g251) & (g302) & (g198) & (!g200)) + ((sk[34]) & (!g301) & (!g251) & (g302) & (g198) & (g200)) + ((sk[34]) & (!g301) & (g251) & (!g302) & (!g198) & (!g200)) + ((sk[34]) & (!g301) & (g251) & (!g302) & (g198) & (!g200)) + ((sk[34]) & (!g301) & (g251) & (g302) & (!g198) & (g200)) + ((sk[34]) & (!g301) & (g251) & (g302) & (g198) & (g200)) + ((sk[34]) & (g301) & (!g251) & (!g302) & (!g198) & (!g200)) + ((sk[34]) & (g301) & (!g251) & (!g302) & (g198) & (!g200)) + ((sk[34]) & (g301) & (!g251) & (g302) & (!g198) & (g200)) + ((sk[34]) & (g301) & (!g251) & (g302) & (g198) & (g200)) + ((sk[34]) & (g301) & (g251) & (!g302) & (!g198) & (!g200)) + ((sk[34]) & (g301) & (g251) & (!g302) & (!g198) & (g200)));
	assign g409 = (((!g406) & (g407) & (!sk[35]) & (!g408)) + ((!g406) & (g407) & (!sk[35]) & (g408)) + ((!g406) & (g407) & (sk[35]) & (g408)) + ((g406) & (!g407) & (sk[35]) & (g408)) + ((g406) & (g407) & (!sk[35]) & (!g408)) + ((g406) & (g407) & (!sk[35]) & (g408)) + ((g406) & (g407) & (sk[35]) & (!g408)) + ((g406) & (g407) & (sk[35]) & (g408)));
	assign g410 = (((!g399) & (!g400) & (!g402) & (!g404) & (!g405) & (!g409)) + ((!g399) & (!g400) & (!g402) & (!g404) & (!g405) & (g409)) + ((!g399) & (!g400) & (!g402) & (!g404) & (g405) & (!g409)) + ((!g399) & (!g400) & (!g402) & (g404) & (!g405) & (!g409)) + ((!g399) & (!g400) & (g402) & (!g404) & (!g405) & (!g409)) + ((!g399) & (!g400) & (g402) & (g404) & (!g405) & (!g409)) + ((!g399) & (g400) & (!g402) & (!g404) & (!g405) & (!g409)) + ((!g399) & (g400) & (!g402) & (!g404) & (!g405) & (g409)) + ((!g399) & (g400) & (!g402) & (!g404) & (g405) & (!g409)) + ((!g399) & (g400) & (!g402) & (!g404) & (g405) & (g409)) + ((!g399) & (g400) & (!g402) & (g404) & (!g405) & (!g409)) + ((!g399) & (g400) & (!g402) & (g404) & (!g405) & (g409)) + ((!g399) & (g400) & (!g402) & (g404) & (g405) & (!g409)) + ((!g399) & (g400) & (!g402) & (g404) & (g405) & (g409)) + ((!g399) & (g400) & (g402) & (!g404) & (!g405) & (!g409)) + ((!g399) & (g400) & (g402) & (!g404) & (!g405) & (g409)) + ((!g399) & (g400) & (g402) & (!g404) & (g405) & (!g409)) + ((!g399) & (g400) & (g402) & (!g404) & (g405) & (g409)) + ((!g399) & (g400) & (g402) & (g404) & (!g405) & (!g409)) + ((!g399) & (g400) & (g402) & (g404) & (!g405) & (g409)) + ((!g399) & (g400) & (g402) & (g404) & (g405) & (!g409)) + ((!g399) & (g400) & (g402) & (g404) & (g405) & (g409)) + ((g399) & (g400) & (!g402) & (!g404) & (!g405) & (!g409)) + ((g399) & (g400) & (!g402) & (!g404) & (!g405) & (g409)) + ((g399) & (g400) & (!g402) & (!g404) & (g405) & (!g409)) + ((g399) & (g400) & (!g402) & (g404) & (!g405) & (!g409)) + ((g399) & (g400) & (g402) & (!g404) & (!g405) & (!g409)) + ((g399) & (g400) & (g402) & (g404) & (!g405) & (!g409)));
	assign g411 = (((!g381) & (!g382) & (sk[37]) & (g383)) + ((!g381) & (g382) & (!sk[37]) & (!g383)) + ((!g381) & (g382) & (!sk[37]) & (g383)) + ((!g381) & (g382) & (sk[37]) & (!g383)) + ((g381) & (!g382) & (sk[37]) & (!g383)) + ((g381) & (g382) & (!sk[37]) & (!g383)) + ((g381) & (g382) & (!sk[37]) & (g383)) + ((g381) & (g382) & (sk[37]) & (g383)));
	assign g412 = (((!g384) & (!g385) & (g386) & (!g395) & (!g410) & (!g411)) + ((!g384) & (!g385) & (g386) & (!g395) & (!g410) & (g411)) + ((!g384) & (!g385) & (g386) & (!g395) & (g410) & (g411)) + ((!g384) & (!g385) & (g386) & (g395) & (!g410) & (g411)) + ((!g384) & (g385) & (!g386) & (!g395) & (!g410) & (!g411)) + ((!g384) & (g385) & (!g386) & (!g395) & (!g410) & (g411)) + ((!g384) & (g385) & (!g386) & (!g395) & (g410) & (g411)) + ((!g384) & (g385) & (!g386) & (g395) & (!g410) & (g411)) + ((g384) & (!g385) & (!g386) & (!g395) & (!g410) & (!g411)) + ((g384) & (!g385) & (!g386) & (!g395) & (!g410) & (g411)) + ((g384) & (!g385) & (!g386) & (!g395) & (g410) & (g411)) + ((g384) & (!g385) & (!g386) & (g395) & (!g410) & (g411)) + ((g384) & (g385) & (g386) & (!g395) & (!g410) & (!g411)) + ((g384) & (g385) & (g386) & (!g395) & (!g410) & (g411)) + ((g384) & (g385) & (g386) & (!g395) & (g410) & (g411)) + ((g384) & (g385) & (g386) & (g395) & (!g410) & (g411)));
	assign g413 = (((!g384) & (!g385) & (!g386) & (!g395) & (!g410) & (!g411)) + ((!g384) & (!g385) & (!g386) & (!g395) & (!g410) & (g411)) + ((!g384) & (!g385) & (!g386) & (!g395) & (g410) & (g411)) + ((!g384) & (!g385) & (!g386) & (g395) & (!g410) & (g411)) + ((!g384) & (!g385) & (g386) & (!g395) & (g410) & (!g411)) + ((!g384) & (!g385) & (g386) & (g395) & (!g410) & (!g411)) + ((!g384) & (!g385) & (g386) & (g395) & (g410) & (!g411)) + ((!g384) & (!g385) & (g386) & (g395) & (g410) & (g411)) + ((!g384) & (g385) & (!g386) & (!g395) & (g410) & (!g411)) + ((!g384) & (g385) & (!g386) & (g395) & (!g410) & (!g411)) + ((!g384) & (g385) & (!g386) & (g395) & (g410) & (!g411)) + ((!g384) & (g385) & (!g386) & (g395) & (g410) & (g411)) + ((!g384) & (g385) & (g386) & (!g395) & (!g410) & (!g411)) + ((!g384) & (g385) & (g386) & (!g395) & (!g410) & (g411)) + ((!g384) & (g385) & (g386) & (!g395) & (g410) & (g411)) + ((!g384) & (g385) & (g386) & (g395) & (!g410) & (g411)) + ((g384) & (!g385) & (!g386) & (!g395) & (g410) & (!g411)) + ((g384) & (!g385) & (!g386) & (g395) & (!g410) & (!g411)) + ((g384) & (!g385) & (!g386) & (g395) & (g410) & (!g411)) + ((g384) & (!g385) & (!g386) & (g395) & (g410) & (g411)) + ((g384) & (!g385) & (g386) & (!g395) & (!g410) & (!g411)) + ((g384) & (!g385) & (g386) & (!g395) & (!g410) & (g411)) + ((g384) & (!g385) & (g386) & (!g395) & (g410) & (g411)) + ((g384) & (!g385) & (g386) & (g395) & (!g410) & (g411)) + ((g384) & (g385) & (!g386) & (!g395) & (!g410) & (!g411)) + ((g384) & (g385) & (!g386) & (!g395) & (!g410) & (g411)) + ((g384) & (g385) & (!g386) & (!g395) & (g410) & (g411)) + ((g384) & (g385) & (!g386) & (g395) & (!g410) & (g411)) + ((g384) & (g385) & (g386) & (!g395) & (g410) & (!g411)) + ((g384) & (g385) & (g386) & (g395) & (!g410) & (!g411)) + ((g384) & (g385) & (g386) & (g395) & (g410) & (!g411)) + ((g384) & (g385) & (g386) & (g395) & (g410) & (g411)));
	assign g414 = (((!ax22x) & (!sk[40]) & (!ax3x) & (!ax2x) & (ax0x) & (!ax1x)) + ((!ax22x) & (!sk[40]) & (!ax3x) & (!ax2x) & (ax0x) & (ax1x)) + ((!ax22x) & (!sk[40]) & (!ax3x) & (ax2x) & (!ax0x) & (!ax1x)) + ((!ax22x) & (!sk[40]) & (!ax3x) & (ax2x) & (!ax0x) & (ax1x)) + ((!ax22x) & (!sk[40]) & (!ax3x) & (ax2x) & (ax0x) & (!ax1x)) + ((!ax22x) & (!sk[40]) & (!ax3x) & (ax2x) & (ax0x) & (ax1x)) + ((!ax22x) & (!sk[40]) & (ax3x) & (!ax2x) & (!ax0x) & (!ax1x)) + ((!ax22x) & (!sk[40]) & (ax3x) & (!ax2x) & (!ax0x) & (ax1x)) + ((!ax22x) & (!sk[40]) & (ax3x) & (!ax2x) & (ax0x) & (!ax1x)) + ((!ax22x) & (!sk[40]) & (ax3x) & (!ax2x) & (ax0x) & (ax1x)) + ((!ax22x) & (!sk[40]) & (ax3x) & (ax2x) & (!ax0x) & (!ax1x)) + ((!ax22x) & (!sk[40]) & (ax3x) & (ax2x) & (!ax0x) & (ax1x)) + ((!ax22x) & (!sk[40]) & (ax3x) & (ax2x) & (ax0x) & (!ax1x)) + ((!ax22x) & (!sk[40]) & (ax3x) & (ax2x) & (ax0x) & (ax1x)) + ((!ax22x) & (sk[40]) & (!ax3x) & (!ax2x) & (!ax0x) & (ax1x)) + ((!ax22x) & (sk[40]) & (!ax3x) & (!ax2x) & (ax0x) & (!ax1x)) + ((!ax22x) & (sk[40]) & (!ax3x) & (!ax2x) & (ax0x) & (ax1x)) + ((!ax22x) & (sk[40]) & (!ax3x) & (ax2x) & (!ax0x) & (!ax1x)) + ((!ax22x) & (sk[40]) & (!ax3x) & (ax2x) & (!ax0x) & (ax1x)) + ((!ax22x) & (sk[40]) & (!ax3x) & (ax2x) & (ax0x) & (!ax1x)) + ((!ax22x) & (sk[40]) & (!ax3x) & (ax2x) & (ax0x) & (ax1x)) + ((!ax22x) & (sk[40]) & (ax3x) & (!ax2x) & (!ax0x) & (!ax1x)) + ((ax22x) & (!sk[40]) & (!ax3x) & (!ax2x) & (ax0x) & (!ax1x)) + ((ax22x) & (!sk[40]) & (!ax3x) & (!ax2x) & (ax0x) & (ax1x)) + ((ax22x) & (!sk[40]) & (!ax3x) & (ax2x) & (!ax0x) & (!ax1x)) + ((ax22x) & (!sk[40]) & (!ax3x) & (ax2x) & (!ax0x) & (ax1x)) + ((ax22x) & (!sk[40]) & (!ax3x) & (ax2x) & (ax0x) & (!ax1x)) + ((ax22x) & (!sk[40]) & (!ax3x) & (ax2x) & (ax0x) & (ax1x)) + ((ax22x) & (!sk[40]) & (ax3x) & (!ax2x) & (!ax0x) & (!ax1x)) + ((ax22x) & (!sk[40]) & (ax3x) & (!ax2x) & (!ax0x) & (ax1x)) + ((ax22x) & (!sk[40]) & (ax3x) & (!ax2x) & (ax0x) & (!ax1x)) + ((ax22x) & (!sk[40]) & (ax3x) & (!ax2x) & (ax0x) & (ax1x)) + ((ax22x) & (!sk[40]) & (ax3x) & (ax2x) & (!ax0x) & (!ax1x)) + ((ax22x) & (!sk[40]) & (ax3x) & (ax2x) & (!ax0x) & (ax1x)) + ((ax22x) & (!sk[40]) & (ax3x) & (ax2x) & (ax0x) & (!ax1x)) + ((ax22x) & (!sk[40]) & (ax3x) & (ax2x) & (ax0x) & (ax1x)) + ((ax22x) & (sk[40]) & (ax3x) & (!ax2x) & (!ax0x) & (!ax1x)) + ((ax22x) & (sk[40]) & (ax3x) & (!ax2x) & (!ax0x) & (ax1x)) + ((ax22x) & (sk[40]) & (ax3x) & (!ax2x) & (ax0x) & (!ax1x)) + ((ax22x) & (sk[40]) & (ax3x) & (!ax2x) & (ax0x) & (ax1x)) + ((ax22x) & (sk[40]) & (ax3x) & (ax2x) & (!ax0x) & (!ax1x)) + ((ax22x) & (sk[40]) & (ax3x) & (ax2x) & (!ax0x) & (ax1x)) + ((ax22x) & (sk[40]) & (ax3x) & (ax2x) & (ax0x) & (!ax1x)) + ((ax22x) & (sk[40]) & (ax3x) & (ax2x) & (ax0x) & (ax1x)));
	assign g415 = (((!sk[41]) & (!g70) & (!g17) & (!g99) & (g40)) + ((!sk[41]) & (!g70) & (!g17) & (g99) & (g40)) + ((!sk[41]) & (!g70) & (g17) & (!g99) & (g40)) + ((!sk[41]) & (!g70) & (g17) & (g99) & (g40)) + ((!sk[41]) & (g70) & (!g17) & (!g99) & (!g40)) + ((!sk[41]) & (g70) & (!g17) & (!g99) & (g40)) + ((!sk[41]) & (g70) & (!g17) & (g99) & (!g40)) + ((!sk[41]) & (g70) & (!g17) & (g99) & (g40)) + ((!sk[41]) & (g70) & (g17) & (!g99) & (!g40)) + ((!sk[41]) & (g70) & (g17) & (!g99) & (g40)) + ((!sk[41]) & (g70) & (g17) & (g99) & (!g40)) + ((!sk[41]) & (g70) & (g17) & (g99) & (g40)) + ((sk[41]) & (!g70) & (!g17) & (g99) & (g40)) + ((sk[41]) & (!g70) & (g17) & (g99) & (g40)) + ((sk[41]) & (g70) & (!g17) & (g99) & (g40)) + ((sk[41]) & (g70) & (g17) & (!g99) & (!g40)) + ((sk[41]) & (g70) & (g17) & (!g99) & (g40)) + ((sk[41]) & (g70) & (g17) & (g99) & (!g40)) + ((sk[41]) & (g70) & (g17) & (g99) & (g40)));
	assign g416 = (((!g114) & (!g115) & (!g8) & (g40) & (!g25) & (!g27)) + ((!g114) & (!g115) & (!g8) & (g40) & (!g25) & (g27)) + ((!g114) & (!g115) & (!g8) & (g40) & (g25) & (!g27)) + ((!g114) & (!g115) & (!g8) & (g40) & (g25) & (g27)) + ((!g114) & (!g115) & (g8) & (!g40) & (g25) & (!g27)) + ((!g114) & (!g115) & (g8) & (!g40) & (g25) & (g27)) + ((!g114) & (!g115) & (g8) & (g40) & (g25) & (!g27)) + ((!g114) & (!g115) & (g8) & (g40) & (g25) & (g27)) + ((!g114) & (g115) & (g8) & (g40) & (!g25) & (!g27)) + ((!g114) & (g115) & (g8) & (g40) & (!g25) & (g27)) + ((!g114) & (g115) & (g8) & (g40) & (g25) & (!g27)) + ((!g114) & (g115) & (g8) & (g40) & (g25) & (g27)) + ((g114) & (!g115) & (g8) & (!g40) & (!g25) & (g27)) + ((g114) & (!g115) & (g8) & (!g40) & (g25) & (g27)) + ((g114) & (!g115) & (g8) & (g40) & (!g25) & (!g27)) + ((g114) & (!g115) & (g8) & (g40) & (!g25) & (g27)) + ((g114) & (!g115) & (g8) & (g40) & (g25) & (!g27)) + ((g114) & (!g115) & (g8) & (g40) & (g25) & (g27)));
	assign g417 = (((!g99) & (!sk[43]) & (!g12) & (!g32) & (g415) & (!g416)) + ((!g99) & (!sk[43]) & (!g12) & (!g32) & (g415) & (g416)) + ((!g99) & (!sk[43]) & (!g12) & (g32) & (!g415) & (!g416)) + ((!g99) & (!sk[43]) & (!g12) & (g32) & (!g415) & (g416)) + ((!g99) & (!sk[43]) & (!g12) & (g32) & (g415) & (!g416)) + ((!g99) & (!sk[43]) & (!g12) & (g32) & (g415) & (g416)) + ((!g99) & (!sk[43]) & (g12) & (!g32) & (!g415) & (!g416)) + ((!g99) & (!sk[43]) & (g12) & (!g32) & (!g415) & (g416)) + ((!g99) & (!sk[43]) & (g12) & (!g32) & (g415) & (!g416)) + ((!g99) & (!sk[43]) & (g12) & (!g32) & (g415) & (g416)) + ((!g99) & (!sk[43]) & (g12) & (g32) & (!g415) & (!g416)) + ((!g99) & (!sk[43]) & (g12) & (g32) & (!g415) & (g416)) + ((!g99) & (!sk[43]) & (g12) & (g32) & (g415) & (!g416)) + ((!g99) & (!sk[43]) & (g12) & (g32) & (g415) & (g416)) + ((!g99) & (sk[43]) & (!g12) & (!g32) & (!g415) & (!g416)) + ((!g99) & (sk[43]) & (!g12) & (g32) & (!g415) & (!g416)) + ((!g99) & (sk[43]) & (g12) & (!g32) & (!g415) & (!g416)) + ((!g99) & (sk[43]) & (g12) & (g32) & (!g415) & (!g416)) + ((g99) & (!sk[43]) & (!g12) & (!g32) & (g415) & (!g416)) + ((g99) & (!sk[43]) & (!g12) & (!g32) & (g415) & (g416)) + ((g99) & (!sk[43]) & (!g12) & (g32) & (!g415) & (!g416)) + ((g99) & (!sk[43]) & (!g12) & (g32) & (!g415) & (g416)) + ((g99) & (!sk[43]) & (!g12) & (g32) & (g415) & (!g416)) + ((g99) & (!sk[43]) & (!g12) & (g32) & (g415) & (g416)) + ((g99) & (!sk[43]) & (g12) & (!g32) & (!g415) & (!g416)) + ((g99) & (!sk[43]) & (g12) & (!g32) & (!g415) & (g416)) + ((g99) & (!sk[43]) & (g12) & (!g32) & (g415) & (!g416)) + ((g99) & (!sk[43]) & (g12) & (!g32) & (g415) & (g416)) + ((g99) & (!sk[43]) & (g12) & (g32) & (!g415) & (!g416)) + ((g99) & (!sk[43]) & (g12) & (g32) & (!g415) & (g416)) + ((g99) & (!sk[43]) & (g12) & (g32) & (g415) & (!g416)) + ((g99) & (!sk[43]) & (g12) & (g32) & (g415) & (g416)) + ((g99) & (sk[43]) & (!g12) & (!g32) & (!g415) & (!g416)));
	assign g418 = (((!g38) & (!sk[44]) & (!g104) & (!g41) & (g193) & (!g84)) + ((!g38) & (!sk[44]) & (!g104) & (!g41) & (g193) & (g84)) + ((!g38) & (!sk[44]) & (!g104) & (g41) & (!g193) & (!g84)) + ((!g38) & (!sk[44]) & (!g104) & (g41) & (!g193) & (g84)) + ((!g38) & (!sk[44]) & (!g104) & (g41) & (g193) & (!g84)) + ((!g38) & (!sk[44]) & (!g104) & (g41) & (g193) & (g84)) + ((!g38) & (!sk[44]) & (g104) & (!g41) & (!g193) & (!g84)) + ((!g38) & (!sk[44]) & (g104) & (!g41) & (!g193) & (g84)) + ((!g38) & (!sk[44]) & (g104) & (!g41) & (g193) & (!g84)) + ((!g38) & (!sk[44]) & (g104) & (!g41) & (g193) & (g84)) + ((!g38) & (!sk[44]) & (g104) & (g41) & (!g193) & (!g84)) + ((!g38) & (!sk[44]) & (g104) & (g41) & (!g193) & (g84)) + ((!g38) & (!sk[44]) & (g104) & (g41) & (g193) & (!g84)) + ((!g38) & (!sk[44]) & (g104) & (g41) & (g193) & (g84)) + ((!g38) & (sk[44]) & (!g104) & (!g41) & (!g193) & (!g84)) + ((!g38) & (sk[44]) & (!g104) & (g41) & (!g193) & (!g84)) + ((!g38) & (sk[44]) & (g104) & (!g41) & (!g193) & (!g84)) + ((g38) & (!sk[44]) & (!g104) & (!g41) & (g193) & (!g84)) + ((g38) & (!sk[44]) & (!g104) & (!g41) & (g193) & (g84)) + ((g38) & (!sk[44]) & (!g104) & (g41) & (!g193) & (!g84)) + ((g38) & (!sk[44]) & (!g104) & (g41) & (!g193) & (g84)) + ((g38) & (!sk[44]) & (!g104) & (g41) & (g193) & (!g84)) + ((g38) & (!sk[44]) & (!g104) & (g41) & (g193) & (g84)) + ((g38) & (!sk[44]) & (g104) & (!g41) & (!g193) & (!g84)) + ((g38) & (!sk[44]) & (g104) & (!g41) & (!g193) & (g84)) + ((g38) & (!sk[44]) & (g104) & (!g41) & (g193) & (!g84)) + ((g38) & (!sk[44]) & (g104) & (!g41) & (g193) & (g84)) + ((g38) & (!sk[44]) & (g104) & (g41) & (!g193) & (!g84)) + ((g38) & (!sk[44]) & (g104) & (g41) & (!g193) & (g84)) + ((g38) & (!sk[44]) & (g104) & (g41) & (g193) & (!g84)) + ((g38) & (!sk[44]) & (g104) & (g41) & (g193) & (g84)) + ((g38) & (sk[44]) & (!g104) & (!g41) & (!g193) & (!g84)) + ((g38) & (sk[44]) & (!g104) & (g41) & (!g193) & (!g84)));
	assign g419 = (((!g114) & (!g115) & (!g8) & (!g49) & (g18) & (!g25)) + ((!g114) & (!g115) & (!g8) & (!g49) & (g18) & (g25)) + ((!g114) & (!g115) & (!g8) & (g49) & (g18) & (!g25)) + ((!g114) & (!g115) & (!g8) & (g49) & (g18) & (g25)) + ((!g114) & (!g115) & (g8) & (!g49) & (g18) & (!g25)) + ((!g114) & (!g115) & (g8) & (!g49) & (g18) & (g25)) + ((!g114) & (!g115) & (g8) & (g49) & (g18) & (!g25)) + ((!g114) & (!g115) & (g8) & (g49) & (g18) & (g25)) + ((!g114) & (g115) & (g8) & (g49) & (!g18) & (!g25)) + ((!g114) & (g115) & (g8) & (g49) & (!g18) & (g25)) + ((!g114) & (g115) & (g8) & (g49) & (g18) & (!g25)) + ((!g114) & (g115) & (g8) & (g49) & (g18) & (g25)) + ((g114) & (g115) & (!g8) & (!g49) & (!g18) & (g25)) + ((g114) & (g115) & (!g8) & (!g49) & (g18) & (g25)) + ((g114) & (g115) & (!g8) & (g49) & (!g18) & (!g25)) + ((g114) & (g115) & (!g8) & (g49) & (!g18) & (g25)) + ((g114) & (g115) & (!g8) & (g49) & (g18) & (!g25)) + ((g114) & (g115) & (!g8) & (g49) & (g18) & (g25)));
	assign g420 = (((!sk[46]) & (!g153) & (!g19) & (!g50) & (g233)) + ((!sk[46]) & (!g153) & (!g19) & (g50) & (g233)) + ((!sk[46]) & (!g153) & (g19) & (!g50) & (g233)) + ((!sk[46]) & (!g153) & (g19) & (g50) & (g233)) + ((!sk[46]) & (g153) & (!g19) & (!g50) & (!g233)) + ((!sk[46]) & (g153) & (!g19) & (!g50) & (g233)) + ((!sk[46]) & (g153) & (!g19) & (g50) & (!g233)) + ((!sk[46]) & (g153) & (!g19) & (g50) & (g233)) + ((!sk[46]) & (g153) & (g19) & (!g50) & (!g233)) + ((!sk[46]) & (g153) & (g19) & (!g50) & (g233)) + ((!sk[46]) & (g153) & (g19) & (g50) & (!g233)) + ((!sk[46]) & (g153) & (g19) & (g50) & (g233)) + ((sk[46]) & (!g153) & (!g19) & (!g50) & (!g233)));
	assign g421 = (((!sk[47]) & (!g62) & (!g66) & (!g243) & (g268) & (!g420)) + ((!sk[47]) & (!g62) & (!g66) & (!g243) & (g268) & (g420)) + ((!sk[47]) & (!g62) & (!g66) & (g243) & (!g268) & (!g420)) + ((!sk[47]) & (!g62) & (!g66) & (g243) & (!g268) & (g420)) + ((!sk[47]) & (!g62) & (!g66) & (g243) & (g268) & (!g420)) + ((!sk[47]) & (!g62) & (!g66) & (g243) & (g268) & (g420)) + ((!sk[47]) & (!g62) & (g66) & (!g243) & (!g268) & (!g420)) + ((!sk[47]) & (!g62) & (g66) & (!g243) & (!g268) & (g420)) + ((!sk[47]) & (!g62) & (g66) & (!g243) & (g268) & (!g420)) + ((!sk[47]) & (!g62) & (g66) & (!g243) & (g268) & (g420)) + ((!sk[47]) & (!g62) & (g66) & (g243) & (!g268) & (!g420)) + ((!sk[47]) & (!g62) & (g66) & (g243) & (!g268) & (g420)) + ((!sk[47]) & (!g62) & (g66) & (g243) & (g268) & (!g420)) + ((!sk[47]) & (!g62) & (g66) & (g243) & (g268) & (g420)) + ((!sk[47]) & (g62) & (!g66) & (!g243) & (g268) & (!g420)) + ((!sk[47]) & (g62) & (!g66) & (!g243) & (g268) & (g420)) + ((!sk[47]) & (g62) & (!g66) & (g243) & (!g268) & (!g420)) + ((!sk[47]) & (g62) & (!g66) & (g243) & (!g268) & (g420)) + ((!sk[47]) & (g62) & (!g66) & (g243) & (g268) & (!g420)) + ((!sk[47]) & (g62) & (!g66) & (g243) & (g268) & (g420)) + ((!sk[47]) & (g62) & (g66) & (!g243) & (!g268) & (!g420)) + ((!sk[47]) & (g62) & (g66) & (!g243) & (!g268) & (g420)) + ((!sk[47]) & (g62) & (g66) & (!g243) & (g268) & (!g420)) + ((!sk[47]) & (g62) & (g66) & (!g243) & (g268) & (g420)) + ((!sk[47]) & (g62) & (g66) & (g243) & (!g268) & (!g420)) + ((!sk[47]) & (g62) & (g66) & (g243) & (!g268) & (g420)) + ((!sk[47]) & (g62) & (g66) & (g243) & (g268) & (!g420)) + ((!sk[47]) & (g62) & (g66) & (g243) & (g268) & (g420)) + ((sk[47]) & (!g62) & (!g66) & (g243) & (!g268) & (g420)) + ((sk[47]) & (!g62) & (g66) & (g243) & (!g268) & (g420)) + ((sk[47]) & (g62) & (!g66) & (g243) & (!g268) & (g420)));
	assign g422 = (((!g38) & (!g10) & (!g16) & (!g41) & (!g244) & (!g55)) + ((!g38) & (!g10) & (!g16) & (g41) & (!g244) & (!g55)) + ((!g38) & (!g10) & (g16) & (!g41) & (!g244) & (!g55)) + ((!g38) & (g10) & (!g16) & (!g41) & (!g244) & (!g55)) + ((!g38) & (g10) & (!g16) & (g41) & (!g244) & (!g55)) + ((g38) & (!g10) & (!g16) & (!g41) & (!g244) & (!g55)) + ((g38) & (!g10) & (!g16) & (g41) & (!g244) & (!g55)) + ((g38) & (g10) & (!g16) & (!g41) & (!g244) & (!g55)) + ((g38) & (g10) & (!g16) & (g41) & (!g244) & (!g55)));
	assign g423 = (((!sk[49]) & (!g16) & (!g46) & (!g40) & (g20) & (!g247)) + ((!sk[49]) & (!g16) & (!g46) & (!g40) & (g20) & (g247)) + ((!sk[49]) & (!g16) & (!g46) & (g40) & (!g20) & (!g247)) + ((!sk[49]) & (!g16) & (!g46) & (g40) & (!g20) & (g247)) + ((!sk[49]) & (!g16) & (!g46) & (g40) & (g20) & (!g247)) + ((!sk[49]) & (!g16) & (!g46) & (g40) & (g20) & (g247)) + ((!sk[49]) & (!g16) & (g46) & (!g40) & (!g20) & (!g247)) + ((!sk[49]) & (!g16) & (g46) & (!g40) & (!g20) & (g247)) + ((!sk[49]) & (!g16) & (g46) & (!g40) & (g20) & (!g247)) + ((!sk[49]) & (!g16) & (g46) & (!g40) & (g20) & (g247)) + ((!sk[49]) & (!g16) & (g46) & (g40) & (!g20) & (!g247)) + ((!sk[49]) & (!g16) & (g46) & (g40) & (!g20) & (g247)) + ((!sk[49]) & (!g16) & (g46) & (g40) & (g20) & (!g247)) + ((!sk[49]) & (!g16) & (g46) & (g40) & (g20) & (g247)) + ((!sk[49]) & (g16) & (!g46) & (!g40) & (g20) & (!g247)) + ((!sk[49]) & (g16) & (!g46) & (!g40) & (g20) & (g247)) + ((!sk[49]) & (g16) & (!g46) & (g40) & (!g20) & (!g247)) + ((!sk[49]) & (g16) & (!g46) & (g40) & (!g20) & (g247)) + ((!sk[49]) & (g16) & (!g46) & (g40) & (g20) & (!g247)) + ((!sk[49]) & (g16) & (!g46) & (g40) & (g20) & (g247)) + ((!sk[49]) & (g16) & (g46) & (!g40) & (!g20) & (!g247)) + ((!sk[49]) & (g16) & (g46) & (!g40) & (!g20) & (g247)) + ((!sk[49]) & (g16) & (g46) & (!g40) & (g20) & (!g247)) + ((!sk[49]) & (g16) & (g46) & (!g40) & (g20) & (g247)) + ((!sk[49]) & (g16) & (g46) & (g40) & (!g20) & (!g247)) + ((!sk[49]) & (g16) & (g46) & (g40) & (!g20) & (g247)) + ((!sk[49]) & (g16) & (g46) & (g40) & (g20) & (!g247)) + ((!sk[49]) & (g16) & (g46) & (g40) & (g20) & (g247)) + ((sk[49]) & (!g16) & (!g46) & (!g40) & (!g20) & (!g247)) + ((sk[49]) & (!g16) & (!g46) & (!g40) & (!g20) & (g247)) + ((sk[49]) & (!g16) & (!g46) & (!g40) & (g20) & (!g247)) + ((sk[49]) & (!g16) & (!g46) & (!g40) & (g20) & (g247)) + ((sk[49]) & (!g16) & (!g46) & (g40) & (!g20) & (!g247)) + ((sk[49]) & (!g16) & (!g46) & (g40) & (!g20) & (g247)) + ((sk[49]) & (!g16) & (!g46) & (g40) & (g20) & (!g247)) + ((sk[49]) & (!g16) & (!g46) & (g40) & (g20) & (g247)) + ((sk[49]) & (!g16) & (g46) & (!g40) & (!g20) & (!g247)) + ((sk[49]) & (g16) & (!g46) & (!g40) & (!g20) & (!g247)) + ((sk[49]) & (g16) & (!g46) & (!g40) & (!g20) & (g247)) + ((sk[49]) & (g16) & (!g46) & (!g40) & (g20) & (!g247)) + ((sk[49]) & (g16) & (!g46) & (!g40) & (g20) & (g247)) + ((sk[49]) & (g16) & (g46) & (!g40) & (!g20) & (!g247)));
	assign g424 = (((!g141) & (!g86) & (!g154) & (g264) & (g422) & (g423)));
	assign g425 = (((g34) & (g417) & (g418) & (!g419) & (g421) & (g424)));
	assign g426 = (((!sk[52]) & (!g69) & (!g252) & (!g347) & (g414) & (!g425)) + ((!sk[52]) & (!g69) & (!g252) & (!g347) & (g414) & (g425)) + ((!sk[52]) & (!g69) & (!g252) & (g347) & (!g414) & (!g425)) + ((!sk[52]) & (!g69) & (!g252) & (g347) & (!g414) & (g425)) + ((!sk[52]) & (!g69) & (!g252) & (g347) & (g414) & (!g425)) + ((!sk[52]) & (!g69) & (!g252) & (g347) & (g414) & (g425)) + ((!sk[52]) & (!g69) & (g252) & (!g347) & (!g414) & (!g425)) + ((!sk[52]) & (!g69) & (g252) & (!g347) & (!g414) & (g425)) + ((!sk[52]) & (!g69) & (g252) & (!g347) & (g414) & (!g425)) + ((!sk[52]) & (!g69) & (g252) & (!g347) & (g414) & (g425)) + ((!sk[52]) & (!g69) & (g252) & (g347) & (!g414) & (!g425)) + ((!sk[52]) & (!g69) & (g252) & (g347) & (!g414) & (g425)) + ((!sk[52]) & (!g69) & (g252) & (g347) & (g414) & (!g425)) + ((!sk[52]) & (!g69) & (g252) & (g347) & (g414) & (g425)) + ((!sk[52]) & (g69) & (!g252) & (!g347) & (g414) & (!g425)) + ((!sk[52]) & (g69) & (!g252) & (!g347) & (g414) & (g425)) + ((!sk[52]) & (g69) & (!g252) & (g347) & (!g414) & (!g425)) + ((!sk[52]) & (g69) & (!g252) & (g347) & (!g414) & (g425)) + ((!sk[52]) & (g69) & (!g252) & (g347) & (g414) & (!g425)) + ((!sk[52]) & (g69) & (!g252) & (g347) & (g414) & (g425)) + ((!sk[52]) & (g69) & (g252) & (!g347) & (!g414) & (!g425)) + ((!sk[52]) & (g69) & (g252) & (!g347) & (!g414) & (g425)) + ((!sk[52]) & (g69) & (g252) & (!g347) & (g414) & (!g425)) + ((!sk[52]) & (g69) & (g252) & (!g347) & (g414) & (g425)) + ((!sk[52]) & (g69) & (g252) & (g347) & (!g414) & (!g425)) + ((!sk[52]) & (g69) & (g252) & (g347) & (!g414) & (g425)) + ((!sk[52]) & (g69) & (g252) & (g347) & (g414) & (!g425)) + ((!sk[52]) & (g69) & (g252) & (g347) & (g414) & (g425)) + ((sk[52]) & (!g69) & (!g252) & (!g347) & (g414) & (!g425)) + ((sk[52]) & (!g69) & (!g252) & (!g347) & (g414) & (g425)) + ((sk[52]) & (!g69) & (g252) & (!g347) & (g414) & (!g425)));
	assign g427 = (((!sk[53]) & (!g69) & (!g252) & (!g347) & (g414) & (!g425)) + ((!sk[53]) & (!g69) & (!g252) & (!g347) & (g414) & (g425)) + ((!sk[53]) & (!g69) & (!g252) & (g347) & (!g414) & (!g425)) + ((!sk[53]) & (!g69) & (!g252) & (g347) & (!g414) & (g425)) + ((!sk[53]) & (!g69) & (!g252) & (g347) & (g414) & (!g425)) + ((!sk[53]) & (!g69) & (!g252) & (g347) & (g414) & (g425)) + ((!sk[53]) & (!g69) & (g252) & (!g347) & (!g414) & (!g425)) + ((!sk[53]) & (!g69) & (g252) & (!g347) & (!g414) & (g425)) + ((!sk[53]) & (!g69) & (g252) & (!g347) & (g414) & (!g425)) + ((!sk[53]) & (!g69) & (g252) & (!g347) & (g414) & (g425)) + ((!sk[53]) & (!g69) & (g252) & (g347) & (!g414) & (!g425)) + ((!sk[53]) & (!g69) & (g252) & (g347) & (!g414) & (g425)) + ((!sk[53]) & (!g69) & (g252) & (g347) & (g414) & (!g425)) + ((!sk[53]) & (!g69) & (g252) & (g347) & (g414) & (g425)) + ((!sk[53]) & (g69) & (!g252) & (!g347) & (g414) & (!g425)) + ((!sk[53]) & (g69) & (!g252) & (!g347) & (g414) & (g425)) + ((!sk[53]) & (g69) & (!g252) & (g347) & (!g414) & (!g425)) + ((!sk[53]) & (g69) & (!g252) & (g347) & (!g414) & (g425)) + ((!sk[53]) & (g69) & (!g252) & (g347) & (g414) & (!g425)) + ((!sk[53]) & (g69) & (!g252) & (g347) & (g414) & (g425)) + ((!sk[53]) & (g69) & (g252) & (!g347) & (!g414) & (!g425)) + ((!sk[53]) & (g69) & (g252) & (!g347) & (!g414) & (g425)) + ((!sk[53]) & (g69) & (g252) & (!g347) & (g414) & (!g425)) + ((!sk[53]) & (g69) & (g252) & (!g347) & (g414) & (g425)) + ((!sk[53]) & (g69) & (g252) & (g347) & (!g414) & (!g425)) + ((!sk[53]) & (g69) & (g252) & (g347) & (!g414) & (g425)) + ((!sk[53]) & (g69) & (g252) & (g347) & (g414) & (!g425)) + ((!sk[53]) & (g69) & (g252) & (g347) & (g414) & (g425)) + ((sk[53]) & (!g69) & (!g252) & (!g347) & (!g414) & (!g425)) + ((sk[53]) & (!g69) & (!g252) & (!g347) & (!g414) & (g425)) + ((sk[53]) & (!g69) & (!g252) & (g347) & (g414) & (!g425)) + ((sk[53]) & (!g69) & (!g252) & (g347) & (g414) & (g425)) + ((sk[53]) & (!g69) & (g252) & (!g347) & (!g414) & (!g425)) + ((sk[53]) & (!g69) & (g252) & (!g347) & (g414) & (g425)) + ((sk[53]) & (!g69) & (g252) & (g347) & (g414) & (!g425)) + ((sk[53]) & (!g69) & (g252) & (g347) & (g414) & (g425)) + ((sk[53]) & (g69) & (!g252) & (!g347) & (!g414) & (!g425)) + ((sk[53]) & (g69) & (!g252) & (!g347) & (!g414) & (g425)) + ((sk[53]) & (g69) & (!g252) & (!g347) & (g414) & (!g425)) + ((sk[53]) & (g69) & (!g252) & (!g347) & (g414) & (g425)) + ((sk[53]) & (g69) & (g252) & (!g347) & (!g414) & (!g425)) + ((sk[53]) & (g69) & (g252) & (!g347) & (g414) & (!g425)));
	assign g428 = (((!g253) & (!g303) & (!g196) & (!g347) & (g365) & (!g393)) + ((!g253) & (!g303) & (!g196) & (!g347) & (g365) & (g393)) + ((!g253) & (!g303) & (!g196) & (g347) & (!g365) & (!g393)) + ((!g253) & (!g303) & (!g196) & (g347) & (!g365) & (g393)) + ((!g253) & (!g303) & (!g196) & (g347) & (g365) & (!g393)) + ((!g253) & (!g303) & (!g196) & (g347) & (g365) & (g393)) + ((!g253) & (g303) & (!g196) & (!g347) & (g365) & (!g393)) + ((!g253) & (g303) & (!g196) & (!g347) & (g365) & (g393)) + ((!g253) & (g303) & (!g196) & (g347) & (!g365) & (!g393)) + ((!g253) & (g303) & (!g196) & (g347) & (!g365) & (g393)) + ((!g253) & (g303) & (g196) & (!g347) & (!g365) & (!g393)) + ((!g253) & (g303) & (g196) & (g347) & (g365) & (!g393)) + ((g253) & (!g303) & (!g196) & (g347) & (g365) & (!g393)) + ((g253) & (!g303) & (!g196) & (g347) & (g365) & (g393)) + ((g253) & (!g303) & (g196) & (!g347) & (g365) & (!g393)) + ((g253) & (!g303) & (g196) & (g347) & (!g365) & (!g393)) + ((g253) & (g303) & (g196) & (!g347) & (!g365) & (!g393)) + ((g253) & (g303) & (g196) & (!g347) & (g365) & (!g393)) + ((g253) & (g303) & (g196) & (g347) & (!g365) & (!g393)) + ((g253) & (g303) & (g196) & (g347) & (g365) & (!g393)));
	assign g429 = (((g427) & (!sk[55]) & (g428)) + ((g427) & (sk[55]) & (g428)));
	assign g430 = (((!g2) & (!g218) & (!g220) & (g221) & (!sk[56]) & (!g367)) + ((!g2) & (!g218) & (!g220) & (g221) & (!sk[56]) & (g367)) + ((!g2) & (!g218) & (!g220) & (g221) & (sk[56]) & (!g367)) + ((!g2) & (!g218) & (!g220) & (g221) & (sk[56]) & (g367)) + ((!g2) & (!g218) & (g220) & (!g221) & (!sk[56]) & (!g367)) + ((!g2) & (!g218) & (g220) & (!g221) & (!sk[56]) & (g367)) + ((!g2) & (!g218) & (g220) & (g221) & (!sk[56]) & (!g367)) + ((!g2) & (!g218) & (g220) & (g221) & (!sk[56]) & (g367)) + ((!g2) & (!g218) & (g220) & (g221) & (sk[56]) & (!g367)) + ((!g2) & (g218) & (!g220) & (!g221) & (!sk[56]) & (!g367)) + ((!g2) & (g218) & (!g220) & (!g221) & (!sk[56]) & (g367)) + ((!g2) & (g218) & (!g220) & (g221) & (!sk[56]) & (!g367)) + ((!g2) & (g218) & (!g220) & (g221) & (!sk[56]) & (g367)) + ((!g2) & (g218) & (!g220) & (g221) & (sk[56]) & (!g367)) + ((!g2) & (g218) & (!g220) & (g221) & (sk[56]) & (g367)) + ((!g2) & (g218) & (g220) & (!g221) & (!sk[56]) & (!g367)) + ((!g2) & (g218) & (g220) & (!g221) & (!sk[56]) & (g367)) + ((!g2) & (g218) & (g220) & (!g221) & (sk[56]) & (g367)) + ((!g2) & (g218) & (g220) & (g221) & (!sk[56]) & (!g367)) + ((!g2) & (g218) & (g220) & (g221) & (!sk[56]) & (g367)) + ((!g2) & (g218) & (g220) & (g221) & (sk[56]) & (!g367)) + ((!g2) & (g218) & (g220) & (g221) & (sk[56]) & (g367)) + ((g2) & (!g218) & (!g220) & (g221) & (!sk[56]) & (!g367)) + ((g2) & (!g218) & (!g220) & (g221) & (!sk[56]) & (g367)) + ((g2) & (!g218) & (g220) & (!g221) & (!sk[56]) & (!g367)) + ((g2) & (!g218) & (g220) & (!g221) & (!sk[56]) & (g367)) + ((g2) & (!g218) & (g220) & (g221) & (!sk[56]) & (!g367)) + ((g2) & (!g218) & (g220) & (g221) & (!sk[56]) & (g367)) + ((g2) & (!g218) & (g220) & (g221) & (sk[56]) & (!g367)) + ((g2) & (g218) & (!g220) & (!g221) & (!sk[56]) & (!g367)) + ((g2) & (g218) & (!g220) & (!g221) & (!sk[56]) & (g367)) + ((g2) & (g218) & (!g220) & (!g221) & (sk[56]) & (!g367)) + ((g2) & (g218) & (!g220) & (!g221) & (sk[56]) & (g367)) + ((g2) & (g218) & (!g220) & (g221) & (!sk[56]) & (!g367)) + ((g2) & (g218) & (!g220) & (g221) & (!sk[56]) & (g367)) + ((g2) & (g218) & (!g220) & (g221) & (sk[56]) & (!g367)) + ((g2) & (g218) & (!g220) & (g221) & (sk[56]) & (g367)) + ((g2) & (g218) & (g220) & (!g221) & (!sk[56]) & (!g367)) + ((g2) & (g218) & (g220) & (!g221) & (!sk[56]) & (g367)) + ((g2) & (g218) & (g220) & (!g221) & (sk[56]) & (g367)) + ((g2) & (g218) & (g220) & (g221) & (!sk[56]) & (!g367)) + ((g2) & (g218) & (g220) & (g221) & (!sk[56]) & (g367)) + ((g2) & (g218) & (g220) & (g221) & (sk[56]) & (!g367)) + ((g2) & (g218) & (g220) & (g221) & (sk[56]) & (g367)));
	assign g431 = (((!sk[57]) & (!g251) & (!g305) & (!g122) & (g280) & (!g200)) + ((!sk[57]) & (!g251) & (!g305) & (!g122) & (g280) & (g200)) + ((!sk[57]) & (!g251) & (!g305) & (g122) & (!g280) & (!g200)) + ((!sk[57]) & (!g251) & (!g305) & (g122) & (!g280) & (g200)) + ((!sk[57]) & (!g251) & (!g305) & (g122) & (g280) & (!g200)) + ((!sk[57]) & (!g251) & (!g305) & (g122) & (g280) & (g200)) + ((!sk[57]) & (!g251) & (g305) & (!g122) & (!g280) & (!g200)) + ((!sk[57]) & (!g251) & (g305) & (!g122) & (!g280) & (g200)) + ((!sk[57]) & (!g251) & (g305) & (!g122) & (g280) & (!g200)) + ((!sk[57]) & (!g251) & (g305) & (!g122) & (g280) & (g200)) + ((!sk[57]) & (!g251) & (g305) & (g122) & (!g280) & (!g200)) + ((!sk[57]) & (!g251) & (g305) & (g122) & (!g280) & (g200)) + ((!sk[57]) & (!g251) & (g305) & (g122) & (g280) & (!g200)) + ((!sk[57]) & (!g251) & (g305) & (g122) & (g280) & (g200)) + ((!sk[57]) & (g251) & (!g305) & (!g122) & (g280) & (!g200)) + ((!sk[57]) & (g251) & (!g305) & (!g122) & (g280) & (g200)) + ((!sk[57]) & (g251) & (!g305) & (g122) & (!g280) & (!g200)) + ((!sk[57]) & (g251) & (!g305) & (g122) & (!g280) & (g200)) + ((!sk[57]) & (g251) & (!g305) & (g122) & (g280) & (!g200)) + ((!sk[57]) & (g251) & (!g305) & (g122) & (g280) & (g200)) + ((!sk[57]) & (g251) & (g305) & (!g122) & (!g280) & (!g200)) + ((!sk[57]) & (g251) & (g305) & (!g122) & (!g280) & (g200)) + ((!sk[57]) & (g251) & (g305) & (!g122) & (g280) & (!g200)) + ((!sk[57]) & (g251) & (g305) & (!g122) & (g280) & (g200)) + ((!sk[57]) & (g251) & (g305) & (g122) & (!g280) & (!g200)) + ((!sk[57]) & (g251) & (g305) & (g122) & (!g280) & (g200)) + ((!sk[57]) & (g251) & (g305) & (g122) & (g280) & (!g200)) + ((!sk[57]) & (g251) & (g305) & (g122) & (g280) & (g200)) + ((sk[57]) & (!g251) & (!g305) & (!g122) & (g280) & (!g200)) + ((sk[57]) & (!g251) & (!g305) & (!g122) & (g280) & (g200)) + ((sk[57]) & (!g251) & (!g305) & (g122) & (!g280) & (!g200)) + ((sk[57]) & (!g251) & (!g305) & (g122) & (!g280) & (g200)) + ((sk[57]) & (!g251) & (!g305) & (g122) & (g280) & (!g200)) + ((sk[57]) & (!g251) & (g305) & (g122) & (g280) & (!g200)) + ((sk[57]) & (g251) & (!g305) & (!g122) & (!g280) & (g200)) + ((sk[57]) & (g251) & (g305) & (!g122) & (!g280) & (g200)) + ((sk[57]) & (g251) & (g305) & (!g122) & (g280) & (!g200)) + ((sk[57]) & (g251) & (g305) & (!g122) & (g280) & (g200)) + ((sk[57]) & (g251) & (g305) & (g122) & (!g280) & (!g200)) + ((sk[57]) & (g251) & (g305) & (g122) & (!g280) & (g200)));
	assign g432 = (((!g202) & (!g122) & (!g222) & (!g159) & (sk[58]) & (g196)) + ((!g202) & (!g122) & (!g222) & (g159) & (!sk[58]) & (!g196)) + ((!g202) & (!g122) & (!g222) & (g159) & (!sk[58]) & (g196)) + ((!g202) & (!g122) & (!g222) & (g159) & (sk[58]) & (!g196)) + ((!g202) & (!g122) & (!g222) & (g159) & (sk[58]) & (g196)) + ((!g202) & (!g122) & (g222) & (!g159) & (!sk[58]) & (!g196)) + ((!g202) & (!g122) & (g222) & (!g159) & (!sk[58]) & (g196)) + ((!g202) & (!g122) & (g222) & (!g159) & (sk[58]) & (g196)) + ((!g202) & (!g122) & (g222) & (g159) & (!sk[58]) & (!g196)) + ((!g202) & (!g122) & (g222) & (g159) & (!sk[58]) & (g196)) + ((!g202) & (!g122) & (g222) & (g159) & (sk[58]) & (!g196)) + ((!g202) & (g122) & (!g222) & (!g159) & (!sk[58]) & (!g196)) + ((!g202) & (g122) & (!g222) & (!g159) & (!sk[58]) & (g196)) + ((!g202) & (g122) & (!g222) & (g159) & (!sk[58]) & (!g196)) + ((!g202) & (g122) & (!g222) & (g159) & (!sk[58]) & (g196)) + ((!g202) & (g122) & (g222) & (!g159) & (!sk[58]) & (!g196)) + ((!g202) & (g122) & (g222) & (!g159) & (!sk[58]) & (g196)) + ((!g202) & (g122) & (g222) & (!g159) & (sk[58]) & (!g196)) + ((!g202) & (g122) & (g222) & (g159) & (!sk[58]) & (!g196)) + ((!g202) & (g122) & (g222) & (g159) & (!sk[58]) & (g196)) + ((g202) & (!g122) & (!g222) & (g159) & (!sk[58]) & (!g196)) + ((g202) & (!g122) & (!g222) & (g159) & (!sk[58]) & (g196)) + ((g202) & (!g122) & (!g222) & (g159) & (sk[58]) & (g196)) + ((g202) & (!g122) & (g222) & (!g159) & (!sk[58]) & (!g196)) + ((g202) & (!g122) & (g222) & (!g159) & (!sk[58]) & (g196)) + ((g202) & (!g122) & (g222) & (g159) & (!sk[58]) & (!g196)) + ((g202) & (!g122) & (g222) & (g159) & (!sk[58]) & (g196)) + ((g202) & (g122) & (!g222) & (!g159) & (!sk[58]) & (!g196)) + ((g202) & (g122) & (!g222) & (!g159) & (!sk[58]) & (g196)) + ((g202) & (g122) & (!g222) & (!g159) & (sk[58]) & (g196)) + ((g202) & (g122) & (!g222) & (g159) & (!sk[58]) & (!g196)) + ((g202) & (g122) & (!g222) & (g159) & (!sk[58]) & (g196)) + ((g202) & (g122) & (!g222) & (g159) & (sk[58]) & (!g196)) + ((g202) & (g122) & (g222) & (!g159) & (!sk[58]) & (!g196)) + ((g202) & (g122) & (g222) & (!g159) & (!sk[58]) & (g196)) + ((g202) & (g122) & (g222) & (!g159) & (sk[58]) & (!g196)) + ((g202) & (g122) & (g222) & (!g159) & (sk[58]) & (g196)) + ((g202) & (g122) & (g222) & (g159) & (!sk[58]) & (!g196)) + ((g202) & (g122) & (g222) & (g159) & (!sk[58]) & (g196)) + ((g202) & (g122) & (g222) & (g159) & (sk[58]) & (!g196)));
	assign g433 = (((!sk[59]) & (!g301) & (!g251) & (!g302) & (g198) & (!g367)) + ((!sk[59]) & (!g301) & (!g251) & (!g302) & (g198) & (g367)) + ((!sk[59]) & (!g301) & (!g251) & (g302) & (!g198) & (!g367)) + ((!sk[59]) & (!g301) & (!g251) & (g302) & (!g198) & (g367)) + ((!sk[59]) & (!g301) & (!g251) & (g302) & (g198) & (!g367)) + ((!sk[59]) & (!g301) & (!g251) & (g302) & (g198) & (g367)) + ((!sk[59]) & (!g301) & (g251) & (!g302) & (!g198) & (!g367)) + ((!sk[59]) & (!g301) & (g251) & (!g302) & (!g198) & (g367)) + ((!sk[59]) & (!g301) & (g251) & (!g302) & (g198) & (!g367)) + ((!sk[59]) & (!g301) & (g251) & (!g302) & (g198) & (g367)) + ((!sk[59]) & (!g301) & (g251) & (g302) & (!g198) & (!g367)) + ((!sk[59]) & (!g301) & (g251) & (g302) & (!g198) & (g367)) + ((!sk[59]) & (!g301) & (g251) & (g302) & (g198) & (!g367)) + ((!sk[59]) & (!g301) & (g251) & (g302) & (g198) & (g367)) + ((!sk[59]) & (g301) & (!g251) & (!g302) & (g198) & (!g367)) + ((!sk[59]) & (g301) & (!g251) & (!g302) & (g198) & (g367)) + ((!sk[59]) & (g301) & (!g251) & (g302) & (!g198) & (!g367)) + ((!sk[59]) & (g301) & (!g251) & (g302) & (!g198) & (g367)) + ((!sk[59]) & (g301) & (!g251) & (g302) & (g198) & (!g367)) + ((!sk[59]) & (g301) & (!g251) & (g302) & (g198) & (g367)) + ((!sk[59]) & (g301) & (g251) & (!g302) & (!g198) & (!g367)) + ((!sk[59]) & (g301) & (g251) & (!g302) & (!g198) & (g367)) + ((!sk[59]) & (g301) & (g251) & (!g302) & (g198) & (!g367)) + ((!sk[59]) & (g301) & (g251) & (!g302) & (g198) & (g367)) + ((!sk[59]) & (g301) & (g251) & (g302) & (!g198) & (!g367)) + ((!sk[59]) & (g301) & (g251) & (g302) & (!g198) & (g367)) + ((!sk[59]) & (g301) & (g251) & (g302) & (g198) & (!g367)) + ((!sk[59]) & (g301) & (g251) & (g302) & (g198) & (g367)) + ((sk[59]) & (!g301) & (!g251) & (g302) & (!g198) & (g367)) + ((sk[59]) & (!g301) & (!g251) & (g302) & (g198) & (g367)) + ((sk[59]) & (!g301) & (g251) & (!g302) & (!g198) & (!g367)) + ((sk[59]) & (!g301) & (g251) & (!g302) & (!g198) & (g367)) + ((sk[59]) & (!g301) & (g251) & (g302) & (g198) & (!g367)) + ((sk[59]) & (!g301) & (g251) & (g302) & (g198) & (g367)) + ((sk[59]) & (g301) & (!g251) & (!g302) & (!g198) & (!g367)) + ((sk[59]) & (g301) & (!g251) & (!g302) & (!g198) & (g367)) + ((sk[59]) & (g301) & (!g251) & (g302) & (g198) & (!g367)) + ((sk[59]) & (g301) & (!g251) & (g302) & (g198) & (g367)) + ((sk[59]) & (g301) & (g251) & (!g302) & (!g198) & (!g367)) + ((sk[59]) & (g301) & (g251) & (!g302) & (g198) & (!g367)));
	assign g434 = (((!sk[60]) & (!g431) & (g432) & (!g433)) + ((!sk[60]) & (!g431) & (g432) & (g433)) + ((!sk[60]) & (g431) & (g432) & (!g433)) + ((!sk[60]) & (g431) & (g432) & (g433)) + ((sk[60]) & (!g431) & (g432) & (g433)) + ((sk[60]) & (g431) & (!g432) & (g433)) + ((sk[60]) & (g431) & (g432) & (!g433)) + ((sk[60]) & (g431) & (g432) & (g433)));
	assign g435 = (((!g391) & (!sk[61]) & (g392) & (!g394)) + ((!g391) & (!sk[61]) & (g392) & (g394)) + ((!g391) & (sk[61]) & (!g392) & (!g394)) + ((!g391) & (sk[61]) & (g392) & (g394)) + ((g391) & (!sk[61]) & (g392) & (!g394)) + ((g391) & (!sk[61]) & (g392) & (g394)) + ((g391) & (sk[61]) & (!g392) & (g394)) + ((g391) & (sk[61]) & (g392) & (g394)));
	assign g436 = (((!g396) & (!sk[62]) & (g397) & (!g398)) + ((!g396) & (!sk[62]) & (g397) & (g398)) + ((!g396) & (sk[62]) & (!g397) & (!g398)) + ((!g396) & (sk[62]) & (g397) & (g398)) + ((g396) & (!sk[62]) & (g397) & (!g398)) + ((g396) & (!sk[62]) & (g397) & (g398)) + ((g396) & (sk[62]) & (!g397) & (g398)) + ((g396) & (sk[62]) & (g397) & (!g398)));
	assign g437 = (((!g426) & (!g429) & (!g430) & (!g434) & (!g435) & (!g436)) + ((!g426) & (!g429) & (!g430) & (!g434) & (!g435) & (g436)) + ((!g426) & (!g429) & (!g430) & (!g434) & (g435) & (g436)) + ((!g426) & (!g429) & (!g430) & (g434) & (!g435) & (!g436)) + ((!g426) & (!g429) & (!g430) & (g434) & (!g435) & (g436)) + ((!g426) & (!g429) & (!g430) & (g434) & (g435) & (g436)) + ((!g426) & (!g429) & (g430) & (!g434) & (!g435) & (!g436)) + ((!g426) & (!g429) & (g430) & (!g434) & (!g435) & (g436)) + ((!g426) & (!g429) & (g430) & (!g434) & (g435) & (g436)) + ((!g426) & (!g429) & (g430) & (g434) & (!g435) & (g436)) + ((!g426) & (g429) & (!g430) & (!g434) & (!g435) & (!g436)) + ((!g426) & (g429) & (!g430) & (!g434) & (!g435) & (g436)) + ((!g426) & (g429) & (!g430) & (!g434) & (g435) & (g436)) + ((!g426) & (g429) & (!g430) & (g434) & (!g435) & (g436)) + ((!g426) & (g429) & (g430) & (!g434) & (!g435) & (g436)) + ((!g426) & (g429) & (g430) & (g434) & (!g435) & (g436)) + ((g426) & (!g429) & (!g430) & (!g434) & (!g435) & (!g436)) + ((g426) & (!g429) & (!g430) & (!g434) & (!g435) & (g436)) + ((g426) & (!g429) & (!g430) & (!g434) & (g435) & (g436)) + ((g426) & (!g429) & (!g430) & (g434) & (!g435) & (g436)) + ((g426) & (!g429) & (g430) & (!g434) & (!g435) & (g436)) + ((g426) & (!g429) & (g430) & (g434) & (!g435) & (g436)) + ((g426) & (g429) & (!g430) & (!g434) & (!g435) & (!g436)) + ((g426) & (g429) & (!g430) & (!g434) & (!g435) & (g436)) + ((g426) & (g429) & (!g430) & (!g434) & (g435) & (g436)) + ((g426) & (g429) & (!g430) & (g434) & (!g435) & (g436)) + ((g426) & (g429) & (g430) & (!g434) & (!g435) & (g436)) + ((g426) & (g429) & (g430) & (g434) & (!g435) & (g436)));
	assign g438 = (((!sk[64]) & (!g389) & (!g390) & (!g391) & (g392) & (!g394)) + ((!sk[64]) & (!g389) & (!g390) & (!g391) & (g392) & (g394)) + ((!sk[64]) & (!g389) & (!g390) & (g391) & (!g392) & (!g394)) + ((!sk[64]) & (!g389) & (!g390) & (g391) & (!g392) & (g394)) + ((!sk[64]) & (!g389) & (!g390) & (g391) & (g392) & (!g394)) + ((!sk[64]) & (!g389) & (!g390) & (g391) & (g392) & (g394)) + ((!sk[64]) & (!g389) & (g390) & (!g391) & (!g392) & (!g394)) + ((!sk[64]) & (!g389) & (g390) & (!g391) & (!g392) & (g394)) + ((!sk[64]) & (!g389) & (g390) & (!g391) & (g392) & (!g394)) + ((!sk[64]) & (!g389) & (g390) & (!g391) & (g392) & (g394)) + ((!sk[64]) & (!g389) & (g390) & (g391) & (!g392) & (!g394)) + ((!sk[64]) & (!g389) & (g390) & (g391) & (!g392) & (g394)) + ((!sk[64]) & (!g389) & (g390) & (g391) & (g392) & (!g394)) + ((!sk[64]) & (!g389) & (g390) & (g391) & (g392) & (g394)) + ((!sk[64]) & (g389) & (!g390) & (!g391) & (g392) & (!g394)) + ((!sk[64]) & (g389) & (!g390) & (!g391) & (g392) & (g394)) + ((!sk[64]) & (g389) & (!g390) & (g391) & (!g392) & (!g394)) + ((!sk[64]) & (g389) & (!g390) & (g391) & (!g392) & (g394)) + ((!sk[64]) & (g389) & (!g390) & (g391) & (g392) & (!g394)) + ((!sk[64]) & (g389) & (!g390) & (g391) & (g392) & (g394)) + ((!sk[64]) & (g389) & (g390) & (!g391) & (!g392) & (!g394)) + ((!sk[64]) & (g389) & (g390) & (!g391) & (!g392) & (g394)) + ((!sk[64]) & (g389) & (g390) & (!g391) & (g392) & (!g394)) + ((!sk[64]) & (g389) & (g390) & (!g391) & (g392) & (g394)) + ((!sk[64]) & (g389) & (g390) & (g391) & (!g392) & (!g394)) + ((!sk[64]) & (g389) & (g390) & (g391) & (!g392) & (g394)) + ((!sk[64]) & (g389) & (g390) & (g391) & (g392) & (!g394)) + ((!sk[64]) & (g389) & (g390) & (g391) & (g392) & (g394)) + ((sk[64]) & (!g389) & (!g390) & (!g391) & (!g392) & (g394)) + ((sk[64]) & (!g389) & (!g390) & (g391) & (!g392) & (!g394)) + ((sk[64]) & (!g389) & (!g390) & (g391) & (!g392) & (g394)) + ((sk[64]) & (!g389) & (!g390) & (g391) & (g392) & (!g394)) + ((sk[64]) & (!g389) & (!g390) & (g391) & (g392) & (g394)) + ((sk[64]) & (!g389) & (g390) & (!g391) & (!g392) & (!g394)) + ((sk[64]) & (!g389) & (g390) & (!g391) & (g392) & (!g394)) + ((sk[64]) & (!g389) & (g390) & (!g391) & (g392) & (g394)) + ((sk[64]) & (g389) & (!g390) & (!g391) & (!g392) & (!g394)) + ((sk[64]) & (g389) & (!g390) & (!g391) & (g392) & (!g394)) + ((sk[64]) & (g389) & (!g390) & (!g391) & (g392) & (g394)) + ((sk[64]) & (g389) & (g390) & (!g391) & (!g392) & (g394)) + ((sk[64]) & (g389) & (g390) & (g391) & (!g392) & (!g394)) + ((sk[64]) & (g389) & (g390) & (g391) & (!g392) & (g394)) + ((sk[64]) & (g389) & (g390) & (g391) & (g392) & (!g394)) + ((sk[64]) & (g389) & (g390) & (g391) & (g392) & (g394)));
	assign g439 = (((!g399) & (!g400) & (!g402) & (!g404) & (g405) & (g409)) + ((!g399) & (!g400) & (!g402) & (g404) & (!g405) & (g409)) + ((!g399) & (!g400) & (!g402) & (g404) & (g405) & (!g409)) + ((!g399) & (!g400) & (!g402) & (g404) & (g405) & (g409)) + ((!g399) & (!g400) & (g402) & (!g404) & (!g405) & (g409)) + ((!g399) & (!g400) & (g402) & (!g404) & (g405) & (!g409)) + ((!g399) & (!g400) & (g402) & (!g404) & (g405) & (g409)) + ((!g399) & (!g400) & (g402) & (g404) & (!g405) & (g409)) + ((!g399) & (!g400) & (g402) & (g404) & (g405) & (!g409)) + ((!g399) & (!g400) & (g402) & (g404) & (g405) & (g409)) + ((!g399) & (g400) & (!g402) & (!g404) & (!g405) & (!g409)) + ((!g399) & (g400) & (!g402) & (!g404) & (!g405) & (g409)) + ((!g399) & (g400) & (!g402) & (!g404) & (g405) & (!g409)) + ((!g399) & (g400) & (!g402) & (g404) & (!g405) & (!g409)) + ((!g399) & (g400) & (g402) & (!g404) & (!g405) & (!g409)) + ((!g399) & (g400) & (g402) & (g404) & (!g405) & (!g409)) + ((g399) & (!g400) & (!g402) & (!g404) & (!g405) & (!g409)) + ((g399) & (!g400) & (!g402) & (!g404) & (!g405) & (g409)) + ((g399) & (!g400) & (!g402) & (!g404) & (g405) & (!g409)) + ((g399) & (!g400) & (!g402) & (g404) & (!g405) & (!g409)) + ((g399) & (!g400) & (g402) & (!g404) & (!g405) & (!g409)) + ((g399) & (!g400) & (g402) & (g404) & (!g405) & (!g409)) + ((g399) & (g400) & (!g402) & (!g404) & (g405) & (g409)) + ((g399) & (g400) & (!g402) & (g404) & (!g405) & (g409)) + ((g399) & (g400) & (!g402) & (g404) & (g405) & (!g409)) + ((g399) & (g400) & (!g402) & (g404) & (g405) & (g409)) + ((g399) & (g400) & (g402) & (!g404) & (!g405) & (g409)) + ((g399) & (g400) & (g402) & (!g404) & (g405) & (!g409)) + ((g399) & (g400) & (g402) & (!g404) & (g405) & (g409)) + ((g399) & (g400) & (g402) & (g404) & (!g405) & (g409)) + ((g399) & (g400) & (g402) & (g404) & (g405) & (!g409)) + ((g399) & (g400) & (g402) & (g404) & (g405) & (g409)));
	assign g440 = (((!g437) & (!g438) & (sk[66]) & (!g439)) + ((!g437) & (!g438) & (sk[66]) & (g439)) + ((!g437) & (g438) & (!sk[66]) & (!g439)) + ((!g437) & (g438) & (!sk[66]) & (g439)) + ((!g437) & (g438) & (sk[66]) & (!g439)) + ((g437) & (!g438) & (sk[66]) & (!g439)) + ((g437) & (g438) & (!sk[66]) & (!g439)) + ((g437) & (g438) & (!sk[66]) & (g439)));
	assign g441 = (((!sk[67]) & (!g395) & (g410) & (!g411)) + ((!sk[67]) & (!g395) & (g410) & (g411)) + ((!sk[67]) & (g395) & (g410) & (!g411)) + ((!sk[67]) & (g395) & (g410) & (g411)) + ((sk[67]) & (!g395) & (!g410) & (g411)) + ((sk[67]) & (!g395) & (g410) & (!g411)) + ((sk[67]) & (g395) & (!g410) & (!g411)) + ((sk[67]) & (g395) & (g410) & (g411)));
	assign g442 = (((!g218) & (!sk[68]) & (!g220) & (!g221) & (g414)) + ((!g218) & (!sk[68]) & (!g220) & (g221) & (g414)) + ((!g218) & (!sk[68]) & (g220) & (!g221) & (g414)) + ((!g218) & (!sk[68]) & (g220) & (g221) & (g414)) + ((!g218) & (sk[68]) & (!g220) & (g221) & (!g414)) + ((!g218) & (sk[68]) & (!g220) & (g221) & (g414)) + ((!g218) & (sk[68]) & (g220) & (g221) & (!g414)) + ((g218) & (!sk[68]) & (!g220) & (!g221) & (!g414)) + ((g218) & (!sk[68]) & (!g220) & (!g221) & (g414)) + ((g218) & (!sk[68]) & (!g220) & (g221) & (!g414)) + ((g218) & (!sk[68]) & (!g220) & (g221) & (g414)) + ((g218) & (!sk[68]) & (g220) & (!g221) & (!g414)) + ((g218) & (!sk[68]) & (g220) & (!g221) & (g414)) + ((g218) & (!sk[68]) & (g220) & (g221) & (!g414)) + ((g218) & (!sk[68]) & (g220) & (g221) & (g414)) + ((g218) & (sk[68]) & (!g220) & (g221) & (!g414)) + ((g218) & (sk[68]) & (!g220) & (g221) & (g414)) + ((g218) & (sk[68]) & (g220) & (g221) & (!g414)) + ((g218) & (sk[68]) & (g220) & (g221) & (g414)));
	assign g443 = (((!sk[69]) & (!g252) & (!g253) & (!g347) & (g425)) + ((!sk[69]) & (!g252) & (!g253) & (g347) & (g425)) + ((!sk[69]) & (!g252) & (g253) & (!g347) & (g425)) + ((!sk[69]) & (!g252) & (g253) & (g347) & (g425)) + ((!sk[69]) & (g252) & (!g253) & (!g347) & (!g425)) + ((!sk[69]) & (g252) & (!g253) & (!g347) & (g425)) + ((!sk[69]) & (g252) & (!g253) & (g347) & (!g425)) + ((!sk[69]) & (g252) & (!g253) & (g347) & (g425)) + ((!sk[69]) & (g252) & (g253) & (!g347) & (!g425)) + ((!sk[69]) & (g252) & (g253) & (!g347) & (g425)) + ((!sk[69]) & (g252) & (g253) & (g347) & (!g425)) + ((!sk[69]) & (g252) & (g253) & (g347) & (g425)) + ((sk[69]) & (!g252) & (!g253) & (!g347) & (!g425)) + ((sk[69]) & (!g252) & (!g253) & (!g347) & (g425)) + ((sk[69]) & (!g252) & (g253) & (!g347) & (!g425)) + ((sk[69]) & (g252) & (!g253) & (!g347) & (g425)) + ((sk[69]) & (g252) & (!g253) & (g347) & (!g425)) + ((sk[69]) & (g252) & (g253) & (g347) & (!g425)));
	assign g444 = (((!g2) & (!g218) & (!g220) & (!sk[70]) & (g221) & (!g401)) + ((!g2) & (!g218) & (!g220) & (!sk[70]) & (g221) & (g401)) + ((!g2) & (!g218) & (!g220) & (sk[70]) & (g221) & (!g401)) + ((!g2) & (!g218) & (g220) & (!sk[70]) & (!g221) & (!g401)) + ((!g2) & (!g218) & (g220) & (!sk[70]) & (!g221) & (g401)) + ((!g2) & (!g218) & (g220) & (!sk[70]) & (g221) & (!g401)) + ((!g2) & (!g218) & (g220) & (!sk[70]) & (g221) & (g401)) + ((!g2) & (!g218) & (g220) & (sk[70]) & (g221) & (!g401)) + ((!g2) & (!g218) & (g220) & (sk[70]) & (g221) & (g401)) + ((!g2) & (g218) & (!g220) & (!sk[70]) & (!g221) & (!g401)) + ((!g2) & (g218) & (!g220) & (!sk[70]) & (!g221) & (g401)) + ((!g2) & (g218) & (!g220) & (!sk[70]) & (g221) & (!g401)) + ((!g2) & (g218) & (!g220) & (!sk[70]) & (g221) & (g401)) + ((!g2) & (g218) & (!g220) & (sk[70]) & (!g221) & (g401)) + ((!g2) & (g218) & (!g220) & (sk[70]) & (g221) & (!g401)) + ((!g2) & (g218) & (!g220) & (sk[70]) & (g221) & (g401)) + ((!g2) & (g218) & (g220) & (!sk[70]) & (!g221) & (!g401)) + ((!g2) & (g218) & (g220) & (!sk[70]) & (!g221) & (g401)) + ((!g2) & (g218) & (g220) & (!sk[70]) & (g221) & (!g401)) + ((!g2) & (g218) & (g220) & (!sk[70]) & (g221) & (g401)) + ((!g2) & (g218) & (g220) & (sk[70]) & (g221) & (!g401)) + ((!g2) & (g218) & (g220) & (sk[70]) & (g221) & (g401)) + ((g2) & (!g218) & (!g220) & (!sk[70]) & (g221) & (!g401)) + ((g2) & (!g218) & (!g220) & (!sk[70]) & (g221) & (g401)) + ((g2) & (!g218) & (!g220) & (sk[70]) & (g221) & (!g401)) + ((g2) & (!g218) & (g220) & (!sk[70]) & (!g221) & (!g401)) + ((g2) & (!g218) & (g220) & (!sk[70]) & (!g221) & (g401)) + ((g2) & (!g218) & (g220) & (!sk[70]) & (g221) & (!g401)) + ((g2) & (!g218) & (g220) & (!sk[70]) & (g221) & (g401)) + ((g2) & (g218) & (!g220) & (!sk[70]) & (!g221) & (!g401)) + ((g2) & (g218) & (!g220) & (!sk[70]) & (!g221) & (g401)) + ((g2) & (g218) & (!g220) & (!sk[70]) & (g221) & (!g401)) + ((g2) & (g218) & (!g220) & (!sk[70]) & (g221) & (g401)) + ((g2) & (g218) & (!g220) & (sk[70]) & (!g221) & (g401)) + ((g2) & (g218) & (!g220) & (sk[70]) & (g221) & (!g401)) + ((g2) & (g218) & (!g220) & (sk[70]) & (g221) & (g401)) + ((g2) & (g218) & (g220) & (!sk[70]) & (!g221) & (!g401)) + ((g2) & (g218) & (g220) & (!sk[70]) & (!g221) & (g401)) + ((g2) & (g218) & (g220) & (!sk[70]) & (g221) & (!g401)) + ((g2) & (g218) & (g220) & (!sk[70]) & (g221) & (g401)) + ((g2) & (g218) & (g220) & (sk[70]) & (!g221) & (!g401)) + ((g2) & (g218) & (g220) & (sk[70]) & (!g221) & (g401)) + ((g2) & (g218) & (g220) & (sk[70]) & (g221) & (!g401)) + ((g2) & (g218) & (g220) & (sk[70]) & (g221) & (g401)));
	assign g445 = (((!g251) & (!g122) & (!g280) & (!sk[71]) & (g198) & (!g200)) + ((!g251) & (!g122) & (!g280) & (!sk[71]) & (g198) & (g200)) + ((!g251) & (!g122) & (g280) & (!sk[71]) & (!g198) & (!g200)) + ((!g251) & (!g122) & (g280) & (!sk[71]) & (!g198) & (g200)) + ((!g251) & (!g122) & (g280) & (!sk[71]) & (g198) & (!g200)) + ((!g251) & (!g122) & (g280) & (!sk[71]) & (g198) & (g200)) + ((!g251) & (!g122) & (g280) & (sk[71]) & (!g198) & (!g200)) + ((!g251) & (!g122) & (g280) & (sk[71]) & (g198) & (!g200)) + ((!g251) & (g122) & (!g280) & (!sk[71]) & (!g198) & (!g200)) + ((!g251) & (g122) & (!g280) & (!sk[71]) & (!g198) & (g200)) + ((!g251) & (g122) & (!g280) & (!sk[71]) & (g198) & (!g200)) + ((!g251) & (g122) & (!g280) & (!sk[71]) & (g198) & (g200)) + ((!g251) & (g122) & (!g280) & (sk[71]) & (!g198) & (!g200)) + ((!g251) & (g122) & (!g280) & (sk[71]) & (g198) & (!g200)) + ((!g251) & (g122) & (g280) & (!sk[71]) & (!g198) & (!g200)) + ((!g251) & (g122) & (g280) & (!sk[71]) & (!g198) & (g200)) + ((!g251) & (g122) & (g280) & (!sk[71]) & (g198) & (!g200)) + ((!g251) & (g122) & (g280) & (!sk[71]) & (g198) & (g200)) + ((!g251) & (g122) & (g280) & (sk[71]) & (!g198) & (!g200)) + ((!g251) & (g122) & (g280) & (sk[71]) & (!g198) & (g200)) + ((g251) & (!g122) & (!g280) & (!sk[71]) & (g198) & (!g200)) + ((g251) & (!g122) & (!g280) & (!sk[71]) & (g198) & (g200)) + ((g251) & (!g122) & (!g280) & (sk[71]) & (g198) & (!g200)) + ((g251) & (!g122) & (!g280) & (sk[71]) & (g198) & (g200)) + ((g251) & (!g122) & (g280) & (!sk[71]) & (!g198) & (!g200)) + ((g251) & (!g122) & (g280) & (!sk[71]) & (!g198) & (g200)) + ((g251) & (!g122) & (g280) & (!sk[71]) & (g198) & (!g200)) + ((g251) & (!g122) & (g280) & (!sk[71]) & (g198) & (g200)) + ((g251) & (!g122) & (g280) & (sk[71]) & (!g198) & (g200)) + ((g251) & (!g122) & (g280) & (sk[71]) & (g198) & (g200)) + ((g251) & (g122) & (!g280) & (!sk[71]) & (!g198) & (!g200)) + ((g251) & (g122) & (!g280) & (!sk[71]) & (!g198) & (g200)) + ((g251) & (g122) & (!g280) & (!sk[71]) & (g198) & (!g200)) + ((g251) & (g122) & (!g280) & (!sk[71]) & (g198) & (g200)) + ((g251) & (g122) & (!g280) & (sk[71]) & (!g198) & (g200)) + ((g251) & (g122) & (!g280) & (sk[71]) & (g198) & (g200)) + ((g251) & (g122) & (g280) & (!sk[71]) & (!g198) & (!g200)) + ((g251) & (g122) & (g280) & (!sk[71]) & (!g198) & (g200)) + ((g251) & (g122) & (g280) & (!sk[71]) & (g198) & (!g200)) + ((g251) & (g122) & (g280) & (!sk[71]) & (g198) & (g200)));
	assign g446 = (((!sk[72]) & (!g2) & (!g301) & (!g251) & (g302) & (!g367)) + ((!sk[72]) & (!g2) & (!g301) & (!g251) & (g302) & (g367)) + ((!sk[72]) & (!g2) & (!g301) & (g251) & (!g302) & (!g367)) + ((!sk[72]) & (!g2) & (!g301) & (g251) & (!g302) & (g367)) + ((!sk[72]) & (!g2) & (!g301) & (g251) & (g302) & (!g367)) + ((!sk[72]) & (!g2) & (!g301) & (g251) & (g302) & (g367)) + ((!sk[72]) & (!g2) & (g301) & (!g251) & (!g302) & (!g367)) + ((!sk[72]) & (!g2) & (g301) & (!g251) & (!g302) & (g367)) + ((!sk[72]) & (!g2) & (g301) & (!g251) & (g302) & (!g367)) + ((!sk[72]) & (!g2) & (g301) & (!g251) & (g302) & (g367)) + ((!sk[72]) & (!g2) & (g301) & (g251) & (!g302) & (!g367)) + ((!sk[72]) & (!g2) & (g301) & (g251) & (!g302) & (g367)) + ((!sk[72]) & (!g2) & (g301) & (g251) & (g302) & (!g367)) + ((!sk[72]) & (!g2) & (g301) & (g251) & (g302) & (g367)) + ((!sk[72]) & (g2) & (!g301) & (!g251) & (g302) & (!g367)) + ((!sk[72]) & (g2) & (!g301) & (!g251) & (g302) & (g367)) + ((!sk[72]) & (g2) & (!g301) & (g251) & (!g302) & (!g367)) + ((!sk[72]) & (g2) & (!g301) & (g251) & (!g302) & (g367)) + ((!sk[72]) & (g2) & (!g301) & (g251) & (g302) & (!g367)) + ((!sk[72]) & (g2) & (!g301) & (g251) & (g302) & (g367)) + ((!sk[72]) & (g2) & (g301) & (!g251) & (!g302) & (!g367)) + ((!sk[72]) & (g2) & (g301) & (!g251) & (!g302) & (g367)) + ((!sk[72]) & (g2) & (g301) & (!g251) & (g302) & (!g367)) + ((!sk[72]) & (g2) & (g301) & (!g251) & (g302) & (g367)) + ((!sk[72]) & (g2) & (g301) & (g251) & (!g302) & (!g367)) + ((!sk[72]) & (g2) & (g301) & (g251) & (!g302) & (g367)) + ((!sk[72]) & (g2) & (g301) & (g251) & (g302) & (!g367)) + ((!sk[72]) & (g2) & (g301) & (g251) & (g302) & (g367)) + ((sk[72]) & (!g2) & (!g301) & (g251) & (!g302) & (!g367)) + ((sk[72]) & (!g2) & (!g301) & (g251) & (g302) & (g367)) + ((sk[72]) & (!g2) & (g301) & (!g251) & (!g302) & (!g367)) + ((sk[72]) & (!g2) & (g301) & (!g251) & (g302) & (g367)) + ((sk[72]) & (!g2) & (g301) & (g251) & (!g302) & (!g367)) + ((sk[72]) & (!g2) & (g301) & (g251) & (!g302) & (g367)) + ((sk[72]) & (g2) & (!g301) & (!g251) & (g302) & (!g367)) + ((sk[72]) & (g2) & (!g301) & (!g251) & (g302) & (g367)) + ((sk[72]) & (g2) & (!g301) & (g251) & (!g302) & (!g367)) + ((sk[72]) & (g2) & (!g301) & (g251) & (g302) & (g367)) + ((sk[72]) & (g2) & (g301) & (!g251) & (!g302) & (!g367)) + ((sk[72]) & (g2) & (g301) & (!g251) & (g302) & (g367)));
	assign g447 = (((!g305) & (!g122) & (!g222) & (!g159) & (sk[73]) & (g196)) + ((!g305) & (!g122) & (!g222) & (g159) & (!sk[73]) & (!g196)) + ((!g305) & (!g122) & (!g222) & (g159) & (!sk[73]) & (g196)) + ((!g305) & (!g122) & (!g222) & (g159) & (sk[73]) & (!g196)) + ((!g305) & (!g122) & (!g222) & (g159) & (sk[73]) & (g196)) + ((!g305) & (!g122) & (g222) & (!g159) & (!sk[73]) & (!g196)) + ((!g305) & (!g122) & (g222) & (!g159) & (!sk[73]) & (g196)) + ((!g305) & (!g122) & (g222) & (g159) & (!sk[73]) & (!g196)) + ((!g305) & (!g122) & (g222) & (g159) & (!sk[73]) & (g196)) + ((!g305) & (!g122) & (g222) & (g159) & (sk[73]) & (g196)) + ((!g305) & (g122) & (!g222) & (!g159) & (!sk[73]) & (!g196)) + ((!g305) & (g122) & (!g222) & (!g159) & (!sk[73]) & (g196)) + ((!g305) & (g122) & (!g222) & (g159) & (!sk[73]) & (!g196)) + ((!g305) & (g122) & (!g222) & (g159) & (!sk[73]) & (g196)) + ((!g305) & (g122) & (g222) & (!g159) & (!sk[73]) & (!g196)) + ((!g305) & (g122) & (g222) & (!g159) & (!sk[73]) & (g196)) + ((!g305) & (g122) & (g222) & (!g159) & (sk[73]) & (g196)) + ((!g305) & (g122) & (g222) & (g159) & (!sk[73]) & (!g196)) + ((!g305) & (g122) & (g222) & (g159) & (!sk[73]) & (g196)) + ((!g305) & (g122) & (g222) & (g159) & (sk[73]) & (!g196)) + ((g305) & (!g122) & (!g222) & (!g159) & (sk[73]) & (g196)) + ((g305) & (!g122) & (!g222) & (g159) & (!sk[73]) & (!g196)) + ((g305) & (!g122) & (!g222) & (g159) & (!sk[73]) & (g196)) + ((g305) & (!g122) & (!g222) & (g159) & (sk[73]) & (!g196)) + ((g305) & (!g122) & (g222) & (!g159) & (!sk[73]) & (!g196)) + ((g305) & (!g122) & (g222) & (!g159) & (!sk[73]) & (g196)) + ((g305) & (!g122) & (g222) & (g159) & (!sk[73]) & (!g196)) + ((g305) & (!g122) & (g222) & (g159) & (!sk[73]) & (g196)) + ((g305) & (g122) & (!g222) & (!g159) & (!sk[73]) & (!g196)) + ((g305) & (g122) & (!g222) & (!g159) & (!sk[73]) & (g196)) + ((g305) & (g122) & (!g222) & (!g159) & (sk[73]) & (!g196)) + ((g305) & (g122) & (!g222) & (g159) & (!sk[73]) & (!g196)) + ((g305) & (g122) & (!g222) & (g159) & (!sk[73]) & (g196)) + ((g305) & (g122) & (g222) & (!g159) & (!sk[73]) & (!g196)) + ((g305) & (g122) & (g222) & (!g159) & (!sk[73]) & (g196)) + ((g305) & (g122) & (g222) & (!g159) & (sk[73]) & (!g196)) + ((g305) & (g122) & (g222) & (!g159) & (sk[73]) & (g196)) + ((g305) & (g122) & (g222) & (g159) & (!sk[73]) & (!g196)) + ((g305) & (g122) & (g222) & (g159) & (!sk[73]) & (g196)) + ((g305) & (g122) & (g222) & (g159) & (sk[73]) & (!g196)));
	assign g448 = (((!g442) & (!g443) & (g444) & (!g445) & (g446) & (g447)) + ((!g442) & (!g443) & (g444) & (g445) & (!g446) & (g447)) + ((!g442) & (!g443) & (g444) & (g445) & (g446) & (!g447)) + ((!g442) & (!g443) & (g444) & (g445) & (g446) & (g447)) + ((!g442) & (g443) & (g444) & (!g445) & (g446) & (g447)) + ((!g442) & (g443) & (g444) & (g445) & (!g446) & (g447)) + ((!g442) & (g443) & (g444) & (g445) & (g446) & (!g447)) + ((!g442) & (g443) & (g444) & (g445) & (g446) & (g447)) + ((g442) & (!g443) & (g444) & (!g445) & (g446) & (g447)) + ((g442) & (!g443) & (g444) & (g445) & (!g446) & (g447)) + ((g442) & (!g443) & (g444) & (g445) & (g446) & (!g447)) + ((g442) & (!g443) & (g444) & (g445) & (g446) & (g447)) + ((g442) & (g443) & (!g444) & (!g445) & (g446) & (g447)) + ((g442) & (g443) & (!g444) & (g445) & (!g446) & (g447)) + ((g442) & (g443) & (!g444) & (g445) & (g446) & (!g447)) + ((g442) & (g443) & (!g444) & (g445) & (g446) & (g447)) + ((g442) & (g443) & (g444) & (!g445) & (!g446) & (!g447)) + ((g442) & (g443) & (g444) & (!g445) & (!g446) & (g447)) + ((g442) & (g443) & (g444) & (!g445) & (g446) & (!g447)) + ((g442) & (g443) & (g444) & (!g445) & (g446) & (g447)) + ((g442) & (g443) & (g444) & (g445) & (!g446) & (!g447)) + ((g442) & (g443) & (g444) & (g445) & (!g446) & (g447)) + ((g442) & (g443) & (g444) & (g445) & (g446) & (!g447)) + ((g442) & (g443) & (g444) & (g445) & (g446) & (g447)));
	assign g449 = (((!g69) & (!sk[75]) & (!g347) & (!g401) & (g403)) + ((!g69) & (!sk[75]) & (!g347) & (g401) & (g403)) + ((!g69) & (!sk[75]) & (g347) & (!g401) & (g403)) + ((!g69) & (!sk[75]) & (g347) & (g401) & (g403)) + ((!g69) & (sk[75]) & (!g347) & (!g401) & (g403)) + ((!g69) & (sk[75]) & (!g347) & (g401) & (!g403)) + ((!g69) & (sk[75]) & (g347) & (!g401) & (!g403)) + ((!g69) & (sk[75]) & (g347) & (g401) & (g403)) + ((g69) & (!sk[75]) & (!g347) & (!g401) & (!g403)) + ((g69) & (!sk[75]) & (!g347) & (!g401) & (g403)) + ((g69) & (!sk[75]) & (!g347) & (g401) & (!g403)) + ((g69) & (!sk[75]) & (!g347) & (g401) & (g403)) + ((g69) & (!sk[75]) & (g347) & (!g401) & (!g403)) + ((g69) & (!sk[75]) & (g347) & (!g401) & (g403)) + ((g69) & (!sk[75]) & (g347) & (g401) & (!g403)) + ((g69) & (!sk[75]) & (g347) & (g401) & (g403)) + ((g69) & (sk[75]) & (!g347) & (!g401) & (g403)) + ((g69) & (sk[75]) & (!g347) & (g401) & (g403)) + ((g69) & (sk[75]) & (g347) & (!g401) & (!g403)) + ((g69) & (sk[75]) & (g347) & (g401) & (!g403)));
	assign g450 = (((!sk[76]) & (!g406) & (g407) & (!g408)) + ((!sk[76]) & (!g406) & (g407) & (g408)) + ((!sk[76]) & (g406) & (g407) & (!g408)) + ((!sk[76]) & (g406) & (g407) & (g408)) + ((sk[76]) & (!g406) & (!g407) & (!g408)) + ((sk[76]) & (!g406) & (g407) & (g408)) + ((sk[76]) & (g406) & (!g407) & (g408)) + ((sk[76]) & (g406) & (g407) & (!g408)));
	assign g451 = (((!g448) & (!sk[77]) & (g449) & (!g450)) + ((!g448) & (!sk[77]) & (g449) & (g450)) + ((!g448) & (sk[77]) & (!g449) & (!g450)) + ((g448) & (!sk[77]) & (g449) & (!g450)) + ((g448) & (!sk[77]) & (g449) & (g450)) + ((g448) & (sk[77]) & (!g449) & (!g450)) + ((g448) & (sk[77]) & (!g449) & (g450)) + ((g448) & (sk[77]) & (g449) & (!g450)));
	assign g452 = (((!sk[78]) & (!g402) & (!g404) & (!g405) & (g409)) + ((!sk[78]) & (!g402) & (!g404) & (g405) & (g409)) + ((!sk[78]) & (!g402) & (g404) & (!g405) & (g409)) + ((!sk[78]) & (!g402) & (g404) & (g405) & (g409)) + ((!sk[78]) & (g402) & (!g404) & (!g405) & (!g409)) + ((!sk[78]) & (g402) & (!g404) & (!g405) & (g409)) + ((!sk[78]) & (g402) & (!g404) & (g405) & (!g409)) + ((!sk[78]) & (g402) & (!g404) & (g405) & (g409)) + ((!sk[78]) & (g402) & (g404) & (!g405) & (!g409)) + ((!sk[78]) & (g402) & (g404) & (!g405) & (g409)) + ((!sk[78]) & (g402) & (g404) & (g405) & (!g409)) + ((!sk[78]) & (g402) & (g404) & (g405) & (g409)) + ((sk[78]) & (!g402) & (!g404) & (!g405) & (g409)) + ((sk[78]) & (!g402) & (!g404) & (g405) & (!g409)) + ((sk[78]) & (!g402) & (g404) & (!g405) & (!g409)) + ((sk[78]) & (!g402) & (g404) & (g405) & (g409)) + ((sk[78]) & (g402) & (!g404) & (!g405) & (!g409)) + ((sk[78]) & (g402) & (!g404) & (g405) & (g409)) + ((sk[78]) & (g402) & (g404) & (!g405) & (!g409)) + ((sk[78]) & (g402) & (g404) & (g405) & (g409)));
	assign g453 = (((!g426) & (!g429) & (!g430) & (!g434) & (!g435) & (!g436)) + ((!g426) & (!g429) & (!g430) & (!g434) & (g435) & (g436)) + ((!g426) & (!g429) & (!g430) & (g434) & (!g435) & (!g436)) + ((!g426) & (!g429) & (!g430) & (g434) & (g435) & (g436)) + ((!g426) & (!g429) & (g430) & (!g434) & (!g435) & (!g436)) + ((!g426) & (!g429) & (g430) & (!g434) & (g435) & (g436)) + ((!g426) & (!g429) & (g430) & (g434) & (!g435) & (g436)) + ((!g426) & (!g429) & (g430) & (g434) & (g435) & (!g436)) + ((!g426) & (g429) & (!g430) & (!g434) & (!g435) & (!g436)) + ((!g426) & (g429) & (!g430) & (!g434) & (g435) & (g436)) + ((!g426) & (g429) & (!g430) & (g434) & (!g435) & (g436)) + ((!g426) & (g429) & (!g430) & (g434) & (g435) & (!g436)) + ((!g426) & (g429) & (g430) & (!g434) & (!g435) & (g436)) + ((!g426) & (g429) & (g430) & (!g434) & (g435) & (!g436)) + ((!g426) & (g429) & (g430) & (g434) & (!g435) & (g436)) + ((!g426) & (g429) & (g430) & (g434) & (g435) & (!g436)) + ((g426) & (!g429) & (!g430) & (!g434) & (!g435) & (!g436)) + ((g426) & (!g429) & (!g430) & (!g434) & (g435) & (g436)) + ((g426) & (!g429) & (!g430) & (g434) & (!g435) & (g436)) + ((g426) & (!g429) & (!g430) & (g434) & (g435) & (!g436)) + ((g426) & (!g429) & (g430) & (!g434) & (!g435) & (g436)) + ((g426) & (!g429) & (g430) & (!g434) & (g435) & (!g436)) + ((g426) & (!g429) & (g430) & (g434) & (!g435) & (g436)) + ((g426) & (!g429) & (g430) & (g434) & (g435) & (!g436)) + ((g426) & (g429) & (!g430) & (!g434) & (!g435) & (!g436)) + ((g426) & (g429) & (!g430) & (!g434) & (g435) & (g436)) + ((g426) & (g429) & (!g430) & (g434) & (!g435) & (g436)) + ((g426) & (g429) & (!g430) & (g434) & (g435) & (!g436)) + ((g426) & (g429) & (g430) & (!g434) & (!g435) & (g436)) + ((g426) & (g429) & (g430) & (!g434) & (g435) & (!g436)) + ((g426) & (g429) & (g430) & (g434) & (!g435) & (g436)) + ((g426) & (g429) & (g430) & (g434) & (g435) & (!g436)));
	assign g454 = (((!sk[80]) & (!g451) & (g452) & (!g453)) + ((!sk[80]) & (!g451) & (g452) & (g453)) + ((!sk[80]) & (g451) & (g452) & (!g453)) + ((!sk[80]) & (g451) & (g452) & (g453)) + ((sk[80]) & (!g451) & (g452) & (g453)) + ((sk[80]) & (g451) & (!g452) & (g453)) + ((sk[80]) & (g451) & (g452) & (!g453)) + ((sk[80]) & (g451) & (g452) & (g453)));
	assign g455 = (((!g437) & (!sk[81]) & (g438) & (!g439)) + ((!g437) & (!sk[81]) & (g438) & (g439)) + ((!g437) & (sk[81]) & (!g438) & (!g439)) + ((!g437) & (sk[81]) & (g438) & (g439)) + ((g437) & (!sk[81]) & (g438) & (!g439)) + ((g437) & (!sk[81]) & (g438) & (g439)) + ((g437) & (sk[81]) & (!g438) & (g439)) + ((g437) & (sk[81]) & (g438) & (!g439)));
	assign g456 = (((!g218) & (!g220) & (!g221) & (g401) & (!sk[82]) & (!g414)) + ((!g218) & (!g220) & (!g221) & (g401) & (!sk[82]) & (g414)) + ((!g218) & (!g220) & (g221) & (!g401) & (!sk[82]) & (!g414)) + ((!g218) & (!g220) & (g221) & (!g401) & (!sk[82]) & (g414)) + ((!g218) & (!g220) & (g221) & (!g401) & (sk[82]) & (!g414)) + ((!g218) & (!g220) & (g221) & (g401) & (!sk[82]) & (!g414)) + ((!g218) & (!g220) & (g221) & (g401) & (!sk[82]) & (g414)) + ((!g218) & (!g220) & (g221) & (g401) & (sk[82]) & (!g414)) + ((!g218) & (g220) & (!g221) & (!g401) & (!sk[82]) & (!g414)) + ((!g218) & (g220) & (!g221) & (!g401) & (!sk[82]) & (g414)) + ((!g218) & (g220) & (!g221) & (g401) & (!sk[82]) & (!g414)) + ((!g218) & (g220) & (!g221) & (g401) & (!sk[82]) & (g414)) + ((!g218) & (g220) & (g221) & (!g401) & (!sk[82]) & (!g414)) + ((!g218) & (g220) & (g221) & (!g401) & (!sk[82]) & (g414)) + ((!g218) & (g220) & (g221) & (!g401) & (sk[82]) & (!g414)) + ((!g218) & (g220) & (g221) & (!g401) & (sk[82]) & (g414)) + ((!g218) & (g220) & (g221) & (g401) & (!sk[82]) & (!g414)) + ((!g218) & (g220) & (g221) & (g401) & (!sk[82]) & (g414)) + ((g218) & (!g220) & (!g221) & (!g401) & (sk[82]) & (g414)) + ((g218) & (!g220) & (!g221) & (g401) & (!sk[82]) & (!g414)) + ((g218) & (!g220) & (!g221) & (g401) & (!sk[82]) & (g414)) + ((g218) & (!g220) & (!g221) & (g401) & (sk[82]) & (g414)) + ((g218) & (!g220) & (g221) & (!g401) & (!sk[82]) & (!g414)) + ((g218) & (!g220) & (g221) & (!g401) & (!sk[82]) & (g414)) + ((g218) & (!g220) & (g221) & (!g401) & (sk[82]) & (!g414)) + ((g218) & (!g220) & (g221) & (!g401) & (sk[82]) & (g414)) + ((g218) & (!g220) & (g221) & (g401) & (!sk[82]) & (!g414)) + ((g218) & (!g220) & (g221) & (g401) & (!sk[82]) & (g414)) + ((g218) & (!g220) & (g221) & (g401) & (sk[82]) & (!g414)) + ((g218) & (!g220) & (g221) & (g401) & (sk[82]) & (g414)) + ((g218) & (g220) & (!g221) & (!g401) & (!sk[82]) & (!g414)) + ((g218) & (g220) & (!g221) & (!g401) & (!sk[82]) & (g414)) + ((g218) & (g220) & (!g221) & (g401) & (!sk[82]) & (!g414)) + ((g218) & (g220) & (!g221) & (g401) & (!sk[82]) & (g414)) + ((g218) & (g220) & (!g221) & (g401) & (sk[82]) & (!g414)) + ((g218) & (g220) & (!g221) & (g401) & (sk[82]) & (g414)) + ((g218) & (g220) & (g221) & (!g401) & (!sk[82]) & (!g414)) + ((g218) & (g220) & (g221) & (!g401) & (!sk[82]) & (g414)) + ((g218) & (g220) & (g221) & (!g401) & (sk[82]) & (!g414)) + ((g218) & (g220) & (g221) & (!g401) & (sk[82]) & (g414)) + ((g218) & (g220) & (g221) & (g401) & (!sk[82]) & (!g414)) + ((g218) & (g220) & (g221) & (g401) & (!sk[82]) & (g414)) + ((g218) & (g220) & (g221) & (g401) & (sk[82]) & (!g414)) + ((g218) & (g220) & (g221) & (g401) & (sk[82]) & (g414)));
	assign g457 = (((!g202) & (!g303) & (!g196) & (!g347) & (g365) & (!g393)) + ((!g202) & (!g303) & (!g196) & (!g347) & (g365) & (g393)) + ((!g202) & (!g303) & (!g196) & (g347) & (!g365) & (!g393)) + ((!g202) & (!g303) & (!g196) & (g347) & (!g365) & (g393)) + ((!g202) & (!g303) & (!g196) & (g347) & (g365) & (!g393)) + ((!g202) & (!g303) & (!g196) & (g347) & (g365) & (g393)) + ((!g202) & (g303) & (!g196) & (g347) & (g365) & (!g393)) + ((!g202) & (g303) & (!g196) & (g347) & (g365) & (g393)) + ((!g202) & (g303) & (g196) & (!g347) & (g365) & (!g393)) + ((!g202) & (g303) & (g196) & (g347) & (!g365) & (!g393)) + ((g202) & (!g303) & (!g196) & (!g347) & (g365) & (!g393)) + ((g202) & (!g303) & (!g196) & (!g347) & (g365) & (g393)) + ((g202) & (!g303) & (!g196) & (g347) & (!g365) & (!g393)) + ((g202) & (!g303) & (!g196) & (g347) & (!g365) & (g393)) + ((g202) & (!g303) & (g196) & (!g347) & (!g365) & (!g393)) + ((g202) & (!g303) & (g196) & (g347) & (g365) & (!g393)) + ((g202) & (g303) & (g196) & (!g347) & (!g365) & (!g393)) + ((g202) & (g303) & (g196) & (!g347) & (g365) & (!g393)) + ((g202) & (g303) & (g196) & (g347) & (!g365) & (!g393)) + ((g202) & (g303) & (g196) & (g347) & (g365) & (!g393)));
	assign g458 = (((!g442) & (!sk[84]) & (!g443) & (!g456) & (g457)) + ((!g442) & (!sk[84]) & (!g443) & (g456) & (g457)) + ((!g442) & (!sk[84]) & (g443) & (!g456) & (g457)) + ((!g442) & (!sk[84]) & (g443) & (g456) & (g457)) + ((!g442) & (sk[84]) & (!g443) & (g456) & (g457)) + ((!g442) & (sk[84]) & (g443) & (!g456) & (g457)) + ((!g442) & (sk[84]) & (g443) & (g456) & (!g457)) + ((!g442) & (sk[84]) & (g443) & (g456) & (g457)) + ((g442) & (!sk[84]) & (!g443) & (!g456) & (!g457)) + ((g442) & (!sk[84]) & (!g443) & (!g456) & (g457)) + ((g442) & (!sk[84]) & (!g443) & (g456) & (!g457)) + ((g442) & (!sk[84]) & (!g443) & (g456) & (g457)) + ((g442) & (!sk[84]) & (g443) & (!g456) & (!g457)) + ((g442) & (!sk[84]) & (g443) & (!g456) & (g457)) + ((g442) & (!sk[84]) & (g443) & (g456) & (!g457)) + ((g442) & (!sk[84]) & (g443) & (g456) & (g457)) + ((g442) & (sk[84]) & (!g443) & (!g456) & (g457)) + ((g442) & (sk[84]) & (!g443) & (g456) & (!g457)) + ((g442) & (sk[84]) & (!g443) & (g456) & (g457)) + ((g442) & (sk[84]) & (g443) & (g456) & (g457)));
	assign g459 = (((!g431) & (!g432) & (sk[85]) & (!g433)) + ((!g431) & (g432) & (!sk[85]) & (!g433)) + ((!g431) & (g432) & (!sk[85]) & (g433)) + ((!g431) & (g432) & (sk[85]) & (g433)) + ((g431) & (!g432) & (sk[85]) & (g433)) + ((g431) & (g432) & (!sk[85]) & (!g433)) + ((g431) & (g432) & (!sk[85]) & (g433)) + ((g431) & (g432) & (sk[85]) & (!g433)));
	assign g460 = (((!g427) & (!sk[86]) & (!g428) & (!g458) & (g459)) + ((!g427) & (!sk[86]) & (!g428) & (g458) & (g459)) + ((!g427) & (!sk[86]) & (g428) & (!g458) & (g459)) + ((!g427) & (!sk[86]) & (g428) & (g458) & (g459)) + ((!g427) & (sk[86]) & (!g428) & (g458) & (!g459)) + ((!g427) & (sk[86]) & (g428) & (!g458) & (!g459)) + ((!g427) & (sk[86]) & (g428) & (g458) & (!g459)) + ((!g427) & (sk[86]) & (g428) & (g458) & (g459)) + ((g427) & (!sk[86]) & (!g428) & (!g458) & (!g459)) + ((g427) & (!sk[86]) & (!g428) & (!g458) & (g459)) + ((g427) & (!sk[86]) & (!g428) & (g458) & (!g459)) + ((g427) & (!sk[86]) & (!g428) & (g458) & (g459)) + ((g427) & (!sk[86]) & (g428) & (!g458) & (!g459)) + ((g427) & (!sk[86]) & (g428) & (!g458) & (g459)) + ((g427) & (!sk[86]) & (g428) & (g458) & (!g459)) + ((g427) & (!sk[86]) & (g428) & (g458) & (g459)) + ((g427) & (sk[86]) & (!g428) & (!g458) & (!g459)) + ((g427) & (sk[86]) & (!g428) & (g458) & (!g459)) + ((g427) & (sk[86]) & (!g428) & (g458) & (g459)) + ((g427) & (sk[86]) & (g428) & (g458) & (!g459)));
	assign g461 = (((!sk[87]) & (!g426) & (!g429) & (!g430) & (g434)) + ((!sk[87]) & (!g426) & (!g429) & (g430) & (g434)) + ((!sk[87]) & (!g426) & (g429) & (!g430) & (g434)) + ((!sk[87]) & (!g426) & (g429) & (g430) & (g434)) + ((!sk[87]) & (g426) & (!g429) & (!g430) & (!g434)) + ((!sk[87]) & (g426) & (!g429) & (!g430) & (g434)) + ((!sk[87]) & (g426) & (!g429) & (g430) & (!g434)) + ((!sk[87]) & (g426) & (!g429) & (g430) & (g434)) + ((!sk[87]) & (g426) & (g429) & (!g430) & (!g434)) + ((!sk[87]) & (g426) & (g429) & (!g430) & (g434)) + ((!sk[87]) & (g426) & (g429) & (g430) & (!g434)) + ((!sk[87]) & (g426) & (g429) & (g430) & (g434)) + ((sk[87]) & (!g426) & (!g429) & (!g430) & (g434)) + ((sk[87]) & (!g426) & (!g429) & (g430) & (!g434)) + ((sk[87]) & (!g426) & (g429) & (!g430) & (!g434)) + ((sk[87]) & (!g426) & (g429) & (g430) & (g434)) + ((sk[87]) & (g426) & (!g429) & (!g430) & (!g434)) + ((sk[87]) & (g426) & (!g429) & (g430) & (g434)) + ((sk[87]) & (g426) & (g429) & (!g430) & (!g434)) + ((sk[87]) & (g426) & (g429) & (g430) & (g434)));
	assign g462 = (((!sk[88]) & (!g448) & (g449) & (!g450)) + ((!sk[88]) & (!g448) & (g449) & (g450)) + ((!sk[88]) & (g448) & (g449) & (!g450)) + ((!sk[88]) & (g448) & (g449) & (g450)) + ((sk[88]) & (!g448) & (!g449) & (g450)) + ((sk[88]) & (!g448) & (g449) & (!g450)) + ((sk[88]) & (g448) & (!g449) & (!g450)) + ((sk[88]) & (g448) & (g449) & (g450)));
	assign g463 = (((!g460) & (!sk[89]) & (g461) & (!g462)) + ((!g460) & (!sk[89]) & (g461) & (g462)) + ((!g460) & (sk[89]) & (g461) & (g462)) + ((g460) & (!sk[89]) & (g461) & (!g462)) + ((g460) & (!sk[89]) & (g461) & (g462)) + ((g460) & (sk[89]) & (!g461) & (g462)) + ((g460) & (sk[89]) & (g461) & (!g462)) + ((g460) & (sk[89]) & (g461) & (g462)));
	assign g464 = (((!sk[90]) & (!g451) & (g452) & (!g453)) + ((!sk[90]) & (!g451) & (g452) & (g453)) + ((!sk[90]) & (g451) & (g452) & (!g453)) + ((!sk[90]) & (g451) & (g452) & (g453)) + ((sk[90]) & (!g451) & (!g452) & (g453)) + ((sk[90]) & (!g451) & (g452) & (!g453)) + ((sk[90]) & (g451) & (!g452) & (!g453)) + ((sk[90]) & (g451) & (g452) & (g453)));
	assign g465 = (((!g427) & (!g428) & (!g442) & (!g443) & (!g456) & (!g457)) + ((!g427) & (!g428) & (!g442) & (!g443) & (!g456) & (g457)) + ((!g427) & (!g428) & (!g442) & (!g443) & (g456) & (!g457)) + ((!g427) & (!g428) & (!g442) & (g443) & (!g456) & (!g457)) + ((!g427) & (!g428) & (g442) & (!g443) & (!g456) & (!g457)) + ((!g427) & (!g428) & (g442) & (g443) & (!g456) & (!g457)) + ((!g427) & (!g428) & (g442) & (g443) & (!g456) & (g457)) + ((!g427) & (!g428) & (g442) & (g443) & (g456) & (!g457)) + ((!g427) & (g428) & (!g442) & (!g443) & (g456) & (g457)) + ((!g427) & (g428) & (!g442) & (g443) & (!g456) & (g457)) + ((!g427) & (g428) & (!g442) & (g443) & (g456) & (!g457)) + ((!g427) & (g428) & (!g442) & (g443) & (g456) & (g457)) + ((!g427) & (g428) & (g442) & (!g443) & (!g456) & (g457)) + ((!g427) & (g428) & (g442) & (!g443) & (g456) & (!g457)) + ((!g427) & (g428) & (g442) & (!g443) & (g456) & (g457)) + ((!g427) & (g428) & (g442) & (g443) & (g456) & (g457)) + ((g427) & (!g428) & (!g442) & (!g443) & (g456) & (g457)) + ((g427) & (!g428) & (!g442) & (g443) & (!g456) & (g457)) + ((g427) & (!g428) & (!g442) & (g443) & (g456) & (!g457)) + ((g427) & (!g428) & (!g442) & (g443) & (g456) & (g457)) + ((g427) & (!g428) & (g442) & (!g443) & (!g456) & (g457)) + ((g427) & (!g428) & (g442) & (!g443) & (g456) & (!g457)) + ((g427) & (!g428) & (g442) & (!g443) & (g456) & (g457)) + ((g427) & (!g428) & (g442) & (g443) & (g456) & (g457)) + ((g427) & (g428) & (!g442) & (!g443) & (!g456) & (!g457)) + ((g427) & (g428) & (!g442) & (!g443) & (!g456) & (g457)) + ((g427) & (g428) & (!g442) & (!g443) & (g456) & (!g457)) + ((g427) & (g428) & (!g442) & (g443) & (!g456) & (!g457)) + ((g427) & (g428) & (g442) & (!g443) & (!g456) & (!g457)) + ((g427) & (g428) & (g442) & (g443) & (!g456) & (!g457)) + ((g427) & (g428) & (g442) & (g443) & (!g456) & (g457)) + ((g427) & (g428) & (g442) & (g443) & (g456) & (!g457)));
	assign g466 = (((!g301) & (!g251) & (!sk[92]) & (!g302) & (g414)) + ((!g301) & (!g251) & (!sk[92]) & (g302) & (g414)) + ((!g301) & (g251) & (!sk[92]) & (!g302) & (g414)) + ((!g301) & (g251) & (!sk[92]) & (g302) & (g414)) + ((!g301) & (g251) & (sk[92]) & (!g302) & (!g414)) + ((g301) & (!g251) & (!sk[92]) & (!g302) & (!g414)) + ((g301) & (!g251) & (!sk[92]) & (!g302) & (g414)) + ((g301) & (!g251) & (!sk[92]) & (g302) & (!g414)) + ((g301) & (!g251) & (!sk[92]) & (g302) & (g414)) + ((g301) & (!g251) & (sk[92]) & (!g302) & (!g414)) + ((g301) & (g251) & (!sk[92]) & (!g302) & (!g414)) + ((g301) & (g251) & (!sk[92]) & (!g302) & (g414)) + ((g301) & (g251) & (!sk[92]) & (g302) & (!g414)) + ((g301) & (g251) & (!sk[92]) & (g302) & (g414)) + ((g301) & (g251) & (sk[92]) & (!g302) & (!g414)) + ((g301) & (g251) & (sk[92]) & (!g302) & (g414)));
	assign g467 = (((!g202) & (!g303) & (!sk[93]) & (!g347) & (g425)) + ((!g202) & (!g303) & (!sk[93]) & (g347) & (g425)) + ((!g202) & (!g303) & (sk[93]) & (!g347) & (!g425)) + ((!g202) & (!g303) & (sk[93]) & (!g347) & (g425)) + ((!g202) & (g303) & (!sk[93]) & (!g347) & (g425)) + ((!g202) & (g303) & (!sk[93]) & (g347) & (g425)) + ((!g202) & (g303) & (sk[93]) & (!g347) & (g425)) + ((!g202) & (g303) & (sk[93]) & (g347) & (!g425)) + ((g202) & (!g303) & (!sk[93]) & (!g347) & (!g425)) + ((g202) & (!g303) & (!sk[93]) & (!g347) & (g425)) + ((g202) & (!g303) & (!sk[93]) & (g347) & (!g425)) + ((g202) & (!g303) & (!sk[93]) & (g347) & (g425)) + ((g202) & (!g303) & (sk[93]) & (!g347) & (!g425)) + ((g202) & (g303) & (!sk[93]) & (!g347) & (!g425)) + ((g202) & (g303) & (!sk[93]) & (!g347) & (g425)) + ((g202) & (g303) & (!sk[93]) & (g347) & (!g425)) + ((g202) & (g303) & (!sk[93]) & (g347) & (g425)) + ((g202) & (g303) & (sk[93]) & (g347) & (!g425)));
	assign g468 = (((!g305) & (!g122) & (!g159) & (!sk[94]) & (g196) & (!g200)) + ((!g305) & (!g122) & (!g159) & (!sk[94]) & (g196) & (g200)) + ((!g305) & (!g122) & (!g159) & (sk[94]) & (g196) & (!g200)) + ((!g305) & (!g122) & (!g159) & (sk[94]) & (g196) & (g200)) + ((!g305) & (!g122) & (g159) & (!sk[94]) & (!g196) & (!g200)) + ((!g305) & (!g122) & (g159) & (!sk[94]) & (!g196) & (g200)) + ((!g305) & (!g122) & (g159) & (!sk[94]) & (g196) & (!g200)) + ((!g305) & (!g122) & (g159) & (!sk[94]) & (g196) & (g200)) + ((!g305) & (!g122) & (g159) & (sk[94]) & (!g196) & (!g200)) + ((!g305) & (!g122) & (g159) & (sk[94]) & (!g196) & (g200)) + ((!g305) & (!g122) & (g159) & (sk[94]) & (g196) & (!g200)) + ((!g305) & (g122) & (!g159) & (!sk[94]) & (!g196) & (!g200)) + ((!g305) & (g122) & (!g159) & (!sk[94]) & (!g196) & (g200)) + ((!g305) & (g122) & (!g159) & (!sk[94]) & (g196) & (!g200)) + ((!g305) & (g122) & (!g159) & (!sk[94]) & (g196) & (g200)) + ((!g305) & (g122) & (!g159) & (sk[94]) & (!g196) & (g200)) + ((!g305) & (g122) & (g159) & (!sk[94]) & (!g196) & (!g200)) + ((!g305) & (g122) & (g159) & (!sk[94]) & (!g196) & (g200)) + ((!g305) & (g122) & (g159) & (!sk[94]) & (g196) & (!g200)) + ((!g305) & (g122) & (g159) & (!sk[94]) & (g196) & (g200)) + ((g305) & (!g122) & (!g159) & (!sk[94]) & (g196) & (!g200)) + ((g305) & (!g122) & (!g159) & (!sk[94]) & (g196) & (g200)) + ((g305) & (!g122) & (g159) & (!sk[94]) & (!g196) & (!g200)) + ((g305) & (!g122) & (g159) & (!sk[94]) & (!g196) & (g200)) + ((g305) & (!g122) & (g159) & (!sk[94]) & (g196) & (!g200)) + ((g305) & (!g122) & (g159) & (!sk[94]) & (g196) & (g200)) + ((g305) & (!g122) & (g159) & (sk[94]) & (g196) & (!g200)) + ((g305) & (g122) & (!g159) & (!sk[94]) & (!g196) & (!g200)) + ((g305) & (g122) & (!g159) & (!sk[94]) & (!g196) & (g200)) + ((g305) & (g122) & (!g159) & (!sk[94]) & (g196) & (!g200)) + ((g305) & (g122) & (!g159) & (!sk[94]) & (g196) & (g200)) + ((g305) & (g122) & (!g159) & (sk[94]) & (!g196) & (g200)) + ((g305) & (g122) & (!g159) & (sk[94]) & (g196) & (!g200)) + ((g305) & (g122) & (!g159) & (sk[94]) & (g196) & (g200)) + ((g305) & (g122) & (g159) & (!sk[94]) & (!g196) & (!g200)) + ((g305) & (g122) & (g159) & (!sk[94]) & (!g196) & (g200)) + ((g305) & (g122) & (g159) & (!sk[94]) & (g196) & (!g200)) + ((g305) & (g122) & (g159) & (!sk[94]) & (g196) & (g200)) + ((g305) & (g122) & (g159) & (sk[94]) & (!g196) & (!g200)) + ((g305) & (g122) & (g159) & (sk[94]) & (!g196) & (g200)));
	assign g469 = (((!g251) & (!g122) & (!sk[95]) & (!g280) & (g198) & (!g367)) + ((!g251) & (!g122) & (!sk[95]) & (!g280) & (g198) & (g367)) + ((!g251) & (!g122) & (!sk[95]) & (g280) & (!g198) & (!g367)) + ((!g251) & (!g122) & (!sk[95]) & (g280) & (!g198) & (g367)) + ((!g251) & (!g122) & (!sk[95]) & (g280) & (g198) & (!g367)) + ((!g251) & (!g122) & (!sk[95]) & (g280) & (g198) & (g367)) + ((!g251) & (!g122) & (sk[95]) & (g280) & (!g198) & (!g367)) + ((!g251) & (!g122) & (sk[95]) & (g280) & (!g198) & (g367)) + ((!g251) & (g122) & (!sk[95]) & (!g280) & (!g198) & (!g367)) + ((!g251) & (g122) & (!sk[95]) & (!g280) & (!g198) & (g367)) + ((!g251) & (g122) & (!sk[95]) & (!g280) & (g198) & (!g367)) + ((!g251) & (g122) & (!sk[95]) & (!g280) & (g198) & (g367)) + ((!g251) & (g122) & (!sk[95]) & (g280) & (!g198) & (!g367)) + ((!g251) & (g122) & (!sk[95]) & (g280) & (!g198) & (g367)) + ((!g251) & (g122) & (!sk[95]) & (g280) & (g198) & (!g367)) + ((!g251) & (g122) & (!sk[95]) & (g280) & (g198) & (g367)) + ((!g251) & (g122) & (sk[95]) & (!g280) & (!g198) & (!g367)) + ((!g251) & (g122) & (sk[95]) & (!g280) & (!g198) & (g367)) + ((!g251) & (g122) & (sk[95]) & (g280) & (!g198) & (!g367)) + ((!g251) & (g122) & (sk[95]) & (g280) & (g198) & (!g367)) + ((g251) & (!g122) & (!sk[95]) & (!g280) & (g198) & (!g367)) + ((g251) & (!g122) & (!sk[95]) & (!g280) & (g198) & (g367)) + ((g251) & (!g122) & (!sk[95]) & (g280) & (!g198) & (!g367)) + ((g251) & (!g122) & (!sk[95]) & (g280) & (!g198) & (g367)) + ((g251) & (!g122) & (!sk[95]) & (g280) & (g198) & (!g367)) + ((g251) & (!g122) & (!sk[95]) & (g280) & (g198) & (g367)) + ((g251) & (!g122) & (sk[95]) & (!g280) & (!g198) & (g367)) + ((g251) & (!g122) & (sk[95]) & (!g280) & (g198) & (g367)) + ((g251) & (!g122) & (sk[95]) & (g280) & (g198) & (!g367)) + ((g251) & (!g122) & (sk[95]) & (g280) & (g198) & (g367)) + ((g251) & (g122) & (!sk[95]) & (!g280) & (!g198) & (!g367)) + ((g251) & (g122) & (!sk[95]) & (!g280) & (!g198) & (g367)) + ((g251) & (g122) & (!sk[95]) & (!g280) & (g198) & (!g367)) + ((g251) & (g122) & (!sk[95]) & (!g280) & (g198) & (g367)) + ((g251) & (g122) & (!sk[95]) & (g280) & (!g198) & (!g367)) + ((g251) & (g122) & (!sk[95]) & (g280) & (!g198) & (g367)) + ((g251) & (g122) & (!sk[95]) & (g280) & (g198) & (!g367)) + ((g251) & (g122) & (!sk[95]) & (g280) & (g198) & (g367)) + ((g251) & (g122) & (sk[95]) & (!g280) & (g198) & (!g367)) + ((g251) & (g122) & (sk[95]) & (!g280) & (g198) & (g367)));
	assign g470 = (((!g466) & (!sk[96]) & (!g467) & (!g468) & (g469)) + ((!g466) & (!sk[96]) & (!g467) & (g468) & (g469)) + ((!g466) & (!sk[96]) & (g467) & (!g468) & (g469)) + ((!g466) & (!sk[96]) & (g467) & (g468) & (g469)) + ((!g466) & (sk[96]) & (!g467) & (g468) & (g469)) + ((!g466) & (sk[96]) & (g467) & (g468) & (g469)) + ((g466) & (!sk[96]) & (!g467) & (!g468) & (!g469)) + ((g466) & (!sk[96]) & (!g467) & (!g468) & (g469)) + ((g466) & (!sk[96]) & (!g467) & (g468) & (!g469)) + ((g466) & (!sk[96]) & (!g467) & (g468) & (g469)) + ((g466) & (!sk[96]) & (g467) & (!g468) & (!g469)) + ((g466) & (!sk[96]) & (g467) & (!g468) & (g469)) + ((g466) & (!sk[96]) & (g467) & (g468) & (!g469)) + ((g466) & (!sk[96]) & (g467) & (g468) & (g469)) + ((g466) & (sk[96]) & (!g467) & (g468) & (g469)) + ((g466) & (sk[96]) & (g467) & (!g468) & (g469)) + ((g466) & (sk[96]) & (g467) & (g468) & (!g469)) + ((g466) & (sk[96]) & (g467) & (g468) & (g469)));
	assign g471 = (((!g253) & (!g303) & (!g347) & (!sk[97]) & (g425)) + ((!g253) & (!g303) & (!g347) & (sk[97]) & (!g425)) + ((!g253) & (!g303) & (!g347) & (sk[97]) & (g425)) + ((!g253) & (!g303) & (g347) & (!sk[97]) & (g425)) + ((!g253) & (g303) & (!g347) & (!sk[97]) & (g425)) + ((!g253) & (g303) & (!g347) & (sk[97]) & (!g425)) + ((!g253) & (g303) & (g347) & (!sk[97]) & (g425)) + ((g253) & (!g303) & (!g347) & (!sk[97]) & (!g425)) + ((g253) & (!g303) & (!g347) & (!sk[97]) & (g425)) + ((g253) & (!g303) & (!g347) & (sk[97]) & (g425)) + ((g253) & (!g303) & (g347) & (!sk[97]) & (!g425)) + ((g253) & (!g303) & (g347) & (!sk[97]) & (g425)) + ((g253) & (!g303) & (g347) & (sk[97]) & (!g425)) + ((g253) & (g303) & (!g347) & (!sk[97]) & (!g425)) + ((g253) & (g303) & (!g347) & (!sk[97]) & (g425)) + ((g253) & (g303) & (g347) & (!sk[97]) & (!g425)) + ((g253) & (g303) & (g347) & (!sk[97]) & (g425)) + ((g253) & (g303) & (g347) & (sk[97]) & (!g425)));
	assign g472 = (((!g202) & (!g222) & (!g196) & (!g347) & (g365) & (!g393)) + ((!g202) & (!g222) & (!g196) & (!g347) & (g365) & (g393)) + ((!g202) & (!g222) & (!g196) & (g347) & (!g365) & (!g393)) + ((!g202) & (!g222) & (!g196) & (g347) & (!g365) & (g393)) + ((!g202) & (!g222) & (!g196) & (g347) & (g365) & (!g393)) + ((!g202) & (!g222) & (!g196) & (g347) & (g365) & (g393)) + ((!g202) & (g222) & (!g196) & (!g347) & (g365) & (!g393)) + ((!g202) & (g222) & (!g196) & (!g347) & (g365) & (g393)) + ((!g202) & (g222) & (!g196) & (g347) & (!g365) & (!g393)) + ((!g202) & (g222) & (!g196) & (g347) & (!g365) & (g393)) + ((!g202) & (g222) & (g196) & (!g347) & (!g365) & (!g393)) + ((!g202) & (g222) & (g196) & (g347) & (g365) & (!g393)) + ((g202) & (!g222) & (!g196) & (g347) & (g365) & (!g393)) + ((g202) & (!g222) & (!g196) & (g347) & (g365) & (g393)) + ((g202) & (!g222) & (g196) & (!g347) & (g365) & (!g393)) + ((g202) & (!g222) & (g196) & (g347) & (!g365) & (!g393)) + ((g202) & (g222) & (g196) & (!g347) & (!g365) & (!g393)) + ((g202) & (g222) & (g196) & (!g347) & (g365) & (!g393)) + ((g202) & (g222) & (g196) & (g347) & (!g365) & (!g393)) + ((g202) & (g222) & (g196) & (g347) & (g365) & (!g393)));
	assign g473 = (((!g2) & (!g301) & (!g251) & (!sk[99]) & (g302) & (!g401)) + ((!g2) & (!g301) & (!g251) & (!sk[99]) & (g302) & (g401)) + ((!g2) & (!g301) & (!g251) & (sk[99]) & (g302) & (g401)) + ((!g2) & (!g301) & (g251) & (!sk[99]) & (!g302) & (!g401)) + ((!g2) & (!g301) & (g251) & (!sk[99]) & (!g302) & (g401)) + ((!g2) & (!g301) & (g251) & (!sk[99]) & (g302) & (!g401)) + ((!g2) & (!g301) & (g251) & (!sk[99]) & (g302) & (g401)) + ((!g2) & (!g301) & (g251) & (sk[99]) & (!g302) & (!g401)) + ((!g2) & (!g301) & (g251) & (sk[99]) & (!g302) & (g401)) + ((!g2) & (g301) & (!g251) & (!sk[99]) & (!g302) & (!g401)) + ((!g2) & (g301) & (!g251) & (!sk[99]) & (!g302) & (g401)) + ((!g2) & (g301) & (!g251) & (!sk[99]) & (g302) & (!g401)) + ((!g2) & (g301) & (!g251) & (!sk[99]) & (g302) & (g401)) + ((!g2) & (g301) & (!g251) & (sk[99]) & (!g302) & (!g401)) + ((!g2) & (g301) & (!g251) & (sk[99]) & (!g302) & (g401)) + ((!g2) & (g301) & (g251) & (!sk[99]) & (!g302) & (!g401)) + ((!g2) & (g301) & (g251) & (!sk[99]) & (!g302) & (g401)) + ((!g2) & (g301) & (g251) & (!sk[99]) & (g302) & (!g401)) + ((!g2) & (g301) & (g251) & (!sk[99]) & (g302) & (g401)) + ((!g2) & (g301) & (g251) & (sk[99]) & (!g302) & (!g401)) + ((g2) & (!g301) & (!g251) & (!sk[99]) & (g302) & (!g401)) + ((g2) & (!g301) & (!g251) & (!sk[99]) & (g302) & (g401)) + ((g2) & (!g301) & (!g251) & (sk[99]) & (g302) & (g401)) + ((g2) & (!g301) & (g251) & (!sk[99]) & (!g302) & (!g401)) + ((g2) & (!g301) & (g251) & (!sk[99]) & (!g302) & (g401)) + ((g2) & (!g301) & (g251) & (!sk[99]) & (g302) & (!g401)) + ((g2) & (!g301) & (g251) & (!sk[99]) & (g302) & (g401)) + ((g2) & (!g301) & (g251) & (sk[99]) & (g302) & (!g401)) + ((g2) & (!g301) & (g251) & (sk[99]) & (g302) & (g401)) + ((g2) & (g301) & (!g251) & (!sk[99]) & (!g302) & (!g401)) + ((g2) & (g301) & (!g251) & (!sk[99]) & (!g302) & (g401)) + ((g2) & (g301) & (!g251) & (!sk[99]) & (g302) & (!g401)) + ((g2) & (g301) & (!g251) & (!sk[99]) & (g302) & (g401)) + ((g2) & (g301) & (!g251) & (sk[99]) & (g302) & (!g401)) + ((g2) & (g301) & (!g251) & (sk[99]) & (g302) & (g401)) + ((g2) & (g301) & (g251) & (!sk[99]) & (!g302) & (!g401)) + ((g2) & (g301) & (g251) & (!sk[99]) & (!g302) & (g401)) + ((g2) & (g301) & (g251) & (!sk[99]) & (g302) & (!g401)) + ((g2) & (g301) & (g251) & (!sk[99]) & (g302) & (g401)) + ((g2) & (g301) & (g251) & (sk[99]) & (!g302) & (!g401)));
	assign g474 = (((!g471) & (g472) & (!sk[100]) & (!g473)) + ((!g471) & (g472) & (!sk[100]) & (g473)) + ((!g471) & (g472) & (sk[100]) & (g473)) + ((g471) & (!g472) & (sk[100]) & (g473)) + ((g471) & (g472) & (!sk[100]) & (!g473)) + ((g471) & (g472) & (!sk[100]) & (g473)) + ((g471) & (g472) & (sk[100]) & (!g473)) + ((g471) & (g472) & (sk[100]) & (g473)));
	assign g475 = (((!sk[101]) & (!g445) & (g446) & (!g447)) + ((!sk[101]) & (!g445) & (g446) & (g447)) + ((!sk[101]) & (g445) & (g446) & (!g447)) + ((!sk[101]) & (g445) & (g446) & (g447)) + ((sk[101]) & (!g445) & (!g446) & (!g447)) + ((sk[101]) & (!g445) & (g446) & (g447)) + ((sk[101]) & (g445) & (!g446) & (g447)) + ((sk[101]) & (g445) & (g446) & (!g447)));
	assign g476 = (((!g442) & (!g443) & (!g444) & (!g445) & (g446) & (g447)) + ((!g442) & (!g443) & (!g444) & (g445) & (!g446) & (g447)) + ((!g442) & (!g443) & (!g444) & (g445) & (g446) & (!g447)) + ((!g442) & (!g443) & (!g444) & (g445) & (g446) & (g447)) + ((!g442) & (!g443) & (g444) & (!g445) & (!g446) & (!g447)) + ((!g442) & (!g443) & (g444) & (!g445) & (!g446) & (g447)) + ((!g442) & (!g443) & (g444) & (!g445) & (g446) & (!g447)) + ((!g442) & (!g443) & (g444) & (g445) & (!g446) & (!g447)) + ((!g442) & (g443) & (!g444) & (!g445) & (g446) & (g447)) + ((!g442) & (g443) & (!g444) & (g445) & (!g446) & (g447)) + ((!g442) & (g443) & (!g444) & (g445) & (g446) & (!g447)) + ((!g442) & (g443) & (!g444) & (g445) & (g446) & (g447)) + ((!g442) & (g443) & (g444) & (!g445) & (!g446) & (!g447)) + ((!g442) & (g443) & (g444) & (!g445) & (!g446) & (g447)) + ((!g442) & (g443) & (g444) & (!g445) & (g446) & (!g447)) + ((!g442) & (g443) & (g444) & (g445) & (!g446) & (!g447)) + ((g442) & (!g443) & (!g444) & (!g445) & (g446) & (g447)) + ((g442) & (!g443) & (!g444) & (g445) & (!g446) & (g447)) + ((g442) & (!g443) & (!g444) & (g445) & (g446) & (!g447)) + ((g442) & (!g443) & (!g444) & (g445) & (g446) & (g447)) + ((g442) & (!g443) & (g444) & (!g445) & (!g446) & (!g447)) + ((g442) & (!g443) & (g444) & (!g445) & (!g446) & (g447)) + ((g442) & (!g443) & (g444) & (!g445) & (g446) & (!g447)) + ((g442) & (!g443) & (g444) & (g445) & (!g446) & (!g447)) + ((g442) & (g443) & (!g444) & (!g445) & (!g446) & (!g447)) + ((g442) & (g443) & (!g444) & (!g445) & (!g446) & (g447)) + ((g442) & (g443) & (!g444) & (!g445) & (g446) & (!g447)) + ((g442) & (g443) & (!g444) & (g445) & (!g446) & (!g447)) + ((g442) & (g443) & (g444) & (!g445) & (g446) & (g447)) + ((g442) & (g443) & (g444) & (g445) & (!g446) & (g447)) + ((g442) & (g443) & (g444) & (g445) & (g446) & (!g447)) + ((g442) & (g443) & (g444) & (g445) & (g446) & (g447)));
	assign g477 = (((!g459) & (!g465) & (!g470) & (g474) & (!g475) & (g476)) + ((!g459) & (!g465) & (g470) & (!g474) & (!g475) & (g476)) + ((!g459) & (!g465) & (g470) & (g474) & (!g475) & (g476)) + ((!g459) & (!g465) & (g470) & (g474) & (g475) & (g476)) + ((!g459) & (g465) & (!g470) & (!g474) & (!g475) & (g476)) + ((!g459) & (g465) & (!g470) & (!g474) & (g475) & (g476)) + ((!g459) & (g465) & (!g470) & (g474) & (!g475) & (!g476)) + ((!g459) & (g465) & (!g470) & (g474) & (!g475) & (g476)) + ((!g459) & (g465) & (!g470) & (g474) & (g475) & (g476)) + ((!g459) & (g465) & (g470) & (!g474) & (!g475) & (!g476)) + ((!g459) & (g465) & (g470) & (!g474) & (!g475) & (g476)) + ((!g459) & (g465) & (g470) & (!g474) & (g475) & (g476)) + ((!g459) & (g465) & (g470) & (g474) & (!g475) & (!g476)) + ((!g459) & (g465) & (g470) & (g474) & (!g475) & (g476)) + ((!g459) & (g465) & (g470) & (g474) & (g475) & (!g476)) + ((!g459) & (g465) & (g470) & (g474) & (g475) & (g476)) + ((g459) & (!g465) & (!g470) & (!g474) & (!g475) & (g476)) + ((g459) & (!g465) & (!g470) & (!g474) & (g475) & (g476)) + ((g459) & (!g465) & (!g470) & (g474) & (!g475) & (!g476)) + ((g459) & (!g465) & (!g470) & (g474) & (!g475) & (g476)) + ((g459) & (!g465) & (!g470) & (g474) & (g475) & (g476)) + ((g459) & (!g465) & (g470) & (!g474) & (!g475) & (!g476)) + ((g459) & (!g465) & (g470) & (!g474) & (!g475) & (g476)) + ((g459) & (!g465) & (g470) & (!g474) & (g475) & (g476)) + ((g459) & (!g465) & (g470) & (g474) & (!g475) & (!g476)) + ((g459) & (!g465) & (g470) & (g474) & (!g475) & (g476)) + ((g459) & (!g465) & (g470) & (g474) & (g475) & (!g476)) + ((g459) & (!g465) & (g470) & (g474) & (g475) & (g476)) + ((g459) & (g465) & (!g470) & (g474) & (!g475) & (g476)) + ((g459) & (g465) & (g470) & (!g474) & (!g475) & (g476)) + ((g459) & (g465) & (g470) & (g474) & (!g475) & (g476)) + ((g459) & (g465) & (g470) & (g474) & (g475) & (g476)));
	assign g478 = (((!sk[104]) & (!g460) & (g461) & (!g462)) + ((!sk[104]) & (!g460) & (g461) & (g462)) + ((!sk[104]) & (g460) & (g461) & (!g462)) + ((!sk[104]) & (g460) & (g461) & (g462)) + ((sk[104]) & (!g460) & (!g461) & (g462)) + ((sk[104]) & (!g460) & (g461) & (!g462)) + ((sk[104]) & (g460) & (!g461) & (!g462)) + ((sk[104]) & (g460) & (g461) & (g462)));
	assign g479 = (((!sk[105]) & (!g466) & (!g467) & (!g468) & (g469)) + ((!sk[105]) & (!g466) & (!g467) & (g468) & (g469)) + ((!sk[105]) & (!g466) & (g467) & (!g468) & (g469)) + ((!sk[105]) & (!g466) & (g467) & (g468) & (g469)) + ((!sk[105]) & (g466) & (!g467) & (!g468) & (!g469)) + ((!sk[105]) & (g466) & (!g467) & (!g468) & (g469)) + ((!sk[105]) & (g466) & (!g467) & (g468) & (!g469)) + ((!sk[105]) & (g466) & (!g467) & (g468) & (g469)) + ((!sk[105]) & (g466) & (g467) & (!g468) & (!g469)) + ((!sk[105]) & (g466) & (g467) & (!g468) & (g469)) + ((!sk[105]) & (g466) & (g467) & (g468) & (!g469)) + ((!sk[105]) & (g466) & (g467) & (g468) & (g469)) + ((sk[105]) & (!g466) & (!g467) & (!g468) & (!g469)) + ((sk[105]) & (!g466) & (!g467) & (g468) & (g469)) + ((sk[105]) & (!g466) & (g467) & (!g468) & (!g469)) + ((sk[105]) & (!g466) & (g467) & (g468) & (g469)) + ((sk[105]) & (g466) & (!g467) & (!g468) & (!g469)) + ((sk[105]) & (g466) & (!g467) & (g468) & (g469)) + ((sk[105]) & (g466) & (g467) & (!g468) & (g469)) + ((sk[105]) & (g466) & (g467) & (g468) & (!g469)));
	assign g480 = (((!sk[106]) & (!g2) & (!g251) & (!g122) & (g280) & (!g367)) + ((!sk[106]) & (!g2) & (!g251) & (!g122) & (g280) & (g367)) + ((!sk[106]) & (!g2) & (!g251) & (g122) & (!g280) & (!g367)) + ((!sk[106]) & (!g2) & (!g251) & (g122) & (!g280) & (g367)) + ((!sk[106]) & (!g2) & (!g251) & (g122) & (g280) & (!g367)) + ((!sk[106]) & (!g2) & (!g251) & (g122) & (g280) & (g367)) + ((!sk[106]) & (!g2) & (g251) & (!g122) & (!g280) & (!g367)) + ((!sk[106]) & (!g2) & (g251) & (!g122) & (!g280) & (g367)) + ((!sk[106]) & (!g2) & (g251) & (!g122) & (g280) & (!g367)) + ((!sk[106]) & (!g2) & (g251) & (!g122) & (g280) & (g367)) + ((!sk[106]) & (!g2) & (g251) & (g122) & (!g280) & (!g367)) + ((!sk[106]) & (!g2) & (g251) & (g122) & (!g280) & (g367)) + ((!sk[106]) & (!g2) & (g251) & (g122) & (g280) & (!g367)) + ((!sk[106]) & (!g2) & (g251) & (g122) & (g280) & (g367)) + ((!sk[106]) & (g2) & (!g251) & (!g122) & (g280) & (!g367)) + ((!sk[106]) & (g2) & (!g251) & (!g122) & (g280) & (g367)) + ((!sk[106]) & (g2) & (!g251) & (g122) & (!g280) & (!g367)) + ((!sk[106]) & (g2) & (!g251) & (g122) & (!g280) & (g367)) + ((!sk[106]) & (g2) & (!g251) & (g122) & (g280) & (!g367)) + ((!sk[106]) & (g2) & (!g251) & (g122) & (g280) & (g367)) + ((!sk[106]) & (g2) & (g251) & (!g122) & (!g280) & (!g367)) + ((!sk[106]) & (g2) & (g251) & (!g122) & (!g280) & (g367)) + ((!sk[106]) & (g2) & (g251) & (!g122) & (g280) & (!g367)) + ((!sk[106]) & (g2) & (g251) & (!g122) & (g280) & (g367)) + ((!sk[106]) & (g2) & (g251) & (g122) & (!g280) & (!g367)) + ((!sk[106]) & (g2) & (g251) & (g122) & (!g280) & (g367)) + ((!sk[106]) & (g2) & (g251) & (g122) & (g280) & (!g367)) + ((!sk[106]) & (g2) & (g251) & (g122) & (g280) & (g367)) + ((sk[106]) & (!g2) & (!g251) & (!g122) & (g280) & (!g367)) + ((sk[106]) & (!g2) & (!g251) & (g122) & (!g280) & (!g367)) + ((sk[106]) & (!g2) & (!g251) & (g122) & (g280) & (!g367)) + ((sk[106]) & (!g2) & (!g251) & (g122) & (g280) & (g367)) + ((sk[106]) & (!g2) & (g251) & (!g122) & (g280) & (g367)) + ((sk[106]) & (!g2) & (g251) & (g122) & (!g280) & (g367)) + ((sk[106]) & (g2) & (!g251) & (!g122) & (g280) & (!g367)) + ((sk[106]) & (g2) & (!g251) & (g122) & (!g280) & (!g367)) + ((sk[106]) & (g2) & (g251) & (!g122) & (!g280) & (!g367)) + ((sk[106]) & (g2) & (g251) & (!g122) & (!g280) & (g367)) + ((sk[106]) & (g2) & (g251) & (!g122) & (g280) & (g367)) + ((sk[106]) & (g2) & (g251) & (g122) & (!g280) & (g367)));
	assign g481 = (((!g305) & (!g222) & (!g196) & (!g347) & (g365) & (!g393)) + ((!g305) & (!g222) & (!g196) & (!g347) & (g365) & (g393)) + ((!g305) & (!g222) & (!g196) & (g347) & (!g365) & (!g393)) + ((!g305) & (!g222) & (!g196) & (g347) & (!g365) & (g393)) + ((!g305) & (!g222) & (!g196) & (g347) & (g365) & (!g393)) + ((!g305) & (!g222) & (!g196) & (g347) & (g365) & (g393)) + ((!g305) & (g222) & (!g196) & (g347) & (g365) & (!g393)) + ((!g305) & (g222) & (!g196) & (g347) & (g365) & (g393)) + ((!g305) & (g222) & (g196) & (!g347) & (g365) & (!g393)) + ((!g305) & (g222) & (g196) & (g347) & (!g365) & (!g393)) + ((g305) & (!g222) & (!g196) & (!g347) & (g365) & (!g393)) + ((g305) & (!g222) & (!g196) & (!g347) & (g365) & (g393)) + ((g305) & (!g222) & (!g196) & (g347) & (!g365) & (!g393)) + ((g305) & (!g222) & (!g196) & (g347) & (!g365) & (g393)) + ((g305) & (!g222) & (g196) & (!g347) & (!g365) & (!g393)) + ((g305) & (!g222) & (g196) & (g347) & (g365) & (!g393)) + ((g305) & (g222) & (g196) & (!g347) & (!g365) & (!g393)) + ((g305) & (g222) & (g196) & (!g347) & (g365) & (!g393)) + ((g305) & (g222) & (g196) & (g347) & (!g365) & (!g393)) + ((g305) & (g222) & (g196) & (g347) & (g365) & (!g393)));
	assign g482 = (((!sk[108]) & (!g122) & (!g159) & (!g196) & (g198) & (!g200)) + ((!sk[108]) & (!g122) & (!g159) & (!g196) & (g198) & (g200)) + ((!sk[108]) & (!g122) & (!g159) & (g196) & (!g198) & (!g200)) + ((!sk[108]) & (!g122) & (!g159) & (g196) & (!g198) & (g200)) + ((!sk[108]) & (!g122) & (!g159) & (g196) & (g198) & (!g200)) + ((!sk[108]) & (!g122) & (!g159) & (g196) & (g198) & (g200)) + ((!sk[108]) & (!g122) & (g159) & (!g196) & (!g198) & (!g200)) + ((!sk[108]) & (!g122) & (g159) & (!g196) & (!g198) & (g200)) + ((!sk[108]) & (!g122) & (g159) & (!g196) & (g198) & (!g200)) + ((!sk[108]) & (!g122) & (g159) & (!g196) & (g198) & (g200)) + ((!sk[108]) & (!g122) & (g159) & (g196) & (!g198) & (!g200)) + ((!sk[108]) & (!g122) & (g159) & (g196) & (!g198) & (g200)) + ((!sk[108]) & (!g122) & (g159) & (g196) & (g198) & (!g200)) + ((!sk[108]) & (!g122) & (g159) & (g196) & (g198) & (g200)) + ((!sk[108]) & (g122) & (!g159) & (!g196) & (g198) & (!g200)) + ((!sk[108]) & (g122) & (!g159) & (!g196) & (g198) & (g200)) + ((!sk[108]) & (g122) & (!g159) & (g196) & (!g198) & (!g200)) + ((!sk[108]) & (g122) & (!g159) & (g196) & (!g198) & (g200)) + ((!sk[108]) & (g122) & (!g159) & (g196) & (g198) & (!g200)) + ((!sk[108]) & (g122) & (!g159) & (g196) & (g198) & (g200)) + ((!sk[108]) & (g122) & (g159) & (!g196) & (!g198) & (!g200)) + ((!sk[108]) & (g122) & (g159) & (!g196) & (!g198) & (g200)) + ((!sk[108]) & (g122) & (g159) & (!g196) & (g198) & (!g200)) + ((!sk[108]) & (g122) & (g159) & (!g196) & (g198) & (g200)) + ((!sk[108]) & (g122) & (g159) & (g196) & (!g198) & (!g200)) + ((!sk[108]) & (g122) & (g159) & (g196) & (!g198) & (g200)) + ((!sk[108]) & (g122) & (g159) & (g196) & (g198) & (!g200)) + ((!sk[108]) & (g122) & (g159) & (g196) & (g198) & (g200)) + ((sk[108]) & (!g122) & (!g159) & (g196) & (!g198) & (!g200)) + ((sk[108]) & (!g122) & (!g159) & (g196) & (g198) & (!g200)) + ((sk[108]) & (!g122) & (g159) & (!g196) & (!g198) & (!g200)) + ((sk[108]) & (!g122) & (g159) & (!g196) & (g198) & (!g200)) + ((sk[108]) & (!g122) & (g159) & (g196) & (!g198) & (!g200)) + ((sk[108]) & (!g122) & (g159) & (g196) & (!g198) & (g200)) + ((sk[108]) & (g122) & (!g159) & (!g196) & (g198) & (!g200)) + ((sk[108]) & (g122) & (!g159) & (!g196) & (g198) & (g200)) + ((sk[108]) & (g122) & (!g159) & (g196) & (!g198) & (g200)) + ((sk[108]) & (g122) & (!g159) & (g196) & (g198) & (g200)) + ((sk[108]) & (g122) & (g159) & (!g196) & (!g198) & (g200)) + ((sk[108]) & (g122) & (g159) & (!g196) & (g198) & (g200)));
	assign g483 = (((!g480) & (!sk[109]) & (g481) & (!g482)) + ((!g480) & (!sk[109]) & (g481) & (g482)) + ((!g480) & (sk[109]) & (g481) & (g482)) + ((g480) & (!sk[109]) & (g481) & (!g482)) + ((g480) & (!sk[109]) & (g481) & (g482)) + ((g480) & (sk[109]) & (!g481) & (g482)) + ((g480) & (sk[109]) & (g481) & (!g482)) + ((g480) & (sk[109]) & (g481) & (g482)));
	assign g484 = (((!g218) & (!sk[110]) & (!g220) & (!g221) & (g414)) + ((!g218) & (!sk[110]) & (!g220) & (g221) & (g414)) + ((!g218) & (!sk[110]) & (g220) & (!g221) & (g414)) + ((!g218) & (!sk[110]) & (g220) & (g221) & (g414)) + ((!g218) & (sk[110]) & (g220) & (g221) & (g414)) + ((g218) & (!sk[110]) & (!g220) & (!g221) & (!g414)) + ((g218) & (!sk[110]) & (!g220) & (!g221) & (g414)) + ((g218) & (!sk[110]) & (!g220) & (g221) & (!g414)) + ((g218) & (!sk[110]) & (!g220) & (g221) & (g414)) + ((g218) & (!sk[110]) & (g220) & (!g221) & (!g414)) + ((g218) & (!sk[110]) & (g220) & (!g221) & (g414)) + ((g218) & (!sk[110]) & (g220) & (g221) & (!g414)) + ((g218) & (!sk[110]) & (g220) & (g221) & (g414)) + ((g218) & (sk[110]) & (g220) & (!g221) & (g414)));
	assign g485 = (((!sk[111]) & (!g479) & (g483) & (!g484)) + ((!sk[111]) & (!g479) & (g483) & (g484)) + ((!sk[111]) & (g479) & (g483) & (!g484)) + ((!sk[111]) & (g479) & (g483) & (g484)) + ((sk[111]) & (!g479) & (!g483) & (g484)) + ((sk[111]) & (!g479) & (g483) & (!g484)) + ((sk[111]) & (!g479) & (g483) & (g484)) + ((sk[111]) & (g479) & (g483) & (g484)));
	assign g486 = (((!g442) & (!g443) & (!sk[112]) & (!g456) & (g457)) + ((!g442) & (!g443) & (!sk[112]) & (g456) & (g457)) + ((!g442) & (!g443) & (sk[112]) & (!g456) & (!g457)) + ((!g442) & (!g443) & (sk[112]) & (g456) & (g457)) + ((!g442) & (g443) & (!sk[112]) & (!g456) & (g457)) + ((!g442) & (g443) & (!sk[112]) & (g456) & (g457)) + ((!g442) & (g443) & (sk[112]) & (!g456) & (g457)) + ((!g442) & (g443) & (sk[112]) & (g456) & (!g457)) + ((g442) & (!g443) & (!sk[112]) & (!g456) & (!g457)) + ((g442) & (!g443) & (!sk[112]) & (!g456) & (g457)) + ((g442) & (!g443) & (!sk[112]) & (g456) & (!g457)) + ((g442) & (!g443) & (!sk[112]) & (g456) & (g457)) + ((g442) & (!g443) & (sk[112]) & (!g456) & (g457)) + ((g442) & (!g443) & (sk[112]) & (g456) & (!g457)) + ((g442) & (g443) & (!sk[112]) & (!g456) & (!g457)) + ((g442) & (g443) & (!sk[112]) & (!g456) & (g457)) + ((g442) & (g443) & (!sk[112]) & (g456) & (!g457)) + ((g442) & (g443) & (!sk[112]) & (g456) & (g457)) + ((g442) & (g443) & (sk[112]) & (!g456) & (!g457)) + ((g442) & (g443) & (sk[112]) & (g456) & (g457)));
	assign g487 = (((!g470) & (!g474) & (sk[113]) & (g475)) + ((!g470) & (g474) & (!sk[113]) & (!g475)) + ((!g470) & (g474) & (!sk[113]) & (g475)) + ((!g470) & (g474) & (sk[113]) & (!g475)) + ((g470) & (!g474) & (sk[113]) & (!g475)) + ((g470) & (g474) & (!sk[113]) & (!g475)) + ((g470) & (g474) & (!sk[113]) & (g475)) + ((g470) & (g474) & (sk[113]) & (g475)));
	assign g488 = (((!g459) & (!g465) & (!g470) & (!g474) & (!g475) & (g476)) + ((!g459) & (!g465) & (!g470) & (!g474) & (g475) & (g476)) + ((!g459) & (!g465) & (!g470) & (g474) & (!g475) & (!g476)) + ((!g459) & (!g465) & (!g470) & (g474) & (g475) & (g476)) + ((!g459) & (!g465) & (g470) & (!g474) & (!g475) & (!g476)) + ((!g459) & (!g465) & (g470) & (!g474) & (g475) & (g476)) + ((!g459) & (!g465) & (g470) & (g474) & (!g475) & (!g476)) + ((!g459) & (!g465) & (g470) & (g474) & (g475) & (!g476)) + ((!g459) & (g465) & (!g470) & (!g474) & (!g475) & (!g476)) + ((!g459) & (g465) & (!g470) & (!g474) & (g475) & (!g476)) + ((!g459) & (g465) & (!g470) & (g474) & (!g475) & (g476)) + ((!g459) & (g465) & (!g470) & (g474) & (g475) & (!g476)) + ((!g459) & (g465) & (g470) & (!g474) & (!g475) & (g476)) + ((!g459) & (g465) & (g470) & (!g474) & (g475) & (!g476)) + ((!g459) & (g465) & (g470) & (g474) & (!g475) & (g476)) + ((!g459) & (g465) & (g470) & (g474) & (g475) & (g476)) + ((g459) & (!g465) & (!g470) & (!g474) & (!g475) & (!g476)) + ((g459) & (!g465) & (!g470) & (!g474) & (g475) & (!g476)) + ((g459) & (!g465) & (!g470) & (g474) & (!g475) & (g476)) + ((g459) & (!g465) & (!g470) & (g474) & (g475) & (!g476)) + ((g459) & (!g465) & (g470) & (!g474) & (!g475) & (g476)) + ((g459) & (!g465) & (g470) & (!g474) & (g475) & (!g476)) + ((g459) & (!g465) & (g470) & (g474) & (!g475) & (g476)) + ((g459) & (!g465) & (g470) & (g474) & (g475) & (g476)) + ((g459) & (g465) & (!g470) & (!g474) & (!g475) & (g476)) + ((g459) & (g465) & (!g470) & (!g474) & (g475) & (g476)) + ((g459) & (g465) & (!g470) & (g474) & (!g475) & (!g476)) + ((g459) & (g465) & (!g470) & (g474) & (g475) & (g476)) + ((g459) & (g465) & (g470) & (!g474) & (!g475) & (!g476)) + ((g459) & (g465) & (g470) & (!g474) & (g475) & (g476)) + ((g459) & (g465) & (g470) & (g474) & (!g475) & (!g476)) + ((g459) & (g465) & (g470) & (g474) & (g475) & (!g476)));
	assign g489 = (((!g485) & (!sk[115]) & (!g486) & (!g487) & (g488)) + ((!g485) & (!sk[115]) & (!g486) & (g487) & (g488)) + ((!g485) & (!sk[115]) & (g486) & (!g487) & (g488)) + ((!g485) & (!sk[115]) & (g486) & (g487) & (g488)) + ((!g485) & (sk[115]) & (!g486) & (!g487) & (g488)) + ((g485) & (!sk[115]) & (!g486) & (!g487) & (!g488)) + ((g485) & (!sk[115]) & (!g486) & (!g487) & (g488)) + ((g485) & (!sk[115]) & (!g486) & (g487) & (!g488)) + ((g485) & (!sk[115]) & (!g486) & (g487) & (g488)) + ((g485) & (!sk[115]) & (g486) & (!g487) & (!g488)) + ((g485) & (!sk[115]) & (g486) & (!g487) & (g488)) + ((g485) & (!sk[115]) & (g486) & (g487) & (!g488)) + ((g485) & (!sk[115]) & (g486) & (g487) & (g488)) + ((g485) & (sk[115]) & (!g486) & (!g487) & (g488)) + ((g485) & (sk[115]) & (!g486) & (g487) & (g488)) + ((g485) & (sk[115]) & (g486) & (!g487) & (g488)));
	assign g490 = (((!sk[116]) & (!g485) & (!g486) & (!g487) & (g488)) + ((!sk[116]) & (!g485) & (!g486) & (g487) & (g488)) + ((!sk[116]) & (!g485) & (g486) & (!g487) & (g488)) + ((!sk[116]) & (!g485) & (g486) & (g487) & (g488)) + ((!sk[116]) & (g485) & (!g486) & (!g487) & (!g488)) + ((!sk[116]) & (g485) & (!g486) & (!g487) & (g488)) + ((!sk[116]) & (g485) & (!g486) & (g487) & (!g488)) + ((!sk[116]) & (g485) & (!g486) & (g487) & (g488)) + ((!sk[116]) & (g485) & (g486) & (!g487) & (!g488)) + ((!sk[116]) & (g485) & (g486) & (!g487) & (g488)) + ((!sk[116]) & (g485) & (g486) & (g487) & (!g488)) + ((!sk[116]) & (g485) & (g486) & (g487) & (g488)) + ((sk[116]) & (!g485) & (!g486) & (!g487) & (!g488)) + ((sk[116]) & (!g485) & (!g486) & (g487) & (g488)) + ((sk[116]) & (!g485) & (g486) & (!g487) & (g488)) + ((sk[116]) & (!g485) & (g486) & (g487) & (g488)) + ((sk[116]) & (g485) & (!g486) & (!g487) & (!g488)) + ((sk[116]) & (g485) & (!g486) & (g487) & (!g488)) + ((sk[116]) & (g485) & (g486) & (!g487) & (!g488)) + ((sk[116]) & (g485) & (g486) & (g487) & (g488)));
	assign g491 = (((!g480) & (sk[117]) & (g481)) + ((g480) & (!sk[117]) & (g481)) + ((g480) & (sk[117]) & (!g481)));
	assign g492 = (((!g301) & (sk[118]) & (g251)) + ((g301) & (!sk[118]) & (g251)) + ((g301) & (sk[118]) & (!g251)));
	assign g493 = (((!g251) & (!sk[119]) & (!g122) & (!g280) & (g414)) + ((!g251) & (!sk[119]) & (!g122) & (g280) & (g414)) + ((!g251) & (!sk[119]) & (g122) & (!g280) & (g414)) + ((!g251) & (!sk[119]) & (g122) & (g280) & (g414)) + ((!g251) & (sk[119]) & (!g122) & (g280) & (!g414)) + ((!g251) & (sk[119]) & (g122) & (!g280) & (!g414)) + ((!g251) & (sk[119]) & (g122) & (g280) & (!g414)) + ((!g251) & (sk[119]) & (g122) & (g280) & (g414)) + ((g251) & (!sk[119]) & (!g122) & (!g280) & (!g414)) + ((g251) & (!sk[119]) & (!g122) & (!g280) & (g414)) + ((g251) & (!sk[119]) & (!g122) & (g280) & (!g414)) + ((g251) & (!sk[119]) & (!g122) & (g280) & (g414)) + ((g251) & (!sk[119]) & (g122) & (!g280) & (!g414)) + ((g251) & (!sk[119]) & (g122) & (!g280) & (g414)) + ((g251) & (!sk[119]) & (g122) & (g280) & (!g414)) + ((g251) & (!sk[119]) & (g122) & (g280) & (g414)));
	assign g494 = (((!sk[120]) & (!g305) & (!g222) & (!g347) & (g425)) + ((!sk[120]) & (!g305) & (!g222) & (g347) & (g425)) + ((!sk[120]) & (!g305) & (g222) & (!g347) & (g425)) + ((!sk[120]) & (!g305) & (g222) & (g347) & (g425)) + ((!sk[120]) & (g305) & (!g222) & (!g347) & (!g425)) + ((!sk[120]) & (g305) & (!g222) & (!g347) & (g425)) + ((!sk[120]) & (g305) & (!g222) & (g347) & (!g425)) + ((!sk[120]) & (g305) & (!g222) & (g347) & (g425)) + ((!sk[120]) & (g305) & (g222) & (!g347) & (!g425)) + ((!sk[120]) & (g305) & (g222) & (!g347) & (g425)) + ((!sk[120]) & (g305) & (g222) & (g347) & (!g425)) + ((!sk[120]) & (g305) & (g222) & (g347) & (g425)) + ((sk[120]) & (!g305) & (!g222) & (!g347) & (!g425)) + ((sk[120]) & (!g305) & (!g222) & (!g347) & (g425)) + ((sk[120]) & (!g305) & (g222) & (!g347) & (g425)) + ((sk[120]) & (!g305) & (g222) & (g347) & (!g425)) + ((sk[120]) & (g305) & (!g222) & (!g347) & (!g425)) + ((sk[120]) & (g305) & (g222) & (g347) & (!g425)));
	assign g495 = (((!g2) & (!g251) & (!sk[121]) & (!g122) & (g280) & (!g401)) + ((!g2) & (!g251) & (!sk[121]) & (!g122) & (g280) & (g401)) + ((!g2) & (!g251) & (!sk[121]) & (g122) & (!g280) & (!g401)) + ((!g2) & (!g251) & (!sk[121]) & (g122) & (!g280) & (g401)) + ((!g2) & (!g251) & (!sk[121]) & (g122) & (g280) & (!g401)) + ((!g2) & (!g251) & (!sk[121]) & (g122) & (g280) & (g401)) + ((!g2) & (!g251) & (sk[121]) & (!g122) & (g280) & (!g401)) + ((!g2) & (!g251) & (sk[121]) & (!g122) & (g280) & (g401)) + ((!g2) & (!g251) & (sk[121]) & (g122) & (!g280) & (!g401)) + ((!g2) & (!g251) & (sk[121]) & (g122) & (!g280) & (g401)) + ((!g2) & (!g251) & (sk[121]) & (g122) & (g280) & (!g401)) + ((!g2) & (g251) & (!sk[121]) & (!g122) & (!g280) & (!g401)) + ((!g2) & (g251) & (!sk[121]) & (!g122) & (!g280) & (g401)) + ((!g2) & (g251) & (!sk[121]) & (!g122) & (g280) & (!g401)) + ((!g2) & (g251) & (!sk[121]) & (!g122) & (g280) & (g401)) + ((!g2) & (g251) & (!sk[121]) & (g122) & (!g280) & (!g401)) + ((!g2) & (g251) & (!sk[121]) & (g122) & (!g280) & (g401)) + ((!g2) & (g251) & (!sk[121]) & (g122) & (g280) & (!g401)) + ((!g2) & (g251) & (!sk[121]) & (g122) & (g280) & (g401)) + ((!g2) & (g251) & (sk[121]) & (!g122) & (!g280) & (g401)) + ((g2) & (!g251) & (!sk[121]) & (!g122) & (g280) & (!g401)) + ((g2) & (!g251) & (!sk[121]) & (!g122) & (g280) & (g401)) + ((g2) & (!g251) & (!sk[121]) & (g122) & (!g280) & (!g401)) + ((g2) & (!g251) & (!sk[121]) & (g122) & (!g280) & (g401)) + ((g2) & (!g251) & (!sk[121]) & (g122) & (g280) & (!g401)) + ((g2) & (!g251) & (!sk[121]) & (g122) & (g280) & (g401)) + ((g2) & (!g251) & (sk[121]) & (g122) & (g280) & (!g401)) + ((g2) & (g251) & (!sk[121]) & (!g122) & (!g280) & (!g401)) + ((g2) & (g251) & (!sk[121]) & (!g122) & (!g280) & (g401)) + ((g2) & (g251) & (!sk[121]) & (!g122) & (g280) & (!g401)) + ((g2) & (g251) & (!sk[121]) & (!g122) & (g280) & (g401)) + ((g2) & (g251) & (!sk[121]) & (g122) & (!g280) & (!g401)) + ((g2) & (g251) & (!sk[121]) & (g122) & (!g280) & (g401)) + ((g2) & (g251) & (!sk[121]) & (g122) & (g280) & (!g401)) + ((g2) & (g251) & (!sk[121]) & (g122) & (g280) & (g401)) + ((g2) & (g251) & (sk[121]) & (!g122) & (!g280) & (g401)) + ((g2) & (g251) & (sk[121]) & (!g122) & (g280) & (!g401)) + ((g2) & (g251) & (sk[121]) & (!g122) & (g280) & (g401)) + ((g2) & (g251) & (sk[121]) & (g122) & (!g280) & (!g401)) + ((g2) & (g251) & (sk[121]) & (g122) & (!g280) & (g401)));
	assign g496 = (((!g492) & (!g414) & (!sk[122]) & (!g493) & (g494) & (!g495)) + ((!g492) & (!g414) & (!sk[122]) & (!g493) & (g494) & (g495)) + ((!g492) & (!g414) & (!sk[122]) & (g493) & (!g494) & (!g495)) + ((!g492) & (!g414) & (!sk[122]) & (g493) & (!g494) & (g495)) + ((!g492) & (!g414) & (!sk[122]) & (g493) & (g494) & (!g495)) + ((!g492) & (!g414) & (!sk[122]) & (g493) & (g494) & (g495)) + ((!g492) & (!g414) & (sk[122]) & (g493) & (g494) & (g495)) + ((!g492) & (g414) & (!sk[122]) & (!g493) & (!g494) & (!g495)) + ((!g492) & (g414) & (!sk[122]) & (!g493) & (!g494) & (g495)) + ((!g492) & (g414) & (!sk[122]) & (!g493) & (g494) & (!g495)) + ((!g492) & (g414) & (!sk[122]) & (!g493) & (g494) & (g495)) + ((!g492) & (g414) & (!sk[122]) & (g493) & (!g494) & (!g495)) + ((!g492) & (g414) & (!sk[122]) & (g493) & (!g494) & (g495)) + ((!g492) & (g414) & (!sk[122]) & (g493) & (g494) & (!g495)) + ((!g492) & (g414) & (!sk[122]) & (g493) & (g494) & (g495)) + ((!g492) & (g414) & (sk[122]) & (g493) & (g494) & (g495)) + ((g492) & (!g414) & (!sk[122]) & (!g493) & (g494) & (!g495)) + ((g492) & (!g414) & (!sk[122]) & (!g493) & (g494) & (g495)) + ((g492) & (!g414) & (!sk[122]) & (g493) & (!g494) & (!g495)) + ((g492) & (!g414) & (!sk[122]) & (g493) & (!g494) & (g495)) + ((g492) & (!g414) & (!sk[122]) & (g493) & (g494) & (!g495)) + ((g492) & (!g414) & (!sk[122]) & (g493) & (g494) & (g495)) + ((g492) & (!g414) & (sk[122]) & (g493) & (g494) & (g495)) + ((g492) & (g414) & (!sk[122]) & (!g493) & (!g494) & (!g495)) + ((g492) & (g414) & (!sk[122]) & (!g493) & (!g494) & (g495)) + ((g492) & (g414) & (!sk[122]) & (!g493) & (g494) & (!g495)) + ((g492) & (g414) & (!sk[122]) & (!g493) & (g494) & (g495)) + ((g492) & (g414) & (!sk[122]) & (g493) & (!g494) & (!g495)) + ((g492) & (g414) & (!sk[122]) & (g493) & (!g494) & (g495)) + ((g492) & (g414) & (!sk[122]) & (g493) & (g494) & (!g495)) + ((g492) & (g414) & (!sk[122]) & (g493) & (g494) & (g495)) + ((g492) & (g414) & (sk[122]) & (!g493) & (!g494) & (g495)) + ((g492) & (g414) & (sk[122]) & (!g493) & (g494) & (g495)) + ((g492) & (g414) & (sk[122]) & (g493) & (!g494) & (g495)) + ((g492) & (g414) & (sk[122]) & (g493) & (g494) & (!g495)) + ((g492) & (g414) & (sk[122]) & (g493) & (g494) & (g495)));
	assign g497 = (((!sk[123]) & (!g202) & (!g222) & (!g347) & (g425)) + ((!sk[123]) & (!g202) & (!g222) & (g347) & (g425)) + ((!sk[123]) & (!g202) & (g222) & (!g347) & (g425)) + ((!sk[123]) & (!g202) & (g222) & (g347) & (g425)) + ((!sk[123]) & (g202) & (!g222) & (!g347) & (!g425)) + ((!sk[123]) & (g202) & (!g222) & (!g347) & (g425)) + ((!sk[123]) & (g202) & (!g222) & (g347) & (!g425)) + ((!sk[123]) & (g202) & (!g222) & (g347) & (g425)) + ((!sk[123]) & (g202) & (g222) & (!g347) & (!g425)) + ((!sk[123]) & (g202) & (g222) & (!g347) & (g425)) + ((!sk[123]) & (g202) & (g222) & (g347) & (!g425)) + ((!sk[123]) & (g202) & (g222) & (g347) & (g425)) + ((sk[123]) & (!g202) & (!g222) & (!g347) & (!g425)) + ((sk[123]) & (!g202) & (!g222) & (!g347) & (g425)) + ((sk[123]) & (!g202) & (g222) & (!g347) & (!g425)) + ((sk[123]) & (g202) & (!g222) & (!g347) & (g425)) + ((sk[123]) & (g202) & (!g222) & (g347) & (!g425)) + ((sk[123]) & (g202) & (g222) & (g347) & (!g425)));
	assign g498 = (((!g305) & (!g196) & (!g200) & (!g347) & (g365) & (!g393)) + ((!g305) & (!g196) & (!g200) & (!g347) & (g365) & (g393)) + ((!g305) & (!g196) & (!g200) & (g347) & (!g365) & (!g393)) + ((!g305) & (!g196) & (!g200) & (g347) & (!g365) & (g393)) + ((!g305) & (!g196) & (!g200) & (g347) & (g365) & (!g393)) + ((!g305) & (!g196) & (!g200) & (g347) & (g365) & (g393)) + ((!g305) & (!g196) & (g200) & (!g347) & (g365) & (!g393)) + ((!g305) & (!g196) & (g200) & (!g347) & (g365) & (g393)) + ((!g305) & (!g196) & (g200) & (g347) & (!g365) & (!g393)) + ((!g305) & (!g196) & (g200) & (g347) & (!g365) & (g393)) + ((!g305) & (g196) & (g200) & (!g347) & (!g365) & (!g393)) + ((!g305) & (g196) & (g200) & (g347) & (g365) & (!g393)) + ((g305) & (!g196) & (!g200) & (g347) & (g365) & (!g393)) + ((g305) & (!g196) & (!g200) & (g347) & (g365) & (g393)) + ((g305) & (g196) & (!g200) & (!g347) & (g365) & (!g393)) + ((g305) & (g196) & (!g200) & (g347) & (!g365) & (!g393)) + ((g305) & (g196) & (g200) & (!g347) & (!g365) & (!g393)) + ((g305) & (g196) & (g200) & (!g347) & (g365) & (!g393)) + ((g305) & (g196) & (g200) & (g347) & (!g365) & (!g393)) + ((g305) & (g196) & (g200) & (g347) & (g365) & (!g393)));
	assign g499 = (((!g122) & (!g159) & (!sk[125]) & (!g196) & (g198) & (!g367)) + ((!g122) & (!g159) & (!sk[125]) & (!g196) & (g198) & (g367)) + ((!g122) & (!g159) & (!sk[125]) & (g196) & (!g198) & (!g367)) + ((!g122) & (!g159) & (!sk[125]) & (g196) & (!g198) & (g367)) + ((!g122) & (!g159) & (!sk[125]) & (g196) & (g198) & (!g367)) + ((!g122) & (!g159) & (!sk[125]) & (g196) & (g198) & (g367)) + ((!g122) & (!g159) & (sk[125]) & (g196) & (!g198) & (!g367)) + ((!g122) & (!g159) & (sk[125]) & (g196) & (!g198) & (g367)) + ((!g122) & (g159) & (!sk[125]) & (!g196) & (!g198) & (!g367)) + ((!g122) & (g159) & (!sk[125]) & (!g196) & (!g198) & (g367)) + ((!g122) & (g159) & (!sk[125]) & (!g196) & (g198) & (!g367)) + ((!g122) & (g159) & (!sk[125]) & (!g196) & (g198) & (g367)) + ((!g122) & (g159) & (!sk[125]) & (g196) & (!g198) & (!g367)) + ((!g122) & (g159) & (!sk[125]) & (g196) & (!g198) & (g367)) + ((!g122) & (g159) & (!sk[125]) & (g196) & (g198) & (!g367)) + ((!g122) & (g159) & (!sk[125]) & (g196) & (g198) & (g367)) + ((!g122) & (g159) & (sk[125]) & (!g196) & (!g198) & (!g367)) + ((!g122) & (g159) & (sk[125]) & (!g196) & (!g198) & (g367)) + ((!g122) & (g159) & (sk[125]) & (g196) & (!g198) & (!g367)) + ((!g122) & (g159) & (sk[125]) & (g196) & (g198) & (!g367)) + ((g122) & (!g159) & (!sk[125]) & (!g196) & (g198) & (!g367)) + ((g122) & (!g159) & (!sk[125]) & (!g196) & (g198) & (g367)) + ((g122) & (!g159) & (!sk[125]) & (g196) & (!g198) & (!g367)) + ((g122) & (!g159) & (!sk[125]) & (g196) & (!g198) & (g367)) + ((g122) & (!g159) & (!sk[125]) & (g196) & (g198) & (!g367)) + ((g122) & (!g159) & (!sk[125]) & (g196) & (g198) & (g367)) + ((g122) & (!g159) & (sk[125]) & (!g196) & (!g198) & (g367)) + ((g122) & (!g159) & (sk[125]) & (!g196) & (g198) & (g367)) + ((g122) & (!g159) & (sk[125]) & (g196) & (g198) & (!g367)) + ((g122) & (!g159) & (sk[125]) & (g196) & (g198) & (g367)) + ((g122) & (g159) & (!sk[125]) & (!g196) & (!g198) & (!g367)) + ((g122) & (g159) & (!sk[125]) & (!g196) & (!g198) & (g367)) + ((g122) & (g159) & (!sk[125]) & (!g196) & (g198) & (!g367)) + ((g122) & (g159) & (!sk[125]) & (!g196) & (g198) & (g367)) + ((g122) & (g159) & (!sk[125]) & (g196) & (!g198) & (!g367)) + ((g122) & (g159) & (!sk[125]) & (g196) & (!g198) & (g367)) + ((g122) & (g159) & (!sk[125]) & (g196) & (g198) & (!g367)) + ((g122) & (g159) & (!sk[125]) & (g196) & (g198) & (g367)) + ((g122) & (g159) & (sk[125]) & (!g196) & (g198) & (!g367)) + ((g122) & (g159) & (sk[125]) & (!g196) & (g198) & (g367)));
	assign g500 = (((!g497) & (!sk[126]) & (g498) & (!g499)) + ((!g497) & (!sk[126]) & (g498) & (g499)) + ((!g497) & (sk[126]) & (g498) & (g499)) + ((g497) & (!sk[126]) & (g498) & (!g499)) + ((g497) & (!sk[126]) & (g498) & (g499)) + ((g497) & (sk[126]) & (!g498) & (g499)) + ((g497) & (sk[126]) & (g498) & (!g499)) + ((g497) & (sk[126]) & (g498) & (g499)));
	assign g501 = (((!g301) & (!g251) & (!g302) & (!sk[127]) & (g401) & (!g414)) + ((!g301) & (!g251) & (!g302) & (!sk[127]) & (g401) & (g414)) + ((!g301) & (!g251) & (g302) & (!sk[127]) & (!g401) & (!g414)) + ((!g301) & (!g251) & (g302) & (!sk[127]) & (!g401) & (g414)) + ((!g301) & (!g251) & (g302) & (!sk[127]) & (g401) & (!g414)) + ((!g301) & (!g251) & (g302) & (!sk[127]) & (g401) & (g414)) + ((!g301) & (!g251) & (g302) & (sk[127]) & (!g401) & (g414)) + ((!g301) & (!g251) & (g302) & (sk[127]) & (g401) & (g414)) + ((!g301) & (g251) & (!g302) & (!sk[127]) & (!g401) & (!g414)) + ((!g301) & (g251) & (!g302) & (!sk[127]) & (!g401) & (g414)) + ((!g301) & (g251) & (!g302) & (!sk[127]) & (g401) & (!g414)) + ((!g301) & (g251) & (!g302) & (!sk[127]) & (g401) & (g414)) + ((!g301) & (g251) & (!g302) & (sk[127]) & (!g401) & (!g414)) + ((!g301) & (g251) & (!g302) & (sk[127]) & (!g401) & (g414)) + ((!g301) & (g251) & (g302) & (!sk[127]) & (!g401) & (!g414)) + ((!g301) & (g251) & (g302) & (!sk[127]) & (!g401) & (g414)) + ((!g301) & (g251) & (g302) & (!sk[127]) & (g401) & (!g414)) + ((!g301) & (g251) & (g302) & (!sk[127]) & (g401) & (g414)) + ((!g301) & (g251) & (g302) & (sk[127]) & (g401) & (!g414)) + ((!g301) & (g251) & (g302) & (sk[127]) & (g401) & (g414)) + ((g301) & (!g251) & (!g302) & (!sk[127]) & (g401) & (!g414)) + ((g301) & (!g251) & (!g302) & (!sk[127]) & (g401) & (g414)) + ((g301) & (!g251) & (!g302) & (sk[127]) & (!g401) & (!g414)) + ((g301) & (!g251) & (!g302) & (sk[127]) & (!g401) & (g414)) + ((g301) & (!g251) & (g302) & (!sk[127]) & (!g401) & (!g414)) + ((g301) & (!g251) & (g302) & (!sk[127]) & (!g401) & (g414)) + ((g301) & (!g251) & (g302) & (!sk[127]) & (g401) & (!g414)) + ((g301) & (!g251) & (g302) & (!sk[127]) & (g401) & (g414)) + ((g301) & (!g251) & (g302) & (sk[127]) & (g401) & (!g414)) + ((g301) & (!g251) & (g302) & (sk[127]) & (g401) & (g414)) + ((g301) & (g251) & (!g302) & (!sk[127]) & (!g401) & (!g414)) + ((g301) & (g251) & (!g302) & (!sk[127]) & (!g401) & (g414)) + ((g301) & (g251) & (!g302) & (!sk[127]) & (g401) & (!g414)) + ((g301) & (g251) & (!g302) & (!sk[127]) & (g401) & (g414)) + ((g301) & (g251) & (!g302) & (sk[127]) & (!g401) & (!g414)) + ((g301) & (g251) & (!g302) & (sk[127]) & (g401) & (!g414)) + ((g301) & (g251) & (g302) & (!sk[127]) & (!g401) & (!g414)) + ((g301) & (g251) & (g302) & (!sk[127]) & (!g401) & (g414)) + ((g301) & (g251) & (g302) & (!sk[127]) & (g401) & (!g414)) + ((g301) & (g251) & (g302) & (!sk[127]) & (g401) & (g414)));
	assign g502 = (((!g466) & (!sk[0]) & (g467) & (!g501)) + ((!g466) & (!sk[0]) & (g467) & (g501)) + ((!g466) & (sk[0]) & (!g467) & (!g501)) + ((!g466) & (sk[0]) & (g467) & (g501)) + ((g466) & (!sk[0]) & (g467) & (!g501)) + ((g466) & (!sk[0]) & (g467) & (g501)) + ((g466) & (sk[0]) & (!g467) & (g501)) + ((g466) & (sk[0]) & (g467) & (!g501)));
	assign g503 = (((!g491) & (!g482) & (!sk[1]) & (!g496) & (g500) & (!g502)) + ((!g491) & (!g482) & (!sk[1]) & (!g496) & (g500) & (g502)) + ((!g491) & (!g482) & (!sk[1]) & (g496) & (!g500) & (!g502)) + ((!g491) & (!g482) & (!sk[1]) & (g496) & (!g500) & (g502)) + ((!g491) & (!g482) & (!sk[1]) & (g496) & (g500) & (!g502)) + ((!g491) & (!g482) & (!sk[1]) & (g496) & (g500) & (g502)) + ((!g491) & (!g482) & (sk[1]) & (g496) & (!g500) & (!g502)) + ((!g491) & (!g482) & (sk[1]) & (g496) & (g500) & (g502)) + ((!g491) & (g482) & (!sk[1]) & (!g496) & (!g500) & (!g502)) + ((!g491) & (g482) & (!sk[1]) & (!g496) & (!g500) & (g502)) + ((!g491) & (g482) & (!sk[1]) & (!g496) & (g500) & (!g502)) + ((!g491) & (g482) & (!sk[1]) & (!g496) & (g500) & (g502)) + ((!g491) & (g482) & (!sk[1]) & (g496) & (!g500) & (!g502)) + ((!g491) & (g482) & (!sk[1]) & (g496) & (!g500) & (g502)) + ((!g491) & (g482) & (!sk[1]) & (g496) & (g500) & (!g502)) + ((!g491) & (g482) & (!sk[1]) & (g496) & (g500) & (g502)) + ((!g491) & (g482) & (sk[1]) & (!g496) & (!g500) & (!g502)) + ((!g491) & (g482) & (sk[1]) & (!g496) & (g500) & (g502)) + ((!g491) & (g482) & (sk[1]) & (g496) & (!g500) & (!g502)) + ((!g491) & (g482) & (sk[1]) & (g496) & (!g500) & (g502)) + ((!g491) & (g482) & (sk[1]) & (g496) & (g500) & (!g502)) + ((!g491) & (g482) & (sk[1]) & (g496) & (g500) & (g502)) + ((g491) & (!g482) & (!sk[1]) & (!g496) & (g500) & (!g502)) + ((g491) & (!g482) & (!sk[1]) & (!g496) & (g500) & (g502)) + ((g491) & (!g482) & (!sk[1]) & (g496) & (!g500) & (!g502)) + ((g491) & (!g482) & (!sk[1]) & (g496) & (!g500) & (g502)) + ((g491) & (!g482) & (!sk[1]) & (g496) & (g500) & (!g502)) + ((g491) & (!g482) & (!sk[1]) & (g496) & (g500) & (g502)) + ((g491) & (!g482) & (sk[1]) & (!g496) & (!g500) & (!g502)) + ((g491) & (!g482) & (sk[1]) & (!g496) & (g500) & (g502)) + ((g491) & (!g482) & (sk[1]) & (g496) & (!g500) & (!g502)) + ((g491) & (!g482) & (sk[1]) & (g496) & (!g500) & (g502)) + ((g491) & (!g482) & (sk[1]) & (g496) & (g500) & (!g502)) + ((g491) & (!g482) & (sk[1]) & (g496) & (g500) & (g502)) + ((g491) & (g482) & (!sk[1]) & (!g496) & (!g500) & (!g502)) + ((g491) & (g482) & (!sk[1]) & (!g496) & (!g500) & (g502)) + ((g491) & (g482) & (!sk[1]) & (!g496) & (g500) & (!g502)) + ((g491) & (g482) & (!sk[1]) & (!g496) & (g500) & (g502)) + ((g491) & (g482) & (!sk[1]) & (g496) & (!g500) & (!g502)) + ((g491) & (g482) & (!sk[1]) & (g496) & (!g500) & (g502)) + ((g491) & (g482) & (!sk[1]) & (g496) & (g500) & (!g502)) + ((g491) & (g482) & (!sk[1]) & (g496) & (g500) & (g502)) + ((g491) & (g482) & (sk[1]) & (g496) & (!g500) & (!g502)) + ((g491) & (g482) & (sk[1]) & (g496) & (g500) & (g502)));
	assign g504 = (((!g305) & (!g200) & (!sk[2]) & (!g347) & (g425)) + ((!g305) & (!g200) & (!sk[2]) & (g347) & (g425)) + ((!g305) & (!g200) & (sk[2]) & (!g347) & (!g425)) + ((!g305) & (!g200) & (sk[2]) & (!g347) & (g425)) + ((!g305) & (g200) & (!sk[2]) & (!g347) & (g425)) + ((!g305) & (g200) & (!sk[2]) & (g347) & (g425)) + ((!g305) & (g200) & (sk[2]) & (!g347) & (!g425)) + ((g305) & (!g200) & (!sk[2]) & (!g347) & (!g425)) + ((g305) & (!g200) & (!sk[2]) & (!g347) & (g425)) + ((g305) & (!g200) & (!sk[2]) & (g347) & (!g425)) + ((g305) & (!g200) & (!sk[2]) & (g347) & (g425)) + ((g305) & (!g200) & (sk[2]) & (!g347) & (g425)) + ((g305) & (!g200) & (sk[2]) & (g347) & (!g425)) + ((g305) & (g200) & (!sk[2]) & (!g347) & (!g425)) + ((g305) & (g200) & (!sk[2]) & (!g347) & (g425)) + ((g305) & (g200) & (!sk[2]) & (g347) & (!g425)) + ((g305) & (g200) & (!sk[2]) & (g347) & (g425)) + ((g305) & (g200) & (sk[2]) & (g347) & (!g425)));
	assign g505 = (((!g196) & (!g198) & (!g347) & (g365) & (!g367) & (!g393)) + ((!g196) & (!g198) & (!g347) & (g365) & (!g367) & (g393)) + ((!g196) & (!g198) & (!g347) & (g365) & (g367) & (!g393)) + ((!g196) & (!g198) & (!g347) & (g365) & (g367) & (g393)) + ((!g196) & (!g198) & (g347) & (!g365) & (!g367) & (!g393)) + ((!g196) & (!g198) & (g347) & (!g365) & (!g367) & (g393)) + ((!g196) & (!g198) & (g347) & (!g365) & (g367) & (!g393)) + ((!g196) & (!g198) & (g347) & (!g365) & (g367) & (g393)) + ((!g196) & (!g198) & (g347) & (g365) & (!g367) & (!g393)) + ((!g196) & (!g198) & (g347) & (g365) & (!g367) & (g393)) + ((!g196) & (g198) & (g347) & (g365) & (!g367) & (!g393)) + ((!g196) & (g198) & (g347) & (g365) & (!g367) & (g393)) + ((g196) & (!g198) & (!g347) & (!g365) & (g367) & (!g393)) + ((g196) & (!g198) & (g347) & (g365) & (g367) & (!g393)) + ((g196) & (g198) & (!g347) & (!g365) & (g367) & (!g393)) + ((g196) & (g198) & (!g347) & (g365) & (!g367) & (!g393)) + ((g196) & (g198) & (!g347) & (g365) & (g367) & (!g393)) + ((g196) & (g198) & (g347) & (!g365) & (!g367) & (!g393)) + ((g196) & (g198) & (g347) & (!g365) & (g367) & (!g393)) + ((g196) & (g198) & (g347) & (g365) & (g367) & (!g393)));
	assign g506 = (((!g2) & (!g122) & (!g159) & (g196) & (!sk[4]) & (!g401)) + ((!g2) & (!g122) & (!g159) & (g196) & (!sk[4]) & (g401)) + ((!g2) & (!g122) & (!g159) & (g196) & (sk[4]) & (!g401)) + ((!g2) & (!g122) & (!g159) & (g196) & (sk[4]) & (g401)) + ((!g2) & (!g122) & (g159) & (!g196) & (!sk[4]) & (!g401)) + ((!g2) & (!g122) & (g159) & (!g196) & (!sk[4]) & (g401)) + ((!g2) & (!g122) & (g159) & (!g196) & (sk[4]) & (!g401)) + ((!g2) & (!g122) & (g159) & (!g196) & (sk[4]) & (g401)) + ((!g2) & (!g122) & (g159) & (g196) & (!sk[4]) & (!g401)) + ((!g2) & (!g122) & (g159) & (g196) & (!sk[4]) & (g401)) + ((!g2) & (!g122) & (g159) & (g196) & (sk[4]) & (!g401)) + ((!g2) & (g122) & (!g159) & (!g196) & (!sk[4]) & (!g401)) + ((!g2) & (g122) & (!g159) & (!g196) & (!sk[4]) & (g401)) + ((!g2) & (g122) & (!g159) & (!g196) & (sk[4]) & (g401)) + ((!g2) & (g122) & (!g159) & (g196) & (!sk[4]) & (!g401)) + ((!g2) & (g122) & (!g159) & (g196) & (!sk[4]) & (g401)) + ((!g2) & (g122) & (g159) & (!g196) & (!sk[4]) & (!g401)) + ((!g2) & (g122) & (g159) & (!g196) & (!sk[4]) & (g401)) + ((!g2) & (g122) & (g159) & (g196) & (!sk[4]) & (!g401)) + ((!g2) & (g122) & (g159) & (g196) & (!sk[4]) & (g401)) + ((g2) & (!g122) & (!g159) & (g196) & (!sk[4]) & (!g401)) + ((g2) & (!g122) & (!g159) & (g196) & (!sk[4]) & (g401)) + ((g2) & (!g122) & (g159) & (!g196) & (!sk[4]) & (!g401)) + ((g2) & (!g122) & (g159) & (!g196) & (!sk[4]) & (g401)) + ((g2) & (!g122) & (g159) & (g196) & (!sk[4]) & (!g401)) + ((g2) & (!g122) & (g159) & (g196) & (!sk[4]) & (g401)) + ((g2) & (!g122) & (g159) & (g196) & (sk[4]) & (!g401)) + ((g2) & (g122) & (!g159) & (!g196) & (!sk[4]) & (!g401)) + ((g2) & (g122) & (!g159) & (!g196) & (!sk[4]) & (g401)) + ((g2) & (g122) & (!g159) & (!g196) & (sk[4]) & (g401)) + ((g2) & (g122) & (!g159) & (g196) & (!sk[4]) & (!g401)) + ((g2) & (g122) & (!g159) & (g196) & (!sk[4]) & (g401)) + ((g2) & (g122) & (!g159) & (g196) & (sk[4]) & (!g401)) + ((g2) & (g122) & (!g159) & (g196) & (sk[4]) & (g401)) + ((g2) & (g122) & (g159) & (!g196) & (!sk[4]) & (!g401)) + ((g2) & (g122) & (g159) & (!g196) & (!sk[4]) & (g401)) + ((g2) & (g122) & (g159) & (!g196) & (sk[4]) & (!g401)) + ((g2) & (g122) & (g159) & (!g196) & (sk[4]) & (g401)) + ((g2) & (g122) & (g159) & (g196) & (!sk[4]) & (!g401)) + ((g2) & (g122) & (g159) & (g196) & (!sk[4]) & (g401)));
	assign g507 = (((!g493) & (sk[5]) & (!g494)) + ((g493) & (!sk[5]) & (g494)) + ((g493) & (sk[5]) & (g494)));
	assign g508 = (((!g2) & (!g122) & (!g159) & (g196) & (!sk[6]) & (!g367)) + ((!g2) & (!g122) & (!g159) & (g196) & (!sk[6]) & (g367)) + ((!g2) & (!g122) & (!g159) & (g196) & (sk[6]) & (!g367)) + ((!g2) & (!g122) & (g159) & (!g196) & (!sk[6]) & (!g367)) + ((!g2) & (!g122) & (g159) & (!g196) & (!sk[6]) & (g367)) + ((!g2) & (!g122) & (g159) & (!g196) & (sk[6]) & (!g367)) + ((!g2) & (!g122) & (g159) & (g196) & (!sk[6]) & (!g367)) + ((!g2) & (!g122) & (g159) & (g196) & (!sk[6]) & (g367)) + ((!g2) & (!g122) & (g159) & (g196) & (sk[6]) & (!g367)) + ((!g2) & (!g122) & (g159) & (g196) & (sk[6]) & (g367)) + ((!g2) & (g122) & (!g159) & (!g196) & (!sk[6]) & (!g367)) + ((!g2) & (g122) & (!g159) & (!g196) & (!sk[6]) & (g367)) + ((!g2) & (g122) & (!g159) & (g196) & (!sk[6]) & (!g367)) + ((!g2) & (g122) & (!g159) & (g196) & (!sk[6]) & (g367)) + ((!g2) & (g122) & (!g159) & (g196) & (sk[6]) & (g367)) + ((!g2) & (g122) & (g159) & (!g196) & (!sk[6]) & (!g367)) + ((!g2) & (g122) & (g159) & (!g196) & (!sk[6]) & (g367)) + ((!g2) & (g122) & (g159) & (!g196) & (sk[6]) & (g367)) + ((!g2) & (g122) & (g159) & (g196) & (!sk[6]) & (!g367)) + ((!g2) & (g122) & (g159) & (g196) & (!sk[6]) & (g367)) + ((g2) & (!g122) & (!g159) & (g196) & (!sk[6]) & (!g367)) + ((g2) & (!g122) & (!g159) & (g196) & (!sk[6]) & (g367)) + ((g2) & (!g122) & (!g159) & (g196) & (sk[6]) & (!g367)) + ((g2) & (!g122) & (g159) & (!g196) & (!sk[6]) & (!g367)) + ((g2) & (!g122) & (g159) & (!g196) & (!sk[6]) & (g367)) + ((g2) & (!g122) & (g159) & (!g196) & (sk[6]) & (!g367)) + ((g2) & (!g122) & (g159) & (g196) & (!sk[6]) & (!g367)) + ((g2) & (!g122) & (g159) & (g196) & (!sk[6]) & (g367)) + ((g2) & (g122) & (!g159) & (!g196) & (!sk[6]) & (!g367)) + ((g2) & (g122) & (!g159) & (!g196) & (!sk[6]) & (g367)) + ((g2) & (g122) & (!g159) & (!g196) & (sk[6]) & (!g367)) + ((g2) & (g122) & (!g159) & (!g196) & (sk[6]) & (g367)) + ((g2) & (g122) & (!g159) & (g196) & (!sk[6]) & (!g367)) + ((g2) & (g122) & (!g159) & (g196) & (!sk[6]) & (g367)) + ((g2) & (g122) & (!g159) & (g196) & (sk[6]) & (g367)) + ((g2) & (g122) & (g159) & (!g196) & (!sk[6]) & (!g367)) + ((g2) & (g122) & (g159) & (!g196) & (!sk[6]) & (g367)) + ((g2) & (g122) & (g159) & (!g196) & (sk[6]) & (g367)) + ((g2) & (g122) & (g159) & (g196) & (!sk[6]) & (!g367)) + ((g2) & (g122) & (g159) & (g196) & (!sk[6]) & (g367)));
	assign g509 = (((!g196) & (!g198) & (!g200) & (!g347) & (g365) & (!g393)) + ((!g196) & (!g198) & (!g200) & (!g347) & (g365) & (g393)) + ((!g196) & (!g198) & (!g200) & (g347) & (!g365) & (!g393)) + ((!g196) & (!g198) & (!g200) & (g347) & (!g365) & (g393)) + ((!g196) & (!g198) & (!g200) & (g347) & (g365) & (!g393)) + ((!g196) & (!g198) & (!g200) & (g347) & (g365) & (g393)) + ((!g196) & (!g198) & (g200) & (g347) & (g365) & (!g393)) + ((!g196) & (!g198) & (g200) & (g347) & (g365) & (g393)) + ((!g196) & (g198) & (!g200) & (!g347) & (g365) & (!g393)) + ((!g196) & (g198) & (!g200) & (!g347) & (g365) & (g393)) + ((!g196) & (g198) & (!g200) & (g347) & (!g365) & (!g393)) + ((!g196) & (g198) & (!g200) & (g347) & (!g365) & (g393)) + ((g196) & (!g198) & (g200) & (!g347) & (g365) & (!g393)) + ((g196) & (!g198) & (g200) & (g347) & (!g365) & (!g393)) + ((g196) & (g198) & (!g200) & (!g347) & (!g365) & (!g393)) + ((g196) & (g198) & (!g200) & (g347) & (g365) & (!g393)) + ((g196) & (g198) & (g200) & (!g347) & (!g365) & (!g393)) + ((g196) & (g198) & (g200) & (!g347) & (g365) & (!g393)) + ((g196) & (g198) & (g200) & (g347) & (!g365) & (!g393)) + ((g196) & (g198) & (g200) & (g347) & (g365) & (!g393)));
	assign g510 = (((!sk[8]) & (g508) & (g509)) + ((sk[8]) & (!g508) & (!g509)) + ((sk[8]) & (g508) & (g509)));
	assign g511 = (((!sk[9]) & (!g251) & (!g122) & (!g280) & (g401) & (!g414)) + ((!sk[9]) & (!g251) & (!g122) & (!g280) & (g401) & (g414)) + ((!sk[9]) & (!g251) & (!g122) & (g280) & (!g401) & (!g414)) + ((!sk[9]) & (!g251) & (!g122) & (g280) & (!g401) & (g414)) + ((!sk[9]) & (!g251) & (!g122) & (g280) & (g401) & (!g414)) + ((!sk[9]) & (!g251) & (!g122) & (g280) & (g401) & (g414)) + ((!sk[9]) & (!g251) & (g122) & (!g280) & (!g401) & (!g414)) + ((!sk[9]) & (!g251) & (g122) & (!g280) & (!g401) & (g414)) + ((!sk[9]) & (!g251) & (g122) & (!g280) & (g401) & (!g414)) + ((!sk[9]) & (!g251) & (g122) & (!g280) & (g401) & (g414)) + ((!sk[9]) & (!g251) & (g122) & (g280) & (!g401) & (!g414)) + ((!sk[9]) & (!g251) & (g122) & (g280) & (!g401) & (g414)) + ((!sk[9]) & (!g251) & (g122) & (g280) & (g401) & (!g414)) + ((!sk[9]) & (!g251) & (g122) & (g280) & (g401) & (g414)) + ((!sk[9]) & (g251) & (!g122) & (!g280) & (g401) & (!g414)) + ((!sk[9]) & (g251) & (!g122) & (!g280) & (g401) & (g414)) + ((!sk[9]) & (g251) & (!g122) & (g280) & (!g401) & (!g414)) + ((!sk[9]) & (g251) & (!g122) & (g280) & (!g401) & (g414)) + ((!sk[9]) & (g251) & (!g122) & (g280) & (g401) & (!g414)) + ((!sk[9]) & (g251) & (!g122) & (g280) & (g401) & (g414)) + ((!sk[9]) & (g251) & (g122) & (!g280) & (!g401) & (!g414)) + ((!sk[9]) & (g251) & (g122) & (!g280) & (!g401) & (g414)) + ((!sk[9]) & (g251) & (g122) & (!g280) & (g401) & (!g414)) + ((!sk[9]) & (g251) & (g122) & (!g280) & (g401) & (g414)) + ((!sk[9]) & (g251) & (g122) & (g280) & (!g401) & (!g414)) + ((!sk[9]) & (g251) & (g122) & (g280) & (!g401) & (g414)) + ((!sk[9]) & (g251) & (g122) & (g280) & (g401) & (!g414)) + ((!sk[9]) & (g251) & (g122) & (g280) & (g401) & (g414)) + ((sk[9]) & (!g251) & (!g122) & (g280) & (!g401) & (!g414)) + ((sk[9]) & (!g251) & (!g122) & (g280) & (!g401) & (g414)) + ((sk[9]) & (!g251) & (g122) & (!g280) & (!g401) & (!g414)) + ((sk[9]) & (!g251) & (g122) & (!g280) & (!g401) & (g414)) + ((sk[9]) & (!g251) & (g122) & (g280) & (!g401) & (!g414)) + ((sk[9]) & (!g251) & (g122) & (g280) & (g401) & (!g414)) + ((sk[9]) & (g251) & (!g122) & (!g280) & (!g401) & (g414)) + ((sk[9]) & (g251) & (!g122) & (!g280) & (g401) & (g414)) + ((sk[9]) & (g251) & (!g122) & (g280) & (g401) & (!g414)) + ((sk[9]) & (g251) & (!g122) & (g280) & (g401) & (g414)) + ((sk[9]) & (g251) & (g122) & (!g280) & (g401) & (!g414)) + ((sk[9]) & (g251) & (g122) & (!g280) & (g401) & (g414)));
	assign g512 = (((!g504) & (!g505) & (!g506) & (!g507) & (!g510) & (!g511)) + ((!g504) & (!g505) & (!g506) & (!g507) & (g510) & (g511)) + ((!g504) & (!g505) & (g506) & (!g507) & (!g510) & (!g511)) + ((!g504) & (!g505) & (g506) & (!g507) & (g510) & (g511)) + ((!g504) & (g505) & (!g506) & (!g507) & (!g510) & (!g511)) + ((!g504) & (g505) & (!g506) & (!g507) & (g510) & (g511)) + ((!g504) & (g505) & (g506) & (!g507) & (!g510) & (!g511)) + ((!g504) & (g505) & (g506) & (!g507) & (!g510) & (g511)) + ((!g504) & (g505) & (g506) & (!g507) & (g510) & (!g511)) + ((!g504) & (g505) & (g506) & (!g507) & (g510) & (g511)) + ((!g504) & (g505) & (g506) & (g507) & (!g510) & (!g511)) + ((!g504) & (g505) & (g506) & (g507) & (g510) & (g511)) + ((g504) & (!g505) & (!g506) & (!g507) & (!g510) & (!g511)) + ((g504) & (!g505) & (!g506) & (!g507) & (g510) & (g511)) + ((g504) & (!g505) & (g506) & (!g507) & (!g510) & (!g511)) + ((g504) & (!g505) & (g506) & (!g507) & (!g510) & (g511)) + ((g504) & (!g505) & (g506) & (!g507) & (g510) & (!g511)) + ((g504) & (!g505) & (g506) & (!g507) & (g510) & (g511)) + ((g504) & (!g505) & (g506) & (g507) & (!g510) & (!g511)) + ((g504) & (!g505) & (g506) & (g507) & (g510) & (g511)) + ((g504) & (g505) & (!g506) & (!g507) & (!g510) & (!g511)) + ((g504) & (g505) & (!g506) & (!g507) & (!g510) & (g511)) + ((g504) & (g505) & (!g506) & (!g507) & (g510) & (!g511)) + ((g504) & (g505) & (!g506) & (!g507) & (g510) & (g511)) + ((g504) & (g505) & (!g506) & (g507) & (!g510) & (!g511)) + ((g504) & (g505) & (!g506) & (g507) & (g510) & (g511)) + ((g504) & (g505) & (g506) & (!g507) & (!g510) & (!g511)) + ((g504) & (g505) & (g506) & (!g507) & (!g510) & (g511)) + ((g504) & (g505) & (g506) & (!g507) & (g510) & (!g511)) + ((g504) & (g505) & (g506) & (!g507) & (g510) & (g511)) + ((g504) & (g505) & (g506) & (g507) & (!g510) & (!g511)) + ((g504) & (g505) & (g506) & (g507) & (g510) & (g511)));
	assign g513 = (((!g122) & (!sk[11]) & (!g159) & (!g196) & (g401) & (!g414)) + ((!g122) & (!sk[11]) & (!g159) & (!g196) & (g401) & (g414)) + ((!g122) & (!sk[11]) & (!g159) & (g196) & (!g401) & (!g414)) + ((!g122) & (!sk[11]) & (!g159) & (g196) & (!g401) & (g414)) + ((!g122) & (!sk[11]) & (!g159) & (g196) & (g401) & (!g414)) + ((!g122) & (!sk[11]) & (!g159) & (g196) & (g401) & (g414)) + ((!g122) & (!sk[11]) & (g159) & (!g196) & (!g401) & (!g414)) + ((!g122) & (!sk[11]) & (g159) & (!g196) & (!g401) & (g414)) + ((!g122) & (!sk[11]) & (g159) & (!g196) & (g401) & (!g414)) + ((!g122) & (!sk[11]) & (g159) & (!g196) & (g401) & (g414)) + ((!g122) & (!sk[11]) & (g159) & (g196) & (!g401) & (!g414)) + ((!g122) & (!sk[11]) & (g159) & (g196) & (!g401) & (g414)) + ((!g122) & (!sk[11]) & (g159) & (g196) & (g401) & (!g414)) + ((!g122) & (!sk[11]) & (g159) & (g196) & (g401) & (g414)) + ((!g122) & (sk[11]) & (!g159) & (g196) & (!g401) & (!g414)) + ((!g122) & (sk[11]) & (!g159) & (g196) & (!g401) & (g414)) + ((!g122) & (sk[11]) & (g159) & (!g196) & (!g401) & (!g414)) + ((!g122) & (sk[11]) & (g159) & (!g196) & (!g401) & (g414)) + ((!g122) & (sk[11]) & (g159) & (g196) & (!g401) & (!g414)) + ((!g122) & (sk[11]) & (g159) & (g196) & (g401) & (!g414)) + ((g122) & (!sk[11]) & (!g159) & (!g196) & (g401) & (!g414)) + ((g122) & (!sk[11]) & (!g159) & (!g196) & (g401) & (g414)) + ((g122) & (!sk[11]) & (!g159) & (g196) & (!g401) & (!g414)) + ((g122) & (!sk[11]) & (!g159) & (g196) & (!g401) & (g414)) + ((g122) & (!sk[11]) & (!g159) & (g196) & (g401) & (!g414)) + ((g122) & (!sk[11]) & (!g159) & (g196) & (g401) & (g414)) + ((g122) & (!sk[11]) & (g159) & (!g196) & (!g401) & (!g414)) + ((g122) & (!sk[11]) & (g159) & (!g196) & (!g401) & (g414)) + ((g122) & (!sk[11]) & (g159) & (!g196) & (g401) & (!g414)) + ((g122) & (!sk[11]) & (g159) & (!g196) & (g401) & (g414)) + ((g122) & (!sk[11]) & (g159) & (g196) & (!g401) & (!g414)) + ((g122) & (!sk[11]) & (g159) & (g196) & (!g401) & (g414)) + ((g122) & (!sk[11]) & (g159) & (g196) & (g401) & (!g414)) + ((g122) & (!sk[11]) & (g159) & (g196) & (g401) & (g414)) + ((g122) & (sk[11]) & (!g159) & (!g196) & (!g401) & (g414)) + ((g122) & (sk[11]) & (!g159) & (!g196) & (g401) & (g414)) + ((g122) & (sk[11]) & (!g159) & (g196) & (g401) & (!g414)) + ((g122) & (sk[11]) & (!g159) & (g196) & (g401) & (g414)) + ((g122) & (sk[11]) & (g159) & (!g196) & (g401) & (!g414)) + ((g122) & (sk[11]) & (g159) & (!g196) & (g401) & (g414)));
	assign g514 = (((!g2) & (!g196) & (!g347) & (g365) & (!g367) & (!g393)) + ((!g2) & (!g196) & (!g347) & (g365) & (!g367) & (g393)) + ((!g2) & (!g196) & (g347) & (!g365) & (!g367) & (!g393)) + ((!g2) & (!g196) & (g347) & (!g365) & (!g367) & (g393)) + ((!g2) & (!g196) & (g347) & (g365) & (!g367) & (!g393)) + ((!g2) & (!g196) & (g347) & (g365) & (!g367) & (g393)) + ((!g2) & (!g196) & (g347) & (g365) & (g367) & (!g393)) + ((!g2) & (!g196) & (g347) & (g365) & (g367) & (g393)) + ((!g2) & (g196) & (!g347) & (g365) & (g367) & (!g393)) + ((!g2) & (g196) & (g347) & (!g365) & (g367) & (!g393)) + ((g2) & (!g196) & (!g347) & (g365) & (!g367) & (!g393)) + ((g2) & (!g196) & (!g347) & (g365) & (!g367) & (g393)) + ((g2) & (!g196) & (g347) & (!g365) & (!g367) & (!g393)) + ((g2) & (!g196) & (g347) & (!g365) & (!g367) & (g393)) + ((g2) & (g196) & (!g347) & (!g365) & (!g367) & (!g393)) + ((g2) & (g196) & (!g347) & (!g365) & (g367) & (!g393)) + ((g2) & (g196) & (!g347) & (g365) & (g367) & (!g393)) + ((g2) & (g196) & (g347) & (!g365) & (g367) & (!g393)) + ((g2) & (g196) & (g347) & (g365) & (!g367) & (!g393)) + ((g2) & (g196) & (g347) & (g365) & (g367) & (!g393)));
	assign g515 = (((!sk[13]) & (!g198) & (!g200) & (!g347) & (g425)) + ((!sk[13]) & (!g198) & (!g200) & (g347) & (g425)) + ((!sk[13]) & (!g198) & (g200) & (!g347) & (g425)) + ((!sk[13]) & (!g198) & (g200) & (g347) & (g425)) + ((!sk[13]) & (g198) & (!g200) & (!g347) & (!g425)) + ((!sk[13]) & (g198) & (!g200) & (!g347) & (g425)) + ((!sk[13]) & (g198) & (!g200) & (g347) & (!g425)) + ((!sk[13]) & (g198) & (!g200) & (g347) & (g425)) + ((!sk[13]) & (g198) & (g200) & (!g347) & (!g425)) + ((!sk[13]) & (g198) & (g200) & (!g347) & (g425)) + ((!sk[13]) & (g198) & (g200) & (g347) & (!g425)) + ((!sk[13]) & (g198) & (g200) & (g347) & (g425)) + ((sk[13]) & (!g198) & (!g200) & (!g347) & (!g425)) + ((sk[13]) & (!g198) & (!g200) & (!g347) & (g425)) + ((sk[13]) & (!g198) & (g200) & (!g347) & (g425)) + ((sk[13]) & (!g198) & (g200) & (g347) & (!g425)) + ((sk[13]) & (g198) & (!g200) & (!g347) & (!g425)) + ((sk[13]) & (g198) & (g200) & (g347) & (!g425)));
	assign g516 = (((!sk[14]) & (!g159) & (g196) & (!g414)) + ((!sk[14]) & (!g159) & (g196) & (g414)) + ((!sk[14]) & (g159) & (g196) & (!g414)) + ((!sk[14]) & (g159) & (g196) & (g414)) + ((sk[14]) & (!g159) & (g196) & (g414)) + ((sk[14]) & (g159) & (!g196) & (g414)));
	assign g517 = (((!g197) & (!g513) & (!sk[15]) & (!g514) & (g515) & (!g516)) + ((!g197) & (!g513) & (!sk[15]) & (!g514) & (g515) & (g516)) + ((!g197) & (!g513) & (!sk[15]) & (g514) & (!g515) & (!g516)) + ((!g197) & (!g513) & (!sk[15]) & (g514) & (!g515) & (g516)) + ((!g197) & (!g513) & (!sk[15]) & (g514) & (g515) & (!g516)) + ((!g197) & (!g513) & (!sk[15]) & (g514) & (g515) & (g516)) + ((!g197) & (!g513) & (sk[15]) & (g514) & (g515) & (!g516)) + ((!g197) & (!g513) & (sk[15]) & (g514) & (g515) & (g516)) + ((!g197) & (g513) & (!sk[15]) & (!g514) & (!g515) & (!g516)) + ((!g197) & (g513) & (!sk[15]) & (!g514) & (!g515) & (g516)) + ((!g197) & (g513) & (!sk[15]) & (!g514) & (g515) & (!g516)) + ((!g197) & (g513) & (!sk[15]) & (!g514) & (g515) & (g516)) + ((!g197) & (g513) & (!sk[15]) & (g514) & (!g515) & (!g516)) + ((!g197) & (g513) & (!sk[15]) & (g514) & (!g515) & (g516)) + ((!g197) & (g513) & (!sk[15]) & (g514) & (g515) & (!g516)) + ((!g197) & (g513) & (!sk[15]) & (g514) & (g515) & (g516)) + ((!g197) & (g513) & (sk[15]) & (!g514) & (g515) & (!g516)) + ((!g197) & (g513) & (sk[15]) & (!g514) & (g515) & (g516)) + ((!g197) & (g513) & (sk[15]) & (g514) & (!g515) & (!g516)) + ((!g197) & (g513) & (sk[15]) & (g514) & (!g515) & (g516)) + ((!g197) & (g513) & (sk[15]) & (g514) & (g515) & (!g516)) + ((!g197) & (g513) & (sk[15]) & (g514) & (g515) & (g516)) + ((g197) & (!g513) & (!sk[15]) & (!g514) & (g515) & (!g516)) + ((g197) & (!g513) & (!sk[15]) & (!g514) & (g515) & (g516)) + ((g197) & (!g513) & (!sk[15]) & (g514) & (!g515) & (!g516)) + ((g197) & (!g513) & (!sk[15]) & (g514) & (!g515) & (g516)) + ((g197) & (!g513) & (!sk[15]) & (g514) & (g515) & (!g516)) + ((g197) & (!g513) & (!sk[15]) & (g514) & (g515) & (g516)) + ((g197) & (!g513) & (sk[15]) & (g514) & (!g515) & (!g516)) + ((g197) & (!g513) & (sk[15]) & (g514) & (g515) & (g516)) + ((g197) & (g513) & (!sk[15]) & (!g514) & (!g515) & (!g516)) + ((g197) & (g513) & (!sk[15]) & (!g514) & (!g515) & (g516)) + ((g197) & (g513) & (!sk[15]) & (!g514) & (g515) & (!g516)) + ((g197) & (g513) & (!sk[15]) & (!g514) & (g515) & (g516)) + ((g197) & (g513) & (!sk[15]) & (g514) & (!g515) & (!g516)) + ((g197) & (g513) & (!sk[15]) & (g514) & (!g515) & (g516)) + ((g197) & (g513) & (!sk[15]) & (g514) & (g515) & (!g516)) + ((g197) & (g513) & (!sk[15]) & (g514) & (g515) & (g516)) + ((g197) & (g513) & (sk[15]) & (!g514) & (!g515) & (!g516)) + ((g197) & (g513) & (sk[15]) & (!g514) & (g515) & (g516)) + ((g197) & (g513) & (sk[15]) & (g514) & (!g515) & (!g516)) + ((g197) & (g513) & (sk[15]) & (g514) & (!g515) & (g516)) + ((g197) & (g513) & (sk[15]) & (g514) & (g515) & (!g516)) + ((g197) & (g513) & (sk[15]) & (g514) & (g515) & (g516)));
	assign g518 = (((!sk[16]) & (!g122) & (g280) & (!g414)) + ((!sk[16]) & (!g122) & (g280) & (g414)) + ((!sk[16]) & (g122) & (g280) & (!g414)) + ((!sk[16]) & (g122) & (g280) & (g414)) + ((sk[16]) & (!g122) & (g280) & (g414)) + ((sk[16]) & (g122) & (!g280) & (g414)));
	assign g519 = (((!sk[17]) & (!g197) & (g515) & (!g516)) + ((!sk[17]) & (!g197) & (g515) & (g516)) + ((!sk[17]) & (g197) & (g515) & (!g516)) + ((!sk[17]) & (g197) & (g515) & (g516)) + ((sk[17]) & (g197) & (g515) & (!g516)));
	assign g520 = (((!sk[18]) & (!g196) & (g347) & (!g365)) + ((!sk[18]) & (!g196) & (g347) & (g365)) + ((!sk[18]) & (g196) & (g347) & (!g365)) + ((!sk[18]) & (g196) & (g347) & (g365)) + ((sk[18]) & (!g196) & (!g347) & (g365)) + ((sk[18]) & (!g196) & (g347) & (!g365)) + ((sk[18]) & (!g196) & (g347) & (g365)));
	assign g521 = (((!g196) & (!g347) & (!g365) & (g393) & (!sk[19]) & (!g414)) + ((!g196) & (!g347) & (!g365) & (g393) & (!sk[19]) & (g414)) + ((!g196) & (!g347) & (g365) & (!g393) & (!sk[19]) & (!g414)) + ((!g196) & (!g347) & (g365) & (!g393) & (!sk[19]) & (g414)) + ((!g196) & (!g347) & (g365) & (!g393) & (sk[19]) & (!g414)) + ((!g196) & (!g347) & (g365) & (g393) & (!sk[19]) & (!g414)) + ((!g196) & (!g347) & (g365) & (g393) & (!sk[19]) & (g414)) + ((!g196) & (!g347) & (g365) & (g393) & (sk[19]) & (!g414)) + ((!g196) & (g347) & (!g365) & (!g393) & (!sk[19]) & (!g414)) + ((!g196) & (g347) & (!g365) & (!g393) & (!sk[19]) & (g414)) + ((!g196) & (g347) & (!g365) & (!g393) & (sk[19]) & (!g414)) + ((!g196) & (g347) & (!g365) & (g393) & (!sk[19]) & (!g414)) + ((!g196) & (g347) & (!g365) & (g393) & (!sk[19]) & (g414)) + ((!g196) & (g347) & (!g365) & (g393) & (sk[19]) & (!g414)) + ((!g196) & (g347) & (g365) & (!g393) & (!sk[19]) & (!g414)) + ((!g196) & (g347) & (g365) & (!g393) & (!sk[19]) & (g414)) + ((!g196) & (g347) & (g365) & (!g393) & (sk[19]) & (!g414)) + ((!g196) & (g347) & (g365) & (!g393) & (sk[19]) & (g414)) + ((!g196) & (g347) & (g365) & (g393) & (!sk[19]) & (!g414)) + ((!g196) & (g347) & (g365) & (g393) & (!sk[19]) & (g414)) + ((!g196) & (g347) & (g365) & (g393) & (sk[19]) & (!g414)) + ((!g196) & (g347) & (g365) & (g393) & (sk[19]) & (g414)) + ((g196) & (!g347) & (!g365) & (g393) & (!sk[19]) & (!g414)) + ((g196) & (!g347) & (!g365) & (g393) & (!sk[19]) & (g414)) + ((g196) & (!g347) & (g365) & (!g393) & (!sk[19]) & (!g414)) + ((g196) & (!g347) & (g365) & (!g393) & (!sk[19]) & (g414)) + ((g196) & (!g347) & (g365) & (!g393) & (sk[19]) & (g414)) + ((g196) & (!g347) & (g365) & (g393) & (!sk[19]) & (!g414)) + ((g196) & (!g347) & (g365) & (g393) & (!sk[19]) & (g414)) + ((g196) & (g347) & (!g365) & (!g393) & (!sk[19]) & (!g414)) + ((g196) & (g347) & (!g365) & (!g393) & (!sk[19]) & (g414)) + ((g196) & (g347) & (!g365) & (!g393) & (sk[19]) & (g414)) + ((g196) & (g347) & (!g365) & (g393) & (!sk[19]) & (!g414)) + ((g196) & (g347) & (!g365) & (g393) & (!sk[19]) & (g414)) + ((g196) & (g347) & (g365) & (!g393) & (!sk[19]) & (!g414)) + ((g196) & (g347) & (g365) & (!g393) & (!sk[19]) & (g414)) + ((g196) & (g347) & (g365) & (g393) & (!sk[19]) & (!g414)) + ((g196) & (g347) & (g365) & (g393) & (!sk[19]) & (g414)));
	assign g522 = (((!g2) & (!sk[20]) & (!g347) & (!g367) & (g425)) + ((!g2) & (!sk[20]) & (!g347) & (g367) & (g425)) + ((!g2) & (!sk[20]) & (g347) & (!g367) & (g425)) + ((!g2) & (!sk[20]) & (g347) & (g367) & (g425)) + ((!g2) & (sk[20]) & (!g347) & (!g367) & (!g425)) + ((!g2) & (sk[20]) & (!g347) & (!g367) & (g425)) + ((!g2) & (sk[20]) & (!g347) & (g367) & (g425)) + ((!g2) & (sk[20]) & (g347) & (g367) & (!g425)) + ((g2) & (!sk[20]) & (!g347) & (!g367) & (!g425)) + ((g2) & (!sk[20]) & (!g347) & (!g367) & (g425)) + ((g2) & (!sk[20]) & (!g347) & (g367) & (!g425)) + ((g2) & (!sk[20]) & (!g347) & (g367) & (g425)) + ((g2) & (!sk[20]) & (g347) & (!g367) & (!g425)) + ((g2) & (!sk[20]) & (g347) & (!g367) & (g425)) + ((g2) & (!sk[20]) & (g347) & (g367) & (!g425)) + ((g2) & (!sk[20]) & (g347) & (g367) & (g425)) + ((g2) & (sk[20]) & (!g347) & (!g367) & (!g425)) + ((g2) & (sk[20]) & (g347) & (g367) & (!g425)));
	assign g523 = (((!g2) & (!sk[21]) & (!g347) & (!g401) & (g425)) + ((!g2) & (!sk[21]) & (!g347) & (g401) & (g425)) + ((!g2) & (!sk[21]) & (g347) & (!g401) & (g425)) + ((!g2) & (!sk[21]) & (g347) & (g401) & (g425)) + ((!g2) & (sk[21]) & (!g347) & (!g401) & (!g425)) + ((!g2) & (sk[21]) & (!g347) & (!g401) & (g425)) + ((!g2) & (sk[21]) & (!g347) & (g401) & (!g425)) + ((g2) & (!sk[21]) & (!g347) & (!g401) & (!g425)) + ((g2) & (!sk[21]) & (!g347) & (!g401) & (g425)) + ((g2) & (!sk[21]) & (!g347) & (g401) & (!g425)) + ((g2) & (!sk[21]) & (!g347) & (g401) & (g425)) + ((g2) & (!sk[21]) & (g347) & (!g401) & (!g425)) + ((g2) & (!sk[21]) & (g347) & (!g401) & (g425)) + ((g2) & (!sk[21]) & (g347) & (g401) & (!g425)) + ((g2) & (!sk[21]) & (g347) & (g401) & (g425)) + ((g2) & (sk[21]) & (!g347) & (!g401) & (g425)) + ((g2) & (sk[21]) & (g347) & (!g401) & (!g425)) + ((g2) & (sk[21]) & (g347) & (g401) & (!g425)));
	assign g524 = (((!g347) & (!g401) & (!g414) & (!sk[22]) & (g425)) + ((!g347) & (!g401) & (!g414) & (sk[22]) & (!g425)) + ((!g347) & (!g401) & (!g414) & (sk[22]) & (g425)) + ((!g347) & (!g401) & (g414) & (!sk[22]) & (g425)) + ((!g347) & (g401) & (!g414) & (!sk[22]) & (g425)) + ((!g347) & (g401) & (!g414) & (sk[22]) & (g425)) + ((!g347) & (g401) & (g414) & (!sk[22]) & (g425)) + ((g347) & (!g401) & (!g414) & (!sk[22]) & (!g425)) + ((g347) & (!g401) & (!g414) & (!sk[22]) & (g425)) + ((g347) & (!g401) & (g414) & (!sk[22]) & (!g425)) + ((g347) & (!g401) & (g414) & (!sk[22]) & (g425)) + ((g347) & (g401) & (!g414) & (!sk[22]) & (!g425)) + ((g347) & (g401) & (!g414) & (!sk[22]) & (g425)) + ((g347) & (g401) & (g414) & (!sk[22]) & (!g425)) + ((g347) & (g401) & (g414) & (!sk[22]) & (g425)));
	assign g525 = (((!g196) & (!g347) & (g365) & (!g393) & (!g401) & (!g414)) + ((!g196) & (!g347) & (g365) & (!g393) & (!g401) & (g414)) + ((!g196) & (!g347) & (g365) & (g393) & (!g401) & (!g414)) + ((!g196) & (!g347) & (g365) & (g393) & (!g401) & (g414)) + ((!g196) & (g347) & (!g365) & (!g393) & (!g401) & (!g414)) + ((!g196) & (g347) & (!g365) & (!g393) & (!g401) & (g414)) + ((!g196) & (g347) & (!g365) & (g393) & (!g401) & (!g414)) + ((!g196) & (g347) & (!g365) & (g393) & (!g401) & (g414)) + ((!g196) & (g347) & (g365) & (!g393) & (!g401) & (!g414)) + ((!g196) & (g347) & (g365) & (!g393) & (g401) & (!g414)) + ((!g196) & (g347) & (g365) & (g393) & (!g401) & (!g414)) + ((!g196) & (g347) & (g365) & (g393) & (g401) & (!g414)) + ((g196) & (!g347) & (!g365) & (!g393) & (!g401) & (g414)) + ((g196) & (!g347) & (!g365) & (!g393) & (g401) & (g414)) + ((g196) & (!g347) & (g365) & (!g393) & (g401) & (!g414)) + ((g196) & (!g347) & (g365) & (!g393) & (g401) & (g414)) + ((g196) & (g347) & (!g365) & (!g393) & (g401) & (!g414)) + ((g196) & (g347) & (!g365) & (!g393) & (g401) & (g414)) + ((g196) & (g347) & (g365) & (!g393) & (!g401) & (g414)) + ((g196) & (g347) & (g365) & (!g393) & (g401) & (g414)));
	assign g526 = (((!g520) & (!g521) & (!g522) & (!g523) & (!g524) & (!g525)) + ((!g520) & (!g521) & (!g522) & (!g523) & (!g524) & (g525)) + ((!g520) & (!g521) & (!g522) & (!g523) & (g524) & (!g525)) + ((!g520) & (!g521) & (!g522) & (!g523) & (g524) & (g525)) + ((!g520) & (!g521) & (!g522) & (g523) & (!g524) & (!g525)) + ((!g520) & (!g521) & (!g522) & (g523) & (!g524) & (g525)) + ((!g520) & (!g521) & (!g522) & (g523) & (g524) & (!g525)) + ((!g520) & (!g521) & (g522) & (!g523) & (!g524) & (!g525)) + ((!g520) & (!g521) & (g522) & (!g523) & (g524) & (!g525)) + ((!g520) & (!g521) & (g522) & (g523) & (!g524) & (!g525)) + ((!g520) & (g521) & (!g522) & (!g523) & (!g524) & (!g525)) + ((!g520) & (g521) & (!g522) & (!g523) & (!g524) & (g525)) + ((!g520) & (g521) & (!g522) & (!g523) & (g524) & (!g525)) + ((!g520) & (g521) & (!g522) & (g523) & (!g524) & (!g525)) + ((!g520) & (g521) & (!g522) & (g523) & (g524) & (!g525)) + ((!g520) & (g521) & (g522) & (!g523) & (!g524) & (!g525)) + ((g520) & (!g521) & (!g522) & (!g523) & (!g524) & (!g525)) + ((g520) & (!g521) & (!g522) & (!g523) & (!g524) & (g525)) + ((g520) & (!g521) & (!g522) & (!g523) & (g524) & (!g525)) + ((g520) & (!g521) & (!g522) & (g523) & (!g524) & (!g525)) + ((g520) & (!g521) & (!g522) & (g523) & (g524) & (!g525)) + ((g520) & (!g521) & (g522) & (!g523) & (!g524) & (!g525)) + ((g520) & (g521) & (!g522) & (!g523) & (!g524) & (!g525)) + ((g520) & (g521) & (!g522) & (!g523) & (g524) & (!g525)) + ((g520) & (g521) & (!g522) & (g523) & (!g524) & (!g525)) + ((g520) & (g521) & (g522) & (!g523) & (!g524) & (!g525)) + ((g520) & (g521) & (g522) & (!g523) & (!g524) & (g525)) + ((g520) & (g521) & (g522) & (!g523) & (g524) & (!g525)) + ((g520) & (g521) & (g522) & (!g523) & (g524) & (g525)) + ((g520) & (g521) & (g522) & (g523) & (!g524) & (!g525)) + ((g520) & (g521) & (g522) & (g523) & (!g524) & (g525)) + ((g520) & (g521) & (g522) & (g523) & (g524) & (!g525)));
	assign g527 = (((!g198) & (!g347) & (!sk[25]) & (!g367) & (g425)) + ((!g198) & (!g347) & (!sk[25]) & (g367) & (g425)) + ((!g198) & (!g347) & (sk[25]) & (!g367) & (!g425)) + ((!g198) & (!g347) & (sk[25]) & (!g367) & (g425)) + ((!g198) & (!g347) & (sk[25]) & (g367) & (!g425)) + ((!g198) & (g347) & (!sk[25]) & (!g367) & (g425)) + ((!g198) & (g347) & (!sk[25]) & (g367) & (g425)) + ((g198) & (!g347) & (!sk[25]) & (!g367) & (!g425)) + ((g198) & (!g347) & (!sk[25]) & (!g367) & (g425)) + ((g198) & (!g347) & (!sk[25]) & (g367) & (!g425)) + ((g198) & (!g347) & (!sk[25]) & (g367) & (g425)) + ((g198) & (!g347) & (sk[25]) & (!g367) & (g425)) + ((g198) & (g347) & (!sk[25]) & (!g367) & (!g425)) + ((g198) & (g347) & (!sk[25]) & (!g367) & (g425)) + ((g198) & (g347) & (!sk[25]) & (g367) & (!g425)) + ((g198) & (g347) & (!sk[25]) & (g367) & (g425)) + ((g198) & (g347) & (sk[25]) & (!g367) & (!g425)) + ((g198) & (g347) & (sk[25]) & (g367) & (!g425)));
	assign g528 = (((!g2) & (!g196) & (!g347) & (g365) & (!g393) & (!g401)) + ((!g2) & (!g196) & (!g347) & (g365) & (!g393) & (g401)) + ((!g2) & (!g196) & (!g347) & (g365) & (g393) & (!g401)) + ((!g2) & (!g196) & (!g347) & (g365) & (g393) & (g401)) + ((!g2) & (!g196) & (g347) & (!g365) & (!g393) & (!g401)) + ((!g2) & (!g196) & (g347) & (!g365) & (!g393) & (g401)) + ((!g2) & (!g196) & (g347) & (!g365) & (g393) & (!g401)) + ((!g2) & (!g196) & (g347) & (!g365) & (g393) & (g401)) + ((!g2) & (!g196) & (g347) & (g365) & (!g393) & (!g401)) + ((!g2) & (!g196) & (g347) & (g365) & (g393) & (!g401)) + ((!g2) & (g196) & (!g347) & (!g365) & (!g393) & (g401)) + ((!g2) & (g196) & (g347) & (g365) & (!g393) & (g401)) + ((g2) & (!g196) & (g347) & (g365) & (!g393) & (!g401)) + ((g2) & (!g196) & (g347) & (g365) & (g393) & (!g401)) + ((g2) & (g196) & (!g347) & (!g365) & (!g393) & (g401)) + ((g2) & (g196) & (!g347) & (g365) & (!g393) & (!g401)) + ((g2) & (g196) & (!g347) & (g365) & (!g393) & (g401)) + ((g2) & (g196) & (g347) & (!g365) & (!g393) & (!g401)) + ((g2) & (g196) & (g347) & (!g365) & (!g393) & (g401)) + ((g2) & (g196) & (g347) & (g365) & (!g393) & (g401)));
	assign g529 = (((!g520) & (!sk[27]) & (g521) & (!g522)) + ((!g520) & (!sk[27]) & (g521) & (g522)) + ((g520) & (!sk[27]) & (g521) & (!g522)) + ((g520) & (!sk[27]) & (g521) & (g522)) + ((g520) & (sk[27]) & (g521) & (g522)));
	assign g530 = (((!g197) & (!sk[28]) & (!g513) & (!g514) & (g515) & (!g516)) + ((!g197) & (!sk[28]) & (!g513) & (!g514) & (g515) & (g516)) + ((!g197) & (!sk[28]) & (!g513) & (g514) & (!g515) & (!g516)) + ((!g197) & (!sk[28]) & (!g513) & (g514) & (!g515) & (g516)) + ((!g197) & (!sk[28]) & (!g513) & (g514) & (g515) & (!g516)) + ((!g197) & (!sk[28]) & (!g513) & (g514) & (g515) & (g516)) + ((!g197) & (!sk[28]) & (g513) & (!g514) & (!g515) & (!g516)) + ((!g197) & (!sk[28]) & (g513) & (!g514) & (!g515) & (g516)) + ((!g197) & (!sk[28]) & (g513) & (!g514) & (g515) & (!g516)) + ((!g197) & (!sk[28]) & (g513) & (!g514) & (g515) & (g516)) + ((!g197) & (!sk[28]) & (g513) & (g514) & (!g515) & (!g516)) + ((!g197) & (!sk[28]) & (g513) & (g514) & (!g515) & (g516)) + ((!g197) & (!sk[28]) & (g513) & (g514) & (g515) & (!g516)) + ((!g197) & (!sk[28]) & (g513) & (g514) & (g515) & (g516)) + ((!g197) & (sk[28]) & (!g513) & (!g514) & (!g515) & (!g516)) + ((!g197) & (sk[28]) & (!g513) & (!g514) & (!g515) & (g516)) + ((!g197) & (sk[28]) & (!g513) & (g514) & (g515) & (!g516)) + ((!g197) & (sk[28]) & (!g513) & (g514) & (g515) & (g516)) + ((!g197) & (sk[28]) & (g513) & (!g514) & (g515) & (!g516)) + ((!g197) & (sk[28]) & (g513) & (!g514) & (g515) & (g516)) + ((!g197) & (sk[28]) & (g513) & (g514) & (!g515) & (!g516)) + ((!g197) & (sk[28]) & (g513) & (g514) & (!g515) & (g516)) + ((g197) & (!sk[28]) & (!g513) & (!g514) & (g515) & (!g516)) + ((g197) & (!sk[28]) & (!g513) & (!g514) & (g515) & (g516)) + ((g197) & (!sk[28]) & (!g513) & (g514) & (!g515) & (!g516)) + ((g197) & (!sk[28]) & (!g513) & (g514) & (!g515) & (g516)) + ((g197) & (!sk[28]) & (!g513) & (g514) & (g515) & (!g516)) + ((g197) & (!sk[28]) & (!g513) & (g514) & (g515) & (g516)) + ((g197) & (!sk[28]) & (g513) & (!g514) & (!g515) & (!g516)) + ((g197) & (!sk[28]) & (g513) & (!g514) & (!g515) & (g516)) + ((g197) & (!sk[28]) & (g513) & (!g514) & (g515) & (!g516)) + ((g197) & (!sk[28]) & (g513) & (!g514) & (g515) & (g516)) + ((g197) & (!sk[28]) & (g513) & (g514) & (!g515) & (!g516)) + ((g197) & (!sk[28]) & (g513) & (g514) & (!g515) & (g516)) + ((g197) & (!sk[28]) & (g513) & (g514) & (g515) & (!g516)) + ((g197) & (!sk[28]) & (g513) & (g514) & (g515) & (g516)) + ((g197) & (sk[28]) & (!g513) & (!g514) & (!g515) & (g516)) + ((g197) & (sk[28]) & (!g513) & (!g514) & (g515) & (!g516)) + ((g197) & (sk[28]) & (!g513) & (g514) & (!g515) & (!g516)) + ((g197) & (sk[28]) & (!g513) & (g514) & (g515) & (g516)) + ((g197) & (sk[28]) & (g513) & (!g514) & (!g515) & (!g516)) + ((g197) & (sk[28]) & (g513) & (!g514) & (g515) & (g516)) + ((g197) & (sk[28]) & (g513) & (g514) & (!g515) & (g516)) + ((g197) & (sk[28]) & (g513) & (g514) & (g515) & (!g516)));
	assign g531 = (((!g516) & (!g526) & (!g527) & (!g528) & (!g529) & (!g530)) + ((!g516) & (!g526) & (!g527) & (!g528) & (!g529) & (g530)) + ((!g516) & (!g526) & (!g527) & (!g528) & (g529) & (g530)) + ((!g516) & (!g526) & (!g527) & (g528) & (!g529) & (g530)) + ((!g516) & (!g526) & (!g527) & (g528) & (g529) & (g530)) + ((!g516) & (!g526) & (g527) & (!g528) & (!g529) & (g530)) + ((!g516) & (!g526) & (g527) & (!g528) & (g529) & (g530)) + ((!g516) & (!g526) & (g527) & (g528) & (!g529) & (g530)) + ((!g516) & (g526) & (!g527) & (!g528) & (!g529) & (!g530)) + ((!g516) & (g526) & (!g527) & (!g528) & (!g529) & (g530)) + ((!g516) & (g526) & (!g527) & (!g528) & (g529) & (!g530)) + ((!g516) & (g526) & (!g527) & (!g528) & (g529) & (g530)) + ((!g516) & (g526) & (!g527) & (g528) & (!g529) & (!g530)) + ((!g516) & (g526) & (!g527) & (g528) & (!g529) & (g530)) + ((!g516) & (g526) & (!g527) & (g528) & (g529) & (g530)) + ((!g516) & (g526) & (g527) & (!g528) & (!g529) & (!g530)) + ((!g516) & (g526) & (g527) & (!g528) & (!g529) & (g530)) + ((!g516) & (g526) & (g527) & (!g528) & (g529) & (g530)) + ((!g516) & (g526) & (g527) & (g528) & (!g529) & (g530)) + ((!g516) & (g526) & (g527) & (g528) & (g529) & (g530)) + ((g516) & (!g526) & (!g527) & (!g528) & (!g529) & (g530)) + ((g516) & (!g526) & (!g527) & (!g528) & (g529) & (g530)) + ((g516) & (!g526) & (!g527) & (g528) & (!g529) & (g530)) + ((g516) & (!g526) & (g527) & (!g528) & (!g529) & (g530)) + ((g516) & (g526) & (!g527) & (!g528) & (!g529) & (!g530)) + ((g516) & (g526) & (!g527) & (!g528) & (!g529) & (g530)) + ((g516) & (g526) & (!g527) & (!g528) & (g529) & (g530)) + ((g516) & (g526) & (!g527) & (g528) & (!g529) & (g530)) + ((g516) & (g526) & (!g527) & (g528) & (g529) & (g530)) + ((g516) & (g526) & (g527) & (!g528) & (!g529) & (g530)) + ((g516) & (g526) & (g527) & (!g528) & (g529) & (g530)) + ((g516) & (g526) & (g527) & (g528) & (!g529) & (g530)));
	assign g532 = (((!g504) & (!g505) & (sk[30]) & (!g506)) + ((!g504) & (g505) & (!sk[30]) & (!g506)) + ((!g504) & (g505) & (!sk[30]) & (g506)) + ((!g504) & (g505) & (sk[30]) & (g506)) + ((g504) & (!g505) & (sk[30]) & (g506)) + ((g504) & (g505) & (!sk[30]) & (!g506)) + ((g504) & (g505) & (!sk[30]) & (g506)) + ((g504) & (g505) & (sk[30]) & (!g506)));
	assign g533 = (((!g504) & (!g505) & (!g506) & (!g507) & (!g510) & (!g511)) + ((!g504) & (!g505) & (!g506) & (!g507) & (g510) & (g511)) + ((!g504) & (!g505) & (!g506) & (g507) & (!g510) & (g511)) + ((!g504) & (!g505) & (!g506) & (g507) & (g510) & (!g511)) + ((!g504) & (!g505) & (g506) & (!g507) & (!g510) & (!g511)) + ((!g504) & (!g505) & (g506) & (!g507) & (g510) & (g511)) + ((!g504) & (!g505) & (g506) & (g507) & (!g510) & (g511)) + ((!g504) & (!g505) & (g506) & (g507) & (g510) & (!g511)) + ((!g504) & (g505) & (!g506) & (!g507) & (!g510) & (!g511)) + ((!g504) & (g505) & (!g506) & (!g507) & (g510) & (g511)) + ((!g504) & (g505) & (!g506) & (g507) & (!g510) & (g511)) + ((!g504) & (g505) & (!g506) & (g507) & (g510) & (!g511)) + ((!g504) & (g505) & (g506) & (!g507) & (!g510) & (g511)) + ((!g504) & (g505) & (g506) & (!g507) & (g510) & (!g511)) + ((!g504) & (g505) & (g506) & (g507) & (!g510) & (!g511)) + ((!g504) & (g505) & (g506) & (g507) & (g510) & (g511)) + ((g504) & (!g505) & (!g506) & (!g507) & (!g510) & (!g511)) + ((g504) & (!g505) & (!g506) & (!g507) & (g510) & (g511)) + ((g504) & (!g505) & (!g506) & (g507) & (!g510) & (g511)) + ((g504) & (!g505) & (!g506) & (g507) & (g510) & (!g511)) + ((g504) & (!g505) & (g506) & (!g507) & (!g510) & (g511)) + ((g504) & (!g505) & (g506) & (!g507) & (g510) & (!g511)) + ((g504) & (!g505) & (g506) & (g507) & (!g510) & (!g511)) + ((g504) & (!g505) & (g506) & (g507) & (g510) & (g511)) + ((g504) & (g505) & (!g506) & (!g507) & (!g510) & (g511)) + ((g504) & (g505) & (!g506) & (!g507) & (g510) & (!g511)) + ((g504) & (g505) & (!g506) & (g507) & (!g510) & (!g511)) + ((g504) & (g505) & (!g506) & (g507) & (g510) & (g511)) + ((g504) & (g505) & (g506) & (!g507) & (!g510) & (g511)) + ((g504) & (g505) & (g506) & (!g507) & (g510) & (!g511)) + ((g504) & (g505) & (g506) & (g507) & (!g510) & (!g511)) + ((g504) & (g505) & (g506) & (g507) & (g510) & (g511)));
	assign g534 = (((!g517) & (!g518) & (!g519) & (!g531) & (!g532) & (g533)) + ((!g517) & (!g518) & (!g519) & (!g531) & (g532) & (!g533)) + ((!g517) & (!g518) & (!g519) & (!g531) & (g532) & (g533)) + ((!g517) & (!g518) & (!g519) & (g531) & (!g532) & (!g533)) + ((!g517) & (!g518) & (!g519) & (g531) & (!g532) & (g533)) + ((!g517) & (!g518) & (!g519) & (g531) & (g532) & (!g533)) + ((!g517) & (!g518) & (!g519) & (g531) & (g532) & (g533)) + ((!g517) & (!g518) & (g519) & (!g531) & (!g532) & (g533)) + ((!g517) & (!g518) & (g519) & (!g531) & (g532) & (g533)) + ((!g517) & (!g518) & (g519) & (g531) & (!g532) & (g533)) + ((!g517) & (!g518) & (g519) & (g531) & (g532) & (!g533)) + ((!g517) & (!g518) & (g519) & (g531) & (g532) & (g533)) + ((!g517) & (g518) & (!g519) & (!g531) & (!g532) & (g533)) + ((!g517) & (g518) & (!g519) & (!g531) & (g532) & (g533)) + ((!g517) & (g518) & (!g519) & (g531) & (!g532) & (g533)) + ((!g517) & (g518) & (!g519) & (g531) & (g532) & (!g533)) + ((!g517) & (g518) & (!g519) & (g531) & (g532) & (g533)) + ((!g517) & (g518) & (g519) & (!g531) & (g532) & (g533)) + ((!g517) & (g518) & (g519) & (g531) & (!g532) & (g533)) + ((!g517) & (g518) & (g519) & (g531) & (g532) & (g533)) + ((g517) & (!g518) & (!g519) & (!g531) & (!g532) & (g533)) + ((g517) & (!g518) & (!g519) & (!g531) & (g532) & (g533)) + ((g517) & (!g518) & (!g519) & (g531) & (!g532) & (g533)) + ((g517) & (!g518) & (!g519) & (g531) & (g532) & (!g533)) + ((g517) & (!g518) & (!g519) & (g531) & (g532) & (g533)) + ((g517) & (!g518) & (g519) & (!g531) & (g532) & (g533)) + ((g517) & (!g518) & (g519) & (g531) & (!g532) & (g533)) + ((g517) & (!g518) & (g519) & (g531) & (g532) & (g533)) + ((g517) & (g518) & (!g519) & (!g531) & (g532) & (g533)) + ((g517) & (g518) & (!g519) & (g531) & (!g532) & (g533)) + ((g517) & (g518) & (!g519) & (g531) & (g532) & (g533)) + ((g517) & (g518) & (g519) & (g531) & (g532) & (g533)));
	assign g535 = (((!sk[33]) & (!g492) & (!g414) & (!g493) & (g494) & (!g495)) + ((!sk[33]) & (!g492) & (!g414) & (!g493) & (g494) & (g495)) + ((!sk[33]) & (!g492) & (!g414) & (g493) & (!g494) & (!g495)) + ((!sk[33]) & (!g492) & (!g414) & (g493) & (!g494) & (g495)) + ((!sk[33]) & (!g492) & (!g414) & (g493) & (g494) & (!g495)) + ((!sk[33]) & (!g492) & (!g414) & (g493) & (g494) & (g495)) + ((!sk[33]) & (!g492) & (g414) & (!g493) & (!g494) & (!g495)) + ((!sk[33]) & (!g492) & (g414) & (!g493) & (!g494) & (g495)) + ((!sk[33]) & (!g492) & (g414) & (!g493) & (g494) & (!g495)) + ((!sk[33]) & (!g492) & (g414) & (!g493) & (g494) & (g495)) + ((!sk[33]) & (!g492) & (g414) & (g493) & (!g494) & (!g495)) + ((!sk[33]) & (!g492) & (g414) & (g493) & (!g494) & (g495)) + ((!sk[33]) & (!g492) & (g414) & (g493) & (g494) & (!g495)) + ((!sk[33]) & (!g492) & (g414) & (g493) & (g494) & (g495)) + ((!sk[33]) & (g492) & (!g414) & (!g493) & (g494) & (!g495)) + ((!sk[33]) & (g492) & (!g414) & (!g493) & (g494) & (g495)) + ((!sk[33]) & (g492) & (!g414) & (g493) & (!g494) & (!g495)) + ((!sk[33]) & (g492) & (!g414) & (g493) & (!g494) & (g495)) + ((!sk[33]) & (g492) & (!g414) & (g493) & (g494) & (!g495)) + ((!sk[33]) & (g492) & (!g414) & (g493) & (g494) & (g495)) + ((!sk[33]) & (g492) & (g414) & (!g493) & (!g494) & (!g495)) + ((!sk[33]) & (g492) & (g414) & (!g493) & (!g494) & (g495)) + ((!sk[33]) & (g492) & (g414) & (!g493) & (g494) & (!g495)) + ((!sk[33]) & (g492) & (g414) & (!g493) & (g494) & (g495)) + ((!sk[33]) & (g492) & (g414) & (g493) & (!g494) & (!g495)) + ((!sk[33]) & (g492) & (g414) & (g493) & (!g494) & (g495)) + ((!sk[33]) & (g492) & (g414) & (g493) & (g494) & (!g495)) + ((!sk[33]) & (g492) & (g414) & (g493) & (g494) & (g495)) + ((sk[33]) & (!g492) & (!g414) & (!g493) & (!g494) & (g495)) + ((sk[33]) & (!g492) & (!g414) & (!g493) & (g494) & (g495)) + ((sk[33]) & (!g492) & (!g414) & (g493) & (!g494) & (g495)) + ((sk[33]) & (!g492) & (!g414) & (g493) & (g494) & (!g495)) + ((sk[33]) & (!g492) & (g414) & (!g493) & (!g494) & (g495)) + ((sk[33]) & (!g492) & (g414) & (!g493) & (g494) & (g495)) + ((sk[33]) & (!g492) & (g414) & (g493) & (!g494) & (g495)) + ((sk[33]) & (!g492) & (g414) & (g493) & (g494) & (!g495)) + ((sk[33]) & (g492) & (!g414) & (!g493) & (!g494) & (g495)) + ((sk[33]) & (g492) & (!g414) & (!g493) & (g494) & (g495)) + ((sk[33]) & (g492) & (!g414) & (g493) & (!g494) & (g495)) + ((sk[33]) & (g492) & (!g414) & (g493) & (g494) & (!g495)) + ((sk[33]) & (g492) & (g414) & (!g493) & (!g494) & (!g495)) + ((sk[33]) & (g492) & (g414) & (!g493) & (g494) & (!g495)) + ((sk[33]) & (g492) & (g414) & (g493) & (!g494) & (!g495)) + ((sk[33]) & (g492) & (g414) & (g493) & (g494) & (g495)));
	assign g536 = (((!g508) & (!sk[34]) & (g509) & (!g511)) + ((!g508) & (!sk[34]) & (g509) & (g511)) + ((!g508) & (sk[34]) & (g509) & (g511)) + ((g508) & (!sk[34]) & (g509) & (!g511)) + ((g508) & (!sk[34]) & (g509) & (g511)) + ((g508) & (sk[34]) & (!g509) & (g511)) + ((g508) & (sk[34]) & (g509) & (!g511)) + ((g508) & (sk[34]) & (g509) & (g511)));
	assign g537 = (((!g497) & (!g498) & (sk[35]) & (g499)) + ((!g497) & (g498) & (!sk[35]) & (!g499)) + ((!g497) & (g498) & (!sk[35]) & (g499)) + ((!g497) & (g498) & (sk[35]) & (!g499)) + ((g497) & (!g498) & (sk[35]) & (!g499)) + ((g497) & (g498) & (!sk[35]) & (!g499)) + ((g497) & (g498) & (!sk[35]) & (g499)) + ((g497) & (g498) & (sk[35]) & (g499)));
	assign g538 = (((!sk[36]) & (!g491) & (!g482) & (!g496) & (g500) & (!g502)) + ((!sk[36]) & (!g491) & (!g482) & (!g496) & (g500) & (g502)) + ((!sk[36]) & (!g491) & (!g482) & (g496) & (!g500) & (!g502)) + ((!sk[36]) & (!g491) & (!g482) & (g496) & (!g500) & (g502)) + ((!sk[36]) & (!g491) & (!g482) & (g496) & (g500) & (!g502)) + ((!sk[36]) & (!g491) & (!g482) & (g496) & (g500) & (g502)) + ((!sk[36]) & (!g491) & (g482) & (!g496) & (!g500) & (!g502)) + ((!sk[36]) & (!g491) & (g482) & (!g496) & (!g500) & (g502)) + ((!sk[36]) & (!g491) & (g482) & (!g496) & (g500) & (!g502)) + ((!sk[36]) & (!g491) & (g482) & (!g496) & (g500) & (g502)) + ((!sk[36]) & (!g491) & (g482) & (g496) & (!g500) & (!g502)) + ((!sk[36]) & (!g491) & (g482) & (g496) & (!g500) & (g502)) + ((!sk[36]) & (!g491) & (g482) & (g496) & (g500) & (!g502)) + ((!sk[36]) & (!g491) & (g482) & (g496) & (g500) & (g502)) + ((!sk[36]) & (g491) & (!g482) & (!g496) & (g500) & (!g502)) + ((!sk[36]) & (g491) & (!g482) & (!g496) & (g500) & (g502)) + ((!sk[36]) & (g491) & (!g482) & (g496) & (!g500) & (!g502)) + ((!sk[36]) & (g491) & (!g482) & (g496) & (!g500) & (g502)) + ((!sk[36]) & (g491) & (!g482) & (g496) & (g500) & (!g502)) + ((!sk[36]) & (g491) & (!g482) & (g496) & (g500) & (g502)) + ((!sk[36]) & (g491) & (g482) & (!g496) & (!g500) & (!g502)) + ((!sk[36]) & (g491) & (g482) & (!g496) & (!g500) & (g502)) + ((!sk[36]) & (g491) & (g482) & (!g496) & (g500) & (!g502)) + ((!sk[36]) & (g491) & (g482) & (!g496) & (g500) & (g502)) + ((!sk[36]) & (g491) & (g482) & (g496) & (!g500) & (!g502)) + ((!sk[36]) & (g491) & (g482) & (g496) & (!g500) & (g502)) + ((!sk[36]) & (g491) & (g482) & (g496) & (g500) & (!g502)) + ((!sk[36]) & (g491) & (g482) & (g496) & (g500) & (g502)) + ((sk[36]) & (!g491) & (!g482) & (!g496) & (!g500) & (g502)) + ((sk[36]) & (!g491) & (!g482) & (!g496) & (g500) & (!g502)) + ((sk[36]) & (!g491) & (!g482) & (g496) & (!g500) & (!g502)) + ((sk[36]) & (!g491) & (!g482) & (g496) & (g500) & (g502)) + ((sk[36]) & (!g491) & (g482) & (!g496) & (!g500) & (!g502)) + ((sk[36]) & (!g491) & (g482) & (!g496) & (g500) & (g502)) + ((sk[36]) & (!g491) & (g482) & (g496) & (!g500) & (g502)) + ((sk[36]) & (!g491) & (g482) & (g496) & (g500) & (!g502)) + ((sk[36]) & (g491) & (!g482) & (!g496) & (!g500) & (!g502)) + ((sk[36]) & (g491) & (!g482) & (!g496) & (g500) & (g502)) + ((sk[36]) & (g491) & (!g482) & (g496) & (!g500) & (g502)) + ((sk[36]) & (g491) & (!g482) & (g496) & (g500) & (!g502)) + ((sk[36]) & (g491) & (g482) & (!g496) & (!g500) & (g502)) + ((sk[36]) & (g491) & (g482) & (!g496) & (g500) & (!g502)) + ((sk[36]) & (g491) & (g482) & (g496) & (!g500) & (!g502)) + ((sk[36]) & (g491) & (g482) & (g496) & (g500) & (g502)));
	assign g539 = (((!g512) & (!g534) & (!g535) & (!g536) & (!g537) & (!g538)) + ((!g512) & (!g534) & (!g535) & (!g536) & (!g537) & (g538)) + ((!g512) & (!g534) & (!g535) & (!g536) & (g537) & (g538)) + ((!g512) & (!g534) & (!g535) & (g536) & (!g537) & (g538)) + ((!g512) & (!g534) & (!g535) & (g536) & (g537) & (g538)) + ((!g512) & (!g534) & (g535) & (!g536) & (!g537) & (g538)) + ((!g512) & (!g534) & (g535) & (!g536) & (g537) & (g538)) + ((!g512) & (!g534) & (g535) & (g536) & (!g537) & (g538)) + ((!g512) & (g534) & (!g535) & (!g536) & (!g537) & (!g538)) + ((!g512) & (g534) & (!g535) & (!g536) & (!g537) & (g538)) + ((!g512) & (g534) & (!g535) & (!g536) & (g537) & (!g538)) + ((!g512) & (g534) & (!g535) & (!g536) & (g537) & (g538)) + ((!g512) & (g534) & (!g535) & (g536) & (!g537) & (!g538)) + ((!g512) & (g534) & (!g535) & (g536) & (!g537) & (g538)) + ((!g512) & (g534) & (!g535) & (g536) & (g537) & (g538)) + ((!g512) & (g534) & (g535) & (!g536) & (!g537) & (!g538)) + ((!g512) & (g534) & (g535) & (!g536) & (!g537) & (g538)) + ((!g512) & (g534) & (g535) & (!g536) & (g537) & (g538)) + ((!g512) & (g534) & (g535) & (g536) & (!g537) & (g538)) + ((!g512) & (g534) & (g535) & (g536) & (g537) & (g538)) + ((g512) & (!g534) & (!g535) & (!g536) & (!g537) & (g538)) + ((g512) & (!g534) & (!g535) & (!g536) & (g537) & (g538)) + ((g512) & (!g534) & (!g535) & (g536) & (!g537) & (g538)) + ((g512) & (!g534) & (g535) & (!g536) & (!g537) & (g538)) + ((g512) & (g534) & (!g535) & (!g536) & (!g537) & (!g538)) + ((g512) & (g534) & (!g535) & (!g536) & (!g537) & (g538)) + ((g512) & (g534) & (!g535) & (!g536) & (g537) & (g538)) + ((g512) & (g534) & (!g535) & (g536) & (!g537) & (g538)) + ((g512) & (g534) & (!g535) & (g536) & (g537) & (g538)) + ((g512) & (g534) & (g535) & (!g536) & (!g537) & (g538)) + ((g512) & (g534) & (g535) & (!g536) & (g537) & (g538)) + ((g512) & (g534) & (g535) & (g536) & (!g537) & (g538)));
	assign g540 = (((!g466) & (!g467) & (!g497) & (g498) & (g499) & (g501)) + ((!g466) & (!g467) & (g497) & (!g498) & (g499) & (g501)) + ((!g466) & (!g467) & (g497) & (g498) & (!g499) & (g501)) + ((!g466) & (!g467) & (g497) & (g498) & (g499) & (g501)) + ((!g466) & (g467) & (!g497) & (!g498) & (!g499) & (g501)) + ((!g466) & (g467) & (!g497) & (!g498) & (g499) & (g501)) + ((!g466) & (g467) & (!g497) & (g498) & (!g499) & (g501)) + ((!g466) & (g467) & (!g497) & (g498) & (g499) & (!g501)) + ((!g466) & (g467) & (!g497) & (g498) & (g499) & (g501)) + ((!g466) & (g467) & (g497) & (!g498) & (!g499) & (g501)) + ((!g466) & (g467) & (g497) & (!g498) & (g499) & (!g501)) + ((!g466) & (g467) & (g497) & (!g498) & (g499) & (g501)) + ((!g466) & (g467) & (g497) & (g498) & (!g499) & (!g501)) + ((!g466) & (g467) & (g497) & (g498) & (!g499) & (g501)) + ((!g466) & (g467) & (g497) & (g498) & (g499) & (!g501)) + ((!g466) & (g467) & (g497) & (g498) & (g499) & (g501)) + ((g466) & (!g467) & (!g497) & (!g498) & (!g499) & (g501)) + ((g466) & (!g467) & (!g497) & (!g498) & (g499) & (g501)) + ((g466) & (!g467) & (!g497) & (g498) & (!g499) & (g501)) + ((g466) & (!g467) & (!g497) & (g498) & (g499) & (!g501)) + ((g466) & (!g467) & (!g497) & (g498) & (g499) & (g501)) + ((g466) & (!g467) & (g497) & (!g498) & (!g499) & (g501)) + ((g466) & (!g467) & (g497) & (!g498) & (g499) & (!g501)) + ((g466) & (!g467) & (g497) & (!g498) & (g499) & (g501)) + ((g466) & (!g467) & (g497) & (g498) & (!g499) & (!g501)) + ((g466) & (!g467) & (g497) & (g498) & (!g499) & (g501)) + ((g466) & (!g467) & (g497) & (g498) & (g499) & (!g501)) + ((g466) & (!g467) & (g497) & (g498) & (g499) & (g501)) + ((g466) & (g467) & (!g497) & (g498) & (g499) & (g501)) + ((g466) & (g467) & (g497) & (!g498) & (g499) & (g501)) + ((g466) & (g467) & (g497) & (g498) & (!g499) & (g501)) + ((g466) & (g467) & (g497) & (g498) & (g499) & (g501)));
	assign g541 = (((!g471) & (!g472) & (sk[39]) & (g473)) + ((!g471) & (g472) & (!sk[39]) & (!g473)) + ((!g471) & (g472) & (!sk[39]) & (g473)) + ((!g471) & (g472) & (sk[39]) & (!g473)) + ((g471) & (!g472) & (sk[39]) & (!g473)) + ((g471) & (g472) & (!sk[39]) & (!g473)) + ((g471) & (g472) & (!sk[39]) & (g473)) + ((g471) & (g472) & (sk[39]) & (g473)));
	assign g542 = (((!g479) & (!g483) & (!g484) & (!g540) & (sk[40]) & (g541)) + ((!g479) & (!g483) & (!g484) & (g540) & (!sk[40]) & (!g541)) + ((!g479) & (!g483) & (!g484) & (g540) & (!sk[40]) & (g541)) + ((!g479) & (!g483) & (!g484) & (g540) & (sk[40]) & (!g541)) + ((!g479) & (!g483) & (g484) & (!g540) & (!sk[40]) & (!g541)) + ((!g479) & (!g483) & (g484) & (!g540) & (!sk[40]) & (g541)) + ((!g479) & (!g483) & (g484) & (!g540) & (sk[40]) & (!g541)) + ((!g479) & (!g483) & (g484) & (g540) & (!sk[40]) & (!g541)) + ((!g479) & (!g483) & (g484) & (g540) & (!sk[40]) & (g541)) + ((!g479) & (!g483) & (g484) & (g540) & (sk[40]) & (g541)) + ((!g479) & (g483) & (!g484) & (!g540) & (!sk[40]) & (!g541)) + ((!g479) & (g483) & (!g484) & (!g540) & (!sk[40]) & (g541)) + ((!g479) & (g483) & (!g484) & (!g540) & (sk[40]) & (!g541)) + ((!g479) & (g483) & (!g484) & (g540) & (!sk[40]) & (!g541)) + ((!g479) & (g483) & (!g484) & (g540) & (!sk[40]) & (g541)) + ((!g479) & (g483) & (!g484) & (g540) & (sk[40]) & (g541)) + ((!g479) & (g483) & (g484) & (!g540) & (!sk[40]) & (!g541)) + ((!g479) & (g483) & (g484) & (!g540) & (!sk[40]) & (g541)) + ((!g479) & (g483) & (g484) & (!g540) & (sk[40]) & (g541)) + ((!g479) & (g483) & (g484) & (g540) & (!sk[40]) & (!g541)) + ((!g479) & (g483) & (g484) & (g540) & (!sk[40]) & (g541)) + ((!g479) & (g483) & (g484) & (g540) & (sk[40]) & (!g541)) + ((g479) & (!g483) & (!g484) & (!g540) & (sk[40]) & (!g541)) + ((g479) & (!g483) & (!g484) & (g540) & (!sk[40]) & (!g541)) + ((g479) & (!g483) & (!g484) & (g540) & (!sk[40]) & (g541)) + ((g479) & (!g483) & (!g484) & (g540) & (sk[40]) & (g541)) + ((g479) & (!g483) & (g484) & (!g540) & (!sk[40]) & (!g541)) + ((g479) & (!g483) & (g484) & (!g540) & (!sk[40]) & (g541)) + ((g479) & (!g483) & (g484) & (!g540) & (sk[40]) & (g541)) + ((g479) & (!g483) & (g484) & (g540) & (!sk[40]) & (!g541)) + ((g479) & (!g483) & (g484) & (g540) & (!sk[40]) & (g541)) + ((g479) & (!g483) & (g484) & (g540) & (sk[40]) & (!g541)) + ((g479) & (g483) & (!g484) & (!g540) & (!sk[40]) & (!g541)) + ((g479) & (g483) & (!g484) & (!g540) & (!sk[40]) & (g541)) + ((g479) & (g483) & (!g484) & (!g540) & (sk[40]) & (g541)) + ((g479) & (g483) & (!g484) & (g540) & (!sk[40]) & (!g541)) + ((g479) & (g483) & (!g484) & (g540) & (!sk[40]) & (g541)) + ((g479) & (g483) & (!g484) & (g540) & (sk[40]) & (!g541)) + ((g479) & (g483) & (g484) & (!g540) & (!sk[40]) & (!g541)) + ((g479) & (g483) & (g484) & (!g540) & (!sk[40]) & (g541)) + ((g479) & (g483) & (g484) & (!g540) & (sk[40]) & (!g541)) + ((g479) & (g483) & (g484) & (g540) & (!sk[40]) & (!g541)) + ((g479) & (g483) & (g484) & (g540) & (!sk[40]) & (g541)) + ((g479) & (g483) & (g484) & (g540) & (sk[40]) & (g541)));
	assign g543 = (((!g479) & (!g483) & (!g484) & (!g540) & (sk[41]) & (!g541)) + ((!g479) & (!g483) & (!g484) & (g540) & (!sk[41]) & (!g541)) + ((!g479) & (!g483) & (!g484) & (g540) & (!sk[41]) & (g541)) + ((!g479) & (!g483) & (g484) & (!g540) & (!sk[41]) & (!g541)) + ((!g479) & (!g483) & (g484) & (!g540) & (!sk[41]) & (g541)) + ((!g479) & (!g483) & (g484) & (!g540) & (sk[41]) & (!g541)) + ((!g479) & (!g483) & (g484) & (!g540) & (sk[41]) & (g541)) + ((!g479) & (!g483) & (g484) & (g540) & (!sk[41]) & (!g541)) + ((!g479) & (!g483) & (g484) & (g540) & (!sk[41]) & (g541)) + ((!g479) & (!g483) & (g484) & (g540) & (sk[41]) & (!g541)) + ((!g479) & (g483) & (!g484) & (!g540) & (!sk[41]) & (!g541)) + ((!g479) & (g483) & (!g484) & (!g540) & (!sk[41]) & (g541)) + ((!g479) & (g483) & (!g484) & (!g540) & (sk[41]) & (!g541)) + ((!g479) & (g483) & (!g484) & (!g540) & (sk[41]) & (g541)) + ((!g479) & (g483) & (!g484) & (g540) & (!sk[41]) & (!g541)) + ((!g479) & (g483) & (!g484) & (g540) & (!sk[41]) & (g541)) + ((!g479) & (g483) & (!g484) & (g540) & (sk[41]) & (!g541)) + ((!g479) & (g483) & (g484) & (!g540) & (!sk[41]) & (!g541)) + ((!g479) & (g483) & (g484) & (!g540) & (!sk[41]) & (g541)) + ((!g479) & (g483) & (g484) & (!g540) & (sk[41]) & (!g541)) + ((!g479) & (g483) & (g484) & (g540) & (!sk[41]) & (!g541)) + ((!g479) & (g483) & (g484) & (g540) & (!sk[41]) & (g541)) + ((g479) & (!g483) & (!g484) & (!g540) & (sk[41]) & (!g541)) + ((g479) & (!g483) & (!g484) & (!g540) & (sk[41]) & (g541)) + ((g479) & (!g483) & (!g484) & (g540) & (!sk[41]) & (!g541)) + ((g479) & (!g483) & (!g484) & (g540) & (!sk[41]) & (g541)) + ((g479) & (!g483) & (!g484) & (g540) & (sk[41]) & (!g541)) + ((g479) & (!g483) & (g484) & (!g540) & (!sk[41]) & (!g541)) + ((g479) & (!g483) & (g484) & (!g540) & (!sk[41]) & (g541)) + ((g479) & (!g483) & (g484) & (!g540) & (sk[41]) & (!g541)) + ((g479) & (!g483) & (g484) & (g540) & (!sk[41]) & (!g541)) + ((g479) & (!g483) & (g484) & (g540) & (!sk[41]) & (g541)) + ((g479) & (g483) & (!g484) & (!g540) & (!sk[41]) & (!g541)) + ((g479) & (g483) & (!g484) & (!g540) & (!sk[41]) & (g541)) + ((g479) & (g483) & (!g484) & (!g540) & (sk[41]) & (!g541)) + ((g479) & (g483) & (!g484) & (g540) & (!sk[41]) & (!g541)) + ((g479) & (g483) & (!g484) & (g540) & (!sk[41]) & (g541)) + ((g479) & (g483) & (g484) & (!g540) & (!sk[41]) & (!g541)) + ((g479) & (g483) & (g484) & (!g540) & (!sk[41]) & (g541)) + ((g479) & (g483) & (g484) & (!g540) & (sk[41]) & (!g541)) + ((g479) & (g483) & (g484) & (!g540) & (sk[41]) & (g541)) + ((g479) & (g483) & (g484) & (g540) & (!sk[41]) & (!g541)) + ((g479) & (g483) & (g484) & (g540) & (!sk[41]) & (g541)) + ((g479) & (g483) & (g484) & (g540) & (sk[41]) & (!g541)));
	assign g544 = (((!g485) & (!g486) & (sk[42]) & (!g487)) + ((!g485) & (g486) & (!sk[42]) & (!g487)) + ((!g485) & (g486) & (!sk[42]) & (g487)) + ((!g485) & (g486) & (sk[42]) & (g487)) + ((g485) & (!g486) & (sk[42]) & (g487)) + ((g485) & (g486) & (!sk[42]) & (!g487)) + ((g485) & (g486) & (!sk[42]) & (g487)) + ((g485) & (g486) & (sk[42]) & (!g487)));
	assign g545 = (((g490) & (!g503) & (!g539) & (!g542) & (!g543) & (!g544)) + ((g490) & (!g503) & (!g539) & (!g542) & (!g543) & (g544)) + ((g490) & (!g503) & (!g539) & (!g542) & (g543) & (!g544)) + ((g490) & (!g503) & (!g539) & (g542) & (!g543) & (!g544)) + ((g490) & (!g503) & (g539) & (!g542) & (!g543) & (!g544)) + ((g490) & (!g503) & (g539) & (g542) & (!g543) & (!g544)) + ((g490) & (g503) & (!g539) & (!g542) & (!g543) & (!g544)) + ((g490) & (g503) & (!g539) & (!g542) & (!g543) & (g544)) + ((g490) & (g503) & (!g539) & (!g542) & (g543) & (!g544)) + ((g490) & (g503) & (!g539) & (g542) & (!g543) & (!g544)) + ((g490) & (g503) & (!g539) & (g542) & (!g543) & (g544)) + ((g490) & (g503) & (!g539) & (g542) & (g543) & (!g544)) + ((g490) & (g503) & (g539) & (!g542) & (!g543) & (!g544)) + ((g490) & (g503) & (g539) & (!g542) & (!g543) & (g544)) + ((g490) & (g503) & (g539) & (!g542) & (g543) & (!g544)) + ((g490) & (g503) & (g539) & (g542) & (!g543) & (!g544)));
	assign g546 = (((!g463) & (!g464) & (!g477) & (!g478) & (!g489) & (!g545)) + ((!g463) & (!g464) & (!g477) & (!g478) & (!g489) & (g545)) + ((!g463) & (!g464) & (!g477) & (!g478) & (g489) & (!g545)) + ((!g463) & (!g464) & (!g477) & (!g478) & (g489) & (g545)) + ((!g463) & (!g464) & (!g477) & (g478) & (!g489) & (!g545)) + ((!g463) & (!g464) & (!g477) & (g478) & (!g489) & (g545)) + ((!g463) & (!g464) & (!g477) & (g478) & (g489) & (!g545)) + ((!g463) & (!g464) & (!g477) & (g478) & (g489) & (g545)) + ((!g463) & (!g464) & (g477) & (!g478) & (!g489) & (!g545)) + ((!g463) & (!g464) & (g477) & (!g478) & (!g489) & (g545)) + ((!g463) & (!g464) & (g477) & (!g478) & (g489) & (!g545)) + ((!g463) & (!g464) & (g477) & (!g478) & (g489) & (g545)) + ((!g463) & (!g464) & (g477) & (g478) & (!g489) & (!g545)) + ((!g463) & (!g464) & (g477) & (g478) & (!g489) & (g545)) + ((!g463) & (!g464) & (g477) & (g478) & (g489) & (!g545)) + ((!g463) & (!g464) & (g477) & (g478) & (g489) & (g545)) + ((!g463) & (g464) & (!g477) & (!g478) & (!g489) & (!g545)) + ((!g463) & (g464) & (!g477) & (!g478) & (!g489) & (g545)) + ((!g463) & (g464) & (!g477) & (!g478) & (g489) & (!g545)) + ((!g463) & (g464) & (!g477) & (!g478) & (g489) & (g545)) + ((!g463) & (g464) & (!g477) & (g478) & (!g489) & (!g545)) + ((!g463) & (g464) & (g477) & (!g478) & (!g489) & (!g545)) + ((g463) & (!g464) & (!g477) & (!g478) & (!g489) & (!g545)) + ((g463) & (!g464) & (!g477) & (!g478) & (!g489) & (g545)) + ((g463) & (!g464) & (!g477) & (!g478) & (g489) & (!g545)) + ((g463) & (!g464) & (!g477) & (!g478) & (g489) & (g545)) + ((g463) & (!g464) & (!g477) & (g478) & (!g489) & (!g545)) + ((g463) & (!g464) & (g477) & (!g478) & (!g489) & (!g545)));
	assign g547 = (((g413) & (!g440) & (g441) & (!g454) & (g455) & (!g546)) + ((g413) & (!g440) & (g441) & (g454) & (!g455) & (!g546)) + ((g413) & (!g440) & (g441) & (g454) & (g455) & (!g546)) + ((g413) & (!g440) & (g441) & (g454) & (g455) & (g546)) + ((g413) & (g440) & (!g441) & (!g454) & (g455) & (!g546)) + ((g413) & (g440) & (!g441) & (g454) & (!g455) & (!g546)) + ((g413) & (g440) & (!g441) & (g454) & (g455) & (!g546)) + ((g413) & (g440) & (!g441) & (g454) & (g455) & (g546)) + ((g413) & (g440) & (g441) & (!g454) & (!g455) & (!g546)) + ((g413) & (g440) & (g441) & (!g454) & (!g455) & (g546)) + ((g413) & (g440) & (g441) & (!g454) & (g455) & (!g546)) + ((g413) & (g440) & (g441) & (!g454) & (g455) & (g546)) + ((g413) & (g440) & (g441) & (g454) & (!g455) & (!g546)) + ((g413) & (g440) & (g441) & (g454) & (!g455) & (g546)) + ((g413) & (g440) & (g441) & (g454) & (g455) & (!g546)) + ((g413) & (g440) & (g441) & (g454) & (g455) & (g546)));
	assign g548 = (((!g376) & (!g377) & (!g387) & (!g388) & (!g412) & (!g547)) + ((!g376) & (!g377) & (!g387) & (!g388) & (!g412) & (g547)) + ((!g376) & (!g377) & (!g387) & (!g388) & (g412) & (!g547)) + ((!g376) & (!g377) & (!g387) & (!g388) & (g412) & (g547)) + ((!g376) & (!g377) & (!g387) & (g388) & (!g412) & (!g547)) + ((!g376) & (!g377) & (g387) & (!g388) & (!g412) & (!g547)) + ((!g376) & (g377) & (!g387) & (!g388) & (!g412) & (!g547)) + ((!g376) & (g377) & (!g387) & (!g388) & (!g412) & (g547)) + ((!g376) & (g377) & (!g387) & (!g388) & (g412) & (!g547)) + ((!g376) & (g377) & (!g387) & (!g388) & (g412) & (g547)) + ((!g376) & (g377) & (!g387) & (g388) & (!g412) & (!g547)) + ((!g376) & (g377) & (!g387) & (g388) & (!g412) & (g547)) + ((!g376) & (g377) & (!g387) & (g388) & (g412) & (!g547)) + ((!g376) & (g377) & (!g387) & (g388) & (g412) & (g547)) + ((!g376) & (g377) & (g387) & (!g388) & (!g412) & (!g547)) + ((!g376) & (g377) & (g387) & (!g388) & (!g412) & (g547)) + ((!g376) & (g377) & (g387) & (!g388) & (g412) & (!g547)) + ((!g376) & (g377) & (g387) & (!g388) & (g412) & (g547)) + ((!g376) & (g377) & (g387) & (g388) & (!g412) & (!g547)) + ((!g376) & (g377) & (g387) & (g388) & (!g412) & (g547)) + ((!g376) & (g377) & (g387) & (g388) & (g412) & (!g547)) + ((!g376) & (g377) & (g387) & (g388) & (g412) & (g547)) + ((g376) & (g377) & (!g387) & (!g388) & (!g412) & (!g547)) + ((g376) & (g377) & (!g387) & (!g388) & (!g412) & (g547)) + ((g376) & (g377) & (!g387) & (!g388) & (g412) & (!g547)) + ((g376) & (g377) & (!g387) & (!g388) & (g412) & (g547)) + ((g376) & (g377) & (!g387) & (g388) & (!g412) & (!g547)) + ((g376) & (g377) & (g387) & (!g388) & (!g412) & (!g547)));
	assign g549 = (((!sk[47]) & (!g316) & (g322) & (!g548)) + ((!sk[47]) & (!g316) & (g322) & (g548)) + ((!sk[47]) & (g316) & (g322) & (!g548)) + ((!sk[47]) & (g316) & (g322) & (g548)) + ((sk[47]) & (!g316) & (!g322) & (g548)) + ((sk[47]) & (!g316) & (g322) & (!g548)) + ((sk[47]) & (g316) & (!g322) & (!g548)) + ((sk[47]) & (g316) & (g322) & (g548)));
	assign g550 = (((!g50) & (!sk[48]) & (g29) & (!g31)) + ((!g50) & (!sk[48]) & (g29) & (g31)) + ((!g50) & (sk[48]) & (!g29) & (!g31)) + ((g50) & (!sk[48]) & (g29) & (!g31)) + ((g50) & (!sk[48]) & (g29) & (g31)));
	assign g551 = (((!sk[49]) & (g49) & (g71)) + ((sk[49]) & (g49) & (g71)));
	assign g552 = (((!g38) & (!g99) & (!g62) & (!sk[50]) & (g74) & (!g551)) + ((!g38) & (!g99) & (!g62) & (!sk[50]) & (g74) & (g551)) + ((!g38) & (!g99) & (!g62) & (sk[50]) & (!g74) & (!g551)) + ((!g38) & (!g99) & (g62) & (!sk[50]) & (!g74) & (!g551)) + ((!g38) & (!g99) & (g62) & (!sk[50]) & (!g74) & (g551)) + ((!g38) & (!g99) & (g62) & (!sk[50]) & (g74) & (!g551)) + ((!g38) & (!g99) & (g62) & (!sk[50]) & (g74) & (g551)) + ((!g38) & (!g99) & (g62) & (sk[50]) & (!g74) & (!g551)) + ((!g38) & (g99) & (!g62) & (!sk[50]) & (!g74) & (!g551)) + ((!g38) & (g99) & (!g62) & (!sk[50]) & (!g74) & (g551)) + ((!g38) & (g99) & (!g62) & (!sk[50]) & (g74) & (!g551)) + ((!g38) & (g99) & (!g62) & (!sk[50]) & (g74) & (g551)) + ((!g38) & (g99) & (!g62) & (sk[50]) & (!g74) & (!g551)) + ((!g38) & (g99) & (g62) & (!sk[50]) & (!g74) & (!g551)) + ((!g38) & (g99) & (g62) & (!sk[50]) & (!g74) & (g551)) + ((!g38) & (g99) & (g62) & (!sk[50]) & (g74) & (!g551)) + ((!g38) & (g99) & (g62) & (!sk[50]) & (g74) & (g551)) + ((!g38) & (g99) & (g62) & (sk[50]) & (!g74) & (!g551)) + ((g38) & (!g99) & (!g62) & (!sk[50]) & (g74) & (!g551)) + ((g38) & (!g99) & (!g62) & (!sk[50]) & (g74) & (g551)) + ((g38) & (!g99) & (!g62) & (sk[50]) & (!g74) & (!g551)) + ((g38) & (!g99) & (g62) & (!sk[50]) & (!g74) & (!g551)) + ((g38) & (!g99) & (g62) & (!sk[50]) & (!g74) & (g551)) + ((g38) & (!g99) & (g62) & (!sk[50]) & (g74) & (!g551)) + ((g38) & (!g99) & (g62) & (!sk[50]) & (g74) & (g551)) + ((g38) & (g99) & (!g62) & (!sk[50]) & (!g74) & (!g551)) + ((g38) & (g99) & (!g62) & (!sk[50]) & (!g74) & (g551)) + ((g38) & (g99) & (!g62) & (!sk[50]) & (g74) & (!g551)) + ((g38) & (g99) & (!g62) & (!sk[50]) & (g74) & (g551)) + ((g38) & (g99) & (g62) & (!sk[50]) & (!g74) & (!g551)) + ((g38) & (g99) & (g62) & (!sk[50]) & (!g74) & (g551)) + ((g38) & (g99) & (g62) & (!sk[50]) & (g74) & (!g551)) + ((g38) & (g99) & (g62) & (!sk[50]) & (g74) & (g551)));
	assign g553 = (((!g9) & (!sk[51]) & (g66) & (!g43)) + ((!g9) & (!sk[51]) & (g66) & (g43)) + ((!g9) & (sk[51]) & (!g66) & (!g43)) + ((!g9) & (sk[51]) & (g66) & (!g43)) + ((g9) & (!sk[51]) & (g66) & (!g43)) + ((g9) & (!sk[51]) & (g66) & (g43)) + ((g9) & (sk[51]) & (!g66) & (!g43)));
	assign g554 = (((!g16) & (!sk[52]) & (!g12) & (!g42) & (g84) & (!g187)) + ((!g16) & (!sk[52]) & (!g12) & (!g42) & (g84) & (g187)) + ((!g16) & (!sk[52]) & (!g12) & (g42) & (!g84) & (!g187)) + ((!g16) & (!sk[52]) & (!g12) & (g42) & (!g84) & (g187)) + ((!g16) & (!sk[52]) & (!g12) & (g42) & (g84) & (!g187)) + ((!g16) & (!sk[52]) & (!g12) & (g42) & (g84) & (g187)) + ((!g16) & (!sk[52]) & (g12) & (!g42) & (!g84) & (!g187)) + ((!g16) & (!sk[52]) & (g12) & (!g42) & (!g84) & (g187)) + ((!g16) & (!sk[52]) & (g12) & (!g42) & (g84) & (!g187)) + ((!g16) & (!sk[52]) & (g12) & (!g42) & (g84) & (g187)) + ((!g16) & (!sk[52]) & (g12) & (g42) & (!g84) & (!g187)) + ((!g16) & (!sk[52]) & (g12) & (g42) & (!g84) & (g187)) + ((!g16) & (!sk[52]) & (g12) & (g42) & (g84) & (!g187)) + ((!g16) & (!sk[52]) & (g12) & (g42) & (g84) & (g187)) + ((!g16) & (sk[52]) & (!g12) & (!g42) & (!g84) & (!g187)) + ((!g16) & (sk[52]) & (!g12) & (g42) & (!g84) & (!g187)) + ((!g16) & (sk[52]) & (g12) & (!g42) & (!g84) & (!g187)) + ((!g16) & (sk[52]) & (g12) & (g42) & (!g84) & (!g187)) + ((g16) & (!sk[52]) & (!g12) & (!g42) & (g84) & (!g187)) + ((g16) & (!sk[52]) & (!g12) & (!g42) & (g84) & (g187)) + ((g16) & (!sk[52]) & (!g12) & (g42) & (!g84) & (!g187)) + ((g16) & (!sk[52]) & (!g12) & (g42) & (!g84) & (g187)) + ((g16) & (!sk[52]) & (!g12) & (g42) & (g84) & (!g187)) + ((g16) & (!sk[52]) & (!g12) & (g42) & (g84) & (g187)) + ((g16) & (!sk[52]) & (g12) & (!g42) & (!g84) & (!g187)) + ((g16) & (!sk[52]) & (g12) & (!g42) & (!g84) & (g187)) + ((g16) & (!sk[52]) & (g12) & (!g42) & (g84) & (!g187)) + ((g16) & (!sk[52]) & (g12) & (!g42) & (g84) & (g187)) + ((g16) & (!sk[52]) & (g12) & (g42) & (!g84) & (!g187)) + ((g16) & (!sk[52]) & (g12) & (g42) & (!g84) & (g187)) + ((g16) & (!sk[52]) & (g12) & (g42) & (g84) & (!g187)) + ((g16) & (!sk[52]) & (g12) & (g42) & (g84) & (g187)) + ((g16) & (sk[52]) & (!g12) & (!g42) & (!g84) & (!g187)));
	assign g555 = (((!sk[53]) & (!g70) & (!g105) & (!g20) & (g141)) + ((!sk[53]) & (!g70) & (!g105) & (g20) & (g141)) + ((!sk[53]) & (!g70) & (g105) & (!g20) & (g141)) + ((!sk[53]) & (!g70) & (g105) & (g20) & (g141)) + ((!sk[53]) & (g70) & (!g105) & (!g20) & (!g141)) + ((!sk[53]) & (g70) & (!g105) & (!g20) & (g141)) + ((!sk[53]) & (g70) & (!g105) & (g20) & (!g141)) + ((!sk[53]) & (g70) & (!g105) & (g20) & (g141)) + ((!sk[53]) & (g70) & (g105) & (!g20) & (!g141)) + ((!sk[53]) & (g70) & (g105) & (!g20) & (g141)) + ((!sk[53]) & (g70) & (g105) & (g20) & (!g141)) + ((!sk[53]) & (g70) & (g105) & (g20) & (g141)) + ((sk[53]) & (!g70) & (!g105) & (!g20) & (!g141)) + ((sk[53]) & (!g70) & (!g105) & (g20) & (!g141)) + ((sk[53]) & (g70) & (!g105) & (!g20) & (!g141)));
	assign g556 = (((!g49) & (!g46) & (!g553) & (g554) & (!sk[54]) & (!g555)) + ((!g49) & (!g46) & (!g553) & (g554) & (!sk[54]) & (g555)) + ((!g49) & (!g46) & (g553) & (!g554) & (!sk[54]) & (!g555)) + ((!g49) & (!g46) & (g553) & (!g554) & (!sk[54]) & (g555)) + ((!g49) & (!g46) & (g553) & (g554) & (!sk[54]) & (!g555)) + ((!g49) & (!g46) & (g553) & (g554) & (!sk[54]) & (g555)) + ((!g49) & (!g46) & (g553) & (g554) & (sk[54]) & (g555)) + ((!g49) & (g46) & (!g553) & (!g554) & (!sk[54]) & (!g555)) + ((!g49) & (g46) & (!g553) & (!g554) & (!sk[54]) & (g555)) + ((!g49) & (g46) & (!g553) & (g554) & (!sk[54]) & (!g555)) + ((!g49) & (g46) & (!g553) & (g554) & (!sk[54]) & (g555)) + ((!g49) & (g46) & (g553) & (!g554) & (!sk[54]) & (!g555)) + ((!g49) & (g46) & (g553) & (!g554) & (!sk[54]) & (g555)) + ((!g49) & (g46) & (g553) & (g554) & (!sk[54]) & (!g555)) + ((!g49) & (g46) & (g553) & (g554) & (!sk[54]) & (g555)) + ((!g49) & (g46) & (g553) & (g554) & (sk[54]) & (g555)) + ((g49) & (!g46) & (!g553) & (g554) & (!sk[54]) & (!g555)) + ((g49) & (!g46) & (!g553) & (g554) & (!sk[54]) & (g555)) + ((g49) & (!g46) & (g553) & (!g554) & (!sk[54]) & (!g555)) + ((g49) & (!g46) & (g553) & (!g554) & (!sk[54]) & (g555)) + ((g49) & (!g46) & (g553) & (g554) & (!sk[54]) & (!g555)) + ((g49) & (!g46) & (g553) & (g554) & (!sk[54]) & (g555)) + ((g49) & (!g46) & (g553) & (g554) & (sk[54]) & (g555)) + ((g49) & (g46) & (!g553) & (!g554) & (!sk[54]) & (!g555)) + ((g49) & (g46) & (!g553) & (!g554) & (!sk[54]) & (g555)) + ((g49) & (g46) & (!g553) & (g554) & (!sk[54]) & (!g555)) + ((g49) & (g46) & (!g553) & (g554) & (!sk[54]) & (g555)) + ((g49) & (g46) & (g553) & (!g554) & (!sk[54]) & (!g555)) + ((g49) & (g46) & (g553) & (!g554) & (!sk[54]) & (g555)) + ((g49) & (g46) & (g553) & (g554) & (!sk[54]) & (!g555)) + ((g49) & (g46) & (g553) & (g554) & (!sk[54]) & (g555)));
	assign g557 = (((!g550) & (!g552) & (!sk[55]) & (!g294) & (g246) & (!g556)) + ((!g550) & (!g552) & (!sk[55]) & (!g294) & (g246) & (g556)) + ((!g550) & (!g552) & (!sk[55]) & (g294) & (!g246) & (!g556)) + ((!g550) & (!g552) & (!sk[55]) & (g294) & (!g246) & (g556)) + ((!g550) & (!g552) & (!sk[55]) & (g294) & (g246) & (!g556)) + ((!g550) & (!g552) & (!sk[55]) & (g294) & (g246) & (g556)) + ((!g550) & (g552) & (!sk[55]) & (!g294) & (!g246) & (!g556)) + ((!g550) & (g552) & (!sk[55]) & (!g294) & (!g246) & (g556)) + ((!g550) & (g552) & (!sk[55]) & (!g294) & (g246) & (!g556)) + ((!g550) & (g552) & (!sk[55]) & (!g294) & (g246) & (g556)) + ((!g550) & (g552) & (!sk[55]) & (g294) & (!g246) & (!g556)) + ((!g550) & (g552) & (!sk[55]) & (g294) & (!g246) & (g556)) + ((!g550) & (g552) & (!sk[55]) & (g294) & (g246) & (!g556)) + ((!g550) & (g552) & (!sk[55]) & (g294) & (g246) & (g556)) + ((g550) & (!g552) & (!sk[55]) & (!g294) & (g246) & (!g556)) + ((g550) & (!g552) & (!sk[55]) & (!g294) & (g246) & (g556)) + ((g550) & (!g552) & (!sk[55]) & (g294) & (!g246) & (!g556)) + ((g550) & (!g552) & (!sk[55]) & (g294) & (!g246) & (g556)) + ((g550) & (!g552) & (!sk[55]) & (g294) & (g246) & (!g556)) + ((g550) & (!g552) & (!sk[55]) & (g294) & (g246) & (g556)) + ((g550) & (g552) & (!sk[55]) & (!g294) & (!g246) & (!g556)) + ((g550) & (g552) & (!sk[55]) & (!g294) & (!g246) & (g556)) + ((g550) & (g552) & (!sk[55]) & (!g294) & (g246) & (!g556)) + ((g550) & (g552) & (!sk[55]) & (!g294) & (g246) & (g556)) + ((g550) & (g552) & (!sk[55]) & (g294) & (!g246) & (!g556)) + ((g550) & (g552) & (!sk[55]) & (g294) & (!g246) & (g556)) + ((g550) & (g552) & (!sk[55]) & (g294) & (g246) & (!g556)) + ((g550) & (g552) & (!sk[55]) & (g294) & (g246) & (g556)) + ((g550) & (g552) & (sk[55]) & (g294) & (g246) & (g556)));
	assign g558 = (((!g17) & (!g62) & (!g58) & (!g27) & (!g11) & (g557)) + ((!g17) & (!g62) & (!g58) & (g27) & (!g11) & (g557)) + ((!g17) & (!g62) & (g58) & (!g27) & (!g11) & (g557)) + ((!g17) & (!g62) & (g58) & (g27) & (!g11) & (g557)) + ((!g17) & (g62) & (!g58) & (!g27) & (!g11) & (g557)) + ((g17) & (!g62) & (!g58) & (!g27) & (!g11) & (g557)) + ((g17) & (!g62) & (!g58) & (g27) & (!g11) & (g557)) + ((g17) & (!g62) & (g58) & (!g27) & (!g11) & (g557)) + ((g17) & (!g62) & (g58) & (g27) & (!g11) & (g557)));
	assign g559 = (((!g78) & (!g71) & (!g58) & (!g46) & (!g41) & (g176)) + ((!g78) & (!g71) & (!g58) & (!g46) & (g41) & (g176)) + ((!g78) & (!g71) & (!g58) & (g46) & (!g41) & (g176)) + ((!g78) & (!g71) & (g58) & (!g46) & (!g41) & (g176)) + ((!g78) & (!g71) & (g58) & (!g46) & (g41) & (g176)) + ((!g78) & (!g71) & (g58) & (g46) & (!g41) & (g176)) + ((!g78) & (g71) & (!g58) & (!g46) & (!g41) & (g176)) + ((!g78) & (g71) & (!g58) & (!g46) & (g41) & (g176)) + ((!g78) & (g71) & (!g58) & (g46) & (!g41) & (g176)));
	assign g560 = (((!g19) & (!sk[58]) & (g36) & (!g242)) + ((!g19) & (!sk[58]) & (g36) & (g242)) + ((!g19) & (sk[58]) & (!g36) & (g242)) + ((g19) & (!sk[58]) & (g36) & (!g242)) + ((g19) & (!sk[58]) & (g36) & (g242)));
	assign g561 = (((!g163) & (!g99) & (!sk[59]) & (!g12) & (g59) & (!g64)) + ((!g163) & (!g99) & (!sk[59]) & (!g12) & (g59) & (g64)) + ((!g163) & (!g99) & (!sk[59]) & (g12) & (!g59) & (!g64)) + ((!g163) & (!g99) & (!sk[59]) & (g12) & (!g59) & (g64)) + ((!g163) & (!g99) & (!sk[59]) & (g12) & (g59) & (!g64)) + ((!g163) & (!g99) & (!sk[59]) & (g12) & (g59) & (g64)) + ((!g163) & (!g99) & (sk[59]) & (!g12) & (!g59) & (!g64)) + ((!g163) & (!g99) & (sk[59]) & (g12) & (!g59) & (!g64)) + ((!g163) & (g99) & (!sk[59]) & (!g12) & (!g59) & (!g64)) + ((!g163) & (g99) & (!sk[59]) & (!g12) & (!g59) & (g64)) + ((!g163) & (g99) & (!sk[59]) & (!g12) & (g59) & (!g64)) + ((!g163) & (g99) & (!sk[59]) & (!g12) & (g59) & (g64)) + ((!g163) & (g99) & (!sk[59]) & (g12) & (!g59) & (!g64)) + ((!g163) & (g99) & (!sk[59]) & (g12) & (!g59) & (g64)) + ((!g163) & (g99) & (!sk[59]) & (g12) & (g59) & (!g64)) + ((!g163) & (g99) & (!sk[59]) & (g12) & (g59) & (g64)) + ((!g163) & (g99) & (sk[59]) & (!g12) & (!g59) & (!g64)) + ((g163) & (!g99) & (!sk[59]) & (!g12) & (g59) & (!g64)) + ((g163) & (!g99) & (!sk[59]) & (!g12) & (g59) & (g64)) + ((g163) & (!g99) & (!sk[59]) & (g12) & (!g59) & (!g64)) + ((g163) & (!g99) & (!sk[59]) & (g12) & (!g59) & (g64)) + ((g163) & (!g99) & (!sk[59]) & (g12) & (g59) & (!g64)) + ((g163) & (!g99) & (!sk[59]) & (g12) & (g59) & (g64)) + ((g163) & (g99) & (!sk[59]) & (!g12) & (!g59) & (!g64)) + ((g163) & (g99) & (!sk[59]) & (!g12) & (!g59) & (g64)) + ((g163) & (g99) & (!sk[59]) & (!g12) & (g59) & (!g64)) + ((g163) & (g99) & (!sk[59]) & (!g12) & (g59) & (g64)) + ((g163) & (g99) & (!sk[59]) & (g12) & (!g59) & (!g64)) + ((g163) & (g99) & (!sk[59]) & (g12) & (!g59) & (g64)) + ((g163) & (g99) & (!sk[59]) & (g12) & (g59) & (!g64)) + ((g163) & (g99) & (!sk[59]) & (g12) & (g59) & (g64)));
	assign g562 = (((!g101) & (!sk[60]) & (!g290) & (!g559) & (g560) & (!g561)) + ((!g101) & (!sk[60]) & (!g290) & (!g559) & (g560) & (g561)) + ((!g101) & (!sk[60]) & (!g290) & (g559) & (!g560) & (!g561)) + ((!g101) & (!sk[60]) & (!g290) & (g559) & (!g560) & (g561)) + ((!g101) & (!sk[60]) & (!g290) & (g559) & (g560) & (!g561)) + ((!g101) & (!sk[60]) & (!g290) & (g559) & (g560) & (g561)) + ((!g101) & (!sk[60]) & (g290) & (!g559) & (!g560) & (!g561)) + ((!g101) & (!sk[60]) & (g290) & (!g559) & (!g560) & (g561)) + ((!g101) & (!sk[60]) & (g290) & (!g559) & (g560) & (!g561)) + ((!g101) & (!sk[60]) & (g290) & (!g559) & (g560) & (g561)) + ((!g101) & (!sk[60]) & (g290) & (g559) & (!g560) & (!g561)) + ((!g101) & (!sk[60]) & (g290) & (g559) & (!g560) & (g561)) + ((!g101) & (!sk[60]) & (g290) & (g559) & (g560) & (!g561)) + ((!g101) & (!sk[60]) & (g290) & (g559) & (g560) & (g561)) + ((!g101) & (sk[60]) & (g290) & (g559) & (g560) & (g561)) + ((g101) & (!sk[60]) & (!g290) & (!g559) & (g560) & (!g561)) + ((g101) & (!sk[60]) & (!g290) & (!g559) & (g560) & (g561)) + ((g101) & (!sk[60]) & (!g290) & (g559) & (!g560) & (!g561)) + ((g101) & (!sk[60]) & (!g290) & (g559) & (!g560) & (g561)) + ((g101) & (!sk[60]) & (!g290) & (g559) & (g560) & (!g561)) + ((g101) & (!sk[60]) & (!g290) & (g559) & (g560) & (g561)) + ((g101) & (!sk[60]) & (g290) & (!g559) & (!g560) & (!g561)) + ((g101) & (!sk[60]) & (g290) & (!g559) & (!g560) & (g561)) + ((g101) & (!sk[60]) & (g290) & (!g559) & (g560) & (!g561)) + ((g101) & (!sk[60]) & (g290) & (!g559) & (g560) & (g561)) + ((g101) & (!sk[60]) & (g290) & (g559) & (!g560) & (!g561)) + ((g101) & (!sk[60]) & (g290) & (g559) & (!g560) & (g561)) + ((g101) & (!sk[60]) & (g290) & (g559) & (g560) & (!g561)) + ((g101) & (!sk[60]) & (g290) & (g559) & (g560) & (g561)));
	assign g563 = (((!sk[61]) & (!g38) & (!g70) & (!g16) & (g17)) + ((!sk[61]) & (!g38) & (!g70) & (g16) & (g17)) + ((!sk[61]) & (!g38) & (g70) & (!g16) & (g17)) + ((!sk[61]) & (!g38) & (g70) & (g16) & (g17)) + ((!sk[61]) & (g38) & (!g70) & (!g16) & (!g17)) + ((!sk[61]) & (g38) & (!g70) & (!g16) & (g17)) + ((!sk[61]) & (g38) & (!g70) & (g16) & (!g17)) + ((!sk[61]) & (g38) & (!g70) & (g16) & (g17)) + ((!sk[61]) & (g38) & (g70) & (!g16) & (!g17)) + ((!sk[61]) & (g38) & (g70) & (!g16) & (g17)) + ((!sk[61]) & (g38) & (g70) & (g16) & (!g17)) + ((!sk[61]) & (g38) & (g70) & (g16) & (g17)) + ((sk[61]) & (!g38) & (g70) & (!g16) & (g17)) + ((sk[61]) & (!g38) & (g70) & (g16) & (g17)) + ((sk[61]) & (g38) & (!g70) & (g16) & (!g17)) + ((sk[61]) & (g38) & (!g70) & (g16) & (g17)) + ((sk[61]) & (g38) & (g70) & (!g16) & (g17)) + ((sk[61]) & (g38) & (g70) & (g16) & (!g17)) + ((sk[61]) & (g38) & (g70) & (g16) & (g17)));
	assign g564 = (((!sk[62]) & (!g9) & (!g62) & (!g18) & (g25)) + ((!sk[62]) & (!g9) & (!g62) & (g18) & (g25)) + ((!sk[62]) & (!g9) & (g62) & (!g18) & (g25)) + ((!sk[62]) & (!g9) & (g62) & (g18) & (g25)) + ((!sk[62]) & (g9) & (!g62) & (!g18) & (!g25)) + ((!sk[62]) & (g9) & (!g62) & (!g18) & (g25)) + ((!sk[62]) & (g9) & (!g62) & (g18) & (!g25)) + ((!sk[62]) & (g9) & (!g62) & (g18) & (g25)) + ((!sk[62]) & (g9) & (g62) & (!g18) & (!g25)) + ((!sk[62]) & (g9) & (g62) & (!g18) & (g25)) + ((!sk[62]) & (g9) & (g62) & (g18) & (!g25)) + ((!sk[62]) & (g9) & (g62) & (g18) & (g25)) + ((sk[62]) & (!g9) & (g62) & (g18) & (!g25)) + ((sk[62]) & (!g9) & (g62) & (g18) & (g25)) + ((sk[62]) & (g9) & (!g62) & (!g18) & (g25)) + ((sk[62]) & (g9) & (!g62) & (g18) & (g25)) + ((sk[62]) & (g9) & (g62) & (!g18) & (g25)) + ((sk[62]) & (g9) & (g62) & (g18) & (!g25)) + ((sk[62]) & (g9) & (g62) & (g18) & (g25)));
	assign g565 = (((!sk[63]) & (!g16) & (!g563) & (!g66) & (g152) & (!g564)) + ((!sk[63]) & (!g16) & (!g563) & (!g66) & (g152) & (g564)) + ((!sk[63]) & (!g16) & (!g563) & (g66) & (!g152) & (!g564)) + ((!sk[63]) & (!g16) & (!g563) & (g66) & (!g152) & (g564)) + ((!sk[63]) & (!g16) & (!g563) & (g66) & (g152) & (!g564)) + ((!sk[63]) & (!g16) & (!g563) & (g66) & (g152) & (g564)) + ((!sk[63]) & (!g16) & (g563) & (!g66) & (!g152) & (!g564)) + ((!sk[63]) & (!g16) & (g563) & (!g66) & (!g152) & (g564)) + ((!sk[63]) & (!g16) & (g563) & (!g66) & (g152) & (!g564)) + ((!sk[63]) & (!g16) & (g563) & (!g66) & (g152) & (g564)) + ((!sk[63]) & (!g16) & (g563) & (g66) & (!g152) & (!g564)) + ((!sk[63]) & (!g16) & (g563) & (g66) & (!g152) & (g564)) + ((!sk[63]) & (!g16) & (g563) & (g66) & (g152) & (!g564)) + ((!sk[63]) & (!g16) & (g563) & (g66) & (g152) & (g564)) + ((!sk[63]) & (g16) & (!g563) & (!g66) & (g152) & (!g564)) + ((!sk[63]) & (g16) & (!g563) & (!g66) & (g152) & (g564)) + ((!sk[63]) & (g16) & (!g563) & (g66) & (!g152) & (!g564)) + ((!sk[63]) & (g16) & (!g563) & (g66) & (!g152) & (g564)) + ((!sk[63]) & (g16) & (!g563) & (g66) & (g152) & (!g564)) + ((!sk[63]) & (g16) & (!g563) & (g66) & (g152) & (g564)) + ((!sk[63]) & (g16) & (g563) & (!g66) & (!g152) & (!g564)) + ((!sk[63]) & (g16) & (g563) & (!g66) & (!g152) & (g564)) + ((!sk[63]) & (g16) & (g563) & (!g66) & (g152) & (!g564)) + ((!sk[63]) & (g16) & (g563) & (!g66) & (g152) & (g564)) + ((!sk[63]) & (g16) & (g563) & (g66) & (!g152) & (!g564)) + ((!sk[63]) & (g16) & (g563) & (g66) & (!g152) & (g564)) + ((!sk[63]) & (g16) & (g563) & (g66) & (g152) & (!g564)) + ((!sk[63]) & (g16) & (g563) & (g66) & (g152) & (g564)) + ((sk[63]) & (!g16) & (!g563) & (!g66) & (!g152) & (!g564)) + ((sk[63]) & (!g16) & (!g563) & (g66) & (!g152) & (!g564)) + ((sk[63]) & (g16) & (!g563) & (!g66) & (!g152) & (!g564)));
	assign g566 = (((!g10) & (!g99) & (!sk[64]) & (!g104) & (g25) & (!g85)) + ((!g10) & (!g99) & (!sk[64]) & (!g104) & (g25) & (g85)) + ((!g10) & (!g99) & (!sk[64]) & (g104) & (!g25) & (!g85)) + ((!g10) & (!g99) & (!sk[64]) & (g104) & (!g25) & (g85)) + ((!g10) & (!g99) & (!sk[64]) & (g104) & (g25) & (!g85)) + ((!g10) & (!g99) & (!sk[64]) & (g104) & (g25) & (g85)) + ((!g10) & (!g99) & (sk[64]) & (!g104) & (!g25) & (!g85)) + ((!g10) & (!g99) & (sk[64]) & (!g104) & (g25) & (!g85)) + ((!g10) & (!g99) & (sk[64]) & (g104) & (!g25) & (!g85)) + ((!g10) & (g99) & (!sk[64]) & (!g104) & (!g25) & (!g85)) + ((!g10) & (g99) & (!sk[64]) & (!g104) & (!g25) & (g85)) + ((!g10) & (g99) & (!sk[64]) & (!g104) & (g25) & (!g85)) + ((!g10) & (g99) & (!sk[64]) & (!g104) & (g25) & (g85)) + ((!g10) & (g99) & (!sk[64]) & (g104) & (!g25) & (!g85)) + ((!g10) & (g99) & (!sk[64]) & (g104) & (!g25) & (g85)) + ((!g10) & (g99) & (!sk[64]) & (g104) & (g25) & (!g85)) + ((!g10) & (g99) & (!sk[64]) & (g104) & (g25) & (g85)) + ((!g10) & (g99) & (sk[64]) & (!g104) & (!g25) & (!g85)) + ((!g10) & (g99) & (sk[64]) & (!g104) & (g25) & (!g85)) + ((!g10) & (g99) & (sk[64]) & (g104) & (!g25) & (!g85)) + ((g10) & (!g99) & (!sk[64]) & (!g104) & (g25) & (!g85)) + ((g10) & (!g99) & (!sk[64]) & (!g104) & (g25) & (g85)) + ((g10) & (!g99) & (!sk[64]) & (g104) & (!g25) & (!g85)) + ((g10) & (!g99) & (!sk[64]) & (g104) & (!g25) & (g85)) + ((g10) & (!g99) & (!sk[64]) & (g104) & (g25) & (!g85)) + ((g10) & (!g99) & (!sk[64]) & (g104) & (g25) & (g85)) + ((g10) & (!g99) & (sk[64]) & (!g104) & (!g25) & (!g85)) + ((g10) & (!g99) & (sk[64]) & (!g104) & (g25) & (!g85)) + ((g10) & (g99) & (!sk[64]) & (!g104) & (!g25) & (!g85)) + ((g10) & (g99) & (!sk[64]) & (!g104) & (!g25) & (g85)) + ((g10) & (g99) & (!sk[64]) & (!g104) & (g25) & (!g85)) + ((g10) & (g99) & (!sk[64]) & (!g104) & (g25) & (g85)) + ((g10) & (g99) & (!sk[64]) & (g104) & (!g25) & (!g85)) + ((g10) & (g99) & (!sk[64]) & (g104) & (!g25) & (g85)) + ((g10) & (g99) & (!sk[64]) & (g104) & (g25) & (!g85)) + ((g10) & (g99) & (!sk[64]) & (g104) & (g25) & (g85)));
	assign g567 = (((!g46) & (!sk[65]) & (!g40) & (!g275) & (g566)) + ((!g46) & (!sk[65]) & (!g40) & (g275) & (g566)) + ((!g46) & (!sk[65]) & (g40) & (!g275) & (g566)) + ((!g46) & (!sk[65]) & (g40) & (g275) & (g566)) + ((!g46) & (sk[65]) & (!g40) & (!g275) & (g566)) + ((!g46) & (sk[65]) & (g40) & (!g275) & (g566)) + ((g46) & (!sk[65]) & (!g40) & (!g275) & (!g566)) + ((g46) & (!sk[65]) & (!g40) & (!g275) & (g566)) + ((g46) & (!sk[65]) & (!g40) & (g275) & (!g566)) + ((g46) & (!sk[65]) & (!g40) & (g275) & (g566)) + ((g46) & (!sk[65]) & (g40) & (!g275) & (!g566)) + ((g46) & (!sk[65]) & (g40) & (!g275) & (g566)) + ((g46) & (!sk[65]) & (g40) & (g275) & (!g566)) + ((g46) & (!sk[65]) & (g40) & (g275) & (g566)) + ((g46) & (sk[65]) & (!g40) & (!g275) & (g566)));
	assign g568 = (((!g55) & (!g73) & (sk[66]) & (!g211)) + ((!g55) & (g73) & (!sk[66]) & (!g211)) + ((!g55) & (g73) & (!sk[66]) & (g211)) + ((g55) & (g73) & (!sk[66]) & (!g211)) + ((g55) & (g73) & (!sk[66]) & (g211)));
	assign g569 = (((!g558) & (!g562) & (!sk[67]) & (!g565) & (g567) & (!g568)) + ((!g558) & (!g562) & (!sk[67]) & (!g565) & (g567) & (g568)) + ((!g558) & (!g562) & (!sk[67]) & (g565) & (!g567) & (!g568)) + ((!g558) & (!g562) & (!sk[67]) & (g565) & (!g567) & (g568)) + ((!g558) & (!g562) & (!sk[67]) & (g565) & (g567) & (!g568)) + ((!g558) & (!g562) & (!sk[67]) & (g565) & (g567) & (g568)) + ((!g558) & (g562) & (!sk[67]) & (!g565) & (!g567) & (!g568)) + ((!g558) & (g562) & (!sk[67]) & (!g565) & (!g567) & (g568)) + ((!g558) & (g562) & (!sk[67]) & (!g565) & (g567) & (!g568)) + ((!g558) & (g562) & (!sk[67]) & (!g565) & (g567) & (g568)) + ((!g558) & (g562) & (!sk[67]) & (g565) & (!g567) & (!g568)) + ((!g558) & (g562) & (!sk[67]) & (g565) & (!g567) & (g568)) + ((!g558) & (g562) & (!sk[67]) & (g565) & (g567) & (!g568)) + ((!g558) & (g562) & (!sk[67]) & (g565) & (g567) & (g568)) + ((g558) & (!g562) & (!sk[67]) & (!g565) & (g567) & (!g568)) + ((g558) & (!g562) & (!sk[67]) & (!g565) & (g567) & (g568)) + ((g558) & (!g562) & (!sk[67]) & (g565) & (!g567) & (!g568)) + ((g558) & (!g562) & (!sk[67]) & (g565) & (!g567) & (g568)) + ((g558) & (!g562) & (!sk[67]) & (g565) & (g567) & (!g568)) + ((g558) & (!g562) & (!sk[67]) & (g565) & (g567) & (g568)) + ((g558) & (g562) & (!sk[67]) & (!g565) & (!g567) & (!g568)) + ((g558) & (g562) & (!sk[67]) & (!g565) & (!g567) & (g568)) + ((g558) & (g562) & (!sk[67]) & (!g565) & (g567) & (!g568)) + ((g558) & (g562) & (!sk[67]) & (!g565) & (g567) & (g568)) + ((g558) & (g562) & (!sk[67]) & (g565) & (!g567) & (!g568)) + ((g558) & (g562) & (!sk[67]) & (g565) & (!g567) & (g568)) + ((g558) & (g562) & (!sk[67]) & (g565) & (g567) & (!g568)) + ((g558) & (g562) & (!sk[67]) & (g565) & (g567) & (g568)) + ((g558) & (g562) & (sk[67]) & (g565) & (g567) & (g568)));
	assign g570 = (((!g376) & (sk[68]) & (g377)) + ((g376) & (!sk[68]) & (g377)) + ((g376) & (sk[68]) & (!g377)));
	assign g571 = (((!g387) & (!g388) & (!g412) & (!sk[69]) & (g547)) + ((!g387) & (!g388) & (!g412) & (sk[69]) & (!g547)) + ((!g387) & (!g388) & (!g412) & (sk[69]) & (g547)) + ((!g387) & (!g388) & (g412) & (!sk[69]) & (g547)) + ((!g387) & (!g388) & (g412) & (sk[69]) & (!g547)) + ((!g387) & (!g388) & (g412) & (sk[69]) & (g547)) + ((!g387) & (g388) & (!g412) & (!sk[69]) & (g547)) + ((!g387) & (g388) & (!g412) & (sk[69]) & (!g547)) + ((!g387) & (g388) & (g412) & (!sk[69]) & (g547)) + ((g387) & (!g388) & (!g412) & (!sk[69]) & (!g547)) + ((g387) & (!g388) & (!g412) & (!sk[69]) & (g547)) + ((g387) & (!g388) & (!g412) & (sk[69]) & (!g547)) + ((g387) & (!g388) & (g412) & (!sk[69]) & (!g547)) + ((g387) & (!g388) & (g412) & (!sk[69]) & (g547)) + ((g387) & (g388) & (!g412) & (!sk[69]) & (!g547)) + ((g387) & (g388) & (!g412) & (!sk[69]) & (g547)) + ((g387) & (g388) & (g412) & (!sk[69]) & (!g547)) + ((g387) & (g388) & (g412) & (!sk[69]) & (g547)));
	assign g572 = (((!sk[70]) & (g62) & (g41)) + ((sk[70]) & (g62) & (g41)));
	assign g573 = (((!g9) & (!g10) & (!sk[71]) & (!g17) & (g99)) + ((!g9) & (!g10) & (!sk[71]) & (g17) & (g99)) + ((!g9) & (!g10) & (sk[71]) & (g17) & (g99)) + ((!g9) & (g10) & (!sk[71]) & (!g17) & (g99)) + ((!g9) & (g10) & (!sk[71]) & (g17) & (g99)) + ((!g9) & (g10) & (sk[71]) & (g17) & (g99)) + ((g9) & (!g10) & (!sk[71]) & (!g17) & (!g99)) + ((g9) & (!g10) & (!sk[71]) & (!g17) & (g99)) + ((g9) & (!g10) & (!sk[71]) & (g17) & (!g99)) + ((g9) & (!g10) & (!sk[71]) & (g17) & (g99)) + ((g9) & (!g10) & (sk[71]) & (g17) & (g99)) + ((g9) & (g10) & (!sk[71]) & (!g17) & (!g99)) + ((g9) & (g10) & (!sk[71]) & (!g17) & (g99)) + ((g9) & (g10) & (!sk[71]) & (g17) & (!g99)) + ((g9) & (g10) & (!sk[71]) & (g17) & (g99)) + ((g9) & (g10) & (sk[71]) & (!g17) & (!g99)) + ((g9) & (g10) & (sk[71]) & (!g17) & (g99)) + ((g9) & (g10) & (sk[71]) & (g17) & (!g99)) + ((g9) & (g10) & (sk[71]) & (g17) & (g99)));
	assign g574 = (((!sk[72]) & (!g572) & (!g233) & (!g160) & (g263) & (!g573)) + ((!sk[72]) & (!g572) & (!g233) & (!g160) & (g263) & (g573)) + ((!sk[72]) & (!g572) & (!g233) & (g160) & (!g263) & (!g573)) + ((!sk[72]) & (!g572) & (!g233) & (g160) & (!g263) & (g573)) + ((!sk[72]) & (!g572) & (!g233) & (g160) & (g263) & (!g573)) + ((!sk[72]) & (!g572) & (!g233) & (g160) & (g263) & (g573)) + ((!sk[72]) & (!g572) & (g233) & (!g160) & (!g263) & (!g573)) + ((!sk[72]) & (!g572) & (g233) & (!g160) & (!g263) & (g573)) + ((!sk[72]) & (!g572) & (g233) & (!g160) & (g263) & (!g573)) + ((!sk[72]) & (!g572) & (g233) & (!g160) & (g263) & (g573)) + ((!sk[72]) & (!g572) & (g233) & (g160) & (!g263) & (!g573)) + ((!sk[72]) & (!g572) & (g233) & (g160) & (!g263) & (g573)) + ((!sk[72]) & (!g572) & (g233) & (g160) & (g263) & (!g573)) + ((!sk[72]) & (!g572) & (g233) & (g160) & (g263) & (g573)) + ((!sk[72]) & (g572) & (!g233) & (!g160) & (g263) & (!g573)) + ((!sk[72]) & (g572) & (!g233) & (!g160) & (g263) & (g573)) + ((!sk[72]) & (g572) & (!g233) & (g160) & (!g263) & (!g573)) + ((!sk[72]) & (g572) & (!g233) & (g160) & (!g263) & (g573)) + ((!sk[72]) & (g572) & (!g233) & (g160) & (g263) & (!g573)) + ((!sk[72]) & (g572) & (!g233) & (g160) & (g263) & (g573)) + ((!sk[72]) & (g572) & (g233) & (!g160) & (!g263) & (!g573)) + ((!sk[72]) & (g572) & (g233) & (!g160) & (!g263) & (g573)) + ((!sk[72]) & (g572) & (g233) & (!g160) & (g263) & (!g573)) + ((!sk[72]) & (g572) & (g233) & (!g160) & (g263) & (g573)) + ((!sk[72]) & (g572) & (g233) & (g160) & (!g263) & (!g573)) + ((!sk[72]) & (g572) & (g233) & (g160) & (!g263) & (g573)) + ((!sk[72]) & (g572) & (g233) & (g160) & (g263) & (!g573)) + ((!sk[72]) & (g572) & (g233) & (g160) & (g263) & (g573)) + ((sk[72]) & (!g572) & (!g233) & (g160) & (!g263) & (!g573)));
	assign g575 = (((!sk[73]) & (!g38) & (!g9) & (!g25) & (g27)) + ((!sk[73]) & (!g38) & (!g9) & (g25) & (g27)) + ((!sk[73]) & (!g38) & (g9) & (!g25) & (g27)) + ((!sk[73]) & (!g38) & (g9) & (g25) & (g27)) + ((!sk[73]) & (g38) & (!g9) & (!g25) & (!g27)) + ((!sk[73]) & (g38) & (!g9) & (!g25) & (g27)) + ((!sk[73]) & (g38) & (!g9) & (g25) & (!g27)) + ((!sk[73]) & (g38) & (!g9) & (g25) & (g27)) + ((!sk[73]) & (g38) & (g9) & (!g25) & (!g27)) + ((!sk[73]) & (g38) & (g9) & (!g25) & (g27)) + ((!sk[73]) & (g38) & (g9) & (g25) & (!g27)) + ((!sk[73]) & (g38) & (g9) & (g25) & (g27)) + ((sk[73]) & (!g38) & (g9) & (!g25) & (g27)) + ((sk[73]) & (!g38) & (g9) & (g25) & (!g27)) + ((sk[73]) & (!g38) & (g9) & (g25) & (g27)) + ((sk[73]) & (g38) & (g9) & (!g25) & (!g27)) + ((sk[73]) & (g38) & (g9) & (!g25) & (g27)) + ((sk[73]) & (g38) & (g9) & (g25) & (!g27)) + ((sk[73]) & (g38) & (g9) & (g25) & (g27)));
	assign g576 = (((!g99) & (!g18) & (!g104) & (!sk[74]) & (g41) & (!g575)) + ((!g99) & (!g18) & (!g104) & (!sk[74]) & (g41) & (g575)) + ((!g99) & (!g18) & (!g104) & (sk[74]) & (!g41) & (!g575)) + ((!g99) & (!g18) & (!g104) & (sk[74]) & (g41) & (!g575)) + ((!g99) & (!g18) & (g104) & (!sk[74]) & (!g41) & (!g575)) + ((!g99) & (!g18) & (g104) & (!sk[74]) & (!g41) & (g575)) + ((!g99) & (!g18) & (g104) & (!sk[74]) & (g41) & (!g575)) + ((!g99) & (!g18) & (g104) & (!sk[74]) & (g41) & (g575)) + ((!g99) & (!g18) & (g104) & (sk[74]) & (!g41) & (!g575)) + ((!g99) & (!g18) & (g104) & (sk[74]) & (g41) & (!g575)) + ((!g99) & (g18) & (!g104) & (!sk[74]) & (!g41) & (!g575)) + ((!g99) & (g18) & (!g104) & (!sk[74]) & (!g41) & (g575)) + ((!g99) & (g18) & (!g104) & (!sk[74]) & (g41) & (!g575)) + ((!g99) & (g18) & (!g104) & (!sk[74]) & (g41) & (g575)) + ((!g99) & (g18) & (!g104) & (sk[74]) & (!g41) & (!g575)) + ((!g99) & (g18) & (!g104) & (sk[74]) & (g41) & (!g575)) + ((!g99) & (g18) & (g104) & (!sk[74]) & (!g41) & (!g575)) + ((!g99) & (g18) & (g104) & (!sk[74]) & (!g41) & (g575)) + ((!g99) & (g18) & (g104) & (!sk[74]) & (g41) & (!g575)) + ((!g99) & (g18) & (g104) & (!sk[74]) & (g41) & (g575)) + ((g99) & (!g18) & (!g104) & (!sk[74]) & (g41) & (!g575)) + ((g99) & (!g18) & (!g104) & (!sk[74]) & (g41) & (g575)) + ((g99) & (!g18) & (!g104) & (sk[74]) & (!g41) & (!g575)) + ((g99) & (!g18) & (g104) & (!sk[74]) & (!g41) & (!g575)) + ((g99) & (!g18) & (g104) & (!sk[74]) & (!g41) & (g575)) + ((g99) & (!g18) & (g104) & (!sk[74]) & (g41) & (!g575)) + ((g99) & (!g18) & (g104) & (!sk[74]) & (g41) & (g575)) + ((g99) & (!g18) & (g104) & (sk[74]) & (!g41) & (!g575)) + ((g99) & (g18) & (!g104) & (!sk[74]) & (!g41) & (!g575)) + ((g99) & (g18) & (!g104) & (!sk[74]) & (!g41) & (g575)) + ((g99) & (g18) & (!g104) & (!sk[74]) & (g41) & (!g575)) + ((g99) & (g18) & (!g104) & (!sk[74]) & (g41) & (g575)) + ((g99) & (g18) & (g104) & (!sk[74]) & (!g41) & (!g575)) + ((g99) & (g18) & (g104) & (!sk[74]) & (!g41) & (g575)) + ((g99) & (g18) & (g104) & (!sk[74]) & (g41) & (!g575)) + ((g99) & (g18) & (g104) & (!sk[74]) & (g41) & (g575)));
	assign g577 = (((!g70) & (!g42) & (!sk[75]) & (!g103) & (g576)) + ((!g70) & (!g42) & (!sk[75]) & (g103) & (g576)) + ((!g70) & (!g42) & (sk[75]) & (g103) & (g576)) + ((!g70) & (g42) & (!sk[75]) & (!g103) & (g576)) + ((!g70) & (g42) & (!sk[75]) & (g103) & (g576)) + ((!g70) & (g42) & (sk[75]) & (g103) & (g576)) + ((g70) & (!g42) & (!sk[75]) & (!g103) & (!g576)) + ((g70) & (!g42) & (!sk[75]) & (!g103) & (g576)) + ((g70) & (!g42) & (!sk[75]) & (g103) & (!g576)) + ((g70) & (!g42) & (!sk[75]) & (g103) & (g576)) + ((g70) & (!g42) & (sk[75]) & (g103) & (g576)) + ((g70) & (g42) & (!sk[75]) & (!g103) & (!g576)) + ((g70) & (g42) & (!sk[75]) & (!g103) & (g576)) + ((g70) & (g42) & (!sk[75]) & (g103) & (!g576)) + ((g70) & (g42) & (!sk[75]) & (g103) & (g576)));
	assign g578 = (((!g153) & (!g154) & (!sk[76]) & (!g358) & (g577)) + ((!g153) & (!g154) & (!sk[76]) & (g358) & (g577)) + ((!g153) & (!g154) & (sk[76]) & (g358) & (g577)) + ((!g153) & (g154) & (!sk[76]) & (!g358) & (g577)) + ((!g153) & (g154) & (!sk[76]) & (g358) & (g577)) + ((g153) & (!g154) & (!sk[76]) & (!g358) & (!g577)) + ((g153) & (!g154) & (!sk[76]) & (!g358) & (g577)) + ((g153) & (!g154) & (!sk[76]) & (g358) & (!g577)) + ((g153) & (!g154) & (!sk[76]) & (g358) & (g577)) + ((g153) & (g154) & (!sk[76]) & (!g358) & (!g577)) + ((g153) & (g154) & (!sk[76]) & (!g358) & (g577)) + ((g153) & (g154) & (!sk[76]) & (g358) & (!g577)) + ((g153) & (g154) & (!sk[76]) & (g358) & (g577)));
	assign g579 = (((!g9) & (!g58) & (sk[77]) & (!g288)) + ((!g9) & (g58) & (!sk[77]) & (!g288)) + ((!g9) & (g58) & (!sk[77]) & (g288)) + ((!g9) & (g58) & (sk[77]) & (!g288)) + ((g9) & (!g58) & (sk[77]) & (!g288)) + ((g9) & (g58) & (!sk[77]) & (!g288)) + ((g9) & (g58) & (!sk[77]) & (g288)));
	assign g580 = (((!g9) & (!g16) & (!sk[78]) & (!g30) & (g133)) + ((!g9) & (!g16) & (!sk[78]) & (g30) & (g133)) + ((!g9) & (g16) & (!sk[78]) & (!g30) & (g133)) + ((!g9) & (g16) & (!sk[78]) & (g30) & (g133)) + ((!g9) & (g16) & (sk[78]) & (g30) & (!g133)) + ((!g9) & (g16) & (sk[78]) & (g30) & (g133)) + ((g9) & (!g16) & (!sk[78]) & (!g30) & (!g133)) + ((g9) & (!g16) & (!sk[78]) & (!g30) & (g133)) + ((g9) & (!g16) & (!sk[78]) & (g30) & (!g133)) + ((g9) & (!g16) & (!sk[78]) & (g30) & (g133)) + ((g9) & (!g16) & (sk[78]) & (!g30) & (g133)) + ((g9) & (!g16) & (sk[78]) & (g30) & (g133)) + ((g9) & (g16) & (!sk[78]) & (!g30) & (!g133)) + ((g9) & (g16) & (!sk[78]) & (!g30) & (g133)) + ((g9) & (g16) & (!sk[78]) & (g30) & (!g133)) + ((g9) & (g16) & (!sk[78]) & (g30) & (g133)) + ((g9) & (g16) & (sk[78]) & (!g30) & (g133)) + ((g9) & (g16) & (sk[78]) & (g30) & (!g133)) + ((g9) & (g16) & (sk[78]) & (g30) & (g133)));
	assign g581 = (((!g147) & (!g81) & (!sk[79]) & (!g579) & (g580)) + ((!g147) & (!g81) & (!sk[79]) & (g579) & (g580)) + ((!g147) & (!g81) & (sk[79]) & (g579) & (!g580)) + ((!g147) & (g81) & (!sk[79]) & (!g579) & (g580)) + ((!g147) & (g81) & (!sk[79]) & (g579) & (g580)) + ((g147) & (!g81) & (!sk[79]) & (!g579) & (!g580)) + ((g147) & (!g81) & (!sk[79]) & (!g579) & (g580)) + ((g147) & (!g81) & (!sk[79]) & (g579) & (!g580)) + ((g147) & (!g81) & (!sk[79]) & (g579) & (g580)) + ((g147) & (g81) & (!sk[79]) & (!g579) & (!g580)) + ((g147) & (g81) & (!sk[79]) & (!g579) & (g580)) + ((g147) & (g81) & (!sk[79]) & (g579) & (!g580)) + ((g147) & (g81) & (!sk[79]) & (g579) & (g580)));
	assign g582 = (((!sk[80]) & (!g70) & (g27) & (!g87)) + ((!sk[80]) & (!g70) & (g27) & (g87)) + ((!sk[80]) & (g70) & (g27) & (!g87)) + ((!sk[80]) & (g70) & (g27) & (g87)) + ((sk[80]) & (!g70) & (!g27) & (!g87)) + ((sk[80]) & (!g70) & (g27) & (!g87)) + ((sk[80]) & (g70) & (!g27) & (!g87)));
	assign g583 = (((!g70) & (!sk[81]) & (!g71) & (!g58) & (g18) & (!g582)) + ((!g70) & (!sk[81]) & (!g71) & (!g58) & (g18) & (g582)) + ((!g70) & (!sk[81]) & (!g71) & (g58) & (!g18) & (!g582)) + ((!g70) & (!sk[81]) & (!g71) & (g58) & (!g18) & (g582)) + ((!g70) & (!sk[81]) & (!g71) & (g58) & (g18) & (!g582)) + ((!g70) & (!sk[81]) & (!g71) & (g58) & (g18) & (g582)) + ((!g70) & (!sk[81]) & (g71) & (!g58) & (!g18) & (!g582)) + ((!g70) & (!sk[81]) & (g71) & (!g58) & (!g18) & (g582)) + ((!g70) & (!sk[81]) & (g71) & (!g58) & (g18) & (!g582)) + ((!g70) & (!sk[81]) & (g71) & (!g58) & (g18) & (g582)) + ((!g70) & (!sk[81]) & (g71) & (g58) & (!g18) & (!g582)) + ((!g70) & (!sk[81]) & (g71) & (g58) & (!g18) & (g582)) + ((!g70) & (!sk[81]) & (g71) & (g58) & (g18) & (!g582)) + ((!g70) & (!sk[81]) & (g71) & (g58) & (g18) & (g582)) + ((!g70) & (sk[81]) & (!g71) & (!g58) & (!g18) & (g582)) + ((!g70) & (sk[81]) & (!g71) & (!g58) & (g18) & (g582)) + ((!g70) & (sk[81]) & (!g71) & (g58) & (!g18) & (g582)) + ((!g70) & (sk[81]) & (!g71) & (g58) & (g18) & (g582)) + ((!g70) & (sk[81]) & (g71) & (!g58) & (!g18) & (g582)) + ((!g70) & (sk[81]) & (g71) & (!g58) & (g18) & (g582)) + ((g70) & (!sk[81]) & (!g71) & (!g58) & (g18) & (!g582)) + ((g70) & (!sk[81]) & (!g71) & (!g58) & (g18) & (g582)) + ((g70) & (!sk[81]) & (!g71) & (g58) & (!g18) & (!g582)) + ((g70) & (!sk[81]) & (!g71) & (g58) & (!g18) & (g582)) + ((g70) & (!sk[81]) & (!g71) & (g58) & (g18) & (!g582)) + ((g70) & (!sk[81]) & (!g71) & (g58) & (g18) & (g582)) + ((g70) & (!sk[81]) & (g71) & (!g58) & (!g18) & (!g582)) + ((g70) & (!sk[81]) & (g71) & (!g58) & (!g18) & (g582)) + ((g70) & (!sk[81]) & (g71) & (!g58) & (g18) & (!g582)) + ((g70) & (!sk[81]) & (g71) & (!g58) & (g18) & (g582)) + ((g70) & (!sk[81]) & (g71) & (g58) & (!g18) & (!g582)) + ((g70) & (!sk[81]) & (g71) & (g58) & (!g18) & (g582)) + ((g70) & (!sk[81]) & (g71) & (g58) & (g18) & (!g582)) + ((g70) & (!sk[81]) & (g71) & (g58) & (g18) & (g582)) + ((g70) & (sk[81]) & (!g71) & (!g58) & (!g18) & (g582)) + ((g70) & (sk[81]) & (g71) & (!g58) & (!g18) & (g582)));
	assign g584 = (((g345) & (g574) & (g558) & (g578) & (g581) & (g583)));
	assign g585 = (((!g387) & (!sk[83]) & (!g388) & (!g412) & (g547)) + ((!g387) & (!sk[83]) & (!g388) & (g412) & (g547)) + ((!g387) & (!sk[83]) & (g388) & (!g412) & (g547)) + ((!g387) & (!sk[83]) & (g388) & (g412) & (g547)) + ((!g387) & (sk[83]) & (!g388) & (!g412) & (!g547)) + ((!g387) & (sk[83]) & (g388) & (!g412) & (g547)) + ((!g387) & (sk[83]) & (g388) & (g412) & (!g547)) + ((!g387) & (sk[83]) & (g388) & (g412) & (g547)) + ((g387) & (!sk[83]) & (!g388) & (!g412) & (!g547)) + ((g387) & (!sk[83]) & (!g388) & (!g412) & (g547)) + ((g387) & (!sk[83]) & (!g388) & (g412) & (!g547)) + ((g387) & (!sk[83]) & (!g388) & (g412) & (g547)) + ((g387) & (!sk[83]) & (g388) & (!g412) & (!g547)) + ((g387) & (!sk[83]) & (g388) & (!g412) & (g547)) + ((g387) & (!sk[83]) & (g388) & (g412) & (!g547)) + ((g387) & (!sk[83]) & (g388) & (g412) & (g547)) + ((g387) & (sk[83]) & (!g388) & (!g412) & (g547)) + ((g387) & (sk[83]) & (!g388) & (g412) & (!g547)) + ((g387) & (sk[83]) & (!g388) & (g412) & (g547)) + ((g387) & (sk[83]) & (g388) & (!g412) & (!g547)));
	assign g586 = (((!g38) & (!g49) & (!g104) & (g173) & (!sk[84]) & (!g180)) + ((!g38) & (!g49) & (!g104) & (g173) & (!sk[84]) & (g180)) + ((!g38) & (!g49) & (!g104) & (g173) & (sk[84]) & (g180)) + ((!g38) & (!g49) & (g104) & (!g173) & (!sk[84]) & (!g180)) + ((!g38) & (!g49) & (g104) & (!g173) & (!sk[84]) & (g180)) + ((!g38) & (!g49) & (g104) & (g173) & (!sk[84]) & (!g180)) + ((!g38) & (!g49) & (g104) & (g173) & (!sk[84]) & (g180)) + ((!g38) & (!g49) & (g104) & (g173) & (sk[84]) & (g180)) + ((!g38) & (g49) & (!g104) & (!g173) & (!sk[84]) & (!g180)) + ((!g38) & (g49) & (!g104) & (!g173) & (!sk[84]) & (g180)) + ((!g38) & (g49) & (!g104) & (g173) & (!sk[84]) & (!g180)) + ((!g38) & (g49) & (!g104) & (g173) & (!sk[84]) & (g180)) + ((!g38) & (g49) & (!g104) & (g173) & (sk[84]) & (g180)) + ((!g38) & (g49) & (g104) & (!g173) & (!sk[84]) & (!g180)) + ((!g38) & (g49) & (g104) & (!g173) & (!sk[84]) & (g180)) + ((!g38) & (g49) & (g104) & (g173) & (!sk[84]) & (!g180)) + ((!g38) & (g49) & (g104) & (g173) & (!sk[84]) & (g180)) + ((g38) & (!g49) & (!g104) & (g173) & (!sk[84]) & (!g180)) + ((g38) & (!g49) & (!g104) & (g173) & (!sk[84]) & (g180)) + ((g38) & (!g49) & (!g104) & (g173) & (sk[84]) & (g180)) + ((g38) & (!g49) & (g104) & (!g173) & (!sk[84]) & (!g180)) + ((g38) & (!g49) & (g104) & (!g173) & (!sk[84]) & (g180)) + ((g38) & (!g49) & (g104) & (g173) & (!sk[84]) & (!g180)) + ((g38) & (!g49) & (g104) & (g173) & (!sk[84]) & (g180)) + ((g38) & (g49) & (!g104) & (!g173) & (!sk[84]) & (!g180)) + ((g38) & (g49) & (!g104) & (!g173) & (!sk[84]) & (g180)) + ((g38) & (g49) & (!g104) & (g173) & (!sk[84]) & (!g180)) + ((g38) & (g49) & (!g104) & (g173) & (!sk[84]) & (g180)) + ((g38) & (g49) & (!g104) & (g173) & (sk[84]) & (g180)) + ((g38) & (g49) & (g104) & (!g173) & (!sk[84]) & (!g180)) + ((g38) & (g49) & (g104) & (!g173) & (!sk[84]) & (g180)) + ((g38) & (g49) & (g104) & (g173) & (!sk[84]) & (!g180)) + ((g38) & (g49) & (g104) & (g173) & (!sk[84]) & (g180)));
	assign g587 = (((!g16) & (g104) & (!sk[85]) & (!g32)) + ((!g16) & (g104) & (!sk[85]) & (g32)) + ((!g16) & (g104) & (sk[85]) & (g32)) + ((g16) & (!g104) & (sk[85]) & (g32)) + ((g16) & (g104) & (!sk[85]) & (!g32)) + ((g16) & (g104) & (!sk[85]) & (g32)) + ((g16) & (g104) & (sk[85]) & (g32)));
	assign g588 = (((!g71) & (!g58) & (!g56) & (!sk[86]) & (g340) & (!g587)) + ((!g71) & (!g58) & (!g56) & (!sk[86]) & (g340) & (g587)) + ((!g71) & (!g58) & (g56) & (!sk[86]) & (!g340) & (!g587)) + ((!g71) & (!g58) & (g56) & (!sk[86]) & (!g340) & (g587)) + ((!g71) & (!g58) & (g56) & (!sk[86]) & (g340) & (!g587)) + ((!g71) & (!g58) & (g56) & (!sk[86]) & (g340) & (g587)) + ((!g71) & (!g58) & (g56) & (sk[86]) & (!g340) & (!g587)) + ((!g71) & (g58) & (!g56) & (!sk[86]) & (!g340) & (!g587)) + ((!g71) & (g58) & (!g56) & (!sk[86]) & (!g340) & (g587)) + ((!g71) & (g58) & (!g56) & (!sk[86]) & (g340) & (!g587)) + ((!g71) & (g58) & (!g56) & (!sk[86]) & (g340) & (g587)) + ((!g71) & (g58) & (g56) & (!sk[86]) & (!g340) & (!g587)) + ((!g71) & (g58) & (g56) & (!sk[86]) & (!g340) & (g587)) + ((!g71) & (g58) & (g56) & (!sk[86]) & (g340) & (!g587)) + ((!g71) & (g58) & (g56) & (!sk[86]) & (g340) & (g587)) + ((!g71) & (g58) & (g56) & (sk[86]) & (!g340) & (!g587)) + ((g71) & (!g58) & (!g56) & (!sk[86]) & (g340) & (!g587)) + ((g71) & (!g58) & (!g56) & (!sk[86]) & (g340) & (g587)) + ((g71) & (!g58) & (g56) & (!sk[86]) & (!g340) & (!g587)) + ((g71) & (!g58) & (g56) & (!sk[86]) & (!g340) & (g587)) + ((g71) & (!g58) & (g56) & (!sk[86]) & (g340) & (!g587)) + ((g71) & (!g58) & (g56) & (!sk[86]) & (g340) & (g587)) + ((g71) & (!g58) & (g56) & (sk[86]) & (!g340) & (!g587)) + ((g71) & (g58) & (!g56) & (!sk[86]) & (!g340) & (!g587)) + ((g71) & (g58) & (!g56) & (!sk[86]) & (!g340) & (g587)) + ((g71) & (g58) & (!g56) & (!sk[86]) & (g340) & (!g587)) + ((g71) & (g58) & (!g56) & (!sk[86]) & (g340) & (g587)) + ((g71) & (g58) & (g56) & (!sk[86]) & (!g340) & (!g587)) + ((g71) & (g58) & (g56) & (!sk[86]) & (!g340) & (g587)) + ((g71) & (g58) & (g56) & (!sk[86]) & (g340) & (!g587)) + ((g71) & (g58) & (g56) & (!sk[86]) & (g340) & (g587)));
	assign g589 = (((!g86) & (!g572) & (!sk[87]) & (!g204) & (g183) & (!g588)) + ((!g86) & (!g572) & (!sk[87]) & (!g204) & (g183) & (g588)) + ((!g86) & (!g572) & (!sk[87]) & (g204) & (!g183) & (!g588)) + ((!g86) & (!g572) & (!sk[87]) & (g204) & (!g183) & (g588)) + ((!g86) & (!g572) & (!sk[87]) & (g204) & (g183) & (!g588)) + ((!g86) & (!g572) & (!sk[87]) & (g204) & (g183) & (g588)) + ((!g86) & (!g572) & (sk[87]) & (!g204) & (g183) & (g588)) + ((!g86) & (g572) & (!sk[87]) & (!g204) & (!g183) & (!g588)) + ((!g86) & (g572) & (!sk[87]) & (!g204) & (!g183) & (g588)) + ((!g86) & (g572) & (!sk[87]) & (!g204) & (g183) & (!g588)) + ((!g86) & (g572) & (!sk[87]) & (!g204) & (g183) & (g588)) + ((!g86) & (g572) & (!sk[87]) & (g204) & (!g183) & (!g588)) + ((!g86) & (g572) & (!sk[87]) & (g204) & (!g183) & (g588)) + ((!g86) & (g572) & (!sk[87]) & (g204) & (g183) & (!g588)) + ((!g86) & (g572) & (!sk[87]) & (g204) & (g183) & (g588)) + ((g86) & (!g572) & (!sk[87]) & (!g204) & (g183) & (!g588)) + ((g86) & (!g572) & (!sk[87]) & (!g204) & (g183) & (g588)) + ((g86) & (!g572) & (!sk[87]) & (g204) & (!g183) & (!g588)) + ((g86) & (!g572) & (!sk[87]) & (g204) & (!g183) & (g588)) + ((g86) & (!g572) & (!sk[87]) & (g204) & (g183) & (!g588)) + ((g86) & (!g572) & (!sk[87]) & (g204) & (g183) & (g588)) + ((g86) & (g572) & (!sk[87]) & (!g204) & (!g183) & (!g588)) + ((g86) & (g572) & (!sk[87]) & (!g204) & (!g183) & (g588)) + ((g86) & (g572) & (!sk[87]) & (!g204) & (g183) & (!g588)) + ((g86) & (g572) & (!sk[87]) & (!g204) & (g183) & (g588)) + ((g86) & (g572) & (!sk[87]) & (g204) & (!g183) & (!g588)) + ((g86) & (g572) & (!sk[87]) & (g204) & (!g183) & (g588)) + ((g86) & (g572) & (!sk[87]) & (g204) & (g183) & (!g588)) + ((g86) & (g572) & (!sk[87]) & (g204) & (g183) & (g588)));
	assign g590 = (((!g99) & (!sk[88]) & (g32) & (!g141)) + ((!g99) & (!sk[88]) & (g32) & (g141)) + ((!g99) & (sk[88]) & (!g32) & (!g141)) + ((!g99) & (sk[88]) & (g32) & (!g141)) + ((g99) & (!sk[88]) & (g32) & (!g141)) + ((g99) & (!sk[88]) & (g32) & (g141)) + ((g99) & (sk[88]) & (!g32) & (!g141)));
	assign g591 = (((!g17) & (!sk[89]) & (g99) & (!g64)) + ((!g17) & (!sk[89]) & (g99) & (g64)) + ((!g17) & (sk[89]) & (!g99) & (!g64)) + ((!g17) & (sk[89]) & (g99) & (!g64)) + ((g17) & (!sk[89]) & (g99) & (!g64)) + ((g17) & (!sk[89]) & (g99) & (g64)) + ((g17) & (sk[89]) & (!g99) & (!g64)));
	assign g592 = (((!g79) & (!sk[90]) & (!g230) & (!g19) & (g590) & (!g591)) + ((!g79) & (!sk[90]) & (!g230) & (!g19) & (g590) & (g591)) + ((!g79) & (!sk[90]) & (!g230) & (g19) & (!g590) & (!g591)) + ((!g79) & (!sk[90]) & (!g230) & (g19) & (!g590) & (g591)) + ((!g79) & (!sk[90]) & (!g230) & (g19) & (g590) & (!g591)) + ((!g79) & (!sk[90]) & (!g230) & (g19) & (g590) & (g591)) + ((!g79) & (!sk[90]) & (g230) & (!g19) & (!g590) & (!g591)) + ((!g79) & (!sk[90]) & (g230) & (!g19) & (!g590) & (g591)) + ((!g79) & (!sk[90]) & (g230) & (!g19) & (g590) & (!g591)) + ((!g79) & (!sk[90]) & (g230) & (!g19) & (g590) & (g591)) + ((!g79) & (!sk[90]) & (g230) & (g19) & (!g590) & (!g591)) + ((!g79) & (!sk[90]) & (g230) & (g19) & (!g590) & (g591)) + ((!g79) & (!sk[90]) & (g230) & (g19) & (g590) & (!g591)) + ((!g79) & (!sk[90]) & (g230) & (g19) & (g590) & (g591)) + ((!g79) & (sk[90]) & (g230) & (!g19) & (g590) & (g591)) + ((g79) & (!sk[90]) & (!g230) & (!g19) & (g590) & (!g591)) + ((g79) & (!sk[90]) & (!g230) & (!g19) & (g590) & (g591)) + ((g79) & (!sk[90]) & (!g230) & (g19) & (!g590) & (!g591)) + ((g79) & (!sk[90]) & (!g230) & (g19) & (!g590) & (g591)) + ((g79) & (!sk[90]) & (!g230) & (g19) & (g590) & (!g591)) + ((g79) & (!sk[90]) & (!g230) & (g19) & (g590) & (g591)) + ((g79) & (!sk[90]) & (g230) & (!g19) & (!g590) & (!g591)) + ((g79) & (!sk[90]) & (g230) & (!g19) & (!g590) & (g591)) + ((g79) & (!sk[90]) & (g230) & (!g19) & (g590) & (!g591)) + ((g79) & (!sk[90]) & (g230) & (!g19) & (g590) & (g591)) + ((g79) & (!sk[90]) & (g230) & (g19) & (!g590) & (!g591)) + ((g79) & (!sk[90]) & (g230) & (g19) & (!g590) & (g591)) + ((g79) & (!sk[90]) & (g230) & (g19) & (g590) & (!g591)) + ((g79) & (!sk[90]) & (g230) & (g19) & (g590) & (g591)));
	assign g593 = (((!sk[91]) & (g16) & (g41)) + ((sk[91]) & (g16) & (g41)));
	assign g594 = (((!g9) & (!sk[92]) & (!g18) & (!g593) & (g73)) + ((!g9) & (!sk[92]) & (!g18) & (g593) & (g73)) + ((!g9) & (!sk[92]) & (g18) & (!g593) & (g73)) + ((!g9) & (!sk[92]) & (g18) & (g593) & (g73)) + ((!g9) & (sk[92]) & (!g18) & (!g593) & (!g73)) + ((!g9) & (sk[92]) & (g18) & (!g593) & (!g73)) + ((g9) & (!sk[92]) & (!g18) & (!g593) & (!g73)) + ((g9) & (!sk[92]) & (!g18) & (!g593) & (g73)) + ((g9) & (!sk[92]) & (!g18) & (g593) & (!g73)) + ((g9) & (!sk[92]) & (!g18) & (g593) & (g73)) + ((g9) & (!sk[92]) & (g18) & (!g593) & (!g73)) + ((g9) & (!sk[92]) & (g18) & (!g593) & (g73)) + ((g9) & (!sk[92]) & (g18) & (g593) & (!g73)) + ((g9) & (!sk[92]) & (g18) & (g593) & (g73)) + ((g9) & (sk[92]) & (!g18) & (!g593) & (!g73)));
	assign g595 = (((!g112) & (!g113) & (!g97) & (!g98) & (!g71) & (g594)) + ((!g112) & (!g113) & (!g97) & (!g98) & (g71) & (g594)) + ((!g112) & (!g113) & (!g97) & (g98) & (!g71) & (g594)) + ((!g112) & (!g113) & (!g97) & (g98) & (g71) & (g594)) + ((!g112) & (!g113) & (g97) & (!g98) & (!g71) & (g594)) + ((!g112) & (!g113) & (g97) & (!g98) & (g71) & (g594)) + ((!g112) & (!g113) & (g97) & (g98) & (!g71) & (g594)) + ((!g112) & (!g113) & (g97) & (g98) & (g71) & (g594)) + ((!g112) & (g113) & (!g97) & (!g98) & (!g71) & (g594)) + ((!g112) & (g113) & (!g97) & (!g98) & (g71) & (g594)) + ((!g112) & (g113) & (!g97) & (g98) & (!g71) & (g594)) + ((!g112) & (g113) & (!g97) & (g98) & (g71) & (g594)) + ((!g112) & (g113) & (g97) & (!g98) & (!g71) & (g594)) + ((!g112) & (g113) & (g97) & (!g98) & (g71) & (g594)) + ((!g112) & (g113) & (g97) & (g98) & (!g71) & (g594)) + ((!g112) & (g113) & (g97) & (g98) & (g71) & (g594)) + ((g112) & (!g113) & (!g97) & (!g98) & (!g71) & (g594)) + ((g112) & (!g113) & (!g97) & (g98) & (!g71) & (g594)) + ((g112) & (!g113) & (!g97) & (g98) & (g71) & (g594)) + ((g112) & (!g113) & (g97) & (!g98) & (!g71) & (g594)) + ((g112) & (!g113) & (g97) & (!g98) & (g71) & (g594)) + ((g112) & (!g113) & (g97) & (g98) & (!g71) & (g594)) + ((g112) & (!g113) & (g97) & (g98) & (g71) & (g594)) + ((g112) & (g113) & (!g97) & (!g98) & (!g71) & (g594)) + ((g112) & (g113) & (!g97) & (g98) & (!g71) & (g594)) + ((g112) & (g113) & (g97) & (!g98) & (!g71) & (g594)) + ((g112) & (g113) & (g97) & (g98) & (!g71) & (g594)) + ((g112) & (g113) & (g97) & (g98) & (g71) & (g594)));
	assign g596 = (((!g70) & (!g49) & (!g62) & (!g32) & (sk[94]) & (!g60)) + ((!g70) & (!g49) & (!g62) & (g32) & (!sk[94]) & (!g60)) + ((!g70) & (!g49) & (!g62) & (g32) & (!sk[94]) & (g60)) + ((!g70) & (!g49) & (!g62) & (g32) & (sk[94]) & (!g60)) + ((!g70) & (!g49) & (g62) & (!g32) & (!sk[94]) & (!g60)) + ((!g70) & (!g49) & (g62) & (!g32) & (!sk[94]) & (g60)) + ((!g70) & (!g49) & (g62) & (!g32) & (sk[94]) & (!g60)) + ((!g70) & (!g49) & (g62) & (g32) & (!sk[94]) & (!g60)) + ((!g70) & (!g49) & (g62) & (g32) & (!sk[94]) & (g60)) + ((!g70) & (!g49) & (g62) & (g32) & (sk[94]) & (!g60)) + ((!g70) & (g49) & (!g62) & (!g32) & (!sk[94]) & (!g60)) + ((!g70) & (g49) & (!g62) & (!g32) & (!sk[94]) & (g60)) + ((!g70) & (g49) & (!g62) & (!g32) & (sk[94]) & (!g60)) + ((!g70) & (g49) & (!g62) & (g32) & (!sk[94]) & (!g60)) + ((!g70) & (g49) & (!g62) & (g32) & (!sk[94]) & (g60)) + ((!g70) & (g49) & (!g62) & (g32) & (sk[94]) & (!g60)) + ((!g70) & (g49) & (g62) & (!g32) & (!sk[94]) & (!g60)) + ((!g70) & (g49) & (g62) & (!g32) & (!sk[94]) & (g60)) + ((!g70) & (g49) & (g62) & (g32) & (!sk[94]) & (!g60)) + ((!g70) & (g49) & (g62) & (g32) & (!sk[94]) & (g60)) + ((g70) & (!g49) & (!g62) & (!g32) & (sk[94]) & (!g60)) + ((g70) & (!g49) & (!g62) & (g32) & (!sk[94]) & (!g60)) + ((g70) & (!g49) & (!g62) & (g32) & (!sk[94]) & (g60)) + ((g70) & (!g49) & (g62) & (!g32) & (!sk[94]) & (!g60)) + ((g70) & (!g49) & (g62) & (!g32) & (!sk[94]) & (g60)) + ((g70) & (!g49) & (g62) & (!g32) & (sk[94]) & (!g60)) + ((g70) & (!g49) & (g62) & (g32) & (!sk[94]) & (!g60)) + ((g70) & (!g49) & (g62) & (g32) & (!sk[94]) & (g60)) + ((g70) & (g49) & (!g62) & (!g32) & (!sk[94]) & (!g60)) + ((g70) & (g49) & (!g62) & (!g32) & (!sk[94]) & (g60)) + ((g70) & (g49) & (!g62) & (g32) & (!sk[94]) & (!g60)) + ((g70) & (g49) & (!g62) & (g32) & (!sk[94]) & (g60)) + ((g70) & (g49) & (g62) & (!g32) & (!sk[94]) & (!g60)) + ((g70) & (g49) & (g62) & (!g32) & (!sk[94]) & (g60)) + ((g70) & (g49) & (g62) & (g32) & (!sk[94]) & (!g60)) + ((g70) & (g49) & (g62) & (g32) & (!sk[94]) & (g60)));
	assign g597 = (((g261) & (g586) & (g589) & (g592) & (g595) & (g596)));
	assign g598 = (((!g413) & (!g440) & (!g441) & (!g454) & (!g455) & (!g546)) + ((!g413) & (!g440) & (!g441) & (!g454) & (!g455) & (g546)) + ((!g413) & (!g440) & (!g441) & (!g454) & (g455) & (!g546)) + ((!g413) & (!g440) & (!g441) & (!g454) & (g455) & (g546)) + ((!g413) & (!g440) & (!g441) & (g454) & (!g455) & (!g546)) + ((!g413) & (!g440) & (!g441) & (g454) & (!g455) & (g546)) + ((!g413) & (!g440) & (!g441) & (g454) & (g455) & (!g546)) + ((!g413) & (!g440) & (!g441) & (g454) & (g455) & (g546)) + ((!g413) & (!g440) & (g441) & (!g454) & (!g455) & (!g546)) + ((!g413) & (!g440) & (g441) & (!g454) & (!g455) & (g546)) + ((!g413) & (!g440) & (g441) & (!g454) & (g455) & (g546)) + ((!g413) & (!g440) & (g441) & (g454) & (!g455) & (g546)) + ((!g413) & (g440) & (!g441) & (!g454) & (!g455) & (!g546)) + ((!g413) & (g440) & (!g441) & (!g454) & (!g455) & (g546)) + ((!g413) & (g440) & (!g441) & (!g454) & (g455) & (g546)) + ((!g413) & (g440) & (!g441) & (g454) & (!g455) & (g546)) + ((g413) & (!g440) & (g441) & (!g454) & (g455) & (!g546)) + ((g413) & (!g440) & (g441) & (g454) & (!g455) & (!g546)) + ((g413) & (!g440) & (g441) & (g454) & (g455) & (!g546)) + ((g413) & (!g440) & (g441) & (g454) & (g455) & (g546)) + ((g413) & (g440) & (!g441) & (!g454) & (g455) & (!g546)) + ((g413) & (g440) & (!g441) & (g454) & (!g455) & (!g546)) + ((g413) & (g440) & (!g441) & (g454) & (g455) & (!g546)) + ((g413) & (g440) & (!g441) & (g454) & (g455) & (g546)) + ((g413) & (g440) & (g441) & (!g454) & (!g455) & (!g546)) + ((g413) & (g440) & (g441) & (!g454) & (!g455) & (g546)) + ((g413) & (g440) & (g441) & (!g454) & (g455) & (!g546)) + ((g413) & (g440) & (g441) & (!g454) & (g455) & (g546)) + ((g413) & (g440) & (g441) & (g454) & (!g455) & (!g546)) + ((g413) & (g440) & (g441) & (g454) & (!g455) & (g546)) + ((g413) & (g440) & (g441) & (g454) & (g455) & (!g546)) + ((g413) & (g440) & (g441) & (g454) & (g455) & (g546)));
	assign g599 = (((!sk[97]) & (g126) & (g135)) + ((sk[97]) & (g126) & (g135)));
	assign g600 = (((!g57) & (!g32) & (!g193) & (!sk[98]) & (g187)) + ((!g57) & (!g32) & (!g193) & (sk[98]) & (!g187)) + ((!g57) & (!g32) & (g193) & (!sk[98]) & (g187)) + ((!g57) & (g32) & (!g193) & (!sk[98]) & (g187)) + ((!g57) & (g32) & (!g193) & (sk[98]) & (!g187)) + ((!g57) & (g32) & (g193) & (!sk[98]) & (g187)) + ((g57) & (!g32) & (!g193) & (!sk[98]) & (!g187)) + ((g57) & (!g32) & (!g193) & (!sk[98]) & (g187)) + ((g57) & (!g32) & (!g193) & (sk[98]) & (!g187)) + ((g57) & (!g32) & (g193) & (!sk[98]) & (!g187)) + ((g57) & (!g32) & (g193) & (!sk[98]) & (g187)) + ((g57) & (g32) & (!g193) & (!sk[98]) & (!g187)) + ((g57) & (g32) & (!g193) & (!sk[98]) & (g187)) + ((g57) & (g32) & (g193) & (!sk[98]) & (!g187)) + ((g57) & (g32) & (g193) & (!sk[98]) & (g187)));
	assign g601 = (((g71) & (!sk[99]) & (g41)) + ((g71) & (sk[99]) & (g41)));
	assign g602 = (((!g70) & (!g238) & (!g32) & (!sk[100]) & (g354)) + ((!g70) & (!g238) & (!g32) & (sk[100]) & (!g354)) + ((!g70) & (!g238) & (g32) & (!sk[100]) & (g354)) + ((!g70) & (!g238) & (g32) & (sk[100]) & (!g354)) + ((!g70) & (g238) & (!g32) & (!sk[100]) & (g354)) + ((!g70) & (g238) & (g32) & (!sk[100]) & (g354)) + ((g70) & (!g238) & (!g32) & (!sk[100]) & (!g354)) + ((g70) & (!g238) & (!g32) & (!sk[100]) & (g354)) + ((g70) & (!g238) & (!g32) & (sk[100]) & (!g354)) + ((g70) & (!g238) & (g32) & (!sk[100]) & (!g354)) + ((g70) & (!g238) & (g32) & (!sk[100]) & (g354)) + ((g70) & (g238) & (!g32) & (!sk[100]) & (!g354)) + ((g70) & (g238) & (!g32) & (!sk[100]) & (g354)) + ((g70) & (g238) & (g32) & (!sk[100]) & (!g354)) + ((g70) & (g238) & (g32) & (!sk[100]) & (g354)));
	assign g603 = (((!sk[101]) & (!g70) & (!g99) & (!g18) & (g20)) + ((!sk[101]) & (!g70) & (!g99) & (g18) & (g20)) + ((!sk[101]) & (!g70) & (g99) & (!g18) & (g20)) + ((!sk[101]) & (!g70) & (g99) & (g18) & (g20)) + ((!sk[101]) & (g70) & (!g99) & (!g18) & (!g20)) + ((!sk[101]) & (g70) & (!g99) & (!g18) & (g20)) + ((!sk[101]) & (g70) & (!g99) & (g18) & (!g20)) + ((!sk[101]) & (g70) & (!g99) & (g18) & (g20)) + ((!sk[101]) & (g70) & (g99) & (!g18) & (!g20)) + ((!sk[101]) & (g70) & (g99) & (!g18) & (g20)) + ((!sk[101]) & (g70) & (g99) & (g18) & (!g20)) + ((!sk[101]) & (g70) & (g99) & (g18) & (g20)) + ((sk[101]) & (!g70) & (g99) & (!g18) & (g20)) + ((sk[101]) & (!g70) & (g99) & (g18) & (g20)) + ((sk[101]) & (g70) & (!g99) & (g18) & (!g20)) + ((sk[101]) & (g70) & (!g99) & (g18) & (g20)) + ((sk[101]) & (g70) & (g99) & (!g18) & (g20)) + ((sk[101]) & (g70) & (g99) & (g18) & (!g20)) + ((sk[101]) & (g70) & (g99) & (g18) & (g20)));
	assign g604 = (((!g162) & (!sk[102]) & (!g337) & (!g602) & (g603)) + ((!g162) & (!sk[102]) & (!g337) & (g602) & (g603)) + ((!g162) & (!sk[102]) & (g337) & (!g602) & (g603)) + ((!g162) & (!sk[102]) & (g337) & (g602) & (g603)) + ((!g162) & (sk[102]) & (g337) & (g602) & (!g603)) + ((g162) & (!sk[102]) & (!g337) & (!g602) & (!g603)) + ((g162) & (!sk[102]) & (!g337) & (!g602) & (g603)) + ((g162) & (!sk[102]) & (!g337) & (g602) & (!g603)) + ((g162) & (!sk[102]) & (!g337) & (g602) & (g603)) + ((g162) & (!sk[102]) & (g337) & (!g602) & (!g603)) + ((g162) & (!sk[102]) & (g337) & (!g602) & (g603)) + ((g162) & (!sk[102]) & (g337) & (g602) & (!g603)) + ((g162) & (!sk[102]) & (g337) & (g602) & (g603)));
	assign g605 = (((!g601) & (!g80) & (sk[103]) & (g604)) + ((!g601) & (g80) & (!sk[103]) & (!g604)) + ((!g601) & (g80) & (!sk[103]) & (g604)) + ((g601) & (g80) & (!sk[103]) & (!g604)) + ((g601) & (g80) & (!sk[103]) & (g604)));
	assign g606 = (((!g79) & (!g267) & (!sk[104]) & (!g52) & (g255)) + ((!g79) & (!g267) & (!sk[104]) & (g52) & (g255)) + ((!g79) & (!g267) & (sk[104]) & (g52) & (g255)) + ((!g79) & (g267) & (!sk[104]) & (!g52) & (g255)) + ((!g79) & (g267) & (!sk[104]) & (g52) & (g255)) + ((g79) & (!g267) & (!sk[104]) & (!g52) & (!g255)) + ((g79) & (!g267) & (!sk[104]) & (!g52) & (g255)) + ((g79) & (!g267) & (!sk[104]) & (g52) & (!g255)) + ((g79) & (!g267) & (!sk[104]) & (g52) & (g255)) + ((g79) & (g267) & (!sk[104]) & (!g52) & (!g255)) + ((g79) & (g267) & (!sk[104]) & (!g52) & (g255)) + ((g79) & (g267) & (!sk[104]) & (g52) & (!g255)) + ((g79) & (g267) & (!sk[104]) & (g52) & (g255)));
	assign g607 = (((!g70) & (!sk[105]) & (!g46) & (!g40) & (g41)) + ((!g70) & (!sk[105]) & (!g46) & (g40) & (g41)) + ((!g70) & (!sk[105]) & (g46) & (!g40) & (g41)) + ((!g70) & (!sk[105]) & (g46) & (g40) & (g41)) + ((!g70) & (sk[105]) & (g46) & (g40) & (!g41)) + ((!g70) & (sk[105]) & (g46) & (g40) & (g41)) + ((g70) & (!sk[105]) & (!g46) & (!g40) & (!g41)) + ((g70) & (!sk[105]) & (!g46) & (!g40) & (g41)) + ((g70) & (!sk[105]) & (!g46) & (g40) & (!g41)) + ((g70) & (!sk[105]) & (!g46) & (g40) & (g41)) + ((g70) & (!sk[105]) & (g46) & (!g40) & (!g41)) + ((g70) & (!sk[105]) & (g46) & (!g40) & (g41)) + ((g70) & (!sk[105]) & (g46) & (g40) & (!g41)) + ((g70) & (!sk[105]) & (g46) & (g40) & (g41)) + ((g70) & (sk[105]) & (!g46) & (!g40) & (g41)) + ((g70) & (sk[105]) & (!g46) & (g40) & (!g41)) + ((g70) & (sk[105]) & (!g46) & (g40) & (g41)) + ((g70) & (sk[105]) & (g46) & (!g40) & (g41)) + ((g70) & (sk[105]) & (g46) & (g40) & (!g41)) + ((g70) & (sk[105]) & (g46) & (g40) & (g41)));
	assign g608 = (((!sk[106]) & (!g10) & (!g17) & (!g99) & (g551) & (!g607)) + ((!sk[106]) & (!g10) & (!g17) & (!g99) & (g551) & (g607)) + ((!sk[106]) & (!g10) & (!g17) & (g99) & (!g551) & (!g607)) + ((!sk[106]) & (!g10) & (!g17) & (g99) & (!g551) & (g607)) + ((!sk[106]) & (!g10) & (!g17) & (g99) & (g551) & (!g607)) + ((!sk[106]) & (!g10) & (!g17) & (g99) & (g551) & (g607)) + ((!sk[106]) & (!g10) & (g17) & (!g99) & (!g551) & (!g607)) + ((!sk[106]) & (!g10) & (g17) & (!g99) & (!g551) & (g607)) + ((!sk[106]) & (!g10) & (g17) & (!g99) & (g551) & (!g607)) + ((!sk[106]) & (!g10) & (g17) & (!g99) & (g551) & (g607)) + ((!sk[106]) & (!g10) & (g17) & (g99) & (!g551) & (!g607)) + ((!sk[106]) & (!g10) & (g17) & (g99) & (!g551) & (g607)) + ((!sk[106]) & (!g10) & (g17) & (g99) & (g551) & (!g607)) + ((!sk[106]) & (!g10) & (g17) & (g99) & (g551) & (g607)) + ((!sk[106]) & (g10) & (!g17) & (!g99) & (g551) & (!g607)) + ((!sk[106]) & (g10) & (!g17) & (!g99) & (g551) & (g607)) + ((!sk[106]) & (g10) & (!g17) & (g99) & (!g551) & (!g607)) + ((!sk[106]) & (g10) & (!g17) & (g99) & (!g551) & (g607)) + ((!sk[106]) & (g10) & (!g17) & (g99) & (g551) & (!g607)) + ((!sk[106]) & (g10) & (!g17) & (g99) & (g551) & (g607)) + ((!sk[106]) & (g10) & (g17) & (!g99) & (!g551) & (!g607)) + ((!sk[106]) & (g10) & (g17) & (!g99) & (!g551) & (g607)) + ((!sk[106]) & (g10) & (g17) & (!g99) & (g551) & (!g607)) + ((!sk[106]) & (g10) & (g17) & (!g99) & (g551) & (g607)) + ((!sk[106]) & (g10) & (g17) & (g99) & (!g551) & (!g607)) + ((!sk[106]) & (g10) & (g17) & (g99) & (!g551) & (g607)) + ((!sk[106]) & (g10) & (g17) & (g99) & (g551) & (!g607)) + ((!sk[106]) & (g10) & (g17) & (g99) & (g551) & (g607)) + ((sk[106]) & (!g10) & (!g17) & (!g99) & (!g551) & (!g607)) + ((sk[106]) & (!g10) & (!g17) & (g99) & (!g551) & (!g607)) + ((sk[106]) & (!g10) & (g17) & (!g99) & (!g551) & (!g607)) + ((sk[106]) & (g10) & (!g17) & (!g99) & (!g551) & (!g607)) + ((sk[106]) & (g10) & (g17) & (!g99) & (!g551) & (!g607)));
	assign g609 = (((!g38) & (!g70) & (!g104) & (!g25) & (sk[107]) & (!g66)) + ((!g38) & (!g70) & (!g104) & (!g25) & (sk[107]) & (g66)) + ((!g38) & (!g70) & (!g104) & (g25) & (!sk[107]) & (!g66)) + ((!g38) & (!g70) & (!g104) & (g25) & (!sk[107]) & (g66)) + ((!g38) & (!g70) & (!g104) & (g25) & (sk[107]) & (!g66)) + ((!g38) & (!g70) & (!g104) & (g25) & (sk[107]) & (g66)) + ((!g38) & (!g70) & (g104) & (!g25) & (!sk[107]) & (!g66)) + ((!g38) & (!g70) & (g104) & (!g25) & (!sk[107]) & (g66)) + ((!g38) & (!g70) & (g104) & (!g25) & (sk[107]) & (!g66)) + ((!g38) & (!g70) & (g104) & (!g25) & (sk[107]) & (g66)) + ((!g38) & (!g70) & (g104) & (g25) & (!sk[107]) & (!g66)) + ((!g38) & (!g70) & (g104) & (g25) & (!sk[107]) & (g66)) + ((!g38) & (!g70) & (g104) & (g25) & (sk[107]) & (!g66)) + ((!g38) & (!g70) & (g104) & (g25) & (sk[107]) & (g66)) + ((!g38) & (g70) & (!g104) & (!g25) & (!sk[107]) & (!g66)) + ((!g38) & (g70) & (!g104) & (!g25) & (!sk[107]) & (g66)) + ((!g38) & (g70) & (!g104) & (!g25) & (sk[107]) & (!g66)) + ((!g38) & (g70) & (!g104) & (g25) & (!sk[107]) & (!g66)) + ((!g38) & (g70) & (!g104) & (g25) & (!sk[107]) & (g66)) + ((!g38) & (g70) & (g104) & (!g25) & (!sk[107]) & (!g66)) + ((!g38) & (g70) & (g104) & (!g25) & (!sk[107]) & (g66)) + ((!g38) & (g70) & (g104) & (!g25) & (sk[107]) & (!g66)) + ((!g38) & (g70) & (g104) & (g25) & (!sk[107]) & (!g66)) + ((!g38) & (g70) & (g104) & (g25) & (!sk[107]) & (g66)) + ((g38) & (!g70) & (!g104) & (!g25) & (sk[107]) & (!g66)) + ((g38) & (!g70) & (!g104) & (!g25) & (sk[107]) & (g66)) + ((g38) & (!g70) & (!g104) & (g25) & (!sk[107]) & (!g66)) + ((g38) & (!g70) & (!g104) & (g25) & (!sk[107]) & (g66)) + ((g38) & (!g70) & (!g104) & (g25) & (sk[107]) & (!g66)) + ((g38) & (!g70) & (!g104) & (g25) & (sk[107]) & (g66)) + ((g38) & (!g70) & (g104) & (!g25) & (!sk[107]) & (!g66)) + ((g38) & (!g70) & (g104) & (!g25) & (!sk[107]) & (g66)) + ((g38) & (!g70) & (g104) & (g25) & (!sk[107]) & (!g66)) + ((g38) & (!g70) & (g104) & (g25) & (!sk[107]) & (g66)) + ((g38) & (g70) & (!g104) & (!g25) & (!sk[107]) & (!g66)) + ((g38) & (g70) & (!g104) & (!g25) & (!sk[107]) & (g66)) + ((g38) & (g70) & (!g104) & (!g25) & (sk[107]) & (!g66)) + ((g38) & (g70) & (!g104) & (g25) & (!sk[107]) & (!g66)) + ((g38) & (g70) & (!g104) & (g25) & (!sk[107]) & (g66)) + ((g38) & (g70) & (g104) & (!g25) & (!sk[107]) & (!g66)) + ((g38) & (g70) & (g104) & (!g25) & (!sk[107]) & (g66)) + ((g38) & (g70) & (g104) & (g25) & (!sk[107]) & (!g66)) + ((g38) & (g70) & (g104) & (g25) & (!sk[107]) & (g66)));
	assign g610 = (((!g165) & (!g579) & (!g608) & (!sk[108]) & (g609)) + ((!g165) & (!g579) & (g608) & (!sk[108]) & (g609)) + ((!g165) & (g579) & (!g608) & (!sk[108]) & (g609)) + ((!g165) & (g579) & (g608) & (!sk[108]) & (g609)) + ((g165) & (!g579) & (!g608) & (!sk[108]) & (!g609)) + ((g165) & (!g579) & (!g608) & (!sk[108]) & (g609)) + ((g165) & (!g579) & (g608) & (!sk[108]) & (!g609)) + ((g165) & (!g579) & (g608) & (!sk[108]) & (g609)) + ((g165) & (g579) & (!g608) & (!sk[108]) & (!g609)) + ((g165) & (g579) & (!g608) & (!sk[108]) & (g609)) + ((g165) & (g579) & (g608) & (!sk[108]) & (!g609)) + ((g165) & (g579) & (g608) & (!sk[108]) & (g609)) + ((g165) & (g579) & (g608) & (sk[108]) & (g609)));
	assign g611 = (((!g599) & (!g600) & (!g605) & (g606) & (!sk[109]) & (!g610)) + ((!g599) & (!g600) & (!g605) & (g606) & (!sk[109]) & (g610)) + ((!g599) & (!g600) & (g605) & (!g606) & (!sk[109]) & (!g610)) + ((!g599) & (!g600) & (g605) & (!g606) & (!sk[109]) & (g610)) + ((!g599) & (!g600) & (g605) & (g606) & (!sk[109]) & (!g610)) + ((!g599) & (!g600) & (g605) & (g606) & (!sk[109]) & (g610)) + ((!g599) & (g600) & (!g605) & (!g606) & (!sk[109]) & (!g610)) + ((!g599) & (g600) & (!g605) & (!g606) & (!sk[109]) & (g610)) + ((!g599) & (g600) & (!g605) & (g606) & (!sk[109]) & (!g610)) + ((!g599) & (g600) & (!g605) & (g606) & (!sk[109]) & (g610)) + ((!g599) & (g600) & (g605) & (!g606) & (!sk[109]) & (!g610)) + ((!g599) & (g600) & (g605) & (!g606) & (!sk[109]) & (g610)) + ((!g599) & (g600) & (g605) & (g606) & (!sk[109]) & (!g610)) + ((!g599) & (g600) & (g605) & (g606) & (!sk[109]) & (g610)) + ((g599) & (!g600) & (!g605) & (g606) & (!sk[109]) & (!g610)) + ((g599) & (!g600) & (!g605) & (g606) & (!sk[109]) & (g610)) + ((g599) & (!g600) & (g605) & (!g606) & (!sk[109]) & (!g610)) + ((g599) & (!g600) & (g605) & (!g606) & (!sk[109]) & (g610)) + ((g599) & (!g600) & (g605) & (g606) & (!sk[109]) & (!g610)) + ((g599) & (!g600) & (g605) & (g606) & (!sk[109]) & (g610)) + ((g599) & (g600) & (!g605) & (!g606) & (!sk[109]) & (!g610)) + ((g599) & (g600) & (!g605) & (!g606) & (!sk[109]) & (g610)) + ((g599) & (g600) & (!g605) & (g606) & (!sk[109]) & (!g610)) + ((g599) & (g600) & (!g605) & (g606) & (!sk[109]) & (g610)) + ((g599) & (g600) & (g605) & (!g606) & (!sk[109]) & (!g610)) + ((g599) & (g600) & (g605) & (!g606) & (!sk[109]) & (g610)) + ((g599) & (g600) & (g605) & (g606) & (!sk[109]) & (!g610)) + ((g599) & (g600) & (g605) & (g606) & (!sk[109]) & (g610)) + ((g599) & (g600) & (g605) & (g606) & (sk[109]) & (g610)));
	assign g612 = (((!g440) & (!sk[110]) & (!g441) & (!g454) & (g455) & (!g546)) + ((!g440) & (!sk[110]) & (!g441) & (!g454) & (g455) & (g546)) + ((!g440) & (!sk[110]) & (!g441) & (g454) & (!g455) & (!g546)) + ((!g440) & (!sk[110]) & (!g441) & (g454) & (!g455) & (g546)) + ((!g440) & (!sk[110]) & (!g441) & (g454) & (g455) & (!g546)) + ((!g440) & (!sk[110]) & (!g441) & (g454) & (g455) & (g546)) + ((!g440) & (!sk[110]) & (g441) & (!g454) & (!g455) & (!g546)) + ((!g440) & (!sk[110]) & (g441) & (!g454) & (!g455) & (g546)) + ((!g440) & (!sk[110]) & (g441) & (!g454) & (g455) & (!g546)) + ((!g440) & (!sk[110]) & (g441) & (!g454) & (g455) & (g546)) + ((!g440) & (!sk[110]) & (g441) & (g454) & (!g455) & (!g546)) + ((!g440) & (!sk[110]) & (g441) & (g454) & (!g455) & (g546)) + ((!g440) & (!sk[110]) & (g441) & (g454) & (g455) & (!g546)) + ((!g440) & (!sk[110]) & (g441) & (g454) & (g455) & (g546)) + ((!g440) & (sk[110]) & (!g441) & (!g454) & (!g455) & (!g546)) + ((!g440) & (sk[110]) & (!g441) & (!g454) & (!g455) & (g546)) + ((!g440) & (sk[110]) & (!g441) & (!g454) & (g455) & (g546)) + ((!g440) & (sk[110]) & (!g441) & (g454) & (!g455) & (g546)) + ((!g440) & (sk[110]) & (g441) & (!g454) & (g455) & (!g546)) + ((!g440) & (sk[110]) & (g441) & (g454) & (!g455) & (!g546)) + ((!g440) & (sk[110]) & (g441) & (g454) & (g455) & (!g546)) + ((!g440) & (sk[110]) & (g441) & (g454) & (g455) & (g546)) + ((g440) & (!sk[110]) & (!g441) & (!g454) & (g455) & (!g546)) + ((g440) & (!sk[110]) & (!g441) & (!g454) & (g455) & (g546)) + ((g440) & (!sk[110]) & (!g441) & (g454) & (!g455) & (!g546)) + ((g440) & (!sk[110]) & (!g441) & (g454) & (!g455) & (g546)) + ((g440) & (!sk[110]) & (!g441) & (g454) & (g455) & (!g546)) + ((g440) & (!sk[110]) & (!g441) & (g454) & (g455) & (g546)) + ((g440) & (!sk[110]) & (g441) & (!g454) & (!g455) & (!g546)) + ((g440) & (!sk[110]) & (g441) & (!g454) & (!g455) & (g546)) + ((g440) & (!sk[110]) & (g441) & (!g454) & (g455) & (!g546)) + ((g440) & (!sk[110]) & (g441) & (!g454) & (g455) & (g546)) + ((g440) & (!sk[110]) & (g441) & (g454) & (!g455) & (!g546)) + ((g440) & (!sk[110]) & (g441) & (g454) & (!g455) & (g546)) + ((g440) & (!sk[110]) & (g441) & (g454) & (g455) & (!g546)) + ((g440) & (!sk[110]) & (g441) & (g454) & (g455) & (g546)) + ((g440) & (sk[110]) & (!g441) & (!g454) & (g455) & (!g546)) + ((g440) & (sk[110]) & (!g441) & (g454) & (!g455) & (!g546)) + ((g440) & (sk[110]) & (!g441) & (g454) & (g455) & (!g546)) + ((g440) & (sk[110]) & (!g441) & (g454) & (g455) & (g546)) + ((g440) & (sk[110]) & (g441) & (!g454) & (!g455) & (!g546)) + ((g440) & (sk[110]) & (g441) & (!g454) & (!g455) & (g546)) + ((g440) & (sk[110]) & (g441) & (!g454) & (g455) & (g546)) + ((g440) & (sk[110]) & (g441) & (g454) & (!g455) & (g546)));
	assign g613 = (((!g70) & (!g18) & (!g154) & (!sk[111]) & (g131) & (!g587)) + ((!g70) & (!g18) & (!g154) & (!sk[111]) & (g131) & (g587)) + ((!g70) & (!g18) & (!g154) & (sk[111]) & (!g131) & (!g587)) + ((!g70) & (!g18) & (g154) & (!sk[111]) & (!g131) & (!g587)) + ((!g70) & (!g18) & (g154) & (!sk[111]) & (!g131) & (g587)) + ((!g70) & (!g18) & (g154) & (!sk[111]) & (g131) & (!g587)) + ((!g70) & (!g18) & (g154) & (!sk[111]) & (g131) & (g587)) + ((!g70) & (g18) & (!g154) & (!sk[111]) & (!g131) & (!g587)) + ((!g70) & (g18) & (!g154) & (!sk[111]) & (!g131) & (g587)) + ((!g70) & (g18) & (!g154) & (!sk[111]) & (g131) & (!g587)) + ((!g70) & (g18) & (!g154) & (!sk[111]) & (g131) & (g587)) + ((!g70) & (g18) & (!g154) & (sk[111]) & (!g131) & (!g587)) + ((!g70) & (g18) & (g154) & (!sk[111]) & (!g131) & (!g587)) + ((!g70) & (g18) & (g154) & (!sk[111]) & (!g131) & (g587)) + ((!g70) & (g18) & (g154) & (!sk[111]) & (g131) & (!g587)) + ((!g70) & (g18) & (g154) & (!sk[111]) & (g131) & (g587)) + ((g70) & (!g18) & (!g154) & (!sk[111]) & (g131) & (!g587)) + ((g70) & (!g18) & (!g154) & (!sk[111]) & (g131) & (g587)) + ((g70) & (!g18) & (!g154) & (sk[111]) & (!g131) & (!g587)) + ((g70) & (!g18) & (g154) & (!sk[111]) & (!g131) & (!g587)) + ((g70) & (!g18) & (g154) & (!sk[111]) & (!g131) & (g587)) + ((g70) & (!g18) & (g154) & (!sk[111]) & (g131) & (!g587)) + ((g70) & (!g18) & (g154) & (!sk[111]) & (g131) & (g587)) + ((g70) & (g18) & (!g154) & (!sk[111]) & (!g131) & (!g587)) + ((g70) & (g18) & (!g154) & (!sk[111]) & (!g131) & (g587)) + ((g70) & (g18) & (!g154) & (!sk[111]) & (g131) & (!g587)) + ((g70) & (g18) & (!g154) & (!sk[111]) & (g131) & (g587)) + ((g70) & (g18) & (g154) & (!sk[111]) & (!g131) & (!g587)) + ((g70) & (g18) & (g154) & (!sk[111]) & (!g131) & (g587)) + ((g70) & (g18) & (g154) & (!sk[111]) & (g131) & (!g587)) + ((g70) & (g18) & (g154) & (!sk[111]) & (g131) & (g587)));
	assign g614 = (((!g38) & (!g114) & (!g115) & (g8) & (g12) & (!g58)) + ((!g38) & (!g114) & (!g115) & (g8) & (g12) & (g58)) + ((!g38) & (g114) & (!g115) & (!g8) & (!g12) & (g58)) + ((!g38) & (g114) & (!g115) & (!g8) & (g12) & (g58)) + ((g38) & (!g114) & (!g115) & (!g8) & (!g12) & (!g58)) + ((g38) & (!g114) & (!g115) & (!g8) & (!g12) & (g58)) + ((g38) & (!g114) & (!g115) & (!g8) & (g12) & (!g58)) + ((g38) & (!g114) & (!g115) & (!g8) & (g12) & (g58)) + ((g38) & (!g114) & (!g115) & (g8) & (g12) & (!g58)) + ((g38) & (!g114) & (!g115) & (g8) & (g12) & (g58)) + ((g38) & (!g114) & (g115) & (g8) & (!g12) & (!g58)) + ((g38) & (!g114) & (g115) & (g8) & (!g12) & (g58)) + ((g38) & (!g114) & (g115) & (g8) & (g12) & (!g58)) + ((g38) & (!g114) & (g115) & (g8) & (g12) & (g58)) + ((g38) & (g114) & (!g115) & (!g8) & (!g12) & (g58)) + ((g38) & (g114) & (!g115) & (!g8) & (g12) & (g58)) + ((g38) & (g114) & (!g115) & (g8) & (!g12) & (!g58)) + ((g38) & (g114) & (!g115) & (g8) & (!g12) & (g58)) + ((g38) & (g114) & (!g115) & (g8) & (g12) & (!g58)) + ((g38) & (g114) & (!g115) & (g8) & (g12) & (g58)));
	assign g615 = (((!g297) & (!g246) & (!g360) & (g613) & (!sk[113]) & (!g614)) + ((!g297) & (!g246) & (!g360) & (g613) & (!sk[113]) & (g614)) + ((!g297) & (!g246) & (g360) & (!g613) & (!sk[113]) & (!g614)) + ((!g297) & (!g246) & (g360) & (!g613) & (!sk[113]) & (g614)) + ((!g297) & (!g246) & (g360) & (g613) & (!sk[113]) & (!g614)) + ((!g297) & (!g246) & (g360) & (g613) & (!sk[113]) & (g614)) + ((!g297) & (g246) & (!g360) & (!g613) & (!sk[113]) & (!g614)) + ((!g297) & (g246) & (!g360) & (!g613) & (!sk[113]) & (g614)) + ((!g297) & (g246) & (!g360) & (g613) & (!sk[113]) & (!g614)) + ((!g297) & (g246) & (!g360) & (g613) & (!sk[113]) & (g614)) + ((!g297) & (g246) & (!g360) & (g613) & (sk[113]) & (!g614)) + ((!g297) & (g246) & (g360) & (!g613) & (!sk[113]) & (!g614)) + ((!g297) & (g246) & (g360) & (!g613) & (!sk[113]) & (g614)) + ((!g297) & (g246) & (g360) & (g613) & (!sk[113]) & (!g614)) + ((!g297) & (g246) & (g360) & (g613) & (!sk[113]) & (g614)) + ((g297) & (!g246) & (!g360) & (g613) & (!sk[113]) & (!g614)) + ((g297) & (!g246) & (!g360) & (g613) & (!sk[113]) & (g614)) + ((g297) & (!g246) & (g360) & (!g613) & (!sk[113]) & (!g614)) + ((g297) & (!g246) & (g360) & (!g613) & (!sk[113]) & (g614)) + ((g297) & (!g246) & (g360) & (g613) & (!sk[113]) & (!g614)) + ((g297) & (!g246) & (g360) & (g613) & (!sk[113]) & (g614)) + ((g297) & (g246) & (!g360) & (!g613) & (!sk[113]) & (!g614)) + ((g297) & (g246) & (!g360) & (!g613) & (!sk[113]) & (g614)) + ((g297) & (g246) & (!g360) & (g613) & (!sk[113]) & (!g614)) + ((g297) & (g246) & (!g360) & (g613) & (!sk[113]) & (g614)) + ((g297) & (g246) & (g360) & (!g613) & (!sk[113]) & (!g614)) + ((g297) & (g246) & (g360) & (!g613) & (!sk[113]) & (g614)) + ((g297) & (g246) & (g360) & (g613) & (!sk[113]) & (!g614)) + ((g297) & (g246) & (g360) & (g613) & (!sk[113]) & (g614)));
	assign g616 = (((!g99) & (!g42) & (!sk[114]) & (!g81) & (g615)) + ((!g99) & (!g42) & (!sk[114]) & (g81) & (g615)) + ((!g99) & (!g42) & (sk[114]) & (!g81) & (g615)) + ((!g99) & (g42) & (!sk[114]) & (!g81) & (g615)) + ((!g99) & (g42) & (!sk[114]) & (g81) & (g615)) + ((!g99) & (g42) & (sk[114]) & (!g81) & (g615)) + ((g99) & (!g42) & (!sk[114]) & (!g81) & (!g615)) + ((g99) & (!g42) & (!sk[114]) & (!g81) & (g615)) + ((g99) & (!g42) & (!sk[114]) & (g81) & (!g615)) + ((g99) & (!g42) & (!sk[114]) & (g81) & (g615)) + ((g99) & (!g42) & (sk[114]) & (!g81) & (g615)) + ((g99) & (g42) & (!sk[114]) & (!g81) & (!g615)) + ((g99) & (g42) & (!sk[114]) & (!g81) & (g615)) + ((g99) & (g42) & (!sk[114]) & (g81) & (!g615)) + ((g99) & (g42) & (!sk[114]) & (g81) & (g615)));
	assign g617 = (((!g70) & (!sk[115]) & (g58) & (!g244)) + ((!g70) & (!sk[115]) & (g58) & (g244)) + ((!g70) & (sk[115]) & (!g58) & (!g244)) + ((!g70) & (sk[115]) & (g58) & (!g244)) + ((g70) & (!sk[115]) & (g58) & (!g244)) + ((g70) & (!sk[115]) & (g58) & (g244)) + ((g70) & (sk[115]) & (!g58) & (!g244)));
	assign g618 = (((!sk[116]) & (!g70) & (g593) & (!g27)) + ((!sk[116]) & (!g70) & (g593) & (g27)) + ((!sk[116]) & (g70) & (g593) & (!g27)) + ((!sk[116]) & (g70) & (g593) & (g27)) + ((sk[116]) & (!g70) & (!g593) & (!g27)) + ((sk[116]) & (!g70) & (!g593) & (g27)) + ((sk[116]) & (g70) & (!g593) & (!g27)));
	assign g619 = (((!g43) & (!g236) & (!g617) & (!sk[117]) & (g618)) + ((!g43) & (!g236) & (g617) & (!sk[117]) & (g618)) + ((!g43) & (!g236) & (g617) & (sk[117]) & (g618)) + ((!g43) & (g236) & (!g617) & (!sk[117]) & (g618)) + ((!g43) & (g236) & (g617) & (!sk[117]) & (g618)) + ((g43) & (!g236) & (!g617) & (!sk[117]) & (!g618)) + ((g43) & (!g236) & (!g617) & (!sk[117]) & (g618)) + ((g43) & (!g236) & (g617) & (!sk[117]) & (!g618)) + ((g43) & (!g236) & (g617) & (!sk[117]) & (g618)) + ((g43) & (g236) & (!g617) & (!sk[117]) & (!g618)) + ((g43) & (g236) & (!g617) & (!sk[117]) & (g618)) + ((g43) & (g236) & (g617) & (!sk[117]) & (!g618)) + ((g43) & (g236) & (g617) & (!sk[117]) & (g618)));
	assign g620 = (((!g127) & (!g93) & (!g77) & (g140) & (!sk[118]) & (!g619)) + ((!g127) & (!g93) & (!g77) & (g140) & (!sk[118]) & (g619)) + ((!g127) & (!g93) & (g77) & (!g140) & (!sk[118]) & (!g619)) + ((!g127) & (!g93) & (g77) & (!g140) & (!sk[118]) & (g619)) + ((!g127) & (!g93) & (g77) & (g140) & (!sk[118]) & (!g619)) + ((!g127) & (!g93) & (g77) & (g140) & (!sk[118]) & (g619)) + ((!g127) & (!g93) & (g77) & (g140) & (sk[118]) & (g619)) + ((!g127) & (g93) & (!g77) & (!g140) & (!sk[118]) & (!g619)) + ((!g127) & (g93) & (!g77) & (!g140) & (!sk[118]) & (g619)) + ((!g127) & (g93) & (!g77) & (g140) & (!sk[118]) & (!g619)) + ((!g127) & (g93) & (!g77) & (g140) & (!sk[118]) & (g619)) + ((!g127) & (g93) & (g77) & (!g140) & (!sk[118]) & (!g619)) + ((!g127) & (g93) & (g77) & (!g140) & (!sk[118]) & (g619)) + ((!g127) & (g93) & (g77) & (g140) & (!sk[118]) & (!g619)) + ((!g127) & (g93) & (g77) & (g140) & (!sk[118]) & (g619)) + ((g127) & (!g93) & (!g77) & (g140) & (!sk[118]) & (!g619)) + ((g127) & (!g93) & (!g77) & (g140) & (!sk[118]) & (g619)) + ((g127) & (!g93) & (g77) & (!g140) & (!sk[118]) & (!g619)) + ((g127) & (!g93) & (g77) & (!g140) & (!sk[118]) & (g619)) + ((g127) & (!g93) & (g77) & (g140) & (!sk[118]) & (!g619)) + ((g127) & (!g93) & (g77) & (g140) & (!sk[118]) & (g619)) + ((g127) & (g93) & (!g77) & (!g140) & (!sk[118]) & (!g619)) + ((g127) & (g93) & (!g77) & (!g140) & (!sk[118]) & (g619)) + ((g127) & (g93) & (!g77) & (g140) & (!sk[118]) & (!g619)) + ((g127) & (g93) & (!g77) & (g140) & (!sk[118]) & (g619)) + ((g127) & (g93) & (g77) & (!g140) & (!sk[118]) & (!g619)) + ((g127) & (g93) & (g77) & (!g140) & (!sk[118]) & (g619)) + ((g127) & (g93) & (g77) & (g140) & (!sk[118]) & (!g619)) + ((g127) & (g93) & (g77) & (g140) & (!sk[118]) & (g619)));
	assign g621 = (((!sk[119]) & (!g71) & (g32) & (!g187)) + ((!sk[119]) & (!g71) & (g32) & (g187)) + ((!sk[119]) & (g71) & (g32) & (!g187)) + ((!sk[119]) & (g71) & (g32) & (g187)) + ((sk[119]) & (!g71) & (!g32) & (!g187)) + ((sk[119]) & (!g71) & (g32) & (!g187)) + ((sk[119]) & (g71) & (!g32) & (!g187)));
	assign g622 = (((!sk[120]) & (!g38) & (g16) & (!g171)) + ((!sk[120]) & (!g38) & (g16) & (g171)) + ((!sk[120]) & (g38) & (g16) & (!g171)) + ((!sk[120]) & (g38) & (g16) & (g171)) + ((sk[120]) & (!g38) & (!g16) & (!g171)) + ((sk[120]) & (!g38) & (g16) & (!g171)) + ((sk[120]) & (g38) & (!g16) & (!g171)));
	assign g623 = (((!g54) & (g621) & (!g233) & (!g51) & (!g36) & (g622)));
	assign g624 = (((!g9) & (!g70) & (!g16) & (!g17) & (sk[122]) & (!g42)) + ((!g9) & (!g70) & (!g16) & (!g17) & (sk[122]) & (g42)) + ((!g9) & (!g70) & (!g16) & (g17) & (!sk[122]) & (!g42)) + ((!g9) & (!g70) & (!g16) & (g17) & (!sk[122]) & (g42)) + ((!g9) & (!g70) & (!g16) & (g17) & (sk[122]) & (!g42)) + ((!g9) & (!g70) & (!g16) & (g17) & (sk[122]) & (g42)) + ((!g9) & (!g70) & (g16) & (!g17) & (!sk[122]) & (!g42)) + ((!g9) & (!g70) & (g16) & (!g17) & (!sk[122]) & (g42)) + ((!g9) & (!g70) & (g16) & (!g17) & (sk[122]) & (!g42)) + ((!g9) & (!g70) & (g16) & (g17) & (!sk[122]) & (!g42)) + ((!g9) & (!g70) & (g16) & (g17) & (!sk[122]) & (g42)) + ((!g9) & (!g70) & (g16) & (g17) & (sk[122]) & (!g42)) + ((!g9) & (g70) & (!g16) & (!g17) & (!sk[122]) & (!g42)) + ((!g9) & (g70) & (!g16) & (!g17) & (!sk[122]) & (g42)) + ((!g9) & (g70) & (!g16) & (!g17) & (sk[122]) & (!g42)) + ((!g9) & (g70) & (!g16) & (!g17) & (sk[122]) & (g42)) + ((!g9) & (g70) & (!g16) & (g17) & (!sk[122]) & (!g42)) + ((!g9) & (g70) & (!g16) & (g17) & (!sk[122]) & (g42)) + ((!g9) & (g70) & (g16) & (!g17) & (!sk[122]) & (!g42)) + ((!g9) & (g70) & (g16) & (!g17) & (!sk[122]) & (g42)) + ((!g9) & (g70) & (g16) & (!g17) & (sk[122]) & (!g42)) + ((!g9) & (g70) & (g16) & (g17) & (!sk[122]) & (!g42)) + ((!g9) & (g70) & (g16) & (g17) & (!sk[122]) & (g42)) + ((g9) & (!g70) & (!g16) & (!g17) & (sk[122]) & (!g42)) + ((g9) & (!g70) & (!g16) & (g17) & (!sk[122]) & (!g42)) + ((g9) & (!g70) & (!g16) & (g17) & (!sk[122]) & (g42)) + ((g9) & (!g70) & (!g16) & (g17) & (sk[122]) & (!g42)) + ((g9) & (!g70) & (g16) & (!g17) & (!sk[122]) & (!g42)) + ((g9) & (!g70) & (g16) & (!g17) & (!sk[122]) & (g42)) + ((g9) & (!g70) & (g16) & (!g17) & (sk[122]) & (!g42)) + ((g9) & (!g70) & (g16) & (g17) & (!sk[122]) & (!g42)) + ((g9) & (!g70) & (g16) & (g17) & (!sk[122]) & (g42)) + ((g9) & (!g70) & (g16) & (g17) & (sk[122]) & (!g42)) + ((g9) & (g70) & (!g16) & (!g17) & (!sk[122]) & (!g42)) + ((g9) & (g70) & (!g16) & (!g17) & (!sk[122]) & (g42)) + ((g9) & (g70) & (!g16) & (!g17) & (sk[122]) & (!g42)) + ((g9) & (g70) & (!g16) & (g17) & (!sk[122]) & (!g42)) + ((g9) & (g70) & (!g16) & (g17) & (!sk[122]) & (g42)) + ((g9) & (g70) & (g16) & (!g17) & (!sk[122]) & (!g42)) + ((g9) & (g70) & (g16) & (!g17) & (!sk[122]) & (g42)) + ((g9) & (g70) & (g16) & (!g17) & (sk[122]) & (!g42)) + ((g9) & (g70) & (g16) & (g17) & (!sk[122]) & (!g42)) + ((g9) & (g70) & (g16) & (g17) & (!sk[122]) & (g42)));
	assign g625 = (((!g184) & (!sk[123]) & (!g50) & (!g86) & (g207) & (!g624)) + ((!g184) & (!sk[123]) & (!g50) & (!g86) & (g207) & (g624)) + ((!g184) & (!sk[123]) & (!g50) & (g86) & (!g207) & (!g624)) + ((!g184) & (!sk[123]) & (!g50) & (g86) & (!g207) & (g624)) + ((!g184) & (!sk[123]) & (!g50) & (g86) & (g207) & (!g624)) + ((!g184) & (!sk[123]) & (!g50) & (g86) & (g207) & (g624)) + ((!g184) & (!sk[123]) & (g50) & (!g86) & (!g207) & (!g624)) + ((!g184) & (!sk[123]) & (g50) & (!g86) & (!g207) & (g624)) + ((!g184) & (!sk[123]) & (g50) & (!g86) & (g207) & (!g624)) + ((!g184) & (!sk[123]) & (g50) & (!g86) & (g207) & (g624)) + ((!g184) & (!sk[123]) & (g50) & (g86) & (!g207) & (!g624)) + ((!g184) & (!sk[123]) & (g50) & (g86) & (!g207) & (g624)) + ((!g184) & (!sk[123]) & (g50) & (g86) & (g207) & (!g624)) + ((!g184) & (!sk[123]) & (g50) & (g86) & (g207) & (g624)) + ((!g184) & (sk[123]) & (!g50) & (!g86) & (!g207) & (g624)) + ((g184) & (!sk[123]) & (!g50) & (!g86) & (g207) & (!g624)) + ((g184) & (!sk[123]) & (!g50) & (!g86) & (g207) & (g624)) + ((g184) & (!sk[123]) & (!g50) & (g86) & (!g207) & (!g624)) + ((g184) & (!sk[123]) & (!g50) & (g86) & (!g207) & (g624)) + ((g184) & (!sk[123]) & (!g50) & (g86) & (g207) & (!g624)) + ((g184) & (!sk[123]) & (!g50) & (g86) & (g207) & (g624)) + ((g184) & (!sk[123]) & (g50) & (!g86) & (!g207) & (!g624)) + ((g184) & (!sk[123]) & (g50) & (!g86) & (!g207) & (g624)) + ((g184) & (!sk[123]) & (g50) & (!g86) & (g207) & (!g624)) + ((g184) & (!sk[123]) & (g50) & (!g86) & (g207) & (g624)) + ((g184) & (!sk[123]) & (g50) & (g86) & (!g207) & (!g624)) + ((g184) & (!sk[123]) & (g50) & (g86) & (!g207) & (g624)) + ((g184) & (!sk[123]) & (g50) & (g86) & (g207) & (!g624)) + ((g184) & (!sk[123]) & (g50) & (g86) & (g207) & (g624)));
	assign g626 = (((!g72) & (!sk[124]) & (!g616) & (!g620) & (g623) & (!g625)) + ((!g72) & (!sk[124]) & (!g616) & (!g620) & (g623) & (g625)) + ((!g72) & (!sk[124]) & (!g616) & (g620) & (!g623) & (!g625)) + ((!g72) & (!sk[124]) & (!g616) & (g620) & (!g623) & (g625)) + ((!g72) & (!sk[124]) & (!g616) & (g620) & (g623) & (!g625)) + ((!g72) & (!sk[124]) & (!g616) & (g620) & (g623) & (g625)) + ((!g72) & (!sk[124]) & (g616) & (!g620) & (!g623) & (!g625)) + ((!g72) & (!sk[124]) & (g616) & (!g620) & (!g623) & (g625)) + ((!g72) & (!sk[124]) & (g616) & (!g620) & (g623) & (!g625)) + ((!g72) & (!sk[124]) & (g616) & (!g620) & (g623) & (g625)) + ((!g72) & (!sk[124]) & (g616) & (g620) & (!g623) & (!g625)) + ((!g72) & (!sk[124]) & (g616) & (g620) & (!g623) & (g625)) + ((!g72) & (!sk[124]) & (g616) & (g620) & (g623) & (!g625)) + ((!g72) & (!sk[124]) & (g616) & (g620) & (g623) & (g625)) + ((!g72) & (sk[124]) & (g616) & (g620) & (g623) & (g625)) + ((g72) & (!sk[124]) & (!g616) & (!g620) & (g623) & (!g625)) + ((g72) & (!sk[124]) & (!g616) & (!g620) & (g623) & (g625)) + ((g72) & (!sk[124]) & (!g616) & (g620) & (!g623) & (!g625)) + ((g72) & (!sk[124]) & (!g616) & (g620) & (!g623) & (g625)) + ((g72) & (!sk[124]) & (!g616) & (g620) & (g623) & (!g625)) + ((g72) & (!sk[124]) & (!g616) & (g620) & (g623) & (g625)) + ((g72) & (!sk[124]) & (g616) & (!g620) & (!g623) & (!g625)) + ((g72) & (!sk[124]) & (g616) & (!g620) & (!g623) & (g625)) + ((g72) & (!sk[124]) & (g616) & (!g620) & (g623) & (!g625)) + ((g72) & (!sk[124]) & (g616) & (!g620) & (g623) & (g625)) + ((g72) & (!sk[124]) & (g616) & (g620) & (!g623) & (!g625)) + ((g72) & (!sk[124]) & (g616) & (g620) & (!g623) & (g625)) + ((g72) & (!sk[124]) & (g616) & (g620) & (g623) & (!g625)) + ((g72) & (!sk[124]) & (g616) & (g620) & (g623) & (g625)));
	assign g627 = (((!g437) & (!g438) & (!g439) & (!g451) & (!g452) & (!g453)) + ((!g437) & (!g438) & (!g439) & (!g451) & (!g452) & (g453)) + ((!g437) & (!g438) & (!g439) & (!g451) & (g452) & (!g453)) + ((!g437) & (!g438) & (!g439) & (g451) & (!g452) & (!g453)) + ((!g437) & (!g438) & (g439) & (!g451) & (g452) & (g453)) + ((!g437) & (!g438) & (g439) & (g451) & (!g452) & (g453)) + ((!g437) & (!g438) & (g439) & (g451) & (g452) & (!g453)) + ((!g437) & (!g438) & (g439) & (g451) & (g452) & (g453)) + ((!g437) & (g438) & (!g439) & (!g451) & (g452) & (g453)) + ((!g437) & (g438) & (!g439) & (g451) & (!g452) & (g453)) + ((!g437) & (g438) & (!g439) & (g451) & (g452) & (!g453)) + ((!g437) & (g438) & (!g439) & (g451) & (g452) & (g453)) + ((!g437) & (g438) & (g439) & (!g451) & (!g452) & (!g453)) + ((!g437) & (g438) & (g439) & (!g451) & (!g452) & (g453)) + ((!g437) & (g438) & (g439) & (!g451) & (g452) & (!g453)) + ((!g437) & (g438) & (g439) & (g451) & (!g452) & (!g453)) + ((g437) & (!g438) & (!g439) & (!g451) & (g452) & (g453)) + ((g437) & (!g438) & (!g439) & (g451) & (!g452) & (g453)) + ((g437) & (!g438) & (!g439) & (g451) & (g452) & (!g453)) + ((g437) & (!g438) & (!g439) & (g451) & (g452) & (g453)) + ((g437) & (!g438) & (g439) & (!g451) & (!g452) & (!g453)) + ((g437) & (!g438) & (g439) & (!g451) & (!g452) & (g453)) + ((g437) & (!g438) & (g439) & (!g451) & (g452) & (!g453)) + ((g437) & (!g438) & (g439) & (g451) & (!g452) & (!g453)) + ((g437) & (g438) & (!g439) & (!g451) & (!g452) & (!g453)) + ((g437) & (g438) & (!g439) & (!g451) & (!g452) & (g453)) + ((g437) & (g438) & (!g439) & (!g451) & (g452) & (!g453)) + ((g437) & (g438) & (!g439) & (g451) & (!g452) & (!g453)) + ((g437) & (g438) & (g439) & (!g451) & (g452) & (g453)) + ((g437) & (g438) & (g439) & (g451) & (!g452) & (g453)) + ((g437) & (g438) & (g439) & (g451) & (g452) & (!g453)) + ((g437) & (g438) & (g439) & (g451) & (g452) & (g453)));
	assign g628 = (((!g78) & (!g71) & (sk[126]) & (!g32)) + ((!g78) & (!g71) & (sk[126]) & (g32)) + ((!g78) & (g71) & (!sk[126]) & (!g32)) + ((!g78) & (g71) & (!sk[126]) & (g32)) + ((!g78) & (g71) & (sk[126]) & (!g32)) + ((g78) & (g71) & (!sk[126]) & (!g32)) + ((g78) & (g71) & (!sk[126]) & (g32)));
	assign g629 = (((!g104) & (!g27) & (sk[127]) & (g107)) + ((!g104) & (g27) & (!sk[127]) & (!g107)) + ((!g104) & (g27) & (!sk[127]) & (g107)) + ((!g104) & (g27) & (sk[127]) & (g107)) + ((g104) & (!g27) & (sk[127]) & (g107)) + ((g104) & (g27) & (!sk[127]) & (!g107)) + ((g104) & (g27) & (!sk[127]) & (g107)));
	assign g630 = (((!g26) & (sk[0]) & (!g141)) + ((g26) & (!sk[0]) & (g141)));
	assign g631 = (((!sk[1]) & (g354) & (g51)) + ((sk[1]) & (!g354) & (!g51)));
	assign g632 = (((!g114) & (!g115) & (!g8) & (g12) & (!g20) & (!g234)) + ((!g114) & (!g115) & (!g8) & (g12) & (!g20) & (g234)) + ((!g114) & (!g115) & (!g8) & (g12) & (g20) & (!g234)) + ((!g114) & (!g115) & (!g8) & (g12) & (g20) & (g234)) + ((!g114) & (!g115) & (g8) & (g12) & (!g20) & (!g234)) + ((!g114) & (!g115) & (g8) & (g12) & (!g20) & (g234)) + ((!g114) & (!g115) & (g8) & (g12) & (g20) & (!g234)) + ((!g114) & (!g115) & (g8) & (g12) & (g20) & (g234)) + ((!g114) & (g115) & (!g8) & (!g12) & (g20) & (!g234)) + ((!g114) & (g115) & (!g8) & (!g12) & (g20) & (g234)) + ((!g114) & (g115) & (!g8) & (g12) & (g20) & (!g234)) + ((!g114) & (g115) & (!g8) & (g12) & (g20) & (g234)) + ((g114) & (g115) & (g8) & (!g12) & (!g20) & (g234)) + ((g114) & (g115) & (g8) & (!g12) & (g20) & (g234)) + ((g114) & (g115) & (g8) & (g12) & (!g20) & (g234)) + ((g114) & (g115) & (g8) & (g12) & (g20) & (g234)));
	assign g633 = (((!g62) & (!g40) & (!sk[3]) & (!g27) & (g632)) + ((!g62) & (!g40) & (!sk[3]) & (g27) & (g632)) + ((!g62) & (!g40) & (sk[3]) & (!g27) & (!g632)) + ((!g62) & (!g40) & (sk[3]) & (g27) & (!g632)) + ((!g62) & (g40) & (!sk[3]) & (!g27) & (g632)) + ((!g62) & (g40) & (!sk[3]) & (g27) & (g632)) + ((!g62) & (g40) & (sk[3]) & (!g27) & (!g632)) + ((!g62) & (g40) & (sk[3]) & (g27) & (!g632)) + ((g62) & (!g40) & (!sk[3]) & (!g27) & (!g632)) + ((g62) & (!g40) & (!sk[3]) & (!g27) & (g632)) + ((g62) & (!g40) & (!sk[3]) & (g27) & (!g632)) + ((g62) & (!g40) & (!sk[3]) & (g27) & (g632)) + ((g62) & (!g40) & (sk[3]) & (!g27) & (!g632)) + ((g62) & (g40) & (!sk[3]) & (!g27) & (!g632)) + ((g62) & (g40) & (!sk[3]) & (!g27) & (g632)) + ((g62) & (g40) & (!sk[3]) & (g27) & (!g632)) + ((g62) & (g40) & (!sk[3]) & (g27) & (g632)));
	assign g634 = (((!g127) & (!sk[4]) & (!g15) & (!g152) & (g631) & (!g633)) + ((!g127) & (!sk[4]) & (!g15) & (!g152) & (g631) & (g633)) + ((!g127) & (!sk[4]) & (!g15) & (g152) & (!g631) & (!g633)) + ((!g127) & (!sk[4]) & (!g15) & (g152) & (!g631) & (g633)) + ((!g127) & (!sk[4]) & (!g15) & (g152) & (g631) & (!g633)) + ((!g127) & (!sk[4]) & (!g15) & (g152) & (g631) & (g633)) + ((!g127) & (!sk[4]) & (g15) & (!g152) & (!g631) & (!g633)) + ((!g127) & (!sk[4]) & (g15) & (!g152) & (!g631) & (g633)) + ((!g127) & (!sk[4]) & (g15) & (!g152) & (g631) & (!g633)) + ((!g127) & (!sk[4]) & (g15) & (!g152) & (g631) & (g633)) + ((!g127) & (!sk[4]) & (g15) & (g152) & (!g631) & (!g633)) + ((!g127) & (!sk[4]) & (g15) & (g152) & (!g631) & (g633)) + ((!g127) & (!sk[4]) & (g15) & (g152) & (g631) & (!g633)) + ((!g127) & (!sk[4]) & (g15) & (g152) & (g631) & (g633)) + ((!g127) & (sk[4]) & (g15) & (!g152) & (g631) & (g633)) + ((g127) & (!sk[4]) & (!g15) & (!g152) & (g631) & (!g633)) + ((g127) & (!sk[4]) & (!g15) & (!g152) & (g631) & (g633)) + ((g127) & (!sk[4]) & (!g15) & (g152) & (!g631) & (!g633)) + ((g127) & (!sk[4]) & (!g15) & (g152) & (!g631) & (g633)) + ((g127) & (!sk[4]) & (!g15) & (g152) & (g631) & (!g633)) + ((g127) & (!sk[4]) & (!g15) & (g152) & (g631) & (g633)) + ((g127) & (!sk[4]) & (g15) & (!g152) & (!g631) & (!g633)) + ((g127) & (!sk[4]) & (g15) & (!g152) & (!g631) & (g633)) + ((g127) & (!sk[4]) & (g15) & (!g152) & (g631) & (!g633)) + ((g127) & (!sk[4]) & (g15) & (!g152) & (g631) & (g633)) + ((g127) & (!sk[4]) & (g15) & (g152) & (!g631) & (!g633)) + ((g127) & (!sk[4]) & (g15) & (g152) & (!g631) & (g633)) + ((g127) & (!sk[4]) & (g15) & (g152) & (g631) & (!g633)) + ((g127) & (!sk[4]) & (g15) & (g152) & (g631) & (g633)));
	assign g635 = (((!sk[5]) & (!g29) & (g60) & (!g154)) + ((!sk[5]) & (!g29) & (g60) & (g154)) + ((!sk[5]) & (g29) & (g60) & (!g154)) + ((!sk[5]) & (g29) & (g60) & (g154)) + ((sk[5]) & (!g29) & (!g60) & (!g154)));
	assign g636 = (((!g70) & (!g25) & (sk[6]) & (!g124)) + ((!g70) & (g25) & (!sk[6]) & (!g124)) + ((!g70) & (g25) & (!sk[6]) & (g124)) + ((!g70) & (g25) & (sk[6]) & (!g124)) + ((g70) & (!g25) & (sk[6]) & (!g124)) + ((g70) & (g25) & (!sk[6]) & (!g124)) + ((g70) & (g25) & (!sk[6]) & (g124)));
	assign g637 = (((!g38) & (!g9) & (!g71) & (!g40) & (!g20) & (!g43)) + ((!g38) & (!g9) & (!g71) & (!g40) & (g20) & (!g43)) + ((!g38) & (!g9) & (!g71) & (g40) & (!g20) & (!g43)) + ((!g38) & (!g9) & (!g71) & (g40) & (g20) & (!g43)) + ((!g38) & (!g9) & (g71) & (!g40) & (!g20) & (!g43)) + ((!g38) & (!g9) & (g71) & (g40) & (!g20) & (!g43)) + ((!g38) & (g9) & (!g71) & (!g40) & (!g20) & (!g43)) + ((!g38) & (g9) & (!g71) & (!g40) & (g20) & (!g43)) + ((!g38) & (g9) & (g71) & (!g40) & (!g20) & (!g43)) + ((g38) & (!g9) & (!g71) & (!g40) & (!g20) & (!g43)) + ((g38) & (!g9) & (!g71) & (!g40) & (g20) & (!g43)) + ((g38) & (!g9) & (!g71) & (g40) & (!g20) & (!g43)) + ((g38) & (!g9) & (!g71) & (g40) & (g20) & (!g43)) + ((g38) & (g9) & (!g71) & (!g40) & (!g20) & (!g43)) + ((g38) & (g9) & (!g71) & (!g40) & (g20) & (!g43)));
	assign g638 = (((!g185) & (!g236) & (sk[8]) & (!g210)) + ((!g185) & (g236) & (!sk[8]) & (!g210)) + ((!g185) & (g236) & (!sk[8]) & (g210)) + ((g185) & (g236) & (!sk[8]) & (!g210)) + ((g185) & (g236) & (!sk[8]) & (g210)));
	assign g639 = (((!sk[9]) & (!g635) & (!g276) & (!g636) & (g637) & (!g638)) + ((!sk[9]) & (!g635) & (!g276) & (!g636) & (g637) & (g638)) + ((!sk[9]) & (!g635) & (!g276) & (g636) & (!g637) & (!g638)) + ((!sk[9]) & (!g635) & (!g276) & (g636) & (!g637) & (g638)) + ((!sk[9]) & (!g635) & (!g276) & (g636) & (g637) & (!g638)) + ((!sk[9]) & (!g635) & (!g276) & (g636) & (g637) & (g638)) + ((!sk[9]) & (!g635) & (g276) & (!g636) & (!g637) & (!g638)) + ((!sk[9]) & (!g635) & (g276) & (!g636) & (!g637) & (g638)) + ((!sk[9]) & (!g635) & (g276) & (!g636) & (g637) & (!g638)) + ((!sk[9]) & (!g635) & (g276) & (!g636) & (g637) & (g638)) + ((!sk[9]) & (!g635) & (g276) & (g636) & (!g637) & (!g638)) + ((!sk[9]) & (!g635) & (g276) & (g636) & (!g637) & (g638)) + ((!sk[9]) & (!g635) & (g276) & (g636) & (g637) & (!g638)) + ((!sk[9]) & (!g635) & (g276) & (g636) & (g637) & (g638)) + ((!sk[9]) & (g635) & (!g276) & (!g636) & (g637) & (!g638)) + ((!sk[9]) & (g635) & (!g276) & (!g636) & (g637) & (g638)) + ((!sk[9]) & (g635) & (!g276) & (g636) & (!g637) & (!g638)) + ((!sk[9]) & (g635) & (!g276) & (g636) & (!g637) & (g638)) + ((!sk[9]) & (g635) & (!g276) & (g636) & (g637) & (!g638)) + ((!sk[9]) & (g635) & (!g276) & (g636) & (g637) & (g638)) + ((!sk[9]) & (g635) & (g276) & (!g636) & (!g637) & (!g638)) + ((!sk[9]) & (g635) & (g276) & (!g636) & (!g637) & (g638)) + ((!sk[9]) & (g635) & (g276) & (!g636) & (g637) & (!g638)) + ((!sk[9]) & (g635) & (g276) & (!g636) & (g637) & (g638)) + ((!sk[9]) & (g635) & (g276) & (g636) & (!g637) & (!g638)) + ((!sk[9]) & (g635) & (g276) & (g636) & (!g637) & (g638)) + ((!sk[9]) & (g635) & (g276) & (g636) & (g637) & (!g638)) + ((!sk[9]) & (g635) & (g276) & (g636) & (g637) & (g638)) + ((sk[9]) & (g635) & (g276) & (g636) & (g637) & (g638)));
	assign g640 = (((!g129) & (g628) & (g629) & (g630) & (g634) & (g639)));
	assign g641 = (((!g463) & (!g464) & (!g477) & (!g478) & (!g489) & (!g545)) + ((!g463) & (!g464) & (!g477) & (!g478) & (!g489) & (g545)) + ((!g463) & (!g464) & (!g477) & (!g478) & (g489) & (!g545)) + ((!g463) & (!g464) & (!g477) & (!g478) & (g489) & (g545)) + ((!g463) & (!g464) & (!g477) & (g478) & (!g489) & (!g545)) + ((!g463) & (!g464) & (g477) & (!g478) & (!g489) & (!g545)) + ((!g463) & (g464) & (!g477) & (g478) & (!g489) & (g545)) + ((!g463) & (g464) & (!g477) & (g478) & (g489) & (!g545)) + ((!g463) & (g464) & (!g477) & (g478) & (g489) & (g545)) + ((!g463) & (g464) & (g477) & (!g478) & (!g489) & (g545)) + ((!g463) & (g464) & (g477) & (!g478) & (g489) & (!g545)) + ((!g463) & (g464) & (g477) & (!g478) & (g489) & (g545)) + ((!g463) & (g464) & (g477) & (g478) & (!g489) & (!g545)) + ((!g463) & (g464) & (g477) & (g478) & (!g489) & (g545)) + ((!g463) & (g464) & (g477) & (g478) & (g489) & (!g545)) + ((!g463) & (g464) & (g477) & (g478) & (g489) & (g545)) + ((g463) & (!g464) & (!g477) & (g478) & (!g489) & (g545)) + ((g463) & (!g464) & (!g477) & (g478) & (g489) & (!g545)) + ((g463) & (!g464) & (!g477) & (g478) & (g489) & (g545)) + ((g463) & (!g464) & (g477) & (!g478) & (!g489) & (g545)) + ((g463) & (!g464) & (g477) & (!g478) & (g489) & (!g545)) + ((g463) & (!g464) & (g477) & (!g478) & (g489) & (g545)) + ((g463) & (!g464) & (g477) & (g478) & (!g489) & (!g545)) + ((g463) & (!g464) & (g477) & (g478) & (!g489) & (g545)) + ((g463) & (!g464) & (g477) & (g478) & (g489) & (!g545)) + ((g463) & (!g464) & (g477) & (g478) & (g489) & (g545)) + ((g463) & (g464) & (!g477) & (!g478) & (!g489) & (!g545)) + ((g463) & (g464) & (!g477) & (!g478) & (!g489) & (g545)) + ((g463) & (g464) & (!g477) & (!g478) & (g489) & (!g545)) + ((g463) & (g464) & (!g477) & (!g478) & (g489) & (g545)) + ((g463) & (g464) & (!g477) & (g478) & (!g489) & (!g545)) + ((g463) & (g464) & (g477) & (!g478) & (!g489) & (!g545)));
	assign g642 = (((!sk[12]) & (g104) & (g149)) + ((sk[12]) & (g104) & (g149)));
	assign g643 = (((!g70) & (!g99) & (!g30) & (!g25) & (!g41) & (!g642)) + ((!g70) & (!g99) & (!g30) & (!g25) & (g41) & (!g642)) + ((!g70) & (!g99) & (!g30) & (g25) & (!g41) & (!g642)) + ((!g70) & (!g99) & (!g30) & (g25) & (g41) & (!g642)) + ((!g70) & (!g99) & (g30) & (!g25) & (!g41) & (!g642)) + ((!g70) & (!g99) & (g30) & (!g25) & (g41) & (!g642)) + ((!g70) & (!g99) & (g30) & (g25) & (!g41) & (!g642)) + ((!g70) & (!g99) & (g30) & (g25) & (g41) & (!g642)) + ((!g70) & (g99) & (!g30) & (!g25) & (!g41) & (!g642)) + ((!g70) & (g99) & (g30) & (!g25) & (!g41) & (!g642)) + ((g70) & (!g99) & (!g30) & (!g25) & (!g41) & (!g642)) + ((g70) & (!g99) & (!g30) & (!g25) & (g41) & (!g642)) + ((g70) & (!g99) & (!g30) & (g25) & (!g41) & (!g642)) + ((g70) & (!g99) & (!g30) & (g25) & (g41) & (!g642)) + ((g70) & (g99) & (!g30) & (!g25) & (!g41) & (!g642)));
	assign g644 = (((!g38) & (!g30) & (!sk[14]) & (!g104) & (g272)) + ((!g38) & (!g30) & (!sk[14]) & (g104) & (g272)) + ((!g38) & (!g30) & (sk[14]) & (!g104) & (!g272)) + ((!g38) & (!g30) & (sk[14]) & (g104) & (!g272)) + ((!g38) & (g30) & (!sk[14]) & (!g104) & (g272)) + ((!g38) & (g30) & (!sk[14]) & (g104) & (g272)) + ((!g38) & (g30) & (sk[14]) & (!g104) & (!g272)) + ((g38) & (!g30) & (!sk[14]) & (!g104) & (!g272)) + ((g38) & (!g30) & (!sk[14]) & (!g104) & (g272)) + ((g38) & (!g30) & (!sk[14]) & (g104) & (!g272)) + ((g38) & (!g30) & (!sk[14]) & (g104) & (g272)) + ((g38) & (!g30) & (sk[14]) & (!g104) & (!g272)) + ((g38) & (g30) & (!sk[14]) & (!g104) & (!g272)) + ((g38) & (g30) & (!sk[14]) & (!g104) & (g272)) + ((g38) & (g30) & (!sk[14]) & (g104) & (!g272)) + ((g38) & (g30) & (!sk[14]) & (g104) & (g272)) + ((g38) & (g30) & (sk[14]) & (!g104) & (!g272)));
	assign g645 = (((!g70) & (!sk[15]) & (!g12) & (!g244) & (g155)) + ((!g70) & (!sk[15]) & (!g12) & (g244) & (g155)) + ((!g70) & (!sk[15]) & (g12) & (!g244) & (g155)) + ((!g70) & (!sk[15]) & (g12) & (g244) & (g155)) + ((!g70) & (sk[15]) & (!g12) & (!g244) & (!g155)) + ((!g70) & (sk[15]) & (!g12) & (!g244) & (g155)) + ((!g70) & (sk[15]) & (g12) & (!g244) & (!g155)) + ((!g70) & (sk[15]) & (g12) & (!g244) & (g155)) + ((g70) & (!sk[15]) & (!g12) & (!g244) & (!g155)) + ((g70) & (!sk[15]) & (!g12) & (!g244) & (g155)) + ((g70) & (!sk[15]) & (!g12) & (g244) & (!g155)) + ((g70) & (!sk[15]) & (!g12) & (g244) & (g155)) + ((g70) & (!sk[15]) & (g12) & (!g244) & (!g155)) + ((g70) & (!sk[15]) & (g12) & (!g244) & (g155)) + ((g70) & (!sk[15]) & (g12) & (g244) & (!g155)) + ((g70) & (!sk[15]) & (g12) & (g244) & (g155)) + ((g70) & (sk[15]) & (!g12) & (!g244) & (!g155)));
	assign g646 = (((!g99) & (!sk[16]) & (!g18) & (!g644) & (g645)) + ((!g99) & (!sk[16]) & (!g18) & (g644) & (g645)) + ((!g99) & (!sk[16]) & (g18) & (!g644) & (g645)) + ((!g99) & (!sk[16]) & (g18) & (g644) & (g645)) + ((!g99) & (sk[16]) & (!g18) & (g644) & (g645)) + ((!g99) & (sk[16]) & (g18) & (g644) & (g645)) + ((g99) & (!sk[16]) & (!g18) & (!g644) & (!g645)) + ((g99) & (!sk[16]) & (!g18) & (!g644) & (g645)) + ((g99) & (!sk[16]) & (!g18) & (g644) & (!g645)) + ((g99) & (!sk[16]) & (!g18) & (g644) & (g645)) + ((g99) & (!sk[16]) & (g18) & (!g644) & (!g645)) + ((g99) & (!sk[16]) & (g18) & (!g644) & (g645)) + ((g99) & (!sk[16]) & (g18) & (g644) & (!g645)) + ((g99) & (!sk[16]) & (g18) & (g644) & (g645)) + ((g99) & (sk[16]) & (!g18) & (g644) & (g645)));
	assign g647 = (((!g132) & (!g583) & (!g608) & (!sk[17]) & (g643) & (!g646)) + ((!g132) & (!g583) & (!g608) & (!sk[17]) & (g643) & (g646)) + ((!g132) & (!g583) & (g608) & (!sk[17]) & (!g643) & (!g646)) + ((!g132) & (!g583) & (g608) & (!sk[17]) & (!g643) & (g646)) + ((!g132) & (!g583) & (g608) & (!sk[17]) & (g643) & (!g646)) + ((!g132) & (!g583) & (g608) & (!sk[17]) & (g643) & (g646)) + ((!g132) & (g583) & (!g608) & (!sk[17]) & (!g643) & (!g646)) + ((!g132) & (g583) & (!g608) & (!sk[17]) & (!g643) & (g646)) + ((!g132) & (g583) & (!g608) & (!sk[17]) & (g643) & (!g646)) + ((!g132) & (g583) & (!g608) & (!sk[17]) & (g643) & (g646)) + ((!g132) & (g583) & (g608) & (!sk[17]) & (!g643) & (!g646)) + ((!g132) & (g583) & (g608) & (!sk[17]) & (!g643) & (g646)) + ((!g132) & (g583) & (g608) & (!sk[17]) & (g643) & (!g646)) + ((!g132) & (g583) & (g608) & (!sk[17]) & (g643) & (g646)) + ((g132) & (!g583) & (!g608) & (!sk[17]) & (g643) & (!g646)) + ((g132) & (!g583) & (!g608) & (!sk[17]) & (g643) & (g646)) + ((g132) & (!g583) & (g608) & (!sk[17]) & (!g643) & (!g646)) + ((g132) & (!g583) & (g608) & (!sk[17]) & (!g643) & (g646)) + ((g132) & (!g583) & (g608) & (!sk[17]) & (g643) & (!g646)) + ((g132) & (!g583) & (g608) & (!sk[17]) & (g643) & (g646)) + ((g132) & (g583) & (!g608) & (!sk[17]) & (!g643) & (!g646)) + ((g132) & (g583) & (!g608) & (!sk[17]) & (!g643) & (g646)) + ((g132) & (g583) & (!g608) & (!sk[17]) & (g643) & (!g646)) + ((g132) & (g583) & (!g608) & (!sk[17]) & (g643) & (g646)) + ((g132) & (g583) & (g608) & (!sk[17]) & (!g643) & (!g646)) + ((g132) & (g583) & (g608) & (!sk[17]) & (!g643) & (g646)) + ((g132) & (g583) & (g608) & (!sk[17]) & (g643) & (!g646)) + ((g132) & (g583) & (g608) & (!sk[17]) & (g643) & (g646)) + ((g132) & (g583) & (g608) & (sk[17]) & (g643) & (g646)));
	assign g648 = (((!sk[18]) & (!g154) & (g93) & (!g647)) + ((!sk[18]) & (!g154) & (g93) & (g647)) + ((!sk[18]) & (g154) & (g93) & (!g647)) + ((!sk[18]) & (g154) & (g93) & (g647)) + ((sk[18]) & (!g154) & (!g93) & (g647)));
	assign g649 = (((g345) & (!sk[19]) & (g173)) + ((g345) & (sk[19]) & (g173)));
	assign g650 = (((!g9) & (!sk[20]) & (!g58) & (!g46) & (g66) & (!g20)) + ((!g9) & (!sk[20]) & (!g58) & (!g46) & (g66) & (g20)) + ((!g9) & (!sk[20]) & (!g58) & (g46) & (!g66) & (!g20)) + ((!g9) & (!sk[20]) & (!g58) & (g46) & (!g66) & (g20)) + ((!g9) & (!sk[20]) & (!g58) & (g46) & (g66) & (!g20)) + ((!g9) & (!sk[20]) & (!g58) & (g46) & (g66) & (g20)) + ((!g9) & (!sk[20]) & (g58) & (!g46) & (!g66) & (!g20)) + ((!g9) & (!sk[20]) & (g58) & (!g46) & (!g66) & (g20)) + ((!g9) & (!sk[20]) & (g58) & (!g46) & (g66) & (!g20)) + ((!g9) & (!sk[20]) & (g58) & (!g46) & (g66) & (g20)) + ((!g9) & (!sk[20]) & (g58) & (g46) & (!g66) & (!g20)) + ((!g9) & (!sk[20]) & (g58) & (g46) & (!g66) & (g20)) + ((!g9) & (!sk[20]) & (g58) & (g46) & (g66) & (!g20)) + ((!g9) & (!sk[20]) & (g58) & (g46) & (g66) & (g20)) + ((!g9) & (sk[20]) & (!g58) & (!g46) & (!g66) & (!g20)) + ((!g9) & (sk[20]) & (!g58) & (!g46) & (!g66) & (g20)) + ((!g9) & (sk[20]) & (!g58) & (!g46) & (g66) & (!g20)) + ((!g9) & (sk[20]) & (!g58) & (!g46) & (g66) & (g20)) + ((!g9) & (sk[20]) & (!g58) & (g46) & (!g66) & (!g20)) + ((!g9) & (sk[20]) & (!g58) & (g46) & (g66) & (!g20)) + ((!g9) & (sk[20]) & (g58) & (!g46) & (!g66) & (!g20)) + ((!g9) & (sk[20]) & (g58) & (!g46) & (!g66) & (g20)) + ((!g9) & (sk[20]) & (g58) & (!g46) & (g66) & (!g20)) + ((!g9) & (sk[20]) & (g58) & (!g46) & (g66) & (g20)) + ((g9) & (!sk[20]) & (!g58) & (!g46) & (g66) & (!g20)) + ((g9) & (!sk[20]) & (!g58) & (!g46) & (g66) & (g20)) + ((g9) & (!sk[20]) & (!g58) & (g46) & (!g66) & (!g20)) + ((g9) & (!sk[20]) & (!g58) & (g46) & (!g66) & (g20)) + ((g9) & (!sk[20]) & (!g58) & (g46) & (g66) & (!g20)) + ((g9) & (!sk[20]) & (!g58) & (g46) & (g66) & (g20)) + ((g9) & (!sk[20]) & (g58) & (!g46) & (!g66) & (!g20)) + ((g9) & (!sk[20]) & (g58) & (!g46) & (!g66) & (g20)) + ((g9) & (!sk[20]) & (g58) & (!g46) & (g66) & (!g20)) + ((g9) & (!sk[20]) & (g58) & (!g46) & (g66) & (g20)) + ((g9) & (!sk[20]) & (g58) & (g46) & (!g66) & (!g20)) + ((g9) & (!sk[20]) & (g58) & (g46) & (!g66) & (g20)) + ((g9) & (!sk[20]) & (g58) & (g46) & (g66) & (!g20)) + ((g9) & (!sk[20]) & (g58) & (g46) & (g66) & (g20)) + ((g9) & (sk[20]) & (!g58) & (!g46) & (!g66) & (!g20)) + ((g9) & (sk[20]) & (!g58) & (g46) & (!g66) & (!g20)) + ((g9) & (sk[20]) & (g58) & (!g46) & (!g66) & (!g20)));
	assign g651 = (((!g112) & (!g113) & (g97) & (g98) & (g62) & (!g71)) + ((!g112) & (!g113) & (g97) & (g98) & (g62) & (g71)) + ((!g112) & (g113) & (!g97) & (!g98) & (!g62) & (g71)) + ((!g112) & (g113) & (!g97) & (!g98) & (g62) & (g71)) + ((g112) & (!g113) & (g97) & (!g98) & (!g62) & (g71)) + ((g112) & (!g113) & (g97) & (!g98) & (g62) & (g71)) + ((g112) & (g113) & (!g97) & (g98) & (g62) & (!g71)) + ((g112) & (g113) & (!g97) & (g98) & (g62) & (g71)) + ((g112) & (g113) & (g97) & (g98) & (g62) & (!g71)) + ((g112) & (g113) & (g97) & (g98) & (g62) & (g71)));
	assign g652 = (((!g9) & (!g16) & (!sk[22]) & (!g40) & (g651)) + ((!g9) & (!g16) & (!sk[22]) & (g40) & (g651)) + ((!g9) & (!g16) & (sk[22]) & (!g40) & (!g651)) + ((!g9) & (!g16) & (sk[22]) & (g40) & (!g651)) + ((!g9) & (g16) & (!sk[22]) & (!g40) & (g651)) + ((!g9) & (g16) & (!sk[22]) & (g40) & (g651)) + ((!g9) & (g16) & (sk[22]) & (!g40) & (!g651)) + ((g9) & (!g16) & (!sk[22]) & (!g40) & (!g651)) + ((g9) & (!g16) & (!sk[22]) & (!g40) & (g651)) + ((g9) & (!g16) & (!sk[22]) & (g40) & (!g651)) + ((g9) & (!g16) & (!sk[22]) & (g40) & (g651)) + ((g9) & (!g16) & (sk[22]) & (!g40) & (!g651)) + ((g9) & (g16) & (!sk[22]) & (!g40) & (!g651)) + ((g9) & (g16) & (!sk[22]) & (!g40) & (g651)) + ((g9) & (g16) & (!sk[22]) & (g40) & (!g651)) + ((g9) & (g16) & (!sk[22]) & (g40) & (g651)) + ((g9) & (g16) & (sk[22]) & (!g40) & (!g651)));
	assign g653 = (((!sk[23]) & (!g228) & (!g335) & (!g650) & (g652)) + ((!sk[23]) & (!g228) & (!g335) & (g650) & (g652)) + ((!sk[23]) & (!g228) & (g335) & (!g650) & (g652)) + ((!sk[23]) & (!g228) & (g335) & (g650) & (g652)) + ((!sk[23]) & (g228) & (!g335) & (!g650) & (!g652)) + ((!sk[23]) & (g228) & (!g335) & (!g650) & (g652)) + ((!sk[23]) & (g228) & (!g335) & (g650) & (!g652)) + ((!sk[23]) & (g228) & (!g335) & (g650) & (g652)) + ((!sk[23]) & (g228) & (g335) & (!g650) & (!g652)) + ((!sk[23]) & (g228) & (g335) & (!g650) & (g652)) + ((!sk[23]) & (g228) & (g335) & (g650) & (!g652)) + ((!sk[23]) & (g228) & (g335) & (g650) & (g652)) + ((sk[23]) & (g228) & (g335) & (g650) & (g652)));
	assign g654 = (((!sk[24]) & (!g210) & (g96) & (!g134)) + ((!sk[24]) & (!g210) & (g96) & (g134)) + ((!sk[24]) & (g210) & (g96) & (!g134)) + ((!sk[24]) & (g210) & (g96) & (g134)) + ((sk[24]) & (!g210) & (g96) & (g134)));
	assign g655 = (((!g648) & (!sk[25]) & (!g649) & (!g653) & (g654)) + ((!g648) & (!sk[25]) & (!g649) & (g653) & (g654)) + ((!g648) & (!sk[25]) & (g649) & (!g653) & (g654)) + ((!g648) & (!sk[25]) & (g649) & (g653) & (g654)) + ((g648) & (!sk[25]) & (!g649) & (!g653) & (!g654)) + ((g648) & (!sk[25]) & (!g649) & (!g653) & (g654)) + ((g648) & (!sk[25]) & (!g649) & (g653) & (!g654)) + ((g648) & (!sk[25]) & (!g649) & (g653) & (g654)) + ((g648) & (!sk[25]) & (g649) & (!g653) & (!g654)) + ((g648) & (!sk[25]) & (g649) & (!g653) & (g654)) + ((g648) & (!sk[25]) & (g649) & (g653) & (!g654)) + ((g648) & (!sk[25]) & (g649) & (g653) & (g654)) + ((g648) & (sk[25]) & (g649) & (g653) & (g654)));
	assign g656 = (((!g460) & (!g461) & (!g462) & (!sk[26]) & (g477)) + ((!g460) & (!g461) & (!g462) & (sk[26]) & (g477)) + ((!g460) & (!g461) & (g462) & (!sk[26]) & (g477)) + ((!g460) & (!g461) & (g462) & (sk[26]) & (!g477)) + ((!g460) & (g461) & (!g462) & (!sk[26]) & (g477)) + ((!g460) & (g461) & (!g462) & (sk[26]) & (!g477)) + ((!g460) & (g461) & (g462) & (!sk[26]) & (g477)) + ((!g460) & (g461) & (g462) & (sk[26]) & (g477)) + ((g460) & (!g461) & (!g462) & (!sk[26]) & (!g477)) + ((g460) & (!g461) & (!g462) & (!sk[26]) & (g477)) + ((g460) & (!g461) & (!g462) & (sk[26]) & (!g477)) + ((g460) & (!g461) & (g462) & (!sk[26]) & (!g477)) + ((g460) & (!g461) & (g462) & (!sk[26]) & (g477)) + ((g460) & (!g461) & (g462) & (sk[26]) & (g477)) + ((g460) & (g461) & (!g462) & (!sk[26]) & (!g477)) + ((g460) & (g461) & (!g462) & (!sk[26]) & (g477)) + ((g460) & (g461) & (!g462) & (sk[26]) & (g477)) + ((g460) & (g461) & (g462) & (!sk[26]) & (!g477)) + ((g460) & (g461) & (g462) & (!sk[26]) & (g477)) + ((g460) & (g461) & (g462) & (sk[26]) & (!g477)));
	assign g657 = (((!g485) & (!sk[27]) & (g486) & (!g487)) + ((!g485) & (!sk[27]) & (g486) & (g487)) + ((!g485) & (sk[27]) & (!g486) & (!g487)) + ((g485) & (!sk[27]) & (g486) & (!g487)) + ((g485) & (!sk[27]) & (g486) & (g487)) + ((g485) & (sk[27]) & (!g486) & (!g487)) + ((g485) & (sk[27]) & (!g486) & (g487)) + ((g485) & (sk[27]) & (g486) & (!g487)));
	assign g658 = (((!g503) & (!g539) & (!g542) & (g543) & (!sk[28]) & (!g544)) + ((!g503) & (!g539) & (!g542) & (g543) & (!sk[28]) & (g544)) + ((!g503) & (!g539) & (!g542) & (g543) & (sk[28]) & (g544)) + ((!g503) & (!g539) & (g542) & (!g543) & (!sk[28]) & (!g544)) + ((!g503) & (!g539) & (g542) & (!g543) & (!sk[28]) & (g544)) + ((!g503) & (!g539) & (g542) & (!g543) & (sk[28]) & (g544)) + ((!g503) & (!g539) & (g542) & (g543) & (!sk[28]) & (!g544)) + ((!g503) & (!g539) & (g542) & (g543) & (!sk[28]) & (g544)) + ((!g503) & (!g539) & (g542) & (g543) & (sk[28]) & (!g544)) + ((!g503) & (!g539) & (g542) & (g543) & (sk[28]) & (g544)) + ((!g503) & (g539) & (!g542) & (!g543) & (!sk[28]) & (!g544)) + ((!g503) & (g539) & (!g542) & (!g543) & (!sk[28]) & (g544)) + ((!g503) & (g539) & (!g542) & (!g543) & (sk[28]) & (g544)) + ((!g503) & (g539) & (!g542) & (g543) & (!sk[28]) & (!g544)) + ((!g503) & (g539) & (!g542) & (g543) & (!sk[28]) & (g544)) + ((!g503) & (g539) & (!g542) & (g543) & (sk[28]) & (!g544)) + ((!g503) & (g539) & (!g542) & (g543) & (sk[28]) & (g544)) + ((!g503) & (g539) & (g542) & (!g543) & (!sk[28]) & (!g544)) + ((!g503) & (g539) & (g542) & (!g543) & (!sk[28]) & (g544)) + ((!g503) & (g539) & (g542) & (!g543) & (sk[28]) & (g544)) + ((!g503) & (g539) & (g542) & (g543) & (!sk[28]) & (!g544)) + ((!g503) & (g539) & (g542) & (g543) & (!sk[28]) & (g544)) + ((!g503) & (g539) & (g542) & (g543) & (sk[28]) & (!g544)) + ((!g503) & (g539) & (g542) & (g543) & (sk[28]) & (g544)) + ((g503) & (!g539) & (!g542) & (g543) & (!sk[28]) & (!g544)) + ((g503) & (!g539) & (!g542) & (g543) & (!sk[28]) & (g544)) + ((g503) & (!g539) & (!g542) & (g543) & (sk[28]) & (g544)) + ((g503) & (!g539) & (g542) & (!g543) & (!sk[28]) & (!g544)) + ((g503) & (!g539) & (g542) & (!g543) & (!sk[28]) & (g544)) + ((g503) & (!g539) & (g542) & (g543) & (!sk[28]) & (!g544)) + ((g503) & (!g539) & (g542) & (g543) & (!sk[28]) & (g544)) + ((g503) & (!g539) & (g542) & (g543) & (sk[28]) & (g544)) + ((g503) & (g539) & (!g542) & (!g543) & (!sk[28]) & (!g544)) + ((g503) & (g539) & (!g542) & (!g543) & (!sk[28]) & (g544)) + ((g503) & (g539) & (!g542) & (g543) & (!sk[28]) & (!g544)) + ((g503) & (g539) & (!g542) & (g543) & (!sk[28]) & (g544)) + ((g503) & (g539) & (!g542) & (g543) & (sk[28]) & (g544)) + ((g503) & (g539) & (g542) & (!g543) & (!sk[28]) & (!g544)) + ((g503) & (g539) & (g542) & (!g543) & (!sk[28]) & (g544)) + ((g503) & (g539) & (g542) & (!g543) & (sk[28]) & (g544)) + ((g503) & (g539) & (g542) & (g543) & (!sk[28]) & (!g544)) + ((g503) & (g539) & (g542) & (g543) & (!sk[28]) & (g544)) + ((g503) & (g539) & (g542) & (g543) & (sk[28]) & (!g544)) + ((g503) & (g539) & (g542) & (g543) & (sk[28]) & (g544)));
	assign g659 = (((!g16) & (!g12) & (sk[29]) & (!g59)) + ((!g16) & (g12) & (!sk[29]) & (!g59)) + ((!g16) & (g12) & (!sk[29]) & (g59)) + ((!g16) & (g12) & (sk[29]) & (!g59)) + ((g16) & (!g12) & (sk[29]) & (!g59)) + ((g16) & (g12) & (!sk[29]) & (!g59)) + ((g16) & (g12) & (!sk[29]) & (g59)));
	assign g660 = (((!g46) & (!sk[30]) & (!g41) & (!g19) & (g43)) + ((!g46) & (!sk[30]) & (!g41) & (g19) & (g43)) + ((!g46) & (!sk[30]) & (g41) & (!g19) & (g43)) + ((!g46) & (!sk[30]) & (g41) & (g19) & (g43)) + ((!g46) & (sk[30]) & (!g41) & (!g19) & (!g43)) + ((!g46) & (sk[30]) & (g41) & (!g19) & (!g43)) + ((g46) & (!sk[30]) & (!g41) & (!g19) & (!g43)) + ((g46) & (!sk[30]) & (!g41) & (!g19) & (g43)) + ((g46) & (!sk[30]) & (!g41) & (g19) & (!g43)) + ((g46) & (!sk[30]) & (!g41) & (g19) & (g43)) + ((g46) & (!sk[30]) & (g41) & (!g19) & (!g43)) + ((g46) & (!sk[30]) & (g41) & (!g19) & (g43)) + ((g46) & (!sk[30]) & (g41) & (g19) & (!g43)) + ((g46) & (!sk[30]) & (g41) & (g19) & (g43)) + ((g46) & (sk[30]) & (!g41) & (!g19) & (!g43)));
	assign g661 = (((!g17) & (!sk[31]) & (g99) & (!g40)) + ((!g17) & (!sk[31]) & (g99) & (g40)) + ((!g17) & (sk[31]) & (g99) & (g40)) + ((g17) & (!sk[31]) & (g99) & (!g40)) + ((g17) & (!sk[31]) & (g99) & (g40)) + ((g17) & (sk[31]) & (g99) & (!g40)) + ((g17) & (sk[31]) & (g99) & (g40)));
	assign g662 = (((!g62) & (!g32) & (!g621) & (!sk[32]) & (g661)) + ((!g62) & (!g32) & (g621) & (!sk[32]) & (g661)) + ((!g62) & (!g32) & (g621) & (sk[32]) & (!g661)) + ((!g62) & (g32) & (!g621) & (!sk[32]) & (g661)) + ((!g62) & (g32) & (g621) & (!sk[32]) & (g661)) + ((!g62) & (g32) & (g621) & (sk[32]) & (!g661)) + ((g62) & (!g32) & (!g621) & (!sk[32]) & (!g661)) + ((g62) & (!g32) & (!g621) & (!sk[32]) & (g661)) + ((g62) & (!g32) & (g621) & (!sk[32]) & (!g661)) + ((g62) & (!g32) & (g621) & (!sk[32]) & (g661)) + ((g62) & (!g32) & (g621) & (sk[32]) & (!g661)) + ((g62) & (g32) & (!g621) & (!sk[32]) & (!g661)) + ((g62) & (g32) & (!g621) & (!sk[32]) & (g661)) + ((g62) & (g32) & (g621) & (!sk[32]) & (!g661)) + ((g62) & (g32) & (g621) & (!sk[32]) & (g661)));
	assign g663 = (((!g55) & (!g73) & (!g278) & (g660) & (!sk[33]) & (!g662)) + ((!g55) & (!g73) & (!g278) & (g660) & (!sk[33]) & (g662)) + ((!g55) & (!g73) & (g278) & (!g660) & (!sk[33]) & (!g662)) + ((!g55) & (!g73) & (g278) & (!g660) & (!sk[33]) & (g662)) + ((!g55) & (!g73) & (g278) & (g660) & (!sk[33]) & (!g662)) + ((!g55) & (!g73) & (g278) & (g660) & (!sk[33]) & (g662)) + ((!g55) & (!g73) & (g278) & (g660) & (sk[33]) & (g662)) + ((!g55) & (g73) & (!g278) & (!g660) & (!sk[33]) & (!g662)) + ((!g55) & (g73) & (!g278) & (!g660) & (!sk[33]) & (g662)) + ((!g55) & (g73) & (!g278) & (g660) & (!sk[33]) & (!g662)) + ((!g55) & (g73) & (!g278) & (g660) & (!sk[33]) & (g662)) + ((!g55) & (g73) & (g278) & (!g660) & (!sk[33]) & (!g662)) + ((!g55) & (g73) & (g278) & (!g660) & (!sk[33]) & (g662)) + ((!g55) & (g73) & (g278) & (g660) & (!sk[33]) & (!g662)) + ((!g55) & (g73) & (g278) & (g660) & (!sk[33]) & (g662)) + ((g55) & (!g73) & (!g278) & (g660) & (!sk[33]) & (!g662)) + ((g55) & (!g73) & (!g278) & (g660) & (!sk[33]) & (g662)) + ((g55) & (!g73) & (g278) & (!g660) & (!sk[33]) & (!g662)) + ((g55) & (!g73) & (g278) & (!g660) & (!sk[33]) & (g662)) + ((g55) & (!g73) & (g278) & (g660) & (!sk[33]) & (!g662)) + ((g55) & (!g73) & (g278) & (g660) & (!sk[33]) & (g662)) + ((g55) & (g73) & (!g278) & (!g660) & (!sk[33]) & (!g662)) + ((g55) & (g73) & (!g278) & (!g660) & (!sk[33]) & (g662)) + ((g55) & (g73) & (!g278) & (g660) & (!sk[33]) & (!g662)) + ((g55) & (g73) & (!g278) & (g660) & (!sk[33]) & (g662)) + ((g55) & (g73) & (g278) & (!g660) & (!sk[33]) & (!g662)) + ((g55) & (g73) & (g278) & (!g660) & (!sk[33]) & (g662)) + ((g55) & (g73) & (g278) & (g660) & (!sk[33]) & (!g662)) + ((g55) & (g73) & (g278) & (g660) & (!sk[33]) & (g662)));
	assign g664 = (((!g70) & (!g10) & (!g551) & (!g171) & (sk[34]) & (g260)) + ((!g70) & (!g10) & (!g551) & (g171) & (!sk[34]) & (!g260)) + ((!g70) & (!g10) & (!g551) & (g171) & (!sk[34]) & (g260)) + ((!g70) & (!g10) & (g551) & (!g171) & (!sk[34]) & (!g260)) + ((!g70) & (!g10) & (g551) & (!g171) & (!sk[34]) & (g260)) + ((!g70) & (!g10) & (g551) & (g171) & (!sk[34]) & (!g260)) + ((!g70) & (!g10) & (g551) & (g171) & (!sk[34]) & (g260)) + ((!g70) & (g10) & (!g551) & (!g171) & (!sk[34]) & (!g260)) + ((!g70) & (g10) & (!g551) & (!g171) & (!sk[34]) & (g260)) + ((!g70) & (g10) & (!g551) & (!g171) & (sk[34]) & (g260)) + ((!g70) & (g10) & (!g551) & (g171) & (!sk[34]) & (!g260)) + ((!g70) & (g10) & (!g551) & (g171) & (!sk[34]) & (g260)) + ((!g70) & (g10) & (g551) & (!g171) & (!sk[34]) & (!g260)) + ((!g70) & (g10) & (g551) & (!g171) & (!sk[34]) & (g260)) + ((!g70) & (g10) & (g551) & (g171) & (!sk[34]) & (!g260)) + ((!g70) & (g10) & (g551) & (g171) & (!sk[34]) & (g260)) + ((g70) & (!g10) & (!g551) & (!g171) & (sk[34]) & (g260)) + ((g70) & (!g10) & (!g551) & (g171) & (!sk[34]) & (!g260)) + ((g70) & (!g10) & (!g551) & (g171) & (!sk[34]) & (g260)) + ((g70) & (!g10) & (g551) & (!g171) & (!sk[34]) & (!g260)) + ((g70) & (!g10) & (g551) & (!g171) & (!sk[34]) & (g260)) + ((g70) & (!g10) & (g551) & (g171) & (!sk[34]) & (!g260)) + ((g70) & (!g10) & (g551) & (g171) & (!sk[34]) & (g260)) + ((g70) & (g10) & (!g551) & (!g171) & (!sk[34]) & (!g260)) + ((g70) & (g10) & (!g551) & (!g171) & (!sk[34]) & (g260)) + ((g70) & (g10) & (!g551) & (g171) & (!sk[34]) & (!g260)) + ((g70) & (g10) & (!g551) & (g171) & (!sk[34]) & (g260)) + ((g70) & (g10) & (g551) & (!g171) & (!sk[34]) & (!g260)) + ((g70) & (g10) & (g551) & (!g171) & (!sk[34]) & (g260)) + ((g70) & (g10) & (g551) & (g171) & (!sk[34]) & (!g260)) + ((g70) & (g10) & (g551) & (g171) & (!sk[34]) & (g260)));
	assign g665 = (((!g9) & (!g10) & (!sk[35]) & (!g99) & (g42)) + ((!g9) & (!g10) & (!sk[35]) & (g99) & (g42)) + ((!g9) & (!g10) & (sk[35]) & (g99) & (g42)) + ((!g9) & (g10) & (!sk[35]) & (!g99) & (g42)) + ((!g9) & (g10) & (!sk[35]) & (g99) & (g42)) + ((!g9) & (g10) & (sk[35]) & (g99) & (g42)) + ((g9) & (!g10) & (!sk[35]) & (!g99) & (!g42)) + ((g9) & (!g10) & (!sk[35]) & (!g99) & (g42)) + ((g9) & (!g10) & (!sk[35]) & (g99) & (!g42)) + ((g9) & (!g10) & (!sk[35]) & (g99) & (g42)) + ((g9) & (!g10) & (sk[35]) & (g99) & (g42)) + ((g9) & (g10) & (!sk[35]) & (!g99) & (!g42)) + ((g9) & (g10) & (!sk[35]) & (!g99) & (g42)) + ((g9) & (g10) & (!sk[35]) & (g99) & (!g42)) + ((g9) & (g10) & (!sk[35]) & (g99) & (g42)) + ((g9) & (g10) & (sk[35]) & (!g99) & (!g42)) + ((g9) & (g10) & (sk[35]) & (!g99) & (g42)) + ((g9) & (g10) & (sk[35]) & (g99) & (!g42)) + ((g9) & (g10) & (sk[35]) & (g99) & (g42)));
	assign g666 = (((!g275) & (sk[36]) & (!g665)) + ((g275) & (!sk[36]) & (g665)));
	assign g667 = (((!g9) & (!g16) & (!g58) & (!g236) & (sk[37]) & (g666)) + ((!g9) & (!g16) & (!g58) & (g236) & (!sk[37]) & (!g666)) + ((!g9) & (!g16) & (!g58) & (g236) & (!sk[37]) & (g666)) + ((!g9) & (!g16) & (g58) & (!g236) & (!sk[37]) & (!g666)) + ((!g9) & (!g16) & (g58) & (!g236) & (!sk[37]) & (g666)) + ((!g9) & (!g16) & (g58) & (!g236) & (sk[37]) & (g666)) + ((!g9) & (!g16) & (g58) & (g236) & (!sk[37]) & (!g666)) + ((!g9) & (!g16) & (g58) & (g236) & (!sk[37]) & (g666)) + ((!g9) & (g16) & (!g58) & (!g236) & (!sk[37]) & (!g666)) + ((!g9) & (g16) & (!g58) & (!g236) & (!sk[37]) & (g666)) + ((!g9) & (g16) & (!g58) & (!g236) & (sk[37]) & (g666)) + ((!g9) & (g16) & (!g58) & (g236) & (!sk[37]) & (!g666)) + ((!g9) & (g16) & (!g58) & (g236) & (!sk[37]) & (g666)) + ((!g9) & (g16) & (g58) & (!g236) & (!sk[37]) & (!g666)) + ((!g9) & (g16) & (g58) & (!g236) & (!sk[37]) & (g666)) + ((!g9) & (g16) & (g58) & (g236) & (!sk[37]) & (!g666)) + ((!g9) & (g16) & (g58) & (g236) & (!sk[37]) & (g666)) + ((g9) & (!g16) & (!g58) & (!g236) & (sk[37]) & (g666)) + ((g9) & (!g16) & (!g58) & (g236) & (!sk[37]) & (!g666)) + ((g9) & (!g16) & (!g58) & (g236) & (!sk[37]) & (g666)) + ((g9) & (!g16) & (g58) & (!g236) & (!sk[37]) & (!g666)) + ((g9) & (!g16) & (g58) & (!g236) & (!sk[37]) & (g666)) + ((g9) & (!g16) & (g58) & (g236) & (!sk[37]) & (!g666)) + ((g9) & (!g16) & (g58) & (g236) & (!sk[37]) & (g666)) + ((g9) & (g16) & (!g58) & (!g236) & (!sk[37]) & (!g666)) + ((g9) & (g16) & (!g58) & (!g236) & (!sk[37]) & (g666)) + ((g9) & (g16) & (!g58) & (!g236) & (sk[37]) & (g666)) + ((g9) & (g16) & (!g58) & (g236) & (!sk[37]) & (!g666)) + ((g9) & (g16) & (!g58) & (g236) & (!sk[37]) & (g666)) + ((g9) & (g16) & (g58) & (!g236) & (!sk[37]) & (!g666)) + ((g9) & (g16) & (g58) & (!g236) & (!sk[37]) & (g666)) + ((g9) & (g16) & (g58) & (g236) & (!sk[37]) & (!g666)) + ((g9) & (g16) & (g58) & (g236) & (!sk[37]) & (g666)));
	assign g668 = (((!g70) & (!g17) & (!g104) & (!sk[38]) & (g572) & (!g288)) + ((!g70) & (!g17) & (!g104) & (!sk[38]) & (g572) & (g288)) + ((!g70) & (!g17) & (!g104) & (sk[38]) & (!g572) & (!g288)) + ((!g70) & (!g17) & (g104) & (!sk[38]) & (!g572) & (!g288)) + ((!g70) & (!g17) & (g104) & (!sk[38]) & (!g572) & (g288)) + ((!g70) & (!g17) & (g104) & (!sk[38]) & (g572) & (!g288)) + ((!g70) & (!g17) & (g104) & (!sk[38]) & (g572) & (g288)) + ((!g70) & (!g17) & (g104) & (sk[38]) & (!g572) & (!g288)) + ((!g70) & (g17) & (!g104) & (!sk[38]) & (!g572) & (!g288)) + ((!g70) & (g17) & (!g104) & (!sk[38]) & (!g572) & (g288)) + ((!g70) & (g17) & (!g104) & (!sk[38]) & (g572) & (!g288)) + ((!g70) & (g17) & (!g104) & (!sk[38]) & (g572) & (g288)) + ((!g70) & (g17) & (!g104) & (sk[38]) & (!g572) & (!g288)) + ((!g70) & (g17) & (g104) & (!sk[38]) & (!g572) & (!g288)) + ((!g70) & (g17) & (g104) & (!sk[38]) & (!g572) & (g288)) + ((!g70) & (g17) & (g104) & (!sk[38]) & (g572) & (!g288)) + ((!g70) & (g17) & (g104) & (!sk[38]) & (g572) & (g288)) + ((g70) & (!g17) & (!g104) & (!sk[38]) & (g572) & (!g288)) + ((g70) & (!g17) & (!g104) & (!sk[38]) & (g572) & (g288)) + ((g70) & (!g17) & (!g104) & (sk[38]) & (!g572) & (!g288)) + ((g70) & (!g17) & (g104) & (!sk[38]) & (!g572) & (!g288)) + ((g70) & (!g17) & (g104) & (!sk[38]) & (!g572) & (g288)) + ((g70) & (!g17) & (g104) & (!sk[38]) & (g572) & (!g288)) + ((g70) & (!g17) & (g104) & (!sk[38]) & (g572) & (g288)) + ((g70) & (!g17) & (g104) & (sk[38]) & (!g572) & (!g288)) + ((g70) & (g17) & (!g104) & (!sk[38]) & (!g572) & (!g288)) + ((g70) & (g17) & (!g104) & (!sk[38]) & (!g572) & (g288)) + ((g70) & (g17) & (!g104) & (!sk[38]) & (g572) & (!g288)) + ((g70) & (g17) & (!g104) & (!sk[38]) & (g572) & (g288)) + ((g70) & (g17) & (g104) & (!sk[38]) & (!g572) & (!g288)) + ((g70) & (g17) & (g104) & (!sk[38]) & (!g572) & (g288)) + ((g70) & (g17) & (g104) & (!sk[38]) & (g572) & (!g288)) + ((g70) & (g17) & (g104) & (!sk[38]) & (g572) & (g288)));
	assign g669 = (((!sk[39]) & (!g99) & (!g18) & (!g664) & (g667) & (!g668)) + ((!sk[39]) & (!g99) & (!g18) & (!g664) & (g667) & (g668)) + ((!sk[39]) & (!g99) & (!g18) & (g664) & (!g667) & (!g668)) + ((!sk[39]) & (!g99) & (!g18) & (g664) & (!g667) & (g668)) + ((!sk[39]) & (!g99) & (!g18) & (g664) & (g667) & (!g668)) + ((!sk[39]) & (!g99) & (!g18) & (g664) & (g667) & (g668)) + ((!sk[39]) & (!g99) & (g18) & (!g664) & (!g667) & (!g668)) + ((!sk[39]) & (!g99) & (g18) & (!g664) & (!g667) & (g668)) + ((!sk[39]) & (!g99) & (g18) & (!g664) & (g667) & (!g668)) + ((!sk[39]) & (!g99) & (g18) & (!g664) & (g667) & (g668)) + ((!sk[39]) & (!g99) & (g18) & (g664) & (!g667) & (!g668)) + ((!sk[39]) & (!g99) & (g18) & (g664) & (!g667) & (g668)) + ((!sk[39]) & (!g99) & (g18) & (g664) & (g667) & (!g668)) + ((!sk[39]) & (!g99) & (g18) & (g664) & (g667) & (g668)) + ((!sk[39]) & (g99) & (!g18) & (!g664) & (g667) & (!g668)) + ((!sk[39]) & (g99) & (!g18) & (!g664) & (g667) & (g668)) + ((!sk[39]) & (g99) & (!g18) & (g664) & (!g667) & (!g668)) + ((!sk[39]) & (g99) & (!g18) & (g664) & (!g667) & (g668)) + ((!sk[39]) & (g99) & (!g18) & (g664) & (g667) & (!g668)) + ((!sk[39]) & (g99) & (!g18) & (g664) & (g667) & (g668)) + ((!sk[39]) & (g99) & (g18) & (!g664) & (!g667) & (!g668)) + ((!sk[39]) & (g99) & (g18) & (!g664) & (!g667) & (g668)) + ((!sk[39]) & (g99) & (g18) & (!g664) & (g667) & (!g668)) + ((!sk[39]) & (g99) & (g18) & (!g664) & (g667) & (g668)) + ((!sk[39]) & (g99) & (g18) & (g664) & (!g667) & (!g668)) + ((!sk[39]) & (g99) & (g18) & (g664) & (!g667) & (g668)) + ((!sk[39]) & (g99) & (g18) & (g664) & (g667) & (!g668)) + ((!sk[39]) & (g99) & (g18) & (g664) & (g667) & (g668)) + ((sk[39]) & (!g99) & (!g18) & (g664) & (g667) & (g668)) + ((sk[39]) & (!g99) & (g18) & (g664) & (g667) & (g668)) + ((sk[39]) & (g99) & (!g18) & (g664) & (g667) & (g668)));
	assign g670 = (((!sk[40]) & (!g604) & (!g617) & (!g659) & (g663) & (!g669)) + ((!sk[40]) & (!g604) & (!g617) & (!g659) & (g663) & (g669)) + ((!sk[40]) & (!g604) & (!g617) & (g659) & (!g663) & (!g669)) + ((!sk[40]) & (!g604) & (!g617) & (g659) & (!g663) & (g669)) + ((!sk[40]) & (!g604) & (!g617) & (g659) & (g663) & (!g669)) + ((!sk[40]) & (!g604) & (!g617) & (g659) & (g663) & (g669)) + ((!sk[40]) & (!g604) & (g617) & (!g659) & (!g663) & (!g669)) + ((!sk[40]) & (!g604) & (g617) & (!g659) & (!g663) & (g669)) + ((!sk[40]) & (!g604) & (g617) & (!g659) & (g663) & (!g669)) + ((!sk[40]) & (!g604) & (g617) & (!g659) & (g663) & (g669)) + ((!sk[40]) & (!g604) & (g617) & (g659) & (!g663) & (!g669)) + ((!sk[40]) & (!g604) & (g617) & (g659) & (!g663) & (g669)) + ((!sk[40]) & (!g604) & (g617) & (g659) & (g663) & (!g669)) + ((!sk[40]) & (!g604) & (g617) & (g659) & (g663) & (g669)) + ((!sk[40]) & (g604) & (!g617) & (!g659) & (g663) & (!g669)) + ((!sk[40]) & (g604) & (!g617) & (!g659) & (g663) & (g669)) + ((!sk[40]) & (g604) & (!g617) & (g659) & (!g663) & (!g669)) + ((!sk[40]) & (g604) & (!g617) & (g659) & (!g663) & (g669)) + ((!sk[40]) & (g604) & (!g617) & (g659) & (g663) & (!g669)) + ((!sk[40]) & (g604) & (!g617) & (g659) & (g663) & (g669)) + ((!sk[40]) & (g604) & (g617) & (!g659) & (!g663) & (!g669)) + ((!sk[40]) & (g604) & (g617) & (!g659) & (!g663) & (g669)) + ((!sk[40]) & (g604) & (g617) & (!g659) & (g663) & (!g669)) + ((!sk[40]) & (g604) & (g617) & (!g659) & (g663) & (g669)) + ((!sk[40]) & (g604) & (g617) & (g659) & (!g663) & (!g669)) + ((!sk[40]) & (g604) & (g617) & (g659) & (!g663) & (g669)) + ((!sk[40]) & (g604) & (g617) & (g659) & (g663) & (!g669)) + ((!sk[40]) & (g604) & (g617) & (g659) & (g663) & (g669)) + ((sk[40]) & (g604) & (g617) & (g659) & (g663) & (g669)));
	assign g671 = (((!g194) & (!sk[41]) & (!g129) & (!g92) & (g415) & (!g94)) + ((!g194) & (!sk[41]) & (!g129) & (!g92) & (g415) & (g94)) + ((!g194) & (!sk[41]) & (!g129) & (g92) & (!g415) & (!g94)) + ((!g194) & (!sk[41]) & (!g129) & (g92) & (!g415) & (g94)) + ((!g194) & (!sk[41]) & (!g129) & (g92) & (g415) & (!g94)) + ((!g194) & (!sk[41]) & (!g129) & (g92) & (g415) & (g94)) + ((!g194) & (!sk[41]) & (g129) & (!g92) & (!g415) & (!g94)) + ((!g194) & (!sk[41]) & (g129) & (!g92) & (!g415) & (g94)) + ((!g194) & (!sk[41]) & (g129) & (!g92) & (g415) & (!g94)) + ((!g194) & (!sk[41]) & (g129) & (!g92) & (g415) & (g94)) + ((!g194) & (!sk[41]) & (g129) & (g92) & (!g415) & (!g94)) + ((!g194) & (!sk[41]) & (g129) & (g92) & (!g415) & (g94)) + ((!g194) & (!sk[41]) & (g129) & (g92) & (g415) & (!g94)) + ((!g194) & (!sk[41]) & (g129) & (g92) & (g415) & (g94)) + ((!g194) & (sk[41]) & (!g129) & (g92) & (!g415) & (g94)) + ((g194) & (!sk[41]) & (!g129) & (!g92) & (g415) & (!g94)) + ((g194) & (!sk[41]) & (!g129) & (!g92) & (g415) & (g94)) + ((g194) & (!sk[41]) & (!g129) & (g92) & (!g415) & (!g94)) + ((g194) & (!sk[41]) & (!g129) & (g92) & (!g415) & (g94)) + ((g194) & (!sk[41]) & (!g129) & (g92) & (g415) & (!g94)) + ((g194) & (!sk[41]) & (!g129) & (g92) & (g415) & (g94)) + ((g194) & (!sk[41]) & (g129) & (!g92) & (!g415) & (!g94)) + ((g194) & (!sk[41]) & (g129) & (!g92) & (!g415) & (g94)) + ((g194) & (!sk[41]) & (g129) & (!g92) & (g415) & (!g94)) + ((g194) & (!sk[41]) & (g129) & (!g92) & (g415) & (g94)) + ((g194) & (!sk[41]) & (g129) & (g92) & (!g415) & (!g94)) + ((g194) & (!sk[41]) & (g129) & (g92) & (!g415) & (g94)) + ((g194) & (!sk[41]) & (g129) & (g92) & (g415) & (!g94)) + ((g194) & (!sk[41]) & (g129) & (g92) & (g415) & (g94)));
	assign g672 = (((!g59) & (!g72) & (!g236) & (g348) & (g552) & (g671)));
	assign g673 = (((!g62) & (!sk[43]) & (g146) & (!g32)) + ((!g62) & (!sk[43]) & (g146) & (g32)) + ((!g62) & (sk[43]) & (!g146) & (!g32)) + ((!g62) & (sk[43]) & (!g146) & (g32)) + ((g62) & (!sk[43]) & (g146) & (!g32)) + ((g62) & (!sk[43]) & (g146) & (g32)) + ((g62) & (sk[43]) & (!g146) & (!g32)));
	assign g674 = (((!g70) & (!sk[44]) & (!g18) & (!g104) & (g36)) + ((!g70) & (!sk[44]) & (!g18) & (g104) & (g36)) + ((!g70) & (!sk[44]) & (g18) & (!g104) & (g36)) + ((!g70) & (!sk[44]) & (g18) & (g104) & (g36)) + ((!g70) & (sk[44]) & (!g18) & (!g104) & (!g36)) + ((!g70) & (sk[44]) & (!g18) & (g104) & (!g36)) + ((!g70) & (sk[44]) & (g18) & (!g104) & (!g36)) + ((g70) & (!sk[44]) & (!g18) & (!g104) & (!g36)) + ((g70) & (!sk[44]) & (!g18) & (!g104) & (g36)) + ((g70) & (!sk[44]) & (!g18) & (g104) & (!g36)) + ((g70) & (!sk[44]) & (!g18) & (g104) & (g36)) + ((g70) & (!sk[44]) & (g18) & (!g104) & (!g36)) + ((g70) & (!sk[44]) & (g18) & (!g104) & (g36)) + ((g70) & (!sk[44]) & (g18) & (g104) & (!g36)) + ((g70) & (!sk[44]) & (g18) & (g104) & (g36)) + ((g70) & (sk[44]) & (!g18) & (!g104) & (!g36)) + ((g70) & (sk[44]) & (!g18) & (g104) & (!g36)));
	assign g675 = (((!g673) & (!g118) & (!g328) & (!sk[45]) & (g644) & (!g674)) + ((!g673) & (!g118) & (!g328) & (!sk[45]) & (g644) & (g674)) + ((!g673) & (!g118) & (g328) & (!sk[45]) & (!g644) & (!g674)) + ((!g673) & (!g118) & (g328) & (!sk[45]) & (!g644) & (g674)) + ((!g673) & (!g118) & (g328) & (!sk[45]) & (g644) & (!g674)) + ((!g673) & (!g118) & (g328) & (!sk[45]) & (g644) & (g674)) + ((!g673) & (g118) & (!g328) & (!sk[45]) & (!g644) & (!g674)) + ((!g673) & (g118) & (!g328) & (!sk[45]) & (!g644) & (g674)) + ((!g673) & (g118) & (!g328) & (!sk[45]) & (g644) & (!g674)) + ((!g673) & (g118) & (!g328) & (!sk[45]) & (g644) & (g674)) + ((!g673) & (g118) & (g328) & (!sk[45]) & (!g644) & (!g674)) + ((!g673) & (g118) & (g328) & (!sk[45]) & (!g644) & (g674)) + ((!g673) & (g118) & (g328) & (!sk[45]) & (g644) & (!g674)) + ((!g673) & (g118) & (g328) & (!sk[45]) & (g644) & (g674)) + ((g673) & (!g118) & (!g328) & (!sk[45]) & (g644) & (!g674)) + ((g673) & (!g118) & (!g328) & (!sk[45]) & (g644) & (g674)) + ((g673) & (!g118) & (g328) & (!sk[45]) & (!g644) & (!g674)) + ((g673) & (!g118) & (g328) & (!sk[45]) & (!g644) & (g674)) + ((g673) & (!g118) & (g328) & (!sk[45]) & (g644) & (!g674)) + ((g673) & (!g118) & (g328) & (!sk[45]) & (g644) & (g674)) + ((g673) & (g118) & (!g328) & (!sk[45]) & (!g644) & (!g674)) + ((g673) & (g118) & (!g328) & (!sk[45]) & (!g644) & (g674)) + ((g673) & (g118) & (!g328) & (!sk[45]) & (g644) & (!g674)) + ((g673) & (g118) & (!g328) & (!sk[45]) & (g644) & (g674)) + ((g673) & (g118) & (g328) & (!sk[45]) & (!g644) & (!g674)) + ((g673) & (g118) & (g328) & (!sk[45]) & (!g644) & (g674)) + ((g673) & (g118) & (g328) & (!sk[45]) & (g644) & (!g674)) + ((g673) & (g118) & (g328) & (!sk[45]) & (g644) & (g674)) + ((g673) & (g118) & (g328) & (sk[45]) & (g644) & (g674)));
	assign g676 = (((!sk[46]) & (!g672) & (!g102) & (!g178) & (g634) & (!g675)) + ((!sk[46]) & (!g672) & (!g102) & (!g178) & (g634) & (g675)) + ((!sk[46]) & (!g672) & (!g102) & (g178) & (!g634) & (!g675)) + ((!sk[46]) & (!g672) & (!g102) & (g178) & (!g634) & (g675)) + ((!sk[46]) & (!g672) & (!g102) & (g178) & (g634) & (!g675)) + ((!sk[46]) & (!g672) & (!g102) & (g178) & (g634) & (g675)) + ((!sk[46]) & (!g672) & (g102) & (!g178) & (!g634) & (!g675)) + ((!sk[46]) & (!g672) & (g102) & (!g178) & (!g634) & (g675)) + ((!sk[46]) & (!g672) & (g102) & (!g178) & (g634) & (!g675)) + ((!sk[46]) & (!g672) & (g102) & (!g178) & (g634) & (g675)) + ((!sk[46]) & (!g672) & (g102) & (g178) & (!g634) & (!g675)) + ((!sk[46]) & (!g672) & (g102) & (g178) & (!g634) & (g675)) + ((!sk[46]) & (!g672) & (g102) & (g178) & (g634) & (!g675)) + ((!sk[46]) & (!g672) & (g102) & (g178) & (g634) & (g675)) + ((!sk[46]) & (g672) & (!g102) & (!g178) & (g634) & (!g675)) + ((!sk[46]) & (g672) & (!g102) & (!g178) & (g634) & (g675)) + ((!sk[46]) & (g672) & (!g102) & (g178) & (!g634) & (!g675)) + ((!sk[46]) & (g672) & (!g102) & (g178) & (!g634) & (g675)) + ((!sk[46]) & (g672) & (!g102) & (g178) & (g634) & (!g675)) + ((!sk[46]) & (g672) & (!g102) & (g178) & (g634) & (g675)) + ((!sk[46]) & (g672) & (g102) & (!g178) & (!g634) & (!g675)) + ((!sk[46]) & (g672) & (g102) & (!g178) & (!g634) & (g675)) + ((!sk[46]) & (g672) & (g102) & (!g178) & (g634) & (!g675)) + ((!sk[46]) & (g672) & (g102) & (!g178) & (g634) & (g675)) + ((!sk[46]) & (g672) & (g102) & (g178) & (!g634) & (!g675)) + ((!sk[46]) & (g672) & (g102) & (g178) & (!g634) & (g675)) + ((!sk[46]) & (g672) & (g102) & (g178) & (g634) & (!g675)) + ((!sk[46]) & (g672) & (g102) & (g178) & (g634) & (g675)) + ((sk[46]) & (g672) & (g102) & (g178) & (g634) & (g675)));
	assign g677 = (((!g656) & (!g657) & (!g488) & (!g658) & (g670) & (g676)) + ((!g656) & (!g657) & (g488) & (!g658) & (g670) & (!g676)) + ((!g656) & (!g657) & (g488) & (!g658) & (g670) & (g676)) + ((!g656) & (!g657) & (g488) & (g658) & (g670) & (g676)) + ((!g656) & (g657) & (!g488) & (!g658) & (g670) & (!g676)) + ((!g656) & (g657) & (!g488) & (!g658) & (g670) & (g676)) + ((!g656) & (g657) & (!g488) & (g658) & (g670) & (g676)) + ((!g656) & (g657) & (g488) & (!g658) & (!g670) & (g676)) + ((!g656) & (g657) & (g488) & (!g658) & (g670) & (!g676)) + ((!g656) & (g657) & (g488) & (!g658) & (g670) & (g676)) + ((!g656) & (g657) & (g488) & (g658) & (g670) & (!g676)) + ((!g656) & (g657) & (g488) & (g658) & (g670) & (g676)) + ((g656) & (!g657) & (!g488) & (!g658) & (!g670) & (g676)) + ((g656) & (!g657) & (!g488) & (!g658) & (g670) & (!g676)) + ((g656) & (!g657) & (!g488) & (!g658) & (g670) & (g676)) + ((g656) & (!g657) & (!g488) & (g658) & (g670) & (!g676)) + ((g656) & (!g657) & (!g488) & (g658) & (g670) & (g676)) + ((g656) & (!g657) & (g488) & (g658) & (!g670) & (g676)) + ((g656) & (!g657) & (g488) & (g658) & (g670) & (!g676)) + ((g656) & (!g657) & (g488) & (g658) & (g670) & (g676)) + ((g656) & (g657) & (!g488) & (g658) & (!g670) & (g676)) + ((g656) & (g657) & (!g488) & (g658) & (g670) & (!g676)) + ((g656) & (g657) & (!g488) & (g658) & (g670) & (g676)) + ((g656) & (g657) & (g488) & (!g658) & (g670) & (g676)));
	assign g678 = (((!g627) & (!g546) & (!g640) & (!g641) & (!g655) & (g677)) + ((!g627) & (!g546) & (!g640) & (!g641) & (g655) & (!g677)) + ((!g627) & (!g546) & (!g640) & (!g641) & (g655) & (g677)) + ((!g627) & (!g546) & (!g640) & (g641) & (g655) & (g677)) + ((!g627) & (!g546) & (g640) & (!g641) & (!g655) & (!g677)) + ((!g627) & (!g546) & (g640) & (!g641) & (!g655) & (g677)) + ((!g627) & (!g546) & (g640) & (!g641) & (g655) & (!g677)) + ((!g627) & (!g546) & (g640) & (!g641) & (g655) & (g677)) + ((!g627) & (!g546) & (g640) & (g641) & (!g655) & (!g677)) + ((!g627) & (!g546) & (g640) & (g641) & (!g655) & (g677)) + ((!g627) & (!g546) & (g640) & (g641) & (g655) & (!g677)) + ((!g627) & (!g546) & (g640) & (g641) & (g655) & (g677)) + ((!g627) & (g546) & (g640) & (!g641) & (!g655) & (g677)) + ((!g627) & (g546) & (g640) & (!g641) & (g655) & (!g677)) + ((!g627) & (g546) & (g640) & (!g641) & (g655) & (g677)) + ((!g627) & (g546) & (g640) & (g641) & (g655) & (g677)) + ((g627) & (!g546) & (g640) & (!g641) & (!g655) & (g677)) + ((g627) & (!g546) & (g640) & (!g641) & (g655) & (!g677)) + ((g627) & (!g546) & (g640) & (!g641) & (g655) & (g677)) + ((g627) & (!g546) & (g640) & (g641) & (g655) & (g677)) + ((g627) & (g546) & (!g640) & (!g641) & (!g655) & (g677)) + ((g627) & (g546) & (!g640) & (!g641) & (g655) & (!g677)) + ((g627) & (g546) & (!g640) & (!g641) & (g655) & (g677)) + ((g627) & (g546) & (!g640) & (g641) & (g655) & (g677)) + ((g627) & (g546) & (g640) & (!g641) & (!g655) & (!g677)) + ((g627) & (g546) & (g640) & (!g641) & (!g655) & (g677)) + ((g627) & (g546) & (g640) & (!g641) & (g655) & (!g677)) + ((g627) & (g546) & (g640) & (!g641) & (g655) & (g677)) + ((g627) & (g546) & (g640) & (g641) & (!g655) & (!g677)) + ((g627) & (g546) & (g640) & (g641) & (!g655) & (g677)) + ((g627) & (g546) & (g640) & (g641) & (g655) & (!g677)) + ((g627) & (g546) & (g640) & (g641) & (g655) & (g677)));
	assign g679 = (((!g598) & (!g611) & (!sk[49]) & (!g612) & (g626) & (!g678)) + ((!g598) & (!g611) & (!sk[49]) & (!g612) & (g626) & (g678)) + ((!g598) & (!g611) & (!sk[49]) & (g612) & (!g626) & (!g678)) + ((!g598) & (!g611) & (!sk[49]) & (g612) & (!g626) & (g678)) + ((!g598) & (!g611) & (!sk[49]) & (g612) & (g626) & (!g678)) + ((!g598) & (!g611) & (!sk[49]) & (g612) & (g626) & (g678)) + ((!g598) & (!g611) & (sk[49]) & (!g612) & (!g626) & (g678)) + ((!g598) & (!g611) & (sk[49]) & (!g612) & (g626) & (!g678)) + ((!g598) & (!g611) & (sk[49]) & (!g612) & (g626) & (g678)) + ((!g598) & (!g611) & (sk[49]) & (g612) & (g626) & (g678)) + ((!g598) & (g611) & (!sk[49]) & (!g612) & (!g626) & (!g678)) + ((!g598) & (g611) & (!sk[49]) & (!g612) & (!g626) & (g678)) + ((!g598) & (g611) & (!sk[49]) & (!g612) & (g626) & (!g678)) + ((!g598) & (g611) & (!sk[49]) & (!g612) & (g626) & (g678)) + ((!g598) & (g611) & (!sk[49]) & (g612) & (!g626) & (!g678)) + ((!g598) & (g611) & (!sk[49]) & (g612) & (!g626) & (g678)) + ((!g598) & (g611) & (!sk[49]) & (g612) & (g626) & (!g678)) + ((!g598) & (g611) & (!sk[49]) & (g612) & (g626) & (g678)) + ((!g598) & (g611) & (sk[49]) & (!g612) & (!g626) & (!g678)) + ((!g598) & (g611) & (sk[49]) & (!g612) & (!g626) & (g678)) + ((!g598) & (g611) & (sk[49]) & (!g612) & (g626) & (!g678)) + ((!g598) & (g611) & (sk[49]) & (!g612) & (g626) & (g678)) + ((!g598) & (g611) & (sk[49]) & (g612) & (!g626) & (!g678)) + ((!g598) & (g611) & (sk[49]) & (g612) & (!g626) & (g678)) + ((!g598) & (g611) & (sk[49]) & (g612) & (g626) & (!g678)) + ((!g598) & (g611) & (sk[49]) & (g612) & (g626) & (g678)) + ((g598) & (!g611) & (!sk[49]) & (!g612) & (g626) & (!g678)) + ((g598) & (!g611) & (!sk[49]) & (!g612) & (g626) & (g678)) + ((g598) & (!g611) & (!sk[49]) & (g612) & (!g626) & (!g678)) + ((g598) & (!g611) & (!sk[49]) & (g612) & (!g626) & (g678)) + ((g598) & (!g611) & (!sk[49]) & (g612) & (g626) & (!g678)) + ((g598) & (!g611) & (!sk[49]) & (g612) & (g626) & (g678)) + ((g598) & (g611) & (!sk[49]) & (!g612) & (!g626) & (!g678)) + ((g598) & (g611) & (!sk[49]) & (!g612) & (!g626) & (g678)) + ((g598) & (g611) & (!sk[49]) & (!g612) & (g626) & (!g678)) + ((g598) & (g611) & (!sk[49]) & (!g612) & (g626) & (g678)) + ((g598) & (g611) & (!sk[49]) & (g612) & (!g626) & (!g678)) + ((g598) & (g611) & (!sk[49]) & (g612) & (!g626) & (g678)) + ((g598) & (g611) & (!sk[49]) & (g612) & (g626) & (!g678)) + ((g598) & (g611) & (!sk[49]) & (g612) & (g626) & (g678)) + ((g598) & (g611) & (sk[49]) & (!g612) & (!g626) & (g678)) + ((g598) & (g611) & (sk[49]) & (!g612) & (g626) & (!g678)) + ((g598) & (g611) & (sk[49]) & (!g612) & (g626) & (g678)) + ((g598) & (g611) & (sk[49]) & (g612) & (g626) & (g678)));
	assign g680 = (((!g570) & (!g571) & (g584) & (!g585) & (!g597) & (g679)) + ((!g570) & (!g571) & (g584) & (!g585) & (g597) & (!g679)) + ((!g570) & (!g571) & (g584) & (!g585) & (g597) & (g679)) + ((!g570) & (!g571) & (g584) & (g585) & (g597) & (g679)) + ((!g570) & (g571) & (!g584) & (!g585) & (!g597) & (g679)) + ((!g570) & (g571) & (!g584) & (!g585) & (g597) & (!g679)) + ((!g570) & (g571) & (!g584) & (!g585) & (g597) & (g679)) + ((!g570) & (g571) & (!g584) & (g585) & (g597) & (g679)) + ((!g570) & (g571) & (g584) & (!g585) & (!g597) & (!g679)) + ((!g570) & (g571) & (g584) & (!g585) & (!g597) & (g679)) + ((!g570) & (g571) & (g584) & (!g585) & (g597) & (!g679)) + ((!g570) & (g571) & (g584) & (!g585) & (g597) & (g679)) + ((!g570) & (g571) & (g584) & (g585) & (!g597) & (!g679)) + ((!g570) & (g571) & (g584) & (g585) & (!g597) & (g679)) + ((!g570) & (g571) & (g584) & (g585) & (g597) & (!g679)) + ((!g570) & (g571) & (g584) & (g585) & (g597) & (g679)) + ((g570) & (!g571) & (!g584) & (!g585) & (!g597) & (g679)) + ((g570) & (!g571) & (!g584) & (!g585) & (g597) & (!g679)) + ((g570) & (!g571) & (!g584) & (!g585) & (g597) & (g679)) + ((g570) & (!g571) & (!g584) & (g585) & (g597) & (g679)) + ((g570) & (!g571) & (g584) & (!g585) & (!g597) & (!g679)) + ((g570) & (!g571) & (g584) & (!g585) & (!g597) & (g679)) + ((g570) & (!g571) & (g584) & (!g585) & (g597) & (!g679)) + ((g570) & (!g571) & (g584) & (!g585) & (g597) & (g679)) + ((g570) & (!g571) & (g584) & (g585) & (!g597) & (!g679)) + ((g570) & (!g571) & (g584) & (g585) & (!g597) & (g679)) + ((g570) & (!g571) & (g584) & (g585) & (g597) & (!g679)) + ((g570) & (!g571) & (g584) & (g585) & (g597) & (g679)) + ((g570) & (g571) & (g584) & (!g585) & (!g597) & (g679)) + ((g570) & (g571) & (g584) & (!g585) & (g597) & (!g679)) + ((g570) & (g571) & (g584) & (!g585) & (g597) & (g679)) + ((g570) & (g571) & (g584) & (g585) & (g597) & (g679)));
	assign g681 = (((!g549) & (!sk[51]) & (g569) & (!g680)) + ((!g549) & (!sk[51]) & (g569) & (g680)) + ((!g549) & (sk[51]) & (!g569) & (!g680)) + ((!g549) & (sk[51]) & (g569) & (g680)) + ((g549) & (!sk[51]) & (g569) & (!g680)) + ((g549) & (!sk[51]) & (g569) & (g680)) + ((g549) & (sk[51]) & (!g569) & (g680)) + ((g549) & (sk[51]) & (g569) & (!g680)));
	assign g682 = (((!g2) & (sk[52]) & (g401)) + ((g2) & (!sk[52]) & (g401)) + ((g2) & (sk[52]) & (!g401)));
	assign g683 = (((!sk[53]) & (!ax22x) & (!ax2x) & (!ax0x) & (ax1x)) + ((!sk[53]) & (!ax22x) & (!ax2x) & (ax0x) & (ax1x)) + ((!sk[53]) & (!ax22x) & (ax2x) & (!ax0x) & (ax1x)) + ((!sk[53]) & (!ax22x) & (ax2x) & (ax0x) & (ax1x)) + ((!sk[53]) & (ax22x) & (!ax2x) & (!ax0x) & (!ax1x)) + ((!sk[53]) & (ax22x) & (!ax2x) & (!ax0x) & (ax1x)) + ((!sk[53]) & (ax22x) & (!ax2x) & (ax0x) & (!ax1x)) + ((!sk[53]) & (ax22x) & (!ax2x) & (ax0x) & (ax1x)) + ((!sk[53]) & (ax22x) & (ax2x) & (!ax0x) & (!ax1x)) + ((!sk[53]) & (ax22x) & (ax2x) & (!ax0x) & (ax1x)) + ((!sk[53]) & (ax22x) & (ax2x) & (ax0x) & (!ax1x)) + ((!sk[53]) & (ax22x) & (ax2x) & (ax0x) & (ax1x)) + ((sk[53]) & (!ax22x) & (!ax2x) & (!ax0x) & (ax1x)) + ((sk[53]) & (!ax22x) & (!ax2x) & (ax0x) & (!ax1x)) + ((sk[53]) & (!ax22x) & (!ax2x) & (ax0x) & (ax1x)) + ((sk[53]) & (!ax22x) & (ax2x) & (!ax0x) & (!ax1x)) + ((sk[53]) & (ax22x) & (ax2x) & (!ax0x) & (!ax1x)) + ((sk[53]) & (ax22x) & (ax2x) & (!ax0x) & (ax1x)) + ((sk[53]) & (ax22x) & (ax2x) & (ax0x) & (!ax1x)) + ((sk[53]) & (ax22x) & (ax2x) & (ax0x) & (ax1x)));
	assign g684 = (((!sk[54]) & (g414) & (g683)) + ((sk[54]) & (!g414) & (g683)) + ((sk[54]) & (g414) & (!g683)));
	assign g685 = (((!g401) & (sk[55]) & (g414)) + ((g401) & (!sk[55]) & (g414)) + ((g401) & (sk[55]) & (!g414)));
	assign g686 = (((!sk[56]) & (!g682) & (g684) & (!g685)) + ((!sk[56]) & (!g682) & (g684) & (g685)) + ((!sk[56]) & (g682) & (g684) & (!g685)) + ((!sk[56]) & (g682) & (g684) & (g685)) + ((sk[56]) & (g682) & (!g684) & (!g685)));
	assign g687 = (((!g202) & (!g69) & (!g319) & (!sk[57]) & (g320)) + ((!g202) & (!g69) & (!g319) & (sk[57]) & (!g320)) + ((!g202) & (!g69) & (g319) & (!sk[57]) & (g320)) + ((!g202) & (g69) & (!g319) & (!sk[57]) & (g320)) + ((!g202) & (g69) & (!g319) & (sk[57]) & (!g320)) + ((!g202) & (g69) & (g319) & (!sk[57]) & (g320)) + ((g202) & (!g69) & (!g319) & (!sk[57]) & (!g320)) + ((g202) & (!g69) & (!g319) & (!sk[57]) & (g320)) + ((g202) & (!g69) & (!g319) & (sk[57]) & (!g320)) + ((g202) & (!g69) & (!g319) & (sk[57]) & (g320)) + ((g202) & (!g69) & (g319) & (!sk[57]) & (!g320)) + ((g202) & (!g69) & (g319) & (!sk[57]) & (g320)) + ((g202) & (!g69) & (g319) & (sk[57]) & (!g320)) + ((g202) & (g69) & (!g319) & (!sk[57]) & (!g320)) + ((g202) & (g69) & (!g319) & (!sk[57]) & (g320)) + ((g202) & (g69) & (!g319) & (sk[57]) & (!g320)) + ((g202) & (g69) & (g319) & (!sk[57]) & (!g320)) + ((g202) & (g69) & (g319) & (!sk[57]) & (g320)));
	assign g688 = (((!g252) & (!sk[58]) & (!g218) & (!g253) & (g220) & (!g221)) + ((!g252) & (!sk[58]) & (!g218) & (!g253) & (g220) & (g221)) + ((!g252) & (!sk[58]) & (!g218) & (g253) & (!g220) & (!g221)) + ((!g252) & (!sk[58]) & (!g218) & (g253) & (!g220) & (g221)) + ((!g252) & (!sk[58]) & (!g218) & (g253) & (g220) & (!g221)) + ((!g252) & (!sk[58]) & (!g218) & (g253) & (g220) & (g221)) + ((!g252) & (!sk[58]) & (g218) & (!g253) & (!g220) & (!g221)) + ((!g252) & (!sk[58]) & (g218) & (!g253) & (!g220) & (g221)) + ((!g252) & (!sk[58]) & (g218) & (!g253) & (g220) & (!g221)) + ((!g252) & (!sk[58]) & (g218) & (!g253) & (g220) & (g221)) + ((!g252) & (!sk[58]) & (g218) & (g253) & (!g220) & (!g221)) + ((!g252) & (!sk[58]) & (g218) & (g253) & (!g220) & (g221)) + ((!g252) & (!sk[58]) & (g218) & (g253) & (g220) & (!g221)) + ((!g252) & (!sk[58]) & (g218) & (g253) & (g220) & (g221)) + ((!g252) & (sk[58]) & (!g218) & (!g253) & (!g220) & (g221)) + ((!g252) & (sk[58]) & (!g218) & (!g253) & (g220) & (g221)) + ((!g252) & (sk[58]) & (!g218) & (g253) & (g220) & (g221)) + ((!g252) & (sk[58]) & (g218) & (!g253) & (!g220) & (g221)) + ((!g252) & (sk[58]) & (g218) & (!g253) & (g220) & (g221)) + ((!g252) & (sk[58]) & (g218) & (g253) & (!g220) & (!g221)) + ((!g252) & (sk[58]) & (g218) & (g253) & (!g220) & (g221)) + ((!g252) & (sk[58]) & (g218) & (g253) & (g220) & (g221)) + ((g252) & (!sk[58]) & (!g218) & (!g253) & (g220) & (!g221)) + ((g252) & (!sk[58]) & (!g218) & (!g253) & (g220) & (g221)) + ((g252) & (!sk[58]) & (!g218) & (g253) & (!g220) & (!g221)) + ((g252) & (!sk[58]) & (!g218) & (g253) & (!g220) & (g221)) + ((g252) & (!sk[58]) & (!g218) & (g253) & (g220) & (!g221)) + ((g252) & (!sk[58]) & (!g218) & (g253) & (g220) & (g221)) + ((g252) & (!sk[58]) & (g218) & (!g253) & (!g220) & (!g221)) + ((g252) & (!sk[58]) & (g218) & (!g253) & (!g220) & (g221)) + ((g252) & (!sk[58]) & (g218) & (!g253) & (g220) & (!g221)) + ((g252) & (!sk[58]) & (g218) & (!g253) & (g220) & (g221)) + ((g252) & (!sk[58]) & (g218) & (g253) & (!g220) & (!g221)) + ((g252) & (!sk[58]) & (g218) & (g253) & (!g220) & (g221)) + ((g252) & (!sk[58]) & (g218) & (g253) & (g220) & (!g221)) + ((g252) & (!sk[58]) & (g218) & (g253) & (g220) & (g221)) + ((g252) & (sk[58]) & (!g218) & (!g253) & (!g220) & (g221)) + ((g252) & (sk[58]) & (g218) & (!g253) & (!g220) & (g221)) + ((g252) & (sk[58]) & (g218) & (!g253) & (g220) & (!g221)) + ((g252) & (sk[58]) & (g218) & (!g253) & (g220) & (g221)) + ((g252) & (sk[58]) & (g218) & (g253) & (!g220) & (!g221)) + ((g252) & (sk[58]) & (g218) & (g253) & (!g220) & (g221)) + ((g252) & (sk[58]) & (g218) & (g253) & (g220) & (!g221)) + ((g252) & (sk[58]) & (g218) & (g253) & (g220) & (g221)));
	assign g689 = (((!g301) & (g251) & (!sk[59]) & (!g302)) + ((!g301) & (g251) & (!sk[59]) & (g302)) + ((!g301) & (g251) & (sk[59]) & (!g302)) + ((g301) & (!g251) & (sk[59]) & (!g302)) + ((g301) & (g251) & (!sk[59]) & (!g302)) + ((g301) & (g251) & (!sk[59]) & (g302)) + ((g301) & (g251) & (sk[59]) & (!g302)));
	assign g690 = (((!sk[60]) & (!g202) & (!g69) & (!g689) & (g303)) + ((!sk[60]) & (!g202) & (!g69) & (g689) & (g303)) + ((!sk[60]) & (!g202) & (g69) & (!g689) & (g303)) + ((!sk[60]) & (!g202) & (g69) & (g689) & (g303)) + ((!sk[60]) & (g202) & (!g69) & (!g689) & (!g303)) + ((!sk[60]) & (g202) & (!g69) & (!g689) & (g303)) + ((!sk[60]) & (g202) & (!g69) & (g689) & (!g303)) + ((!sk[60]) & (g202) & (!g69) & (g689) & (g303)) + ((!sk[60]) & (g202) & (g69) & (!g689) & (!g303)) + ((!sk[60]) & (g202) & (g69) & (!g689) & (g303)) + ((!sk[60]) & (g202) & (g69) & (g689) & (!g303)) + ((!sk[60]) & (g202) & (g69) & (g689) & (g303)) + ((sk[60]) & (!g202) & (!g69) & (!g689) & (g303)) + ((sk[60]) & (!g202) & (!g69) & (g689) & (!g303)) + ((sk[60]) & (!g202) & (g69) & (g689) & (!g303)) + ((sk[60]) & (!g202) & (g69) & (g689) & (g303)) + ((sk[60]) & (g202) & (!g69) & (!g689) & (!g303)) + ((sk[60]) & (g202) & (!g69) & (g689) & (g303)) + ((sk[60]) & (g202) & (g69) & (g689) & (!g303)) + ((sk[60]) & (g202) & (g69) & (g689) & (g303)));
	assign g691 = (((!sk[61]) & (!g687) & (g688) & (!g690)) + ((!sk[61]) & (!g687) & (g688) & (g690)) + ((!sk[61]) & (g687) & (g688) & (!g690)) + ((!sk[61]) & (g687) & (g688) & (g690)) + ((sk[61]) & (!g687) & (!g688) & (!g690)) + ((sk[61]) & (!g687) & (g688) & (!g690)) + ((sk[61]) & (!g687) & (g688) & (g690)) + ((sk[61]) & (g687) & (g688) & (!g690)));
	assign g692 = (((!sk[62]) & (!g252) & (!g218) & (!g220) & (g221)) + ((!sk[62]) & (!g252) & (!g218) & (g220) & (g221)) + ((!sk[62]) & (!g252) & (g218) & (!g220) & (g221)) + ((!sk[62]) & (!g252) & (g218) & (g220) & (g221)) + ((!sk[62]) & (g252) & (!g218) & (!g220) & (!g221)) + ((!sk[62]) & (g252) & (!g218) & (!g220) & (g221)) + ((!sk[62]) & (g252) & (!g218) & (g220) & (!g221)) + ((!sk[62]) & (g252) & (!g218) & (g220) & (g221)) + ((!sk[62]) & (g252) & (g218) & (!g220) & (!g221)) + ((!sk[62]) & (g252) & (g218) & (!g220) & (g221)) + ((!sk[62]) & (g252) & (g218) & (g220) & (!g221)) + ((!sk[62]) & (g252) & (g218) & (g220) & (g221)) + ((sk[62]) & (!g252) & (!g218) & (!g220) & (g221)) + ((sk[62]) & (!g252) & (!g218) & (g220) & (g221)) + ((sk[62]) & (!g252) & (g218) & (!g220) & (g221)) + ((sk[62]) & (!g252) & (g218) & (g220) & (g221)) + ((sk[62]) & (g252) & (!g218) & (g220) & (g221)) + ((sk[62]) & (g252) & (g218) & (!g220) & (!g221)) + ((sk[62]) & (g252) & (g218) & (!g220) & (g221)) + ((sk[62]) & (g252) & (g218) & (g220) & (g221)));
	assign g693 = (((!g202) & (!sk[63]) & (!g69) & (!g689) & (g303)) + ((!g202) & (!sk[63]) & (!g69) & (g689) & (g303)) + ((!g202) & (!sk[63]) & (g69) & (!g689) & (g303)) + ((!g202) & (!sk[63]) & (g69) & (g689) & (g303)) + ((!g202) & (sk[63]) & (!g69) & (!g689) & (g303)) + ((g202) & (!sk[63]) & (!g69) & (!g689) & (!g303)) + ((g202) & (!sk[63]) & (!g69) & (!g689) & (g303)) + ((g202) & (!sk[63]) & (!g69) & (g689) & (!g303)) + ((g202) & (!sk[63]) & (!g69) & (g689) & (g303)) + ((g202) & (!sk[63]) & (g69) & (!g689) & (!g303)) + ((g202) & (!sk[63]) & (g69) & (!g689) & (g303)) + ((g202) & (!sk[63]) & (g69) & (g689) & (!g303)) + ((g202) & (!sk[63]) & (g69) & (g689) & (g303)) + ((g202) & (sk[63]) & (!g69) & (!g689) & (!g303)) + ((g202) & (sk[63]) & (!g69) & (!g689) & (g303)) + ((g202) & (sk[63]) & (!g69) & (g689) & (g303)));
	assign g694 = (((!sk[64]) & (!g69) & (!g253) & (!g692) & (g693)) + ((!sk[64]) & (!g69) & (!g253) & (g692) & (g693)) + ((!sk[64]) & (!g69) & (g253) & (!g692) & (g693)) + ((!sk[64]) & (!g69) & (g253) & (g692) & (g693)) + ((!sk[64]) & (g69) & (!g253) & (!g692) & (!g693)) + ((!sk[64]) & (g69) & (!g253) & (!g692) & (g693)) + ((!sk[64]) & (g69) & (!g253) & (g692) & (!g693)) + ((!sk[64]) & (g69) & (!g253) & (g692) & (g693)) + ((!sk[64]) & (g69) & (g253) & (!g692) & (!g693)) + ((!sk[64]) & (g69) & (g253) & (!g692) & (g693)) + ((!sk[64]) & (g69) & (g253) & (g692) & (!g693)) + ((!sk[64]) & (g69) & (g253) & (g692) & (g693)) + ((sk[64]) & (!g69) & (!g253) & (!g692) & (g693)) + ((sk[64]) & (!g69) & (!g253) & (g692) & (!g693)) + ((sk[64]) & (!g69) & (g253) & (!g692) & (!g693)) + ((sk[64]) & (!g69) & (g253) & (g692) & (g693)) + ((sk[64]) & (g69) & (!g253) & (!g692) & (g693)) + ((sk[64]) & (g69) & (!g253) & (g692) & (!g693)) + ((sk[64]) & (g69) & (g253) & (!g692) & (g693)) + ((sk[64]) & (g69) & (g253) & (g692) & (!g693)));
	assign g695 = (((!g691) & (sk[65]) & (g694)) + ((g691) & (!sk[65]) & (g694)) + ((g691) & (sk[65]) & (!g694)));
	assign g696 = (((!sk[66]) & (!g317) & (g318) & (!g321)) + ((!sk[66]) & (!g317) & (g318) & (g321)) + ((!sk[66]) & (g317) & (g318) & (!g321)) + ((!sk[66]) & (g317) & (g318) & (g321)) + ((sk[66]) & (!g317) & (g318) & (!g321)) + ((sk[66]) & (g317) & (!g318) & (!g321)) + ((sk[66]) & (g317) & (g318) & (!g321)) + ((sk[66]) & (g317) & (g318) & (g321)));
	assign g697 = (((!g687) & (!g688) & (sk[67]) & (!g690)) + ((!g687) & (g688) & (!sk[67]) & (!g690)) + ((!g687) & (g688) & (!sk[67]) & (g690)) + ((!g687) & (g688) & (sk[67]) & (g690)) + ((g687) & (!g688) & (sk[67]) & (g690)) + ((g687) & (g688) & (!sk[67]) & (!g690)) + ((g687) & (g688) & (!sk[67]) & (g690)) + ((g687) & (g688) & (sk[67]) & (!g690)));
	assign g698 = (((!g695) & (!g696) & (!g697) & (!g316) & (!g322) & (!g548)) + ((!g695) & (!g696) & (!g697) & (!g316) & (!g322) & (g548)) + ((!g695) & (!g696) & (!g697) & (!g316) & (g322) & (g548)) + ((!g695) & (!g696) & (!g697) & (g316) & (!g322) & (g548)) + ((!g695) & (!g696) & (g697) & (!g316) & (!g322) & (!g548)) + ((!g695) & (!g696) & (g697) & (!g316) & (!g322) & (g548)) + ((!g695) & (!g696) & (g697) & (!g316) & (g322) & (!g548)) + ((!g695) & (!g696) & (g697) & (!g316) & (g322) & (g548)) + ((!g695) & (!g696) & (g697) & (g316) & (!g322) & (!g548)) + ((!g695) & (!g696) & (g697) & (g316) & (!g322) & (g548)) + ((!g695) & (!g696) & (g697) & (g316) & (g322) & (!g548)) + ((!g695) & (!g696) & (g697) & (g316) & (g322) & (g548)) + ((!g695) & (g696) & (g697) & (!g316) & (!g322) & (!g548)) + ((!g695) & (g696) & (g697) & (!g316) & (!g322) & (g548)) + ((!g695) & (g696) & (g697) & (!g316) & (g322) & (g548)) + ((!g695) & (g696) & (g697) & (g316) & (!g322) & (g548)) + ((g695) & (!g696) & (!g697) & (!g316) & (g322) & (!g548)) + ((g695) & (!g696) & (!g697) & (g316) & (!g322) & (!g548)) + ((g695) & (!g696) & (!g697) & (g316) & (g322) & (!g548)) + ((g695) & (!g696) & (!g697) & (g316) & (g322) & (g548)) + ((g695) & (g696) & (!g697) & (!g316) & (!g322) & (!g548)) + ((g695) & (g696) & (!g697) & (!g316) & (!g322) & (g548)) + ((g695) & (g696) & (!g697) & (!g316) & (g322) & (!g548)) + ((g695) & (g696) & (!g697) & (!g316) & (g322) & (g548)) + ((g695) & (g696) & (!g697) & (g316) & (!g322) & (!g548)) + ((g695) & (g696) & (!g697) & (g316) & (!g322) & (g548)) + ((g695) & (g696) & (!g697) & (g316) & (g322) & (!g548)) + ((g695) & (g696) & (!g697) & (g316) & (g322) & (g548)) + ((g695) & (g696) & (g697) & (!g316) & (g322) & (!g548)) + ((g695) & (g696) & (g697) & (g316) & (!g322) & (!g548)) + ((g695) & (g696) & (g697) & (g316) & (g322) & (!g548)) + ((g695) & (g696) & (g697) & (g316) & (g322) & (g548)));
	assign g699 = (((!sk[69]) & (g275) & (g672)) + ((sk[69]) & (!g275) & (g672)));
	assign g700 = (((!g112) & (!g97) & (!sk[70]) & (!g98) & (g46)) + ((!g112) & (!g97) & (!sk[70]) & (g98) & (g46)) + ((!g112) & (!g97) & (sk[70]) & (g98) & (g46)) + ((!g112) & (g97) & (!sk[70]) & (!g98) & (g46)) + ((!g112) & (g97) & (!sk[70]) & (g98) & (g46)) + ((g112) & (!g97) & (!sk[70]) & (!g98) & (!g46)) + ((g112) & (!g97) & (!sk[70]) & (!g98) & (g46)) + ((g112) & (!g97) & (!sk[70]) & (g98) & (!g46)) + ((g112) & (!g97) & (!sk[70]) & (g98) & (g46)) + ((g112) & (g97) & (!sk[70]) & (!g98) & (!g46)) + ((g112) & (g97) & (!sk[70]) & (!g98) & (g46)) + ((g112) & (g97) & (!sk[70]) & (g98) & (!g46)) + ((g112) & (g97) & (!sk[70]) & (g98) & (g46)));
	assign g701 = (((!g70) & (!g25) & (!g354) & (!g272) & (sk[71]) & (!g700)) + ((!g70) & (!g25) & (!g354) & (g272) & (!sk[71]) & (!g700)) + ((!g70) & (!g25) & (!g354) & (g272) & (!sk[71]) & (g700)) + ((!g70) & (!g25) & (g354) & (!g272) & (!sk[71]) & (!g700)) + ((!g70) & (!g25) & (g354) & (!g272) & (!sk[71]) & (g700)) + ((!g70) & (!g25) & (g354) & (g272) & (!sk[71]) & (!g700)) + ((!g70) & (!g25) & (g354) & (g272) & (!sk[71]) & (g700)) + ((!g70) & (g25) & (!g354) & (!g272) & (!sk[71]) & (!g700)) + ((!g70) & (g25) & (!g354) & (!g272) & (!sk[71]) & (g700)) + ((!g70) & (g25) & (!g354) & (!g272) & (sk[71]) & (!g700)) + ((!g70) & (g25) & (!g354) & (g272) & (!sk[71]) & (!g700)) + ((!g70) & (g25) & (!g354) & (g272) & (!sk[71]) & (g700)) + ((!g70) & (g25) & (g354) & (!g272) & (!sk[71]) & (!g700)) + ((!g70) & (g25) & (g354) & (!g272) & (!sk[71]) & (g700)) + ((!g70) & (g25) & (g354) & (g272) & (!sk[71]) & (!g700)) + ((!g70) & (g25) & (g354) & (g272) & (!sk[71]) & (g700)) + ((g70) & (!g25) & (!g354) & (!g272) & (sk[71]) & (!g700)) + ((g70) & (!g25) & (!g354) & (g272) & (!sk[71]) & (!g700)) + ((g70) & (!g25) & (!g354) & (g272) & (!sk[71]) & (g700)) + ((g70) & (!g25) & (g354) & (!g272) & (!sk[71]) & (!g700)) + ((g70) & (!g25) & (g354) & (!g272) & (!sk[71]) & (g700)) + ((g70) & (!g25) & (g354) & (g272) & (!sk[71]) & (!g700)) + ((g70) & (!g25) & (g354) & (g272) & (!sk[71]) & (g700)) + ((g70) & (g25) & (!g354) & (!g272) & (!sk[71]) & (!g700)) + ((g70) & (g25) & (!g354) & (!g272) & (!sk[71]) & (g700)) + ((g70) & (g25) & (!g354) & (g272) & (!sk[71]) & (!g700)) + ((g70) & (g25) & (!g354) & (g272) & (!sk[71]) & (g700)) + ((g70) & (g25) & (g354) & (!g272) & (!sk[71]) & (!g700)) + ((g70) & (g25) & (g354) & (!g272) & (!sk[71]) & (g700)) + ((g70) & (g25) & (g354) & (g272) & (!sk[71]) & (!g700)) + ((g70) & (g25) & (g354) & (g272) & (!sk[71]) & (g700)));
	assign g702 = (((!g184) & (!g104) & (!g146) & (!sk[72]) & (g27)) + ((!g184) & (!g104) & (!g146) & (sk[72]) & (!g27)) + ((!g184) & (!g104) & (!g146) & (sk[72]) & (g27)) + ((!g184) & (!g104) & (g146) & (!sk[72]) & (g27)) + ((!g184) & (g104) & (!g146) & (!sk[72]) & (g27)) + ((!g184) & (g104) & (!g146) & (sk[72]) & (!g27)) + ((!g184) & (g104) & (g146) & (!sk[72]) & (g27)) + ((g184) & (!g104) & (!g146) & (!sk[72]) & (!g27)) + ((g184) & (!g104) & (!g146) & (!sk[72]) & (g27)) + ((g184) & (!g104) & (g146) & (!sk[72]) & (!g27)) + ((g184) & (!g104) & (g146) & (!sk[72]) & (g27)) + ((g184) & (g104) & (!g146) & (!sk[72]) & (!g27)) + ((g184) & (g104) & (!g146) & (!sk[72]) & (g27)) + ((g184) & (g104) & (g146) & (!sk[72]) & (!g27)) + ((g184) & (g104) & (g146) & (!sk[72]) & (g27)));
	assign g703 = (((!g105) & (!sk[73]) & (!g326) & (!g181) & (g701) & (!g702)) + ((!g105) & (!sk[73]) & (!g326) & (!g181) & (g701) & (g702)) + ((!g105) & (!sk[73]) & (!g326) & (g181) & (!g701) & (!g702)) + ((!g105) & (!sk[73]) & (!g326) & (g181) & (!g701) & (g702)) + ((!g105) & (!sk[73]) & (!g326) & (g181) & (g701) & (!g702)) + ((!g105) & (!sk[73]) & (!g326) & (g181) & (g701) & (g702)) + ((!g105) & (!sk[73]) & (g326) & (!g181) & (!g701) & (!g702)) + ((!g105) & (!sk[73]) & (g326) & (!g181) & (!g701) & (g702)) + ((!g105) & (!sk[73]) & (g326) & (!g181) & (g701) & (!g702)) + ((!g105) & (!sk[73]) & (g326) & (!g181) & (g701) & (g702)) + ((!g105) & (!sk[73]) & (g326) & (g181) & (!g701) & (!g702)) + ((!g105) & (!sk[73]) & (g326) & (g181) & (!g701) & (g702)) + ((!g105) & (!sk[73]) & (g326) & (g181) & (g701) & (!g702)) + ((!g105) & (!sk[73]) & (g326) & (g181) & (g701) & (g702)) + ((!g105) & (sk[73]) & (g326) & (g181) & (g701) & (g702)) + ((g105) & (!sk[73]) & (!g326) & (!g181) & (g701) & (!g702)) + ((g105) & (!sk[73]) & (!g326) & (!g181) & (g701) & (g702)) + ((g105) & (!sk[73]) & (!g326) & (g181) & (!g701) & (!g702)) + ((g105) & (!sk[73]) & (!g326) & (g181) & (!g701) & (g702)) + ((g105) & (!sk[73]) & (!g326) & (g181) & (g701) & (!g702)) + ((g105) & (!sk[73]) & (!g326) & (g181) & (g701) & (g702)) + ((g105) & (!sk[73]) & (g326) & (!g181) & (!g701) & (!g702)) + ((g105) & (!sk[73]) & (g326) & (!g181) & (!g701) & (g702)) + ((g105) & (!sk[73]) & (g326) & (!g181) & (g701) & (!g702)) + ((g105) & (!sk[73]) & (g326) & (!g181) & (g701) & (g702)) + ((g105) & (!sk[73]) & (g326) & (g181) & (!g701) & (!g702)) + ((g105) & (!sk[73]) & (g326) & (g181) & (!g701) & (g702)) + ((g105) & (!sk[73]) & (g326) & (g181) & (g701) & (!g702)) + ((g105) & (!sk[73]) & (g326) & (g181) & (g701) & (g702)));
	assign g704 = (((!g9) & (!g70) & (!sk[74]) & (!g18) & (g66)) + ((!g9) & (!g70) & (!sk[74]) & (g18) & (g66)) + ((!g9) & (g70) & (!sk[74]) & (!g18) & (g66)) + ((!g9) & (g70) & (!sk[74]) & (g18) & (g66)) + ((!g9) & (g70) & (sk[74]) & (g18) & (!g66)) + ((!g9) & (g70) & (sk[74]) & (g18) & (g66)) + ((g9) & (!g70) & (!sk[74]) & (!g18) & (!g66)) + ((g9) & (!g70) & (!sk[74]) & (!g18) & (g66)) + ((g9) & (!g70) & (!sk[74]) & (g18) & (!g66)) + ((g9) & (!g70) & (!sk[74]) & (g18) & (g66)) + ((g9) & (!g70) & (sk[74]) & (!g18) & (g66)) + ((g9) & (!g70) & (sk[74]) & (g18) & (g66)) + ((g9) & (g70) & (!sk[74]) & (!g18) & (!g66)) + ((g9) & (g70) & (!sk[74]) & (!g18) & (g66)) + ((g9) & (g70) & (!sk[74]) & (g18) & (!g66)) + ((g9) & (g70) & (!sk[74]) & (g18) & (g66)) + ((g9) & (g70) & (sk[74]) & (!g18) & (g66)) + ((g9) & (g70) & (sk[74]) & (g18) & (!g66)) + ((g9) & (g70) & (sk[74]) & (g18) & (g66)));
	assign g705 = (((!sk[75]) & (!g48) & (!g296) & (!g331) & (g225) & (!g704)) + ((!sk[75]) & (!g48) & (!g296) & (!g331) & (g225) & (g704)) + ((!sk[75]) & (!g48) & (!g296) & (g331) & (!g225) & (!g704)) + ((!sk[75]) & (!g48) & (!g296) & (g331) & (!g225) & (g704)) + ((!sk[75]) & (!g48) & (!g296) & (g331) & (g225) & (!g704)) + ((!sk[75]) & (!g48) & (!g296) & (g331) & (g225) & (g704)) + ((!sk[75]) & (!g48) & (g296) & (!g331) & (!g225) & (!g704)) + ((!sk[75]) & (!g48) & (g296) & (!g331) & (!g225) & (g704)) + ((!sk[75]) & (!g48) & (g296) & (!g331) & (g225) & (!g704)) + ((!sk[75]) & (!g48) & (g296) & (!g331) & (g225) & (g704)) + ((!sk[75]) & (!g48) & (g296) & (g331) & (!g225) & (!g704)) + ((!sk[75]) & (!g48) & (g296) & (g331) & (!g225) & (g704)) + ((!sk[75]) & (!g48) & (g296) & (g331) & (g225) & (!g704)) + ((!sk[75]) & (!g48) & (g296) & (g331) & (g225) & (g704)) + ((!sk[75]) & (g48) & (!g296) & (!g331) & (g225) & (!g704)) + ((!sk[75]) & (g48) & (!g296) & (!g331) & (g225) & (g704)) + ((!sk[75]) & (g48) & (!g296) & (g331) & (!g225) & (!g704)) + ((!sk[75]) & (g48) & (!g296) & (g331) & (!g225) & (g704)) + ((!sk[75]) & (g48) & (!g296) & (g331) & (g225) & (!g704)) + ((!sk[75]) & (g48) & (!g296) & (g331) & (g225) & (g704)) + ((!sk[75]) & (g48) & (g296) & (!g331) & (!g225) & (!g704)) + ((!sk[75]) & (g48) & (g296) & (!g331) & (!g225) & (g704)) + ((!sk[75]) & (g48) & (g296) & (!g331) & (g225) & (!g704)) + ((!sk[75]) & (g48) & (g296) & (!g331) & (g225) & (g704)) + ((!sk[75]) & (g48) & (g296) & (g331) & (!g225) & (!g704)) + ((!sk[75]) & (g48) & (g296) & (g331) & (!g225) & (g704)) + ((!sk[75]) & (g48) & (g296) & (g331) & (g225) & (!g704)) + ((!sk[75]) & (g48) & (g296) & (g331) & (g225) & (g704)) + ((sk[75]) & (g48) & (g296) & (!g331) & (g225) & (!g704)));
	assign g706 = (((!g699) & (!g117) & (!sk[76]) & (!g703) & (g574) & (!g705)) + ((!g699) & (!g117) & (!sk[76]) & (!g703) & (g574) & (g705)) + ((!g699) & (!g117) & (!sk[76]) & (g703) & (!g574) & (!g705)) + ((!g699) & (!g117) & (!sk[76]) & (g703) & (!g574) & (g705)) + ((!g699) & (!g117) & (!sk[76]) & (g703) & (g574) & (!g705)) + ((!g699) & (!g117) & (!sk[76]) & (g703) & (g574) & (g705)) + ((!g699) & (g117) & (!sk[76]) & (!g703) & (!g574) & (!g705)) + ((!g699) & (g117) & (!sk[76]) & (!g703) & (!g574) & (g705)) + ((!g699) & (g117) & (!sk[76]) & (!g703) & (g574) & (!g705)) + ((!g699) & (g117) & (!sk[76]) & (!g703) & (g574) & (g705)) + ((!g699) & (g117) & (!sk[76]) & (g703) & (!g574) & (!g705)) + ((!g699) & (g117) & (!sk[76]) & (g703) & (!g574) & (g705)) + ((!g699) & (g117) & (!sk[76]) & (g703) & (g574) & (!g705)) + ((!g699) & (g117) & (!sk[76]) & (g703) & (g574) & (g705)) + ((g699) & (!g117) & (!sk[76]) & (!g703) & (g574) & (!g705)) + ((g699) & (!g117) & (!sk[76]) & (!g703) & (g574) & (g705)) + ((g699) & (!g117) & (!sk[76]) & (g703) & (!g574) & (!g705)) + ((g699) & (!g117) & (!sk[76]) & (g703) & (!g574) & (g705)) + ((g699) & (!g117) & (!sk[76]) & (g703) & (g574) & (!g705)) + ((g699) & (!g117) & (!sk[76]) & (g703) & (g574) & (g705)) + ((g699) & (!g117) & (sk[76]) & (g703) & (g574) & (g705)) + ((g699) & (g117) & (!sk[76]) & (!g703) & (!g574) & (!g705)) + ((g699) & (g117) & (!sk[76]) & (!g703) & (!g574) & (g705)) + ((g699) & (g117) & (!sk[76]) & (!g703) & (g574) & (!g705)) + ((g699) & (g117) & (!sk[76]) & (!g703) & (g574) & (g705)) + ((g699) & (g117) & (!sk[76]) & (g703) & (!g574) & (!g705)) + ((g699) & (g117) & (!sk[76]) & (g703) & (!g574) & (g705)) + ((g699) & (g117) & (!sk[76]) & (g703) & (g574) & (!g705)) + ((g699) & (g117) & (!sk[76]) & (g703) & (g574) & (g705)));
	assign g707 = (((!g698) & (sk[77]) & (!g706)) + ((g698) & (!sk[77]) & (g706)) + ((g698) & (sk[77]) & (g706)));
	assign g708 = (((!g696) & (!g697) & (!g316) & (!sk[78]) & (g322) & (!g548)) + ((!g696) & (!g697) & (!g316) & (!sk[78]) & (g322) & (g548)) + ((!g696) & (!g697) & (!g316) & (sk[78]) & (!g322) & (!g548)) + ((!g696) & (!g697) & (!g316) & (sk[78]) & (!g322) & (g548)) + ((!g696) & (!g697) & (!g316) & (sk[78]) & (g322) & (g548)) + ((!g696) & (!g697) & (g316) & (!sk[78]) & (!g322) & (!g548)) + ((!g696) & (!g697) & (g316) & (!sk[78]) & (!g322) & (g548)) + ((!g696) & (!g697) & (g316) & (!sk[78]) & (g322) & (!g548)) + ((!g696) & (!g697) & (g316) & (!sk[78]) & (g322) & (g548)) + ((!g696) & (!g697) & (g316) & (sk[78]) & (!g322) & (g548)) + ((!g696) & (g697) & (!g316) & (!sk[78]) & (!g322) & (!g548)) + ((!g696) & (g697) & (!g316) & (!sk[78]) & (!g322) & (g548)) + ((!g696) & (g697) & (!g316) & (!sk[78]) & (g322) & (!g548)) + ((!g696) & (g697) & (!g316) & (!sk[78]) & (g322) & (g548)) + ((!g696) & (g697) & (!g316) & (sk[78]) & (g322) & (!g548)) + ((!g696) & (g697) & (g316) & (!sk[78]) & (!g322) & (!g548)) + ((!g696) & (g697) & (g316) & (!sk[78]) & (!g322) & (g548)) + ((!g696) & (g697) & (g316) & (!sk[78]) & (g322) & (!g548)) + ((!g696) & (g697) & (g316) & (!sk[78]) & (g322) & (g548)) + ((!g696) & (g697) & (g316) & (sk[78]) & (!g322) & (!g548)) + ((!g696) & (g697) & (g316) & (sk[78]) & (g322) & (!g548)) + ((!g696) & (g697) & (g316) & (sk[78]) & (g322) & (g548)) + ((g696) & (!g697) & (!g316) & (!sk[78]) & (g322) & (!g548)) + ((g696) & (!g697) & (!g316) & (!sk[78]) & (g322) & (g548)) + ((g696) & (!g697) & (!g316) & (sk[78]) & (g322) & (!g548)) + ((g696) & (!g697) & (g316) & (!sk[78]) & (!g322) & (!g548)) + ((g696) & (!g697) & (g316) & (!sk[78]) & (!g322) & (g548)) + ((g696) & (!g697) & (g316) & (!sk[78]) & (g322) & (!g548)) + ((g696) & (!g697) & (g316) & (!sk[78]) & (g322) & (g548)) + ((g696) & (!g697) & (g316) & (sk[78]) & (!g322) & (!g548)) + ((g696) & (!g697) & (g316) & (sk[78]) & (g322) & (!g548)) + ((g696) & (!g697) & (g316) & (sk[78]) & (g322) & (g548)) + ((g696) & (g697) & (!g316) & (!sk[78]) & (!g322) & (!g548)) + ((g696) & (g697) & (!g316) & (!sk[78]) & (!g322) & (g548)) + ((g696) & (g697) & (!g316) & (!sk[78]) & (g322) & (!g548)) + ((g696) & (g697) & (!g316) & (!sk[78]) & (g322) & (g548)) + ((g696) & (g697) & (!g316) & (sk[78]) & (!g322) & (!g548)) + ((g696) & (g697) & (!g316) & (sk[78]) & (!g322) & (g548)) + ((g696) & (g697) & (!g316) & (sk[78]) & (g322) & (g548)) + ((g696) & (g697) & (g316) & (!sk[78]) & (!g322) & (!g548)) + ((g696) & (g697) & (g316) & (!sk[78]) & (!g322) & (g548)) + ((g696) & (g697) & (g316) & (!sk[78]) & (g322) & (!g548)) + ((g696) & (g697) & (g316) & (!sk[78]) & (g322) & (g548)) + ((g696) & (g697) & (g316) & (sk[78]) & (!g322) & (g548)));
	assign g709 = (((!g572) & (!g171) & (sk[79]) & (g330)) + ((!g572) & (g171) & (!sk[79]) & (!g330)) + ((!g572) & (g171) & (!sk[79]) & (g330)) + ((g572) & (g171) & (!sk[79]) & (!g330)) + ((g572) & (g171) & (!sk[79]) & (g330)));
	assign g710 = (((!g70) & (!g71) & (!sk[80]) & (!g25) & (g27)) + ((!g70) & (!g71) & (!sk[80]) & (g25) & (g27)) + ((!g70) & (g71) & (!sk[80]) & (!g25) & (g27)) + ((!g70) & (g71) & (!sk[80]) & (g25) & (g27)) + ((!g70) & (g71) & (sk[80]) & (g25) & (!g27)) + ((!g70) & (g71) & (sk[80]) & (g25) & (g27)) + ((g70) & (!g71) & (!sk[80]) & (!g25) & (!g27)) + ((g70) & (!g71) & (!sk[80]) & (!g25) & (g27)) + ((g70) & (!g71) & (!sk[80]) & (g25) & (!g27)) + ((g70) & (!g71) & (!sk[80]) & (g25) & (g27)) + ((g70) & (!g71) & (sk[80]) & (!g25) & (g27)) + ((g70) & (!g71) & (sk[80]) & (g25) & (g27)) + ((g70) & (g71) & (!sk[80]) & (!g25) & (!g27)) + ((g70) & (g71) & (!sk[80]) & (!g25) & (g27)) + ((g70) & (g71) & (!sk[80]) & (g25) & (!g27)) + ((g70) & (g71) & (!sk[80]) & (g25) & (g27)) + ((g70) & (g71) & (sk[80]) & (!g25) & (g27)) + ((g70) & (g71) & (sk[80]) & (g25) & (!g27)) + ((g70) & (g71) & (sk[80]) & (g25) & (g27)));
	assign g711 = (((!g16) & (!g99) & (!g25) & (!g47) & (!g66) & (!g187)) + ((!g16) & (!g99) & (!g25) & (!g47) & (g66) & (!g187)) + ((!g16) & (!g99) & (g25) & (!g47) & (!g66) & (!g187)) + ((!g16) & (!g99) & (g25) & (!g47) & (g66) & (!g187)) + ((!g16) & (g99) & (!g25) & (!g47) & (!g66) & (!g187)) + ((!g16) & (g99) & (!g25) & (!g47) & (g66) & (!g187)) + ((g16) & (!g99) & (!g25) & (!g47) & (!g66) & (!g187)) + ((g16) & (!g99) & (g25) & (!g47) & (!g66) & (!g187)) + ((g16) & (g99) & (!g25) & (!g47) & (!g66) & (!g187)));
	assign g712 = (((!g38) & (!g9) & (!g99) & (!g40) & (sk[82]) & (!g66)) + ((!g38) & (!g9) & (!g99) & (!g40) & (sk[82]) & (g66)) + ((!g38) & (!g9) & (!g99) & (g40) & (!sk[82]) & (!g66)) + ((!g38) & (!g9) & (!g99) & (g40) & (!sk[82]) & (g66)) + ((!g38) & (!g9) & (!g99) & (g40) & (sk[82]) & (!g66)) + ((!g38) & (!g9) & (!g99) & (g40) & (sk[82]) & (g66)) + ((!g38) & (!g9) & (g99) & (!g40) & (!sk[82]) & (!g66)) + ((!g38) & (!g9) & (g99) & (!g40) & (!sk[82]) & (g66)) + ((!g38) & (!g9) & (g99) & (!g40) & (sk[82]) & (!g66)) + ((!g38) & (!g9) & (g99) & (g40) & (!sk[82]) & (!g66)) + ((!g38) & (!g9) & (g99) & (g40) & (!sk[82]) & (g66)) + ((!g38) & (g9) & (!g99) & (!g40) & (!sk[82]) & (!g66)) + ((!g38) & (g9) & (!g99) & (!g40) & (!sk[82]) & (g66)) + ((!g38) & (g9) & (!g99) & (!g40) & (sk[82]) & (!g66)) + ((!g38) & (g9) & (!g99) & (!g40) & (sk[82]) & (g66)) + ((!g38) & (g9) & (!g99) & (g40) & (!sk[82]) & (!g66)) + ((!g38) & (g9) & (!g99) & (g40) & (!sk[82]) & (g66)) + ((!g38) & (g9) & (g99) & (!g40) & (!sk[82]) & (!g66)) + ((!g38) & (g9) & (g99) & (!g40) & (!sk[82]) & (g66)) + ((!g38) & (g9) & (g99) & (!g40) & (sk[82]) & (!g66)) + ((!g38) & (g9) & (g99) & (g40) & (!sk[82]) & (!g66)) + ((!g38) & (g9) & (g99) & (g40) & (!sk[82]) & (g66)) + ((g38) & (!g9) & (!g99) & (!g40) & (sk[82]) & (!g66)) + ((g38) & (!g9) & (!g99) & (!g40) & (sk[82]) & (g66)) + ((g38) & (!g9) & (!g99) & (g40) & (!sk[82]) & (!g66)) + ((g38) & (!g9) & (!g99) & (g40) & (!sk[82]) & (g66)) + ((g38) & (!g9) & (!g99) & (g40) & (sk[82]) & (!g66)) + ((g38) & (!g9) & (!g99) & (g40) & (sk[82]) & (g66)) + ((g38) & (!g9) & (g99) & (!g40) & (!sk[82]) & (!g66)) + ((g38) & (!g9) & (g99) & (!g40) & (!sk[82]) & (g66)) + ((g38) & (!g9) & (g99) & (g40) & (!sk[82]) & (!g66)) + ((g38) & (!g9) & (g99) & (g40) & (!sk[82]) & (g66)) + ((g38) & (g9) & (!g99) & (!g40) & (!sk[82]) & (!g66)) + ((g38) & (g9) & (!g99) & (!g40) & (!sk[82]) & (g66)) + ((g38) & (g9) & (!g99) & (!g40) & (sk[82]) & (!g66)) + ((g38) & (g9) & (!g99) & (!g40) & (sk[82]) & (g66)) + ((g38) & (g9) & (!g99) & (g40) & (!sk[82]) & (!g66)) + ((g38) & (g9) & (!g99) & (g40) & (!sk[82]) & (g66)) + ((g38) & (g9) & (g99) & (!g40) & (!sk[82]) & (!g66)) + ((g38) & (g9) & (g99) & (!g40) & (!sk[82]) & (g66)) + ((g38) & (g9) & (g99) & (g40) & (!sk[82]) & (!g66)) + ((g38) & (g9) & (g99) & (g40) & (!sk[82]) & (g66)));
	assign g713 = (((!sk[83]) & (!g98) & (!g99) & (!g100) & (g62) & (!g32)) + ((!sk[83]) & (!g98) & (!g99) & (!g100) & (g62) & (g32)) + ((!sk[83]) & (!g98) & (!g99) & (g100) & (!g62) & (!g32)) + ((!sk[83]) & (!g98) & (!g99) & (g100) & (!g62) & (g32)) + ((!sk[83]) & (!g98) & (!g99) & (g100) & (g62) & (!g32)) + ((!sk[83]) & (!g98) & (!g99) & (g100) & (g62) & (g32)) + ((!sk[83]) & (!g98) & (g99) & (!g100) & (!g62) & (!g32)) + ((!sk[83]) & (!g98) & (g99) & (!g100) & (!g62) & (g32)) + ((!sk[83]) & (!g98) & (g99) & (!g100) & (g62) & (!g32)) + ((!sk[83]) & (!g98) & (g99) & (!g100) & (g62) & (g32)) + ((!sk[83]) & (!g98) & (g99) & (g100) & (!g62) & (!g32)) + ((!sk[83]) & (!g98) & (g99) & (g100) & (!g62) & (g32)) + ((!sk[83]) & (!g98) & (g99) & (g100) & (g62) & (!g32)) + ((!sk[83]) & (!g98) & (g99) & (g100) & (g62) & (g32)) + ((!sk[83]) & (g98) & (!g99) & (!g100) & (g62) & (!g32)) + ((!sk[83]) & (g98) & (!g99) & (!g100) & (g62) & (g32)) + ((!sk[83]) & (g98) & (!g99) & (g100) & (!g62) & (!g32)) + ((!sk[83]) & (g98) & (!g99) & (g100) & (!g62) & (g32)) + ((!sk[83]) & (g98) & (!g99) & (g100) & (g62) & (!g32)) + ((!sk[83]) & (g98) & (!g99) & (g100) & (g62) & (g32)) + ((!sk[83]) & (g98) & (g99) & (!g100) & (!g62) & (!g32)) + ((!sk[83]) & (g98) & (g99) & (!g100) & (!g62) & (g32)) + ((!sk[83]) & (g98) & (g99) & (!g100) & (g62) & (!g32)) + ((!sk[83]) & (g98) & (g99) & (!g100) & (g62) & (g32)) + ((!sk[83]) & (g98) & (g99) & (g100) & (!g62) & (!g32)) + ((!sk[83]) & (g98) & (g99) & (g100) & (!g62) & (g32)) + ((!sk[83]) & (g98) & (g99) & (g100) & (g62) & (!g32)) + ((!sk[83]) & (g98) & (g99) & (g100) & (g62) & (g32)) + ((sk[83]) & (!g98) & (g99) & (!g100) & (!g62) & (g32)) + ((sk[83]) & (!g98) & (g99) & (!g100) & (g62) & (g32)) + ((sk[83]) & (!g98) & (g99) & (g100) & (!g62) & (g32)) + ((sk[83]) & (!g98) & (g99) & (g100) & (g62) & (g32)) + ((sk[83]) & (g98) & (!g99) & (g100) & (g62) & (!g32)) + ((sk[83]) & (g98) & (!g99) & (g100) & (g62) & (g32)) + ((sk[83]) & (g98) & (g99) & (!g100) & (!g62) & (g32)) + ((sk[83]) & (g98) & (g99) & (!g100) & (g62) & (g32)) + ((sk[83]) & (g98) & (g99) & (g100) & (!g62) & (g32)) + ((sk[83]) & (g98) & (g99) & (g100) & (g62) & (!g32)) + ((sk[83]) & (g98) & (g99) & (g100) & (g62) & (g32)));
	assign g714 = (((!g58) & (!sk[84]) & (!g104) & (!g25) & (g101) & (!g713)) + ((!g58) & (!sk[84]) & (!g104) & (!g25) & (g101) & (g713)) + ((!g58) & (!sk[84]) & (!g104) & (g25) & (!g101) & (!g713)) + ((!g58) & (!sk[84]) & (!g104) & (g25) & (!g101) & (g713)) + ((!g58) & (!sk[84]) & (!g104) & (g25) & (g101) & (!g713)) + ((!g58) & (!sk[84]) & (!g104) & (g25) & (g101) & (g713)) + ((!g58) & (!sk[84]) & (g104) & (!g25) & (!g101) & (!g713)) + ((!g58) & (!sk[84]) & (g104) & (!g25) & (!g101) & (g713)) + ((!g58) & (!sk[84]) & (g104) & (!g25) & (g101) & (!g713)) + ((!g58) & (!sk[84]) & (g104) & (!g25) & (g101) & (g713)) + ((!g58) & (!sk[84]) & (g104) & (g25) & (!g101) & (!g713)) + ((!g58) & (!sk[84]) & (g104) & (g25) & (!g101) & (g713)) + ((!g58) & (!sk[84]) & (g104) & (g25) & (g101) & (!g713)) + ((!g58) & (!sk[84]) & (g104) & (g25) & (g101) & (g713)) + ((!g58) & (sk[84]) & (!g104) & (!g25) & (!g101) & (!g713)) + ((!g58) & (sk[84]) & (!g104) & (g25) & (!g101) & (!g713)) + ((!g58) & (sk[84]) & (g104) & (!g25) & (!g101) & (!g713)) + ((g58) & (!sk[84]) & (!g104) & (!g25) & (g101) & (!g713)) + ((g58) & (!sk[84]) & (!g104) & (!g25) & (g101) & (g713)) + ((g58) & (!sk[84]) & (!g104) & (g25) & (!g101) & (!g713)) + ((g58) & (!sk[84]) & (!g104) & (g25) & (!g101) & (g713)) + ((g58) & (!sk[84]) & (!g104) & (g25) & (g101) & (!g713)) + ((g58) & (!sk[84]) & (!g104) & (g25) & (g101) & (g713)) + ((g58) & (!sk[84]) & (g104) & (!g25) & (!g101) & (!g713)) + ((g58) & (!sk[84]) & (g104) & (!g25) & (!g101) & (g713)) + ((g58) & (!sk[84]) & (g104) & (!g25) & (g101) & (!g713)) + ((g58) & (!sk[84]) & (g104) & (!g25) & (g101) & (g713)) + ((g58) & (!sk[84]) & (g104) & (g25) & (!g101) & (!g713)) + ((g58) & (!sk[84]) & (g104) & (g25) & (!g101) & (g713)) + ((g58) & (!sk[84]) & (g104) & (g25) & (g101) & (!g713)) + ((g58) & (!sk[84]) & (g104) & (g25) & (g101) & (g713)) + ((g58) & (sk[84]) & (!g104) & (!g25) & (!g101) & (!g713)) + ((g58) & (sk[84]) & (!g104) & (g25) & (!g101) & (!g713)));
	assign g715 = (((!g39) & (!g710) & (!g711) & (g712) & (!sk[85]) & (!g714)) + ((!g39) & (!g710) & (!g711) & (g712) & (!sk[85]) & (g714)) + ((!g39) & (!g710) & (g711) & (!g712) & (!sk[85]) & (!g714)) + ((!g39) & (!g710) & (g711) & (!g712) & (!sk[85]) & (g714)) + ((!g39) & (!g710) & (g711) & (g712) & (!sk[85]) & (!g714)) + ((!g39) & (!g710) & (g711) & (g712) & (!sk[85]) & (g714)) + ((!g39) & (g710) & (!g711) & (!g712) & (!sk[85]) & (!g714)) + ((!g39) & (g710) & (!g711) & (!g712) & (!sk[85]) & (g714)) + ((!g39) & (g710) & (!g711) & (g712) & (!sk[85]) & (!g714)) + ((!g39) & (g710) & (!g711) & (g712) & (!sk[85]) & (g714)) + ((!g39) & (g710) & (g711) & (!g712) & (!sk[85]) & (!g714)) + ((!g39) & (g710) & (g711) & (!g712) & (!sk[85]) & (g714)) + ((!g39) & (g710) & (g711) & (g712) & (!sk[85]) & (!g714)) + ((!g39) & (g710) & (g711) & (g712) & (!sk[85]) & (g714)) + ((g39) & (!g710) & (!g711) & (g712) & (!sk[85]) & (!g714)) + ((g39) & (!g710) & (!g711) & (g712) & (!sk[85]) & (g714)) + ((g39) & (!g710) & (g711) & (!g712) & (!sk[85]) & (!g714)) + ((g39) & (!g710) & (g711) & (!g712) & (!sk[85]) & (g714)) + ((g39) & (!g710) & (g711) & (g712) & (!sk[85]) & (!g714)) + ((g39) & (!g710) & (g711) & (g712) & (!sk[85]) & (g714)) + ((g39) & (!g710) & (g711) & (g712) & (sk[85]) & (g714)) + ((g39) & (g710) & (!g711) & (!g712) & (!sk[85]) & (!g714)) + ((g39) & (g710) & (!g711) & (!g712) & (!sk[85]) & (g714)) + ((g39) & (g710) & (!g711) & (g712) & (!sk[85]) & (!g714)) + ((g39) & (g710) & (!g711) & (g712) & (!sk[85]) & (g714)) + ((g39) & (g710) & (g711) & (!g712) & (!sk[85]) & (!g714)) + ((g39) & (g710) & (g711) & (!g712) & (!sk[85]) & (g714)) + ((g39) & (g710) & (g711) & (g712) & (!sk[85]) & (!g714)) + ((g39) & (g710) & (g711) & (g712) & (!sk[85]) & (g714)));
	assign g716 = (((!g286) & (!g145) & (!g709) & (!sk[86]) & (g715)) + ((!g286) & (!g145) & (g709) & (!sk[86]) & (g715)) + ((!g286) & (g145) & (!g709) & (!sk[86]) & (g715)) + ((!g286) & (g145) & (g709) & (!sk[86]) & (g715)) + ((g286) & (!g145) & (!g709) & (!sk[86]) & (!g715)) + ((g286) & (!g145) & (!g709) & (!sk[86]) & (g715)) + ((g286) & (!g145) & (g709) & (!sk[86]) & (!g715)) + ((g286) & (!g145) & (g709) & (!sk[86]) & (g715)) + ((g286) & (g145) & (!g709) & (!sk[86]) & (!g715)) + ((g286) & (g145) & (!g709) & (!sk[86]) & (g715)) + ((g286) & (g145) & (g709) & (!sk[86]) & (!g715)) + ((g286) & (g145) & (g709) & (!sk[86]) & (g715)) + ((g286) & (g145) & (g709) & (sk[86]) & (g715)));
	assign g717 = (((!g708) & (!sk[87]) & (!g716) & (!g549) & (g569) & (!g680)) + ((!g708) & (!sk[87]) & (!g716) & (!g549) & (g569) & (g680)) + ((!g708) & (!sk[87]) & (!g716) & (g549) & (!g569) & (!g680)) + ((!g708) & (!sk[87]) & (!g716) & (g549) & (!g569) & (g680)) + ((!g708) & (!sk[87]) & (!g716) & (g549) & (g569) & (!g680)) + ((!g708) & (!sk[87]) & (!g716) & (g549) & (g569) & (g680)) + ((!g708) & (!sk[87]) & (g716) & (!g549) & (!g569) & (!g680)) + ((!g708) & (!sk[87]) & (g716) & (!g549) & (!g569) & (g680)) + ((!g708) & (!sk[87]) & (g716) & (!g549) & (g569) & (!g680)) + ((!g708) & (!sk[87]) & (g716) & (!g549) & (g569) & (g680)) + ((!g708) & (!sk[87]) & (g716) & (g549) & (!g569) & (!g680)) + ((!g708) & (!sk[87]) & (g716) & (g549) & (!g569) & (g680)) + ((!g708) & (!sk[87]) & (g716) & (g549) & (g569) & (!g680)) + ((!g708) & (!sk[87]) & (g716) & (g549) & (g569) & (g680)) + ((!g708) & (sk[87]) & (g716) & (!g549) & (!g569) & (g680)) + ((!g708) & (sk[87]) & (g716) & (!g549) & (g569) & (!g680)) + ((!g708) & (sk[87]) & (g716) & (!g549) & (g569) & (g680)) + ((!g708) & (sk[87]) & (g716) & (g549) & (g569) & (g680)) + ((g708) & (!sk[87]) & (!g716) & (!g549) & (g569) & (!g680)) + ((g708) & (!sk[87]) & (!g716) & (!g549) & (g569) & (g680)) + ((g708) & (!sk[87]) & (!g716) & (g549) & (!g569) & (!g680)) + ((g708) & (!sk[87]) & (!g716) & (g549) & (!g569) & (g680)) + ((g708) & (!sk[87]) & (!g716) & (g549) & (g569) & (!g680)) + ((g708) & (!sk[87]) & (!g716) & (g549) & (g569) & (g680)) + ((g708) & (!sk[87]) & (g716) & (!g549) & (!g569) & (!g680)) + ((g708) & (!sk[87]) & (g716) & (!g549) & (!g569) & (g680)) + ((g708) & (!sk[87]) & (g716) & (!g549) & (g569) & (!g680)) + ((g708) & (!sk[87]) & (g716) & (!g549) & (g569) & (g680)) + ((g708) & (!sk[87]) & (g716) & (g549) & (!g569) & (!g680)) + ((g708) & (!sk[87]) & (g716) & (g549) & (!g569) & (g680)) + ((g708) & (!sk[87]) & (g716) & (g549) & (g569) & (!g680)) + ((g708) & (!sk[87]) & (g716) & (g549) & (g569) & (g680)) + ((g708) & (sk[87]) & (!g716) & (!g549) & (!g569) & (g680)) + ((g708) & (sk[87]) & (!g716) & (!g549) & (g569) & (!g680)) + ((g708) & (sk[87]) & (!g716) & (!g549) & (g569) & (g680)) + ((g708) & (sk[87]) & (!g716) & (g549) & (g569) & (g680)) + ((g708) & (sk[87]) & (g716) & (!g549) & (!g569) & (!g680)) + ((g708) & (sk[87]) & (g716) & (!g549) & (!g569) & (g680)) + ((g708) & (sk[87]) & (g716) & (!g549) & (g569) & (!g680)) + ((g708) & (sk[87]) & (g716) & (!g549) & (g569) & (g680)) + ((g708) & (sk[87]) & (g716) & (g549) & (!g569) & (!g680)) + ((g708) & (sk[87]) & (g716) & (g549) & (!g569) & (g680)) + ((g708) & (sk[87]) & (g716) & (g549) & (g569) & (!g680)) + ((g708) & (sk[87]) & (g716) & (g549) & (g569) & (g680)));
	assign g718 = (((!g708) & (!g716) & (!g549) & (!g569) & (sk[88]) & (!g680)) + ((!g708) & (!g716) & (!g549) & (g569) & (!sk[88]) & (!g680)) + ((!g708) & (!g716) & (!g549) & (g569) & (!sk[88]) & (g680)) + ((!g708) & (!g716) & (g549) & (!g569) & (!sk[88]) & (!g680)) + ((!g708) & (!g716) & (g549) & (!g569) & (!sk[88]) & (g680)) + ((!g708) & (!g716) & (g549) & (!g569) & (sk[88]) & (!g680)) + ((!g708) & (!g716) & (g549) & (!g569) & (sk[88]) & (g680)) + ((!g708) & (!g716) & (g549) & (g569) & (!sk[88]) & (!g680)) + ((!g708) & (!g716) & (g549) & (g569) & (!sk[88]) & (g680)) + ((!g708) & (!g716) & (g549) & (g569) & (sk[88]) & (!g680)) + ((!g708) & (g716) & (!g549) & (!g569) & (!sk[88]) & (!g680)) + ((!g708) & (g716) & (!g549) & (!g569) & (!sk[88]) & (g680)) + ((!g708) & (g716) & (!g549) & (!g569) & (sk[88]) & (g680)) + ((!g708) & (g716) & (!g549) & (g569) & (!sk[88]) & (!g680)) + ((!g708) & (g716) & (!g549) & (g569) & (!sk[88]) & (g680)) + ((!g708) & (g716) & (!g549) & (g569) & (sk[88]) & (!g680)) + ((!g708) & (g716) & (!g549) & (g569) & (sk[88]) & (g680)) + ((!g708) & (g716) & (g549) & (!g569) & (!sk[88]) & (!g680)) + ((!g708) & (g716) & (g549) & (!g569) & (!sk[88]) & (g680)) + ((!g708) & (g716) & (g549) & (g569) & (!sk[88]) & (!g680)) + ((!g708) & (g716) & (g549) & (g569) & (!sk[88]) & (g680)) + ((!g708) & (g716) & (g549) & (g569) & (sk[88]) & (g680)) + ((g708) & (!g716) & (!g549) & (!g569) & (sk[88]) & (g680)) + ((g708) & (!g716) & (!g549) & (g569) & (!sk[88]) & (!g680)) + ((g708) & (!g716) & (!g549) & (g569) & (!sk[88]) & (g680)) + ((g708) & (!g716) & (!g549) & (g569) & (sk[88]) & (!g680)) + ((g708) & (!g716) & (!g549) & (g569) & (sk[88]) & (g680)) + ((g708) & (!g716) & (g549) & (!g569) & (!sk[88]) & (!g680)) + ((g708) & (!g716) & (g549) & (!g569) & (!sk[88]) & (g680)) + ((g708) & (!g716) & (g549) & (g569) & (!sk[88]) & (!g680)) + ((g708) & (!g716) & (g549) & (g569) & (!sk[88]) & (g680)) + ((g708) & (!g716) & (g549) & (g569) & (sk[88]) & (g680)) + ((g708) & (g716) & (!g549) & (!g569) & (!sk[88]) & (!g680)) + ((g708) & (g716) & (!g549) & (!g569) & (!sk[88]) & (g680)) + ((g708) & (g716) & (!g549) & (!g569) & (sk[88]) & (!g680)) + ((g708) & (g716) & (!g549) & (g569) & (!sk[88]) & (!g680)) + ((g708) & (g716) & (!g549) & (g569) & (!sk[88]) & (g680)) + ((g708) & (g716) & (g549) & (!g569) & (!sk[88]) & (!g680)) + ((g708) & (g716) & (g549) & (!g569) & (!sk[88]) & (g680)) + ((g708) & (g716) & (g549) & (!g569) & (sk[88]) & (!g680)) + ((g708) & (g716) & (g549) & (!g569) & (sk[88]) & (g680)) + ((g708) & (g716) & (g549) & (g569) & (!sk[88]) & (!g680)) + ((g708) & (g716) & (g549) & (g569) & (!sk[88]) & (g680)) + ((g708) & (g716) & (g549) & (g569) & (sk[88]) & (!g680)));
	assign g719 = (((!g585) & (!g597) & (sk[89]) & (!g679)) + ((!g585) & (g597) & (!sk[89]) & (!g679)) + ((!g585) & (g597) & (!sk[89]) & (g679)) + ((!g585) & (g597) & (sk[89]) & (g679)) + ((g585) & (!g597) & (sk[89]) & (g679)) + ((g585) & (g597) & (!sk[89]) & (!g679)) + ((g585) & (g597) & (!sk[89]) & (g679)) + ((g585) & (g597) & (sk[89]) & (!g679)));
	assign g720 = (((!g598) & (!g611) & (!sk[90]) & (!g612) & (g626) & (!g678)) + ((!g598) & (!g611) & (!sk[90]) & (!g612) & (g626) & (g678)) + ((!g598) & (!g611) & (!sk[90]) & (g612) & (!g626) & (!g678)) + ((!g598) & (!g611) & (!sk[90]) & (g612) & (!g626) & (g678)) + ((!g598) & (!g611) & (!sk[90]) & (g612) & (g626) & (!g678)) + ((!g598) & (!g611) & (!sk[90]) & (g612) & (g626) & (g678)) + ((!g598) & (!g611) & (sk[90]) & (!g612) & (!g626) & (g678)) + ((!g598) & (!g611) & (sk[90]) & (!g612) & (g626) & (!g678)) + ((!g598) & (!g611) & (sk[90]) & (!g612) & (g626) & (g678)) + ((!g598) & (!g611) & (sk[90]) & (g612) & (g626) & (g678)) + ((!g598) & (g611) & (!sk[90]) & (!g612) & (!g626) & (!g678)) + ((!g598) & (g611) & (!sk[90]) & (!g612) & (!g626) & (g678)) + ((!g598) & (g611) & (!sk[90]) & (!g612) & (g626) & (!g678)) + ((!g598) & (g611) & (!sk[90]) & (!g612) & (g626) & (g678)) + ((!g598) & (g611) & (!sk[90]) & (g612) & (!g626) & (!g678)) + ((!g598) & (g611) & (!sk[90]) & (g612) & (!g626) & (g678)) + ((!g598) & (g611) & (!sk[90]) & (g612) & (g626) & (!g678)) + ((!g598) & (g611) & (!sk[90]) & (g612) & (g626) & (g678)) + ((!g598) & (g611) & (sk[90]) & (!g612) & (!g626) & (!g678)) + ((!g598) & (g611) & (sk[90]) & (g612) & (!g626) & (!g678)) + ((!g598) & (g611) & (sk[90]) & (g612) & (!g626) & (g678)) + ((!g598) & (g611) & (sk[90]) & (g612) & (g626) & (!g678)) + ((g598) & (!g611) & (!sk[90]) & (!g612) & (g626) & (!g678)) + ((g598) & (!g611) & (!sk[90]) & (!g612) & (g626) & (g678)) + ((g598) & (!g611) & (!sk[90]) & (g612) & (!g626) & (!g678)) + ((g598) & (!g611) & (!sk[90]) & (g612) & (!g626) & (g678)) + ((g598) & (!g611) & (!sk[90]) & (g612) & (g626) & (!g678)) + ((g598) & (!g611) & (!sk[90]) & (g612) & (g626) & (g678)) + ((g598) & (!g611) & (sk[90]) & (!g612) & (!g626) & (!g678)) + ((g598) & (!g611) & (sk[90]) & (g612) & (!g626) & (!g678)) + ((g598) & (!g611) & (sk[90]) & (g612) & (!g626) & (g678)) + ((g598) & (!g611) & (sk[90]) & (g612) & (g626) & (!g678)) + ((g598) & (g611) & (!sk[90]) & (!g612) & (!g626) & (!g678)) + ((g598) & (g611) & (!sk[90]) & (!g612) & (!g626) & (g678)) + ((g598) & (g611) & (!sk[90]) & (!g612) & (g626) & (!g678)) + ((g598) & (g611) & (!sk[90]) & (!g612) & (g626) & (g678)) + ((g598) & (g611) & (!sk[90]) & (g612) & (!g626) & (!g678)) + ((g598) & (g611) & (!sk[90]) & (g612) & (!g626) & (g678)) + ((g598) & (g611) & (!sk[90]) & (g612) & (g626) & (!g678)) + ((g598) & (g611) & (!sk[90]) & (g612) & (g626) & (g678)) + ((g598) & (g611) & (sk[90]) & (!g612) & (!g626) & (g678)) + ((g598) & (g611) & (sk[90]) & (!g612) & (g626) & (!g678)) + ((g598) & (g611) & (sk[90]) & (!g612) & (g626) & (g678)) + ((g598) & (g611) & (sk[90]) & (g612) & (g626) & (g678)));
	assign g721 = (((!g440) & (!g441) & (!g454) & (!g455) & (!g546) & (g626)) + ((!g440) & (!g441) & (!g454) & (!g455) & (g546) & (g626)) + ((!g440) & (!g441) & (!g454) & (g455) & (!g546) & (!g626)) + ((!g440) & (!g441) & (!g454) & (g455) & (g546) & (g626)) + ((!g440) & (!g441) & (g454) & (!g455) & (!g546) & (!g626)) + ((!g440) & (!g441) & (g454) & (!g455) & (g546) & (g626)) + ((!g440) & (!g441) & (g454) & (g455) & (!g546) & (!g626)) + ((!g440) & (!g441) & (g454) & (g455) & (g546) & (!g626)) + ((!g440) & (g441) & (!g454) & (!g455) & (!g546) & (!g626)) + ((!g440) & (g441) & (!g454) & (!g455) & (g546) & (!g626)) + ((!g440) & (g441) & (!g454) & (g455) & (!g546) & (g626)) + ((!g440) & (g441) & (!g454) & (g455) & (g546) & (!g626)) + ((!g440) & (g441) & (g454) & (!g455) & (!g546) & (g626)) + ((!g440) & (g441) & (g454) & (!g455) & (g546) & (!g626)) + ((!g440) & (g441) & (g454) & (g455) & (!g546) & (g626)) + ((!g440) & (g441) & (g454) & (g455) & (g546) & (g626)) + ((g440) & (!g441) & (!g454) & (!g455) & (!g546) & (!g626)) + ((g440) & (!g441) & (!g454) & (!g455) & (g546) & (!g626)) + ((g440) & (!g441) & (!g454) & (g455) & (!g546) & (g626)) + ((g440) & (!g441) & (!g454) & (g455) & (g546) & (!g626)) + ((g440) & (!g441) & (g454) & (!g455) & (!g546) & (g626)) + ((g440) & (!g441) & (g454) & (!g455) & (g546) & (!g626)) + ((g440) & (!g441) & (g454) & (g455) & (!g546) & (g626)) + ((g440) & (!g441) & (g454) & (g455) & (g546) & (g626)) + ((g440) & (g441) & (!g454) & (!g455) & (!g546) & (g626)) + ((g440) & (g441) & (!g454) & (!g455) & (g546) & (g626)) + ((g440) & (g441) & (!g454) & (g455) & (!g546) & (!g626)) + ((g440) & (g441) & (!g454) & (g455) & (g546) & (g626)) + ((g440) & (g441) & (g454) & (!g455) & (!g546) & (!g626)) + ((g440) & (g441) & (g454) & (!g455) & (g546) & (g626)) + ((g440) & (g441) & (g454) & (g455) & (!g546) & (!g626)) + ((g440) & (g441) & (g454) & (g455) & (g546) & (!g626)));
	assign g722 = (((!sk[92]) & (g721) & (g678)) + ((sk[92]) & (!g721) & (g678)) + ((sk[92]) & (g721) & (!g678)));
	assign g723 = (((!g627) & (!g546) & (!g640) & (!g641) & (!g655) & (!g677)) + ((!g627) & (!g546) & (!g640) & (g641) & (!g655) & (!g677)) + ((!g627) & (!g546) & (!g640) & (g641) & (!g655) & (g677)) + ((!g627) & (!g546) & (!g640) & (g641) & (g655) & (!g677)) + ((!g627) & (!g546) & (g640) & (!g641) & (!g655) & (g677)) + ((!g627) & (!g546) & (g640) & (!g641) & (g655) & (!g677)) + ((!g627) & (!g546) & (g640) & (!g641) & (g655) & (g677)) + ((!g627) & (!g546) & (g640) & (g641) & (g655) & (g677)) + ((!g627) & (g546) & (!g640) & (!g641) & (!g655) & (g677)) + ((!g627) & (g546) & (!g640) & (!g641) & (g655) & (!g677)) + ((!g627) & (g546) & (!g640) & (!g641) & (g655) & (g677)) + ((!g627) & (g546) & (!g640) & (g641) & (g655) & (g677)) + ((!g627) & (g546) & (g640) & (!g641) & (!g655) & (!g677)) + ((!g627) & (g546) & (g640) & (g641) & (!g655) & (!g677)) + ((!g627) & (g546) & (g640) & (g641) & (!g655) & (g677)) + ((!g627) & (g546) & (g640) & (g641) & (g655) & (!g677)) + ((g627) & (!g546) & (!g640) & (!g641) & (!g655) & (g677)) + ((g627) & (!g546) & (!g640) & (!g641) & (g655) & (!g677)) + ((g627) & (!g546) & (!g640) & (!g641) & (g655) & (g677)) + ((g627) & (!g546) & (!g640) & (g641) & (g655) & (g677)) + ((g627) & (!g546) & (g640) & (!g641) & (!g655) & (!g677)) + ((g627) & (!g546) & (g640) & (g641) & (!g655) & (!g677)) + ((g627) & (!g546) & (g640) & (g641) & (!g655) & (g677)) + ((g627) & (!g546) & (g640) & (g641) & (g655) & (!g677)) + ((g627) & (g546) & (!g640) & (!g641) & (!g655) & (!g677)) + ((g627) & (g546) & (!g640) & (g641) & (!g655) & (!g677)) + ((g627) & (g546) & (!g640) & (g641) & (!g655) & (g677)) + ((g627) & (g546) & (!g640) & (g641) & (g655) & (!g677)) + ((g627) & (g546) & (g640) & (!g641) & (!g655) & (g677)) + ((g627) & (g546) & (g640) & (!g641) & (g655) & (!g677)) + ((g627) & (g546) & (g640) & (!g641) & (g655) & (g677)) + ((g627) & (g546) & (g640) & (g641) & (g655) & (g677)));
	assign g724 = (((!sk[94]) & (!g641) & (g655) & (!g677)) + ((!sk[94]) & (!g641) & (g655) & (g677)) + ((!sk[94]) & (g641) & (g655) & (!g677)) + ((!sk[94]) & (g641) & (g655) & (g677)) + ((sk[94]) & (!g641) & (!g655) & (!g677)) + ((sk[94]) & (!g641) & (g655) & (g677)) + ((sk[94]) & (g641) & (!g655) & (g677)) + ((sk[94]) & (g641) & (g655) & (!g677)));
	assign g725 = (((!sk[95]) & (!g490) & (g658) & (!g676)) + ((!sk[95]) & (!g490) & (g658) & (g676)) + ((!sk[95]) & (g490) & (g658) & (!g676)) + ((!sk[95]) & (g490) & (g658) & (g676)) + ((sk[95]) & (!g490) & (!g658) & (!g676)) + ((sk[95]) & (!g490) & (g658) & (g676)) + ((sk[95]) & (g490) & (!g658) & (g676)) + ((sk[95]) & (g490) & (g658) & (!g676)));
	assign g726 = (((!g656) & (!g657) & (!g488) & (!g658) & (!g670) & (!g676)) + ((!g656) & (!g657) & (!g488) & (!g658) & (g670) & (g676)) + ((!g656) & (!g657) & (!g488) & (g658) & (!g670) & (!g676)) + ((!g656) & (!g657) & (!g488) & (g658) & (!g670) & (g676)) + ((!g656) & (!g657) & (g488) & (!g658) & (g670) & (!g676)) + ((!g656) & (!g657) & (g488) & (!g658) & (g670) & (g676)) + ((!g656) & (!g657) & (g488) & (g658) & (!g670) & (!g676)) + ((!g656) & (!g657) & (g488) & (g658) & (g670) & (g676)) + ((!g656) & (g657) & (!g488) & (!g658) & (g670) & (!g676)) + ((!g656) & (g657) & (!g488) & (!g658) & (g670) & (g676)) + ((!g656) & (g657) & (!g488) & (g658) & (!g670) & (!g676)) + ((!g656) & (g657) & (!g488) & (g658) & (g670) & (g676)) + ((!g656) & (g657) & (g488) & (!g658) & (!g670) & (g676)) + ((!g656) & (g657) & (g488) & (!g658) & (g670) & (!g676)) + ((!g656) & (g657) & (g488) & (g658) & (g670) & (!g676)) + ((!g656) & (g657) & (g488) & (g658) & (g670) & (g676)) + ((g656) & (!g657) & (!g488) & (!g658) & (!g670) & (g676)) + ((g656) & (!g657) & (!g488) & (!g658) & (g670) & (!g676)) + ((g656) & (!g657) & (!g488) & (g658) & (g670) & (!g676)) + ((g656) & (!g657) & (!g488) & (g658) & (g670) & (g676)) + ((g656) & (!g657) & (g488) & (!g658) & (!g670) & (!g676)) + ((g656) & (!g657) & (g488) & (!g658) & (!g670) & (g676)) + ((g656) & (!g657) & (g488) & (g658) & (!g670) & (g676)) + ((g656) & (!g657) & (g488) & (g658) & (g670) & (!g676)) + ((g656) & (g657) & (!g488) & (!g658) & (!g670) & (!g676)) + ((g656) & (g657) & (!g488) & (!g658) & (!g670) & (g676)) + ((g656) & (g657) & (!g488) & (g658) & (!g670) & (g676)) + ((g656) & (g657) & (!g488) & (g658) & (g670) & (!g676)) + ((g656) & (g657) & (g488) & (!g658) & (!g670) & (!g676)) + ((g656) & (g657) & (g488) & (!g658) & (g670) & (g676)) + ((g656) & (g657) & (g488) & (g658) & (!g670) & (!g676)) + ((g656) & (g657) & (g488) & (g658) & (!g670) & (g676)));
	assign g727 = (((!g721) & (!g678) & (!g723) & (!g724) & (!g725) & (!g726)) + ((!g721) & (!g678) & (!g723) & (!g724) & (!g725) & (g726)) + ((!g721) & (!g678) & (!g723) & (!g724) & (g725) & (!g726)) + ((!g721) & (!g678) & (!g723) & (!g724) & (g725) & (g726)) + ((!g721) & (!g678) & (!g723) & (g724) & (!g725) & (!g726)) + ((!g721) & (!g678) & (!g723) & (g724) & (!g725) & (g726)) + ((!g721) & (!g678) & (!g723) & (g724) & (g725) & (!g726)) + ((!g721) & (!g678) & (!g723) & (g724) & (g725) & (g726)) + ((!g721) & (!g678) & (g723) & (!g724) & (!g725) & (g726)) + ((!g721) & (!g678) & (g723) & (!g724) & (g725) & (g726)) + ((!g721) & (g678) & (!g723) & (!g724) & (!g725) & (!g726)) + ((!g721) & (g678) & (!g723) & (!g724) & (!g725) & (g726)) + ((!g721) & (g678) & (!g723) & (!g724) & (g725) & (!g726)) + ((!g721) & (g678) & (!g723) & (!g724) & (g725) & (g726)) + ((!g721) & (g678) & (!g723) & (g724) & (!g725) & (g726)) + ((g721) & (!g678) & (!g723) & (!g724) & (!g725) & (!g726)) + ((g721) & (!g678) & (!g723) & (!g724) & (!g725) & (g726)) + ((g721) & (!g678) & (!g723) & (!g724) & (g725) & (!g726)) + ((g721) & (!g678) & (!g723) & (!g724) & (g725) & (g726)) + ((g721) & (!g678) & (!g723) & (g724) & (!g725) & (g726)) + ((g721) & (g678) & (!g723) & (!g724) & (!g725) & (!g726)) + ((g721) & (g678) & (!g723) & (!g724) & (!g725) & (g726)) + ((g721) & (g678) & (!g723) & (!g724) & (g725) & (!g726)) + ((g721) & (g678) & (!g723) & (!g724) & (g725) & (g726)) + ((g721) & (g678) & (!g723) & (g724) & (!g725) & (!g726)) + ((g721) & (g678) & (!g723) & (g724) & (!g725) & (g726)) + ((g721) & (g678) & (!g723) & (g724) & (g725) & (!g726)) + ((g721) & (g678) & (!g723) & (g724) & (g725) & (g726)) + ((g721) & (g678) & (g723) & (!g724) & (!g725) & (g726)) + ((g721) & (g678) & (g723) & (!g724) & (g725) & (g726)));
	assign g728 = (((!g585) & (!g597) & (!g679) & (g720) & (!g722) & (!g727)) + ((!g585) & (!g597) & (!g679) & (g720) & (!g722) & (g727)) + ((!g585) & (!g597) & (!g679) & (g720) & (g722) & (g727)) + ((!g585) & (!g597) & (g679) & (!g720) & (!g722) & (g727)) + ((!g585) & (!g597) & (g679) & (g720) & (!g722) & (!g727)) + ((!g585) & (!g597) & (g679) & (g720) & (!g722) & (g727)) + ((!g585) & (!g597) & (g679) & (g720) & (g722) & (!g727)) + ((!g585) & (!g597) & (g679) & (g720) & (g722) & (g727)) + ((!g585) & (g597) & (!g679) & (!g720) & (!g722) & (g727)) + ((!g585) & (g597) & (!g679) & (g720) & (!g722) & (!g727)) + ((!g585) & (g597) & (!g679) & (g720) & (!g722) & (g727)) + ((!g585) & (g597) & (!g679) & (g720) & (g722) & (!g727)) + ((!g585) & (g597) & (!g679) & (g720) & (g722) & (g727)) + ((!g585) & (g597) & (g679) & (g720) & (!g722) & (!g727)) + ((!g585) & (g597) & (g679) & (g720) & (!g722) & (g727)) + ((!g585) & (g597) & (g679) & (g720) & (g722) & (g727)) + ((g585) & (!g597) & (!g679) & (!g720) & (!g722) & (g727)) + ((g585) & (!g597) & (!g679) & (g720) & (!g722) & (!g727)) + ((g585) & (!g597) & (!g679) & (g720) & (!g722) & (g727)) + ((g585) & (!g597) & (!g679) & (g720) & (g722) & (!g727)) + ((g585) & (!g597) & (!g679) & (g720) & (g722) & (g727)) + ((g585) & (!g597) & (g679) & (g720) & (!g722) & (!g727)) + ((g585) & (!g597) & (g679) & (g720) & (!g722) & (g727)) + ((g585) & (!g597) & (g679) & (g720) & (g722) & (g727)) + ((g585) & (g597) & (!g679) & (g720) & (!g722) & (!g727)) + ((g585) & (g597) & (!g679) & (g720) & (!g722) & (g727)) + ((g585) & (g597) & (!g679) & (g720) & (g722) & (g727)) + ((g585) & (g597) & (g679) & (!g720) & (!g722) & (g727)) + ((g585) & (g597) & (g679) & (g720) & (!g722) & (!g727)) + ((g585) & (g597) & (g679) & (g720) & (!g722) & (g727)) + ((g585) & (g597) & (g679) & (g720) & (g722) & (!g727)) + ((g585) & (g597) & (g679) & (g720) & (g722) & (g727)));
	assign g729 = (((!g570) & (!g571) & (!g584) & (!g585) & (!g597) & (g679)) + ((!g570) & (!g571) & (!g584) & (!g585) & (g597) & (!g679)) + ((!g570) & (!g571) & (!g584) & (!g585) & (g597) & (g679)) + ((!g570) & (!g571) & (!g584) & (g585) & (g597) & (g679)) + ((!g570) & (!g571) & (g584) & (!g585) & (!g597) & (!g679)) + ((!g570) & (!g571) & (g584) & (g585) & (!g597) & (!g679)) + ((!g570) & (!g571) & (g584) & (g585) & (!g597) & (g679)) + ((!g570) & (!g571) & (g584) & (g585) & (g597) & (!g679)) + ((!g570) & (g571) & (!g584) & (!g585) & (!g597) & (!g679)) + ((!g570) & (g571) & (!g584) & (g585) & (!g597) & (!g679)) + ((!g570) & (g571) & (!g584) & (g585) & (!g597) & (g679)) + ((!g570) & (g571) & (!g584) & (g585) & (g597) & (!g679)) + ((!g570) & (g571) & (g584) & (!g585) & (!g597) & (g679)) + ((!g570) & (g571) & (g584) & (!g585) & (g597) & (!g679)) + ((!g570) & (g571) & (g584) & (!g585) & (g597) & (g679)) + ((!g570) & (g571) & (g584) & (g585) & (g597) & (g679)) + ((g570) & (!g571) & (!g584) & (!g585) & (!g597) & (!g679)) + ((g570) & (!g571) & (!g584) & (g585) & (!g597) & (!g679)) + ((g570) & (!g571) & (!g584) & (g585) & (!g597) & (g679)) + ((g570) & (!g571) & (!g584) & (g585) & (g597) & (!g679)) + ((g570) & (!g571) & (g584) & (!g585) & (!g597) & (g679)) + ((g570) & (!g571) & (g584) & (!g585) & (g597) & (!g679)) + ((g570) & (!g571) & (g584) & (!g585) & (g597) & (g679)) + ((g570) & (!g571) & (g584) & (g585) & (g597) & (g679)) + ((g570) & (g571) & (!g584) & (!g585) & (!g597) & (g679)) + ((g570) & (g571) & (!g584) & (!g585) & (g597) & (!g679)) + ((g570) & (g571) & (!g584) & (!g585) & (g597) & (g679)) + ((g570) & (g571) & (!g584) & (g585) & (g597) & (g679)) + ((g570) & (g571) & (g584) & (!g585) & (!g597) & (!g679)) + ((g570) & (g571) & (g584) & (g585) & (!g597) & (!g679)) + ((g570) & (g571) & (g584) & (g585) & (!g597) & (g679)) + ((g570) & (g571) & (g584) & (g585) & (g597) & (!g679)));
	assign g730 = (((!g549) & (!g569) & (!g680) & (!g719) & (!g728) & (!g729)) + ((!g549) & (!g569) & (!g680) & (!g719) & (g728) & (!g729)) + ((!g549) & (!g569) & (!g680) & (g719) & (g728) & (!g729)) + ((!g549) & (!g569) & (g680) & (!g719) & (!g728) & (!g729)) + ((!g549) & (!g569) & (g680) & (!g719) & (g728) & (!g729)) + ((!g549) & (!g569) & (g680) & (!g719) & (g728) & (g729)) + ((!g549) & (!g569) & (g680) & (g719) & (!g728) & (!g729)) + ((!g549) & (!g569) & (g680) & (g719) & (g728) & (!g729)) + ((!g549) & (g569) & (!g680) & (!g719) & (!g728) & (!g729)) + ((!g549) & (g569) & (!g680) & (!g719) & (g728) & (!g729)) + ((!g549) & (g569) & (!g680) & (!g719) & (g728) & (g729)) + ((!g549) & (g569) & (!g680) & (g719) & (!g728) & (!g729)) + ((!g549) & (g569) & (!g680) & (g719) & (g728) & (!g729)) + ((!g549) & (g569) & (g680) & (!g719) & (!g728) & (!g729)) + ((!g549) & (g569) & (g680) & (!g719) & (g728) & (!g729)) + ((!g549) & (g569) & (g680) & (g719) & (g728) & (!g729)) + ((g549) & (!g569) & (!g680) & (!g719) & (!g728) & (!g729)) + ((g549) & (!g569) & (!g680) & (!g719) & (g728) & (!g729)) + ((g549) & (!g569) & (!g680) & (!g719) & (g728) & (g729)) + ((g549) & (!g569) & (!g680) & (g719) & (!g728) & (!g729)) + ((g549) & (!g569) & (!g680) & (g719) & (g728) & (!g729)) + ((g549) & (!g569) & (g680) & (!g719) & (!g728) & (!g729)) + ((g549) & (!g569) & (g680) & (!g719) & (g728) & (!g729)) + ((g549) & (!g569) & (g680) & (g719) & (g728) & (!g729)) + ((g549) & (g569) & (!g680) & (!g719) & (!g728) & (!g729)) + ((g549) & (g569) & (!g680) & (!g719) & (g728) & (!g729)) + ((g549) & (g569) & (!g680) & (g719) & (g728) & (!g729)) + ((g549) & (g569) & (g680) & (!g719) & (!g728) & (!g729)) + ((g549) & (g569) & (g680) & (!g719) & (g728) & (!g729)) + ((g549) & (g569) & (g680) & (!g719) & (g728) & (g729)) + ((g549) & (g569) & (g680) & (g719) & (!g728) & (!g729)) + ((g549) & (g569) & (g680) & (g719) & (g728) & (!g729)));
	assign g731 = (((!g707) & (!g717) & (!sk[101]) & (!g681) & (g718) & (!g730)) + ((!g707) & (!g717) & (!sk[101]) & (!g681) & (g718) & (g730)) + ((!g707) & (!g717) & (!sk[101]) & (g681) & (!g718) & (!g730)) + ((!g707) & (!g717) & (!sk[101]) & (g681) & (!g718) & (g730)) + ((!g707) & (!g717) & (!sk[101]) & (g681) & (g718) & (!g730)) + ((!g707) & (!g717) & (!sk[101]) & (g681) & (g718) & (g730)) + ((!g707) & (!g717) & (sk[101]) & (!g681) & (!g718) & (g730)) + ((!g707) & (!g717) & (sk[101]) & (g681) & (g718) & (!g730)) + ((!g707) & (g717) & (!sk[101]) & (!g681) & (!g718) & (!g730)) + ((!g707) & (g717) & (!sk[101]) & (!g681) & (!g718) & (g730)) + ((!g707) & (g717) & (!sk[101]) & (!g681) & (g718) & (!g730)) + ((!g707) & (g717) & (!sk[101]) & (!g681) & (g718) & (g730)) + ((!g707) & (g717) & (!sk[101]) & (g681) & (!g718) & (!g730)) + ((!g707) & (g717) & (!sk[101]) & (g681) & (!g718) & (g730)) + ((!g707) & (g717) & (!sk[101]) & (g681) & (g718) & (!g730)) + ((!g707) & (g717) & (!sk[101]) & (g681) & (g718) & (g730)) + ((!g707) & (g717) & (sk[101]) & (!g681) & (!g718) & (!g730)) + ((!g707) & (g717) & (sk[101]) & (!g681) & (g718) & (!g730)) + ((!g707) & (g717) & (sk[101]) & (!g681) & (g718) & (g730)) + ((!g707) & (g717) & (sk[101]) & (g681) & (!g718) & (!g730)) + ((!g707) & (g717) & (sk[101]) & (g681) & (!g718) & (g730)) + ((!g707) & (g717) & (sk[101]) & (g681) & (g718) & (g730)) + ((g707) & (!g717) & (!sk[101]) & (!g681) & (g718) & (!g730)) + ((g707) & (!g717) & (!sk[101]) & (!g681) & (g718) & (g730)) + ((g707) & (!g717) & (!sk[101]) & (g681) & (!g718) & (!g730)) + ((g707) & (!g717) & (!sk[101]) & (g681) & (!g718) & (g730)) + ((g707) & (!g717) & (!sk[101]) & (g681) & (g718) & (!g730)) + ((g707) & (!g717) & (!sk[101]) & (g681) & (g718) & (g730)) + ((g707) & (!g717) & (sk[101]) & (!g681) & (!g718) & (!g730)) + ((g707) & (!g717) & (sk[101]) & (!g681) & (g718) & (!g730)) + ((g707) & (!g717) & (sk[101]) & (!g681) & (g718) & (g730)) + ((g707) & (!g717) & (sk[101]) & (g681) & (!g718) & (!g730)) + ((g707) & (!g717) & (sk[101]) & (g681) & (!g718) & (g730)) + ((g707) & (!g717) & (sk[101]) & (g681) & (g718) & (g730)) + ((g707) & (g717) & (!sk[101]) & (!g681) & (!g718) & (!g730)) + ((g707) & (g717) & (!sk[101]) & (!g681) & (!g718) & (g730)) + ((g707) & (g717) & (!sk[101]) & (!g681) & (g718) & (!g730)) + ((g707) & (g717) & (!sk[101]) & (!g681) & (g718) & (g730)) + ((g707) & (g717) & (!sk[101]) & (g681) & (!g718) & (!g730)) + ((g707) & (g717) & (!sk[101]) & (g681) & (!g718) & (g730)) + ((g707) & (g717) & (!sk[101]) & (g681) & (g718) & (!g730)) + ((g707) & (g717) & (!sk[101]) & (g681) & (g718) & (g730)) + ((g707) & (g717) & (sk[101]) & (!g681) & (!g718) & (g730)) + ((g707) & (g717) & (sk[101]) & (g681) & (g718) & (!g730)));
	assign g732 = (((!sk[102]) & (g682) & (g684)) + ((sk[102]) & (g682) & (g684)));
	assign g733 = (((!sk[103]) & (g682) & (g684)) + ((sk[103]) & (!g682) & (g684)));
	assign g734 = (((!sk[104]) & (g684) & (g685)) + ((sk[104]) & (!g684) & (g685)));
	assign g735 = (((!g707) & (!g717) & (!g733) & (!sk[105]) & (g734) & (!g718)) + ((!g707) & (!g717) & (!g733) & (!sk[105]) & (g734) & (g718)) + ((!g707) & (!g717) & (!g733) & (sk[105]) & (g734) & (g718)) + ((!g707) & (!g717) & (g733) & (!sk[105]) & (!g734) & (!g718)) + ((!g707) & (!g717) & (g733) & (!sk[105]) & (!g734) & (g718)) + ((!g707) & (!g717) & (g733) & (!sk[105]) & (g734) & (!g718)) + ((!g707) & (!g717) & (g733) & (!sk[105]) & (g734) & (g718)) + ((!g707) & (!g717) & (g733) & (sk[105]) & (g734) & (g718)) + ((!g707) & (g717) & (!g733) & (!sk[105]) & (!g734) & (!g718)) + ((!g707) & (g717) & (!g733) & (!sk[105]) & (!g734) & (g718)) + ((!g707) & (g717) & (!g733) & (!sk[105]) & (g734) & (!g718)) + ((!g707) & (g717) & (!g733) & (!sk[105]) & (g734) & (g718)) + ((!g707) & (g717) & (!g733) & (sk[105]) & (g734) & (g718)) + ((!g707) & (g717) & (g733) & (!sk[105]) & (!g734) & (!g718)) + ((!g707) & (g717) & (g733) & (!sk[105]) & (!g734) & (g718)) + ((!g707) & (g717) & (g733) & (!sk[105]) & (g734) & (!g718)) + ((!g707) & (g717) & (g733) & (!sk[105]) & (g734) & (g718)) + ((!g707) & (g717) & (g733) & (sk[105]) & (!g734) & (!g718)) + ((!g707) & (g717) & (g733) & (sk[105]) & (!g734) & (g718)) + ((!g707) & (g717) & (g733) & (sk[105]) & (g734) & (!g718)) + ((!g707) & (g717) & (g733) & (sk[105]) & (g734) & (g718)) + ((g707) & (!g717) & (!g733) & (!sk[105]) & (g734) & (!g718)) + ((g707) & (!g717) & (!g733) & (!sk[105]) & (g734) & (g718)) + ((g707) & (!g717) & (!g733) & (sk[105]) & (g734) & (g718)) + ((g707) & (!g717) & (g733) & (!sk[105]) & (!g734) & (!g718)) + ((g707) & (!g717) & (g733) & (!sk[105]) & (!g734) & (g718)) + ((g707) & (!g717) & (g733) & (!sk[105]) & (g734) & (!g718)) + ((g707) & (!g717) & (g733) & (!sk[105]) & (g734) & (g718)) + ((g707) & (!g717) & (g733) & (sk[105]) & (!g734) & (!g718)) + ((g707) & (!g717) & (g733) & (sk[105]) & (!g734) & (g718)) + ((g707) & (!g717) & (g733) & (sk[105]) & (g734) & (!g718)) + ((g707) & (!g717) & (g733) & (sk[105]) & (g734) & (g718)) + ((g707) & (g717) & (!g733) & (!sk[105]) & (!g734) & (!g718)) + ((g707) & (g717) & (!g733) & (!sk[105]) & (!g734) & (g718)) + ((g707) & (g717) & (!g733) & (!sk[105]) & (g734) & (!g718)) + ((g707) & (g717) & (!g733) & (!sk[105]) & (g734) & (g718)) + ((g707) & (g717) & (!g733) & (sk[105]) & (g734) & (g718)) + ((g707) & (g717) & (g733) & (!sk[105]) & (!g734) & (!g718)) + ((g707) & (g717) & (g733) & (!sk[105]) & (!g734) & (g718)) + ((g707) & (g717) & (g733) & (!sk[105]) & (g734) & (!g718)) + ((g707) & (g717) & (g733) & (!sk[105]) & (g734) & (g718)) + ((g707) & (g717) & (g733) & (sk[105]) & (g734) & (g718)));
	assign g736 = (((!g2) & (!g681) & (!g686) & (!g731) & (!g732) & (!g735)) + ((!g2) & (!g681) & (!g686) & (!g731) & (g732) & (!g735)) + ((!g2) & (!g681) & (!g686) & (g731) & (!g732) & (!g735)) + ((!g2) & (g681) & (!g686) & (!g731) & (!g732) & (!g735)) + ((!g2) & (g681) & (!g686) & (!g731) & (g732) & (!g735)) + ((!g2) & (g681) & (!g686) & (g731) & (!g732) & (!g735)) + ((!g2) & (g681) & (g686) & (!g731) & (!g732) & (!g735)) + ((!g2) & (g681) & (g686) & (!g731) & (g732) & (!g735)) + ((!g2) & (g681) & (g686) & (g731) & (!g732) & (!g735)) + ((g2) & (!g681) & (!g686) & (!g731) & (!g732) & (g735)) + ((g2) & (!g681) & (!g686) & (!g731) & (g732) & (g735)) + ((g2) & (!g681) & (!g686) & (g731) & (!g732) & (g735)) + ((g2) & (!g681) & (!g686) & (g731) & (g732) & (!g735)) + ((g2) & (!g681) & (!g686) & (g731) & (g732) & (g735)) + ((g2) & (!g681) & (g686) & (!g731) & (!g732) & (!g735)) + ((g2) & (!g681) & (g686) & (!g731) & (!g732) & (g735)) + ((g2) & (!g681) & (g686) & (!g731) & (g732) & (!g735)) + ((g2) & (!g681) & (g686) & (!g731) & (g732) & (g735)) + ((g2) & (!g681) & (g686) & (g731) & (!g732) & (!g735)) + ((g2) & (!g681) & (g686) & (g731) & (!g732) & (g735)) + ((g2) & (!g681) & (g686) & (g731) & (g732) & (!g735)) + ((g2) & (!g681) & (g686) & (g731) & (g732) & (g735)) + ((g2) & (g681) & (!g686) & (!g731) & (!g732) & (g735)) + ((g2) & (g681) & (!g686) & (!g731) & (g732) & (g735)) + ((g2) & (g681) & (!g686) & (g731) & (!g732) & (g735)) + ((g2) & (g681) & (!g686) & (g731) & (g732) & (!g735)) + ((g2) & (g681) & (!g686) & (g731) & (g732) & (g735)) + ((g2) & (g681) & (g686) & (!g731) & (!g732) & (g735)) + ((g2) & (g681) & (g686) & (!g731) & (g732) & (g735)) + ((g2) & (g681) & (g686) & (g731) & (!g732) & (g735)) + ((g2) & (g681) & (g686) & (g731) & (g732) & (!g735)) + ((g2) & (g681) & (g686) & (g731) & (g732) & (g735)));
	assign g737 = (((!sk[107]) & (g305) & (g200)) + ((sk[107]) & (!g305) & (g200)) + ((sk[107]) & (g305) & (!g200)));
	assign g738 = (((!sk[108]) & (!g490) & (!g658) & (!g676) & (g737)) + ((!sk[108]) & (!g490) & (!g658) & (g676) & (g737)) + ((!sk[108]) & (!g490) & (g658) & (!g676) & (g737)) + ((!sk[108]) & (!g490) & (g658) & (g676) & (g737)) + ((!sk[108]) & (g490) & (!g658) & (!g676) & (!g737)) + ((!sk[108]) & (g490) & (!g658) & (!g676) & (g737)) + ((!sk[108]) & (g490) & (!g658) & (g676) & (!g737)) + ((!sk[108]) & (g490) & (!g658) & (g676) & (g737)) + ((!sk[108]) & (g490) & (g658) & (!g676) & (!g737)) + ((!sk[108]) & (g490) & (g658) & (!g676) & (g737)) + ((!sk[108]) & (g490) & (g658) & (g676) & (!g737)) + ((!sk[108]) & (g490) & (g658) & (g676) & (g737)) + ((sk[108]) & (!g490) & (!g658) & (g676) & (g737)) + ((sk[108]) & (!g490) & (g658) & (!g676) & (g737)) + ((sk[108]) & (g490) & (!g658) & (!g676) & (g737)) + ((sk[108]) & (g490) & (g658) & (g676) & (g737)));
	assign g739 = (((!g2) & (!g198) & (g200) & (!g367) & (!g725) & (!g726)) + ((!g2) & (!g198) & (g200) & (!g367) & (!g725) & (g726)) + ((!g2) & (!g198) & (g200) & (!g367) & (g725) & (!g726)) + ((!g2) & (!g198) & (g200) & (!g367) & (g725) & (g726)) + ((!g2) & (!g198) & (g200) & (g367) & (g725) & (!g726)) + ((!g2) & (g198) & (g200) & (!g367) & (g725) & (!g726)) + ((!g2) & (g198) & (g200) & (!g367) & (g725) & (g726)) + ((!g2) & (g198) & (g200) & (g367) & (g725) & (!g726)) + ((g2) & (!g198) & (g200) & (!g367) & (g725) & (!g726)) + ((g2) & (!g198) & (g200) & (g367) & (g725) & (!g726)) + ((g2) & (!g198) & (g200) & (g367) & (g725) & (g726)) + ((g2) & (g198) & (g200) & (!g367) & (g725) & (!g726)) + ((g2) & (g198) & (g200) & (g367) & (!g725) & (!g726)) + ((g2) & (g198) & (g200) & (g367) & (!g725) & (g726)) + ((g2) & (g198) & (g200) & (g367) & (g725) & (!g726)) + ((g2) & (g198) & (g200) & (g367) & (g725) & (g726)));
	assign g740 = (((!sk[110]) & (g198) & (g200)) + ((sk[110]) & (!g198) & (g200)) + ((sk[110]) & (g198) & (!g200)));
	assign g741 = (((!sk[111]) & (g2) & (g367)) + ((sk[111]) & (!g2) & (g367)) + ((sk[111]) & (g2) & (!g367)));
	assign g742 = (((g740) & (!sk[112]) & (g741)) + ((g740) & (sk[112]) & (g741)));
	assign g743 = (((!sk[113]) & (g198) & (g367)) + ((sk[113]) & (!g198) & (g367)) + ((sk[113]) & (g198) & (!g367)));
	assign g744 = (((!sk[114]) & (g741) & (g743)) + ((sk[114]) & (!g741) & (g743)));
	assign g745 = (((!sk[115]) & (g726) & (g744)) + ((sk[115]) & (g726) & (g744)));
	assign g746 = (((!g641) & (!g655) & (!sk[116]) & (!g677) & (g725) & (!g726)) + ((!g641) & (!g655) & (!sk[116]) & (!g677) & (g725) & (g726)) + ((!g641) & (!g655) & (!sk[116]) & (g677) & (!g725) & (!g726)) + ((!g641) & (!g655) & (!sk[116]) & (g677) & (!g725) & (g726)) + ((!g641) & (!g655) & (!sk[116]) & (g677) & (g725) & (!g726)) + ((!g641) & (!g655) & (!sk[116]) & (g677) & (g725) & (g726)) + ((!g641) & (!g655) & (sk[116]) & (!g677) & (!g725) & (!g726)) + ((!g641) & (!g655) & (sk[116]) & (!g677) & (!g725) & (g726)) + ((!g641) & (!g655) & (sk[116]) & (!g677) & (g725) & (!g726)) + ((!g641) & (!g655) & (sk[116]) & (g677) & (g725) & (g726)) + ((!g641) & (g655) & (!sk[116]) & (!g677) & (!g725) & (!g726)) + ((!g641) & (g655) & (!sk[116]) & (!g677) & (!g725) & (g726)) + ((!g641) & (g655) & (!sk[116]) & (!g677) & (g725) & (!g726)) + ((!g641) & (g655) & (!sk[116]) & (!g677) & (g725) & (g726)) + ((!g641) & (g655) & (!sk[116]) & (g677) & (!g725) & (!g726)) + ((!g641) & (g655) & (!sk[116]) & (g677) & (!g725) & (g726)) + ((!g641) & (g655) & (!sk[116]) & (g677) & (g725) & (!g726)) + ((!g641) & (g655) & (!sk[116]) & (g677) & (g725) & (g726)) + ((!g641) & (g655) & (sk[116]) & (!g677) & (g725) & (g726)) + ((!g641) & (g655) & (sk[116]) & (g677) & (!g725) & (!g726)) + ((!g641) & (g655) & (sk[116]) & (g677) & (!g725) & (g726)) + ((!g641) & (g655) & (sk[116]) & (g677) & (g725) & (!g726)) + ((g641) & (!g655) & (!sk[116]) & (!g677) & (g725) & (!g726)) + ((g641) & (!g655) & (!sk[116]) & (!g677) & (g725) & (g726)) + ((g641) & (!g655) & (!sk[116]) & (g677) & (!g725) & (!g726)) + ((g641) & (!g655) & (!sk[116]) & (g677) & (!g725) & (g726)) + ((g641) & (!g655) & (!sk[116]) & (g677) & (g725) & (!g726)) + ((g641) & (!g655) & (!sk[116]) & (g677) & (g725) & (g726)) + ((g641) & (!g655) & (sk[116]) & (!g677) & (g725) & (g726)) + ((g641) & (!g655) & (sk[116]) & (g677) & (!g725) & (!g726)) + ((g641) & (!g655) & (sk[116]) & (g677) & (!g725) & (g726)) + ((g641) & (!g655) & (sk[116]) & (g677) & (g725) & (!g726)) + ((g641) & (g655) & (!sk[116]) & (!g677) & (!g725) & (!g726)) + ((g641) & (g655) & (!sk[116]) & (!g677) & (!g725) & (g726)) + ((g641) & (g655) & (!sk[116]) & (!g677) & (g725) & (!g726)) + ((g641) & (g655) & (!sk[116]) & (!g677) & (g725) & (g726)) + ((g641) & (g655) & (!sk[116]) & (g677) & (!g725) & (!g726)) + ((g641) & (g655) & (!sk[116]) & (g677) & (!g725) & (g726)) + ((g641) & (g655) & (!sk[116]) & (g677) & (g725) & (!g726)) + ((g641) & (g655) & (!sk[116]) & (g677) & (g725) & (g726)) + ((g641) & (g655) & (sk[116]) & (!g677) & (!g725) & (!g726)) + ((g641) & (g655) & (sk[116]) & (!g677) & (!g725) & (g726)) + ((g641) & (g655) & (sk[116]) & (!g677) & (g725) & (!g726)) + ((g641) & (g655) & (sk[116]) & (g677) & (g725) & (g726)));
	assign g747 = (((!sk[117]) & (g740) & (g741)) + ((sk[117]) & (!g740) & (g741)));
	assign g748 = (((!sk[118]) & (!g740) & (g741) & (!g743)) + ((!sk[118]) & (!g740) & (g741) & (g743)) + ((!sk[118]) & (g740) & (g741) & (!g743)) + ((!sk[118]) & (g740) & (g741) & (g743)) + ((sk[118]) & (g740) & (!g741) & (!g743)));
	assign g749 = (((!g641) & (!g655) & (!g677) & (!g725) & (!g747) & (g748)) + ((!g641) & (!g655) & (!g677) & (!g725) & (g747) & (g748)) + ((!g641) & (!g655) & (g677) & (!g725) & (!g747) & (g748)) + ((!g641) & (!g655) & (g677) & (!g725) & (g747) & (!g748)) + ((!g641) & (!g655) & (g677) & (!g725) & (g747) & (g748)) + ((!g641) & (!g655) & (g677) & (g725) & (g747) & (!g748)) + ((!g641) & (!g655) & (g677) & (g725) & (g747) & (g748)) + ((!g641) & (g655) & (!g677) & (!g725) & (!g747) & (g748)) + ((!g641) & (g655) & (!g677) & (!g725) & (g747) & (!g748)) + ((!g641) & (g655) & (!g677) & (!g725) & (g747) & (g748)) + ((!g641) & (g655) & (!g677) & (g725) & (g747) & (!g748)) + ((!g641) & (g655) & (!g677) & (g725) & (g747) & (g748)) + ((!g641) & (g655) & (g677) & (!g725) & (!g747) & (g748)) + ((!g641) & (g655) & (g677) & (!g725) & (g747) & (g748)) + ((g641) & (!g655) & (!g677) & (!g725) & (!g747) & (g748)) + ((g641) & (!g655) & (!g677) & (!g725) & (g747) & (!g748)) + ((g641) & (!g655) & (!g677) & (!g725) & (g747) & (g748)) + ((g641) & (!g655) & (!g677) & (g725) & (g747) & (!g748)) + ((g641) & (!g655) & (!g677) & (g725) & (g747) & (g748)) + ((g641) & (!g655) & (g677) & (!g725) & (!g747) & (g748)) + ((g641) & (!g655) & (g677) & (!g725) & (g747) & (g748)) + ((g641) & (g655) & (!g677) & (!g725) & (!g747) & (g748)) + ((g641) & (g655) & (!g677) & (!g725) & (g747) & (g748)) + ((g641) & (g655) & (g677) & (!g725) & (!g747) & (g748)) + ((g641) & (g655) & (g677) & (!g725) & (g747) & (!g748)) + ((g641) & (g655) & (g677) & (!g725) & (g747) & (g748)) + ((g641) & (g655) & (g677) & (g725) & (g747) & (!g748)) + ((g641) & (g655) & (g677) & (g725) & (g747) & (g748)));
	assign g750 = (((!g742) & (!g745) & (!g746) & (!sk[120]) & (g749)) + ((!g742) & (!g745) & (!g746) & (sk[120]) & (!g749)) + ((!g742) & (!g745) & (g746) & (!sk[120]) & (g749)) + ((!g742) & (!g745) & (g746) & (sk[120]) & (!g749)) + ((!g742) & (g745) & (!g746) & (!sk[120]) & (g749)) + ((!g742) & (g745) & (g746) & (!sk[120]) & (g749)) + ((g742) & (!g745) & (!g746) & (!sk[120]) & (!g749)) + ((g742) & (!g745) & (!g746) & (!sk[120]) & (g749)) + ((g742) & (!g745) & (g746) & (!sk[120]) & (!g749)) + ((g742) & (!g745) & (g746) & (!sk[120]) & (g749)) + ((g742) & (!g745) & (g746) & (sk[120]) & (!g749)) + ((g742) & (g745) & (!g746) & (!sk[120]) & (!g749)) + ((g742) & (g745) & (!g746) & (!sk[120]) & (g749)) + ((g742) & (g745) & (g746) & (!sk[120]) & (!g749)) + ((g742) & (g745) & (g746) & (!sk[120]) & (g749)));
	assign g751 = (((!g723) & (!g724) & (!g725) & (!sk[121]) & (g726) & (!g742)) + ((!g723) & (!g724) & (!g725) & (!sk[121]) & (g726) & (g742)) + ((!g723) & (!g724) & (!g725) & (sk[121]) & (g726) & (g742)) + ((!g723) & (!g724) & (g725) & (!sk[121]) & (!g726) & (!g742)) + ((!g723) & (!g724) & (g725) & (!sk[121]) & (!g726) & (g742)) + ((!g723) & (!g724) & (g725) & (!sk[121]) & (g726) & (!g742)) + ((!g723) & (!g724) & (g725) & (!sk[121]) & (g726) & (g742)) + ((!g723) & (!g724) & (g725) & (sk[121]) & (g726) & (g742)) + ((!g723) & (g724) & (!g725) & (!sk[121]) & (!g726) & (!g742)) + ((!g723) & (g724) & (!g725) & (!sk[121]) & (!g726) & (g742)) + ((!g723) & (g724) & (!g725) & (!sk[121]) & (g726) & (!g742)) + ((!g723) & (g724) & (!g725) & (!sk[121]) & (g726) & (g742)) + ((!g723) & (g724) & (!g725) & (sk[121]) & (!g726) & (g742)) + ((!g723) & (g724) & (g725) & (!sk[121]) & (!g726) & (!g742)) + ((!g723) & (g724) & (g725) & (!sk[121]) & (!g726) & (g742)) + ((!g723) & (g724) & (g725) & (!sk[121]) & (g726) & (!g742)) + ((!g723) & (g724) & (g725) & (!sk[121]) & (g726) & (g742)) + ((!g723) & (g724) & (g725) & (sk[121]) & (!g726) & (g742)) + ((!g723) & (g724) & (g725) & (sk[121]) & (g726) & (g742)) + ((g723) & (!g724) & (!g725) & (!sk[121]) & (g726) & (!g742)) + ((g723) & (!g724) & (!g725) & (!sk[121]) & (g726) & (g742)) + ((g723) & (!g724) & (!g725) & (sk[121]) & (!g726) & (g742)) + ((g723) & (!g724) & (g725) & (!sk[121]) & (!g726) & (!g742)) + ((g723) & (!g724) & (g725) & (!sk[121]) & (!g726) & (g742)) + ((g723) & (!g724) & (g725) & (!sk[121]) & (g726) & (!g742)) + ((g723) & (!g724) & (g725) & (!sk[121]) & (g726) & (g742)) + ((g723) & (!g724) & (g725) & (sk[121]) & (!g726) & (g742)) + ((g723) & (g724) & (!g725) & (!sk[121]) & (!g726) & (!g742)) + ((g723) & (g724) & (!g725) & (!sk[121]) & (!g726) & (g742)) + ((g723) & (g724) & (!g725) & (!sk[121]) & (g726) & (!g742)) + ((g723) & (g724) & (!g725) & (!sk[121]) & (g726) & (g742)) + ((g723) & (g724) & (!g725) & (sk[121]) & (g726) & (g742)) + ((g723) & (g724) & (g725) & (!sk[121]) & (!g726) & (!g742)) + ((g723) & (g724) & (g725) & (!sk[121]) & (!g726) & (g742)) + ((g723) & (g724) & (g725) & (!sk[121]) & (g726) & (!g742)) + ((g723) & (g724) & (g725) & (!sk[121]) & (g726) & (g742)));
	assign g752 = (((!g723) & (!g724) & (!g726) & (!g747) & (!g744) & (!g748)) + ((!g723) & (!g724) & (!g726) & (!g747) & (!g744) & (g748)) + ((!g723) & (!g724) & (g726) & (!g747) & (!g744) & (!g748)) + ((!g723) & (g724) & (!g726) & (!g747) & (!g744) & (!g748)) + ((!g723) & (g724) & (!g726) & (!g747) & (!g744) & (g748)) + ((!g723) & (g724) & (!g726) & (!g747) & (g744) & (!g748)) + ((!g723) & (g724) & (!g726) & (!g747) & (g744) & (g748)) + ((!g723) & (g724) & (g726) & (!g747) & (!g744) & (!g748)) + ((!g723) & (g724) & (g726) & (!g747) & (g744) & (!g748)) + ((g723) & (!g724) & (!g726) & (!g747) & (!g744) & (!g748)) + ((g723) & (!g724) & (!g726) & (!g747) & (!g744) & (g748)) + ((g723) & (!g724) & (!g726) & (g747) & (!g744) & (!g748)) + ((g723) & (!g724) & (!g726) & (g747) & (!g744) & (g748)) + ((g723) & (!g724) & (g726) & (!g747) & (!g744) & (!g748)) + ((g723) & (!g724) & (g726) & (g747) & (!g744) & (!g748)) + ((g723) & (g724) & (!g726) & (!g747) & (!g744) & (!g748)) + ((g723) & (g724) & (!g726) & (!g747) & (!g744) & (g748)) + ((g723) & (g724) & (!g726) & (!g747) & (g744) & (!g748)) + ((g723) & (g724) & (!g726) & (!g747) & (g744) & (g748)) + ((g723) & (g724) & (!g726) & (g747) & (!g744) & (!g748)) + ((g723) & (g724) & (!g726) & (g747) & (!g744) & (g748)) + ((g723) & (g724) & (!g726) & (g747) & (g744) & (!g748)) + ((g723) & (g724) & (!g726) & (g747) & (g744) & (g748)) + ((g723) & (g724) & (g726) & (!g747) & (!g744) & (!g748)) + ((g723) & (g724) & (g726) & (!g747) & (g744) & (!g748)) + ((g723) & (g724) & (g726) & (g747) & (!g744) & (!g748)) + ((g723) & (g724) & (g726) & (g747) & (g744) & (!g748)));
	assign g753 = (((!g200) & (!g738) & (g739) & (!g750) & (!g751) & (!g752)) + ((!g200) & (!g738) & (g739) & (!g750) & (g751) & (!g752)) + ((!g200) & (!g738) & (g739) & (!g750) & (g751) & (g752)) + ((!g200) & (g738) & (!g739) & (!g750) & (!g751) & (!g752)) + ((!g200) & (g738) & (!g739) & (!g750) & (g751) & (!g752)) + ((!g200) & (g738) & (!g739) & (!g750) & (g751) & (g752)) + ((!g200) & (g738) & (!g739) & (g750) & (!g751) & (!g752)) + ((!g200) & (g738) & (!g739) & (g750) & (g751) & (!g752)) + ((!g200) & (g738) & (!g739) & (g750) & (g751) & (g752)) + ((!g200) & (g738) & (g739) & (!g750) & (!g751) & (!g752)) + ((!g200) & (g738) & (g739) & (!g750) & (!g751) & (g752)) + ((!g200) & (g738) & (g739) & (!g750) & (g751) & (!g752)) + ((!g200) & (g738) & (g739) & (!g750) & (g751) & (g752)) + ((!g200) & (g738) & (g739) & (g750) & (!g751) & (!g752)) + ((!g200) & (g738) & (g739) & (g750) & (g751) & (!g752)) + ((!g200) & (g738) & (g739) & (g750) & (g751) & (g752)) + ((g200) & (!g738) & (g739) & (g750) & (!g751) & (g752)) + ((g200) & (g738) & (!g739) & (!g750) & (!g751) & (g752)) + ((g200) & (g738) & (!g739) & (g750) & (!g751) & (g752)) + ((g200) & (g738) & (g739) & (!g750) & (!g751) & (g752)) + ((g200) & (g738) & (g739) & (g750) & (!g751) & (!g752)) + ((g200) & (g738) & (g739) & (g750) & (!g751) & (g752)) + ((g200) & (g738) & (g739) & (g750) & (g751) & (!g752)) + ((g200) & (g738) & (g739) & (g750) & (g751) & (g752)));
	assign g754 = (((!g721) & (!g678) & (!g723) & (!g724) & (!g725) & (!g726)) + ((!g721) & (!g678) & (!g723) & (!g724) & (!g725) & (g726)) + ((!g721) & (!g678) & (!g723) & (!g724) & (g725) & (!g726)) + ((!g721) & (!g678) & (!g723) & (!g724) & (g725) & (g726)) + ((!g721) & (!g678) & (!g723) & (g724) & (!g725) & (g726)) + ((!g721) & (!g678) & (g723) & (!g724) & (!g725) & (!g726)) + ((!g721) & (!g678) & (g723) & (!g724) & (g725) & (!g726)) + ((!g721) & (!g678) & (g723) & (g724) & (!g725) & (!g726)) + ((!g721) & (!g678) & (g723) & (g724) & (!g725) & (g726)) + ((!g721) & (!g678) & (g723) & (g724) & (g725) & (!g726)) + ((!g721) & (!g678) & (g723) & (g724) & (g725) & (g726)) + ((!g721) & (g678) & (!g723) & (g724) & (!g725) & (!g726)) + ((!g721) & (g678) & (!g723) & (g724) & (g725) & (!g726)) + ((!g721) & (g678) & (!g723) & (g724) & (g725) & (g726)) + ((!g721) & (g678) & (g723) & (!g724) & (!g725) & (g726)) + ((!g721) & (g678) & (g723) & (!g724) & (g725) & (g726)) + ((g721) & (!g678) & (!g723) & (g724) & (!g725) & (!g726)) + ((g721) & (!g678) & (!g723) & (g724) & (g725) & (!g726)) + ((g721) & (!g678) & (!g723) & (g724) & (g725) & (g726)) + ((g721) & (!g678) & (g723) & (!g724) & (!g725) & (g726)) + ((g721) & (!g678) & (g723) & (!g724) & (g725) & (g726)) + ((g721) & (g678) & (!g723) & (!g724) & (!g725) & (!g726)) + ((g721) & (g678) & (!g723) & (!g724) & (!g725) & (g726)) + ((g721) & (g678) & (!g723) & (!g724) & (g725) & (!g726)) + ((g721) & (g678) & (!g723) & (!g724) & (g725) & (g726)) + ((g721) & (g678) & (!g723) & (g724) & (!g725) & (g726)) + ((g721) & (g678) & (g723) & (!g724) & (!g725) & (!g726)) + ((g721) & (g678) & (g723) & (!g724) & (g725) & (!g726)) + ((g721) & (g678) & (g723) & (g724) & (!g725) & (!g726)) + ((g721) & (g678) & (g723) & (g724) & (!g725) & (g726)) + ((g721) & (g678) & (g723) & (g724) & (g725) & (!g726)) + ((g721) & (g678) & (g723) & (g724) & (g725) & (g726)));
	assign g755 = (((!sk[125]) & (!g723) & (!g724) & (!g744) & (g748)) + ((!sk[125]) & (!g723) & (!g724) & (g744) & (g748)) + ((!sk[125]) & (!g723) & (g724) & (!g744) & (g748)) + ((!sk[125]) & (!g723) & (g724) & (g744) & (g748)) + ((!sk[125]) & (g723) & (!g724) & (!g744) & (!g748)) + ((!sk[125]) & (g723) & (!g724) & (!g744) & (g748)) + ((!sk[125]) & (g723) & (!g724) & (g744) & (!g748)) + ((!sk[125]) & (g723) & (!g724) & (g744) & (g748)) + ((!sk[125]) & (g723) & (g724) & (!g744) & (!g748)) + ((!sk[125]) & (g723) & (g724) & (!g744) & (g748)) + ((!sk[125]) & (g723) & (g724) & (g744) & (!g748)) + ((!sk[125]) & (g723) & (g724) & (g744) & (g748)) + ((sk[125]) & (!g723) & (!g724) & (!g744) & (g748)) + ((sk[125]) & (!g723) & (!g724) & (g744) & (!g748)) + ((sk[125]) & (!g723) & (!g724) & (g744) & (g748)) + ((sk[125]) & (!g723) & (g724) & (g744) & (!g748)) + ((sk[125]) & (!g723) & (g724) & (g744) & (g748)) + ((sk[125]) & (g723) & (!g724) & (!g744) & (g748)) + ((sk[125]) & (g723) & (!g724) & (g744) & (g748)));
	assign g756 = (((!g198) & (!g200) & (!g722) & (!g741) & (!g754) & (!g755)) + ((!g198) & (!g200) & (!g722) & (!g741) & (g754) & (!g755)) + ((!g198) & (!g200) & (g722) & (!g741) & (!g754) & (!g755)) + ((!g198) & (!g200) & (g722) & (!g741) & (g754) & (!g755)) + ((!g198) & (!g200) & (g722) & (g741) & (!g754) & (!g755)) + ((!g198) & (!g200) & (g722) & (g741) & (g754) & (!g755)) + ((!g198) & (g200) & (!g722) & (!g741) & (!g754) & (g755)) + ((!g198) & (g200) & (!g722) & (!g741) & (g754) & (g755)) + ((!g198) & (g200) & (!g722) & (g741) & (!g754) & (g755)) + ((!g198) & (g200) & (!g722) & (g741) & (g754) & (!g755)) + ((!g198) & (g200) & (!g722) & (g741) & (g754) & (g755)) + ((!g198) & (g200) & (g722) & (!g741) & (!g754) & (g755)) + ((!g198) & (g200) & (g722) & (!g741) & (g754) & (g755)) + ((!g198) & (g200) & (g722) & (g741) & (!g754) & (g755)) + ((!g198) & (g200) & (g722) & (g741) & (g754) & (!g755)) + ((!g198) & (g200) & (g722) & (g741) & (g754) & (g755)) + ((g198) & (!g200) & (!g722) & (!g741) & (!g754) & (!g755)) + ((g198) & (!g200) & (!g722) & (!g741) & (g754) & (!g755)) + ((g198) & (!g200) & (!g722) & (g741) & (!g754) & (!g755)) + ((g198) & (!g200) & (g722) & (!g741) & (!g754) & (!g755)) + ((g198) & (!g200) & (g722) & (!g741) & (g754) & (!g755)) + ((g198) & (!g200) & (g722) & (g741) & (!g754) & (!g755)) + ((g198) & (g200) & (!g722) & (!g741) & (!g754) & (g755)) + ((g198) & (g200) & (!g722) & (!g741) & (g754) & (g755)) + ((g198) & (g200) & (!g722) & (g741) & (!g754) & (!g755)) + ((g198) & (g200) & (!g722) & (g741) & (!g754) & (g755)) + ((g198) & (g200) & (!g722) & (g741) & (g754) & (!g755)) + ((g198) & (g200) & (!g722) & (g741) & (g754) & (g755)) + ((g198) & (g200) & (g722) & (!g741) & (!g754) & (g755)) + ((g198) & (g200) & (g722) & (!g741) & (g754) & (g755)) + ((g198) & (g200) & (g722) & (g741) & (!g754) & (g755)) + ((g198) & (g200) & (g722) & (g741) & (g754) & (g755)));
	assign g757 = (((!g305) & (!g222) & (!g200) & (!sk[127]) & (g725) & (!g726)) + ((!g305) & (!g222) & (!g200) & (!sk[127]) & (g725) & (g726)) + ((!g305) & (!g222) & (g200) & (!sk[127]) & (!g725) & (!g726)) + ((!g305) & (!g222) & (g200) & (!sk[127]) & (!g725) & (g726)) + ((!g305) & (!g222) & (g200) & (!sk[127]) & (g725) & (!g726)) + ((!g305) & (!g222) & (g200) & (!sk[127]) & (g725) & (g726)) + ((!g305) & (!g222) & (g200) & (sk[127]) & (!g725) & (g726)) + ((!g305) & (!g222) & (g200) & (sk[127]) & (g725) & (g726)) + ((!g305) & (g222) & (!g200) & (!sk[127]) & (!g725) & (!g726)) + ((!g305) & (g222) & (!g200) & (!sk[127]) & (!g725) & (g726)) + ((!g305) & (g222) & (!g200) & (!sk[127]) & (g725) & (!g726)) + ((!g305) & (g222) & (!g200) & (!sk[127]) & (g725) & (g726)) + ((!g305) & (g222) & (!g200) & (sk[127]) & (!g725) & (!g726)) + ((!g305) & (g222) & (!g200) & (sk[127]) & (!g725) & (g726)) + ((!g305) & (g222) & (g200) & (!sk[127]) & (!g725) & (!g726)) + ((!g305) & (g222) & (g200) & (!sk[127]) & (!g725) & (g726)) + ((!g305) & (g222) & (g200) & (!sk[127]) & (g725) & (!g726)) + ((!g305) & (g222) & (g200) & (!sk[127]) & (g725) & (g726)) + ((!g305) & (g222) & (g200) & (sk[127]) & (!g725) & (!g726)) + ((!g305) & (g222) & (g200) & (sk[127]) & (g725) & (g726)) + ((g305) & (!g222) & (!g200) & (!sk[127]) & (g725) & (!g726)) + ((g305) & (!g222) & (!g200) & (!sk[127]) & (g725) & (g726)) + ((g305) & (!g222) & (!g200) & (sk[127]) & (!g725) & (g726)) + ((g305) & (!g222) & (!g200) & (sk[127]) & (g725) & (g726)) + ((g305) & (!g222) & (g200) & (!sk[127]) & (!g725) & (!g726)) + ((g305) & (!g222) & (g200) & (!sk[127]) & (!g725) & (g726)) + ((g305) & (!g222) & (g200) & (!sk[127]) & (g725) & (!g726)) + ((g305) & (!g222) & (g200) & (!sk[127]) & (g725) & (g726)) + ((g305) & (!g222) & (g200) & (sk[127]) & (!g725) & (!g726)) + ((g305) & (!g222) & (g200) & (sk[127]) & (!g725) & (g726)) + ((g305) & (g222) & (!g200) & (!sk[127]) & (!g725) & (!g726)) + ((g305) & (g222) & (!g200) & (!sk[127]) & (!g725) & (g726)) + ((g305) & (g222) & (!g200) & (!sk[127]) & (g725) & (!g726)) + ((g305) & (g222) & (!g200) & (!sk[127]) & (g725) & (g726)) + ((g305) & (g222) & (!g200) & (sk[127]) & (!g725) & (!g726)) + ((g305) & (g222) & (!g200) & (sk[127]) & (g725) & (g726)) + ((g305) & (g222) & (g200) & (!sk[127]) & (!g725) & (!g726)) + ((g305) & (g222) & (g200) & (!sk[127]) & (!g725) & (g726)) + ((g305) & (g222) & (g200) & (!sk[127]) & (g725) & (!g726)) + ((g305) & (g222) & (g200) & (!sk[127]) & (g725) & (g726)));
	assign g758 = (((!sk[0]) & (g202) & (g222)) + ((sk[0]) & (!g202) & (g222)) + ((sk[0]) & (g202) & (!g222)));
	assign g759 = (((g737) & (!sk[1]) & (g758)) + ((g737) & (sk[1]) & (g758)));
	assign g760 = (((g202) & (!g305) & (!g222) & (!g200) & (!g725) & (!g726)) + ((g202) & (!g305) & (!g222) & (!g200) & (!g725) & (g726)) + ((g202) & (!g305) & (!g222) & (!g200) & (g725) & (!g726)) + ((g202) & (!g305) & (!g222) & (!g200) & (g725) & (g726)) + ((g202) & (!g305) & (!g222) & (g200) & (g725) & (!g726)) + ((g202) & (!g305) & (g222) & (!g200) & (g725) & (!g726)) + ((g202) & (!g305) & (g222) & (!g200) & (g725) & (g726)) + ((g202) & (!g305) & (g222) & (g200) & (g725) & (!g726)) + ((g202) & (g305) & (!g222) & (!g200) & (g725) & (!g726)) + ((g202) & (g305) & (!g222) & (g200) & (g725) & (!g726)) + ((g202) & (g305) & (!g222) & (g200) & (g725) & (g726)) + ((g202) & (g305) & (g222) & (!g200) & (g725) & (!g726)) + ((g202) & (g305) & (g222) & (g200) & (!g725) & (!g726)) + ((g202) & (g305) & (g222) & (g200) & (!g725) & (g726)) + ((g202) & (g305) & (g222) & (g200) & (g725) & (!g726)) + ((g202) & (g305) & (g222) & (g200) & (g725) & (g726)));
	assign g761 = (((!g305) & (sk[3]) & (g222)) + ((g305) & (!sk[3]) & (g222)) + ((g305) & (sk[3]) & (!g222)));
	assign g762 = (((!sk[4]) & (g737) & (g761)) + ((sk[4]) & (!g737) & (g761)));
	assign g763 = (((g726) & (!sk[5]) & (g762)) + ((g726) & (sk[5]) & (g762)));
	assign g764 = (((!sk[6]) & (g737) & (g758)) + ((sk[6]) & (g737) & (!g758)));
	assign g765 = (((!g737) & (!sk[7]) & (g758) & (!g761)) + ((!g737) & (!sk[7]) & (g758) & (g761)) + ((!g737) & (sk[7]) & (g758) & (!g761)) + ((g737) & (!sk[7]) & (g758) & (!g761)) + ((g737) & (!sk[7]) & (g758) & (g761)));
	assign g766 = (((!g641) & (!g655) & (!g677) & (!g725) & (!g764) & (g765)) + ((!g641) & (!g655) & (!g677) & (!g725) & (g764) & (g765)) + ((!g641) & (!g655) & (g677) & (!g725) & (!g764) & (g765)) + ((!g641) & (!g655) & (g677) & (!g725) & (g764) & (!g765)) + ((!g641) & (!g655) & (g677) & (!g725) & (g764) & (g765)) + ((!g641) & (!g655) & (g677) & (g725) & (g764) & (!g765)) + ((!g641) & (!g655) & (g677) & (g725) & (g764) & (g765)) + ((!g641) & (g655) & (!g677) & (!g725) & (!g764) & (g765)) + ((!g641) & (g655) & (!g677) & (!g725) & (g764) & (!g765)) + ((!g641) & (g655) & (!g677) & (!g725) & (g764) & (g765)) + ((!g641) & (g655) & (!g677) & (g725) & (g764) & (!g765)) + ((!g641) & (g655) & (!g677) & (g725) & (g764) & (g765)) + ((!g641) & (g655) & (g677) & (!g725) & (!g764) & (g765)) + ((!g641) & (g655) & (g677) & (!g725) & (g764) & (g765)) + ((g641) & (!g655) & (!g677) & (!g725) & (!g764) & (g765)) + ((g641) & (!g655) & (!g677) & (!g725) & (g764) & (!g765)) + ((g641) & (!g655) & (!g677) & (!g725) & (g764) & (g765)) + ((g641) & (!g655) & (!g677) & (g725) & (g764) & (!g765)) + ((g641) & (!g655) & (!g677) & (g725) & (g764) & (g765)) + ((g641) & (!g655) & (g677) & (!g725) & (!g764) & (g765)) + ((g641) & (!g655) & (g677) & (!g725) & (g764) & (g765)) + ((g641) & (g655) & (!g677) & (!g725) & (!g764) & (g765)) + ((g641) & (g655) & (!g677) & (!g725) & (g764) & (g765)) + ((g641) & (g655) & (g677) & (!g725) & (!g764) & (g765)) + ((g641) & (g655) & (g677) & (!g725) & (g764) & (!g765)) + ((g641) & (g655) & (g677) & (!g725) & (g764) & (g765)) + ((g641) & (g655) & (g677) & (g725) & (g764) & (!g765)) + ((g641) & (g655) & (g677) & (g725) & (g764) & (g765)));
	assign g767 = (((!g202) & (!g746) & (!g759) & (!g760) & (!g763) & (g766)) + ((!g202) & (!g746) & (!g759) & (!g760) & (g763) & (!g766)) + ((!g202) & (!g746) & (!g759) & (!g760) & (g763) & (g766)) + ((!g202) & (!g746) & (!g759) & (g760) & (!g763) & (!g766)) + ((!g202) & (!g746) & (g759) & (!g760) & (!g763) & (!g766)) + ((!g202) & (!g746) & (g759) & (!g760) & (!g763) & (g766)) + ((!g202) & (!g746) & (g759) & (!g760) & (g763) & (!g766)) + ((!g202) & (!g746) & (g759) & (!g760) & (g763) & (g766)) + ((!g202) & (g746) & (!g759) & (!g760) & (!g763) & (g766)) + ((!g202) & (g746) & (!g759) & (!g760) & (g763) & (!g766)) + ((!g202) & (g746) & (!g759) & (!g760) & (g763) & (g766)) + ((!g202) & (g746) & (!g759) & (g760) & (!g763) & (!g766)) + ((!g202) & (g746) & (g759) & (!g760) & (!g763) & (g766)) + ((!g202) & (g746) & (g759) & (!g760) & (g763) & (!g766)) + ((!g202) & (g746) & (g759) & (!g760) & (g763) & (g766)) + ((!g202) & (g746) & (g759) & (g760) & (!g763) & (!g766)) + ((g202) & (!g746) & (!g759) & (!g760) & (!g763) & (!g766)) + ((g202) & (!g746) & (!g759) & (g760) & (!g763) & (g766)) + ((g202) & (!g746) & (!g759) & (g760) & (g763) & (!g766)) + ((g202) & (!g746) & (!g759) & (g760) & (g763) & (g766)) + ((g202) & (!g746) & (g759) & (g760) & (!g763) & (!g766)) + ((g202) & (!g746) & (g759) & (g760) & (!g763) & (g766)) + ((g202) & (!g746) & (g759) & (g760) & (g763) & (!g766)) + ((g202) & (!g746) & (g759) & (g760) & (g763) & (g766)) + ((g202) & (g746) & (!g759) & (!g760) & (!g763) & (!g766)) + ((g202) & (g746) & (!g759) & (g760) & (!g763) & (g766)) + ((g202) & (g746) & (!g759) & (g760) & (g763) & (!g766)) + ((g202) & (g746) & (!g759) & (g760) & (g763) & (g766)) + ((g202) & (g746) & (g759) & (!g760) & (!g763) & (!g766)) + ((g202) & (g746) & (g759) & (g760) & (!g763) & (g766)) + ((g202) & (g746) & (g759) & (g760) & (g763) & (!g766)) + ((g202) & (g746) & (g759) & (g760) & (g763) & (g766)));
	assign g768 = (((!g721) & (!g678) & (!g723) & (!sk[10]) & (g744) & (!g748)) + ((!g721) & (!g678) & (!g723) & (!sk[10]) & (g744) & (g748)) + ((!g721) & (!g678) & (!g723) & (sk[10]) & (!g744) & (g748)) + ((!g721) & (!g678) & (!g723) & (sk[10]) & (g744) & (!g748)) + ((!g721) & (!g678) & (!g723) & (sk[10]) & (g744) & (g748)) + ((!g721) & (!g678) & (g723) & (!sk[10]) & (!g744) & (!g748)) + ((!g721) & (!g678) & (g723) & (!sk[10]) & (!g744) & (g748)) + ((!g721) & (!g678) & (g723) & (!sk[10]) & (g744) & (!g748)) + ((!g721) & (!g678) & (g723) & (!sk[10]) & (g744) & (g748)) + ((!g721) & (!g678) & (g723) & (sk[10]) & (g744) & (!g748)) + ((!g721) & (!g678) & (g723) & (sk[10]) & (g744) & (g748)) + ((!g721) & (g678) & (!g723) & (!sk[10]) & (!g744) & (!g748)) + ((!g721) & (g678) & (!g723) & (!sk[10]) & (!g744) & (g748)) + ((!g721) & (g678) & (!g723) & (!sk[10]) & (g744) & (!g748)) + ((!g721) & (g678) & (!g723) & (!sk[10]) & (g744) & (g748)) + ((!g721) & (g678) & (!g723) & (sk[10]) & (!g744) & (g748)) + ((!g721) & (g678) & (!g723) & (sk[10]) & (g744) & (g748)) + ((!g721) & (g678) & (g723) & (!sk[10]) & (!g744) & (!g748)) + ((!g721) & (g678) & (g723) & (!sk[10]) & (!g744) & (g748)) + ((!g721) & (g678) & (g723) & (!sk[10]) & (g744) & (!g748)) + ((!g721) & (g678) & (g723) & (!sk[10]) & (g744) & (g748)) + ((g721) & (!g678) & (!g723) & (!sk[10]) & (g744) & (!g748)) + ((g721) & (!g678) & (!g723) & (!sk[10]) & (g744) & (g748)) + ((g721) & (!g678) & (!g723) & (sk[10]) & (!g744) & (g748)) + ((g721) & (!g678) & (!g723) & (sk[10]) & (g744) & (g748)) + ((g721) & (!g678) & (g723) & (!sk[10]) & (!g744) & (!g748)) + ((g721) & (!g678) & (g723) & (!sk[10]) & (!g744) & (g748)) + ((g721) & (!g678) & (g723) & (!sk[10]) & (g744) & (!g748)) + ((g721) & (!g678) & (g723) & (!sk[10]) & (g744) & (g748)) + ((g721) & (g678) & (!g723) & (!sk[10]) & (!g744) & (!g748)) + ((g721) & (g678) & (!g723) & (!sk[10]) & (!g744) & (g748)) + ((g721) & (g678) & (!g723) & (!sk[10]) & (g744) & (!g748)) + ((g721) & (g678) & (!g723) & (!sk[10]) & (g744) & (g748)) + ((g721) & (g678) & (!g723) & (sk[10]) & (!g744) & (g748)) + ((g721) & (g678) & (!g723) & (sk[10]) & (g744) & (!g748)) + ((g721) & (g678) & (!g723) & (sk[10]) & (g744) & (g748)) + ((g721) & (g678) & (g723) & (!sk[10]) & (!g744) & (!g748)) + ((g721) & (g678) & (g723) & (!sk[10]) & (!g744) & (g748)) + ((g721) & (g678) & (g723) & (!sk[10]) & (g744) & (!g748)) + ((g721) & (g678) & (g723) & (!sk[10]) & (g744) & (g748)) + ((g721) & (g678) & (g723) & (sk[10]) & (g744) & (!g748)) + ((g721) & (g678) & (g723) & (sk[10]) & (g744) & (g748)));
	assign g769 = (((!g720) & (!g722) & (!g727) & (!g747) & (!g742) & (!g768)) + ((!g720) & (!g722) & (!g727) & (g747) & (!g742) & (!g768)) + ((!g720) & (!g722) & (g727) & (!g747) & (!g742) & (!g768)) + ((!g720) & (!g722) & (g727) & (!g747) & (g742) & (!g768)) + ((!g720) & (!g722) & (g727) & (g747) & (!g742) & (!g768)) + ((!g720) & (!g722) & (g727) & (g747) & (g742) & (!g768)) + ((!g720) & (g722) & (!g727) & (!g747) & (!g742) & (!g768)) + ((!g720) & (g722) & (!g727) & (!g747) & (g742) & (!g768)) + ((!g720) & (g722) & (!g727) & (g747) & (!g742) & (!g768)) + ((!g720) & (g722) & (!g727) & (g747) & (g742) & (!g768)) + ((!g720) & (g722) & (g727) & (!g747) & (!g742) & (!g768)) + ((!g720) & (g722) & (g727) & (g747) & (!g742) & (!g768)) + ((g720) & (!g722) & (!g727) & (!g747) & (!g742) & (!g768)) + ((g720) & (!g722) & (!g727) & (!g747) & (g742) & (!g768)) + ((g720) & (!g722) & (g727) & (!g747) & (!g742) & (!g768)) + ((g720) & (g722) & (!g727) & (!g747) & (!g742) & (!g768)) + ((g720) & (g722) & (g727) & (!g747) & (!g742) & (!g768)) + ((g720) & (g722) & (g727) & (!g747) & (g742) & (!g768)));
	assign g770 = (((!g200) & (!g753) & (!g756) & (!g757) & (g767) & (!g769)) + ((!g200) & (!g753) & (!g756) & (g757) & (!g767) & (!g769)) + ((!g200) & (!g753) & (!g756) & (g757) & (g767) & (!g769)) + ((!g200) & (!g753) & (!g756) & (g757) & (g767) & (g769)) + ((!g200) & (!g753) & (g756) & (!g757) & (g767) & (!g769)) + ((!g200) & (!g753) & (g756) & (g757) & (g767) & (!g769)) + ((!g200) & (g753) & (!g756) & (!g757) & (!g767) & (!g769)) + ((!g200) & (g753) & (!g756) & (!g757) & (g767) & (!g769)) + ((!g200) & (g753) & (!g756) & (!g757) & (g767) & (g769)) + ((!g200) & (g753) & (!g756) & (g757) & (!g767) & (!g769)) + ((!g200) & (g753) & (!g756) & (g757) & (g767) & (!g769)) + ((!g200) & (g753) & (!g756) & (g757) & (g767) & (g769)) + ((!g200) & (g753) & (g756) & (!g757) & (g767) & (!g769)) + ((!g200) & (g753) & (g756) & (g757) & (!g767) & (!g769)) + ((!g200) & (g753) & (g756) & (g757) & (g767) & (!g769)) + ((!g200) & (g753) & (g756) & (g757) & (g767) & (g769)) + ((g200) & (!g753) & (!g756) & (!g757) & (g767) & (g769)) + ((g200) & (!g753) & (!g756) & (g757) & (!g767) & (g769)) + ((g200) & (!g753) & (!g756) & (g757) & (g767) & (!g769)) + ((g200) & (!g753) & (!g756) & (g757) & (g767) & (g769)) + ((g200) & (!g753) & (g756) & (!g757) & (g767) & (g769)) + ((g200) & (!g753) & (g756) & (g757) & (g767) & (g769)) + ((g200) & (g753) & (!g756) & (!g757) & (!g767) & (g769)) + ((g200) & (g753) & (!g756) & (!g757) & (g767) & (!g769)) + ((g200) & (g753) & (!g756) & (!g757) & (g767) & (g769)) + ((g200) & (g753) & (!g756) & (g757) & (!g767) & (g769)) + ((g200) & (g753) & (!g756) & (g757) & (g767) & (!g769)) + ((g200) & (g753) & (!g756) & (g757) & (g767) & (g769)) + ((g200) & (g753) & (g756) & (!g757) & (g767) & (g769)) + ((g200) & (g753) & (g756) & (g757) & (!g767) & (g769)) + ((g200) & (g753) & (g756) & (g757) & (g767) & (!g769)) + ((g200) & (g753) & (g756) & (g757) & (g767) & (g769)));
	assign g771 = (((!g585) & (!g597) & (!g679) & (!g720) & (!g722) & (!g727)) + ((!g585) & (!g597) & (!g679) & (!g720) & (g722) & (!g727)) + ((!g585) & (!g597) & (!g679) & (!g720) & (g722) & (g727)) + ((!g585) & (!g597) & (!g679) & (g720) & (!g722) & (!g727)) + ((!g585) & (!g597) & (!g679) & (g720) & (!g722) & (g727)) + ((!g585) & (!g597) & (!g679) & (g720) & (g722) & (g727)) + ((!g585) & (!g597) & (g679) & (!g720) & (!g722) & (g727)) + ((!g585) & (!g597) & (g679) & (g720) & (g722) & (!g727)) + ((!g585) & (g597) & (!g679) & (!g720) & (!g722) & (g727)) + ((!g585) & (g597) & (!g679) & (g720) & (g722) & (!g727)) + ((!g585) & (g597) & (g679) & (!g720) & (!g722) & (!g727)) + ((!g585) & (g597) & (g679) & (!g720) & (g722) & (!g727)) + ((!g585) & (g597) & (g679) & (!g720) & (g722) & (g727)) + ((!g585) & (g597) & (g679) & (g720) & (!g722) & (!g727)) + ((!g585) & (g597) & (g679) & (g720) & (!g722) & (g727)) + ((!g585) & (g597) & (g679) & (g720) & (g722) & (g727)) + ((g585) & (!g597) & (!g679) & (!g720) & (!g722) & (g727)) + ((g585) & (!g597) & (!g679) & (g720) & (g722) & (!g727)) + ((g585) & (!g597) & (g679) & (!g720) & (!g722) & (!g727)) + ((g585) & (!g597) & (g679) & (!g720) & (g722) & (!g727)) + ((g585) & (!g597) & (g679) & (!g720) & (g722) & (g727)) + ((g585) & (!g597) & (g679) & (g720) & (!g722) & (!g727)) + ((g585) & (!g597) & (g679) & (g720) & (!g722) & (g727)) + ((g585) & (!g597) & (g679) & (g720) & (g722) & (g727)) + ((g585) & (g597) & (!g679) & (!g720) & (!g722) & (!g727)) + ((g585) & (g597) & (!g679) & (!g720) & (g722) & (!g727)) + ((g585) & (g597) & (!g679) & (!g720) & (g722) & (g727)) + ((g585) & (g597) & (!g679) & (g720) & (!g722) & (!g727)) + ((g585) & (g597) & (!g679) & (g720) & (!g722) & (g727)) + ((g585) & (g597) & (!g679) & (g720) & (g722) & (g727)) + ((g585) & (g597) & (g679) & (!g720) & (!g722) & (g727)) + ((g585) & (g597) & (g679) & (g720) & (g722) & (!g727)));
	assign g772 = (((!g585) & (!g597) & (!g679) & (g720) & (!g747) & (g744)) + ((!g585) & (!g597) & (!g679) & (g720) & (g747) & (g744)) + ((!g585) & (!g597) & (g679) & (!g720) & (g747) & (!g744)) + ((!g585) & (!g597) & (g679) & (!g720) & (g747) & (g744)) + ((!g585) & (!g597) & (g679) & (g720) & (!g747) & (g744)) + ((!g585) & (!g597) & (g679) & (g720) & (g747) & (!g744)) + ((!g585) & (!g597) & (g679) & (g720) & (g747) & (g744)) + ((!g585) & (g597) & (!g679) & (!g720) & (g747) & (!g744)) + ((!g585) & (g597) & (!g679) & (!g720) & (g747) & (g744)) + ((!g585) & (g597) & (!g679) & (g720) & (!g747) & (g744)) + ((!g585) & (g597) & (!g679) & (g720) & (g747) & (!g744)) + ((!g585) & (g597) & (!g679) & (g720) & (g747) & (g744)) + ((!g585) & (g597) & (g679) & (g720) & (!g747) & (g744)) + ((!g585) & (g597) & (g679) & (g720) & (g747) & (g744)) + ((g585) & (!g597) & (!g679) & (!g720) & (g747) & (!g744)) + ((g585) & (!g597) & (!g679) & (!g720) & (g747) & (g744)) + ((g585) & (!g597) & (!g679) & (g720) & (!g747) & (g744)) + ((g585) & (!g597) & (!g679) & (g720) & (g747) & (!g744)) + ((g585) & (!g597) & (!g679) & (g720) & (g747) & (g744)) + ((g585) & (!g597) & (g679) & (g720) & (!g747) & (g744)) + ((g585) & (!g597) & (g679) & (g720) & (g747) & (g744)) + ((g585) & (g597) & (!g679) & (g720) & (!g747) & (g744)) + ((g585) & (g597) & (!g679) & (g720) & (g747) & (g744)) + ((g585) & (g597) & (g679) & (!g720) & (g747) & (!g744)) + ((g585) & (g597) & (g679) & (!g720) & (g747) & (g744)) + ((g585) & (g597) & (g679) & (g720) & (!g747) & (g744)) + ((g585) & (g597) & (g679) & (g720) & (g747) & (!g744)) + ((g585) & (g597) & (g679) & (g720) & (g747) & (g744)));
	assign g773 = (((!g200) & (!g722) & (!g742) & (!g748) & (!g771) & (!g772)) + ((!g200) & (!g722) & (!g742) & (!g748) & (g771) & (!g772)) + ((!g200) & (!g722) & (g742) & (!g748) & (g771) & (!g772)) + ((!g200) & (g722) & (!g742) & (!g748) & (!g771) & (!g772)) + ((!g200) & (g722) & (!g742) & (!g748) & (g771) & (!g772)) + ((!g200) & (g722) & (!g742) & (g748) & (!g771) & (!g772)) + ((!g200) & (g722) & (!g742) & (g748) & (g771) & (!g772)) + ((!g200) & (g722) & (g742) & (!g748) & (g771) & (!g772)) + ((!g200) & (g722) & (g742) & (g748) & (g771) & (!g772)) + ((g200) & (!g722) & (!g742) & (!g748) & (!g771) & (g772)) + ((g200) & (!g722) & (!g742) & (!g748) & (g771) & (g772)) + ((g200) & (!g722) & (!g742) & (g748) & (!g771) & (!g772)) + ((g200) & (!g722) & (!g742) & (g748) & (!g771) & (g772)) + ((g200) & (!g722) & (!g742) & (g748) & (g771) & (!g772)) + ((g200) & (!g722) & (!g742) & (g748) & (g771) & (g772)) + ((g200) & (!g722) & (g742) & (!g748) & (!g771) & (!g772)) + ((g200) & (!g722) & (g742) & (!g748) & (!g771) & (g772)) + ((g200) & (!g722) & (g742) & (!g748) & (g771) & (g772)) + ((g200) & (!g722) & (g742) & (g748) & (!g771) & (!g772)) + ((g200) & (!g722) & (g742) & (g748) & (!g771) & (g772)) + ((g200) & (!g722) & (g742) & (g748) & (g771) & (!g772)) + ((g200) & (!g722) & (g742) & (g748) & (g771) & (g772)) + ((g200) & (g722) & (!g742) & (!g748) & (!g771) & (g772)) + ((g200) & (g722) & (!g742) & (!g748) & (g771) & (g772)) + ((g200) & (g722) & (!g742) & (g748) & (!g771) & (g772)) + ((g200) & (g722) & (!g742) & (g748) & (g771) & (g772)) + ((g200) & (g722) & (g742) & (!g748) & (!g771) & (!g772)) + ((g200) & (g722) & (g742) & (!g748) & (!g771) & (g772)) + ((g200) & (g722) & (g742) & (!g748) & (g771) & (g772)) + ((g200) & (g722) & (g742) & (g748) & (!g771) & (!g772)) + ((g200) & (g722) & (g742) & (g748) & (!g771) & (g772)) + ((g200) & (g722) & (g742) & (g748) & (g771) & (g772)));
	assign g774 = (((!sk[16]) & (!g746) & (!g759) & (!g763) & (g766)) + ((!sk[16]) & (!g746) & (!g759) & (g763) & (g766)) + ((!sk[16]) & (!g746) & (g759) & (!g763) & (g766)) + ((!sk[16]) & (!g746) & (g759) & (g763) & (g766)) + ((!sk[16]) & (g746) & (!g759) & (!g763) & (!g766)) + ((!sk[16]) & (g746) & (!g759) & (!g763) & (g766)) + ((!sk[16]) & (g746) & (!g759) & (g763) & (!g766)) + ((!sk[16]) & (g746) & (!g759) & (g763) & (g766)) + ((!sk[16]) & (g746) & (g759) & (!g763) & (!g766)) + ((!sk[16]) & (g746) & (g759) & (!g763) & (g766)) + ((!sk[16]) & (g746) & (g759) & (g763) & (!g766)) + ((!sk[16]) & (g746) & (g759) & (g763) & (g766)) + ((sk[16]) & (!g746) & (!g759) & (!g763) & (!g766)) + ((sk[16]) & (g746) & (!g759) & (!g763) & (!g766)) + ((sk[16]) & (g746) & (g759) & (!g763) & (!g766)));
	assign g775 = (((!g723) & (!sk[17]) & (!g724) & (!g725) & (g726) & (!g759)) + ((!g723) & (!sk[17]) & (!g724) & (!g725) & (g726) & (g759)) + ((!g723) & (!sk[17]) & (!g724) & (g725) & (!g726) & (!g759)) + ((!g723) & (!sk[17]) & (!g724) & (g725) & (!g726) & (g759)) + ((!g723) & (!sk[17]) & (!g724) & (g725) & (g726) & (!g759)) + ((!g723) & (!sk[17]) & (!g724) & (g725) & (g726) & (g759)) + ((!g723) & (!sk[17]) & (g724) & (!g725) & (!g726) & (!g759)) + ((!g723) & (!sk[17]) & (g724) & (!g725) & (!g726) & (g759)) + ((!g723) & (!sk[17]) & (g724) & (!g725) & (g726) & (!g759)) + ((!g723) & (!sk[17]) & (g724) & (!g725) & (g726) & (g759)) + ((!g723) & (!sk[17]) & (g724) & (g725) & (!g726) & (!g759)) + ((!g723) & (!sk[17]) & (g724) & (g725) & (!g726) & (g759)) + ((!g723) & (!sk[17]) & (g724) & (g725) & (g726) & (!g759)) + ((!g723) & (!sk[17]) & (g724) & (g725) & (g726) & (g759)) + ((!g723) & (sk[17]) & (!g724) & (!g725) & (g726) & (g759)) + ((!g723) & (sk[17]) & (!g724) & (g725) & (g726) & (g759)) + ((!g723) & (sk[17]) & (g724) & (!g725) & (!g726) & (g759)) + ((!g723) & (sk[17]) & (g724) & (g725) & (!g726) & (g759)) + ((!g723) & (sk[17]) & (g724) & (g725) & (g726) & (g759)) + ((g723) & (!sk[17]) & (!g724) & (!g725) & (g726) & (!g759)) + ((g723) & (!sk[17]) & (!g724) & (!g725) & (g726) & (g759)) + ((g723) & (!sk[17]) & (!g724) & (g725) & (!g726) & (!g759)) + ((g723) & (!sk[17]) & (!g724) & (g725) & (!g726) & (g759)) + ((g723) & (!sk[17]) & (!g724) & (g725) & (g726) & (!g759)) + ((g723) & (!sk[17]) & (!g724) & (g725) & (g726) & (g759)) + ((g723) & (!sk[17]) & (g724) & (!g725) & (!g726) & (!g759)) + ((g723) & (!sk[17]) & (g724) & (!g725) & (!g726) & (g759)) + ((g723) & (!sk[17]) & (g724) & (!g725) & (g726) & (!g759)) + ((g723) & (!sk[17]) & (g724) & (!g725) & (g726) & (g759)) + ((g723) & (!sk[17]) & (g724) & (g725) & (!g726) & (!g759)) + ((g723) & (!sk[17]) & (g724) & (g725) & (!g726) & (g759)) + ((g723) & (!sk[17]) & (g724) & (g725) & (g726) & (!g759)) + ((g723) & (!sk[17]) & (g724) & (g725) & (g726) & (g759)) + ((g723) & (sk[17]) & (!g724) & (!g725) & (!g726) & (g759)) + ((g723) & (sk[17]) & (!g724) & (g725) & (!g726) & (g759)) + ((g723) & (sk[17]) & (g724) & (!g725) & (g726) & (g759)));
	assign g776 = (((!g723) & (!g724) & (!g726) & (!g764) & (!g762) & (!g765)) + ((!g723) & (!g724) & (!g726) & (!g764) & (!g762) & (g765)) + ((!g723) & (!g724) & (g726) & (!g764) & (!g762) & (!g765)) + ((!g723) & (g724) & (!g726) & (!g764) & (!g762) & (!g765)) + ((!g723) & (g724) & (!g726) & (!g764) & (!g762) & (g765)) + ((!g723) & (g724) & (!g726) & (!g764) & (g762) & (!g765)) + ((!g723) & (g724) & (!g726) & (!g764) & (g762) & (g765)) + ((!g723) & (g724) & (g726) & (!g764) & (!g762) & (!g765)) + ((!g723) & (g724) & (g726) & (!g764) & (g762) & (!g765)) + ((g723) & (!g724) & (!g726) & (!g764) & (!g762) & (!g765)) + ((g723) & (!g724) & (!g726) & (!g764) & (!g762) & (g765)) + ((g723) & (!g724) & (!g726) & (g764) & (!g762) & (!g765)) + ((g723) & (!g724) & (!g726) & (g764) & (!g762) & (g765)) + ((g723) & (!g724) & (g726) & (!g764) & (!g762) & (!g765)) + ((g723) & (!g724) & (g726) & (g764) & (!g762) & (!g765)) + ((g723) & (g724) & (!g726) & (!g764) & (!g762) & (!g765)) + ((g723) & (g724) & (!g726) & (!g764) & (!g762) & (g765)) + ((g723) & (g724) & (!g726) & (!g764) & (g762) & (!g765)) + ((g723) & (g724) & (!g726) & (!g764) & (g762) & (g765)) + ((g723) & (g724) & (!g726) & (g764) & (!g762) & (!g765)) + ((g723) & (g724) & (!g726) & (g764) & (!g762) & (g765)) + ((g723) & (g724) & (!g726) & (g764) & (g762) & (!g765)) + ((g723) & (g724) & (!g726) & (g764) & (g762) & (g765)) + ((g723) & (g724) & (g726) & (!g764) & (!g762) & (!g765)) + ((g723) & (g724) & (g726) & (!g764) & (g762) & (!g765)) + ((g723) & (g724) & (g726) & (g764) & (!g762) & (!g765)) + ((g723) & (g724) & (g726) & (g764) & (g762) & (!g765)));
	assign g777 = (((!sk[19]) & (g202) & (g303)) + ((sk[19]) & (!g202) & (g303)) + ((sk[19]) & (g202) & (!g303)));
	assign g778 = (((!g490) & (!g658) & (!sk[20]) & (!g676) & (g777)) + ((!g490) & (!g658) & (!sk[20]) & (g676) & (g777)) + ((!g490) & (!g658) & (sk[20]) & (g676) & (g777)) + ((!g490) & (g658) & (!sk[20]) & (!g676) & (g777)) + ((!g490) & (g658) & (!sk[20]) & (g676) & (g777)) + ((!g490) & (g658) & (sk[20]) & (!g676) & (g777)) + ((g490) & (!g658) & (!sk[20]) & (!g676) & (!g777)) + ((g490) & (!g658) & (!sk[20]) & (!g676) & (g777)) + ((g490) & (!g658) & (!sk[20]) & (g676) & (!g777)) + ((g490) & (!g658) & (!sk[20]) & (g676) & (g777)) + ((g490) & (!g658) & (sk[20]) & (!g676) & (g777)) + ((g490) & (g658) & (!sk[20]) & (!g676) & (!g777)) + ((g490) & (g658) & (!sk[20]) & (!g676) & (g777)) + ((g490) & (g658) & (!sk[20]) & (g676) & (!g777)) + ((g490) & (g658) & (!sk[20]) & (g676) & (g777)) + ((g490) & (g658) & (sk[20]) & (g676) & (g777)));
	assign g779 = (((!g202) & (!g760) & (!g774) & (!g775) & (!g776) & (g778)) + ((!g202) & (!g760) & (!g774) & (!g775) & (g776) & (!g778)) + ((!g202) & (!g760) & (!g774) & (g775) & (!g776) & (g778)) + ((!g202) & (!g760) & (!g774) & (g775) & (g776) & (g778)) + ((!g202) & (!g760) & (g774) & (!g775) & (!g776) & (g778)) + ((!g202) & (!g760) & (g774) & (!g775) & (g776) & (!g778)) + ((!g202) & (!g760) & (g774) & (g775) & (!g776) & (g778)) + ((!g202) & (!g760) & (g774) & (g775) & (g776) & (g778)) + ((!g202) & (g760) & (!g774) & (!g775) & (!g776) & (!g778)) + ((!g202) & (g760) & (!g774) & (!g775) & (g776) & (g778)) + ((!g202) & (g760) & (!g774) & (g775) & (!g776) & (!g778)) + ((!g202) & (g760) & (!g774) & (g775) & (g776) & (!g778)) + ((!g202) & (g760) & (g774) & (!g775) & (!g776) & (g778)) + ((!g202) & (g760) & (g774) & (!g775) & (g776) & (!g778)) + ((!g202) & (g760) & (g774) & (g775) & (!g776) & (g778)) + ((!g202) & (g760) & (g774) & (g775) & (g776) & (g778)) + ((g202) & (!g760) & (!g774) & (!g775) & (!g776) & (!g778)) + ((g202) & (!g760) & (!g774) & (!g775) & (g776) & (g778)) + ((g202) & (!g760) & (!g774) & (g775) & (!g776) & (!g778)) + ((g202) & (!g760) & (!g774) & (g775) & (g776) & (!g778)) + ((g202) & (!g760) & (g774) & (!g775) & (!g776) & (!g778)) + ((g202) & (!g760) & (g774) & (!g775) & (g776) & (g778)) + ((g202) & (!g760) & (g774) & (g775) & (!g776) & (!g778)) + ((g202) & (!g760) & (g774) & (g775) & (g776) & (!g778)) + ((g202) & (g760) & (!g774) & (!g775) & (!g776) & (!g778)) + ((g202) & (g760) & (!g774) & (!g775) & (g776) & (g778)) + ((g202) & (g760) & (!g774) & (g775) & (!g776) & (!g778)) + ((g202) & (g760) & (!g774) & (g775) & (g776) & (!g778)) + ((g202) & (g760) & (g774) & (!g775) & (!g776) & (g778)) + ((g202) & (g760) & (g774) & (!g775) & (g776) & (!g778)) + ((g202) & (g760) & (g774) & (g775) & (!g776) & (g778)) + ((g202) & (g760) & (g774) & (g775) & (g776) & (g778)));
	assign g780 = (((!g770) & (!sk[22]) & (g773) & (!g779)) + ((!g770) & (!sk[22]) & (g773) & (g779)) + ((!g770) & (sk[22]) & (!g773) & (!g779)) + ((g770) & (!sk[22]) & (g773) & (!g779)) + ((g770) & (!sk[22]) & (g773) & (g779)) + ((g770) & (sk[22]) & (!g773) & (!g779)) + ((g770) & (sk[22]) & (!g773) & (g779)) + ((g770) & (sk[22]) & (g773) & (!g779)));
	assign g781 = (((!g202) & (!g760) & (!g774) & (!g775) & (!g776) & (g778)) + ((!g202) & (!g760) & (!g774) & (g775) & (!g776) & (g778)) + ((!g202) & (!g760) & (!g774) & (g775) & (g776) & (g778)) + ((!g202) & (!g760) & (g774) & (!g775) & (!g776) & (g778)) + ((!g202) & (!g760) & (g774) & (g775) & (!g776) & (g778)) + ((!g202) & (!g760) & (g774) & (g775) & (g776) & (g778)) + ((!g202) & (g760) & (!g774) & (!g775) & (!g776) & (!g778)) + ((!g202) & (g760) & (!g774) & (!g775) & (!g776) & (g778)) + ((!g202) & (g760) & (!g774) & (!g775) & (g776) & (g778)) + ((!g202) & (g760) & (!g774) & (g775) & (!g776) & (!g778)) + ((!g202) & (g760) & (!g774) & (g775) & (!g776) & (g778)) + ((!g202) & (g760) & (!g774) & (g775) & (g776) & (!g778)) + ((!g202) & (g760) & (!g774) & (g775) & (g776) & (g778)) + ((!g202) & (g760) & (g774) & (!g775) & (!g776) & (g778)) + ((!g202) & (g760) & (g774) & (g775) & (!g776) & (g778)) + ((!g202) & (g760) & (g774) & (g775) & (g776) & (g778)) + ((g202) & (!g760) & (!g774) & (!g775) & (g776) & (g778)) + ((g202) & (!g760) & (g774) & (!g775) & (g776) & (g778)) + ((g202) & (g760) & (!g774) & (!g775) & (g776) & (g778)) + ((g202) & (g760) & (g774) & (!g775) & (!g776) & (g778)) + ((g202) & (g760) & (g774) & (!g775) & (g776) & (!g778)) + ((g202) & (g760) & (g774) & (!g775) & (g776) & (g778)) + ((g202) & (g760) & (g774) & (g775) & (!g776) & (g778)) + ((g202) & (g760) & (g774) & (g775) & (g776) & (g778)));
	assign g782 = (((!g723) & (!g724) & (!sk[24]) & (!g762) & (g765)) + ((!g723) & (!g724) & (!sk[24]) & (g762) & (g765)) + ((!g723) & (!g724) & (sk[24]) & (!g762) & (g765)) + ((!g723) & (!g724) & (sk[24]) & (g762) & (!g765)) + ((!g723) & (!g724) & (sk[24]) & (g762) & (g765)) + ((!g723) & (g724) & (!sk[24]) & (!g762) & (g765)) + ((!g723) & (g724) & (!sk[24]) & (g762) & (g765)) + ((!g723) & (g724) & (sk[24]) & (g762) & (!g765)) + ((!g723) & (g724) & (sk[24]) & (g762) & (g765)) + ((g723) & (!g724) & (!sk[24]) & (!g762) & (!g765)) + ((g723) & (!g724) & (!sk[24]) & (!g762) & (g765)) + ((g723) & (!g724) & (!sk[24]) & (g762) & (!g765)) + ((g723) & (!g724) & (!sk[24]) & (g762) & (g765)) + ((g723) & (!g724) & (sk[24]) & (!g762) & (g765)) + ((g723) & (!g724) & (sk[24]) & (g762) & (g765)) + ((g723) & (g724) & (!sk[24]) & (!g762) & (!g765)) + ((g723) & (g724) & (!sk[24]) & (!g762) & (g765)) + ((g723) & (g724) & (!sk[24]) & (g762) & (!g765)) + ((g723) & (g724) & (!sk[24]) & (g762) & (g765)));
	assign g783 = (((!g202) & (!g222) & (!g722) & (!g737) & (!g754) & (!g782)) + ((!g202) & (!g222) & (!g722) & (!g737) & (g754) & (!g782)) + ((!g202) & (!g222) & (g722) & (!g737) & (!g754) & (!g782)) + ((!g202) & (!g222) & (g722) & (!g737) & (g754) & (!g782)) + ((!g202) & (!g222) & (g722) & (g737) & (!g754) & (!g782)) + ((!g202) & (!g222) & (g722) & (g737) & (g754) & (!g782)) + ((!g202) & (g222) & (!g722) & (!g737) & (!g754) & (!g782)) + ((!g202) & (g222) & (!g722) & (!g737) & (g754) & (!g782)) + ((!g202) & (g222) & (!g722) & (g737) & (!g754) & (!g782)) + ((!g202) & (g222) & (g722) & (!g737) & (!g754) & (!g782)) + ((!g202) & (g222) & (g722) & (!g737) & (g754) & (!g782)) + ((!g202) & (g222) & (g722) & (g737) & (!g754) & (!g782)) + ((g202) & (!g222) & (!g722) & (!g737) & (!g754) & (g782)) + ((g202) & (!g222) & (!g722) & (!g737) & (g754) & (g782)) + ((g202) & (!g222) & (!g722) & (g737) & (!g754) & (g782)) + ((g202) & (!g222) & (!g722) & (g737) & (g754) & (!g782)) + ((g202) & (!g222) & (!g722) & (g737) & (g754) & (g782)) + ((g202) & (!g222) & (g722) & (!g737) & (!g754) & (g782)) + ((g202) & (!g222) & (g722) & (!g737) & (g754) & (g782)) + ((g202) & (!g222) & (g722) & (g737) & (!g754) & (g782)) + ((g202) & (!g222) & (g722) & (g737) & (g754) & (!g782)) + ((g202) & (!g222) & (g722) & (g737) & (g754) & (g782)) + ((g202) & (g222) & (!g722) & (!g737) & (!g754) & (g782)) + ((g202) & (g222) & (!g722) & (!g737) & (g754) & (g782)) + ((g202) & (g222) & (!g722) & (g737) & (!g754) & (!g782)) + ((g202) & (g222) & (!g722) & (g737) & (!g754) & (g782)) + ((g202) & (g222) & (!g722) & (g737) & (g754) & (!g782)) + ((g202) & (g222) & (!g722) & (g737) & (g754) & (g782)) + ((g202) & (g222) & (g722) & (!g737) & (!g754) & (g782)) + ((g202) & (g222) & (g722) & (!g737) & (g754) & (g782)) + ((g202) & (g222) & (g722) & (g737) & (!g754) & (g782)) + ((g202) & (g222) & (g722) & (g737) & (g754) & (g782)));
	assign g784 = (((!g202) & (!sk[26]) & (!g253) & (!g303) & (g725) & (!g726)) + ((!g202) & (!sk[26]) & (!g253) & (!g303) & (g725) & (g726)) + ((!g202) & (!sk[26]) & (!g253) & (g303) & (!g725) & (!g726)) + ((!g202) & (!sk[26]) & (!g253) & (g303) & (!g725) & (g726)) + ((!g202) & (!sk[26]) & (!g253) & (g303) & (g725) & (!g726)) + ((!g202) & (!sk[26]) & (!g253) & (g303) & (g725) & (g726)) + ((!g202) & (!sk[26]) & (g253) & (!g303) & (!g725) & (!g726)) + ((!g202) & (!sk[26]) & (g253) & (!g303) & (!g725) & (g726)) + ((!g202) & (!sk[26]) & (g253) & (!g303) & (g725) & (!g726)) + ((!g202) & (!sk[26]) & (g253) & (!g303) & (g725) & (g726)) + ((!g202) & (!sk[26]) & (g253) & (g303) & (!g725) & (!g726)) + ((!g202) & (!sk[26]) & (g253) & (g303) & (!g725) & (g726)) + ((!g202) & (!sk[26]) & (g253) & (g303) & (g725) & (!g726)) + ((!g202) & (!sk[26]) & (g253) & (g303) & (g725) & (g726)) + ((!g202) & (sk[26]) & (!g253) & (g303) & (!g725) & (g726)) + ((!g202) & (sk[26]) & (!g253) & (g303) & (g725) & (g726)) + ((!g202) & (sk[26]) & (g253) & (!g303) & (!g725) & (!g726)) + ((!g202) & (sk[26]) & (g253) & (!g303) & (!g725) & (g726)) + ((!g202) & (sk[26]) & (g253) & (g303) & (!g725) & (!g726)) + ((!g202) & (sk[26]) & (g253) & (g303) & (g725) & (g726)) + ((g202) & (!sk[26]) & (!g253) & (!g303) & (g725) & (!g726)) + ((g202) & (!sk[26]) & (!g253) & (!g303) & (g725) & (g726)) + ((g202) & (!sk[26]) & (!g253) & (g303) & (!g725) & (!g726)) + ((g202) & (!sk[26]) & (!g253) & (g303) & (!g725) & (g726)) + ((g202) & (!sk[26]) & (!g253) & (g303) & (g725) & (!g726)) + ((g202) & (!sk[26]) & (!g253) & (g303) & (g725) & (g726)) + ((g202) & (!sk[26]) & (g253) & (!g303) & (!g725) & (!g726)) + ((g202) & (!sk[26]) & (g253) & (!g303) & (!g725) & (g726)) + ((g202) & (!sk[26]) & (g253) & (!g303) & (g725) & (!g726)) + ((g202) & (!sk[26]) & (g253) & (!g303) & (g725) & (g726)) + ((g202) & (!sk[26]) & (g253) & (g303) & (!g725) & (!g726)) + ((g202) & (!sk[26]) & (g253) & (g303) & (!g725) & (g726)) + ((g202) & (!sk[26]) & (g253) & (g303) & (g725) & (!g726)) + ((g202) & (!sk[26]) & (g253) & (g303) & (g725) & (g726)) + ((g202) & (sk[26]) & (!g253) & (!g303) & (!g725) & (g726)) + ((g202) & (sk[26]) & (!g253) & (!g303) & (g725) & (g726)) + ((g202) & (sk[26]) & (!g253) & (g303) & (!g725) & (!g726)) + ((g202) & (sk[26]) & (!g253) & (g303) & (!g725) & (g726)) + ((g202) & (sk[26]) & (g253) & (!g303) & (!g725) & (!g726)) + ((g202) & (sk[26]) & (g253) & (!g303) & (g725) & (g726)));
	assign g785 = (((!sk[27]) & (!g781) & (g783) & (!g784)) + ((!sk[27]) & (!g781) & (g783) & (g784)) + ((!sk[27]) & (g781) & (g783) & (!g784)) + ((!sk[27]) & (g781) & (g783) & (g784)) + ((sk[27]) & (!g781) & (!g783) & (g784)) + ((sk[27]) & (!g781) & (g783) & (!g784)) + ((sk[27]) & (g781) & (!g783) & (!g784)) + ((sk[27]) & (g781) & (g783) & (g784)));
	assign g786 = (((!g585) & (!g597) & (!g679) & (g720) & (!g744) & (g748)) + ((!g585) & (!g597) & (!g679) & (g720) & (g744) & (g748)) + ((!g585) & (!g597) & (g679) & (!g720) & (g744) & (!g748)) + ((!g585) & (!g597) & (g679) & (!g720) & (g744) & (g748)) + ((!g585) & (!g597) & (g679) & (g720) & (!g744) & (g748)) + ((!g585) & (!g597) & (g679) & (g720) & (g744) & (!g748)) + ((!g585) & (!g597) & (g679) & (g720) & (g744) & (g748)) + ((!g585) & (g597) & (!g679) & (!g720) & (g744) & (!g748)) + ((!g585) & (g597) & (!g679) & (!g720) & (g744) & (g748)) + ((!g585) & (g597) & (!g679) & (g720) & (!g744) & (g748)) + ((!g585) & (g597) & (!g679) & (g720) & (g744) & (!g748)) + ((!g585) & (g597) & (!g679) & (g720) & (g744) & (g748)) + ((!g585) & (g597) & (g679) & (g720) & (!g744) & (g748)) + ((!g585) & (g597) & (g679) & (g720) & (g744) & (g748)) + ((g585) & (!g597) & (!g679) & (!g720) & (g744) & (!g748)) + ((g585) & (!g597) & (!g679) & (!g720) & (g744) & (g748)) + ((g585) & (!g597) & (!g679) & (g720) & (!g744) & (g748)) + ((g585) & (!g597) & (!g679) & (g720) & (g744) & (!g748)) + ((g585) & (!g597) & (!g679) & (g720) & (g744) & (g748)) + ((g585) & (!g597) & (g679) & (g720) & (!g744) & (g748)) + ((g585) & (!g597) & (g679) & (g720) & (g744) & (g748)) + ((g585) & (g597) & (!g679) & (g720) & (!g744) & (g748)) + ((g585) & (g597) & (!g679) & (g720) & (g744) & (g748)) + ((g585) & (g597) & (g679) & (!g720) & (g744) & (!g748)) + ((g585) & (g597) & (g679) & (!g720) & (g744) & (g748)) + ((g585) & (g597) & (g679) & (g720) & (!g744) & (g748)) + ((g585) & (g597) & (g679) & (g720) & (g744) & (!g748)) + ((g585) & (g597) & (g679) & (g720) & (g744) & (g748)));
	assign g787 = (((!g719) & (!g728) & (!g729) & (!g747) & (!g742) & (!g786)) + ((!g719) & (!g728) & (!g729) & (!g747) & (g742) & (!g786)) + ((!g719) & (!g728) & (g729) & (!g747) & (!g742) & (!g786)) + ((!g719) & (!g728) & (g729) & (g747) & (!g742) & (!g786)) + ((!g719) & (g728) & (!g729) & (!g747) & (!g742) & (!g786)) + ((!g719) & (g728) & (g729) & (!g747) & (!g742) & (!g786)) + ((!g719) & (g728) & (g729) & (!g747) & (g742) & (!g786)) + ((!g719) & (g728) & (g729) & (g747) & (!g742) & (!g786)) + ((!g719) & (g728) & (g729) & (g747) & (g742) & (!g786)) + ((g719) & (!g728) & (!g729) & (!g747) & (!g742) & (!g786)) + ((g719) & (!g728) & (g729) & (!g747) & (!g742) & (!g786)) + ((g719) & (!g728) & (g729) & (!g747) & (g742) & (!g786)) + ((g719) & (!g728) & (g729) & (g747) & (!g742) & (!g786)) + ((g719) & (!g728) & (g729) & (g747) & (g742) & (!g786)) + ((g719) & (g728) & (!g729) & (!g747) & (!g742) & (!g786)) + ((g719) & (g728) & (!g729) & (!g747) & (g742) & (!g786)) + ((g719) & (g728) & (g729) & (!g747) & (!g742) & (!g786)) + ((g719) & (g728) & (g729) & (g747) & (!g742) & (!g786)));
	assign g788 = (((!sk[30]) & (!g200) & (g785) & (!g787)) + ((!sk[30]) & (!g200) & (g785) & (g787)) + ((!sk[30]) & (g200) & (g785) & (!g787)) + ((!sk[30]) & (g200) & (g785) & (g787)) + ((sk[30]) & (!g200) & (!g785) & (!g787)) + ((sk[30]) & (!g200) & (g785) & (g787)) + ((sk[30]) & (g200) & (!g785) & (g787)) + ((sk[30]) & (g200) & (g785) & (!g787)));
	assign g789 = (((!g753) & (!g756) & (sk[31]) & (g757)) + ((!g753) & (g756) & (!sk[31]) & (!g757)) + ((!g753) & (g756) & (!sk[31]) & (g757)) + ((g753) & (!g756) & (sk[31]) & (!g757)) + ((g753) & (!g756) & (sk[31]) & (g757)) + ((g753) & (g756) & (!sk[31]) & (!g757)) + ((g753) & (g756) & (!sk[31]) & (g757)) + ((g753) & (g756) & (sk[31]) & (g757)));
	assign g790 = (((!g200) & (!g767) & (sk[32]) & (!g769)) + ((!g200) & (g767) & (!sk[32]) & (!g769)) + ((!g200) & (g767) & (!sk[32]) & (g769)) + ((!g200) & (g767) & (sk[32]) & (g769)) + ((g200) & (!g767) & (sk[32]) & (g769)) + ((g200) & (g767) & (!sk[32]) & (!g769)) + ((g200) & (g767) & (!sk[32]) & (g769)) + ((g200) & (g767) & (sk[32]) & (!g769)));
	assign g791 = (((!g549) & (!g569) & (!g680) & (!g719) & (g728) & (g729)) + ((!g549) & (!g569) & (!g680) & (g719) & (!g728) & (!g729)) + ((!g549) & (!g569) & (g680) & (!g719) & (!g728) & (!g729)) + ((!g549) & (!g569) & (g680) & (!g719) & (!g728) & (g729)) + ((!g549) & (!g569) & (g680) & (!g719) & (g728) & (!g729)) + ((!g549) & (!g569) & (g680) & (g719) & (!g728) & (g729)) + ((!g549) & (!g569) & (g680) & (g719) & (g728) & (!g729)) + ((!g549) & (!g569) & (g680) & (g719) & (g728) & (g729)) + ((!g549) & (g569) & (!g680) & (!g719) & (!g728) & (!g729)) + ((!g549) & (g569) & (!g680) & (!g719) & (!g728) & (g729)) + ((!g549) & (g569) & (!g680) & (!g719) & (g728) & (!g729)) + ((!g549) & (g569) & (!g680) & (g719) & (!g728) & (g729)) + ((!g549) & (g569) & (!g680) & (g719) & (g728) & (!g729)) + ((!g549) & (g569) & (!g680) & (g719) & (g728) & (g729)) + ((!g549) & (g569) & (g680) & (!g719) & (g728) & (g729)) + ((!g549) & (g569) & (g680) & (g719) & (!g728) & (!g729)) + ((g549) & (!g569) & (!g680) & (!g719) & (!g728) & (!g729)) + ((g549) & (!g569) & (!g680) & (!g719) & (!g728) & (g729)) + ((g549) & (!g569) & (!g680) & (!g719) & (g728) & (!g729)) + ((g549) & (!g569) & (!g680) & (g719) & (!g728) & (g729)) + ((g549) & (!g569) & (!g680) & (g719) & (g728) & (!g729)) + ((g549) & (!g569) & (!g680) & (g719) & (g728) & (g729)) + ((g549) & (!g569) & (g680) & (!g719) & (g728) & (g729)) + ((g549) & (!g569) & (g680) & (g719) & (!g728) & (!g729)) + ((g549) & (g569) & (!g680) & (!g719) & (g728) & (g729)) + ((g549) & (g569) & (!g680) & (g719) & (!g728) & (!g729)) + ((g549) & (g569) & (g680) & (!g719) & (!g728) & (!g729)) + ((g549) & (g569) & (g680) & (!g719) & (!g728) & (g729)) + ((g549) & (g569) & (g680) & (!g719) & (g728) & (!g729)) + ((g549) & (g569) & (g680) & (g719) & (!g728) & (g729)) + ((g549) & (g569) & (g680) & (g719) & (g728) & (!g729)) + ((g549) & (g569) & (g680) & (g719) & (g728) & (g729)));
	assign g792 = (((!g549) & (!g569) & (!g680) & (!g733) & (g734) & (!g729)) + ((!g549) & (!g569) & (!g680) & (g733) & (g734) & (!g729)) + ((!g549) & (!g569) & (g680) & (!g733) & (g734) & (!g729)) + ((!g549) & (!g569) & (g680) & (g733) & (!g734) & (!g729)) + ((!g549) & (!g569) & (g680) & (g733) & (!g734) & (g729)) + ((!g549) & (!g569) & (g680) & (g733) & (g734) & (!g729)) + ((!g549) & (!g569) & (g680) & (g733) & (g734) & (g729)) + ((!g549) & (g569) & (!g680) & (!g733) & (g734) & (!g729)) + ((!g549) & (g569) & (!g680) & (g733) & (!g734) & (!g729)) + ((!g549) & (g569) & (!g680) & (g733) & (!g734) & (g729)) + ((!g549) & (g569) & (!g680) & (g733) & (g734) & (!g729)) + ((!g549) & (g569) & (!g680) & (g733) & (g734) & (g729)) + ((!g549) & (g569) & (g680) & (!g733) & (g734) & (!g729)) + ((!g549) & (g569) & (g680) & (g733) & (g734) & (!g729)) + ((g549) & (!g569) & (!g680) & (!g733) & (g734) & (!g729)) + ((g549) & (!g569) & (!g680) & (g733) & (!g734) & (!g729)) + ((g549) & (!g569) & (!g680) & (g733) & (!g734) & (g729)) + ((g549) & (!g569) & (!g680) & (g733) & (g734) & (!g729)) + ((g549) & (!g569) & (!g680) & (g733) & (g734) & (g729)) + ((g549) & (!g569) & (g680) & (!g733) & (g734) & (!g729)) + ((g549) & (!g569) & (g680) & (g733) & (g734) & (!g729)) + ((g549) & (g569) & (!g680) & (!g733) & (g734) & (!g729)) + ((g549) & (g569) & (!g680) & (g733) & (g734) & (!g729)) + ((g549) & (g569) & (g680) & (!g733) & (g734) & (!g729)) + ((g549) & (g569) & (g680) & (g733) & (!g734) & (!g729)) + ((g549) & (g569) & (g680) & (g733) & (!g734) & (g729)) + ((g549) & (g569) & (g680) & (g733) & (g734) & (!g729)) + ((g549) & (g569) & (g680) & (g733) & (g734) & (g729)));
	assign g793 = (((!g2) & (!g686) & (!g719) & (!g732) & (!g791) & (!g792)) + ((!g2) & (!g686) & (!g719) & (!g732) & (g791) & (!g792)) + ((!g2) & (!g686) & (!g719) & (g732) & (!g791) & (!g792)) + ((!g2) & (!g686) & (g719) & (!g732) & (!g791) & (!g792)) + ((!g2) & (!g686) & (g719) & (!g732) & (g791) & (!g792)) + ((!g2) & (!g686) & (g719) & (g732) & (!g791) & (!g792)) + ((!g2) & (g686) & (g719) & (!g732) & (!g791) & (!g792)) + ((!g2) & (g686) & (g719) & (!g732) & (g791) & (!g792)) + ((!g2) & (g686) & (g719) & (g732) & (!g791) & (!g792)) + ((g2) & (!g686) & (!g719) & (!g732) & (!g791) & (g792)) + ((g2) & (!g686) & (!g719) & (!g732) & (g791) & (g792)) + ((g2) & (!g686) & (!g719) & (g732) & (!g791) & (g792)) + ((g2) & (!g686) & (!g719) & (g732) & (g791) & (!g792)) + ((g2) & (!g686) & (!g719) & (g732) & (g791) & (g792)) + ((g2) & (!g686) & (g719) & (!g732) & (!g791) & (g792)) + ((g2) & (!g686) & (g719) & (!g732) & (g791) & (g792)) + ((g2) & (!g686) & (g719) & (g732) & (!g791) & (g792)) + ((g2) & (!g686) & (g719) & (g732) & (g791) & (!g792)) + ((g2) & (!g686) & (g719) & (g732) & (g791) & (g792)) + ((g2) & (g686) & (!g719) & (!g732) & (!g791) & (!g792)) + ((g2) & (g686) & (!g719) & (!g732) & (!g791) & (g792)) + ((g2) & (g686) & (!g719) & (!g732) & (g791) & (!g792)) + ((g2) & (g686) & (!g719) & (!g732) & (g791) & (g792)) + ((g2) & (g686) & (!g719) & (g732) & (!g791) & (!g792)) + ((g2) & (g686) & (!g719) & (g732) & (!g791) & (g792)) + ((g2) & (g686) & (!g719) & (g732) & (g791) & (!g792)) + ((g2) & (g686) & (!g719) & (g732) & (g791) & (g792)) + ((g2) & (g686) & (g719) & (!g732) & (!g791) & (g792)) + ((g2) & (g686) & (g719) & (!g732) & (g791) & (g792)) + ((g2) & (g686) & (g719) & (g732) & (!g791) & (g792)) + ((g2) & (g686) & (g719) & (g732) & (g791) & (!g792)) + ((g2) & (g686) & (g719) & (g732) & (g791) & (g792)));
	assign g794 = (((!sk[36]) & (!g686) & (!g734) & (!g723) & (g724)) + ((!sk[36]) & (!g686) & (!g734) & (g723) & (g724)) + ((!sk[36]) & (!g686) & (g734) & (!g723) & (g724)) + ((!sk[36]) & (!g686) & (g734) & (g723) & (g724)) + ((!sk[36]) & (g686) & (!g734) & (!g723) & (!g724)) + ((!sk[36]) & (g686) & (!g734) & (!g723) & (g724)) + ((!sk[36]) & (g686) & (!g734) & (g723) & (!g724)) + ((!sk[36]) & (g686) & (!g734) & (g723) & (g724)) + ((!sk[36]) & (g686) & (g734) & (!g723) & (!g724)) + ((!sk[36]) & (g686) & (g734) & (!g723) & (g724)) + ((!sk[36]) & (g686) & (g734) & (g723) & (!g724)) + ((!sk[36]) & (g686) & (g734) & (g723) & (g724)) + ((sk[36]) & (!g686) & (g734) & (!g723) & (!g724)) + ((sk[36]) & (!g686) & (g734) & (!g723) & (g724)) + ((sk[36]) & (g686) & (!g734) & (!g723) & (!g724)) + ((sk[36]) & (g686) & (!g734) & (g723) & (!g724)) + ((sk[36]) & (g686) & (g734) & (!g723) & (!g724)) + ((sk[36]) & (g686) & (g734) & (!g723) & (g724)) + ((sk[36]) & (g686) & (g734) & (g723) & (!g724)));
	assign g795 = (((!g2) & (!g401) & (!g684) & (!g722) & (!g754) & (!g794)) + ((!g2) & (!g401) & (!g684) & (!g722) & (g754) & (!g794)) + ((!g2) & (!g401) & (!g684) & (g722) & (!g754) & (!g794)) + ((!g2) & (!g401) & (!g684) & (g722) & (g754) & (!g794)) + ((!g2) & (!g401) & (g684) & (g722) & (!g754) & (!g794)) + ((!g2) & (!g401) & (g684) & (g722) & (g754) & (!g794)) + ((!g2) & (g401) & (!g684) & (!g722) & (!g754) & (!g794)) + ((!g2) & (g401) & (!g684) & (!g722) & (g754) & (!g794)) + ((!g2) & (g401) & (!g684) & (g722) & (!g754) & (!g794)) + ((!g2) & (g401) & (!g684) & (g722) & (g754) & (!g794)) + ((!g2) & (g401) & (g684) & (!g722) & (!g754) & (!g794)) + ((!g2) & (g401) & (g684) & (g722) & (!g754) & (!g794)) + ((g2) & (!g401) & (!g684) & (!g722) & (!g754) & (g794)) + ((g2) & (!g401) & (!g684) & (!g722) & (g754) & (g794)) + ((g2) & (!g401) & (!g684) & (g722) & (!g754) & (g794)) + ((g2) & (!g401) & (!g684) & (g722) & (g754) & (g794)) + ((g2) & (!g401) & (g684) & (!g722) & (!g754) & (g794)) + ((g2) & (!g401) & (g684) & (!g722) & (g754) & (!g794)) + ((g2) & (!g401) & (g684) & (!g722) & (g754) & (g794)) + ((g2) & (!g401) & (g684) & (g722) & (!g754) & (g794)) + ((g2) & (!g401) & (g684) & (g722) & (g754) & (!g794)) + ((g2) & (!g401) & (g684) & (g722) & (g754) & (g794)) + ((g2) & (g401) & (!g684) & (!g722) & (!g754) & (g794)) + ((g2) & (g401) & (!g684) & (!g722) & (g754) & (g794)) + ((g2) & (g401) & (!g684) & (g722) & (!g754) & (g794)) + ((g2) & (g401) & (!g684) & (g722) & (g754) & (g794)) + ((g2) & (g401) & (g684) & (!g722) & (!g754) & (!g794)) + ((g2) & (g401) & (g684) & (!g722) & (!g754) & (g794)) + ((g2) & (g401) & (g684) & (!g722) & (g754) & (!g794)) + ((g2) & (g401) & (g684) & (!g722) & (g754) & (g794)) + ((g2) & (g401) & (g684) & (g722) & (!g754) & (g794)) + ((g2) & (g401) & (g684) & (g722) & (g754) & (g794)));
	assign g796 = (((!g2) & (!g198) & (!sk[38]) & (!g367) & (g725) & (!g726)) + ((!g2) & (!g198) & (!sk[38]) & (!g367) & (g725) & (g726)) + ((!g2) & (!g198) & (!sk[38]) & (g367) & (!g725) & (!g726)) + ((!g2) & (!g198) & (!sk[38]) & (g367) & (!g725) & (g726)) + ((!g2) & (!g198) & (!sk[38]) & (g367) & (g725) & (!g726)) + ((!g2) & (!g198) & (!sk[38]) & (g367) & (g725) & (g726)) + ((!g2) & (!g198) & (sk[38]) & (g367) & (!g725) & (g726)) + ((!g2) & (!g198) & (sk[38]) & (g367) & (g725) & (g726)) + ((!g2) & (g198) & (!sk[38]) & (!g367) & (!g725) & (!g726)) + ((!g2) & (g198) & (!sk[38]) & (!g367) & (!g725) & (g726)) + ((!g2) & (g198) & (!sk[38]) & (!g367) & (g725) & (!g726)) + ((!g2) & (g198) & (!sk[38]) & (!g367) & (g725) & (g726)) + ((!g2) & (g198) & (!sk[38]) & (g367) & (!g725) & (!g726)) + ((!g2) & (g198) & (!sk[38]) & (g367) & (!g725) & (g726)) + ((!g2) & (g198) & (!sk[38]) & (g367) & (g725) & (!g726)) + ((!g2) & (g198) & (!sk[38]) & (g367) & (g725) & (g726)) + ((!g2) & (g198) & (sk[38]) & (!g367) & (!g725) & (!g726)) + ((!g2) & (g198) & (sk[38]) & (!g367) & (!g725) & (g726)) + ((!g2) & (g198) & (sk[38]) & (g367) & (!g725) & (!g726)) + ((!g2) & (g198) & (sk[38]) & (g367) & (g725) & (g726)) + ((g2) & (!g198) & (!sk[38]) & (!g367) & (g725) & (!g726)) + ((g2) & (!g198) & (!sk[38]) & (!g367) & (g725) & (g726)) + ((g2) & (!g198) & (!sk[38]) & (g367) & (!g725) & (!g726)) + ((g2) & (!g198) & (!sk[38]) & (g367) & (!g725) & (g726)) + ((g2) & (!g198) & (!sk[38]) & (g367) & (g725) & (!g726)) + ((g2) & (!g198) & (!sk[38]) & (g367) & (g725) & (g726)) + ((g2) & (!g198) & (sk[38]) & (!g367) & (!g725) & (g726)) + ((g2) & (!g198) & (sk[38]) & (!g367) & (g725) & (g726)) + ((g2) & (!g198) & (sk[38]) & (g367) & (!g725) & (!g726)) + ((g2) & (!g198) & (sk[38]) & (g367) & (!g725) & (g726)) + ((g2) & (g198) & (!sk[38]) & (!g367) & (!g725) & (!g726)) + ((g2) & (g198) & (!sk[38]) & (!g367) & (!g725) & (g726)) + ((g2) & (g198) & (!sk[38]) & (!g367) & (g725) & (!g726)) + ((g2) & (g198) & (!sk[38]) & (!g367) & (g725) & (g726)) + ((g2) & (g198) & (!sk[38]) & (g367) & (!g725) & (!g726)) + ((g2) & (g198) & (!sk[38]) & (g367) & (!g725) & (g726)) + ((g2) & (g198) & (!sk[38]) & (g367) & (g725) & (!g726)) + ((g2) & (g198) & (!sk[38]) & (g367) & (g725) & (g726)) + ((g2) & (g198) & (sk[38]) & (!g367) & (!g725) & (!g726)) + ((g2) & (g198) & (sk[38]) & (!g367) & (g725) & (g726)));
	assign g797 = (((!g490) & (!g658) & (!sk[39]) & (!g676) & (g741)) + ((!g490) & (!g658) & (!sk[39]) & (g676) & (g741)) + ((!g490) & (!g658) & (sk[39]) & (g676) & (g741)) + ((!g490) & (g658) & (!sk[39]) & (!g676) & (g741)) + ((!g490) & (g658) & (!sk[39]) & (g676) & (g741)) + ((!g490) & (g658) & (sk[39]) & (!g676) & (g741)) + ((g490) & (!g658) & (!sk[39]) & (!g676) & (!g741)) + ((g490) & (!g658) & (!sk[39]) & (!g676) & (g741)) + ((g490) & (!g658) & (!sk[39]) & (g676) & (!g741)) + ((g490) & (!g658) & (!sk[39]) & (g676) & (g741)) + ((g490) & (!g658) & (sk[39]) & (!g676) & (g741)) + ((g490) & (g658) & (!sk[39]) & (!g676) & (!g741)) + ((g490) & (g658) & (!sk[39]) & (!g676) & (g741)) + ((g490) & (g658) & (!sk[39]) & (g676) & (!g741)) + ((g490) & (g658) & (!sk[39]) & (g676) & (g741)) + ((g490) & (g658) & (sk[39]) & (g676) & (g741)));
	assign g798 = (((!sk[40]) & (g734) & (g726)) + ((sk[40]) & (g734) & (g726)));
	assign g799 = (((!g641) & (!g655) & (!g677) & (!g733) & (g686) & (!g725)) + ((!g641) & (!g655) & (!g677) & (g733) & (g686) & (!g725)) + ((!g641) & (!g655) & (g677) & (!g733) & (g686) & (!g725)) + ((!g641) & (!g655) & (g677) & (g733) & (!g686) & (!g725)) + ((!g641) & (!g655) & (g677) & (g733) & (!g686) & (g725)) + ((!g641) & (!g655) & (g677) & (g733) & (g686) & (!g725)) + ((!g641) & (!g655) & (g677) & (g733) & (g686) & (g725)) + ((!g641) & (g655) & (!g677) & (!g733) & (g686) & (!g725)) + ((!g641) & (g655) & (!g677) & (g733) & (!g686) & (!g725)) + ((!g641) & (g655) & (!g677) & (g733) & (!g686) & (g725)) + ((!g641) & (g655) & (!g677) & (g733) & (g686) & (!g725)) + ((!g641) & (g655) & (!g677) & (g733) & (g686) & (g725)) + ((!g641) & (g655) & (g677) & (!g733) & (g686) & (!g725)) + ((!g641) & (g655) & (g677) & (g733) & (g686) & (!g725)) + ((g641) & (!g655) & (!g677) & (!g733) & (g686) & (!g725)) + ((g641) & (!g655) & (!g677) & (g733) & (!g686) & (!g725)) + ((g641) & (!g655) & (!g677) & (g733) & (!g686) & (g725)) + ((g641) & (!g655) & (!g677) & (g733) & (g686) & (!g725)) + ((g641) & (!g655) & (!g677) & (g733) & (g686) & (g725)) + ((g641) & (!g655) & (g677) & (!g733) & (g686) & (!g725)) + ((g641) & (!g655) & (g677) & (g733) & (g686) & (!g725)) + ((g641) & (g655) & (!g677) & (!g733) & (g686) & (!g725)) + ((g641) & (g655) & (!g677) & (g733) & (g686) & (!g725)) + ((g641) & (g655) & (g677) & (!g733) & (g686) & (!g725)) + ((g641) & (g655) & (g677) & (g733) & (!g686) & (!g725)) + ((g641) & (g655) & (g677) & (g733) & (!g686) & (g725)) + ((g641) & (g655) & (g677) & (g733) & (g686) & (!g725)) + ((g641) & (g655) & (g677) & (g733) & (g686) & (g725)));
	assign g800 = (((!g732) & (!sk[42]) & (!g746) & (!g798) & (g799)) + ((!g732) & (!sk[42]) & (!g746) & (g798) & (g799)) + ((!g732) & (!sk[42]) & (g746) & (!g798) & (g799)) + ((!g732) & (!sk[42]) & (g746) & (g798) & (g799)) + ((!g732) & (sk[42]) & (!g746) & (!g798) & (!g799)) + ((!g732) & (sk[42]) & (g746) & (!g798) & (!g799)) + ((g732) & (!sk[42]) & (!g746) & (!g798) & (!g799)) + ((g732) & (!sk[42]) & (!g746) & (!g798) & (g799)) + ((g732) & (!sk[42]) & (!g746) & (g798) & (!g799)) + ((g732) & (!sk[42]) & (!g746) & (g798) & (g799)) + ((g732) & (!sk[42]) & (g746) & (!g798) & (!g799)) + ((g732) & (!sk[42]) & (g746) & (!g798) & (g799)) + ((g732) & (!sk[42]) & (g746) & (g798) & (!g799)) + ((g732) & (!sk[42]) & (g746) & (g798) & (g799)) + ((g732) & (sk[42]) & (g746) & (!g798) & (!g799)));
	assign g801 = (((g2) & (!g401) & (!g414) & (!g683) & (!g725) & (!g726)) + ((g2) & (!g401) & (!g414) & (!g683) & (!g725) & (g726)) + ((g2) & (!g401) & (!g414) & (!g683) & (g725) & (!g726)) + ((g2) & (!g401) & (!g414) & (!g683) & (g725) & (g726)) + ((g2) & (!g401) & (!g414) & (g683) & (g725) & (!g726)) + ((g2) & (!g401) & (g414) & (!g683) & (g725) & (!g726)) + ((g2) & (!g401) & (g414) & (g683) & (g725) & (!g726)) + ((g2) & (!g401) & (g414) & (g683) & (g725) & (g726)) + ((g2) & (g401) & (!g414) & (!g683) & (g725) & (!g726)) + ((g2) & (g401) & (!g414) & (!g683) & (g725) & (g726)) + ((g2) & (g401) & (!g414) & (g683) & (g725) & (!g726)) + ((g2) & (g401) & (g414) & (!g683) & (g725) & (!g726)) + ((g2) & (g401) & (g414) & (g683) & (!g725) & (!g726)) + ((g2) & (g401) & (g414) & (g683) & (!g725) & (g726)) + ((g2) & (g401) & (g414) & (g683) & (g725) & (!g726)) + ((g2) & (g401) & (g414) & (g683) & (g725) & (g726)));
	assign g802 = (((!g723) & (!g724) & (!g725) & (!sk[44]) & (g726) & (!g732)) + ((!g723) & (!g724) & (!g725) & (!sk[44]) & (g726) & (g732)) + ((!g723) & (!g724) & (!g725) & (sk[44]) & (g726) & (g732)) + ((!g723) & (!g724) & (g725) & (!sk[44]) & (!g726) & (!g732)) + ((!g723) & (!g724) & (g725) & (!sk[44]) & (!g726) & (g732)) + ((!g723) & (!g724) & (g725) & (!sk[44]) & (g726) & (!g732)) + ((!g723) & (!g724) & (g725) & (!sk[44]) & (g726) & (g732)) + ((!g723) & (!g724) & (g725) & (sk[44]) & (g726) & (g732)) + ((!g723) & (g724) & (!g725) & (!sk[44]) & (!g726) & (!g732)) + ((!g723) & (g724) & (!g725) & (!sk[44]) & (!g726) & (g732)) + ((!g723) & (g724) & (!g725) & (!sk[44]) & (g726) & (!g732)) + ((!g723) & (g724) & (!g725) & (!sk[44]) & (g726) & (g732)) + ((!g723) & (g724) & (!g725) & (sk[44]) & (!g726) & (g732)) + ((!g723) & (g724) & (g725) & (!sk[44]) & (!g726) & (!g732)) + ((!g723) & (g724) & (g725) & (!sk[44]) & (!g726) & (g732)) + ((!g723) & (g724) & (g725) & (!sk[44]) & (g726) & (!g732)) + ((!g723) & (g724) & (g725) & (!sk[44]) & (g726) & (g732)) + ((!g723) & (g724) & (g725) & (sk[44]) & (!g726) & (g732)) + ((!g723) & (g724) & (g725) & (sk[44]) & (g726) & (g732)) + ((g723) & (!g724) & (!g725) & (!sk[44]) & (g726) & (!g732)) + ((g723) & (!g724) & (!g725) & (!sk[44]) & (g726) & (g732)) + ((g723) & (!g724) & (!g725) & (sk[44]) & (!g726) & (g732)) + ((g723) & (!g724) & (g725) & (!sk[44]) & (!g726) & (!g732)) + ((g723) & (!g724) & (g725) & (!sk[44]) & (!g726) & (g732)) + ((g723) & (!g724) & (g725) & (!sk[44]) & (g726) & (!g732)) + ((g723) & (!g724) & (g725) & (!sk[44]) & (g726) & (g732)) + ((g723) & (!g724) & (g725) & (sk[44]) & (!g726) & (g732)) + ((g723) & (g724) & (!g725) & (!sk[44]) & (!g726) & (!g732)) + ((g723) & (g724) & (!g725) & (!sk[44]) & (!g726) & (g732)) + ((g723) & (g724) & (!g725) & (!sk[44]) & (g726) & (!g732)) + ((g723) & (g724) & (!g725) & (!sk[44]) & (g726) & (g732)) + ((g723) & (g724) & (!g725) & (sk[44]) & (g726) & (g732)) + ((g723) & (g724) & (g725) & (!sk[44]) & (!g726) & (!g732)) + ((g723) & (g724) & (g725) & (!sk[44]) & (!g726) & (g732)) + ((g723) & (g724) & (g725) & (!sk[44]) & (g726) & (!g732)) + ((g723) & (g724) & (g725) & (!sk[44]) & (g726) & (g732)));
	assign g803 = (((!g733) & (!g686) & (!g734) & (!g723) & (!g724) & (!g726)) + ((!g733) & (!g686) & (!g734) & (!g723) & (!g724) & (g726)) + ((!g733) & (!g686) & (!g734) & (!g723) & (g724) & (!g726)) + ((!g733) & (!g686) & (!g734) & (!g723) & (g724) & (g726)) + ((!g733) & (!g686) & (!g734) & (g723) & (!g724) & (!g726)) + ((!g733) & (!g686) & (!g734) & (g723) & (!g724) & (g726)) + ((!g733) & (!g686) & (!g734) & (g723) & (g724) & (!g726)) + ((!g733) & (!g686) & (!g734) & (g723) & (g724) & (g726)) + ((!g733) & (!g686) & (g734) & (!g723) & (g724) & (!g726)) + ((!g733) & (!g686) & (g734) & (!g723) & (g724) & (g726)) + ((!g733) & (!g686) & (g734) & (g723) & (g724) & (!g726)) + ((!g733) & (!g686) & (g734) & (g723) & (g724) & (g726)) + ((!g733) & (g686) & (!g734) & (!g723) & (!g724) & (!g726)) + ((!g733) & (g686) & (!g734) & (!g723) & (g724) & (!g726)) + ((!g733) & (g686) & (!g734) & (g723) & (!g724) & (!g726)) + ((!g733) & (g686) & (!g734) & (g723) & (g724) & (!g726)) + ((!g733) & (g686) & (g734) & (!g723) & (g724) & (!g726)) + ((!g733) & (g686) & (g734) & (g723) & (g724) & (!g726)) + ((g733) & (!g686) & (!g734) & (g723) & (!g724) & (!g726)) + ((g733) & (!g686) & (!g734) & (g723) & (!g724) & (g726)) + ((g733) & (!g686) & (!g734) & (g723) & (g724) & (!g726)) + ((g733) & (!g686) & (!g734) & (g723) & (g724) & (g726)) + ((g733) & (!g686) & (g734) & (g723) & (g724) & (!g726)) + ((g733) & (!g686) & (g734) & (g723) & (g724) & (g726)) + ((g733) & (g686) & (!g734) & (g723) & (!g724) & (!g726)) + ((g733) & (g686) & (!g734) & (g723) & (g724) & (!g726)) + ((g733) & (g686) & (g734) & (g723) & (g724) & (!g726)));
	assign g804 = (((!g2) & (!g797) & (!g800) & (g801) & (!g802) & (!g803)) + ((!g2) & (!g797) & (!g800) & (g801) & (g802) & (!g803)) + ((!g2) & (!g797) & (!g800) & (g801) & (g802) & (g803)) + ((!g2) & (g797) & (!g800) & (!g801) & (!g802) & (!g803)) + ((!g2) & (g797) & (!g800) & (!g801) & (g802) & (!g803)) + ((!g2) & (g797) & (!g800) & (!g801) & (g802) & (g803)) + ((!g2) & (g797) & (!g800) & (g801) & (!g802) & (!g803)) + ((!g2) & (g797) & (!g800) & (g801) & (!g802) & (g803)) + ((!g2) & (g797) & (!g800) & (g801) & (g802) & (!g803)) + ((!g2) & (g797) & (!g800) & (g801) & (g802) & (g803)) + ((!g2) & (g797) & (g800) & (!g801) & (!g802) & (!g803)) + ((!g2) & (g797) & (g800) & (!g801) & (g802) & (!g803)) + ((!g2) & (g797) & (g800) & (!g801) & (g802) & (g803)) + ((!g2) & (g797) & (g800) & (g801) & (!g802) & (!g803)) + ((!g2) & (g797) & (g800) & (g801) & (g802) & (!g803)) + ((!g2) & (g797) & (g800) & (g801) & (g802) & (g803)) + ((g2) & (!g797) & (g800) & (g801) & (!g802) & (g803)) + ((g2) & (g797) & (!g800) & (!g801) & (!g802) & (g803)) + ((g2) & (g797) & (!g800) & (g801) & (!g802) & (g803)) + ((g2) & (g797) & (g800) & (!g801) & (!g802) & (g803)) + ((g2) & (g797) & (g800) & (g801) & (!g802) & (!g803)) + ((g2) & (g797) & (g800) & (g801) & (!g802) & (g803)) + ((g2) & (g797) & (g800) & (g801) & (g802) & (!g803)) + ((g2) & (g797) & (g800) & (g801) & (g802) & (g803)));
	assign g805 = (((!g721) & (!sk[47]) & (!g678) & (!g686) & (g734) & (!g723)) + ((!g721) & (!sk[47]) & (!g678) & (!g686) & (g734) & (g723)) + ((!g721) & (!sk[47]) & (!g678) & (g686) & (!g734) & (!g723)) + ((!g721) & (!sk[47]) & (!g678) & (g686) & (!g734) & (g723)) + ((!g721) & (!sk[47]) & (!g678) & (g686) & (g734) & (!g723)) + ((!g721) & (!sk[47]) & (!g678) & (g686) & (g734) & (g723)) + ((!g721) & (!sk[47]) & (g678) & (!g686) & (!g734) & (!g723)) + ((!g721) & (!sk[47]) & (g678) & (!g686) & (!g734) & (g723)) + ((!g721) & (!sk[47]) & (g678) & (!g686) & (g734) & (!g723)) + ((!g721) & (!sk[47]) & (g678) & (!g686) & (g734) & (g723)) + ((!g721) & (!sk[47]) & (g678) & (g686) & (!g734) & (!g723)) + ((!g721) & (!sk[47]) & (g678) & (g686) & (!g734) & (g723)) + ((!g721) & (!sk[47]) & (g678) & (g686) & (g734) & (!g723)) + ((!g721) & (!sk[47]) & (g678) & (g686) & (g734) & (g723)) + ((!g721) & (sk[47]) & (!g678) & (!g686) & (g734) & (!g723)) + ((!g721) & (sk[47]) & (!g678) & (!g686) & (g734) & (g723)) + ((!g721) & (sk[47]) & (!g678) & (g686) & (!g734) & (!g723)) + ((!g721) & (sk[47]) & (!g678) & (g686) & (g734) & (!g723)) + ((!g721) & (sk[47]) & (!g678) & (g686) & (g734) & (g723)) + ((!g721) & (sk[47]) & (g678) & (g686) & (!g734) & (!g723)) + ((!g721) & (sk[47]) & (g678) & (g686) & (g734) & (!g723)) + ((g721) & (!sk[47]) & (!g678) & (!g686) & (g734) & (!g723)) + ((g721) & (!sk[47]) & (!g678) & (!g686) & (g734) & (g723)) + ((g721) & (!sk[47]) & (!g678) & (g686) & (!g734) & (!g723)) + ((g721) & (!sk[47]) & (!g678) & (g686) & (!g734) & (g723)) + ((g721) & (!sk[47]) & (!g678) & (g686) & (g734) & (!g723)) + ((g721) & (!sk[47]) & (!g678) & (g686) & (g734) & (g723)) + ((g721) & (!sk[47]) & (g678) & (!g686) & (!g734) & (!g723)) + ((g721) & (!sk[47]) & (g678) & (!g686) & (!g734) & (g723)) + ((g721) & (!sk[47]) & (g678) & (!g686) & (g734) & (!g723)) + ((g721) & (!sk[47]) & (g678) & (!g686) & (g734) & (g723)) + ((g721) & (!sk[47]) & (g678) & (g686) & (!g734) & (!g723)) + ((g721) & (!sk[47]) & (g678) & (g686) & (!g734) & (g723)) + ((g721) & (!sk[47]) & (g678) & (g686) & (g734) & (!g723)) + ((g721) & (!sk[47]) & (g678) & (g686) & (g734) & (g723)) + ((g721) & (sk[47]) & (!g678) & (g686) & (!g734) & (!g723)) + ((g721) & (sk[47]) & (!g678) & (g686) & (g734) & (!g723)) + ((g721) & (sk[47]) & (g678) & (!g686) & (g734) & (!g723)) + ((g721) & (sk[47]) & (g678) & (!g686) & (g734) & (g723)) + ((g721) & (sk[47]) & (g678) & (g686) & (!g734) & (!g723)) + ((g721) & (sk[47]) & (g678) & (g686) & (g734) & (!g723)) + ((g721) & (sk[47]) & (g678) & (g686) & (g734) & (g723)));
	assign g806 = (((!g733) & (!g720) & (!g722) & (!g727) & (!g732) & (!g805)) + ((!g733) & (!g720) & (!g722) & (g727) & (!g732) & (!g805)) + ((!g733) & (!g720) & (!g722) & (g727) & (g732) & (!g805)) + ((!g733) & (!g720) & (g722) & (!g727) & (!g732) & (!g805)) + ((!g733) & (!g720) & (g722) & (!g727) & (g732) & (!g805)) + ((!g733) & (!g720) & (g722) & (g727) & (!g732) & (!g805)) + ((!g733) & (g720) & (!g722) & (!g727) & (!g732) & (!g805)) + ((!g733) & (g720) & (!g722) & (!g727) & (g732) & (!g805)) + ((!g733) & (g720) & (!g722) & (g727) & (!g732) & (!g805)) + ((!g733) & (g720) & (g722) & (!g727) & (!g732) & (!g805)) + ((!g733) & (g720) & (g722) & (g727) & (!g732) & (!g805)) + ((!g733) & (g720) & (g722) & (g727) & (g732) & (!g805)) + ((g733) & (!g720) & (!g722) & (!g727) & (!g732) & (!g805)) + ((g733) & (!g720) & (!g722) & (g727) & (!g732) & (!g805)) + ((g733) & (!g720) & (!g722) & (g727) & (g732) & (!g805)) + ((g733) & (!g720) & (g722) & (!g727) & (!g732) & (!g805)) + ((g733) & (!g720) & (g722) & (!g727) & (g732) & (!g805)) + ((g733) & (!g720) & (g722) & (g727) & (!g732) & (!g805)));
	assign g807 = (((!g200) & (!g742) & (!g739) & (!g745) & (!g746) & (g749)) + ((!g200) & (!g742) & (!g739) & (!g745) & (g746) & (g749)) + ((!g200) & (!g742) & (!g739) & (g745) & (!g746) & (!g749)) + ((!g200) & (!g742) & (!g739) & (g745) & (!g746) & (g749)) + ((!g200) & (!g742) & (!g739) & (g745) & (g746) & (!g749)) + ((!g200) & (!g742) & (!g739) & (g745) & (g746) & (g749)) + ((!g200) & (!g742) & (g739) & (!g745) & (!g746) & (!g749)) + ((!g200) & (!g742) & (g739) & (!g745) & (g746) & (!g749)) + ((!g200) & (g742) & (!g739) & (!g745) & (!g746) & (!g749)) + ((!g200) & (g742) & (!g739) & (!g745) & (!g746) & (g749)) + ((!g200) & (g742) & (!g739) & (!g745) & (g746) & (g749)) + ((!g200) & (g742) & (!g739) & (g745) & (!g746) & (!g749)) + ((!g200) & (g742) & (!g739) & (g745) & (!g746) & (g749)) + ((!g200) & (g742) & (!g739) & (g745) & (g746) & (!g749)) + ((!g200) & (g742) & (!g739) & (g745) & (g746) & (g749)) + ((!g200) & (g742) & (g739) & (!g745) & (g746) & (!g749)) + ((g200) & (!g742) & (!g739) & (!g745) & (!g746) & (!g749)) + ((g200) & (!g742) & (!g739) & (!g745) & (g746) & (!g749)) + ((g200) & (!g742) & (g739) & (!g745) & (!g746) & (g749)) + ((g200) & (!g742) & (g739) & (!g745) & (g746) & (g749)) + ((g200) & (!g742) & (g739) & (g745) & (!g746) & (!g749)) + ((g200) & (!g742) & (g739) & (g745) & (!g746) & (g749)) + ((g200) & (!g742) & (g739) & (g745) & (g746) & (!g749)) + ((g200) & (!g742) & (g739) & (g745) & (g746) & (g749)) + ((g200) & (g742) & (!g739) & (!g745) & (g746) & (!g749)) + ((g200) & (g742) & (g739) & (!g745) & (!g746) & (!g749)) + ((g200) & (g742) & (g739) & (!g745) & (!g746) & (g749)) + ((g200) & (g742) & (g739) & (!g745) & (g746) & (g749)) + ((g200) & (g742) & (g739) & (g745) & (!g746) & (!g749)) + ((g200) & (g742) & (g739) & (g745) & (!g746) & (g749)) + ((g200) & (g742) & (g739) & (g745) & (g746) & (!g749)) + ((g200) & (g742) & (g739) & (g745) & (g746) & (g749)));
	assign g808 = (((!g2) & (!g795) & (!g796) & (!g804) & (!g806) & (g807)) + ((!g2) & (!g795) & (!g796) & (g804) & (!g806) & (!g807)) + ((!g2) & (!g795) & (!g796) & (g804) & (!g806) & (g807)) + ((!g2) & (!g795) & (!g796) & (g804) & (g806) & (g807)) + ((!g2) & (!g795) & (g796) & (!g804) & (!g806) & (!g807)) + ((!g2) & (!g795) & (g796) & (!g804) & (!g806) & (g807)) + ((!g2) & (!g795) & (g796) & (!g804) & (g806) & (g807)) + ((!g2) & (!g795) & (g796) & (g804) & (!g806) & (!g807)) + ((!g2) & (!g795) & (g796) & (g804) & (!g806) & (g807)) + ((!g2) & (!g795) & (g796) & (g804) & (g806) & (g807)) + ((!g2) & (g795) & (!g796) & (!g804) & (!g806) & (g807)) + ((!g2) & (g795) & (!g796) & (g804) & (!g806) & (g807)) + ((!g2) & (g795) & (g796) & (!g804) & (!g806) & (g807)) + ((!g2) & (g795) & (g796) & (g804) & (!g806) & (!g807)) + ((!g2) & (g795) & (g796) & (g804) & (!g806) & (g807)) + ((!g2) & (g795) & (g796) & (g804) & (g806) & (g807)) + ((g2) & (!g795) & (!g796) & (!g804) & (g806) & (g807)) + ((g2) & (!g795) & (!g796) & (g804) & (!g806) & (g807)) + ((g2) & (!g795) & (!g796) & (g804) & (g806) & (!g807)) + ((g2) & (!g795) & (!g796) & (g804) & (g806) & (g807)) + ((g2) & (!g795) & (g796) & (!g804) & (!g806) & (g807)) + ((g2) & (!g795) & (g796) & (!g804) & (g806) & (!g807)) + ((g2) & (!g795) & (g796) & (!g804) & (g806) & (g807)) + ((g2) & (!g795) & (g796) & (g804) & (!g806) & (g807)) + ((g2) & (!g795) & (g796) & (g804) & (g806) & (!g807)) + ((g2) & (!g795) & (g796) & (g804) & (g806) & (g807)) + ((g2) & (g795) & (!g796) & (!g804) & (g806) & (g807)) + ((g2) & (g795) & (!g796) & (g804) & (g806) & (g807)) + ((g2) & (g795) & (g796) & (!g804) & (g806) & (g807)) + ((g2) & (g795) & (g796) & (g804) & (!g806) & (g807)) + ((g2) & (g795) & (g796) & (g804) & (g806) & (!g807)) + ((g2) & (g795) & (g796) & (g804) & (g806) & (g807)));
	assign g809 = (((!g585) & (!g597) & (!g679) & (!g733) & (g734) & (g720)) + ((!g585) & (!g597) & (!g679) & (g733) & (g734) & (g720)) + ((!g585) & (!g597) & (g679) & (!g733) & (g734) & (g720)) + ((!g585) & (!g597) & (g679) & (g733) & (!g734) & (!g720)) + ((!g585) & (!g597) & (g679) & (g733) & (!g734) & (g720)) + ((!g585) & (!g597) & (g679) & (g733) & (g734) & (!g720)) + ((!g585) & (!g597) & (g679) & (g733) & (g734) & (g720)) + ((!g585) & (g597) & (!g679) & (!g733) & (g734) & (g720)) + ((!g585) & (g597) & (!g679) & (g733) & (!g734) & (!g720)) + ((!g585) & (g597) & (!g679) & (g733) & (!g734) & (g720)) + ((!g585) & (g597) & (!g679) & (g733) & (g734) & (!g720)) + ((!g585) & (g597) & (!g679) & (g733) & (g734) & (g720)) + ((!g585) & (g597) & (g679) & (!g733) & (g734) & (g720)) + ((!g585) & (g597) & (g679) & (g733) & (g734) & (g720)) + ((g585) & (!g597) & (!g679) & (!g733) & (g734) & (g720)) + ((g585) & (!g597) & (!g679) & (g733) & (!g734) & (!g720)) + ((g585) & (!g597) & (!g679) & (g733) & (!g734) & (g720)) + ((g585) & (!g597) & (!g679) & (g733) & (g734) & (!g720)) + ((g585) & (!g597) & (!g679) & (g733) & (g734) & (g720)) + ((g585) & (!g597) & (g679) & (!g733) & (g734) & (g720)) + ((g585) & (!g597) & (g679) & (g733) & (g734) & (g720)) + ((g585) & (g597) & (!g679) & (!g733) & (g734) & (g720)) + ((g585) & (g597) & (!g679) & (g733) & (g734) & (g720)) + ((g585) & (g597) & (g679) & (!g733) & (g734) & (g720)) + ((g585) & (g597) & (g679) & (g733) & (!g734) & (!g720)) + ((g585) & (g597) & (g679) & (g733) & (!g734) & (g720)) + ((g585) & (g597) & (g679) & (g733) & (g734) & (!g720)) + ((g585) & (g597) & (g679) & (g733) & (g734) & (g720)));
	assign g810 = (((!g2) & (!g686) & (!g722) & (!g732) & (!g771) & (!g809)) + ((!g2) & (!g686) & (!g722) & (!g732) & (g771) & (!g809)) + ((!g2) & (!g686) & (!g722) & (g732) & (g771) & (!g809)) + ((!g2) & (!g686) & (g722) & (!g732) & (!g771) & (!g809)) + ((!g2) & (!g686) & (g722) & (!g732) & (g771) & (!g809)) + ((!g2) & (!g686) & (g722) & (g732) & (g771) & (!g809)) + ((!g2) & (g686) & (g722) & (!g732) & (!g771) & (!g809)) + ((!g2) & (g686) & (g722) & (!g732) & (g771) & (!g809)) + ((!g2) & (g686) & (g722) & (g732) & (g771) & (!g809)) + ((g2) & (!g686) & (!g722) & (!g732) & (!g771) & (g809)) + ((g2) & (!g686) & (!g722) & (!g732) & (g771) & (g809)) + ((g2) & (!g686) & (!g722) & (g732) & (!g771) & (!g809)) + ((g2) & (!g686) & (!g722) & (g732) & (!g771) & (g809)) + ((g2) & (!g686) & (!g722) & (g732) & (g771) & (g809)) + ((g2) & (!g686) & (g722) & (!g732) & (!g771) & (g809)) + ((g2) & (!g686) & (g722) & (!g732) & (g771) & (g809)) + ((g2) & (!g686) & (g722) & (g732) & (!g771) & (!g809)) + ((g2) & (!g686) & (g722) & (g732) & (!g771) & (g809)) + ((g2) & (!g686) & (g722) & (g732) & (g771) & (g809)) + ((g2) & (g686) & (!g722) & (!g732) & (!g771) & (!g809)) + ((g2) & (g686) & (!g722) & (!g732) & (!g771) & (g809)) + ((g2) & (g686) & (!g722) & (!g732) & (g771) & (!g809)) + ((g2) & (g686) & (!g722) & (!g732) & (g771) & (g809)) + ((g2) & (g686) & (!g722) & (g732) & (!g771) & (!g809)) + ((g2) & (g686) & (!g722) & (g732) & (!g771) & (g809)) + ((g2) & (g686) & (!g722) & (g732) & (g771) & (!g809)) + ((g2) & (g686) & (!g722) & (g732) & (g771) & (g809)) + ((g2) & (g686) & (g722) & (!g732) & (!g771) & (g809)) + ((g2) & (g686) & (g722) & (!g732) & (g771) & (g809)) + ((g2) & (g686) & (g722) & (g732) & (!g771) & (!g809)) + ((g2) & (g686) & (g722) & (g732) & (!g771) & (g809)) + ((g2) & (g686) & (g722) & (g732) & (g771) & (g809)));
	assign g811 = (((!g200) & (!g738) & (!g739) & (!g750) & (!g751) & (g752)) + ((!g200) & (!g738) & (!g739) & (g750) & (!g751) & (g752)) + ((!g200) & (!g738) & (g739) & (!g750) & (!g751) & (!g752)) + ((!g200) & (!g738) & (g739) & (!g750) & (g751) & (!g752)) + ((!g200) & (!g738) & (g739) & (!g750) & (g751) & (g752)) + ((!g200) & (!g738) & (g739) & (g750) & (!g751) & (g752)) + ((!g200) & (g738) & (!g739) & (!g750) & (!g751) & (!g752)) + ((!g200) & (g738) & (!g739) & (!g750) & (g751) & (!g752)) + ((!g200) & (g738) & (!g739) & (!g750) & (g751) & (g752)) + ((!g200) & (g738) & (!g739) & (g750) & (!g751) & (!g752)) + ((!g200) & (g738) & (!g739) & (g750) & (g751) & (!g752)) + ((!g200) & (g738) & (!g739) & (g750) & (g751) & (g752)) + ((!g200) & (g738) & (g739) & (!g750) & (!g751) & (g752)) + ((!g200) & (g738) & (g739) & (g750) & (!g751) & (!g752)) + ((!g200) & (g738) & (g739) & (g750) & (g751) & (!g752)) + ((!g200) & (g738) & (g739) & (g750) & (g751) & (g752)) + ((g200) & (!g738) & (!g739) & (!g750) & (!g751) & (!g752)) + ((g200) & (!g738) & (!g739) & (!g750) & (g751) & (!g752)) + ((g200) & (!g738) & (!g739) & (!g750) & (g751) & (g752)) + ((g200) & (!g738) & (!g739) & (g750) & (!g751) & (!g752)) + ((g200) & (!g738) & (!g739) & (g750) & (g751) & (!g752)) + ((g200) & (!g738) & (!g739) & (g750) & (g751) & (g752)) + ((g200) & (!g738) & (g739) & (!g750) & (!g751) & (!g752)) + ((g200) & (!g738) & (g739) & (!g750) & (g751) & (!g752)) + ((g200) & (!g738) & (g739) & (!g750) & (g751) & (g752)) + ((g200) & (!g738) & (g739) & (g750) & (!g751) & (g752)) + ((g200) & (g738) & (!g739) & (!g750) & (!g751) & (g752)) + ((g200) & (g738) & (!g739) & (g750) & (!g751) & (g752)) + ((g200) & (g738) & (g739) & (!g750) & (!g751) & (g752)) + ((g200) & (g738) & (g739) & (g750) & (!g751) & (!g752)) + ((g200) & (g738) & (g739) & (g750) & (g751) & (!g752)) + ((g200) & (g738) & (g739) & (g750) & (g751) & (g752)));
	assign g812 = (((!g585) & (!g597) & (!g679) & (g686) & (!g734) & (g720)) + ((!g585) & (!g597) & (!g679) & (g686) & (g734) & (g720)) + ((!g585) & (!g597) & (g679) & (!g686) & (g734) & (!g720)) + ((!g585) & (!g597) & (g679) & (!g686) & (g734) & (g720)) + ((!g585) & (!g597) & (g679) & (g686) & (!g734) & (g720)) + ((!g585) & (!g597) & (g679) & (g686) & (g734) & (!g720)) + ((!g585) & (!g597) & (g679) & (g686) & (g734) & (g720)) + ((!g585) & (g597) & (!g679) & (!g686) & (g734) & (!g720)) + ((!g585) & (g597) & (!g679) & (!g686) & (g734) & (g720)) + ((!g585) & (g597) & (!g679) & (g686) & (!g734) & (g720)) + ((!g585) & (g597) & (!g679) & (g686) & (g734) & (!g720)) + ((!g585) & (g597) & (!g679) & (g686) & (g734) & (g720)) + ((!g585) & (g597) & (g679) & (g686) & (!g734) & (g720)) + ((!g585) & (g597) & (g679) & (g686) & (g734) & (g720)) + ((g585) & (!g597) & (!g679) & (!g686) & (g734) & (!g720)) + ((g585) & (!g597) & (!g679) & (!g686) & (g734) & (g720)) + ((g585) & (!g597) & (!g679) & (g686) & (!g734) & (g720)) + ((g585) & (!g597) & (!g679) & (g686) & (g734) & (!g720)) + ((g585) & (!g597) & (!g679) & (g686) & (g734) & (g720)) + ((g585) & (!g597) & (g679) & (g686) & (!g734) & (g720)) + ((g585) & (!g597) & (g679) & (g686) & (g734) & (g720)) + ((g585) & (g597) & (!g679) & (g686) & (!g734) & (g720)) + ((g585) & (g597) & (!g679) & (g686) & (g734) & (g720)) + ((g585) & (g597) & (g679) & (!g686) & (g734) & (!g720)) + ((g585) & (g597) & (g679) & (!g686) & (g734) & (g720)) + ((g585) & (g597) & (g679) & (g686) & (!g734) & (g720)) + ((g585) & (g597) & (g679) & (g686) & (g734) & (!g720)) + ((g585) & (g597) & (g679) & (g686) & (g734) & (g720)));
	assign g813 = (((!g733) & (!g719) & (!g728) & (!g729) & (!g732) & (!g812)) + ((!g733) & (!g719) & (!g728) & (!g729) & (g732) & (!g812)) + ((!g733) & (!g719) & (!g728) & (g729) & (!g732) & (!g812)) + ((!g733) & (!g719) & (g728) & (!g729) & (!g732) & (!g812)) + ((!g733) & (!g719) & (g728) & (g729) & (!g732) & (!g812)) + ((!g733) & (!g719) & (g728) & (g729) & (g732) & (!g812)) + ((!g733) & (g719) & (!g728) & (!g729) & (!g732) & (!g812)) + ((!g733) & (g719) & (!g728) & (g729) & (!g732) & (!g812)) + ((!g733) & (g719) & (!g728) & (g729) & (g732) & (!g812)) + ((!g733) & (g719) & (g728) & (!g729) & (!g732) & (!g812)) + ((!g733) & (g719) & (g728) & (!g729) & (g732) & (!g812)) + ((!g733) & (g719) & (g728) & (g729) & (!g732) & (!g812)) + ((g733) & (!g719) & (!g728) & (g729) & (!g732) & (!g812)) + ((g733) & (!g719) & (g728) & (g729) & (!g732) & (!g812)) + ((g733) & (!g719) & (g728) & (g729) & (g732) & (!g812)) + ((g733) & (g719) & (!g728) & (g729) & (!g732) & (!g812)) + ((g733) & (g719) & (!g728) & (g729) & (g732) & (!g812)) + ((g733) & (g719) & (g728) & (g729) & (!g732) & (!g812)));
	assign g814 = (((!g753) & (!g756) & (sk[56]) & (g757)) + ((!g753) & (g756) & (!sk[56]) & (!g757)) + ((!g753) & (g756) & (!sk[56]) & (g757)) + ((!g753) & (g756) & (sk[56]) & (!g757)) + ((g753) & (!g756) & (sk[56]) & (!g757)) + ((g753) & (g756) & (!sk[56]) & (!g757)) + ((g753) & (g756) & (!sk[56]) & (g757)) + ((g753) & (g756) & (sk[56]) & (g757)));
	assign g815 = (((!g2) & (!g808) & (!g810) & (!g811) & (!g813) & (!g814)) + ((!g2) & (!g808) & (!g810) & (!g811) & (!g813) & (g814)) + ((!g2) & (!g808) & (!g810) & (!g811) & (g813) & (!g814)) + ((!g2) & (!g808) & (!g810) & (g811) & (!g813) & (!g814)) + ((!g2) & (!g808) & (g810) & (!g811) & (!g813) & (!g814)) + ((!g2) & (!g808) & (g810) & (g811) & (!g813) & (!g814)) + ((!g2) & (g808) & (!g810) & (!g811) & (!g813) & (!g814)) + ((!g2) & (g808) & (!g810) & (!g811) & (!g813) & (g814)) + ((!g2) & (g808) & (!g810) & (!g811) & (g813) & (!g814)) + ((!g2) & (g808) & (!g810) & (g811) & (!g813) & (!g814)) + ((!g2) & (g808) & (!g810) & (g811) & (!g813) & (g814)) + ((!g2) & (g808) & (!g810) & (g811) & (g813) & (!g814)) + ((!g2) & (g808) & (g810) & (!g811) & (!g813) & (!g814)) + ((!g2) & (g808) & (g810) & (!g811) & (!g813) & (g814)) + ((!g2) & (g808) & (g810) & (!g811) & (g813) & (!g814)) + ((!g2) & (g808) & (g810) & (g811) & (!g813) & (!g814)) + ((g2) & (!g808) & (!g810) & (!g811) & (!g813) & (!g814)) + ((g2) & (!g808) & (!g810) & (!g811) & (g813) & (!g814)) + ((g2) & (!g808) & (!g810) & (!g811) & (g813) & (g814)) + ((g2) & (!g808) & (!g810) & (g811) & (g813) & (!g814)) + ((g2) & (!g808) & (g810) & (!g811) & (g813) & (!g814)) + ((g2) & (!g808) & (g810) & (g811) & (g813) & (!g814)) + ((g2) & (g808) & (!g810) & (!g811) & (!g813) & (!g814)) + ((g2) & (g808) & (!g810) & (!g811) & (g813) & (!g814)) + ((g2) & (g808) & (!g810) & (!g811) & (g813) & (g814)) + ((g2) & (g808) & (!g810) & (g811) & (!g813) & (!g814)) + ((g2) & (g808) & (!g810) & (g811) & (g813) & (!g814)) + ((g2) & (g808) & (!g810) & (g811) & (g813) & (g814)) + ((g2) & (g808) & (g810) & (!g811) & (!g813) & (!g814)) + ((g2) & (g808) & (g810) & (!g811) & (g813) & (!g814)) + ((g2) & (g808) & (g810) & (!g811) & (g813) & (g814)) + ((g2) & (g808) & (g810) & (g811) & (g813) & (!g814)));
	assign g816 = (((!g708) & (!sk[58]) & (!g716) & (!g549) & (g569) & (!g680)) + ((!g708) & (!sk[58]) & (!g716) & (!g549) & (g569) & (g680)) + ((!g708) & (!sk[58]) & (!g716) & (g549) & (!g569) & (!g680)) + ((!g708) & (!sk[58]) & (!g716) & (g549) & (!g569) & (g680)) + ((!g708) & (!sk[58]) & (!g716) & (g549) & (g569) & (!g680)) + ((!g708) & (!sk[58]) & (!g716) & (g549) & (g569) & (g680)) + ((!g708) & (!sk[58]) & (g716) & (!g549) & (!g569) & (!g680)) + ((!g708) & (!sk[58]) & (g716) & (!g549) & (!g569) & (g680)) + ((!g708) & (!sk[58]) & (g716) & (!g549) & (g569) & (!g680)) + ((!g708) & (!sk[58]) & (g716) & (!g549) & (g569) & (g680)) + ((!g708) & (!sk[58]) & (g716) & (g549) & (!g569) & (!g680)) + ((!g708) & (!sk[58]) & (g716) & (g549) & (!g569) & (g680)) + ((!g708) & (!sk[58]) & (g716) & (g549) & (g569) & (!g680)) + ((!g708) & (!sk[58]) & (g716) & (g549) & (g569) & (g680)) + ((!g708) & (sk[58]) & (!g716) & (!g549) & (g569) & (g680)) + ((!g708) & (sk[58]) & (!g716) & (g549) & (!g569) & (!g680)) + ((!g708) & (sk[58]) & (g716) & (!g549) & (!g569) & (!g680)) + ((!g708) & (sk[58]) & (g716) & (!g549) & (!g569) & (g680)) + ((!g708) & (sk[58]) & (g716) & (!g549) & (g569) & (!g680)) + ((!g708) & (sk[58]) & (g716) & (g549) & (!g569) & (g680)) + ((!g708) & (sk[58]) & (g716) & (g549) & (g569) & (!g680)) + ((!g708) & (sk[58]) & (g716) & (g549) & (g569) & (g680)) + ((g708) & (!sk[58]) & (!g716) & (!g549) & (g569) & (!g680)) + ((g708) & (!sk[58]) & (!g716) & (!g549) & (g569) & (g680)) + ((g708) & (!sk[58]) & (!g716) & (g549) & (!g569) & (!g680)) + ((g708) & (!sk[58]) & (!g716) & (g549) & (!g569) & (g680)) + ((g708) & (!sk[58]) & (!g716) & (g549) & (g569) & (!g680)) + ((g708) & (!sk[58]) & (!g716) & (g549) & (g569) & (g680)) + ((g708) & (!sk[58]) & (g716) & (!g549) & (!g569) & (!g680)) + ((g708) & (!sk[58]) & (g716) & (!g549) & (!g569) & (g680)) + ((g708) & (!sk[58]) & (g716) & (!g549) & (g569) & (!g680)) + ((g708) & (!sk[58]) & (g716) & (!g549) & (g569) & (g680)) + ((g708) & (!sk[58]) & (g716) & (g549) & (!g569) & (!g680)) + ((g708) & (!sk[58]) & (g716) & (g549) & (!g569) & (g680)) + ((g708) & (!sk[58]) & (g716) & (g549) & (g569) & (!g680)) + ((g708) & (!sk[58]) & (g716) & (g549) & (g569) & (g680)) + ((g708) & (sk[58]) & (!g716) & (!g549) & (!g569) & (!g680)) + ((g708) & (sk[58]) & (!g716) & (!g549) & (!g569) & (g680)) + ((g708) & (sk[58]) & (!g716) & (!g549) & (g569) & (!g680)) + ((g708) & (sk[58]) & (!g716) & (g549) & (!g569) & (g680)) + ((g708) & (sk[58]) & (!g716) & (g549) & (g569) & (!g680)) + ((g708) & (sk[58]) & (!g716) & (g549) & (g569) & (g680)) + ((g708) & (sk[58]) & (g716) & (!g549) & (g569) & (g680)) + ((g708) & (sk[58]) & (g716) & (g549) & (!g569) & (!g680)));
	assign g817 = (((!g708) & (!g716) & (!g549) & (!g569) & (!g680) & (g733)) + ((!g708) & (!g716) & (g549) & (!g569) & (!g680) & (g733)) + ((!g708) & (!g716) & (g549) & (!g569) & (g680) & (g733)) + ((!g708) & (!g716) & (g549) & (g569) & (!g680) & (g733)) + ((!g708) & (g716) & (!g549) & (!g569) & (g680) & (g733)) + ((!g708) & (g716) & (!g549) & (g569) & (!g680) & (g733)) + ((!g708) & (g716) & (!g549) & (g569) & (g680) & (g733)) + ((!g708) & (g716) & (g549) & (g569) & (g680) & (g733)) + ((g708) & (!g716) & (!g549) & (!g569) & (g680) & (g733)) + ((g708) & (!g716) & (!g549) & (g569) & (!g680) & (g733)) + ((g708) & (!g716) & (!g549) & (g569) & (g680) & (g733)) + ((g708) & (!g716) & (g549) & (g569) & (g680) & (g733)) + ((g708) & (g716) & (!g549) & (!g569) & (!g680) & (g733)) + ((g708) & (g716) & (g549) & (!g569) & (!g680) & (g733)) + ((g708) & (g716) & (g549) & (!g569) & (g680) & (g733)) + ((g708) & (g716) & (g549) & (g569) & (!g680) & (g733)));
	assign g818 = (((!g549) & (!g569) & (!g680) & (g686) & (!g734) & (!g729)) + ((!g549) & (!g569) & (!g680) & (g686) & (g734) & (!g729)) + ((!g549) & (!g569) & (g680) & (!g686) & (g734) & (!g729)) + ((!g549) & (!g569) & (g680) & (!g686) & (g734) & (g729)) + ((!g549) & (!g569) & (g680) & (g686) & (!g734) & (!g729)) + ((!g549) & (!g569) & (g680) & (g686) & (g734) & (!g729)) + ((!g549) & (!g569) & (g680) & (g686) & (g734) & (g729)) + ((!g549) & (g569) & (!g680) & (!g686) & (g734) & (!g729)) + ((!g549) & (g569) & (!g680) & (!g686) & (g734) & (g729)) + ((!g549) & (g569) & (!g680) & (g686) & (!g734) & (!g729)) + ((!g549) & (g569) & (!g680) & (g686) & (g734) & (!g729)) + ((!g549) & (g569) & (!g680) & (g686) & (g734) & (g729)) + ((!g549) & (g569) & (g680) & (g686) & (!g734) & (!g729)) + ((!g549) & (g569) & (g680) & (g686) & (g734) & (!g729)) + ((g549) & (!g569) & (!g680) & (!g686) & (g734) & (!g729)) + ((g549) & (!g569) & (!g680) & (!g686) & (g734) & (g729)) + ((g549) & (!g569) & (!g680) & (g686) & (!g734) & (!g729)) + ((g549) & (!g569) & (!g680) & (g686) & (g734) & (!g729)) + ((g549) & (!g569) & (!g680) & (g686) & (g734) & (g729)) + ((g549) & (!g569) & (g680) & (g686) & (!g734) & (!g729)) + ((g549) & (!g569) & (g680) & (g686) & (g734) & (!g729)) + ((g549) & (g569) & (!g680) & (g686) & (!g734) & (!g729)) + ((g549) & (g569) & (!g680) & (g686) & (g734) & (!g729)) + ((g549) & (g569) & (g680) & (!g686) & (g734) & (!g729)) + ((g549) & (g569) & (g680) & (!g686) & (g734) & (g729)) + ((g549) & (g569) & (g680) & (g686) & (!g734) & (!g729)) + ((g549) & (g569) & (g680) & (g686) & (g734) & (!g729)) + ((g549) & (g569) & (g680) & (g686) & (g734) & (g729)));
	assign g819 = (((!g2) & (!g730) & (!g816) & (!g732) & (!g817) & (!g818)) + ((!g2) & (!g730) & (g816) & (!g732) & (!g817) & (!g818)) + ((!g2) & (!g730) & (g816) & (g732) & (!g817) & (!g818)) + ((!g2) & (g730) & (!g816) & (!g732) & (!g817) & (!g818)) + ((!g2) & (g730) & (!g816) & (g732) & (!g817) & (!g818)) + ((!g2) & (g730) & (g816) & (!g732) & (!g817) & (!g818)) + ((g2) & (!g730) & (!g816) & (!g732) & (!g817) & (g818)) + ((g2) & (!g730) & (!g816) & (!g732) & (g817) & (!g818)) + ((g2) & (!g730) & (!g816) & (!g732) & (g817) & (g818)) + ((g2) & (!g730) & (!g816) & (g732) & (!g817) & (!g818)) + ((g2) & (!g730) & (!g816) & (g732) & (!g817) & (g818)) + ((g2) & (!g730) & (!g816) & (g732) & (g817) & (!g818)) + ((g2) & (!g730) & (!g816) & (g732) & (g817) & (g818)) + ((g2) & (!g730) & (g816) & (!g732) & (!g817) & (g818)) + ((g2) & (!g730) & (g816) & (!g732) & (g817) & (!g818)) + ((g2) & (!g730) & (g816) & (!g732) & (g817) & (g818)) + ((g2) & (!g730) & (g816) & (g732) & (!g817) & (g818)) + ((g2) & (!g730) & (g816) & (g732) & (g817) & (!g818)) + ((g2) & (!g730) & (g816) & (g732) & (g817) & (g818)) + ((g2) & (g730) & (!g816) & (!g732) & (!g817) & (g818)) + ((g2) & (g730) & (!g816) & (!g732) & (g817) & (!g818)) + ((g2) & (g730) & (!g816) & (!g732) & (g817) & (g818)) + ((g2) & (g730) & (!g816) & (g732) & (!g817) & (g818)) + ((g2) & (g730) & (!g816) & (g732) & (g817) & (!g818)) + ((g2) & (g730) & (!g816) & (g732) & (g817) & (g818)) + ((g2) & (g730) & (g816) & (!g732) & (!g817) & (g818)) + ((g2) & (g730) & (g816) & (!g732) & (g817) & (!g818)) + ((g2) & (g730) & (g816) & (!g732) & (g817) & (g818)) + ((g2) & (g730) & (g816) & (g732) & (!g817) & (!g818)) + ((g2) & (g730) & (g816) & (g732) & (!g817) & (g818)) + ((g2) & (g730) & (g816) & (g732) & (g817) & (!g818)) + ((g2) & (g730) & (g816) & (g732) & (g817) & (g818)));
	assign g820 = (((!g770) & (!g773) & (sk[62]) & (g779)) + ((!g770) & (g773) & (!sk[62]) & (!g779)) + ((!g770) & (g773) & (!sk[62]) & (g779)) + ((!g770) & (g773) & (sk[62]) & (!g779)) + ((g770) & (!g773) & (sk[62]) & (!g779)) + ((g770) & (g773) & (!sk[62]) & (!g779)) + ((g770) & (g773) & (!sk[62]) & (g779)) + ((g770) & (g773) & (sk[62]) & (g779)));
	assign g821 = (((!g789) & (!g790) & (!g793) & (!g815) & (!g819) & (!g820)) + ((!g789) & (!g790) & (!g793) & (!g815) & (g819) & (!g820)) + ((!g789) & (!g790) & (!g793) & (!g815) & (g819) & (g820)) + ((!g789) & (!g790) & (!g793) & (g815) & (g819) & (!g820)) + ((!g789) & (!g790) & (g793) & (!g815) & (!g819) & (!g820)) + ((!g789) & (!g790) & (g793) & (!g815) & (g819) & (!g820)) + ((!g789) & (!g790) & (g793) & (!g815) & (g819) & (g820)) + ((!g789) & (!g790) & (g793) & (g815) & (!g819) & (!g820)) + ((!g789) & (!g790) & (g793) & (g815) & (g819) & (!g820)) + ((!g789) & (!g790) & (g793) & (g815) & (g819) & (g820)) + ((!g789) & (g790) & (!g793) & (!g815) & (g819) & (!g820)) + ((!g789) & (g790) & (!g793) & (g815) & (g819) & (!g820)) + ((!g789) & (g790) & (g793) & (!g815) & (!g819) & (!g820)) + ((!g789) & (g790) & (g793) & (!g815) & (g819) & (!g820)) + ((!g789) & (g790) & (g793) & (!g815) & (g819) & (g820)) + ((!g789) & (g790) & (g793) & (g815) & (g819) & (!g820)) + ((g789) & (!g790) & (!g793) & (!g815) & (g819) & (!g820)) + ((g789) & (!g790) & (!g793) & (g815) & (g819) & (!g820)) + ((g789) & (!g790) & (g793) & (!g815) & (!g819) & (!g820)) + ((g789) & (!g790) & (g793) & (!g815) & (g819) & (!g820)) + ((g789) & (!g790) & (g793) & (!g815) & (g819) & (g820)) + ((g789) & (!g790) & (g793) & (g815) & (g819) & (!g820)) + ((g789) & (g790) & (!g793) & (!g815) & (!g819) & (!g820)) + ((g789) & (g790) & (!g793) & (!g815) & (g819) & (!g820)) + ((g789) & (g790) & (!g793) & (!g815) & (g819) & (g820)) + ((g789) & (g790) & (!g793) & (g815) & (g819) & (!g820)) + ((g789) & (g790) & (g793) & (!g815) & (!g819) & (!g820)) + ((g789) & (g790) & (g793) & (!g815) & (g819) & (!g820)) + ((g789) & (g790) & (g793) & (!g815) & (g819) & (g820)) + ((g789) & (g790) & (g793) & (g815) & (!g819) & (!g820)) + ((g789) & (g790) & (g793) & (g815) & (g819) & (!g820)) + ((g789) & (g790) & (g793) & (g815) & (g819) & (g820)));
	assign g822 = (((!g696) & (!g697) & (!g316) & (!g322) & (sk[64]) & (!g548)) + ((!g696) & (!g697) & (!g316) & (!g322) & (sk[64]) & (g548)) + ((!g696) & (!g697) & (!g316) & (g322) & (!sk[64]) & (!g548)) + ((!g696) & (!g697) & (!g316) & (g322) & (!sk[64]) & (g548)) + ((!g696) & (!g697) & (!g316) & (g322) & (sk[64]) & (g548)) + ((!g696) & (!g697) & (g316) & (!g322) & (!sk[64]) & (!g548)) + ((!g696) & (!g697) & (g316) & (!g322) & (!sk[64]) & (g548)) + ((!g696) & (!g697) & (g316) & (!g322) & (sk[64]) & (g548)) + ((!g696) & (!g697) & (g316) & (g322) & (!sk[64]) & (!g548)) + ((!g696) & (!g697) & (g316) & (g322) & (!sk[64]) & (g548)) + ((!g696) & (g697) & (!g316) & (!g322) & (!sk[64]) & (!g548)) + ((!g696) & (g697) & (!g316) & (!g322) & (!sk[64]) & (g548)) + ((!g696) & (g697) & (!g316) & (!g322) & (sk[64]) & (!g548)) + ((!g696) & (g697) & (!g316) & (!g322) & (sk[64]) & (g548)) + ((!g696) & (g697) & (!g316) & (g322) & (!sk[64]) & (!g548)) + ((!g696) & (g697) & (!g316) & (g322) & (!sk[64]) & (g548)) + ((!g696) & (g697) & (!g316) & (g322) & (sk[64]) & (!g548)) + ((!g696) & (g697) & (!g316) & (g322) & (sk[64]) & (g548)) + ((!g696) & (g697) & (g316) & (!g322) & (!sk[64]) & (!g548)) + ((!g696) & (g697) & (g316) & (!g322) & (!sk[64]) & (g548)) + ((!g696) & (g697) & (g316) & (!g322) & (sk[64]) & (!g548)) + ((!g696) & (g697) & (g316) & (!g322) & (sk[64]) & (g548)) + ((!g696) & (g697) & (g316) & (g322) & (!sk[64]) & (!g548)) + ((!g696) & (g697) & (g316) & (g322) & (!sk[64]) & (g548)) + ((!g696) & (g697) & (g316) & (g322) & (sk[64]) & (!g548)) + ((!g696) & (g697) & (g316) & (g322) & (sk[64]) & (g548)) + ((g696) & (!g697) & (!g316) & (g322) & (!sk[64]) & (!g548)) + ((g696) & (!g697) & (!g316) & (g322) & (!sk[64]) & (g548)) + ((g696) & (!g697) & (g316) & (!g322) & (!sk[64]) & (!g548)) + ((g696) & (!g697) & (g316) & (!g322) & (!sk[64]) & (g548)) + ((g696) & (!g697) & (g316) & (g322) & (!sk[64]) & (!g548)) + ((g696) & (!g697) & (g316) & (g322) & (!sk[64]) & (g548)) + ((g696) & (g697) & (!g316) & (!g322) & (!sk[64]) & (!g548)) + ((g696) & (g697) & (!g316) & (!g322) & (!sk[64]) & (g548)) + ((g696) & (g697) & (!g316) & (!g322) & (sk[64]) & (!g548)) + ((g696) & (g697) & (!g316) & (!g322) & (sk[64]) & (g548)) + ((g696) & (g697) & (!g316) & (g322) & (!sk[64]) & (!g548)) + ((g696) & (g697) & (!g316) & (g322) & (!sk[64]) & (g548)) + ((g696) & (g697) & (!g316) & (g322) & (sk[64]) & (g548)) + ((g696) & (g697) & (g316) & (!g322) & (!sk[64]) & (!g548)) + ((g696) & (g697) & (g316) & (!g322) & (!sk[64]) & (g548)) + ((g696) & (g697) & (g316) & (!g322) & (sk[64]) & (g548)) + ((g696) & (g697) & (g316) & (g322) & (!sk[64]) & (!g548)) + ((g696) & (g697) & (g316) & (g322) & (!sk[64]) & (g548)));
	assign g823 = (((!g209) & (!g215) & (!g216) & (!sk[65]) & (g219)) + ((!g209) & (!g215) & (g216) & (!sk[65]) & (g219)) + ((!g209) & (g215) & (!g216) & (!sk[65]) & (g219)) + ((!g209) & (g215) & (g216) & (!sk[65]) & (g219)) + ((g209) & (!g215) & (!g216) & (!sk[65]) & (!g219)) + ((g209) & (!g215) & (!g216) & (!sk[65]) & (g219)) + ((g209) & (!g215) & (!g216) & (sk[65]) & (g219)) + ((g209) & (!g215) & (g216) & (!sk[65]) & (!g219)) + ((g209) & (!g215) & (g216) & (!sk[65]) & (g219)) + ((g209) & (g215) & (!g216) & (!sk[65]) & (!g219)) + ((g209) & (g215) & (!g216) & (!sk[65]) & (g219)) + ((g209) & (g215) & (!g216) & (sk[65]) & (!g219)) + ((g209) & (g215) & (!g216) & (sk[65]) & (g219)) + ((g209) & (g215) & (g216) & (!sk[65]) & (!g219)) + ((g209) & (g215) & (g216) & (!sk[65]) & (g219)) + ((g209) & (g215) & (g216) & (sk[65]) & (!g219)) + ((g209) & (g215) & (g216) & (sk[65]) & (g219)));
	assign g824 = (((!g69) & (!g252) & (!g253) & (!g823) & (!g692) & (!g693)) + ((!g69) & (!g252) & (!g253) & (g823) & (!g692) & (g693)) + ((!g69) & (!g252) & (!g253) & (g823) & (g692) & (!g693)) + ((!g69) & (!g252) & (!g253) & (g823) & (g692) & (g693)) + ((!g69) & (!g252) & (g253) & (!g823) & (g692) & (g693)) + ((!g69) & (!g252) & (g253) & (g823) & (!g692) & (!g693)) + ((!g69) & (!g252) & (g253) & (g823) & (!g692) & (g693)) + ((!g69) & (!g252) & (g253) & (g823) & (g692) & (!g693)) + ((!g69) & (g252) & (!g253) & (!g823) & (!g692) & (g693)) + ((!g69) & (g252) & (!g253) & (!g823) & (g692) & (!g693)) + ((!g69) & (g252) & (!g253) & (!g823) & (g692) & (g693)) + ((!g69) & (g252) & (!g253) & (g823) & (!g692) & (!g693)) + ((!g69) & (g252) & (g253) & (!g823) & (!g692) & (!g693)) + ((!g69) & (g252) & (g253) & (!g823) & (!g692) & (g693)) + ((!g69) & (g252) & (g253) & (!g823) & (g692) & (!g693)) + ((!g69) & (g252) & (g253) & (g823) & (g692) & (g693)) + ((g69) & (!g252) & (!g253) & (!g823) & (!g692) & (!g693)) + ((g69) & (!g252) & (!g253) & (g823) & (!g692) & (!g693)) + ((g69) & (!g252) & (g253) & (!g823) & (!g692) & (!g693)) + ((g69) & (!g252) & (g253) & (g823) & (!g692) & (!g693)) + ((g69) & (g252) & (!g253) & (!g823) & (!g692) & (!g693)) + ((g69) & (g252) & (!g253) & (g823) & (!g692) & (!g693)) + ((g69) & (g252) & (g253) & (!g823) & (!g692) & (!g693)) + ((g69) & (g252) & (g253) & (g823) & (!g692) & (!g693)));
	assign g825 = (((!g691) & (!g694) & (!g822) & (!sk[67]) & (g824)) + ((!g691) & (!g694) & (!g822) & (sk[67]) & (!g824)) + ((!g691) & (!g694) & (g822) & (!sk[67]) & (g824)) + ((!g691) & (!g694) & (g822) & (sk[67]) & (g824)) + ((!g691) & (g694) & (!g822) & (!sk[67]) & (g824)) + ((!g691) & (g694) & (!g822) & (sk[67]) & (g824)) + ((!g691) & (g694) & (g822) & (!sk[67]) & (g824)) + ((!g691) & (g694) & (g822) & (sk[67]) & (g824)) + ((g691) & (!g694) & (!g822) & (!sk[67]) & (!g824)) + ((g691) & (!g694) & (!g822) & (!sk[67]) & (g824)) + ((g691) & (!g694) & (!g822) & (sk[67]) & (!g824)) + ((g691) & (!g694) & (g822) & (!sk[67]) & (!g824)) + ((g691) & (!g694) & (g822) & (!sk[67]) & (g824)) + ((g691) & (!g694) & (g822) & (sk[67]) & (!g824)) + ((g691) & (g694) & (!g822) & (!sk[67]) & (!g824)) + ((g691) & (g694) & (!g822) & (!sk[67]) & (g824)) + ((g691) & (g694) & (!g822) & (sk[67]) & (!g824)) + ((g691) & (g694) & (g822) & (!sk[67]) & (!g824)) + ((g691) & (g694) & (g822) & (!sk[67]) & (g824)) + ((g691) & (g694) & (g822) & (sk[67]) & (g824)));
	assign g826 = (((!g9) & (!g16) & (!g25) & (!g275) & (!g194) & (!g169)) + ((!g9) & (!g16) & (!g25) & (!g275) & (!g194) & (g169)) + ((!g9) & (!g16) & (g25) & (!g275) & (!g194) & (!g169)) + ((!g9) & (!g16) & (g25) & (!g275) & (!g194) & (g169)) + ((!g9) & (g16) & (!g25) & (!g275) & (!g194) & (!g169)) + ((!g9) & (g16) & (!g25) & (!g275) & (!g194) & (g169)) + ((g9) & (!g16) & (!g25) & (!g275) & (!g194) & (!g169)) + ((g9) & (!g16) & (g25) & (!g275) & (!g194) & (!g169)) + ((g9) & (g16) & (!g25) & (!g275) & (!g194) & (!g169)));
	assign g827 = (((!sk[69]) & (!g9) & (g32) & (!g826)) + ((!sk[69]) & (!g9) & (g32) & (g826)) + ((!sk[69]) & (g9) & (g32) & (!g826)) + ((!sk[69]) & (g9) & (g32) & (g826)) + ((sk[69]) & (!g9) & (!g32) & (g826)) + ((sk[69]) & (!g9) & (g32) & (g826)) + ((sk[69]) & (g9) & (!g32) & (g826)));
	assign g828 = (((!g334) & (!g335) & (!sk[70]) & (!g336) & (g337)) + ((!g334) & (!g335) & (!sk[70]) & (g336) & (g337)) + ((!g334) & (g335) & (!sk[70]) & (!g336) & (g337)) + ((!g334) & (g335) & (!sk[70]) & (g336) & (g337)) + ((g334) & (!g335) & (!sk[70]) & (!g336) & (!g337)) + ((g334) & (!g335) & (!sk[70]) & (!g336) & (g337)) + ((g334) & (!g335) & (!sk[70]) & (g336) & (!g337)) + ((g334) & (!g335) & (!sk[70]) & (g336) & (g337)) + ((g334) & (g335) & (!sk[70]) & (!g336) & (!g337)) + ((g334) & (g335) & (!sk[70]) & (!g336) & (g337)) + ((g334) & (g335) & (!sk[70]) & (g336) & (!g337)) + ((g334) & (g335) & (!sk[70]) & (g336) & (g337)) + ((g334) & (g335) & (sk[70]) & (g336) & (g337)));
	assign g829 = (((!g563) & (!g74) & (!g185) & (!g288) & (sk[71]) & (g828)) + ((!g563) & (!g74) & (!g185) & (g288) & (!sk[71]) & (!g828)) + ((!g563) & (!g74) & (!g185) & (g288) & (!sk[71]) & (g828)) + ((!g563) & (!g74) & (g185) & (!g288) & (!sk[71]) & (!g828)) + ((!g563) & (!g74) & (g185) & (!g288) & (!sk[71]) & (g828)) + ((!g563) & (!g74) & (g185) & (g288) & (!sk[71]) & (!g828)) + ((!g563) & (!g74) & (g185) & (g288) & (!sk[71]) & (g828)) + ((!g563) & (g74) & (!g185) & (!g288) & (!sk[71]) & (!g828)) + ((!g563) & (g74) & (!g185) & (!g288) & (!sk[71]) & (g828)) + ((!g563) & (g74) & (!g185) & (g288) & (!sk[71]) & (!g828)) + ((!g563) & (g74) & (!g185) & (g288) & (!sk[71]) & (g828)) + ((!g563) & (g74) & (g185) & (!g288) & (!sk[71]) & (!g828)) + ((!g563) & (g74) & (g185) & (!g288) & (!sk[71]) & (g828)) + ((!g563) & (g74) & (g185) & (g288) & (!sk[71]) & (!g828)) + ((!g563) & (g74) & (g185) & (g288) & (!sk[71]) & (g828)) + ((g563) & (!g74) & (!g185) & (g288) & (!sk[71]) & (!g828)) + ((g563) & (!g74) & (!g185) & (g288) & (!sk[71]) & (g828)) + ((g563) & (!g74) & (g185) & (!g288) & (!sk[71]) & (!g828)) + ((g563) & (!g74) & (g185) & (!g288) & (!sk[71]) & (g828)) + ((g563) & (!g74) & (g185) & (g288) & (!sk[71]) & (!g828)) + ((g563) & (!g74) & (g185) & (g288) & (!sk[71]) & (g828)) + ((g563) & (g74) & (!g185) & (!g288) & (!sk[71]) & (!g828)) + ((g563) & (g74) & (!g185) & (!g288) & (!sk[71]) & (g828)) + ((g563) & (g74) & (!g185) & (g288) & (!sk[71]) & (!g828)) + ((g563) & (g74) & (!g185) & (g288) & (!sk[71]) & (g828)) + ((g563) & (g74) & (g185) & (!g288) & (!sk[71]) & (!g828)) + ((g563) & (g74) & (g185) & (!g288) & (!sk[71]) & (g828)) + ((g563) & (g74) & (g185) & (g288) & (!sk[71]) & (!g828)) + ((g563) & (g74) & (g185) & (g288) & (!sk[71]) & (g828)));
	assign g830 = (((!g17) & (!g49) & (!g58) & (!g46) & (!g104) & (g553)) + ((!g17) & (!g49) & (!g58) & (!g46) & (g104) & (g553)) + ((!g17) & (!g49) & (!g58) & (g46) & (!g104) & (g553)) + ((!g17) & (!g49) & (!g58) & (g46) & (g104) & (g553)) + ((!g17) & (!g49) & (g58) & (!g46) & (!g104) & (g553)) + ((!g17) & (!g49) & (g58) & (g46) & (!g104) & (g553)) + ((!g17) & (g49) & (!g58) & (!g46) & (!g104) & (g553)) + ((!g17) & (g49) & (g58) & (!g46) & (!g104) & (g553)) + ((g17) & (!g49) & (!g58) & (!g46) & (!g104) & (g553)) + ((g17) & (!g49) & (!g58) & (!g46) & (g104) & (g553)) + ((g17) & (!g49) & (g58) & (!g46) & (!g104) & (g553)) + ((g17) & (g49) & (!g58) & (!g46) & (!g104) & (g553)) + ((g17) & (g49) & (g58) & (!g46) & (!g104) & (g553)));
	assign g831 = (((!g70) & (!g40) & (!g25) & (!g80) & (g659) & (g830)) + ((!g70) & (!g40) & (g25) & (!g80) & (g659) & (g830)) + ((!g70) & (g40) & (!g25) & (!g80) & (g659) & (g830)) + ((!g70) & (g40) & (g25) & (!g80) & (g659) & (g830)) + ((g70) & (!g40) & (!g25) & (!g80) & (g659) & (g830)));
	assign g832 = (((!g616) & (!g649) & (!g827) & (!sk[74]) & (g829) & (!g831)) + ((!g616) & (!g649) & (!g827) & (!sk[74]) & (g829) & (g831)) + ((!g616) & (!g649) & (g827) & (!sk[74]) & (!g829) & (!g831)) + ((!g616) & (!g649) & (g827) & (!sk[74]) & (!g829) & (g831)) + ((!g616) & (!g649) & (g827) & (!sk[74]) & (g829) & (!g831)) + ((!g616) & (!g649) & (g827) & (!sk[74]) & (g829) & (g831)) + ((!g616) & (g649) & (!g827) & (!sk[74]) & (!g829) & (!g831)) + ((!g616) & (g649) & (!g827) & (!sk[74]) & (!g829) & (g831)) + ((!g616) & (g649) & (!g827) & (!sk[74]) & (g829) & (!g831)) + ((!g616) & (g649) & (!g827) & (!sk[74]) & (g829) & (g831)) + ((!g616) & (g649) & (g827) & (!sk[74]) & (!g829) & (!g831)) + ((!g616) & (g649) & (g827) & (!sk[74]) & (!g829) & (g831)) + ((!g616) & (g649) & (g827) & (!sk[74]) & (g829) & (!g831)) + ((!g616) & (g649) & (g827) & (!sk[74]) & (g829) & (g831)) + ((g616) & (!g649) & (!g827) & (!sk[74]) & (g829) & (!g831)) + ((g616) & (!g649) & (!g827) & (!sk[74]) & (g829) & (g831)) + ((g616) & (!g649) & (g827) & (!sk[74]) & (!g829) & (!g831)) + ((g616) & (!g649) & (g827) & (!sk[74]) & (!g829) & (g831)) + ((g616) & (!g649) & (g827) & (!sk[74]) & (g829) & (!g831)) + ((g616) & (!g649) & (g827) & (!sk[74]) & (g829) & (g831)) + ((g616) & (g649) & (!g827) & (!sk[74]) & (!g829) & (!g831)) + ((g616) & (g649) & (!g827) & (!sk[74]) & (!g829) & (g831)) + ((g616) & (g649) & (!g827) & (!sk[74]) & (g829) & (!g831)) + ((g616) & (g649) & (!g827) & (!sk[74]) & (g829) & (g831)) + ((g616) & (g649) & (g827) & (!sk[74]) & (!g829) & (!g831)) + ((g616) & (g649) & (g827) & (!sk[74]) & (!g829) & (g831)) + ((g616) & (g649) & (g827) & (!sk[74]) & (g829) & (!g831)) + ((g616) & (g649) & (g827) & (!sk[74]) & (g829) & (g831)) + ((g616) & (g649) & (g827) & (sk[74]) & (g829) & (g831)));
	assign g833 = (((!g698) & (!g706) & (!g717) & (g733) & (!g825) & (!g832)) + ((!g698) & (!g706) & (!g717) & (g733) & (g825) & (g832)) + ((!g698) & (!g706) & (g717) & (g733) & (!g825) & (!g832)) + ((!g698) & (!g706) & (g717) & (g733) & (g825) & (g832)) + ((!g698) & (g706) & (!g717) & (g733) & (!g825) & (!g832)) + ((!g698) & (g706) & (!g717) & (g733) & (g825) & (g832)) + ((!g698) & (g706) & (g717) & (g733) & (!g825) & (g832)) + ((!g698) & (g706) & (g717) & (g733) & (g825) & (!g832)) + ((g698) & (!g706) & (!g717) & (g733) & (!g825) & (!g832)) + ((g698) & (!g706) & (!g717) & (g733) & (g825) & (g832)) + ((g698) & (!g706) & (g717) & (g733) & (!g825) & (g832)) + ((g698) & (!g706) & (g717) & (g733) & (g825) & (!g832)) + ((g698) & (g706) & (!g717) & (g733) & (!g825) & (g832)) + ((g698) & (g706) & (!g717) & (g733) & (g825) & (!g832)) + ((g698) & (g706) & (g717) & (g733) & (!g825) & (g832)) + ((g698) & (g706) & (g717) & (g733) & (g825) & (!g832)));
	assign g834 = (((!sk[76]) & (!g707) & (!g717) & (!g681) & (g718) & (!g730)) + ((!sk[76]) & (!g707) & (!g717) & (!g681) & (g718) & (g730)) + ((!sk[76]) & (!g707) & (!g717) & (g681) & (!g718) & (!g730)) + ((!sk[76]) & (!g707) & (!g717) & (g681) & (!g718) & (g730)) + ((!sk[76]) & (!g707) & (!g717) & (g681) & (g718) & (!g730)) + ((!sk[76]) & (!g707) & (!g717) & (g681) & (g718) & (g730)) + ((!sk[76]) & (!g707) & (g717) & (!g681) & (!g718) & (!g730)) + ((!sk[76]) & (!g707) & (g717) & (!g681) & (!g718) & (g730)) + ((!sk[76]) & (!g707) & (g717) & (!g681) & (g718) & (!g730)) + ((!sk[76]) & (!g707) & (g717) & (!g681) & (g718) & (g730)) + ((!sk[76]) & (!g707) & (g717) & (g681) & (!g718) & (!g730)) + ((!sk[76]) & (!g707) & (g717) & (g681) & (!g718) & (g730)) + ((!sk[76]) & (!g707) & (g717) & (g681) & (g718) & (!g730)) + ((!sk[76]) & (!g707) & (g717) & (g681) & (g718) & (g730)) + ((!sk[76]) & (g707) & (!g717) & (!g681) & (g718) & (!g730)) + ((!sk[76]) & (g707) & (!g717) & (!g681) & (g718) & (g730)) + ((!sk[76]) & (g707) & (!g717) & (g681) & (!g718) & (!g730)) + ((!sk[76]) & (g707) & (!g717) & (g681) & (!g718) & (g730)) + ((!sk[76]) & (g707) & (!g717) & (g681) & (g718) & (!g730)) + ((!sk[76]) & (g707) & (!g717) & (g681) & (g718) & (g730)) + ((!sk[76]) & (g707) & (g717) & (!g681) & (!g718) & (!g730)) + ((!sk[76]) & (g707) & (g717) & (!g681) & (!g718) & (g730)) + ((!sk[76]) & (g707) & (g717) & (!g681) & (g718) & (!g730)) + ((!sk[76]) & (g707) & (g717) & (!g681) & (g718) & (g730)) + ((!sk[76]) & (g707) & (g717) & (g681) & (!g718) & (!g730)) + ((!sk[76]) & (g707) & (g717) & (g681) & (!g718) & (g730)) + ((!sk[76]) & (g707) & (g717) & (g681) & (g718) & (!g730)) + ((!sk[76]) & (g707) & (g717) & (g681) & (g718) & (g730)) + ((sk[76]) & (!g707) & (!g717) & (!g681) & (g718) & (!g730)) + ((sk[76]) & (!g707) & (!g717) & (!g681) & (g718) & (g730)) + ((sk[76]) & (!g707) & (!g717) & (g681) & (g718) & (g730)) + ((sk[76]) & (!g707) & (g717) & (!g681) & (!g718) & (g730)) + ((sk[76]) & (!g707) & (g717) & (!g681) & (g718) & (!g730)) + ((sk[76]) & (!g707) & (g717) & (!g681) & (g718) & (g730)) + ((sk[76]) & (!g707) & (g717) & (g681) & (g718) & (!g730)) + ((sk[76]) & (!g707) & (g717) & (g681) & (g718) & (g730)) + ((sk[76]) & (g707) & (!g717) & (!g681) & (!g718) & (g730)) + ((sk[76]) & (g707) & (!g717) & (!g681) & (g718) & (!g730)) + ((sk[76]) & (g707) & (!g717) & (!g681) & (g718) & (g730)) + ((sk[76]) & (g707) & (!g717) & (g681) & (g718) & (!g730)) + ((sk[76]) & (g707) & (!g717) & (g681) & (g718) & (g730)) + ((sk[76]) & (g707) & (g717) & (!g681) & (g718) & (!g730)) + ((sk[76]) & (g707) & (g717) & (!g681) & (g718) & (g730)) + ((sk[76]) & (g707) & (g717) & (g681) & (g718) & (g730)));
	assign g835 = (((!g698) & (!sk[77]) & (!g706) & (!g717) & (g825) & (!g832)) + ((!g698) & (!sk[77]) & (!g706) & (!g717) & (g825) & (g832)) + ((!g698) & (!sk[77]) & (!g706) & (g717) & (!g825) & (!g832)) + ((!g698) & (!sk[77]) & (!g706) & (g717) & (!g825) & (g832)) + ((!g698) & (!sk[77]) & (!g706) & (g717) & (g825) & (!g832)) + ((!g698) & (!sk[77]) & (!g706) & (g717) & (g825) & (g832)) + ((!g698) & (!sk[77]) & (g706) & (!g717) & (!g825) & (!g832)) + ((!g698) & (!sk[77]) & (g706) & (!g717) & (!g825) & (g832)) + ((!g698) & (!sk[77]) & (g706) & (!g717) & (g825) & (!g832)) + ((!g698) & (!sk[77]) & (g706) & (!g717) & (g825) & (g832)) + ((!g698) & (!sk[77]) & (g706) & (g717) & (!g825) & (!g832)) + ((!g698) & (!sk[77]) & (g706) & (g717) & (!g825) & (g832)) + ((!g698) & (!sk[77]) & (g706) & (g717) & (g825) & (!g832)) + ((!g698) & (!sk[77]) & (g706) & (g717) & (g825) & (g832)) + ((!g698) & (sk[77]) & (!g706) & (!g717) & (!g825) & (!g832)) + ((!g698) & (sk[77]) & (!g706) & (!g717) & (g825) & (g832)) + ((!g698) & (sk[77]) & (!g706) & (g717) & (!g825) & (g832)) + ((!g698) & (sk[77]) & (!g706) & (g717) & (g825) & (!g832)) + ((!g698) & (sk[77]) & (g706) & (!g717) & (!g825) & (g832)) + ((!g698) & (sk[77]) & (g706) & (!g717) & (g825) & (!g832)) + ((!g698) & (sk[77]) & (g706) & (g717) & (!g825) & (g832)) + ((!g698) & (sk[77]) & (g706) & (g717) & (g825) & (!g832)) + ((g698) & (!sk[77]) & (!g706) & (!g717) & (g825) & (!g832)) + ((g698) & (!sk[77]) & (!g706) & (!g717) & (g825) & (g832)) + ((g698) & (!sk[77]) & (!g706) & (g717) & (!g825) & (!g832)) + ((g698) & (!sk[77]) & (!g706) & (g717) & (!g825) & (g832)) + ((g698) & (!sk[77]) & (!g706) & (g717) & (g825) & (!g832)) + ((g698) & (!sk[77]) & (!g706) & (g717) & (g825) & (g832)) + ((g698) & (!sk[77]) & (g706) & (!g717) & (!g825) & (!g832)) + ((g698) & (!sk[77]) & (g706) & (!g717) & (!g825) & (g832)) + ((g698) & (!sk[77]) & (g706) & (!g717) & (g825) & (!g832)) + ((g698) & (!sk[77]) & (g706) & (!g717) & (g825) & (g832)) + ((g698) & (!sk[77]) & (g706) & (g717) & (!g825) & (!g832)) + ((g698) & (!sk[77]) & (g706) & (g717) & (!g825) & (g832)) + ((g698) & (!sk[77]) & (g706) & (g717) & (g825) & (!g832)) + ((g698) & (!sk[77]) & (g706) & (g717) & (g825) & (g832)) + ((g698) & (sk[77]) & (!g706) & (!g717) & (!g825) & (g832)) + ((g698) & (sk[77]) & (!g706) & (!g717) & (g825) & (!g832)) + ((g698) & (sk[77]) & (!g706) & (g717) & (!g825) & (g832)) + ((g698) & (sk[77]) & (!g706) & (g717) & (g825) & (!g832)) + ((g698) & (sk[77]) & (g706) & (!g717) & (!g825) & (g832)) + ((g698) & (sk[77]) & (g706) & (!g717) & (g825) & (!g832)) + ((g698) & (sk[77]) & (g706) & (g717) & (!g825) & (!g832)) + ((g698) & (sk[77]) & (g706) & (g717) & (g825) & (g832)));
	assign g836 = (((!g707) & (!g717) & (!sk[78]) & (!g686) & (g734) & (!g718)) + ((!g707) & (!g717) & (!sk[78]) & (!g686) & (g734) & (g718)) + ((!g707) & (!g717) & (!sk[78]) & (g686) & (!g734) & (!g718)) + ((!g707) & (!g717) & (!sk[78]) & (g686) & (!g734) & (g718)) + ((!g707) & (!g717) & (!sk[78]) & (g686) & (g734) & (!g718)) + ((!g707) & (!g717) & (!sk[78]) & (g686) & (g734) & (g718)) + ((!g707) & (!g717) & (sk[78]) & (g686) & (!g734) & (g718)) + ((!g707) & (!g717) & (sk[78]) & (g686) & (g734) & (g718)) + ((!g707) & (g717) & (!sk[78]) & (!g686) & (!g734) & (!g718)) + ((!g707) & (g717) & (!sk[78]) & (!g686) & (!g734) & (g718)) + ((!g707) & (g717) & (!sk[78]) & (!g686) & (g734) & (!g718)) + ((!g707) & (g717) & (!sk[78]) & (!g686) & (g734) & (g718)) + ((!g707) & (g717) & (!sk[78]) & (g686) & (!g734) & (!g718)) + ((!g707) & (g717) & (!sk[78]) & (g686) & (!g734) & (g718)) + ((!g707) & (g717) & (!sk[78]) & (g686) & (g734) & (!g718)) + ((!g707) & (g717) & (!sk[78]) & (g686) & (g734) & (g718)) + ((!g707) & (g717) & (sk[78]) & (!g686) & (g734) & (!g718)) + ((!g707) & (g717) & (sk[78]) & (!g686) & (g734) & (g718)) + ((!g707) & (g717) & (sk[78]) & (g686) & (!g734) & (g718)) + ((!g707) & (g717) & (sk[78]) & (g686) & (g734) & (!g718)) + ((!g707) & (g717) & (sk[78]) & (g686) & (g734) & (g718)) + ((g707) & (!g717) & (!sk[78]) & (!g686) & (g734) & (!g718)) + ((g707) & (!g717) & (!sk[78]) & (!g686) & (g734) & (g718)) + ((g707) & (!g717) & (!sk[78]) & (g686) & (!g734) & (!g718)) + ((g707) & (!g717) & (!sk[78]) & (g686) & (!g734) & (g718)) + ((g707) & (!g717) & (!sk[78]) & (g686) & (g734) & (!g718)) + ((g707) & (!g717) & (!sk[78]) & (g686) & (g734) & (g718)) + ((g707) & (!g717) & (sk[78]) & (!g686) & (g734) & (!g718)) + ((g707) & (!g717) & (sk[78]) & (!g686) & (g734) & (g718)) + ((g707) & (!g717) & (sk[78]) & (g686) & (!g734) & (g718)) + ((g707) & (!g717) & (sk[78]) & (g686) & (g734) & (!g718)) + ((g707) & (!g717) & (sk[78]) & (g686) & (g734) & (g718)) + ((g707) & (g717) & (!sk[78]) & (!g686) & (!g734) & (!g718)) + ((g707) & (g717) & (!sk[78]) & (!g686) & (!g734) & (g718)) + ((g707) & (g717) & (!sk[78]) & (!g686) & (g734) & (!g718)) + ((g707) & (g717) & (!sk[78]) & (!g686) & (g734) & (g718)) + ((g707) & (g717) & (!sk[78]) & (g686) & (!g734) & (!g718)) + ((g707) & (g717) & (!sk[78]) & (g686) & (!g734) & (g718)) + ((g707) & (g717) & (!sk[78]) & (g686) & (g734) & (!g718)) + ((g707) & (g717) & (!sk[78]) & (g686) & (g734) & (g718)) + ((g707) & (g717) & (sk[78]) & (g686) & (!g734) & (g718)) + ((g707) & (g717) & (sk[78]) & (g686) & (g734) & (g718)));
	assign g837 = (((!g2) & (!g732) & (!g833) & (!g834) & (!g835) & (g836)) + ((!g2) & (!g732) & (!g833) & (!g834) & (g835) & (g836)) + ((!g2) & (!g732) & (!g833) & (g834) & (!g835) & (g836)) + ((!g2) & (!g732) & (!g833) & (g834) & (g835) & (g836)) + ((!g2) & (!g732) & (g833) & (!g834) & (!g835) & (!g836)) + ((!g2) & (!g732) & (g833) & (!g834) & (!g835) & (g836)) + ((!g2) & (!g732) & (g833) & (!g834) & (g835) & (!g836)) + ((!g2) & (!g732) & (g833) & (!g834) & (g835) & (g836)) + ((!g2) & (!g732) & (g833) & (g834) & (!g835) & (!g836)) + ((!g2) & (!g732) & (g833) & (g834) & (!g835) & (g836)) + ((!g2) & (!g732) & (g833) & (g834) & (g835) & (!g836)) + ((!g2) & (!g732) & (g833) & (g834) & (g835) & (g836)) + ((!g2) & (g732) & (!g833) & (!g834) & (!g835) & (!g836)) + ((!g2) & (g732) & (!g833) & (!g834) & (!g835) & (g836)) + ((!g2) & (g732) & (!g833) & (!g834) & (g835) & (g836)) + ((!g2) & (g732) & (!g833) & (g834) & (!g835) & (g836)) + ((!g2) & (g732) & (!g833) & (g834) & (g835) & (!g836)) + ((!g2) & (g732) & (!g833) & (g834) & (g835) & (g836)) + ((!g2) & (g732) & (g833) & (!g834) & (!g835) & (!g836)) + ((!g2) & (g732) & (g833) & (!g834) & (!g835) & (g836)) + ((!g2) & (g732) & (g833) & (!g834) & (g835) & (!g836)) + ((!g2) & (g732) & (g833) & (!g834) & (g835) & (g836)) + ((!g2) & (g732) & (g833) & (g834) & (!g835) & (!g836)) + ((!g2) & (g732) & (g833) & (g834) & (!g835) & (g836)) + ((!g2) & (g732) & (g833) & (g834) & (g835) & (!g836)) + ((!g2) & (g732) & (g833) & (g834) & (g835) & (g836)) + ((g2) & (!g732) & (!g833) & (!g834) & (!g835) & (!g836)) + ((g2) & (!g732) & (!g833) & (!g834) & (g835) & (!g836)) + ((g2) & (!g732) & (!g833) & (g834) & (!g835) & (!g836)) + ((g2) & (!g732) & (!g833) & (g834) & (g835) & (!g836)) + ((g2) & (g732) & (!g833) & (!g834) & (g835) & (!g836)) + ((g2) & (g732) & (!g833) & (g834) & (!g835) & (!g836)));
	assign g838 = (((!g200) & (!g770) & (!g773) & (!g779) & (!g785) & (!g787)) + ((!g200) & (!g770) & (!g773) & (!g779) & (!g785) & (g787)) + ((!g200) & (!g770) & (!g773) & (!g779) & (g785) & (!g787)) + ((!g200) & (!g770) & (!g773) & (g779) & (!g785) & (!g787)) + ((!g200) & (!g770) & (g773) & (!g779) & (!g785) & (!g787)) + ((!g200) & (!g770) & (g773) & (g779) & (!g785) & (!g787)) + ((!g200) & (g770) & (!g773) & (!g779) & (!g785) & (!g787)) + ((!g200) & (g770) & (!g773) & (!g779) & (!g785) & (g787)) + ((!g200) & (g770) & (!g773) & (!g779) & (g785) & (!g787)) + ((!g200) & (g770) & (!g773) & (g779) & (!g785) & (!g787)) + ((!g200) & (g770) & (!g773) & (g779) & (!g785) & (g787)) + ((!g200) & (g770) & (!g773) & (g779) & (g785) & (!g787)) + ((!g200) & (g770) & (g773) & (!g779) & (!g785) & (!g787)) + ((!g200) & (g770) & (g773) & (!g779) & (!g785) & (g787)) + ((!g200) & (g770) & (g773) & (!g779) & (g785) & (!g787)) + ((!g200) & (g770) & (g773) & (g779) & (!g785) & (!g787)) + ((g200) & (!g770) & (!g773) & (!g779) & (!g785) & (!g787)) + ((g200) & (!g770) & (!g773) & (!g779) & (!g785) & (g787)) + ((g200) & (!g770) & (!g773) & (!g779) & (g785) & (g787)) + ((g200) & (!g770) & (!g773) & (g779) & (!g785) & (g787)) + ((g200) & (!g770) & (g773) & (!g779) & (!g785) & (g787)) + ((g200) & (!g770) & (g773) & (g779) & (!g785) & (g787)) + ((g200) & (g770) & (!g773) & (!g779) & (!g785) & (!g787)) + ((g200) & (g770) & (!g773) & (!g779) & (!g785) & (g787)) + ((g200) & (g770) & (!g773) & (!g779) & (g785) & (g787)) + ((g200) & (g770) & (!g773) & (g779) & (!g785) & (!g787)) + ((g200) & (g770) & (!g773) & (g779) & (!g785) & (g787)) + ((g200) & (g770) & (!g773) & (g779) & (g785) & (g787)) + ((g200) & (g770) & (g773) & (!g779) & (!g785) & (!g787)) + ((g200) & (g770) & (g773) & (!g779) & (!g785) & (g787)) + ((g200) & (g770) & (g773) & (!g779) & (g785) & (g787)) + ((g200) & (g770) & (g773) & (g779) & (!g785) & (g787)));
	assign g839 = (((!g781) & (!sk[81]) & (g783) & (!g784)) + ((!g781) & (!sk[81]) & (g783) & (g784)) + ((!g781) & (sk[81]) & (!g783) & (g784)) + ((g781) & (!sk[81]) & (g783) & (!g784)) + ((g781) & (!sk[81]) & (g783) & (g784)) + ((g781) & (sk[81]) & (!g783) & (!g784)) + ((g781) & (sk[81]) & (!g783) & (g784)) + ((g781) & (sk[81]) & (g783) & (g784)));
	assign g840 = (((!sk[82]) & (!g721) & (!g678) & (!g723) & (g762) & (!g765)) + ((!sk[82]) & (!g721) & (!g678) & (!g723) & (g762) & (g765)) + ((!sk[82]) & (!g721) & (!g678) & (g723) & (!g762) & (!g765)) + ((!sk[82]) & (!g721) & (!g678) & (g723) & (!g762) & (g765)) + ((!sk[82]) & (!g721) & (!g678) & (g723) & (g762) & (!g765)) + ((!sk[82]) & (!g721) & (!g678) & (g723) & (g762) & (g765)) + ((!sk[82]) & (!g721) & (g678) & (!g723) & (!g762) & (!g765)) + ((!sk[82]) & (!g721) & (g678) & (!g723) & (!g762) & (g765)) + ((!sk[82]) & (!g721) & (g678) & (!g723) & (g762) & (!g765)) + ((!sk[82]) & (!g721) & (g678) & (!g723) & (g762) & (g765)) + ((!sk[82]) & (!g721) & (g678) & (g723) & (!g762) & (!g765)) + ((!sk[82]) & (!g721) & (g678) & (g723) & (!g762) & (g765)) + ((!sk[82]) & (!g721) & (g678) & (g723) & (g762) & (!g765)) + ((!sk[82]) & (!g721) & (g678) & (g723) & (g762) & (g765)) + ((!sk[82]) & (g721) & (!g678) & (!g723) & (g762) & (!g765)) + ((!sk[82]) & (g721) & (!g678) & (!g723) & (g762) & (g765)) + ((!sk[82]) & (g721) & (!g678) & (g723) & (!g762) & (!g765)) + ((!sk[82]) & (g721) & (!g678) & (g723) & (!g762) & (g765)) + ((!sk[82]) & (g721) & (!g678) & (g723) & (g762) & (!g765)) + ((!sk[82]) & (g721) & (!g678) & (g723) & (g762) & (g765)) + ((!sk[82]) & (g721) & (g678) & (!g723) & (!g762) & (!g765)) + ((!sk[82]) & (g721) & (g678) & (!g723) & (!g762) & (g765)) + ((!sk[82]) & (g721) & (g678) & (!g723) & (g762) & (!g765)) + ((!sk[82]) & (g721) & (g678) & (!g723) & (g762) & (g765)) + ((!sk[82]) & (g721) & (g678) & (g723) & (!g762) & (!g765)) + ((!sk[82]) & (g721) & (g678) & (g723) & (!g762) & (g765)) + ((!sk[82]) & (g721) & (g678) & (g723) & (g762) & (!g765)) + ((!sk[82]) & (g721) & (g678) & (g723) & (g762) & (g765)) + ((sk[82]) & (!g721) & (!g678) & (!g723) & (!g762) & (g765)) + ((sk[82]) & (!g721) & (!g678) & (!g723) & (g762) & (!g765)) + ((sk[82]) & (!g721) & (!g678) & (!g723) & (g762) & (g765)) + ((sk[82]) & (!g721) & (!g678) & (g723) & (g762) & (!g765)) + ((sk[82]) & (!g721) & (!g678) & (g723) & (g762) & (g765)) + ((sk[82]) & (!g721) & (g678) & (!g723) & (!g762) & (g765)) + ((sk[82]) & (!g721) & (g678) & (!g723) & (g762) & (g765)) + ((sk[82]) & (g721) & (!g678) & (!g723) & (!g762) & (g765)) + ((sk[82]) & (g721) & (!g678) & (!g723) & (g762) & (g765)) + ((sk[82]) & (g721) & (g678) & (!g723) & (!g762) & (g765)) + ((sk[82]) & (g721) & (g678) & (!g723) & (g762) & (!g765)) + ((sk[82]) & (g721) & (g678) & (!g723) & (g762) & (g765)) + ((sk[82]) & (g721) & (g678) & (g723) & (g762) & (!g765)) + ((sk[82]) & (g721) & (g678) & (g723) & (g762) & (g765)));
	assign g841 = (((!g720) & (!g722) & (!g727) & (!g764) & (!g759) & (!g840)) + ((!g720) & (!g722) & (!g727) & (g764) & (!g759) & (!g840)) + ((!g720) & (!g722) & (g727) & (!g764) & (!g759) & (!g840)) + ((!g720) & (!g722) & (g727) & (!g764) & (g759) & (!g840)) + ((!g720) & (!g722) & (g727) & (g764) & (!g759) & (!g840)) + ((!g720) & (!g722) & (g727) & (g764) & (g759) & (!g840)) + ((!g720) & (g722) & (!g727) & (!g764) & (!g759) & (!g840)) + ((!g720) & (g722) & (!g727) & (!g764) & (g759) & (!g840)) + ((!g720) & (g722) & (!g727) & (g764) & (!g759) & (!g840)) + ((!g720) & (g722) & (!g727) & (g764) & (g759) & (!g840)) + ((!g720) & (g722) & (g727) & (!g764) & (!g759) & (!g840)) + ((!g720) & (g722) & (g727) & (g764) & (!g759) & (!g840)) + ((g720) & (!g722) & (!g727) & (!g764) & (!g759) & (!g840)) + ((g720) & (!g722) & (!g727) & (!g764) & (g759) & (!g840)) + ((g720) & (!g722) & (g727) & (!g764) & (!g759) & (!g840)) + ((g720) & (g722) & (!g727) & (!g764) & (!g759) & (!g840)) + ((g720) & (g722) & (g727) & (!g764) & (!g759) & (!g840)) + ((g720) & (g722) & (g727) & (!g764) & (g759) & (!g840)));
	assign g842 = (((!sk[84]) & (g252) & (g253)) + ((sk[84]) & (!g252) & (g253)) + ((sk[84]) & (g252) & (!g253)));
	assign g843 = (((!sk[85]) & (g777) & (g842)) + ((sk[85]) & (g777) & (g842)));
	assign g844 = (((!g253) & (sk[86]) & (g303)) + ((g253) & (!sk[86]) & (g303)) + ((g253) & (sk[86]) & (!g303)));
	assign g845 = (((!sk[87]) & (g777) & (g844)) + ((sk[87]) & (!g777) & (g844)));
	assign g846 = (((g726) & (!sk[88]) & (g845)) + ((g726) & (sk[88]) & (g845)));
	assign g847 = (((g777) & (!sk[89]) & (g842)) + ((g777) & (sk[89]) & (!g842)));
	assign g848 = (((!g777) & (!sk[90]) & (g842) & (!g844)) + ((!g777) & (!sk[90]) & (g842) & (g844)) + ((!g777) & (sk[90]) & (g842) & (!g844)) + ((g777) & (!sk[90]) & (g842) & (!g844)) + ((g777) & (!sk[90]) & (g842) & (g844)));
	assign g849 = (((!g641) & (!g655) & (!g677) & (!g725) & (!g847) & (g848)) + ((!g641) & (!g655) & (!g677) & (!g725) & (g847) & (g848)) + ((!g641) & (!g655) & (g677) & (!g725) & (!g847) & (g848)) + ((!g641) & (!g655) & (g677) & (!g725) & (g847) & (!g848)) + ((!g641) & (!g655) & (g677) & (!g725) & (g847) & (g848)) + ((!g641) & (!g655) & (g677) & (g725) & (g847) & (!g848)) + ((!g641) & (!g655) & (g677) & (g725) & (g847) & (g848)) + ((!g641) & (g655) & (!g677) & (!g725) & (!g847) & (g848)) + ((!g641) & (g655) & (!g677) & (!g725) & (g847) & (!g848)) + ((!g641) & (g655) & (!g677) & (!g725) & (g847) & (g848)) + ((!g641) & (g655) & (!g677) & (g725) & (g847) & (!g848)) + ((!g641) & (g655) & (!g677) & (g725) & (g847) & (g848)) + ((!g641) & (g655) & (g677) & (!g725) & (!g847) & (g848)) + ((!g641) & (g655) & (g677) & (!g725) & (g847) & (g848)) + ((g641) & (!g655) & (!g677) & (!g725) & (!g847) & (g848)) + ((g641) & (!g655) & (!g677) & (!g725) & (g847) & (!g848)) + ((g641) & (!g655) & (!g677) & (!g725) & (g847) & (g848)) + ((g641) & (!g655) & (!g677) & (g725) & (g847) & (!g848)) + ((g641) & (!g655) & (!g677) & (g725) & (g847) & (g848)) + ((g641) & (!g655) & (g677) & (!g725) & (!g847) & (g848)) + ((g641) & (!g655) & (g677) & (!g725) & (g847) & (g848)) + ((g641) & (g655) & (!g677) & (!g725) & (!g847) & (g848)) + ((g641) & (g655) & (!g677) & (!g725) & (g847) & (g848)) + ((g641) & (g655) & (g677) & (!g725) & (!g847) & (g848)) + ((g641) & (g655) & (g677) & (!g725) & (g847) & (!g848)) + ((g641) & (g655) & (g677) & (!g725) & (g847) & (g848)) + ((g641) & (g655) & (g677) & (g725) & (g847) & (!g848)) + ((g641) & (g655) & (g677) & (g725) & (g847) & (g848)));
	assign g850 = (((!g202) & (g252) & (!g253) & (!g303) & (!g725) & (!g726)) + ((!g202) & (g252) & (!g253) & (!g303) & (!g725) & (g726)) + ((!g202) & (g252) & (!g253) & (!g303) & (g725) & (!g726)) + ((!g202) & (g252) & (!g253) & (!g303) & (g725) & (g726)) + ((!g202) & (g252) & (!g253) & (g303) & (g725) & (!g726)) + ((!g202) & (g252) & (g253) & (!g303) & (g725) & (!g726)) + ((!g202) & (g252) & (g253) & (!g303) & (g725) & (g726)) + ((!g202) & (g252) & (g253) & (g303) & (g725) & (!g726)) + ((g202) & (g252) & (!g253) & (!g303) & (g725) & (!g726)) + ((g202) & (g252) & (!g253) & (g303) & (g725) & (!g726)) + ((g202) & (g252) & (!g253) & (g303) & (g725) & (g726)) + ((g202) & (g252) & (g253) & (!g303) & (g725) & (!g726)) + ((g202) & (g252) & (g253) & (g303) & (!g725) & (!g726)) + ((g202) & (g252) & (g253) & (g303) & (!g725) & (g726)) + ((g202) & (g252) & (g253) & (g303) & (g725) & (!g726)) + ((g202) & (g252) & (g253) & (g303) & (g725) & (g726)));
	assign g851 = (((!g252) & (!g746) & (!g843) & (!g846) & (!g849) & (g850)) + ((!g252) & (!g746) & (!g843) & (!g846) & (g849) & (!g850)) + ((!g252) & (!g746) & (!g843) & (g846) & (!g849) & (!g850)) + ((!g252) & (!g746) & (!g843) & (g846) & (g849) & (!g850)) + ((!g252) & (!g746) & (g843) & (!g846) & (!g849) & (!g850)) + ((!g252) & (!g746) & (g843) & (!g846) & (g849) & (!g850)) + ((!g252) & (!g746) & (g843) & (g846) & (!g849) & (!g850)) + ((!g252) & (!g746) & (g843) & (g846) & (g849) & (!g850)) + ((!g252) & (g746) & (!g843) & (!g846) & (!g849) & (g850)) + ((!g252) & (g746) & (!g843) & (!g846) & (g849) & (!g850)) + ((!g252) & (g746) & (!g843) & (g846) & (!g849) & (!g850)) + ((!g252) & (g746) & (!g843) & (g846) & (g849) & (!g850)) + ((!g252) & (g746) & (g843) & (!g846) & (!g849) & (g850)) + ((!g252) & (g746) & (g843) & (!g846) & (g849) & (!g850)) + ((!g252) & (g746) & (g843) & (g846) & (!g849) & (!g850)) + ((!g252) & (g746) & (g843) & (g846) & (g849) & (!g850)) + ((g252) & (!g746) & (!g843) & (!g846) & (!g849) & (!g850)) + ((g252) & (!g746) & (!g843) & (!g846) & (g849) & (g850)) + ((g252) & (!g746) & (!g843) & (g846) & (!g849) & (g850)) + ((g252) & (!g746) & (!g843) & (g846) & (g849) & (g850)) + ((g252) & (!g746) & (g843) & (!g846) & (!g849) & (g850)) + ((g252) & (!g746) & (g843) & (!g846) & (g849) & (g850)) + ((g252) & (!g746) & (g843) & (g846) & (!g849) & (g850)) + ((g252) & (!g746) & (g843) & (g846) & (g849) & (g850)) + ((g252) & (g746) & (!g843) & (!g846) & (!g849) & (!g850)) + ((g252) & (g746) & (!g843) & (!g846) & (g849) & (g850)) + ((g252) & (g746) & (!g843) & (g846) & (!g849) & (g850)) + ((g252) & (g746) & (!g843) & (g846) & (g849) & (g850)) + ((g252) & (g746) & (g843) & (!g846) & (!g849) & (!g850)) + ((g252) & (g746) & (g843) & (!g846) & (g849) & (g850)) + ((g252) & (g746) & (g843) & (g846) & (!g849) & (g850)) + ((g252) & (g746) & (g843) & (g846) & (g849) & (g850)));
	assign g852 = (((!sk[94]) & (!g202) & (g841) & (!g851)) + ((!sk[94]) & (!g202) & (g841) & (g851)) + ((!sk[94]) & (g202) & (g841) & (!g851)) + ((!sk[94]) & (g202) & (g841) & (g851)) + ((sk[94]) & (!g202) & (!g841) & (!g851)) + ((sk[94]) & (!g202) & (g841) & (g851)) + ((sk[94]) & (g202) & (!g841) & (g851)) + ((sk[94]) & (g202) & (g841) & (!g851)));
	assign g853 = (((!g549) & (!g569) & (!g680) & (!g729) & (!g747) & (g744)) + ((!g549) & (!g569) & (!g680) & (!g729) & (g747) & (g744)) + ((!g549) & (!g569) & (g680) & (!g729) & (!g747) & (g744)) + ((!g549) & (!g569) & (g680) & (!g729) & (g747) & (!g744)) + ((!g549) & (!g569) & (g680) & (!g729) & (g747) & (g744)) + ((!g549) & (!g569) & (g680) & (g729) & (g747) & (!g744)) + ((!g549) & (!g569) & (g680) & (g729) & (g747) & (g744)) + ((!g549) & (g569) & (!g680) & (!g729) & (!g747) & (g744)) + ((!g549) & (g569) & (!g680) & (!g729) & (g747) & (!g744)) + ((!g549) & (g569) & (!g680) & (!g729) & (g747) & (g744)) + ((!g549) & (g569) & (!g680) & (g729) & (g747) & (!g744)) + ((!g549) & (g569) & (!g680) & (g729) & (g747) & (g744)) + ((!g549) & (g569) & (g680) & (!g729) & (!g747) & (g744)) + ((!g549) & (g569) & (g680) & (!g729) & (g747) & (g744)) + ((g549) & (!g569) & (!g680) & (!g729) & (!g747) & (g744)) + ((g549) & (!g569) & (!g680) & (!g729) & (g747) & (!g744)) + ((g549) & (!g569) & (!g680) & (!g729) & (g747) & (g744)) + ((g549) & (!g569) & (!g680) & (g729) & (g747) & (!g744)) + ((g549) & (!g569) & (!g680) & (g729) & (g747) & (g744)) + ((g549) & (!g569) & (g680) & (!g729) & (!g747) & (g744)) + ((g549) & (!g569) & (g680) & (!g729) & (g747) & (g744)) + ((g549) & (g569) & (!g680) & (!g729) & (!g747) & (g744)) + ((g549) & (g569) & (!g680) & (!g729) & (g747) & (g744)) + ((g549) & (g569) & (g680) & (!g729) & (!g747) & (g744)) + ((g549) & (g569) & (g680) & (!g729) & (g747) & (!g744)) + ((g549) & (g569) & (g680) & (!g729) & (g747) & (g744)) + ((g549) & (g569) & (g680) & (g729) & (g747) & (!g744)) + ((g549) & (g569) & (g680) & (g729) & (g747) & (g744)));
	assign g854 = (((!g200) & (!g719) & (!g742) & (!g748) & (!g791) & (!g853)) + ((!g200) & (!g719) & (!g742) & (!g748) & (g791) & (!g853)) + ((!g200) & (!g719) & (g742) & (!g748) & (!g791) & (!g853)) + ((!g200) & (g719) & (!g742) & (!g748) & (!g791) & (!g853)) + ((!g200) & (g719) & (!g742) & (!g748) & (g791) & (!g853)) + ((!g200) & (g719) & (!g742) & (g748) & (!g791) & (!g853)) + ((!g200) & (g719) & (!g742) & (g748) & (g791) & (!g853)) + ((!g200) & (g719) & (g742) & (!g748) & (!g791) & (!g853)) + ((!g200) & (g719) & (g742) & (g748) & (!g791) & (!g853)) + ((g200) & (!g719) & (!g742) & (!g748) & (!g791) & (g853)) + ((g200) & (!g719) & (!g742) & (!g748) & (g791) & (g853)) + ((g200) & (!g719) & (!g742) & (g748) & (!g791) & (!g853)) + ((g200) & (!g719) & (!g742) & (g748) & (!g791) & (g853)) + ((g200) & (!g719) & (!g742) & (g748) & (g791) & (!g853)) + ((g200) & (!g719) & (!g742) & (g748) & (g791) & (g853)) + ((g200) & (!g719) & (g742) & (!g748) & (!g791) & (g853)) + ((g200) & (!g719) & (g742) & (!g748) & (g791) & (!g853)) + ((g200) & (!g719) & (g742) & (!g748) & (g791) & (g853)) + ((g200) & (!g719) & (g742) & (g748) & (!g791) & (!g853)) + ((g200) & (!g719) & (g742) & (g748) & (!g791) & (g853)) + ((g200) & (!g719) & (g742) & (g748) & (g791) & (!g853)) + ((g200) & (!g719) & (g742) & (g748) & (g791) & (g853)) + ((g200) & (g719) & (!g742) & (!g748) & (!g791) & (g853)) + ((g200) & (g719) & (!g742) & (!g748) & (g791) & (g853)) + ((g200) & (g719) & (!g742) & (g748) & (!g791) & (g853)) + ((g200) & (g719) & (!g742) & (g748) & (g791) & (g853)) + ((g200) & (g719) & (g742) & (!g748) & (!g791) & (g853)) + ((g200) & (g719) & (g742) & (!g748) & (g791) & (!g853)) + ((g200) & (g719) & (g742) & (!g748) & (g791) & (g853)) + ((g200) & (g719) & (g742) & (g748) & (!g791) & (g853)) + ((g200) & (g719) & (g742) & (g748) & (g791) & (!g853)) + ((g200) & (g719) & (g742) & (g748) & (g791) & (g853)));
	assign g855 = (((!sk[97]) & (!g838) & (!g839) & (!g852) & (g854)) + ((!sk[97]) & (!g838) & (!g839) & (g852) & (g854)) + ((!sk[97]) & (!g838) & (g839) & (!g852) & (g854)) + ((!sk[97]) & (!g838) & (g839) & (g852) & (g854)) + ((!sk[97]) & (g838) & (!g839) & (!g852) & (!g854)) + ((!sk[97]) & (g838) & (!g839) & (!g852) & (g854)) + ((!sk[97]) & (g838) & (!g839) & (g852) & (!g854)) + ((!sk[97]) & (g838) & (!g839) & (g852) & (g854)) + ((!sk[97]) & (g838) & (g839) & (!g852) & (!g854)) + ((!sk[97]) & (g838) & (g839) & (!g852) & (g854)) + ((!sk[97]) & (g838) & (g839) & (g852) & (!g854)) + ((!sk[97]) & (g838) & (g839) & (g852) & (g854)) + ((sk[97]) & (!g838) & (!g839) & (!g852) & (g854)) + ((sk[97]) & (!g838) & (!g839) & (g852) & (!g854)) + ((sk[97]) & (!g838) & (g839) & (!g852) & (!g854)) + ((sk[97]) & (!g838) & (g839) & (g852) & (g854)) + ((sk[97]) & (g838) & (!g839) & (!g852) & (!g854)) + ((sk[97]) & (g838) & (!g839) & (g852) & (g854)) + ((sk[97]) & (g838) & (g839) & (!g852) & (g854)) + ((sk[97]) & (g838) & (g839) & (g852) & (!g854)));
	assign g856 = (((!g736) & (!g780) & (!g788) & (!g821) & (!g837) & (!g855)) + ((!g736) & (!g780) & (!g788) & (!g821) & (g837) & (g855)) + ((!g736) & (!g780) & (!g788) & (g821) & (!g837) & (!g855)) + ((!g736) & (!g780) & (!g788) & (g821) & (g837) & (g855)) + ((!g736) & (!g780) & (g788) & (!g821) & (!g837) & (!g855)) + ((!g736) & (!g780) & (g788) & (!g821) & (g837) & (g855)) + ((!g736) & (!g780) & (g788) & (g821) & (!g837) & (g855)) + ((!g736) & (!g780) & (g788) & (g821) & (g837) & (!g855)) + ((!g736) & (g780) & (!g788) & (!g821) & (!g837) & (!g855)) + ((!g736) & (g780) & (!g788) & (!g821) & (g837) & (g855)) + ((!g736) & (g780) & (!g788) & (g821) & (!g837) & (g855)) + ((!g736) & (g780) & (!g788) & (g821) & (g837) & (!g855)) + ((!g736) & (g780) & (g788) & (!g821) & (!g837) & (!g855)) + ((!g736) & (g780) & (g788) & (!g821) & (g837) & (g855)) + ((!g736) & (g780) & (g788) & (g821) & (!g837) & (!g855)) + ((!g736) & (g780) & (g788) & (g821) & (g837) & (g855)) + ((g736) & (!g780) & (!g788) & (!g821) & (!g837) & (!g855)) + ((g736) & (!g780) & (!g788) & (!g821) & (g837) & (g855)) + ((g736) & (!g780) & (!g788) & (g821) & (!g837) & (g855)) + ((g736) & (!g780) & (!g788) & (g821) & (g837) & (!g855)) + ((g736) & (!g780) & (g788) & (!g821) & (!g837) & (g855)) + ((g736) & (!g780) & (g788) & (!g821) & (g837) & (!g855)) + ((g736) & (!g780) & (g788) & (g821) & (!g837) & (g855)) + ((g736) & (!g780) & (g788) & (g821) & (g837) & (!g855)) + ((g736) & (g780) & (!g788) & (!g821) & (!g837) & (g855)) + ((g736) & (g780) & (!g788) & (!g821) & (g837) & (!g855)) + ((g736) & (g780) & (!g788) & (g821) & (!g837) & (g855)) + ((g736) & (g780) & (!g788) & (g821) & (g837) & (!g855)) + ((g736) & (g780) & (g788) & (!g821) & (!g837) & (!g855)) + ((g736) & (g780) & (g788) & (!g821) & (g837) & (g855)) + ((g736) & (g780) & (g788) & (g821) & (!g837) & (g855)) + ((g736) & (g780) & (g788) & (g821) & (g837) & (!g855)));
	assign g857 = (((!sk[99]) & (!g267) & (g186) & (!g424)) + ((!sk[99]) & (!g267) & (g186) & (g424)) + ((!sk[99]) & (g267) & (g186) & (!g424)) + ((!sk[99]) & (g267) & (g186) & (g424)) + ((sk[99]) & (!g267) & (g186) & (g424)));
	assign g858 = (((!g153) & (!sk[100]) & (!g104) & (!g32) & (g64)) + ((!g153) & (!sk[100]) & (!g104) & (g32) & (g64)) + ((!g153) & (!sk[100]) & (g104) & (!g32) & (g64)) + ((!g153) & (!sk[100]) & (g104) & (g32) & (g64)) + ((!g153) & (sk[100]) & (!g104) & (!g32) & (!g64)) + ((!g153) & (sk[100]) & (!g104) & (g32) & (!g64)) + ((!g153) & (sk[100]) & (g104) & (!g32) & (!g64)) + ((g153) & (!sk[100]) & (!g104) & (!g32) & (!g64)) + ((g153) & (!sk[100]) & (!g104) & (!g32) & (g64)) + ((g153) & (!sk[100]) & (!g104) & (g32) & (!g64)) + ((g153) & (!sk[100]) & (!g104) & (g32) & (g64)) + ((g153) & (!sk[100]) & (g104) & (!g32) & (!g64)) + ((g153) & (!sk[100]) & (g104) & (!g32) & (g64)) + ((g153) & (!sk[100]) & (g104) & (g32) & (!g64)) + ((g153) & (!sk[100]) & (g104) & (g32) & (g64)));
	assign g859 = (((!g9) & (!g18) & (!g27) & (g262) & (!sk[101]) & (!g858)) + ((!g9) & (!g18) & (!g27) & (g262) & (!sk[101]) & (g858)) + ((!g9) & (!g18) & (!g27) & (g262) & (sk[101]) & (g858)) + ((!g9) & (!g18) & (g27) & (!g262) & (!sk[101]) & (!g858)) + ((!g9) & (!g18) & (g27) & (!g262) & (!sk[101]) & (g858)) + ((!g9) & (!g18) & (g27) & (g262) & (!sk[101]) & (!g858)) + ((!g9) & (!g18) & (g27) & (g262) & (!sk[101]) & (g858)) + ((!g9) & (!g18) & (g27) & (g262) & (sk[101]) & (g858)) + ((!g9) & (g18) & (!g27) & (!g262) & (!sk[101]) & (!g858)) + ((!g9) & (g18) & (!g27) & (!g262) & (!sk[101]) & (g858)) + ((!g9) & (g18) & (!g27) & (g262) & (!sk[101]) & (!g858)) + ((!g9) & (g18) & (!g27) & (g262) & (!sk[101]) & (g858)) + ((!g9) & (g18) & (!g27) & (g262) & (sk[101]) & (g858)) + ((!g9) & (g18) & (g27) & (!g262) & (!sk[101]) & (!g858)) + ((!g9) & (g18) & (g27) & (!g262) & (!sk[101]) & (g858)) + ((!g9) & (g18) & (g27) & (g262) & (!sk[101]) & (!g858)) + ((!g9) & (g18) & (g27) & (g262) & (!sk[101]) & (g858)) + ((!g9) & (g18) & (g27) & (g262) & (sk[101]) & (g858)) + ((g9) & (!g18) & (!g27) & (g262) & (!sk[101]) & (!g858)) + ((g9) & (!g18) & (!g27) & (g262) & (!sk[101]) & (g858)) + ((g9) & (!g18) & (!g27) & (g262) & (sk[101]) & (g858)) + ((g9) & (!g18) & (g27) & (!g262) & (!sk[101]) & (!g858)) + ((g9) & (!g18) & (g27) & (!g262) & (!sk[101]) & (g858)) + ((g9) & (!g18) & (g27) & (g262) & (!sk[101]) & (!g858)) + ((g9) & (!g18) & (g27) & (g262) & (!sk[101]) & (g858)) + ((g9) & (g18) & (!g27) & (!g262) & (!sk[101]) & (!g858)) + ((g9) & (g18) & (!g27) & (!g262) & (!sk[101]) & (g858)) + ((g9) & (g18) & (!g27) & (g262) & (!sk[101]) & (!g858)) + ((g9) & (g18) & (!g27) & (g262) & (!sk[101]) & (g858)) + ((g9) & (g18) & (g27) & (!g262) & (!sk[101]) & (!g858)) + ((g9) & (g18) & (g27) & (!g262) & (!sk[101]) & (g858)) + ((g9) & (g18) & (g27) & (g262) & (!sk[101]) & (!g858)) + ((g9) & (g18) & (g27) & (g262) & (!sk[101]) & (g858)));
	assign g860 = (((!sk[102]) & (!g128) & (!g97) & (!g70) & (g12)) + ((!sk[102]) & (!g128) & (!g97) & (g70) & (g12)) + ((!sk[102]) & (!g128) & (g97) & (!g70) & (g12)) + ((!sk[102]) & (!g128) & (g97) & (g70) & (g12)) + ((!sk[102]) & (g128) & (!g97) & (!g70) & (!g12)) + ((!sk[102]) & (g128) & (!g97) & (!g70) & (g12)) + ((!sk[102]) & (g128) & (!g97) & (g70) & (!g12)) + ((!sk[102]) & (g128) & (!g97) & (g70) & (g12)) + ((!sk[102]) & (g128) & (g97) & (!g70) & (!g12)) + ((!sk[102]) & (g128) & (g97) & (!g70) & (g12)) + ((!sk[102]) & (g128) & (g97) & (g70) & (!g12)) + ((!sk[102]) & (g128) & (g97) & (g70) & (g12)) + ((sk[102]) & (!g128) & (!g97) & (g70) & (g12)) + ((sk[102]) & (!g128) & (g97) & (g70) & (g12)) + ((sk[102]) & (g128) & (!g97) & (g70) & (!g12)) + ((sk[102]) & (g128) & (!g97) & (g70) & (g12)) + ((sk[102]) & (g128) & (g97) & (g70) & (g12)));
	assign g861 = (((!sk[103]) & (!g160) & (!g194) & (!g236) & (g860)) + ((!sk[103]) & (!g160) & (!g194) & (g236) & (g860)) + ((!sk[103]) & (!g160) & (g194) & (!g236) & (g860)) + ((!sk[103]) & (!g160) & (g194) & (g236) & (g860)) + ((!sk[103]) & (g160) & (!g194) & (!g236) & (!g860)) + ((!sk[103]) & (g160) & (!g194) & (!g236) & (g860)) + ((!sk[103]) & (g160) & (!g194) & (g236) & (!g860)) + ((!sk[103]) & (g160) & (!g194) & (g236) & (g860)) + ((!sk[103]) & (g160) & (g194) & (!g236) & (!g860)) + ((!sk[103]) & (g160) & (g194) & (!g236) & (g860)) + ((!sk[103]) & (g160) & (g194) & (g236) & (!g860)) + ((!sk[103]) & (g160) & (g194) & (g236) & (g860)) + ((sk[103]) & (g160) & (!g194) & (!g236) & (!g860)));
	assign g862 = (((!g283) & (!g605) & (!sk[104]) & (!g857) & (g859) & (!g861)) + ((!g283) & (!g605) & (!sk[104]) & (!g857) & (g859) & (g861)) + ((!g283) & (!g605) & (!sk[104]) & (g857) & (!g859) & (!g861)) + ((!g283) & (!g605) & (!sk[104]) & (g857) & (!g859) & (g861)) + ((!g283) & (!g605) & (!sk[104]) & (g857) & (g859) & (!g861)) + ((!g283) & (!g605) & (!sk[104]) & (g857) & (g859) & (g861)) + ((!g283) & (g605) & (!sk[104]) & (!g857) & (!g859) & (!g861)) + ((!g283) & (g605) & (!sk[104]) & (!g857) & (!g859) & (g861)) + ((!g283) & (g605) & (!sk[104]) & (!g857) & (g859) & (!g861)) + ((!g283) & (g605) & (!sk[104]) & (!g857) & (g859) & (g861)) + ((!g283) & (g605) & (!sk[104]) & (g857) & (!g859) & (!g861)) + ((!g283) & (g605) & (!sk[104]) & (g857) & (!g859) & (g861)) + ((!g283) & (g605) & (!sk[104]) & (g857) & (g859) & (!g861)) + ((!g283) & (g605) & (!sk[104]) & (g857) & (g859) & (g861)) + ((g283) & (!g605) & (!sk[104]) & (!g857) & (g859) & (!g861)) + ((g283) & (!g605) & (!sk[104]) & (!g857) & (g859) & (g861)) + ((g283) & (!g605) & (!sk[104]) & (g857) & (!g859) & (!g861)) + ((g283) & (!g605) & (!sk[104]) & (g857) & (!g859) & (g861)) + ((g283) & (!g605) & (!sk[104]) & (g857) & (g859) & (!g861)) + ((g283) & (!g605) & (!sk[104]) & (g857) & (g859) & (g861)) + ((g283) & (g605) & (!sk[104]) & (!g857) & (!g859) & (!g861)) + ((g283) & (g605) & (!sk[104]) & (!g857) & (!g859) & (g861)) + ((g283) & (g605) & (!sk[104]) & (!g857) & (g859) & (!g861)) + ((g283) & (g605) & (!sk[104]) & (!g857) & (g859) & (g861)) + ((g283) & (g605) & (!sk[104]) & (g857) & (!g859) & (!g861)) + ((g283) & (g605) & (!sk[104]) & (g857) & (!g859) & (g861)) + ((g283) & (g605) & (!sk[104]) & (g857) & (g859) & (!g861)) + ((g283) & (g605) & (!sk[104]) & (g857) & (g859) & (g861)) + ((g283) & (g605) & (sk[104]) & (g857) & (g859) & (g861)));
	assign g863 = (((!g698) & (!g706) & (!g717) & (!g825) & (!g832) & (!g862)) + ((!g698) & (!g706) & (!g717) & (!g825) & (g832) & (!g862)) + ((!g698) & (!g706) & (!g717) & (g825) & (!g832) & (!g862)) + ((!g698) & (!g706) & (!g717) & (g825) & (g832) & (g862)) + ((!g698) & (!g706) & (g717) & (!g825) & (!g832) & (!g862)) + ((!g698) & (!g706) & (g717) & (!g825) & (g832) & (!g862)) + ((!g698) & (!g706) & (g717) & (g825) & (!g832) & (!g862)) + ((!g698) & (!g706) & (g717) & (g825) & (g832) & (g862)) + ((!g698) & (g706) & (!g717) & (!g825) & (!g832) & (!g862)) + ((!g698) & (g706) & (!g717) & (!g825) & (g832) & (!g862)) + ((!g698) & (g706) & (!g717) & (g825) & (!g832) & (!g862)) + ((!g698) & (g706) & (!g717) & (g825) & (g832) & (g862)) + ((!g698) & (g706) & (g717) & (!g825) & (!g832) & (!g862)) + ((!g698) & (g706) & (g717) & (!g825) & (g832) & (g862)) + ((!g698) & (g706) & (g717) & (g825) & (!g832) & (g862)) + ((!g698) & (g706) & (g717) & (g825) & (g832) & (g862)) + ((g698) & (!g706) & (!g717) & (!g825) & (!g832) & (!g862)) + ((g698) & (!g706) & (!g717) & (!g825) & (g832) & (!g862)) + ((g698) & (!g706) & (!g717) & (g825) & (!g832) & (!g862)) + ((g698) & (!g706) & (!g717) & (g825) & (g832) & (g862)) + ((g698) & (!g706) & (g717) & (!g825) & (!g832) & (!g862)) + ((g698) & (!g706) & (g717) & (!g825) & (g832) & (g862)) + ((g698) & (!g706) & (g717) & (g825) & (!g832) & (g862)) + ((g698) & (!g706) & (g717) & (g825) & (g832) & (g862)) + ((g698) & (g706) & (!g717) & (!g825) & (!g832) & (!g862)) + ((g698) & (g706) & (!g717) & (!g825) & (g832) & (g862)) + ((g698) & (g706) & (!g717) & (g825) & (!g832) & (g862)) + ((g698) & (g706) & (!g717) & (g825) & (g832) & (g862)) + ((g698) & (g706) & (g717) & (!g825) & (!g832) & (!g862)) + ((g698) & (g706) & (g717) & (!g825) & (g832) & (g862)) + ((g698) & (g706) & (g717) & (g825) & (!g832) & (g862)) + ((g698) & (g706) & (g717) & (g825) & (g832) & (g862)));
	assign g864 = (((!ax2x) & (!sk[106]) & (ax0x) & (!ax1x)) + ((!ax2x) & (!sk[106]) & (ax0x) & (ax1x)) + ((ax2x) & (!sk[106]) & (ax0x) & (!ax1x)) + ((ax2x) & (!sk[106]) & (ax0x) & (ax1x)) + ((ax2x) & (sk[106]) & (!ax0x) & (!ax1x)));
	assign g865 = (((g863) & (!sk[107]) & (g864)) + ((g863) & (sk[107]) & (g864)));
	assign g866 = (((!sk[108]) & (!ax22x) & (ax0x) & (!ax1x)) + ((!sk[108]) & (!ax22x) & (ax0x) & (ax1x)) + ((!sk[108]) & (ax22x) & (ax0x) & (!ax1x)) + ((!sk[108]) & (ax22x) & (ax0x) & (ax1x)) + ((sk[108]) & (!ax22x) & (!ax0x) & (ax1x)) + ((sk[108]) & (!ax22x) & (ax0x) & (!ax1x)) + ((sk[108]) & (ax22x) & (!ax0x) & (ax1x)) + ((sk[108]) & (ax22x) & (ax0x) & (ax1x)));
	assign g867 = (((!g683) & (sk[109]) & (g866)) + ((g683) & (!sk[109]) & (g866)) + ((g683) & (sk[109]) & (!g866)));
	assign g868 = (((!sk[110]) & (ax0x) & (g867)) + ((sk[110]) & (ax0x) & (g867)));
	assign g869 = (((!sk[111]) & (g707) & (g717)) + ((sk[111]) & (!g707) & (g717)) + ((sk[111]) & (g707) & (!g717)));
	assign g870 = (((!g698) & (!g706) & (!g717) & (!g825) & (sk[112]) & (g832)) + ((!g698) & (!g706) & (!g717) & (g825) & (!sk[112]) & (!g832)) + ((!g698) & (!g706) & (!g717) & (g825) & (!sk[112]) & (g832)) + ((!g698) & (!g706) & (!g717) & (g825) & (sk[112]) & (!g832)) + ((!g698) & (!g706) & (g717) & (!g825) & (!sk[112]) & (!g832)) + ((!g698) & (!g706) & (g717) & (!g825) & (!sk[112]) & (g832)) + ((!g698) & (!g706) & (g717) & (!g825) & (sk[112]) & (g832)) + ((!g698) & (!g706) & (g717) & (g825) & (!sk[112]) & (!g832)) + ((!g698) & (!g706) & (g717) & (g825) & (!sk[112]) & (g832)) + ((!g698) & (!g706) & (g717) & (g825) & (sk[112]) & (!g832)) + ((!g698) & (g706) & (!g717) & (!g825) & (!sk[112]) & (!g832)) + ((!g698) & (g706) & (!g717) & (!g825) & (!sk[112]) & (g832)) + ((!g698) & (g706) & (!g717) & (!g825) & (sk[112]) & (g832)) + ((!g698) & (g706) & (!g717) & (g825) & (!sk[112]) & (!g832)) + ((!g698) & (g706) & (!g717) & (g825) & (!sk[112]) & (g832)) + ((!g698) & (g706) & (!g717) & (g825) & (sk[112]) & (!g832)) + ((!g698) & (g706) & (g717) & (!g825) & (!sk[112]) & (!g832)) + ((!g698) & (g706) & (g717) & (!g825) & (!sk[112]) & (g832)) + ((!g698) & (g706) & (g717) & (!g825) & (sk[112]) & (!g832)) + ((!g698) & (g706) & (g717) & (g825) & (!sk[112]) & (!g832)) + ((!g698) & (g706) & (g717) & (g825) & (!sk[112]) & (g832)) + ((!g698) & (g706) & (g717) & (g825) & (sk[112]) & (g832)) + ((g698) & (!g706) & (!g717) & (!g825) & (sk[112]) & (g832)) + ((g698) & (!g706) & (!g717) & (g825) & (!sk[112]) & (!g832)) + ((g698) & (!g706) & (!g717) & (g825) & (!sk[112]) & (g832)) + ((g698) & (!g706) & (!g717) & (g825) & (sk[112]) & (!g832)) + ((g698) & (!g706) & (g717) & (!g825) & (!sk[112]) & (!g832)) + ((g698) & (!g706) & (g717) & (!g825) & (!sk[112]) & (g832)) + ((g698) & (!g706) & (g717) & (!g825) & (sk[112]) & (!g832)) + ((g698) & (!g706) & (g717) & (g825) & (!sk[112]) & (!g832)) + ((g698) & (!g706) & (g717) & (g825) & (!sk[112]) & (g832)) + ((g698) & (!g706) & (g717) & (g825) & (sk[112]) & (g832)) + ((g698) & (g706) & (!g717) & (!g825) & (!sk[112]) & (!g832)) + ((g698) & (g706) & (!g717) & (!g825) & (!sk[112]) & (g832)) + ((g698) & (g706) & (!g717) & (!g825) & (sk[112]) & (!g832)) + ((g698) & (g706) & (!g717) & (g825) & (!sk[112]) & (!g832)) + ((g698) & (g706) & (!g717) & (g825) & (!sk[112]) & (g832)) + ((g698) & (g706) & (!g717) & (g825) & (sk[112]) & (g832)) + ((g698) & (g706) & (g717) & (!g825) & (!sk[112]) & (!g832)) + ((g698) & (g706) & (g717) & (!g825) & (!sk[112]) & (g832)) + ((g698) & (g706) & (g717) & (!g825) & (sk[112]) & (!g832)) + ((g698) & (g706) & (g717) & (g825) & (!sk[112]) & (!g832)) + ((g698) & (g706) & (g717) & (g825) & (!sk[112]) & (g832)) + ((g698) & (g706) & (g717) & (g825) & (sk[112]) & (g832)));
	assign g871 = (((!g698) & (!g706) & (!g717) & (g825) & (g832) & (g862)) + ((!g698) & (!g706) & (g717) & (g825) & (g832) & (g862)) + ((!g698) & (g706) & (!g717) & (g825) & (g832) & (g862)) + ((!g698) & (g706) & (g717) & (!g825) & (g832) & (g862)) + ((!g698) & (g706) & (g717) & (g825) & (!g832) & (g862)) + ((!g698) & (g706) & (g717) & (g825) & (g832) & (g862)) + ((g698) & (!g706) & (!g717) & (g825) & (g832) & (g862)) + ((g698) & (!g706) & (g717) & (!g825) & (g832) & (g862)) + ((g698) & (!g706) & (g717) & (g825) & (!g832) & (g862)) + ((g698) & (!g706) & (g717) & (g825) & (g832) & (g862)) + ((g698) & (g706) & (!g717) & (!g825) & (g832) & (g862)) + ((g698) & (g706) & (!g717) & (g825) & (!g832) & (g862)) + ((g698) & (g706) & (!g717) & (g825) & (g832) & (g862)) + ((g698) & (g706) & (g717) & (!g825) & (g832) & (g862)) + ((g698) & (g706) & (g717) & (g825) & (!g832) & (g862)) + ((g698) & (g706) & (g717) & (g825) & (g832) & (g862)));
	assign g872 = (((!sk[114]) & (!g9) & (!g40) & (!g29) & (g131)) + ((!sk[114]) & (!g9) & (!g40) & (g29) & (g131)) + ((!sk[114]) & (!g9) & (g40) & (!g29) & (g131)) + ((!sk[114]) & (!g9) & (g40) & (g29) & (g131)) + ((!sk[114]) & (g9) & (!g40) & (!g29) & (!g131)) + ((!sk[114]) & (g9) & (!g40) & (!g29) & (g131)) + ((!sk[114]) & (g9) & (!g40) & (g29) & (!g131)) + ((!sk[114]) & (g9) & (!g40) & (g29) & (g131)) + ((!sk[114]) & (g9) & (g40) & (!g29) & (!g131)) + ((!sk[114]) & (g9) & (g40) & (!g29) & (g131)) + ((!sk[114]) & (g9) & (g40) & (g29) & (!g131)) + ((!sk[114]) & (g9) & (g40) & (g29) & (g131)) + ((sk[114]) & (!g9) & (!g40) & (!g29) & (!g131)) + ((sk[114]) & (!g9) & (g40) & (!g29) & (!g131)) + ((sk[114]) & (g9) & (!g40) & (!g29) & (!g131)));
	assign g873 = (((!g62) & (!g18) & (!sk[115]) & (!g593) & (g241) & (!g673)) + ((!g62) & (!g18) & (!sk[115]) & (!g593) & (g241) & (g673)) + ((!g62) & (!g18) & (!sk[115]) & (g593) & (!g241) & (!g673)) + ((!g62) & (!g18) & (!sk[115]) & (g593) & (!g241) & (g673)) + ((!g62) & (!g18) & (!sk[115]) & (g593) & (g241) & (!g673)) + ((!g62) & (!g18) & (!sk[115]) & (g593) & (g241) & (g673)) + ((!g62) & (!g18) & (sk[115]) & (!g593) & (!g241) & (g673)) + ((!g62) & (g18) & (!sk[115]) & (!g593) & (!g241) & (!g673)) + ((!g62) & (g18) & (!sk[115]) & (!g593) & (!g241) & (g673)) + ((!g62) & (g18) & (!sk[115]) & (!g593) & (g241) & (!g673)) + ((!g62) & (g18) & (!sk[115]) & (!g593) & (g241) & (g673)) + ((!g62) & (g18) & (!sk[115]) & (g593) & (!g241) & (!g673)) + ((!g62) & (g18) & (!sk[115]) & (g593) & (!g241) & (g673)) + ((!g62) & (g18) & (!sk[115]) & (g593) & (g241) & (!g673)) + ((!g62) & (g18) & (!sk[115]) & (g593) & (g241) & (g673)) + ((!g62) & (g18) & (sk[115]) & (!g593) & (!g241) & (g673)) + ((g62) & (!g18) & (!sk[115]) & (!g593) & (g241) & (!g673)) + ((g62) & (!g18) & (!sk[115]) & (!g593) & (g241) & (g673)) + ((g62) & (!g18) & (!sk[115]) & (g593) & (!g241) & (!g673)) + ((g62) & (!g18) & (!sk[115]) & (g593) & (!g241) & (g673)) + ((g62) & (!g18) & (!sk[115]) & (g593) & (g241) & (!g673)) + ((g62) & (!g18) & (!sk[115]) & (g593) & (g241) & (g673)) + ((g62) & (!g18) & (sk[115]) & (!g593) & (!g241) & (g673)) + ((g62) & (g18) & (!sk[115]) & (!g593) & (!g241) & (!g673)) + ((g62) & (g18) & (!sk[115]) & (!g593) & (!g241) & (g673)) + ((g62) & (g18) & (!sk[115]) & (!g593) & (g241) & (!g673)) + ((g62) & (g18) & (!sk[115]) & (!g593) & (g241) & (g673)) + ((g62) & (g18) & (!sk[115]) & (g593) & (!g241) & (!g673)) + ((g62) & (g18) & (!sk[115]) & (g593) & (!g241) & (g673)) + ((g62) & (g18) & (!sk[115]) & (g593) & (g241) & (!g673)) + ((g62) & (g18) & (!sk[115]) & (g593) & (g241) & (g673)));
	assign g874 = (((!g71) & (!g58) & (!sk[116]) & (!g272) & (g194)) + ((!g71) & (!g58) & (!sk[116]) & (g272) & (g194)) + ((!g71) & (!g58) & (sk[116]) & (!g272) & (!g194)) + ((!g71) & (g58) & (!sk[116]) & (!g272) & (g194)) + ((!g71) & (g58) & (!sk[116]) & (g272) & (g194)) + ((!g71) & (g58) & (sk[116]) & (!g272) & (!g194)) + ((g71) & (!g58) & (!sk[116]) & (!g272) & (!g194)) + ((g71) & (!g58) & (!sk[116]) & (!g272) & (g194)) + ((g71) & (!g58) & (!sk[116]) & (g272) & (!g194)) + ((g71) & (!g58) & (!sk[116]) & (g272) & (g194)) + ((g71) & (!g58) & (sk[116]) & (!g272) & (!g194)) + ((g71) & (g58) & (!sk[116]) & (!g272) & (!g194)) + ((g71) & (g58) & (!sk[116]) & (!g272) & (g194)) + ((g71) & (g58) & (!sk[116]) & (g272) & (!g194)) + ((g71) & (g58) & (!sk[116]) & (g272) & (g194)));
	assign g875 = (((!g114) & (!g115) & (!g8) & (!g40) & (!g20) & (g874)) + ((!g114) & (!g115) & (!g8) & (!g40) & (g20) & (g874)) + ((!g114) & (!g115) & (!g8) & (g40) & (!g20) & (g874)) + ((!g114) & (!g115) & (!g8) & (g40) & (g20) & (g874)) + ((!g114) & (!g115) & (g8) & (!g40) & (!g20) & (g874)) + ((!g114) & (!g115) & (g8) & (g40) & (!g20) & (g874)) + ((!g114) & (g115) & (!g8) & (!g40) & (!g20) & (g874)) + ((!g114) & (g115) & (!g8) & (g40) & (!g20) & (g874)) + ((!g114) & (g115) & (g8) & (!g40) & (!g20) & (g874)) + ((!g114) & (g115) & (g8) & (!g40) & (g20) & (g874)) + ((!g114) & (g115) & (g8) & (g40) & (!g20) & (g874)) + ((!g114) & (g115) & (g8) & (g40) & (g20) & (g874)) + ((g114) & (!g115) & (!g8) & (!g40) & (!g20) & (g874)) + ((g114) & (!g115) & (!g8) & (!g40) & (g20) & (g874)) + ((g114) & (!g115) & (g8) & (!g40) & (!g20) & (g874)) + ((g114) & (!g115) & (g8) & (!g40) & (g20) & (g874)) + ((g114) & (!g115) & (g8) & (g40) & (!g20) & (g874)) + ((g114) & (!g115) & (g8) & (g40) & (g20) & (g874)) + ((g114) & (g115) & (!g8) & (!g40) & (!g20) & (g874)) + ((g114) & (g115) & (!g8) & (!g40) & (g20) & (g874)) + ((g114) & (g115) & (!g8) & (g40) & (!g20) & (g874)) + ((g114) & (g115) & (!g8) & (g40) & (g20) & (g874)) + ((g114) & (g115) & (g8) & (!g40) & (!g20) & (g874)) + ((g114) & (g115) & (g8) & (!g40) & (g20) & (g874)) + ((g114) & (g115) & (g8) & (g40) & (!g20) & (g874)) + ((g114) & (g115) & (g8) & (g40) & (g20) & (g874)));
	assign g876 = (((!g9) & (!g30) & (!g62) & (!g66) & (!g20) & (!g354)) + ((!g9) & (!g30) & (!g62) & (!g66) & (g20) & (!g354)) + ((!g9) & (!g30) & (!g62) & (g66) & (!g20) & (!g354)) + ((!g9) & (!g30) & (!g62) & (g66) & (g20) & (!g354)) + ((!g9) & (!g30) & (g62) & (!g66) & (!g20) & (!g354)) + ((!g9) & (g30) & (!g62) & (!g66) & (!g20) & (!g354)) + ((!g9) & (g30) & (!g62) & (!g66) & (g20) & (!g354)) + ((!g9) & (g30) & (!g62) & (g66) & (!g20) & (!g354)) + ((!g9) & (g30) & (!g62) & (g66) & (g20) & (!g354)) + ((!g9) & (g30) & (g62) & (!g66) & (!g20) & (!g354)) + ((g9) & (!g30) & (!g62) & (!g66) & (!g20) & (!g354)) + ((g9) & (!g30) & (!g62) & (!g66) & (g20) & (!g354)) + ((g9) & (!g30) & (!g62) & (g66) & (!g20) & (!g354)) + ((g9) & (!g30) & (!g62) & (g66) & (g20) & (!g354)) + ((g9) & (!g30) & (g62) & (!g66) & (!g20) & (!g354)));
	assign g877 = (((!g284) & (g636) & (g872) & (g873) & (g875) & (g876)));
	assign g878 = (((!sk[120]) & (g563) & (g877)) + ((sk[120]) & (!g563) & (g877)));
	assign g879 = (((!g47) & (!g105) & (sk[121]) & (!g59)) + ((!g47) & (g105) & (!sk[121]) & (!g59)) + ((!g47) & (g105) & (!sk[121]) & (g59)) + ((g47) & (g105) & (!sk[121]) & (!g59)) + ((g47) & (g105) & (!sk[121]) & (g59)));
	assign g880 = (((!g9) & (!g10) & (!g99) & (!g104) & (sk[122]) & (!g32)) + ((!g9) & (!g10) & (!g99) & (!g104) & (sk[122]) & (g32)) + ((!g9) & (!g10) & (!g99) & (g104) & (!sk[122]) & (!g32)) + ((!g9) & (!g10) & (!g99) & (g104) & (!sk[122]) & (g32)) + ((!g9) & (!g10) & (!g99) & (g104) & (sk[122]) & (!g32)) + ((!g9) & (!g10) & (!g99) & (g104) & (sk[122]) & (g32)) + ((!g9) & (!g10) & (g99) & (!g104) & (!sk[122]) & (!g32)) + ((!g9) & (!g10) & (g99) & (!g104) & (!sk[122]) & (g32)) + ((!g9) & (!g10) & (g99) & (!g104) & (sk[122]) & (!g32)) + ((!g9) & (!g10) & (g99) & (!g104) & (sk[122]) & (g32)) + ((!g9) & (!g10) & (g99) & (g104) & (!sk[122]) & (!g32)) + ((!g9) & (!g10) & (g99) & (g104) & (!sk[122]) & (g32)) + ((!g9) & (!g10) & (g99) & (g104) & (sk[122]) & (!g32)) + ((!g9) & (!g10) & (g99) & (g104) & (sk[122]) & (g32)) + ((!g9) & (g10) & (!g99) & (!g104) & (!sk[122]) & (!g32)) + ((!g9) & (g10) & (!g99) & (!g104) & (!sk[122]) & (g32)) + ((!g9) & (g10) & (!g99) & (!g104) & (sk[122]) & (!g32)) + ((!g9) & (g10) & (!g99) & (!g104) & (sk[122]) & (g32)) + ((!g9) & (g10) & (!g99) & (g104) & (!sk[122]) & (!g32)) + ((!g9) & (g10) & (!g99) & (g104) & (!sk[122]) & (g32)) + ((!g9) & (g10) & (g99) & (!g104) & (!sk[122]) & (!g32)) + ((!g9) & (g10) & (g99) & (!g104) & (!sk[122]) & (g32)) + ((!g9) & (g10) & (g99) & (g104) & (!sk[122]) & (!g32)) + ((!g9) & (g10) & (g99) & (g104) & (!sk[122]) & (g32)) + ((g9) & (!g10) & (!g99) & (!g104) & (sk[122]) & (!g32)) + ((g9) & (!g10) & (!g99) & (g104) & (!sk[122]) & (!g32)) + ((g9) & (!g10) & (!g99) & (g104) & (!sk[122]) & (g32)) + ((g9) & (!g10) & (!g99) & (g104) & (sk[122]) & (!g32)) + ((g9) & (!g10) & (g99) & (!g104) & (!sk[122]) & (!g32)) + ((g9) & (!g10) & (g99) & (!g104) & (!sk[122]) & (g32)) + ((g9) & (!g10) & (g99) & (!g104) & (sk[122]) & (!g32)) + ((g9) & (!g10) & (g99) & (g104) & (!sk[122]) & (!g32)) + ((g9) & (!g10) & (g99) & (g104) & (!sk[122]) & (g32)) + ((g9) & (!g10) & (g99) & (g104) & (sk[122]) & (!g32)) + ((g9) & (g10) & (!g99) & (!g104) & (!sk[122]) & (!g32)) + ((g9) & (g10) & (!g99) & (!g104) & (!sk[122]) & (g32)) + ((g9) & (g10) & (!g99) & (!g104) & (sk[122]) & (!g32)) + ((g9) & (g10) & (!g99) & (g104) & (!sk[122]) & (!g32)) + ((g9) & (g10) & (!g99) & (g104) & (!sk[122]) & (g32)) + ((g9) & (g10) & (g99) & (!g104) & (!sk[122]) & (!g32)) + ((g9) & (g10) & (g99) & (!g104) & (!sk[122]) & (g32)) + ((g9) & (g10) & (g99) & (g104) & (!sk[122]) & (!g32)) + ((g9) & (g10) & (g99) & (g104) & (!sk[122]) & (g32)));
	assign g881 = (((!g70) & (!g16) & (!g30) & (!sk[123]) & (g551) & (!g880)) + ((!g70) & (!g16) & (!g30) & (!sk[123]) & (g551) & (g880)) + ((!g70) & (!g16) & (!g30) & (sk[123]) & (!g551) & (g880)) + ((!g70) & (!g16) & (g30) & (!sk[123]) & (!g551) & (!g880)) + ((!g70) & (!g16) & (g30) & (!sk[123]) & (!g551) & (g880)) + ((!g70) & (!g16) & (g30) & (!sk[123]) & (g551) & (!g880)) + ((!g70) & (!g16) & (g30) & (!sk[123]) & (g551) & (g880)) + ((!g70) & (!g16) & (g30) & (sk[123]) & (!g551) & (g880)) + ((!g70) & (g16) & (!g30) & (!sk[123]) & (!g551) & (!g880)) + ((!g70) & (g16) & (!g30) & (!sk[123]) & (!g551) & (g880)) + ((!g70) & (g16) & (!g30) & (!sk[123]) & (g551) & (!g880)) + ((!g70) & (g16) & (!g30) & (!sk[123]) & (g551) & (g880)) + ((!g70) & (g16) & (!g30) & (sk[123]) & (!g551) & (g880)) + ((!g70) & (g16) & (g30) & (!sk[123]) & (!g551) & (!g880)) + ((!g70) & (g16) & (g30) & (!sk[123]) & (!g551) & (g880)) + ((!g70) & (g16) & (g30) & (!sk[123]) & (g551) & (!g880)) + ((!g70) & (g16) & (g30) & (!sk[123]) & (g551) & (g880)) + ((g70) & (!g16) & (!g30) & (!sk[123]) & (g551) & (!g880)) + ((g70) & (!g16) & (!g30) & (!sk[123]) & (g551) & (g880)) + ((g70) & (!g16) & (!g30) & (sk[123]) & (!g551) & (g880)) + ((g70) & (!g16) & (g30) & (!sk[123]) & (!g551) & (!g880)) + ((g70) & (!g16) & (g30) & (!sk[123]) & (!g551) & (g880)) + ((g70) & (!g16) & (g30) & (!sk[123]) & (g551) & (!g880)) + ((g70) & (!g16) & (g30) & (!sk[123]) & (g551) & (g880)) + ((g70) & (g16) & (!g30) & (!sk[123]) & (!g551) & (!g880)) + ((g70) & (g16) & (!g30) & (!sk[123]) & (!g551) & (g880)) + ((g70) & (g16) & (!g30) & (!sk[123]) & (g551) & (!g880)) + ((g70) & (g16) & (!g30) & (!sk[123]) & (g551) & (g880)) + ((g70) & (g16) & (!g30) & (sk[123]) & (!g551) & (g880)) + ((g70) & (g16) & (g30) & (!sk[123]) & (!g551) & (!g880)) + ((g70) & (g16) & (g30) & (!sk[123]) & (!g551) & (g880)) + ((g70) & (g16) & (g30) & (!sk[123]) & (g551) & (!g880)) + ((g70) & (g16) & (g30) & (!sk[123]) & (g551) & (g880)));
	assign g882 = (((g879) & (!g43) & (!g187) & (!g601) & (!g137) & (g881)));
	assign g883 = (((!g64) & (!g95) & (g245) & (g89) & (g878) & (g882)));
	assign g884 = (((!g869) & (!g870) & (!g834) & (!g871) & (!g883) & (g863)) + ((!g869) & (!g870) & (!g834) & (!g871) & (g883) & (g863)) + ((!g869) & (!g870) & (!g834) & (g871) & (!g883) & (g863)) + ((!g869) & (!g870) & (!g834) & (g871) & (g883) & (g863)) + ((!g869) & (!g870) & (g834) & (!g871) & (!g883) & (!g863)) + ((!g869) & (!g870) & (g834) & (!g871) & (!g883) & (g863)) + ((!g869) & (!g870) & (g834) & (!g871) & (g883) & (g863)) + ((!g869) & (!g870) & (g834) & (g871) & (!g883) & (g863)) + ((!g869) & (!g870) & (g834) & (g871) & (g883) & (!g863)) + ((!g869) & (!g870) & (g834) & (g871) & (g883) & (g863)) + ((!g869) & (g870) & (!g834) & (!g871) & (!g883) & (g863)) + ((!g869) & (g870) & (!g834) & (g871) & (g883) & (g863)) + ((!g869) & (g870) & (g834) & (!g871) & (!g883) & (g863)) + ((!g869) & (g870) & (g834) & (g871) & (g883) & (g863)) + ((g869) & (!g870) & (!g834) & (!g871) & (!g883) & (!g863)) + ((g869) & (!g870) & (!g834) & (!g871) & (!g883) & (g863)) + ((g869) & (!g870) & (!g834) & (!g871) & (g883) & (g863)) + ((g869) & (!g870) & (!g834) & (g871) & (!g883) & (g863)) + ((g869) & (!g870) & (!g834) & (g871) & (g883) & (!g863)) + ((g869) & (!g870) & (!g834) & (g871) & (g883) & (g863)) + ((g869) & (!g870) & (g834) & (!g871) & (!g883) & (!g863)) + ((g869) & (!g870) & (g834) & (!g871) & (!g883) & (g863)) + ((g869) & (!g870) & (g834) & (!g871) & (g883) & (g863)) + ((g869) & (!g870) & (g834) & (g871) & (!g883) & (g863)) + ((g869) & (!g870) & (g834) & (g871) & (g883) & (!g863)) + ((g869) & (!g870) & (g834) & (g871) & (g883) & (g863)) + ((g869) & (g870) & (!g834) & (!g871) & (!g883) & (g863)) + ((g869) & (g870) & (!g834) & (g871) & (g883) & (g863)) + ((g869) & (g870) & (g834) & (!g871) & (!g883) & (g863)) + ((g869) & (g870) & (g834) & (!g871) & (g883) & (g863)) + ((g869) & (g870) & (g834) & (g871) & (!g883) & (g863)) + ((g869) & (g870) & (g834) & (g871) & (g883) & (g863)));
	assign g885 = (((!g92) & (!g210) & (!g211) & (!sk[127]) & (g212)) + ((!g92) & (!g210) & (g211) & (!sk[127]) & (g212)) + ((!g92) & (g210) & (!g211) & (!sk[127]) & (g212)) + ((!g92) & (g210) & (g211) & (!sk[127]) & (g212)) + ((g92) & (!g210) & (!g211) & (!sk[127]) & (!g212)) + ((g92) & (!g210) & (!g211) & (!sk[127]) & (g212)) + ((g92) & (!g210) & (!g211) & (sk[127]) & (g212)) + ((g92) & (!g210) & (g211) & (!sk[127]) & (!g212)) + ((g92) & (!g210) & (g211) & (!sk[127]) & (g212)) + ((g92) & (g210) & (!g211) & (!sk[127]) & (!g212)) + ((g92) & (g210) & (!g211) & (!sk[127]) & (g212)) + ((g92) & (g210) & (g211) & (!sk[127]) & (!g212)) + ((g92) & (g210) & (g211) & (!sk[127]) & (g212)));
	assign g886 = (((!g146) & (!g152) & (!sk[0]) & (!g268) & (g710)) + ((!g146) & (!g152) & (!sk[0]) & (g268) & (g710)) + ((!g146) & (!g152) & (sk[0]) & (!g268) & (!g710)) + ((!g146) & (g152) & (!sk[0]) & (!g268) & (g710)) + ((!g146) & (g152) & (!sk[0]) & (g268) & (g710)) + ((g146) & (!g152) & (!sk[0]) & (!g268) & (!g710)) + ((g146) & (!g152) & (!sk[0]) & (!g268) & (g710)) + ((g146) & (!g152) & (!sk[0]) & (g268) & (!g710)) + ((g146) & (!g152) & (!sk[0]) & (g268) & (g710)) + ((g146) & (g152) & (!sk[0]) & (!g268) & (!g710)) + ((g146) & (g152) & (!sk[0]) & (!g268) & (g710)) + ((g146) & (g152) & (!sk[0]) & (g268) & (!g710)) + ((g146) & (g152) & (!sk[0]) & (g268) & (g710)));
	assign g887 = (((!g112) & (!g113) & (!g97) & (!g98) & (!g71) & (g104)) + ((!g112) & (!g113) & (!g97) & (!g98) & (g71) & (g104)) + ((!g112) & (!g113) & (!g97) & (g98) & (!g71) & (g104)) + ((!g112) & (!g113) & (!g97) & (g98) & (g71) & (g104)) + ((!g112) & (!g113) & (g97) & (!g98) & (!g71) & (g104)) + ((!g112) & (!g113) & (g97) & (!g98) & (g71) & (g104)) + ((!g112) & (g113) & (!g97) & (!g98) & (!g71) & (g104)) + ((!g112) & (g113) & (!g97) & (!g98) & (g71) & (g104)) + ((!g112) & (g113) & (g97) & (g98) & (g71) & (!g104)) + ((!g112) & (g113) & (g97) & (g98) & (g71) & (g104)) + ((g112) & (g113) & (g97) & (g98) & (g71) & (!g104)) + ((g112) & (g113) & (g97) & (g98) & (g71) & (g104)));
	assign g888 = (((!g45) & (!sk[2]) & (!g559) & (!g608) & (g886) & (!g887)) + ((!g45) & (!sk[2]) & (!g559) & (!g608) & (g886) & (g887)) + ((!g45) & (!sk[2]) & (!g559) & (g608) & (!g886) & (!g887)) + ((!g45) & (!sk[2]) & (!g559) & (g608) & (!g886) & (g887)) + ((!g45) & (!sk[2]) & (!g559) & (g608) & (g886) & (!g887)) + ((!g45) & (!sk[2]) & (!g559) & (g608) & (g886) & (g887)) + ((!g45) & (!sk[2]) & (g559) & (!g608) & (!g886) & (!g887)) + ((!g45) & (!sk[2]) & (g559) & (!g608) & (!g886) & (g887)) + ((!g45) & (!sk[2]) & (g559) & (!g608) & (g886) & (!g887)) + ((!g45) & (!sk[2]) & (g559) & (!g608) & (g886) & (g887)) + ((!g45) & (!sk[2]) & (g559) & (g608) & (!g886) & (!g887)) + ((!g45) & (!sk[2]) & (g559) & (g608) & (!g886) & (g887)) + ((!g45) & (!sk[2]) & (g559) & (g608) & (g886) & (!g887)) + ((!g45) & (!sk[2]) & (g559) & (g608) & (g886) & (g887)) + ((g45) & (!sk[2]) & (!g559) & (!g608) & (g886) & (!g887)) + ((g45) & (!sk[2]) & (!g559) & (!g608) & (g886) & (g887)) + ((g45) & (!sk[2]) & (!g559) & (g608) & (!g886) & (!g887)) + ((g45) & (!sk[2]) & (!g559) & (g608) & (!g886) & (g887)) + ((g45) & (!sk[2]) & (!g559) & (g608) & (g886) & (!g887)) + ((g45) & (!sk[2]) & (!g559) & (g608) & (g886) & (g887)) + ((g45) & (!sk[2]) & (g559) & (!g608) & (!g886) & (!g887)) + ((g45) & (!sk[2]) & (g559) & (!g608) & (!g886) & (g887)) + ((g45) & (!sk[2]) & (g559) & (!g608) & (g886) & (!g887)) + ((g45) & (!sk[2]) & (g559) & (!g608) & (g886) & (g887)) + ((g45) & (!sk[2]) & (g559) & (g608) & (!g886) & (!g887)) + ((g45) & (!sk[2]) & (g559) & (g608) & (!g886) & (g887)) + ((g45) & (!sk[2]) & (g559) & (g608) & (g886) & (!g887)) + ((g45) & (!sk[2]) & (g559) & (g608) & (g886) & (g887)) + ((g45) & (sk[2]) & (g559) & (g608) & (g886) & (!g887)));
	assign g889 = (((!sk[3]) & (g885) & (g888)) + ((sk[3]) & (g885) & (g888)));
	assign g890 = (((!sk[4]) & (!g889) & (g871) & (!g883)) + ((!sk[4]) & (!g889) & (g871) & (g883)) + ((!sk[4]) & (g889) & (g871) & (!g883)) + ((!sk[4]) & (g889) & (g871) & (g883)) + ((sk[4]) & (!g889) & (!g871) & (!g883)) + ((sk[4]) & (g889) & (!g871) & (g883)) + ((sk[4]) & (g889) & (g871) & (!g883)) + ((sk[4]) & (g889) & (g871) & (g883)));
	assign g891 = (((!sk[5]) & (ax0x) & (g867)) + ((sk[5]) & (ax0x) & (!g867)));
	assign g892 = (((!sk[6]) & (ax0x) & (ax1x)) + ((sk[6]) & (!ax0x) & (ax1x)));
	assign g893 = (((!g891) & (!g889) & (!sk[7]) & (!g871) & (g883) & (!g892)) + ((!g891) & (!g889) & (!sk[7]) & (!g871) & (g883) & (g892)) + ((!g891) & (!g889) & (!sk[7]) & (g871) & (!g883) & (!g892)) + ((!g891) & (!g889) & (!sk[7]) & (g871) & (!g883) & (g892)) + ((!g891) & (!g889) & (!sk[7]) & (g871) & (g883) & (!g892)) + ((!g891) & (!g889) & (!sk[7]) & (g871) & (g883) & (g892)) + ((!g891) & (!g889) & (sk[7]) & (!g871) & (!g883) & (g892)) + ((!g891) & (!g889) & (sk[7]) & (g871) & (g883) & (g892)) + ((!g891) & (g889) & (!sk[7]) & (!g871) & (!g883) & (!g892)) + ((!g891) & (g889) & (!sk[7]) & (!g871) & (!g883) & (g892)) + ((!g891) & (g889) & (!sk[7]) & (!g871) & (g883) & (!g892)) + ((!g891) & (g889) & (!sk[7]) & (!g871) & (g883) & (g892)) + ((!g891) & (g889) & (!sk[7]) & (g871) & (!g883) & (!g892)) + ((!g891) & (g889) & (!sk[7]) & (g871) & (!g883) & (g892)) + ((!g891) & (g889) & (!sk[7]) & (g871) & (g883) & (!g892)) + ((!g891) & (g889) & (!sk[7]) & (g871) & (g883) & (g892)) + ((!g891) & (g889) & (sk[7]) & (!g871) & (!g883) & (g892)) + ((!g891) & (g889) & (sk[7]) & (g871) & (g883) & (g892)) + ((g891) & (!g889) & (!sk[7]) & (!g871) & (g883) & (!g892)) + ((g891) & (!g889) & (!sk[7]) & (!g871) & (g883) & (g892)) + ((g891) & (!g889) & (!sk[7]) & (g871) & (!g883) & (!g892)) + ((g891) & (!g889) & (!sk[7]) & (g871) & (!g883) & (g892)) + ((g891) & (!g889) & (!sk[7]) & (g871) & (g883) & (!g892)) + ((g891) & (!g889) & (!sk[7]) & (g871) & (g883) & (g892)) + ((g891) & (!g889) & (sk[7]) & (!g871) & (!g883) & (!g892)) + ((g891) & (!g889) & (sk[7]) & (!g871) & (!g883) & (g892)) + ((g891) & (!g889) & (sk[7]) & (!g871) & (g883) & (!g892)) + ((g891) & (!g889) & (sk[7]) & (!g871) & (g883) & (g892)) + ((g891) & (!g889) & (sk[7]) & (g871) & (!g883) & (!g892)) + ((g891) & (!g889) & (sk[7]) & (g871) & (!g883) & (g892)) + ((g891) & (!g889) & (sk[7]) & (g871) & (g883) & (g892)) + ((g891) & (g889) & (!sk[7]) & (!g871) & (!g883) & (!g892)) + ((g891) & (g889) & (!sk[7]) & (!g871) & (!g883) & (g892)) + ((g891) & (g889) & (!sk[7]) & (!g871) & (g883) & (!g892)) + ((g891) & (g889) & (!sk[7]) & (!g871) & (g883) & (g892)) + ((g891) & (g889) & (!sk[7]) & (g871) & (!g883) & (!g892)) + ((g891) & (g889) & (!sk[7]) & (g871) & (!g883) & (g892)) + ((g891) & (g889) & (!sk[7]) & (g871) & (g883) & (!g892)) + ((g891) & (g889) & (!sk[7]) & (g871) & (g883) & (g892)) + ((g891) & (g889) & (sk[7]) & (!g871) & (!g883) & (g892)) + ((g891) & (g889) & (sk[7]) & (g871) & (g883) & (!g892)) + ((g891) & (g889) & (sk[7]) & (g871) & (g883) & (g892)));
	assign g894 = (((!g683) & (!g865) & (!g868) & (!g884) & (!g890) & (!g893)) + ((!g683) & (!g865) & (!g868) & (!g884) & (g890) & (!g893)) + ((!g683) & (!g865) & (!g868) & (g884) & (!g890) & (!g893)) + ((!g683) & (!g865) & (!g868) & (g884) & (g890) & (!g893)) + ((!g683) & (!g865) & (g868) & (!g884) & (g890) & (!g893)) + ((!g683) & (!g865) & (g868) & (g884) & (!g890) & (!g893)) + ((g683) & (!g865) & (!g868) & (!g884) & (!g890) & (g893)) + ((g683) & (!g865) & (!g868) & (!g884) & (g890) & (g893)) + ((g683) & (!g865) & (!g868) & (g884) & (!g890) & (g893)) + ((g683) & (!g865) & (!g868) & (g884) & (g890) & (g893)) + ((g683) & (!g865) & (g868) & (!g884) & (!g890) & (!g893)) + ((g683) & (!g865) & (g868) & (!g884) & (!g890) & (g893)) + ((g683) & (!g865) & (g868) & (!g884) & (g890) & (g893)) + ((g683) & (!g865) & (g868) & (g884) & (!g890) & (g893)) + ((g683) & (!g865) & (g868) & (g884) & (g890) & (!g893)) + ((g683) & (!g865) & (g868) & (g884) & (g890) & (g893)) + ((g683) & (g865) & (!g868) & (!g884) & (!g890) & (!g893)) + ((g683) & (g865) & (!g868) & (!g884) & (!g890) & (g893)) + ((g683) & (g865) & (!g868) & (!g884) & (g890) & (!g893)) + ((g683) & (g865) & (!g868) & (!g884) & (g890) & (g893)) + ((g683) & (g865) & (!g868) & (g884) & (!g890) & (!g893)) + ((g683) & (g865) & (!g868) & (g884) & (!g890) & (g893)) + ((g683) & (g865) & (!g868) & (g884) & (g890) & (!g893)) + ((g683) & (g865) & (!g868) & (g884) & (g890) & (g893)) + ((g683) & (g865) & (g868) & (!g884) & (!g890) & (!g893)) + ((g683) & (g865) & (g868) & (!g884) & (!g890) & (g893)) + ((g683) & (g865) & (g868) & (!g884) & (g890) & (!g893)) + ((g683) & (g865) & (g868) & (!g884) & (g890) & (g893)) + ((g683) & (g865) & (g868) & (g884) & (!g890) & (!g893)) + ((g683) & (g865) & (g868) & (g884) & (!g890) & (g893)) + ((g683) & (g865) & (g868) & (g884) & (g890) & (!g893)) + ((g683) & (g865) & (g868) & (g884) & (g890) & (g893)));
	assign g895 = (((!g869) & (!g870) & (!g834) & (!g871) & (!g883) & (!g863)) + ((!g869) & (!g870) & (!g834) & (!g871) & (!g883) & (g863)) + ((!g869) & (!g870) & (!g834) & (g871) & (g883) & (!g863)) + ((!g869) & (!g870) & (!g834) & (g871) & (g883) & (g863)) + ((!g869) & (!g870) & (g834) & (!g871) & (!g883) & (g863)) + ((!g869) & (!g870) & (g834) & (!g871) & (g883) & (!g863)) + ((!g869) & (!g870) & (g834) & (g871) & (!g883) & (!g863)) + ((!g869) & (!g870) & (g834) & (g871) & (g883) & (g863)) + ((!g869) & (g870) & (!g834) & (!g871) & (!g883) & (!g863)) + ((!g869) & (g870) & (!g834) & (!g871) & (g883) & (g863)) + ((!g869) & (g870) & (!g834) & (g871) & (!g883) & (g863)) + ((!g869) & (g870) & (!g834) & (g871) & (g883) & (!g863)) + ((!g869) & (g870) & (g834) & (!g871) & (!g883) & (!g863)) + ((!g869) & (g870) & (g834) & (!g871) & (g883) & (g863)) + ((!g869) & (g870) & (g834) & (g871) & (!g883) & (g863)) + ((!g869) & (g870) & (g834) & (g871) & (g883) & (!g863)) + ((g869) & (!g870) & (!g834) & (!g871) & (!g883) & (g863)) + ((g869) & (!g870) & (!g834) & (!g871) & (g883) & (!g863)) + ((g869) & (!g870) & (!g834) & (g871) & (!g883) & (!g863)) + ((g869) & (!g870) & (!g834) & (g871) & (g883) & (g863)) + ((g869) & (!g870) & (g834) & (!g871) & (!g883) & (g863)) + ((g869) & (!g870) & (g834) & (!g871) & (g883) & (!g863)) + ((g869) & (!g870) & (g834) & (g871) & (!g883) & (!g863)) + ((g869) & (!g870) & (g834) & (g871) & (g883) & (g863)) + ((g869) & (g870) & (!g834) & (!g871) & (!g883) & (!g863)) + ((g869) & (g870) & (!g834) & (!g871) & (g883) & (g863)) + ((g869) & (g870) & (!g834) & (g871) & (!g883) & (g863)) + ((g869) & (g870) & (!g834) & (g871) & (g883) & (!g863)) + ((g869) & (g870) & (g834) & (!g871) & (!g883) & (!g863)) + ((g869) & (g870) & (g834) & (!g871) & (!g883) & (g863)) + ((g869) & (g870) & (g834) & (g871) & (g883) & (!g863)) + ((g869) & (g870) & (g834) & (g871) & (g883) & (g863)));
	assign g896 = (((!sk[10]) & (!g870) & (!g891) & (!g871) & (g883) & (!g864)) + ((!sk[10]) & (!g870) & (!g891) & (!g871) & (g883) & (g864)) + ((!sk[10]) & (!g870) & (!g891) & (g871) & (!g883) & (!g864)) + ((!sk[10]) & (!g870) & (!g891) & (g871) & (!g883) & (g864)) + ((!sk[10]) & (!g870) & (!g891) & (g871) & (g883) & (!g864)) + ((!sk[10]) & (!g870) & (!g891) & (g871) & (g883) & (g864)) + ((!sk[10]) & (!g870) & (g891) & (!g871) & (!g883) & (!g864)) + ((!sk[10]) & (!g870) & (g891) & (!g871) & (!g883) & (g864)) + ((!sk[10]) & (!g870) & (g891) & (!g871) & (g883) & (!g864)) + ((!sk[10]) & (!g870) & (g891) & (!g871) & (g883) & (g864)) + ((!sk[10]) & (!g870) & (g891) & (g871) & (!g883) & (!g864)) + ((!sk[10]) & (!g870) & (g891) & (g871) & (!g883) & (g864)) + ((!sk[10]) & (!g870) & (g891) & (g871) & (g883) & (!g864)) + ((!sk[10]) & (!g870) & (g891) & (g871) & (g883) & (g864)) + ((!sk[10]) & (g870) & (!g891) & (!g871) & (g883) & (!g864)) + ((!sk[10]) & (g870) & (!g891) & (!g871) & (g883) & (g864)) + ((!sk[10]) & (g870) & (!g891) & (g871) & (!g883) & (!g864)) + ((!sk[10]) & (g870) & (!g891) & (g871) & (!g883) & (g864)) + ((!sk[10]) & (g870) & (!g891) & (g871) & (g883) & (!g864)) + ((!sk[10]) & (g870) & (!g891) & (g871) & (g883) & (g864)) + ((!sk[10]) & (g870) & (g891) & (!g871) & (!g883) & (!g864)) + ((!sk[10]) & (g870) & (g891) & (!g871) & (!g883) & (g864)) + ((!sk[10]) & (g870) & (g891) & (!g871) & (g883) & (!g864)) + ((!sk[10]) & (g870) & (g891) & (!g871) & (g883) & (g864)) + ((!sk[10]) & (g870) & (g891) & (g871) & (!g883) & (!g864)) + ((!sk[10]) & (g870) & (g891) & (g871) & (!g883) & (g864)) + ((!sk[10]) & (g870) & (g891) & (g871) & (g883) & (!g864)) + ((!sk[10]) & (g870) & (g891) & (g871) & (g883) & (g864)) + ((sk[10]) & (!g870) & (!g891) & (!g871) & (!g883) & (g864)) + ((sk[10]) & (!g870) & (!g891) & (!g871) & (g883) & (g864)) + ((sk[10]) & (!g870) & (!g891) & (g871) & (!g883) & (g864)) + ((sk[10]) & (!g870) & (!g891) & (g871) & (g883) & (g864)) + ((sk[10]) & (!g870) & (g891) & (!g871) & (!g883) & (!g864)) + ((sk[10]) & (!g870) & (g891) & (!g871) & (!g883) & (g864)) + ((sk[10]) & (!g870) & (g891) & (!g871) & (g883) & (g864)) + ((sk[10]) & (!g870) & (g891) & (g871) & (!g883) & (g864)) + ((sk[10]) & (!g870) & (g891) & (g871) & (g883) & (!g864)) + ((sk[10]) & (!g870) & (g891) & (g871) & (g883) & (g864)) + ((sk[10]) & (g870) & (g891) & (!g871) & (!g883) & (!g864)) + ((sk[10]) & (g870) & (g891) & (!g871) & (!g883) & (g864)) + ((sk[10]) & (g870) & (g891) & (g871) & (g883) & (!g864)) + ((sk[10]) & (g870) & (g891) & (g871) & (g883) & (g864)));
	assign g897 = (((!sk[11]) & (!g863) & (!g892) & (!g868) & (g895) & (!g896)) + ((!sk[11]) & (!g863) & (!g892) & (!g868) & (g895) & (g896)) + ((!sk[11]) & (!g863) & (!g892) & (g868) & (!g895) & (!g896)) + ((!sk[11]) & (!g863) & (!g892) & (g868) & (!g895) & (g896)) + ((!sk[11]) & (!g863) & (!g892) & (g868) & (g895) & (!g896)) + ((!sk[11]) & (!g863) & (!g892) & (g868) & (g895) & (g896)) + ((!sk[11]) & (!g863) & (g892) & (!g868) & (!g895) & (!g896)) + ((!sk[11]) & (!g863) & (g892) & (!g868) & (!g895) & (g896)) + ((!sk[11]) & (!g863) & (g892) & (!g868) & (g895) & (!g896)) + ((!sk[11]) & (!g863) & (g892) & (!g868) & (g895) & (g896)) + ((!sk[11]) & (!g863) & (g892) & (g868) & (!g895) & (!g896)) + ((!sk[11]) & (!g863) & (g892) & (g868) & (!g895) & (g896)) + ((!sk[11]) & (!g863) & (g892) & (g868) & (g895) & (!g896)) + ((!sk[11]) & (!g863) & (g892) & (g868) & (g895) & (g896)) + ((!sk[11]) & (g863) & (!g892) & (!g868) & (g895) & (!g896)) + ((!sk[11]) & (g863) & (!g892) & (!g868) & (g895) & (g896)) + ((!sk[11]) & (g863) & (!g892) & (g868) & (!g895) & (!g896)) + ((!sk[11]) & (g863) & (!g892) & (g868) & (!g895) & (g896)) + ((!sk[11]) & (g863) & (!g892) & (g868) & (g895) & (!g896)) + ((!sk[11]) & (g863) & (!g892) & (g868) & (g895) & (g896)) + ((!sk[11]) & (g863) & (g892) & (!g868) & (!g895) & (!g896)) + ((!sk[11]) & (g863) & (g892) & (!g868) & (!g895) & (g896)) + ((!sk[11]) & (g863) & (g892) & (!g868) & (g895) & (!g896)) + ((!sk[11]) & (g863) & (g892) & (!g868) & (g895) & (g896)) + ((!sk[11]) & (g863) & (g892) & (g868) & (!g895) & (!g896)) + ((!sk[11]) & (g863) & (g892) & (g868) & (!g895) & (g896)) + ((!sk[11]) & (g863) & (g892) & (g868) & (g895) & (!g896)) + ((!sk[11]) & (g863) & (g892) & (g868) & (g895) & (g896)) + ((sk[11]) & (!g863) & (!g892) & (!g868) & (!g895) & (!g896)) + ((sk[11]) & (!g863) & (!g892) & (!g868) & (g895) & (!g896)) + ((sk[11]) & (!g863) & (!g892) & (g868) & (!g895) & (!g896)) + ((sk[11]) & (!g863) & (g892) & (!g868) & (!g895) & (!g896)) + ((sk[11]) & (!g863) & (g892) & (!g868) & (g895) & (!g896)) + ((sk[11]) & (!g863) & (g892) & (g868) & (!g895) & (!g896)) + ((sk[11]) & (g863) & (!g892) & (!g868) & (!g895) & (!g896)) + ((sk[11]) & (g863) & (!g892) & (!g868) & (g895) & (!g896)) + ((sk[11]) & (g863) & (!g892) & (g868) & (!g895) & (!g896)));
	assign g898 = (((!g789) & (!g790) & (!g793) & (!g815) & (!g819) & (g820)) + ((!g789) & (!g790) & (!g793) & (!g815) & (g819) & (!g820)) + ((!g789) & (!g790) & (!g793) & (g815) & (!g819) & (!g820)) + ((!g789) & (!g790) & (!g793) & (g815) & (g819) & (g820)) + ((!g789) & (!g790) & (g793) & (!g815) & (!g819) & (g820)) + ((!g789) & (!g790) & (g793) & (!g815) & (g819) & (!g820)) + ((!g789) & (!g790) & (g793) & (g815) & (!g819) & (g820)) + ((!g789) & (!g790) & (g793) & (g815) & (g819) & (!g820)) + ((!g789) & (g790) & (!g793) & (!g815) & (!g819) & (!g820)) + ((!g789) & (g790) & (!g793) & (!g815) & (g819) & (g820)) + ((!g789) & (g790) & (!g793) & (g815) & (!g819) & (!g820)) + ((!g789) & (g790) & (!g793) & (g815) & (g819) & (g820)) + ((!g789) & (g790) & (g793) & (!g815) & (!g819) & (g820)) + ((!g789) & (g790) & (g793) & (!g815) & (g819) & (!g820)) + ((!g789) & (g790) & (g793) & (g815) & (!g819) & (!g820)) + ((!g789) & (g790) & (g793) & (g815) & (g819) & (g820)) + ((g789) & (!g790) & (!g793) & (!g815) & (!g819) & (!g820)) + ((g789) & (!g790) & (!g793) & (!g815) & (g819) & (g820)) + ((g789) & (!g790) & (!g793) & (g815) & (!g819) & (!g820)) + ((g789) & (!g790) & (!g793) & (g815) & (g819) & (g820)) + ((g789) & (!g790) & (g793) & (!g815) & (!g819) & (g820)) + ((g789) & (!g790) & (g793) & (!g815) & (g819) & (!g820)) + ((g789) & (!g790) & (g793) & (g815) & (!g819) & (!g820)) + ((g789) & (!g790) & (g793) & (g815) & (g819) & (g820)) + ((g789) & (g790) & (!g793) & (!g815) & (!g819) & (g820)) + ((g789) & (g790) & (!g793) & (!g815) & (g819) & (!g820)) + ((g789) & (g790) & (!g793) & (g815) & (!g819) & (!g820)) + ((g789) & (g790) & (!g793) & (g815) & (g819) & (g820)) + ((g789) & (g790) & (g793) & (!g815) & (!g819) & (g820)) + ((g789) & (g790) & (g793) & (!g815) & (g819) & (!g820)) + ((g789) & (g790) & (g793) & (g815) & (!g819) & (g820)) + ((g789) & (g790) & (g793) & (g815) & (g819) & (!g820)));
	assign g899 = (((!g869) & (!g870) & (!g834) & (!sk[13]) & (g863)) + ((!g869) & (!g870) & (!g834) & (sk[13]) & (g863)) + ((!g869) & (!g870) & (g834) & (!sk[13]) & (g863)) + ((!g869) & (!g870) & (g834) & (sk[13]) & (!g863)) + ((!g869) & (g870) & (!g834) & (!sk[13]) & (g863)) + ((!g869) & (g870) & (!g834) & (sk[13]) & (!g863)) + ((!g869) & (g870) & (g834) & (!sk[13]) & (g863)) + ((!g869) & (g870) & (g834) & (sk[13]) & (!g863)) + ((g869) & (!g870) & (!g834) & (!sk[13]) & (!g863)) + ((g869) & (!g870) & (!g834) & (!sk[13]) & (g863)) + ((g869) & (!g870) & (!g834) & (sk[13]) & (!g863)) + ((g869) & (!g870) & (g834) & (!sk[13]) & (!g863)) + ((g869) & (!g870) & (g834) & (!sk[13]) & (g863)) + ((g869) & (!g870) & (g834) & (sk[13]) & (!g863)) + ((g869) & (g870) & (!g834) & (!sk[13]) & (!g863)) + ((g869) & (g870) & (!g834) & (!sk[13]) & (g863)) + ((g869) & (g870) & (!g834) & (sk[13]) & (!g863)) + ((g869) & (g870) & (g834) & (!sk[13]) & (!g863)) + ((g869) & (g870) & (g834) & (!sk[13]) & (g863)) + ((g869) & (g870) & (g834) & (sk[13]) & (g863)));
	assign g900 = (((!sk[14]) & (!g870) & (!g891) & (!g863) & (g892)) + ((!sk[14]) & (!g870) & (!g891) & (g863) & (g892)) + ((!sk[14]) & (!g870) & (g891) & (!g863) & (g892)) + ((!sk[14]) & (!g870) & (g891) & (g863) & (g892)) + ((!sk[14]) & (g870) & (!g891) & (!g863) & (!g892)) + ((!sk[14]) & (g870) & (!g891) & (!g863) & (g892)) + ((!sk[14]) & (g870) & (!g891) & (g863) & (!g892)) + ((!sk[14]) & (g870) & (!g891) & (g863) & (g892)) + ((!sk[14]) & (g870) & (g891) & (!g863) & (!g892)) + ((!sk[14]) & (g870) & (g891) & (!g863) & (g892)) + ((!sk[14]) & (g870) & (g891) & (g863) & (!g892)) + ((!sk[14]) & (g870) & (g891) & (g863) & (g892)) + ((sk[14]) & (!g870) & (!g891) & (!g863) & (g892)) + ((sk[14]) & (!g870) & (!g891) & (g863) & (g892)) + ((sk[14]) & (!g870) & (g891) & (!g863) & (g892)) + ((sk[14]) & (!g870) & (g891) & (g863) & (!g892)) + ((sk[14]) & (!g870) & (g891) & (g863) & (g892)) + ((sk[14]) & (g870) & (g891) & (g863) & (!g892)) + ((sk[14]) & (g870) & (g891) & (g863) & (g892)));
	assign g901 = (((!sk[15]) & (!g869) & (!g864) & (!g868) & (g899) & (!g900)) + ((!sk[15]) & (!g869) & (!g864) & (!g868) & (g899) & (g900)) + ((!sk[15]) & (!g869) & (!g864) & (g868) & (!g899) & (!g900)) + ((!sk[15]) & (!g869) & (!g864) & (g868) & (!g899) & (g900)) + ((!sk[15]) & (!g869) & (!g864) & (g868) & (g899) & (!g900)) + ((!sk[15]) & (!g869) & (!g864) & (g868) & (g899) & (g900)) + ((!sk[15]) & (!g869) & (g864) & (!g868) & (!g899) & (!g900)) + ((!sk[15]) & (!g869) & (g864) & (!g868) & (!g899) & (g900)) + ((!sk[15]) & (!g869) & (g864) & (!g868) & (g899) & (!g900)) + ((!sk[15]) & (!g869) & (g864) & (!g868) & (g899) & (g900)) + ((!sk[15]) & (!g869) & (g864) & (g868) & (!g899) & (!g900)) + ((!sk[15]) & (!g869) & (g864) & (g868) & (!g899) & (g900)) + ((!sk[15]) & (!g869) & (g864) & (g868) & (g899) & (!g900)) + ((!sk[15]) & (!g869) & (g864) & (g868) & (g899) & (g900)) + ((!sk[15]) & (g869) & (!g864) & (!g868) & (g899) & (!g900)) + ((!sk[15]) & (g869) & (!g864) & (!g868) & (g899) & (g900)) + ((!sk[15]) & (g869) & (!g864) & (g868) & (!g899) & (!g900)) + ((!sk[15]) & (g869) & (!g864) & (g868) & (!g899) & (g900)) + ((!sk[15]) & (g869) & (!g864) & (g868) & (g899) & (!g900)) + ((!sk[15]) & (g869) & (!g864) & (g868) & (g899) & (g900)) + ((!sk[15]) & (g869) & (g864) & (!g868) & (!g899) & (!g900)) + ((!sk[15]) & (g869) & (g864) & (!g868) & (!g899) & (g900)) + ((!sk[15]) & (g869) & (g864) & (!g868) & (g899) & (!g900)) + ((!sk[15]) & (g869) & (g864) & (!g868) & (g899) & (g900)) + ((!sk[15]) & (g869) & (g864) & (g868) & (!g899) & (!g900)) + ((!sk[15]) & (g869) & (g864) & (g868) & (!g899) & (g900)) + ((!sk[15]) & (g869) & (g864) & (g868) & (g899) & (!g900)) + ((!sk[15]) & (g869) & (g864) & (g868) & (g899) & (g900)) + ((sk[15]) & (!g869) & (!g864) & (!g868) & (!g899) & (!g900)) + ((sk[15]) & (!g869) & (!g864) & (!g868) & (g899) & (!g900)) + ((sk[15]) & (!g869) & (!g864) & (g868) & (g899) & (!g900)) + ((sk[15]) & (!g869) & (g864) & (!g868) & (!g899) & (!g900)) + ((sk[15]) & (!g869) & (g864) & (!g868) & (g899) & (!g900)) + ((sk[15]) & (!g869) & (g864) & (g868) & (g899) & (!g900)) + ((sk[15]) & (g869) & (!g864) & (!g868) & (!g899) & (!g900)) + ((sk[15]) & (g869) & (!g864) & (!g868) & (g899) & (!g900)) + ((sk[15]) & (g869) & (!g864) & (g868) & (g899) & (!g900)));
	assign g902 = (((!g789) & (!g790) & (!sk[16]) & (!g793) & (g815)) + ((!g789) & (!g790) & (!sk[16]) & (g793) & (g815)) + ((!g789) & (!g790) & (sk[16]) & (!g793) & (g815)) + ((!g789) & (!g790) & (sk[16]) & (g793) & (!g815)) + ((!g789) & (g790) & (!sk[16]) & (!g793) & (g815)) + ((!g789) & (g790) & (!sk[16]) & (g793) & (g815)) + ((!g789) & (g790) & (sk[16]) & (!g793) & (!g815)) + ((!g789) & (g790) & (sk[16]) & (g793) & (g815)) + ((g789) & (!g790) & (!sk[16]) & (!g793) & (!g815)) + ((g789) & (!g790) & (!sk[16]) & (!g793) & (g815)) + ((g789) & (!g790) & (!sk[16]) & (g793) & (!g815)) + ((g789) & (!g790) & (!sk[16]) & (g793) & (g815)) + ((g789) & (!g790) & (sk[16]) & (!g793) & (!g815)) + ((g789) & (!g790) & (sk[16]) & (g793) & (g815)) + ((g789) & (g790) & (!sk[16]) & (!g793) & (!g815)) + ((g789) & (g790) & (!sk[16]) & (!g793) & (g815)) + ((g789) & (g790) & (!sk[16]) & (g793) & (!g815)) + ((g789) & (g790) & (!sk[16]) & (g793) & (g815)) + ((g789) & (g790) & (sk[16]) & (!g793) & (g815)) + ((g789) & (g790) & (sk[16]) & (g793) & (!g815)));
	assign g903 = (((!g707) & (!g717) & (!g718) & (!sk[17]) & (g864) & (!g892)) + ((!g707) & (!g717) & (!g718) & (!sk[17]) & (g864) & (g892)) + ((!g707) & (!g717) & (g718) & (!sk[17]) & (!g864) & (!g892)) + ((!g707) & (!g717) & (g718) & (!sk[17]) & (!g864) & (g892)) + ((!g707) & (!g717) & (g718) & (!sk[17]) & (g864) & (!g892)) + ((!g707) & (!g717) & (g718) & (!sk[17]) & (g864) & (g892)) + ((!g707) & (!g717) & (g718) & (sk[17]) & (g864) & (!g892)) + ((!g707) & (!g717) & (g718) & (sk[17]) & (g864) & (g892)) + ((!g707) & (g717) & (!g718) & (!sk[17]) & (!g864) & (!g892)) + ((!g707) & (g717) & (!g718) & (!sk[17]) & (!g864) & (g892)) + ((!g707) & (g717) & (!g718) & (!sk[17]) & (g864) & (!g892)) + ((!g707) & (g717) & (!g718) & (!sk[17]) & (g864) & (g892)) + ((!g707) & (g717) & (!g718) & (sk[17]) & (!g864) & (g892)) + ((!g707) & (g717) & (!g718) & (sk[17]) & (g864) & (g892)) + ((!g707) & (g717) & (g718) & (!sk[17]) & (!g864) & (!g892)) + ((!g707) & (g717) & (g718) & (!sk[17]) & (!g864) & (g892)) + ((!g707) & (g717) & (g718) & (!sk[17]) & (g864) & (!g892)) + ((!g707) & (g717) & (g718) & (!sk[17]) & (g864) & (g892)) + ((!g707) & (g717) & (g718) & (sk[17]) & (!g864) & (g892)) + ((!g707) & (g717) & (g718) & (sk[17]) & (g864) & (!g892)) + ((!g707) & (g717) & (g718) & (sk[17]) & (g864) & (g892)) + ((g707) & (!g717) & (!g718) & (!sk[17]) & (g864) & (!g892)) + ((g707) & (!g717) & (!g718) & (!sk[17]) & (g864) & (g892)) + ((g707) & (!g717) & (!g718) & (sk[17]) & (!g864) & (g892)) + ((g707) & (!g717) & (!g718) & (sk[17]) & (g864) & (g892)) + ((g707) & (!g717) & (g718) & (!sk[17]) & (!g864) & (!g892)) + ((g707) & (!g717) & (g718) & (!sk[17]) & (!g864) & (g892)) + ((g707) & (!g717) & (g718) & (!sk[17]) & (g864) & (!g892)) + ((g707) & (!g717) & (g718) & (!sk[17]) & (g864) & (g892)) + ((g707) & (!g717) & (g718) & (sk[17]) & (!g864) & (g892)) + ((g707) & (!g717) & (g718) & (sk[17]) & (g864) & (!g892)) + ((g707) & (!g717) & (g718) & (sk[17]) & (g864) & (g892)) + ((g707) & (g717) & (!g718) & (!sk[17]) & (!g864) & (!g892)) + ((g707) & (g717) & (!g718) & (!sk[17]) & (!g864) & (g892)) + ((g707) & (g717) & (!g718) & (!sk[17]) & (g864) & (!g892)) + ((g707) & (g717) & (!g718) & (!sk[17]) & (g864) & (g892)) + ((g707) & (g717) & (g718) & (!sk[17]) & (!g864) & (!g892)) + ((g707) & (g717) & (g718) & (!sk[17]) & (!g864) & (g892)) + ((g707) & (g717) & (g718) & (!sk[17]) & (g864) & (!g892)) + ((g707) & (g717) & (g718) & (!sk[17]) & (g864) & (g892)) + ((g707) & (g717) & (g718) & (sk[17]) & (g864) & (!g892)) + ((g707) & (g717) & (g718) & (sk[17]) & (g864) & (g892)));
	assign g904 = (((!ax0x) & (!g869) & (!g870) & (!g834) & (!g867) & (!g903)) + ((!ax0x) & (!g869) & (!g870) & (!g834) & (g867) & (!g903)) + ((!ax0x) & (!g869) & (!g870) & (g834) & (!g867) & (!g903)) + ((!ax0x) & (!g869) & (!g870) & (g834) & (g867) & (!g903)) + ((!ax0x) & (!g869) & (g870) & (!g834) & (!g867) & (!g903)) + ((!ax0x) & (!g869) & (g870) & (!g834) & (g867) & (!g903)) + ((!ax0x) & (!g869) & (g870) & (g834) & (!g867) & (!g903)) + ((!ax0x) & (!g869) & (g870) & (g834) & (g867) & (!g903)) + ((!ax0x) & (g869) & (!g870) & (!g834) & (!g867) & (!g903)) + ((!ax0x) & (g869) & (!g870) & (!g834) & (g867) & (!g903)) + ((!ax0x) & (g869) & (!g870) & (g834) & (!g867) & (!g903)) + ((!ax0x) & (g869) & (!g870) & (g834) & (g867) & (!g903)) + ((!ax0x) & (g869) & (g870) & (!g834) & (!g867) & (!g903)) + ((!ax0x) & (g869) & (g870) & (!g834) & (g867) & (!g903)) + ((!ax0x) & (g869) & (g870) & (g834) & (!g867) & (!g903)) + ((!ax0x) & (g869) & (g870) & (g834) & (g867) & (!g903)) + ((ax0x) & (!g869) & (!g870) & (g834) & (g867) & (!g903)) + ((ax0x) & (!g869) & (g870) & (!g834) & (!g867) & (!g903)) + ((ax0x) & (!g869) & (g870) & (!g834) & (g867) & (!g903)) + ((ax0x) & (!g869) & (g870) & (g834) & (!g867) & (!g903)) + ((ax0x) & (g869) & (!g870) & (!g834) & (g867) & (!g903)) + ((ax0x) & (g869) & (g870) & (!g834) & (!g867) & (!g903)) + ((ax0x) & (g869) & (g870) & (g834) & (!g867) & (!g903)) + ((ax0x) & (g869) & (g870) & (g834) & (g867) & (!g903)));
	assign g905 = (((!g2) & (!g808) & (!g810) & (!g811) & (!g813) & (g814)) + ((!g2) & (!g808) & (!g810) & (!g811) & (g813) & (!g814)) + ((!g2) & (!g808) & (!g810) & (g811) & (!g813) & (!g814)) + ((!g2) & (!g808) & (!g810) & (g811) & (g813) & (g814)) + ((!g2) & (!g808) & (g810) & (!g811) & (!g813) & (!g814)) + ((!g2) & (!g808) & (g810) & (!g811) & (g813) & (g814)) + ((!g2) & (!g808) & (g810) & (g811) & (!g813) & (!g814)) + ((!g2) & (!g808) & (g810) & (g811) & (g813) & (g814)) + ((!g2) & (g808) & (!g810) & (!g811) & (!g813) & (g814)) + ((!g2) & (g808) & (!g810) & (!g811) & (g813) & (!g814)) + ((!g2) & (g808) & (!g810) & (g811) & (!g813) & (g814)) + ((!g2) & (g808) & (!g810) & (g811) & (g813) & (!g814)) + ((!g2) & (g808) & (g810) & (!g811) & (!g813) & (g814)) + ((!g2) & (g808) & (g810) & (!g811) & (g813) & (!g814)) + ((!g2) & (g808) & (g810) & (g811) & (!g813) & (!g814)) + ((!g2) & (g808) & (g810) & (g811) & (g813) & (g814)) + ((g2) & (!g808) & (!g810) & (!g811) & (!g813) & (!g814)) + ((g2) & (!g808) & (!g810) & (!g811) & (g813) & (g814)) + ((g2) & (!g808) & (!g810) & (g811) & (!g813) & (g814)) + ((g2) & (!g808) & (!g810) & (g811) & (g813) & (!g814)) + ((g2) & (!g808) & (g810) & (!g811) & (!g813) & (g814)) + ((g2) & (!g808) & (g810) & (!g811) & (g813) & (!g814)) + ((g2) & (!g808) & (g810) & (g811) & (!g813) & (g814)) + ((g2) & (!g808) & (g810) & (g811) & (g813) & (!g814)) + ((g2) & (g808) & (!g810) & (!g811) & (!g813) & (!g814)) + ((g2) & (g808) & (!g810) & (!g811) & (g813) & (g814)) + ((g2) & (g808) & (!g810) & (g811) & (!g813) & (!g814)) + ((g2) & (g808) & (!g810) & (g811) & (g813) & (g814)) + ((g2) & (g808) & (g810) & (!g811) & (!g813) & (!g814)) + ((g2) & (g808) & (g810) & (!g811) & (g813) & (g814)) + ((g2) & (g808) & (g810) & (g811) & (!g813) & (g814)) + ((g2) & (g808) & (g810) & (g811) & (g813) & (!g814)));
	assign g906 = (((!g549) & (!g569) & (!sk[20]) & (!g680) & (g864)) + ((!g549) & (!g569) & (!sk[20]) & (g680) & (g864)) + ((!g549) & (!g569) & (sk[20]) & (g680) & (g864)) + ((!g549) & (g569) & (!sk[20]) & (!g680) & (g864)) + ((!g549) & (g569) & (!sk[20]) & (g680) & (g864)) + ((!g549) & (g569) & (sk[20]) & (!g680) & (g864)) + ((g549) & (!g569) & (!sk[20]) & (!g680) & (!g864)) + ((g549) & (!g569) & (!sk[20]) & (!g680) & (g864)) + ((g549) & (!g569) & (!sk[20]) & (g680) & (!g864)) + ((g549) & (!g569) & (!sk[20]) & (g680) & (g864)) + ((g549) & (!g569) & (sk[20]) & (!g680) & (g864)) + ((g549) & (g569) & (!sk[20]) & (!g680) & (!g864)) + ((g549) & (g569) & (!sk[20]) & (!g680) & (g864)) + ((g549) & (g569) & (!sk[20]) & (g680) & (!g864)) + ((g549) & (g569) & (!sk[20]) & (g680) & (g864)) + ((g549) & (g569) & (sk[20]) & (g680) & (g864)));
	assign g907 = (((!g707) & (!g717) & (!g718) & (g891) & (!sk[21]) & (!g892)) + ((!g707) & (!g717) & (!g718) & (g891) & (!sk[21]) & (g892)) + ((!g707) & (!g717) & (g718) & (!g891) & (!sk[21]) & (!g892)) + ((!g707) & (!g717) & (g718) & (!g891) & (!sk[21]) & (g892)) + ((!g707) & (!g717) & (g718) & (!g891) & (sk[21]) & (g892)) + ((!g707) & (!g717) & (g718) & (g891) & (!sk[21]) & (!g892)) + ((!g707) & (!g717) & (g718) & (g891) & (!sk[21]) & (g892)) + ((!g707) & (!g717) & (g718) & (g891) & (sk[21]) & (g892)) + ((!g707) & (g717) & (!g718) & (!g891) & (!sk[21]) & (!g892)) + ((!g707) & (g717) & (!g718) & (!g891) & (!sk[21]) & (g892)) + ((!g707) & (g717) & (!g718) & (g891) & (!sk[21]) & (!g892)) + ((!g707) & (g717) & (!g718) & (g891) & (!sk[21]) & (g892)) + ((!g707) & (g717) & (!g718) & (g891) & (sk[21]) & (!g892)) + ((!g707) & (g717) & (!g718) & (g891) & (sk[21]) & (g892)) + ((!g707) & (g717) & (g718) & (!g891) & (!sk[21]) & (!g892)) + ((!g707) & (g717) & (g718) & (!g891) & (!sk[21]) & (g892)) + ((!g707) & (g717) & (g718) & (!g891) & (sk[21]) & (g892)) + ((!g707) & (g717) & (g718) & (g891) & (!sk[21]) & (!g892)) + ((!g707) & (g717) & (g718) & (g891) & (!sk[21]) & (g892)) + ((!g707) & (g717) & (g718) & (g891) & (sk[21]) & (!g892)) + ((!g707) & (g717) & (g718) & (g891) & (sk[21]) & (g892)) + ((g707) & (!g717) & (!g718) & (g891) & (!sk[21]) & (!g892)) + ((g707) & (!g717) & (!g718) & (g891) & (!sk[21]) & (g892)) + ((g707) & (!g717) & (!g718) & (g891) & (sk[21]) & (!g892)) + ((g707) & (!g717) & (!g718) & (g891) & (sk[21]) & (g892)) + ((g707) & (!g717) & (g718) & (!g891) & (!sk[21]) & (!g892)) + ((g707) & (!g717) & (g718) & (!g891) & (!sk[21]) & (g892)) + ((g707) & (!g717) & (g718) & (!g891) & (sk[21]) & (g892)) + ((g707) & (!g717) & (g718) & (g891) & (!sk[21]) & (!g892)) + ((g707) & (!g717) & (g718) & (g891) & (!sk[21]) & (g892)) + ((g707) & (!g717) & (g718) & (g891) & (sk[21]) & (!g892)) + ((g707) & (!g717) & (g718) & (g891) & (sk[21]) & (g892)) + ((g707) & (g717) & (!g718) & (!g891) & (!sk[21]) & (!g892)) + ((g707) & (g717) & (!g718) & (!g891) & (!sk[21]) & (g892)) + ((g707) & (g717) & (!g718) & (g891) & (!sk[21]) & (!g892)) + ((g707) & (g717) & (!g718) & (g891) & (!sk[21]) & (g892)) + ((g707) & (g717) & (g718) & (!g891) & (!sk[21]) & (!g892)) + ((g707) & (g717) & (g718) & (!g891) & (!sk[21]) & (g892)) + ((g707) & (g717) & (g718) & (!g891) & (sk[21]) & (g892)) + ((g707) & (g717) & (g718) & (g891) & (!sk[21]) & (!g892)) + ((g707) & (g717) & (g718) & (g891) & (!sk[21]) & (g892)) + ((g707) & (g717) & (g718) & (g891) & (sk[21]) & (g892)));
	assign g908 = (((!ax0x) & (!g683) & (!g731) & (!g866) & (!g906) & (g907)) + ((!ax0x) & (!g683) & (!g731) & (!g866) & (g906) & (!g907)) + ((!ax0x) & (!g683) & (!g731) & (!g866) & (g906) & (g907)) + ((!ax0x) & (!g683) & (!g731) & (g866) & (!g906) & (g907)) + ((!ax0x) & (!g683) & (!g731) & (g866) & (g906) & (!g907)) + ((!ax0x) & (!g683) & (!g731) & (g866) & (g906) & (g907)) + ((!ax0x) & (!g683) & (g731) & (!g866) & (!g906) & (g907)) + ((!ax0x) & (!g683) & (g731) & (!g866) & (g906) & (!g907)) + ((!ax0x) & (!g683) & (g731) & (!g866) & (g906) & (g907)) + ((!ax0x) & (!g683) & (g731) & (g866) & (!g906) & (g907)) + ((!ax0x) & (!g683) & (g731) & (g866) & (g906) & (!g907)) + ((!ax0x) & (!g683) & (g731) & (g866) & (g906) & (g907)) + ((!ax0x) & (g683) & (!g731) & (!g866) & (!g906) & (!g907)) + ((!ax0x) & (g683) & (!g731) & (g866) & (!g906) & (!g907)) + ((!ax0x) & (g683) & (g731) & (!g866) & (!g906) & (!g907)) + ((!ax0x) & (g683) & (g731) & (g866) & (!g906) & (!g907)) + ((ax0x) & (!g683) & (!g731) & (!g866) & (!g906) & (g907)) + ((ax0x) & (!g683) & (!g731) & (!g866) & (g906) & (!g907)) + ((ax0x) & (!g683) & (!g731) & (!g866) & (g906) & (g907)) + ((ax0x) & (!g683) & (!g731) & (g866) & (!g906) & (g907)) + ((ax0x) & (!g683) & (!g731) & (g866) & (g906) & (!g907)) + ((ax0x) & (!g683) & (!g731) & (g866) & (g906) & (g907)) + ((ax0x) & (!g683) & (g731) & (!g866) & (!g906) & (g907)) + ((ax0x) & (!g683) & (g731) & (!g866) & (g906) & (!g907)) + ((ax0x) & (!g683) & (g731) & (!g866) & (g906) & (g907)) + ((ax0x) & (!g683) & (g731) & (g866) & (!g906) & (!g907)) + ((ax0x) & (!g683) & (g731) & (g866) & (!g906) & (g907)) + ((ax0x) & (!g683) & (g731) & (g866) & (g906) & (!g907)) + ((ax0x) & (!g683) & (g731) & (g866) & (g906) & (g907)) + ((ax0x) & (g683) & (!g731) & (!g866) & (!g906) & (!g907)) + ((ax0x) & (g683) & (!g731) & (g866) & (!g906) & (!g907)) + ((ax0x) & (g683) & (g731) & (g866) & (!g906) & (!g907)));
	assign g909 = (((!sk[23]) & (!g808) & (g810) & (!g811)) + ((!sk[23]) & (!g808) & (g810) & (g811)) + ((!sk[23]) & (g808) & (g810) & (!g811)) + ((!sk[23]) & (g808) & (g810) & (g811)) + ((sk[23]) & (!g808) & (!g810) & (g811)) + ((sk[23]) & (!g808) & (g810) & (!g811)) + ((sk[23]) & (g808) & (!g810) & (!g811)) + ((sk[23]) & (g808) & (g810) & (g811)));
	assign g910 = (((!g708) & (!g716) & (!g549) & (!g569) & (!g680) & (g891)) + ((!g708) & (!g716) & (g549) & (!g569) & (!g680) & (g891)) + ((!g708) & (!g716) & (g549) & (!g569) & (g680) & (g891)) + ((!g708) & (!g716) & (g549) & (g569) & (!g680) & (g891)) + ((!g708) & (g716) & (!g549) & (!g569) & (g680) & (g891)) + ((!g708) & (g716) & (!g549) & (g569) & (!g680) & (g891)) + ((!g708) & (g716) & (!g549) & (g569) & (g680) & (g891)) + ((!g708) & (g716) & (g549) & (g569) & (g680) & (g891)) + ((g708) & (!g716) & (!g549) & (!g569) & (g680) & (g891)) + ((g708) & (!g716) & (!g549) & (g569) & (!g680) & (g891)) + ((g708) & (!g716) & (!g549) & (g569) & (g680) & (g891)) + ((g708) & (!g716) & (g549) & (g569) & (g680) & (g891)) + ((g708) & (g716) & (!g549) & (!g569) & (!g680) & (g891)) + ((g708) & (g716) & (g549) & (!g569) & (!g680) & (g891)) + ((g708) & (g716) & (g549) & (!g569) & (g680) & (g891)) + ((g708) & (g716) & (g549) & (g569) & (!g680) & (g891)));
	assign g911 = (((!g549) & (!g569) & (!g680) & (!g729) & (g864) & (!g892)) + ((!g549) & (!g569) & (!g680) & (!g729) & (g864) & (g892)) + ((!g549) & (!g569) & (g680) & (!g729) & (!g864) & (g892)) + ((!g549) & (!g569) & (g680) & (!g729) & (g864) & (!g892)) + ((!g549) & (!g569) & (g680) & (!g729) & (g864) & (g892)) + ((!g549) & (!g569) & (g680) & (g729) & (!g864) & (g892)) + ((!g549) & (!g569) & (g680) & (g729) & (g864) & (g892)) + ((!g549) & (g569) & (!g680) & (!g729) & (!g864) & (g892)) + ((!g549) & (g569) & (!g680) & (!g729) & (g864) & (!g892)) + ((!g549) & (g569) & (!g680) & (!g729) & (g864) & (g892)) + ((!g549) & (g569) & (!g680) & (g729) & (!g864) & (g892)) + ((!g549) & (g569) & (!g680) & (g729) & (g864) & (g892)) + ((!g549) & (g569) & (g680) & (!g729) & (g864) & (!g892)) + ((!g549) & (g569) & (g680) & (!g729) & (g864) & (g892)) + ((g549) & (!g569) & (!g680) & (!g729) & (!g864) & (g892)) + ((g549) & (!g569) & (!g680) & (!g729) & (g864) & (!g892)) + ((g549) & (!g569) & (!g680) & (!g729) & (g864) & (g892)) + ((g549) & (!g569) & (!g680) & (g729) & (!g864) & (g892)) + ((g549) & (!g569) & (!g680) & (g729) & (g864) & (g892)) + ((g549) & (!g569) & (g680) & (!g729) & (g864) & (!g892)) + ((g549) & (!g569) & (g680) & (!g729) & (g864) & (g892)) + ((g549) & (g569) & (!g680) & (!g729) & (g864) & (!g892)) + ((g549) & (g569) & (!g680) & (!g729) & (g864) & (g892)) + ((g549) & (g569) & (g680) & (!g729) & (!g864) & (g892)) + ((g549) & (g569) & (g680) & (!g729) & (g864) & (!g892)) + ((g549) & (g569) & (g680) & (!g729) & (g864) & (g892)) + ((g549) & (g569) & (g680) & (g729) & (!g864) & (g892)) + ((g549) & (g569) & (g680) & (g729) & (g864) & (g892)));
	assign g912 = (((!ax0x) & (g683) & (!g730) & (!g816) & (!g910) & (!g911)) + ((!ax0x) & (g683) & (!g730) & (g816) & (!g910) & (!g911)) + ((!ax0x) & (g683) & (g730) & (!g816) & (!g910) & (!g911)) + ((!ax0x) & (g683) & (g730) & (g816) & (!g910) & (!g911)) + ((ax0x) & (g683) & (!g730) & (g816) & (!g910) & (!g911)) + ((ax0x) & (g683) & (g730) & (!g816) & (!g910) & (!g911)));
	assign g913 = (((ax0x) & (!sk[27]) & (g866)) + ((ax0x) & (sk[27]) & (g866)));
	assign g914 = (((!g683) & (!g730) & (!g816) & (!g913) & (!g910) & (g911)) + ((!g683) & (!g730) & (!g816) & (!g913) & (g910) & (!g911)) + ((!g683) & (!g730) & (!g816) & (!g913) & (g910) & (g911)) + ((!g683) & (!g730) & (!g816) & (g913) & (!g910) & (!g911)) + ((!g683) & (!g730) & (!g816) & (g913) & (!g910) & (g911)) + ((!g683) & (!g730) & (!g816) & (g913) & (g910) & (!g911)) + ((!g683) & (!g730) & (!g816) & (g913) & (g910) & (g911)) + ((!g683) & (!g730) & (g816) & (!g913) & (!g910) & (g911)) + ((!g683) & (!g730) & (g816) & (!g913) & (g910) & (!g911)) + ((!g683) & (!g730) & (g816) & (!g913) & (g910) & (g911)) + ((!g683) & (!g730) & (g816) & (g913) & (!g910) & (g911)) + ((!g683) & (!g730) & (g816) & (g913) & (g910) & (!g911)) + ((!g683) & (!g730) & (g816) & (g913) & (g910) & (g911)) + ((!g683) & (g730) & (!g816) & (!g913) & (!g910) & (g911)) + ((!g683) & (g730) & (!g816) & (!g913) & (g910) & (!g911)) + ((!g683) & (g730) & (!g816) & (!g913) & (g910) & (g911)) + ((!g683) & (g730) & (!g816) & (g913) & (!g910) & (g911)) + ((!g683) & (g730) & (!g816) & (g913) & (g910) & (!g911)) + ((!g683) & (g730) & (!g816) & (g913) & (g910) & (g911)) + ((!g683) & (g730) & (g816) & (!g913) & (!g910) & (g911)) + ((!g683) & (g730) & (g816) & (!g913) & (g910) & (!g911)) + ((!g683) & (g730) & (g816) & (!g913) & (g910) & (g911)) + ((!g683) & (g730) & (g816) & (g913) & (!g910) & (!g911)) + ((!g683) & (g730) & (g816) & (g913) & (!g910) & (g911)) + ((!g683) & (g730) & (g816) & (g913) & (g910) & (!g911)) + ((!g683) & (g730) & (g816) & (g913) & (g910) & (g911)) + ((g683) & (!g730) & (!g816) & (g913) & (!g910) & (!g911)) + ((g683) & (g730) & (g816) & (g913) & (!g910) & (!g911)));
	assign g915 = (((!g2) & (!g795) & (!g796) & (!g804) & (!g806) & (!g807)) + ((!g2) & (!g795) & (!g796) & (!g804) & (g806) & (g807)) + ((!g2) & (!g795) & (!g796) & (g804) & (!g806) & (g807)) + ((!g2) & (!g795) & (!g796) & (g804) & (g806) & (!g807)) + ((!g2) & (!g795) & (g796) & (!g804) & (!g806) & (g807)) + ((!g2) & (!g795) & (g796) & (!g804) & (g806) & (!g807)) + ((!g2) & (!g795) & (g796) & (g804) & (!g806) & (g807)) + ((!g2) & (!g795) & (g796) & (g804) & (g806) & (!g807)) + ((!g2) & (g795) & (!g796) & (!g804) & (!g806) & (!g807)) + ((!g2) & (g795) & (!g796) & (!g804) & (g806) & (g807)) + ((!g2) & (g795) & (!g796) & (g804) & (!g806) & (!g807)) + ((!g2) & (g795) & (!g796) & (g804) & (g806) & (g807)) + ((!g2) & (g795) & (g796) & (!g804) & (!g806) & (!g807)) + ((!g2) & (g795) & (g796) & (!g804) & (g806) & (g807)) + ((!g2) & (g795) & (g796) & (g804) & (!g806) & (g807)) + ((!g2) & (g795) & (g796) & (g804) & (g806) & (!g807)) + ((g2) & (!g795) & (!g796) & (!g804) & (!g806) & (g807)) + ((g2) & (!g795) & (!g796) & (!g804) & (g806) & (!g807)) + ((g2) & (!g795) & (!g796) & (g804) & (!g806) & (!g807)) + ((g2) & (!g795) & (!g796) & (g804) & (g806) & (g807)) + ((g2) & (!g795) & (g796) & (!g804) & (!g806) & (!g807)) + ((g2) & (!g795) & (g796) & (!g804) & (g806) & (g807)) + ((g2) & (!g795) & (g796) & (g804) & (!g806) & (!g807)) + ((g2) & (!g795) & (g796) & (g804) & (g806) & (g807)) + ((g2) & (g795) & (!g796) & (!g804) & (!g806) & (g807)) + ((g2) & (g795) & (!g796) & (!g804) & (g806) & (!g807)) + ((g2) & (g795) & (!g796) & (g804) & (!g806) & (g807)) + ((g2) & (g795) & (!g796) & (g804) & (g806) & (!g807)) + ((g2) & (g795) & (g796) & (!g804) & (!g806) & (g807)) + ((g2) & (g795) & (g796) & (!g804) & (g806) & (!g807)) + ((g2) & (g795) & (g796) & (g804) & (!g806) & (!g807)) + ((g2) & (g795) & (g796) & (g804) & (g806) & (g807)));
	assign g916 = (((!g585) & (!sk[30]) & (!g597) & (!g679) & (g864)) + ((!g585) & (!sk[30]) & (!g597) & (g679) & (g864)) + ((!g585) & (!sk[30]) & (g597) & (!g679) & (g864)) + ((!g585) & (!sk[30]) & (g597) & (g679) & (g864)) + ((!g585) & (sk[30]) & (!g597) & (g679) & (g864)) + ((!g585) & (sk[30]) & (g597) & (!g679) & (g864)) + ((g585) & (!sk[30]) & (!g597) & (!g679) & (!g864)) + ((g585) & (!sk[30]) & (!g597) & (!g679) & (g864)) + ((g585) & (!sk[30]) & (!g597) & (g679) & (!g864)) + ((g585) & (!sk[30]) & (!g597) & (g679) & (g864)) + ((g585) & (!sk[30]) & (g597) & (!g679) & (!g864)) + ((g585) & (!sk[30]) & (g597) & (!g679) & (g864)) + ((g585) & (!sk[30]) & (g597) & (g679) & (!g864)) + ((g585) & (!sk[30]) & (g597) & (g679) & (g864)) + ((g585) & (sk[30]) & (!g597) & (!g679) & (g864)) + ((g585) & (sk[30]) & (g597) & (g679) & (g864)));
	assign g917 = (((!g549) & (!g569) & (!g680) & (!g729) & (!g891) & (g892)) + ((!g549) & (!g569) & (!g680) & (!g729) & (g891) & (g892)) + ((!g549) & (!g569) & (g680) & (!g729) & (!g891) & (g892)) + ((!g549) & (!g569) & (g680) & (!g729) & (g891) & (!g892)) + ((!g549) & (!g569) & (g680) & (!g729) & (g891) & (g892)) + ((!g549) & (!g569) & (g680) & (g729) & (g891) & (!g892)) + ((!g549) & (!g569) & (g680) & (g729) & (g891) & (g892)) + ((!g549) & (g569) & (!g680) & (!g729) & (!g891) & (g892)) + ((!g549) & (g569) & (!g680) & (!g729) & (g891) & (!g892)) + ((!g549) & (g569) & (!g680) & (!g729) & (g891) & (g892)) + ((!g549) & (g569) & (!g680) & (g729) & (g891) & (!g892)) + ((!g549) & (g569) & (!g680) & (g729) & (g891) & (g892)) + ((!g549) & (g569) & (g680) & (!g729) & (!g891) & (g892)) + ((!g549) & (g569) & (g680) & (!g729) & (g891) & (g892)) + ((g549) & (!g569) & (!g680) & (!g729) & (!g891) & (g892)) + ((g549) & (!g569) & (!g680) & (!g729) & (g891) & (!g892)) + ((g549) & (!g569) & (!g680) & (!g729) & (g891) & (g892)) + ((g549) & (!g569) & (!g680) & (g729) & (g891) & (!g892)) + ((g549) & (!g569) & (!g680) & (g729) & (g891) & (g892)) + ((g549) & (!g569) & (g680) & (!g729) & (!g891) & (g892)) + ((g549) & (!g569) & (g680) & (!g729) & (g891) & (g892)) + ((g549) & (g569) & (!g680) & (!g729) & (!g891) & (g892)) + ((g549) & (g569) & (!g680) & (!g729) & (g891) & (g892)) + ((g549) & (g569) & (g680) & (!g729) & (!g891) & (g892)) + ((g549) & (g569) & (g680) & (!g729) & (g891) & (!g892)) + ((g549) & (g569) & (g680) & (!g729) & (g891) & (g892)) + ((g549) & (g569) & (g680) & (g729) & (g891) & (!g892)) + ((g549) & (g569) & (g680) & (g729) & (g891) & (g892)));
	assign g918 = (((!ax0x) & (!g683) & (!g791) & (!g866) & (!g916) & (g917)) + ((!ax0x) & (!g683) & (!g791) & (!g866) & (g916) & (!g917)) + ((!ax0x) & (!g683) & (!g791) & (!g866) & (g916) & (g917)) + ((!ax0x) & (!g683) & (!g791) & (g866) & (!g916) & (g917)) + ((!ax0x) & (!g683) & (!g791) & (g866) & (g916) & (!g917)) + ((!ax0x) & (!g683) & (!g791) & (g866) & (g916) & (g917)) + ((!ax0x) & (!g683) & (g791) & (!g866) & (!g916) & (g917)) + ((!ax0x) & (!g683) & (g791) & (!g866) & (g916) & (!g917)) + ((!ax0x) & (!g683) & (g791) & (!g866) & (g916) & (g917)) + ((!ax0x) & (!g683) & (g791) & (g866) & (!g916) & (g917)) + ((!ax0x) & (!g683) & (g791) & (g866) & (g916) & (!g917)) + ((!ax0x) & (!g683) & (g791) & (g866) & (g916) & (g917)) + ((!ax0x) & (g683) & (!g791) & (!g866) & (!g916) & (!g917)) + ((!ax0x) & (g683) & (!g791) & (g866) & (!g916) & (!g917)) + ((!ax0x) & (g683) & (g791) & (!g866) & (!g916) & (!g917)) + ((!ax0x) & (g683) & (g791) & (g866) & (!g916) & (!g917)) + ((ax0x) & (!g683) & (!g791) & (!g866) & (!g916) & (g917)) + ((ax0x) & (!g683) & (!g791) & (!g866) & (g916) & (!g917)) + ((ax0x) & (!g683) & (!g791) & (!g866) & (g916) & (g917)) + ((ax0x) & (!g683) & (!g791) & (g866) & (!g916) & (g917)) + ((ax0x) & (!g683) & (!g791) & (g866) & (g916) & (!g917)) + ((ax0x) & (!g683) & (!g791) & (g866) & (g916) & (g917)) + ((ax0x) & (!g683) & (g791) & (!g866) & (!g916) & (g917)) + ((ax0x) & (!g683) & (g791) & (!g866) & (g916) & (!g917)) + ((ax0x) & (!g683) & (g791) & (!g866) & (g916) & (g917)) + ((ax0x) & (!g683) & (g791) & (g866) & (!g916) & (!g917)) + ((ax0x) & (!g683) & (g791) & (g866) & (!g916) & (g917)) + ((ax0x) & (!g683) & (g791) & (g866) & (g916) & (!g917)) + ((ax0x) & (!g683) & (g791) & (g866) & (g916) & (g917)) + ((ax0x) & (g683) & (!g791) & (!g866) & (!g916) & (!g917)) + ((ax0x) & (g683) & (!g791) & (g866) & (!g916) & (!g917)) + ((ax0x) & (g683) & (g791) & (g866) & (!g916) & (!g917)));
	assign g919 = (((!g585) & (!g597) & (!g679) & (g720) & (g864) & (!g892)) + ((!g585) & (!g597) & (!g679) & (g720) & (g864) & (g892)) + ((!g585) & (!g597) & (g679) & (!g720) & (!g864) & (g892)) + ((!g585) & (!g597) & (g679) & (!g720) & (g864) & (g892)) + ((!g585) & (!g597) & (g679) & (g720) & (!g864) & (g892)) + ((!g585) & (!g597) & (g679) & (g720) & (g864) & (!g892)) + ((!g585) & (!g597) & (g679) & (g720) & (g864) & (g892)) + ((!g585) & (g597) & (!g679) & (!g720) & (!g864) & (g892)) + ((!g585) & (g597) & (!g679) & (!g720) & (g864) & (g892)) + ((!g585) & (g597) & (!g679) & (g720) & (!g864) & (g892)) + ((!g585) & (g597) & (!g679) & (g720) & (g864) & (!g892)) + ((!g585) & (g597) & (!g679) & (g720) & (g864) & (g892)) + ((!g585) & (g597) & (g679) & (g720) & (g864) & (!g892)) + ((!g585) & (g597) & (g679) & (g720) & (g864) & (g892)) + ((g585) & (!g597) & (!g679) & (!g720) & (!g864) & (g892)) + ((g585) & (!g597) & (!g679) & (!g720) & (g864) & (g892)) + ((g585) & (!g597) & (!g679) & (g720) & (!g864) & (g892)) + ((g585) & (!g597) & (!g679) & (g720) & (g864) & (!g892)) + ((g585) & (!g597) & (!g679) & (g720) & (g864) & (g892)) + ((g585) & (!g597) & (g679) & (g720) & (g864) & (!g892)) + ((g585) & (!g597) & (g679) & (g720) & (g864) & (g892)) + ((g585) & (g597) & (!g679) & (g720) & (g864) & (!g892)) + ((g585) & (g597) & (!g679) & (g720) & (g864) & (g892)) + ((g585) & (g597) & (g679) & (!g720) & (!g864) & (g892)) + ((g585) & (g597) & (g679) & (!g720) & (g864) & (g892)) + ((g585) & (g597) & (g679) & (g720) & (!g864) & (g892)) + ((g585) & (g597) & (g679) & (g720) & (g864) & (!g892)) + ((g585) & (g597) & (g679) & (g720) & (g864) & (g892)));
	assign g920 = (((!ax0x) & (!g719) & (!g728) & (!g729) & (!g867) & (!g919)) + ((!ax0x) & (!g719) & (!g728) & (!g729) & (g867) & (!g919)) + ((!ax0x) & (!g719) & (!g728) & (g729) & (!g867) & (!g919)) + ((!ax0x) & (!g719) & (!g728) & (g729) & (g867) & (!g919)) + ((!ax0x) & (!g719) & (g728) & (!g729) & (!g867) & (!g919)) + ((!ax0x) & (!g719) & (g728) & (!g729) & (g867) & (!g919)) + ((!ax0x) & (!g719) & (g728) & (g729) & (!g867) & (!g919)) + ((!ax0x) & (!g719) & (g728) & (g729) & (g867) & (!g919)) + ((!ax0x) & (g719) & (!g728) & (!g729) & (!g867) & (!g919)) + ((!ax0x) & (g719) & (!g728) & (!g729) & (g867) & (!g919)) + ((!ax0x) & (g719) & (!g728) & (g729) & (!g867) & (!g919)) + ((!ax0x) & (g719) & (!g728) & (g729) & (g867) & (!g919)) + ((!ax0x) & (g719) & (g728) & (!g729) & (!g867) & (!g919)) + ((!ax0x) & (g719) & (g728) & (!g729) & (g867) & (!g919)) + ((!ax0x) & (g719) & (g728) & (g729) & (!g867) & (!g919)) + ((!ax0x) & (g719) & (g728) & (g729) & (g867) & (!g919)) + ((ax0x) & (!g719) & (!g728) & (!g729) & (g867) & (!g919)) + ((ax0x) & (!g719) & (!g728) & (g729) & (!g867) & (!g919)) + ((ax0x) & (!g719) & (g728) & (g729) & (!g867) & (!g919)) + ((ax0x) & (!g719) & (g728) & (g729) & (g867) & (!g919)) + ((ax0x) & (g719) & (!g728) & (g729) & (!g867) & (!g919)) + ((ax0x) & (g719) & (!g728) & (g729) & (g867) & (!g919)) + ((ax0x) & (g719) & (g728) & (!g729) & (g867) & (!g919)) + ((ax0x) & (g719) & (g728) & (g729) & (!g867) & (!g919)));
	assign g921 = (((!g2) & (!g797) & (!g800) & (!g801) & (!g802) & (g803)) + ((!g2) & (!g797) & (!g800) & (g801) & (!g802) & (!g803)) + ((!g2) & (!g797) & (!g800) & (g801) & (g802) & (!g803)) + ((!g2) & (!g797) & (!g800) & (g801) & (g802) & (g803)) + ((!g2) & (!g797) & (g800) & (!g801) & (!g802) & (g803)) + ((!g2) & (!g797) & (g800) & (g801) & (!g802) & (g803)) + ((!g2) & (g797) & (!g800) & (!g801) & (!g802) & (!g803)) + ((!g2) & (g797) & (!g800) & (!g801) & (g802) & (!g803)) + ((!g2) & (g797) & (!g800) & (!g801) & (g802) & (g803)) + ((!g2) & (g797) & (!g800) & (g801) & (!g802) & (g803)) + ((!g2) & (g797) & (g800) & (!g801) & (!g802) & (!g803)) + ((!g2) & (g797) & (g800) & (!g801) & (g802) & (!g803)) + ((!g2) & (g797) & (g800) & (!g801) & (g802) & (g803)) + ((!g2) & (g797) & (g800) & (g801) & (!g802) & (!g803)) + ((!g2) & (g797) & (g800) & (g801) & (g802) & (!g803)) + ((!g2) & (g797) & (g800) & (g801) & (g802) & (g803)) + ((g2) & (!g797) & (!g800) & (!g801) & (!g802) & (!g803)) + ((g2) & (!g797) & (!g800) & (!g801) & (g802) & (!g803)) + ((g2) & (!g797) & (!g800) & (!g801) & (g802) & (g803)) + ((g2) & (!g797) & (!g800) & (g801) & (!g802) & (!g803)) + ((g2) & (!g797) & (!g800) & (g801) & (g802) & (!g803)) + ((g2) & (!g797) & (!g800) & (g801) & (g802) & (g803)) + ((g2) & (!g797) & (g800) & (!g801) & (!g802) & (!g803)) + ((g2) & (!g797) & (g800) & (!g801) & (g802) & (!g803)) + ((g2) & (!g797) & (g800) & (!g801) & (g802) & (g803)) + ((g2) & (!g797) & (g800) & (g801) & (!g802) & (g803)) + ((g2) & (g797) & (!g800) & (!g801) & (!g802) & (g803)) + ((g2) & (g797) & (!g800) & (g801) & (!g802) & (g803)) + ((g2) & (g797) & (g800) & (!g801) & (!g802) & (g803)) + ((g2) & (g797) & (g800) & (g801) & (!g802) & (!g803)) + ((g2) & (g797) & (g800) & (g801) & (g802) & (!g803)) + ((g2) & (g797) & (g800) & (g801) & (g802) & (g803)));
	assign g922 = (((!sk[36]) & (!g721) & (g678) & (!g864)) + ((!sk[36]) & (!g721) & (g678) & (g864)) + ((!sk[36]) & (g721) & (g678) & (!g864)) + ((!sk[36]) & (g721) & (g678) & (g864)) + ((sk[36]) & (!g721) & (!g678) & (g864)) + ((sk[36]) & (g721) & (g678) & (g864)));
	assign g923 = (((!g585) & (!g597) & (!g679) & (g720) & (!g891) & (g892)) + ((!g585) & (!g597) & (!g679) & (g720) & (g891) & (g892)) + ((!g585) & (!g597) & (g679) & (!g720) & (g891) & (!g892)) + ((!g585) & (!g597) & (g679) & (!g720) & (g891) & (g892)) + ((!g585) & (!g597) & (g679) & (g720) & (!g891) & (g892)) + ((!g585) & (!g597) & (g679) & (g720) & (g891) & (!g892)) + ((!g585) & (!g597) & (g679) & (g720) & (g891) & (g892)) + ((!g585) & (g597) & (!g679) & (!g720) & (g891) & (!g892)) + ((!g585) & (g597) & (!g679) & (!g720) & (g891) & (g892)) + ((!g585) & (g597) & (!g679) & (g720) & (!g891) & (g892)) + ((!g585) & (g597) & (!g679) & (g720) & (g891) & (!g892)) + ((!g585) & (g597) & (!g679) & (g720) & (g891) & (g892)) + ((!g585) & (g597) & (g679) & (g720) & (!g891) & (g892)) + ((!g585) & (g597) & (g679) & (g720) & (g891) & (g892)) + ((g585) & (!g597) & (!g679) & (!g720) & (g891) & (!g892)) + ((g585) & (!g597) & (!g679) & (!g720) & (g891) & (g892)) + ((g585) & (!g597) & (!g679) & (g720) & (!g891) & (g892)) + ((g585) & (!g597) & (!g679) & (g720) & (g891) & (!g892)) + ((g585) & (!g597) & (!g679) & (g720) & (g891) & (g892)) + ((g585) & (!g597) & (g679) & (g720) & (!g891) & (g892)) + ((g585) & (!g597) & (g679) & (g720) & (g891) & (g892)) + ((g585) & (g597) & (!g679) & (g720) & (!g891) & (g892)) + ((g585) & (g597) & (!g679) & (g720) & (g891) & (g892)) + ((g585) & (g597) & (g679) & (!g720) & (g891) & (!g892)) + ((g585) & (g597) & (g679) & (!g720) & (g891) & (g892)) + ((g585) & (g597) & (g679) & (g720) & (!g891) & (g892)) + ((g585) & (g597) & (g679) & (g720) & (g891) & (!g892)) + ((g585) & (g597) & (g679) & (g720) & (g891) & (g892)));
	assign g924 = (((!ax0x) & (!g683) & (!g771) & (!g866) & (!g922) & (g923)) + ((!ax0x) & (!g683) & (!g771) & (!g866) & (g922) & (!g923)) + ((!ax0x) & (!g683) & (!g771) & (!g866) & (g922) & (g923)) + ((!ax0x) & (!g683) & (!g771) & (g866) & (!g922) & (g923)) + ((!ax0x) & (!g683) & (!g771) & (g866) & (g922) & (!g923)) + ((!ax0x) & (!g683) & (!g771) & (g866) & (g922) & (g923)) + ((!ax0x) & (!g683) & (g771) & (!g866) & (!g922) & (g923)) + ((!ax0x) & (!g683) & (g771) & (!g866) & (g922) & (!g923)) + ((!ax0x) & (!g683) & (g771) & (!g866) & (g922) & (g923)) + ((!ax0x) & (!g683) & (g771) & (g866) & (!g922) & (g923)) + ((!ax0x) & (!g683) & (g771) & (g866) & (g922) & (!g923)) + ((!ax0x) & (!g683) & (g771) & (g866) & (g922) & (g923)) + ((!ax0x) & (g683) & (!g771) & (!g866) & (!g922) & (!g923)) + ((!ax0x) & (g683) & (!g771) & (g866) & (!g922) & (!g923)) + ((!ax0x) & (g683) & (g771) & (!g866) & (!g922) & (!g923)) + ((!ax0x) & (g683) & (g771) & (g866) & (!g922) & (!g923)) + ((ax0x) & (!g683) & (!g771) & (!g866) & (!g922) & (g923)) + ((ax0x) & (!g683) & (!g771) & (!g866) & (g922) & (!g923)) + ((ax0x) & (!g683) & (!g771) & (!g866) & (g922) & (g923)) + ((ax0x) & (!g683) & (!g771) & (g866) & (!g922) & (!g923)) + ((ax0x) & (!g683) & (!g771) & (g866) & (!g922) & (g923)) + ((ax0x) & (!g683) & (!g771) & (g866) & (g922) & (!g923)) + ((ax0x) & (!g683) & (!g771) & (g866) & (g922) & (g923)) + ((ax0x) & (!g683) & (g771) & (!g866) & (!g922) & (g923)) + ((ax0x) & (!g683) & (g771) & (!g866) & (g922) & (!g923)) + ((ax0x) & (!g683) & (g771) & (!g866) & (g922) & (g923)) + ((ax0x) & (!g683) & (g771) & (g866) & (!g922) & (g923)) + ((ax0x) & (!g683) & (g771) & (g866) & (g922) & (!g923)) + ((ax0x) & (!g683) & (g771) & (g866) & (g922) & (g923)) + ((ax0x) & (g683) & (!g771) & (g866) & (!g922) & (!g923)) + ((ax0x) & (g683) & (g771) & (!g866) & (!g922) & (!g923)) + ((ax0x) & (g683) & (g771) & (g866) & (!g922) & (!g923)));
	assign g925 = (((!g721) & (!sk[39]) & (!g678) & (!g723) & (g864) & (!g892)) + ((!g721) & (!sk[39]) & (!g678) & (!g723) & (g864) & (g892)) + ((!g721) & (!sk[39]) & (!g678) & (g723) & (!g864) & (!g892)) + ((!g721) & (!sk[39]) & (!g678) & (g723) & (!g864) & (g892)) + ((!g721) & (!sk[39]) & (!g678) & (g723) & (g864) & (!g892)) + ((!g721) & (!sk[39]) & (!g678) & (g723) & (g864) & (g892)) + ((!g721) & (!sk[39]) & (g678) & (!g723) & (!g864) & (!g892)) + ((!g721) & (!sk[39]) & (g678) & (!g723) & (!g864) & (g892)) + ((!g721) & (!sk[39]) & (g678) & (!g723) & (g864) & (!g892)) + ((!g721) & (!sk[39]) & (g678) & (!g723) & (g864) & (g892)) + ((!g721) & (!sk[39]) & (g678) & (g723) & (!g864) & (!g892)) + ((!g721) & (!sk[39]) & (g678) & (g723) & (!g864) & (g892)) + ((!g721) & (!sk[39]) & (g678) & (g723) & (g864) & (!g892)) + ((!g721) & (!sk[39]) & (g678) & (g723) & (g864) & (g892)) + ((!g721) & (sk[39]) & (!g678) & (!g723) & (!g864) & (g892)) + ((!g721) & (sk[39]) & (!g678) & (!g723) & (g864) & (!g892)) + ((!g721) & (sk[39]) & (!g678) & (!g723) & (g864) & (g892)) + ((!g721) & (sk[39]) & (!g678) & (g723) & (!g864) & (g892)) + ((!g721) & (sk[39]) & (!g678) & (g723) & (g864) & (g892)) + ((!g721) & (sk[39]) & (g678) & (!g723) & (g864) & (!g892)) + ((!g721) & (sk[39]) & (g678) & (!g723) & (g864) & (g892)) + ((g721) & (!sk[39]) & (!g678) & (!g723) & (g864) & (!g892)) + ((g721) & (!sk[39]) & (!g678) & (!g723) & (g864) & (g892)) + ((g721) & (!sk[39]) & (!g678) & (g723) & (!g864) & (!g892)) + ((g721) & (!sk[39]) & (!g678) & (g723) & (!g864) & (g892)) + ((g721) & (!sk[39]) & (!g678) & (g723) & (g864) & (!g892)) + ((g721) & (!sk[39]) & (!g678) & (g723) & (g864) & (g892)) + ((g721) & (!sk[39]) & (g678) & (!g723) & (!g864) & (!g892)) + ((g721) & (!sk[39]) & (g678) & (!g723) & (!g864) & (g892)) + ((g721) & (!sk[39]) & (g678) & (!g723) & (g864) & (!g892)) + ((g721) & (!sk[39]) & (g678) & (!g723) & (g864) & (g892)) + ((g721) & (!sk[39]) & (g678) & (g723) & (!g864) & (!g892)) + ((g721) & (!sk[39]) & (g678) & (g723) & (!g864) & (g892)) + ((g721) & (!sk[39]) & (g678) & (g723) & (g864) & (!g892)) + ((g721) & (!sk[39]) & (g678) & (g723) & (g864) & (g892)) + ((g721) & (sk[39]) & (!g678) & (!g723) & (g864) & (!g892)) + ((g721) & (sk[39]) & (!g678) & (!g723) & (g864) & (g892)) + ((g721) & (sk[39]) & (g678) & (!g723) & (!g864) & (g892)) + ((g721) & (sk[39]) & (g678) & (!g723) & (g864) & (!g892)) + ((g721) & (sk[39]) & (g678) & (!g723) & (g864) & (g892)) + ((g721) & (sk[39]) & (g678) & (g723) & (!g864) & (g892)) + ((g721) & (sk[39]) & (g678) & (g723) & (g864) & (g892)));
	assign g926 = (((!ax0x) & (!g720) & (!g722) & (!g727) & (!g867) & (!g925)) + ((!ax0x) & (!g720) & (!g722) & (!g727) & (g867) & (!g925)) + ((!ax0x) & (!g720) & (!g722) & (g727) & (!g867) & (!g925)) + ((!ax0x) & (!g720) & (!g722) & (g727) & (g867) & (!g925)) + ((!ax0x) & (!g720) & (g722) & (!g727) & (!g867) & (!g925)) + ((!ax0x) & (!g720) & (g722) & (!g727) & (g867) & (!g925)) + ((!ax0x) & (!g720) & (g722) & (g727) & (!g867) & (!g925)) + ((!ax0x) & (!g720) & (g722) & (g727) & (g867) & (!g925)) + ((!ax0x) & (g720) & (!g722) & (!g727) & (!g867) & (!g925)) + ((!ax0x) & (g720) & (!g722) & (!g727) & (g867) & (!g925)) + ((!ax0x) & (g720) & (!g722) & (g727) & (!g867) & (!g925)) + ((!ax0x) & (g720) & (!g722) & (g727) & (g867) & (!g925)) + ((!ax0x) & (g720) & (g722) & (!g727) & (!g867) & (!g925)) + ((!ax0x) & (g720) & (g722) & (!g727) & (g867) & (!g925)) + ((!ax0x) & (g720) & (g722) & (g727) & (!g867) & (!g925)) + ((!ax0x) & (g720) & (g722) & (g727) & (g867) & (!g925)) + ((ax0x) & (!g720) & (!g722) & (!g727) & (!g867) & (!g925)) + ((ax0x) & (!g720) & (!g722) & (g727) & (!g867) & (!g925)) + ((ax0x) & (!g720) & (!g722) & (g727) & (g867) & (!g925)) + ((ax0x) & (!g720) & (g722) & (!g727) & (!g867) & (!g925)) + ((ax0x) & (!g720) & (g722) & (!g727) & (g867) & (!g925)) + ((ax0x) & (!g720) & (g722) & (g727) & (!g867) & (!g925)) + ((ax0x) & (g720) & (!g722) & (!g727) & (g867) & (!g925)) + ((ax0x) & (g720) & (g722) & (g727) & (g867) & (!g925)));
	assign g927 = (((!sk[41]) & (!g641) & (!g655) & (!g677) & (g725) & (!g726)) + ((!sk[41]) & (!g641) & (!g655) & (!g677) & (g725) & (g726)) + ((!sk[41]) & (!g641) & (!g655) & (g677) & (!g725) & (!g726)) + ((!sk[41]) & (!g641) & (!g655) & (g677) & (!g725) & (g726)) + ((!sk[41]) & (!g641) & (!g655) & (g677) & (g725) & (!g726)) + ((!sk[41]) & (!g641) & (!g655) & (g677) & (g725) & (g726)) + ((!sk[41]) & (!g641) & (g655) & (!g677) & (!g725) & (!g726)) + ((!sk[41]) & (!g641) & (g655) & (!g677) & (!g725) & (g726)) + ((!sk[41]) & (!g641) & (g655) & (!g677) & (g725) & (!g726)) + ((!sk[41]) & (!g641) & (g655) & (!g677) & (g725) & (g726)) + ((!sk[41]) & (!g641) & (g655) & (g677) & (!g725) & (!g726)) + ((!sk[41]) & (!g641) & (g655) & (g677) & (!g725) & (g726)) + ((!sk[41]) & (!g641) & (g655) & (g677) & (g725) & (!g726)) + ((!sk[41]) & (!g641) & (g655) & (g677) & (g725) & (g726)) + ((!sk[41]) & (g641) & (!g655) & (!g677) & (g725) & (!g726)) + ((!sk[41]) & (g641) & (!g655) & (!g677) & (g725) & (g726)) + ((!sk[41]) & (g641) & (!g655) & (g677) & (!g725) & (!g726)) + ((!sk[41]) & (g641) & (!g655) & (g677) & (!g725) & (g726)) + ((!sk[41]) & (g641) & (!g655) & (g677) & (g725) & (!g726)) + ((!sk[41]) & (g641) & (!g655) & (g677) & (g725) & (g726)) + ((!sk[41]) & (g641) & (g655) & (!g677) & (!g725) & (!g726)) + ((!sk[41]) & (g641) & (g655) & (!g677) & (!g725) & (g726)) + ((!sk[41]) & (g641) & (g655) & (!g677) & (g725) & (!g726)) + ((!sk[41]) & (g641) & (g655) & (!g677) & (g725) & (g726)) + ((!sk[41]) & (g641) & (g655) & (g677) & (!g725) & (!g726)) + ((!sk[41]) & (g641) & (g655) & (g677) & (!g725) & (g726)) + ((!sk[41]) & (g641) & (g655) & (g677) & (g725) & (!g726)) + ((!sk[41]) & (g641) & (g655) & (g677) & (g725) & (g726)) + ((sk[41]) & (!g641) & (!g655) & (!g677) & (!g725) & (g726)) + ((sk[41]) & (!g641) & (!g655) & (!g677) & (g725) & (!g726)) + ((sk[41]) & (!g641) & (g655) & (g677) & (!g725) & (g726)) + ((sk[41]) & (!g641) & (g655) & (g677) & (g725) & (!g726)) + ((sk[41]) & (g641) & (!g655) & (g677) & (!g725) & (g726)) + ((sk[41]) & (g641) & (!g655) & (g677) & (g725) & (!g726)) + ((sk[41]) & (g641) & (g655) & (!g677) & (!g725) & (g726)) + ((sk[41]) & (g641) & (g655) & (!g677) & (g725) & (!g726)));
	assign g928 = (((!ax0x) & (!ax1x) & (!g490) & (!g658) & (!g676) & (!g867)) + ((!ax0x) & (!ax1x) & (!g490) & (!g658) & (!g676) & (g867)) + ((!ax0x) & (!ax1x) & (!g490) & (!g658) & (g676) & (!g867)) + ((!ax0x) & (!ax1x) & (!g490) & (g658) & (!g676) & (!g867)) + ((!ax0x) & (!ax1x) & (!g490) & (g658) & (g676) & (!g867)) + ((!ax0x) & (!ax1x) & (!g490) & (g658) & (g676) & (g867)) + ((!ax0x) & (!ax1x) & (g490) & (!g658) & (!g676) & (!g867)) + ((!ax0x) & (!ax1x) & (g490) & (!g658) & (g676) & (!g867)) + ((!ax0x) & (!ax1x) & (g490) & (!g658) & (g676) & (g867)) + ((!ax0x) & (!ax1x) & (g490) & (g658) & (!g676) & (!g867)) + ((!ax0x) & (!ax1x) & (g490) & (g658) & (!g676) & (g867)) + ((!ax0x) & (!ax1x) & (g490) & (g658) & (g676) & (!g867)) + ((ax0x) & (!ax1x) & (!g490) & (!g658) & (!g676) & (g867)) + ((ax0x) & (!ax1x) & (!g490) & (g658) & (g676) & (g867)) + ((ax0x) & (!ax1x) & (g490) & (!g658) & (g676) & (g867)) + ((ax0x) & (!ax1x) & (g490) & (g658) & (!g676) & (g867)) + ((ax0x) & (ax1x) & (!g490) & (!g658) & (!g676) & (g867)) + ((ax0x) & (ax1x) & (!g490) & (g658) & (g676) & (g867)) + ((ax0x) & (ax1x) & (g490) & (!g658) & (g676) & (g867)) + ((ax0x) & (ax1x) & (g490) & (g658) & (!g676) & (g867)));
	assign g929 = (((!g656) & (!g489) & (!g545) & (!sk[43]) & (g670)) + ((!g656) & (!g489) & (!g545) & (sk[43]) & (g670)) + ((!g656) & (!g489) & (g545) & (!sk[43]) & (g670)) + ((!g656) & (!g489) & (g545) & (sk[43]) & (!g670)) + ((!g656) & (g489) & (!g545) & (!sk[43]) & (g670)) + ((!g656) & (g489) & (!g545) & (sk[43]) & (!g670)) + ((!g656) & (g489) & (g545) & (!sk[43]) & (g670)) + ((!g656) & (g489) & (g545) & (sk[43]) & (!g670)) + ((g656) & (!g489) & (!g545) & (!sk[43]) & (!g670)) + ((g656) & (!g489) & (!g545) & (!sk[43]) & (g670)) + ((g656) & (!g489) & (!g545) & (sk[43]) & (!g670)) + ((g656) & (!g489) & (g545) & (!sk[43]) & (!g670)) + ((g656) & (!g489) & (g545) & (!sk[43]) & (g670)) + ((g656) & (!g489) & (g545) & (sk[43]) & (g670)) + ((g656) & (g489) & (!g545) & (!sk[43]) & (!g670)) + ((g656) & (g489) & (!g545) & (!sk[43]) & (g670)) + ((g656) & (g489) & (!g545) & (sk[43]) & (g670)) + ((g656) & (g489) & (g545) & (!sk[43]) & (!g670)) + ((g656) & (g489) & (g545) & (!sk[43]) & (g670)) + ((g656) & (g489) & (g545) & (sk[43]) & (g670)));
	assign g930 = (((!g641) & (!g655) & (g929) & (!g677) & (g725) & (!g891)) + ((!g641) & (!g655) & (g929) & (!g677) & (g725) & (g891)) + ((!g641) & (!g655) & (g929) & (g677) & (g725) & (!g891)) + ((!g641) & (g655) & (g929) & (!g677) & (g725) & (!g891)) + ((!g641) & (g655) & (g929) & (g677) & (g725) & (!g891)) + ((!g641) & (g655) & (g929) & (g677) & (g725) & (g891)) + ((g641) & (!g655) & (g929) & (!g677) & (g725) & (!g891)) + ((g641) & (!g655) & (g929) & (g677) & (g725) & (!g891)) + ((g641) & (!g655) & (g929) & (g677) & (g725) & (g891)) + ((g641) & (g655) & (g929) & (!g677) & (g725) & (!g891)) + ((g641) & (g655) & (g929) & (!g677) & (g725) & (g891)) + ((g641) & (g655) & (g929) & (g677) & (g725) & (!g891)));
	assign g931 = (((!ax0x) & (g683) & (!g866) & (!g927) & (!g928) & (g930)) + ((!ax0x) & (g683) & (!g866) & (!g927) & (g928) & (!g930)) + ((!ax0x) & (g683) & (!g866) & (!g927) & (g928) & (g930)) + ((!ax0x) & (g683) & (!g866) & (g927) & (!g928) & (g930)) + ((!ax0x) & (g683) & (!g866) & (g927) & (g928) & (!g930)) + ((!ax0x) & (g683) & (!g866) & (g927) & (g928) & (g930)) + ((!ax0x) & (g683) & (g866) & (!g927) & (!g928) & (g930)) + ((!ax0x) & (g683) & (g866) & (!g927) & (g928) & (!g930)) + ((!ax0x) & (g683) & (g866) & (!g927) & (g928) & (g930)) + ((!ax0x) & (g683) & (g866) & (g927) & (!g928) & (g930)) + ((!ax0x) & (g683) & (g866) & (g927) & (g928) & (!g930)) + ((!ax0x) & (g683) & (g866) & (g927) & (g928) & (g930)) + ((ax0x) & (g683) & (!g866) & (g927) & (!g928) & (g930)) + ((ax0x) & (g683) & (!g866) & (g927) & (g928) & (!g930)) + ((ax0x) & (g683) & (!g866) & (g927) & (g928) & (g930)) + ((ax0x) & (g683) & (g866) & (!g927) & (!g928) & (g930)) + ((ax0x) & (g683) & (g866) & (!g927) & (g928) & (!g930)) + ((ax0x) & (g683) & (g866) & (!g927) & (g928) & (g930)) + ((ax0x) & (g683) & (g866) & (g927) & (!g928) & (g930)) + ((ax0x) & (g683) & (g866) & (g927) & (g928) & (!g930)) + ((ax0x) & (g683) & (g866) & (g927) & (g928) & (g930)));
	assign g932 = (((!g723) & (!g724) & (!g725) & (g726) & (!sk[46]) & (!g868)) + ((!g723) & (!g724) & (!g725) & (g726) & (!sk[46]) & (g868)) + ((!g723) & (!g724) & (!g725) & (g726) & (sk[46]) & (g868)) + ((!g723) & (!g724) & (g725) & (!g726) & (!sk[46]) & (!g868)) + ((!g723) & (!g724) & (g725) & (!g726) & (!sk[46]) & (g868)) + ((!g723) & (!g724) & (g725) & (g726) & (!sk[46]) & (!g868)) + ((!g723) & (!g724) & (g725) & (g726) & (!sk[46]) & (g868)) + ((!g723) & (!g724) & (g725) & (g726) & (sk[46]) & (g868)) + ((!g723) & (g724) & (!g725) & (!g726) & (!sk[46]) & (!g868)) + ((!g723) & (g724) & (!g725) & (!g726) & (!sk[46]) & (g868)) + ((!g723) & (g724) & (!g725) & (!g726) & (sk[46]) & (g868)) + ((!g723) & (g724) & (!g725) & (g726) & (!sk[46]) & (!g868)) + ((!g723) & (g724) & (!g725) & (g726) & (!sk[46]) & (g868)) + ((!g723) & (g724) & (g725) & (!g726) & (!sk[46]) & (!g868)) + ((!g723) & (g724) & (g725) & (!g726) & (!sk[46]) & (g868)) + ((!g723) & (g724) & (g725) & (!g726) & (sk[46]) & (g868)) + ((!g723) & (g724) & (g725) & (g726) & (!sk[46]) & (!g868)) + ((!g723) & (g724) & (g725) & (g726) & (!sk[46]) & (g868)) + ((!g723) & (g724) & (g725) & (g726) & (sk[46]) & (g868)) + ((g723) & (!g724) & (!g725) & (!g726) & (sk[46]) & (g868)) + ((g723) & (!g724) & (!g725) & (g726) & (!sk[46]) & (!g868)) + ((g723) & (!g724) & (!g725) & (g726) & (!sk[46]) & (g868)) + ((g723) & (!g724) & (g725) & (!g726) & (!sk[46]) & (!g868)) + ((g723) & (!g724) & (g725) & (!g726) & (!sk[46]) & (g868)) + ((g723) & (!g724) & (g725) & (!g726) & (sk[46]) & (g868)) + ((g723) & (!g724) & (g725) & (g726) & (!sk[46]) & (!g868)) + ((g723) & (!g724) & (g725) & (g726) & (!sk[46]) & (g868)) + ((g723) & (g724) & (!g725) & (!g726) & (!sk[46]) & (!g868)) + ((g723) & (g724) & (!g725) & (!g726) & (!sk[46]) & (g868)) + ((g723) & (g724) & (!g725) & (g726) & (!sk[46]) & (!g868)) + ((g723) & (g724) & (!g725) & (g726) & (!sk[46]) & (g868)) + ((g723) & (g724) & (!g725) & (g726) & (sk[46]) & (g868)) + ((g723) & (g724) & (g725) & (!g726) & (!sk[46]) & (!g868)) + ((g723) & (g724) & (g725) & (!g726) & (!sk[46]) & (g868)) + ((g723) & (g724) & (g725) & (g726) & (!sk[46]) & (!g868)) + ((g723) & (g724) & (g725) & (g726) & (!sk[46]) & (g868)));
	assign g933 = (((!g723) & (!g724) & (!g726) & (!g891) & (!g864) & (!g892)) + ((!g723) & (!g724) & (!g726) & (!g891) & (g864) & (!g892)) + ((!g723) & (!g724) & (g726) & (!g891) & (!g864) & (!g892)) + ((!g723) & (g724) & (!g726) & (!g891) & (!g864) & (!g892)) + ((!g723) & (g724) & (!g726) & (!g891) & (!g864) & (g892)) + ((!g723) & (g724) & (!g726) & (!g891) & (g864) & (!g892)) + ((!g723) & (g724) & (!g726) & (!g891) & (g864) & (g892)) + ((!g723) & (g724) & (g726) & (!g891) & (!g864) & (!g892)) + ((!g723) & (g724) & (g726) & (!g891) & (!g864) & (g892)) + ((g723) & (!g724) & (!g726) & (!g891) & (!g864) & (!g892)) + ((g723) & (!g724) & (!g726) & (!g891) & (g864) & (!g892)) + ((g723) & (!g724) & (!g726) & (g891) & (!g864) & (!g892)) + ((g723) & (!g724) & (!g726) & (g891) & (g864) & (!g892)) + ((g723) & (!g724) & (g726) & (!g891) & (!g864) & (!g892)) + ((g723) & (!g724) & (g726) & (g891) & (!g864) & (!g892)) + ((g723) & (g724) & (!g726) & (!g891) & (!g864) & (!g892)) + ((g723) & (g724) & (!g726) & (!g891) & (!g864) & (g892)) + ((g723) & (g724) & (!g726) & (!g891) & (g864) & (!g892)) + ((g723) & (g724) & (!g726) & (!g891) & (g864) & (g892)) + ((g723) & (g724) & (!g726) & (g891) & (!g864) & (!g892)) + ((g723) & (g724) & (!g726) & (g891) & (!g864) & (g892)) + ((g723) & (g724) & (!g726) & (g891) & (g864) & (!g892)) + ((g723) & (g724) & (!g726) & (g891) & (g864) & (g892)) + ((g723) & (g724) & (g726) & (!g891) & (!g864) & (!g892)) + ((g723) & (g724) & (g726) & (!g891) & (!g864) & (g892)) + ((g723) & (g724) & (g726) & (g891) & (!g864) & (!g892)) + ((g723) & (g724) & (g726) & (g891) & (!g864) & (g892)));
	assign g934 = (((!g414) & (!g683) & (!g725) & (g931) & (!g932) & (!g933)) + ((!g414) & (!g683) & (!g725) & (g931) & (g932) & (!g933)) + ((!g414) & (!g683) & (!g725) & (g931) & (g932) & (g933)) + ((!g414) & (!g683) & (g725) & (g931) & (!g932) & (!g933)) + ((!g414) & (!g683) & (g725) & (g931) & (g932) & (!g933)) + ((!g414) & (!g683) & (g725) & (g931) & (g932) & (g933)) + ((!g414) & (g683) & (!g725) & (!g931) & (!g932) & (g933)) + ((!g414) & (g683) & (!g725) & (g931) & (!g932) & (!g933)) + ((!g414) & (g683) & (!g725) & (g931) & (!g932) & (g933)) + ((!g414) & (g683) & (!g725) & (g931) & (g932) & (!g933)) + ((!g414) & (g683) & (!g725) & (g931) & (g932) & (g933)) + ((!g414) & (g683) & (g725) & (g931) & (!g932) & (g933)) + ((g414) & (!g683) & (!g725) & (!g931) & (!g932) & (!g933)) + ((g414) & (!g683) & (!g725) & (!g931) & (g932) & (!g933)) + ((g414) & (!g683) & (!g725) & (!g931) & (g932) & (g933)) + ((g414) & (!g683) & (!g725) & (g931) & (!g932) & (!g933)) + ((g414) & (!g683) & (!g725) & (g931) & (!g932) & (g933)) + ((g414) & (!g683) & (!g725) & (g931) & (g932) & (!g933)) + ((g414) & (!g683) & (!g725) & (g931) & (g932) & (g933)) + ((g414) & (!g683) & (g725) & (g931) & (!g932) & (!g933)) + ((g414) & (!g683) & (g725) & (g931) & (g932) & (!g933)) + ((g414) & (!g683) & (g725) & (g931) & (g932) & (g933)) + ((g414) & (g683) & (!g725) & (g931) & (!g932) & (g933)) + ((g414) & (g683) & (g725) & (g931) & (!g932) & (g933)));
	assign g935 = (((!g401) & (!g414) & (!g683) & (g725) & (!sk[49]) & (!g726)) + ((!g401) & (!g414) & (!g683) & (g725) & (!sk[49]) & (g726)) + ((!g401) & (!g414) & (g683) & (!g725) & (!sk[49]) & (!g726)) + ((!g401) & (!g414) & (g683) & (!g725) & (!sk[49]) & (g726)) + ((!g401) & (!g414) & (g683) & (!g725) & (sk[49]) & (g726)) + ((!g401) & (!g414) & (g683) & (g725) & (!sk[49]) & (!g726)) + ((!g401) & (!g414) & (g683) & (g725) & (!sk[49]) & (g726)) + ((!g401) & (!g414) & (g683) & (g725) & (sk[49]) & (g726)) + ((!g401) & (g414) & (!g683) & (!g725) & (!sk[49]) & (!g726)) + ((!g401) & (g414) & (!g683) & (!g725) & (!sk[49]) & (g726)) + ((!g401) & (g414) & (!g683) & (!g725) & (sk[49]) & (g726)) + ((!g401) & (g414) & (!g683) & (g725) & (!sk[49]) & (!g726)) + ((!g401) & (g414) & (!g683) & (g725) & (!sk[49]) & (g726)) + ((!g401) & (g414) & (!g683) & (g725) & (sk[49]) & (g726)) + ((!g401) & (g414) & (g683) & (!g725) & (!sk[49]) & (!g726)) + ((!g401) & (g414) & (g683) & (!g725) & (!sk[49]) & (g726)) + ((!g401) & (g414) & (g683) & (!g725) & (sk[49]) & (!g726)) + ((!g401) & (g414) & (g683) & (!g725) & (sk[49]) & (g726)) + ((!g401) & (g414) & (g683) & (g725) & (!sk[49]) & (!g726)) + ((!g401) & (g414) & (g683) & (g725) & (!sk[49]) & (g726)) + ((g401) & (!g414) & (!g683) & (!g725) & (sk[49]) & (!g726)) + ((g401) & (!g414) & (!g683) & (!g725) & (sk[49]) & (g726)) + ((g401) & (!g414) & (!g683) & (g725) & (!sk[49]) & (!g726)) + ((g401) & (!g414) & (!g683) & (g725) & (!sk[49]) & (g726)) + ((g401) & (!g414) & (g683) & (!g725) & (!sk[49]) & (!g726)) + ((g401) & (!g414) & (g683) & (!g725) & (!sk[49]) & (g726)) + ((g401) & (!g414) & (g683) & (!g725) & (sk[49]) & (!g726)) + ((g401) & (!g414) & (g683) & (g725) & (!sk[49]) & (!g726)) + ((g401) & (!g414) & (g683) & (g725) & (!sk[49]) & (g726)) + ((g401) & (!g414) & (g683) & (g725) & (sk[49]) & (g726)) + ((g401) & (g414) & (!g683) & (!g725) & (!sk[49]) & (!g726)) + ((g401) & (g414) & (!g683) & (!g725) & (!sk[49]) & (g726)) + ((g401) & (g414) & (!g683) & (!g725) & (sk[49]) & (!g726)) + ((g401) & (g414) & (!g683) & (g725) & (!sk[49]) & (!g726)) + ((g401) & (g414) & (!g683) & (g725) & (!sk[49]) & (g726)) + ((g401) & (g414) & (!g683) & (g725) & (sk[49]) & (g726)) + ((g401) & (g414) & (g683) & (!g725) & (!sk[49]) & (!g726)) + ((g401) & (g414) & (g683) & (!g725) & (!sk[49]) & (g726)) + ((g401) & (g414) & (g683) & (g725) & (!sk[49]) & (!g726)) + ((g401) & (g414) & (g683) & (g725) & (!sk[49]) & (g726)));
	assign g936 = (((!g723) & (!sk[50]) & (!g724) & (!g864) & (g892)) + ((!g723) & (!sk[50]) & (!g724) & (g864) & (g892)) + ((!g723) & (!sk[50]) & (g724) & (!g864) & (g892)) + ((!g723) & (!sk[50]) & (g724) & (g864) & (g892)) + ((!g723) & (sk[50]) & (!g724) & (!g864) & (g892)) + ((!g723) & (sk[50]) & (!g724) & (g864) & (!g892)) + ((!g723) & (sk[50]) & (!g724) & (g864) & (g892)) + ((!g723) & (sk[50]) & (g724) & (!g864) & (g892)) + ((!g723) & (sk[50]) & (g724) & (g864) & (g892)) + ((g723) & (!sk[50]) & (!g724) & (!g864) & (!g892)) + ((g723) & (!sk[50]) & (!g724) & (!g864) & (g892)) + ((g723) & (!sk[50]) & (!g724) & (g864) & (!g892)) + ((g723) & (!sk[50]) & (!g724) & (g864) & (g892)) + ((g723) & (!sk[50]) & (g724) & (!g864) & (!g892)) + ((g723) & (!sk[50]) & (g724) & (!g864) & (g892)) + ((g723) & (!sk[50]) & (g724) & (g864) & (!g892)) + ((g723) & (!sk[50]) & (g724) & (g864) & (g892)) + ((g723) & (sk[50]) & (!g724) & (g864) & (!g892)) + ((g723) & (sk[50]) & (!g724) & (g864) & (g892)));
	assign g937 = (((!ax0x) & (!g683) & (!g722) & (!g754) & (!g866) & (g936)) + ((!ax0x) & (!g683) & (!g722) & (!g754) & (g866) & (g936)) + ((!ax0x) & (!g683) & (!g722) & (g754) & (!g866) & (g936)) + ((!ax0x) & (!g683) & (!g722) & (g754) & (g866) & (g936)) + ((!ax0x) & (!g683) & (g722) & (!g754) & (!g866) & (g936)) + ((!ax0x) & (!g683) & (g722) & (!g754) & (g866) & (g936)) + ((!ax0x) & (!g683) & (g722) & (g754) & (!g866) & (g936)) + ((!ax0x) & (!g683) & (g722) & (g754) & (g866) & (g936)) + ((!ax0x) & (g683) & (!g722) & (!g754) & (!g866) & (!g936)) + ((!ax0x) & (g683) & (!g722) & (!g754) & (g866) & (!g936)) + ((!ax0x) & (g683) & (!g722) & (g754) & (!g866) & (!g936)) + ((!ax0x) & (g683) & (!g722) & (g754) & (g866) & (!g936)) + ((!ax0x) & (g683) & (g722) & (!g754) & (!g866) & (!g936)) + ((!ax0x) & (g683) & (g722) & (!g754) & (g866) & (!g936)) + ((!ax0x) & (g683) & (g722) & (g754) & (!g866) & (!g936)) + ((!ax0x) & (g683) & (g722) & (g754) & (g866) & (!g936)) + ((ax0x) & (!g683) & (!g722) & (!g754) & (!g866) & (!g936)) + ((ax0x) & (!g683) & (!g722) & (!g754) & (!g866) & (g936)) + ((ax0x) & (!g683) & (!g722) & (!g754) & (g866) & (g936)) + ((ax0x) & (!g683) & (!g722) & (g754) & (!g866) & (!g936)) + ((ax0x) & (!g683) & (!g722) & (g754) & (!g866) & (g936)) + ((ax0x) & (!g683) & (!g722) & (g754) & (g866) & (!g936)) + ((ax0x) & (!g683) & (!g722) & (g754) & (g866) & (g936)) + ((ax0x) & (!g683) & (g722) & (!g754) & (!g866) & (g936)) + ((ax0x) & (!g683) & (g722) & (!g754) & (g866) & (g936)) + ((ax0x) & (!g683) & (g722) & (g754) & (!g866) & (g936)) + ((ax0x) & (!g683) & (g722) & (g754) & (g866) & (!g936)) + ((ax0x) & (!g683) & (g722) & (g754) & (g866) & (g936)) + ((ax0x) & (g683) & (!g722) & (!g754) & (!g866) & (!g936)) + ((ax0x) & (g683) & (g722) & (!g754) & (!g866) & (!g936)) + ((ax0x) & (g683) & (g722) & (!g754) & (g866) & (!g936)) + ((ax0x) & (g683) & (g722) & (g754) & (g866) & (!g936)));
	assign g938 = (((!g2) & (!g732) & (!g746) & (!g798) & (!g799) & (g801)) + ((!g2) & (!g732) & (!g746) & (!g798) & (g799) & (!g801)) + ((!g2) & (!g732) & (!g746) & (g798) & (!g799) & (!g801)) + ((!g2) & (!g732) & (!g746) & (g798) & (g799) & (!g801)) + ((!g2) & (!g732) & (g746) & (!g798) & (!g799) & (g801)) + ((!g2) & (!g732) & (g746) & (!g798) & (g799) & (!g801)) + ((!g2) & (!g732) & (g746) & (g798) & (!g799) & (!g801)) + ((!g2) & (!g732) & (g746) & (g798) & (g799) & (!g801)) + ((!g2) & (g732) & (!g746) & (!g798) & (!g799) & (!g801)) + ((!g2) & (g732) & (!g746) & (!g798) & (g799) & (!g801)) + ((!g2) & (g732) & (!g746) & (g798) & (!g799) & (!g801)) + ((!g2) & (g732) & (!g746) & (g798) & (g799) & (!g801)) + ((!g2) & (g732) & (g746) & (!g798) & (!g799) & (g801)) + ((!g2) & (g732) & (g746) & (!g798) & (g799) & (!g801)) + ((!g2) & (g732) & (g746) & (g798) & (!g799) & (!g801)) + ((!g2) & (g732) & (g746) & (g798) & (g799) & (!g801)) + ((g2) & (!g732) & (!g746) & (!g798) & (!g799) & (!g801)) + ((g2) & (!g732) & (!g746) & (!g798) & (g799) & (g801)) + ((g2) & (!g732) & (!g746) & (g798) & (!g799) & (g801)) + ((g2) & (!g732) & (!g746) & (g798) & (g799) & (g801)) + ((g2) & (!g732) & (g746) & (!g798) & (!g799) & (!g801)) + ((g2) & (!g732) & (g746) & (!g798) & (g799) & (g801)) + ((g2) & (!g732) & (g746) & (g798) & (!g799) & (g801)) + ((g2) & (!g732) & (g746) & (g798) & (g799) & (g801)) + ((g2) & (g732) & (!g746) & (!g798) & (!g799) & (g801)) + ((g2) & (g732) & (!g746) & (!g798) & (g799) & (g801)) + ((g2) & (g732) & (!g746) & (g798) & (!g799) & (g801)) + ((g2) & (g732) & (!g746) & (g798) & (g799) & (g801)) + ((g2) & (g732) & (g746) & (!g798) & (!g799) & (!g801)) + ((g2) & (g732) & (g746) & (!g798) & (g799) & (g801)) + ((g2) & (g732) & (g746) & (g798) & (!g799) & (g801)) + ((g2) & (g732) & (g746) & (g798) & (g799) & (g801)));
	assign g939 = (((!g683) & (!g926) & (!g934) & (!g935) & (!g937) & (g938)) + ((!g683) & (!g926) & (!g934) & (!g935) & (g937) & (g938)) + ((!g683) & (!g926) & (!g934) & (g935) & (!g937) & (g938)) + ((!g683) & (!g926) & (!g934) & (g935) & (g937) & (!g938)) + ((!g683) & (!g926) & (!g934) & (g935) & (g937) & (g938)) + ((!g683) & (!g926) & (g934) & (!g935) & (!g937) & (g938)) + ((!g683) & (!g926) & (g934) & (!g935) & (g937) & (!g938)) + ((!g683) & (!g926) & (g934) & (!g935) & (g937) & (g938)) + ((!g683) & (!g926) & (g934) & (g935) & (!g937) & (!g938)) + ((!g683) & (!g926) & (g934) & (g935) & (!g937) & (g938)) + ((!g683) & (!g926) & (g934) & (g935) & (g937) & (!g938)) + ((!g683) & (!g926) & (g934) & (g935) & (g937) & (g938)) + ((!g683) & (g926) & (!g934) & (g935) & (g937) & (g938)) + ((!g683) & (g926) & (g934) & (!g935) & (g937) & (g938)) + ((!g683) & (g926) & (g934) & (g935) & (!g937) & (g938)) + ((!g683) & (g926) & (g934) & (g935) & (g937) & (g938)) + ((g683) & (!g926) & (!g934) & (g935) & (g937) & (g938)) + ((g683) & (!g926) & (g934) & (!g935) & (g937) & (g938)) + ((g683) & (!g926) & (g934) & (g935) & (!g937) & (g938)) + ((g683) & (!g926) & (g934) & (g935) & (g937) & (g938)) + ((g683) & (g926) & (!g934) & (!g935) & (!g937) & (g938)) + ((g683) & (g926) & (!g934) & (!g935) & (g937) & (g938)) + ((g683) & (g926) & (!g934) & (g935) & (!g937) & (g938)) + ((g683) & (g926) & (!g934) & (g935) & (g937) & (!g938)) + ((g683) & (g926) & (!g934) & (g935) & (g937) & (g938)) + ((g683) & (g926) & (g934) & (!g935) & (!g937) & (g938)) + ((g683) & (g926) & (g934) & (!g935) & (g937) & (!g938)) + ((g683) & (g926) & (g934) & (!g935) & (g937) & (g938)) + ((g683) & (g926) & (g934) & (g935) & (!g937) & (!g938)) + ((g683) & (g926) & (g934) & (g935) & (!g937) & (g938)) + ((g683) & (g926) & (g934) & (g935) & (g937) & (!g938)) + ((g683) & (g926) & (g934) & (g935) & (g937) & (g938)));
	assign g940 = (((!sk[54]) & (!g795) & (g796) & (!g804)) + ((!sk[54]) & (!g795) & (g796) & (g804)) + ((!sk[54]) & (g795) & (g796) & (!g804)) + ((!sk[54]) & (g795) & (g796) & (g804)) + ((sk[54]) & (!g795) & (!g796) & (!g804)) + ((sk[54]) & (!g795) & (g796) & (g804)) + ((sk[54]) & (g795) & (!g796) & (g804)) + ((sk[54]) & (g795) & (g796) & (!g804)));
	assign g941 = (((!g683) & (!g920) & (!g921) & (!g924) & (!g939) & (g940)) + ((!g683) & (!g920) & (!g921) & (!g924) & (g939) & (!g940)) + ((!g683) & (!g920) & (!g921) & (!g924) & (g939) & (g940)) + ((!g683) & (!g920) & (!g921) & (g924) & (!g939) & (!g940)) + ((!g683) & (!g920) & (!g921) & (g924) & (!g939) & (g940)) + ((!g683) & (!g920) & (!g921) & (g924) & (g939) & (!g940)) + ((!g683) & (!g920) & (!g921) & (g924) & (g939) & (g940)) + ((!g683) & (!g920) & (g921) & (!g924) & (!g939) & (g940)) + ((!g683) & (!g920) & (g921) & (!g924) & (g939) & (g940)) + ((!g683) & (!g920) & (g921) & (g924) & (!g939) & (g940)) + ((!g683) & (!g920) & (g921) & (g924) & (g939) & (!g940)) + ((!g683) & (!g920) & (g921) & (g924) & (g939) & (g940)) + ((!g683) & (g920) & (!g921) & (!g924) & (g939) & (g940)) + ((!g683) & (g920) & (!g921) & (g924) & (!g939) & (g940)) + ((!g683) & (g920) & (!g921) & (g924) & (g939) & (g940)) + ((!g683) & (g920) & (g921) & (g924) & (g939) & (g940)) + ((g683) & (!g920) & (!g921) & (!g924) & (g939) & (g940)) + ((g683) & (!g920) & (!g921) & (g924) & (!g939) & (g940)) + ((g683) & (!g920) & (!g921) & (g924) & (g939) & (g940)) + ((g683) & (!g920) & (g921) & (g924) & (g939) & (g940)) + ((g683) & (g920) & (!g921) & (!g924) & (!g939) & (g940)) + ((g683) & (g920) & (!g921) & (!g924) & (g939) & (!g940)) + ((g683) & (g920) & (!g921) & (!g924) & (g939) & (g940)) + ((g683) & (g920) & (!g921) & (g924) & (!g939) & (!g940)) + ((g683) & (g920) & (!g921) & (g924) & (!g939) & (g940)) + ((g683) & (g920) & (!g921) & (g924) & (g939) & (!g940)) + ((g683) & (g920) & (!g921) & (g924) & (g939) & (g940)) + ((g683) & (g920) & (g921) & (!g924) & (!g939) & (g940)) + ((g683) & (g920) & (g921) & (!g924) & (g939) & (g940)) + ((g683) & (g920) & (g921) & (g924) & (!g939) & (g940)) + ((g683) & (g920) & (g921) & (g924) & (g939) & (!g940)) + ((g683) & (g920) & (g921) & (g924) & (g939) & (g940)));
	assign g942 = (((!g909) & (!g912) & (!g914) & (!g915) & (!g918) & (!g941)) + ((!g909) & (!g912) & (!g914) & (!g915) & (!g918) & (g941)) + ((!g909) & (!g912) & (!g914) & (!g915) & (g918) & (!g941)) + ((!g909) & (!g912) & (!g914) & (!g915) & (g918) & (g941)) + ((!g909) & (!g912) & (!g914) & (g915) & (!g918) & (!g941)) + ((!g909) & (!g912) & (!g914) & (g915) & (!g918) & (g941)) + ((!g909) & (!g912) & (!g914) & (g915) & (g918) & (!g941)) + ((!g909) & (!g912) & (!g914) & (g915) & (g918) & (g941)) + ((!g909) & (!g912) & (g914) & (!g915) & (!g918) & (!g941)) + ((!g909) & (!g912) & (g914) & (!g915) & (!g918) & (g941)) + ((!g909) & (!g912) & (g914) & (!g915) & (g918) & (!g941)) + ((!g909) & (!g912) & (g914) & (g915) & (!g918) & (!g941)) + ((!g909) & (g912) & (!g914) & (!g915) & (!g918) & (!g941)) + ((!g909) & (g912) & (!g914) & (!g915) & (!g918) & (g941)) + ((!g909) & (g912) & (!g914) & (!g915) & (g918) & (!g941)) + ((!g909) & (g912) & (!g914) & (g915) & (!g918) & (!g941)) + ((!g909) & (g912) & (g914) & (!g915) & (!g918) & (!g941)) + ((!g909) & (g912) & (g914) & (!g915) & (!g918) & (g941)) + ((!g909) & (g912) & (g914) & (!g915) & (g918) & (!g941)) + ((!g909) & (g912) & (g914) & (g915) & (!g918) & (!g941)) + ((g909) & (!g912) & (!g914) & (!g915) & (!g918) & (!g941)) + ((g909) & (!g912) & (!g914) & (!g915) & (!g918) & (g941)) + ((g909) & (!g912) & (!g914) & (!g915) & (g918) & (!g941)) + ((g909) & (!g912) & (!g914) & (g915) & (!g918) & (!g941)));
	assign g943 = (((!g683) & (!g902) & (!g904) & (!g905) & (!g908) & (!g942)) + ((!g683) & (!g902) & (!g904) & (!g905) & (!g908) & (g942)) + ((!g683) & (!g902) & (!g904) & (!g905) & (g908) & (!g942)) + ((!g683) & (!g902) & (!g904) & (!g905) & (g908) & (g942)) + ((!g683) & (!g902) & (!g904) & (g905) & (!g908) & (!g942)) + ((!g683) & (!g902) & (!g904) & (g905) & (!g908) & (g942)) + ((!g683) & (!g902) & (!g904) & (g905) & (g908) & (!g942)) + ((!g683) & (!g902) & (!g904) & (g905) & (g908) & (g942)) + ((!g683) & (!g902) & (g904) & (!g905) & (!g908) & (!g942)) + ((!g683) & (!g902) & (g904) & (!g905) & (g908) & (!g942)) + ((!g683) & (!g902) & (g904) & (!g905) & (g908) & (g942)) + ((!g683) & (!g902) & (g904) & (g905) & (g908) & (!g942)) + ((!g683) & (g902) & (!g904) & (!g905) & (!g908) & (!g942)) + ((!g683) & (g902) & (!g904) & (!g905) & (g908) & (!g942)) + ((!g683) & (g902) & (!g904) & (!g905) & (g908) & (g942)) + ((!g683) & (g902) & (!g904) & (g905) & (g908) & (!g942)) + ((g683) & (!g902) & (!g904) & (!g905) & (!g908) & (!g942)) + ((g683) & (!g902) & (!g904) & (!g905) & (g908) & (!g942)) + ((g683) & (!g902) & (!g904) & (!g905) & (g908) & (g942)) + ((g683) & (!g902) & (!g904) & (g905) & (g908) & (!g942)) + ((g683) & (!g902) & (g904) & (!g905) & (!g908) & (!g942)) + ((g683) & (!g902) & (g904) & (!g905) & (!g908) & (g942)) + ((g683) & (!g902) & (g904) & (!g905) & (g908) & (!g942)) + ((g683) & (!g902) & (g904) & (!g905) & (g908) & (g942)) + ((g683) & (!g902) & (g904) & (g905) & (!g908) & (!g942)) + ((g683) & (!g902) & (g904) & (g905) & (!g908) & (g942)) + ((g683) & (!g902) & (g904) & (g905) & (g908) & (!g942)) + ((g683) & (!g902) & (g904) & (g905) & (g908) & (g942)) + ((g683) & (g902) & (g904) & (!g905) & (!g908) & (!g942)) + ((g683) & (g902) & (g904) & (!g905) & (g908) & (!g942)) + ((g683) & (g902) & (g904) & (!g905) & (g908) & (g942)) + ((g683) & (g902) & (g904) & (g905) & (g908) & (!g942)));
	assign g944 = (((!g736) & (!sk[58]) & (!g780) & (!g788) & (g821)) + ((!g736) & (!sk[58]) & (!g780) & (g788) & (g821)) + ((!g736) & (!sk[58]) & (g780) & (!g788) & (g821)) + ((!g736) & (!sk[58]) & (g780) & (g788) & (g821)) + ((!g736) & (sk[58]) & (!g780) & (!g788) & (!g821)) + ((!g736) & (sk[58]) & (!g780) & (g788) & (g821)) + ((!g736) & (sk[58]) & (g780) & (!g788) & (g821)) + ((!g736) & (sk[58]) & (g780) & (g788) & (!g821)) + ((g736) & (!sk[58]) & (!g780) & (!g788) & (!g821)) + ((g736) & (!sk[58]) & (!g780) & (!g788) & (g821)) + ((g736) & (!sk[58]) & (!g780) & (g788) & (!g821)) + ((g736) & (!sk[58]) & (!g780) & (g788) & (g821)) + ((g736) & (!sk[58]) & (g780) & (!g788) & (!g821)) + ((g736) & (!sk[58]) & (g780) & (!g788) & (g821)) + ((g736) & (!sk[58]) & (g780) & (g788) & (!g821)) + ((g736) & (!sk[58]) & (g780) & (g788) & (g821)) + ((g736) & (sk[58]) & (!g780) & (!g788) & (g821)) + ((g736) & (sk[58]) & (!g780) & (g788) & (!g821)) + ((g736) & (sk[58]) & (g780) & (!g788) & (!g821)) + ((g736) & (sk[58]) & (g780) & (g788) & (g821)));
	assign g945 = (((!g683) & (!g897) & (!g898) & (!g901) & (!g943) & (!g944)) + ((!g683) & (!g897) & (!g898) & (!g901) & (!g943) & (g944)) + ((!g683) & (!g897) & (!g898) & (!g901) & (g943) & (!g944)) + ((!g683) & (!g897) & (!g898) & (!g901) & (g943) & (g944)) + ((!g683) & (!g897) & (!g898) & (g901) & (!g943) & (g944)) + ((!g683) & (!g897) & (!g898) & (g901) & (g943) & (!g944)) + ((!g683) & (!g897) & (!g898) & (g901) & (g943) & (g944)) + ((!g683) & (!g897) & (g898) & (!g901) & (!g943) & (g944)) + ((!g683) & (!g897) & (g898) & (!g901) & (g943) & (!g944)) + ((!g683) & (!g897) & (g898) & (!g901) & (g943) & (g944)) + ((!g683) & (!g897) & (g898) & (g901) & (!g943) & (g944)) + ((!g683) & (!g897) & (g898) & (g901) & (g943) & (g944)) + ((!g683) & (g897) & (!g898) & (!g901) & (!g943) & (g944)) + ((!g683) & (g897) & (!g898) & (!g901) & (g943) & (g944)) + ((!g683) & (g897) & (!g898) & (g901) & (g943) & (g944)) + ((!g683) & (g897) & (g898) & (!g901) & (g943) & (g944)) + ((g683) & (!g897) & (!g898) & (!g901) & (g943) & (g944)) + ((g683) & (!g897) & (!g898) & (g901) & (!g943) & (g944)) + ((g683) & (!g897) & (!g898) & (g901) & (g943) & (g944)) + ((g683) & (!g897) & (g898) & (g901) & (g943) & (g944)) + ((g683) & (g897) & (!g898) & (!g901) & (!g943) & (g944)) + ((g683) & (g897) & (!g898) & (!g901) & (g943) & (!g944)) + ((g683) & (g897) & (!g898) & (!g901) & (g943) & (g944)) + ((g683) & (g897) & (!g898) & (g901) & (!g943) & (!g944)) + ((g683) & (g897) & (!g898) & (g901) & (!g943) & (g944)) + ((g683) & (g897) & (!g898) & (g901) & (g943) & (!g944)) + ((g683) & (g897) & (!g898) & (g901) & (g943) & (g944)) + ((g683) & (g897) & (g898) & (!g901) & (!g943) & (g944)) + ((g683) & (g897) & (g898) & (!g901) & (g943) & (g944)) + ((g683) & (g897) & (g898) & (g901) & (!g943) & (g944)) + ((g683) & (g897) & (g898) & (g901) & (g943) & (!g944)) + ((g683) & (g897) & (g898) & (g901) & (g943) & (g944)));
	assign g946 = (((!g736) & (!g780) & (!g788) & (!g821) & (!g837) & (!g855)) + ((!g736) & (!g780) & (!g788) & (!g821) & (g837) & (!g855)) + ((!g736) & (!g780) & (!g788) & (!g821) & (g837) & (g855)) + ((!g736) & (!g780) & (!g788) & (g821) & (!g837) & (!g855)) + ((!g736) & (!g780) & (!g788) & (g821) & (g837) & (!g855)) + ((!g736) & (!g780) & (!g788) & (g821) & (g837) & (g855)) + ((!g736) & (!g780) & (g788) & (!g821) & (!g837) & (!g855)) + ((!g736) & (!g780) & (g788) & (!g821) & (g837) & (!g855)) + ((!g736) & (!g780) & (g788) & (!g821) & (g837) & (g855)) + ((!g736) & (!g780) & (g788) & (g821) & (g837) & (!g855)) + ((!g736) & (g780) & (!g788) & (!g821) & (!g837) & (!g855)) + ((!g736) & (g780) & (!g788) & (!g821) & (g837) & (!g855)) + ((!g736) & (g780) & (!g788) & (!g821) & (g837) & (g855)) + ((!g736) & (g780) & (!g788) & (g821) & (g837) & (!g855)) + ((!g736) & (g780) & (g788) & (!g821) & (!g837) & (!g855)) + ((!g736) & (g780) & (g788) & (!g821) & (g837) & (!g855)) + ((!g736) & (g780) & (g788) & (!g821) & (g837) & (g855)) + ((!g736) & (g780) & (g788) & (g821) & (!g837) & (!g855)) + ((!g736) & (g780) & (g788) & (g821) & (g837) & (!g855)) + ((!g736) & (g780) & (g788) & (g821) & (g837) & (g855)) + ((g736) & (!g780) & (!g788) & (!g821) & (!g837) & (!g855)) + ((g736) & (!g780) & (!g788) & (!g821) & (g837) & (!g855)) + ((g736) & (!g780) & (!g788) & (!g821) & (g837) & (g855)) + ((g736) & (!g780) & (!g788) & (g821) & (g837) & (!g855)) + ((g736) & (!g780) & (g788) & (!g821) & (g837) & (!g855)) + ((g736) & (!g780) & (g788) & (g821) & (g837) & (!g855)) + ((g736) & (g780) & (!g788) & (!g821) & (g837) & (!g855)) + ((g736) & (g780) & (!g788) & (g821) & (g837) & (!g855)) + ((g736) & (g780) & (g788) & (!g821) & (!g837) & (!g855)) + ((g736) & (g780) & (g788) & (!g821) & (g837) & (!g855)) + ((g736) & (g780) & (g788) & (!g821) & (g837) & (g855)) + ((g736) & (g780) & (g788) & (g821) & (g837) & (!g855)));
	assign g947 = (((!g869) & (!g733) & (!g686) & (!g734) & (!g870) & (!g863)) + ((!g869) & (!g733) & (!g686) & (!g734) & (!g870) & (g863)) + ((!g869) & (!g733) & (!g686) & (!g734) & (g870) & (!g863)) + ((!g869) & (!g733) & (!g686) & (!g734) & (g870) & (g863)) + ((!g869) & (!g733) & (!g686) & (g734) & (g870) & (!g863)) + ((!g869) & (!g733) & (!g686) & (g734) & (g870) & (g863)) + ((!g869) & (!g733) & (g686) & (!g734) & (!g870) & (!g863)) + ((!g869) & (!g733) & (g686) & (!g734) & (!g870) & (g863)) + ((!g869) & (!g733) & (g686) & (!g734) & (g870) & (!g863)) + ((!g869) & (!g733) & (g686) & (!g734) & (g870) & (g863)) + ((!g869) & (!g733) & (g686) & (g734) & (g870) & (!g863)) + ((!g869) & (!g733) & (g686) & (g734) & (g870) & (g863)) + ((!g869) & (g733) & (!g686) & (!g734) & (!g870) & (!g863)) + ((!g869) & (g733) & (!g686) & (!g734) & (g870) & (!g863)) + ((!g869) & (g733) & (!g686) & (g734) & (g870) & (!g863)) + ((!g869) & (g733) & (g686) & (!g734) & (!g870) & (!g863)) + ((!g869) & (g733) & (g686) & (!g734) & (g870) & (!g863)) + ((!g869) & (g733) & (g686) & (g734) & (g870) & (!g863)) + ((g869) & (!g733) & (!g686) & (!g734) & (!g870) & (!g863)) + ((g869) & (!g733) & (!g686) & (!g734) & (!g870) & (g863)) + ((g869) & (!g733) & (!g686) & (!g734) & (g870) & (!g863)) + ((g869) & (!g733) & (!g686) & (!g734) & (g870) & (g863)) + ((g869) & (!g733) & (!g686) & (g734) & (g870) & (!g863)) + ((g869) & (!g733) & (!g686) & (g734) & (g870) & (g863)) + ((g869) & (g733) & (!g686) & (!g734) & (!g870) & (!g863)) + ((g869) & (g733) & (!g686) & (!g734) & (g870) & (!g863)) + ((g869) & (g733) & (!g686) & (g734) & (g870) & (!g863)));
	assign g948 = (((!g838) & (!g839) & (!sk[62]) & (!g852) & (g854)) + ((!g838) & (!g839) & (!sk[62]) & (g852) & (g854)) + ((!g838) & (!g839) & (sk[62]) & (g852) & (!g854)) + ((!g838) & (g839) & (!sk[62]) & (!g852) & (g854)) + ((!g838) & (g839) & (!sk[62]) & (g852) & (g854)) + ((!g838) & (g839) & (sk[62]) & (!g852) & (!g854)) + ((g838) & (!g839) & (!sk[62]) & (!g852) & (!g854)) + ((g838) & (!g839) & (!sk[62]) & (!g852) & (g854)) + ((g838) & (!g839) & (!sk[62]) & (g852) & (!g854)) + ((g838) & (!g839) & (!sk[62]) & (g852) & (g854)) + ((g838) & (!g839) & (sk[62]) & (!g852) & (!g854)) + ((g838) & (!g839) & (sk[62]) & (g852) & (!g854)) + ((g838) & (!g839) & (sk[62]) & (g852) & (g854)) + ((g838) & (g839) & (!sk[62]) & (!g852) & (!g854)) + ((g838) & (g839) & (!sk[62]) & (!g852) & (g854)) + ((g838) & (g839) & (!sk[62]) & (g852) & (!g854)) + ((g838) & (g839) & (!sk[62]) & (g852) & (g854)) + ((g838) & (g839) & (sk[62]) & (!g852) & (!g854)) + ((g838) & (g839) & (sk[62]) & (!g852) & (g854)) + ((g838) & (g839) & (sk[62]) & (g852) & (!g854)));
	assign g949 = (((!g202) & (!g781) & (!g783) & (!g784) & (!g841) & (g851)) + ((!g202) & (!g781) & (!g783) & (g784) & (!g841) & (!g851)) + ((!g202) & (!g781) & (!g783) & (g784) & (!g841) & (g851)) + ((!g202) & (!g781) & (!g783) & (g784) & (g841) & (g851)) + ((!g202) & (!g781) & (g783) & (!g784) & (!g841) & (g851)) + ((!g202) & (!g781) & (g783) & (g784) & (!g841) & (g851)) + ((!g202) & (g781) & (!g783) & (!g784) & (!g841) & (!g851)) + ((!g202) & (g781) & (!g783) & (!g784) & (!g841) & (g851)) + ((!g202) & (g781) & (!g783) & (!g784) & (g841) & (g851)) + ((!g202) & (g781) & (!g783) & (g784) & (!g841) & (!g851)) + ((!g202) & (g781) & (!g783) & (g784) & (!g841) & (g851)) + ((!g202) & (g781) & (!g783) & (g784) & (g841) & (g851)) + ((!g202) & (g781) & (g783) & (!g784) & (!g841) & (g851)) + ((!g202) & (g781) & (g783) & (g784) & (!g841) & (!g851)) + ((!g202) & (g781) & (g783) & (g784) & (!g841) & (g851)) + ((!g202) & (g781) & (g783) & (g784) & (g841) & (g851)) + ((g202) & (!g781) & (!g783) & (!g784) & (g841) & (g851)) + ((g202) & (!g781) & (!g783) & (g784) & (!g841) & (g851)) + ((g202) & (!g781) & (!g783) & (g784) & (g841) & (!g851)) + ((g202) & (!g781) & (!g783) & (g784) & (g841) & (g851)) + ((g202) & (!g781) & (g783) & (!g784) & (g841) & (g851)) + ((g202) & (!g781) & (g783) & (g784) & (g841) & (g851)) + ((g202) & (g781) & (!g783) & (!g784) & (!g841) & (g851)) + ((g202) & (g781) & (!g783) & (!g784) & (g841) & (!g851)) + ((g202) & (g781) & (!g783) & (!g784) & (g841) & (g851)) + ((g202) & (g781) & (!g783) & (g784) & (!g841) & (g851)) + ((g202) & (g781) & (!g783) & (g784) & (g841) & (!g851)) + ((g202) & (g781) & (!g783) & (g784) & (g841) & (g851)) + ((g202) & (g781) & (g783) & (!g784) & (g841) & (g851)) + ((g202) & (g781) & (g783) & (g784) & (!g841) & (g851)) + ((g202) & (g781) & (g783) & (g784) & (g841) & (!g851)) + ((g202) & (g781) & (g783) & (g784) & (g841) & (g851)));
	assign g950 = (((!g585) & (!g597) & (!g679) & (g720) & (!g764) & (g762)) + ((!g585) & (!g597) & (!g679) & (g720) & (g764) & (g762)) + ((!g585) & (!g597) & (g679) & (!g720) & (g764) & (!g762)) + ((!g585) & (!g597) & (g679) & (!g720) & (g764) & (g762)) + ((!g585) & (!g597) & (g679) & (g720) & (!g764) & (g762)) + ((!g585) & (!g597) & (g679) & (g720) & (g764) & (!g762)) + ((!g585) & (!g597) & (g679) & (g720) & (g764) & (g762)) + ((!g585) & (g597) & (!g679) & (!g720) & (g764) & (!g762)) + ((!g585) & (g597) & (!g679) & (!g720) & (g764) & (g762)) + ((!g585) & (g597) & (!g679) & (g720) & (!g764) & (g762)) + ((!g585) & (g597) & (!g679) & (g720) & (g764) & (!g762)) + ((!g585) & (g597) & (!g679) & (g720) & (g764) & (g762)) + ((!g585) & (g597) & (g679) & (g720) & (!g764) & (g762)) + ((!g585) & (g597) & (g679) & (g720) & (g764) & (g762)) + ((g585) & (!g597) & (!g679) & (!g720) & (g764) & (!g762)) + ((g585) & (!g597) & (!g679) & (!g720) & (g764) & (g762)) + ((g585) & (!g597) & (!g679) & (g720) & (!g764) & (g762)) + ((g585) & (!g597) & (!g679) & (g720) & (g764) & (!g762)) + ((g585) & (!g597) & (!g679) & (g720) & (g764) & (g762)) + ((g585) & (!g597) & (g679) & (g720) & (!g764) & (g762)) + ((g585) & (!g597) & (g679) & (g720) & (g764) & (g762)) + ((g585) & (g597) & (!g679) & (g720) & (!g764) & (g762)) + ((g585) & (g597) & (!g679) & (g720) & (g764) & (g762)) + ((g585) & (g597) & (g679) & (!g720) & (g764) & (!g762)) + ((g585) & (g597) & (g679) & (!g720) & (g764) & (g762)) + ((g585) & (g597) & (g679) & (g720) & (!g764) & (g762)) + ((g585) & (g597) & (g679) & (g720) & (g764) & (!g762)) + ((g585) & (g597) & (g679) & (g720) & (g764) & (g762)));
	assign g951 = (((!g202) & (!g722) & (!g759) & (!g765) & (!g771) & (g950)) + ((!g202) & (!g722) & (!g759) & (!g765) & (g771) & (g950)) + ((!g202) & (!g722) & (!g759) & (g765) & (!g771) & (!g950)) + ((!g202) & (!g722) & (!g759) & (g765) & (!g771) & (g950)) + ((!g202) & (!g722) & (!g759) & (g765) & (g771) & (!g950)) + ((!g202) & (!g722) & (!g759) & (g765) & (g771) & (g950)) + ((!g202) & (!g722) & (g759) & (!g765) & (!g771) & (!g950)) + ((!g202) & (!g722) & (g759) & (!g765) & (!g771) & (g950)) + ((!g202) & (!g722) & (g759) & (!g765) & (g771) & (g950)) + ((!g202) & (!g722) & (g759) & (g765) & (!g771) & (!g950)) + ((!g202) & (!g722) & (g759) & (g765) & (!g771) & (g950)) + ((!g202) & (!g722) & (g759) & (g765) & (g771) & (!g950)) + ((!g202) & (!g722) & (g759) & (g765) & (g771) & (g950)) + ((!g202) & (g722) & (!g759) & (!g765) & (!g771) & (g950)) + ((!g202) & (g722) & (!g759) & (!g765) & (g771) & (g950)) + ((!g202) & (g722) & (!g759) & (g765) & (!g771) & (g950)) + ((!g202) & (g722) & (!g759) & (g765) & (g771) & (g950)) + ((!g202) & (g722) & (g759) & (!g765) & (!g771) & (!g950)) + ((!g202) & (g722) & (g759) & (!g765) & (!g771) & (g950)) + ((!g202) & (g722) & (g759) & (!g765) & (g771) & (g950)) + ((!g202) & (g722) & (g759) & (g765) & (!g771) & (!g950)) + ((!g202) & (g722) & (g759) & (g765) & (!g771) & (g950)) + ((!g202) & (g722) & (g759) & (g765) & (g771) & (g950)) + ((g202) & (!g722) & (!g759) & (!g765) & (!g771) & (!g950)) + ((g202) & (!g722) & (!g759) & (!g765) & (g771) & (!g950)) + ((g202) & (!g722) & (g759) & (!g765) & (g771) & (!g950)) + ((g202) & (g722) & (!g759) & (!g765) & (!g771) & (!g950)) + ((g202) & (g722) & (!g759) & (!g765) & (g771) & (!g950)) + ((g202) & (g722) & (!g759) & (g765) & (!g771) & (!g950)) + ((g202) & (g722) & (!g759) & (g765) & (g771) & (!g950)) + ((g202) & (g722) & (g759) & (!g765) & (g771) & (!g950)) + ((g202) & (g722) & (g759) & (g765) & (g771) & (!g950)));
	assign g952 = (((!sk[66]) & (!g746) & (!g843) & (!g846) & (g849)) + ((!sk[66]) & (!g746) & (!g843) & (g846) & (g849)) + ((!sk[66]) & (!g746) & (g843) & (!g846) & (g849)) + ((!sk[66]) & (!g746) & (g843) & (g846) & (g849)) + ((!sk[66]) & (g746) & (!g843) & (!g846) & (!g849)) + ((!sk[66]) & (g746) & (!g843) & (!g846) & (g849)) + ((!sk[66]) & (g746) & (!g843) & (g846) & (!g849)) + ((!sk[66]) & (g746) & (!g843) & (g846) & (g849)) + ((!sk[66]) & (g746) & (g843) & (!g846) & (!g849)) + ((!sk[66]) & (g746) & (g843) & (!g846) & (g849)) + ((!sk[66]) & (g746) & (g843) & (g846) & (!g849)) + ((!sk[66]) & (g746) & (g843) & (g846) & (g849)) + ((sk[66]) & (!g746) & (!g843) & (!g846) & (!g849)) + ((sk[66]) & (g746) & (!g843) & (!g846) & (!g849)) + ((sk[66]) & (g746) & (g843) & (!g846) & (!g849)));
	assign g953 = (((!g723) & (!g724) & (!g725) & (!sk[67]) & (g726) & (!g843)) + ((!g723) & (!g724) & (!g725) & (!sk[67]) & (g726) & (g843)) + ((!g723) & (!g724) & (!g725) & (sk[67]) & (g726) & (g843)) + ((!g723) & (!g724) & (g725) & (!sk[67]) & (!g726) & (!g843)) + ((!g723) & (!g724) & (g725) & (!sk[67]) & (!g726) & (g843)) + ((!g723) & (!g724) & (g725) & (!sk[67]) & (g726) & (!g843)) + ((!g723) & (!g724) & (g725) & (!sk[67]) & (g726) & (g843)) + ((!g723) & (!g724) & (g725) & (sk[67]) & (g726) & (g843)) + ((!g723) & (g724) & (!g725) & (!sk[67]) & (!g726) & (!g843)) + ((!g723) & (g724) & (!g725) & (!sk[67]) & (!g726) & (g843)) + ((!g723) & (g724) & (!g725) & (!sk[67]) & (g726) & (!g843)) + ((!g723) & (g724) & (!g725) & (!sk[67]) & (g726) & (g843)) + ((!g723) & (g724) & (!g725) & (sk[67]) & (!g726) & (g843)) + ((!g723) & (g724) & (g725) & (!sk[67]) & (!g726) & (!g843)) + ((!g723) & (g724) & (g725) & (!sk[67]) & (!g726) & (g843)) + ((!g723) & (g724) & (g725) & (!sk[67]) & (g726) & (!g843)) + ((!g723) & (g724) & (g725) & (!sk[67]) & (g726) & (g843)) + ((!g723) & (g724) & (g725) & (sk[67]) & (!g726) & (g843)) + ((!g723) & (g724) & (g725) & (sk[67]) & (g726) & (g843)) + ((g723) & (!g724) & (!g725) & (!sk[67]) & (g726) & (!g843)) + ((g723) & (!g724) & (!g725) & (!sk[67]) & (g726) & (g843)) + ((g723) & (!g724) & (!g725) & (sk[67]) & (!g726) & (g843)) + ((g723) & (!g724) & (g725) & (!sk[67]) & (!g726) & (!g843)) + ((g723) & (!g724) & (g725) & (!sk[67]) & (!g726) & (g843)) + ((g723) & (!g724) & (g725) & (!sk[67]) & (g726) & (!g843)) + ((g723) & (!g724) & (g725) & (!sk[67]) & (g726) & (g843)) + ((g723) & (!g724) & (g725) & (sk[67]) & (!g726) & (g843)) + ((g723) & (g724) & (!g725) & (!sk[67]) & (!g726) & (!g843)) + ((g723) & (g724) & (!g725) & (!sk[67]) & (!g726) & (g843)) + ((g723) & (g724) & (!g725) & (!sk[67]) & (g726) & (!g843)) + ((g723) & (g724) & (!g725) & (!sk[67]) & (g726) & (g843)) + ((g723) & (g724) & (!g725) & (sk[67]) & (g726) & (g843)) + ((g723) & (g724) & (g725) & (!sk[67]) & (!g726) & (!g843)) + ((g723) & (g724) & (g725) & (!sk[67]) & (!g726) & (g843)) + ((g723) & (g724) & (g725) & (!sk[67]) & (g726) & (!g843)) + ((g723) & (g724) & (g725) & (!sk[67]) & (g726) & (g843)));
	assign g954 = (((!g723) & (!g724) & (!g726) & (!g847) & (!g845) & (!g848)) + ((!g723) & (!g724) & (!g726) & (!g847) & (!g845) & (g848)) + ((!g723) & (!g724) & (g726) & (!g847) & (!g845) & (!g848)) + ((!g723) & (g724) & (!g726) & (!g847) & (!g845) & (!g848)) + ((!g723) & (g724) & (!g726) & (!g847) & (!g845) & (g848)) + ((!g723) & (g724) & (!g726) & (!g847) & (g845) & (!g848)) + ((!g723) & (g724) & (!g726) & (!g847) & (g845) & (g848)) + ((!g723) & (g724) & (g726) & (!g847) & (!g845) & (!g848)) + ((!g723) & (g724) & (g726) & (!g847) & (g845) & (!g848)) + ((g723) & (!g724) & (!g726) & (!g847) & (!g845) & (!g848)) + ((g723) & (!g724) & (!g726) & (!g847) & (!g845) & (g848)) + ((g723) & (!g724) & (!g726) & (g847) & (!g845) & (!g848)) + ((g723) & (!g724) & (!g726) & (g847) & (!g845) & (g848)) + ((g723) & (!g724) & (g726) & (!g847) & (!g845) & (!g848)) + ((g723) & (!g724) & (g726) & (g847) & (!g845) & (!g848)) + ((g723) & (g724) & (!g726) & (!g847) & (!g845) & (!g848)) + ((g723) & (g724) & (!g726) & (!g847) & (!g845) & (g848)) + ((g723) & (g724) & (!g726) & (!g847) & (g845) & (!g848)) + ((g723) & (g724) & (!g726) & (!g847) & (g845) & (g848)) + ((g723) & (g724) & (!g726) & (g847) & (!g845) & (!g848)) + ((g723) & (g724) & (!g726) & (g847) & (!g845) & (g848)) + ((g723) & (g724) & (!g726) & (g847) & (g845) & (!g848)) + ((g723) & (g724) & (!g726) & (g847) & (g845) & (g848)) + ((g723) & (g724) & (g726) & (!g847) & (!g845) & (!g848)) + ((g723) & (g724) & (g726) & (!g847) & (g845) & (!g848)) + ((g723) & (g724) & (g726) & (g847) & (!g845) & (!g848)) + ((g723) & (g724) & (g726) & (g847) & (g845) & (!g848)));
	assign g955 = (((!g252) & (!g725) & (!g952) & (!g850) & (!g953) & (g954)) + ((!g252) & (!g725) & (!g952) & (g850) & (!g953) & (g954)) + ((!g252) & (!g725) & (g952) & (!g850) & (!g953) & (g954)) + ((!g252) & (!g725) & (g952) & (g850) & (!g953) & (g954)) + ((!g252) & (g725) & (!g952) & (!g850) & (!g953) & (g954)) + ((!g252) & (g725) & (!g952) & (g850) & (!g953) & (!g954)) + ((!g252) & (g725) & (!g952) & (g850) & (g953) & (!g954)) + ((!g252) & (g725) & (!g952) & (g850) & (g953) & (g954)) + ((!g252) & (g725) & (g952) & (!g850) & (!g953) & (g954)) + ((!g252) & (g725) & (g952) & (g850) & (!g953) & (g954)) + ((g252) & (!g725) & (!g952) & (!g850) & (!g953) & (g954)) + ((g252) & (!g725) & (!g952) & (g850) & (!g953) & (g954)) + ((g252) & (!g725) & (g952) & (!g850) & (!g953) & (g954)) + ((g252) & (!g725) & (g952) & (g850) & (!g953) & (!g954)) + ((g252) & (!g725) & (g952) & (g850) & (g953) & (!g954)) + ((g252) & (!g725) & (g952) & (g850) & (g953) & (g954)) + ((g252) & (g725) & (!g952) & (!g850) & (!g953) & (!g954)) + ((g252) & (g725) & (!g952) & (!g850) & (g953) & (!g954)) + ((g252) & (g725) & (!g952) & (!g850) & (g953) & (g954)) + ((g252) & (g725) & (!g952) & (g850) & (!g953) & (!g954)) + ((g252) & (g725) & (!g952) & (g850) & (g953) & (!g954)) + ((g252) & (g725) & (!g952) & (g850) & (g953) & (g954)) + ((g252) & (g725) & (g952) & (!g850) & (!g953) & (!g954)) + ((g252) & (g725) & (g952) & (!g850) & (g953) & (!g954)) + ((g252) & (g725) & (g952) & (!g850) & (g953) & (g954)) + ((g252) & (g725) & (g952) & (g850) & (!g953) & (g954)));
	assign g956 = (((!g949) & (!g951) & (sk[70]) & (!g955)) + ((!g949) & (g951) & (!sk[70]) & (!g955)) + ((!g949) & (g951) & (!sk[70]) & (g955)) + ((!g949) & (g951) & (sk[70]) & (g955)) + ((g949) & (!g951) & (sk[70]) & (g955)) + ((g949) & (g951) & (!sk[70]) & (!g955)) + ((g949) & (g951) & (!sk[70]) & (g955)) + ((g949) & (g951) & (sk[70]) & (!g955)));
	assign g957 = (((!g708) & (!g716) & (!g549) & (!g569) & (!g680) & (g747)) + ((!g708) & (!g716) & (g549) & (!g569) & (!g680) & (g747)) + ((!g708) & (!g716) & (g549) & (!g569) & (g680) & (g747)) + ((!g708) & (!g716) & (g549) & (g569) & (!g680) & (g747)) + ((!g708) & (g716) & (!g549) & (!g569) & (g680) & (g747)) + ((!g708) & (g716) & (!g549) & (g569) & (!g680) & (g747)) + ((!g708) & (g716) & (!g549) & (g569) & (g680) & (g747)) + ((!g708) & (g716) & (g549) & (g569) & (g680) & (g747)) + ((g708) & (!g716) & (!g549) & (!g569) & (g680) & (g747)) + ((g708) & (!g716) & (!g549) & (g569) & (!g680) & (g747)) + ((g708) & (!g716) & (!g549) & (g569) & (g680) & (g747)) + ((g708) & (!g716) & (g549) & (g569) & (g680) & (g747)) + ((g708) & (g716) & (!g549) & (!g569) & (!g680) & (g747)) + ((g708) & (g716) & (g549) & (!g569) & (!g680) & (g747)) + ((g708) & (g716) & (g549) & (!g569) & (g680) & (g747)) + ((g708) & (g716) & (g549) & (g569) & (!g680) & (g747)));
	assign g958 = (((!g549) & (!g569) & (!g680) & (!g729) & (!g744) & (g748)) + ((!g549) & (!g569) & (!g680) & (!g729) & (g744) & (g748)) + ((!g549) & (!g569) & (g680) & (!g729) & (!g744) & (g748)) + ((!g549) & (!g569) & (g680) & (!g729) & (g744) & (!g748)) + ((!g549) & (!g569) & (g680) & (!g729) & (g744) & (g748)) + ((!g549) & (!g569) & (g680) & (g729) & (g744) & (!g748)) + ((!g549) & (!g569) & (g680) & (g729) & (g744) & (g748)) + ((!g549) & (g569) & (!g680) & (!g729) & (!g744) & (g748)) + ((!g549) & (g569) & (!g680) & (!g729) & (g744) & (!g748)) + ((!g549) & (g569) & (!g680) & (!g729) & (g744) & (g748)) + ((!g549) & (g569) & (!g680) & (g729) & (g744) & (!g748)) + ((!g549) & (g569) & (!g680) & (g729) & (g744) & (g748)) + ((!g549) & (g569) & (g680) & (!g729) & (!g744) & (g748)) + ((!g549) & (g569) & (g680) & (!g729) & (g744) & (g748)) + ((g549) & (!g569) & (!g680) & (!g729) & (!g744) & (g748)) + ((g549) & (!g569) & (!g680) & (!g729) & (g744) & (!g748)) + ((g549) & (!g569) & (!g680) & (!g729) & (g744) & (g748)) + ((g549) & (!g569) & (!g680) & (g729) & (g744) & (!g748)) + ((g549) & (!g569) & (!g680) & (g729) & (g744) & (g748)) + ((g549) & (!g569) & (g680) & (!g729) & (!g744) & (g748)) + ((g549) & (!g569) & (g680) & (!g729) & (g744) & (g748)) + ((g549) & (g569) & (!g680) & (!g729) & (!g744) & (g748)) + ((g549) & (g569) & (!g680) & (!g729) & (g744) & (g748)) + ((g549) & (g569) & (g680) & (!g729) & (!g744) & (g748)) + ((g549) & (g569) & (g680) & (!g729) & (g744) & (!g748)) + ((g549) & (g569) & (g680) & (!g729) & (g744) & (g748)) + ((g549) & (g569) & (g680) & (g729) & (g744) & (!g748)) + ((g549) & (g569) & (g680) & (g729) & (g744) & (g748)));
	assign g959 = (((!g200) & (!g730) & (!g816) & (!g742) & (!g957) & (!g958)) + ((!g200) & (!g730) & (g816) & (!g742) & (!g957) & (!g958)) + ((!g200) & (!g730) & (g816) & (g742) & (!g957) & (!g958)) + ((!g200) & (g730) & (!g816) & (!g742) & (!g957) & (!g958)) + ((!g200) & (g730) & (!g816) & (g742) & (!g957) & (!g958)) + ((!g200) & (g730) & (g816) & (!g742) & (!g957) & (!g958)) + ((g200) & (!g730) & (!g816) & (!g742) & (!g957) & (g958)) + ((g200) & (!g730) & (!g816) & (!g742) & (g957) & (!g958)) + ((g200) & (!g730) & (!g816) & (!g742) & (g957) & (g958)) + ((g200) & (!g730) & (!g816) & (g742) & (!g957) & (!g958)) + ((g200) & (!g730) & (!g816) & (g742) & (!g957) & (g958)) + ((g200) & (!g730) & (!g816) & (g742) & (g957) & (!g958)) + ((g200) & (!g730) & (!g816) & (g742) & (g957) & (g958)) + ((g200) & (!g730) & (g816) & (!g742) & (!g957) & (g958)) + ((g200) & (!g730) & (g816) & (!g742) & (g957) & (!g958)) + ((g200) & (!g730) & (g816) & (!g742) & (g957) & (g958)) + ((g200) & (!g730) & (g816) & (g742) & (!g957) & (g958)) + ((g200) & (!g730) & (g816) & (g742) & (g957) & (!g958)) + ((g200) & (!g730) & (g816) & (g742) & (g957) & (g958)) + ((g200) & (g730) & (!g816) & (!g742) & (!g957) & (g958)) + ((g200) & (g730) & (!g816) & (!g742) & (g957) & (!g958)) + ((g200) & (g730) & (!g816) & (!g742) & (g957) & (g958)) + ((g200) & (g730) & (!g816) & (g742) & (!g957) & (g958)) + ((g200) & (g730) & (!g816) & (g742) & (g957) & (!g958)) + ((g200) & (g730) & (!g816) & (g742) & (g957) & (g958)) + ((g200) & (g730) & (g816) & (!g742) & (!g957) & (g958)) + ((g200) & (g730) & (g816) & (!g742) & (g957) & (!g958)) + ((g200) & (g730) & (g816) & (!g742) & (g957) & (g958)) + ((g200) & (g730) & (g816) & (g742) & (!g957) & (!g958)) + ((g200) & (g730) & (g816) & (g742) & (!g957) & (g958)) + ((g200) & (g730) & (g816) & (g742) & (g957) & (!g958)) + ((g200) & (g730) & (g816) & (g742) & (g957) & (g958)));
	assign g960 = (((!g956) & (sk[74]) & (g959)) + ((g956) & (!sk[74]) & (g959)) + ((g956) & (sk[74]) & (!g959)));
	assign g961 = (((!g2) & (!g732) & (!g899) & (!g947) & (!g948) & (!g960)) + ((!g2) & (!g732) & (!g899) & (!g947) & (g948) & (g960)) + ((!g2) & (!g732) & (!g899) & (g947) & (!g948) & (g960)) + ((!g2) & (!g732) & (!g899) & (g947) & (g948) & (!g960)) + ((!g2) & (!g732) & (g899) & (!g947) & (!g948) & (!g960)) + ((!g2) & (!g732) & (g899) & (!g947) & (g948) & (g960)) + ((!g2) & (!g732) & (g899) & (g947) & (!g948) & (g960)) + ((!g2) & (!g732) & (g899) & (g947) & (g948) & (!g960)) + ((!g2) & (g732) & (!g899) & (!g947) & (!g948) & (!g960)) + ((!g2) & (g732) & (!g899) & (!g947) & (g948) & (g960)) + ((!g2) & (g732) & (!g899) & (g947) & (!g948) & (!g960)) + ((!g2) & (g732) & (!g899) & (g947) & (g948) & (g960)) + ((!g2) & (g732) & (g899) & (!g947) & (!g948) & (!g960)) + ((!g2) & (g732) & (g899) & (!g947) & (g948) & (g960)) + ((!g2) & (g732) & (g899) & (g947) & (!g948) & (g960)) + ((!g2) & (g732) & (g899) & (g947) & (g948) & (!g960)) + ((g2) & (!g732) & (!g899) & (!g947) & (!g948) & (g960)) + ((g2) & (!g732) & (!g899) & (!g947) & (g948) & (!g960)) + ((g2) & (!g732) & (!g899) & (g947) & (!g948) & (!g960)) + ((g2) & (!g732) & (!g899) & (g947) & (g948) & (g960)) + ((g2) & (!g732) & (g899) & (!g947) & (!g948) & (g960)) + ((g2) & (!g732) & (g899) & (!g947) & (g948) & (!g960)) + ((g2) & (!g732) & (g899) & (g947) & (!g948) & (!g960)) + ((g2) & (!g732) & (g899) & (g947) & (g948) & (g960)) + ((g2) & (g732) & (!g899) & (!g947) & (!g948) & (g960)) + ((g2) & (g732) & (!g899) & (!g947) & (g948) & (!g960)) + ((g2) & (g732) & (!g899) & (g947) & (!g948) & (g960)) + ((g2) & (g732) & (!g899) & (g947) & (g948) & (!g960)) + ((g2) & (g732) & (g899) & (!g947) & (!g948) & (g960)) + ((g2) & (g732) & (g899) & (!g947) & (g948) & (!g960)) + ((g2) & (g732) & (g899) & (g947) & (!g948) & (!g960)) + ((g2) & (g732) & (g899) & (g947) & (g948) & (g960)));
	assign g962 = (((!sk[76]) & (!g889) & (g871) & (!g883)) + ((!sk[76]) & (!g889) & (g871) & (g883)) + ((!sk[76]) & (g889) & (g871) & (!g883)) + ((!sk[76]) & (g889) & (g871) & (g883)) + ((sk[76]) & (!g889) & (g871) & (g883)) + ((sk[76]) & (g889) & (!g871) & (!g883)) + ((sk[76]) & (g889) & (!g871) & (g883)) + ((sk[76]) & (g889) & (g871) & (!g883)));
	assign g963 = (((!sk[77]) & (g871) & (g883)) + ((sk[77]) & (!g871) & (!g883)) + ((sk[77]) & (g871) & (g883)));
	assign g964 = (((!sk[78]) & (!g193) & (!g272) & (!g147) & (g194) & (!g601)) + ((!sk[78]) & (!g193) & (!g272) & (!g147) & (g194) & (g601)) + ((!sk[78]) & (!g193) & (!g272) & (g147) & (!g194) & (!g601)) + ((!sk[78]) & (!g193) & (!g272) & (g147) & (!g194) & (g601)) + ((!sk[78]) & (!g193) & (!g272) & (g147) & (g194) & (!g601)) + ((!sk[78]) & (!g193) & (!g272) & (g147) & (g194) & (g601)) + ((!sk[78]) & (!g193) & (g272) & (!g147) & (!g194) & (!g601)) + ((!sk[78]) & (!g193) & (g272) & (!g147) & (!g194) & (g601)) + ((!sk[78]) & (!g193) & (g272) & (!g147) & (g194) & (!g601)) + ((!sk[78]) & (!g193) & (g272) & (!g147) & (g194) & (g601)) + ((!sk[78]) & (!g193) & (g272) & (g147) & (!g194) & (!g601)) + ((!sk[78]) & (!g193) & (g272) & (g147) & (!g194) & (g601)) + ((!sk[78]) & (!g193) & (g272) & (g147) & (g194) & (!g601)) + ((!sk[78]) & (!g193) & (g272) & (g147) & (g194) & (g601)) + ((!sk[78]) & (g193) & (!g272) & (!g147) & (g194) & (!g601)) + ((!sk[78]) & (g193) & (!g272) & (!g147) & (g194) & (g601)) + ((!sk[78]) & (g193) & (!g272) & (g147) & (!g194) & (!g601)) + ((!sk[78]) & (g193) & (!g272) & (g147) & (!g194) & (g601)) + ((!sk[78]) & (g193) & (!g272) & (g147) & (g194) & (!g601)) + ((!sk[78]) & (g193) & (!g272) & (g147) & (g194) & (g601)) + ((!sk[78]) & (g193) & (g272) & (!g147) & (!g194) & (!g601)) + ((!sk[78]) & (g193) & (g272) & (!g147) & (!g194) & (g601)) + ((!sk[78]) & (g193) & (g272) & (!g147) & (g194) & (!g601)) + ((!sk[78]) & (g193) & (g272) & (!g147) & (g194) & (g601)) + ((!sk[78]) & (g193) & (g272) & (g147) & (!g194) & (!g601)) + ((!sk[78]) & (g193) & (g272) & (g147) & (!g194) & (g601)) + ((!sk[78]) & (g193) & (g272) & (g147) & (g194) & (!g601)) + ((!sk[78]) & (g193) & (g272) & (g147) & (g194) & (g601)) + ((sk[78]) & (!g193) & (!g272) & (!g147) & (!g194) & (!g601)));
	assign g965 = (((!g99) & (!g18) & (!sk[79]) & (!g105) & (g141) & (!g964)) + ((!g99) & (!g18) & (!sk[79]) & (!g105) & (g141) & (g964)) + ((!g99) & (!g18) & (!sk[79]) & (g105) & (!g141) & (!g964)) + ((!g99) & (!g18) & (!sk[79]) & (g105) & (!g141) & (g964)) + ((!g99) & (!g18) & (!sk[79]) & (g105) & (g141) & (!g964)) + ((!g99) & (!g18) & (!sk[79]) & (g105) & (g141) & (g964)) + ((!g99) & (!g18) & (sk[79]) & (!g105) & (!g141) & (g964)) + ((!g99) & (g18) & (!sk[79]) & (!g105) & (!g141) & (!g964)) + ((!g99) & (g18) & (!sk[79]) & (!g105) & (!g141) & (g964)) + ((!g99) & (g18) & (!sk[79]) & (!g105) & (g141) & (!g964)) + ((!g99) & (g18) & (!sk[79]) & (!g105) & (g141) & (g964)) + ((!g99) & (g18) & (!sk[79]) & (g105) & (!g141) & (!g964)) + ((!g99) & (g18) & (!sk[79]) & (g105) & (!g141) & (g964)) + ((!g99) & (g18) & (!sk[79]) & (g105) & (g141) & (!g964)) + ((!g99) & (g18) & (!sk[79]) & (g105) & (g141) & (g964)) + ((!g99) & (g18) & (sk[79]) & (!g105) & (!g141) & (g964)) + ((g99) & (!g18) & (!sk[79]) & (!g105) & (g141) & (!g964)) + ((g99) & (!g18) & (!sk[79]) & (!g105) & (g141) & (g964)) + ((g99) & (!g18) & (!sk[79]) & (g105) & (!g141) & (!g964)) + ((g99) & (!g18) & (!sk[79]) & (g105) & (!g141) & (g964)) + ((g99) & (!g18) & (!sk[79]) & (g105) & (g141) & (!g964)) + ((g99) & (!g18) & (!sk[79]) & (g105) & (g141) & (g964)) + ((g99) & (!g18) & (sk[79]) & (!g105) & (!g141) & (g964)) + ((g99) & (g18) & (!sk[79]) & (!g105) & (!g141) & (!g964)) + ((g99) & (g18) & (!sk[79]) & (!g105) & (!g141) & (g964)) + ((g99) & (g18) & (!sk[79]) & (!g105) & (g141) & (!g964)) + ((g99) & (g18) & (!sk[79]) & (!g105) & (g141) & (g964)) + ((g99) & (g18) & (!sk[79]) & (g105) & (!g141) & (!g964)) + ((g99) & (g18) & (!sk[79]) & (g105) & (!g141) & (g964)) + ((g99) & (g18) & (!sk[79]) & (g105) & (g141) & (!g964)) + ((g99) & (g18) & (!sk[79]) & (g105) & (g141) & (g964)));
	assign g966 = (((!g80) & (g885) & (!sk[80]) & (!g965)) + ((!g80) & (g885) & (!sk[80]) & (g965)) + ((!g80) & (g885) & (sk[80]) & (g965)) + ((g80) & (g885) & (!sk[80]) & (!g965)) + ((g80) & (g885) & (!sk[80]) & (g965)));
	assign g967 = (((!g16) & (g12) & (!sk[81]) & (!g18)) + ((!g16) & (g12) & (!sk[81]) & (g18)) + ((g16) & (!g12) & (sk[81]) & (g18)) + ((g16) & (g12) & (!sk[81]) & (!g18)) + ((g16) & (g12) & (!sk[81]) & (g18)) + ((g16) & (g12) & (sk[81]) & (!g18)) + ((g16) & (g12) & (sk[81]) & (g18)));
	assign g968 = (((!sk[82]) & (!g203) & (!g359) & (!g665) & (g967)) + ((!sk[82]) & (!g203) & (!g359) & (g665) & (g967)) + ((!sk[82]) & (!g203) & (g359) & (!g665) & (g967)) + ((!sk[82]) & (!g203) & (g359) & (g665) & (g967)) + ((!sk[82]) & (g203) & (!g359) & (!g665) & (!g967)) + ((!sk[82]) & (g203) & (!g359) & (!g665) & (g967)) + ((!sk[82]) & (g203) & (!g359) & (g665) & (!g967)) + ((!sk[82]) & (g203) & (!g359) & (g665) & (g967)) + ((!sk[82]) & (g203) & (g359) & (!g665) & (!g967)) + ((!sk[82]) & (g203) & (g359) & (!g665) & (g967)) + ((!sk[82]) & (g203) & (g359) & (g665) & (!g967)) + ((!sk[82]) & (g203) & (g359) & (g665) & (g967)) + ((sk[82]) & (!g203) & (!g359) & (!g665) & (!g967)));
	assign g969 = (((!g48) & (!g52) & (!g34) & (g37) & (!sk[83]) & (!g65)) + ((!g48) & (!g52) & (!g34) & (g37) & (!sk[83]) & (g65)) + ((!g48) & (!g52) & (g34) & (!g37) & (!sk[83]) & (!g65)) + ((!g48) & (!g52) & (g34) & (!g37) & (!sk[83]) & (g65)) + ((!g48) & (!g52) & (g34) & (g37) & (!sk[83]) & (!g65)) + ((!g48) & (!g52) & (g34) & (g37) & (!sk[83]) & (g65)) + ((!g48) & (g52) & (!g34) & (!g37) & (!sk[83]) & (!g65)) + ((!g48) & (g52) & (!g34) & (!g37) & (!sk[83]) & (g65)) + ((!g48) & (g52) & (!g34) & (g37) & (!sk[83]) & (!g65)) + ((!g48) & (g52) & (!g34) & (g37) & (!sk[83]) & (g65)) + ((!g48) & (g52) & (g34) & (!g37) & (!sk[83]) & (!g65)) + ((!g48) & (g52) & (g34) & (!g37) & (!sk[83]) & (g65)) + ((!g48) & (g52) & (g34) & (g37) & (!sk[83]) & (!g65)) + ((!g48) & (g52) & (g34) & (g37) & (!sk[83]) & (g65)) + ((g48) & (!g52) & (!g34) & (g37) & (!sk[83]) & (!g65)) + ((g48) & (!g52) & (!g34) & (g37) & (!sk[83]) & (g65)) + ((g48) & (!g52) & (g34) & (!g37) & (!sk[83]) & (!g65)) + ((g48) & (!g52) & (g34) & (!g37) & (!sk[83]) & (g65)) + ((g48) & (!g52) & (g34) & (g37) & (!sk[83]) & (!g65)) + ((g48) & (!g52) & (g34) & (g37) & (!sk[83]) & (g65)) + ((g48) & (g52) & (!g34) & (!g37) & (!sk[83]) & (!g65)) + ((g48) & (g52) & (!g34) & (!g37) & (!sk[83]) & (g65)) + ((g48) & (g52) & (!g34) & (g37) & (!sk[83]) & (!g65)) + ((g48) & (g52) & (!g34) & (g37) & (!sk[83]) & (g65)) + ((g48) & (g52) & (g34) & (!g37) & (!sk[83]) & (!g65)) + ((g48) & (g52) & (g34) & (!g37) & (!sk[83]) & (g65)) + ((g48) & (g52) & (g34) & (g37) & (!sk[83]) & (!g65)) + ((g48) & (g52) & (g34) & (g37) & (!sk[83]) & (g65)) + ((g48) & (g52) & (g34) & (g37) & (sk[83]) & (g65)));
	assign g970 = (((!g208) & (!g966) & (!sk[84]) & (!g968) & (g969)) + ((!g208) & (!g966) & (!sk[84]) & (g968) & (g969)) + ((!g208) & (g966) & (!sk[84]) & (!g968) & (g969)) + ((!g208) & (g966) & (!sk[84]) & (g968) & (g969)) + ((g208) & (!g966) & (!sk[84]) & (!g968) & (!g969)) + ((g208) & (!g966) & (!sk[84]) & (!g968) & (g969)) + ((g208) & (!g966) & (!sk[84]) & (g968) & (!g969)) + ((g208) & (!g966) & (!sk[84]) & (g968) & (g969)) + ((g208) & (g966) & (!sk[84]) & (!g968) & (!g969)) + ((g208) & (g966) & (!sk[84]) & (!g968) & (g969)) + ((g208) & (g966) & (!sk[84]) & (g968) & (!g969)) + ((g208) & (g966) & (!sk[84]) & (g968) & (g969)) + ((g208) & (g966) & (sk[84]) & (g968) & (g969)));
	assign g971 = (((!sk[85]) & (!g889) & (!g871) & (!g883) & (g970)) + ((!sk[85]) & (!g889) & (!g871) & (g883) & (g970)) + ((!sk[85]) & (!g889) & (g871) & (!g883) & (g970)) + ((!sk[85]) & (!g889) & (g871) & (g883) & (g970)) + ((!sk[85]) & (g889) & (!g871) & (!g883) & (!g970)) + ((!sk[85]) & (g889) & (!g871) & (!g883) & (g970)) + ((!sk[85]) & (g889) & (!g871) & (g883) & (!g970)) + ((!sk[85]) & (g889) & (!g871) & (g883) & (g970)) + ((!sk[85]) & (g889) & (g871) & (!g883) & (!g970)) + ((!sk[85]) & (g889) & (g871) & (!g883) & (g970)) + ((!sk[85]) & (g889) & (g871) & (g883) & (!g970)) + ((!sk[85]) & (g889) & (g871) & (g883) & (g970)) + ((sk[85]) & (!g889) & (!g871) & (!g883) & (!g970)) + ((sk[85]) & (!g889) & (!g871) & (g883) & (!g970)) + ((sk[85]) & (!g889) & (g871) & (!g883) & (!g970)) + ((sk[85]) & (!g889) & (g871) & (g883) & (!g970)) + ((sk[85]) & (g889) & (!g871) & (!g883) & (!g970)) + ((sk[85]) & (g889) & (!g871) & (g883) & (!g970)) + ((sk[85]) & (g889) & (g871) & (!g883) & (!g970)) + ((sk[85]) & (g889) & (g871) & (g883) & (g970)));
	assign g972 = (((!g962) & (!g963) & (!g884) & (!sk[86]) & (g971)) + ((!g962) & (!g963) & (!g884) & (sk[86]) & (g971)) + ((!g962) & (!g963) & (g884) & (!sk[86]) & (g971)) + ((!g962) & (!g963) & (g884) & (sk[86]) & (!g971)) + ((!g962) & (g963) & (!g884) & (!sk[86]) & (g971)) + ((!g962) & (g963) & (!g884) & (sk[86]) & (!g971)) + ((!g962) & (g963) & (g884) & (!sk[86]) & (g971)) + ((!g962) & (g963) & (g884) & (sk[86]) & (!g971)) + ((g962) & (!g963) & (!g884) & (!sk[86]) & (!g971)) + ((g962) & (!g963) & (!g884) & (!sk[86]) & (g971)) + ((g962) & (!g963) & (!g884) & (sk[86]) & (!g971)) + ((g962) & (!g963) & (g884) & (!sk[86]) & (!g971)) + ((g962) & (!g963) & (g884) & (!sk[86]) & (g971)) + ((g962) & (!g963) & (g884) & (sk[86]) & (!g971)) + ((g962) & (g963) & (!g884) & (!sk[86]) & (!g971)) + ((g962) & (g963) & (!g884) & (!sk[86]) & (g971)) + ((g962) & (g963) & (!g884) & (sk[86]) & (!g971)) + ((g962) & (g963) & (g884) & (!sk[86]) & (!g971)) + ((g962) & (g963) & (g884) & (!sk[86]) & (g971)) + ((g962) & (g963) & (g884) & (sk[86]) & (g971)));
	assign g973 = (((!g891) & (!g962) & (!g864) & (!g892) & (!g963) & (!g971)) + ((!g891) & (!g962) & (!g864) & (!g892) & (!g963) & (g971)) + ((!g891) & (!g962) & (!g864) & (!g892) & (g963) & (!g971)) + ((!g891) & (!g962) & (!g864) & (!g892) & (g963) & (g971)) + ((!g891) & (!g962) & (g864) & (!g892) & (!g963) & (!g971)) + ((!g891) & (!g962) & (g864) & (!g892) & (!g963) & (g971)) + ((!g891) & (g962) & (!g864) & (!g892) & (!g963) & (!g971)) + ((!g891) & (g962) & (!g864) & (!g892) & (!g963) & (g971)) + ((!g891) & (g962) & (!g864) & (!g892) & (g963) & (!g971)) + ((!g891) & (g962) & (!g864) & (!g892) & (g963) & (g971)) + ((!g891) & (g962) & (!g864) & (g892) & (!g963) & (!g971)) + ((!g891) & (g962) & (!g864) & (g892) & (!g963) & (g971)) + ((!g891) & (g962) & (!g864) & (g892) & (g963) & (!g971)) + ((!g891) & (g962) & (!g864) & (g892) & (g963) & (g971)) + ((!g891) & (g962) & (g864) & (!g892) & (!g963) & (!g971)) + ((!g891) & (g962) & (g864) & (!g892) & (!g963) & (g971)) + ((!g891) & (g962) & (g864) & (g892) & (!g963) & (!g971)) + ((!g891) & (g962) & (g864) & (g892) & (!g963) & (g971)) + ((g891) & (!g962) & (!g864) & (!g892) & (!g963) & (!g971)) + ((g891) & (!g962) & (!g864) & (!g892) & (g963) & (!g971)) + ((g891) & (!g962) & (g864) & (!g892) & (!g963) & (!g971)) + ((g891) & (g962) & (!g864) & (!g892) & (!g963) & (!g971)) + ((g891) & (g962) & (!g864) & (!g892) & (g963) & (!g971)) + ((g891) & (g962) & (!g864) & (g892) & (!g963) & (!g971)) + ((g891) & (g962) & (!g864) & (g892) & (g963) & (!g971)) + ((g891) & (g962) & (g864) & (!g892) & (!g963) & (!g971)) + ((g891) & (g962) & (g864) & (g892) & (!g963) & (!g971)));
	assign g974 = (((!sk[88]) & (!g683) & (!g868) & (!g972) & (g973)) + ((!sk[88]) & (!g683) & (!g868) & (g972) & (g973)) + ((!sk[88]) & (!g683) & (g868) & (!g972) & (g973)) + ((!sk[88]) & (!g683) & (g868) & (g972) & (g973)) + ((!sk[88]) & (g683) & (!g868) & (!g972) & (!g973)) + ((!sk[88]) & (g683) & (!g868) & (!g972) & (g973)) + ((!sk[88]) & (g683) & (!g868) & (g972) & (!g973)) + ((!sk[88]) & (g683) & (!g868) & (g972) & (g973)) + ((!sk[88]) & (g683) & (g868) & (!g972) & (!g973)) + ((!sk[88]) & (g683) & (g868) & (!g972) & (g973)) + ((!sk[88]) & (g683) & (g868) & (g972) & (!g973)) + ((!sk[88]) & (g683) & (g868) & (g972) & (g973)) + ((sk[88]) & (!g683) & (!g868) & (!g972) & (g973)) + ((sk[88]) & (!g683) & (!g868) & (g972) & (g973)) + ((sk[88]) & (!g683) & (g868) & (g972) & (g973)) + ((sk[88]) & (g683) & (!g868) & (!g972) & (!g973)) + ((sk[88]) & (g683) & (!g868) & (g972) & (!g973)) + ((sk[88]) & (g683) & (g868) & (!g972) & (!g973)) + ((sk[88]) & (g683) & (g868) & (!g972) & (g973)) + ((sk[88]) & (g683) & (g868) & (g972) & (!g973)));
	assign g975 = (((!g856) & (!g894) & (!g945) & (!g946) & (!g961) & (!g974)) + ((!g856) & (!g894) & (!g945) & (!g946) & (!g961) & (g974)) + ((!g856) & (!g894) & (!g945) & (!g946) & (g961) & (!g974)) + ((!g856) & (!g894) & (!g945) & (g946) & (!g961) & (!g974)) + ((!g856) & (!g894) & (!g945) & (g946) & (g961) & (!g974)) + ((!g856) & (!g894) & (!g945) & (g946) & (g961) & (g974)) + ((!g856) & (!g894) & (g945) & (!g946) & (!g961) & (!g974)) + ((!g856) & (!g894) & (g945) & (!g946) & (!g961) & (g974)) + ((!g856) & (!g894) & (g945) & (!g946) & (g961) & (!g974)) + ((!g856) & (!g894) & (g945) & (g946) & (!g961) & (!g974)) + ((!g856) & (!g894) & (g945) & (g946) & (g961) & (!g974)) + ((!g856) & (!g894) & (g945) & (g946) & (g961) & (g974)) + ((!g856) & (g894) & (!g945) & (!g946) & (!g961) & (!g974)) + ((!g856) & (g894) & (!g945) & (g946) & (g961) & (!g974)) + ((!g856) & (g894) & (g945) & (!g946) & (!g961) & (!g974)) + ((!g856) & (g894) & (g945) & (!g946) & (!g961) & (g974)) + ((!g856) & (g894) & (g945) & (!g946) & (g961) & (!g974)) + ((!g856) & (g894) & (g945) & (g946) & (!g961) & (!g974)) + ((!g856) & (g894) & (g945) & (g946) & (g961) & (!g974)) + ((!g856) & (g894) & (g945) & (g946) & (g961) & (g974)) + ((g856) & (!g894) & (!g945) & (!g946) & (!g961) & (!g974)) + ((g856) & (!g894) & (!g945) & (g946) & (g961) & (!g974)) + ((g856) & (!g894) & (g945) & (!g946) & (!g961) & (!g974)) + ((g856) & (!g894) & (g945) & (!g946) & (!g961) & (g974)) + ((g856) & (!g894) & (g945) & (!g946) & (g961) & (!g974)) + ((g856) & (!g894) & (g945) & (g946) & (!g961) & (!g974)) + ((g856) & (!g894) & (g945) & (g946) & (g961) & (!g974)) + ((g856) & (!g894) & (g945) & (g946) & (g961) & (g974)) + ((g856) & (g894) & (!g945) & (!g946) & (!g961) & (!g974)) + ((g856) & (g894) & (!g945) & (g946) & (g961) & (!g974)) + ((g856) & (g894) & (g945) & (!g946) & (!g961) & (!g974)) + ((g856) & (g894) & (g945) & (g946) & (g961) & (!g974)));
	assign g976 = (((!g2) & (!g732) & (!g899) & (!sk[90]) & (g947)) + ((!g2) & (!g732) & (!g899) & (sk[90]) & (!g947)) + ((!g2) & (!g732) & (g899) & (!sk[90]) & (g947)) + ((!g2) & (!g732) & (g899) & (sk[90]) & (!g947)) + ((!g2) & (g732) & (!g899) & (!sk[90]) & (g947)) + ((!g2) & (g732) & (!g899) & (sk[90]) & (!g947)) + ((!g2) & (g732) & (!g899) & (sk[90]) & (g947)) + ((!g2) & (g732) & (g899) & (!sk[90]) & (g947)) + ((!g2) & (g732) & (g899) & (sk[90]) & (!g947)) + ((g2) & (!g732) & (!g899) & (!sk[90]) & (!g947)) + ((g2) & (!g732) & (!g899) & (!sk[90]) & (g947)) + ((g2) & (!g732) & (!g899) & (sk[90]) & (g947)) + ((g2) & (!g732) & (g899) & (!sk[90]) & (!g947)) + ((g2) & (!g732) & (g899) & (!sk[90]) & (g947)) + ((g2) & (!g732) & (g899) & (sk[90]) & (g947)) + ((g2) & (g732) & (!g899) & (!sk[90]) & (!g947)) + ((g2) & (g732) & (!g899) & (!sk[90]) & (g947)) + ((g2) & (g732) & (g899) & (!sk[90]) & (!g947)) + ((g2) & (g732) & (g899) & (!sk[90]) & (g947)) + ((g2) & (g732) & (g899) & (sk[90]) & (g947)));
	assign g977 = (((!g733) & (!sk[91]) & (!g686) & (!g870) & (g871) & (!g883)) + ((!g733) & (!sk[91]) & (!g686) & (!g870) & (g871) & (g883)) + ((!g733) & (!sk[91]) & (!g686) & (g870) & (!g871) & (!g883)) + ((!g733) & (!sk[91]) & (!g686) & (g870) & (!g871) & (g883)) + ((!g733) & (!sk[91]) & (!g686) & (g870) & (g871) & (!g883)) + ((!g733) & (!sk[91]) & (!g686) & (g870) & (g871) & (g883)) + ((!g733) & (!sk[91]) & (g686) & (!g870) & (!g871) & (!g883)) + ((!g733) & (!sk[91]) & (g686) & (!g870) & (!g871) & (g883)) + ((!g733) & (!sk[91]) & (g686) & (!g870) & (g871) & (!g883)) + ((!g733) & (!sk[91]) & (g686) & (!g870) & (g871) & (g883)) + ((!g733) & (!sk[91]) & (g686) & (g870) & (!g871) & (!g883)) + ((!g733) & (!sk[91]) & (g686) & (g870) & (!g871) & (g883)) + ((!g733) & (!sk[91]) & (g686) & (g870) & (g871) & (!g883)) + ((!g733) & (!sk[91]) & (g686) & (g870) & (g871) & (g883)) + ((!g733) & (sk[91]) & (g686) & (!g870) & (!g871) & (!g883)) + ((!g733) & (sk[91]) & (g686) & (!g870) & (!g871) & (g883)) + ((!g733) & (sk[91]) & (g686) & (!g870) & (g871) & (!g883)) + ((!g733) & (sk[91]) & (g686) & (!g870) & (g871) & (g883)) + ((g733) & (!sk[91]) & (!g686) & (!g870) & (g871) & (!g883)) + ((g733) & (!sk[91]) & (!g686) & (!g870) & (g871) & (g883)) + ((g733) & (!sk[91]) & (!g686) & (g870) & (!g871) & (!g883)) + ((g733) & (!sk[91]) & (!g686) & (g870) & (!g871) & (g883)) + ((g733) & (!sk[91]) & (!g686) & (g870) & (g871) & (!g883)) + ((g733) & (!sk[91]) & (!g686) & (g870) & (g871) & (g883)) + ((g733) & (!sk[91]) & (g686) & (!g870) & (!g871) & (!g883)) + ((g733) & (!sk[91]) & (g686) & (!g870) & (!g871) & (g883)) + ((g733) & (!sk[91]) & (g686) & (!g870) & (g871) & (!g883)) + ((g733) & (!sk[91]) & (g686) & (!g870) & (g871) & (g883)) + ((g733) & (!sk[91]) & (g686) & (g870) & (!g871) & (!g883)) + ((g733) & (!sk[91]) & (g686) & (g870) & (!g871) & (g883)) + ((g733) & (!sk[91]) & (g686) & (g870) & (g871) & (!g883)) + ((g733) & (!sk[91]) & (g686) & (g870) & (g871) & (g883)) + ((g733) & (sk[91]) & (!g686) & (!g870) & (!g871) & (!g883)) + ((g733) & (sk[91]) & (!g686) & (!g870) & (g871) & (g883)) + ((g733) & (sk[91]) & (!g686) & (g870) & (!g871) & (!g883)) + ((g733) & (sk[91]) & (!g686) & (g870) & (g871) & (g883)) + ((g733) & (sk[91]) & (g686) & (!g870) & (!g871) & (!g883)) + ((g733) & (sk[91]) & (g686) & (!g870) & (!g871) & (g883)) + ((g733) & (sk[91]) & (g686) & (!g870) & (g871) & (!g883)) + ((g733) & (sk[91]) & (g686) & (!g870) & (g871) & (g883)) + ((g733) & (sk[91]) & (g686) & (g870) & (!g871) & (!g883)) + ((g733) & (sk[91]) & (g686) & (g870) & (g871) & (g883)));
	assign g978 = (((!g2) & (!g734) & (!g732) & (!g863) & (!g895) & (g977)) + ((!g2) & (!g734) & (!g732) & (!g863) & (g895) & (g977)) + ((!g2) & (!g734) & (!g732) & (g863) & (!g895) & (g977)) + ((!g2) & (!g734) & (!g732) & (g863) & (g895) & (g977)) + ((!g2) & (!g734) & (g732) & (!g863) & (!g895) & (g977)) + ((!g2) & (!g734) & (g732) & (!g863) & (g895) & (!g977)) + ((!g2) & (!g734) & (g732) & (!g863) & (g895) & (g977)) + ((!g2) & (!g734) & (g732) & (g863) & (!g895) & (g977)) + ((!g2) & (!g734) & (g732) & (g863) & (g895) & (!g977)) + ((!g2) & (!g734) & (g732) & (g863) & (g895) & (g977)) + ((!g2) & (g734) & (!g732) & (!g863) & (!g895) & (g977)) + ((!g2) & (g734) & (!g732) & (!g863) & (g895) & (g977)) + ((!g2) & (g734) & (!g732) & (g863) & (!g895) & (!g977)) + ((!g2) & (g734) & (!g732) & (g863) & (!g895) & (g977)) + ((!g2) & (g734) & (!g732) & (g863) & (g895) & (!g977)) + ((!g2) & (g734) & (!g732) & (g863) & (g895) & (g977)) + ((!g2) & (g734) & (g732) & (!g863) & (!g895) & (g977)) + ((!g2) & (g734) & (g732) & (!g863) & (g895) & (!g977)) + ((!g2) & (g734) & (g732) & (!g863) & (g895) & (g977)) + ((!g2) & (g734) & (g732) & (g863) & (!g895) & (!g977)) + ((!g2) & (g734) & (g732) & (g863) & (!g895) & (g977)) + ((!g2) & (g734) & (g732) & (g863) & (g895) & (!g977)) + ((!g2) & (g734) & (g732) & (g863) & (g895) & (g977)) + ((g2) & (!g734) & (!g732) & (!g863) & (!g895) & (!g977)) + ((g2) & (!g734) & (!g732) & (!g863) & (g895) & (!g977)) + ((g2) & (!g734) & (!g732) & (g863) & (!g895) & (!g977)) + ((g2) & (!g734) & (!g732) & (g863) & (g895) & (!g977)) + ((g2) & (!g734) & (g732) & (!g863) & (!g895) & (!g977)) + ((g2) & (!g734) & (g732) & (g863) & (!g895) & (!g977)) + ((g2) & (g734) & (!g732) & (!g863) & (!g895) & (!g977)) + ((g2) & (g734) & (!g732) & (!g863) & (g895) & (!g977)) + ((g2) & (g734) & (g732) & (!g863) & (!g895) & (!g977)));
	assign g979 = (((!g838) & (!g839) & (!g852) & (!g854) & (g956) & (!g959)) + ((!g838) & (!g839) & (!g852) & (g854) & (g956) & (!g959)) + ((!g838) & (!g839) & (g852) & (!g854) & (!g956) & (!g959)) + ((!g838) & (!g839) & (g852) & (!g854) & (g956) & (!g959)) + ((!g838) & (!g839) & (g852) & (!g854) & (g956) & (g959)) + ((!g838) & (!g839) & (g852) & (g854) & (g956) & (!g959)) + ((!g838) & (g839) & (!g852) & (!g854) & (!g956) & (!g959)) + ((!g838) & (g839) & (!g852) & (!g854) & (g956) & (!g959)) + ((!g838) & (g839) & (!g852) & (!g854) & (g956) & (g959)) + ((!g838) & (g839) & (!g852) & (g854) & (g956) & (!g959)) + ((!g838) & (g839) & (g852) & (!g854) & (g956) & (!g959)) + ((!g838) & (g839) & (g852) & (g854) & (g956) & (!g959)) + ((g838) & (!g839) & (!g852) & (!g854) & (!g956) & (!g959)) + ((g838) & (!g839) & (!g852) & (!g854) & (g956) & (!g959)) + ((g838) & (!g839) & (!g852) & (!g854) & (g956) & (g959)) + ((g838) & (!g839) & (!g852) & (g854) & (g956) & (!g959)) + ((g838) & (!g839) & (g852) & (!g854) & (!g956) & (!g959)) + ((g838) & (!g839) & (g852) & (!g854) & (g956) & (!g959)) + ((g838) & (!g839) & (g852) & (!g854) & (g956) & (g959)) + ((g838) & (!g839) & (g852) & (g854) & (!g956) & (!g959)) + ((g838) & (!g839) & (g852) & (g854) & (g956) & (!g959)) + ((g838) & (!g839) & (g852) & (g854) & (g956) & (g959)) + ((g838) & (g839) & (!g852) & (!g854) & (!g956) & (!g959)) + ((g838) & (g839) & (!g852) & (!g854) & (g956) & (!g959)) + ((g838) & (g839) & (!g852) & (!g854) & (g956) & (g959)) + ((g838) & (g839) & (!g852) & (g854) & (!g956) & (!g959)) + ((g838) & (g839) & (!g852) & (g854) & (g956) & (!g959)) + ((g838) & (g839) & (!g852) & (g854) & (g956) & (g959)) + ((g838) & (g839) & (g852) & (!g854) & (!g956) & (!g959)) + ((g838) & (g839) & (g852) & (!g854) & (g956) & (!g959)) + ((g838) & (g839) & (g852) & (!g854) & (g956) & (g959)) + ((g838) & (g839) & (g852) & (g854) & (g956) & (!g959)));
	assign g980 = (((!g707) & (!g717) & (!sk[94]) & (!g718) & (g747) & (!g744)) + ((!g707) & (!g717) & (!sk[94]) & (!g718) & (g747) & (g744)) + ((!g707) & (!g717) & (!sk[94]) & (g718) & (!g747) & (!g744)) + ((!g707) & (!g717) & (!sk[94]) & (g718) & (!g747) & (g744)) + ((!g707) & (!g717) & (!sk[94]) & (g718) & (g747) & (!g744)) + ((!g707) & (!g717) & (!sk[94]) & (g718) & (g747) & (g744)) + ((!g707) & (!g717) & (sk[94]) & (g718) & (!g747) & (g744)) + ((!g707) & (!g717) & (sk[94]) & (g718) & (g747) & (g744)) + ((!g707) & (g717) & (!sk[94]) & (!g718) & (!g747) & (!g744)) + ((!g707) & (g717) & (!sk[94]) & (!g718) & (!g747) & (g744)) + ((!g707) & (g717) & (!sk[94]) & (!g718) & (g747) & (!g744)) + ((!g707) & (g717) & (!sk[94]) & (!g718) & (g747) & (g744)) + ((!g707) & (g717) & (!sk[94]) & (g718) & (!g747) & (!g744)) + ((!g707) & (g717) & (!sk[94]) & (g718) & (!g747) & (g744)) + ((!g707) & (g717) & (!sk[94]) & (g718) & (g747) & (!g744)) + ((!g707) & (g717) & (!sk[94]) & (g718) & (g747) & (g744)) + ((!g707) & (g717) & (sk[94]) & (!g718) & (g747) & (!g744)) + ((!g707) & (g717) & (sk[94]) & (!g718) & (g747) & (g744)) + ((!g707) & (g717) & (sk[94]) & (g718) & (!g747) & (g744)) + ((!g707) & (g717) & (sk[94]) & (g718) & (g747) & (!g744)) + ((!g707) & (g717) & (sk[94]) & (g718) & (g747) & (g744)) + ((g707) & (!g717) & (!sk[94]) & (!g718) & (g747) & (!g744)) + ((g707) & (!g717) & (!sk[94]) & (!g718) & (g747) & (g744)) + ((g707) & (!g717) & (!sk[94]) & (g718) & (!g747) & (!g744)) + ((g707) & (!g717) & (!sk[94]) & (g718) & (!g747) & (g744)) + ((g707) & (!g717) & (!sk[94]) & (g718) & (g747) & (!g744)) + ((g707) & (!g717) & (!sk[94]) & (g718) & (g747) & (g744)) + ((g707) & (!g717) & (sk[94]) & (!g718) & (g747) & (!g744)) + ((g707) & (!g717) & (sk[94]) & (!g718) & (g747) & (g744)) + ((g707) & (!g717) & (sk[94]) & (g718) & (!g747) & (g744)) + ((g707) & (!g717) & (sk[94]) & (g718) & (g747) & (!g744)) + ((g707) & (!g717) & (sk[94]) & (g718) & (g747) & (g744)) + ((g707) & (g717) & (!sk[94]) & (!g718) & (!g747) & (!g744)) + ((g707) & (g717) & (!sk[94]) & (!g718) & (!g747) & (g744)) + ((g707) & (g717) & (!sk[94]) & (!g718) & (g747) & (!g744)) + ((g707) & (g717) & (!sk[94]) & (!g718) & (g747) & (g744)) + ((g707) & (g717) & (!sk[94]) & (g718) & (!g747) & (!g744)) + ((g707) & (g717) & (!sk[94]) & (g718) & (!g747) & (g744)) + ((g707) & (g717) & (!sk[94]) & (g718) & (g747) & (!g744)) + ((g707) & (g717) & (!sk[94]) & (g718) & (g747) & (g744)) + ((g707) & (g717) & (sk[94]) & (g718) & (!g747) & (g744)) + ((g707) & (g717) & (sk[94]) & (g718) & (g747) & (g744)));
	assign g981 = (((!g200) & (!g681) & (!g731) & (!g742) & (!g748) & (!g980)) + ((!g200) & (!g681) & (!g731) & (g742) & (!g748) & (!g980)) + ((!g200) & (!g681) & (g731) & (!g742) & (!g748) & (!g980)) + ((!g200) & (g681) & (!g731) & (!g742) & (!g748) & (!g980)) + ((!g200) & (g681) & (!g731) & (!g742) & (g748) & (!g980)) + ((!g200) & (g681) & (!g731) & (g742) & (!g748) & (!g980)) + ((!g200) & (g681) & (!g731) & (g742) & (g748) & (!g980)) + ((!g200) & (g681) & (g731) & (!g742) & (!g748) & (!g980)) + ((!g200) & (g681) & (g731) & (!g742) & (g748) & (!g980)) + ((g200) & (!g681) & (!g731) & (!g742) & (!g748) & (g980)) + ((g200) & (!g681) & (!g731) & (!g742) & (g748) & (!g980)) + ((g200) & (!g681) & (!g731) & (!g742) & (g748) & (g980)) + ((g200) & (!g681) & (!g731) & (g742) & (!g748) & (g980)) + ((g200) & (!g681) & (!g731) & (g742) & (g748) & (!g980)) + ((g200) & (!g681) & (!g731) & (g742) & (g748) & (g980)) + ((g200) & (!g681) & (g731) & (!g742) & (!g748) & (g980)) + ((g200) & (!g681) & (g731) & (!g742) & (g748) & (!g980)) + ((g200) & (!g681) & (g731) & (!g742) & (g748) & (g980)) + ((g200) & (!g681) & (g731) & (g742) & (!g748) & (!g980)) + ((g200) & (!g681) & (g731) & (g742) & (!g748) & (g980)) + ((g200) & (!g681) & (g731) & (g742) & (g748) & (!g980)) + ((g200) & (!g681) & (g731) & (g742) & (g748) & (g980)) + ((g200) & (g681) & (!g731) & (!g742) & (!g748) & (g980)) + ((g200) & (g681) & (!g731) & (!g742) & (g748) & (g980)) + ((g200) & (g681) & (!g731) & (g742) & (!g748) & (g980)) + ((g200) & (g681) & (!g731) & (g742) & (g748) & (g980)) + ((g200) & (g681) & (g731) & (!g742) & (!g748) & (g980)) + ((g200) & (g681) & (g731) & (!g742) & (g748) & (g980)) + ((g200) & (g681) & (g731) & (g742) & (!g748) & (!g980)) + ((g200) & (g681) & (g731) & (g742) & (!g748) & (g980)) + ((g200) & (g681) & (g731) & (g742) & (g748) & (!g980)) + ((g200) & (g681) & (g731) & (g742) & (g748) & (g980)));
	assign g982 = (((!g949) & (g951) & (!sk[96]) & (!g955)) + ((!g949) & (g951) & (!sk[96]) & (g955)) + ((!g949) & (g951) & (sk[96]) & (!g955)) + ((g949) & (!g951) & (sk[96]) & (!g955)) + ((g949) & (g951) & (!sk[96]) & (!g955)) + ((g949) & (g951) & (!sk[96]) & (g955)) + ((g949) & (g951) & (sk[96]) & (!g955)) + ((g949) & (g951) & (sk[96]) & (g955)));
	assign g983 = (((!g585) & (!g597) & (!g679) & (g720) & (!g762) & (g765)) + ((!g585) & (!g597) & (!g679) & (g720) & (g762) & (g765)) + ((!g585) & (!g597) & (g679) & (!g720) & (g762) & (!g765)) + ((!g585) & (!g597) & (g679) & (!g720) & (g762) & (g765)) + ((!g585) & (!g597) & (g679) & (g720) & (!g762) & (g765)) + ((!g585) & (!g597) & (g679) & (g720) & (g762) & (!g765)) + ((!g585) & (!g597) & (g679) & (g720) & (g762) & (g765)) + ((!g585) & (g597) & (!g679) & (!g720) & (g762) & (!g765)) + ((!g585) & (g597) & (!g679) & (!g720) & (g762) & (g765)) + ((!g585) & (g597) & (!g679) & (g720) & (!g762) & (g765)) + ((!g585) & (g597) & (!g679) & (g720) & (g762) & (!g765)) + ((!g585) & (g597) & (!g679) & (g720) & (g762) & (g765)) + ((!g585) & (g597) & (g679) & (g720) & (!g762) & (g765)) + ((!g585) & (g597) & (g679) & (g720) & (g762) & (g765)) + ((g585) & (!g597) & (!g679) & (!g720) & (g762) & (!g765)) + ((g585) & (!g597) & (!g679) & (!g720) & (g762) & (g765)) + ((g585) & (!g597) & (!g679) & (g720) & (!g762) & (g765)) + ((g585) & (!g597) & (!g679) & (g720) & (g762) & (!g765)) + ((g585) & (!g597) & (!g679) & (g720) & (g762) & (g765)) + ((g585) & (!g597) & (g679) & (g720) & (!g762) & (g765)) + ((g585) & (!g597) & (g679) & (g720) & (g762) & (g765)) + ((g585) & (g597) & (!g679) & (g720) & (!g762) & (g765)) + ((g585) & (g597) & (!g679) & (g720) & (g762) & (g765)) + ((g585) & (g597) & (g679) & (!g720) & (g762) & (!g765)) + ((g585) & (g597) & (g679) & (!g720) & (g762) & (g765)) + ((g585) & (g597) & (g679) & (g720) & (!g762) & (g765)) + ((g585) & (g597) & (g679) & (g720) & (g762) & (!g765)) + ((g585) & (g597) & (g679) & (g720) & (g762) & (g765)));
	assign g984 = (((!g719) & (!g728) & (!g729) & (!g764) & (!g759) & (!g983)) + ((!g719) & (!g728) & (!g729) & (!g764) & (g759) & (!g983)) + ((!g719) & (!g728) & (g729) & (!g764) & (!g759) & (!g983)) + ((!g719) & (!g728) & (g729) & (g764) & (!g759) & (!g983)) + ((!g719) & (g728) & (!g729) & (!g764) & (!g759) & (!g983)) + ((!g719) & (g728) & (g729) & (!g764) & (!g759) & (!g983)) + ((!g719) & (g728) & (g729) & (!g764) & (g759) & (!g983)) + ((!g719) & (g728) & (g729) & (g764) & (!g759) & (!g983)) + ((!g719) & (g728) & (g729) & (g764) & (g759) & (!g983)) + ((g719) & (!g728) & (!g729) & (!g764) & (!g759) & (!g983)) + ((g719) & (!g728) & (g729) & (!g764) & (!g759) & (!g983)) + ((g719) & (!g728) & (g729) & (!g764) & (g759) & (!g983)) + ((g719) & (!g728) & (g729) & (g764) & (!g759) & (!g983)) + ((g719) & (!g728) & (g729) & (g764) & (g759) & (!g983)) + ((g719) & (g728) & (!g729) & (!g764) & (!g759) & (!g983)) + ((g719) & (g728) & (!g729) & (!g764) & (g759) & (!g983)) + ((g719) & (g728) & (g729) & (!g764) & (!g759) & (!g983)) + ((g719) & (g728) & (g729) & (g764) & (!g759) & (!g983)));
	assign g985 = (((!g252) & (!g725) & (!g952) & (g850) & (!g953) & (!g954)) + ((!g252) & (!g725) & (!g952) & (g850) & (!g953) & (g954)) + ((!g252) & (!g725) & (!g952) & (g850) & (g953) & (!g954)) + ((!g252) & (!g725) & (!g952) & (g850) & (g953) & (g954)) + ((!g252) & (g725) & (!g952) & (g850) & (!g953) & (!g954)) + ((!g252) & (g725) & (!g952) & (g850) & (g953) & (!g954)) + ((!g252) & (g725) & (!g952) & (g850) & (g953) & (g954)) + ((g252) & (!g725) & (!g952) & (!g850) & (!g953) & (g954)) + ((g252) & (!g725) & (!g952) & (g850) & (!g953) & (g954)) + ((g252) & (!g725) & (g952) & (!g850) & (!g953) & (g954)) + ((g252) & (!g725) & (g952) & (g850) & (!g953) & (!g954)) + ((g252) & (!g725) & (g952) & (g850) & (!g953) & (g954)) + ((g252) & (!g725) & (g952) & (g850) & (g953) & (!g954)) + ((g252) & (!g725) & (g952) & (g850) & (g953) & (g954)) + ((g252) & (g725) & (g952) & (g850) & (!g953) & (g954)));
	assign g986 = (((g252) & (!sk[100]) & (g726)) + ((g252) & (sk[100]) & (g726)));
	assign g987 = (((!g252) & (!sk[101]) & (!g985) & (!g986) & (g1447)) + ((!g252) & (!sk[101]) & (!g985) & (g986) & (g1447)) + ((!g252) & (!sk[101]) & (g985) & (!g986) & (g1447)) + ((!g252) & (!sk[101]) & (g985) & (g986) & (g1447)) + ((!g252) & (sk[101]) & (!g985) & (!g986) & (!g1447)) + ((!g252) & (sk[101]) & (!g985) & (g986) & (!g1447)) + ((!g252) & (sk[101]) & (g985) & (!g986) & (g1447)) + ((!g252) & (sk[101]) & (g985) & (g986) & (g1447)) + ((g252) & (!sk[101]) & (!g985) & (!g986) & (!g1447)) + ((g252) & (!sk[101]) & (!g985) & (!g986) & (g1447)) + ((g252) & (!sk[101]) & (!g985) & (g986) & (!g1447)) + ((g252) & (!sk[101]) & (!g985) & (g986) & (g1447)) + ((g252) & (!sk[101]) & (g985) & (!g986) & (!g1447)) + ((g252) & (!sk[101]) & (g985) & (!g986) & (g1447)) + ((g252) & (!sk[101]) & (g985) & (g986) & (!g1447)) + ((g252) & (!sk[101]) & (g985) & (g986) & (g1447)) + ((g252) & (sk[101]) & (!g985) & (!g986) & (g1447)) + ((g252) & (sk[101]) & (!g985) & (g986) & (!g1447)) + ((g252) & (sk[101]) & (g985) & (!g986) & (!g1447)) + ((g252) & (sk[101]) & (g985) & (g986) & (g1447)));
	assign g988 = (((!sk[102]) & (!g202) & (g984) & (!g987)) + ((!sk[102]) & (!g202) & (g984) & (g987)) + ((!sk[102]) & (g202) & (g984) & (!g987)) + ((!sk[102]) & (g202) & (g984) & (g987)) + ((sk[102]) & (!g202) & (!g984) & (!g987)) + ((sk[102]) & (!g202) & (g984) & (g987)) + ((sk[102]) & (g202) & (!g984) & (g987)) + ((sk[102]) & (g202) & (g984) & (!g987)));
	assign g989 = (((!g979) & (!sk[103]) & (!g981) & (!g982) & (g988)) + ((!g979) & (!sk[103]) & (!g981) & (g982) & (g988)) + ((!g979) & (!sk[103]) & (g981) & (!g982) & (g988)) + ((!g979) & (!sk[103]) & (g981) & (g982) & (g988)) + ((!g979) & (sk[103]) & (!g981) & (!g982) & (g988)) + ((!g979) & (sk[103]) & (!g981) & (g982) & (!g988)) + ((!g979) & (sk[103]) & (g981) & (!g982) & (!g988)) + ((!g979) & (sk[103]) & (g981) & (g982) & (g988)) + ((g979) & (!sk[103]) & (!g981) & (!g982) & (!g988)) + ((g979) & (!sk[103]) & (!g981) & (!g982) & (g988)) + ((g979) & (!sk[103]) & (!g981) & (g982) & (!g988)) + ((g979) & (!sk[103]) & (!g981) & (g982) & (g988)) + ((g979) & (!sk[103]) & (g981) & (!g982) & (!g988)) + ((g979) & (!sk[103]) & (g981) & (!g982) & (g988)) + ((g979) & (!sk[103]) & (g981) & (g982) & (!g988)) + ((g979) & (!sk[103]) & (g981) & (g982) & (g988)) + ((g979) & (sk[103]) & (!g981) & (!g982) & (!g988)) + ((g979) & (sk[103]) & (!g981) & (g982) & (g988)) + ((g979) & (sk[103]) & (g981) & (!g982) & (g988)) + ((g979) & (sk[103]) & (g981) & (g982) & (!g988)));
	assign g990 = (((!g946) & (!g976) & (!g948) & (!g960) & (!g978) & (g989)) + ((!g946) & (!g976) & (!g948) & (!g960) & (g978) & (!g989)) + ((!g946) & (!g976) & (!g948) & (g960) & (!g978) & (g989)) + ((!g946) & (!g976) & (!g948) & (g960) & (g978) & (!g989)) + ((!g946) & (!g976) & (g948) & (!g960) & (!g978) & (g989)) + ((!g946) & (!g976) & (g948) & (!g960) & (g978) & (!g989)) + ((!g946) & (!g976) & (g948) & (g960) & (!g978) & (g989)) + ((!g946) & (!g976) & (g948) & (g960) & (g978) & (!g989)) + ((!g946) & (g976) & (!g948) & (!g960) & (!g978) & (!g989)) + ((!g946) & (g976) & (!g948) & (!g960) & (g978) & (g989)) + ((!g946) & (g976) & (!g948) & (g960) & (!g978) & (g989)) + ((!g946) & (g976) & (!g948) & (g960) & (g978) & (!g989)) + ((!g946) & (g976) & (g948) & (!g960) & (!g978) & (g989)) + ((!g946) & (g976) & (g948) & (!g960) & (g978) & (!g989)) + ((!g946) & (g976) & (g948) & (g960) & (!g978) & (!g989)) + ((!g946) & (g976) & (g948) & (g960) & (g978) & (g989)) + ((g946) & (!g976) & (!g948) & (!g960) & (!g978) & (!g989)) + ((g946) & (!g976) & (!g948) & (!g960) & (g978) & (g989)) + ((g946) & (!g976) & (!g948) & (g960) & (!g978) & (g989)) + ((g946) & (!g976) & (!g948) & (g960) & (g978) & (!g989)) + ((g946) & (!g976) & (g948) & (!g960) & (!g978) & (g989)) + ((g946) & (!g976) & (g948) & (!g960) & (g978) & (!g989)) + ((g946) & (!g976) & (g948) & (g960) & (!g978) & (!g989)) + ((g946) & (!g976) & (g948) & (g960) & (g978) & (g989)) + ((g946) & (g976) & (!g948) & (!g960) & (!g978) & (!g989)) + ((g946) & (g976) & (!g948) & (!g960) & (g978) & (g989)) + ((g946) & (g976) & (!g948) & (g960) & (!g978) & (!g989)) + ((g946) & (g976) & (!g948) & (g960) & (g978) & (g989)) + ((g946) & (g976) & (g948) & (!g960) & (!g978) & (!g989)) + ((g946) & (g976) & (g948) & (!g960) & (g978) & (g989)) + ((g946) & (g976) & (g948) & (g960) & (!g978) & (!g989)) + ((g946) & (g976) & (g948) & (g960) & (g978) & (g989)));
	assign g991 = (((!g48) & (!sk[105]) & (!g52) & (!g56) & (g61)) + ((!g48) & (!sk[105]) & (!g52) & (g56) & (g61)) + ((!g48) & (!sk[105]) & (g52) & (!g56) & (g61)) + ((!g48) & (!sk[105]) & (g52) & (g56) & (g61)) + ((g48) & (!sk[105]) & (!g52) & (!g56) & (!g61)) + ((g48) & (!sk[105]) & (!g52) & (!g56) & (g61)) + ((g48) & (!sk[105]) & (!g52) & (g56) & (!g61)) + ((g48) & (!sk[105]) & (!g52) & (g56) & (g61)) + ((g48) & (!sk[105]) & (g52) & (!g56) & (!g61)) + ((g48) & (!sk[105]) & (g52) & (!g56) & (g61)) + ((g48) & (!sk[105]) & (g52) & (g56) & (!g61)) + ((g48) & (!sk[105]) & (g52) & (g56) & (g61)) + ((g48) & (sk[105]) & (g52) & (g56) & (g61)));
	assign g992 = (((!g28) & (!sk[106]) & (g29) & (!g628)) + ((!g28) & (!sk[106]) & (g29) & (g628)) + ((!g28) & (sk[106]) & (!g29) & (g628)) + ((g28) & (!sk[106]) & (g29) & (!g628)) + ((g28) & (!sk[106]) & (g29) & (g628)));
	assign g993 = (((g15) & (g22) & (g991) & (!g217) & (g966) & (g992)));
	assign g994 = (((!g889) & (!g871) & (!g883) & (!sk[108]) & (g970) & (!g993)) + ((!g889) & (!g871) & (!g883) & (!sk[108]) & (g970) & (g993)) + ((!g889) & (!g871) & (!g883) & (sk[108]) & (!g970) & (!g993)) + ((!g889) & (!g871) & (!g883) & (sk[108]) & (g970) & (!g993)) + ((!g889) & (!g871) & (g883) & (!sk[108]) & (!g970) & (!g993)) + ((!g889) & (!g871) & (g883) & (!sk[108]) & (!g970) & (g993)) + ((!g889) & (!g871) & (g883) & (!sk[108]) & (g970) & (!g993)) + ((!g889) & (!g871) & (g883) & (!sk[108]) & (g970) & (g993)) + ((!g889) & (!g871) & (g883) & (sk[108]) & (!g970) & (!g993)) + ((!g889) & (!g871) & (g883) & (sk[108]) & (g970) & (!g993)) + ((!g889) & (g871) & (!g883) & (!sk[108]) & (!g970) & (!g993)) + ((!g889) & (g871) & (!g883) & (!sk[108]) & (!g970) & (g993)) + ((!g889) & (g871) & (!g883) & (!sk[108]) & (g970) & (!g993)) + ((!g889) & (g871) & (!g883) & (!sk[108]) & (g970) & (g993)) + ((!g889) & (g871) & (!g883) & (sk[108]) & (!g970) & (!g993)) + ((!g889) & (g871) & (!g883) & (sk[108]) & (g970) & (!g993)) + ((!g889) & (g871) & (g883) & (!sk[108]) & (!g970) & (!g993)) + ((!g889) & (g871) & (g883) & (!sk[108]) & (!g970) & (g993)) + ((!g889) & (g871) & (g883) & (!sk[108]) & (g970) & (!g993)) + ((!g889) & (g871) & (g883) & (!sk[108]) & (g970) & (g993)) + ((!g889) & (g871) & (g883) & (sk[108]) & (!g970) & (!g993)) + ((!g889) & (g871) & (g883) & (sk[108]) & (g970) & (!g993)) + ((g889) & (!g871) & (!g883) & (!sk[108]) & (g970) & (!g993)) + ((g889) & (!g871) & (!g883) & (!sk[108]) & (g970) & (g993)) + ((g889) & (!g871) & (!g883) & (sk[108]) & (!g970) & (!g993)) + ((g889) & (!g871) & (!g883) & (sk[108]) & (g970) & (!g993)) + ((g889) & (!g871) & (g883) & (!sk[108]) & (!g970) & (!g993)) + ((g889) & (!g871) & (g883) & (!sk[108]) & (!g970) & (g993)) + ((g889) & (!g871) & (g883) & (!sk[108]) & (g970) & (!g993)) + ((g889) & (!g871) & (g883) & (!sk[108]) & (g970) & (g993)) + ((g889) & (!g871) & (g883) & (sk[108]) & (!g970) & (!g993)) + ((g889) & (!g871) & (g883) & (sk[108]) & (g970) & (!g993)) + ((g889) & (g871) & (!g883) & (!sk[108]) & (!g970) & (!g993)) + ((g889) & (g871) & (!g883) & (!sk[108]) & (!g970) & (g993)) + ((g889) & (g871) & (!g883) & (!sk[108]) & (g970) & (!g993)) + ((g889) & (g871) & (!g883) & (!sk[108]) & (g970) & (g993)) + ((g889) & (g871) & (!g883) & (sk[108]) & (!g970) & (!g993)) + ((g889) & (g871) & (!g883) & (sk[108]) & (g970) & (!g993)) + ((g889) & (g871) & (g883) & (!sk[108]) & (!g970) & (!g993)) + ((g889) & (g871) & (g883) & (!sk[108]) & (!g970) & (g993)) + ((g889) & (g871) & (g883) & (!sk[108]) & (g970) & (!g993)) + ((g889) & (g871) & (g883) & (!sk[108]) & (g970) & (g993)) + ((g889) & (g871) & (g883) & (sk[108]) & (!g970) & (!g993)) + ((g889) & (g871) & (g883) & (sk[108]) & (g970) & (g993)));
	assign g995 = (((!g962) & (!sk[109]) & (!g963) & (!g884) & (g971) & (!g994)) + ((!g962) & (!sk[109]) & (!g963) & (!g884) & (g971) & (g994)) + ((!g962) & (!sk[109]) & (!g963) & (g884) & (!g971) & (!g994)) + ((!g962) & (!sk[109]) & (!g963) & (g884) & (!g971) & (g994)) + ((!g962) & (!sk[109]) & (!g963) & (g884) & (g971) & (!g994)) + ((!g962) & (!sk[109]) & (!g963) & (g884) & (g971) & (g994)) + ((!g962) & (!sk[109]) & (g963) & (!g884) & (!g971) & (!g994)) + ((!g962) & (!sk[109]) & (g963) & (!g884) & (!g971) & (g994)) + ((!g962) & (!sk[109]) & (g963) & (!g884) & (g971) & (!g994)) + ((!g962) & (!sk[109]) & (g963) & (!g884) & (g971) & (g994)) + ((!g962) & (!sk[109]) & (g963) & (g884) & (!g971) & (!g994)) + ((!g962) & (!sk[109]) & (g963) & (g884) & (!g971) & (g994)) + ((!g962) & (!sk[109]) & (g963) & (g884) & (g971) & (!g994)) + ((!g962) & (!sk[109]) & (g963) & (g884) & (g971) & (g994)) + ((!g962) & (sk[109]) & (!g963) & (!g884) & (!g971) & (g994)) + ((!g962) & (sk[109]) & (!g963) & (!g884) & (g971) & (g994)) + ((!g962) & (sk[109]) & (!g963) & (g884) & (!g971) & (!g994)) + ((!g962) & (sk[109]) & (!g963) & (g884) & (g971) & (g994)) + ((!g962) & (sk[109]) & (g963) & (!g884) & (!g971) & (!g994)) + ((!g962) & (sk[109]) & (g963) & (!g884) & (g971) & (g994)) + ((!g962) & (sk[109]) & (g963) & (g884) & (!g971) & (!g994)) + ((!g962) & (sk[109]) & (g963) & (g884) & (g971) & (g994)) + ((g962) & (!sk[109]) & (!g963) & (!g884) & (g971) & (!g994)) + ((g962) & (!sk[109]) & (!g963) & (!g884) & (g971) & (g994)) + ((g962) & (!sk[109]) & (!g963) & (g884) & (!g971) & (!g994)) + ((g962) & (!sk[109]) & (!g963) & (g884) & (!g971) & (g994)) + ((g962) & (!sk[109]) & (!g963) & (g884) & (g971) & (!g994)) + ((g962) & (!sk[109]) & (!g963) & (g884) & (g971) & (g994)) + ((g962) & (!sk[109]) & (g963) & (!g884) & (!g971) & (!g994)) + ((g962) & (!sk[109]) & (g963) & (!g884) & (!g971) & (g994)) + ((g962) & (!sk[109]) & (g963) & (!g884) & (g971) & (!g994)) + ((g962) & (!sk[109]) & (g963) & (!g884) & (g971) & (g994)) + ((g962) & (!sk[109]) & (g963) & (g884) & (!g971) & (!g994)) + ((g962) & (!sk[109]) & (g963) & (g884) & (!g971) & (g994)) + ((g962) & (!sk[109]) & (g963) & (g884) & (g971) & (!g994)) + ((g962) & (!sk[109]) & (g963) & (g884) & (g971) & (g994)) + ((g962) & (sk[109]) & (!g963) & (!g884) & (!g971) & (g994)) + ((g962) & (sk[109]) & (!g963) & (!g884) & (g971) & (!g994)) + ((g962) & (sk[109]) & (!g963) & (g884) & (!g971) & (g994)) + ((g962) & (sk[109]) & (!g963) & (g884) & (g971) & (!g994)) + ((g962) & (sk[109]) & (g963) & (!g884) & (!g971) & (g994)) + ((g962) & (sk[109]) & (g963) & (!g884) & (g971) & (!g994)) + ((g962) & (sk[109]) & (g963) & (g884) & (!g971) & (g994)) + ((g962) & (sk[109]) & (g963) & (g884) & (g971) & (g994)));
	assign g996 = (((!g891) & (!g962) & (!g864) & (!g892) & (!g971) & (!g994)) + ((!g891) & (!g962) & (!g864) & (!g892) & (!g971) & (g994)) + ((!g891) & (!g962) & (!g864) & (!g892) & (g971) & (!g994)) + ((!g891) & (!g962) & (!g864) & (!g892) & (g971) & (g994)) + ((!g891) & (!g962) & (!g864) & (g892) & (!g971) & (!g994)) + ((!g891) & (!g962) & (!g864) & (g892) & (!g971) & (g994)) + ((!g891) & (g962) & (!g864) & (!g892) & (!g971) & (!g994)) + ((!g891) & (g962) & (!g864) & (!g892) & (!g971) & (g994)) + ((!g891) & (g962) & (!g864) & (!g892) & (g971) & (!g994)) + ((!g891) & (g962) & (!g864) & (!g892) & (g971) & (g994)) + ((!g891) & (g962) & (!g864) & (g892) & (!g971) & (!g994)) + ((!g891) & (g962) & (!g864) & (g892) & (!g971) & (g994)) + ((!g891) & (g962) & (g864) & (!g892) & (!g971) & (!g994)) + ((!g891) & (g962) & (g864) & (!g892) & (!g971) & (g994)) + ((!g891) & (g962) & (g864) & (!g892) & (g971) & (!g994)) + ((!g891) & (g962) & (g864) & (!g892) & (g971) & (g994)) + ((!g891) & (g962) & (g864) & (g892) & (!g971) & (!g994)) + ((!g891) & (g962) & (g864) & (g892) & (!g971) & (g994)) + ((g891) & (!g962) & (!g864) & (!g892) & (!g971) & (!g994)) + ((g891) & (!g962) & (!g864) & (!g892) & (g971) & (!g994)) + ((g891) & (!g962) & (!g864) & (g892) & (!g971) & (!g994)) + ((g891) & (g962) & (!g864) & (!g892) & (!g971) & (!g994)) + ((g891) & (g962) & (!g864) & (!g892) & (g971) & (!g994)) + ((g891) & (g962) & (!g864) & (g892) & (!g971) & (!g994)) + ((g891) & (g962) & (g864) & (!g892) & (!g971) & (!g994)) + ((g891) & (g962) & (g864) & (!g892) & (g971) & (!g994)) + ((g891) & (g962) & (g864) & (g892) & (!g971) & (!g994)));
	assign g997 = (((!g683) & (!sk[111]) & (!g868) & (!g995) & (g996)) + ((!g683) & (!sk[111]) & (!g868) & (g995) & (g996)) + ((!g683) & (!sk[111]) & (g868) & (!g995) & (g996)) + ((!g683) & (!sk[111]) & (g868) & (g995) & (g996)) + ((!g683) & (sk[111]) & (!g868) & (!g995) & (g996)) + ((!g683) & (sk[111]) & (!g868) & (g995) & (g996)) + ((!g683) & (sk[111]) & (g868) & (!g995) & (g996)) + ((g683) & (!sk[111]) & (!g868) & (!g995) & (!g996)) + ((g683) & (!sk[111]) & (!g868) & (!g995) & (g996)) + ((g683) & (!sk[111]) & (!g868) & (g995) & (!g996)) + ((g683) & (!sk[111]) & (!g868) & (g995) & (g996)) + ((g683) & (!sk[111]) & (g868) & (!g995) & (!g996)) + ((g683) & (!sk[111]) & (g868) & (!g995) & (g996)) + ((g683) & (!sk[111]) & (g868) & (g995) & (!g996)) + ((g683) & (!sk[111]) & (g868) & (g995) & (g996)) + ((g683) & (sk[111]) & (!g868) & (!g995) & (!g996)) + ((g683) & (sk[111]) & (!g868) & (g995) & (!g996)) + ((g683) & (sk[111]) & (g868) & (!g995) & (!g996)) + ((g683) & (sk[111]) & (g868) & (g995) & (!g996)) + ((g683) & (sk[111]) & (g868) & (g995) & (g996)));
	assign g998 = (((!sk[112]) & (g990) & (g997)) + ((sk[112]) & (!g990) & (g997)) + ((sk[112]) & (g990) & (!g997)));
	assign g999 = (((!g9) & (!g70) & (!g12) & (!g41) & (sk[113]) & (!g35)) + ((!g9) & (!g70) & (!g12) & (g41) & (!sk[113]) & (!g35)) + ((!g9) & (!g70) & (!g12) & (g41) & (!sk[113]) & (g35)) + ((!g9) & (!g70) & (!g12) & (g41) & (sk[113]) & (!g35)) + ((!g9) & (!g70) & (g12) & (!g41) & (!sk[113]) & (!g35)) + ((!g9) & (!g70) & (g12) & (!g41) & (!sk[113]) & (g35)) + ((!g9) & (!g70) & (g12) & (!g41) & (sk[113]) & (!g35)) + ((!g9) & (!g70) & (g12) & (g41) & (!sk[113]) & (!g35)) + ((!g9) & (!g70) & (g12) & (g41) & (!sk[113]) & (g35)) + ((!g9) & (!g70) & (g12) & (g41) & (sk[113]) & (!g35)) + ((!g9) & (g70) & (!g12) & (!g41) & (!sk[113]) & (!g35)) + ((!g9) & (g70) & (!g12) & (!g41) & (!sk[113]) & (g35)) + ((!g9) & (g70) & (!g12) & (!g41) & (sk[113]) & (!g35)) + ((!g9) & (g70) & (!g12) & (g41) & (!sk[113]) & (!g35)) + ((!g9) & (g70) & (!g12) & (g41) & (!sk[113]) & (g35)) + ((!g9) & (g70) & (!g12) & (g41) & (sk[113]) & (!g35)) + ((!g9) & (g70) & (g12) & (!g41) & (!sk[113]) & (!g35)) + ((!g9) & (g70) & (g12) & (!g41) & (!sk[113]) & (g35)) + ((!g9) & (g70) & (g12) & (g41) & (!sk[113]) & (!g35)) + ((!g9) & (g70) & (g12) & (g41) & (!sk[113]) & (g35)) + ((g9) & (!g70) & (!g12) & (!g41) & (sk[113]) & (!g35)) + ((g9) & (!g70) & (!g12) & (g41) & (!sk[113]) & (!g35)) + ((g9) & (!g70) & (!g12) & (g41) & (!sk[113]) & (g35)) + ((g9) & (!g70) & (g12) & (!g41) & (!sk[113]) & (!g35)) + ((g9) & (!g70) & (g12) & (!g41) & (!sk[113]) & (g35)) + ((g9) & (!g70) & (g12) & (!g41) & (sk[113]) & (!g35)) + ((g9) & (!g70) & (g12) & (g41) & (!sk[113]) & (!g35)) + ((g9) & (!g70) & (g12) & (g41) & (!sk[113]) & (g35)) + ((g9) & (g70) & (!g12) & (!g41) & (!sk[113]) & (!g35)) + ((g9) & (g70) & (!g12) & (!g41) & (!sk[113]) & (g35)) + ((g9) & (g70) & (!g12) & (!g41) & (sk[113]) & (!g35)) + ((g9) & (g70) & (!g12) & (g41) & (!sk[113]) & (!g35)) + ((g9) & (g70) & (!g12) & (g41) & (!sk[113]) & (g35)) + ((g9) & (g70) & (g12) & (!g41) & (!sk[113]) & (!g35)) + ((g9) & (g70) & (g12) & (!g41) & (!sk[113]) & (g35)) + ((g9) & (g70) & (g12) & (g41) & (!sk[113]) & (!g35)) + ((g9) & (g70) & (g12) & (g41) & (!sk[113]) & (g35)));
	assign g1000 = (((!g112) & (!sk[114]) & (!g113) & (!g97) & (g70)) + ((!g112) & (!sk[114]) & (!g113) & (g97) & (g70)) + ((!g112) & (!sk[114]) & (g113) & (!g97) & (g70)) + ((!g112) & (!sk[114]) & (g113) & (g97) & (g70)) + ((!g112) & (sk[114]) & (!g113) & (g97) & (g70)) + ((g112) & (!sk[114]) & (!g113) & (!g97) & (!g70)) + ((g112) & (!sk[114]) & (!g113) & (!g97) & (g70)) + ((g112) & (!sk[114]) & (!g113) & (g97) & (!g70)) + ((g112) & (!sk[114]) & (!g113) & (g97) & (g70)) + ((g112) & (!sk[114]) & (g113) & (!g97) & (!g70)) + ((g112) & (!sk[114]) & (g113) & (!g97) & (g70)) + ((g112) & (!sk[114]) & (g113) & (g97) & (!g70)) + ((g112) & (!sk[114]) & (g113) & (g97) & (g70)));
	assign g1001 = (((!sk[115]) & (!g11) & (g124) & (!g1000)) + ((!sk[115]) & (!g11) & (g124) & (g1000)) + ((!sk[115]) & (g11) & (g124) & (!g1000)) + ((!sk[115]) & (g11) & (g124) & (g1000)) + ((sk[115]) & (!g11) & (!g124) & (!g1000)));
	assign g1002 = (((!g70) & (!sk[116]) & (!g49) & (!g62) & (g18)) + ((!g70) & (!sk[116]) & (!g49) & (g62) & (g18)) + ((!g70) & (!sk[116]) & (g49) & (!g62) & (g18)) + ((!g70) & (!sk[116]) & (g49) & (g62) & (g18)) + ((!g70) & (sk[116]) & (g49) & (g62) & (!g18)) + ((!g70) & (sk[116]) & (g49) & (g62) & (g18)) + ((g70) & (!sk[116]) & (!g49) & (!g62) & (!g18)) + ((g70) & (!sk[116]) & (!g49) & (!g62) & (g18)) + ((g70) & (!sk[116]) & (!g49) & (g62) & (!g18)) + ((g70) & (!sk[116]) & (!g49) & (g62) & (g18)) + ((g70) & (!sk[116]) & (g49) & (!g62) & (!g18)) + ((g70) & (!sk[116]) & (g49) & (!g62) & (g18)) + ((g70) & (!sk[116]) & (g49) & (g62) & (!g18)) + ((g70) & (!sk[116]) & (g49) & (g62) & (g18)) + ((g70) & (sk[116]) & (!g49) & (!g62) & (g18)) + ((g70) & (sk[116]) & (!g49) & (g62) & (g18)) + ((g70) & (sk[116]) & (g49) & (!g62) & (g18)) + ((g70) & (sk[116]) & (g49) & (g62) & (!g18)) + ((g70) & (sk[116]) & (g49) & (g62) & (g18)));
	assign g1003 = (((!g97) & (!g98) & (!g16) & (!g100) & (sk[117]) & (!g1002)) + ((!g97) & (!g98) & (!g16) & (g100) & (!sk[117]) & (!g1002)) + ((!g97) & (!g98) & (!g16) & (g100) & (!sk[117]) & (g1002)) + ((!g97) & (!g98) & (!g16) & (g100) & (sk[117]) & (!g1002)) + ((!g97) & (!g98) & (g16) & (!g100) & (!sk[117]) & (!g1002)) + ((!g97) & (!g98) & (g16) & (!g100) & (!sk[117]) & (g1002)) + ((!g97) & (!g98) & (g16) & (!g100) & (sk[117]) & (!g1002)) + ((!g97) & (!g98) & (g16) & (g100) & (!sk[117]) & (!g1002)) + ((!g97) & (!g98) & (g16) & (g100) & (!sk[117]) & (g1002)) + ((!g97) & (g98) & (!g16) & (!g100) & (!sk[117]) & (!g1002)) + ((!g97) & (g98) & (!g16) & (!g100) & (!sk[117]) & (g1002)) + ((!g97) & (g98) & (!g16) & (!g100) & (sk[117]) & (!g1002)) + ((!g97) & (g98) & (!g16) & (g100) & (!sk[117]) & (!g1002)) + ((!g97) & (g98) & (!g16) & (g100) & (!sk[117]) & (g1002)) + ((!g97) & (g98) & (!g16) & (g100) & (sk[117]) & (!g1002)) + ((!g97) & (g98) & (g16) & (!g100) & (!sk[117]) & (!g1002)) + ((!g97) & (g98) & (g16) & (!g100) & (!sk[117]) & (g1002)) + ((!g97) & (g98) & (g16) & (!g100) & (sk[117]) & (!g1002)) + ((!g97) & (g98) & (g16) & (g100) & (!sk[117]) & (!g1002)) + ((!g97) & (g98) & (g16) & (g100) & (!sk[117]) & (g1002)) + ((!g97) & (g98) & (g16) & (g100) & (sk[117]) & (!g1002)) + ((g97) & (!g98) & (!g16) & (!g100) & (sk[117]) & (!g1002)) + ((g97) & (!g98) & (!g16) & (g100) & (!sk[117]) & (!g1002)) + ((g97) & (!g98) & (!g16) & (g100) & (!sk[117]) & (g1002)) + ((g97) & (!g98) & (!g16) & (g100) & (sk[117]) & (!g1002)) + ((g97) & (!g98) & (g16) & (!g100) & (!sk[117]) & (!g1002)) + ((g97) & (!g98) & (g16) & (!g100) & (!sk[117]) & (g1002)) + ((g97) & (!g98) & (g16) & (!g100) & (sk[117]) & (!g1002)) + ((g97) & (!g98) & (g16) & (g100) & (!sk[117]) & (!g1002)) + ((g97) & (!g98) & (g16) & (g100) & (!sk[117]) & (g1002)) + ((g97) & (!g98) & (g16) & (g100) & (sk[117]) & (!g1002)) + ((g97) & (g98) & (!g16) & (!g100) & (!sk[117]) & (!g1002)) + ((g97) & (g98) & (!g16) & (!g100) & (!sk[117]) & (g1002)) + ((g97) & (g98) & (!g16) & (!g100) & (sk[117]) & (!g1002)) + ((g97) & (g98) & (!g16) & (g100) & (!sk[117]) & (!g1002)) + ((g97) & (g98) & (!g16) & (g100) & (!sk[117]) & (g1002)) + ((g97) & (g98) & (!g16) & (g100) & (sk[117]) & (!g1002)) + ((g97) & (g98) & (g16) & (!g100) & (!sk[117]) & (!g1002)) + ((g97) & (g98) & (g16) & (!g100) & (!sk[117]) & (g1002)) + ((g97) & (g98) & (g16) & (!g100) & (sk[117]) & (!g1002)) + ((g97) & (g98) & (g16) & (g100) & (!sk[117]) & (!g1002)) + ((g97) & (g98) & (g16) & (g100) & (!sk[117]) & (g1002)));
	assign g1004 = (((g550) & (g590) & (g621) & (g999) & (g1001) & (g1003)));
	assign g1005 = (((!g16) & (!g40) & (!g85) & (!sk[119]) & (g1004)) + ((!g16) & (!g40) & (!g85) & (sk[119]) & (g1004)) + ((!g16) & (!g40) & (g85) & (!sk[119]) & (g1004)) + ((!g16) & (g40) & (!g85) & (!sk[119]) & (g1004)) + ((!g16) & (g40) & (!g85) & (sk[119]) & (g1004)) + ((!g16) & (g40) & (g85) & (!sk[119]) & (g1004)) + ((g16) & (!g40) & (!g85) & (!sk[119]) & (!g1004)) + ((g16) & (!g40) & (!g85) & (!sk[119]) & (g1004)) + ((g16) & (!g40) & (!g85) & (sk[119]) & (g1004)) + ((g16) & (!g40) & (g85) & (!sk[119]) & (!g1004)) + ((g16) & (!g40) & (g85) & (!sk[119]) & (g1004)) + ((g16) & (g40) & (!g85) & (!sk[119]) & (!g1004)) + ((g16) & (g40) & (!g85) & (!sk[119]) & (g1004)) + ((g16) & (g40) & (g85) & (!sk[119]) & (!g1004)) + ((g16) & (g40) & (g85) & (!sk[119]) & (g1004)));
	assign g1006 = (((!g26) & (sk[120]) & (!g28)) + ((g26) & (!sk[120]) & (g28)));
	assign g1007 = (((!g127) & (!g184) & (g230) & (g1006) & (g239) & (g873)));
	assign g1008 = (((!g38) & (!g114) & (g115) & (!g8) & (!g40) & (g20)) + ((!g38) & (!g114) & (g115) & (!g8) & (g40) & (g20)) + ((!g38) & (g114) & (!g115) & (!g8) & (!g40) & (g20)) + ((!g38) & (g114) & (!g115) & (!g8) & (g40) & (!g20)) + ((!g38) & (g114) & (!g115) & (!g8) & (g40) & (g20)) + ((g38) & (!g114) & (g115) & (!g8) & (!g40) & (g20)) + ((g38) & (!g114) & (g115) & (!g8) & (g40) & (g20)) + ((g38) & (g114) & (!g115) & (!g8) & (!g40) & (g20)) + ((g38) & (g114) & (!g115) & (!g8) & (g40) & (!g20)) + ((g38) & (g114) & (!g115) & (!g8) & (g40) & (g20)) + ((g38) & (g114) & (g115) & (!g8) & (!g40) & (!g20)) + ((g38) & (g114) & (g115) & (!g8) & (!g40) & (g20)) + ((g38) & (g114) & (g115) & (!g8) & (g40) & (!g20)) + ((g38) & (g114) & (g115) & (!g8) & (g40) & (g20)));
	assign g1009 = (((!g99) & (!g25) & (g879) & (!g33) & (g660) & (!g1008)) + ((!g99) & (g25) & (g879) & (!g33) & (g660) & (!g1008)) + ((g99) & (!g25) & (g879) & (!g33) & (g660) & (!g1008)));
	assign g1010 = (((!g228) & (!g418) & (!sk[124]) & (!g1005) & (g1007) & (!g1009)) + ((!g228) & (!g418) & (!sk[124]) & (!g1005) & (g1007) & (g1009)) + ((!g228) & (!g418) & (!sk[124]) & (g1005) & (!g1007) & (!g1009)) + ((!g228) & (!g418) & (!sk[124]) & (g1005) & (!g1007) & (g1009)) + ((!g228) & (!g418) & (!sk[124]) & (g1005) & (g1007) & (!g1009)) + ((!g228) & (!g418) & (!sk[124]) & (g1005) & (g1007) & (g1009)) + ((!g228) & (g418) & (!sk[124]) & (!g1005) & (!g1007) & (!g1009)) + ((!g228) & (g418) & (!sk[124]) & (!g1005) & (!g1007) & (g1009)) + ((!g228) & (g418) & (!sk[124]) & (!g1005) & (g1007) & (!g1009)) + ((!g228) & (g418) & (!sk[124]) & (!g1005) & (g1007) & (g1009)) + ((!g228) & (g418) & (!sk[124]) & (g1005) & (!g1007) & (!g1009)) + ((!g228) & (g418) & (!sk[124]) & (g1005) & (!g1007) & (g1009)) + ((!g228) & (g418) & (!sk[124]) & (g1005) & (g1007) & (!g1009)) + ((!g228) & (g418) & (!sk[124]) & (g1005) & (g1007) & (g1009)) + ((g228) & (!g418) & (!sk[124]) & (!g1005) & (g1007) & (!g1009)) + ((g228) & (!g418) & (!sk[124]) & (!g1005) & (g1007) & (g1009)) + ((g228) & (!g418) & (!sk[124]) & (g1005) & (!g1007) & (!g1009)) + ((g228) & (!g418) & (!sk[124]) & (g1005) & (!g1007) & (g1009)) + ((g228) & (!g418) & (!sk[124]) & (g1005) & (g1007) & (!g1009)) + ((g228) & (!g418) & (!sk[124]) & (g1005) & (g1007) & (g1009)) + ((g228) & (g418) & (!sk[124]) & (!g1005) & (!g1007) & (!g1009)) + ((g228) & (g418) & (!sk[124]) & (!g1005) & (!g1007) & (g1009)) + ((g228) & (g418) & (!sk[124]) & (!g1005) & (g1007) & (!g1009)) + ((g228) & (g418) & (!sk[124]) & (!g1005) & (g1007) & (g1009)) + ((g228) & (g418) & (!sk[124]) & (g1005) & (!g1007) & (!g1009)) + ((g228) & (g418) & (!sk[124]) & (g1005) & (!g1007) & (g1009)) + ((g228) & (g418) & (!sk[124]) & (g1005) & (g1007) & (!g1009)) + ((g228) & (g418) & (!sk[124]) & (g1005) & (g1007) & (g1009)) + ((g228) & (g418) & (sk[124]) & (g1005) & (g1007) & (g1009)));
	assign g1011 = (((!g683) & (!g868) & (!g946) & (!g961) & (!g972) & (g973)) + ((!g683) & (!g868) & (!g946) & (!g961) & (g972) & (g973)) + ((!g683) & (!g868) & (!g946) & (g961) & (!g972) & (!g973)) + ((!g683) & (!g868) & (!g946) & (g961) & (g972) & (!g973)) + ((!g683) & (!g868) & (g946) & (!g961) & (!g972) & (!g973)) + ((!g683) & (!g868) & (g946) & (!g961) & (g972) & (!g973)) + ((!g683) & (!g868) & (g946) & (g961) & (!g972) & (g973)) + ((!g683) & (!g868) & (g946) & (g961) & (g972) & (g973)) + ((!g683) & (g868) & (!g946) & (!g961) & (g972) & (g973)) + ((!g683) & (g868) & (!g946) & (g961) & (!g972) & (!g973)) + ((!g683) & (g868) & (!g946) & (g961) & (!g972) & (g973)) + ((!g683) & (g868) & (!g946) & (g961) & (g972) & (!g973)) + ((!g683) & (g868) & (g946) & (!g961) & (!g972) & (!g973)) + ((!g683) & (g868) & (g946) & (!g961) & (!g972) & (g973)) + ((!g683) & (g868) & (g946) & (!g961) & (g972) & (!g973)) + ((!g683) & (g868) & (g946) & (g961) & (g972) & (g973)) + ((g683) & (!g868) & (!g946) & (!g961) & (!g972) & (!g973)) + ((g683) & (!g868) & (!g946) & (!g961) & (g972) & (!g973)) + ((g683) & (!g868) & (!g946) & (g961) & (!g972) & (g973)) + ((g683) & (!g868) & (!g946) & (g961) & (g972) & (g973)) + ((g683) & (!g868) & (g946) & (!g961) & (!g972) & (g973)) + ((g683) & (!g868) & (g946) & (!g961) & (g972) & (g973)) + ((g683) & (!g868) & (g946) & (g961) & (!g972) & (!g973)) + ((g683) & (!g868) & (g946) & (g961) & (g972) & (!g973)) + ((g683) & (g868) & (!g946) & (!g961) & (!g972) & (!g973)) + ((g683) & (g868) & (!g946) & (!g961) & (!g972) & (g973)) + ((g683) & (g868) & (!g946) & (!g961) & (g972) & (!g973)) + ((g683) & (g868) & (!g946) & (g961) & (g972) & (g973)) + ((g683) & (g868) & (g946) & (!g961) & (g972) & (g973)) + ((g683) & (g868) & (g946) & (g961) & (!g972) & (!g973)) + ((g683) & (g868) & (g946) & (g961) & (!g972) & (g973)) + ((g683) & (g868) & (g946) & (g961) & (g972) & (!g973)));
	assign g1012 = (((!g70) & (!g49) & (!sk[126]) & (!g62) & (g42) & (!g233)) + ((!g70) & (!g49) & (!sk[126]) & (!g62) & (g42) & (g233)) + ((!g70) & (!g49) & (!sk[126]) & (g62) & (!g42) & (!g233)) + ((!g70) & (!g49) & (!sk[126]) & (g62) & (!g42) & (g233)) + ((!g70) & (!g49) & (!sk[126]) & (g62) & (g42) & (!g233)) + ((!g70) & (!g49) & (!sk[126]) & (g62) & (g42) & (g233)) + ((!g70) & (!g49) & (sk[126]) & (!g62) & (!g42) & (!g233)) + ((!g70) & (!g49) & (sk[126]) & (!g62) & (g42) & (!g233)) + ((!g70) & (!g49) & (sk[126]) & (g62) & (!g42) & (!g233)) + ((!g70) & (g49) & (!sk[126]) & (!g62) & (!g42) & (!g233)) + ((!g70) & (g49) & (!sk[126]) & (!g62) & (!g42) & (g233)) + ((!g70) & (g49) & (!sk[126]) & (!g62) & (g42) & (!g233)) + ((!g70) & (g49) & (!sk[126]) & (!g62) & (g42) & (g233)) + ((!g70) & (g49) & (!sk[126]) & (g62) & (!g42) & (!g233)) + ((!g70) & (g49) & (!sk[126]) & (g62) & (!g42) & (g233)) + ((!g70) & (g49) & (!sk[126]) & (g62) & (g42) & (!g233)) + ((!g70) & (g49) & (!sk[126]) & (g62) & (g42) & (g233)) + ((!g70) & (g49) & (sk[126]) & (!g62) & (!g42) & (!g233)) + ((!g70) & (g49) & (sk[126]) & (!g62) & (g42) & (!g233)) + ((g70) & (!g49) & (!sk[126]) & (!g62) & (g42) & (!g233)) + ((g70) & (!g49) & (!sk[126]) & (!g62) & (g42) & (g233)) + ((g70) & (!g49) & (!sk[126]) & (g62) & (!g42) & (!g233)) + ((g70) & (!g49) & (!sk[126]) & (g62) & (!g42) & (g233)) + ((g70) & (!g49) & (!sk[126]) & (g62) & (g42) & (!g233)) + ((g70) & (!g49) & (!sk[126]) & (g62) & (g42) & (g233)) + ((g70) & (!g49) & (sk[126]) & (!g62) & (!g42) & (!g233)) + ((g70) & (!g49) & (sk[126]) & (g62) & (!g42) & (!g233)) + ((g70) & (g49) & (!sk[126]) & (!g62) & (!g42) & (!g233)) + ((g70) & (g49) & (!sk[126]) & (!g62) & (!g42) & (g233)) + ((g70) & (g49) & (!sk[126]) & (!g62) & (g42) & (!g233)) + ((g70) & (g49) & (!sk[126]) & (!g62) & (g42) & (g233)) + ((g70) & (g49) & (!sk[126]) & (g62) & (!g42) & (!g233)) + ((g70) & (g49) & (!sk[126]) & (g62) & (!g42) & (g233)) + ((g70) & (g49) & (!sk[126]) & (g62) & (g42) & (!g233)) + ((g70) & (g49) & (!sk[126]) & (g62) & (g42) & (g233)) + ((g70) & (g49) & (sk[126]) & (!g62) & (!g42) & (!g233)));
	assign g1013 = (((!g601) & (!sk[127]) & (g73) & (!g613)) + ((!g601) & (!sk[127]) & (g73) & (g613)) + ((!g601) & (sk[127]) & (!g73) & (g613)) + ((g601) & (!sk[127]) & (g73) & (!g613)) + ((g601) & (!sk[127]) & (g73) & (g613)));
	assign g1014 = (((!g254) & (!g340) & (!sk[0]) & (!g353) & (g1012) & (!g1013)) + ((!g254) & (!g340) & (!sk[0]) & (!g353) & (g1012) & (g1013)) + ((!g254) & (!g340) & (!sk[0]) & (g353) & (!g1012) & (!g1013)) + ((!g254) & (!g340) & (!sk[0]) & (g353) & (!g1012) & (g1013)) + ((!g254) & (!g340) & (!sk[0]) & (g353) & (g1012) & (!g1013)) + ((!g254) & (!g340) & (!sk[0]) & (g353) & (g1012) & (g1013)) + ((!g254) & (!g340) & (sk[0]) & (!g353) & (g1012) & (g1013)) + ((!g254) & (g340) & (!sk[0]) & (!g353) & (!g1012) & (!g1013)) + ((!g254) & (g340) & (!sk[0]) & (!g353) & (!g1012) & (g1013)) + ((!g254) & (g340) & (!sk[0]) & (!g353) & (g1012) & (!g1013)) + ((!g254) & (g340) & (!sk[0]) & (!g353) & (g1012) & (g1013)) + ((!g254) & (g340) & (!sk[0]) & (g353) & (!g1012) & (!g1013)) + ((!g254) & (g340) & (!sk[0]) & (g353) & (!g1012) & (g1013)) + ((!g254) & (g340) & (!sk[0]) & (g353) & (g1012) & (!g1013)) + ((!g254) & (g340) & (!sk[0]) & (g353) & (g1012) & (g1013)) + ((g254) & (!g340) & (!sk[0]) & (!g353) & (g1012) & (!g1013)) + ((g254) & (!g340) & (!sk[0]) & (!g353) & (g1012) & (g1013)) + ((g254) & (!g340) & (!sk[0]) & (g353) & (!g1012) & (!g1013)) + ((g254) & (!g340) & (!sk[0]) & (g353) & (!g1012) & (g1013)) + ((g254) & (!g340) & (!sk[0]) & (g353) & (g1012) & (!g1013)) + ((g254) & (!g340) & (!sk[0]) & (g353) & (g1012) & (g1013)) + ((g254) & (g340) & (!sk[0]) & (!g353) & (!g1012) & (!g1013)) + ((g254) & (g340) & (!sk[0]) & (!g353) & (!g1012) & (g1013)) + ((g254) & (g340) & (!sk[0]) & (!g353) & (g1012) & (!g1013)) + ((g254) & (g340) & (!sk[0]) & (!g353) & (g1012) & (g1013)) + ((g254) & (g340) & (!sk[0]) & (g353) & (!g1012) & (!g1013)) + ((g254) & (g340) & (!sk[0]) & (g353) & (!g1012) & (g1013)) + ((g254) & (g340) & (!sk[0]) & (g353) & (g1012) & (!g1013)) + ((g254) & (g340) & (!sk[0]) & (g353) & (g1012) & (g1013)));
	assign g1015 = (((!g71) & (!g20) & (!sk[1]) & (!g36) & (g278) & (!g1014)) + ((!g71) & (!g20) & (!sk[1]) & (!g36) & (g278) & (g1014)) + ((!g71) & (!g20) & (!sk[1]) & (g36) & (!g278) & (!g1014)) + ((!g71) & (!g20) & (!sk[1]) & (g36) & (!g278) & (g1014)) + ((!g71) & (!g20) & (!sk[1]) & (g36) & (g278) & (!g1014)) + ((!g71) & (!g20) & (!sk[1]) & (g36) & (g278) & (g1014)) + ((!g71) & (!g20) & (sk[1]) & (!g36) & (g278) & (g1014)) + ((!g71) & (g20) & (!sk[1]) & (!g36) & (!g278) & (!g1014)) + ((!g71) & (g20) & (!sk[1]) & (!g36) & (!g278) & (g1014)) + ((!g71) & (g20) & (!sk[1]) & (!g36) & (g278) & (!g1014)) + ((!g71) & (g20) & (!sk[1]) & (!g36) & (g278) & (g1014)) + ((!g71) & (g20) & (!sk[1]) & (g36) & (!g278) & (!g1014)) + ((!g71) & (g20) & (!sk[1]) & (g36) & (!g278) & (g1014)) + ((!g71) & (g20) & (!sk[1]) & (g36) & (g278) & (!g1014)) + ((!g71) & (g20) & (!sk[1]) & (g36) & (g278) & (g1014)) + ((!g71) & (g20) & (sk[1]) & (!g36) & (g278) & (g1014)) + ((g71) & (!g20) & (!sk[1]) & (!g36) & (g278) & (!g1014)) + ((g71) & (!g20) & (!sk[1]) & (!g36) & (g278) & (g1014)) + ((g71) & (!g20) & (!sk[1]) & (g36) & (!g278) & (!g1014)) + ((g71) & (!g20) & (!sk[1]) & (g36) & (!g278) & (g1014)) + ((g71) & (!g20) & (!sk[1]) & (g36) & (g278) & (!g1014)) + ((g71) & (!g20) & (!sk[1]) & (g36) & (g278) & (g1014)) + ((g71) & (!g20) & (sk[1]) & (!g36) & (g278) & (g1014)) + ((g71) & (g20) & (!sk[1]) & (!g36) & (!g278) & (!g1014)) + ((g71) & (g20) & (!sk[1]) & (!g36) & (!g278) & (g1014)) + ((g71) & (g20) & (!sk[1]) & (!g36) & (g278) & (!g1014)) + ((g71) & (g20) & (!sk[1]) & (!g36) & (g278) & (g1014)) + ((g71) & (g20) & (!sk[1]) & (g36) & (!g278) & (!g1014)) + ((g71) & (g20) & (!sk[1]) & (g36) & (!g278) & (g1014)) + ((g71) & (g20) & (!sk[1]) & (g36) & (g278) & (!g1014)) + ((g71) & (g20) & (!sk[1]) & (g36) & (g278) & (g1014)));
	assign g1016 = (((!g38) & (!sk[2]) & (!g99) & (!g62) & (g18) & (!g104)) + ((!g38) & (!sk[2]) & (!g99) & (!g62) & (g18) & (g104)) + ((!g38) & (!sk[2]) & (!g99) & (g62) & (!g18) & (!g104)) + ((!g38) & (!sk[2]) & (!g99) & (g62) & (!g18) & (g104)) + ((!g38) & (!sk[2]) & (!g99) & (g62) & (g18) & (!g104)) + ((!g38) & (!sk[2]) & (!g99) & (g62) & (g18) & (g104)) + ((!g38) & (!sk[2]) & (g99) & (!g62) & (!g18) & (!g104)) + ((!g38) & (!sk[2]) & (g99) & (!g62) & (!g18) & (g104)) + ((!g38) & (!sk[2]) & (g99) & (!g62) & (g18) & (!g104)) + ((!g38) & (!sk[2]) & (g99) & (!g62) & (g18) & (g104)) + ((!g38) & (!sk[2]) & (g99) & (g62) & (!g18) & (!g104)) + ((!g38) & (!sk[2]) & (g99) & (g62) & (!g18) & (g104)) + ((!g38) & (!sk[2]) & (g99) & (g62) & (g18) & (!g104)) + ((!g38) & (!sk[2]) & (g99) & (g62) & (g18) & (g104)) + ((!g38) & (sk[2]) & (!g99) & (!g62) & (!g18) & (!g104)) + ((!g38) & (sk[2]) & (!g99) & (!g62) & (!g18) & (g104)) + ((!g38) & (sk[2]) & (!g99) & (!g62) & (g18) & (!g104)) + ((!g38) & (sk[2]) & (!g99) & (!g62) & (g18) & (g104)) + ((!g38) & (sk[2]) & (!g99) & (g62) & (!g18) & (!g104)) + ((!g38) & (sk[2]) & (!g99) & (g62) & (!g18) & (g104)) + ((!g38) & (sk[2]) & (!g99) & (g62) & (g18) & (!g104)) + ((!g38) & (sk[2]) & (!g99) & (g62) & (g18) & (g104)) + ((!g38) & (sk[2]) & (g99) & (!g62) & (!g18) & (!g104)) + ((!g38) & (sk[2]) & (g99) & (!g62) & (!g18) & (g104)) + ((!g38) & (sk[2]) & (g99) & (g62) & (!g18) & (!g104)) + ((!g38) & (sk[2]) & (g99) & (g62) & (!g18) & (g104)) + ((g38) & (!sk[2]) & (!g99) & (!g62) & (g18) & (!g104)) + ((g38) & (!sk[2]) & (!g99) & (!g62) & (g18) & (g104)) + ((g38) & (!sk[2]) & (!g99) & (g62) & (!g18) & (!g104)) + ((g38) & (!sk[2]) & (!g99) & (g62) & (!g18) & (g104)) + ((g38) & (!sk[2]) & (!g99) & (g62) & (g18) & (!g104)) + ((g38) & (!sk[2]) & (!g99) & (g62) & (g18) & (g104)) + ((g38) & (!sk[2]) & (g99) & (!g62) & (!g18) & (!g104)) + ((g38) & (!sk[2]) & (g99) & (!g62) & (!g18) & (g104)) + ((g38) & (!sk[2]) & (g99) & (!g62) & (g18) & (!g104)) + ((g38) & (!sk[2]) & (g99) & (!g62) & (g18) & (g104)) + ((g38) & (!sk[2]) & (g99) & (g62) & (!g18) & (!g104)) + ((g38) & (!sk[2]) & (g99) & (g62) & (!g18) & (g104)) + ((g38) & (!sk[2]) & (g99) & (g62) & (g18) & (!g104)) + ((g38) & (!sk[2]) & (g99) & (g62) & (g18) & (g104)) + ((g38) & (sk[2]) & (!g99) & (!g62) & (!g18) & (!g104)) + ((g38) & (sk[2]) & (!g99) & (!g62) & (g18) & (!g104)));
	assign g1017 = (((!g9) & (!g12) & (!g32) & (!sk[3]) & (g1016)) + ((!g9) & (!g12) & (!g32) & (sk[3]) & (g1016)) + ((!g9) & (!g12) & (g32) & (!sk[3]) & (g1016)) + ((!g9) & (!g12) & (g32) & (sk[3]) & (g1016)) + ((!g9) & (g12) & (!g32) & (!sk[3]) & (g1016)) + ((!g9) & (g12) & (!g32) & (sk[3]) & (g1016)) + ((!g9) & (g12) & (g32) & (!sk[3]) & (g1016)) + ((!g9) & (g12) & (g32) & (sk[3]) & (g1016)) + ((g9) & (!g12) & (!g32) & (!sk[3]) & (!g1016)) + ((g9) & (!g12) & (!g32) & (!sk[3]) & (g1016)) + ((g9) & (!g12) & (!g32) & (sk[3]) & (g1016)) + ((g9) & (!g12) & (g32) & (!sk[3]) & (!g1016)) + ((g9) & (!g12) & (g32) & (!sk[3]) & (g1016)) + ((g9) & (g12) & (!g32) & (!sk[3]) & (!g1016)) + ((g9) & (g12) & (!g32) & (!sk[3]) & (g1016)) + ((g9) & (g12) & (g32) & (!sk[3]) & (!g1016)) + ((g9) & (g12) & (g32) & (!sk[3]) & (g1016)));
	assign g1018 = (((!g10) & (!sk[4]) & (!g99) & (!g20) & (g101) & (!g174)) + ((!g10) & (!sk[4]) & (!g99) & (!g20) & (g101) & (g174)) + ((!g10) & (!sk[4]) & (!g99) & (g20) & (!g101) & (!g174)) + ((!g10) & (!sk[4]) & (!g99) & (g20) & (!g101) & (g174)) + ((!g10) & (!sk[4]) & (!g99) & (g20) & (g101) & (!g174)) + ((!g10) & (!sk[4]) & (!g99) & (g20) & (g101) & (g174)) + ((!g10) & (!sk[4]) & (g99) & (!g20) & (!g101) & (!g174)) + ((!g10) & (!sk[4]) & (g99) & (!g20) & (!g101) & (g174)) + ((!g10) & (!sk[4]) & (g99) & (!g20) & (g101) & (!g174)) + ((!g10) & (!sk[4]) & (g99) & (!g20) & (g101) & (g174)) + ((!g10) & (!sk[4]) & (g99) & (g20) & (!g101) & (!g174)) + ((!g10) & (!sk[4]) & (g99) & (g20) & (!g101) & (g174)) + ((!g10) & (!sk[4]) & (g99) & (g20) & (g101) & (!g174)) + ((!g10) & (!sk[4]) & (g99) & (g20) & (g101) & (g174)) + ((!g10) & (sk[4]) & (!g99) & (!g20) & (!g101) & (!g174)) + ((!g10) & (sk[4]) & (!g99) & (g20) & (!g101) & (!g174)) + ((!g10) & (sk[4]) & (g99) & (!g20) & (!g101) & (!g174)) + ((g10) & (!sk[4]) & (!g99) & (!g20) & (g101) & (!g174)) + ((g10) & (!sk[4]) & (!g99) & (!g20) & (g101) & (g174)) + ((g10) & (!sk[4]) & (!g99) & (g20) & (!g101) & (!g174)) + ((g10) & (!sk[4]) & (!g99) & (g20) & (!g101) & (g174)) + ((g10) & (!sk[4]) & (!g99) & (g20) & (g101) & (!g174)) + ((g10) & (!sk[4]) & (!g99) & (g20) & (g101) & (g174)) + ((g10) & (!sk[4]) & (g99) & (!g20) & (!g101) & (!g174)) + ((g10) & (!sk[4]) & (g99) & (!g20) & (!g101) & (g174)) + ((g10) & (!sk[4]) & (g99) & (!g20) & (g101) & (!g174)) + ((g10) & (!sk[4]) & (g99) & (!g20) & (g101) & (g174)) + ((g10) & (!sk[4]) & (g99) & (g20) & (!g101) & (!g174)) + ((g10) & (!sk[4]) & (g99) & (g20) & (!g101) & (g174)) + ((g10) & (!sk[4]) & (g99) & (g20) & (g101) & (!g174)) + ((g10) & (!sk[4]) & (g99) & (g20) & (g101) & (g174)) + ((g10) & (sk[4]) & (!g99) & (!g20) & (!g101) & (!g174)) + ((g10) & (sk[4]) & (!g99) & (g20) & (!g101) & (!g174)));
	assign g1019 = (((!g26) & (!sk[5]) & (!g51) & (!g274) & (g1017) & (!g1018)) + ((!g26) & (!sk[5]) & (!g51) & (!g274) & (g1017) & (g1018)) + ((!g26) & (!sk[5]) & (!g51) & (g274) & (!g1017) & (!g1018)) + ((!g26) & (!sk[5]) & (!g51) & (g274) & (!g1017) & (g1018)) + ((!g26) & (!sk[5]) & (!g51) & (g274) & (g1017) & (!g1018)) + ((!g26) & (!sk[5]) & (!g51) & (g274) & (g1017) & (g1018)) + ((!g26) & (!sk[5]) & (g51) & (!g274) & (!g1017) & (!g1018)) + ((!g26) & (!sk[5]) & (g51) & (!g274) & (!g1017) & (g1018)) + ((!g26) & (!sk[5]) & (g51) & (!g274) & (g1017) & (!g1018)) + ((!g26) & (!sk[5]) & (g51) & (!g274) & (g1017) & (g1018)) + ((!g26) & (!sk[5]) & (g51) & (g274) & (!g1017) & (!g1018)) + ((!g26) & (!sk[5]) & (g51) & (g274) & (!g1017) & (g1018)) + ((!g26) & (!sk[5]) & (g51) & (g274) & (g1017) & (!g1018)) + ((!g26) & (!sk[5]) & (g51) & (g274) & (g1017) & (g1018)) + ((!g26) & (sk[5]) & (!g51) & (g274) & (g1017) & (g1018)) + ((g26) & (!sk[5]) & (!g51) & (!g274) & (g1017) & (!g1018)) + ((g26) & (!sk[5]) & (!g51) & (!g274) & (g1017) & (g1018)) + ((g26) & (!sk[5]) & (!g51) & (g274) & (!g1017) & (!g1018)) + ((g26) & (!sk[5]) & (!g51) & (g274) & (!g1017) & (g1018)) + ((g26) & (!sk[5]) & (!g51) & (g274) & (g1017) & (!g1018)) + ((g26) & (!sk[5]) & (!g51) & (g274) & (g1017) & (g1018)) + ((g26) & (!sk[5]) & (g51) & (!g274) & (!g1017) & (!g1018)) + ((g26) & (!sk[5]) & (g51) & (!g274) & (!g1017) & (g1018)) + ((g26) & (!sk[5]) & (g51) & (!g274) & (g1017) & (!g1018)) + ((g26) & (!sk[5]) & (g51) & (!g274) & (g1017) & (g1018)) + ((g26) & (!sk[5]) & (g51) & (g274) & (!g1017) & (!g1018)) + ((g26) & (!sk[5]) & (g51) & (g274) & (!g1017) & (g1018)) + ((g26) & (!sk[5]) & (g51) & (g274) & (g1017) & (!g1018)) + ((g26) & (!sk[5]) & (g51) & (g274) & (g1017) & (g1018)));
	assign g1020 = (((!g38) & (!g9) & (!g71) & (!g25) & (!g137) & (!g133)) + ((!g38) & (!g9) & (!g71) & (!g25) & (!g137) & (g133)) + ((!g38) & (!g9) & (!g71) & (g25) & (!g137) & (!g133)) + ((!g38) & (!g9) & (!g71) & (g25) & (!g137) & (g133)) + ((!g38) & (!g9) & (g71) & (!g25) & (!g137) & (!g133)) + ((!g38) & (!g9) & (g71) & (!g25) & (!g137) & (g133)) + ((!g38) & (g9) & (!g71) & (!g25) & (!g137) & (!g133)) + ((!g38) & (g9) & (!g71) & (g25) & (!g137) & (!g133)) + ((!g38) & (g9) & (g71) & (!g25) & (!g137) & (!g133)) + ((g38) & (!g9) & (!g71) & (!g25) & (!g137) & (!g133)) + ((g38) & (!g9) & (!g71) & (!g25) & (!g137) & (g133)) + ((g38) & (!g9) & (!g71) & (g25) & (!g137) & (!g133)) + ((g38) & (!g9) & (!g71) & (g25) & (!g137) & (g133)) + ((g38) & (g9) & (!g71) & (!g25) & (!g137) & (!g133)) + ((g38) & (g9) & (!g71) & (g25) & (!g137) & (!g133)));
	assign g1021 = (((!g114) & (!g115) & (!g8) & (!g17) & (g25) & (!g41)) + ((!g114) & (!g115) & (!g8) & (!g17) & (g25) & (g41)) + ((!g114) & (!g115) & (!g8) & (g17) & (g25) & (!g41)) + ((!g114) & (!g115) & (!g8) & (g17) & (g25) & (g41)) + ((!g114) & (!g115) & (g8) & (!g17) & (g25) & (!g41)) + ((!g114) & (!g115) & (g8) & (!g17) & (g25) & (g41)) + ((!g114) & (!g115) & (g8) & (g17) & (g25) & (!g41)) + ((!g114) & (!g115) & (g8) & (g17) & (g25) & (g41)) + ((!g114) & (g115) & (!g8) & (!g17) & (!g25) & (g41)) + ((!g114) & (g115) & (!g8) & (!g17) & (g25) & (g41)) + ((!g114) & (g115) & (!g8) & (g17) & (!g25) & (g41)) + ((!g114) & (g115) & (!g8) & (g17) & (g25) & (g41)) + ((g114) & (!g115) & (!g8) & (!g17) & (!g25) & (g41)) + ((g114) & (!g115) & (!g8) & (!g17) & (g25) & (g41)) + ((g114) & (!g115) & (!g8) & (g17) & (!g25) & (!g41)) + ((g114) & (!g115) & (!g8) & (g17) & (!g25) & (g41)) + ((g114) & (!g115) & (!g8) & (g17) & (g25) & (!g41)) + ((g114) & (!g115) & (!g8) & (g17) & (g25) & (g41)) + ((g114) & (g115) & (g8) & (g17) & (!g25) & (!g41)) + ((g114) & (g115) & (g8) & (g17) & (!g25) & (g41)) + ((g114) & (g115) & (g8) & (g17) & (g25) & (!g41)) + ((g114) & (g115) & (g8) & (g17) & (g25) & (g41)));
	assign g1022 = (((!g667) & (!g1015) & (!g1019) & (!sk[8]) & (g1020) & (!g1021)) + ((!g667) & (!g1015) & (!g1019) & (!sk[8]) & (g1020) & (g1021)) + ((!g667) & (!g1015) & (g1019) & (!sk[8]) & (!g1020) & (!g1021)) + ((!g667) & (!g1015) & (g1019) & (!sk[8]) & (!g1020) & (g1021)) + ((!g667) & (!g1015) & (g1019) & (!sk[8]) & (g1020) & (!g1021)) + ((!g667) & (!g1015) & (g1019) & (!sk[8]) & (g1020) & (g1021)) + ((!g667) & (g1015) & (!g1019) & (!sk[8]) & (!g1020) & (!g1021)) + ((!g667) & (g1015) & (!g1019) & (!sk[8]) & (!g1020) & (g1021)) + ((!g667) & (g1015) & (!g1019) & (!sk[8]) & (g1020) & (!g1021)) + ((!g667) & (g1015) & (!g1019) & (!sk[8]) & (g1020) & (g1021)) + ((!g667) & (g1015) & (g1019) & (!sk[8]) & (!g1020) & (!g1021)) + ((!g667) & (g1015) & (g1019) & (!sk[8]) & (!g1020) & (g1021)) + ((!g667) & (g1015) & (g1019) & (!sk[8]) & (g1020) & (!g1021)) + ((!g667) & (g1015) & (g1019) & (!sk[8]) & (g1020) & (g1021)) + ((g667) & (!g1015) & (!g1019) & (!sk[8]) & (g1020) & (!g1021)) + ((g667) & (!g1015) & (!g1019) & (!sk[8]) & (g1020) & (g1021)) + ((g667) & (!g1015) & (g1019) & (!sk[8]) & (!g1020) & (!g1021)) + ((g667) & (!g1015) & (g1019) & (!sk[8]) & (!g1020) & (g1021)) + ((g667) & (!g1015) & (g1019) & (!sk[8]) & (g1020) & (!g1021)) + ((g667) & (!g1015) & (g1019) & (!sk[8]) & (g1020) & (g1021)) + ((g667) & (g1015) & (!g1019) & (!sk[8]) & (!g1020) & (!g1021)) + ((g667) & (g1015) & (!g1019) & (!sk[8]) & (!g1020) & (g1021)) + ((g667) & (g1015) & (!g1019) & (!sk[8]) & (g1020) & (!g1021)) + ((g667) & (g1015) & (!g1019) & (!sk[8]) & (g1020) & (g1021)) + ((g667) & (g1015) & (g1019) & (!sk[8]) & (!g1020) & (!g1021)) + ((g667) & (g1015) & (g1019) & (!sk[8]) & (!g1020) & (g1021)) + ((g667) & (g1015) & (g1019) & (!sk[8]) & (g1020) & (!g1021)) + ((g667) & (g1015) & (g1019) & (!sk[8]) & (g1020) & (g1021)) + ((g667) & (g1015) & (g1019) & (sk[8]) & (g1020) & (!g1021)));
	assign g1023 = (((!g16) & (!g66) & (!g289) & (!sk[9]) & (g152)) + ((!g16) & (!g66) & (g289) & (!sk[9]) & (g152)) + ((!g16) & (!g66) & (g289) & (sk[9]) & (!g152)) + ((!g16) & (g66) & (!g289) & (!sk[9]) & (g152)) + ((!g16) & (g66) & (g289) & (!sk[9]) & (g152)) + ((!g16) & (g66) & (g289) & (sk[9]) & (!g152)) + ((g16) & (!g66) & (!g289) & (!sk[9]) & (!g152)) + ((g16) & (!g66) & (!g289) & (!sk[9]) & (g152)) + ((g16) & (!g66) & (g289) & (!sk[9]) & (!g152)) + ((g16) & (!g66) & (g289) & (!sk[9]) & (g152)) + ((g16) & (!g66) & (g289) & (sk[9]) & (!g152)) + ((g16) & (g66) & (!g289) & (!sk[9]) & (!g152)) + ((g16) & (g66) & (!g289) & (!sk[9]) & (g152)) + ((g16) & (g66) & (g289) & (!sk[9]) & (!g152)) + ((g16) & (g66) & (g289) & (!sk[9]) & (g152)));
	assign g1024 = (((!sk[10]) & (!g153) & (g143) & (!g617)) + ((!sk[10]) & (!g153) & (g143) & (g617)) + ((!sk[10]) & (g153) & (g143) & (!g617)) + ((!sk[10]) & (g153) & (g143) & (g617)) + ((sk[10]) & (!g153) & (g143) & (g617)));
	assign g1025 = (((!g96) & (!g827) & (!g872) & (!sk[11]) & (g1023) & (!g1024)) + ((!g96) & (!g827) & (!g872) & (!sk[11]) & (g1023) & (g1024)) + ((!g96) & (!g827) & (g872) & (!sk[11]) & (!g1023) & (!g1024)) + ((!g96) & (!g827) & (g872) & (!sk[11]) & (!g1023) & (g1024)) + ((!g96) & (!g827) & (g872) & (!sk[11]) & (g1023) & (!g1024)) + ((!g96) & (!g827) & (g872) & (!sk[11]) & (g1023) & (g1024)) + ((!g96) & (g827) & (!g872) & (!sk[11]) & (!g1023) & (!g1024)) + ((!g96) & (g827) & (!g872) & (!sk[11]) & (!g1023) & (g1024)) + ((!g96) & (g827) & (!g872) & (!sk[11]) & (g1023) & (!g1024)) + ((!g96) & (g827) & (!g872) & (!sk[11]) & (g1023) & (g1024)) + ((!g96) & (g827) & (g872) & (!sk[11]) & (!g1023) & (!g1024)) + ((!g96) & (g827) & (g872) & (!sk[11]) & (!g1023) & (g1024)) + ((!g96) & (g827) & (g872) & (!sk[11]) & (g1023) & (!g1024)) + ((!g96) & (g827) & (g872) & (!sk[11]) & (g1023) & (g1024)) + ((g96) & (!g827) & (!g872) & (!sk[11]) & (g1023) & (!g1024)) + ((g96) & (!g827) & (!g872) & (!sk[11]) & (g1023) & (g1024)) + ((g96) & (!g827) & (g872) & (!sk[11]) & (!g1023) & (!g1024)) + ((g96) & (!g827) & (g872) & (!sk[11]) & (!g1023) & (g1024)) + ((g96) & (!g827) & (g872) & (!sk[11]) & (g1023) & (!g1024)) + ((g96) & (!g827) & (g872) & (!sk[11]) & (g1023) & (g1024)) + ((g96) & (g827) & (!g872) & (!sk[11]) & (!g1023) & (!g1024)) + ((g96) & (g827) & (!g872) & (!sk[11]) & (!g1023) & (g1024)) + ((g96) & (g827) & (!g872) & (!sk[11]) & (g1023) & (!g1024)) + ((g96) & (g827) & (!g872) & (!sk[11]) & (g1023) & (g1024)) + ((g96) & (g827) & (g872) & (!sk[11]) & (!g1023) & (!g1024)) + ((g96) & (g827) & (g872) & (!sk[11]) & (!g1023) & (g1024)) + ((g96) & (g827) & (g872) & (!sk[11]) & (g1023) & (!g1024)) + ((g96) & (g827) & (g872) & (!sk[11]) & (g1023) & (g1024)) + ((g96) & (g827) & (g872) & (sk[11]) & (g1023) & (g1024)));
	assign g1026 = (((!g70) & (!g99) & (!g12) & (!g30) & (!g71) & (!g58)) + ((!g70) & (!g99) & (!g12) & (!g30) & (!g71) & (g58)) + ((!g70) & (!g99) & (!g12) & (!g30) & (g71) & (!g58)) + ((!g70) & (!g99) & (!g12) & (g30) & (!g71) & (!g58)) + ((!g70) & (!g99) & (!g12) & (g30) & (!g71) & (g58)) + ((!g70) & (!g99) & (!g12) & (g30) & (g71) & (!g58)) + ((!g70) & (!g99) & (g12) & (!g30) & (!g71) & (!g58)) + ((!g70) & (!g99) & (g12) & (!g30) & (!g71) & (g58)) + ((!g70) & (!g99) & (g12) & (!g30) & (g71) & (!g58)) + ((!g70) & (!g99) & (g12) & (g30) & (!g71) & (!g58)) + ((!g70) & (!g99) & (g12) & (g30) & (!g71) & (g58)) + ((!g70) & (!g99) & (g12) & (g30) & (g71) & (!g58)) + ((!g70) & (g99) & (!g12) & (!g30) & (!g71) & (!g58)) + ((!g70) & (g99) & (!g12) & (!g30) & (!g71) & (g58)) + ((!g70) & (g99) & (!g12) & (!g30) & (g71) & (!g58)) + ((!g70) & (g99) & (!g12) & (g30) & (!g71) & (!g58)) + ((!g70) & (g99) & (!g12) & (g30) & (!g71) & (g58)) + ((!g70) & (g99) & (!g12) & (g30) & (g71) & (!g58)) + ((g70) & (!g99) & (!g12) & (!g30) & (!g71) & (!g58)) + ((g70) & (!g99) & (!g12) & (!g30) & (!g71) & (g58)) + ((g70) & (!g99) & (!g12) & (!g30) & (g71) & (!g58)) + ((g70) & (!g99) & (g12) & (!g30) & (!g71) & (!g58)) + ((g70) & (!g99) & (g12) & (!g30) & (!g71) & (g58)) + ((g70) & (!g99) & (g12) & (!g30) & (g71) & (!g58)) + ((g70) & (g99) & (!g12) & (!g30) & (!g71) & (!g58)) + ((g70) & (g99) & (!g12) & (!g30) & (!g71) & (g58)) + ((g70) & (g99) & (!g12) & (!g30) & (g71) & (!g58)));
	assign g1027 = (((!sk[13]) & (!g9) & (!g99) & (!g30) & (g40)) + ((!sk[13]) & (!g9) & (!g99) & (g30) & (g40)) + ((!sk[13]) & (!g9) & (g99) & (!g30) & (g40)) + ((!sk[13]) & (!g9) & (g99) & (g30) & (g40)) + ((!sk[13]) & (g9) & (!g99) & (!g30) & (!g40)) + ((!sk[13]) & (g9) & (!g99) & (!g30) & (g40)) + ((!sk[13]) & (g9) & (!g99) & (g30) & (!g40)) + ((!sk[13]) & (g9) & (!g99) & (g30) & (g40)) + ((!sk[13]) & (g9) & (g99) & (!g30) & (!g40)) + ((!sk[13]) & (g9) & (g99) & (!g30) & (g40)) + ((!sk[13]) & (g9) & (g99) & (g30) & (!g40)) + ((!sk[13]) & (g9) & (g99) & (g30) & (g40)) + ((sk[13]) & (!g9) & (g99) & (!g30) & (g40)) + ((sk[13]) & (!g9) & (g99) & (g30) & (g40)) + ((sk[13]) & (g9) & (!g99) & (g30) & (!g40)) + ((sk[13]) & (g9) & (!g99) & (g30) & (g40)) + ((sk[13]) & (g9) & (g99) & (!g30) & (g40)) + ((sk[13]) & (g9) & (g99) & (g30) & (!g40)) + ((sk[13]) & (g9) & (g99) & (g30) & (g40)));
	assign g1028 = (((!sk[14]) & (!g48) & (!g582) & (!g592) & (g1026) & (!g1027)) + ((!sk[14]) & (!g48) & (!g582) & (!g592) & (g1026) & (g1027)) + ((!sk[14]) & (!g48) & (!g582) & (g592) & (!g1026) & (!g1027)) + ((!sk[14]) & (!g48) & (!g582) & (g592) & (!g1026) & (g1027)) + ((!sk[14]) & (!g48) & (!g582) & (g592) & (g1026) & (!g1027)) + ((!sk[14]) & (!g48) & (!g582) & (g592) & (g1026) & (g1027)) + ((!sk[14]) & (!g48) & (g582) & (!g592) & (!g1026) & (!g1027)) + ((!sk[14]) & (!g48) & (g582) & (!g592) & (!g1026) & (g1027)) + ((!sk[14]) & (!g48) & (g582) & (!g592) & (g1026) & (!g1027)) + ((!sk[14]) & (!g48) & (g582) & (!g592) & (g1026) & (g1027)) + ((!sk[14]) & (!g48) & (g582) & (g592) & (!g1026) & (!g1027)) + ((!sk[14]) & (!g48) & (g582) & (g592) & (!g1026) & (g1027)) + ((!sk[14]) & (!g48) & (g582) & (g592) & (g1026) & (!g1027)) + ((!sk[14]) & (!g48) & (g582) & (g592) & (g1026) & (g1027)) + ((!sk[14]) & (g48) & (!g582) & (!g592) & (g1026) & (!g1027)) + ((!sk[14]) & (g48) & (!g582) & (!g592) & (g1026) & (g1027)) + ((!sk[14]) & (g48) & (!g582) & (g592) & (!g1026) & (!g1027)) + ((!sk[14]) & (g48) & (!g582) & (g592) & (!g1026) & (g1027)) + ((!sk[14]) & (g48) & (!g582) & (g592) & (g1026) & (!g1027)) + ((!sk[14]) & (g48) & (!g582) & (g592) & (g1026) & (g1027)) + ((!sk[14]) & (g48) & (g582) & (!g592) & (!g1026) & (!g1027)) + ((!sk[14]) & (g48) & (g582) & (!g592) & (!g1026) & (g1027)) + ((!sk[14]) & (g48) & (g582) & (!g592) & (g1026) & (!g1027)) + ((!sk[14]) & (g48) & (g582) & (!g592) & (g1026) & (g1027)) + ((!sk[14]) & (g48) & (g582) & (g592) & (!g1026) & (!g1027)) + ((!sk[14]) & (g48) & (g582) & (g592) & (!g1026) & (g1027)) + ((!sk[14]) & (g48) & (g582) & (g592) & (g1026) & (!g1027)) + ((!sk[14]) & (g48) & (g582) & (g592) & (g1026) & (g1027)) + ((sk[14]) & (g48) & (g582) & (g592) & (g1026) & (!g1027)));
	assign g1029 = (((!g270) & (!g623) & (!sk[15]) & (!g1025) & (g1028)) + ((!g270) & (!g623) & (!sk[15]) & (g1025) & (g1028)) + ((!g270) & (g623) & (!sk[15]) & (!g1025) & (g1028)) + ((!g270) & (g623) & (!sk[15]) & (g1025) & (g1028)) + ((g270) & (!g623) & (!sk[15]) & (!g1025) & (!g1028)) + ((g270) & (!g623) & (!sk[15]) & (!g1025) & (g1028)) + ((g270) & (!g623) & (!sk[15]) & (g1025) & (!g1028)) + ((g270) & (!g623) & (!sk[15]) & (g1025) & (g1028)) + ((g270) & (g623) & (!sk[15]) & (!g1025) & (!g1028)) + ((g270) & (g623) & (!sk[15]) & (!g1025) & (g1028)) + ((g270) & (g623) & (!sk[15]) & (g1025) & (!g1028)) + ((g270) & (g623) & (!sk[15]) & (g1025) & (g1028)) + ((g270) & (g623) & (sk[15]) & (g1025) & (g1028)));
	assign g1030 = (((!g856) & (!g894) & (!g945) & (!g1011) & (!g1022) & (!g1029)) + ((!g856) & (!g894) & (!g945) & (!g1011) & (!g1022) & (g1029)) + ((!g856) & (!g894) & (g945) & (!g1011) & (!g1022) & (!g1029)) + ((!g856) & (!g894) & (g945) & (!g1011) & (!g1022) & (g1029)) + ((!g856) & (!g894) & (g945) & (!g1011) & (g1022) & (!g1029)) + ((!g856) & (!g894) & (g945) & (g1011) & (!g1022) & (!g1029)) + ((!g856) & (g894) & (!g945) & (!g1011) & (!g1022) & (!g1029)) + ((!g856) & (g894) & (!g945) & (g1011) & (!g1022) & (!g1029)) + ((!g856) & (g894) & (!g945) & (g1011) & (!g1022) & (g1029)) + ((!g856) & (g894) & (!g945) & (g1011) & (g1022) & (!g1029)) + ((!g856) & (g894) & (g945) & (!g1011) & (!g1022) & (!g1029)) + ((!g856) & (g894) & (g945) & (!g1011) & (!g1022) & (g1029)) + ((g856) & (!g894) & (!g945) & (!g1011) & (!g1022) & (!g1029)) + ((g856) & (!g894) & (!g945) & (g1011) & (!g1022) & (!g1029)) + ((g856) & (!g894) & (!g945) & (g1011) & (!g1022) & (g1029)) + ((g856) & (!g894) & (!g945) & (g1011) & (g1022) & (!g1029)) + ((g856) & (!g894) & (g945) & (!g1011) & (!g1022) & (!g1029)) + ((g856) & (!g894) & (g945) & (!g1011) & (!g1022) & (g1029)) + ((g856) & (g894) & (!g945) & (g1011) & (!g1022) & (!g1029)) + ((g856) & (g894) & (!g945) & (g1011) & (!g1022) & (g1029)) + ((g856) & (g894) & (g945) & (!g1011) & (!g1022) & (!g1029)) + ((g856) & (g894) & (g945) & (g1011) & (!g1022) & (!g1029)) + ((g856) & (g894) & (g945) & (g1011) & (!g1022) & (g1029)) + ((g856) & (g894) & (g945) & (g1011) & (g1022) & (!g1029)));
	assign g1031 = (((!g975) & (!sk[17]) & (!g998) & (!g1010) & (g1030)) + ((!g975) & (!sk[17]) & (!g998) & (g1010) & (g1030)) + ((!g975) & (!sk[17]) & (g998) & (!g1010) & (g1030)) + ((!g975) & (!sk[17]) & (g998) & (g1010) & (g1030)) + ((!g975) & (sk[17]) & (!g998) & (!g1010) & (!g1030)) + ((!g975) & (sk[17]) & (!g998) & (!g1010) & (g1030)) + ((!g975) & (sk[17]) & (!g998) & (g1010) & (g1030)) + ((!g975) & (sk[17]) & (g998) & (!g1010) & (g1030)) + ((g975) & (!sk[17]) & (!g998) & (!g1010) & (!g1030)) + ((g975) & (!sk[17]) & (!g998) & (!g1010) & (g1030)) + ((g975) & (!sk[17]) & (!g998) & (g1010) & (!g1030)) + ((g975) & (!sk[17]) & (!g998) & (g1010) & (g1030)) + ((g975) & (!sk[17]) & (g998) & (!g1010) & (!g1030)) + ((g975) & (!sk[17]) & (g998) & (!g1010) & (g1030)) + ((g975) & (!sk[17]) & (g998) & (g1010) & (!g1030)) + ((g975) & (!sk[17]) & (g998) & (g1010) & (g1030)) + ((g975) & (sk[17]) & (!g998) & (!g1010) & (g1030)) + ((g975) & (sk[17]) & (g998) & (!g1010) & (!g1030)) + ((g975) & (sk[17]) & (g998) & (!g1010) & (g1030)) + ((g975) & (sk[17]) & (g998) & (g1010) & (g1030)));
	assign g1032 = (((!sk[18]) & (!g62) & (!g32) & (!g124) & (g95)) + ((!sk[18]) & (!g62) & (!g32) & (g124) & (g95)) + ((!sk[18]) & (!g62) & (g32) & (!g124) & (g95)) + ((!sk[18]) & (!g62) & (g32) & (g124) & (g95)) + ((!sk[18]) & (g62) & (!g32) & (!g124) & (!g95)) + ((!sk[18]) & (g62) & (!g32) & (!g124) & (g95)) + ((!sk[18]) & (g62) & (!g32) & (g124) & (!g95)) + ((!sk[18]) & (g62) & (!g32) & (g124) & (g95)) + ((!sk[18]) & (g62) & (g32) & (!g124) & (!g95)) + ((!sk[18]) & (g62) & (g32) & (!g124) & (g95)) + ((!sk[18]) & (g62) & (g32) & (g124) & (!g95)) + ((!sk[18]) & (g62) & (g32) & (g124) & (g95)) + ((sk[18]) & (!g62) & (!g32) & (!g124) & (!g95)) + ((sk[18]) & (!g62) & (g32) & (!g124) & (!g95)) + ((sk[18]) & (g62) & (!g32) & (!g124) & (!g95)));
	assign g1033 = (((!g114) & (!g115) & (!g8) & (g12) & (!sk[19]) & (!g32)) + ((!g114) & (!g115) & (!g8) & (g12) & (!sk[19]) & (g32)) + ((!g114) & (!g115) & (!g8) & (g12) & (sk[19]) & (!g32)) + ((!g114) & (!g115) & (!g8) & (g12) & (sk[19]) & (g32)) + ((!g114) & (!g115) & (g8) & (!g12) & (!sk[19]) & (!g32)) + ((!g114) & (!g115) & (g8) & (!g12) & (!sk[19]) & (g32)) + ((!g114) & (!g115) & (g8) & (!g12) & (sk[19]) & (g32)) + ((!g114) & (!g115) & (g8) & (g12) & (!sk[19]) & (!g32)) + ((!g114) & (!g115) & (g8) & (g12) & (!sk[19]) & (g32)) + ((!g114) & (!g115) & (g8) & (g12) & (sk[19]) & (g32)) + ((!g114) & (g115) & (!g8) & (!g12) & (!sk[19]) & (!g32)) + ((!g114) & (g115) & (!g8) & (!g12) & (!sk[19]) & (g32)) + ((!g114) & (g115) & (!g8) & (g12) & (!sk[19]) & (!g32)) + ((!g114) & (g115) & (!g8) & (g12) & (!sk[19]) & (g32)) + ((!g114) & (g115) & (g8) & (!g12) & (!sk[19]) & (!g32)) + ((!g114) & (g115) & (g8) & (!g12) & (!sk[19]) & (g32)) + ((!g114) & (g115) & (g8) & (g12) & (!sk[19]) & (!g32)) + ((!g114) & (g115) & (g8) & (g12) & (!sk[19]) & (g32)) + ((g114) & (!g115) & (!g8) & (!g12) & (sk[19]) & (g32)) + ((g114) & (!g115) & (!g8) & (g12) & (!sk[19]) & (!g32)) + ((g114) & (!g115) & (!g8) & (g12) & (!sk[19]) & (g32)) + ((g114) & (!g115) & (!g8) & (g12) & (sk[19]) & (g32)) + ((g114) & (!g115) & (g8) & (!g12) & (!sk[19]) & (!g32)) + ((g114) & (!g115) & (g8) & (!g12) & (!sk[19]) & (g32)) + ((g114) & (!g115) & (g8) & (g12) & (!sk[19]) & (!g32)) + ((g114) & (!g115) & (g8) & (g12) & (!sk[19]) & (g32)) + ((g114) & (!g115) & (g8) & (g12) & (sk[19]) & (!g32)) + ((g114) & (!g115) & (g8) & (g12) & (sk[19]) & (g32)) + ((g114) & (g115) & (!g8) & (!g12) & (!sk[19]) & (!g32)) + ((g114) & (g115) & (!g8) & (!g12) & (!sk[19]) & (g32)) + ((g114) & (g115) & (!g8) & (g12) & (!sk[19]) & (!g32)) + ((g114) & (g115) & (!g8) & (g12) & (!sk[19]) & (g32)) + ((g114) & (g115) & (g8) & (!g12) & (!sk[19]) & (!g32)) + ((g114) & (g115) & (g8) & (!g12) & (!sk[19]) & (g32)) + ((g114) & (g115) & (g8) & (g12) & (!sk[19]) & (!g32)) + ((g114) & (g115) & (g8) & (g12) & (!sk[19]) & (g32)));
	assign g1034 = (((!g104) & (!g27) & (!sk[20]) & (!g47) & (g1033)) + ((!g104) & (!g27) & (!sk[20]) & (g47) & (g1033)) + ((!g104) & (!g27) & (sk[20]) & (!g47) & (!g1033)) + ((!g104) & (g27) & (!sk[20]) & (!g47) & (g1033)) + ((!g104) & (g27) & (!sk[20]) & (g47) & (g1033)) + ((!g104) & (g27) & (sk[20]) & (!g47) & (!g1033)) + ((g104) & (!g27) & (!sk[20]) & (!g47) & (!g1033)) + ((g104) & (!g27) & (!sk[20]) & (!g47) & (g1033)) + ((g104) & (!g27) & (!sk[20]) & (g47) & (!g1033)) + ((g104) & (!g27) & (!sk[20]) & (g47) & (g1033)) + ((g104) & (!g27) & (sk[20]) & (!g47) & (!g1033)) + ((g104) & (g27) & (!sk[20]) & (!g47) & (!g1033)) + ((g104) & (g27) & (!sk[20]) & (!g47) & (g1033)) + ((g104) & (g27) & (!sk[20]) & (g47) & (!g1033)) + ((g104) & (g27) & (!sk[20]) & (g47) & (g1033)));
	assign g1035 = (((!g26) & (!sk[21]) & (!g51) & (!g1000) & (g1034)) + ((!g26) & (!sk[21]) & (!g51) & (g1000) & (g1034)) + ((!g26) & (!sk[21]) & (g51) & (!g1000) & (g1034)) + ((!g26) & (!sk[21]) & (g51) & (g1000) & (g1034)) + ((!g26) & (sk[21]) & (!g51) & (!g1000) & (g1034)) + ((g26) & (!sk[21]) & (!g51) & (!g1000) & (!g1034)) + ((g26) & (!sk[21]) & (!g51) & (!g1000) & (g1034)) + ((g26) & (!sk[21]) & (!g51) & (g1000) & (!g1034)) + ((g26) & (!sk[21]) & (!g51) & (g1000) & (g1034)) + ((g26) & (!sk[21]) & (g51) & (!g1000) & (!g1034)) + ((g26) & (!sk[21]) & (g51) & (!g1000) & (g1034)) + ((g26) & (!sk[21]) & (g51) & (g1000) & (!g1034)) + ((g26) & (!sk[21]) & (g51) & (g1000) & (g1034)));
	assign g1036 = (((!sk[22]) & (!g70) & (!g10) & (!g16) & (g66) & (!g20)) + ((!sk[22]) & (!g70) & (!g10) & (!g16) & (g66) & (g20)) + ((!sk[22]) & (!g70) & (!g10) & (g16) & (!g66) & (!g20)) + ((!sk[22]) & (!g70) & (!g10) & (g16) & (!g66) & (g20)) + ((!sk[22]) & (!g70) & (!g10) & (g16) & (g66) & (!g20)) + ((!sk[22]) & (!g70) & (!g10) & (g16) & (g66) & (g20)) + ((!sk[22]) & (!g70) & (g10) & (!g16) & (!g66) & (!g20)) + ((!sk[22]) & (!g70) & (g10) & (!g16) & (!g66) & (g20)) + ((!sk[22]) & (!g70) & (g10) & (!g16) & (g66) & (!g20)) + ((!sk[22]) & (!g70) & (g10) & (!g16) & (g66) & (g20)) + ((!sk[22]) & (!g70) & (g10) & (g16) & (!g66) & (!g20)) + ((!sk[22]) & (!g70) & (g10) & (g16) & (!g66) & (g20)) + ((!sk[22]) & (!g70) & (g10) & (g16) & (g66) & (!g20)) + ((!sk[22]) & (!g70) & (g10) & (g16) & (g66) & (g20)) + ((!sk[22]) & (g70) & (!g10) & (!g16) & (g66) & (!g20)) + ((!sk[22]) & (g70) & (!g10) & (!g16) & (g66) & (g20)) + ((!sk[22]) & (g70) & (!g10) & (g16) & (!g66) & (!g20)) + ((!sk[22]) & (g70) & (!g10) & (g16) & (!g66) & (g20)) + ((!sk[22]) & (g70) & (!g10) & (g16) & (g66) & (!g20)) + ((!sk[22]) & (g70) & (!g10) & (g16) & (g66) & (g20)) + ((!sk[22]) & (g70) & (g10) & (!g16) & (!g66) & (!g20)) + ((!sk[22]) & (g70) & (g10) & (!g16) & (!g66) & (g20)) + ((!sk[22]) & (g70) & (g10) & (!g16) & (g66) & (!g20)) + ((!sk[22]) & (g70) & (g10) & (!g16) & (g66) & (g20)) + ((!sk[22]) & (g70) & (g10) & (g16) & (!g66) & (!g20)) + ((!sk[22]) & (g70) & (g10) & (g16) & (!g66) & (g20)) + ((!sk[22]) & (g70) & (g10) & (g16) & (g66) & (!g20)) + ((!sk[22]) & (g70) & (g10) & (g16) & (g66) & (g20)) + ((sk[22]) & (!g70) & (!g10) & (!g16) & (!g66) & (!g20)) + ((sk[22]) & (!g70) & (!g10) & (!g16) & (!g66) & (g20)) + ((sk[22]) & (!g70) & (!g10) & (!g16) & (g66) & (!g20)) + ((sk[22]) & (!g70) & (!g10) & (!g16) & (g66) & (g20)) + ((sk[22]) & (!g70) & (!g10) & (g16) & (!g66) & (!g20)) + ((sk[22]) & (!g70) & (!g10) & (g16) & (!g66) & (g20)) + ((sk[22]) & (!g70) & (g10) & (!g16) & (!g66) & (!g20)) + ((sk[22]) & (!g70) & (g10) & (!g16) & (!g66) & (g20)) + ((sk[22]) & (!g70) & (g10) & (!g16) & (g66) & (!g20)) + ((sk[22]) & (!g70) & (g10) & (!g16) & (g66) & (g20)) + ((sk[22]) & (!g70) & (g10) & (g16) & (!g66) & (!g20)) + ((sk[22]) & (!g70) & (g10) & (g16) & (!g66) & (g20)) + ((sk[22]) & (g70) & (!g10) & (!g16) & (!g66) & (!g20)) + ((sk[22]) & (g70) & (!g10) & (!g16) & (g66) & (!g20)) + ((sk[22]) & (g70) & (!g10) & (g16) & (!g66) & (!g20)));
	assign g1037 = (((!g83) & (!g84) & (g1032) & (g830) & (g1035) & (g1036)));
	assign g1038 = (((!g236) & (!sk[24]) & (g642) & (!g999)) + ((!g236) & (!sk[24]) & (g642) & (g999)) + ((!g236) & (sk[24]) & (!g642) & (g999)) + ((g236) & (!sk[24]) & (g642) & (!g999)) + ((g236) & (!sk[24]) & (g642) & (g999)));
	assign g1039 = (((!g275) & (!g352) & (!g362) & (!sk[25]) & (g1037) & (!g1038)) + ((!g275) & (!g352) & (!g362) & (!sk[25]) & (g1037) & (g1038)) + ((!g275) & (!g352) & (g362) & (!sk[25]) & (!g1037) & (!g1038)) + ((!g275) & (!g352) & (g362) & (!sk[25]) & (!g1037) & (g1038)) + ((!g275) & (!g352) & (g362) & (!sk[25]) & (g1037) & (!g1038)) + ((!g275) & (!g352) & (g362) & (!sk[25]) & (g1037) & (g1038)) + ((!g275) & (g352) & (!g362) & (!sk[25]) & (!g1037) & (!g1038)) + ((!g275) & (g352) & (!g362) & (!sk[25]) & (!g1037) & (g1038)) + ((!g275) & (g352) & (!g362) & (!sk[25]) & (g1037) & (!g1038)) + ((!g275) & (g352) & (!g362) & (!sk[25]) & (g1037) & (g1038)) + ((!g275) & (g352) & (g362) & (!sk[25]) & (!g1037) & (!g1038)) + ((!g275) & (g352) & (g362) & (!sk[25]) & (!g1037) & (g1038)) + ((!g275) & (g352) & (g362) & (!sk[25]) & (g1037) & (!g1038)) + ((!g275) & (g352) & (g362) & (!sk[25]) & (g1037) & (g1038)) + ((!g275) & (g352) & (g362) & (sk[25]) & (g1037) & (g1038)) + ((g275) & (!g352) & (!g362) & (!sk[25]) & (g1037) & (!g1038)) + ((g275) & (!g352) & (!g362) & (!sk[25]) & (g1037) & (g1038)) + ((g275) & (!g352) & (g362) & (!sk[25]) & (!g1037) & (!g1038)) + ((g275) & (!g352) & (g362) & (!sk[25]) & (!g1037) & (g1038)) + ((g275) & (!g352) & (g362) & (!sk[25]) & (g1037) & (!g1038)) + ((g275) & (!g352) & (g362) & (!sk[25]) & (g1037) & (g1038)) + ((g275) & (g352) & (!g362) & (!sk[25]) & (!g1037) & (!g1038)) + ((g275) & (g352) & (!g362) & (!sk[25]) & (!g1037) & (g1038)) + ((g275) & (g352) & (!g362) & (!sk[25]) & (g1037) & (!g1038)) + ((g275) & (g352) & (!g362) & (!sk[25]) & (g1037) & (g1038)) + ((g275) & (g352) & (g362) & (!sk[25]) & (!g1037) & (!g1038)) + ((g275) & (g352) & (g362) & (!sk[25]) & (!g1037) & (g1038)) + ((g275) & (g352) & (g362) & (!sk[25]) & (g1037) & (!g1038)) + ((g275) & (g352) & (g362) & (!sk[25]) & (g1037) & (g1038)));
	assign g1040 = (((!g889) & (!g871) & (!g883) & (!g970) & (!g993) & (g1039)) + ((!g889) & (!g871) & (!g883) & (!g970) & (g993) & (g1039)) + ((!g889) & (!g871) & (!g883) & (g970) & (!g993) & (g1039)) + ((!g889) & (!g871) & (!g883) & (g970) & (g993) & (g1039)) + ((!g889) & (!g871) & (g883) & (!g970) & (!g993) & (g1039)) + ((!g889) & (!g871) & (g883) & (!g970) & (g993) & (g1039)) + ((!g889) & (!g871) & (g883) & (g970) & (!g993) & (g1039)) + ((!g889) & (!g871) & (g883) & (g970) & (g993) & (g1039)) + ((!g889) & (g871) & (!g883) & (!g970) & (!g993) & (g1039)) + ((!g889) & (g871) & (!g883) & (!g970) & (g993) & (g1039)) + ((!g889) & (g871) & (!g883) & (g970) & (!g993) & (g1039)) + ((!g889) & (g871) & (!g883) & (g970) & (g993) & (g1039)) + ((!g889) & (g871) & (g883) & (!g970) & (!g993) & (g1039)) + ((!g889) & (g871) & (g883) & (!g970) & (g993) & (g1039)) + ((!g889) & (g871) & (g883) & (g970) & (!g993) & (g1039)) + ((!g889) & (g871) & (g883) & (g970) & (g993) & (g1039)) + ((g889) & (!g871) & (!g883) & (!g970) & (!g993) & (g1039)) + ((g889) & (!g871) & (!g883) & (!g970) & (g993) & (g1039)) + ((g889) & (!g871) & (!g883) & (g970) & (!g993) & (g1039)) + ((g889) & (!g871) & (!g883) & (g970) & (g993) & (g1039)) + ((g889) & (!g871) & (g883) & (!g970) & (!g993) & (g1039)) + ((g889) & (!g871) & (g883) & (!g970) & (g993) & (g1039)) + ((g889) & (!g871) & (g883) & (g970) & (!g993) & (g1039)) + ((g889) & (!g871) & (g883) & (g970) & (g993) & (g1039)) + ((g889) & (g871) & (!g883) & (!g970) & (!g993) & (g1039)) + ((g889) & (g871) & (!g883) & (!g970) & (g993) & (g1039)) + ((g889) & (g871) & (!g883) & (g970) & (!g993) & (g1039)) + ((g889) & (g871) & (!g883) & (g970) & (g993) & (g1039)) + ((g889) & (g871) & (g883) & (!g970) & (!g993) & (g1039)) + ((g889) & (g871) & (g883) & (!g970) & (g993) & (g1039)) + ((g889) & (g871) & (g883) & (g970) & (!g993) & (g1039)) + ((g889) & (g871) & (g883) & (g970) & (g993) & (!g1039)));
	assign g1041 = (((!g962) & (!g963) & (!g884) & (!g971) & (!g994) & (g1040)) + ((!g962) & (!g963) & (!g884) & (!g971) & (g994) & (!g1040)) + ((!g962) & (!g963) & (!g884) & (g971) & (!g994) & (!g1040)) + ((!g962) & (!g963) & (!g884) & (g971) & (g994) & (g1040)) + ((!g962) & (!g963) & (g884) & (!g971) & (!g994) & (g1040)) + ((!g962) & (!g963) & (g884) & (!g971) & (g994) & (g1040)) + ((!g962) & (!g963) & (g884) & (g971) & (!g994) & (!g1040)) + ((!g962) & (!g963) & (g884) & (g971) & (g994) & (g1040)) + ((!g962) & (g963) & (!g884) & (!g971) & (!g994) & (g1040)) + ((!g962) & (g963) & (!g884) & (!g971) & (g994) & (g1040)) + ((!g962) & (g963) & (!g884) & (g971) & (!g994) & (!g1040)) + ((!g962) & (g963) & (!g884) & (g971) & (g994) & (g1040)) + ((!g962) & (g963) & (g884) & (!g971) & (!g994) & (g1040)) + ((!g962) & (g963) & (g884) & (!g971) & (g994) & (g1040)) + ((!g962) & (g963) & (g884) & (g971) & (!g994) & (!g1040)) + ((!g962) & (g963) & (g884) & (g971) & (g994) & (g1040)) + ((g962) & (!g963) & (!g884) & (!g971) & (!g994) & (g1040)) + ((g962) & (!g963) & (!g884) & (!g971) & (g994) & (!g1040)) + ((g962) & (!g963) & (!g884) & (g971) & (!g994) & (g1040)) + ((g962) & (!g963) & (!g884) & (g971) & (g994) & (g1040)) + ((g962) & (!g963) & (g884) & (!g971) & (!g994) & (g1040)) + ((g962) & (!g963) & (g884) & (!g971) & (g994) & (!g1040)) + ((g962) & (!g963) & (g884) & (g971) & (!g994) & (g1040)) + ((g962) & (!g963) & (g884) & (g971) & (g994) & (g1040)) + ((g962) & (g963) & (!g884) & (!g971) & (!g994) & (g1040)) + ((g962) & (g963) & (!g884) & (!g971) & (g994) & (!g1040)) + ((g962) & (g963) & (!g884) & (g971) & (!g994) & (g1040)) + ((g962) & (g963) & (!g884) & (g971) & (g994) & (g1040)) + ((g962) & (g963) & (g884) & (!g971) & (!g994) & (g1040)) + ((g962) & (g963) & (g884) & (!g971) & (g994) & (!g1040)) + ((g962) & (g963) & (g884) & (g971) & (!g994) & (!g1040)) + ((g962) & (g963) & (g884) & (g971) & (g994) & (g1040)));
	assign g1042 = (((!g891) & (!g892) & (!sk[28]) & (!g994) & (g1040)) + ((!g891) & (!g892) & (!sk[28]) & (g994) & (g1040)) + ((!g891) & (g892) & (!sk[28]) & (!g994) & (g1040)) + ((!g891) & (g892) & (!sk[28]) & (g994) & (g1040)) + ((!g891) & (g892) & (sk[28]) & (g994) & (!g1040)) + ((!g891) & (g892) & (sk[28]) & (g994) & (g1040)) + ((g891) & (!g892) & (!sk[28]) & (!g994) & (!g1040)) + ((g891) & (!g892) & (!sk[28]) & (!g994) & (g1040)) + ((g891) & (!g892) & (!sk[28]) & (g994) & (!g1040)) + ((g891) & (!g892) & (!sk[28]) & (g994) & (g1040)) + ((g891) & (!g892) & (sk[28]) & (!g994) & (!g1040)) + ((g891) & (!g892) & (sk[28]) & (g994) & (!g1040)) + ((g891) & (g892) & (!sk[28]) & (!g994) & (!g1040)) + ((g891) & (g892) & (!sk[28]) & (!g994) & (g1040)) + ((g891) & (g892) & (!sk[28]) & (g994) & (!g1040)) + ((g891) & (g892) & (!sk[28]) & (g994) & (g1040)) + ((g891) & (g892) & (sk[28]) & (!g994) & (!g1040)) + ((g891) & (g892) & (sk[28]) & (g994) & (!g1040)) + ((g891) & (g892) & (sk[28]) & (g994) & (g1040)));
	assign g1043 = (((!g683) & (!g864) & (!g868) & (!g971) & (!g1041) & (g1042)) + ((!g683) & (!g864) & (!g868) & (!g971) & (g1041) & (g1042)) + ((!g683) & (!g864) & (!g868) & (g971) & (!g1041) & (g1042)) + ((!g683) & (!g864) & (!g868) & (g971) & (g1041) & (g1042)) + ((!g683) & (!g864) & (g868) & (!g971) & (!g1041) & (!g1042)) + ((!g683) & (!g864) & (g868) & (!g971) & (!g1041) & (g1042)) + ((!g683) & (!g864) & (g868) & (!g971) & (g1041) & (g1042)) + ((!g683) & (!g864) & (g868) & (g971) & (!g1041) & (!g1042)) + ((!g683) & (!g864) & (g868) & (g971) & (!g1041) & (g1042)) + ((!g683) & (!g864) & (g868) & (g971) & (g1041) & (g1042)) + ((!g683) & (g864) & (!g868) & (!g971) & (!g1041) & (g1042)) + ((!g683) & (g864) & (!g868) & (!g971) & (g1041) & (g1042)) + ((!g683) & (g864) & (!g868) & (g971) & (!g1041) & (!g1042)) + ((!g683) & (g864) & (!g868) & (g971) & (!g1041) & (g1042)) + ((!g683) & (g864) & (!g868) & (g971) & (g1041) & (!g1042)) + ((!g683) & (g864) & (!g868) & (g971) & (g1041) & (g1042)) + ((!g683) & (g864) & (g868) & (!g971) & (!g1041) & (!g1042)) + ((!g683) & (g864) & (g868) & (!g971) & (!g1041) & (g1042)) + ((!g683) & (g864) & (g868) & (!g971) & (g1041) & (g1042)) + ((!g683) & (g864) & (g868) & (g971) & (!g1041) & (!g1042)) + ((!g683) & (g864) & (g868) & (g971) & (!g1041) & (g1042)) + ((!g683) & (g864) & (g868) & (g971) & (g1041) & (!g1042)) + ((!g683) & (g864) & (g868) & (g971) & (g1041) & (g1042)) + ((g683) & (!g864) & (!g868) & (!g971) & (!g1041) & (!g1042)) + ((g683) & (!g864) & (!g868) & (!g971) & (g1041) & (!g1042)) + ((g683) & (!g864) & (!g868) & (g971) & (!g1041) & (!g1042)) + ((g683) & (!g864) & (!g868) & (g971) & (g1041) & (!g1042)) + ((g683) & (!g864) & (g868) & (!g971) & (g1041) & (!g1042)) + ((g683) & (!g864) & (g868) & (g971) & (g1041) & (!g1042)) + ((g683) & (g864) & (!g868) & (!g971) & (!g1041) & (!g1042)) + ((g683) & (g864) & (!g868) & (!g971) & (g1041) & (!g1042)) + ((g683) & (g864) & (g868) & (!g971) & (g1041) & (!g1042)));
	assign g1044 = (((!g946) & (!g976) & (!g948) & (!g960) & (g978) & (g989)) + ((!g946) & (!g976) & (!g948) & (g960) & (g978) & (g989)) + ((!g946) & (!g976) & (g948) & (!g960) & (g978) & (g989)) + ((!g946) & (!g976) & (g948) & (g960) & (g978) & (g989)) + ((!g946) & (g976) & (!g948) & (!g960) & (!g978) & (g989)) + ((!g946) & (g976) & (!g948) & (!g960) & (g978) & (!g989)) + ((!g946) & (g976) & (!g948) & (!g960) & (g978) & (g989)) + ((!g946) & (g976) & (!g948) & (g960) & (g978) & (g989)) + ((!g946) & (g976) & (g948) & (!g960) & (g978) & (g989)) + ((!g946) & (g976) & (g948) & (g960) & (!g978) & (g989)) + ((!g946) & (g976) & (g948) & (g960) & (g978) & (!g989)) + ((!g946) & (g976) & (g948) & (g960) & (g978) & (g989)) + ((g946) & (!g976) & (!g948) & (!g960) & (!g978) & (g989)) + ((g946) & (!g976) & (!g948) & (!g960) & (g978) & (!g989)) + ((g946) & (!g976) & (!g948) & (!g960) & (g978) & (g989)) + ((g946) & (!g976) & (!g948) & (g960) & (g978) & (g989)) + ((g946) & (!g976) & (g948) & (!g960) & (g978) & (g989)) + ((g946) & (!g976) & (g948) & (g960) & (!g978) & (g989)) + ((g946) & (!g976) & (g948) & (g960) & (g978) & (!g989)) + ((g946) & (!g976) & (g948) & (g960) & (g978) & (g989)) + ((g946) & (g976) & (!g948) & (!g960) & (!g978) & (g989)) + ((g946) & (g976) & (!g948) & (!g960) & (g978) & (!g989)) + ((g946) & (g976) & (!g948) & (!g960) & (g978) & (g989)) + ((g946) & (g976) & (!g948) & (g960) & (!g978) & (g989)) + ((g946) & (g976) & (!g948) & (g960) & (g978) & (!g989)) + ((g946) & (g976) & (!g948) & (g960) & (g978) & (g989)) + ((g946) & (g976) & (g948) & (!g960) & (!g978) & (g989)) + ((g946) & (g976) & (g948) & (!g960) & (g978) & (!g989)) + ((g946) & (g976) & (g948) & (!g960) & (g978) & (g989)) + ((g946) & (g976) & (g948) & (g960) & (!g978) & (g989)) + ((g946) & (g976) & (g948) & (g960) & (g978) & (!g989)) + ((g946) & (g976) & (g948) & (g960) & (g978) & (g989)));
	assign g1045 = (((!g698) & (!g706) & (!g717) & (g747) & (!g825) & (!g832)) + ((!g698) & (!g706) & (!g717) & (g747) & (g825) & (g832)) + ((!g698) & (!g706) & (g717) & (g747) & (!g825) & (!g832)) + ((!g698) & (!g706) & (g717) & (g747) & (g825) & (g832)) + ((!g698) & (g706) & (!g717) & (g747) & (!g825) & (!g832)) + ((!g698) & (g706) & (!g717) & (g747) & (g825) & (g832)) + ((!g698) & (g706) & (g717) & (g747) & (!g825) & (g832)) + ((!g698) & (g706) & (g717) & (g747) & (g825) & (!g832)) + ((g698) & (!g706) & (!g717) & (g747) & (!g825) & (!g832)) + ((g698) & (!g706) & (!g717) & (g747) & (g825) & (g832)) + ((g698) & (!g706) & (g717) & (g747) & (!g825) & (g832)) + ((g698) & (!g706) & (g717) & (g747) & (g825) & (!g832)) + ((g698) & (g706) & (!g717) & (g747) & (!g825) & (g832)) + ((g698) & (g706) & (!g717) & (g747) & (g825) & (!g832)) + ((g698) & (g706) & (g717) & (g747) & (!g825) & (g832)) + ((g698) & (g706) & (g717) & (g747) & (g825) & (!g832)));
	assign g1046 = (((!g707) & (!g717) & (!g718) & (g744) & (!sk[32]) & (!g748)) + ((!g707) & (!g717) & (!g718) & (g744) & (!sk[32]) & (g748)) + ((!g707) & (!g717) & (g718) & (!g744) & (!sk[32]) & (!g748)) + ((!g707) & (!g717) & (g718) & (!g744) & (!sk[32]) & (g748)) + ((!g707) & (!g717) & (g718) & (!g744) & (sk[32]) & (g748)) + ((!g707) & (!g717) & (g718) & (g744) & (!sk[32]) & (!g748)) + ((!g707) & (!g717) & (g718) & (g744) & (!sk[32]) & (g748)) + ((!g707) & (!g717) & (g718) & (g744) & (sk[32]) & (g748)) + ((!g707) & (g717) & (!g718) & (!g744) & (!sk[32]) & (!g748)) + ((!g707) & (g717) & (!g718) & (!g744) & (!sk[32]) & (g748)) + ((!g707) & (g717) & (!g718) & (g744) & (!sk[32]) & (!g748)) + ((!g707) & (g717) & (!g718) & (g744) & (!sk[32]) & (g748)) + ((!g707) & (g717) & (!g718) & (g744) & (sk[32]) & (!g748)) + ((!g707) & (g717) & (!g718) & (g744) & (sk[32]) & (g748)) + ((!g707) & (g717) & (g718) & (!g744) & (!sk[32]) & (!g748)) + ((!g707) & (g717) & (g718) & (!g744) & (!sk[32]) & (g748)) + ((!g707) & (g717) & (g718) & (!g744) & (sk[32]) & (g748)) + ((!g707) & (g717) & (g718) & (g744) & (!sk[32]) & (!g748)) + ((!g707) & (g717) & (g718) & (g744) & (!sk[32]) & (g748)) + ((!g707) & (g717) & (g718) & (g744) & (sk[32]) & (!g748)) + ((!g707) & (g717) & (g718) & (g744) & (sk[32]) & (g748)) + ((g707) & (!g717) & (!g718) & (g744) & (!sk[32]) & (!g748)) + ((g707) & (!g717) & (!g718) & (g744) & (!sk[32]) & (g748)) + ((g707) & (!g717) & (!g718) & (g744) & (sk[32]) & (!g748)) + ((g707) & (!g717) & (!g718) & (g744) & (sk[32]) & (g748)) + ((g707) & (!g717) & (g718) & (!g744) & (!sk[32]) & (!g748)) + ((g707) & (!g717) & (g718) & (!g744) & (!sk[32]) & (g748)) + ((g707) & (!g717) & (g718) & (!g744) & (sk[32]) & (g748)) + ((g707) & (!g717) & (g718) & (g744) & (!sk[32]) & (!g748)) + ((g707) & (!g717) & (g718) & (g744) & (!sk[32]) & (g748)) + ((g707) & (!g717) & (g718) & (g744) & (sk[32]) & (!g748)) + ((g707) & (!g717) & (g718) & (g744) & (sk[32]) & (g748)) + ((g707) & (g717) & (!g718) & (!g744) & (!sk[32]) & (!g748)) + ((g707) & (g717) & (!g718) & (!g744) & (!sk[32]) & (g748)) + ((g707) & (g717) & (!g718) & (g744) & (!sk[32]) & (!g748)) + ((g707) & (g717) & (!g718) & (g744) & (!sk[32]) & (g748)) + ((g707) & (g717) & (g718) & (!g744) & (!sk[32]) & (!g748)) + ((g707) & (g717) & (g718) & (!g744) & (!sk[32]) & (g748)) + ((g707) & (g717) & (g718) & (!g744) & (sk[32]) & (g748)) + ((g707) & (g717) & (g718) & (g744) & (!sk[32]) & (!g748)) + ((g707) & (g717) & (g718) & (g744) & (!sk[32]) & (g748)) + ((g707) & (g717) & (g718) & (g744) & (sk[32]) & (g748)));
	assign g1047 = (((!g200) & (!g742) & (!g834) & (!g835) & (!g1045) & (g1046)) + ((!g200) & (!g742) & (!g834) & (!g835) & (g1045) & (!g1046)) + ((!g200) & (!g742) & (!g834) & (!g835) & (g1045) & (g1046)) + ((!g200) & (!g742) & (!g834) & (g835) & (!g1045) & (g1046)) + ((!g200) & (!g742) & (!g834) & (g835) & (g1045) & (!g1046)) + ((!g200) & (!g742) & (!g834) & (g835) & (g1045) & (g1046)) + ((!g200) & (!g742) & (g834) & (!g835) & (!g1045) & (g1046)) + ((!g200) & (!g742) & (g834) & (!g835) & (g1045) & (!g1046)) + ((!g200) & (!g742) & (g834) & (!g835) & (g1045) & (g1046)) + ((!g200) & (!g742) & (g834) & (g835) & (!g1045) & (g1046)) + ((!g200) & (!g742) & (g834) & (g835) & (g1045) & (!g1046)) + ((!g200) & (!g742) & (g834) & (g835) & (g1045) & (g1046)) + ((!g200) & (g742) & (!g834) & (!g835) & (!g1045) & (!g1046)) + ((!g200) & (g742) & (!g834) & (!g835) & (!g1045) & (g1046)) + ((!g200) & (g742) & (!g834) & (!g835) & (g1045) & (!g1046)) + ((!g200) & (g742) & (!g834) & (!g835) & (g1045) & (g1046)) + ((!g200) & (g742) & (!g834) & (g835) & (!g1045) & (g1046)) + ((!g200) & (g742) & (!g834) & (g835) & (g1045) & (!g1046)) + ((!g200) & (g742) & (!g834) & (g835) & (g1045) & (g1046)) + ((!g200) & (g742) & (g834) & (!g835) & (!g1045) & (g1046)) + ((!g200) & (g742) & (g834) & (!g835) & (g1045) & (!g1046)) + ((!g200) & (g742) & (g834) & (!g835) & (g1045) & (g1046)) + ((!g200) & (g742) & (g834) & (g835) & (!g1045) & (!g1046)) + ((!g200) & (g742) & (g834) & (g835) & (!g1045) & (g1046)) + ((!g200) & (g742) & (g834) & (g835) & (g1045) & (!g1046)) + ((!g200) & (g742) & (g834) & (g835) & (g1045) & (g1046)) + ((g200) & (!g742) & (!g834) & (!g835) & (!g1045) & (!g1046)) + ((g200) & (!g742) & (!g834) & (g835) & (!g1045) & (!g1046)) + ((g200) & (!g742) & (g834) & (!g835) & (!g1045) & (!g1046)) + ((g200) & (!g742) & (g834) & (g835) & (!g1045) & (!g1046)) + ((g200) & (g742) & (!g834) & (g835) & (!g1045) & (!g1046)) + ((g200) & (g742) & (g834) & (!g835) & (!g1045) & (!g1046)));
	assign g1048 = (((!g202) & (!g949) & (!g951) & (!g955) & (!g984) & (!g987)) + ((!g202) & (!g949) & (!g951) & (g955) & (!g984) & (!g987)) + ((!g202) & (!g949) & (g951) & (!g955) & (!g984) & (!g987)) + ((!g202) & (!g949) & (g951) & (!g955) & (!g984) & (g987)) + ((!g202) & (!g949) & (g951) & (!g955) & (g984) & (!g987)) + ((!g202) & (!g949) & (g951) & (g955) & (!g984) & (!g987)) + ((!g202) & (g949) & (!g951) & (!g955) & (!g984) & (!g987)) + ((!g202) & (g949) & (!g951) & (!g955) & (!g984) & (g987)) + ((!g202) & (g949) & (!g951) & (!g955) & (g984) & (!g987)) + ((!g202) & (g949) & (!g951) & (g955) & (!g984) & (!g987)) + ((!g202) & (g949) & (g951) & (!g955) & (!g984) & (!g987)) + ((!g202) & (g949) & (g951) & (!g955) & (!g984) & (g987)) + ((!g202) & (g949) & (g951) & (!g955) & (g984) & (!g987)) + ((!g202) & (g949) & (g951) & (g955) & (!g984) & (!g987)) + ((!g202) & (g949) & (g951) & (g955) & (!g984) & (g987)) + ((!g202) & (g949) & (g951) & (g955) & (g984) & (!g987)) + ((g202) & (!g949) & (!g951) & (!g955) & (g984) & (!g987)) + ((g202) & (!g949) & (!g951) & (g955) & (g984) & (!g987)) + ((g202) & (!g949) & (g951) & (!g955) & (!g984) & (!g987)) + ((g202) & (!g949) & (g951) & (!g955) & (g984) & (!g987)) + ((g202) & (!g949) & (g951) & (!g955) & (g984) & (g987)) + ((g202) & (!g949) & (g951) & (g955) & (g984) & (!g987)) + ((g202) & (g949) & (!g951) & (!g955) & (!g984) & (!g987)) + ((g202) & (g949) & (!g951) & (!g955) & (g984) & (!g987)) + ((g202) & (g949) & (!g951) & (!g955) & (g984) & (g987)) + ((g202) & (g949) & (!g951) & (g955) & (g984) & (!g987)) + ((g202) & (g949) & (g951) & (!g955) & (!g984) & (!g987)) + ((g202) & (g949) & (g951) & (!g955) & (g984) & (!g987)) + ((g202) & (g949) & (g951) & (!g955) & (g984) & (g987)) + ((g202) & (g949) & (g951) & (g955) & (!g984) & (!g987)) + ((g202) & (g949) & (g951) & (g955) & (g984) & (!g987)) + ((g202) & (g949) & (g951) & (g955) & (g984) & (g987)));
	assign g1049 = (((!g721) & (!g678) & (!g723) & (!sk[35]) & (g845) & (!g848)) + ((!g721) & (!g678) & (!g723) & (!sk[35]) & (g845) & (g848)) + ((!g721) & (!g678) & (!g723) & (sk[35]) & (!g845) & (g848)) + ((!g721) & (!g678) & (!g723) & (sk[35]) & (g845) & (!g848)) + ((!g721) & (!g678) & (!g723) & (sk[35]) & (g845) & (g848)) + ((!g721) & (!g678) & (g723) & (!sk[35]) & (!g845) & (!g848)) + ((!g721) & (!g678) & (g723) & (!sk[35]) & (!g845) & (g848)) + ((!g721) & (!g678) & (g723) & (!sk[35]) & (g845) & (!g848)) + ((!g721) & (!g678) & (g723) & (!sk[35]) & (g845) & (g848)) + ((!g721) & (!g678) & (g723) & (sk[35]) & (g845) & (!g848)) + ((!g721) & (!g678) & (g723) & (sk[35]) & (g845) & (g848)) + ((!g721) & (g678) & (!g723) & (!sk[35]) & (!g845) & (!g848)) + ((!g721) & (g678) & (!g723) & (!sk[35]) & (!g845) & (g848)) + ((!g721) & (g678) & (!g723) & (!sk[35]) & (g845) & (!g848)) + ((!g721) & (g678) & (!g723) & (!sk[35]) & (g845) & (g848)) + ((!g721) & (g678) & (!g723) & (sk[35]) & (!g845) & (g848)) + ((!g721) & (g678) & (!g723) & (sk[35]) & (g845) & (g848)) + ((!g721) & (g678) & (g723) & (!sk[35]) & (!g845) & (!g848)) + ((!g721) & (g678) & (g723) & (!sk[35]) & (!g845) & (g848)) + ((!g721) & (g678) & (g723) & (!sk[35]) & (g845) & (!g848)) + ((!g721) & (g678) & (g723) & (!sk[35]) & (g845) & (g848)) + ((g721) & (!g678) & (!g723) & (!sk[35]) & (g845) & (!g848)) + ((g721) & (!g678) & (!g723) & (!sk[35]) & (g845) & (g848)) + ((g721) & (!g678) & (!g723) & (sk[35]) & (!g845) & (g848)) + ((g721) & (!g678) & (!g723) & (sk[35]) & (g845) & (g848)) + ((g721) & (!g678) & (g723) & (!sk[35]) & (!g845) & (!g848)) + ((g721) & (!g678) & (g723) & (!sk[35]) & (!g845) & (g848)) + ((g721) & (!g678) & (g723) & (!sk[35]) & (g845) & (!g848)) + ((g721) & (!g678) & (g723) & (!sk[35]) & (g845) & (g848)) + ((g721) & (g678) & (!g723) & (!sk[35]) & (!g845) & (!g848)) + ((g721) & (g678) & (!g723) & (!sk[35]) & (!g845) & (g848)) + ((g721) & (g678) & (!g723) & (!sk[35]) & (g845) & (!g848)) + ((g721) & (g678) & (!g723) & (!sk[35]) & (g845) & (g848)) + ((g721) & (g678) & (!g723) & (sk[35]) & (!g845) & (g848)) + ((g721) & (g678) & (!g723) & (sk[35]) & (g845) & (!g848)) + ((g721) & (g678) & (!g723) & (sk[35]) & (g845) & (g848)) + ((g721) & (g678) & (g723) & (!sk[35]) & (!g845) & (!g848)) + ((g721) & (g678) & (g723) & (!sk[35]) & (!g845) & (g848)) + ((g721) & (g678) & (g723) & (!sk[35]) & (g845) & (!g848)) + ((g721) & (g678) & (g723) & (!sk[35]) & (g845) & (g848)) + ((g721) & (g678) & (g723) & (sk[35]) & (g845) & (!g848)) + ((g721) & (g678) & (g723) & (sk[35]) & (g845) & (g848)));
	assign g1050 = (((!g720) & (!g722) & (!g727) & (!g847) & (!g843) & (!g1049)) + ((!g720) & (!g722) & (!g727) & (g847) & (!g843) & (!g1049)) + ((!g720) & (!g722) & (g727) & (!g847) & (!g843) & (!g1049)) + ((!g720) & (!g722) & (g727) & (!g847) & (g843) & (!g1049)) + ((!g720) & (!g722) & (g727) & (g847) & (!g843) & (!g1049)) + ((!g720) & (!g722) & (g727) & (g847) & (g843) & (!g1049)) + ((!g720) & (g722) & (!g727) & (!g847) & (!g843) & (!g1049)) + ((!g720) & (g722) & (!g727) & (!g847) & (g843) & (!g1049)) + ((!g720) & (g722) & (!g727) & (g847) & (!g843) & (!g1049)) + ((!g720) & (g722) & (!g727) & (g847) & (g843) & (!g1049)) + ((!g720) & (g722) & (g727) & (!g847) & (!g843) & (!g1049)) + ((!g720) & (g722) & (g727) & (g847) & (!g843) & (!g1049)) + ((g720) & (!g722) & (!g727) & (!g847) & (!g843) & (!g1049)) + ((g720) & (!g722) & (!g727) & (!g847) & (g843) & (!g1049)) + ((g720) & (!g722) & (g727) & (!g847) & (!g843) & (!g1049)) + ((g720) & (g722) & (!g727) & (!g847) & (!g843) & (!g1049)) + ((g720) & (g722) & (g727) & (!g847) & (!g843) & (!g1049)) + ((g720) & (g722) & (g727) & (!g847) & (g843) & (!g1049)));
	assign g1051 = (((!g252) & (!g724) & (!g985) & (!g986) & (!g1447) & (!g1050)) + ((!g252) & (!g724) & (!g985) & (!g986) & (g1447) & (!g1050)) + ((!g252) & (!g724) & (!g985) & (g986) & (!g1447) & (g1050)) + ((!g252) & (!g724) & (!g985) & (g986) & (g1447) & (!g1050)) + ((!g252) & (!g724) & (g985) & (!g986) & (!g1447) & (!g1050)) + ((!g252) & (!g724) & (g985) & (!g986) & (g1447) & (g1050)) + ((!g252) & (!g724) & (g985) & (g986) & (!g1447) & (g1050)) + ((!g252) & (!g724) & (g985) & (g986) & (g1447) & (g1050)) + ((!g252) & (g724) & (!g985) & (!g986) & (!g1447) & (!g1050)) + ((!g252) & (g724) & (!g985) & (!g986) & (g1447) & (!g1050)) + ((!g252) & (g724) & (!g985) & (g986) & (!g1447) & (g1050)) + ((!g252) & (g724) & (!g985) & (g986) & (g1447) & (!g1050)) + ((!g252) & (g724) & (g985) & (!g986) & (!g1447) & (!g1050)) + ((!g252) & (g724) & (g985) & (!g986) & (g1447) & (g1050)) + ((!g252) & (g724) & (g985) & (g986) & (!g1447) & (g1050)) + ((!g252) & (g724) & (g985) & (g986) & (g1447) & (g1050)) + ((g252) & (!g724) & (!g985) & (!g986) & (!g1447) & (!g1050)) + ((g252) & (!g724) & (!g985) & (!g986) & (g1447) & (!g1050)) + ((g252) & (!g724) & (!g985) & (g986) & (!g1447) & (g1050)) + ((g252) & (!g724) & (!g985) & (g986) & (g1447) & (!g1050)) + ((g252) & (!g724) & (g985) & (!g986) & (!g1447) & (g1050)) + ((g252) & (!g724) & (g985) & (!g986) & (g1447) & (!g1050)) + ((g252) & (!g724) & (g985) & (g986) & (!g1447) & (g1050)) + ((g252) & (!g724) & (g985) & (g986) & (g1447) & (g1050)) + ((g252) & (g724) & (!g985) & (!g986) & (!g1447) & (g1050)) + ((g252) & (g724) & (!g985) & (!g986) & (g1447) & (g1050)) + ((g252) & (g724) & (!g985) & (g986) & (!g1447) & (!g1050)) + ((g252) & (g724) & (!g985) & (g986) & (g1447) & (g1050)) + ((g252) & (g724) & (g985) & (!g986) & (!g1447) & (!g1050)) + ((g252) & (g724) & (g985) & (!g986) & (g1447) & (g1050)) + ((g252) & (g724) & (g985) & (g986) & (!g1447) & (!g1050)) + ((g252) & (g724) & (g985) & (g986) & (g1447) & (!g1050)));
	assign g1052 = (((!g549) & (!g569) & (!g680) & (!g729) & (!g764) & (g762)) + ((!g549) & (!g569) & (!g680) & (!g729) & (g764) & (g762)) + ((!g549) & (!g569) & (g680) & (!g729) & (!g764) & (g762)) + ((!g549) & (!g569) & (g680) & (!g729) & (g764) & (!g762)) + ((!g549) & (!g569) & (g680) & (!g729) & (g764) & (g762)) + ((!g549) & (!g569) & (g680) & (g729) & (g764) & (!g762)) + ((!g549) & (!g569) & (g680) & (g729) & (g764) & (g762)) + ((!g549) & (g569) & (!g680) & (!g729) & (!g764) & (g762)) + ((!g549) & (g569) & (!g680) & (!g729) & (g764) & (!g762)) + ((!g549) & (g569) & (!g680) & (!g729) & (g764) & (g762)) + ((!g549) & (g569) & (!g680) & (g729) & (g764) & (!g762)) + ((!g549) & (g569) & (!g680) & (g729) & (g764) & (g762)) + ((!g549) & (g569) & (g680) & (!g729) & (!g764) & (g762)) + ((!g549) & (g569) & (g680) & (!g729) & (g764) & (g762)) + ((g549) & (!g569) & (!g680) & (!g729) & (!g764) & (g762)) + ((g549) & (!g569) & (!g680) & (!g729) & (g764) & (!g762)) + ((g549) & (!g569) & (!g680) & (!g729) & (g764) & (g762)) + ((g549) & (!g569) & (!g680) & (g729) & (g764) & (!g762)) + ((g549) & (!g569) & (!g680) & (g729) & (g764) & (g762)) + ((g549) & (!g569) & (g680) & (!g729) & (!g764) & (g762)) + ((g549) & (!g569) & (g680) & (!g729) & (g764) & (g762)) + ((g549) & (g569) & (!g680) & (!g729) & (!g764) & (g762)) + ((g549) & (g569) & (!g680) & (!g729) & (g764) & (g762)) + ((g549) & (g569) & (g680) & (!g729) & (!g764) & (g762)) + ((g549) & (g569) & (g680) & (!g729) & (g764) & (!g762)) + ((g549) & (g569) & (g680) & (!g729) & (g764) & (g762)) + ((g549) & (g569) & (g680) & (g729) & (g764) & (!g762)) + ((g549) & (g569) & (g680) & (g729) & (g764) & (g762)));
	assign g1053 = (((!g202) & (!g719) & (!g759) & (!g765) & (!g791) & (!g1052)) + ((!g202) & (!g719) & (!g759) & (!g765) & (g791) & (!g1052)) + ((!g202) & (!g719) & (g759) & (!g765) & (!g791) & (!g1052)) + ((!g202) & (g719) & (!g759) & (!g765) & (!g791) & (!g1052)) + ((!g202) & (g719) & (!g759) & (!g765) & (g791) & (!g1052)) + ((!g202) & (g719) & (!g759) & (g765) & (!g791) & (!g1052)) + ((!g202) & (g719) & (!g759) & (g765) & (g791) & (!g1052)) + ((!g202) & (g719) & (g759) & (!g765) & (!g791) & (!g1052)) + ((!g202) & (g719) & (g759) & (g765) & (!g791) & (!g1052)) + ((g202) & (!g719) & (!g759) & (!g765) & (!g791) & (g1052)) + ((g202) & (!g719) & (!g759) & (!g765) & (g791) & (g1052)) + ((g202) & (!g719) & (!g759) & (g765) & (!g791) & (!g1052)) + ((g202) & (!g719) & (!g759) & (g765) & (!g791) & (g1052)) + ((g202) & (!g719) & (!g759) & (g765) & (g791) & (!g1052)) + ((g202) & (!g719) & (!g759) & (g765) & (g791) & (g1052)) + ((g202) & (!g719) & (g759) & (!g765) & (!g791) & (g1052)) + ((g202) & (!g719) & (g759) & (!g765) & (g791) & (!g1052)) + ((g202) & (!g719) & (g759) & (!g765) & (g791) & (g1052)) + ((g202) & (!g719) & (g759) & (g765) & (!g791) & (!g1052)) + ((g202) & (!g719) & (g759) & (g765) & (!g791) & (g1052)) + ((g202) & (!g719) & (g759) & (g765) & (g791) & (!g1052)) + ((g202) & (!g719) & (g759) & (g765) & (g791) & (g1052)) + ((g202) & (g719) & (!g759) & (!g765) & (!g791) & (g1052)) + ((g202) & (g719) & (!g759) & (!g765) & (g791) & (g1052)) + ((g202) & (g719) & (!g759) & (g765) & (!g791) & (g1052)) + ((g202) & (g719) & (!g759) & (g765) & (g791) & (g1052)) + ((g202) & (g719) & (g759) & (!g765) & (!g791) & (g1052)) + ((g202) & (g719) & (g759) & (!g765) & (g791) & (!g1052)) + ((g202) & (g719) & (g759) & (!g765) & (g791) & (g1052)) + ((g202) & (g719) & (g759) & (g765) & (!g791) & (g1052)) + ((g202) & (g719) & (g759) & (g765) & (g791) & (!g1052)) + ((g202) & (g719) & (g759) & (g765) & (g791) & (g1052)));
	assign g1054 = (((!g1048) & (!g1051) & (sk[40]) & (g1053)) + ((!g1048) & (g1051) & (!sk[40]) & (!g1053)) + ((!g1048) & (g1051) & (!sk[40]) & (g1053)) + ((!g1048) & (g1051) & (sk[40]) & (!g1053)) + ((g1048) & (!g1051) & (sk[40]) & (!g1053)) + ((g1048) & (g1051) & (!sk[40]) & (!g1053)) + ((g1048) & (g1051) & (!sk[40]) & (g1053)) + ((g1048) & (g1051) & (sk[40]) & (g1053)));
	assign g1055 = (((!g979) & (!g981) & (!g982) & (!g988) & (!g1047) & (!g1054)) + ((!g979) & (!g981) & (!g982) & (!g988) & (g1047) & (g1054)) + ((!g979) & (!g981) & (!g982) & (g988) & (!g1047) & (g1054)) + ((!g979) & (!g981) & (!g982) & (g988) & (g1047) & (!g1054)) + ((!g979) & (!g981) & (g982) & (!g988) & (!g1047) & (g1054)) + ((!g979) & (!g981) & (g982) & (!g988) & (g1047) & (!g1054)) + ((!g979) & (!g981) & (g982) & (g988) & (!g1047) & (!g1054)) + ((!g979) & (!g981) & (g982) & (g988) & (g1047) & (g1054)) + ((!g979) & (g981) & (!g982) & (!g988) & (!g1047) & (g1054)) + ((!g979) & (g981) & (!g982) & (!g988) & (g1047) & (!g1054)) + ((!g979) & (g981) & (!g982) & (g988) & (!g1047) & (g1054)) + ((!g979) & (g981) & (!g982) & (g988) & (g1047) & (!g1054)) + ((!g979) & (g981) & (g982) & (!g988) & (!g1047) & (g1054)) + ((!g979) & (g981) & (g982) & (!g988) & (g1047) & (!g1054)) + ((!g979) & (g981) & (g982) & (g988) & (!g1047) & (g1054)) + ((!g979) & (g981) & (g982) & (g988) & (g1047) & (!g1054)) + ((g979) & (!g981) & (!g982) & (!g988) & (!g1047) & (!g1054)) + ((g979) & (!g981) & (!g982) & (!g988) & (g1047) & (g1054)) + ((g979) & (!g981) & (!g982) & (g988) & (!g1047) & (!g1054)) + ((g979) & (!g981) & (!g982) & (g988) & (g1047) & (g1054)) + ((g979) & (!g981) & (g982) & (!g988) & (!g1047) & (!g1054)) + ((g979) & (!g981) & (g982) & (!g988) & (g1047) & (g1054)) + ((g979) & (!g981) & (g982) & (g988) & (!g1047) & (!g1054)) + ((g979) & (!g981) & (g982) & (g988) & (g1047) & (g1054)) + ((g979) & (g981) & (!g982) & (!g988) & (!g1047) & (!g1054)) + ((g979) & (g981) & (!g982) & (!g988) & (g1047) & (g1054)) + ((g979) & (g981) & (!g982) & (g988) & (!g1047) & (g1054)) + ((g979) & (g981) & (!g982) & (g988) & (g1047) & (!g1054)) + ((g979) & (g981) & (g982) & (!g988) & (!g1047) & (g1054)) + ((g979) & (g981) & (g982) & (!g988) & (g1047) & (!g1054)) + ((g979) & (g981) & (g982) & (g988) & (!g1047) & (!g1054)) + ((g979) & (g981) & (g982) & (g988) & (g1047) & (g1054)));
	assign g1056 = (((g686) & (!sk[42]) & (g863)) + ((g686) & (sk[42]) & (g863)));
	assign g1057 = (((!g733) & (!g734) & (!g889) & (!sk[43]) & (g871) & (!g883)) + ((!g733) & (!g734) & (!g889) & (!sk[43]) & (g871) & (g883)) + ((!g733) & (!g734) & (g889) & (!sk[43]) & (!g871) & (!g883)) + ((!g733) & (!g734) & (g889) & (!sk[43]) & (!g871) & (g883)) + ((!g733) & (!g734) & (g889) & (!sk[43]) & (g871) & (!g883)) + ((!g733) & (!g734) & (g889) & (!sk[43]) & (g871) & (g883)) + ((!g733) & (g734) & (!g889) & (!sk[43]) & (!g871) & (!g883)) + ((!g733) & (g734) & (!g889) & (!sk[43]) & (!g871) & (g883)) + ((!g733) & (g734) & (!g889) & (!sk[43]) & (g871) & (!g883)) + ((!g733) & (g734) & (!g889) & (!sk[43]) & (g871) & (g883)) + ((!g733) & (g734) & (!g889) & (sk[43]) & (!g871) & (!g883)) + ((!g733) & (g734) & (!g889) & (sk[43]) & (g871) & (g883)) + ((!g733) & (g734) & (g889) & (!sk[43]) & (!g871) & (!g883)) + ((!g733) & (g734) & (g889) & (!sk[43]) & (!g871) & (g883)) + ((!g733) & (g734) & (g889) & (!sk[43]) & (g871) & (!g883)) + ((!g733) & (g734) & (g889) & (!sk[43]) & (g871) & (g883)) + ((!g733) & (g734) & (g889) & (sk[43]) & (!g871) & (!g883)) + ((!g733) & (g734) & (g889) & (sk[43]) & (g871) & (g883)) + ((g733) & (!g734) & (!g889) & (!sk[43]) & (g871) & (!g883)) + ((g733) & (!g734) & (!g889) & (!sk[43]) & (g871) & (g883)) + ((g733) & (!g734) & (!g889) & (sk[43]) & (!g871) & (!g883)) + ((g733) & (!g734) & (!g889) & (sk[43]) & (!g871) & (g883)) + ((g733) & (!g734) & (!g889) & (sk[43]) & (g871) & (!g883)) + ((g733) & (!g734) & (g889) & (!sk[43]) & (!g871) & (!g883)) + ((g733) & (!g734) & (g889) & (!sk[43]) & (!g871) & (g883)) + ((g733) & (!g734) & (g889) & (!sk[43]) & (g871) & (!g883)) + ((g733) & (!g734) & (g889) & (!sk[43]) & (g871) & (g883)) + ((g733) & (!g734) & (g889) & (sk[43]) & (g871) & (g883)) + ((g733) & (g734) & (!g889) & (!sk[43]) & (!g871) & (!g883)) + ((g733) & (g734) & (!g889) & (!sk[43]) & (!g871) & (g883)) + ((g733) & (g734) & (!g889) & (!sk[43]) & (g871) & (!g883)) + ((g733) & (g734) & (!g889) & (!sk[43]) & (g871) & (g883)) + ((g733) & (g734) & (!g889) & (sk[43]) & (!g871) & (!g883)) + ((g733) & (g734) & (!g889) & (sk[43]) & (!g871) & (g883)) + ((g733) & (g734) & (!g889) & (sk[43]) & (g871) & (!g883)) + ((g733) & (g734) & (!g889) & (sk[43]) & (g871) & (g883)) + ((g733) & (g734) & (g889) & (!sk[43]) & (!g871) & (!g883)) + ((g733) & (g734) & (g889) & (!sk[43]) & (!g871) & (g883)) + ((g733) & (g734) & (g889) & (!sk[43]) & (g871) & (!g883)) + ((g733) & (g734) & (g889) & (!sk[43]) & (g871) & (g883)) + ((g733) & (g734) & (g889) & (sk[43]) & (!g871) & (!g883)) + ((g733) & (g734) & (g889) & (sk[43]) & (g871) & (g883)));
	assign g1058 = (((!g2) & (!g732) & (!g884) & (!g890) & (!g1056) & (!g1057)) + ((!g2) & (!g732) & (!g884) & (g890) & (!g1056) & (!g1057)) + ((!g2) & (!g732) & (g884) & (!g890) & (!g1056) & (!g1057)) + ((!g2) & (!g732) & (g884) & (g890) & (!g1056) & (!g1057)) + ((!g2) & (g732) & (!g884) & (g890) & (!g1056) & (!g1057)) + ((!g2) & (g732) & (g884) & (!g890) & (!g1056) & (!g1057)) + ((g2) & (!g732) & (!g884) & (!g890) & (!g1056) & (g1057)) + ((g2) & (!g732) & (!g884) & (!g890) & (g1056) & (!g1057)) + ((g2) & (!g732) & (!g884) & (!g890) & (g1056) & (g1057)) + ((g2) & (!g732) & (!g884) & (g890) & (!g1056) & (g1057)) + ((g2) & (!g732) & (!g884) & (g890) & (g1056) & (!g1057)) + ((g2) & (!g732) & (!g884) & (g890) & (g1056) & (g1057)) + ((g2) & (!g732) & (g884) & (!g890) & (!g1056) & (g1057)) + ((g2) & (!g732) & (g884) & (!g890) & (g1056) & (!g1057)) + ((g2) & (!g732) & (g884) & (!g890) & (g1056) & (g1057)) + ((g2) & (!g732) & (g884) & (g890) & (!g1056) & (g1057)) + ((g2) & (!g732) & (g884) & (g890) & (g1056) & (!g1057)) + ((g2) & (!g732) & (g884) & (g890) & (g1056) & (g1057)) + ((g2) & (g732) & (!g884) & (!g890) & (!g1056) & (!g1057)) + ((g2) & (g732) & (!g884) & (!g890) & (!g1056) & (g1057)) + ((g2) & (g732) & (!g884) & (!g890) & (g1056) & (!g1057)) + ((g2) & (g732) & (!g884) & (!g890) & (g1056) & (g1057)) + ((g2) & (g732) & (!g884) & (g890) & (!g1056) & (g1057)) + ((g2) & (g732) & (!g884) & (g890) & (g1056) & (!g1057)) + ((g2) & (g732) & (!g884) & (g890) & (g1056) & (g1057)) + ((g2) & (g732) & (g884) & (!g890) & (!g1056) & (g1057)) + ((g2) & (g732) & (g884) & (!g890) & (g1056) & (!g1057)) + ((g2) & (g732) & (g884) & (!g890) & (g1056) & (g1057)) + ((g2) & (g732) & (g884) & (g890) & (!g1056) & (!g1057)) + ((g2) & (g732) & (g884) & (g890) & (!g1056) & (g1057)) + ((g2) & (g732) & (g884) & (g890) & (g1056) & (!g1057)) + ((g2) & (g732) & (g884) & (g890) & (g1056) & (g1057)));
	assign g1059 = (((!g1044) & (!sk[45]) & (g1055) & (!g1058)) + ((!g1044) & (!sk[45]) & (g1055) & (g1058)) + ((!g1044) & (sk[45]) & (!g1055) & (g1058)) + ((!g1044) & (sk[45]) & (g1055) & (!g1058)) + ((g1044) & (!sk[45]) & (g1055) & (!g1058)) + ((g1044) & (!sk[45]) & (g1055) & (g1058)) + ((g1044) & (sk[45]) & (!g1055) & (!g1058)) + ((g1044) & (sk[45]) & (g1055) & (g1058)));
	assign g1060 = (((!g975) & (!sk[46]) & (!g990) & (!g997) & (g1043) & (!g1059)) + ((!g975) & (!sk[46]) & (!g990) & (!g997) & (g1043) & (g1059)) + ((!g975) & (!sk[46]) & (!g990) & (g997) & (!g1043) & (!g1059)) + ((!g975) & (!sk[46]) & (!g990) & (g997) & (!g1043) & (g1059)) + ((!g975) & (!sk[46]) & (!g990) & (g997) & (g1043) & (!g1059)) + ((!g975) & (!sk[46]) & (!g990) & (g997) & (g1043) & (g1059)) + ((!g975) & (!sk[46]) & (g990) & (!g997) & (!g1043) & (!g1059)) + ((!g975) & (!sk[46]) & (g990) & (!g997) & (!g1043) & (g1059)) + ((!g975) & (!sk[46]) & (g990) & (!g997) & (g1043) & (!g1059)) + ((!g975) & (!sk[46]) & (g990) & (!g997) & (g1043) & (g1059)) + ((!g975) & (!sk[46]) & (g990) & (g997) & (!g1043) & (!g1059)) + ((!g975) & (!sk[46]) & (g990) & (g997) & (!g1043) & (g1059)) + ((!g975) & (!sk[46]) & (g990) & (g997) & (g1043) & (!g1059)) + ((!g975) & (!sk[46]) & (g990) & (g997) & (g1043) & (g1059)) + ((!g975) & (sk[46]) & (!g990) & (!g997) & (!g1043) & (g1059)) + ((!g975) & (sk[46]) & (!g990) & (!g997) & (g1043) & (!g1059)) + ((!g975) & (sk[46]) & (!g990) & (g997) & (!g1043) & (g1059)) + ((!g975) & (sk[46]) & (!g990) & (g997) & (g1043) & (!g1059)) + ((!g975) & (sk[46]) & (g990) & (!g997) & (!g1043) & (!g1059)) + ((!g975) & (sk[46]) & (g990) & (!g997) & (g1043) & (g1059)) + ((!g975) & (sk[46]) & (g990) & (g997) & (!g1043) & (g1059)) + ((!g975) & (sk[46]) & (g990) & (g997) & (g1043) & (!g1059)) + ((g975) & (!sk[46]) & (!g990) & (!g997) & (g1043) & (!g1059)) + ((g975) & (!sk[46]) & (!g990) & (!g997) & (g1043) & (g1059)) + ((g975) & (!sk[46]) & (!g990) & (g997) & (!g1043) & (!g1059)) + ((g975) & (!sk[46]) & (!g990) & (g997) & (!g1043) & (g1059)) + ((g975) & (!sk[46]) & (!g990) & (g997) & (g1043) & (!g1059)) + ((g975) & (!sk[46]) & (!g990) & (g997) & (g1043) & (g1059)) + ((g975) & (!sk[46]) & (g990) & (!g997) & (!g1043) & (!g1059)) + ((g975) & (!sk[46]) & (g990) & (!g997) & (!g1043) & (g1059)) + ((g975) & (!sk[46]) & (g990) & (!g997) & (g1043) & (!g1059)) + ((g975) & (!sk[46]) & (g990) & (!g997) & (g1043) & (g1059)) + ((g975) & (!sk[46]) & (g990) & (g997) & (!g1043) & (!g1059)) + ((g975) & (!sk[46]) & (g990) & (g997) & (!g1043) & (g1059)) + ((g975) & (!sk[46]) & (g990) & (g997) & (g1043) & (!g1059)) + ((g975) & (!sk[46]) & (g990) & (g997) & (g1043) & (g1059)) + ((g975) & (sk[46]) & (!g990) & (!g997) & (!g1043) & (!g1059)) + ((g975) & (sk[46]) & (!g990) & (!g997) & (g1043) & (g1059)) + ((g975) & (sk[46]) & (!g990) & (g997) & (!g1043) & (g1059)) + ((g975) & (sk[46]) & (!g990) & (g997) & (g1043) & (!g1059)) + ((g975) & (sk[46]) & (g990) & (!g997) & (!g1043) & (!g1059)) + ((g975) & (sk[46]) & (g990) & (!g997) & (g1043) & (g1059)) + ((g975) & (sk[46]) & (g990) & (g997) & (!g1043) & (!g1059)) + ((g975) & (sk[46]) & (g990) & (g997) & (g1043) & (g1059)));
	assign g1061 = (((!g254) & (!g255) & (!g256) & (g258) & (!sk[47]) & (!g151)) + ((!g254) & (!g255) & (!g256) & (g258) & (!sk[47]) & (g151)) + ((!g254) & (!g255) & (g256) & (!g258) & (!sk[47]) & (!g151)) + ((!g254) & (!g255) & (g256) & (!g258) & (!sk[47]) & (g151)) + ((!g254) & (!g255) & (g256) & (g258) & (!sk[47]) & (!g151)) + ((!g254) & (!g255) & (g256) & (g258) & (!sk[47]) & (g151)) + ((!g254) & (g255) & (!g256) & (!g258) & (!sk[47]) & (!g151)) + ((!g254) & (g255) & (!g256) & (!g258) & (!sk[47]) & (g151)) + ((!g254) & (g255) & (!g256) & (g258) & (!sk[47]) & (!g151)) + ((!g254) & (g255) & (!g256) & (g258) & (!sk[47]) & (g151)) + ((!g254) & (g255) & (g256) & (!g258) & (!sk[47]) & (!g151)) + ((!g254) & (g255) & (g256) & (!g258) & (!sk[47]) & (g151)) + ((!g254) & (g255) & (g256) & (g258) & (!sk[47]) & (!g151)) + ((!g254) & (g255) & (g256) & (g258) & (!sk[47]) & (g151)) + ((!g254) & (g255) & (g256) & (g258) & (sk[47]) & (g151)) + ((g254) & (!g255) & (!g256) & (g258) & (!sk[47]) & (!g151)) + ((g254) & (!g255) & (!g256) & (g258) & (!sk[47]) & (g151)) + ((g254) & (!g255) & (g256) & (!g258) & (!sk[47]) & (!g151)) + ((g254) & (!g255) & (g256) & (!g258) & (!sk[47]) & (g151)) + ((g254) & (!g255) & (g256) & (g258) & (!sk[47]) & (!g151)) + ((g254) & (!g255) & (g256) & (g258) & (!sk[47]) & (g151)) + ((g254) & (g255) & (!g256) & (!g258) & (!sk[47]) & (!g151)) + ((g254) & (g255) & (!g256) & (!g258) & (!sk[47]) & (g151)) + ((g254) & (g255) & (!g256) & (g258) & (!sk[47]) & (!g151)) + ((g254) & (g255) & (!g256) & (g258) & (!sk[47]) & (g151)) + ((g254) & (g255) & (g256) & (!g258) & (!sk[47]) & (!g151)) + ((g254) & (g255) & (g256) & (!g258) & (!sk[47]) & (g151)) + ((g254) & (g255) & (g256) & (g258) & (!sk[47]) & (!g151)) + ((g254) & (g255) & (g256) & (g258) & (!sk[47]) & (g151)));
	assign g1062 = (((!g147) & (!g137) & (sk[48]) & (!g108)) + ((!g147) & (g137) & (!sk[48]) & (!g108)) + ((!g147) & (g137) & (!sk[48]) & (g108)) + ((g147) & (g137) & (!sk[48]) & (!g108)) + ((g147) & (g137) & (!sk[48]) & (g108)));
	assign g1063 = (((!g43) & (!sk[49]) & (!g233) & (!g160) & (g1062)) + ((!g43) & (!sk[49]) & (!g233) & (g160) & (g1062)) + ((!g43) & (!sk[49]) & (g233) & (!g160) & (g1062)) + ((!g43) & (!sk[49]) & (g233) & (g160) & (g1062)) + ((!g43) & (sk[49]) & (!g233) & (g160) & (g1062)) + ((g43) & (!sk[49]) & (!g233) & (!g160) & (!g1062)) + ((g43) & (!sk[49]) & (!g233) & (!g160) & (g1062)) + ((g43) & (!sk[49]) & (!g233) & (g160) & (!g1062)) + ((g43) & (!sk[49]) & (!g233) & (g160) & (g1062)) + ((g43) & (!sk[49]) & (g233) & (!g160) & (!g1062)) + ((g43) & (!sk[49]) & (g233) & (!g160) & (g1062)) + ((g43) & (!sk[49]) & (g233) & (g160) & (!g1062)) + ((g43) & (!sk[49]) & (g233) & (g160) & (g1062)));
	assign g1064 = (((!g879) & (!g31) & (!sk[50]) & (!g81) & (g1001)) + ((!g879) & (!g31) & (!sk[50]) & (g81) & (g1001)) + ((!g879) & (g31) & (!sk[50]) & (!g81) & (g1001)) + ((!g879) & (g31) & (!sk[50]) & (g81) & (g1001)) + ((g879) & (!g31) & (!sk[50]) & (!g81) & (!g1001)) + ((g879) & (!g31) & (!sk[50]) & (!g81) & (g1001)) + ((g879) & (!g31) & (!sk[50]) & (g81) & (!g1001)) + ((g879) & (!g31) & (!sk[50]) & (g81) & (g1001)) + ((g879) & (!g31) & (sk[50]) & (!g81) & (g1001)) + ((g879) & (g31) & (!sk[50]) & (!g81) & (!g1001)) + ((g879) & (g31) & (!sk[50]) & (!g81) & (g1001)) + ((g879) & (g31) & (!sk[50]) & (g81) & (!g1001)) + ((g879) & (g31) & (!sk[50]) & (g81) & (g1001)));
	assign g1065 = (((!sk[51]) & (!g1061) & (!g295) & (!g589) & (g1063) & (!g1064)) + ((!sk[51]) & (!g1061) & (!g295) & (!g589) & (g1063) & (g1064)) + ((!sk[51]) & (!g1061) & (!g295) & (g589) & (!g1063) & (!g1064)) + ((!sk[51]) & (!g1061) & (!g295) & (g589) & (!g1063) & (g1064)) + ((!sk[51]) & (!g1061) & (!g295) & (g589) & (g1063) & (!g1064)) + ((!sk[51]) & (!g1061) & (!g295) & (g589) & (g1063) & (g1064)) + ((!sk[51]) & (!g1061) & (g295) & (!g589) & (!g1063) & (!g1064)) + ((!sk[51]) & (!g1061) & (g295) & (!g589) & (!g1063) & (g1064)) + ((!sk[51]) & (!g1061) & (g295) & (!g589) & (g1063) & (!g1064)) + ((!sk[51]) & (!g1061) & (g295) & (!g589) & (g1063) & (g1064)) + ((!sk[51]) & (!g1061) & (g295) & (g589) & (!g1063) & (!g1064)) + ((!sk[51]) & (!g1061) & (g295) & (g589) & (!g1063) & (g1064)) + ((!sk[51]) & (!g1061) & (g295) & (g589) & (g1063) & (!g1064)) + ((!sk[51]) & (!g1061) & (g295) & (g589) & (g1063) & (g1064)) + ((!sk[51]) & (g1061) & (!g295) & (!g589) & (g1063) & (!g1064)) + ((!sk[51]) & (g1061) & (!g295) & (!g589) & (g1063) & (g1064)) + ((!sk[51]) & (g1061) & (!g295) & (g589) & (!g1063) & (!g1064)) + ((!sk[51]) & (g1061) & (!g295) & (g589) & (!g1063) & (g1064)) + ((!sk[51]) & (g1061) & (!g295) & (g589) & (g1063) & (!g1064)) + ((!sk[51]) & (g1061) & (!g295) & (g589) & (g1063) & (g1064)) + ((!sk[51]) & (g1061) & (g295) & (!g589) & (!g1063) & (!g1064)) + ((!sk[51]) & (g1061) & (g295) & (!g589) & (!g1063) & (g1064)) + ((!sk[51]) & (g1061) & (g295) & (!g589) & (g1063) & (!g1064)) + ((!sk[51]) & (g1061) & (g295) & (!g589) & (g1063) & (g1064)) + ((!sk[51]) & (g1061) & (g295) & (g589) & (!g1063) & (!g1064)) + ((!sk[51]) & (g1061) & (g295) & (g589) & (!g1063) & (g1064)) + ((!sk[51]) & (g1061) & (g295) & (g589) & (g1063) & (!g1064)) + ((!sk[51]) & (g1061) & (g295) & (g589) & (g1063) & (g1064)) + ((sk[51]) & (g1061) & (g295) & (g589) & (g1063) & (g1064)));
	assign g1066 = (((!g975) & (!sk[52]) & (!g998) & (!g1010) & (g1030)) + ((!g975) & (!sk[52]) & (!g998) & (g1010) & (g1030)) + ((!g975) & (!sk[52]) & (g998) & (!g1010) & (g1030)) + ((!g975) & (!sk[52]) & (g998) & (g1010) & (g1030)) + ((!g975) & (sk[52]) & (!g998) & (!g1010) & (!g1030)) + ((!g975) & (sk[52]) & (!g998) & (g1010) & (g1030)) + ((!g975) & (sk[52]) & (g998) & (!g1010) & (g1030)) + ((!g975) & (sk[52]) & (g998) & (g1010) & (!g1030)) + ((g975) & (!sk[52]) & (!g998) & (!g1010) & (!g1030)) + ((g975) & (!sk[52]) & (!g998) & (!g1010) & (g1030)) + ((g975) & (!sk[52]) & (!g998) & (g1010) & (!g1030)) + ((g975) & (!sk[52]) & (!g998) & (g1010) & (g1030)) + ((g975) & (!sk[52]) & (g998) & (!g1010) & (!g1030)) + ((g975) & (!sk[52]) & (g998) & (!g1010) & (g1030)) + ((g975) & (!sk[52]) & (g998) & (g1010) & (!g1030)) + ((g975) & (!sk[52]) & (g998) & (g1010) & (g1030)) + ((g975) & (sk[52]) & (!g998) & (!g1010) & (g1030)) + ((g975) & (sk[52]) & (!g998) & (g1010) & (!g1030)) + ((g975) & (sk[52]) & (g998) & (!g1010) & (!g1030)) + ((g975) & (sk[52]) & (g998) & (g1010) & (g1030)));
	assign g1067 = (((!g1031) & (!g1060) & (!g1065) & (!sk[53]) & (g1066)) + ((!g1031) & (!g1060) & (!g1065) & (sk[53]) & (!g1066)) + ((!g1031) & (!g1060) & (g1065) & (!sk[53]) & (g1066)) + ((!g1031) & (!g1060) & (g1065) & (sk[53]) & (g1066)) + ((!g1031) & (g1060) & (!g1065) & (!sk[53]) & (g1066)) + ((!g1031) & (g1060) & (!g1065) & (sk[53]) & (g1066)) + ((!g1031) & (g1060) & (g1065) & (!sk[53]) & (g1066)) + ((!g1031) & (g1060) & (g1065) & (sk[53]) & (!g1066)) + ((g1031) & (!g1060) & (!g1065) & (!sk[53]) & (!g1066)) + ((g1031) & (!g1060) & (!g1065) & (!sk[53]) & (g1066)) + ((g1031) & (!g1060) & (!g1065) & (sk[53]) & (g1066)) + ((g1031) & (!g1060) & (g1065) & (!sk[53]) & (!g1066)) + ((g1031) & (!g1060) & (g1065) & (!sk[53]) & (g1066)) + ((g1031) & (!g1060) & (g1065) & (sk[53]) & (!g1066)) + ((g1031) & (g1060) & (!g1065) & (!sk[53]) & (!g1066)) + ((g1031) & (g1060) & (!g1065) & (!sk[53]) & (g1066)) + ((g1031) & (g1060) & (!g1065) & (sk[53]) & (!g1066)) + ((g1031) & (g1060) & (g1065) & (!sk[53]) & (!g1066)) + ((g1031) & (g1060) & (g1065) & (!sk[53]) & (g1066)) + ((g1031) & (g1060) & (g1065) & (sk[53]) & (g1066)));
	assign g1068 = (((!sk[54]) & (ax22x) & (ax23x)) + ((sk[54]) & (!ax22x) & (ax23x)) + ((sk[54]) & (ax22x) & (!ax23x)));
	assign g1069 = (((!g1031) & (!sk[55]) & (!g1060) & (!g1065) & (g1066)) + ((!g1031) & (!sk[55]) & (!g1060) & (g1065) & (g1066)) + ((!g1031) & (!sk[55]) & (g1060) & (!g1065) & (g1066)) + ((!g1031) & (!sk[55]) & (g1060) & (g1065) & (g1066)) + ((!g1031) & (sk[55]) & (!g1060) & (!g1065) & (!g1066)) + ((!g1031) & (sk[55]) & (g1060) & (g1065) & (!g1066)) + ((g1031) & (!sk[55]) & (!g1060) & (!g1065) & (!g1066)) + ((g1031) & (!sk[55]) & (!g1060) & (!g1065) & (g1066)) + ((g1031) & (!sk[55]) & (!g1060) & (g1065) & (!g1066)) + ((g1031) & (!sk[55]) & (!g1060) & (g1065) & (g1066)) + ((g1031) & (!sk[55]) & (g1060) & (!g1065) & (!g1066)) + ((g1031) & (!sk[55]) & (g1060) & (!g1065) & (g1066)) + ((g1031) & (!sk[55]) & (g1060) & (g1065) & (!g1066)) + ((g1031) & (!sk[55]) & (g1060) & (g1065) & (g1066)) + ((g1031) & (sk[55]) & (!g1060) & (g1065) & (!g1066)) + ((g1031) & (sk[55]) & (g1060) & (!g1065) & (!g1066)));
	assign g1070 = (((!sk[56]) & (!g275) & (!g352) & (!g970) & (g993) & (!g1037)) + ((!sk[56]) & (!g275) & (!g352) & (!g970) & (g993) & (g1037)) + ((!sk[56]) & (!g275) & (!g352) & (g970) & (!g993) & (!g1037)) + ((!sk[56]) & (!g275) & (!g352) & (g970) & (!g993) & (g1037)) + ((!sk[56]) & (!g275) & (!g352) & (g970) & (g993) & (!g1037)) + ((!sk[56]) & (!g275) & (!g352) & (g970) & (g993) & (g1037)) + ((!sk[56]) & (!g275) & (g352) & (!g970) & (!g993) & (!g1037)) + ((!sk[56]) & (!g275) & (g352) & (!g970) & (!g993) & (g1037)) + ((!sk[56]) & (!g275) & (g352) & (!g970) & (g993) & (!g1037)) + ((!sk[56]) & (!g275) & (g352) & (!g970) & (g993) & (g1037)) + ((!sk[56]) & (!g275) & (g352) & (g970) & (!g993) & (!g1037)) + ((!sk[56]) & (!g275) & (g352) & (g970) & (!g993) & (g1037)) + ((!sk[56]) & (!g275) & (g352) & (g970) & (g993) & (!g1037)) + ((!sk[56]) & (!g275) & (g352) & (g970) & (g993) & (g1037)) + ((!sk[56]) & (g275) & (!g352) & (!g970) & (g993) & (!g1037)) + ((!sk[56]) & (g275) & (!g352) & (!g970) & (g993) & (g1037)) + ((!sk[56]) & (g275) & (!g352) & (g970) & (!g993) & (!g1037)) + ((!sk[56]) & (g275) & (!g352) & (g970) & (!g993) & (g1037)) + ((!sk[56]) & (g275) & (!g352) & (g970) & (g993) & (!g1037)) + ((!sk[56]) & (g275) & (!g352) & (g970) & (g993) & (g1037)) + ((!sk[56]) & (g275) & (g352) & (!g970) & (!g993) & (!g1037)) + ((!sk[56]) & (g275) & (g352) & (!g970) & (!g993) & (g1037)) + ((!sk[56]) & (g275) & (g352) & (!g970) & (g993) & (!g1037)) + ((!sk[56]) & (g275) & (g352) & (!g970) & (g993) & (g1037)) + ((!sk[56]) & (g275) & (g352) & (g970) & (!g993) & (!g1037)) + ((!sk[56]) & (g275) & (g352) & (g970) & (!g993) & (g1037)) + ((!sk[56]) & (g275) & (g352) & (g970) & (g993) & (!g1037)) + ((!sk[56]) & (g275) & (g352) & (g970) & (g993) & (g1037)) + ((sk[56]) & (!g275) & (g352) & (g970) & (g993) & (g1037)));
	assign g1071 = (((!g146) & (!g152) & (sk[57]) & (!g170)) + ((!g146) & (g152) & (!sk[57]) & (!g170)) + ((!g146) & (g152) & (!sk[57]) & (g170)) + ((g146) & (g152) & (!sk[57]) & (!g170)) + ((g146) & (g152) & (!sk[57]) & (g170)));
	assign g1072 = (((!g354) & (!g601) & (!g236) & (!sk[58]) & (g177)) + ((!g354) & (!g601) & (!g236) & (sk[58]) & (!g177)) + ((!g354) & (!g601) & (g236) & (!sk[58]) & (g177)) + ((!g354) & (g601) & (!g236) & (!sk[58]) & (g177)) + ((!g354) & (g601) & (g236) & (!sk[58]) & (g177)) + ((g354) & (!g601) & (!g236) & (!sk[58]) & (!g177)) + ((g354) & (!g601) & (!g236) & (!sk[58]) & (g177)) + ((g354) & (!g601) & (g236) & (!sk[58]) & (!g177)) + ((g354) & (!g601) & (g236) & (!sk[58]) & (g177)) + ((g354) & (g601) & (!g236) & (!sk[58]) & (!g177)) + ((g354) & (g601) & (!g236) & (!sk[58]) & (g177)) + ((g354) & (g601) & (g236) & (!sk[58]) & (!g177)) + ((g354) & (g601) & (g236) & (!sk[58]) & (g177)));
	assign g1073 = (((!g76) & (!g238) & (!g193) & (!sk[59]) & (g95)) + ((!g76) & (!g238) & (!g193) & (sk[59]) & (!g95)) + ((!g76) & (!g238) & (g193) & (!sk[59]) & (g95)) + ((!g76) & (g238) & (!g193) & (!sk[59]) & (g95)) + ((!g76) & (g238) & (g193) & (!sk[59]) & (g95)) + ((g76) & (!g238) & (!g193) & (!sk[59]) & (!g95)) + ((g76) & (!g238) & (!g193) & (!sk[59]) & (g95)) + ((g76) & (!g238) & (g193) & (!sk[59]) & (!g95)) + ((g76) & (!g238) & (g193) & (!sk[59]) & (g95)) + ((g76) & (g238) & (!g193) & (!sk[59]) & (!g95)) + ((g76) & (g238) & (!g193) & (!sk[59]) & (g95)) + ((g76) & (g238) & (g193) & (!sk[59]) & (!g95)) + ((g76) & (g238) & (g193) & (!sk[59]) & (g95)));
	assign g1074 = (((!sk[60]) & (!g17) & (!g71) & (!g127) & (g27)) + ((!sk[60]) & (!g17) & (!g71) & (g127) & (g27)) + ((!sk[60]) & (!g17) & (g71) & (!g127) & (g27)) + ((!sk[60]) & (!g17) & (g71) & (g127) & (g27)) + ((!sk[60]) & (g17) & (!g71) & (!g127) & (!g27)) + ((!sk[60]) & (g17) & (!g71) & (!g127) & (g27)) + ((!sk[60]) & (g17) & (!g71) & (g127) & (!g27)) + ((!sk[60]) & (g17) & (!g71) & (g127) & (g27)) + ((!sk[60]) & (g17) & (g71) & (!g127) & (!g27)) + ((!sk[60]) & (g17) & (g71) & (!g127) & (g27)) + ((!sk[60]) & (g17) & (g71) & (g127) & (!g27)) + ((!sk[60]) & (g17) & (g71) & (g127) & (g27)) + ((sk[60]) & (!g17) & (!g71) & (!g127) & (!g27)) + ((sk[60]) & (!g17) & (!g71) & (!g127) & (g27)) + ((sk[60]) & (!g17) & (g71) & (!g127) & (!g27)) + ((sk[60]) & (g17) & (!g71) & (!g127) & (!g27)) + ((sk[60]) & (g17) & (!g71) & (!g127) & (g27)));
	assign g1075 = (((!g58) & (!g104) & (!g187) & (!sk[61]) & (g1074)) + ((!g58) & (!g104) & (!g187) & (sk[61]) & (g1074)) + ((!g58) & (!g104) & (g187) & (!sk[61]) & (g1074)) + ((!g58) & (g104) & (!g187) & (!sk[61]) & (g1074)) + ((!g58) & (g104) & (!g187) & (sk[61]) & (g1074)) + ((!g58) & (g104) & (g187) & (!sk[61]) & (g1074)) + ((g58) & (!g104) & (!g187) & (!sk[61]) & (!g1074)) + ((g58) & (!g104) & (!g187) & (!sk[61]) & (g1074)) + ((g58) & (!g104) & (!g187) & (sk[61]) & (g1074)) + ((g58) & (!g104) & (g187) & (!sk[61]) & (!g1074)) + ((g58) & (!g104) & (g187) & (!sk[61]) & (g1074)) + ((g58) & (g104) & (!g187) & (!sk[61]) & (!g1074)) + ((g58) & (g104) & (!g187) & (!sk[61]) & (g1074)) + ((g58) & (g104) & (g187) & (!sk[61]) & (!g1074)) + ((g58) & (g104) & (g187) & (!sk[61]) & (g1074)));
	assign g1076 = (((!sk[62]) & (!g72) & (!g205) & (!g1073) & (g1075)) + ((!sk[62]) & (!g72) & (!g205) & (g1073) & (g1075)) + ((!sk[62]) & (!g72) & (g205) & (!g1073) & (g1075)) + ((!sk[62]) & (!g72) & (g205) & (g1073) & (g1075)) + ((!sk[62]) & (g72) & (!g205) & (!g1073) & (!g1075)) + ((!sk[62]) & (g72) & (!g205) & (!g1073) & (g1075)) + ((!sk[62]) & (g72) & (!g205) & (g1073) & (!g1075)) + ((!sk[62]) & (g72) & (!g205) & (g1073) & (g1075)) + ((!sk[62]) & (g72) & (g205) & (!g1073) & (!g1075)) + ((!sk[62]) & (g72) & (g205) & (!g1073) & (g1075)) + ((!sk[62]) & (g72) & (g205) & (g1073) & (!g1075)) + ((!sk[62]) & (g72) & (g205) & (g1073) & (g1075)) + ((sk[62]) & (!g72) & (!g205) & (g1073) & (g1075)));
	assign g1077 = (((!g270) & (g271) & (!sk[63]) & (!g1076)) + ((!g270) & (g271) & (!sk[63]) & (g1076)) + ((g270) & (!g271) & (sk[63]) & (g1076)) + ((g270) & (g271) & (!sk[63]) & (!g1076)) + ((g270) & (g271) & (!sk[63]) & (g1076)));
	assign g1078 = (((!g417) & (!g648) & (!g1071) & (!sk[64]) & (g1072) & (!g1077)) + ((!g417) & (!g648) & (!g1071) & (!sk[64]) & (g1072) & (g1077)) + ((!g417) & (!g648) & (g1071) & (!sk[64]) & (!g1072) & (!g1077)) + ((!g417) & (!g648) & (g1071) & (!sk[64]) & (!g1072) & (g1077)) + ((!g417) & (!g648) & (g1071) & (!sk[64]) & (g1072) & (!g1077)) + ((!g417) & (!g648) & (g1071) & (!sk[64]) & (g1072) & (g1077)) + ((!g417) & (g648) & (!g1071) & (!sk[64]) & (!g1072) & (!g1077)) + ((!g417) & (g648) & (!g1071) & (!sk[64]) & (!g1072) & (g1077)) + ((!g417) & (g648) & (!g1071) & (!sk[64]) & (g1072) & (!g1077)) + ((!g417) & (g648) & (!g1071) & (!sk[64]) & (g1072) & (g1077)) + ((!g417) & (g648) & (g1071) & (!sk[64]) & (!g1072) & (!g1077)) + ((!g417) & (g648) & (g1071) & (!sk[64]) & (!g1072) & (g1077)) + ((!g417) & (g648) & (g1071) & (!sk[64]) & (g1072) & (!g1077)) + ((!g417) & (g648) & (g1071) & (!sk[64]) & (g1072) & (g1077)) + ((g417) & (!g648) & (!g1071) & (!sk[64]) & (g1072) & (!g1077)) + ((g417) & (!g648) & (!g1071) & (!sk[64]) & (g1072) & (g1077)) + ((g417) & (!g648) & (g1071) & (!sk[64]) & (!g1072) & (!g1077)) + ((g417) & (!g648) & (g1071) & (!sk[64]) & (!g1072) & (g1077)) + ((g417) & (!g648) & (g1071) & (!sk[64]) & (g1072) & (!g1077)) + ((g417) & (!g648) & (g1071) & (!sk[64]) & (g1072) & (g1077)) + ((g417) & (g648) & (!g1071) & (!sk[64]) & (!g1072) & (!g1077)) + ((g417) & (g648) & (!g1071) & (!sk[64]) & (!g1072) & (g1077)) + ((g417) & (g648) & (!g1071) & (!sk[64]) & (g1072) & (!g1077)) + ((g417) & (g648) & (!g1071) & (!sk[64]) & (g1072) & (g1077)) + ((g417) & (g648) & (g1071) & (!sk[64]) & (!g1072) & (!g1077)) + ((g417) & (g648) & (g1071) & (!sk[64]) & (!g1072) & (g1077)) + ((g417) & (g648) & (g1071) & (!sk[64]) & (g1072) & (!g1077)) + ((g417) & (g648) & (g1071) & (!sk[64]) & (g1072) & (g1077)) + ((g417) & (g648) & (g1071) & (sk[64]) & (g1072) & (g1077)));
	assign g1079 = (((!g888) & (!g871) & (!g883) & (!sk[65]) & (g1070) & (!g1078)) + ((!g888) & (!g871) & (!g883) & (!sk[65]) & (g1070) & (g1078)) + ((!g888) & (!g871) & (!g883) & (sk[65]) & (!g1070) & (g1078)) + ((!g888) & (!g871) & (!g883) & (sk[65]) & (g1070) & (g1078)) + ((!g888) & (!g871) & (g883) & (!sk[65]) & (!g1070) & (!g1078)) + ((!g888) & (!g871) & (g883) & (!sk[65]) & (!g1070) & (g1078)) + ((!g888) & (!g871) & (g883) & (!sk[65]) & (g1070) & (!g1078)) + ((!g888) & (!g871) & (g883) & (!sk[65]) & (g1070) & (g1078)) + ((!g888) & (!g871) & (g883) & (sk[65]) & (!g1070) & (g1078)) + ((!g888) & (!g871) & (g883) & (sk[65]) & (g1070) & (g1078)) + ((!g888) & (g871) & (!g883) & (!sk[65]) & (!g1070) & (!g1078)) + ((!g888) & (g871) & (!g883) & (!sk[65]) & (!g1070) & (g1078)) + ((!g888) & (g871) & (!g883) & (!sk[65]) & (g1070) & (!g1078)) + ((!g888) & (g871) & (!g883) & (!sk[65]) & (g1070) & (g1078)) + ((!g888) & (g871) & (!g883) & (sk[65]) & (!g1070) & (g1078)) + ((!g888) & (g871) & (!g883) & (sk[65]) & (g1070) & (g1078)) + ((!g888) & (g871) & (g883) & (!sk[65]) & (!g1070) & (!g1078)) + ((!g888) & (g871) & (g883) & (!sk[65]) & (!g1070) & (g1078)) + ((!g888) & (g871) & (g883) & (!sk[65]) & (g1070) & (!g1078)) + ((!g888) & (g871) & (g883) & (!sk[65]) & (g1070) & (g1078)) + ((!g888) & (g871) & (g883) & (sk[65]) & (!g1070) & (g1078)) + ((!g888) & (g871) & (g883) & (sk[65]) & (g1070) & (g1078)) + ((g888) & (!g871) & (!g883) & (!sk[65]) & (g1070) & (!g1078)) + ((g888) & (!g871) & (!g883) & (!sk[65]) & (g1070) & (g1078)) + ((g888) & (!g871) & (!g883) & (sk[65]) & (!g1070) & (g1078)) + ((g888) & (!g871) & (!g883) & (sk[65]) & (g1070) & (g1078)) + ((g888) & (!g871) & (g883) & (!sk[65]) & (!g1070) & (!g1078)) + ((g888) & (!g871) & (g883) & (!sk[65]) & (!g1070) & (g1078)) + ((g888) & (!g871) & (g883) & (!sk[65]) & (g1070) & (!g1078)) + ((g888) & (!g871) & (g883) & (!sk[65]) & (g1070) & (g1078)) + ((g888) & (!g871) & (g883) & (sk[65]) & (!g1070) & (g1078)) + ((g888) & (!g871) & (g883) & (sk[65]) & (g1070) & (g1078)) + ((g888) & (g871) & (!g883) & (!sk[65]) & (!g1070) & (!g1078)) + ((g888) & (g871) & (!g883) & (!sk[65]) & (!g1070) & (g1078)) + ((g888) & (g871) & (!g883) & (!sk[65]) & (g1070) & (!g1078)) + ((g888) & (g871) & (!g883) & (!sk[65]) & (g1070) & (g1078)) + ((g888) & (g871) & (!g883) & (sk[65]) & (!g1070) & (g1078)) + ((g888) & (g871) & (!g883) & (sk[65]) & (g1070) & (g1078)) + ((g888) & (g871) & (g883) & (!sk[65]) & (!g1070) & (!g1078)) + ((g888) & (g871) & (g883) & (!sk[65]) & (!g1070) & (g1078)) + ((g888) & (g871) & (g883) & (!sk[65]) & (g1070) & (!g1078)) + ((g888) & (g871) & (g883) & (!sk[65]) & (g1070) & (g1078)) + ((g888) & (g871) & (g883) & (sk[65]) & (!g1070) & (g1078)) + ((g888) & (g871) & (g883) & (sk[65]) & (g1070) & (!g1078)));
	assign g1080 = (((!g962) & (!g963) & (!g884) & (!g971) & (g994) & (!g1040)) + ((!g962) & (!g963) & (!g884) & (g971) & (!g994) & (!g1040)) + ((!g962) & (!g963) & (!g884) & (g971) & (g994) & (!g1040)) + ((!g962) & (!g963) & (!g884) & (g971) & (g994) & (g1040)) + ((!g962) & (!g963) & (g884) & (!g971) & (g994) & (!g1040)) + ((!g962) & (!g963) & (g884) & (!g971) & (g994) & (g1040)) + ((!g962) & (!g963) & (g884) & (g971) & (!g994) & (!g1040)) + ((!g962) & (!g963) & (g884) & (g971) & (g994) & (!g1040)) + ((!g962) & (!g963) & (g884) & (g971) & (g994) & (g1040)) + ((!g962) & (g963) & (!g884) & (!g971) & (g994) & (!g1040)) + ((!g962) & (g963) & (!g884) & (!g971) & (g994) & (g1040)) + ((!g962) & (g963) & (!g884) & (g971) & (!g994) & (!g1040)) + ((!g962) & (g963) & (!g884) & (g971) & (g994) & (!g1040)) + ((!g962) & (g963) & (!g884) & (g971) & (g994) & (g1040)) + ((!g962) & (g963) & (g884) & (!g971) & (g994) & (!g1040)) + ((!g962) & (g963) & (g884) & (!g971) & (g994) & (g1040)) + ((!g962) & (g963) & (g884) & (g971) & (!g994) & (!g1040)) + ((!g962) & (g963) & (g884) & (g971) & (g994) & (!g1040)) + ((!g962) & (g963) & (g884) & (g971) & (g994) & (g1040)) + ((g962) & (!g963) & (!g884) & (!g971) & (g994) & (!g1040)) + ((g962) & (!g963) & (!g884) & (g971) & (g994) & (!g1040)) + ((g962) & (!g963) & (!g884) & (g971) & (g994) & (g1040)) + ((g962) & (!g963) & (g884) & (!g971) & (g994) & (!g1040)) + ((g962) & (!g963) & (g884) & (g971) & (g994) & (!g1040)) + ((g962) & (!g963) & (g884) & (g971) & (g994) & (g1040)) + ((g962) & (g963) & (!g884) & (!g971) & (g994) & (!g1040)) + ((g962) & (g963) & (!g884) & (g971) & (g994) & (!g1040)) + ((g962) & (g963) & (!g884) & (g971) & (g994) & (g1040)) + ((g962) & (g963) & (g884) & (!g971) & (g994) & (!g1040)) + ((g962) & (g963) & (g884) & (g971) & (!g994) & (!g1040)) + ((g962) & (g963) & (g884) & (g971) & (g994) & (!g1040)) + ((g962) & (g963) & (g884) & (g971) & (g994) & (g1040)));
	assign g1081 = (((!g891) & (!g864) & (!g892) & (!g994) & (!g1040) & (!g1079)) + ((!g891) & (!g864) & (!g892) & (!g994) & (!g1040) & (g1079)) + ((!g891) & (!g864) & (!g892) & (!g994) & (g1040) & (!g1079)) + ((!g891) & (!g864) & (!g892) & (!g994) & (g1040) & (g1079)) + ((!g891) & (!g864) & (!g892) & (g994) & (!g1040) & (!g1079)) + ((!g891) & (!g864) & (!g892) & (g994) & (!g1040) & (g1079)) + ((!g891) & (!g864) & (!g892) & (g994) & (g1040) & (!g1079)) + ((!g891) & (!g864) & (!g892) & (g994) & (g1040) & (g1079)) + ((!g891) & (!g864) & (g892) & (!g994) & (g1040) & (!g1079)) + ((!g891) & (!g864) & (g892) & (!g994) & (g1040) & (g1079)) + ((!g891) & (!g864) & (g892) & (g994) & (g1040) & (!g1079)) + ((!g891) & (!g864) & (g892) & (g994) & (g1040) & (g1079)) + ((!g891) & (g864) & (!g892) & (!g994) & (!g1040) & (!g1079)) + ((!g891) & (g864) & (!g892) & (!g994) & (!g1040) & (g1079)) + ((!g891) & (g864) & (!g892) & (!g994) & (g1040) & (!g1079)) + ((!g891) & (g864) & (!g892) & (!g994) & (g1040) & (g1079)) + ((!g891) & (g864) & (g892) & (!g994) & (g1040) & (!g1079)) + ((!g891) & (g864) & (g892) & (!g994) & (g1040) & (g1079)) + ((g891) & (!g864) & (!g892) & (!g994) & (!g1040) & (g1079)) + ((g891) & (!g864) & (!g892) & (!g994) & (g1040) & (g1079)) + ((g891) & (!g864) & (!g892) & (g994) & (!g1040) & (g1079)) + ((g891) & (!g864) & (!g892) & (g994) & (g1040) & (g1079)) + ((g891) & (!g864) & (g892) & (!g994) & (g1040) & (g1079)) + ((g891) & (!g864) & (g892) & (g994) & (g1040) & (g1079)) + ((g891) & (g864) & (!g892) & (!g994) & (!g1040) & (g1079)) + ((g891) & (g864) & (!g892) & (!g994) & (g1040) & (g1079)) + ((g891) & (g864) & (g892) & (!g994) & (g1040) & (g1079)));
	assign g1082 = (((!g683) & (!g868) & (!g1040) & (!g1079) & (!g1080) & (!g1081)) + ((!g683) & (!g868) & (!g1040) & (!g1079) & (g1080) & (!g1081)) + ((!g683) & (!g868) & (!g1040) & (g1079) & (!g1080) & (!g1081)) + ((!g683) & (!g868) & (!g1040) & (g1079) & (g1080) & (!g1081)) + ((!g683) & (!g868) & (g1040) & (!g1079) & (!g1080) & (!g1081)) + ((!g683) & (!g868) & (g1040) & (!g1079) & (g1080) & (!g1081)) + ((!g683) & (!g868) & (g1040) & (g1079) & (!g1080) & (!g1081)) + ((!g683) & (!g868) & (g1040) & (g1079) & (g1080) & (!g1081)) + ((!g683) & (g868) & (!g1040) & (!g1079) & (!g1080) & (!g1081)) + ((!g683) & (g868) & (!g1040) & (!g1079) & (g1080) & (!g1081)) + ((!g683) & (g868) & (!g1040) & (!g1079) & (g1080) & (g1081)) + ((!g683) & (g868) & (!g1040) & (g1079) & (!g1080) & (!g1081)) + ((!g683) & (g868) & (!g1040) & (g1079) & (!g1080) & (g1081)) + ((!g683) & (g868) & (!g1040) & (g1079) & (g1080) & (!g1081)) + ((!g683) & (g868) & (g1040) & (!g1079) & (!g1080) & (!g1081)) + ((!g683) & (g868) & (g1040) & (!g1079) & (!g1080) & (g1081)) + ((!g683) & (g868) & (g1040) & (!g1079) & (g1080) & (!g1081)) + ((!g683) & (g868) & (g1040) & (g1079) & (!g1080) & (!g1081)) + ((!g683) & (g868) & (g1040) & (g1079) & (g1080) & (!g1081)) + ((!g683) & (g868) & (g1040) & (g1079) & (g1080) & (g1081)) + ((g683) & (!g868) & (!g1040) & (!g1079) & (!g1080) & (g1081)) + ((g683) & (!g868) & (!g1040) & (!g1079) & (g1080) & (g1081)) + ((g683) & (!g868) & (!g1040) & (g1079) & (!g1080) & (g1081)) + ((g683) & (!g868) & (!g1040) & (g1079) & (g1080) & (g1081)) + ((g683) & (!g868) & (g1040) & (!g1079) & (!g1080) & (g1081)) + ((g683) & (!g868) & (g1040) & (!g1079) & (g1080) & (g1081)) + ((g683) & (!g868) & (g1040) & (g1079) & (!g1080) & (g1081)) + ((g683) & (!g868) & (g1040) & (g1079) & (g1080) & (g1081)) + ((g683) & (g868) & (!g1040) & (!g1079) & (!g1080) & (g1081)) + ((g683) & (g868) & (!g1040) & (g1079) & (g1080) & (g1081)) + ((g683) & (g868) & (g1040) & (!g1079) & (g1080) & (g1081)) + ((g683) & (g868) & (g1040) & (g1079) & (!g1080) & (g1081)));
	assign g1083 = (((!g979) & (!g981) & (!g982) & (!g988) & (!g1047) & (!g1054)) + ((!g979) & (!g981) & (!g982) & (!g988) & (g1047) & (!g1054)) + ((!g979) & (!g981) & (!g982) & (!g988) & (g1047) & (g1054)) + ((!g979) & (!g981) & (!g982) & (g988) & (g1047) & (!g1054)) + ((!g979) & (!g981) & (g982) & (!g988) & (g1047) & (!g1054)) + ((!g979) & (!g981) & (g982) & (g988) & (!g1047) & (!g1054)) + ((!g979) & (!g981) & (g982) & (g988) & (g1047) & (!g1054)) + ((!g979) & (!g981) & (g982) & (g988) & (g1047) & (g1054)) + ((!g979) & (g981) & (!g982) & (!g988) & (g1047) & (!g1054)) + ((!g979) & (g981) & (!g982) & (g988) & (g1047) & (!g1054)) + ((!g979) & (g981) & (g982) & (!g988) & (g1047) & (!g1054)) + ((!g979) & (g981) & (g982) & (g988) & (g1047) & (!g1054)) + ((g979) & (!g981) & (!g982) & (!g988) & (!g1047) & (!g1054)) + ((g979) & (!g981) & (!g982) & (!g988) & (g1047) & (!g1054)) + ((g979) & (!g981) & (!g982) & (!g988) & (g1047) & (g1054)) + ((g979) & (!g981) & (!g982) & (g988) & (!g1047) & (!g1054)) + ((g979) & (!g981) & (!g982) & (g988) & (g1047) & (!g1054)) + ((g979) & (!g981) & (!g982) & (g988) & (g1047) & (g1054)) + ((g979) & (!g981) & (g982) & (!g988) & (!g1047) & (!g1054)) + ((g979) & (!g981) & (g982) & (!g988) & (g1047) & (!g1054)) + ((g979) & (!g981) & (g982) & (!g988) & (g1047) & (g1054)) + ((g979) & (!g981) & (g982) & (g988) & (!g1047) & (!g1054)) + ((g979) & (!g981) & (g982) & (g988) & (g1047) & (!g1054)) + ((g979) & (!g981) & (g982) & (g988) & (g1047) & (g1054)) + ((g979) & (g981) & (!g982) & (!g988) & (!g1047) & (!g1054)) + ((g979) & (g981) & (!g982) & (!g988) & (g1047) & (!g1054)) + ((g979) & (g981) & (!g982) & (!g988) & (g1047) & (g1054)) + ((g979) & (g981) & (!g982) & (g988) & (g1047) & (!g1054)) + ((g979) & (g981) & (g982) & (!g988) & (g1047) & (!g1054)) + ((g979) & (g981) & (g982) & (g988) & (!g1047) & (!g1054)) + ((g979) & (g981) & (g982) & (g988) & (g1047) & (!g1054)) + ((g979) & (g981) & (g982) & (g988) & (g1047) & (g1054)));
	assign g1084 = (((!sk[70]) & (!g747) & (!g744) & (!g870) & (g863)) + ((!sk[70]) & (!g747) & (!g744) & (g870) & (g863)) + ((!sk[70]) & (!g747) & (g744) & (!g870) & (g863)) + ((!sk[70]) & (!g747) & (g744) & (g870) & (g863)) + ((!sk[70]) & (g747) & (!g744) & (!g870) & (!g863)) + ((!sk[70]) & (g747) & (!g744) & (!g870) & (g863)) + ((!sk[70]) & (g747) & (!g744) & (g870) & (!g863)) + ((!sk[70]) & (g747) & (!g744) & (g870) & (g863)) + ((!sk[70]) & (g747) & (g744) & (!g870) & (!g863)) + ((!sk[70]) & (g747) & (g744) & (!g870) & (g863)) + ((!sk[70]) & (g747) & (g744) & (g870) & (!g863)) + ((!sk[70]) & (g747) & (g744) & (g870) & (g863)) + ((sk[70]) & (!g747) & (g744) & (!g870) & (!g863)) + ((sk[70]) & (!g747) & (g744) & (!g870) & (g863)) + ((sk[70]) & (g747) & (!g744) & (!g870) & (g863)) + ((sk[70]) & (g747) & (!g744) & (g870) & (g863)) + ((sk[70]) & (g747) & (g744) & (!g870) & (!g863)) + ((sk[70]) & (g747) & (g744) & (!g870) & (g863)) + ((sk[70]) & (g747) & (g744) & (g870) & (g863)));
	assign g1085 = (((!g200) & (!g869) & (!g742) & (!g748) & (!g899) & (g1084)) + ((!g200) & (!g869) & (!g742) & (!g748) & (g899) & (g1084)) + ((!g200) & (!g869) & (!g742) & (g748) & (!g899) & (g1084)) + ((!g200) & (!g869) & (!g742) & (g748) & (g899) & (g1084)) + ((!g200) & (!g869) & (g742) & (!g748) & (!g899) & (!g1084)) + ((!g200) & (!g869) & (g742) & (!g748) & (!g899) & (g1084)) + ((!g200) & (!g869) & (g742) & (!g748) & (g899) & (g1084)) + ((!g200) & (!g869) & (g742) & (g748) & (!g899) & (!g1084)) + ((!g200) & (!g869) & (g742) & (g748) & (!g899) & (g1084)) + ((!g200) & (!g869) & (g742) & (g748) & (g899) & (g1084)) + ((!g200) & (g869) & (!g742) & (!g748) & (!g899) & (g1084)) + ((!g200) & (g869) & (!g742) & (!g748) & (g899) & (g1084)) + ((!g200) & (g869) & (!g742) & (g748) & (!g899) & (!g1084)) + ((!g200) & (g869) & (!g742) & (g748) & (!g899) & (g1084)) + ((!g200) & (g869) & (!g742) & (g748) & (g899) & (!g1084)) + ((!g200) & (g869) & (!g742) & (g748) & (g899) & (g1084)) + ((!g200) & (g869) & (g742) & (!g748) & (!g899) & (!g1084)) + ((!g200) & (g869) & (g742) & (!g748) & (!g899) & (g1084)) + ((!g200) & (g869) & (g742) & (!g748) & (g899) & (g1084)) + ((!g200) & (g869) & (g742) & (g748) & (!g899) & (!g1084)) + ((!g200) & (g869) & (g742) & (g748) & (!g899) & (g1084)) + ((!g200) & (g869) & (g742) & (g748) & (g899) & (!g1084)) + ((!g200) & (g869) & (g742) & (g748) & (g899) & (g1084)) + ((g200) & (!g869) & (!g742) & (!g748) & (!g899) & (!g1084)) + ((g200) & (!g869) & (!g742) & (!g748) & (g899) & (!g1084)) + ((g200) & (!g869) & (!g742) & (g748) & (!g899) & (!g1084)) + ((g200) & (!g869) & (!g742) & (g748) & (g899) & (!g1084)) + ((g200) & (!g869) & (g742) & (!g748) & (g899) & (!g1084)) + ((g200) & (!g869) & (g742) & (g748) & (g899) & (!g1084)) + ((g200) & (g869) & (!g742) & (!g748) & (!g899) & (!g1084)) + ((g200) & (g869) & (!g742) & (!g748) & (g899) & (!g1084)) + ((g200) & (g869) & (g742) & (!g748) & (g899) & (!g1084)));
	assign g1086 = (((!g1048) & (g1051) & (!sk[72]) & (!g1053)) + ((!g1048) & (g1051) & (!sk[72]) & (g1053)) + ((!g1048) & (g1051) & (sk[72]) & (!g1053)) + ((g1048) & (!g1051) & (sk[72]) & (!g1053)) + ((g1048) & (g1051) & (!sk[72]) & (!g1053)) + ((g1048) & (g1051) & (!sk[72]) & (g1053)) + ((g1048) & (g1051) & (sk[72]) & (!g1053)) + ((g1048) & (g1051) & (sk[72]) & (g1053)));
	assign g1087 = (((!g549) & (!g569) & (!g680) & (!g729) & (!g762) & (g765)) + ((!g549) & (!g569) & (!g680) & (!g729) & (g762) & (g765)) + ((!g549) & (!g569) & (g680) & (!g729) & (!g762) & (g765)) + ((!g549) & (!g569) & (g680) & (!g729) & (g762) & (!g765)) + ((!g549) & (!g569) & (g680) & (!g729) & (g762) & (g765)) + ((!g549) & (!g569) & (g680) & (g729) & (g762) & (!g765)) + ((!g549) & (!g569) & (g680) & (g729) & (g762) & (g765)) + ((!g549) & (g569) & (!g680) & (!g729) & (!g762) & (g765)) + ((!g549) & (g569) & (!g680) & (!g729) & (g762) & (!g765)) + ((!g549) & (g569) & (!g680) & (!g729) & (g762) & (g765)) + ((!g549) & (g569) & (!g680) & (g729) & (g762) & (!g765)) + ((!g549) & (g569) & (!g680) & (g729) & (g762) & (g765)) + ((!g549) & (g569) & (g680) & (!g729) & (!g762) & (g765)) + ((!g549) & (g569) & (g680) & (!g729) & (g762) & (g765)) + ((g549) & (!g569) & (!g680) & (!g729) & (!g762) & (g765)) + ((g549) & (!g569) & (!g680) & (!g729) & (g762) & (!g765)) + ((g549) & (!g569) & (!g680) & (!g729) & (g762) & (g765)) + ((g549) & (!g569) & (!g680) & (g729) & (g762) & (!g765)) + ((g549) & (!g569) & (!g680) & (g729) & (g762) & (g765)) + ((g549) & (!g569) & (g680) & (!g729) & (!g762) & (g765)) + ((g549) & (!g569) & (g680) & (!g729) & (g762) & (g765)) + ((g549) & (g569) & (!g680) & (!g729) & (!g762) & (g765)) + ((g549) & (g569) & (!g680) & (!g729) & (g762) & (g765)) + ((g549) & (g569) & (g680) & (!g729) & (!g762) & (g765)) + ((g549) & (g569) & (g680) & (!g729) & (g762) & (!g765)) + ((g549) & (g569) & (g680) & (!g729) & (g762) & (g765)) + ((g549) & (g569) & (g680) & (g729) & (g762) & (!g765)) + ((g549) & (g569) & (g680) & (g729) & (g762) & (g765)));
	assign g1088 = (((!g681) & (!g718) & (!g730) & (!g764) & (!g759) & (!g1087)) + ((!g681) & (!g718) & (!g730) & (g764) & (!g759) & (!g1087)) + ((!g681) & (!g718) & (g730) & (!g764) & (!g759) & (!g1087)) + ((!g681) & (!g718) & (g730) & (!g764) & (g759) & (!g1087)) + ((!g681) & (!g718) & (g730) & (g764) & (!g759) & (!g1087)) + ((!g681) & (!g718) & (g730) & (g764) & (g759) & (!g1087)) + ((!g681) & (g718) & (!g730) & (!g764) & (!g759) & (!g1087)) + ((!g681) & (g718) & (!g730) & (!g764) & (g759) & (!g1087)) + ((!g681) & (g718) & (g730) & (!g764) & (!g759) & (!g1087)) + ((g681) & (!g718) & (!g730) & (!g764) & (!g759) & (!g1087)) + ((g681) & (!g718) & (!g730) & (!g764) & (g759) & (!g1087)) + ((g681) & (!g718) & (!g730) & (g764) & (!g759) & (!g1087)) + ((g681) & (!g718) & (!g730) & (g764) & (g759) & (!g1087)) + ((g681) & (!g718) & (g730) & (!g764) & (!g759) & (!g1087)) + ((g681) & (!g718) & (g730) & (g764) & (!g759) & (!g1087)) + ((g681) & (g718) & (!g730) & (!g764) & (!g759) & (!g1087)) + ((g681) & (g718) & (g730) & (!g764) & (!g759) & (!g1087)) + ((g681) & (g718) & (g730) & (!g764) & (g759) & (!g1087)));
	assign g1089 = (((!g252) & (!g724) & (!g985) & (g986) & (!g1447) & (!g1050)) + ((!g252) & (!g724) & (g985) & (!g986) & (g1447) & (!g1050)) + ((!g252) & (!g724) & (g985) & (g986) & (!g1447) & (!g1050)) + ((!g252) & (!g724) & (g985) & (g986) & (g1447) & (!g1050)) + ((!g252) & (g724) & (!g985) & (g986) & (!g1447) & (!g1050)) + ((!g252) & (g724) & (g985) & (!g986) & (g1447) & (!g1050)) + ((!g252) & (g724) & (g985) & (g986) & (!g1447) & (!g1050)) + ((!g252) & (g724) & (g985) & (g986) & (g1447) & (!g1050)) + ((g252) & (!g724) & (!g985) & (!g986) & (!g1447) & (g1050)) + ((g252) & (!g724) & (!g985) & (!g986) & (g1447) & (g1050)) + ((g252) & (!g724) & (!g985) & (g986) & (!g1447) & (!g1050)) + ((g252) & (!g724) & (!g985) & (g986) & (!g1447) & (g1050)) + ((g252) & (!g724) & (!g985) & (g986) & (g1447) & (g1050)) + ((g252) & (!g724) & (g985) & (!g986) & (!g1447) & (!g1050)) + ((g252) & (!g724) & (g985) & (!g986) & (!g1447) & (g1050)) + ((g252) & (!g724) & (g985) & (!g986) & (g1447) & (g1050)) + ((g252) & (!g724) & (g985) & (g986) & (!g1447) & (!g1050)) + ((g252) & (!g724) & (g985) & (g986) & (!g1447) & (g1050)) + ((g252) & (!g724) & (g985) & (g986) & (g1447) & (!g1050)) + ((g252) & (!g724) & (g985) & (g986) & (g1447) & (g1050)) + ((g252) & (g724) & (!g985) & (g986) & (!g1447) & (g1050)) + ((g252) & (g724) & (g985) & (!g986) & (!g1447) & (g1050)) + ((g252) & (g724) & (g985) & (g986) & (!g1447) & (g1050)) + ((g252) & (g724) & (g985) & (g986) & (g1447) & (g1050)));
	assign g1090 = (((!g585) & (!g597) & (!g679) & (g720) & (!g847) & (g845)) + ((!g585) & (!g597) & (!g679) & (g720) & (g847) & (g845)) + ((!g585) & (!g597) & (g679) & (!g720) & (g847) & (!g845)) + ((!g585) & (!g597) & (g679) & (!g720) & (g847) & (g845)) + ((!g585) & (!g597) & (g679) & (g720) & (!g847) & (g845)) + ((!g585) & (!g597) & (g679) & (g720) & (g847) & (!g845)) + ((!g585) & (!g597) & (g679) & (g720) & (g847) & (g845)) + ((!g585) & (g597) & (!g679) & (!g720) & (g847) & (!g845)) + ((!g585) & (g597) & (!g679) & (!g720) & (g847) & (g845)) + ((!g585) & (g597) & (!g679) & (g720) & (!g847) & (g845)) + ((!g585) & (g597) & (!g679) & (g720) & (g847) & (!g845)) + ((!g585) & (g597) & (!g679) & (g720) & (g847) & (g845)) + ((!g585) & (g597) & (g679) & (g720) & (!g847) & (g845)) + ((!g585) & (g597) & (g679) & (g720) & (g847) & (g845)) + ((g585) & (!g597) & (!g679) & (!g720) & (g847) & (!g845)) + ((g585) & (!g597) & (!g679) & (!g720) & (g847) & (g845)) + ((g585) & (!g597) & (!g679) & (g720) & (!g847) & (g845)) + ((g585) & (!g597) & (!g679) & (g720) & (g847) & (!g845)) + ((g585) & (!g597) & (!g679) & (g720) & (g847) & (g845)) + ((g585) & (!g597) & (g679) & (g720) & (!g847) & (g845)) + ((g585) & (!g597) & (g679) & (g720) & (g847) & (g845)) + ((g585) & (g597) & (!g679) & (g720) & (!g847) & (g845)) + ((g585) & (g597) & (!g679) & (g720) & (g847) & (g845)) + ((g585) & (g597) & (g679) & (!g720) & (g847) & (!g845)) + ((g585) & (g597) & (g679) & (!g720) & (g847) & (g845)) + ((g585) & (g597) & (g679) & (g720) & (!g847) & (g845)) + ((g585) & (g597) & (g679) & (g720) & (g847) & (!g845)) + ((g585) & (g597) & (g679) & (g720) & (g847) & (g845)));
	assign g1091 = (((!g722) & (!g771) & (!sk[77]) & (!g843) & (g848) & (!g1090)) + ((!g722) & (!g771) & (!sk[77]) & (!g843) & (g848) & (g1090)) + ((!g722) & (!g771) & (!sk[77]) & (g843) & (!g848) & (!g1090)) + ((!g722) & (!g771) & (!sk[77]) & (g843) & (!g848) & (g1090)) + ((!g722) & (!g771) & (!sk[77]) & (g843) & (g848) & (!g1090)) + ((!g722) & (!g771) & (!sk[77]) & (g843) & (g848) & (g1090)) + ((!g722) & (!g771) & (sk[77]) & (!g843) & (!g848) & (!g1090)) + ((!g722) & (g771) & (!sk[77]) & (!g843) & (!g848) & (!g1090)) + ((!g722) & (g771) & (!sk[77]) & (!g843) & (!g848) & (g1090)) + ((!g722) & (g771) & (!sk[77]) & (!g843) & (g848) & (!g1090)) + ((!g722) & (g771) & (!sk[77]) & (!g843) & (g848) & (g1090)) + ((!g722) & (g771) & (!sk[77]) & (g843) & (!g848) & (!g1090)) + ((!g722) & (g771) & (!sk[77]) & (g843) & (!g848) & (g1090)) + ((!g722) & (g771) & (!sk[77]) & (g843) & (g848) & (!g1090)) + ((!g722) & (g771) & (!sk[77]) & (g843) & (g848) & (g1090)) + ((!g722) & (g771) & (sk[77]) & (!g843) & (!g848) & (!g1090)) + ((!g722) & (g771) & (sk[77]) & (g843) & (!g848) & (!g1090)) + ((g722) & (!g771) & (!sk[77]) & (!g843) & (g848) & (!g1090)) + ((g722) & (!g771) & (!sk[77]) & (!g843) & (g848) & (g1090)) + ((g722) & (!g771) & (!sk[77]) & (g843) & (!g848) & (!g1090)) + ((g722) & (!g771) & (!sk[77]) & (g843) & (!g848) & (g1090)) + ((g722) & (!g771) & (!sk[77]) & (g843) & (g848) & (!g1090)) + ((g722) & (!g771) & (!sk[77]) & (g843) & (g848) & (g1090)) + ((g722) & (!g771) & (sk[77]) & (!g843) & (!g848) & (!g1090)) + ((g722) & (!g771) & (sk[77]) & (!g843) & (g848) & (!g1090)) + ((g722) & (g771) & (!sk[77]) & (!g843) & (!g848) & (!g1090)) + ((g722) & (g771) & (!sk[77]) & (!g843) & (!g848) & (g1090)) + ((g722) & (g771) & (!sk[77]) & (!g843) & (g848) & (!g1090)) + ((g722) & (g771) & (!sk[77]) & (!g843) & (g848) & (g1090)) + ((g722) & (g771) & (!sk[77]) & (g843) & (!g848) & (!g1090)) + ((g722) & (g771) & (!sk[77]) & (g843) & (!g848) & (g1090)) + ((g722) & (g771) & (!sk[77]) & (g843) & (g848) & (!g1090)) + ((g722) & (g771) & (!sk[77]) & (g843) & (g848) & (g1090)) + ((g722) & (g771) & (sk[77]) & (!g843) & (!g848) & (!g1090)) + ((g722) & (g771) & (sk[77]) & (!g843) & (g848) & (!g1090)) + ((g722) & (g771) & (sk[77]) & (g843) & (!g848) & (!g1090)) + ((g722) & (g771) & (sk[77]) & (g843) & (g848) & (!g1090)));
	assign g1092 = (((!sk[78]) & (!g252) & (!g723) & (!g1089) & (g1091)) + ((!sk[78]) & (!g252) & (!g723) & (g1089) & (g1091)) + ((!sk[78]) & (!g252) & (g723) & (!g1089) & (g1091)) + ((!sk[78]) & (!g252) & (g723) & (g1089) & (g1091)) + ((!sk[78]) & (g252) & (!g723) & (!g1089) & (!g1091)) + ((!sk[78]) & (g252) & (!g723) & (!g1089) & (g1091)) + ((!sk[78]) & (g252) & (!g723) & (g1089) & (!g1091)) + ((!sk[78]) & (g252) & (!g723) & (g1089) & (g1091)) + ((!sk[78]) & (g252) & (g723) & (!g1089) & (!g1091)) + ((!sk[78]) & (g252) & (g723) & (!g1089) & (g1091)) + ((!sk[78]) & (g252) & (g723) & (g1089) & (!g1091)) + ((!sk[78]) & (g252) & (g723) & (g1089) & (g1091)) + ((sk[78]) & (!g252) & (!g723) & (!g1089) & (!g1091)) + ((sk[78]) & (!g252) & (!g723) & (g1089) & (g1091)) + ((sk[78]) & (!g252) & (g723) & (!g1089) & (!g1091)) + ((sk[78]) & (!g252) & (g723) & (g1089) & (g1091)) + ((sk[78]) & (g252) & (!g723) & (!g1089) & (!g1091)) + ((sk[78]) & (g252) & (!g723) & (g1089) & (g1091)) + ((sk[78]) & (g252) & (g723) & (!g1089) & (g1091)) + ((sk[78]) & (g252) & (g723) & (g1089) & (!g1091)));
	assign g1093 = (((!g202) & (!sk[79]) & (g1088) & (!g1092)) + ((!g202) & (!sk[79]) & (g1088) & (g1092)) + ((!g202) & (sk[79]) & (!g1088) & (g1092)) + ((!g202) & (sk[79]) & (g1088) & (!g1092)) + ((g202) & (!sk[79]) & (g1088) & (!g1092)) + ((g202) & (!sk[79]) & (g1088) & (g1092)) + ((g202) & (sk[79]) & (!g1088) & (!g1092)) + ((g202) & (sk[79]) & (g1088) & (g1092)));
	assign g1094 = (((!g1083) & (!g1085) & (!g1086) & (!sk[80]) & (g1093)) + ((!g1083) & (!g1085) & (!g1086) & (sk[80]) & (g1093)) + ((!g1083) & (!g1085) & (g1086) & (!sk[80]) & (g1093)) + ((!g1083) & (!g1085) & (g1086) & (sk[80]) & (!g1093)) + ((!g1083) & (g1085) & (!g1086) & (!sk[80]) & (g1093)) + ((!g1083) & (g1085) & (!g1086) & (sk[80]) & (!g1093)) + ((!g1083) & (g1085) & (g1086) & (!sk[80]) & (g1093)) + ((!g1083) & (g1085) & (g1086) & (sk[80]) & (g1093)) + ((g1083) & (!g1085) & (!g1086) & (!sk[80]) & (!g1093)) + ((g1083) & (!g1085) & (!g1086) & (!sk[80]) & (g1093)) + ((g1083) & (!g1085) & (!g1086) & (sk[80]) & (!g1093)) + ((g1083) & (!g1085) & (g1086) & (!sk[80]) & (!g1093)) + ((g1083) & (!g1085) & (g1086) & (!sk[80]) & (g1093)) + ((g1083) & (!g1085) & (g1086) & (sk[80]) & (g1093)) + ((g1083) & (g1085) & (!g1086) & (!sk[80]) & (!g1093)) + ((g1083) & (g1085) & (!g1086) & (!sk[80]) & (g1093)) + ((g1083) & (g1085) & (!g1086) & (sk[80]) & (g1093)) + ((g1083) & (g1085) & (g1086) & (!sk[80]) & (!g1093)) + ((g1083) & (g1085) & (g1086) & (!sk[80]) & (g1093)) + ((g1083) & (g1085) & (g1086) & (sk[80]) & (!g1093)));
	assign g1095 = (((!g733) & (!g686) & (!g734) & (!g962) & (!g963) & (!g971)) + ((!g733) & (!g686) & (!g734) & (!g962) & (!g963) & (g971)) + ((!g733) & (!g686) & (!g734) & (!g962) & (g963) & (!g971)) + ((!g733) & (!g686) & (!g734) & (!g962) & (g963) & (g971)) + ((!g733) & (!g686) & (!g734) & (g962) & (!g963) & (!g971)) + ((!g733) & (!g686) & (!g734) & (g962) & (!g963) & (g971)) + ((!g733) & (!g686) & (!g734) & (g962) & (g963) & (!g971)) + ((!g733) & (!g686) & (!g734) & (g962) & (g963) & (g971)) + ((!g733) & (!g686) & (g734) & (g962) & (!g963) & (!g971)) + ((!g733) & (!g686) & (g734) & (g962) & (!g963) & (g971)) + ((!g733) & (!g686) & (g734) & (g962) & (g963) & (!g971)) + ((!g733) & (!g686) & (g734) & (g962) & (g963) & (g971)) + ((!g733) & (g686) & (!g734) & (!g962) & (!g963) & (!g971)) + ((!g733) & (g686) & (!g734) & (!g962) & (!g963) & (g971)) + ((!g733) & (g686) & (!g734) & (g962) & (!g963) & (!g971)) + ((!g733) & (g686) & (!g734) & (g962) & (!g963) & (g971)) + ((!g733) & (g686) & (g734) & (g962) & (!g963) & (!g971)) + ((!g733) & (g686) & (g734) & (g962) & (!g963) & (g971)) + ((g733) & (!g686) & (!g734) & (!g962) & (!g963) & (!g971)) + ((g733) & (!g686) & (!g734) & (!g962) & (g963) & (!g971)) + ((g733) & (!g686) & (!g734) & (g962) & (!g963) & (!g971)) + ((g733) & (!g686) & (!g734) & (g962) & (g963) & (!g971)) + ((g733) & (!g686) & (g734) & (g962) & (!g963) & (!g971)) + ((g733) & (!g686) & (g734) & (g962) & (g963) & (!g971)) + ((g733) & (g686) & (!g734) & (!g962) & (!g963) & (!g971)) + ((g733) & (g686) & (!g734) & (g962) & (!g963) & (!g971)) + ((g733) & (g686) & (g734) & (g962) & (!g963) & (!g971)));
	assign g1096 = (((!g2) & (!g732) & (!sk[82]) & (!g972) & (g1095)) + ((!g2) & (!g732) & (!sk[82]) & (g972) & (g1095)) + ((!g2) & (!g732) & (sk[82]) & (!g972) & (g1095)) + ((!g2) & (!g732) & (sk[82]) & (g972) & (g1095)) + ((!g2) & (g732) & (!sk[82]) & (!g972) & (g1095)) + ((!g2) & (g732) & (!sk[82]) & (g972) & (g1095)) + ((!g2) & (g732) & (sk[82]) & (g972) & (g1095)) + ((g2) & (!g732) & (!sk[82]) & (!g972) & (!g1095)) + ((g2) & (!g732) & (!sk[82]) & (!g972) & (g1095)) + ((g2) & (!g732) & (!sk[82]) & (g972) & (!g1095)) + ((g2) & (!g732) & (!sk[82]) & (g972) & (g1095)) + ((g2) & (!g732) & (sk[82]) & (!g972) & (!g1095)) + ((g2) & (!g732) & (sk[82]) & (g972) & (!g1095)) + ((g2) & (g732) & (!sk[82]) & (!g972) & (!g1095)) + ((g2) & (g732) & (!sk[82]) & (!g972) & (g1095)) + ((g2) & (g732) & (!sk[82]) & (g972) & (!g1095)) + ((g2) & (g732) & (!sk[82]) & (g972) & (g1095)) + ((g2) & (g732) & (sk[82]) & (!g972) & (!g1095)) + ((g2) & (g732) & (sk[82]) & (!g972) & (g1095)) + ((g2) & (g732) & (sk[82]) & (g972) & (!g1095)));
	assign g1097 = (((!g1044) & (!g1055) & (!g1058) & (!g1082) & (!g1094) & (!g1096)) + ((!g1044) & (!g1055) & (!g1058) & (!g1082) & (g1094) & (g1096)) + ((!g1044) & (!g1055) & (!g1058) & (g1082) & (!g1094) & (g1096)) + ((!g1044) & (!g1055) & (!g1058) & (g1082) & (g1094) & (!g1096)) + ((!g1044) & (!g1055) & (g1058) & (!g1082) & (!g1094) & (g1096)) + ((!g1044) & (!g1055) & (g1058) & (!g1082) & (g1094) & (!g1096)) + ((!g1044) & (!g1055) & (g1058) & (g1082) & (!g1094) & (!g1096)) + ((!g1044) & (!g1055) & (g1058) & (g1082) & (g1094) & (g1096)) + ((!g1044) & (g1055) & (!g1058) & (!g1082) & (!g1094) & (g1096)) + ((!g1044) & (g1055) & (!g1058) & (!g1082) & (g1094) & (!g1096)) + ((!g1044) & (g1055) & (!g1058) & (g1082) & (!g1094) & (!g1096)) + ((!g1044) & (g1055) & (!g1058) & (g1082) & (g1094) & (g1096)) + ((!g1044) & (g1055) & (g1058) & (!g1082) & (!g1094) & (g1096)) + ((!g1044) & (g1055) & (g1058) & (!g1082) & (g1094) & (!g1096)) + ((!g1044) & (g1055) & (g1058) & (g1082) & (!g1094) & (!g1096)) + ((!g1044) & (g1055) & (g1058) & (g1082) & (g1094) & (g1096)) + ((g1044) & (!g1055) & (!g1058) & (!g1082) & (!g1094) & (!g1096)) + ((g1044) & (!g1055) & (!g1058) & (!g1082) & (g1094) & (g1096)) + ((g1044) & (!g1055) & (!g1058) & (g1082) & (!g1094) & (g1096)) + ((g1044) & (!g1055) & (!g1058) & (g1082) & (g1094) & (!g1096)) + ((g1044) & (!g1055) & (g1058) & (!g1082) & (!g1094) & (!g1096)) + ((g1044) & (!g1055) & (g1058) & (!g1082) & (g1094) & (g1096)) + ((g1044) & (!g1055) & (g1058) & (g1082) & (!g1094) & (g1096)) + ((g1044) & (!g1055) & (g1058) & (g1082) & (g1094) & (!g1096)) + ((g1044) & (g1055) & (!g1058) & (!g1082) & (!g1094) & (!g1096)) + ((g1044) & (g1055) & (!g1058) & (!g1082) & (g1094) & (g1096)) + ((g1044) & (g1055) & (!g1058) & (g1082) & (!g1094) & (g1096)) + ((g1044) & (g1055) & (!g1058) & (g1082) & (g1094) & (!g1096)) + ((g1044) & (g1055) & (g1058) & (!g1082) & (!g1094) & (g1096)) + ((g1044) & (g1055) & (g1058) & (!g1082) & (g1094) & (!g1096)) + ((g1044) & (g1055) & (g1058) & (g1082) & (!g1094) & (!g1096)) + ((g1044) & (g1055) & (g1058) & (g1082) & (g1094) & (g1096)));
	assign g1098 = (((!g975) & (!g990) & (!g997) & (!g1043) & (!g1059) & (g1097)) + ((!g975) & (!g990) & (!g997) & (!g1043) & (g1059) & (g1097)) + ((!g975) & (!g990) & (!g997) & (g1043) & (!g1059) & (g1097)) + ((!g975) & (!g990) & (!g997) & (g1043) & (g1059) & (!g1097)) + ((!g975) & (!g990) & (g997) & (!g1043) & (!g1059) & (g1097)) + ((!g975) & (!g990) & (g997) & (!g1043) & (g1059) & (g1097)) + ((!g975) & (!g990) & (g997) & (g1043) & (!g1059) & (g1097)) + ((!g975) & (!g990) & (g997) & (g1043) & (g1059) & (!g1097)) + ((!g975) & (g990) & (!g997) & (!g1043) & (!g1059) & (g1097)) + ((!g975) & (g990) & (!g997) & (!g1043) & (g1059) & (!g1097)) + ((!g975) & (g990) & (!g997) & (g1043) & (!g1059) & (!g1097)) + ((!g975) & (g990) & (!g997) & (g1043) & (g1059) & (!g1097)) + ((!g975) & (g990) & (g997) & (!g1043) & (!g1059) & (g1097)) + ((!g975) & (g990) & (g997) & (!g1043) & (g1059) & (g1097)) + ((!g975) & (g990) & (g997) & (g1043) & (!g1059) & (g1097)) + ((!g975) & (g990) & (g997) & (g1043) & (g1059) & (!g1097)) + ((g975) & (!g990) & (!g997) & (!g1043) & (!g1059) & (g1097)) + ((g975) & (!g990) & (!g997) & (!g1043) & (g1059) & (!g1097)) + ((g975) & (!g990) & (!g997) & (g1043) & (!g1059) & (!g1097)) + ((g975) & (!g990) & (!g997) & (g1043) & (g1059) & (!g1097)) + ((g975) & (!g990) & (g997) & (!g1043) & (!g1059) & (g1097)) + ((g975) & (!g990) & (g997) & (!g1043) & (g1059) & (g1097)) + ((g975) & (!g990) & (g997) & (g1043) & (!g1059) & (g1097)) + ((g975) & (!g990) & (g997) & (g1043) & (g1059) & (!g1097)) + ((g975) & (g990) & (!g997) & (!g1043) & (!g1059) & (g1097)) + ((g975) & (g990) & (!g997) & (!g1043) & (g1059) & (!g1097)) + ((g975) & (g990) & (!g997) & (g1043) & (!g1059) & (!g1097)) + ((g975) & (g990) & (!g997) & (g1043) & (g1059) & (!g1097)) + ((g975) & (g990) & (g997) & (!g1043) & (!g1059) & (g1097)) + ((g975) & (g990) & (g997) & (!g1043) & (g1059) & (!g1097)) + ((g975) & (g990) & (g997) & (g1043) & (!g1059) & (!g1097)) + ((g975) & (g990) & (g997) & (g1043) & (g1059) & (!g1097)));
	assign g1099 = (((!g879) & (g72) & (!sk[85]) & (!g73)) + ((!g879) & (g72) & (!sk[85]) & (g73)) + ((g879) & (!g72) & (sk[85]) & (!g73)) + ((g879) & (g72) & (!sk[85]) & (!g73)) + ((g879) & (g72) & (!sk[85]) & (g73)));
	assign g1100 = (((!g16) & (!sk[86]) & (g25) & (!g185)) + ((!g16) & (!sk[86]) & (g25) & (g185)) + ((!g16) & (sk[86]) & (!g25) & (!g185)) + ((!g16) & (sk[86]) & (g25) & (!g185)) + ((g16) & (!sk[86]) & (g25) & (!g185)) + ((g16) & (!sk[86]) & (g25) & (g185)) + ((g16) & (sk[86]) & (!g25) & (!g185)));
	assign g1101 = (((!g9) & (!g10) & (!sk[87]) & (!g267) & (g551)) + ((!g9) & (!g10) & (!sk[87]) & (g267) & (g551)) + ((!g9) & (!g10) & (sk[87]) & (!g267) & (!g551)) + ((!g9) & (g10) & (!sk[87]) & (!g267) & (g551)) + ((!g9) & (g10) & (!sk[87]) & (g267) & (g551)) + ((!g9) & (g10) & (sk[87]) & (!g267) & (!g551)) + ((g9) & (!g10) & (!sk[87]) & (!g267) & (!g551)) + ((g9) & (!g10) & (!sk[87]) & (!g267) & (g551)) + ((g9) & (!g10) & (!sk[87]) & (g267) & (!g551)) + ((g9) & (!g10) & (!sk[87]) & (g267) & (g551)) + ((g9) & (!g10) & (sk[87]) & (!g267) & (!g551)) + ((g9) & (g10) & (!sk[87]) & (!g267) & (!g551)) + ((g9) & (g10) & (!sk[87]) & (!g267) & (g551)) + ((g9) & (g10) & (!sk[87]) & (g267) & (!g551)) + ((g9) & (g10) & (!sk[87]) & (g267) & (g551)));
	assign g1102 = (((!g16) & (!g18) & (!g1100) & (!sk[88]) & (g1101)) + ((!g16) & (!g18) & (g1100) & (!sk[88]) & (g1101)) + ((!g16) & (!g18) & (g1100) & (sk[88]) & (g1101)) + ((!g16) & (g18) & (!g1100) & (!sk[88]) & (g1101)) + ((!g16) & (g18) & (g1100) & (!sk[88]) & (g1101)) + ((!g16) & (g18) & (g1100) & (sk[88]) & (g1101)) + ((g16) & (!g18) & (!g1100) & (!sk[88]) & (!g1101)) + ((g16) & (!g18) & (!g1100) & (!sk[88]) & (g1101)) + ((g16) & (!g18) & (g1100) & (!sk[88]) & (!g1101)) + ((g16) & (!g18) & (g1100) & (!sk[88]) & (g1101)) + ((g16) & (!g18) & (g1100) & (sk[88]) & (g1101)) + ((g16) & (g18) & (!g1100) & (!sk[88]) & (!g1101)) + ((g16) & (g18) & (!g1100) & (!sk[88]) & (g1101)) + ((g16) & (g18) & (g1100) & (!sk[88]) & (!g1101)) + ((g16) & (g18) & (g1100) & (!sk[88]) & (g1101)));
	assign g1103 = (((!g114) & (!g115) & (!sk[89]) & (!g8) & (g17) & (!g18)) + ((!g114) & (!g115) & (!sk[89]) & (!g8) & (g17) & (g18)) + ((!g114) & (!g115) & (!sk[89]) & (g8) & (!g17) & (!g18)) + ((!g114) & (!g115) & (!sk[89]) & (g8) & (!g17) & (g18)) + ((!g114) & (!g115) & (!sk[89]) & (g8) & (g17) & (!g18)) + ((!g114) & (!g115) & (!sk[89]) & (g8) & (g17) & (g18)) + ((!g114) & (g115) & (!sk[89]) & (!g8) & (!g17) & (!g18)) + ((!g114) & (g115) & (!sk[89]) & (!g8) & (!g17) & (g18)) + ((!g114) & (g115) & (!sk[89]) & (!g8) & (g17) & (!g18)) + ((!g114) & (g115) & (!sk[89]) & (!g8) & (g17) & (g18)) + ((!g114) & (g115) & (!sk[89]) & (g8) & (!g17) & (!g18)) + ((!g114) & (g115) & (!sk[89]) & (g8) & (!g17) & (g18)) + ((!g114) & (g115) & (!sk[89]) & (g8) & (g17) & (!g18)) + ((!g114) & (g115) & (!sk[89]) & (g8) & (g17) & (g18)) + ((!g114) & (g115) & (sk[89]) & (g8) & (!g17) & (g18)) + ((!g114) & (g115) & (sk[89]) & (g8) & (g17) & (g18)) + ((g114) & (!g115) & (!sk[89]) & (!g8) & (g17) & (!g18)) + ((g114) & (!g115) & (!sk[89]) & (!g8) & (g17) & (g18)) + ((g114) & (!g115) & (!sk[89]) & (g8) & (!g17) & (!g18)) + ((g114) & (!g115) & (!sk[89]) & (g8) & (!g17) & (g18)) + ((g114) & (!g115) & (!sk[89]) & (g8) & (g17) & (!g18)) + ((g114) & (!g115) & (!sk[89]) & (g8) & (g17) & (g18)) + ((g114) & (!g115) & (sk[89]) & (!g8) & (g17) & (!g18)) + ((g114) & (!g115) & (sk[89]) & (!g8) & (g17) & (g18)) + ((g114) & (!g115) & (sk[89]) & (g8) & (!g17) & (g18)) + ((g114) & (!g115) & (sk[89]) & (g8) & (g17) & (g18)) + ((g114) & (g115) & (!sk[89]) & (!g8) & (!g17) & (!g18)) + ((g114) & (g115) & (!sk[89]) & (!g8) & (!g17) & (g18)) + ((g114) & (g115) & (!sk[89]) & (!g8) & (g17) & (!g18)) + ((g114) & (g115) & (!sk[89]) & (!g8) & (g17) & (g18)) + ((g114) & (g115) & (!sk[89]) & (g8) & (!g17) & (!g18)) + ((g114) & (g115) & (!sk[89]) & (g8) & (!g17) & (g18)) + ((g114) & (g115) & (!sk[89]) & (g8) & (g17) & (!g18)) + ((g114) & (g115) & (!sk[89]) & (g8) & (g17) & (g18)) + ((g114) & (g115) & (sk[89]) & (!g8) & (g17) & (!g18)) + ((g114) & (g115) & (sk[89]) & (!g8) & (g17) & (g18)));
	assign g1104 = (((!g9) & (!g40) & (!g622) & (!sk[90]) & (g876) & (!g1103)) + ((!g9) & (!g40) & (!g622) & (!sk[90]) & (g876) & (g1103)) + ((!g9) & (!g40) & (g622) & (!sk[90]) & (!g876) & (!g1103)) + ((!g9) & (!g40) & (g622) & (!sk[90]) & (!g876) & (g1103)) + ((!g9) & (!g40) & (g622) & (!sk[90]) & (g876) & (!g1103)) + ((!g9) & (!g40) & (g622) & (!sk[90]) & (g876) & (g1103)) + ((!g9) & (!g40) & (g622) & (sk[90]) & (g876) & (!g1103)) + ((!g9) & (g40) & (!g622) & (!sk[90]) & (!g876) & (!g1103)) + ((!g9) & (g40) & (!g622) & (!sk[90]) & (!g876) & (g1103)) + ((!g9) & (g40) & (!g622) & (!sk[90]) & (g876) & (!g1103)) + ((!g9) & (g40) & (!g622) & (!sk[90]) & (g876) & (g1103)) + ((!g9) & (g40) & (g622) & (!sk[90]) & (!g876) & (!g1103)) + ((!g9) & (g40) & (g622) & (!sk[90]) & (!g876) & (g1103)) + ((!g9) & (g40) & (g622) & (!sk[90]) & (g876) & (!g1103)) + ((!g9) & (g40) & (g622) & (!sk[90]) & (g876) & (g1103)) + ((!g9) & (g40) & (g622) & (sk[90]) & (g876) & (!g1103)) + ((g9) & (!g40) & (!g622) & (!sk[90]) & (g876) & (!g1103)) + ((g9) & (!g40) & (!g622) & (!sk[90]) & (g876) & (g1103)) + ((g9) & (!g40) & (g622) & (!sk[90]) & (!g876) & (!g1103)) + ((g9) & (!g40) & (g622) & (!sk[90]) & (!g876) & (g1103)) + ((g9) & (!g40) & (g622) & (!sk[90]) & (g876) & (!g1103)) + ((g9) & (!g40) & (g622) & (!sk[90]) & (g876) & (g1103)) + ((g9) & (!g40) & (g622) & (sk[90]) & (g876) & (!g1103)) + ((g9) & (g40) & (!g622) & (!sk[90]) & (!g876) & (!g1103)) + ((g9) & (g40) & (!g622) & (!sk[90]) & (!g876) & (g1103)) + ((g9) & (g40) & (!g622) & (!sk[90]) & (g876) & (!g1103)) + ((g9) & (g40) & (!g622) & (!sk[90]) & (g876) & (g1103)) + ((g9) & (g40) & (g622) & (!sk[90]) & (!g876) & (!g1103)) + ((g9) & (g40) & (g622) & (!sk[90]) & (!g876) & (g1103)) + ((g9) & (g40) & (g622) & (!sk[90]) & (g876) & (!g1103)) + ((g9) & (g40) & (g622) & (!sk[90]) & (g876) & (g1103)));
	assign g1105 = (((!g578) & (!sk[91]) & (!g1004) & (!g1099) & (g1102) & (!g1104)) + ((!g578) & (!sk[91]) & (!g1004) & (!g1099) & (g1102) & (g1104)) + ((!g578) & (!sk[91]) & (!g1004) & (g1099) & (!g1102) & (!g1104)) + ((!g578) & (!sk[91]) & (!g1004) & (g1099) & (!g1102) & (g1104)) + ((!g578) & (!sk[91]) & (!g1004) & (g1099) & (g1102) & (!g1104)) + ((!g578) & (!sk[91]) & (!g1004) & (g1099) & (g1102) & (g1104)) + ((!g578) & (!sk[91]) & (g1004) & (!g1099) & (!g1102) & (!g1104)) + ((!g578) & (!sk[91]) & (g1004) & (!g1099) & (!g1102) & (g1104)) + ((!g578) & (!sk[91]) & (g1004) & (!g1099) & (g1102) & (!g1104)) + ((!g578) & (!sk[91]) & (g1004) & (!g1099) & (g1102) & (g1104)) + ((!g578) & (!sk[91]) & (g1004) & (g1099) & (!g1102) & (!g1104)) + ((!g578) & (!sk[91]) & (g1004) & (g1099) & (!g1102) & (g1104)) + ((!g578) & (!sk[91]) & (g1004) & (g1099) & (g1102) & (!g1104)) + ((!g578) & (!sk[91]) & (g1004) & (g1099) & (g1102) & (g1104)) + ((g578) & (!sk[91]) & (!g1004) & (!g1099) & (g1102) & (!g1104)) + ((g578) & (!sk[91]) & (!g1004) & (!g1099) & (g1102) & (g1104)) + ((g578) & (!sk[91]) & (!g1004) & (g1099) & (!g1102) & (!g1104)) + ((g578) & (!sk[91]) & (!g1004) & (g1099) & (!g1102) & (g1104)) + ((g578) & (!sk[91]) & (!g1004) & (g1099) & (g1102) & (!g1104)) + ((g578) & (!sk[91]) & (!g1004) & (g1099) & (g1102) & (g1104)) + ((g578) & (!sk[91]) & (g1004) & (!g1099) & (!g1102) & (!g1104)) + ((g578) & (!sk[91]) & (g1004) & (!g1099) & (!g1102) & (g1104)) + ((g578) & (!sk[91]) & (g1004) & (!g1099) & (g1102) & (!g1104)) + ((g578) & (!sk[91]) & (g1004) & (!g1099) & (g1102) & (g1104)) + ((g578) & (!sk[91]) & (g1004) & (g1099) & (!g1102) & (!g1104)) + ((g578) & (!sk[91]) & (g1004) & (g1099) & (!g1102) & (g1104)) + ((g578) & (!sk[91]) & (g1004) & (g1099) & (g1102) & (!g1104)) + ((g578) & (!sk[91]) & (g1004) & (g1099) & (g1102) & (g1104)) + ((g578) & (sk[91]) & (g1004) & (g1099) & (g1102) & (g1104)));
	assign g1106 = (((!g1031) & (!g1060) & (!sk[92]) & (!g1065) & (g1098) & (!g1105)) + ((!g1031) & (!g1060) & (!sk[92]) & (!g1065) & (g1098) & (g1105)) + ((!g1031) & (!g1060) & (!sk[92]) & (g1065) & (!g1098) & (!g1105)) + ((!g1031) & (!g1060) & (!sk[92]) & (g1065) & (!g1098) & (g1105)) + ((!g1031) & (!g1060) & (!sk[92]) & (g1065) & (g1098) & (!g1105)) + ((!g1031) & (!g1060) & (!sk[92]) & (g1065) & (g1098) & (g1105)) + ((!g1031) & (!g1060) & (sk[92]) & (!g1065) & (!g1098) & (!g1105)) + ((!g1031) & (!g1060) & (sk[92]) & (!g1065) & (g1098) & (g1105)) + ((!g1031) & (!g1060) & (sk[92]) & (g1065) & (!g1098) & (!g1105)) + ((!g1031) & (!g1060) & (sk[92]) & (g1065) & (g1098) & (g1105)) + ((!g1031) & (g1060) & (!sk[92]) & (!g1065) & (!g1098) & (!g1105)) + ((!g1031) & (g1060) & (!sk[92]) & (!g1065) & (!g1098) & (g1105)) + ((!g1031) & (g1060) & (!sk[92]) & (!g1065) & (g1098) & (!g1105)) + ((!g1031) & (g1060) & (!sk[92]) & (!g1065) & (g1098) & (g1105)) + ((!g1031) & (g1060) & (!sk[92]) & (g1065) & (!g1098) & (!g1105)) + ((!g1031) & (g1060) & (!sk[92]) & (g1065) & (!g1098) & (g1105)) + ((!g1031) & (g1060) & (!sk[92]) & (g1065) & (g1098) & (!g1105)) + ((!g1031) & (g1060) & (!sk[92]) & (g1065) & (g1098) & (g1105)) + ((!g1031) & (g1060) & (sk[92]) & (!g1065) & (!g1098) & (g1105)) + ((!g1031) & (g1060) & (sk[92]) & (!g1065) & (g1098) & (!g1105)) + ((!g1031) & (g1060) & (sk[92]) & (g1065) & (!g1098) & (!g1105)) + ((!g1031) & (g1060) & (sk[92]) & (g1065) & (g1098) & (g1105)) + ((g1031) & (!g1060) & (!sk[92]) & (!g1065) & (g1098) & (!g1105)) + ((g1031) & (!g1060) & (!sk[92]) & (!g1065) & (g1098) & (g1105)) + ((g1031) & (!g1060) & (!sk[92]) & (g1065) & (!g1098) & (!g1105)) + ((g1031) & (!g1060) & (!sk[92]) & (g1065) & (!g1098) & (g1105)) + ((g1031) & (!g1060) & (!sk[92]) & (g1065) & (g1098) & (!g1105)) + ((g1031) & (!g1060) & (!sk[92]) & (g1065) & (g1098) & (g1105)) + ((g1031) & (!g1060) & (sk[92]) & (!g1065) & (!g1098) & (g1105)) + ((g1031) & (!g1060) & (sk[92]) & (!g1065) & (g1098) & (!g1105)) + ((g1031) & (!g1060) & (sk[92]) & (g1065) & (!g1098) & (!g1105)) + ((g1031) & (!g1060) & (sk[92]) & (g1065) & (g1098) & (g1105)) + ((g1031) & (g1060) & (!sk[92]) & (!g1065) & (!g1098) & (!g1105)) + ((g1031) & (g1060) & (!sk[92]) & (!g1065) & (!g1098) & (g1105)) + ((g1031) & (g1060) & (!sk[92]) & (!g1065) & (g1098) & (!g1105)) + ((g1031) & (g1060) & (!sk[92]) & (!g1065) & (g1098) & (g1105)) + ((g1031) & (g1060) & (!sk[92]) & (g1065) & (!g1098) & (!g1105)) + ((g1031) & (g1060) & (!sk[92]) & (g1065) & (!g1098) & (g1105)) + ((g1031) & (g1060) & (!sk[92]) & (g1065) & (g1098) & (!g1105)) + ((g1031) & (g1060) & (!sk[92]) & (g1065) & (g1098) & (g1105)) + ((g1031) & (g1060) & (sk[92]) & (!g1065) & (!g1098) & (g1105)) + ((g1031) & (g1060) & (sk[92]) & (!g1065) & (g1098) & (!g1105)) + ((g1031) & (g1060) & (sk[92]) & (g1065) & (!g1098) & (g1105)) + ((g1031) & (g1060) & (sk[92]) & (g1065) & (g1098) & (!g1105)));
	assign g1107 = (((!g1067) & (!sk[93]) & (!g1068) & (!g1069) & (g1106)) + ((!g1067) & (!sk[93]) & (!g1068) & (g1069) & (g1106)) + ((!g1067) & (!sk[93]) & (g1068) & (!g1069) & (g1106)) + ((!g1067) & (!sk[93]) & (g1068) & (g1069) & (g1106)) + ((!g1067) & (sk[93]) & (!g1068) & (!g1069) & (!g1106)) + ((!g1067) & (sk[93]) & (!g1068) & (g1069) & (g1106)) + ((!g1067) & (sk[93]) & (g1068) & (!g1069) & (g1106)) + ((!g1067) & (sk[93]) & (g1068) & (g1069) & (!g1106)) + ((g1067) & (!sk[93]) & (!g1068) & (!g1069) & (!g1106)) + ((g1067) & (!sk[93]) & (!g1068) & (!g1069) & (g1106)) + ((g1067) & (!sk[93]) & (!g1068) & (g1069) & (!g1106)) + ((g1067) & (!sk[93]) & (!g1068) & (g1069) & (g1106)) + ((g1067) & (!sk[93]) & (g1068) & (!g1069) & (!g1106)) + ((g1067) & (!sk[93]) & (g1068) & (!g1069) & (g1106)) + ((g1067) & (!sk[93]) & (g1068) & (g1069) & (!g1106)) + ((g1067) & (!sk[93]) & (g1068) & (g1069) & (g1106)) + ((g1067) & (sk[93]) & (!g1068) & (!g1069) & (!g1106)) + ((g1067) & (sk[93]) & (!g1068) & (g1069) & (g1106)) + ((g1067) & (sk[93]) & (g1068) & (!g1069) & (!g1106)) + ((g1067) & (sk[93]) & (g1068) & (g1069) & (g1106)));
	assign g1108 = (((!g975) & (!g990) & (!g997) & (g1043) & (g1059) & (g1097)) + ((!g975) & (!g990) & (g997) & (g1043) & (g1059) & (g1097)) + ((!g975) & (g990) & (!g997) & (!g1043) & (g1059) & (g1097)) + ((!g975) & (g990) & (!g997) & (g1043) & (!g1059) & (g1097)) + ((!g975) & (g990) & (!g997) & (g1043) & (g1059) & (g1097)) + ((!g975) & (g990) & (g997) & (g1043) & (g1059) & (g1097)) + ((g975) & (!g990) & (!g997) & (!g1043) & (g1059) & (g1097)) + ((g975) & (!g990) & (!g997) & (g1043) & (!g1059) & (g1097)) + ((g975) & (!g990) & (!g997) & (g1043) & (g1059) & (g1097)) + ((g975) & (!g990) & (g997) & (g1043) & (g1059) & (g1097)) + ((g975) & (g990) & (!g997) & (!g1043) & (g1059) & (g1097)) + ((g975) & (g990) & (!g997) & (g1043) & (!g1059) & (g1097)) + ((g975) & (g990) & (!g997) & (g1043) & (g1059) & (g1097)) + ((g975) & (g990) & (g997) & (!g1043) & (g1059) & (g1097)) + ((g975) & (g990) & (g997) & (g1043) & (!g1059) & (g1097)) + ((g975) & (g990) & (g997) & (g1043) & (g1059) & (g1097)));
	assign g1109 = (((!g1044) & (!g1055) & (!g1058) & (g1082) & (!g1094) & (!g1096)) + ((!g1044) & (!g1055) & (!g1058) & (g1082) & (g1094) & (g1096)) + ((!g1044) & (!g1055) & (g1058) & (g1082) & (!g1094) & (g1096)) + ((!g1044) & (!g1055) & (g1058) & (g1082) & (g1094) & (!g1096)) + ((!g1044) & (g1055) & (!g1058) & (g1082) & (!g1094) & (g1096)) + ((!g1044) & (g1055) & (!g1058) & (g1082) & (g1094) & (!g1096)) + ((!g1044) & (g1055) & (g1058) & (g1082) & (!g1094) & (g1096)) + ((!g1044) & (g1055) & (g1058) & (g1082) & (g1094) & (!g1096)) + ((g1044) & (!g1055) & (!g1058) & (g1082) & (!g1094) & (!g1096)) + ((g1044) & (!g1055) & (!g1058) & (g1082) & (g1094) & (g1096)) + ((g1044) & (!g1055) & (g1058) & (g1082) & (!g1094) & (!g1096)) + ((g1044) & (!g1055) & (g1058) & (g1082) & (g1094) & (g1096)) + ((g1044) & (g1055) & (!g1058) & (g1082) & (!g1094) & (!g1096)) + ((g1044) & (g1055) & (!g1058) & (g1082) & (g1094) & (g1096)) + ((g1044) & (g1055) & (g1058) & (g1082) & (!g1094) & (g1096)) + ((g1044) & (g1055) & (g1058) & (g1082) & (g1094) & (!g1096)));
	assign g1110 = (((!sk[96]) & (!g864) & (!g892) & (!g1040) & (g1079)) + ((!sk[96]) & (!g864) & (!g892) & (g1040) & (g1079)) + ((!sk[96]) & (!g864) & (g892) & (!g1040) & (g1079)) + ((!sk[96]) & (!g864) & (g892) & (g1040) & (g1079)) + ((!sk[96]) & (g864) & (!g892) & (!g1040) & (!g1079)) + ((!sk[96]) & (g864) & (!g892) & (!g1040) & (g1079)) + ((!sk[96]) & (g864) & (!g892) & (g1040) & (!g1079)) + ((!sk[96]) & (g864) & (!g892) & (g1040) & (g1079)) + ((!sk[96]) & (g864) & (g892) & (!g1040) & (!g1079)) + ((!sk[96]) & (g864) & (g892) & (!g1040) & (g1079)) + ((!sk[96]) & (g864) & (g892) & (g1040) & (!g1079)) + ((!sk[96]) & (g864) & (g892) & (g1040) & (g1079)) + ((sk[96]) & (!g864) & (g892) & (!g1040) & (!g1079)) + ((sk[96]) & (!g864) & (g892) & (g1040) & (!g1079)) + ((sk[96]) & (g864) & (!g892) & (!g1040) & (!g1079)) + ((sk[96]) & (g864) & (!g892) & (!g1040) & (g1079)) + ((sk[96]) & (g864) & (g892) & (!g1040) & (!g1079)) + ((sk[96]) & (g864) & (g892) & (!g1040) & (g1079)) + ((sk[96]) & (g864) & (g892) & (g1040) & (!g1079)));
	assign g1111 = (((!g683) & (!g868) & (!g1040) & (!g1079) & (!g1080) & (g1110)) + ((!g683) & (!g868) & (!g1040) & (!g1079) & (g1080) & (g1110)) + ((!g683) & (!g868) & (!g1040) & (g1079) & (!g1080) & (g1110)) + ((!g683) & (!g868) & (!g1040) & (g1079) & (g1080) & (g1110)) + ((!g683) & (!g868) & (g1040) & (!g1079) & (!g1080) & (g1110)) + ((!g683) & (!g868) & (g1040) & (!g1079) & (g1080) & (g1110)) + ((!g683) & (!g868) & (g1040) & (g1079) & (!g1080) & (g1110)) + ((!g683) & (!g868) & (g1040) & (g1079) & (g1080) & (g1110)) + ((!g683) & (g868) & (!g1040) & (!g1079) & (!g1080) & (g1110)) + ((!g683) & (g868) & (!g1040) & (!g1079) & (g1080) & (g1110)) + ((!g683) & (g868) & (!g1040) & (g1079) & (!g1080) & (g1110)) + ((!g683) & (g868) & (!g1040) & (g1079) & (g1080) & (!g1110)) + ((!g683) & (g868) & (!g1040) & (g1079) & (g1080) & (g1110)) + ((!g683) & (g868) & (g1040) & (!g1079) & (!g1080) & (!g1110)) + ((!g683) & (g868) & (g1040) & (!g1079) & (!g1080) & (g1110)) + ((!g683) & (g868) & (g1040) & (!g1079) & (g1080) & (g1110)) + ((!g683) & (g868) & (g1040) & (g1079) & (!g1080) & (g1110)) + ((!g683) & (g868) & (g1040) & (g1079) & (g1080) & (g1110)) + ((g683) & (!g868) & (!g1040) & (!g1079) & (!g1080) & (!g1110)) + ((g683) & (!g868) & (!g1040) & (!g1079) & (g1080) & (!g1110)) + ((g683) & (!g868) & (!g1040) & (g1079) & (!g1080) & (!g1110)) + ((g683) & (!g868) & (!g1040) & (g1079) & (g1080) & (!g1110)) + ((g683) & (!g868) & (g1040) & (!g1079) & (!g1080) & (!g1110)) + ((g683) & (!g868) & (g1040) & (!g1079) & (g1080) & (!g1110)) + ((g683) & (!g868) & (g1040) & (g1079) & (!g1080) & (!g1110)) + ((g683) & (!g868) & (g1040) & (g1079) & (g1080) & (!g1110)) + ((g683) & (g868) & (!g1040) & (!g1079) & (!g1080) & (!g1110)) + ((g683) & (g868) & (!g1040) & (!g1079) & (g1080) & (!g1110)) + ((g683) & (g868) & (!g1040) & (g1079) & (!g1080) & (!g1110)) + ((g683) & (g868) & (g1040) & (!g1079) & (g1080) & (!g1110)) + ((g683) & (g868) & (g1040) & (g1079) & (!g1080) & (!g1110)) + ((g683) & (g868) & (g1040) & (g1079) & (g1080) & (!g1110)));
	assign g1112 = (((!g1044) & (!g1055) & (!g1058) & (!sk[98]) & (g1094) & (!g1096)) + ((!g1044) & (!g1055) & (!g1058) & (!sk[98]) & (g1094) & (g1096)) + ((!g1044) & (!g1055) & (!g1058) & (sk[98]) & (!g1094) & (!g1096)) + ((!g1044) & (!g1055) & (!g1058) & (sk[98]) & (!g1094) & (g1096)) + ((!g1044) & (!g1055) & (!g1058) & (sk[98]) & (g1094) & (!g1096)) + ((!g1044) & (!g1055) & (g1058) & (!sk[98]) & (!g1094) & (!g1096)) + ((!g1044) & (!g1055) & (g1058) & (!sk[98]) & (!g1094) & (g1096)) + ((!g1044) & (!g1055) & (g1058) & (!sk[98]) & (g1094) & (!g1096)) + ((!g1044) & (!g1055) & (g1058) & (!sk[98]) & (g1094) & (g1096)) + ((!g1044) & (!g1055) & (g1058) & (sk[98]) & (!g1094) & (!g1096)) + ((!g1044) & (g1055) & (!g1058) & (!sk[98]) & (!g1094) & (!g1096)) + ((!g1044) & (g1055) & (!g1058) & (!sk[98]) & (!g1094) & (g1096)) + ((!g1044) & (g1055) & (!g1058) & (!sk[98]) & (g1094) & (!g1096)) + ((!g1044) & (g1055) & (!g1058) & (!sk[98]) & (g1094) & (g1096)) + ((!g1044) & (g1055) & (!g1058) & (sk[98]) & (!g1094) & (!g1096)) + ((!g1044) & (g1055) & (g1058) & (!sk[98]) & (!g1094) & (!g1096)) + ((!g1044) & (g1055) & (g1058) & (!sk[98]) & (!g1094) & (g1096)) + ((!g1044) & (g1055) & (g1058) & (!sk[98]) & (g1094) & (!g1096)) + ((!g1044) & (g1055) & (g1058) & (!sk[98]) & (g1094) & (g1096)) + ((!g1044) & (g1055) & (g1058) & (sk[98]) & (!g1094) & (!g1096)) + ((g1044) & (!g1055) & (!g1058) & (!sk[98]) & (g1094) & (!g1096)) + ((g1044) & (!g1055) & (!g1058) & (!sk[98]) & (g1094) & (g1096)) + ((g1044) & (!g1055) & (!g1058) & (sk[98]) & (!g1094) & (!g1096)) + ((g1044) & (!g1055) & (!g1058) & (sk[98]) & (!g1094) & (g1096)) + ((g1044) & (!g1055) & (!g1058) & (sk[98]) & (g1094) & (!g1096)) + ((g1044) & (!g1055) & (g1058) & (!sk[98]) & (!g1094) & (!g1096)) + ((g1044) & (!g1055) & (g1058) & (!sk[98]) & (!g1094) & (g1096)) + ((g1044) & (!g1055) & (g1058) & (!sk[98]) & (g1094) & (!g1096)) + ((g1044) & (!g1055) & (g1058) & (!sk[98]) & (g1094) & (g1096)) + ((g1044) & (!g1055) & (g1058) & (sk[98]) & (!g1094) & (!g1096)) + ((g1044) & (!g1055) & (g1058) & (sk[98]) & (!g1094) & (g1096)) + ((g1044) & (!g1055) & (g1058) & (sk[98]) & (g1094) & (!g1096)) + ((g1044) & (g1055) & (!g1058) & (!sk[98]) & (!g1094) & (!g1096)) + ((g1044) & (g1055) & (!g1058) & (!sk[98]) & (!g1094) & (g1096)) + ((g1044) & (g1055) & (!g1058) & (!sk[98]) & (g1094) & (!g1096)) + ((g1044) & (g1055) & (!g1058) & (!sk[98]) & (g1094) & (g1096)) + ((g1044) & (g1055) & (!g1058) & (sk[98]) & (!g1094) & (!g1096)) + ((g1044) & (g1055) & (!g1058) & (sk[98]) & (!g1094) & (g1096)) + ((g1044) & (g1055) & (!g1058) & (sk[98]) & (g1094) & (!g1096)) + ((g1044) & (g1055) & (g1058) & (!sk[98]) & (!g1094) & (!g1096)) + ((g1044) & (g1055) & (g1058) & (!sk[98]) & (!g1094) & (g1096)) + ((g1044) & (g1055) & (g1058) & (!sk[98]) & (g1094) & (!g1096)) + ((g1044) & (g1055) & (g1058) & (!sk[98]) & (g1094) & (g1096)) + ((g1044) & (g1055) & (g1058) & (sk[98]) & (!g1094) & (!g1096)));
	assign g1113 = (((!g747) & (!g748) & (!sk[99]) & (!g870) & (g871) & (!g883)) + ((!g747) & (!g748) & (!sk[99]) & (!g870) & (g871) & (g883)) + ((!g747) & (!g748) & (!sk[99]) & (g870) & (!g871) & (!g883)) + ((!g747) & (!g748) & (!sk[99]) & (g870) & (!g871) & (g883)) + ((!g747) & (!g748) & (!sk[99]) & (g870) & (g871) & (!g883)) + ((!g747) & (!g748) & (!sk[99]) & (g870) & (g871) & (g883)) + ((!g747) & (g748) & (!sk[99]) & (!g870) & (!g871) & (!g883)) + ((!g747) & (g748) & (!sk[99]) & (!g870) & (!g871) & (g883)) + ((!g747) & (g748) & (!sk[99]) & (!g870) & (g871) & (!g883)) + ((!g747) & (g748) & (!sk[99]) & (!g870) & (g871) & (g883)) + ((!g747) & (g748) & (!sk[99]) & (g870) & (!g871) & (!g883)) + ((!g747) & (g748) & (!sk[99]) & (g870) & (!g871) & (g883)) + ((!g747) & (g748) & (!sk[99]) & (g870) & (g871) & (!g883)) + ((!g747) & (g748) & (!sk[99]) & (g870) & (g871) & (g883)) + ((!g747) & (g748) & (sk[99]) & (!g870) & (!g871) & (!g883)) + ((!g747) & (g748) & (sk[99]) & (!g870) & (!g871) & (g883)) + ((!g747) & (g748) & (sk[99]) & (!g870) & (g871) & (!g883)) + ((!g747) & (g748) & (sk[99]) & (!g870) & (g871) & (g883)) + ((g747) & (!g748) & (!sk[99]) & (!g870) & (g871) & (!g883)) + ((g747) & (!g748) & (!sk[99]) & (!g870) & (g871) & (g883)) + ((g747) & (!g748) & (!sk[99]) & (g870) & (!g871) & (!g883)) + ((g747) & (!g748) & (!sk[99]) & (g870) & (!g871) & (g883)) + ((g747) & (!g748) & (!sk[99]) & (g870) & (g871) & (!g883)) + ((g747) & (!g748) & (!sk[99]) & (g870) & (g871) & (g883)) + ((g747) & (!g748) & (sk[99]) & (!g870) & (!g871) & (!g883)) + ((g747) & (!g748) & (sk[99]) & (!g870) & (g871) & (g883)) + ((g747) & (!g748) & (sk[99]) & (g870) & (!g871) & (!g883)) + ((g747) & (!g748) & (sk[99]) & (g870) & (g871) & (g883)) + ((g747) & (g748) & (!sk[99]) & (!g870) & (!g871) & (!g883)) + ((g747) & (g748) & (!sk[99]) & (!g870) & (!g871) & (g883)) + ((g747) & (g748) & (!sk[99]) & (!g870) & (g871) & (!g883)) + ((g747) & (g748) & (!sk[99]) & (!g870) & (g871) & (g883)) + ((g747) & (g748) & (!sk[99]) & (g870) & (!g871) & (!g883)) + ((g747) & (g748) & (!sk[99]) & (g870) & (!g871) & (g883)) + ((g747) & (g748) & (!sk[99]) & (g870) & (g871) & (!g883)) + ((g747) & (g748) & (!sk[99]) & (g870) & (g871) & (g883)) + ((g747) & (g748) & (sk[99]) & (!g870) & (!g871) & (!g883)) + ((g747) & (g748) & (sk[99]) & (!g870) & (!g871) & (g883)) + ((g747) & (g748) & (sk[99]) & (!g870) & (g871) & (!g883)) + ((g747) & (g748) & (sk[99]) & (!g870) & (g871) & (g883)) + ((g747) & (g748) & (sk[99]) & (g870) & (!g871) & (!g883)) + ((g747) & (g748) & (sk[99]) & (g870) & (g871) & (g883)));
	assign g1114 = (((!g200) & (!g742) & (!g744) & (!g863) & (!g895) & (g1113)) + ((!g200) & (!g742) & (!g744) & (!g863) & (g895) & (g1113)) + ((!g200) & (!g742) & (!g744) & (g863) & (!g895) & (g1113)) + ((!g200) & (!g742) & (!g744) & (g863) & (g895) & (g1113)) + ((!g200) & (!g742) & (g744) & (!g863) & (!g895) & (g1113)) + ((!g200) & (!g742) & (g744) & (!g863) & (g895) & (g1113)) + ((!g200) & (!g742) & (g744) & (g863) & (!g895) & (!g1113)) + ((!g200) & (!g742) & (g744) & (g863) & (!g895) & (g1113)) + ((!g200) & (!g742) & (g744) & (g863) & (g895) & (!g1113)) + ((!g200) & (!g742) & (g744) & (g863) & (g895) & (g1113)) + ((!g200) & (g742) & (!g744) & (!g863) & (!g895) & (g1113)) + ((!g200) & (g742) & (!g744) & (!g863) & (g895) & (!g1113)) + ((!g200) & (g742) & (!g744) & (!g863) & (g895) & (g1113)) + ((!g200) & (g742) & (!g744) & (g863) & (!g895) & (g1113)) + ((!g200) & (g742) & (!g744) & (g863) & (g895) & (!g1113)) + ((!g200) & (g742) & (!g744) & (g863) & (g895) & (g1113)) + ((!g200) & (g742) & (g744) & (!g863) & (!g895) & (g1113)) + ((!g200) & (g742) & (g744) & (!g863) & (g895) & (!g1113)) + ((!g200) & (g742) & (g744) & (!g863) & (g895) & (g1113)) + ((!g200) & (g742) & (g744) & (g863) & (!g895) & (!g1113)) + ((!g200) & (g742) & (g744) & (g863) & (!g895) & (g1113)) + ((!g200) & (g742) & (g744) & (g863) & (g895) & (!g1113)) + ((!g200) & (g742) & (g744) & (g863) & (g895) & (g1113)) + ((g200) & (!g742) & (!g744) & (!g863) & (!g895) & (!g1113)) + ((g200) & (!g742) & (!g744) & (!g863) & (g895) & (!g1113)) + ((g200) & (!g742) & (!g744) & (g863) & (!g895) & (!g1113)) + ((g200) & (!g742) & (!g744) & (g863) & (g895) & (!g1113)) + ((g200) & (!g742) & (g744) & (!g863) & (!g895) & (!g1113)) + ((g200) & (!g742) & (g744) & (!g863) & (g895) & (!g1113)) + ((g200) & (g742) & (!g744) & (!g863) & (!g895) & (!g1113)) + ((g200) & (g742) & (!g744) & (g863) & (!g895) & (!g1113)) + ((g200) & (g742) & (g744) & (!g863) & (!g895) & (!g1113)));
	assign g1115 = (((!g202) & (!g1048) & (!g1051) & (!g1053) & (!g1088) & (g1092)) + ((!g202) & (!g1048) & (!g1051) & (g1053) & (!g1088) & (g1092)) + ((!g202) & (!g1048) & (g1051) & (!g1053) & (!g1088) & (!g1092)) + ((!g202) & (!g1048) & (g1051) & (!g1053) & (!g1088) & (g1092)) + ((!g202) & (!g1048) & (g1051) & (!g1053) & (g1088) & (g1092)) + ((!g202) & (!g1048) & (g1051) & (g1053) & (!g1088) & (g1092)) + ((!g202) & (g1048) & (!g1051) & (!g1053) & (!g1088) & (!g1092)) + ((!g202) & (g1048) & (!g1051) & (!g1053) & (!g1088) & (g1092)) + ((!g202) & (g1048) & (!g1051) & (!g1053) & (g1088) & (g1092)) + ((!g202) & (g1048) & (!g1051) & (g1053) & (!g1088) & (g1092)) + ((!g202) & (g1048) & (g1051) & (!g1053) & (!g1088) & (!g1092)) + ((!g202) & (g1048) & (g1051) & (!g1053) & (!g1088) & (g1092)) + ((!g202) & (g1048) & (g1051) & (!g1053) & (g1088) & (g1092)) + ((!g202) & (g1048) & (g1051) & (g1053) & (!g1088) & (!g1092)) + ((!g202) & (g1048) & (g1051) & (g1053) & (!g1088) & (g1092)) + ((!g202) & (g1048) & (g1051) & (g1053) & (g1088) & (g1092)) + ((g202) & (!g1048) & (!g1051) & (!g1053) & (g1088) & (g1092)) + ((g202) & (!g1048) & (!g1051) & (g1053) & (g1088) & (g1092)) + ((g202) & (!g1048) & (g1051) & (!g1053) & (!g1088) & (g1092)) + ((g202) & (!g1048) & (g1051) & (!g1053) & (g1088) & (!g1092)) + ((g202) & (!g1048) & (g1051) & (!g1053) & (g1088) & (g1092)) + ((g202) & (!g1048) & (g1051) & (g1053) & (g1088) & (g1092)) + ((g202) & (g1048) & (!g1051) & (!g1053) & (!g1088) & (g1092)) + ((g202) & (g1048) & (!g1051) & (!g1053) & (g1088) & (!g1092)) + ((g202) & (g1048) & (!g1051) & (!g1053) & (g1088) & (g1092)) + ((g202) & (g1048) & (!g1051) & (g1053) & (g1088) & (g1092)) + ((g202) & (g1048) & (g1051) & (!g1053) & (!g1088) & (g1092)) + ((g202) & (g1048) & (g1051) & (!g1053) & (g1088) & (!g1092)) + ((g202) & (g1048) & (g1051) & (!g1053) & (g1088) & (g1092)) + ((g202) & (g1048) & (g1051) & (g1053) & (!g1088) & (g1092)) + ((g202) & (g1048) & (g1051) & (g1053) & (g1088) & (!g1092)) + ((g202) & (g1048) & (g1051) & (g1053) & (g1088) & (g1092)));
	assign g1116 = (((!g707) & (!g717) & (!sk[102]) & (!g718) & (g764) & (!g762)) + ((!g707) & (!g717) & (!sk[102]) & (!g718) & (g764) & (g762)) + ((!g707) & (!g717) & (!sk[102]) & (g718) & (!g764) & (!g762)) + ((!g707) & (!g717) & (!sk[102]) & (g718) & (!g764) & (g762)) + ((!g707) & (!g717) & (!sk[102]) & (g718) & (g764) & (!g762)) + ((!g707) & (!g717) & (!sk[102]) & (g718) & (g764) & (g762)) + ((!g707) & (!g717) & (sk[102]) & (g718) & (!g764) & (g762)) + ((!g707) & (!g717) & (sk[102]) & (g718) & (g764) & (g762)) + ((!g707) & (g717) & (!sk[102]) & (!g718) & (!g764) & (!g762)) + ((!g707) & (g717) & (!sk[102]) & (!g718) & (!g764) & (g762)) + ((!g707) & (g717) & (!sk[102]) & (!g718) & (g764) & (!g762)) + ((!g707) & (g717) & (!sk[102]) & (!g718) & (g764) & (g762)) + ((!g707) & (g717) & (!sk[102]) & (g718) & (!g764) & (!g762)) + ((!g707) & (g717) & (!sk[102]) & (g718) & (!g764) & (g762)) + ((!g707) & (g717) & (!sk[102]) & (g718) & (g764) & (!g762)) + ((!g707) & (g717) & (!sk[102]) & (g718) & (g764) & (g762)) + ((!g707) & (g717) & (sk[102]) & (!g718) & (g764) & (!g762)) + ((!g707) & (g717) & (sk[102]) & (!g718) & (g764) & (g762)) + ((!g707) & (g717) & (sk[102]) & (g718) & (!g764) & (g762)) + ((!g707) & (g717) & (sk[102]) & (g718) & (g764) & (!g762)) + ((!g707) & (g717) & (sk[102]) & (g718) & (g764) & (g762)) + ((g707) & (!g717) & (!sk[102]) & (!g718) & (g764) & (!g762)) + ((g707) & (!g717) & (!sk[102]) & (!g718) & (g764) & (g762)) + ((g707) & (!g717) & (!sk[102]) & (g718) & (!g764) & (!g762)) + ((g707) & (!g717) & (!sk[102]) & (g718) & (!g764) & (g762)) + ((g707) & (!g717) & (!sk[102]) & (g718) & (g764) & (!g762)) + ((g707) & (!g717) & (!sk[102]) & (g718) & (g764) & (g762)) + ((g707) & (!g717) & (sk[102]) & (!g718) & (g764) & (!g762)) + ((g707) & (!g717) & (sk[102]) & (!g718) & (g764) & (g762)) + ((g707) & (!g717) & (sk[102]) & (g718) & (!g764) & (g762)) + ((g707) & (!g717) & (sk[102]) & (g718) & (g764) & (!g762)) + ((g707) & (!g717) & (sk[102]) & (g718) & (g764) & (g762)) + ((g707) & (g717) & (!sk[102]) & (!g718) & (!g764) & (!g762)) + ((g707) & (g717) & (!sk[102]) & (!g718) & (!g764) & (g762)) + ((g707) & (g717) & (!sk[102]) & (!g718) & (g764) & (!g762)) + ((g707) & (g717) & (!sk[102]) & (!g718) & (g764) & (g762)) + ((g707) & (g717) & (!sk[102]) & (g718) & (!g764) & (!g762)) + ((g707) & (g717) & (!sk[102]) & (g718) & (!g764) & (g762)) + ((g707) & (g717) & (!sk[102]) & (g718) & (g764) & (!g762)) + ((g707) & (g717) & (!sk[102]) & (g718) & (g764) & (g762)) + ((g707) & (g717) & (sk[102]) & (g718) & (!g764) & (g762)) + ((g707) & (g717) & (sk[102]) & (g718) & (g764) & (g762)));
	assign g1117 = (((!g202) & (!g681) & (!g731) & (!g759) & (!g765) & (!g1116)) + ((!g202) & (!g681) & (!g731) & (g759) & (!g765) & (!g1116)) + ((!g202) & (!g681) & (g731) & (!g759) & (!g765) & (!g1116)) + ((!g202) & (g681) & (!g731) & (!g759) & (!g765) & (!g1116)) + ((!g202) & (g681) & (!g731) & (!g759) & (g765) & (!g1116)) + ((!g202) & (g681) & (!g731) & (g759) & (!g765) & (!g1116)) + ((!g202) & (g681) & (!g731) & (g759) & (g765) & (!g1116)) + ((!g202) & (g681) & (g731) & (!g759) & (!g765) & (!g1116)) + ((!g202) & (g681) & (g731) & (!g759) & (g765) & (!g1116)) + ((g202) & (!g681) & (!g731) & (!g759) & (!g765) & (g1116)) + ((g202) & (!g681) & (!g731) & (!g759) & (g765) & (!g1116)) + ((g202) & (!g681) & (!g731) & (!g759) & (g765) & (g1116)) + ((g202) & (!g681) & (!g731) & (g759) & (!g765) & (g1116)) + ((g202) & (!g681) & (!g731) & (g759) & (g765) & (!g1116)) + ((g202) & (!g681) & (!g731) & (g759) & (g765) & (g1116)) + ((g202) & (!g681) & (g731) & (!g759) & (!g765) & (g1116)) + ((g202) & (!g681) & (g731) & (!g759) & (g765) & (!g1116)) + ((g202) & (!g681) & (g731) & (!g759) & (g765) & (g1116)) + ((g202) & (!g681) & (g731) & (g759) & (!g765) & (!g1116)) + ((g202) & (!g681) & (g731) & (g759) & (!g765) & (g1116)) + ((g202) & (!g681) & (g731) & (g759) & (g765) & (!g1116)) + ((g202) & (!g681) & (g731) & (g759) & (g765) & (g1116)) + ((g202) & (g681) & (!g731) & (!g759) & (!g765) & (g1116)) + ((g202) & (g681) & (!g731) & (!g759) & (g765) & (g1116)) + ((g202) & (g681) & (!g731) & (g759) & (!g765) & (g1116)) + ((g202) & (g681) & (!g731) & (g759) & (g765) & (g1116)) + ((g202) & (g681) & (g731) & (!g759) & (!g765) & (g1116)) + ((g202) & (g681) & (g731) & (!g759) & (g765) & (g1116)) + ((g202) & (g681) & (g731) & (g759) & (!g765) & (!g1116)) + ((g202) & (g681) & (g731) & (g759) & (!g765) & (g1116)) + ((g202) & (g681) & (g731) & (g759) & (g765) & (!g1116)) + ((g202) & (g681) & (g731) & (g759) & (g765) & (g1116)));
	assign g1118 = (((!g585) & (!g597) & (!g679) & (g720) & (!g845) & (g848)) + ((!g585) & (!g597) & (!g679) & (g720) & (g845) & (g848)) + ((!g585) & (!g597) & (g679) & (!g720) & (g845) & (!g848)) + ((!g585) & (!g597) & (g679) & (!g720) & (g845) & (g848)) + ((!g585) & (!g597) & (g679) & (g720) & (!g845) & (g848)) + ((!g585) & (!g597) & (g679) & (g720) & (g845) & (!g848)) + ((!g585) & (!g597) & (g679) & (g720) & (g845) & (g848)) + ((!g585) & (g597) & (!g679) & (!g720) & (g845) & (!g848)) + ((!g585) & (g597) & (!g679) & (!g720) & (g845) & (g848)) + ((!g585) & (g597) & (!g679) & (g720) & (!g845) & (g848)) + ((!g585) & (g597) & (!g679) & (g720) & (g845) & (!g848)) + ((!g585) & (g597) & (!g679) & (g720) & (g845) & (g848)) + ((!g585) & (g597) & (g679) & (g720) & (!g845) & (g848)) + ((!g585) & (g597) & (g679) & (g720) & (g845) & (g848)) + ((g585) & (!g597) & (!g679) & (!g720) & (g845) & (!g848)) + ((g585) & (!g597) & (!g679) & (!g720) & (g845) & (g848)) + ((g585) & (!g597) & (!g679) & (g720) & (!g845) & (g848)) + ((g585) & (!g597) & (!g679) & (g720) & (g845) & (!g848)) + ((g585) & (!g597) & (!g679) & (g720) & (g845) & (g848)) + ((g585) & (!g597) & (g679) & (g720) & (!g845) & (g848)) + ((g585) & (!g597) & (g679) & (g720) & (g845) & (g848)) + ((g585) & (g597) & (!g679) & (g720) & (!g845) & (g848)) + ((g585) & (g597) & (!g679) & (g720) & (g845) & (g848)) + ((g585) & (g597) & (g679) & (!g720) & (g845) & (!g848)) + ((g585) & (g597) & (g679) & (!g720) & (g845) & (g848)) + ((g585) & (g597) & (g679) & (g720) & (!g845) & (g848)) + ((g585) & (g597) & (g679) & (g720) & (g845) & (!g848)) + ((g585) & (g597) & (g679) & (g720) & (g845) & (g848)));
	assign g1119 = (((!g719) & (!g728) & (!g729) & (!g847) & (!g843) & (!g1118)) + ((!g719) & (!g728) & (!g729) & (!g847) & (g843) & (!g1118)) + ((!g719) & (!g728) & (g729) & (!g847) & (!g843) & (!g1118)) + ((!g719) & (!g728) & (g729) & (g847) & (!g843) & (!g1118)) + ((!g719) & (g728) & (!g729) & (!g847) & (!g843) & (!g1118)) + ((!g719) & (g728) & (g729) & (!g847) & (!g843) & (!g1118)) + ((!g719) & (g728) & (g729) & (!g847) & (g843) & (!g1118)) + ((!g719) & (g728) & (g729) & (g847) & (!g843) & (!g1118)) + ((!g719) & (g728) & (g729) & (g847) & (g843) & (!g1118)) + ((g719) & (!g728) & (!g729) & (!g847) & (!g843) & (!g1118)) + ((g719) & (!g728) & (g729) & (!g847) & (!g843) & (!g1118)) + ((g719) & (!g728) & (g729) & (!g847) & (g843) & (!g1118)) + ((g719) & (!g728) & (g729) & (g847) & (!g843) & (!g1118)) + ((g719) & (!g728) & (g729) & (g847) & (g843) & (!g1118)) + ((g719) & (g728) & (!g729) & (!g847) & (!g843) & (!g1118)) + ((g719) & (g728) & (!g729) & (!g847) & (g843) & (!g1118)) + ((g719) & (g728) & (g729) & (!g847) & (!g843) & (!g1118)) + ((g719) & (g728) & (g729) & (g847) & (!g843) & (!g1118)));
	assign g1120 = (((!g252) & (!g722) & (!g723) & (!g1089) & (!g1091) & (!g1119)) + ((!g252) & (!g722) & (!g723) & (!g1089) & (g1091) & (!g1119)) + ((!g252) & (!g722) & (!g723) & (g1089) & (!g1091) & (g1119)) + ((!g252) & (!g722) & (!g723) & (g1089) & (g1091) & (!g1119)) + ((!g252) & (!g722) & (g723) & (!g1089) & (!g1091) & (!g1119)) + ((!g252) & (!g722) & (g723) & (!g1089) & (g1091) & (!g1119)) + ((!g252) & (!g722) & (g723) & (g1089) & (!g1091) & (g1119)) + ((!g252) & (!g722) & (g723) & (g1089) & (g1091) & (!g1119)) + ((!g252) & (g722) & (!g723) & (!g1089) & (!g1091) & (!g1119)) + ((!g252) & (g722) & (!g723) & (!g1089) & (g1091) & (!g1119)) + ((!g252) & (g722) & (!g723) & (g1089) & (!g1091) & (g1119)) + ((!g252) & (g722) & (!g723) & (g1089) & (g1091) & (!g1119)) + ((!g252) & (g722) & (g723) & (!g1089) & (!g1091) & (!g1119)) + ((!g252) & (g722) & (g723) & (!g1089) & (g1091) & (!g1119)) + ((!g252) & (g722) & (g723) & (g1089) & (!g1091) & (g1119)) + ((!g252) & (g722) & (g723) & (g1089) & (g1091) & (!g1119)) + ((g252) & (!g722) & (!g723) & (!g1089) & (!g1091) & (!g1119)) + ((g252) & (!g722) & (!g723) & (!g1089) & (g1091) & (g1119)) + ((g252) & (!g722) & (!g723) & (g1089) & (!g1091) & (g1119)) + ((g252) & (!g722) & (!g723) & (g1089) & (g1091) & (g1119)) + ((g252) & (!g722) & (g723) & (!g1089) & (!g1091) & (!g1119)) + ((g252) & (!g722) & (g723) & (!g1089) & (g1091) & (!g1119)) + ((g252) & (!g722) & (g723) & (g1089) & (!g1091) & (!g1119)) + ((g252) & (!g722) & (g723) & (g1089) & (g1091) & (g1119)) + ((g252) & (g722) & (!g723) & (!g1089) & (!g1091) & (g1119)) + ((g252) & (g722) & (!g723) & (!g1089) & (g1091) & (!g1119)) + ((g252) & (g722) & (!g723) & (g1089) & (!g1091) & (!g1119)) + ((g252) & (g722) & (!g723) & (g1089) & (g1091) & (!g1119)) + ((g252) & (g722) & (g723) & (!g1089) & (!g1091) & (g1119)) + ((g252) & (g722) & (g723) & (!g1089) & (g1091) & (g1119)) + ((g252) & (g722) & (g723) & (g1089) & (!g1091) & (g1119)) + ((g252) & (g722) & (g723) & (g1089) & (g1091) & (!g1119)));
	assign g1121 = (((!sk[107]) & (!g1115) & (g1117) & (!g1120)) + ((!sk[107]) & (!g1115) & (g1117) & (g1120)) + ((!sk[107]) & (g1115) & (g1117) & (!g1120)) + ((!sk[107]) & (g1115) & (g1117) & (g1120)) + ((sk[107]) & (!g1115) & (!g1117) & (g1120)) + ((sk[107]) & (!g1115) & (g1117) & (!g1120)) + ((sk[107]) & (g1115) & (!g1117) & (!g1120)) + ((sk[107]) & (g1115) & (g1117) & (g1120)));
	assign g1122 = (((!g1083) & (!g1085) & (!g1086) & (!g1093) & (!g1114) & (g1121)) + ((!g1083) & (!g1085) & (!g1086) & (!g1093) & (g1114) & (!g1121)) + ((!g1083) & (!g1085) & (!g1086) & (g1093) & (!g1114) & (g1121)) + ((!g1083) & (!g1085) & (!g1086) & (g1093) & (g1114) & (!g1121)) + ((!g1083) & (!g1085) & (g1086) & (!g1093) & (!g1114) & (g1121)) + ((!g1083) & (!g1085) & (g1086) & (!g1093) & (g1114) & (!g1121)) + ((!g1083) & (!g1085) & (g1086) & (g1093) & (!g1114) & (g1121)) + ((!g1083) & (!g1085) & (g1086) & (g1093) & (g1114) & (!g1121)) + ((!g1083) & (g1085) & (!g1086) & (!g1093) & (!g1114) & (!g1121)) + ((!g1083) & (g1085) & (!g1086) & (!g1093) & (g1114) & (g1121)) + ((!g1083) & (g1085) & (!g1086) & (g1093) & (!g1114) & (g1121)) + ((!g1083) & (g1085) & (!g1086) & (g1093) & (g1114) & (!g1121)) + ((!g1083) & (g1085) & (g1086) & (!g1093) & (!g1114) & (g1121)) + ((!g1083) & (g1085) & (g1086) & (!g1093) & (g1114) & (!g1121)) + ((!g1083) & (g1085) & (g1086) & (g1093) & (!g1114) & (!g1121)) + ((!g1083) & (g1085) & (g1086) & (g1093) & (g1114) & (g1121)) + ((g1083) & (!g1085) & (!g1086) & (!g1093) & (!g1114) & (!g1121)) + ((g1083) & (!g1085) & (!g1086) & (!g1093) & (g1114) & (g1121)) + ((g1083) & (!g1085) & (!g1086) & (g1093) & (!g1114) & (g1121)) + ((g1083) & (!g1085) & (!g1086) & (g1093) & (g1114) & (!g1121)) + ((g1083) & (!g1085) & (g1086) & (!g1093) & (!g1114) & (g1121)) + ((g1083) & (!g1085) & (g1086) & (!g1093) & (g1114) & (!g1121)) + ((g1083) & (!g1085) & (g1086) & (g1093) & (!g1114) & (!g1121)) + ((g1083) & (!g1085) & (g1086) & (g1093) & (g1114) & (g1121)) + ((g1083) & (g1085) & (!g1086) & (!g1093) & (!g1114) & (!g1121)) + ((g1083) & (g1085) & (!g1086) & (!g1093) & (g1114) & (g1121)) + ((g1083) & (g1085) & (!g1086) & (g1093) & (!g1114) & (!g1121)) + ((g1083) & (g1085) & (!g1086) & (g1093) & (g1114) & (g1121)) + ((g1083) & (g1085) & (g1086) & (!g1093) & (!g1114) & (!g1121)) + ((g1083) & (g1085) & (g1086) & (!g1093) & (g1114) & (g1121)) + ((g1083) & (g1085) & (g1086) & (g1093) & (!g1114) & (!g1121)) + ((g1083) & (g1085) & (g1086) & (g1093) & (g1114) & (g1121)));
	assign g1123 = (((!g733) & (!g686) & (!g734) & (!g962) & (!g971) & (!g994)) + ((!g733) & (!g686) & (!g734) & (!g962) & (!g971) & (g994)) + ((!g733) & (!g686) & (!g734) & (!g962) & (g971) & (!g994)) + ((!g733) & (!g686) & (!g734) & (!g962) & (g971) & (g994)) + ((!g733) & (!g686) & (!g734) & (g962) & (!g971) & (!g994)) + ((!g733) & (!g686) & (!g734) & (g962) & (!g971) & (g994)) + ((!g733) & (!g686) & (!g734) & (g962) & (g971) & (!g994)) + ((!g733) & (!g686) & (!g734) & (g962) & (g971) & (g994)) + ((!g733) & (!g686) & (g734) & (!g962) & (!g971) & (!g994)) + ((!g733) & (!g686) & (g734) & (!g962) & (!g971) & (g994)) + ((!g733) & (!g686) & (g734) & (g962) & (!g971) & (!g994)) + ((!g733) & (!g686) & (g734) & (g962) & (!g971) & (g994)) + ((!g733) & (g686) & (!g734) & (g962) & (!g971) & (!g994)) + ((!g733) & (g686) & (!g734) & (g962) & (!g971) & (g994)) + ((!g733) & (g686) & (!g734) & (g962) & (g971) & (!g994)) + ((!g733) & (g686) & (!g734) & (g962) & (g971) & (g994)) + ((!g733) & (g686) & (g734) & (g962) & (!g971) & (!g994)) + ((!g733) & (g686) & (g734) & (g962) & (!g971) & (g994)) + ((g733) & (!g686) & (!g734) & (!g962) & (!g971) & (!g994)) + ((g733) & (!g686) & (!g734) & (!g962) & (g971) & (!g994)) + ((g733) & (!g686) & (!g734) & (g962) & (!g971) & (!g994)) + ((g733) & (!g686) & (!g734) & (g962) & (g971) & (!g994)) + ((g733) & (!g686) & (g734) & (!g962) & (!g971) & (!g994)) + ((g733) & (!g686) & (g734) & (g962) & (!g971) & (!g994)) + ((g733) & (g686) & (!g734) & (g962) & (!g971) & (!g994)) + ((g733) & (g686) & (!g734) & (g962) & (g971) & (!g994)) + ((g733) & (g686) & (g734) & (g962) & (!g971) & (!g994)));
	assign g1124 = (((!sk[110]) & (!g2) & (!g732) & (!g995) & (g1123)) + ((!sk[110]) & (!g2) & (!g732) & (g995) & (g1123)) + ((!sk[110]) & (!g2) & (g732) & (!g995) & (g1123)) + ((!sk[110]) & (!g2) & (g732) & (g995) & (g1123)) + ((!sk[110]) & (g2) & (!g732) & (!g995) & (!g1123)) + ((!sk[110]) & (g2) & (!g732) & (!g995) & (g1123)) + ((!sk[110]) & (g2) & (!g732) & (g995) & (!g1123)) + ((!sk[110]) & (g2) & (!g732) & (g995) & (g1123)) + ((!sk[110]) & (g2) & (g732) & (!g995) & (!g1123)) + ((!sk[110]) & (g2) & (g732) & (!g995) & (g1123)) + ((!sk[110]) & (g2) & (g732) & (g995) & (!g1123)) + ((!sk[110]) & (g2) & (g732) & (g995) & (g1123)) + ((sk[110]) & (!g2) & (!g732) & (!g995) & (g1123)) + ((sk[110]) & (!g2) & (!g732) & (g995) & (g1123)) + ((sk[110]) & (!g2) & (g732) & (!g995) & (g1123)) + ((sk[110]) & (g2) & (!g732) & (!g995) & (!g1123)) + ((sk[110]) & (g2) & (!g732) & (g995) & (!g1123)) + ((sk[110]) & (g2) & (g732) & (!g995) & (!g1123)) + ((sk[110]) & (g2) & (g732) & (g995) & (!g1123)) + ((sk[110]) & (g2) & (g732) & (g995) & (g1123)));
	assign g1125 = (((!g1112) & (!g1122) & (sk[111]) & (g1124)) + ((!g1112) & (g1122) & (!sk[111]) & (!g1124)) + ((!g1112) & (g1122) & (!sk[111]) & (g1124)) + ((!g1112) & (g1122) & (sk[111]) & (!g1124)) + ((g1112) & (!g1122) & (sk[111]) & (!g1124)) + ((g1112) & (g1122) & (!sk[111]) & (!g1124)) + ((g1112) & (g1122) & (!sk[111]) & (g1124)) + ((g1112) & (g1122) & (sk[111]) & (g1124)));
	assign g1126 = (((!sk[112]) & (!g1108) & (!g1109) & (!g1111) & (g1125)) + ((!sk[112]) & (!g1108) & (!g1109) & (g1111) & (g1125)) + ((!sk[112]) & (!g1108) & (g1109) & (!g1111) & (g1125)) + ((!sk[112]) & (!g1108) & (g1109) & (g1111) & (g1125)) + ((!sk[112]) & (g1108) & (!g1109) & (!g1111) & (!g1125)) + ((!sk[112]) & (g1108) & (!g1109) & (!g1111) & (g1125)) + ((!sk[112]) & (g1108) & (!g1109) & (g1111) & (!g1125)) + ((!sk[112]) & (g1108) & (!g1109) & (g1111) & (g1125)) + ((!sk[112]) & (g1108) & (g1109) & (!g1111) & (!g1125)) + ((!sk[112]) & (g1108) & (g1109) & (!g1111) & (g1125)) + ((!sk[112]) & (g1108) & (g1109) & (g1111) & (!g1125)) + ((!sk[112]) & (g1108) & (g1109) & (g1111) & (g1125)) + ((sk[112]) & (!g1108) & (!g1109) & (!g1111) & (g1125)) + ((sk[112]) & (!g1108) & (!g1109) & (g1111) & (!g1125)) + ((sk[112]) & (!g1108) & (g1109) & (!g1111) & (!g1125)) + ((sk[112]) & (!g1108) & (g1109) & (g1111) & (g1125)) + ((sk[112]) & (g1108) & (!g1109) & (!g1111) & (!g1125)) + ((sk[112]) & (g1108) & (!g1109) & (g1111) & (g1125)) + ((sk[112]) & (g1108) & (g1109) & (!g1111) & (!g1125)) + ((sk[112]) & (g1108) & (g1109) & (g1111) & (g1125)));
	assign g1127 = (((!g9) & (!sk[113]) & (!g70) & (!g10) & (g18) & (!g40)) + ((!g9) & (!sk[113]) & (!g70) & (!g10) & (g18) & (g40)) + ((!g9) & (!sk[113]) & (!g70) & (g10) & (!g18) & (!g40)) + ((!g9) & (!sk[113]) & (!g70) & (g10) & (!g18) & (g40)) + ((!g9) & (!sk[113]) & (!g70) & (g10) & (g18) & (!g40)) + ((!g9) & (!sk[113]) & (!g70) & (g10) & (g18) & (g40)) + ((!g9) & (!sk[113]) & (g70) & (!g10) & (!g18) & (!g40)) + ((!g9) & (!sk[113]) & (g70) & (!g10) & (!g18) & (g40)) + ((!g9) & (!sk[113]) & (g70) & (!g10) & (g18) & (!g40)) + ((!g9) & (!sk[113]) & (g70) & (!g10) & (g18) & (g40)) + ((!g9) & (!sk[113]) & (g70) & (g10) & (!g18) & (!g40)) + ((!g9) & (!sk[113]) & (g70) & (g10) & (!g18) & (g40)) + ((!g9) & (!sk[113]) & (g70) & (g10) & (g18) & (!g40)) + ((!g9) & (!sk[113]) & (g70) & (g10) & (g18) & (g40)) + ((!g9) & (sk[113]) & (!g70) & (!g10) & (!g18) & (!g40)) + ((!g9) & (sk[113]) & (!g70) & (!g10) & (!g18) & (g40)) + ((!g9) & (sk[113]) & (!g70) & (!g10) & (g18) & (!g40)) + ((!g9) & (sk[113]) & (!g70) & (!g10) & (g18) & (g40)) + ((!g9) & (sk[113]) & (!g70) & (g10) & (!g18) & (!g40)) + ((!g9) & (sk[113]) & (!g70) & (g10) & (!g18) & (g40)) + ((!g9) & (sk[113]) & (!g70) & (g10) & (g18) & (!g40)) + ((!g9) & (sk[113]) & (!g70) & (g10) & (g18) & (g40)) + ((!g9) & (sk[113]) & (g70) & (!g10) & (!g18) & (!g40)) + ((!g9) & (sk[113]) & (g70) & (!g10) & (g18) & (!g40)) + ((g9) & (!sk[113]) & (!g70) & (!g10) & (g18) & (!g40)) + ((g9) & (!sk[113]) & (!g70) & (!g10) & (g18) & (g40)) + ((g9) & (!sk[113]) & (!g70) & (g10) & (!g18) & (!g40)) + ((g9) & (!sk[113]) & (!g70) & (g10) & (!g18) & (g40)) + ((g9) & (!sk[113]) & (!g70) & (g10) & (g18) & (!g40)) + ((g9) & (!sk[113]) & (!g70) & (g10) & (g18) & (g40)) + ((g9) & (!sk[113]) & (g70) & (!g10) & (!g18) & (!g40)) + ((g9) & (!sk[113]) & (g70) & (!g10) & (!g18) & (g40)) + ((g9) & (!sk[113]) & (g70) & (!g10) & (g18) & (!g40)) + ((g9) & (!sk[113]) & (g70) & (!g10) & (g18) & (g40)) + ((g9) & (!sk[113]) & (g70) & (g10) & (!g18) & (!g40)) + ((g9) & (!sk[113]) & (g70) & (g10) & (!g18) & (g40)) + ((g9) & (!sk[113]) & (g70) & (g10) & (g18) & (!g40)) + ((g9) & (!sk[113]) & (g70) & (g10) & (g18) & (g40)) + ((g9) & (sk[113]) & (!g70) & (!g10) & (!g18) & (!g40)) + ((g9) & (sk[113]) & (!g70) & (!g10) & (!g18) & (g40)) + ((g9) & (sk[113]) & (!g70) & (g10) & (!g18) & (!g40)) + ((g9) & (sk[113]) & (!g70) & (g10) & (!g18) & (g40)) + ((g9) & (sk[113]) & (g70) & (!g10) & (!g18) & (!g40)));
	assign g1128 = (((!g38) & (!g9) & (!g99) & (!g32) & (!g60) & (g1127)) + ((!g38) & (!g9) & (!g99) & (g32) & (!g60) & (g1127)) + ((!g38) & (!g9) & (g99) & (!g32) & (!g60) & (g1127)) + ((!g38) & (!g9) & (g99) & (g32) & (!g60) & (g1127)) + ((!g38) & (g9) & (!g99) & (!g32) & (!g60) & (g1127)) + ((!g38) & (g9) & (g99) & (!g32) & (!g60) & (g1127)) + ((g38) & (!g9) & (!g99) & (!g32) & (!g60) & (g1127)) + ((g38) & (!g9) & (!g99) & (g32) & (!g60) & (g1127)));
	assign g1129 = (((!sk[115]) & (!g10) & (!g17) & (!g99) & (g71) & (!g572)) + ((!sk[115]) & (!g10) & (!g17) & (!g99) & (g71) & (g572)) + ((!sk[115]) & (!g10) & (!g17) & (g99) & (!g71) & (!g572)) + ((!sk[115]) & (!g10) & (!g17) & (g99) & (!g71) & (g572)) + ((!sk[115]) & (!g10) & (!g17) & (g99) & (g71) & (!g572)) + ((!sk[115]) & (!g10) & (!g17) & (g99) & (g71) & (g572)) + ((!sk[115]) & (!g10) & (g17) & (!g99) & (!g71) & (!g572)) + ((!sk[115]) & (!g10) & (g17) & (!g99) & (!g71) & (g572)) + ((!sk[115]) & (!g10) & (g17) & (!g99) & (g71) & (!g572)) + ((!sk[115]) & (!g10) & (g17) & (!g99) & (g71) & (g572)) + ((!sk[115]) & (!g10) & (g17) & (g99) & (!g71) & (!g572)) + ((!sk[115]) & (!g10) & (g17) & (g99) & (!g71) & (g572)) + ((!sk[115]) & (!g10) & (g17) & (g99) & (g71) & (!g572)) + ((!sk[115]) & (!g10) & (g17) & (g99) & (g71) & (g572)) + ((!sk[115]) & (g10) & (!g17) & (!g99) & (g71) & (!g572)) + ((!sk[115]) & (g10) & (!g17) & (!g99) & (g71) & (g572)) + ((!sk[115]) & (g10) & (!g17) & (g99) & (!g71) & (!g572)) + ((!sk[115]) & (g10) & (!g17) & (g99) & (!g71) & (g572)) + ((!sk[115]) & (g10) & (!g17) & (g99) & (g71) & (!g572)) + ((!sk[115]) & (g10) & (!g17) & (g99) & (g71) & (g572)) + ((!sk[115]) & (g10) & (g17) & (!g99) & (!g71) & (!g572)) + ((!sk[115]) & (g10) & (g17) & (!g99) & (!g71) & (g572)) + ((!sk[115]) & (g10) & (g17) & (!g99) & (g71) & (!g572)) + ((!sk[115]) & (g10) & (g17) & (!g99) & (g71) & (g572)) + ((!sk[115]) & (g10) & (g17) & (g99) & (!g71) & (!g572)) + ((!sk[115]) & (g10) & (g17) & (g99) & (!g71) & (g572)) + ((!sk[115]) & (g10) & (g17) & (g99) & (g71) & (!g572)) + ((!sk[115]) & (g10) & (g17) & (g99) & (g71) & (g572)) + ((sk[115]) & (!g10) & (!g17) & (!g99) & (!g71) & (!g572)) + ((sk[115]) & (!g10) & (!g17) & (!g99) & (g71) & (!g572)) + ((sk[115]) & (!g10) & (!g17) & (g99) & (!g71) & (!g572)) + ((sk[115]) & (!g10) & (!g17) & (g99) & (g71) & (!g572)) + ((sk[115]) & (!g10) & (g17) & (!g99) & (!g71) & (!g572)) + ((sk[115]) & (!g10) & (g17) & (g99) & (!g71) & (!g572)) + ((sk[115]) & (g10) & (!g17) & (!g99) & (!g71) & (!g572)) + ((sk[115]) & (g10) & (!g17) & (!g99) & (g71) & (!g572)) + ((sk[115]) & (g10) & (g17) & (!g99) & (!g71) & (!g572)));
	assign g1130 = (((!g287) & (!g631) & (!sk[116]) & (!g637) & (g1129)) + ((!g287) & (!g631) & (!sk[116]) & (g637) & (g1129)) + ((!g287) & (g631) & (!sk[116]) & (!g637) & (g1129)) + ((!g287) & (g631) & (!sk[116]) & (g637) & (g1129)) + ((!g287) & (g631) & (sk[116]) & (g637) & (g1129)) + ((g287) & (!g631) & (!sk[116]) & (!g637) & (!g1129)) + ((g287) & (!g631) & (!sk[116]) & (!g637) & (g1129)) + ((g287) & (!g631) & (!sk[116]) & (g637) & (!g1129)) + ((g287) & (!g631) & (!sk[116]) & (g637) & (g1129)) + ((g287) & (g631) & (!sk[116]) & (!g637) & (!g1129)) + ((g287) & (g631) & (!sk[116]) & (!g637) & (g1129)) + ((g287) & (g631) & (!sk[116]) & (g637) & (!g1129)) + ((g287) & (g631) & (!sk[116]) & (g637) & (g1129)));
	assign g1131 = (((!g266) & (!g1028) & (!g1128) & (!sk[117]) & (g1130)) + ((!g266) & (!g1028) & (g1128) & (!sk[117]) & (g1130)) + ((!g266) & (g1028) & (!g1128) & (!sk[117]) & (g1130)) + ((!g266) & (g1028) & (g1128) & (!sk[117]) & (g1130)) + ((g266) & (!g1028) & (!g1128) & (!sk[117]) & (!g1130)) + ((g266) & (!g1028) & (!g1128) & (!sk[117]) & (g1130)) + ((g266) & (!g1028) & (g1128) & (!sk[117]) & (!g1130)) + ((g266) & (!g1028) & (g1128) & (!sk[117]) & (g1130)) + ((g266) & (g1028) & (!g1128) & (!sk[117]) & (!g1130)) + ((g266) & (g1028) & (!g1128) & (!sk[117]) & (g1130)) + ((g266) & (g1028) & (g1128) & (!sk[117]) & (!g1130)) + ((g266) & (g1028) & (g1128) & (!sk[117]) & (g1130)) + ((g266) & (g1028) & (g1128) & (sk[117]) & (g1130)));
	assign g1132 = (((!g1031) & (!g1060) & (!sk[118]) & (!g1065) & (g1098) & (!g1105)) + ((!g1031) & (!g1060) & (!sk[118]) & (!g1065) & (g1098) & (g1105)) + ((!g1031) & (!g1060) & (!sk[118]) & (g1065) & (!g1098) & (!g1105)) + ((!g1031) & (!g1060) & (!sk[118]) & (g1065) & (!g1098) & (g1105)) + ((!g1031) & (!g1060) & (!sk[118]) & (g1065) & (g1098) & (!g1105)) + ((!g1031) & (!g1060) & (!sk[118]) & (g1065) & (g1098) & (g1105)) + ((!g1031) & (!g1060) & (sk[118]) & (!g1065) & (g1098) & (!g1105)) + ((!g1031) & (!g1060) & (sk[118]) & (g1065) & (g1098) & (!g1105)) + ((!g1031) & (g1060) & (!sk[118]) & (!g1065) & (!g1098) & (!g1105)) + ((!g1031) & (g1060) & (!sk[118]) & (!g1065) & (!g1098) & (g1105)) + ((!g1031) & (g1060) & (!sk[118]) & (!g1065) & (g1098) & (!g1105)) + ((!g1031) & (g1060) & (!sk[118]) & (!g1065) & (g1098) & (g1105)) + ((!g1031) & (g1060) & (!sk[118]) & (g1065) & (!g1098) & (!g1105)) + ((!g1031) & (g1060) & (!sk[118]) & (g1065) & (!g1098) & (g1105)) + ((!g1031) & (g1060) & (!sk[118]) & (g1065) & (g1098) & (!g1105)) + ((!g1031) & (g1060) & (!sk[118]) & (g1065) & (g1098) & (g1105)) + ((!g1031) & (g1060) & (sk[118]) & (!g1065) & (!g1098) & (!g1105)) + ((!g1031) & (g1060) & (sk[118]) & (!g1065) & (g1098) & (!g1105)) + ((!g1031) & (g1060) & (sk[118]) & (!g1065) & (g1098) & (g1105)) + ((!g1031) & (g1060) & (sk[118]) & (g1065) & (g1098) & (!g1105)) + ((g1031) & (!g1060) & (!sk[118]) & (!g1065) & (g1098) & (!g1105)) + ((g1031) & (!g1060) & (!sk[118]) & (!g1065) & (g1098) & (g1105)) + ((g1031) & (!g1060) & (!sk[118]) & (g1065) & (!g1098) & (!g1105)) + ((g1031) & (!g1060) & (!sk[118]) & (g1065) & (!g1098) & (g1105)) + ((g1031) & (!g1060) & (!sk[118]) & (g1065) & (g1098) & (!g1105)) + ((g1031) & (!g1060) & (!sk[118]) & (g1065) & (g1098) & (g1105)) + ((g1031) & (!g1060) & (sk[118]) & (!g1065) & (!g1098) & (!g1105)) + ((g1031) & (!g1060) & (sk[118]) & (!g1065) & (g1098) & (!g1105)) + ((g1031) & (!g1060) & (sk[118]) & (!g1065) & (g1098) & (g1105)) + ((g1031) & (!g1060) & (sk[118]) & (g1065) & (g1098) & (!g1105)) + ((g1031) & (g1060) & (!sk[118]) & (!g1065) & (!g1098) & (!g1105)) + ((g1031) & (g1060) & (!sk[118]) & (!g1065) & (!g1098) & (g1105)) + ((g1031) & (g1060) & (!sk[118]) & (!g1065) & (g1098) & (!g1105)) + ((g1031) & (g1060) & (!sk[118]) & (!g1065) & (g1098) & (g1105)) + ((g1031) & (g1060) & (!sk[118]) & (g1065) & (!g1098) & (!g1105)) + ((g1031) & (g1060) & (!sk[118]) & (g1065) & (!g1098) & (g1105)) + ((g1031) & (g1060) & (!sk[118]) & (g1065) & (g1098) & (!g1105)) + ((g1031) & (g1060) & (!sk[118]) & (g1065) & (g1098) & (g1105)) + ((g1031) & (g1060) & (sk[118]) & (!g1065) & (!g1098) & (!g1105)) + ((g1031) & (g1060) & (sk[118]) & (!g1065) & (g1098) & (!g1105)) + ((g1031) & (g1060) & (sk[118]) & (!g1065) & (g1098) & (g1105)) + ((g1031) & (g1060) & (sk[118]) & (g1065) & (!g1098) & (!g1105)) + ((g1031) & (g1060) & (sk[118]) & (g1065) & (g1098) & (!g1105)) + ((g1031) & (g1060) & (sk[118]) & (g1065) & (g1098) & (g1105)));
	assign g1133 = (((!sk[119]) & (!g1126) & (g1131) & (!g1132)) + ((!sk[119]) & (!g1126) & (g1131) & (g1132)) + ((!sk[119]) & (g1126) & (g1131) & (!g1132)) + ((!sk[119]) & (g1126) & (g1131) & (g1132)) + ((sk[119]) & (!g1126) & (!g1131) & (!g1132)) + ((sk[119]) & (!g1126) & (g1131) & (g1132)) + ((sk[119]) & (g1126) & (!g1131) & (g1132)) + ((sk[119]) & (g1126) & (g1131) & (!g1132)));
	assign g1134 = (((!g1067) & (!g1068) & (!g1069) & (!sk[120]) & (g1106) & (!g1133)) + ((!g1067) & (!g1068) & (!g1069) & (!sk[120]) & (g1106) & (g1133)) + ((!g1067) & (!g1068) & (!g1069) & (sk[120]) & (!g1106) & (!g1133)) + ((!g1067) & (!g1068) & (!g1069) & (sk[120]) & (g1106) & (!g1133)) + ((!g1067) & (!g1068) & (g1069) & (!sk[120]) & (!g1106) & (!g1133)) + ((!g1067) & (!g1068) & (g1069) & (!sk[120]) & (!g1106) & (g1133)) + ((!g1067) & (!g1068) & (g1069) & (!sk[120]) & (g1106) & (!g1133)) + ((!g1067) & (!g1068) & (g1069) & (!sk[120]) & (g1106) & (g1133)) + ((!g1067) & (!g1068) & (g1069) & (sk[120]) & (!g1106) & (!g1133)) + ((!g1067) & (!g1068) & (g1069) & (sk[120]) & (g1106) & (g1133)) + ((!g1067) & (g1068) & (!g1069) & (!sk[120]) & (!g1106) & (!g1133)) + ((!g1067) & (g1068) & (!g1069) & (!sk[120]) & (!g1106) & (g1133)) + ((!g1067) & (g1068) & (!g1069) & (!sk[120]) & (g1106) & (!g1133)) + ((!g1067) & (g1068) & (!g1069) & (!sk[120]) & (g1106) & (g1133)) + ((!g1067) & (g1068) & (!g1069) & (sk[120]) & (!g1106) & (g1133)) + ((!g1067) & (g1068) & (!g1069) & (sk[120]) & (g1106) & (g1133)) + ((!g1067) & (g1068) & (g1069) & (!sk[120]) & (!g1106) & (!g1133)) + ((!g1067) & (g1068) & (g1069) & (!sk[120]) & (!g1106) & (g1133)) + ((!g1067) & (g1068) & (g1069) & (!sk[120]) & (g1106) & (!g1133)) + ((!g1067) & (g1068) & (g1069) & (!sk[120]) & (g1106) & (g1133)) + ((!g1067) & (g1068) & (g1069) & (sk[120]) & (!g1106) & (g1133)) + ((!g1067) & (g1068) & (g1069) & (sk[120]) & (g1106) & (!g1133)) + ((g1067) & (!g1068) & (!g1069) & (!sk[120]) & (g1106) & (!g1133)) + ((g1067) & (!g1068) & (!g1069) & (!sk[120]) & (g1106) & (g1133)) + ((g1067) & (!g1068) & (!g1069) & (sk[120]) & (!g1106) & (!g1133)) + ((g1067) & (!g1068) & (!g1069) & (sk[120]) & (g1106) & (!g1133)) + ((g1067) & (!g1068) & (g1069) & (!sk[120]) & (!g1106) & (!g1133)) + ((g1067) & (!g1068) & (g1069) & (!sk[120]) & (!g1106) & (g1133)) + ((g1067) & (!g1068) & (g1069) & (!sk[120]) & (g1106) & (!g1133)) + ((g1067) & (!g1068) & (g1069) & (!sk[120]) & (g1106) & (g1133)) + ((g1067) & (!g1068) & (g1069) & (sk[120]) & (!g1106) & (!g1133)) + ((g1067) & (!g1068) & (g1069) & (sk[120]) & (g1106) & (g1133)) + ((g1067) & (g1068) & (!g1069) & (!sk[120]) & (!g1106) & (!g1133)) + ((g1067) & (g1068) & (!g1069) & (!sk[120]) & (!g1106) & (g1133)) + ((g1067) & (g1068) & (!g1069) & (!sk[120]) & (g1106) & (!g1133)) + ((g1067) & (g1068) & (!g1069) & (!sk[120]) & (g1106) & (g1133)) + ((g1067) & (g1068) & (!g1069) & (sk[120]) & (!g1106) & (!g1133)) + ((g1067) & (g1068) & (!g1069) & (sk[120]) & (g1106) & (g1133)) + ((g1067) & (g1068) & (g1069) & (!sk[120]) & (!g1106) & (!g1133)) + ((g1067) & (g1068) & (g1069) & (!sk[120]) & (!g1106) & (g1133)) + ((g1067) & (g1068) & (g1069) & (!sk[120]) & (g1106) & (!g1133)) + ((g1067) & (g1068) & (g1069) & (!sk[120]) & (g1106) & (g1133)) + ((g1067) & (g1068) & (g1069) & (sk[120]) & (!g1106) & (g1133)) + ((g1067) & (g1068) & (g1069) & (sk[120]) & (g1106) & (g1133)));
	assign g1135 = (((!sk[121]) & (!g1069) & (!g1106) & (!g1126) & (g1131) & (!g1132)) + ((!sk[121]) & (!g1069) & (!g1106) & (!g1126) & (g1131) & (g1132)) + ((!sk[121]) & (!g1069) & (!g1106) & (g1126) & (!g1131) & (!g1132)) + ((!sk[121]) & (!g1069) & (!g1106) & (g1126) & (!g1131) & (g1132)) + ((!sk[121]) & (!g1069) & (!g1106) & (g1126) & (g1131) & (!g1132)) + ((!sk[121]) & (!g1069) & (!g1106) & (g1126) & (g1131) & (g1132)) + ((!sk[121]) & (!g1069) & (g1106) & (!g1126) & (!g1131) & (!g1132)) + ((!sk[121]) & (!g1069) & (g1106) & (!g1126) & (!g1131) & (g1132)) + ((!sk[121]) & (!g1069) & (g1106) & (!g1126) & (g1131) & (!g1132)) + ((!sk[121]) & (!g1069) & (g1106) & (!g1126) & (g1131) & (g1132)) + ((!sk[121]) & (!g1069) & (g1106) & (g1126) & (!g1131) & (!g1132)) + ((!sk[121]) & (!g1069) & (g1106) & (g1126) & (!g1131) & (g1132)) + ((!sk[121]) & (!g1069) & (g1106) & (g1126) & (g1131) & (!g1132)) + ((!sk[121]) & (!g1069) & (g1106) & (g1126) & (g1131) & (g1132)) + ((!sk[121]) & (g1069) & (!g1106) & (!g1126) & (g1131) & (!g1132)) + ((!sk[121]) & (g1069) & (!g1106) & (!g1126) & (g1131) & (g1132)) + ((!sk[121]) & (g1069) & (!g1106) & (g1126) & (!g1131) & (!g1132)) + ((!sk[121]) & (g1069) & (!g1106) & (g1126) & (!g1131) & (g1132)) + ((!sk[121]) & (g1069) & (!g1106) & (g1126) & (g1131) & (!g1132)) + ((!sk[121]) & (g1069) & (!g1106) & (g1126) & (g1131) & (g1132)) + ((!sk[121]) & (g1069) & (g1106) & (!g1126) & (!g1131) & (!g1132)) + ((!sk[121]) & (g1069) & (g1106) & (!g1126) & (!g1131) & (g1132)) + ((!sk[121]) & (g1069) & (g1106) & (!g1126) & (g1131) & (!g1132)) + ((!sk[121]) & (g1069) & (g1106) & (!g1126) & (g1131) & (g1132)) + ((!sk[121]) & (g1069) & (g1106) & (g1126) & (!g1131) & (!g1132)) + ((!sk[121]) & (g1069) & (g1106) & (g1126) & (!g1131) & (g1132)) + ((!sk[121]) & (g1069) & (g1106) & (g1126) & (g1131) & (!g1132)) + ((!sk[121]) & (g1069) & (g1106) & (g1126) & (g1131) & (g1132)) + ((sk[121]) & (g1069) & (g1106) & (!g1126) & (!g1131) & (!g1132)) + ((sk[121]) & (g1069) & (g1106) & (!g1126) & (g1131) & (g1132)) + ((sk[121]) & (g1069) & (g1106) & (g1126) & (!g1131) & (g1132)) + ((sk[121]) & (g1069) & (g1106) & (g1126) & (g1131) & (!g1132)));
	assign g1136 = (((!sk[122]) & (!g1112) & (g1122) & (!g1124)) + ((!sk[122]) & (!g1112) & (g1122) & (g1124)) + ((!sk[122]) & (g1112) & (g1122) & (!g1124)) + ((!sk[122]) & (g1112) & (g1122) & (g1124)) + ((sk[122]) & (!g1112) & (!g1122) & (!g1124)) + ((sk[122]) & (g1112) & (!g1122) & (!g1124)) + ((sk[122]) & (g1112) & (!g1122) & (g1124)) + ((sk[122]) & (g1112) & (g1122) & (!g1124)));
	assign g1137 = (((!g1083) & (!g1085) & (!g1086) & (!g1093) & (g1114) & (!g1121)) + ((!g1083) & (!g1085) & (!g1086) & (g1093) & (g1114) & (!g1121)) + ((!g1083) & (!g1085) & (g1086) & (!g1093) & (g1114) & (!g1121)) + ((!g1083) & (!g1085) & (g1086) & (g1093) & (g1114) & (!g1121)) + ((!g1083) & (g1085) & (!g1086) & (!g1093) & (!g1114) & (!g1121)) + ((!g1083) & (g1085) & (!g1086) & (!g1093) & (g1114) & (!g1121)) + ((!g1083) & (g1085) & (!g1086) & (!g1093) & (g1114) & (g1121)) + ((!g1083) & (g1085) & (!g1086) & (g1093) & (g1114) & (!g1121)) + ((!g1083) & (g1085) & (g1086) & (!g1093) & (g1114) & (!g1121)) + ((!g1083) & (g1085) & (g1086) & (g1093) & (!g1114) & (!g1121)) + ((!g1083) & (g1085) & (g1086) & (g1093) & (g1114) & (!g1121)) + ((!g1083) & (g1085) & (g1086) & (g1093) & (g1114) & (g1121)) + ((g1083) & (!g1085) & (!g1086) & (!g1093) & (!g1114) & (!g1121)) + ((g1083) & (!g1085) & (!g1086) & (!g1093) & (g1114) & (!g1121)) + ((g1083) & (!g1085) & (!g1086) & (!g1093) & (g1114) & (g1121)) + ((g1083) & (!g1085) & (!g1086) & (g1093) & (g1114) & (!g1121)) + ((g1083) & (!g1085) & (g1086) & (!g1093) & (g1114) & (!g1121)) + ((g1083) & (!g1085) & (g1086) & (g1093) & (!g1114) & (!g1121)) + ((g1083) & (!g1085) & (g1086) & (g1093) & (g1114) & (!g1121)) + ((g1083) & (!g1085) & (g1086) & (g1093) & (g1114) & (g1121)) + ((g1083) & (g1085) & (!g1086) & (!g1093) & (!g1114) & (!g1121)) + ((g1083) & (g1085) & (!g1086) & (!g1093) & (g1114) & (!g1121)) + ((g1083) & (g1085) & (!g1086) & (!g1093) & (g1114) & (g1121)) + ((g1083) & (g1085) & (!g1086) & (g1093) & (!g1114) & (!g1121)) + ((g1083) & (g1085) & (!g1086) & (g1093) & (g1114) & (!g1121)) + ((g1083) & (g1085) & (!g1086) & (g1093) & (g1114) & (g1121)) + ((g1083) & (g1085) & (g1086) & (!g1093) & (!g1114) & (!g1121)) + ((g1083) & (g1085) & (g1086) & (!g1093) & (g1114) & (!g1121)) + ((g1083) & (g1085) & (g1086) & (!g1093) & (g1114) & (g1121)) + ((g1083) & (g1085) & (g1086) & (g1093) & (!g1114) & (!g1121)) + ((g1083) & (g1085) & (g1086) & (g1093) & (g1114) & (!g1121)) + ((g1083) & (g1085) & (g1086) & (g1093) & (g1114) & (g1121)));
	assign g1138 = (((!sk[124]) & (!g707) & (!g717) & (!g718) & (g762) & (!g765)) + ((!sk[124]) & (!g707) & (!g717) & (!g718) & (g762) & (g765)) + ((!sk[124]) & (!g707) & (!g717) & (g718) & (!g762) & (!g765)) + ((!sk[124]) & (!g707) & (!g717) & (g718) & (!g762) & (g765)) + ((!sk[124]) & (!g707) & (!g717) & (g718) & (g762) & (!g765)) + ((!sk[124]) & (!g707) & (!g717) & (g718) & (g762) & (g765)) + ((!sk[124]) & (!g707) & (g717) & (!g718) & (!g762) & (!g765)) + ((!sk[124]) & (!g707) & (g717) & (!g718) & (!g762) & (g765)) + ((!sk[124]) & (!g707) & (g717) & (!g718) & (g762) & (!g765)) + ((!sk[124]) & (!g707) & (g717) & (!g718) & (g762) & (g765)) + ((!sk[124]) & (!g707) & (g717) & (g718) & (!g762) & (!g765)) + ((!sk[124]) & (!g707) & (g717) & (g718) & (!g762) & (g765)) + ((!sk[124]) & (!g707) & (g717) & (g718) & (g762) & (!g765)) + ((!sk[124]) & (!g707) & (g717) & (g718) & (g762) & (g765)) + ((!sk[124]) & (g707) & (!g717) & (!g718) & (g762) & (!g765)) + ((!sk[124]) & (g707) & (!g717) & (!g718) & (g762) & (g765)) + ((!sk[124]) & (g707) & (!g717) & (g718) & (!g762) & (!g765)) + ((!sk[124]) & (g707) & (!g717) & (g718) & (!g762) & (g765)) + ((!sk[124]) & (g707) & (!g717) & (g718) & (g762) & (!g765)) + ((!sk[124]) & (g707) & (!g717) & (g718) & (g762) & (g765)) + ((!sk[124]) & (g707) & (g717) & (!g718) & (!g762) & (!g765)) + ((!sk[124]) & (g707) & (g717) & (!g718) & (!g762) & (g765)) + ((!sk[124]) & (g707) & (g717) & (!g718) & (g762) & (!g765)) + ((!sk[124]) & (g707) & (g717) & (!g718) & (g762) & (g765)) + ((!sk[124]) & (g707) & (g717) & (g718) & (!g762) & (!g765)) + ((!sk[124]) & (g707) & (g717) & (g718) & (!g762) & (g765)) + ((!sk[124]) & (g707) & (g717) & (g718) & (g762) & (!g765)) + ((!sk[124]) & (g707) & (g717) & (g718) & (g762) & (g765)) + ((sk[124]) & (!g707) & (!g717) & (g718) & (!g762) & (g765)) + ((sk[124]) & (!g707) & (!g717) & (g718) & (g762) & (g765)) + ((sk[124]) & (!g707) & (g717) & (!g718) & (g762) & (!g765)) + ((sk[124]) & (!g707) & (g717) & (!g718) & (g762) & (g765)) + ((sk[124]) & (!g707) & (g717) & (g718) & (!g762) & (g765)) + ((sk[124]) & (!g707) & (g717) & (g718) & (g762) & (!g765)) + ((sk[124]) & (!g707) & (g717) & (g718) & (g762) & (g765)) + ((sk[124]) & (g707) & (!g717) & (!g718) & (g762) & (!g765)) + ((sk[124]) & (g707) & (!g717) & (!g718) & (g762) & (g765)) + ((sk[124]) & (g707) & (!g717) & (g718) & (!g762) & (g765)) + ((sk[124]) & (g707) & (!g717) & (g718) & (g762) & (!g765)) + ((sk[124]) & (g707) & (!g717) & (g718) & (g762) & (g765)) + ((sk[124]) & (g707) & (g717) & (g718) & (!g762) & (g765)) + ((sk[124]) & (g707) & (g717) & (g718) & (g762) & (g765)));
	assign g1139 = (((!g869) & (!g764) & (!g759) & (!g870) & (!g834) & (!g1138)) + ((!g869) & (!g764) & (!g759) & (!g870) & (g834) & (!g1138)) + ((!g869) & (!g764) & (!g759) & (g870) & (!g834) & (!g1138)) + ((!g869) & (!g764) & (!g759) & (g870) & (g834) & (!g1138)) + ((!g869) & (!g764) & (g759) & (!g870) & (g834) & (!g1138)) + ((!g869) & (!g764) & (g759) & (g870) & (!g834) & (!g1138)) + ((!g869) & (g764) & (!g759) & (g870) & (!g834) & (!g1138)) + ((!g869) & (g764) & (!g759) & (g870) & (g834) & (!g1138)) + ((!g869) & (g764) & (g759) & (g870) & (!g834) & (!g1138)) + ((g869) & (!g764) & (!g759) & (!g870) & (!g834) & (!g1138)) + ((g869) & (!g764) & (!g759) & (!g870) & (g834) & (!g1138)) + ((g869) & (!g764) & (!g759) & (g870) & (!g834) & (!g1138)) + ((g869) & (!g764) & (!g759) & (g870) & (g834) & (!g1138)) + ((g869) & (!g764) & (g759) & (!g870) & (!g834) & (!g1138)) + ((g869) & (!g764) & (g759) & (g870) & (g834) & (!g1138)) + ((g869) & (g764) & (!g759) & (g870) & (!g834) & (!g1138)) + ((g869) & (g764) & (!g759) & (g870) & (g834) & (!g1138)) + ((g869) & (g764) & (g759) & (g870) & (g834) & (!g1138)));
	assign g1140 = (((!g252) & (!g722) & (!g723) & (g1089) & (!g1091) & (!g1119)) + ((!g252) & (!g722) & (g723) & (g1089) & (!g1091) & (!g1119)) + ((!g252) & (g722) & (!g723) & (g1089) & (!g1091) & (!g1119)) + ((!g252) & (g722) & (g723) & (g1089) & (!g1091) & (!g1119)) + ((g252) & (!g722) & (!g723) & (!g1089) & (!g1091) & (g1119)) + ((g252) & (!g722) & (!g723) & (!g1089) & (g1091) & (!g1119)) + ((g252) & (!g722) & (!g723) & (!g1089) & (g1091) & (g1119)) + ((g252) & (!g722) & (!g723) & (g1089) & (!g1091) & (!g1119)) + ((g252) & (!g722) & (!g723) & (g1089) & (!g1091) & (g1119)) + ((g252) & (!g722) & (!g723) & (g1089) & (g1091) & (!g1119)) + ((g252) & (!g722) & (!g723) & (g1089) & (g1091) & (g1119)) + ((g252) & (!g722) & (g723) & (!g1089) & (!g1091) & (g1119)) + ((g252) & (!g722) & (g723) & (!g1089) & (g1091) & (g1119)) + ((g252) & (!g722) & (g723) & (g1089) & (!g1091) & (g1119)) + ((g252) & (!g722) & (g723) & (g1089) & (g1091) & (!g1119)) + ((g252) & (!g722) & (g723) & (g1089) & (g1091) & (g1119)) + ((g252) & (g722) & (!g723) & (!g1089) & (g1091) & (g1119)) + ((g252) & (g722) & (!g723) & (g1089) & (!g1091) & (g1119)) + ((g252) & (g722) & (!g723) & (g1089) & (g1091) & (g1119)) + ((g252) & (g722) & (g723) & (g1089) & (g1091) & (g1119)));
	assign g1141 = (((!g549) & (!g569) & (!g680) & (!g729) & (!g847) & (g845)) + ((!g549) & (!g569) & (!g680) & (!g729) & (g847) & (g845)) + ((!g549) & (!g569) & (g680) & (!g729) & (!g847) & (g845)) + ((!g549) & (!g569) & (g680) & (!g729) & (g847) & (!g845)) + ((!g549) & (!g569) & (g680) & (!g729) & (g847) & (g845)) + ((!g549) & (!g569) & (g680) & (g729) & (g847) & (!g845)) + ((!g549) & (!g569) & (g680) & (g729) & (g847) & (g845)) + ((!g549) & (g569) & (!g680) & (!g729) & (!g847) & (g845)) + ((!g549) & (g569) & (!g680) & (!g729) & (g847) & (!g845)) + ((!g549) & (g569) & (!g680) & (!g729) & (g847) & (g845)) + ((!g549) & (g569) & (!g680) & (g729) & (g847) & (!g845)) + ((!g549) & (g569) & (!g680) & (g729) & (g847) & (g845)) + ((!g549) & (g569) & (g680) & (!g729) & (!g847) & (g845)) + ((!g549) & (g569) & (g680) & (!g729) & (g847) & (g845)) + ((g549) & (!g569) & (!g680) & (!g729) & (!g847) & (g845)) + ((g549) & (!g569) & (!g680) & (!g729) & (g847) & (!g845)) + ((g549) & (!g569) & (!g680) & (!g729) & (g847) & (g845)) + ((g549) & (!g569) & (!g680) & (g729) & (g847) & (!g845)) + ((g549) & (!g569) & (!g680) & (g729) & (g847) & (g845)) + ((g549) & (!g569) & (g680) & (!g729) & (!g847) & (g845)) + ((g549) & (!g569) & (g680) & (!g729) & (g847) & (g845)) + ((g549) & (g569) & (!g680) & (!g729) & (!g847) & (g845)) + ((g549) & (g569) & (!g680) & (!g729) & (g847) & (g845)) + ((g549) & (g569) & (g680) & (!g729) & (!g847) & (g845)) + ((g549) & (g569) & (g680) & (!g729) & (g847) & (!g845)) + ((g549) & (g569) & (g680) & (!g729) & (g847) & (g845)) + ((g549) & (g569) & (g680) & (g729) & (g847) & (!g845)) + ((g549) & (g569) & (g680) & (g729) & (g847) & (g845)));
	assign g1142 = (((!g719) & (!sk[0]) & (!g843) & (!g791) & (g848) & (!g1141)) + ((!g719) & (!sk[0]) & (!g843) & (!g791) & (g848) & (g1141)) + ((!g719) & (!sk[0]) & (!g843) & (g791) & (!g848) & (!g1141)) + ((!g719) & (!sk[0]) & (!g843) & (g791) & (!g848) & (g1141)) + ((!g719) & (!sk[0]) & (!g843) & (g791) & (g848) & (!g1141)) + ((!g719) & (!sk[0]) & (!g843) & (g791) & (g848) & (g1141)) + ((!g719) & (!sk[0]) & (g843) & (!g791) & (!g848) & (!g1141)) + ((!g719) & (!sk[0]) & (g843) & (!g791) & (!g848) & (g1141)) + ((!g719) & (!sk[0]) & (g843) & (!g791) & (g848) & (!g1141)) + ((!g719) & (!sk[0]) & (g843) & (!g791) & (g848) & (g1141)) + ((!g719) & (!sk[0]) & (g843) & (g791) & (!g848) & (!g1141)) + ((!g719) & (!sk[0]) & (g843) & (g791) & (!g848) & (g1141)) + ((!g719) & (!sk[0]) & (g843) & (g791) & (g848) & (!g1141)) + ((!g719) & (!sk[0]) & (g843) & (g791) & (g848) & (g1141)) + ((!g719) & (sk[0]) & (!g843) & (!g791) & (!g848) & (!g1141)) + ((!g719) & (sk[0]) & (!g843) & (g791) & (!g848) & (!g1141)) + ((!g719) & (sk[0]) & (g843) & (!g791) & (!g848) & (!g1141)) + ((g719) & (!sk[0]) & (!g843) & (!g791) & (g848) & (!g1141)) + ((g719) & (!sk[0]) & (!g843) & (!g791) & (g848) & (g1141)) + ((g719) & (!sk[0]) & (!g843) & (g791) & (!g848) & (!g1141)) + ((g719) & (!sk[0]) & (!g843) & (g791) & (!g848) & (g1141)) + ((g719) & (!sk[0]) & (!g843) & (g791) & (g848) & (!g1141)) + ((g719) & (!sk[0]) & (!g843) & (g791) & (g848) & (g1141)) + ((g719) & (!sk[0]) & (g843) & (!g791) & (!g848) & (!g1141)) + ((g719) & (!sk[0]) & (g843) & (!g791) & (!g848) & (g1141)) + ((g719) & (!sk[0]) & (g843) & (!g791) & (g848) & (!g1141)) + ((g719) & (!sk[0]) & (g843) & (!g791) & (g848) & (g1141)) + ((g719) & (!sk[0]) & (g843) & (g791) & (!g848) & (!g1141)) + ((g719) & (!sk[0]) & (g843) & (g791) & (!g848) & (g1141)) + ((g719) & (!sk[0]) & (g843) & (g791) & (g848) & (!g1141)) + ((g719) & (!sk[0]) & (g843) & (g791) & (g848) & (g1141)) + ((g719) & (sk[0]) & (!g843) & (!g791) & (!g848) & (!g1141)) + ((g719) & (sk[0]) & (!g843) & (!g791) & (g848) & (!g1141)) + ((g719) & (sk[0]) & (!g843) & (g791) & (!g848) & (!g1141)) + ((g719) & (sk[0]) & (!g843) & (g791) & (g848) & (!g1141)) + ((g719) & (sk[0]) & (g843) & (!g791) & (!g848) & (!g1141)) + ((g719) & (sk[0]) & (g843) & (!g791) & (g848) & (!g1141)));
	assign g1143 = (((!g252) & (!sk[1]) & (!g720) & (!g1140) & (g1142)) + ((!g252) & (!sk[1]) & (!g720) & (g1140) & (g1142)) + ((!g252) & (!sk[1]) & (g720) & (!g1140) & (g1142)) + ((!g252) & (!sk[1]) & (g720) & (g1140) & (g1142)) + ((!g252) & (sk[1]) & (!g720) & (!g1140) & (!g1142)) + ((!g252) & (sk[1]) & (!g720) & (g1140) & (g1142)) + ((!g252) & (sk[1]) & (g720) & (!g1140) & (!g1142)) + ((!g252) & (sk[1]) & (g720) & (g1140) & (g1142)) + ((g252) & (!sk[1]) & (!g720) & (!g1140) & (!g1142)) + ((g252) & (!sk[1]) & (!g720) & (!g1140) & (g1142)) + ((g252) & (!sk[1]) & (!g720) & (g1140) & (!g1142)) + ((g252) & (!sk[1]) & (!g720) & (g1140) & (g1142)) + ((g252) & (!sk[1]) & (g720) & (!g1140) & (!g1142)) + ((g252) & (!sk[1]) & (g720) & (!g1140) & (g1142)) + ((g252) & (!sk[1]) & (g720) & (g1140) & (!g1142)) + ((g252) & (!sk[1]) & (g720) & (g1140) & (g1142)) + ((g252) & (sk[1]) & (!g720) & (!g1140) & (g1142)) + ((g252) & (sk[1]) & (!g720) & (g1140) & (!g1142)) + ((g252) & (sk[1]) & (g720) & (!g1140) & (!g1142)) + ((g252) & (sk[1]) & (g720) & (g1140) & (g1142)));
	assign g1144 = (((!g202) & (!g1115) & (!g1117) & (!g1120) & (!g1139) & (g1143)) + ((!g202) & (!g1115) & (!g1117) & (!g1120) & (g1139) & (!g1143)) + ((!g202) & (!g1115) & (!g1117) & (g1120) & (!g1139) & (!g1143)) + ((!g202) & (!g1115) & (!g1117) & (g1120) & (g1139) & (g1143)) + ((!g202) & (!g1115) & (g1117) & (!g1120) & (!g1139) & (g1143)) + ((!g202) & (!g1115) & (g1117) & (!g1120) & (g1139) & (!g1143)) + ((!g202) & (!g1115) & (g1117) & (g1120) & (!g1139) & (g1143)) + ((!g202) & (!g1115) & (g1117) & (g1120) & (g1139) & (!g1143)) + ((!g202) & (g1115) & (!g1117) & (!g1120) & (!g1139) & (!g1143)) + ((!g202) & (g1115) & (!g1117) & (!g1120) & (g1139) & (g1143)) + ((!g202) & (g1115) & (!g1117) & (g1120) & (!g1139) & (!g1143)) + ((!g202) & (g1115) & (!g1117) & (g1120) & (g1139) & (g1143)) + ((!g202) & (g1115) & (g1117) & (!g1120) & (!g1139) & (g1143)) + ((!g202) & (g1115) & (g1117) & (!g1120) & (g1139) & (!g1143)) + ((!g202) & (g1115) & (g1117) & (g1120) & (!g1139) & (!g1143)) + ((!g202) & (g1115) & (g1117) & (g1120) & (g1139) & (g1143)) + ((g202) & (!g1115) & (!g1117) & (!g1120) & (!g1139) & (!g1143)) + ((g202) & (!g1115) & (!g1117) & (!g1120) & (g1139) & (g1143)) + ((g202) & (!g1115) & (!g1117) & (g1120) & (!g1139) & (g1143)) + ((g202) & (!g1115) & (!g1117) & (g1120) & (g1139) & (!g1143)) + ((g202) & (!g1115) & (g1117) & (!g1120) & (!g1139) & (!g1143)) + ((g202) & (!g1115) & (g1117) & (!g1120) & (g1139) & (g1143)) + ((g202) & (!g1115) & (g1117) & (g1120) & (!g1139) & (!g1143)) + ((g202) & (!g1115) & (g1117) & (g1120) & (g1139) & (g1143)) + ((g202) & (g1115) & (!g1117) & (!g1120) & (!g1139) & (g1143)) + ((g202) & (g1115) & (!g1117) & (!g1120) & (g1139) & (!g1143)) + ((g202) & (g1115) & (!g1117) & (g1120) & (!g1139) & (g1143)) + ((g202) & (g1115) & (!g1117) & (g1120) & (g1139) & (!g1143)) + ((g202) & (g1115) & (g1117) & (!g1120) & (!g1139) & (!g1143)) + ((g202) & (g1115) & (g1117) & (!g1120) & (g1139) & (g1143)) + ((g202) & (g1115) & (g1117) & (g1120) & (!g1139) & (g1143)) + ((g202) & (g1115) & (g1117) & (g1120) & (g1139) & (!g1143)));
	assign g1145 = (((!sk[3]) & (g748) & (g863)) + ((sk[3]) & (g748) & (g863)));
	assign g1146 = (((!g747) & (!g744) & (!sk[4]) & (!g889) & (g871) & (!g883)) + ((!g747) & (!g744) & (!sk[4]) & (!g889) & (g871) & (g883)) + ((!g747) & (!g744) & (!sk[4]) & (g889) & (!g871) & (!g883)) + ((!g747) & (!g744) & (!sk[4]) & (g889) & (!g871) & (g883)) + ((!g747) & (!g744) & (!sk[4]) & (g889) & (g871) & (!g883)) + ((!g747) & (!g744) & (!sk[4]) & (g889) & (g871) & (g883)) + ((!g747) & (g744) & (!sk[4]) & (!g889) & (!g871) & (!g883)) + ((!g747) & (g744) & (!sk[4]) & (!g889) & (!g871) & (g883)) + ((!g747) & (g744) & (!sk[4]) & (!g889) & (g871) & (!g883)) + ((!g747) & (g744) & (!sk[4]) & (!g889) & (g871) & (g883)) + ((!g747) & (g744) & (!sk[4]) & (g889) & (!g871) & (!g883)) + ((!g747) & (g744) & (!sk[4]) & (g889) & (!g871) & (g883)) + ((!g747) & (g744) & (!sk[4]) & (g889) & (g871) & (!g883)) + ((!g747) & (g744) & (!sk[4]) & (g889) & (g871) & (g883)) + ((!g747) & (g744) & (sk[4]) & (!g889) & (!g871) & (!g883)) + ((!g747) & (g744) & (sk[4]) & (!g889) & (g871) & (g883)) + ((!g747) & (g744) & (sk[4]) & (g889) & (!g871) & (!g883)) + ((!g747) & (g744) & (sk[4]) & (g889) & (g871) & (g883)) + ((g747) & (!g744) & (!sk[4]) & (!g889) & (g871) & (!g883)) + ((g747) & (!g744) & (!sk[4]) & (!g889) & (g871) & (g883)) + ((g747) & (!g744) & (!sk[4]) & (g889) & (!g871) & (!g883)) + ((g747) & (!g744) & (!sk[4]) & (g889) & (!g871) & (g883)) + ((g747) & (!g744) & (!sk[4]) & (g889) & (g871) & (!g883)) + ((g747) & (!g744) & (!sk[4]) & (g889) & (g871) & (g883)) + ((g747) & (!g744) & (sk[4]) & (!g889) & (!g871) & (!g883)) + ((g747) & (!g744) & (sk[4]) & (!g889) & (!g871) & (g883)) + ((g747) & (!g744) & (sk[4]) & (!g889) & (g871) & (!g883)) + ((g747) & (!g744) & (sk[4]) & (g889) & (g871) & (g883)) + ((g747) & (g744) & (!sk[4]) & (!g889) & (!g871) & (!g883)) + ((g747) & (g744) & (!sk[4]) & (!g889) & (!g871) & (g883)) + ((g747) & (g744) & (!sk[4]) & (!g889) & (g871) & (!g883)) + ((g747) & (g744) & (!sk[4]) & (!g889) & (g871) & (g883)) + ((g747) & (g744) & (!sk[4]) & (g889) & (!g871) & (!g883)) + ((g747) & (g744) & (!sk[4]) & (g889) & (!g871) & (g883)) + ((g747) & (g744) & (!sk[4]) & (g889) & (g871) & (!g883)) + ((g747) & (g744) & (!sk[4]) & (g889) & (g871) & (g883)) + ((g747) & (g744) & (sk[4]) & (!g889) & (!g871) & (!g883)) + ((g747) & (g744) & (sk[4]) & (!g889) & (!g871) & (g883)) + ((g747) & (g744) & (sk[4]) & (!g889) & (g871) & (!g883)) + ((g747) & (g744) & (sk[4]) & (!g889) & (g871) & (g883)) + ((g747) & (g744) & (sk[4]) & (g889) & (!g871) & (!g883)) + ((g747) & (g744) & (sk[4]) & (g889) & (g871) & (g883)));
	assign g1147 = (((!g200) & (!g742) & (!g884) & (!g890) & (!g1145) & (g1146)) + ((!g200) & (!g742) & (!g884) & (!g890) & (g1145) & (!g1146)) + ((!g200) & (!g742) & (!g884) & (!g890) & (g1145) & (g1146)) + ((!g200) & (!g742) & (!g884) & (g890) & (!g1145) & (g1146)) + ((!g200) & (!g742) & (!g884) & (g890) & (g1145) & (!g1146)) + ((!g200) & (!g742) & (!g884) & (g890) & (g1145) & (g1146)) + ((!g200) & (!g742) & (g884) & (!g890) & (!g1145) & (g1146)) + ((!g200) & (!g742) & (g884) & (!g890) & (g1145) & (!g1146)) + ((!g200) & (!g742) & (g884) & (!g890) & (g1145) & (g1146)) + ((!g200) & (!g742) & (g884) & (g890) & (!g1145) & (g1146)) + ((!g200) & (!g742) & (g884) & (g890) & (g1145) & (!g1146)) + ((!g200) & (!g742) & (g884) & (g890) & (g1145) & (g1146)) + ((!g200) & (g742) & (!g884) & (!g890) & (!g1145) & (!g1146)) + ((!g200) & (g742) & (!g884) & (!g890) & (!g1145) & (g1146)) + ((!g200) & (g742) & (!g884) & (!g890) & (g1145) & (!g1146)) + ((!g200) & (g742) & (!g884) & (!g890) & (g1145) & (g1146)) + ((!g200) & (g742) & (!g884) & (g890) & (!g1145) & (g1146)) + ((!g200) & (g742) & (!g884) & (g890) & (g1145) & (!g1146)) + ((!g200) & (g742) & (!g884) & (g890) & (g1145) & (g1146)) + ((!g200) & (g742) & (g884) & (!g890) & (!g1145) & (g1146)) + ((!g200) & (g742) & (g884) & (!g890) & (g1145) & (!g1146)) + ((!g200) & (g742) & (g884) & (!g890) & (g1145) & (g1146)) + ((!g200) & (g742) & (g884) & (g890) & (!g1145) & (!g1146)) + ((!g200) & (g742) & (g884) & (g890) & (!g1145) & (g1146)) + ((!g200) & (g742) & (g884) & (g890) & (g1145) & (!g1146)) + ((!g200) & (g742) & (g884) & (g890) & (g1145) & (g1146)) + ((g200) & (!g742) & (!g884) & (!g890) & (!g1145) & (!g1146)) + ((g200) & (!g742) & (!g884) & (g890) & (!g1145) & (!g1146)) + ((g200) & (!g742) & (g884) & (!g890) & (!g1145) & (!g1146)) + ((g200) & (!g742) & (g884) & (g890) & (!g1145) & (!g1146)) + ((g200) & (g742) & (!g884) & (g890) & (!g1145) & (!g1146)) + ((g200) & (g742) & (g884) & (!g890) & (!g1145) & (!g1146)));
	assign g1148 = (((!g1144) & (sk[6]) & (g1147)) + ((g1144) & (!sk[6]) & (g1147)) + ((g1144) & (sk[6]) & (!g1147)));
	assign g1149 = (((!g733) & (!g734) & (!g994) & (!sk[7]) & (g1040)) + ((!g733) & (!g734) & (g994) & (!sk[7]) & (g1040)) + ((!g733) & (g734) & (!g994) & (!sk[7]) & (g1040)) + ((!g733) & (g734) & (g994) & (!sk[7]) & (g1040)) + ((!g733) & (g734) & (g994) & (sk[7]) & (!g1040)) + ((!g733) & (g734) & (g994) & (sk[7]) & (g1040)) + ((g733) & (!g734) & (!g994) & (!sk[7]) & (!g1040)) + ((g733) & (!g734) & (!g994) & (!sk[7]) & (g1040)) + ((g733) & (!g734) & (!g994) & (sk[7]) & (!g1040)) + ((g733) & (!g734) & (g994) & (!sk[7]) & (!g1040)) + ((g733) & (!g734) & (g994) & (!sk[7]) & (g1040)) + ((g733) & (!g734) & (g994) & (sk[7]) & (!g1040)) + ((g733) & (g734) & (!g994) & (!sk[7]) & (!g1040)) + ((g733) & (g734) & (!g994) & (!sk[7]) & (g1040)) + ((g733) & (g734) & (!g994) & (sk[7]) & (!g1040)) + ((g733) & (g734) & (g994) & (!sk[7]) & (!g1040)) + ((g733) & (g734) & (g994) & (!sk[7]) & (g1040)) + ((g733) & (g734) & (g994) & (sk[7]) & (!g1040)) + ((g733) & (g734) & (g994) & (sk[7]) & (g1040)));
	assign g1150 = (((!g2) & (!g686) & (!g732) & (!g971) & (!g1041) & (!g1149)) + ((!g2) & (!g686) & (!g732) & (!g971) & (g1041) & (!g1149)) + ((!g2) & (!g686) & (!g732) & (g971) & (!g1041) & (!g1149)) + ((!g2) & (!g686) & (!g732) & (g971) & (g1041) & (!g1149)) + ((!g2) & (!g686) & (g732) & (!g971) & (g1041) & (!g1149)) + ((!g2) & (!g686) & (g732) & (g971) & (g1041) & (!g1149)) + ((!g2) & (g686) & (!g732) & (!g971) & (!g1041) & (!g1149)) + ((!g2) & (g686) & (!g732) & (!g971) & (g1041) & (!g1149)) + ((!g2) & (g686) & (g732) & (!g971) & (g1041) & (!g1149)) + ((g2) & (!g686) & (!g732) & (!g971) & (!g1041) & (g1149)) + ((g2) & (!g686) & (!g732) & (!g971) & (g1041) & (g1149)) + ((g2) & (!g686) & (!g732) & (g971) & (!g1041) & (g1149)) + ((g2) & (!g686) & (!g732) & (g971) & (g1041) & (g1149)) + ((g2) & (!g686) & (g732) & (!g971) & (!g1041) & (!g1149)) + ((g2) & (!g686) & (g732) & (!g971) & (!g1041) & (g1149)) + ((g2) & (!g686) & (g732) & (!g971) & (g1041) & (g1149)) + ((g2) & (!g686) & (g732) & (g971) & (!g1041) & (!g1149)) + ((g2) & (!g686) & (g732) & (g971) & (!g1041) & (g1149)) + ((g2) & (!g686) & (g732) & (g971) & (g1041) & (g1149)) + ((g2) & (g686) & (!g732) & (!g971) & (!g1041) & (g1149)) + ((g2) & (g686) & (!g732) & (!g971) & (g1041) & (g1149)) + ((g2) & (g686) & (!g732) & (g971) & (!g1041) & (!g1149)) + ((g2) & (g686) & (!g732) & (g971) & (!g1041) & (g1149)) + ((g2) & (g686) & (!g732) & (g971) & (g1041) & (!g1149)) + ((g2) & (g686) & (!g732) & (g971) & (g1041) & (g1149)) + ((g2) & (g686) & (g732) & (!g971) & (!g1041) & (!g1149)) + ((g2) & (g686) & (g732) & (!g971) & (!g1041) & (g1149)) + ((g2) & (g686) & (g732) & (!g971) & (g1041) & (g1149)) + ((g2) & (g686) & (g732) & (g971) & (!g1041) & (!g1149)) + ((g2) & (g686) & (g732) & (g971) & (!g1041) & (g1149)) + ((g2) & (g686) & (g732) & (g971) & (g1041) & (!g1149)) + ((g2) & (g686) & (g732) & (g971) & (g1041) & (g1149)));
	assign g1151 = (((!g683) & (!g864) & (g868) & (!g1040) & (!g1079) & (!g1080)) + ((!g683) & (!g864) & (g868) & (!g1040) & (!g1079) & (g1080)) + ((!g683) & (!g864) & (g868) & (g1040) & (!g1079) & (g1080)) + ((!g683) & (g864) & (!g868) & (!g1040) & (!g1079) & (!g1080)) + ((!g683) & (g864) & (!g868) & (!g1040) & (!g1079) & (g1080)) + ((!g683) & (g864) & (!g868) & (g1040) & (!g1079) & (!g1080)) + ((!g683) & (g864) & (!g868) & (g1040) & (!g1079) & (g1080)) + ((!g683) & (g864) & (g868) & (!g1040) & (!g1079) & (!g1080)) + ((!g683) & (g864) & (g868) & (!g1040) & (!g1079) & (g1080)) + ((!g683) & (g864) & (g868) & (g1040) & (!g1079) & (!g1080)) + ((!g683) & (g864) & (g868) & (g1040) & (!g1079) & (g1080)) + ((g683) & (!g864) & (!g868) & (!g1040) & (!g1079) & (!g1080)) + ((g683) & (!g864) & (!g868) & (!g1040) & (!g1079) & (g1080)) + ((g683) & (!g864) & (!g868) & (!g1040) & (g1079) & (!g1080)) + ((g683) & (!g864) & (!g868) & (!g1040) & (g1079) & (g1080)) + ((g683) & (!g864) & (!g868) & (g1040) & (!g1079) & (!g1080)) + ((g683) & (!g864) & (!g868) & (g1040) & (!g1079) & (g1080)) + ((g683) & (!g864) & (!g868) & (g1040) & (g1079) & (!g1080)) + ((g683) & (!g864) & (!g868) & (g1040) & (g1079) & (g1080)) + ((g683) & (!g864) & (g868) & (!g1040) & (g1079) & (!g1080)) + ((g683) & (!g864) & (g868) & (!g1040) & (g1079) & (g1080)) + ((g683) & (!g864) & (g868) & (g1040) & (!g1079) & (!g1080)) + ((g683) & (!g864) & (g868) & (g1040) & (g1079) & (!g1080)) + ((g683) & (!g864) & (g868) & (g1040) & (g1079) & (g1080)) + ((g683) & (g864) & (!g868) & (!g1040) & (g1079) & (!g1080)) + ((g683) & (g864) & (!g868) & (!g1040) & (g1079) & (g1080)) + ((g683) & (g864) & (!g868) & (g1040) & (g1079) & (!g1080)) + ((g683) & (g864) & (!g868) & (g1040) & (g1079) & (g1080)) + ((g683) & (g864) & (g868) & (!g1040) & (g1079) & (!g1080)) + ((g683) & (g864) & (g868) & (!g1040) & (g1079) & (g1080)) + ((g683) & (g864) & (g868) & (g1040) & (g1079) & (!g1080)) + ((g683) & (g864) & (g868) & (g1040) & (g1079) & (g1080)));
	assign g1152 = (((!g1137) & (!sk[10]) & (!g1148) & (!g1150) & (g1151)) + ((!g1137) & (!sk[10]) & (!g1148) & (g1150) & (g1151)) + ((!g1137) & (!sk[10]) & (g1148) & (!g1150) & (g1151)) + ((!g1137) & (!sk[10]) & (g1148) & (g1150) & (g1151)) + ((!g1137) & (sk[10]) & (!g1148) & (!g1150) & (g1151)) + ((!g1137) & (sk[10]) & (!g1148) & (g1150) & (!g1151)) + ((!g1137) & (sk[10]) & (g1148) & (!g1150) & (!g1151)) + ((!g1137) & (sk[10]) & (g1148) & (g1150) & (g1151)) + ((g1137) & (!sk[10]) & (!g1148) & (!g1150) & (!g1151)) + ((g1137) & (!sk[10]) & (!g1148) & (!g1150) & (g1151)) + ((g1137) & (!sk[10]) & (!g1148) & (g1150) & (!g1151)) + ((g1137) & (!sk[10]) & (!g1148) & (g1150) & (g1151)) + ((g1137) & (!sk[10]) & (g1148) & (!g1150) & (!g1151)) + ((g1137) & (!sk[10]) & (g1148) & (!g1150) & (g1151)) + ((g1137) & (!sk[10]) & (g1148) & (g1150) & (!g1151)) + ((g1137) & (!sk[10]) & (g1148) & (g1150) & (g1151)) + ((g1137) & (sk[10]) & (!g1148) & (!g1150) & (!g1151)) + ((g1137) & (sk[10]) & (!g1148) & (g1150) & (g1151)) + ((g1137) & (sk[10]) & (g1148) & (!g1150) & (g1151)) + ((g1137) & (sk[10]) & (g1148) & (g1150) & (!g1151)));
	assign g1153 = (((!g1108) & (!g1109) & (!g1111) & (!g1125) & (!g1136) & (g1152)) + ((!g1108) & (!g1109) & (!g1111) & (!g1125) & (g1136) & (!g1152)) + ((!g1108) & (!g1109) & (!g1111) & (g1125) & (!g1136) & (g1152)) + ((!g1108) & (!g1109) & (!g1111) & (g1125) & (g1136) & (!g1152)) + ((!g1108) & (!g1109) & (g1111) & (!g1125) & (!g1136) & (g1152)) + ((!g1108) & (!g1109) & (g1111) & (!g1125) & (g1136) & (!g1152)) + ((!g1108) & (!g1109) & (g1111) & (g1125) & (!g1136) & (!g1152)) + ((!g1108) & (!g1109) & (g1111) & (g1125) & (g1136) & (g1152)) + ((!g1108) & (g1109) & (!g1111) & (!g1125) & (!g1136) & (g1152)) + ((!g1108) & (g1109) & (!g1111) & (!g1125) & (g1136) & (!g1152)) + ((!g1108) & (g1109) & (!g1111) & (g1125) & (!g1136) & (!g1152)) + ((!g1108) & (g1109) & (!g1111) & (g1125) & (g1136) & (g1152)) + ((!g1108) & (g1109) & (g1111) & (!g1125) & (!g1136) & (!g1152)) + ((!g1108) & (g1109) & (g1111) & (!g1125) & (g1136) & (g1152)) + ((!g1108) & (g1109) & (g1111) & (g1125) & (!g1136) & (!g1152)) + ((!g1108) & (g1109) & (g1111) & (g1125) & (g1136) & (g1152)) + ((g1108) & (!g1109) & (!g1111) & (!g1125) & (!g1136) & (g1152)) + ((g1108) & (!g1109) & (!g1111) & (!g1125) & (g1136) & (!g1152)) + ((g1108) & (!g1109) & (!g1111) & (g1125) & (!g1136) & (!g1152)) + ((g1108) & (!g1109) & (!g1111) & (g1125) & (g1136) & (g1152)) + ((g1108) & (!g1109) & (g1111) & (!g1125) & (!g1136) & (!g1152)) + ((g1108) & (!g1109) & (g1111) & (!g1125) & (g1136) & (g1152)) + ((g1108) & (!g1109) & (g1111) & (g1125) & (!g1136) & (!g1152)) + ((g1108) & (!g1109) & (g1111) & (g1125) & (g1136) & (g1152)) + ((g1108) & (g1109) & (!g1111) & (!g1125) & (!g1136) & (g1152)) + ((g1108) & (g1109) & (!g1111) & (!g1125) & (g1136) & (!g1152)) + ((g1108) & (g1109) & (!g1111) & (g1125) & (!g1136) & (!g1152)) + ((g1108) & (g1109) & (!g1111) & (g1125) & (g1136) & (g1152)) + ((g1108) & (g1109) & (g1111) & (!g1125) & (!g1136) & (!g1152)) + ((g1108) & (g1109) & (g1111) & (!g1125) & (g1136) & (g1152)) + ((g1108) & (g1109) & (g1111) & (g1125) & (!g1136) & (!g1152)) + ((g1108) & (g1109) & (g1111) & (g1125) & (g1136) & (g1152)));
	assign g1154 = (((!g114) & (!g115) & (!sk[12]) & (!g8) & (g17) & (!g66)) + ((!g114) & (!g115) & (!sk[12]) & (!g8) & (g17) & (g66)) + ((!g114) & (!g115) & (!sk[12]) & (g8) & (!g17) & (!g66)) + ((!g114) & (!g115) & (!sk[12]) & (g8) & (!g17) & (g66)) + ((!g114) & (!g115) & (!sk[12]) & (g8) & (g17) & (!g66)) + ((!g114) & (!g115) & (!sk[12]) & (g8) & (g17) & (g66)) + ((!g114) & (!g115) & (sk[12]) & (g8) & (!g17) & (g66)) + ((!g114) & (!g115) & (sk[12]) & (g8) & (g17) & (g66)) + ((!g114) & (g115) & (!sk[12]) & (!g8) & (!g17) & (!g66)) + ((!g114) & (g115) & (!sk[12]) & (!g8) & (!g17) & (g66)) + ((!g114) & (g115) & (!sk[12]) & (!g8) & (g17) & (!g66)) + ((!g114) & (g115) & (!sk[12]) & (!g8) & (g17) & (g66)) + ((!g114) & (g115) & (!sk[12]) & (g8) & (!g17) & (!g66)) + ((!g114) & (g115) & (!sk[12]) & (g8) & (!g17) & (g66)) + ((!g114) & (g115) & (!sk[12]) & (g8) & (g17) & (!g66)) + ((!g114) & (g115) & (!sk[12]) & (g8) & (g17) & (g66)) + ((g114) & (!g115) & (!sk[12]) & (!g8) & (g17) & (!g66)) + ((g114) & (!g115) & (!sk[12]) & (!g8) & (g17) & (g66)) + ((g114) & (!g115) & (!sk[12]) & (g8) & (!g17) & (!g66)) + ((g114) & (!g115) & (!sk[12]) & (g8) & (!g17) & (g66)) + ((g114) & (!g115) & (!sk[12]) & (g8) & (g17) & (!g66)) + ((g114) & (!g115) & (!sk[12]) & (g8) & (g17) & (g66)) + ((g114) & (!g115) & (sk[12]) & (!g8) & (!g17) & (g66)) + ((g114) & (!g115) & (sk[12]) & (!g8) & (g17) & (!g66)) + ((g114) & (!g115) & (sk[12]) & (!g8) & (g17) & (g66)) + ((g114) & (g115) & (!sk[12]) & (!g8) & (!g17) & (!g66)) + ((g114) & (g115) & (!sk[12]) & (!g8) & (!g17) & (g66)) + ((g114) & (g115) & (!sk[12]) & (!g8) & (g17) & (!g66)) + ((g114) & (g115) & (!sk[12]) & (!g8) & (g17) & (g66)) + ((g114) & (g115) & (!sk[12]) & (g8) & (!g17) & (!g66)) + ((g114) & (g115) & (!sk[12]) & (g8) & (!g17) & (g66)) + ((g114) & (g115) & (!sk[12]) & (g8) & (g17) & (!g66)) + ((g114) & (g115) & (!sk[12]) & (g8) & (g17) & (g66)) + ((g114) & (g115) & (sk[12]) & (!g8) & (g17) & (!g66)) + ((g114) & (g115) & (sk[12]) & (!g8) & (g17) & (g66)));
	assign g1155 = (((!g246) & (!sk[13]) & (!g1018) & (!g1100) & (g1154)) + ((!g246) & (!sk[13]) & (!g1018) & (g1100) & (g1154)) + ((!g246) & (!sk[13]) & (g1018) & (!g1100) & (g1154)) + ((!g246) & (!sk[13]) & (g1018) & (g1100) & (g1154)) + ((g246) & (!sk[13]) & (!g1018) & (!g1100) & (!g1154)) + ((g246) & (!sk[13]) & (!g1018) & (!g1100) & (g1154)) + ((g246) & (!sk[13]) & (!g1018) & (g1100) & (!g1154)) + ((g246) & (!sk[13]) & (!g1018) & (g1100) & (g1154)) + ((g246) & (!sk[13]) & (g1018) & (!g1100) & (!g1154)) + ((g246) & (!sk[13]) & (g1018) & (!g1100) & (g1154)) + ((g246) & (!sk[13]) & (g1018) & (g1100) & (!g1154)) + ((g246) & (!sk[13]) & (g1018) & (g1100) & (g1154)) + ((g246) & (sk[13]) & (g1018) & (g1100) & (!g1154)));
	assign g1156 = (((!g111) & (!g574) & (!sk[14]) & (!g711) & (g857) & (!g1155)) + ((!g111) & (!g574) & (!sk[14]) & (!g711) & (g857) & (g1155)) + ((!g111) & (!g574) & (!sk[14]) & (g711) & (!g857) & (!g1155)) + ((!g111) & (!g574) & (!sk[14]) & (g711) & (!g857) & (g1155)) + ((!g111) & (!g574) & (!sk[14]) & (g711) & (g857) & (!g1155)) + ((!g111) & (!g574) & (!sk[14]) & (g711) & (g857) & (g1155)) + ((!g111) & (g574) & (!sk[14]) & (!g711) & (!g857) & (!g1155)) + ((!g111) & (g574) & (!sk[14]) & (!g711) & (!g857) & (g1155)) + ((!g111) & (g574) & (!sk[14]) & (!g711) & (g857) & (!g1155)) + ((!g111) & (g574) & (!sk[14]) & (!g711) & (g857) & (g1155)) + ((!g111) & (g574) & (!sk[14]) & (g711) & (!g857) & (!g1155)) + ((!g111) & (g574) & (!sk[14]) & (g711) & (!g857) & (g1155)) + ((!g111) & (g574) & (!sk[14]) & (g711) & (g857) & (!g1155)) + ((!g111) & (g574) & (!sk[14]) & (g711) & (g857) & (g1155)) + ((g111) & (!g574) & (!sk[14]) & (!g711) & (g857) & (!g1155)) + ((g111) & (!g574) & (!sk[14]) & (!g711) & (g857) & (g1155)) + ((g111) & (!g574) & (!sk[14]) & (g711) & (!g857) & (!g1155)) + ((g111) & (!g574) & (!sk[14]) & (g711) & (!g857) & (g1155)) + ((g111) & (!g574) & (!sk[14]) & (g711) & (g857) & (!g1155)) + ((g111) & (!g574) & (!sk[14]) & (g711) & (g857) & (g1155)) + ((g111) & (g574) & (!sk[14]) & (!g711) & (!g857) & (!g1155)) + ((g111) & (g574) & (!sk[14]) & (!g711) & (!g857) & (g1155)) + ((g111) & (g574) & (!sk[14]) & (!g711) & (g857) & (!g1155)) + ((g111) & (g574) & (!sk[14]) & (!g711) & (g857) & (g1155)) + ((g111) & (g574) & (!sk[14]) & (g711) & (!g857) & (!g1155)) + ((g111) & (g574) & (!sk[14]) & (g711) & (!g857) & (g1155)) + ((g111) & (g574) & (!sk[14]) & (g711) & (g857) & (!g1155)) + ((g111) & (g574) & (!sk[14]) & (g711) & (g857) & (g1155)) + ((g111) & (g574) & (sk[14]) & (g711) & (g857) & (g1155)));
	assign g1157 = (((!g1126) & (!g1131) & (!sk[15]) & (!g1132) & (g1153) & (!g1156)) + ((!g1126) & (!g1131) & (!sk[15]) & (!g1132) & (g1153) & (g1156)) + ((!g1126) & (!g1131) & (!sk[15]) & (g1132) & (!g1153) & (!g1156)) + ((!g1126) & (!g1131) & (!sk[15]) & (g1132) & (!g1153) & (g1156)) + ((!g1126) & (!g1131) & (!sk[15]) & (g1132) & (g1153) & (!g1156)) + ((!g1126) & (!g1131) & (!sk[15]) & (g1132) & (g1153) & (g1156)) + ((!g1126) & (!g1131) & (sk[15]) & (!g1132) & (!g1153) & (!g1156)) + ((!g1126) & (!g1131) & (sk[15]) & (!g1132) & (g1153) & (g1156)) + ((!g1126) & (!g1131) & (sk[15]) & (g1132) & (!g1153) & (g1156)) + ((!g1126) & (!g1131) & (sk[15]) & (g1132) & (g1153) & (!g1156)) + ((!g1126) & (g1131) & (!sk[15]) & (!g1132) & (!g1153) & (!g1156)) + ((!g1126) & (g1131) & (!sk[15]) & (!g1132) & (!g1153) & (g1156)) + ((!g1126) & (g1131) & (!sk[15]) & (!g1132) & (g1153) & (!g1156)) + ((!g1126) & (g1131) & (!sk[15]) & (!g1132) & (g1153) & (g1156)) + ((!g1126) & (g1131) & (!sk[15]) & (g1132) & (!g1153) & (!g1156)) + ((!g1126) & (g1131) & (!sk[15]) & (g1132) & (!g1153) & (g1156)) + ((!g1126) & (g1131) & (!sk[15]) & (g1132) & (g1153) & (!g1156)) + ((!g1126) & (g1131) & (!sk[15]) & (g1132) & (g1153) & (g1156)) + ((!g1126) & (g1131) & (sk[15]) & (!g1132) & (!g1153) & (!g1156)) + ((!g1126) & (g1131) & (sk[15]) & (!g1132) & (g1153) & (g1156)) + ((!g1126) & (g1131) & (sk[15]) & (g1132) & (!g1153) & (!g1156)) + ((!g1126) & (g1131) & (sk[15]) & (g1132) & (g1153) & (g1156)) + ((g1126) & (!g1131) & (!sk[15]) & (!g1132) & (g1153) & (!g1156)) + ((g1126) & (!g1131) & (!sk[15]) & (!g1132) & (g1153) & (g1156)) + ((g1126) & (!g1131) & (!sk[15]) & (g1132) & (!g1153) & (!g1156)) + ((g1126) & (!g1131) & (!sk[15]) & (g1132) & (!g1153) & (g1156)) + ((g1126) & (!g1131) & (!sk[15]) & (g1132) & (g1153) & (!g1156)) + ((g1126) & (!g1131) & (!sk[15]) & (g1132) & (g1153) & (g1156)) + ((g1126) & (!g1131) & (sk[15]) & (!g1132) & (!g1153) & (g1156)) + ((g1126) & (!g1131) & (sk[15]) & (!g1132) & (g1153) & (!g1156)) + ((g1126) & (!g1131) & (sk[15]) & (g1132) & (!g1153) & (g1156)) + ((g1126) & (!g1131) & (sk[15]) & (g1132) & (g1153) & (!g1156)) + ((g1126) & (g1131) & (!sk[15]) & (!g1132) & (!g1153) & (!g1156)) + ((g1126) & (g1131) & (!sk[15]) & (!g1132) & (!g1153) & (g1156)) + ((g1126) & (g1131) & (!sk[15]) & (!g1132) & (g1153) & (!g1156)) + ((g1126) & (g1131) & (!sk[15]) & (!g1132) & (g1153) & (g1156)) + ((g1126) & (g1131) & (!sk[15]) & (g1132) & (!g1153) & (!g1156)) + ((g1126) & (g1131) & (!sk[15]) & (g1132) & (!g1153) & (g1156)) + ((g1126) & (g1131) & (!sk[15]) & (g1132) & (g1153) & (!g1156)) + ((g1126) & (g1131) & (!sk[15]) & (g1132) & (g1153) & (g1156)) + ((g1126) & (g1131) & (sk[15]) & (!g1132) & (!g1153) & (!g1156)) + ((g1126) & (g1131) & (sk[15]) & (!g1132) & (g1153) & (g1156)) + ((g1126) & (g1131) & (sk[15]) & (g1132) & (!g1153) & (g1156)) + ((g1126) & (g1131) & (sk[15]) & (g1132) & (g1153) & (!g1156)));
	assign g1158 = (((g1067) & (!g1069) & (!g1106) & (!g1126) & (!g1131) & (g1132)) + ((g1067) & (!g1069) & (!g1106) & (!g1126) & (g1131) & (!g1132)) + ((g1067) & (!g1069) & (!g1106) & (g1126) & (!g1131) & (!g1132)) + ((g1067) & (!g1069) & (!g1106) & (g1126) & (g1131) & (g1132)) + ((g1067) & (g1069) & (g1106) & (!g1126) & (!g1131) & (!g1132)) + ((g1067) & (g1069) & (g1106) & (!g1126) & (g1131) & (g1132)) + ((g1067) & (g1069) & (g1106) & (g1126) & (!g1131) & (g1132)) + ((g1067) & (g1069) & (g1106) & (g1126) & (g1131) & (!g1132)));
	assign sinx3x = (((!g1068) & (!g1135) & (!sk[17]) & (!g1157) & (g1158)) + ((!g1068) & (!g1135) & (!sk[17]) & (g1157) & (g1158)) + ((!g1068) & (!g1135) & (sk[17]) & (g1157) & (!g1158)) + ((!g1068) & (!g1135) & (sk[17]) & (g1157) & (g1158)) + ((!g1068) & (g1135) & (!sk[17]) & (!g1157) & (g1158)) + ((!g1068) & (g1135) & (!sk[17]) & (g1157) & (g1158)) + ((!g1068) & (g1135) & (sk[17]) & (!g1157) & (!g1158)) + ((!g1068) & (g1135) & (sk[17]) & (!g1157) & (g1158)) + ((g1068) & (!g1135) & (!sk[17]) & (!g1157) & (!g1158)) + ((g1068) & (!g1135) & (!sk[17]) & (!g1157) & (g1158)) + ((g1068) & (!g1135) & (!sk[17]) & (g1157) & (!g1158)) + ((g1068) & (!g1135) & (!sk[17]) & (g1157) & (g1158)) + ((g1068) & (!g1135) & (sk[17]) & (!g1157) & (!g1158)) + ((g1068) & (!g1135) & (sk[17]) & (g1157) & (g1158)) + ((g1068) & (g1135) & (!sk[17]) & (!g1157) & (!g1158)) + ((g1068) & (g1135) & (!sk[17]) & (!g1157) & (g1158)) + ((g1068) & (g1135) & (!sk[17]) & (g1157) & (!g1158)) + ((g1068) & (g1135) & (!sk[17]) & (g1157) & (g1158)) + ((g1068) & (g1135) & (sk[17]) & (!g1157) & (g1158)) + ((g1068) & (g1135) & (sk[17]) & (g1157) & (!g1158)));
	assign g1160 = (((!g1126) & (!sk[18]) & (!g1131) & (!g1132) & (g1153) & (!g1156)) + ((!g1126) & (!sk[18]) & (!g1131) & (!g1132) & (g1153) & (g1156)) + ((!g1126) & (!sk[18]) & (!g1131) & (g1132) & (!g1153) & (!g1156)) + ((!g1126) & (!sk[18]) & (!g1131) & (g1132) & (!g1153) & (g1156)) + ((!g1126) & (!sk[18]) & (!g1131) & (g1132) & (g1153) & (!g1156)) + ((!g1126) & (!sk[18]) & (!g1131) & (g1132) & (g1153) & (g1156)) + ((!g1126) & (!sk[18]) & (g1131) & (!g1132) & (!g1153) & (!g1156)) + ((!g1126) & (!sk[18]) & (g1131) & (!g1132) & (!g1153) & (g1156)) + ((!g1126) & (!sk[18]) & (g1131) & (!g1132) & (g1153) & (!g1156)) + ((!g1126) & (!sk[18]) & (g1131) & (!g1132) & (g1153) & (g1156)) + ((!g1126) & (!sk[18]) & (g1131) & (g1132) & (!g1153) & (!g1156)) + ((!g1126) & (!sk[18]) & (g1131) & (g1132) & (!g1153) & (g1156)) + ((!g1126) & (!sk[18]) & (g1131) & (g1132) & (g1153) & (!g1156)) + ((!g1126) & (!sk[18]) & (g1131) & (g1132) & (g1153) & (g1156)) + ((!g1126) & (sk[18]) & (!g1131) & (!g1132) & (g1153) & (!g1156)) + ((!g1126) & (sk[18]) & (!g1131) & (g1132) & (!g1153) & (!g1156)) + ((!g1126) & (sk[18]) & (!g1131) & (g1132) & (g1153) & (!g1156)) + ((!g1126) & (sk[18]) & (!g1131) & (g1132) & (g1153) & (g1156)) + ((!g1126) & (sk[18]) & (g1131) & (!g1132) & (g1153) & (!g1156)) + ((!g1126) & (sk[18]) & (g1131) & (g1132) & (g1153) & (!g1156)) + ((g1126) & (!sk[18]) & (!g1131) & (!g1132) & (g1153) & (!g1156)) + ((g1126) & (!sk[18]) & (!g1131) & (!g1132) & (g1153) & (g1156)) + ((g1126) & (!sk[18]) & (!g1131) & (g1132) & (!g1153) & (!g1156)) + ((g1126) & (!sk[18]) & (!g1131) & (g1132) & (!g1153) & (g1156)) + ((g1126) & (!sk[18]) & (!g1131) & (g1132) & (g1153) & (!g1156)) + ((g1126) & (!sk[18]) & (!g1131) & (g1132) & (g1153) & (g1156)) + ((g1126) & (!sk[18]) & (g1131) & (!g1132) & (!g1153) & (!g1156)) + ((g1126) & (!sk[18]) & (g1131) & (!g1132) & (!g1153) & (g1156)) + ((g1126) & (!sk[18]) & (g1131) & (!g1132) & (g1153) & (!g1156)) + ((g1126) & (!sk[18]) & (g1131) & (!g1132) & (g1153) & (g1156)) + ((g1126) & (!sk[18]) & (g1131) & (g1132) & (!g1153) & (!g1156)) + ((g1126) & (!sk[18]) & (g1131) & (g1132) & (!g1153) & (g1156)) + ((g1126) & (!sk[18]) & (g1131) & (g1132) & (g1153) & (!g1156)) + ((g1126) & (!sk[18]) & (g1131) & (g1132) & (g1153) & (g1156)) + ((g1126) & (sk[18]) & (!g1131) & (!g1132) & (!g1153) & (!g1156)) + ((g1126) & (sk[18]) & (!g1131) & (!g1132) & (g1153) & (!g1156)) + ((g1126) & (sk[18]) & (!g1131) & (!g1132) & (g1153) & (g1156)) + ((g1126) & (sk[18]) & (!g1131) & (g1132) & (!g1153) & (!g1156)) + ((g1126) & (sk[18]) & (!g1131) & (g1132) & (g1153) & (!g1156)) + ((g1126) & (sk[18]) & (!g1131) & (g1132) & (g1153) & (g1156)) + ((g1126) & (sk[18]) & (g1131) & (!g1132) & (g1153) & (!g1156)) + ((g1126) & (sk[18]) & (g1131) & (g1132) & (!g1153) & (!g1156)) + ((g1126) & (sk[18]) & (g1131) & (g1132) & (g1153) & (!g1156)) + ((g1126) & (sk[18]) & (g1131) & (g1132) & (g1153) & (g1156)));
	assign g1161 = (((!g1108) & (!g1109) & (!g1111) & (!g1125) & (!g1136) & (!g1152)) + ((!g1108) & (!g1109) & (!g1111) & (!g1125) & (!g1136) & (g1152)) + ((!g1108) & (!g1109) & (!g1111) & (!g1125) & (g1136) & (!g1152)) + ((!g1108) & (!g1109) & (!g1111) & (g1125) & (!g1136) & (!g1152)) + ((!g1108) & (!g1109) & (!g1111) & (g1125) & (!g1136) & (g1152)) + ((!g1108) & (!g1109) & (!g1111) & (g1125) & (g1136) & (!g1152)) + ((!g1108) & (!g1109) & (g1111) & (!g1125) & (!g1136) & (!g1152)) + ((!g1108) & (!g1109) & (g1111) & (!g1125) & (!g1136) & (g1152)) + ((!g1108) & (!g1109) & (g1111) & (!g1125) & (g1136) & (!g1152)) + ((!g1108) & (!g1109) & (g1111) & (g1125) & (!g1136) & (!g1152)) + ((!g1108) & (g1109) & (!g1111) & (!g1125) & (!g1136) & (!g1152)) + ((!g1108) & (g1109) & (!g1111) & (!g1125) & (!g1136) & (g1152)) + ((!g1108) & (g1109) & (!g1111) & (!g1125) & (g1136) & (!g1152)) + ((!g1108) & (g1109) & (!g1111) & (g1125) & (!g1136) & (!g1152)) + ((!g1108) & (g1109) & (g1111) & (!g1125) & (!g1136) & (!g1152)) + ((!g1108) & (g1109) & (g1111) & (g1125) & (!g1136) & (!g1152)) + ((g1108) & (!g1109) & (!g1111) & (!g1125) & (!g1136) & (!g1152)) + ((g1108) & (!g1109) & (!g1111) & (!g1125) & (!g1136) & (g1152)) + ((g1108) & (!g1109) & (!g1111) & (!g1125) & (g1136) & (!g1152)) + ((g1108) & (!g1109) & (!g1111) & (g1125) & (!g1136) & (!g1152)) + ((g1108) & (!g1109) & (g1111) & (!g1125) & (!g1136) & (!g1152)) + ((g1108) & (!g1109) & (g1111) & (g1125) & (!g1136) & (!g1152)) + ((g1108) & (g1109) & (!g1111) & (!g1125) & (!g1136) & (!g1152)) + ((g1108) & (g1109) & (!g1111) & (!g1125) & (!g1136) & (g1152)) + ((g1108) & (g1109) & (!g1111) & (!g1125) & (g1136) & (!g1152)) + ((g1108) & (g1109) & (!g1111) & (g1125) & (!g1136) & (!g1152)) + ((g1108) & (g1109) & (g1111) & (!g1125) & (!g1136) & (!g1152)) + ((g1108) & (g1109) & (g1111) & (g1125) & (!g1136) & (!g1152)));
	assign g1162 = (((!g1137) & (!g1148) & (!sk[20]) & (!g1150) & (g1151)) + ((!g1137) & (!g1148) & (!sk[20]) & (g1150) & (g1151)) + ((!g1137) & (!g1148) & (sk[20]) & (!g1150) & (!g1151)) + ((!g1137) & (!g1148) & (sk[20]) & (!g1150) & (g1151)) + ((!g1137) & (!g1148) & (sk[20]) & (g1150) & (g1151)) + ((!g1137) & (g1148) & (!sk[20]) & (!g1150) & (g1151)) + ((!g1137) & (g1148) & (!sk[20]) & (g1150) & (g1151)) + ((!g1137) & (g1148) & (sk[20]) & (!g1150) & (g1151)) + ((g1137) & (!g1148) & (!sk[20]) & (!g1150) & (!g1151)) + ((g1137) & (!g1148) & (!sk[20]) & (!g1150) & (g1151)) + ((g1137) & (!g1148) & (!sk[20]) & (g1150) & (!g1151)) + ((g1137) & (!g1148) & (!sk[20]) & (g1150) & (g1151)) + ((g1137) & (!g1148) & (sk[20]) & (!g1150) & (g1151)) + ((g1137) & (g1148) & (!sk[20]) & (!g1150) & (!g1151)) + ((g1137) & (g1148) & (!sk[20]) & (!g1150) & (g1151)) + ((g1137) & (g1148) & (!sk[20]) & (g1150) & (!g1151)) + ((g1137) & (g1148) & (!sk[20]) & (g1150) & (g1151)) + ((g1137) & (g1148) & (sk[20]) & (!g1150) & (!g1151)) + ((g1137) & (g1148) & (sk[20]) & (!g1150) & (g1151)) + ((g1137) & (g1148) & (sk[20]) & (g1150) & (g1151)));
	assign g1163 = (((!g747) & (!g744) & (!g748) & (!g962) & (!g963) & (!g971)) + ((!g747) & (!g744) & (!g748) & (!g962) & (!g963) & (g971)) + ((!g747) & (!g744) & (!g748) & (!g962) & (g963) & (!g971)) + ((!g747) & (!g744) & (!g748) & (!g962) & (g963) & (g971)) + ((!g747) & (!g744) & (!g748) & (g962) & (!g963) & (!g971)) + ((!g747) & (!g744) & (!g748) & (g962) & (!g963) & (g971)) + ((!g747) & (!g744) & (!g748) & (g962) & (g963) & (!g971)) + ((!g747) & (!g744) & (!g748) & (g962) & (g963) & (g971)) + ((!g747) & (!g744) & (g748) & (!g962) & (!g963) & (!g971)) + ((!g747) & (!g744) & (g748) & (!g962) & (!g963) & (g971)) + ((!g747) & (!g744) & (g748) & (g962) & (!g963) & (!g971)) + ((!g747) & (!g744) & (g748) & (g962) & (!g963) & (g971)) + ((!g747) & (g744) & (!g748) & (g962) & (!g963) & (!g971)) + ((!g747) & (g744) & (!g748) & (g962) & (!g963) & (g971)) + ((!g747) & (g744) & (!g748) & (g962) & (g963) & (!g971)) + ((!g747) & (g744) & (!g748) & (g962) & (g963) & (g971)) + ((!g747) & (g744) & (g748) & (g962) & (!g963) & (!g971)) + ((!g747) & (g744) & (g748) & (g962) & (!g963) & (g971)) + ((g747) & (!g744) & (!g748) & (!g962) & (!g963) & (!g971)) + ((g747) & (!g744) & (!g748) & (!g962) & (g963) & (!g971)) + ((g747) & (!g744) & (!g748) & (g962) & (!g963) & (!g971)) + ((g747) & (!g744) & (!g748) & (g962) & (g963) & (!g971)) + ((g747) & (!g744) & (g748) & (!g962) & (!g963) & (!g971)) + ((g747) & (!g744) & (g748) & (g962) & (!g963) & (!g971)) + ((g747) & (g744) & (!g748) & (g962) & (!g963) & (!g971)) + ((g747) & (g744) & (!g748) & (g962) & (g963) & (!g971)) + ((g747) & (g744) & (g748) & (g962) & (!g963) & (!g971)));
	assign g1164 = (((!g202) & (!g1115) & (!g1117) & (!g1120) & (!g1139) & (g1143)) + ((!g202) & (!g1115) & (!g1117) & (g1120) & (!g1139) & (!g1143)) + ((!g202) & (!g1115) & (!g1117) & (g1120) & (!g1139) & (g1143)) + ((!g202) & (!g1115) & (!g1117) & (g1120) & (g1139) & (g1143)) + ((!g202) & (!g1115) & (g1117) & (!g1120) & (!g1139) & (g1143)) + ((!g202) & (!g1115) & (g1117) & (g1120) & (!g1139) & (g1143)) + ((!g202) & (g1115) & (!g1117) & (!g1120) & (!g1139) & (!g1143)) + ((!g202) & (g1115) & (!g1117) & (!g1120) & (!g1139) & (g1143)) + ((!g202) & (g1115) & (!g1117) & (!g1120) & (g1139) & (g1143)) + ((!g202) & (g1115) & (!g1117) & (g1120) & (!g1139) & (!g1143)) + ((!g202) & (g1115) & (!g1117) & (g1120) & (!g1139) & (g1143)) + ((!g202) & (g1115) & (!g1117) & (g1120) & (g1139) & (g1143)) + ((!g202) & (g1115) & (g1117) & (!g1120) & (!g1139) & (g1143)) + ((!g202) & (g1115) & (g1117) & (g1120) & (!g1139) & (!g1143)) + ((!g202) & (g1115) & (g1117) & (g1120) & (!g1139) & (g1143)) + ((!g202) & (g1115) & (g1117) & (g1120) & (g1139) & (g1143)) + ((g202) & (!g1115) & (!g1117) & (!g1120) & (g1139) & (g1143)) + ((g202) & (!g1115) & (!g1117) & (g1120) & (!g1139) & (g1143)) + ((g202) & (!g1115) & (!g1117) & (g1120) & (g1139) & (!g1143)) + ((g202) & (!g1115) & (!g1117) & (g1120) & (g1139) & (g1143)) + ((g202) & (!g1115) & (g1117) & (!g1120) & (g1139) & (g1143)) + ((g202) & (!g1115) & (g1117) & (g1120) & (g1139) & (g1143)) + ((g202) & (g1115) & (!g1117) & (!g1120) & (!g1139) & (g1143)) + ((g202) & (g1115) & (!g1117) & (!g1120) & (g1139) & (!g1143)) + ((g202) & (g1115) & (!g1117) & (!g1120) & (g1139) & (g1143)) + ((g202) & (g1115) & (!g1117) & (g1120) & (!g1139) & (g1143)) + ((g202) & (g1115) & (!g1117) & (g1120) & (g1139) & (!g1143)) + ((g202) & (g1115) & (!g1117) & (g1120) & (g1139) & (g1143)) + ((g202) & (g1115) & (g1117) & (!g1120) & (g1139) & (g1143)) + ((g202) & (g1115) & (g1117) & (g1120) & (!g1139) & (g1143)) + ((g202) & (g1115) & (g1117) & (g1120) & (g1139) & (!g1143)) + ((g202) & (g1115) & (g1117) & (g1120) & (g1139) & (g1143)));
	assign g1165 = (((!g869) & (!g764) & (!g762) & (!g765) & (!g870) & (!g863)) + ((!g869) & (!g764) & (!g762) & (!g765) & (!g870) & (g863)) + ((!g869) & (!g764) & (!g762) & (!g765) & (g870) & (!g863)) + ((!g869) & (!g764) & (!g762) & (!g765) & (g870) & (g863)) + ((!g869) & (!g764) & (!g762) & (g765) & (!g870) & (!g863)) + ((!g869) & (!g764) & (!g762) & (g765) & (!g870) & (g863)) + ((!g869) & (!g764) & (!g762) & (g765) & (g870) & (!g863)) + ((!g869) & (!g764) & (!g762) & (g765) & (g870) & (g863)) + ((!g869) & (!g764) & (g762) & (!g765) & (g870) & (!g863)) + ((!g869) & (!g764) & (g762) & (!g765) & (g870) & (g863)) + ((!g869) & (!g764) & (g762) & (g765) & (g870) & (!g863)) + ((!g869) & (!g764) & (g762) & (g765) & (g870) & (g863)) + ((!g869) & (g764) & (!g762) & (!g765) & (!g870) & (!g863)) + ((!g869) & (g764) & (!g762) & (!g765) & (g870) & (!g863)) + ((!g869) & (g764) & (!g762) & (g765) & (!g870) & (!g863)) + ((!g869) & (g764) & (!g762) & (g765) & (g870) & (!g863)) + ((!g869) & (g764) & (g762) & (!g765) & (g870) & (!g863)) + ((!g869) & (g764) & (g762) & (g765) & (g870) & (!g863)) + ((g869) & (!g764) & (!g762) & (!g765) & (!g870) & (!g863)) + ((g869) & (!g764) & (!g762) & (!g765) & (!g870) & (g863)) + ((g869) & (!g764) & (!g762) & (!g765) & (g870) & (!g863)) + ((g869) & (!g764) & (!g762) & (!g765) & (g870) & (g863)) + ((g869) & (!g764) & (g762) & (!g765) & (g870) & (!g863)) + ((g869) & (!g764) & (g762) & (!g765) & (g870) & (g863)) + ((g869) & (g764) & (!g762) & (!g765) & (!g870) & (!g863)) + ((g869) & (g764) & (!g762) & (!g765) & (g870) & (!g863)) + ((g869) & (g764) & (g762) & (!g765) & (g870) & (!g863)));
	assign g1166 = (((!g252) & (!sk[24]) & (!g720) & (!g1140) & (g1142)) + ((!g252) & (!sk[24]) & (!g720) & (g1140) & (g1142)) + ((!g252) & (!sk[24]) & (g720) & (!g1140) & (g1142)) + ((!g252) & (!sk[24]) & (g720) & (g1140) & (g1142)) + ((!g252) & (sk[24]) & (!g720) & (g1140) & (!g1142)) + ((!g252) & (sk[24]) & (g720) & (g1140) & (!g1142)) + ((g252) & (!sk[24]) & (!g720) & (!g1140) & (!g1142)) + ((g252) & (!sk[24]) & (!g720) & (!g1140) & (g1142)) + ((g252) & (!sk[24]) & (!g720) & (g1140) & (!g1142)) + ((g252) & (!sk[24]) & (!g720) & (g1140) & (g1142)) + ((g252) & (!sk[24]) & (g720) & (!g1140) & (!g1142)) + ((g252) & (!sk[24]) & (g720) & (!g1140) & (g1142)) + ((g252) & (!sk[24]) & (g720) & (g1140) & (!g1142)) + ((g252) & (!sk[24]) & (g720) & (g1140) & (g1142)) + ((g252) & (sk[24]) & (!g720) & (g1140) & (g1142)) + ((g252) & (sk[24]) & (g720) & (!g1140) & (g1142)) + ((g252) & (sk[24]) & (g720) & (g1140) & (!g1142)) + ((g252) & (sk[24]) & (g720) & (g1140) & (g1142)));
	assign g1167 = (((!g549) & (!g569) & (!g680) & (!g729) & (!g845) & (g848)) + ((!g549) & (!g569) & (!g680) & (!g729) & (g845) & (g848)) + ((!g549) & (!g569) & (g680) & (!g729) & (!g845) & (g848)) + ((!g549) & (!g569) & (g680) & (!g729) & (g845) & (!g848)) + ((!g549) & (!g569) & (g680) & (!g729) & (g845) & (g848)) + ((!g549) & (!g569) & (g680) & (g729) & (g845) & (!g848)) + ((!g549) & (!g569) & (g680) & (g729) & (g845) & (g848)) + ((!g549) & (g569) & (!g680) & (!g729) & (!g845) & (g848)) + ((!g549) & (g569) & (!g680) & (!g729) & (g845) & (!g848)) + ((!g549) & (g569) & (!g680) & (!g729) & (g845) & (g848)) + ((!g549) & (g569) & (!g680) & (g729) & (g845) & (!g848)) + ((!g549) & (g569) & (!g680) & (g729) & (g845) & (g848)) + ((!g549) & (g569) & (g680) & (!g729) & (!g845) & (g848)) + ((!g549) & (g569) & (g680) & (!g729) & (g845) & (g848)) + ((g549) & (!g569) & (!g680) & (!g729) & (!g845) & (g848)) + ((g549) & (!g569) & (!g680) & (!g729) & (g845) & (!g848)) + ((g549) & (!g569) & (!g680) & (!g729) & (g845) & (g848)) + ((g549) & (!g569) & (!g680) & (g729) & (g845) & (!g848)) + ((g549) & (!g569) & (!g680) & (g729) & (g845) & (g848)) + ((g549) & (!g569) & (g680) & (!g729) & (!g845) & (g848)) + ((g549) & (!g569) & (g680) & (!g729) & (g845) & (g848)) + ((g549) & (g569) & (!g680) & (!g729) & (!g845) & (g848)) + ((g549) & (g569) & (!g680) & (!g729) & (g845) & (g848)) + ((g549) & (g569) & (g680) & (!g729) & (!g845) & (g848)) + ((g549) & (g569) & (g680) & (!g729) & (g845) & (!g848)) + ((g549) & (g569) & (g680) & (!g729) & (g845) & (g848)) + ((g549) & (g569) & (g680) & (g729) & (g845) & (!g848)) + ((g549) & (g569) & (g680) & (g729) & (g845) & (g848)));
	assign g1168 = (((!g681) & (!g718) & (!g730) & (!g847) & (!g843) & (!g1167)) + ((!g681) & (!g718) & (!g730) & (g847) & (!g843) & (!g1167)) + ((!g681) & (!g718) & (g730) & (!g847) & (!g843) & (!g1167)) + ((!g681) & (!g718) & (g730) & (!g847) & (g843) & (!g1167)) + ((!g681) & (!g718) & (g730) & (g847) & (!g843) & (!g1167)) + ((!g681) & (!g718) & (g730) & (g847) & (g843) & (!g1167)) + ((!g681) & (g718) & (!g730) & (!g847) & (!g843) & (!g1167)) + ((!g681) & (g718) & (!g730) & (!g847) & (g843) & (!g1167)) + ((!g681) & (g718) & (g730) & (!g847) & (!g843) & (!g1167)) + ((g681) & (!g718) & (!g730) & (!g847) & (!g843) & (!g1167)) + ((g681) & (!g718) & (!g730) & (!g847) & (g843) & (!g1167)) + ((g681) & (!g718) & (!g730) & (g847) & (!g843) & (!g1167)) + ((g681) & (!g718) & (!g730) & (g847) & (g843) & (!g1167)) + ((g681) & (!g718) & (g730) & (!g847) & (!g843) & (!g1167)) + ((g681) & (!g718) & (g730) & (g847) & (!g843) & (!g1167)) + ((g681) & (g718) & (!g730) & (!g847) & (!g843) & (!g1167)) + ((g681) & (g718) & (g730) & (!g847) & (!g843) & (!g1167)) + ((g681) & (g718) & (g730) & (!g847) & (g843) & (!g1167)));
	assign g1169 = (((!g252) & (!g683) & (!g719) & (!sk[27]) & (g1168)) + ((!g252) & (!g683) & (!g719) & (sk[27]) & (!g1168)) + ((!g252) & (!g683) & (g719) & (!sk[27]) & (g1168)) + ((!g252) & (!g683) & (g719) & (sk[27]) & (!g1168)) + ((!g252) & (g683) & (!g719) & (!sk[27]) & (g1168)) + ((!g252) & (g683) & (!g719) & (sk[27]) & (g1168)) + ((!g252) & (g683) & (g719) & (!sk[27]) & (g1168)) + ((!g252) & (g683) & (g719) & (sk[27]) & (g1168)) + ((g252) & (!g683) & (!g719) & (!sk[27]) & (!g1168)) + ((g252) & (!g683) & (!g719) & (!sk[27]) & (g1168)) + ((g252) & (!g683) & (!g719) & (sk[27]) & (!g1168)) + ((g252) & (!g683) & (g719) & (!sk[27]) & (!g1168)) + ((g252) & (!g683) & (g719) & (!sk[27]) & (g1168)) + ((g252) & (!g683) & (g719) & (sk[27]) & (g1168)) + ((g252) & (g683) & (!g719) & (!sk[27]) & (!g1168)) + ((g252) & (g683) & (!g719) & (!sk[27]) & (g1168)) + ((g252) & (g683) & (!g719) & (sk[27]) & (g1168)) + ((g252) & (g683) & (g719) & (!sk[27]) & (!g1168)) + ((g252) & (g683) & (g719) & (!sk[27]) & (g1168)) + ((g252) & (g683) & (g719) & (sk[27]) & (!g1168)));
	assign g1170 = (((!g202) & (!g759) & (!g899) & (!g1165) & (!g1166) & (!g1169)) + ((!g202) & (!g759) & (!g899) & (!g1165) & (g1166) & (g1169)) + ((!g202) & (!g759) & (!g899) & (g1165) & (!g1166) & (g1169)) + ((!g202) & (!g759) & (!g899) & (g1165) & (g1166) & (!g1169)) + ((!g202) & (!g759) & (g899) & (!g1165) & (!g1166) & (!g1169)) + ((!g202) & (!g759) & (g899) & (!g1165) & (g1166) & (g1169)) + ((!g202) & (!g759) & (g899) & (g1165) & (!g1166) & (g1169)) + ((!g202) & (!g759) & (g899) & (g1165) & (g1166) & (!g1169)) + ((!g202) & (g759) & (!g899) & (!g1165) & (!g1166) & (!g1169)) + ((!g202) & (g759) & (!g899) & (!g1165) & (g1166) & (g1169)) + ((!g202) & (g759) & (!g899) & (g1165) & (!g1166) & (!g1169)) + ((!g202) & (g759) & (!g899) & (g1165) & (g1166) & (g1169)) + ((!g202) & (g759) & (g899) & (!g1165) & (!g1166) & (!g1169)) + ((!g202) & (g759) & (g899) & (!g1165) & (g1166) & (g1169)) + ((!g202) & (g759) & (g899) & (g1165) & (!g1166) & (g1169)) + ((!g202) & (g759) & (g899) & (g1165) & (g1166) & (!g1169)) + ((g202) & (!g759) & (!g899) & (!g1165) & (!g1166) & (g1169)) + ((g202) & (!g759) & (!g899) & (!g1165) & (g1166) & (!g1169)) + ((g202) & (!g759) & (!g899) & (g1165) & (!g1166) & (!g1169)) + ((g202) & (!g759) & (!g899) & (g1165) & (g1166) & (g1169)) + ((g202) & (!g759) & (g899) & (!g1165) & (!g1166) & (g1169)) + ((g202) & (!g759) & (g899) & (!g1165) & (g1166) & (!g1169)) + ((g202) & (!g759) & (g899) & (g1165) & (!g1166) & (!g1169)) + ((g202) & (!g759) & (g899) & (g1165) & (g1166) & (g1169)) + ((g202) & (g759) & (!g899) & (!g1165) & (!g1166) & (g1169)) + ((g202) & (g759) & (!g899) & (!g1165) & (g1166) & (!g1169)) + ((g202) & (g759) & (!g899) & (g1165) & (!g1166) & (g1169)) + ((g202) & (g759) & (!g899) & (g1165) & (g1166) & (!g1169)) + ((g202) & (g759) & (g899) & (!g1165) & (!g1166) & (g1169)) + ((g202) & (g759) & (g899) & (!g1165) & (g1166) & (!g1169)) + ((g202) & (g759) & (g899) & (g1165) & (!g1166) & (!g1169)) + ((g202) & (g759) & (g899) & (g1165) & (g1166) & (g1169)));
	assign g1171 = (((!g200) & (!g742) & (!g972) & (!g1163) & (!g1164) & (!g1170)) + ((!g200) & (!g742) & (!g972) & (!g1163) & (g1164) & (g1170)) + ((!g200) & (!g742) & (!g972) & (g1163) & (!g1164) & (g1170)) + ((!g200) & (!g742) & (!g972) & (g1163) & (g1164) & (!g1170)) + ((!g200) & (!g742) & (g972) & (!g1163) & (!g1164) & (!g1170)) + ((!g200) & (!g742) & (g972) & (!g1163) & (g1164) & (g1170)) + ((!g200) & (!g742) & (g972) & (g1163) & (!g1164) & (g1170)) + ((!g200) & (!g742) & (g972) & (g1163) & (g1164) & (!g1170)) + ((!g200) & (g742) & (!g972) & (!g1163) & (!g1164) & (!g1170)) + ((!g200) & (g742) & (!g972) & (!g1163) & (g1164) & (g1170)) + ((!g200) & (g742) & (!g972) & (g1163) & (!g1164) & (!g1170)) + ((!g200) & (g742) & (!g972) & (g1163) & (g1164) & (g1170)) + ((!g200) & (g742) & (g972) & (!g1163) & (!g1164) & (!g1170)) + ((!g200) & (g742) & (g972) & (!g1163) & (g1164) & (g1170)) + ((!g200) & (g742) & (g972) & (g1163) & (!g1164) & (g1170)) + ((!g200) & (g742) & (g972) & (g1163) & (g1164) & (!g1170)) + ((g200) & (!g742) & (!g972) & (!g1163) & (!g1164) & (g1170)) + ((g200) & (!g742) & (!g972) & (!g1163) & (g1164) & (!g1170)) + ((g200) & (!g742) & (!g972) & (g1163) & (!g1164) & (!g1170)) + ((g200) & (!g742) & (!g972) & (g1163) & (g1164) & (g1170)) + ((g200) & (!g742) & (g972) & (!g1163) & (!g1164) & (g1170)) + ((g200) & (!g742) & (g972) & (!g1163) & (g1164) & (!g1170)) + ((g200) & (!g742) & (g972) & (g1163) & (!g1164) & (!g1170)) + ((g200) & (!g742) & (g972) & (g1163) & (g1164) & (g1170)) + ((g200) & (g742) & (!g972) & (!g1163) & (!g1164) & (g1170)) + ((g200) & (g742) & (!g972) & (!g1163) & (g1164) & (!g1170)) + ((g200) & (g742) & (!g972) & (g1163) & (!g1164) & (g1170)) + ((g200) & (g742) & (!g972) & (g1163) & (g1164) & (!g1170)) + ((g200) & (g742) & (g972) & (!g1163) & (!g1164) & (g1170)) + ((g200) & (g742) & (g972) & (!g1163) & (g1164) & (!g1170)) + ((g200) & (g742) & (g972) & (g1163) & (!g1164) & (!g1170)) + ((g200) & (g742) & (g972) & (g1163) & (g1164) & (g1170)));
	assign g1172 = (((!g733) & (!g686) & (!g734) & (!g994) & (!g1040) & (!g1079)) + ((!g733) & (!g686) & (!g734) & (!g994) & (!g1040) & (g1079)) + ((!g733) & (!g686) & (!g734) & (!g994) & (g1040) & (!g1079)) + ((!g733) & (!g686) & (!g734) & (!g994) & (g1040) & (g1079)) + ((!g733) & (!g686) & (!g734) & (g994) & (!g1040) & (!g1079)) + ((!g733) & (!g686) & (!g734) & (g994) & (!g1040) & (g1079)) + ((!g733) & (!g686) & (!g734) & (g994) & (g1040) & (!g1079)) + ((!g733) & (!g686) & (!g734) & (g994) & (g1040) & (g1079)) + ((!g733) & (!g686) & (g734) & (!g994) & (g1040) & (!g1079)) + ((!g733) & (!g686) & (g734) & (!g994) & (g1040) & (g1079)) + ((!g733) & (!g686) & (g734) & (g994) & (g1040) & (!g1079)) + ((!g733) & (!g686) & (g734) & (g994) & (g1040) & (g1079)) + ((!g733) & (g686) & (!g734) & (!g994) & (!g1040) & (!g1079)) + ((!g733) & (g686) & (!g734) & (!g994) & (!g1040) & (g1079)) + ((!g733) & (g686) & (!g734) & (!g994) & (g1040) & (!g1079)) + ((!g733) & (g686) & (!g734) & (!g994) & (g1040) & (g1079)) + ((!g733) & (g686) & (g734) & (!g994) & (g1040) & (!g1079)) + ((!g733) & (g686) & (g734) & (!g994) & (g1040) & (g1079)) + ((g733) & (!g686) & (!g734) & (!g994) & (!g1040) & (g1079)) + ((g733) & (!g686) & (!g734) & (!g994) & (g1040) & (g1079)) + ((g733) & (!g686) & (!g734) & (g994) & (!g1040) & (g1079)) + ((g733) & (!g686) & (!g734) & (g994) & (g1040) & (g1079)) + ((g733) & (!g686) & (g734) & (!g994) & (g1040) & (g1079)) + ((g733) & (!g686) & (g734) & (g994) & (g1040) & (g1079)) + ((g733) & (g686) & (!g734) & (!g994) & (!g1040) & (g1079)) + ((g733) & (g686) & (!g734) & (!g994) & (g1040) & (g1079)) + ((g733) & (g686) & (g734) & (!g994) & (g1040) & (g1079)));
	assign g1173 = (((!g2) & (!g732) & (!g1040) & (!g1079) & (!g1080) & (!g1172)) + ((!g2) & (!g732) & (!g1040) & (!g1079) & (g1080) & (!g1172)) + ((!g2) & (!g732) & (!g1040) & (g1079) & (!g1080) & (!g1172)) + ((!g2) & (!g732) & (!g1040) & (g1079) & (g1080) & (!g1172)) + ((!g2) & (!g732) & (g1040) & (!g1079) & (!g1080) & (!g1172)) + ((!g2) & (!g732) & (g1040) & (!g1079) & (g1080) & (!g1172)) + ((!g2) & (!g732) & (g1040) & (g1079) & (!g1080) & (!g1172)) + ((!g2) & (!g732) & (g1040) & (g1079) & (g1080) & (!g1172)) + ((!g2) & (g732) & (!g1040) & (!g1079) & (!g1080) & (!g1172)) + ((!g2) & (g732) & (!g1040) & (!g1079) & (g1080) & (!g1172)) + ((!g2) & (g732) & (!g1040) & (!g1079) & (g1080) & (g1172)) + ((!g2) & (g732) & (!g1040) & (g1079) & (!g1080) & (!g1172)) + ((!g2) & (g732) & (!g1040) & (g1079) & (!g1080) & (g1172)) + ((!g2) & (g732) & (!g1040) & (g1079) & (g1080) & (!g1172)) + ((!g2) & (g732) & (g1040) & (!g1079) & (!g1080) & (!g1172)) + ((!g2) & (g732) & (g1040) & (!g1079) & (!g1080) & (g1172)) + ((!g2) & (g732) & (g1040) & (!g1079) & (g1080) & (!g1172)) + ((!g2) & (g732) & (g1040) & (g1079) & (!g1080) & (!g1172)) + ((!g2) & (g732) & (g1040) & (g1079) & (g1080) & (!g1172)) + ((!g2) & (g732) & (g1040) & (g1079) & (g1080) & (g1172)) + ((g2) & (!g732) & (!g1040) & (!g1079) & (!g1080) & (g1172)) + ((g2) & (!g732) & (!g1040) & (!g1079) & (g1080) & (g1172)) + ((g2) & (!g732) & (!g1040) & (g1079) & (!g1080) & (g1172)) + ((g2) & (!g732) & (!g1040) & (g1079) & (g1080) & (g1172)) + ((g2) & (!g732) & (g1040) & (!g1079) & (!g1080) & (g1172)) + ((g2) & (!g732) & (g1040) & (!g1079) & (g1080) & (g1172)) + ((g2) & (!g732) & (g1040) & (g1079) & (!g1080) & (g1172)) + ((g2) & (!g732) & (g1040) & (g1079) & (g1080) & (g1172)) + ((g2) & (g732) & (!g1040) & (!g1079) & (!g1080) & (g1172)) + ((g2) & (g732) & (!g1040) & (g1079) & (g1080) & (g1172)) + ((g2) & (g732) & (g1040) & (!g1079) & (g1080) & (g1172)) + ((g2) & (g732) & (g1040) & (g1079) & (!g1080) & (g1172)));
	assign g1174 = (((!g1137) & (!g1144) & (!g1147) & (!sk[32]) & (g1171) & (!g1173)) + ((!g1137) & (!g1144) & (!g1147) & (!sk[32]) & (g1171) & (g1173)) + ((!g1137) & (!g1144) & (!g1147) & (sk[32]) & (!g1171) & (g1173)) + ((!g1137) & (!g1144) & (!g1147) & (sk[32]) & (g1171) & (!g1173)) + ((!g1137) & (!g1144) & (g1147) & (!sk[32]) & (!g1171) & (!g1173)) + ((!g1137) & (!g1144) & (g1147) & (!sk[32]) & (!g1171) & (g1173)) + ((!g1137) & (!g1144) & (g1147) & (!sk[32]) & (g1171) & (!g1173)) + ((!g1137) & (!g1144) & (g1147) & (!sk[32]) & (g1171) & (g1173)) + ((!g1137) & (!g1144) & (g1147) & (sk[32]) & (!g1171) & (!g1173)) + ((!g1137) & (!g1144) & (g1147) & (sk[32]) & (g1171) & (g1173)) + ((!g1137) & (g1144) & (!g1147) & (!sk[32]) & (!g1171) & (!g1173)) + ((!g1137) & (g1144) & (!g1147) & (!sk[32]) & (!g1171) & (g1173)) + ((!g1137) & (g1144) & (!g1147) & (!sk[32]) & (g1171) & (!g1173)) + ((!g1137) & (g1144) & (!g1147) & (!sk[32]) & (g1171) & (g1173)) + ((!g1137) & (g1144) & (!g1147) & (sk[32]) & (!g1171) & (g1173)) + ((!g1137) & (g1144) & (!g1147) & (sk[32]) & (g1171) & (!g1173)) + ((!g1137) & (g1144) & (g1147) & (!sk[32]) & (!g1171) & (!g1173)) + ((!g1137) & (g1144) & (g1147) & (!sk[32]) & (!g1171) & (g1173)) + ((!g1137) & (g1144) & (g1147) & (!sk[32]) & (g1171) & (!g1173)) + ((!g1137) & (g1144) & (g1147) & (!sk[32]) & (g1171) & (g1173)) + ((!g1137) & (g1144) & (g1147) & (sk[32]) & (!g1171) & (g1173)) + ((!g1137) & (g1144) & (g1147) & (sk[32]) & (g1171) & (!g1173)) + ((g1137) & (!g1144) & (!g1147) & (!sk[32]) & (g1171) & (!g1173)) + ((g1137) & (!g1144) & (!g1147) & (!sk[32]) & (g1171) & (g1173)) + ((g1137) & (!g1144) & (!g1147) & (sk[32]) & (!g1171) & (!g1173)) + ((g1137) & (!g1144) & (!g1147) & (sk[32]) & (g1171) & (g1173)) + ((g1137) & (!g1144) & (g1147) & (!sk[32]) & (!g1171) & (!g1173)) + ((g1137) & (!g1144) & (g1147) & (!sk[32]) & (!g1171) & (g1173)) + ((g1137) & (!g1144) & (g1147) & (!sk[32]) & (g1171) & (!g1173)) + ((g1137) & (!g1144) & (g1147) & (!sk[32]) & (g1171) & (g1173)) + ((g1137) & (!g1144) & (g1147) & (sk[32]) & (!g1171) & (!g1173)) + ((g1137) & (!g1144) & (g1147) & (sk[32]) & (g1171) & (g1173)) + ((g1137) & (g1144) & (!g1147) & (!sk[32]) & (!g1171) & (!g1173)) + ((g1137) & (g1144) & (!g1147) & (!sk[32]) & (!g1171) & (g1173)) + ((g1137) & (g1144) & (!g1147) & (!sk[32]) & (g1171) & (!g1173)) + ((g1137) & (g1144) & (!g1147) & (!sk[32]) & (g1171) & (g1173)) + ((g1137) & (g1144) & (!g1147) & (sk[32]) & (!g1171) & (g1173)) + ((g1137) & (g1144) & (!g1147) & (sk[32]) & (g1171) & (!g1173)) + ((g1137) & (g1144) & (g1147) & (!sk[32]) & (!g1171) & (!g1173)) + ((g1137) & (g1144) & (g1147) & (!sk[32]) & (!g1171) & (g1173)) + ((g1137) & (g1144) & (g1147) & (!sk[32]) & (g1171) & (!g1173)) + ((g1137) & (g1144) & (g1147) & (!sk[32]) & (g1171) & (g1173)) + ((g1137) & (g1144) & (g1147) & (sk[32]) & (!g1171) & (!g1173)) + ((g1137) & (g1144) & (g1147) & (sk[32]) & (g1171) & (g1173)));
	assign g1175 = (((!g1161) & (!sk[33]) & (g1162) & (!g1174)) + ((!g1161) & (!sk[33]) & (g1162) & (g1174)) + ((!g1161) & (sk[33]) & (!g1162) & (!g1174)) + ((!g1161) & (sk[33]) & (g1162) & (g1174)) + ((g1161) & (!sk[33]) & (g1162) & (!g1174)) + ((g1161) & (!sk[33]) & (g1162) & (g1174)) + ((g1161) & (sk[33]) & (!g1162) & (g1174)) + ((g1161) & (sk[33]) & (g1162) & (!g1174)));
	assign g1176 = (((!g62) & (!sk[34]) & (!g66) & (!g193) & (g194)) + ((!g62) & (!sk[34]) & (!g66) & (g193) & (g194)) + ((!g62) & (!sk[34]) & (g66) & (!g193) & (g194)) + ((!g62) & (!sk[34]) & (g66) & (g193) & (g194)) + ((!g62) & (sk[34]) & (!g66) & (!g193) & (!g194)) + ((!g62) & (sk[34]) & (g66) & (!g193) & (!g194)) + ((g62) & (!sk[34]) & (!g66) & (!g193) & (!g194)) + ((g62) & (!sk[34]) & (!g66) & (!g193) & (g194)) + ((g62) & (!sk[34]) & (!g66) & (g193) & (!g194)) + ((g62) & (!sk[34]) & (!g66) & (g193) & (g194)) + ((g62) & (!sk[34]) & (g66) & (!g193) & (!g194)) + ((g62) & (!sk[34]) & (g66) & (!g193) & (g194)) + ((g62) & (!sk[34]) & (g66) & (g193) & (!g194)) + ((g62) & (!sk[34]) & (g66) & (g193) & (g194)) + ((g62) & (sk[34]) & (!g66) & (!g193) & (!g194)));
	assign g1177 = (((!sk[35]) & (g70) & (g155)) + ((sk[35]) & (g70) & (g155)));
	assign g1178 = (((!g9) & (!g46) & (!g40) & (!g32) & (!g84) & (!g1177)) + ((!g9) & (!g46) & (!g40) & (g32) & (!g84) & (!g1177)) + ((!g9) & (!g46) & (g40) & (!g32) & (!g84) & (!g1177)) + ((!g9) & (!g46) & (g40) & (g32) & (!g84) & (!g1177)) + ((!g9) & (g46) & (!g40) & (!g32) & (!g84) & (!g1177)) + ((!g9) & (g46) & (!g40) & (g32) & (!g84) & (!g1177)) + ((g9) & (!g46) & (!g40) & (!g32) & (!g84) & (!g1177)) + ((g9) & (!g46) & (g40) & (!g32) & (!g84) & (!g1177)) + ((g9) & (g46) & (!g40) & (!g32) & (!g84) & (!g1177)));
	assign g1179 = (((!g9) & (!g30) & (!sk[37]) & (!g104) & (g25)) + ((!g9) & (!g30) & (!sk[37]) & (g104) & (g25)) + ((!g9) & (g30) & (!sk[37]) & (!g104) & (g25)) + ((!g9) & (g30) & (!sk[37]) & (g104) & (g25)) + ((!g9) & (g30) & (sk[37]) & (g104) & (!g25)) + ((!g9) & (g30) & (sk[37]) & (g104) & (g25)) + ((g9) & (!g30) & (!sk[37]) & (!g104) & (!g25)) + ((g9) & (!g30) & (!sk[37]) & (!g104) & (g25)) + ((g9) & (!g30) & (!sk[37]) & (g104) & (!g25)) + ((g9) & (!g30) & (!sk[37]) & (g104) & (g25)) + ((g9) & (!g30) & (sk[37]) & (!g104) & (g25)) + ((g9) & (!g30) & (sk[37]) & (g104) & (g25)) + ((g9) & (g30) & (!sk[37]) & (!g104) & (!g25)) + ((g9) & (g30) & (!sk[37]) & (!g104) & (g25)) + ((g9) & (g30) & (!sk[37]) & (g104) & (!g25)) + ((g9) & (g30) & (!sk[37]) & (g104) & (g25)) + ((g9) & (g30) & (sk[37]) & (!g104) & (!g25)) + ((g9) & (g30) & (sk[37]) & (!g104) & (g25)) + ((g9) & (g30) & (sk[37]) & (g104) & (!g25)) + ((g9) & (g30) & (sk[37]) & (g104) & (g25)));
	assign g1180 = (((!g17) & (!g46) & (!g642) & (!sk[38]) & (g1179)) + ((!g17) & (!g46) & (!g642) & (sk[38]) & (!g1179)) + ((!g17) & (!g46) & (g642) & (!sk[38]) & (g1179)) + ((!g17) & (g46) & (!g642) & (!sk[38]) & (g1179)) + ((!g17) & (g46) & (!g642) & (sk[38]) & (!g1179)) + ((!g17) & (g46) & (g642) & (!sk[38]) & (g1179)) + ((g17) & (!g46) & (!g642) & (!sk[38]) & (!g1179)) + ((g17) & (!g46) & (!g642) & (!sk[38]) & (g1179)) + ((g17) & (!g46) & (!g642) & (sk[38]) & (!g1179)) + ((g17) & (!g46) & (g642) & (!sk[38]) & (!g1179)) + ((g17) & (!g46) & (g642) & (!sk[38]) & (g1179)) + ((g17) & (g46) & (!g642) & (!sk[38]) & (!g1179)) + ((g17) & (g46) & (!g642) & (!sk[38]) & (g1179)) + ((g17) & (g46) & (g642) & (!sk[38]) & (!g1179)) + ((g17) & (g46) & (g642) & (!sk[38]) & (g1179)));
	assign g1181 = (((!sk[39]) & (!g593) & (!g157) & (!g1062) & (g1178) & (!g1180)) + ((!sk[39]) & (!g593) & (!g157) & (!g1062) & (g1178) & (g1180)) + ((!sk[39]) & (!g593) & (!g157) & (g1062) & (!g1178) & (!g1180)) + ((!sk[39]) & (!g593) & (!g157) & (g1062) & (!g1178) & (g1180)) + ((!sk[39]) & (!g593) & (!g157) & (g1062) & (g1178) & (!g1180)) + ((!sk[39]) & (!g593) & (!g157) & (g1062) & (g1178) & (g1180)) + ((!sk[39]) & (!g593) & (g157) & (!g1062) & (!g1178) & (!g1180)) + ((!sk[39]) & (!g593) & (g157) & (!g1062) & (!g1178) & (g1180)) + ((!sk[39]) & (!g593) & (g157) & (!g1062) & (g1178) & (!g1180)) + ((!sk[39]) & (!g593) & (g157) & (!g1062) & (g1178) & (g1180)) + ((!sk[39]) & (!g593) & (g157) & (g1062) & (!g1178) & (!g1180)) + ((!sk[39]) & (!g593) & (g157) & (g1062) & (!g1178) & (g1180)) + ((!sk[39]) & (!g593) & (g157) & (g1062) & (g1178) & (!g1180)) + ((!sk[39]) & (!g593) & (g157) & (g1062) & (g1178) & (g1180)) + ((!sk[39]) & (g593) & (!g157) & (!g1062) & (g1178) & (!g1180)) + ((!sk[39]) & (g593) & (!g157) & (!g1062) & (g1178) & (g1180)) + ((!sk[39]) & (g593) & (!g157) & (g1062) & (!g1178) & (!g1180)) + ((!sk[39]) & (g593) & (!g157) & (g1062) & (!g1178) & (g1180)) + ((!sk[39]) & (g593) & (!g157) & (g1062) & (g1178) & (!g1180)) + ((!sk[39]) & (g593) & (!g157) & (g1062) & (g1178) & (g1180)) + ((!sk[39]) & (g593) & (g157) & (!g1062) & (!g1178) & (!g1180)) + ((!sk[39]) & (g593) & (g157) & (!g1062) & (!g1178) & (g1180)) + ((!sk[39]) & (g593) & (g157) & (!g1062) & (g1178) & (!g1180)) + ((!sk[39]) & (g593) & (g157) & (!g1062) & (g1178) & (g1180)) + ((!sk[39]) & (g593) & (g157) & (g1062) & (!g1178) & (!g1180)) + ((!sk[39]) & (g593) & (g157) & (g1062) & (!g1178) & (g1180)) + ((!sk[39]) & (g593) & (g157) & (g1062) & (g1178) & (!g1180)) + ((!sk[39]) & (g593) & (g157) & (g1062) & (g1178) & (g1180)) + ((sk[39]) & (!g593) & (g157) & (g1062) & (g1178) & (g1180)));
	assign g1182 = (((!g1176) & (!sk[40]) & (!g629) & (!g669) & (g1181)) + ((!g1176) & (!sk[40]) & (!g629) & (g669) & (g1181)) + ((!g1176) & (!sk[40]) & (g629) & (!g669) & (g1181)) + ((!g1176) & (!sk[40]) & (g629) & (g669) & (g1181)) + ((g1176) & (!sk[40]) & (!g629) & (!g669) & (!g1181)) + ((g1176) & (!sk[40]) & (!g629) & (!g669) & (g1181)) + ((g1176) & (!sk[40]) & (!g629) & (g669) & (!g1181)) + ((g1176) & (!sk[40]) & (!g629) & (g669) & (g1181)) + ((g1176) & (!sk[40]) & (g629) & (!g669) & (!g1181)) + ((g1176) & (!sk[40]) & (g629) & (!g669) & (g1181)) + ((g1176) & (!sk[40]) & (g629) & (g669) & (!g1181)) + ((g1176) & (!sk[40]) & (g629) & (g669) & (g1181)) + ((g1176) & (sk[40]) & (g629) & (g669) & (g1181)));
	assign g1183 = (((!g1160) & (!g1175) & (sk[41]) & (!g1182)) + ((!g1160) & (g1175) & (!sk[41]) & (!g1182)) + ((!g1160) & (g1175) & (!sk[41]) & (g1182)) + ((!g1160) & (g1175) & (sk[41]) & (g1182)) + ((g1160) & (!g1175) & (sk[41]) & (g1182)) + ((g1160) & (g1175) & (!sk[41]) & (!g1182)) + ((g1160) & (g1175) & (!sk[41]) & (g1182)) + ((g1160) & (g1175) & (sk[41]) & (!g1182)));
	assign sinx4x = (((!g1068) & (!sk[42]) & (!g1135) & (!g1157) & (g1158) & (!g1183)) + ((!g1068) & (!sk[42]) & (!g1135) & (!g1157) & (g1158) & (g1183)) + ((!g1068) & (!sk[42]) & (!g1135) & (g1157) & (!g1158) & (!g1183)) + ((!g1068) & (!sk[42]) & (!g1135) & (g1157) & (!g1158) & (g1183)) + ((!g1068) & (!sk[42]) & (!g1135) & (g1157) & (g1158) & (!g1183)) + ((!g1068) & (!sk[42]) & (!g1135) & (g1157) & (g1158) & (g1183)) + ((!g1068) & (!sk[42]) & (g1135) & (!g1157) & (!g1158) & (!g1183)) + ((!g1068) & (!sk[42]) & (g1135) & (!g1157) & (!g1158) & (g1183)) + ((!g1068) & (!sk[42]) & (g1135) & (!g1157) & (g1158) & (!g1183)) + ((!g1068) & (!sk[42]) & (g1135) & (!g1157) & (g1158) & (g1183)) + ((!g1068) & (!sk[42]) & (g1135) & (g1157) & (!g1158) & (!g1183)) + ((!g1068) & (!sk[42]) & (g1135) & (g1157) & (!g1158) & (g1183)) + ((!g1068) & (!sk[42]) & (g1135) & (g1157) & (g1158) & (!g1183)) + ((!g1068) & (!sk[42]) & (g1135) & (g1157) & (g1158) & (g1183)) + ((!g1068) & (sk[42]) & (!g1135) & (!g1157) & (!g1158) & (g1183)) + ((!g1068) & (sk[42]) & (!g1135) & (!g1157) & (g1158) & (g1183)) + ((!g1068) & (sk[42]) & (!g1135) & (g1157) & (!g1158) & (g1183)) + ((!g1068) & (sk[42]) & (!g1135) & (g1157) & (g1158) & (g1183)) + ((!g1068) & (sk[42]) & (g1135) & (!g1157) & (!g1158) & (g1183)) + ((!g1068) & (sk[42]) & (g1135) & (!g1157) & (g1158) & (g1183)) + ((!g1068) & (sk[42]) & (g1135) & (g1157) & (!g1158) & (!g1183)) + ((!g1068) & (sk[42]) & (g1135) & (g1157) & (g1158) & (!g1183)) + ((g1068) & (!sk[42]) & (!g1135) & (!g1157) & (g1158) & (!g1183)) + ((g1068) & (!sk[42]) & (!g1135) & (!g1157) & (g1158) & (g1183)) + ((g1068) & (!sk[42]) & (!g1135) & (g1157) & (!g1158) & (!g1183)) + ((g1068) & (!sk[42]) & (!g1135) & (g1157) & (!g1158) & (g1183)) + ((g1068) & (!sk[42]) & (!g1135) & (g1157) & (g1158) & (!g1183)) + ((g1068) & (!sk[42]) & (!g1135) & (g1157) & (g1158) & (g1183)) + ((g1068) & (!sk[42]) & (g1135) & (!g1157) & (!g1158) & (!g1183)) + ((g1068) & (!sk[42]) & (g1135) & (!g1157) & (!g1158) & (g1183)) + ((g1068) & (!sk[42]) & (g1135) & (!g1157) & (g1158) & (!g1183)) + ((g1068) & (!sk[42]) & (g1135) & (!g1157) & (g1158) & (g1183)) + ((g1068) & (!sk[42]) & (g1135) & (g1157) & (!g1158) & (!g1183)) + ((g1068) & (!sk[42]) & (g1135) & (g1157) & (!g1158) & (g1183)) + ((g1068) & (!sk[42]) & (g1135) & (g1157) & (g1158) & (!g1183)) + ((g1068) & (!sk[42]) & (g1135) & (g1157) & (g1158) & (g1183)) + ((g1068) & (sk[42]) & (!g1135) & (!g1157) & (!g1158) & (!g1183)) + ((g1068) & (sk[42]) & (!g1135) & (!g1157) & (g1158) & (g1183)) + ((g1068) & (sk[42]) & (!g1135) & (g1157) & (!g1158) & (!g1183)) + ((g1068) & (sk[42]) & (!g1135) & (g1157) & (g1158) & (!g1183)) + ((g1068) & (sk[42]) & (g1135) & (!g1157) & (!g1158) & (!g1183)) + ((g1068) & (sk[42]) & (g1135) & (!g1157) & (g1158) & (!g1183)) + ((g1068) & (sk[42]) & (g1135) & (g1157) & (!g1158) & (g1183)) + ((g1068) & (sk[42]) & (g1135) & (g1157) & (g1158) & (!g1183)));
	assign g1185 = (((!g1135) & (!g1157) & (g1158) & (!g1160) & (!g1175) & (g1182)) + ((!g1135) & (!g1157) & (g1158) & (!g1160) & (g1175) & (!g1182)) + ((!g1135) & (!g1157) & (g1158) & (g1160) & (!g1175) & (!g1182)) + ((!g1135) & (!g1157) & (g1158) & (g1160) & (g1175) & (g1182)) + ((g1135) & (g1157) & (g1158) & (!g1160) & (!g1175) & (!g1182)) + ((g1135) & (g1157) & (g1158) & (!g1160) & (g1175) & (g1182)) + ((g1135) & (g1157) & (g1158) & (g1160) & (!g1175) & (g1182)) + ((g1135) & (g1157) & (g1158) & (g1160) & (g1175) & (!g1182)));
	assign g1186 = (((!sk[44]) & (!g1135) & (!g1157) & (!g1160) & (g1175) & (!g1182)) + ((!sk[44]) & (!g1135) & (!g1157) & (!g1160) & (g1175) & (g1182)) + ((!sk[44]) & (!g1135) & (!g1157) & (g1160) & (!g1175) & (!g1182)) + ((!sk[44]) & (!g1135) & (!g1157) & (g1160) & (!g1175) & (g1182)) + ((!sk[44]) & (!g1135) & (!g1157) & (g1160) & (g1175) & (!g1182)) + ((!sk[44]) & (!g1135) & (!g1157) & (g1160) & (g1175) & (g1182)) + ((!sk[44]) & (!g1135) & (g1157) & (!g1160) & (!g1175) & (!g1182)) + ((!sk[44]) & (!g1135) & (g1157) & (!g1160) & (!g1175) & (g1182)) + ((!sk[44]) & (!g1135) & (g1157) & (!g1160) & (g1175) & (!g1182)) + ((!sk[44]) & (!g1135) & (g1157) & (!g1160) & (g1175) & (g1182)) + ((!sk[44]) & (!g1135) & (g1157) & (g1160) & (!g1175) & (!g1182)) + ((!sk[44]) & (!g1135) & (g1157) & (g1160) & (!g1175) & (g1182)) + ((!sk[44]) & (!g1135) & (g1157) & (g1160) & (g1175) & (!g1182)) + ((!sk[44]) & (!g1135) & (g1157) & (g1160) & (g1175) & (g1182)) + ((!sk[44]) & (g1135) & (!g1157) & (!g1160) & (g1175) & (!g1182)) + ((!sk[44]) & (g1135) & (!g1157) & (!g1160) & (g1175) & (g1182)) + ((!sk[44]) & (g1135) & (!g1157) & (g1160) & (!g1175) & (!g1182)) + ((!sk[44]) & (g1135) & (!g1157) & (g1160) & (!g1175) & (g1182)) + ((!sk[44]) & (g1135) & (!g1157) & (g1160) & (g1175) & (!g1182)) + ((!sk[44]) & (g1135) & (!g1157) & (g1160) & (g1175) & (g1182)) + ((!sk[44]) & (g1135) & (g1157) & (!g1160) & (!g1175) & (!g1182)) + ((!sk[44]) & (g1135) & (g1157) & (!g1160) & (!g1175) & (g1182)) + ((!sk[44]) & (g1135) & (g1157) & (!g1160) & (g1175) & (!g1182)) + ((!sk[44]) & (g1135) & (g1157) & (!g1160) & (g1175) & (g1182)) + ((!sk[44]) & (g1135) & (g1157) & (g1160) & (!g1175) & (!g1182)) + ((!sk[44]) & (g1135) & (g1157) & (g1160) & (!g1175) & (g1182)) + ((!sk[44]) & (g1135) & (g1157) & (g1160) & (g1175) & (!g1182)) + ((!sk[44]) & (g1135) & (g1157) & (g1160) & (g1175) & (g1182)) + ((sk[44]) & (g1135) & (g1157) & (!g1160) & (!g1175) & (!g1182)) + ((sk[44]) & (g1135) & (g1157) & (!g1160) & (g1175) & (g1182)) + ((sk[44]) & (g1135) & (g1157) & (g1160) & (!g1175) & (g1182)) + ((sk[44]) & (g1135) & (g1157) & (g1160) & (g1175) & (!g1182)));
	assign g1187 = (((!g1137) & (!g1144) & (!g1147) & (!sk[45]) & (g1171) & (!g1173)) + ((!g1137) & (!g1144) & (!g1147) & (!sk[45]) & (g1171) & (g1173)) + ((!g1137) & (!g1144) & (!g1147) & (sk[45]) & (g1171) & (g1173)) + ((!g1137) & (!g1144) & (g1147) & (!sk[45]) & (!g1171) & (!g1173)) + ((!g1137) & (!g1144) & (g1147) & (!sk[45]) & (!g1171) & (g1173)) + ((!g1137) & (!g1144) & (g1147) & (!sk[45]) & (g1171) & (!g1173)) + ((!g1137) & (!g1144) & (g1147) & (!sk[45]) & (g1171) & (g1173)) + ((!g1137) & (!g1144) & (g1147) & (sk[45]) & (!g1171) & (g1173)) + ((!g1137) & (!g1144) & (g1147) & (sk[45]) & (g1171) & (!g1173)) + ((!g1137) & (!g1144) & (g1147) & (sk[45]) & (g1171) & (g1173)) + ((!g1137) & (g1144) & (!g1147) & (!sk[45]) & (!g1171) & (!g1173)) + ((!g1137) & (g1144) & (!g1147) & (!sk[45]) & (!g1171) & (g1173)) + ((!g1137) & (g1144) & (!g1147) & (!sk[45]) & (g1171) & (!g1173)) + ((!g1137) & (g1144) & (!g1147) & (!sk[45]) & (g1171) & (g1173)) + ((!g1137) & (g1144) & (!g1147) & (sk[45]) & (g1171) & (g1173)) + ((!g1137) & (g1144) & (g1147) & (!sk[45]) & (!g1171) & (!g1173)) + ((!g1137) & (g1144) & (g1147) & (!sk[45]) & (!g1171) & (g1173)) + ((!g1137) & (g1144) & (g1147) & (!sk[45]) & (g1171) & (!g1173)) + ((!g1137) & (g1144) & (g1147) & (!sk[45]) & (g1171) & (g1173)) + ((!g1137) & (g1144) & (g1147) & (sk[45]) & (g1171) & (g1173)) + ((g1137) & (!g1144) & (!g1147) & (!sk[45]) & (g1171) & (!g1173)) + ((g1137) & (!g1144) & (!g1147) & (!sk[45]) & (g1171) & (g1173)) + ((g1137) & (!g1144) & (!g1147) & (sk[45]) & (!g1171) & (g1173)) + ((g1137) & (!g1144) & (!g1147) & (sk[45]) & (g1171) & (!g1173)) + ((g1137) & (!g1144) & (!g1147) & (sk[45]) & (g1171) & (g1173)) + ((g1137) & (!g1144) & (g1147) & (!sk[45]) & (!g1171) & (!g1173)) + ((g1137) & (!g1144) & (g1147) & (!sk[45]) & (!g1171) & (g1173)) + ((g1137) & (!g1144) & (g1147) & (!sk[45]) & (g1171) & (!g1173)) + ((g1137) & (!g1144) & (g1147) & (!sk[45]) & (g1171) & (g1173)) + ((g1137) & (!g1144) & (g1147) & (sk[45]) & (!g1171) & (g1173)) + ((g1137) & (!g1144) & (g1147) & (sk[45]) & (g1171) & (!g1173)) + ((g1137) & (!g1144) & (g1147) & (sk[45]) & (g1171) & (g1173)) + ((g1137) & (g1144) & (!g1147) & (!sk[45]) & (!g1171) & (!g1173)) + ((g1137) & (g1144) & (!g1147) & (!sk[45]) & (!g1171) & (g1173)) + ((g1137) & (g1144) & (!g1147) & (!sk[45]) & (g1171) & (!g1173)) + ((g1137) & (g1144) & (!g1147) & (!sk[45]) & (g1171) & (g1173)) + ((g1137) & (g1144) & (!g1147) & (sk[45]) & (g1171) & (g1173)) + ((g1137) & (g1144) & (g1147) & (!sk[45]) & (!g1171) & (!g1173)) + ((g1137) & (g1144) & (g1147) & (!sk[45]) & (!g1171) & (g1173)) + ((g1137) & (g1144) & (g1147) & (!sk[45]) & (g1171) & (!g1173)) + ((g1137) & (g1144) & (g1147) & (!sk[45]) & (g1171) & (g1173)) + ((g1137) & (g1144) & (g1147) & (sk[45]) & (!g1171) & (g1173)) + ((g1137) & (g1144) & (g1147) & (sk[45]) & (g1171) & (!g1173)) + ((g1137) & (g1144) & (g1147) & (sk[45]) & (g1171) & (g1173)));
	assign g1188 = (((!g1040) & (!sk[46]) & (g1079) & (!g1080)) + ((!g1040) & (!sk[46]) & (g1079) & (g1080)) + ((!g1040) & (sk[46]) & (g1079) & (g1080)) + ((g1040) & (!sk[46]) & (g1079) & (!g1080)) + ((g1040) & (!sk[46]) & (g1079) & (g1080)) + ((g1040) & (sk[46]) & (!g1079) & (!g1080)));
	assign g1189 = (((!g686) & (!sk[47]) & (!g734) & (!g1040) & (g1079)) + ((!g686) & (!sk[47]) & (!g734) & (g1040) & (g1079)) + ((!g686) & (!sk[47]) & (g734) & (!g1040) & (g1079)) + ((!g686) & (!sk[47]) & (g734) & (g1040) & (g1079)) + ((!g686) & (sk[47]) & (g734) & (!g1040) & (!g1079)) + ((!g686) & (sk[47]) & (g734) & (g1040) & (!g1079)) + ((g686) & (!sk[47]) & (!g734) & (!g1040) & (!g1079)) + ((g686) & (!sk[47]) & (!g734) & (!g1040) & (g1079)) + ((g686) & (!sk[47]) & (!g734) & (g1040) & (!g1079)) + ((g686) & (!sk[47]) & (!g734) & (g1040) & (g1079)) + ((g686) & (!sk[47]) & (g734) & (!g1040) & (!g1079)) + ((g686) & (!sk[47]) & (g734) & (!g1040) & (g1079)) + ((g686) & (!sk[47]) & (g734) & (g1040) & (!g1079)) + ((g686) & (!sk[47]) & (g734) & (g1040) & (g1079)) + ((g686) & (sk[47]) & (!g734) & (!g1040) & (!g1079)) + ((g686) & (sk[47]) & (!g734) & (!g1040) & (g1079)) + ((g686) & (sk[47]) & (g734) & (!g1040) & (!g1079)) + ((g686) & (sk[47]) & (g734) & (!g1040) & (g1079)) + ((g686) & (sk[47]) & (g734) & (g1040) & (!g1079)));
	assign g1190 = (((!g200) & (!g742) & (!g972) & (!g1163) & (!g1164) & (g1170)) + ((!g200) & (!g742) & (!g972) & (!g1163) & (g1164) & (!g1170)) + ((!g200) & (!g742) & (!g972) & (!g1163) & (g1164) & (g1170)) + ((!g200) & (!g742) & (!g972) & (g1163) & (g1164) & (g1170)) + ((!g200) & (!g742) & (g972) & (!g1163) & (!g1164) & (g1170)) + ((!g200) & (!g742) & (g972) & (!g1163) & (g1164) & (!g1170)) + ((!g200) & (!g742) & (g972) & (!g1163) & (g1164) & (g1170)) + ((!g200) & (!g742) & (g972) & (g1163) & (g1164) & (g1170)) + ((!g200) & (g742) & (!g972) & (!g1163) & (!g1164) & (g1170)) + ((!g200) & (g742) & (!g972) & (!g1163) & (g1164) & (!g1170)) + ((!g200) & (g742) & (!g972) & (!g1163) & (g1164) & (g1170)) + ((!g200) & (g742) & (!g972) & (g1163) & (!g1164) & (g1170)) + ((!g200) & (g742) & (!g972) & (g1163) & (g1164) & (!g1170)) + ((!g200) & (g742) & (!g972) & (g1163) & (g1164) & (g1170)) + ((!g200) & (g742) & (g972) & (!g1163) & (!g1164) & (g1170)) + ((!g200) & (g742) & (g972) & (!g1163) & (g1164) & (!g1170)) + ((!g200) & (g742) & (g972) & (!g1163) & (g1164) & (g1170)) + ((!g200) & (g742) & (g972) & (g1163) & (g1164) & (g1170)) + ((g200) & (!g742) & (!g972) & (!g1163) & (g1164) & (g1170)) + ((g200) & (!g742) & (!g972) & (g1163) & (!g1164) & (g1170)) + ((g200) & (!g742) & (!g972) & (g1163) & (g1164) & (!g1170)) + ((g200) & (!g742) & (!g972) & (g1163) & (g1164) & (g1170)) + ((g200) & (!g742) & (g972) & (!g1163) & (g1164) & (g1170)) + ((g200) & (!g742) & (g972) & (g1163) & (!g1164) & (g1170)) + ((g200) & (!g742) & (g972) & (g1163) & (g1164) & (!g1170)) + ((g200) & (!g742) & (g972) & (g1163) & (g1164) & (g1170)) + ((g200) & (g742) & (!g972) & (!g1163) & (g1164) & (g1170)) + ((g200) & (g742) & (!g972) & (g1163) & (g1164) & (g1170)) + ((g200) & (g742) & (g972) & (!g1163) & (g1164) & (g1170)) + ((g200) & (g742) & (g972) & (g1163) & (!g1164) & (g1170)) + ((g200) & (g742) & (g972) & (g1163) & (g1164) & (!g1170)) + ((g200) & (g742) & (g972) & (g1163) & (g1164) & (g1170)));
	assign g1191 = (((!g747) & (!g744) & (!g748) & (!g962) & (!g971) & (!g994)) + ((!g747) & (!g744) & (!g748) & (!g962) & (!g971) & (g994)) + ((!g747) & (!g744) & (!g748) & (!g962) & (g971) & (!g994)) + ((!g747) & (!g744) & (!g748) & (!g962) & (g971) & (g994)) + ((!g747) & (!g744) & (!g748) & (g962) & (!g971) & (!g994)) + ((!g747) & (!g744) & (!g748) & (g962) & (!g971) & (g994)) + ((!g747) & (!g744) & (!g748) & (g962) & (g971) & (!g994)) + ((!g747) & (!g744) & (!g748) & (g962) & (g971) & (g994)) + ((!g747) & (!g744) & (g748) & (g962) & (!g971) & (!g994)) + ((!g747) & (!g744) & (g748) & (g962) & (!g971) & (g994)) + ((!g747) & (!g744) & (g748) & (g962) & (g971) & (!g994)) + ((!g747) & (!g744) & (g748) & (g962) & (g971) & (g994)) + ((!g747) & (g744) & (!g748) & (!g962) & (!g971) & (!g994)) + ((!g747) & (g744) & (!g748) & (!g962) & (!g971) & (g994)) + ((!g747) & (g744) & (!g748) & (g962) & (!g971) & (!g994)) + ((!g747) & (g744) & (!g748) & (g962) & (!g971) & (g994)) + ((!g747) & (g744) & (g748) & (g962) & (!g971) & (!g994)) + ((!g747) & (g744) & (g748) & (g962) & (!g971) & (g994)) + ((g747) & (!g744) & (!g748) & (!g962) & (!g971) & (!g994)) + ((g747) & (!g744) & (!g748) & (!g962) & (g971) & (!g994)) + ((g747) & (!g744) & (!g748) & (g962) & (!g971) & (!g994)) + ((g747) & (!g744) & (!g748) & (g962) & (g971) & (!g994)) + ((g747) & (!g744) & (g748) & (g962) & (!g971) & (!g994)) + ((g747) & (!g744) & (g748) & (g962) & (g971) & (!g994)) + ((g747) & (g744) & (!g748) & (!g962) & (!g971) & (!g994)) + ((g747) & (g744) & (!g748) & (g962) & (!g971) & (!g994)) + ((g747) & (g744) & (g748) & (g962) & (!g971) & (!g994)));
	assign g1192 = (((!g202) & (!g759) & (!g899) & (!g1165) & (!g1166) & (g1169)) + ((!g202) & (!g759) & (!g899) & (!g1165) & (g1166) & (!g1169)) + ((!g202) & (!g759) & (!g899) & (!g1165) & (g1166) & (g1169)) + ((!g202) & (!g759) & (!g899) & (g1165) & (g1166) & (g1169)) + ((!g202) & (!g759) & (g899) & (!g1165) & (!g1166) & (g1169)) + ((!g202) & (!g759) & (g899) & (!g1165) & (g1166) & (!g1169)) + ((!g202) & (!g759) & (g899) & (!g1165) & (g1166) & (g1169)) + ((!g202) & (!g759) & (g899) & (g1165) & (g1166) & (g1169)) + ((!g202) & (g759) & (!g899) & (!g1165) & (!g1166) & (g1169)) + ((!g202) & (g759) & (!g899) & (!g1165) & (g1166) & (!g1169)) + ((!g202) & (g759) & (!g899) & (!g1165) & (g1166) & (g1169)) + ((!g202) & (g759) & (!g899) & (g1165) & (!g1166) & (g1169)) + ((!g202) & (g759) & (!g899) & (g1165) & (g1166) & (!g1169)) + ((!g202) & (g759) & (!g899) & (g1165) & (g1166) & (g1169)) + ((!g202) & (g759) & (g899) & (!g1165) & (!g1166) & (g1169)) + ((!g202) & (g759) & (g899) & (!g1165) & (g1166) & (!g1169)) + ((!g202) & (g759) & (g899) & (!g1165) & (g1166) & (g1169)) + ((!g202) & (g759) & (g899) & (g1165) & (g1166) & (g1169)) + ((g202) & (!g759) & (!g899) & (!g1165) & (g1166) & (g1169)) + ((g202) & (!g759) & (!g899) & (g1165) & (!g1166) & (g1169)) + ((g202) & (!g759) & (!g899) & (g1165) & (g1166) & (!g1169)) + ((g202) & (!g759) & (!g899) & (g1165) & (g1166) & (g1169)) + ((g202) & (!g759) & (g899) & (!g1165) & (g1166) & (g1169)) + ((g202) & (!g759) & (g899) & (g1165) & (!g1166) & (g1169)) + ((g202) & (!g759) & (g899) & (g1165) & (g1166) & (!g1169)) + ((g202) & (!g759) & (g899) & (g1165) & (g1166) & (g1169)) + ((g202) & (g759) & (!g899) & (!g1165) & (g1166) & (g1169)) + ((g202) & (g759) & (!g899) & (g1165) & (g1166) & (g1169)) + ((g202) & (g759) & (g899) & (!g1165) & (g1166) & (g1169)) + ((g202) & (g759) & (g899) & (g1165) & (!g1166) & (g1169)) + ((g202) & (g759) & (g899) & (g1165) & (g1166) & (!g1169)) + ((g202) & (g759) & (g899) & (g1165) & (g1166) & (g1169)));
	assign g1193 = (((!g698) & (!g706) & (!g717) & (g765) & (!g825) & (!g832)) + ((!g698) & (!g706) & (!g717) & (g765) & (g825) & (g832)) + ((!g698) & (!g706) & (g717) & (g765) & (!g825) & (!g832)) + ((!g698) & (!g706) & (g717) & (g765) & (g825) & (g832)) + ((!g698) & (g706) & (!g717) & (g765) & (!g825) & (!g832)) + ((!g698) & (g706) & (!g717) & (g765) & (g825) & (g832)) + ((!g698) & (g706) & (g717) & (g765) & (!g825) & (g832)) + ((!g698) & (g706) & (g717) & (g765) & (g825) & (!g832)) + ((g698) & (!g706) & (!g717) & (g765) & (!g825) & (!g832)) + ((g698) & (!g706) & (!g717) & (g765) & (g825) & (g832)) + ((g698) & (!g706) & (g717) & (g765) & (!g825) & (g832)) + ((g698) & (!g706) & (g717) & (g765) & (g825) & (!g832)) + ((g698) & (g706) & (!g717) & (g765) & (!g825) & (g832)) + ((g698) & (g706) & (!g717) & (g765) & (g825) & (!g832)) + ((g698) & (g706) & (g717) & (g765) & (!g825) & (g832)) + ((g698) & (g706) & (g717) & (g765) & (g825) & (!g832)));
	assign g1194 = (((!g764) & (!g762) & (!g871) & (!g883) & (!g863) & (!g1193)) + ((!g764) & (!g762) & (!g871) & (!g883) & (g863) & (!g1193)) + ((!g764) & (!g762) & (!g871) & (g883) & (!g863) & (!g1193)) + ((!g764) & (!g762) & (!g871) & (g883) & (g863) & (!g1193)) + ((!g764) & (!g762) & (g871) & (!g883) & (!g863) & (!g1193)) + ((!g764) & (!g762) & (g871) & (!g883) & (g863) & (!g1193)) + ((!g764) & (!g762) & (g871) & (g883) & (!g863) & (!g1193)) + ((!g764) & (!g762) & (g871) & (g883) & (g863) & (!g1193)) + ((!g764) & (g762) & (!g871) & (!g883) & (!g863) & (!g1193)) + ((!g764) & (g762) & (!g871) & (g883) & (!g863) & (!g1193)) + ((!g764) & (g762) & (g871) & (!g883) & (!g863) & (!g1193)) + ((!g764) & (g762) & (g871) & (g883) & (!g863) & (!g1193)) + ((g764) & (!g762) & (!g871) & (g883) & (!g863) & (!g1193)) + ((g764) & (!g762) & (!g871) & (g883) & (g863) & (!g1193)) + ((g764) & (!g762) & (g871) & (!g883) & (!g863) & (!g1193)) + ((g764) & (!g762) & (g871) & (!g883) & (g863) & (!g1193)) + ((g764) & (g762) & (!g871) & (g883) & (!g863) & (!g1193)) + ((g764) & (g762) & (g871) & (!g883) & (!g863) & (!g1193)));
	assign g1195 = (((!g707) & (!g717) & (!g718) & (g847) & (!sk[53]) & (!g845)) + ((!g707) & (!g717) & (!g718) & (g847) & (!sk[53]) & (g845)) + ((!g707) & (!g717) & (g718) & (!g847) & (!sk[53]) & (!g845)) + ((!g707) & (!g717) & (g718) & (!g847) & (!sk[53]) & (g845)) + ((!g707) & (!g717) & (g718) & (!g847) & (sk[53]) & (g845)) + ((!g707) & (!g717) & (g718) & (g847) & (!sk[53]) & (!g845)) + ((!g707) & (!g717) & (g718) & (g847) & (!sk[53]) & (g845)) + ((!g707) & (!g717) & (g718) & (g847) & (sk[53]) & (g845)) + ((!g707) & (g717) & (!g718) & (!g847) & (!sk[53]) & (!g845)) + ((!g707) & (g717) & (!g718) & (!g847) & (!sk[53]) & (g845)) + ((!g707) & (g717) & (!g718) & (g847) & (!sk[53]) & (!g845)) + ((!g707) & (g717) & (!g718) & (g847) & (!sk[53]) & (g845)) + ((!g707) & (g717) & (!g718) & (g847) & (sk[53]) & (!g845)) + ((!g707) & (g717) & (!g718) & (g847) & (sk[53]) & (g845)) + ((!g707) & (g717) & (g718) & (!g847) & (!sk[53]) & (!g845)) + ((!g707) & (g717) & (g718) & (!g847) & (!sk[53]) & (g845)) + ((!g707) & (g717) & (g718) & (!g847) & (sk[53]) & (g845)) + ((!g707) & (g717) & (g718) & (g847) & (!sk[53]) & (!g845)) + ((!g707) & (g717) & (g718) & (g847) & (!sk[53]) & (g845)) + ((!g707) & (g717) & (g718) & (g847) & (sk[53]) & (!g845)) + ((!g707) & (g717) & (g718) & (g847) & (sk[53]) & (g845)) + ((g707) & (!g717) & (!g718) & (g847) & (!sk[53]) & (!g845)) + ((g707) & (!g717) & (!g718) & (g847) & (!sk[53]) & (g845)) + ((g707) & (!g717) & (!g718) & (g847) & (sk[53]) & (!g845)) + ((g707) & (!g717) & (!g718) & (g847) & (sk[53]) & (g845)) + ((g707) & (!g717) & (g718) & (!g847) & (!sk[53]) & (!g845)) + ((g707) & (!g717) & (g718) & (!g847) & (!sk[53]) & (g845)) + ((g707) & (!g717) & (g718) & (!g847) & (sk[53]) & (g845)) + ((g707) & (!g717) & (g718) & (g847) & (!sk[53]) & (!g845)) + ((g707) & (!g717) & (g718) & (g847) & (!sk[53]) & (g845)) + ((g707) & (!g717) & (g718) & (g847) & (sk[53]) & (!g845)) + ((g707) & (!g717) & (g718) & (g847) & (sk[53]) & (g845)) + ((g707) & (g717) & (!g718) & (!g847) & (!sk[53]) & (!g845)) + ((g707) & (g717) & (!g718) & (!g847) & (!sk[53]) & (g845)) + ((g707) & (g717) & (!g718) & (g847) & (!sk[53]) & (!g845)) + ((g707) & (g717) & (!g718) & (g847) & (!sk[53]) & (g845)) + ((g707) & (g717) & (g718) & (!g847) & (!sk[53]) & (!g845)) + ((g707) & (g717) & (g718) & (!g847) & (!sk[53]) & (g845)) + ((g707) & (g717) & (g718) & (!g847) & (sk[53]) & (g845)) + ((g707) & (g717) & (g718) & (g847) & (!sk[53]) & (!g845)) + ((g707) & (g717) & (g718) & (g847) & (!sk[53]) & (g845)) + ((g707) & (g717) & (g718) & (g847) & (sk[53]) & (g845)));
	assign g1196 = (((!g252) & (!g681) & (!g731) & (!g843) & (!g848) & (!g1195)) + ((!g252) & (!g681) & (!g731) & (g843) & (!g848) & (!g1195)) + ((!g252) & (!g681) & (g731) & (!g843) & (!g848) & (!g1195)) + ((!g252) & (g681) & (!g731) & (!g843) & (!g848) & (!g1195)) + ((!g252) & (g681) & (!g731) & (!g843) & (g848) & (!g1195)) + ((!g252) & (g681) & (!g731) & (g843) & (!g848) & (!g1195)) + ((!g252) & (g681) & (!g731) & (g843) & (g848) & (!g1195)) + ((!g252) & (g681) & (g731) & (!g843) & (!g848) & (!g1195)) + ((!g252) & (g681) & (g731) & (!g843) & (g848) & (!g1195)) + ((g252) & (!g681) & (!g731) & (!g843) & (!g848) & (g1195)) + ((g252) & (!g681) & (!g731) & (!g843) & (g848) & (!g1195)) + ((g252) & (!g681) & (!g731) & (!g843) & (g848) & (g1195)) + ((g252) & (!g681) & (!g731) & (g843) & (!g848) & (g1195)) + ((g252) & (!g681) & (!g731) & (g843) & (g848) & (!g1195)) + ((g252) & (!g681) & (!g731) & (g843) & (g848) & (g1195)) + ((g252) & (!g681) & (g731) & (!g843) & (!g848) & (g1195)) + ((g252) & (!g681) & (g731) & (!g843) & (g848) & (!g1195)) + ((g252) & (!g681) & (g731) & (!g843) & (g848) & (g1195)) + ((g252) & (!g681) & (g731) & (g843) & (!g848) & (!g1195)) + ((g252) & (!g681) & (g731) & (g843) & (!g848) & (g1195)) + ((g252) & (!g681) & (g731) & (g843) & (g848) & (!g1195)) + ((g252) & (!g681) & (g731) & (g843) & (g848) & (g1195)) + ((g252) & (g681) & (!g731) & (!g843) & (!g848) & (g1195)) + ((g252) & (g681) & (!g731) & (!g843) & (g848) & (g1195)) + ((g252) & (g681) & (!g731) & (g843) & (!g848) & (g1195)) + ((g252) & (g681) & (!g731) & (g843) & (g848) & (g1195)) + ((g252) & (g681) & (g731) & (!g843) & (!g848) & (g1195)) + ((g252) & (g681) & (g731) & (!g843) & (g848) & (g1195)) + ((g252) & (g681) & (g731) & (g843) & (!g848) & (!g1195)) + ((g252) & (g681) & (g731) & (g843) & (!g848) & (g1195)) + ((g252) & (g681) & (g731) & (g843) & (g848) & (!g1195)) + ((g252) & (g681) & (g731) & (g843) & (g848) & (g1195)));
	assign g1197 = (((!g252) & (!g683) & (!g719) & (!sk[55]) & (g729) & (!g1168)) + ((!g252) & (!g683) & (!g719) & (!sk[55]) & (g729) & (g1168)) + ((!g252) & (!g683) & (g719) & (!sk[55]) & (!g729) & (!g1168)) + ((!g252) & (!g683) & (g719) & (!sk[55]) & (!g729) & (g1168)) + ((!g252) & (!g683) & (g719) & (!sk[55]) & (g729) & (!g1168)) + ((!g252) & (!g683) & (g719) & (!sk[55]) & (g729) & (g1168)) + ((!g252) & (g683) & (!g719) & (!sk[55]) & (!g729) & (!g1168)) + ((!g252) & (g683) & (!g719) & (!sk[55]) & (!g729) & (g1168)) + ((!g252) & (g683) & (!g719) & (!sk[55]) & (g729) & (!g1168)) + ((!g252) & (g683) & (!g719) & (!sk[55]) & (g729) & (g1168)) + ((!g252) & (g683) & (!g719) & (sk[55]) & (!g729) & (g1168)) + ((!g252) & (g683) & (!g719) & (sk[55]) & (g729) & (g1168)) + ((!g252) & (g683) & (g719) & (!sk[55]) & (!g729) & (!g1168)) + ((!g252) & (g683) & (g719) & (!sk[55]) & (!g729) & (g1168)) + ((!g252) & (g683) & (g719) & (!sk[55]) & (g729) & (!g1168)) + ((!g252) & (g683) & (g719) & (!sk[55]) & (g729) & (g1168)) + ((!g252) & (g683) & (g719) & (sk[55]) & (!g729) & (g1168)) + ((!g252) & (g683) & (g719) & (sk[55]) & (g729) & (g1168)) + ((g252) & (!g683) & (!g719) & (!sk[55]) & (g729) & (!g1168)) + ((g252) & (!g683) & (!g719) & (!sk[55]) & (g729) & (g1168)) + ((g252) & (!g683) & (!g719) & (sk[55]) & (!g729) & (!g1168)) + ((g252) & (!g683) & (!g719) & (sk[55]) & (g729) & (g1168)) + ((g252) & (!g683) & (g719) & (!sk[55]) & (!g729) & (!g1168)) + ((g252) & (!g683) & (g719) & (!sk[55]) & (!g729) & (g1168)) + ((g252) & (!g683) & (g719) & (!sk[55]) & (g729) & (!g1168)) + ((g252) & (!g683) & (g719) & (!sk[55]) & (g729) & (g1168)) + ((g252) & (!g683) & (g719) & (sk[55]) & (!g729) & (!g1168)) + ((g252) & (!g683) & (g719) & (sk[55]) & (!g729) & (g1168)) + ((g252) & (g683) & (!g719) & (!sk[55]) & (!g729) & (!g1168)) + ((g252) & (g683) & (!g719) & (!sk[55]) & (!g729) & (g1168)) + ((g252) & (g683) & (!g719) & (!sk[55]) & (g729) & (!g1168)) + ((g252) & (g683) & (!g719) & (!sk[55]) & (g729) & (g1168)) + ((g252) & (g683) & (!g719) & (sk[55]) & (!g729) & (!g1168)) + ((g252) & (g683) & (!g719) & (sk[55]) & (!g729) & (g1168)) + ((g252) & (g683) & (g719) & (!sk[55]) & (!g729) & (!g1168)) + ((g252) & (g683) & (g719) & (!sk[55]) & (!g729) & (g1168)) + ((g252) & (g683) & (g719) & (!sk[55]) & (g729) & (!g1168)) + ((g252) & (g683) & (g719) & (!sk[55]) & (g729) & (g1168)) + ((g252) & (g683) & (g719) & (sk[55]) & (!g729) & (g1168)) + ((g252) & (g683) & (g719) & (sk[55]) & (g729) & (!g1168)));
	assign g1198 = (((!g202) & (!g759) & (!g895) & (!g1194) & (!g1196) & (!g1197)) + ((!g202) & (!g759) & (!g895) & (!g1194) & (g1196) & (g1197)) + ((!g202) & (!g759) & (!g895) & (g1194) & (!g1196) & (g1197)) + ((!g202) & (!g759) & (!g895) & (g1194) & (g1196) & (!g1197)) + ((!g202) & (!g759) & (g895) & (!g1194) & (!g1196) & (!g1197)) + ((!g202) & (!g759) & (g895) & (!g1194) & (g1196) & (g1197)) + ((!g202) & (!g759) & (g895) & (g1194) & (!g1196) & (g1197)) + ((!g202) & (!g759) & (g895) & (g1194) & (g1196) & (!g1197)) + ((!g202) & (g759) & (!g895) & (!g1194) & (!g1196) & (!g1197)) + ((!g202) & (g759) & (!g895) & (!g1194) & (g1196) & (g1197)) + ((!g202) & (g759) & (!g895) & (g1194) & (!g1196) & (g1197)) + ((!g202) & (g759) & (!g895) & (g1194) & (g1196) & (!g1197)) + ((!g202) & (g759) & (g895) & (!g1194) & (!g1196) & (!g1197)) + ((!g202) & (g759) & (g895) & (!g1194) & (g1196) & (g1197)) + ((!g202) & (g759) & (g895) & (g1194) & (!g1196) & (!g1197)) + ((!g202) & (g759) & (g895) & (g1194) & (g1196) & (g1197)) + ((g202) & (!g759) & (!g895) & (!g1194) & (!g1196) & (g1197)) + ((g202) & (!g759) & (!g895) & (!g1194) & (g1196) & (!g1197)) + ((g202) & (!g759) & (!g895) & (g1194) & (!g1196) & (!g1197)) + ((g202) & (!g759) & (!g895) & (g1194) & (g1196) & (g1197)) + ((g202) & (!g759) & (g895) & (!g1194) & (!g1196) & (g1197)) + ((g202) & (!g759) & (g895) & (!g1194) & (g1196) & (!g1197)) + ((g202) & (!g759) & (g895) & (g1194) & (!g1196) & (!g1197)) + ((g202) & (!g759) & (g895) & (g1194) & (g1196) & (g1197)) + ((g202) & (g759) & (!g895) & (!g1194) & (!g1196) & (g1197)) + ((g202) & (g759) & (!g895) & (!g1194) & (g1196) & (!g1197)) + ((g202) & (g759) & (!g895) & (g1194) & (!g1196) & (!g1197)) + ((g202) & (g759) & (!g895) & (g1194) & (g1196) & (g1197)) + ((g202) & (g759) & (g895) & (!g1194) & (!g1196) & (g1197)) + ((g202) & (g759) & (g895) & (!g1194) & (g1196) & (!g1197)) + ((g202) & (g759) & (g895) & (g1194) & (!g1196) & (g1197)) + ((g202) & (g759) & (g895) & (g1194) & (g1196) & (!g1197)));
	assign g1199 = (((!g200) & (!g742) & (!g995) & (!g1191) & (!g1192) & (!g1198)) + ((!g200) & (!g742) & (!g995) & (!g1191) & (g1192) & (g1198)) + ((!g200) & (!g742) & (!g995) & (g1191) & (!g1192) & (g1198)) + ((!g200) & (!g742) & (!g995) & (g1191) & (g1192) & (!g1198)) + ((!g200) & (!g742) & (g995) & (!g1191) & (!g1192) & (!g1198)) + ((!g200) & (!g742) & (g995) & (!g1191) & (g1192) & (g1198)) + ((!g200) & (!g742) & (g995) & (g1191) & (!g1192) & (g1198)) + ((!g200) & (!g742) & (g995) & (g1191) & (g1192) & (!g1198)) + ((!g200) & (g742) & (!g995) & (!g1191) & (!g1192) & (!g1198)) + ((!g200) & (g742) & (!g995) & (!g1191) & (g1192) & (g1198)) + ((!g200) & (g742) & (!g995) & (g1191) & (!g1192) & (g1198)) + ((!g200) & (g742) & (!g995) & (g1191) & (g1192) & (!g1198)) + ((!g200) & (g742) & (g995) & (!g1191) & (!g1192) & (!g1198)) + ((!g200) & (g742) & (g995) & (!g1191) & (g1192) & (g1198)) + ((!g200) & (g742) & (g995) & (g1191) & (!g1192) & (!g1198)) + ((!g200) & (g742) & (g995) & (g1191) & (g1192) & (g1198)) + ((g200) & (!g742) & (!g995) & (!g1191) & (!g1192) & (g1198)) + ((g200) & (!g742) & (!g995) & (!g1191) & (g1192) & (!g1198)) + ((g200) & (!g742) & (!g995) & (g1191) & (!g1192) & (!g1198)) + ((g200) & (!g742) & (!g995) & (g1191) & (g1192) & (g1198)) + ((g200) & (!g742) & (g995) & (!g1191) & (!g1192) & (g1198)) + ((g200) & (!g742) & (g995) & (!g1191) & (g1192) & (!g1198)) + ((g200) & (!g742) & (g995) & (g1191) & (!g1192) & (!g1198)) + ((g200) & (!g742) & (g995) & (g1191) & (g1192) & (g1198)) + ((g200) & (g742) & (!g995) & (!g1191) & (!g1192) & (g1198)) + ((g200) & (g742) & (!g995) & (!g1191) & (g1192) & (!g1198)) + ((g200) & (g742) & (!g995) & (g1191) & (!g1192) & (!g1198)) + ((g200) & (g742) & (!g995) & (g1191) & (g1192) & (g1198)) + ((g200) & (g742) & (g995) & (!g1191) & (!g1192) & (g1198)) + ((g200) & (g742) & (g995) & (!g1191) & (g1192) & (!g1198)) + ((g200) & (g742) & (g995) & (g1191) & (!g1192) & (g1198)) + ((g200) & (g742) & (g995) & (g1191) & (g1192) & (!g1198)));
	assign g1200 = (((!g2) & (!g732) & (!g1188) & (!g1189) & (!g1190) & (g1199)) + ((!g2) & (!g732) & (!g1188) & (!g1189) & (g1190) & (!g1199)) + ((!g2) & (!g732) & (!g1188) & (g1189) & (!g1190) & (!g1199)) + ((!g2) & (!g732) & (!g1188) & (g1189) & (g1190) & (g1199)) + ((!g2) & (!g732) & (g1188) & (!g1189) & (!g1190) & (g1199)) + ((!g2) & (!g732) & (g1188) & (!g1189) & (g1190) & (!g1199)) + ((!g2) & (!g732) & (g1188) & (g1189) & (!g1190) & (!g1199)) + ((!g2) & (!g732) & (g1188) & (g1189) & (g1190) & (g1199)) + ((!g2) & (g732) & (!g1188) & (!g1189) & (!g1190) & (g1199)) + ((!g2) & (g732) & (!g1188) & (!g1189) & (g1190) & (!g1199)) + ((!g2) & (g732) & (!g1188) & (g1189) & (!g1190) & (!g1199)) + ((!g2) & (g732) & (!g1188) & (g1189) & (g1190) & (g1199)) + ((!g2) & (g732) & (g1188) & (!g1189) & (!g1190) & (!g1199)) + ((!g2) & (g732) & (g1188) & (!g1189) & (g1190) & (g1199)) + ((!g2) & (g732) & (g1188) & (g1189) & (!g1190) & (!g1199)) + ((!g2) & (g732) & (g1188) & (g1189) & (g1190) & (g1199)) + ((g2) & (!g732) & (!g1188) & (!g1189) & (!g1190) & (!g1199)) + ((g2) & (!g732) & (!g1188) & (!g1189) & (g1190) & (g1199)) + ((g2) & (!g732) & (!g1188) & (g1189) & (!g1190) & (g1199)) + ((g2) & (!g732) & (!g1188) & (g1189) & (g1190) & (!g1199)) + ((g2) & (!g732) & (g1188) & (!g1189) & (!g1190) & (!g1199)) + ((g2) & (!g732) & (g1188) & (!g1189) & (g1190) & (g1199)) + ((g2) & (!g732) & (g1188) & (g1189) & (!g1190) & (g1199)) + ((g2) & (!g732) & (g1188) & (g1189) & (g1190) & (!g1199)) + ((g2) & (g732) & (!g1188) & (!g1189) & (!g1190) & (!g1199)) + ((g2) & (g732) & (!g1188) & (!g1189) & (g1190) & (g1199)) + ((g2) & (g732) & (!g1188) & (g1189) & (!g1190) & (g1199)) + ((g2) & (g732) & (!g1188) & (g1189) & (g1190) & (!g1199)) + ((g2) & (g732) & (g1188) & (!g1189) & (!g1190) & (g1199)) + ((g2) & (g732) & (g1188) & (!g1189) & (g1190) & (!g1199)) + ((g2) & (g732) & (g1188) & (g1189) & (!g1190) & (g1199)) + ((g2) & (g732) & (g1188) & (g1189) & (g1190) & (!g1199)));
	assign g1201 = (((!g1161) & (!g1162) & (!sk[59]) & (!g1174) & (g1187) & (!g1200)) + ((!g1161) & (!g1162) & (!sk[59]) & (!g1174) & (g1187) & (g1200)) + ((!g1161) & (!g1162) & (!sk[59]) & (g1174) & (!g1187) & (!g1200)) + ((!g1161) & (!g1162) & (!sk[59]) & (g1174) & (!g1187) & (g1200)) + ((!g1161) & (!g1162) & (!sk[59]) & (g1174) & (g1187) & (!g1200)) + ((!g1161) & (!g1162) & (!sk[59]) & (g1174) & (g1187) & (g1200)) + ((!g1161) & (!g1162) & (sk[59]) & (!g1174) & (!g1187) & (g1200)) + ((!g1161) & (!g1162) & (sk[59]) & (!g1174) & (g1187) & (!g1200)) + ((!g1161) & (!g1162) & (sk[59]) & (g1174) & (!g1187) & (!g1200)) + ((!g1161) & (!g1162) & (sk[59]) & (g1174) & (g1187) & (g1200)) + ((!g1161) & (g1162) & (!sk[59]) & (!g1174) & (!g1187) & (!g1200)) + ((!g1161) & (g1162) & (!sk[59]) & (!g1174) & (!g1187) & (g1200)) + ((!g1161) & (g1162) & (!sk[59]) & (!g1174) & (g1187) & (!g1200)) + ((!g1161) & (g1162) & (!sk[59]) & (!g1174) & (g1187) & (g1200)) + ((!g1161) & (g1162) & (!sk[59]) & (g1174) & (!g1187) & (!g1200)) + ((!g1161) & (g1162) & (!sk[59]) & (g1174) & (!g1187) & (g1200)) + ((!g1161) & (g1162) & (!sk[59]) & (g1174) & (g1187) & (!g1200)) + ((!g1161) & (g1162) & (!sk[59]) & (g1174) & (g1187) & (g1200)) + ((!g1161) & (g1162) & (sk[59]) & (!g1174) & (!g1187) & (!g1200)) + ((!g1161) & (g1162) & (sk[59]) & (!g1174) & (g1187) & (g1200)) + ((!g1161) & (g1162) & (sk[59]) & (g1174) & (!g1187) & (!g1200)) + ((!g1161) & (g1162) & (sk[59]) & (g1174) & (g1187) & (g1200)) + ((g1161) & (!g1162) & (!sk[59]) & (!g1174) & (g1187) & (!g1200)) + ((g1161) & (!g1162) & (!sk[59]) & (!g1174) & (g1187) & (g1200)) + ((g1161) & (!g1162) & (!sk[59]) & (g1174) & (!g1187) & (!g1200)) + ((g1161) & (!g1162) & (!sk[59]) & (g1174) & (!g1187) & (g1200)) + ((g1161) & (!g1162) & (!sk[59]) & (g1174) & (g1187) & (!g1200)) + ((g1161) & (!g1162) & (!sk[59]) & (g1174) & (g1187) & (g1200)) + ((g1161) & (!g1162) & (sk[59]) & (!g1174) & (!g1187) & (g1200)) + ((g1161) & (!g1162) & (sk[59]) & (!g1174) & (g1187) & (!g1200)) + ((g1161) & (!g1162) & (sk[59]) & (g1174) & (!g1187) & (g1200)) + ((g1161) & (!g1162) & (sk[59]) & (g1174) & (g1187) & (!g1200)) + ((g1161) & (g1162) & (!sk[59]) & (!g1174) & (!g1187) & (!g1200)) + ((g1161) & (g1162) & (!sk[59]) & (!g1174) & (!g1187) & (g1200)) + ((g1161) & (g1162) & (!sk[59]) & (!g1174) & (g1187) & (!g1200)) + ((g1161) & (g1162) & (!sk[59]) & (!g1174) & (g1187) & (g1200)) + ((g1161) & (g1162) & (!sk[59]) & (g1174) & (!g1187) & (!g1200)) + ((g1161) & (g1162) & (!sk[59]) & (g1174) & (!g1187) & (g1200)) + ((g1161) & (g1162) & (!sk[59]) & (g1174) & (g1187) & (!g1200)) + ((g1161) & (g1162) & (!sk[59]) & (g1174) & (g1187) & (g1200)) + ((g1161) & (g1162) & (sk[59]) & (!g1174) & (!g1187) & (g1200)) + ((g1161) & (g1162) & (sk[59]) & (!g1174) & (g1187) & (!g1200)) + ((g1161) & (g1162) & (sk[59]) & (g1174) & (!g1187) & (!g1200)) + ((g1161) & (g1162) & (sk[59]) & (g1174) & (g1187) & (g1200)));
	assign g1202 = (((!g16) & (!g99) & (!sk[60]) & (!g18) & (g66) & (!g86)) + ((!g16) & (!g99) & (!sk[60]) & (!g18) & (g66) & (g86)) + ((!g16) & (!g99) & (!sk[60]) & (g18) & (!g66) & (!g86)) + ((!g16) & (!g99) & (!sk[60]) & (g18) & (!g66) & (g86)) + ((!g16) & (!g99) & (!sk[60]) & (g18) & (g66) & (!g86)) + ((!g16) & (!g99) & (!sk[60]) & (g18) & (g66) & (g86)) + ((!g16) & (!g99) & (sk[60]) & (!g18) & (!g66) & (!g86)) + ((!g16) & (!g99) & (sk[60]) & (!g18) & (g66) & (!g86)) + ((!g16) & (!g99) & (sk[60]) & (g18) & (!g66) & (!g86)) + ((!g16) & (!g99) & (sk[60]) & (g18) & (g66) & (!g86)) + ((!g16) & (g99) & (!sk[60]) & (!g18) & (!g66) & (!g86)) + ((!g16) & (g99) & (!sk[60]) & (!g18) & (!g66) & (g86)) + ((!g16) & (g99) & (!sk[60]) & (!g18) & (g66) & (!g86)) + ((!g16) & (g99) & (!sk[60]) & (!g18) & (g66) & (g86)) + ((!g16) & (g99) & (!sk[60]) & (g18) & (!g66) & (!g86)) + ((!g16) & (g99) & (!sk[60]) & (g18) & (!g66) & (g86)) + ((!g16) & (g99) & (!sk[60]) & (g18) & (g66) & (!g86)) + ((!g16) & (g99) & (!sk[60]) & (g18) & (g66) & (g86)) + ((!g16) & (g99) & (sk[60]) & (!g18) & (!g66) & (!g86)) + ((!g16) & (g99) & (sk[60]) & (!g18) & (g66) & (!g86)) + ((g16) & (!g99) & (!sk[60]) & (!g18) & (g66) & (!g86)) + ((g16) & (!g99) & (!sk[60]) & (!g18) & (g66) & (g86)) + ((g16) & (!g99) & (!sk[60]) & (g18) & (!g66) & (!g86)) + ((g16) & (!g99) & (!sk[60]) & (g18) & (!g66) & (g86)) + ((g16) & (!g99) & (!sk[60]) & (g18) & (g66) & (!g86)) + ((g16) & (!g99) & (!sk[60]) & (g18) & (g66) & (g86)) + ((g16) & (!g99) & (sk[60]) & (!g18) & (!g66) & (!g86)) + ((g16) & (!g99) & (sk[60]) & (g18) & (!g66) & (!g86)) + ((g16) & (g99) & (!sk[60]) & (!g18) & (!g66) & (!g86)) + ((g16) & (g99) & (!sk[60]) & (!g18) & (!g66) & (g86)) + ((g16) & (g99) & (!sk[60]) & (!g18) & (g66) & (!g86)) + ((g16) & (g99) & (!sk[60]) & (!g18) & (g66) & (g86)) + ((g16) & (g99) & (!sk[60]) & (g18) & (!g66) & (!g86)) + ((g16) & (g99) & (!sk[60]) & (g18) & (!g66) & (g86)) + ((g16) & (g99) & (!sk[60]) & (g18) & (g66) & (!g86)) + ((g16) & (g99) & (!sk[60]) & (g18) & (g66) & (g86)) + ((g16) & (g99) & (sk[60]) & (!g18) & (!g66) & (!g86)));
	assign g1203 = (((!sk[61]) & (!g9) & (!g70) & (!g25) & (g27)) + ((!sk[61]) & (!g9) & (!g70) & (g25) & (g27)) + ((!sk[61]) & (!g9) & (g70) & (!g25) & (g27)) + ((!sk[61]) & (!g9) & (g70) & (g25) & (g27)) + ((!sk[61]) & (g9) & (!g70) & (!g25) & (!g27)) + ((!sk[61]) & (g9) & (!g70) & (!g25) & (g27)) + ((!sk[61]) & (g9) & (!g70) & (g25) & (!g27)) + ((!sk[61]) & (g9) & (!g70) & (g25) & (g27)) + ((!sk[61]) & (g9) & (g70) & (!g25) & (!g27)) + ((!sk[61]) & (g9) & (g70) & (!g25) & (g27)) + ((!sk[61]) & (g9) & (g70) & (g25) & (!g27)) + ((!sk[61]) & (g9) & (g70) & (g25) & (g27)) + ((sk[61]) & (!g9) & (g70) & (!g25) & (g27)) + ((sk[61]) & (!g9) & (g70) & (g25) & (g27)) + ((sk[61]) & (g9) & (!g70) & (g25) & (!g27)) + ((sk[61]) & (g9) & (!g70) & (g25) & (g27)) + ((sk[61]) & (g9) & (g70) & (!g25) & (g27)) + ((sk[61]) & (g9) & (g70) & (g25) & (!g27)) + ((sk[61]) & (g9) & (g70) & (g25) & (g27)));
	assign g1204 = (((!sk[62]) & (!g19) & (!g13) & (!g36) & (g1203)) + ((!sk[62]) & (!g19) & (!g13) & (g36) & (g1203)) + ((!sk[62]) & (!g19) & (g13) & (!g36) & (g1203)) + ((!sk[62]) & (!g19) & (g13) & (g36) & (g1203)) + ((!sk[62]) & (g19) & (!g13) & (!g36) & (!g1203)) + ((!sk[62]) & (g19) & (!g13) & (!g36) & (g1203)) + ((!sk[62]) & (g19) & (!g13) & (g36) & (!g1203)) + ((!sk[62]) & (g19) & (!g13) & (g36) & (g1203)) + ((!sk[62]) & (g19) & (g13) & (!g36) & (!g1203)) + ((!sk[62]) & (g19) & (g13) & (!g36) & (g1203)) + ((!sk[62]) & (g19) & (g13) & (g36) & (!g1203)) + ((!sk[62]) & (g19) & (g13) & (g36) & (g1203)) + ((sk[62]) & (!g19) & (!g13) & (!g36) & (!g1203)));
	assign g1205 = (((!g52) & (!g596) & (!g1102) & (!sk[63]) & (g1204)) + ((!g52) & (!g596) & (g1102) & (!sk[63]) & (g1204)) + ((!g52) & (g596) & (!g1102) & (!sk[63]) & (g1204)) + ((!g52) & (g596) & (g1102) & (!sk[63]) & (g1204)) + ((g52) & (!g596) & (!g1102) & (!sk[63]) & (!g1204)) + ((g52) & (!g596) & (!g1102) & (!sk[63]) & (g1204)) + ((g52) & (!g596) & (g1102) & (!sk[63]) & (!g1204)) + ((g52) & (!g596) & (g1102) & (!sk[63]) & (g1204)) + ((g52) & (g596) & (!g1102) & (!sk[63]) & (!g1204)) + ((g52) & (g596) & (!g1102) & (!sk[63]) & (g1204)) + ((g52) & (g596) & (g1102) & (!sk[63]) & (!g1204)) + ((g52) & (g596) & (g1102) & (!sk[63]) & (g1204)) + ((g52) & (g596) & (g1102) & (sk[63]) & (g1204)));
	assign g1206 = (((g1006) & (!g587) & (g877) & (g1076) & (g1202) & (g1205)));
	assign g1207 = (((!g1160) & (!g1175) & (!sk[65]) & (!g1182) & (g1201) & (!g1206)) + ((!g1160) & (!g1175) & (!sk[65]) & (!g1182) & (g1201) & (g1206)) + ((!g1160) & (!g1175) & (!sk[65]) & (g1182) & (!g1201) & (!g1206)) + ((!g1160) & (!g1175) & (!sk[65]) & (g1182) & (!g1201) & (g1206)) + ((!g1160) & (!g1175) & (!sk[65]) & (g1182) & (g1201) & (!g1206)) + ((!g1160) & (!g1175) & (!sk[65]) & (g1182) & (g1201) & (g1206)) + ((!g1160) & (!g1175) & (sk[65]) & (!g1182) & (!g1201) & (!g1206)) + ((!g1160) & (!g1175) & (sk[65]) & (!g1182) & (g1201) & (g1206)) + ((!g1160) & (!g1175) & (sk[65]) & (g1182) & (!g1201) & (!g1206)) + ((!g1160) & (!g1175) & (sk[65]) & (g1182) & (g1201) & (g1206)) + ((!g1160) & (g1175) & (!sk[65]) & (!g1182) & (!g1201) & (!g1206)) + ((!g1160) & (g1175) & (!sk[65]) & (!g1182) & (!g1201) & (g1206)) + ((!g1160) & (g1175) & (!sk[65]) & (!g1182) & (g1201) & (!g1206)) + ((!g1160) & (g1175) & (!sk[65]) & (!g1182) & (g1201) & (g1206)) + ((!g1160) & (g1175) & (!sk[65]) & (g1182) & (!g1201) & (!g1206)) + ((!g1160) & (g1175) & (!sk[65]) & (g1182) & (!g1201) & (g1206)) + ((!g1160) & (g1175) & (!sk[65]) & (g1182) & (g1201) & (!g1206)) + ((!g1160) & (g1175) & (!sk[65]) & (g1182) & (g1201) & (g1206)) + ((!g1160) & (g1175) & (sk[65]) & (!g1182) & (!g1201) & (g1206)) + ((!g1160) & (g1175) & (sk[65]) & (!g1182) & (g1201) & (!g1206)) + ((!g1160) & (g1175) & (sk[65]) & (g1182) & (!g1201) & (!g1206)) + ((!g1160) & (g1175) & (sk[65]) & (g1182) & (g1201) & (g1206)) + ((g1160) & (!g1175) & (!sk[65]) & (!g1182) & (g1201) & (!g1206)) + ((g1160) & (!g1175) & (!sk[65]) & (!g1182) & (g1201) & (g1206)) + ((g1160) & (!g1175) & (!sk[65]) & (g1182) & (!g1201) & (!g1206)) + ((g1160) & (!g1175) & (!sk[65]) & (g1182) & (!g1201) & (g1206)) + ((g1160) & (!g1175) & (!sk[65]) & (g1182) & (g1201) & (!g1206)) + ((g1160) & (!g1175) & (!sk[65]) & (g1182) & (g1201) & (g1206)) + ((g1160) & (!g1175) & (sk[65]) & (!g1182) & (!g1201) & (g1206)) + ((g1160) & (!g1175) & (sk[65]) & (!g1182) & (g1201) & (!g1206)) + ((g1160) & (!g1175) & (sk[65]) & (g1182) & (!g1201) & (!g1206)) + ((g1160) & (!g1175) & (sk[65]) & (g1182) & (g1201) & (g1206)) + ((g1160) & (g1175) & (!sk[65]) & (!g1182) & (!g1201) & (!g1206)) + ((g1160) & (g1175) & (!sk[65]) & (!g1182) & (!g1201) & (g1206)) + ((g1160) & (g1175) & (!sk[65]) & (!g1182) & (g1201) & (!g1206)) + ((g1160) & (g1175) & (!sk[65]) & (!g1182) & (g1201) & (g1206)) + ((g1160) & (g1175) & (!sk[65]) & (g1182) & (!g1201) & (!g1206)) + ((g1160) & (g1175) & (!sk[65]) & (g1182) & (!g1201) & (g1206)) + ((g1160) & (g1175) & (!sk[65]) & (g1182) & (g1201) & (!g1206)) + ((g1160) & (g1175) & (!sk[65]) & (g1182) & (g1201) & (g1206)) + ((g1160) & (g1175) & (sk[65]) & (!g1182) & (!g1201) & (g1206)) + ((g1160) & (g1175) & (sk[65]) & (!g1182) & (g1201) & (!g1206)) + ((g1160) & (g1175) & (sk[65]) & (g1182) & (!g1201) & (g1206)) + ((g1160) & (g1175) & (sk[65]) & (g1182) & (g1201) & (!g1206)));
	assign g1208 = (((!g1068) & (!g1185) & (!g1186) & (!sk[66]) & (g1207)) + ((!g1068) & (!g1185) & (!g1186) & (sk[66]) & (g1207)) + ((!g1068) & (!g1185) & (g1186) & (!sk[66]) & (g1207)) + ((!g1068) & (!g1185) & (g1186) & (sk[66]) & (!g1207)) + ((!g1068) & (g1185) & (!g1186) & (!sk[66]) & (g1207)) + ((!g1068) & (g1185) & (!g1186) & (sk[66]) & (g1207)) + ((!g1068) & (g1185) & (g1186) & (!sk[66]) & (g1207)) + ((!g1068) & (g1185) & (g1186) & (sk[66]) & (!g1207)) + ((g1068) & (!g1185) & (!g1186) & (!sk[66]) & (!g1207)) + ((g1068) & (!g1185) & (!g1186) & (!sk[66]) & (g1207)) + ((g1068) & (!g1185) & (!g1186) & (sk[66]) & (!g1207)) + ((g1068) & (!g1185) & (g1186) & (!sk[66]) & (!g1207)) + ((g1068) & (!g1185) & (g1186) & (!sk[66]) & (g1207)) + ((g1068) & (!g1185) & (g1186) & (sk[66]) & (g1207)) + ((g1068) & (g1185) & (!g1186) & (!sk[66]) & (!g1207)) + ((g1068) & (g1185) & (!g1186) & (!sk[66]) & (g1207)) + ((g1068) & (g1185) & (!g1186) & (sk[66]) & (g1207)) + ((g1068) & (g1185) & (g1186) & (!sk[66]) & (!g1207)) + ((g1068) & (g1185) & (g1186) & (!sk[66]) & (g1207)) + ((g1068) & (g1185) & (g1186) & (sk[66]) & (!g1207)));
	assign g1209 = (((!g1160) & (!g1175) & (!sk[67]) & (!g1182) & (g1201) & (!g1206)) + ((!g1160) & (!g1175) & (!sk[67]) & (!g1182) & (g1201) & (g1206)) + ((!g1160) & (!g1175) & (!sk[67]) & (g1182) & (!g1201) & (!g1206)) + ((!g1160) & (!g1175) & (!sk[67]) & (g1182) & (!g1201) & (g1206)) + ((!g1160) & (!g1175) & (!sk[67]) & (g1182) & (g1201) & (!g1206)) + ((!g1160) & (!g1175) & (!sk[67]) & (g1182) & (g1201) & (g1206)) + ((!g1160) & (!g1175) & (sk[67]) & (!g1182) & (!g1201) & (!g1206)) + ((!g1160) & (!g1175) & (sk[67]) & (g1182) & (!g1201) & (!g1206)) + ((!g1160) & (g1175) & (!sk[67]) & (!g1182) & (!g1201) & (!g1206)) + ((!g1160) & (g1175) & (!sk[67]) & (!g1182) & (!g1201) & (g1206)) + ((!g1160) & (g1175) & (!sk[67]) & (!g1182) & (g1201) & (!g1206)) + ((!g1160) & (g1175) & (!sk[67]) & (!g1182) & (g1201) & (g1206)) + ((!g1160) & (g1175) & (!sk[67]) & (g1182) & (!g1201) & (!g1206)) + ((!g1160) & (g1175) & (!sk[67]) & (g1182) & (!g1201) & (g1206)) + ((!g1160) & (g1175) & (!sk[67]) & (g1182) & (g1201) & (!g1206)) + ((!g1160) & (g1175) & (!sk[67]) & (g1182) & (g1201) & (g1206)) + ((!g1160) & (g1175) & (sk[67]) & (!g1182) & (!g1201) & (!g1206)) + ((!g1160) & (g1175) & (sk[67]) & (!g1182) & (!g1201) & (g1206)) + ((!g1160) & (g1175) & (sk[67]) & (!g1182) & (g1201) & (!g1206)) + ((!g1160) & (g1175) & (sk[67]) & (g1182) & (!g1201) & (!g1206)) + ((g1160) & (!g1175) & (!sk[67]) & (!g1182) & (g1201) & (!g1206)) + ((g1160) & (!g1175) & (!sk[67]) & (!g1182) & (g1201) & (g1206)) + ((g1160) & (!g1175) & (!sk[67]) & (g1182) & (!g1201) & (!g1206)) + ((g1160) & (!g1175) & (!sk[67]) & (g1182) & (!g1201) & (g1206)) + ((g1160) & (!g1175) & (!sk[67]) & (g1182) & (g1201) & (!g1206)) + ((g1160) & (!g1175) & (!sk[67]) & (g1182) & (g1201) & (g1206)) + ((g1160) & (!g1175) & (sk[67]) & (!g1182) & (!g1201) & (!g1206)) + ((g1160) & (!g1175) & (sk[67]) & (!g1182) & (!g1201) & (g1206)) + ((g1160) & (!g1175) & (sk[67]) & (!g1182) & (g1201) & (!g1206)) + ((g1160) & (!g1175) & (sk[67]) & (g1182) & (!g1201) & (!g1206)) + ((g1160) & (g1175) & (!sk[67]) & (!g1182) & (!g1201) & (!g1206)) + ((g1160) & (g1175) & (!sk[67]) & (!g1182) & (!g1201) & (g1206)) + ((g1160) & (g1175) & (!sk[67]) & (!g1182) & (g1201) & (!g1206)) + ((g1160) & (g1175) & (!sk[67]) & (!g1182) & (g1201) & (g1206)) + ((g1160) & (g1175) & (!sk[67]) & (g1182) & (!g1201) & (!g1206)) + ((g1160) & (g1175) & (!sk[67]) & (g1182) & (!g1201) & (g1206)) + ((g1160) & (g1175) & (!sk[67]) & (g1182) & (g1201) & (!g1206)) + ((g1160) & (g1175) & (!sk[67]) & (g1182) & (g1201) & (g1206)) + ((g1160) & (g1175) & (sk[67]) & (!g1182) & (!g1201) & (!g1206)) + ((g1160) & (g1175) & (sk[67]) & (!g1182) & (!g1201) & (g1206)) + ((g1160) & (g1175) & (sk[67]) & (!g1182) & (g1201) & (!g1206)) + ((g1160) & (g1175) & (sk[67]) & (g1182) & (!g1201) & (!g1206)) + ((g1160) & (g1175) & (sk[67]) & (g1182) & (!g1201) & (g1206)) + ((g1160) & (g1175) & (sk[67]) & (g1182) & (g1201) & (!g1206)));
	assign g1210 = (((!sk[68]) & (!g1161) & (!g1162) & (!g1174) & (g1187) & (!g1200)) + ((!sk[68]) & (!g1161) & (!g1162) & (!g1174) & (g1187) & (g1200)) + ((!sk[68]) & (!g1161) & (!g1162) & (g1174) & (!g1187) & (!g1200)) + ((!sk[68]) & (!g1161) & (!g1162) & (g1174) & (!g1187) & (g1200)) + ((!sk[68]) & (!g1161) & (!g1162) & (g1174) & (g1187) & (!g1200)) + ((!sk[68]) & (!g1161) & (!g1162) & (g1174) & (g1187) & (g1200)) + ((!sk[68]) & (!g1161) & (g1162) & (!g1174) & (!g1187) & (!g1200)) + ((!sk[68]) & (!g1161) & (g1162) & (!g1174) & (!g1187) & (g1200)) + ((!sk[68]) & (!g1161) & (g1162) & (!g1174) & (g1187) & (!g1200)) + ((!sk[68]) & (!g1161) & (g1162) & (!g1174) & (g1187) & (g1200)) + ((!sk[68]) & (!g1161) & (g1162) & (g1174) & (!g1187) & (!g1200)) + ((!sk[68]) & (!g1161) & (g1162) & (g1174) & (!g1187) & (g1200)) + ((!sk[68]) & (!g1161) & (g1162) & (g1174) & (g1187) & (!g1200)) + ((!sk[68]) & (!g1161) & (g1162) & (g1174) & (g1187) & (g1200)) + ((!sk[68]) & (g1161) & (!g1162) & (!g1174) & (g1187) & (!g1200)) + ((!sk[68]) & (g1161) & (!g1162) & (!g1174) & (g1187) & (g1200)) + ((!sk[68]) & (g1161) & (!g1162) & (g1174) & (!g1187) & (!g1200)) + ((!sk[68]) & (g1161) & (!g1162) & (g1174) & (!g1187) & (g1200)) + ((!sk[68]) & (g1161) & (!g1162) & (g1174) & (g1187) & (!g1200)) + ((!sk[68]) & (g1161) & (!g1162) & (g1174) & (g1187) & (g1200)) + ((!sk[68]) & (g1161) & (g1162) & (!g1174) & (!g1187) & (!g1200)) + ((!sk[68]) & (g1161) & (g1162) & (!g1174) & (!g1187) & (g1200)) + ((!sk[68]) & (g1161) & (g1162) & (!g1174) & (g1187) & (!g1200)) + ((!sk[68]) & (g1161) & (g1162) & (!g1174) & (g1187) & (g1200)) + ((!sk[68]) & (g1161) & (g1162) & (g1174) & (!g1187) & (!g1200)) + ((!sk[68]) & (g1161) & (g1162) & (g1174) & (!g1187) & (g1200)) + ((!sk[68]) & (g1161) & (g1162) & (g1174) & (g1187) & (!g1200)) + ((!sk[68]) & (g1161) & (g1162) & (g1174) & (g1187) & (g1200)) + ((sk[68]) & (!g1161) & (!g1162) & (!g1174) & (g1187) & (!g1200)) + ((sk[68]) & (!g1161) & (!g1162) & (g1174) & (!g1187) & (!g1200)) + ((sk[68]) & (!g1161) & (!g1162) & (g1174) & (g1187) & (!g1200)) + ((sk[68]) & (!g1161) & (!g1162) & (g1174) & (g1187) & (g1200)) + ((sk[68]) & (!g1161) & (g1162) & (!g1174) & (!g1187) & (!g1200)) + ((sk[68]) & (!g1161) & (g1162) & (!g1174) & (g1187) & (!g1200)) + ((sk[68]) & (!g1161) & (g1162) & (!g1174) & (g1187) & (g1200)) + ((sk[68]) & (!g1161) & (g1162) & (g1174) & (!g1187) & (!g1200)) + ((sk[68]) & (!g1161) & (g1162) & (g1174) & (g1187) & (!g1200)) + ((sk[68]) & (!g1161) & (g1162) & (g1174) & (g1187) & (g1200)) + ((sk[68]) & (g1161) & (!g1162) & (!g1174) & (g1187) & (!g1200)) + ((sk[68]) & (g1161) & (!g1162) & (g1174) & (g1187) & (!g1200)) + ((sk[68]) & (g1161) & (g1162) & (!g1174) & (g1187) & (!g1200)) + ((sk[68]) & (g1161) & (g1162) & (g1174) & (!g1187) & (!g1200)) + ((sk[68]) & (g1161) & (g1162) & (g1174) & (g1187) & (!g1200)) + ((sk[68]) & (g1161) & (g1162) & (g1174) & (g1187) & (g1200)));
	assign g1211 = (((!g2) & (!g732) & (!g1188) & (!g1189) & (g1190) & (!g1199)) + ((!g2) & (!g732) & (!g1188) & (g1189) & (!g1190) & (!g1199)) + ((!g2) & (!g732) & (!g1188) & (g1189) & (g1190) & (!g1199)) + ((!g2) & (!g732) & (!g1188) & (g1189) & (g1190) & (g1199)) + ((!g2) & (!g732) & (g1188) & (!g1189) & (g1190) & (!g1199)) + ((!g2) & (!g732) & (g1188) & (g1189) & (!g1190) & (!g1199)) + ((!g2) & (!g732) & (g1188) & (g1189) & (g1190) & (!g1199)) + ((!g2) & (!g732) & (g1188) & (g1189) & (g1190) & (g1199)) + ((!g2) & (g732) & (!g1188) & (!g1189) & (g1190) & (!g1199)) + ((!g2) & (g732) & (!g1188) & (g1189) & (!g1190) & (!g1199)) + ((!g2) & (g732) & (!g1188) & (g1189) & (g1190) & (!g1199)) + ((!g2) & (g732) & (!g1188) & (g1189) & (g1190) & (g1199)) + ((!g2) & (g732) & (g1188) & (!g1189) & (!g1190) & (!g1199)) + ((!g2) & (g732) & (g1188) & (!g1189) & (g1190) & (!g1199)) + ((!g2) & (g732) & (g1188) & (!g1189) & (g1190) & (g1199)) + ((!g2) & (g732) & (g1188) & (g1189) & (!g1190) & (!g1199)) + ((!g2) & (g732) & (g1188) & (g1189) & (g1190) & (!g1199)) + ((!g2) & (g732) & (g1188) & (g1189) & (g1190) & (g1199)) + ((g2) & (!g732) & (!g1188) & (!g1189) & (!g1190) & (!g1199)) + ((g2) & (!g732) & (!g1188) & (!g1189) & (g1190) & (!g1199)) + ((g2) & (!g732) & (!g1188) & (!g1189) & (g1190) & (g1199)) + ((g2) & (!g732) & (!g1188) & (g1189) & (g1190) & (!g1199)) + ((g2) & (!g732) & (g1188) & (!g1189) & (!g1190) & (!g1199)) + ((g2) & (!g732) & (g1188) & (!g1189) & (g1190) & (!g1199)) + ((g2) & (!g732) & (g1188) & (!g1189) & (g1190) & (g1199)) + ((g2) & (!g732) & (g1188) & (g1189) & (g1190) & (!g1199)) + ((g2) & (g732) & (!g1188) & (!g1189) & (!g1190) & (!g1199)) + ((g2) & (g732) & (!g1188) & (!g1189) & (g1190) & (!g1199)) + ((g2) & (g732) & (!g1188) & (!g1189) & (g1190) & (g1199)) + ((g2) & (g732) & (!g1188) & (g1189) & (g1190) & (!g1199)) + ((g2) & (g732) & (g1188) & (!g1189) & (g1190) & (!g1199)) + ((g2) & (g732) & (g1188) & (g1189) & (g1190) & (!g1199)));
	assign g1212 = (((!g200) & (!g742) & (!g995) & (!g1191) & (!g1192) & (!g1198)) + ((!g200) & (!g742) & (!g995) & (!g1191) & (g1192) & (!g1198)) + ((!g200) & (!g742) & (!g995) & (!g1191) & (g1192) & (g1198)) + ((!g200) & (!g742) & (!g995) & (g1191) & (g1192) & (!g1198)) + ((!g200) & (!g742) & (g995) & (!g1191) & (!g1192) & (!g1198)) + ((!g200) & (!g742) & (g995) & (!g1191) & (g1192) & (!g1198)) + ((!g200) & (!g742) & (g995) & (!g1191) & (g1192) & (g1198)) + ((!g200) & (!g742) & (g995) & (g1191) & (g1192) & (!g1198)) + ((!g200) & (g742) & (!g995) & (!g1191) & (!g1192) & (!g1198)) + ((!g200) & (g742) & (!g995) & (!g1191) & (g1192) & (!g1198)) + ((!g200) & (g742) & (!g995) & (!g1191) & (g1192) & (g1198)) + ((!g200) & (g742) & (!g995) & (g1191) & (g1192) & (!g1198)) + ((!g200) & (g742) & (g995) & (!g1191) & (!g1192) & (!g1198)) + ((!g200) & (g742) & (g995) & (!g1191) & (g1192) & (!g1198)) + ((!g200) & (g742) & (g995) & (!g1191) & (g1192) & (g1198)) + ((!g200) & (g742) & (g995) & (g1191) & (!g1192) & (!g1198)) + ((!g200) & (g742) & (g995) & (g1191) & (g1192) & (!g1198)) + ((!g200) & (g742) & (g995) & (g1191) & (g1192) & (g1198)) + ((g200) & (!g742) & (!g995) & (!g1191) & (g1192) & (!g1198)) + ((g200) & (!g742) & (!g995) & (g1191) & (!g1192) & (!g1198)) + ((g200) & (!g742) & (!g995) & (g1191) & (g1192) & (!g1198)) + ((g200) & (!g742) & (!g995) & (g1191) & (g1192) & (g1198)) + ((g200) & (!g742) & (g995) & (!g1191) & (g1192) & (!g1198)) + ((g200) & (!g742) & (g995) & (g1191) & (!g1192) & (!g1198)) + ((g200) & (!g742) & (g995) & (g1191) & (g1192) & (!g1198)) + ((g200) & (!g742) & (g995) & (g1191) & (g1192) & (g1198)) + ((g200) & (g742) & (!g995) & (!g1191) & (g1192) & (!g1198)) + ((g200) & (g742) & (!g995) & (g1191) & (!g1192) & (!g1198)) + ((g200) & (g742) & (!g995) & (g1191) & (g1192) & (!g1198)) + ((g200) & (g742) & (!g995) & (g1191) & (g1192) & (g1198)) + ((g200) & (g742) & (g995) & (!g1191) & (g1192) & (!g1198)) + ((g200) & (g742) & (g995) & (g1191) & (g1192) & (!g1198)));
	assign g1213 = (((!g2) & (!g686) & (g732) & (!g1040) & (!g1079) & (!g1080)) + ((!g2) & (!g686) & (g732) & (!g1040) & (!g1079) & (g1080)) + ((!g2) & (!g686) & (g732) & (g1040) & (!g1079) & (g1080)) + ((!g2) & (g686) & (!g732) & (!g1040) & (!g1079) & (!g1080)) + ((!g2) & (g686) & (!g732) & (!g1040) & (!g1079) & (g1080)) + ((!g2) & (g686) & (!g732) & (g1040) & (!g1079) & (!g1080)) + ((!g2) & (g686) & (!g732) & (g1040) & (!g1079) & (g1080)) + ((!g2) & (g686) & (g732) & (!g1040) & (!g1079) & (!g1080)) + ((!g2) & (g686) & (g732) & (!g1040) & (!g1079) & (g1080)) + ((!g2) & (g686) & (g732) & (g1040) & (!g1079) & (!g1080)) + ((!g2) & (g686) & (g732) & (g1040) & (!g1079) & (g1080)) + ((g2) & (!g686) & (!g732) & (!g1040) & (!g1079) & (!g1080)) + ((g2) & (!g686) & (!g732) & (!g1040) & (!g1079) & (g1080)) + ((g2) & (!g686) & (!g732) & (!g1040) & (g1079) & (!g1080)) + ((g2) & (!g686) & (!g732) & (!g1040) & (g1079) & (g1080)) + ((g2) & (!g686) & (!g732) & (g1040) & (!g1079) & (!g1080)) + ((g2) & (!g686) & (!g732) & (g1040) & (!g1079) & (g1080)) + ((g2) & (!g686) & (!g732) & (g1040) & (g1079) & (!g1080)) + ((g2) & (!g686) & (!g732) & (g1040) & (g1079) & (g1080)) + ((g2) & (!g686) & (g732) & (!g1040) & (g1079) & (!g1080)) + ((g2) & (!g686) & (g732) & (!g1040) & (g1079) & (g1080)) + ((g2) & (!g686) & (g732) & (g1040) & (!g1079) & (!g1080)) + ((g2) & (!g686) & (g732) & (g1040) & (g1079) & (!g1080)) + ((g2) & (!g686) & (g732) & (g1040) & (g1079) & (g1080)) + ((g2) & (g686) & (!g732) & (!g1040) & (g1079) & (!g1080)) + ((g2) & (g686) & (!g732) & (!g1040) & (g1079) & (g1080)) + ((g2) & (g686) & (!g732) & (g1040) & (g1079) & (!g1080)) + ((g2) & (g686) & (!g732) & (g1040) & (g1079) & (g1080)) + ((g2) & (g686) & (g732) & (!g1040) & (g1079) & (!g1080)) + ((g2) & (g686) & (g732) & (!g1040) & (g1079) & (g1080)) + ((g2) & (g686) & (g732) & (g1040) & (g1079) & (!g1080)) + ((g2) & (g686) & (g732) & (g1040) & (g1079) & (g1080)));
	assign g1214 = (((!g747) & (!g744) & (!sk[72]) & (!g994) & (g1040)) + ((!g747) & (!g744) & (!sk[72]) & (g994) & (g1040)) + ((!g747) & (g744) & (!sk[72]) & (!g994) & (g1040)) + ((!g747) & (g744) & (!sk[72]) & (g994) & (g1040)) + ((!g747) & (g744) & (sk[72]) & (g994) & (!g1040)) + ((!g747) & (g744) & (sk[72]) & (g994) & (g1040)) + ((g747) & (!g744) & (!sk[72]) & (!g994) & (!g1040)) + ((g747) & (!g744) & (!sk[72]) & (!g994) & (g1040)) + ((g747) & (!g744) & (!sk[72]) & (g994) & (!g1040)) + ((g747) & (!g744) & (!sk[72]) & (g994) & (g1040)) + ((g747) & (!g744) & (sk[72]) & (!g994) & (!g1040)) + ((g747) & (!g744) & (sk[72]) & (g994) & (!g1040)) + ((g747) & (g744) & (!sk[72]) & (!g994) & (!g1040)) + ((g747) & (g744) & (!sk[72]) & (!g994) & (g1040)) + ((g747) & (g744) & (!sk[72]) & (g994) & (!g1040)) + ((g747) & (g744) & (!sk[72]) & (g994) & (g1040)) + ((g747) & (g744) & (sk[72]) & (!g994) & (!g1040)) + ((g747) & (g744) & (sk[72]) & (g994) & (!g1040)) + ((g747) & (g744) & (sk[72]) & (g994) & (g1040)));
	assign g1215 = (((!g200) & (!g742) & (!g748) & (!g971) & (!g1041) & (g1214)) + ((!g200) & (!g742) & (!g748) & (!g971) & (g1041) & (g1214)) + ((!g200) & (!g742) & (!g748) & (g971) & (!g1041) & (g1214)) + ((!g200) & (!g742) & (!g748) & (g971) & (g1041) & (g1214)) + ((!g200) & (!g742) & (g748) & (!g971) & (!g1041) & (g1214)) + ((!g200) & (!g742) & (g748) & (!g971) & (g1041) & (g1214)) + ((!g200) & (!g742) & (g748) & (g971) & (!g1041) & (!g1214)) + ((!g200) & (!g742) & (g748) & (g971) & (!g1041) & (g1214)) + ((!g200) & (!g742) & (g748) & (g971) & (g1041) & (!g1214)) + ((!g200) & (!g742) & (g748) & (g971) & (g1041) & (g1214)) + ((!g200) & (g742) & (!g748) & (!g971) & (!g1041) & (!g1214)) + ((!g200) & (g742) & (!g748) & (!g971) & (!g1041) & (g1214)) + ((!g200) & (g742) & (!g748) & (!g971) & (g1041) & (g1214)) + ((!g200) & (g742) & (!g748) & (g971) & (!g1041) & (!g1214)) + ((!g200) & (g742) & (!g748) & (g971) & (!g1041) & (g1214)) + ((!g200) & (g742) & (!g748) & (g971) & (g1041) & (g1214)) + ((!g200) & (g742) & (g748) & (!g971) & (!g1041) & (!g1214)) + ((!g200) & (g742) & (g748) & (!g971) & (!g1041) & (g1214)) + ((!g200) & (g742) & (g748) & (!g971) & (g1041) & (g1214)) + ((!g200) & (g742) & (g748) & (g971) & (!g1041) & (!g1214)) + ((!g200) & (g742) & (g748) & (g971) & (!g1041) & (g1214)) + ((!g200) & (g742) & (g748) & (g971) & (g1041) & (!g1214)) + ((!g200) & (g742) & (g748) & (g971) & (g1041) & (g1214)) + ((g200) & (!g742) & (!g748) & (!g971) & (!g1041) & (!g1214)) + ((g200) & (!g742) & (!g748) & (!g971) & (g1041) & (!g1214)) + ((g200) & (!g742) & (!g748) & (g971) & (!g1041) & (!g1214)) + ((g200) & (!g742) & (!g748) & (g971) & (g1041) & (!g1214)) + ((g200) & (!g742) & (g748) & (!g971) & (!g1041) & (!g1214)) + ((g200) & (!g742) & (g748) & (!g971) & (g1041) & (!g1214)) + ((g200) & (g742) & (!g748) & (!g971) & (g1041) & (!g1214)) + ((g200) & (g742) & (!g748) & (g971) & (g1041) & (!g1214)) + ((g200) & (g742) & (g748) & (!g971) & (g1041) & (!g1214)));
	assign g1216 = (((!g202) & (!g759) & (!g895) & (!g1194) & (!g1196) & (!g1197)) + ((!g202) & (!g759) & (!g895) & (!g1194) & (!g1196) & (g1197)) + ((!g202) & (!g759) & (!g895) & (!g1194) & (g1196) & (g1197)) + ((!g202) & (!g759) & (!g895) & (g1194) & (!g1196) & (g1197)) + ((!g202) & (!g759) & (g895) & (!g1194) & (!g1196) & (!g1197)) + ((!g202) & (!g759) & (g895) & (!g1194) & (!g1196) & (g1197)) + ((!g202) & (!g759) & (g895) & (!g1194) & (g1196) & (g1197)) + ((!g202) & (!g759) & (g895) & (g1194) & (!g1196) & (g1197)) + ((!g202) & (g759) & (!g895) & (!g1194) & (!g1196) & (!g1197)) + ((!g202) & (g759) & (!g895) & (!g1194) & (!g1196) & (g1197)) + ((!g202) & (g759) & (!g895) & (!g1194) & (g1196) & (g1197)) + ((!g202) & (g759) & (!g895) & (g1194) & (!g1196) & (g1197)) + ((!g202) & (g759) & (g895) & (!g1194) & (!g1196) & (!g1197)) + ((!g202) & (g759) & (g895) & (!g1194) & (!g1196) & (g1197)) + ((!g202) & (g759) & (g895) & (!g1194) & (g1196) & (g1197)) + ((!g202) & (g759) & (g895) & (g1194) & (!g1196) & (!g1197)) + ((!g202) & (g759) & (g895) & (g1194) & (!g1196) & (g1197)) + ((!g202) & (g759) & (g895) & (g1194) & (g1196) & (g1197)) + ((g202) & (!g759) & (!g895) & (!g1194) & (!g1196) & (g1197)) + ((g202) & (!g759) & (!g895) & (g1194) & (!g1196) & (!g1197)) + ((g202) & (!g759) & (!g895) & (g1194) & (!g1196) & (g1197)) + ((g202) & (!g759) & (!g895) & (g1194) & (g1196) & (g1197)) + ((g202) & (!g759) & (g895) & (!g1194) & (!g1196) & (g1197)) + ((g202) & (!g759) & (g895) & (g1194) & (!g1196) & (!g1197)) + ((g202) & (!g759) & (g895) & (g1194) & (!g1196) & (g1197)) + ((g202) & (!g759) & (g895) & (g1194) & (g1196) & (g1197)) + ((g202) & (g759) & (!g895) & (!g1194) & (!g1196) & (g1197)) + ((g202) & (g759) & (!g895) & (g1194) & (!g1196) & (!g1197)) + ((g202) & (g759) & (!g895) & (g1194) & (!g1196) & (g1197)) + ((g202) & (g759) & (!g895) & (g1194) & (g1196) & (g1197)) + ((g202) & (g759) & (g895) & (!g1194) & (!g1196) & (g1197)) + ((g202) & (g759) & (g895) & (g1194) & (!g1196) & (g1197)));
	assign g1217 = (((!g884) & (sk[75]) & (g890)) + ((g884) & (!sk[75]) & (g890)) + ((g884) & (sk[75]) & (!g890)));
	assign g1218 = (((!g764) & (!g762) & (!g765) & (!g962) & (!g863) & (!g963)) + ((!g764) & (!g762) & (!g765) & (!g962) & (!g863) & (g963)) + ((!g764) & (!g762) & (!g765) & (!g962) & (g863) & (!g963)) + ((!g764) & (!g762) & (!g765) & (!g962) & (g863) & (g963)) + ((!g764) & (!g762) & (!g765) & (g962) & (!g863) & (!g963)) + ((!g764) & (!g762) & (!g765) & (g962) & (!g863) & (g963)) + ((!g764) & (!g762) & (!g765) & (g962) & (g863) & (!g963)) + ((!g764) & (!g762) & (!g765) & (g962) & (g863) & (g963)) + ((!g764) & (!g762) & (g765) & (!g962) & (!g863) & (!g963)) + ((!g764) & (!g762) & (g765) & (!g962) & (!g863) & (g963)) + ((!g764) & (!g762) & (g765) & (g962) & (!g863) & (!g963)) + ((!g764) & (!g762) & (g765) & (g962) & (!g863) & (g963)) + ((!g764) & (g762) & (!g765) & (!g962) & (!g863) & (!g963)) + ((!g764) & (g762) & (!g765) & (!g962) & (g863) & (!g963)) + ((!g764) & (g762) & (!g765) & (g962) & (!g863) & (!g963)) + ((!g764) & (g762) & (!g765) & (g962) & (g863) & (!g963)) + ((!g764) & (g762) & (g765) & (!g962) & (!g863) & (!g963)) + ((!g764) & (g762) & (g765) & (g962) & (!g863) & (!g963)) + ((g764) & (!g762) & (!g765) & (g962) & (!g863) & (!g963)) + ((g764) & (!g762) & (!g765) & (g962) & (!g863) & (g963)) + ((g764) & (!g762) & (!g765) & (g962) & (g863) & (!g963)) + ((g764) & (!g762) & (!g765) & (g962) & (g863) & (g963)) + ((g764) & (!g762) & (g765) & (g962) & (!g863) & (!g963)) + ((g764) & (!g762) & (g765) & (g962) & (!g863) & (g963)) + ((g764) & (g762) & (!g765) & (g962) & (!g863) & (!g963)) + ((g764) & (g762) & (!g765) & (g962) & (g863) & (!g963)) + ((g764) & (g762) & (g765) & (g962) & (!g863) & (!g963)));
	assign g1219 = (((!sk[77]) & (!g843) & (g834) & (!g835)) + ((!sk[77]) & (!g843) & (g834) & (g835)) + ((!sk[77]) & (g843) & (g834) & (!g835)) + ((!sk[77]) & (g843) & (g834) & (g835)) + ((sk[77]) & (g843) & (!g834) & (!g835)) + ((sk[77]) & (g843) & (g834) & (g835)));
	assign g1220 = (((!g869) & (!g718) & (!g847) & (!g845) & (!g870) & (!g848)) + ((!g869) & (!g718) & (!g847) & (!g845) & (!g870) & (g848)) + ((!g869) & (!g718) & (!g847) & (!g845) & (g870) & (!g848)) + ((!g869) & (!g718) & (!g847) & (!g845) & (g870) & (g848)) + ((!g869) & (!g718) & (!g847) & (g845) & (!g870) & (!g848)) + ((!g869) & (!g718) & (!g847) & (g845) & (!g870) & (g848)) + ((!g869) & (!g718) & (!g847) & (g845) & (g870) & (!g848)) + ((!g869) & (!g718) & (!g847) & (g845) & (g870) & (g848)) + ((!g869) & (!g718) & (g847) & (!g845) & (g870) & (!g848)) + ((!g869) & (!g718) & (g847) & (!g845) & (g870) & (g848)) + ((!g869) & (!g718) & (g847) & (g845) & (g870) & (!g848)) + ((!g869) & (!g718) & (g847) & (g845) & (g870) & (g848)) + ((!g869) & (g718) & (!g847) & (!g845) & (!g870) & (!g848)) + ((!g869) & (g718) & (!g847) & (!g845) & (g870) & (!g848)) + ((!g869) & (g718) & (!g847) & (g845) & (!g870) & (!g848)) + ((!g869) & (g718) & (!g847) & (g845) & (g870) & (!g848)) + ((!g869) & (g718) & (g847) & (!g845) & (g870) & (!g848)) + ((!g869) & (g718) & (g847) & (g845) & (g870) & (!g848)) + ((g869) & (!g718) & (!g847) & (!g845) & (!g870) & (!g848)) + ((g869) & (!g718) & (!g847) & (!g845) & (!g870) & (g848)) + ((g869) & (!g718) & (!g847) & (!g845) & (g870) & (!g848)) + ((g869) & (!g718) & (!g847) & (!g845) & (g870) & (g848)) + ((g869) & (!g718) & (g847) & (!g845) & (g870) & (!g848)) + ((g869) & (!g718) & (g847) & (!g845) & (g870) & (g848)) + ((g869) & (g718) & (!g847) & (!g845) & (!g870) & (!g848)) + ((g869) & (g718) & (!g847) & (!g845) & (g870) & (!g848)) + ((g869) & (g718) & (g847) & (!g845) & (g870) & (!g848)));
	assign g1221 = (((!g252) & (!g683) & (!sk[79]) & (!g719) & (g729) & (!g1168)) + ((!g252) & (!g683) & (!sk[79]) & (!g719) & (g729) & (g1168)) + ((!g252) & (!g683) & (!sk[79]) & (g719) & (!g729) & (!g1168)) + ((!g252) & (!g683) & (!sk[79]) & (g719) & (!g729) & (g1168)) + ((!g252) & (!g683) & (!sk[79]) & (g719) & (g729) & (!g1168)) + ((!g252) & (!g683) & (!sk[79]) & (g719) & (g729) & (g1168)) + ((!g252) & (g683) & (!sk[79]) & (!g719) & (!g729) & (!g1168)) + ((!g252) & (g683) & (!sk[79]) & (!g719) & (!g729) & (g1168)) + ((!g252) & (g683) & (!sk[79]) & (!g719) & (g729) & (!g1168)) + ((!g252) & (g683) & (!sk[79]) & (!g719) & (g729) & (g1168)) + ((!g252) & (g683) & (!sk[79]) & (g719) & (!g729) & (!g1168)) + ((!g252) & (g683) & (!sk[79]) & (g719) & (!g729) & (g1168)) + ((!g252) & (g683) & (!sk[79]) & (g719) & (g729) & (!g1168)) + ((!g252) & (g683) & (!sk[79]) & (g719) & (g729) & (g1168)) + ((!g252) & (g683) & (sk[79]) & (!g719) & (!g729) & (!g1168)) + ((!g252) & (g683) & (sk[79]) & (!g719) & (g729) & (!g1168)) + ((!g252) & (g683) & (sk[79]) & (g719) & (!g729) & (!g1168)) + ((!g252) & (g683) & (sk[79]) & (g719) & (g729) & (!g1168)) + ((g252) & (!g683) & (!sk[79]) & (!g719) & (g729) & (!g1168)) + ((g252) & (!g683) & (!sk[79]) & (!g719) & (g729) & (g1168)) + ((g252) & (!g683) & (!sk[79]) & (g719) & (!g729) & (!g1168)) + ((g252) & (!g683) & (!sk[79]) & (g719) & (!g729) & (g1168)) + ((g252) & (!g683) & (!sk[79]) & (g719) & (g729) & (!g1168)) + ((g252) & (!g683) & (!sk[79]) & (g719) & (g729) & (g1168)) + ((g252) & (!g683) & (sk[79]) & (!g719) & (!g729) & (g1168)) + ((g252) & (g683) & (!sk[79]) & (!g719) & (!g729) & (!g1168)) + ((g252) & (g683) & (!sk[79]) & (!g719) & (!g729) & (g1168)) + ((g252) & (g683) & (!sk[79]) & (!g719) & (g729) & (!g1168)) + ((g252) & (g683) & (!sk[79]) & (!g719) & (g729) & (g1168)) + ((g252) & (g683) & (!sk[79]) & (g719) & (!g729) & (!g1168)) + ((g252) & (g683) & (!sk[79]) & (g719) & (!g729) & (g1168)) + ((g252) & (g683) & (!sk[79]) & (g719) & (g729) & (!g1168)) + ((g252) & (g683) & (!sk[79]) & (g719) & (g729) & (g1168)) + ((g252) & (g683) & (sk[79]) & (!g719) & (!g729) & (!g1168)) + ((g252) & (g683) & (sk[79]) & (!g719) & (!g729) & (g1168)) + ((g252) & (g683) & (sk[79]) & (!g719) & (g729) & (!g1168)) + ((g252) & (g683) & (sk[79]) & (!g719) & (g729) & (g1168)) + ((g252) & (g683) & (sk[79]) & (g719) & (!g729) & (!g1168)) + ((g252) & (g683) & (sk[79]) & (g719) & (!g729) & (g1168)) + ((g252) & (g683) & (sk[79]) & (g719) & (g729) & (g1168)));
	assign g1222 = (((!g252) & (!g683) & (!g681) & (!g1219) & (!g1220) & (g1221)) + ((!g252) & (!g683) & (!g681) & (!g1219) & (g1220) & (!g1221)) + ((!g252) & (!g683) & (!g681) & (g1219) & (!g1220) & (g1221)) + ((!g252) & (!g683) & (!g681) & (g1219) & (g1220) & (g1221)) + ((!g252) & (!g683) & (g681) & (!g1219) & (!g1220) & (g1221)) + ((!g252) & (!g683) & (g681) & (!g1219) & (g1220) & (!g1221)) + ((!g252) & (!g683) & (g681) & (g1219) & (!g1220) & (g1221)) + ((!g252) & (!g683) & (g681) & (g1219) & (g1220) & (g1221)) + ((!g252) & (g683) & (!g681) & (!g1219) & (!g1220) & (!g1221)) + ((!g252) & (g683) & (!g681) & (!g1219) & (g1220) & (g1221)) + ((!g252) & (g683) & (!g681) & (g1219) & (!g1220) & (!g1221)) + ((!g252) & (g683) & (!g681) & (g1219) & (g1220) & (!g1221)) + ((!g252) & (g683) & (g681) & (!g1219) & (!g1220) & (!g1221)) + ((!g252) & (g683) & (g681) & (!g1219) & (g1220) & (g1221)) + ((!g252) & (g683) & (g681) & (g1219) & (!g1220) & (!g1221)) + ((!g252) & (g683) & (g681) & (g1219) & (g1220) & (!g1221)) + ((g252) & (!g683) & (!g681) & (!g1219) & (!g1220) & (g1221)) + ((g252) & (!g683) & (!g681) & (!g1219) & (g1220) & (!g1221)) + ((g252) & (!g683) & (!g681) & (g1219) & (!g1220) & (g1221)) + ((g252) & (!g683) & (!g681) & (g1219) & (g1220) & (g1221)) + ((g252) & (!g683) & (g681) & (!g1219) & (!g1220) & (!g1221)) + ((g252) & (!g683) & (g681) & (!g1219) & (g1220) & (g1221)) + ((g252) & (!g683) & (g681) & (g1219) & (!g1220) & (!g1221)) + ((g252) & (!g683) & (g681) & (g1219) & (g1220) & (!g1221)) + ((g252) & (g683) & (!g681) & (!g1219) & (!g1220) & (!g1221)) + ((g252) & (g683) & (!g681) & (!g1219) & (g1220) & (g1221)) + ((g252) & (g683) & (!g681) & (g1219) & (!g1220) & (!g1221)) + ((g252) & (g683) & (!g681) & (g1219) & (g1220) & (!g1221)) + ((g252) & (g683) & (g681) & (!g1219) & (!g1220) & (g1221)) + ((g252) & (g683) & (g681) & (!g1219) & (g1220) & (!g1221)) + ((g252) & (g683) & (g681) & (g1219) & (!g1220) & (g1221)) + ((g252) & (g683) & (g681) & (g1219) & (g1220) & (g1221)));
	assign g1223 = (((!g202) & (!g759) & (!g1217) & (!sk[81]) & (g1218) & (!g1222)) + ((!g202) & (!g759) & (!g1217) & (!sk[81]) & (g1218) & (g1222)) + ((!g202) & (!g759) & (!g1217) & (sk[81]) & (!g1218) & (!g1222)) + ((!g202) & (!g759) & (!g1217) & (sk[81]) & (g1218) & (g1222)) + ((!g202) & (!g759) & (g1217) & (!sk[81]) & (!g1218) & (!g1222)) + ((!g202) & (!g759) & (g1217) & (!sk[81]) & (!g1218) & (g1222)) + ((!g202) & (!g759) & (g1217) & (!sk[81]) & (g1218) & (!g1222)) + ((!g202) & (!g759) & (g1217) & (!sk[81]) & (g1218) & (g1222)) + ((!g202) & (!g759) & (g1217) & (sk[81]) & (!g1218) & (!g1222)) + ((!g202) & (!g759) & (g1217) & (sk[81]) & (g1218) & (g1222)) + ((!g202) & (g759) & (!g1217) & (!sk[81]) & (!g1218) & (!g1222)) + ((!g202) & (g759) & (!g1217) & (!sk[81]) & (!g1218) & (g1222)) + ((!g202) & (g759) & (!g1217) & (!sk[81]) & (g1218) & (!g1222)) + ((!g202) & (g759) & (!g1217) & (!sk[81]) & (g1218) & (g1222)) + ((!g202) & (g759) & (!g1217) & (sk[81]) & (!g1218) & (!g1222)) + ((!g202) & (g759) & (!g1217) & (sk[81]) & (g1218) & (!g1222)) + ((!g202) & (g759) & (g1217) & (!sk[81]) & (!g1218) & (!g1222)) + ((!g202) & (g759) & (g1217) & (!sk[81]) & (!g1218) & (g1222)) + ((!g202) & (g759) & (g1217) & (!sk[81]) & (g1218) & (!g1222)) + ((!g202) & (g759) & (g1217) & (!sk[81]) & (g1218) & (g1222)) + ((!g202) & (g759) & (g1217) & (sk[81]) & (!g1218) & (!g1222)) + ((!g202) & (g759) & (g1217) & (sk[81]) & (g1218) & (g1222)) + ((g202) & (!g759) & (!g1217) & (!sk[81]) & (g1218) & (!g1222)) + ((g202) & (!g759) & (!g1217) & (!sk[81]) & (g1218) & (g1222)) + ((g202) & (!g759) & (!g1217) & (sk[81]) & (!g1218) & (g1222)) + ((g202) & (!g759) & (!g1217) & (sk[81]) & (g1218) & (!g1222)) + ((g202) & (!g759) & (g1217) & (!sk[81]) & (!g1218) & (!g1222)) + ((g202) & (!g759) & (g1217) & (!sk[81]) & (!g1218) & (g1222)) + ((g202) & (!g759) & (g1217) & (!sk[81]) & (g1218) & (!g1222)) + ((g202) & (!g759) & (g1217) & (!sk[81]) & (g1218) & (g1222)) + ((g202) & (!g759) & (g1217) & (sk[81]) & (!g1218) & (g1222)) + ((g202) & (!g759) & (g1217) & (sk[81]) & (g1218) & (!g1222)) + ((g202) & (g759) & (!g1217) & (!sk[81]) & (!g1218) & (!g1222)) + ((g202) & (g759) & (!g1217) & (!sk[81]) & (!g1218) & (g1222)) + ((g202) & (g759) & (!g1217) & (!sk[81]) & (g1218) & (!g1222)) + ((g202) & (g759) & (!g1217) & (!sk[81]) & (g1218) & (g1222)) + ((g202) & (g759) & (!g1217) & (sk[81]) & (!g1218) & (g1222)) + ((g202) & (g759) & (!g1217) & (sk[81]) & (g1218) & (g1222)) + ((g202) & (g759) & (g1217) & (!sk[81]) & (!g1218) & (!g1222)) + ((g202) & (g759) & (g1217) & (!sk[81]) & (!g1218) & (g1222)) + ((g202) & (g759) & (g1217) & (!sk[81]) & (g1218) & (!g1222)) + ((g202) & (g759) & (g1217) & (!sk[81]) & (g1218) & (g1222)) + ((g202) & (g759) & (g1217) & (sk[81]) & (!g1218) & (g1222)) + ((g202) & (g759) & (g1217) & (sk[81]) & (g1218) & (!g1222)));
	assign g1224 = (((!g1212) & (!g1213) & (!g1215) & (!sk[82]) & (g1216) & (!g1223)) + ((!g1212) & (!g1213) & (!g1215) & (!sk[82]) & (g1216) & (g1223)) + ((!g1212) & (!g1213) & (!g1215) & (sk[82]) & (!g1216) & (g1223)) + ((!g1212) & (!g1213) & (!g1215) & (sk[82]) & (g1216) & (!g1223)) + ((!g1212) & (!g1213) & (g1215) & (!sk[82]) & (!g1216) & (!g1223)) + ((!g1212) & (!g1213) & (g1215) & (!sk[82]) & (!g1216) & (g1223)) + ((!g1212) & (!g1213) & (g1215) & (!sk[82]) & (g1216) & (!g1223)) + ((!g1212) & (!g1213) & (g1215) & (!sk[82]) & (g1216) & (g1223)) + ((!g1212) & (!g1213) & (g1215) & (sk[82]) & (!g1216) & (!g1223)) + ((!g1212) & (!g1213) & (g1215) & (sk[82]) & (g1216) & (g1223)) + ((!g1212) & (g1213) & (!g1215) & (!sk[82]) & (!g1216) & (!g1223)) + ((!g1212) & (g1213) & (!g1215) & (!sk[82]) & (!g1216) & (g1223)) + ((!g1212) & (g1213) & (!g1215) & (!sk[82]) & (g1216) & (!g1223)) + ((!g1212) & (g1213) & (!g1215) & (!sk[82]) & (g1216) & (g1223)) + ((!g1212) & (g1213) & (!g1215) & (sk[82]) & (!g1216) & (!g1223)) + ((!g1212) & (g1213) & (!g1215) & (sk[82]) & (g1216) & (g1223)) + ((!g1212) & (g1213) & (g1215) & (!sk[82]) & (!g1216) & (!g1223)) + ((!g1212) & (g1213) & (g1215) & (!sk[82]) & (!g1216) & (g1223)) + ((!g1212) & (g1213) & (g1215) & (!sk[82]) & (g1216) & (!g1223)) + ((!g1212) & (g1213) & (g1215) & (!sk[82]) & (g1216) & (g1223)) + ((!g1212) & (g1213) & (g1215) & (sk[82]) & (!g1216) & (g1223)) + ((!g1212) & (g1213) & (g1215) & (sk[82]) & (g1216) & (!g1223)) + ((g1212) & (!g1213) & (!g1215) & (!sk[82]) & (g1216) & (!g1223)) + ((g1212) & (!g1213) & (!g1215) & (!sk[82]) & (g1216) & (g1223)) + ((g1212) & (!g1213) & (!g1215) & (sk[82]) & (!g1216) & (!g1223)) + ((g1212) & (!g1213) & (!g1215) & (sk[82]) & (g1216) & (g1223)) + ((g1212) & (!g1213) & (g1215) & (!sk[82]) & (!g1216) & (!g1223)) + ((g1212) & (!g1213) & (g1215) & (!sk[82]) & (!g1216) & (g1223)) + ((g1212) & (!g1213) & (g1215) & (!sk[82]) & (g1216) & (!g1223)) + ((g1212) & (!g1213) & (g1215) & (!sk[82]) & (g1216) & (g1223)) + ((g1212) & (!g1213) & (g1215) & (sk[82]) & (!g1216) & (g1223)) + ((g1212) & (!g1213) & (g1215) & (sk[82]) & (g1216) & (!g1223)) + ((g1212) & (g1213) & (!g1215) & (!sk[82]) & (!g1216) & (!g1223)) + ((g1212) & (g1213) & (!g1215) & (!sk[82]) & (!g1216) & (g1223)) + ((g1212) & (g1213) & (!g1215) & (!sk[82]) & (g1216) & (!g1223)) + ((g1212) & (g1213) & (!g1215) & (!sk[82]) & (g1216) & (g1223)) + ((g1212) & (g1213) & (!g1215) & (sk[82]) & (!g1216) & (g1223)) + ((g1212) & (g1213) & (!g1215) & (sk[82]) & (g1216) & (!g1223)) + ((g1212) & (g1213) & (g1215) & (!sk[82]) & (!g1216) & (!g1223)) + ((g1212) & (g1213) & (g1215) & (!sk[82]) & (!g1216) & (g1223)) + ((g1212) & (g1213) & (g1215) & (!sk[82]) & (g1216) & (!g1223)) + ((g1212) & (g1213) & (g1215) & (!sk[82]) & (g1216) & (g1223)) + ((g1212) & (g1213) & (g1215) & (sk[82]) & (!g1216) & (!g1223)) + ((g1212) & (g1213) & (g1215) & (sk[82]) & (g1216) & (g1223)));
	assign g1225 = (((!sk[83]) & (g1211) & (g1224)) + ((sk[83]) & (!g1211) & (g1224)) + ((sk[83]) & (g1211) & (!g1224)));
	assign g1226 = (((!g38) & (!g79) & (!g71) & (!g20) & (!g661) & (!g587)) + ((!g38) & (!g79) & (!g71) & (g20) & (!g661) & (!g587)) + ((!g38) & (!g79) & (g71) & (!g20) & (!g661) & (!g587)) + ((g38) & (!g79) & (!g71) & (!g20) & (!g661) & (!g587)) + ((g38) & (!g79) & (!g71) & (g20) & (!g661) & (!g587)));
	assign g1227 = (((!g563) & (!g643) & (!sk[85]) & (!g666) & (g1071) & (!g1226)) + ((!g563) & (!g643) & (!sk[85]) & (!g666) & (g1071) & (g1226)) + ((!g563) & (!g643) & (!sk[85]) & (g666) & (!g1071) & (!g1226)) + ((!g563) & (!g643) & (!sk[85]) & (g666) & (!g1071) & (g1226)) + ((!g563) & (!g643) & (!sk[85]) & (g666) & (g1071) & (!g1226)) + ((!g563) & (!g643) & (!sk[85]) & (g666) & (g1071) & (g1226)) + ((!g563) & (g643) & (!sk[85]) & (!g666) & (!g1071) & (!g1226)) + ((!g563) & (g643) & (!sk[85]) & (!g666) & (!g1071) & (g1226)) + ((!g563) & (g643) & (!sk[85]) & (!g666) & (g1071) & (!g1226)) + ((!g563) & (g643) & (!sk[85]) & (!g666) & (g1071) & (g1226)) + ((!g563) & (g643) & (!sk[85]) & (g666) & (!g1071) & (!g1226)) + ((!g563) & (g643) & (!sk[85]) & (g666) & (!g1071) & (g1226)) + ((!g563) & (g643) & (!sk[85]) & (g666) & (g1071) & (!g1226)) + ((!g563) & (g643) & (!sk[85]) & (g666) & (g1071) & (g1226)) + ((!g563) & (g643) & (sk[85]) & (g666) & (g1071) & (g1226)) + ((g563) & (!g643) & (!sk[85]) & (!g666) & (g1071) & (!g1226)) + ((g563) & (!g643) & (!sk[85]) & (!g666) & (g1071) & (g1226)) + ((g563) & (!g643) & (!sk[85]) & (g666) & (!g1071) & (!g1226)) + ((g563) & (!g643) & (!sk[85]) & (g666) & (!g1071) & (g1226)) + ((g563) & (!g643) & (!sk[85]) & (g666) & (g1071) & (!g1226)) + ((g563) & (!g643) & (!sk[85]) & (g666) & (g1071) & (g1226)) + ((g563) & (g643) & (!sk[85]) & (!g666) & (!g1071) & (!g1226)) + ((g563) & (g643) & (!sk[85]) & (!g666) & (!g1071) & (g1226)) + ((g563) & (g643) & (!sk[85]) & (!g666) & (g1071) & (!g1226)) + ((g563) & (g643) & (!sk[85]) & (!g666) & (g1071) & (g1226)) + ((g563) & (g643) & (!sk[85]) & (g666) & (!g1071) & (!g1226)) + ((g563) & (g643) & (!sk[85]) & (g666) & (!g1071) & (g1226)) + ((g563) & (g643) & (!sk[85]) & (g666) & (g1071) & (!g1226)) + ((g563) & (g643) & (!sk[85]) & (g666) & (g1071) & (g1226)));
	assign g1228 = (((!g78) & (!g90) & (!sk[86]) & (!g55) & (g142) & (!g967)) + ((!g78) & (!g90) & (!sk[86]) & (!g55) & (g142) & (g967)) + ((!g78) & (!g90) & (!sk[86]) & (g55) & (!g142) & (!g967)) + ((!g78) & (!g90) & (!sk[86]) & (g55) & (!g142) & (g967)) + ((!g78) & (!g90) & (!sk[86]) & (g55) & (g142) & (!g967)) + ((!g78) & (!g90) & (!sk[86]) & (g55) & (g142) & (g967)) + ((!g78) & (!g90) & (sk[86]) & (!g55) & (!g142) & (!g967)) + ((!g78) & (g90) & (!sk[86]) & (!g55) & (!g142) & (!g967)) + ((!g78) & (g90) & (!sk[86]) & (!g55) & (!g142) & (g967)) + ((!g78) & (g90) & (!sk[86]) & (!g55) & (g142) & (!g967)) + ((!g78) & (g90) & (!sk[86]) & (!g55) & (g142) & (g967)) + ((!g78) & (g90) & (!sk[86]) & (g55) & (!g142) & (!g967)) + ((!g78) & (g90) & (!sk[86]) & (g55) & (!g142) & (g967)) + ((!g78) & (g90) & (!sk[86]) & (g55) & (g142) & (!g967)) + ((!g78) & (g90) & (!sk[86]) & (g55) & (g142) & (g967)) + ((g78) & (!g90) & (!sk[86]) & (!g55) & (g142) & (!g967)) + ((g78) & (!g90) & (!sk[86]) & (!g55) & (g142) & (g967)) + ((g78) & (!g90) & (!sk[86]) & (g55) & (!g142) & (!g967)) + ((g78) & (!g90) & (!sk[86]) & (g55) & (!g142) & (g967)) + ((g78) & (!g90) & (!sk[86]) & (g55) & (g142) & (!g967)) + ((g78) & (!g90) & (!sk[86]) & (g55) & (g142) & (g967)) + ((g78) & (g90) & (!sk[86]) & (!g55) & (!g142) & (!g967)) + ((g78) & (g90) & (!sk[86]) & (!g55) & (!g142) & (g967)) + ((g78) & (g90) & (!sk[86]) & (!g55) & (g142) & (!g967)) + ((g78) & (g90) & (!sk[86]) & (!g55) & (g142) & (g967)) + ((g78) & (g90) & (!sk[86]) & (g55) & (!g142) & (!g967)) + ((g78) & (g90) & (!sk[86]) & (g55) & (!g142) & (g967)) + ((g78) & (g90) & (!sk[86]) & (g55) & (g142) & (!g967)) + ((g78) & (g90) & (!sk[86]) & (g55) & (g142) & (g967)));
	assign g1229 = (((!g664) & (!g1005) & (!sk[87]) & (!g1178) & (g1227) & (!g1228)) + ((!g664) & (!g1005) & (!sk[87]) & (!g1178) & (g1227) & (g1228)) + ((!g664) & (!g1005) & (!sk[87]) & (g1178) & (!g1227) & (!g1228)) + ((!g664) & (!g1005) & (!sk[87]) & (g1178) & (!g1227) & (g1228)) + ((!g664) & (!g1005) & (!sk[87]) & (g1178) & (g1227) & (!g1228)) + ((!g664) & (!g1005) & (!sk[87]) & (g1178) & (g1227) & (g1228)) + ((!g664) & (g1005) & (!sk[87]) & (!g1178) & (!g1227) & (!g1228)) + ((!g664) & (g1005) & (!sk[87]) & (!g1178) & (!g1227) & (g1228)) + ((!g664) & (g1005) & (!sk[87]) & (!g1178) & (g1227) & (!g1228)) + ((!g664) & (g1005) & (!sk[87]) & (!g1178) & (g1227) & (g1228)) + ((!g664) & (g1005) & (!sk[87]) & (g1178) & (!g1227) & (!g1228)) + ((!g664) & (g1005) & (!sk[87]) & (g1178) & (!g1227) & (g1228)) + ((!g664) & (g1005) & (!sk[87]) & (g1178) & (g1227) & (!g1228)) + ((!g664) & (g1005) & (!sk[87]) & (g1178) & (g1227) & (g1228)) + ((g664) & (!g1005) & (!sk[87]) & (!g1178) & (g1227) & (!g1228)) + ((g664) & (!g1005) & (!sk[87]) & (!g1178) & (g1227) & (g1228)) + ((g664) & (!g1005) & (!sk[87]) & (g1178) & (!g1227) & (!g1228)) + ((g664) & (!g1005) & (!sk[87]) & (g1178) & (!g1227) & (g1228)) + ((g664) & (!g1005) & (!sk[87]) & (g1178) & (g1227) & (!g1228)) + ((g664) & (!g1005) & (!sk[87]) & (g1178) & (g1227) & (g1228)) + ((g664) & (g1005) & (!sk[87]) & (!g1178) & (!g1227) & (!g1228)) + ((g664) & (g1005) & (!sk[87]) & (!g1178) & (!g1227) & (g1228)) + ((g664) & (g1005) & (!sk[87]) & (!g1178) & (g1227) & (!g1228)) + ((g664) & (g1005) & (!sk[87]) & (!g1178) & (g1227) & (g1228)) + ((g664) & (g1005) & (!sk[87]) & (g1178) & (!g1227) & (!g1228)) + ((g664) & (g1005) & (!sk[87]) & (g1178) & (!g1227) & (g1228)) + ((g664) & (g1005) & (!sk[87]) & (g1178) & (g1227) & (!g1228)) + ((g664) & (g1005) & (!sk[87]) & (g1178) & (g1227) & (g1228)) + ((g664) & (g1005) & (sk[87]) & (g1178) & (g1227) & (g1228)));
	assign g1230 = (((!sk[88]) & (!g1210) & (g1225) & (!g1229)) + ((!sk[88]) & (!g1210) & (g1225) & (g1229)) + ((!sk[88]) & (g1210) & (g1225) & (!g1229)) + ((!sk[88]) & (g1210) & (g1225) & (g1229)) + ((sk[88]) & (!g1210) & (!g1225) & (!g1229)) + ((sk[88]) & (!g1210) & (g1225) & (g1229)) + ((sk[88]) & (g1210) & (!g1225) & (g1229)) + ((sk[88]) & (g1210) & (g1225) & (!g1229)));
	assign g1231 = (((!g1068) & (!g1185) & (!g1186) & (!g1207) & (!g1209) & (g1230)) + ((!g1068) & (!g1185) & (!g1186) & (!g1207) & (g1209) & (!g1230)) + ((!g1068) & (!g1185) & (!g1186) & (g1207) & (!g1209) & (g1230)) + ((!g1068) & (!g1185) & (!g1186) & (g1207) & (g1209) & (!g1230)) + ((!g1068) & (!g1185) & (g1186) & (!g1207) & (!g1209) & (!g1230)) + ((!g1068) & (!g1185) & (g1186) & (!g1207) & (g1209) & (g1230)) + ((!g1068) & (!g1185) & (g1186) & (g1207) & (!g1209) & (g1230)) + ((!g1068) & (!g1185) & (g1186) & (g1207) & (g1209) & (!g1230)) + ((!g1068) & (g1185) & (!g1186) & (!g1207) & (!g1209) & (g1230)) + ((!g1068) & (g1185) & (!g1186) & (!g1207) & (g1209) & (!g1230)) + ((!g1068) & (g1185) & (!g1186) & (g1207) & (!g1209) & (g1230)) + ((!g1068) & (g1185) & (!g1186) & (g1207) & (g1209) & (!g1230)) + ((!g1068) & (g1185) & (g1186) & (!g1207) & (!g1209) & (!g1230)) + ((!g1068) & (g1185) & (g1186) & (!g1207) & (g1209) & (g1230)) + ((!g1068) & (g1185) & (g1186) & (g1207) & (!g1209) & (g1230)) + ((!g1068) & (g1185) & (g1186) & (g1207) & (g1209) & (!g1230)) + ((g1068) & (!g1185) & (!g1186) & (!g1207) & (!g1209) & (!g1230)) + ((g1068) & (!g1185) & (!g1186) & (!g1207) & (g1209) & (g1230)) + ((g1068) & (!g1185) & (!g1186) & (g1207) & (!g1209) & (!g1230)) + ((g1068) & (!g1185) & (!g1186) & (g1207) & (g1209) & (g1230)) + ((g1068) & (!g1185) & (g1186) & (!g1207) & (!g1209) & (g1230)) + ((g1068) & (!g1185) & (g1186) & (!g1207) & (g1209) & (!g1230)) + ((g1068) & (!g1185) & (g1186) & (g1207) & (!g1209) & (!g1230)) + ((g1068) & (!g1185) & (g1186) & (g1207) & (g1209) & (g1230)) + ((g1068) & (g1185) & (!g1186) & (!g1207) & (!g1209) & (!g1230)) + ((g1068) & (g1185) & (!g1186) & (!g1207) & (g1209) & (g1230)) + ((g1068) & (g1185) & (!g1186) & (g1207) & (!g1209) & (g1230)) + ((g1068) & (g1185) & (!g1186) & (g1207) & (g1209) & (!g1230)) + ((g1068) & (g1185) & (g1186) & (!g1207) & (!g1209) & (!g1230)) + ((g1068) & (g1185) & (g1186) & (!g1207) & (g1209) & (g1230)) + ((g1068) & (g1185) & (g1186) & (g1207) & (!g1209) & (!g1230)) + ((g1068) & (g1185) & (g1186) & (g1207) & (g1209) & (g1230)));
	assign g1232 = (((!g1186) & (!g1207) & (!g1209) & (!sk[90]) & (g1230)) + ((!g1186) & (!g1207) & (g1209) & (!sk[90]) & (g1230)) + ((!g1186) & (g1207) & (!g1209) & (!sk[90]) & (g1230)) + ((!g1186) & (g1207) & (g1209) & (!sk[90]) & (g1230)) + ((g1186) & (!g1207) & (!g1209) & (!sk[90]) & (!g1230)) + ((g1186) & (!g1207) & (!g1209) & (!sk[90]) & (g1230)) + ((g1186) & (!g1207) & (!g1209) & (sk[90]) & (!g1230)) + ((g1186) & (!g1207) & (g1209) & (!sk[90]) & (!g1230)) + ((g1186) & (!g1207) & (g1209) & (!sk[90]) & (g1230)) + ((g1186) & (!g1207) & (g1209) & (sk[90]) & (g1230)) + ((g1186) & (g1207) & (!g1209) & (!sk[90]) & (!g1230)) + ((g1186) & (g1207) & (!g1209) & (!sk[90]) & (g1230)) + ((g1186) & (g1207) & (g1209) & (!sk[90]) & (!g1230)) + ((g1186) & (g1207) & (g1209) & (!sk[90]) & (g1230)));
	assign g1233 = (((!g1210) & (!g1225) & (sk[91]) & (!g1229)) + ((!g1210) & (g1225) & (!sk[91]) & (!g1229)) + ((!g1210) & (g1225) & (!sk[91]) & (g1229)) + ((g1210) & (g1225) & (!sk[91]) & (!g1229)) + ((g1210) & (g1225) & (!sk[91]) & (g1229)) + ((g1210) & (g1225) & (sk[91]) & (!g1229)));
	assign g1234 = (((!sk[92]) & (g1211) & (g1224)) + ((sk[92]) & (g1211) & (!g1224)));
	assign g1235 = (((!g1161) & (!g1162) & (!g1174) & (g1187) & (!g1200) & (!g1225)) + ((!g1161) & (!g1162) & (g1174) & (!g1187) & (!g1200) & (!g1225)) + ((!g1161) & (!g1162) & (g1174) & (g1187) & (!g1200) & (!g1225)) + ((!g1161) & (!g1162) & (g1174) & (g1187) & (g1200) & (!g1225)) + ((!g1161) & (g1162) & (!g1174) & (!g1187) & (!g1200) & (!g1225)) + ((!g1161) & (g1162) & (!g1174) & (g1187) & (!g1200) & (!g1225)) + ((!g1161) & (g1162) & (!g1174) & (g1187) & (g1200) & (!g1225)) + ((!g1161) & (g1162) & (g1174) & (!g1187) & (!g1200) & (!g1225)) + ((!g1161) & (g1162) & (g1174) & (g1187) & (!g1200) & (!g1225)) + ((!g1161) & (g1162) & (g1174) & (g1187) & (g1200) & (!g1225)) + ((g1161) & (!g1162) & (!g1174) & (g1187) & (!g1200) & (!g1225)) + ((g1161) & (!g1162) & (g1174) & (g1187) & (!g1200) & (!g1225)) + ((g1161) & (g1162) & (!g1174) & (g1187) & (!g1200) & (!g1225)) + ((g1161) & (g1162) & (g1174) & (!g1187) & (!g1200) & (!g1225)) + ((g1161) & (g1162) & (g1174) & (g1187) & (!g1200) & (!g1225)) + ((g1161) & (g1162) & (g1174) & (g1187) & (g1200) & (!g1225)));
	assign g1236 = (((!g1212) & (!g1213) & (!sk[94]) & (!g1215) & (g1216) & (!g1223)) + ((!g1212) & (!g1213) & (!sk[94]) & (!g1215) & (g1216) & (g1223)) + ((!g1212) & (!g1213) & (!sk[94]) & (g1215) & (!g1216) & (!g1223)) + ((!g1212) & (!g1213) & (!sk[94]) & (g1215) & (!g1216) & (g1223)) + ((!g1212) & (!g1213) & (!sk[94]) & (g1215) & (g1216) & (!g1223)) + ((!g1212) & (!g1213) & (!sk[94]) & (g1215) & (g1216) & (g1223)) + ((!g1212) & (g1213) & (!sk[94]) & (!g1215) & (!g1216) & (!g1223)) + ((!g1212) & (g1213) & (!sk[94]) & (!g1215) & (!g1216) & (g1223)) + ((!g1212) & (g1213) & (!sk[94]) & (!g1215) & (g1216) & (!g1223)) + ((!g1212) & (g1213) & (!sk[94]) & (!g1215) & (g1216) & (g1223)) + ((!g1212) & (g1213) & (!sk[94]) & (g1215) & (!g1216) & (!g1223)) + ((!g1212) & (g1213) & (!sk[94]) & (g1215) & (!g1216) & (g1223)) + ((!g1212) & (g1213) & (!sk[94]) & (g1215) & (g1216) & (!g1223)) + ((!g1212) & (g1213) & (!sk[94]) & (g1215) & (g1216) & (g1223)) + ((!g1212) & (g1213) & (sk[94]) & (!g1215) & (!g1216) & (!g1223)) + ((!g1212) & (g1213) & (sk[94]) & (!g1215) & (g1216) & (g1223)) + ((!g1212) & (g1213) & (sk[94]) & (g1215) & (!g1216) & (g1223)) + ((!g1212) & (g1213) & (sk[94]) & (g1215) & (g1216) & (!g1223)) + ((g1212) & (!g1213) & (!sk[94]) & (!g1215) & (g1216) & (!g1223)) + ((g1212) & (!g1213) & (!sk[94]) & (!g1215) & (g1216) & (g1223)) + ((g1212) & (!g1213) & (!sk[94]) & (g1215) & (!g1216) & (!g1223)) + ((g1212) & (!g1213) & (!sk[94]) & (g1215) & (!g1216) & (g1223)) + ((g1212) & (!g1213) & (!sk[94]) & (g1215) & (g1216) & (!g1223)) + ((g1212) & (!g1213) & (!sk[94]) & (g1215) & (g1216) & (g1223)) + ((g1212) & (!g1213) & (sk[94]) & (!g1215) & (!g1216) & (!g1223)) + ((g1212) & (!g1213) & (sk[94]) & (!g1215) & (g1216) & (g1223)) + ((g1212) & (!g1213) & (sk[94]) & (g1215) & (!g1216) & (g1223)) + ((g1212) & (!g1213) & (sk[94]) & (g1215) & (g1216) & (!g1223)) + ((g1212) & (g1213) & (!sk[94]) & (!g1215) & (!g1216) & (!g1223)) + ((g1212) & (g1213) & (!sk[94]) & (!g1215) & (!g1216) & (g1223)) + ((g1212) & (g1213) & (!sk[94]) & (!g1215) & (g1216) & (!g1223)) + ((g1212) & (g1213) & (!sk[94]) & (!g1215) & (g1216) & (g1223)) + ((g1212) & (g1213) & (!sk[94]) & (g1215) & (!g1216) & (!g1223)) + ((g1212) & (g1213) & (!sk[94]) & (g1215) & (!g1216) & (g1223)) + ((g1212) & (g1213) & (!sk[94]) & (g1215) & (g1216) & (!g1223)) + ((g1212) & (g1213) & (!sk[94]) & (g1215) & (g1216) & (g1223)) + ((g1212) & (g1213) & (sk[94]) & (!g1215) & (!g1216) & (!g1223)) + ((g1212) & (g1213) & (sk[94]) & (!g1215) & (!g1216) & (g1223)) + ((g1212) & (g1213) & (sk[94]) & (!g1215) & (g1216) & (!g1223)) + ((g1212) & (g1213) & (sk[94]) & (!g1215) & (g1216) & (g1223)) + ((g1212) & (g1213) & (sk[94]) & (g1215) & (!g1216) & (!g1223)) + ((g1212) & (g1213) & (sk[94]) & (g1215) & (!g1216) & (g1223)) + ((g1212) & (g1213) & (sk[94]) & (g1215) & (g1216) & (!g1223)) + ((g1212) & (g1213) & (sk[94]) & (g1215) & (g1216) & (g1223)));
	assign g1237 = (((!g747) & (!g744) & (!g748) & (!g994) & (!g1040) & (!g1079)) + ((!g747) & (!g744) & (!g748) & (!g994) & (!g1040) & (g1079)) + ((!g747) & (!g744) & (!g748) & (!g994) & (g1040) & (!g1079)) + ((!g747) & (!g744) & (!g748) & (!g994) & (g1040) & (g1079)) + ((!g747) & (!g744) & (!g748) & (g994) & (!g1040) & (!g1079)) + ((!g747) & (!g744) & (!g748) & (g994) & (!g1040) & (g1079)) + ((!g747) & (!g744) & (!g748) & (g994) & (g1040) & (!g1079)) + ((!g747) & (!g744) & (!g748) & (g994) & (g1040) & (g1079)) + ((!g747) & (!g744) & (g748) & (!g994) & (!g1040) & (!g1079)) + ((!g747) & (!g744) & (g748) & (!g994) & (!g1040) & (g1079)) + ((!g747) & (!g744) & (g748) & (!g994) & (g1040) & (!g1079)) + ((!g747) & (!g744) & (g748) & (!g994) & (g1040) & (g1079)) + ((!g747) & (g744) & (!g748) & (!g994) & (g1040) & (!g1079)) + ((!g747) & (g744) & (!g748) & (!g994) & (g1040) & (g1079)) + ((!g747) & (g744) & (!g748) & (g994) & (g1040) & (!g1079)) + ((!g747) & (g744) & (!g748) & (g994) & (g1040) & (g1079)) + ((!g747) & (g744) & (g748) & (!g994) & (g1040) & (!g1079)) + ((!g747) & (g744) & (g748) & (!g994) & (g1040) & (g1079)) + ((g747) & (!g744) & (!g748) & (!g994) & (!g1040) & (g1079)) + ((g747) & (!g744) & (!g748) & (!g994) & (g1040) & (g1079)) + ((g747) & (!g744) & (!g748) & (g994) & (!g1040) & (g1079)) + ((g747) & (!g744) & (!g748) & (g994) & (g1040) & (g1079)) + ((g747) & (!g744) & (g748) & (!g994) & (!g1040) & (g1079)) + ((g747) & (!g744) & (g748) & (!g994) & (g1040) & (g1079)) + ((g747) & (g744) & (!g748) & (!g994) & (g1040) & (g1079)) + ((g747) & (g744) & (!g748) & (g994) & (g1040) & (g1079)) + ((g747) & (g744) & (g748) & (!g994) & (g1040) & (g1079)));
	assign g1238 = (((!g200) & (!g742) & (!g1040) & (!g1079) & (!g1080) & (g1237)) + ((!g200) & (!g742) & (!g1040) & (!g1079) & (g1080) & (g1237)) + ((!g200) & (!g742) & (!g1040) & (g1079) & (!g1080) & (g1237)) + ((!g200) & (!g742) & (!g1040) & (g1079) & (g1080) & (g1237)) + ((!g200) & (!g742) & (g1040) & (!g1079) & (!g1080) & (g1237)) + ((!g200) & (!g742) & (g1040) & (!g1079) & (g1080) & (g1237)) + ((!g200) & (!g742) & (g1040) & (g1079) & (!g1080) & (g1237)) + ((!g200) & (!g742) & (g1040) & (g1079) & (g1080) & (g1237)) + ((!g200) & (g742) & (!g1040) & (!g1079) & (!g1080) & (g1237)) + ((!g200) & (g742) & (!g1040) & (g1079) & (g1080) & (g1237)) + ((!g200) & (g742) & (g1040) & (!g1079) & (g1080) & (g1237)) + ((!g200) & (g742) & (g1040) & (g1079) & (!g1080) & (g1237)) + ((g200) & (!g742) & (!g1040) & (!g1079) & (!g1080) & (!g1237)) + ((g200) & (!g742) & (!g1040) & (!g1079) & (g1080) & (!g1237)) + ((g200) & (!g742) & (!g1040) & (g1079) & (!g1080) & (!g1237)) + ((g200) & (!g742) & (!g1040) & (g1079) & (g1080) & (!g1237)) + ((g200) & (!g742) & (g1040) & (!g1079) & (!g1080) & (!g1237)) + ((g200) & (!g742) & (g1040) & (!g1079) & (g1080) & (!g1237)) + ((g200) & (!g742) & (g1040) & (g1079) & (!g1080) & (!g1237)) + ((g200) & (!g742) & (g1040) & (g1079) & (g1080) & (!g1237)) + ((g200) & (g742) & (!g1040) & (!g1079) & (!g1080) & (!g1237)) + ((g200) & (g742) & (!g1040) & (!g1079) & (g1080) & (!g1237)) + ((g200) & (g742) & (!g1040) & (!g1079) & (g1080) & (g1237)) + ((g200) & (g742) & (!g1040) & (g1079) & (!g1080) & (!g1237)) + ((g200) & (g742) & (!g1040) & (g1079) & (!g1080) & (g1237)) + ((g200) & (g742) & (!g1040) & (g1079) & (g1080) & (!g1237)) + ((g200) & (g742) & (g1040) & (!g1079) & (!g1080) & (!g1237)) + ((g200) & (g742) & (g1040) & (!g1079) & (!g1080) & (g1237)) + ((g200) & (g742) & (g1040) & (!g1079) & (g1080) & (!g1237)) + ((g200) & (g742) & (g1040) & (g1079) & (!g1080) & (!g1237)) + ((g200) & (g742) & (g1040) & (g1079) & (g1080) & (!g1237)) + ((g200) & (g742) & (g1040) & (g1079) & (g1080) & (g1237)));
	assign g1239 = (((!g252) & (!g683) & (!g681) & (!g1219) & (!g1220) & (g1221)) + ((!g252) & (!g683) & (!g681) & (g1219) & (!g1220) & (g1221)) + ((!g252) & (!g683) & (!g681) & (g1219) & (g1220) & (g1221)) + ((!g252) & (!g683) & (g681) & (!g1219) & (!g1220) & (g1221)) + ((!g252) & (!g683) & (g681) & (g1219) & (!g1220) & (g1221)) + ((!g252) & (!g683) & (g681) & (g1219) & (g1220) & (g1221)) + ((!g252) & (g683) & (!g681) & (!g1219) & (!g1220) & (!g1221)) + ((!g252) & (g683) & (!g681) & (g1219) & (!g1220) & (!g1221)) + ((!g252) & (g683) & (!g681) & (g1219) & (g1220) & (!g1221)) + ((!g252) & (g683) & (g681) & (!g1219) & (!g1220) & (!g1221)) + ((!g252) & (g683) & (g681) & (g1219) & (!g1220) & (!g1221)) + ((!g252) & (g683) & (g681) & (g1219) & (g1220) & (!g1221)) + ((g252) & (!g683) & (!g681) & (!g1219) & (g1220) & (!g1221)) + ((g252) & (!g683) & (g681) & (!g1219) & (g1220) & (g1221)) + ((g252) & (g683) & (!g681) & (!g1219) & (g1220) & (g1221)) + ((g252) & (g683) & (g681) & (!g1219) & (g1220) & (!g1221)));
	assign g1240 = (((!g202) & (!g759) & (!g1217) & (!g1218) & (g1222) & (!g1239)) + ((!g202) & (!g759) & (!g1217) & (g1218) & (!g1222) & (!g1239)) + ((!g202) & (!g759) & (!g1217) & (g1218) & (g1222) & (!g1239)) + ((!g202) & (!g759) & (g1217) & (!g1218) & (g1222) & (!g1239)) + ((!g202) & (!g759) & (g1217) & (g1218) & (!g1222) & (!g1239)) + ((!g202) & (!g759) & (g1217) & (g1218) & (g1222) & (!g1239)) + ((!g202) & (g759) & (!g1217) & (!g1218) & (g1222) & (!g1239)) + ((!g202) & (g759) & (!g1217) & (g1218) & (g1222) & (!g1239)) + ((!g202) & (g759) & (g1217) & (!g1218) & (g1222) & (!g1239)) + ((!g202) & (g759) & (g1217) & (g1218) & (!g1222) & (!g1239)) + ((!g202) & (g759) & (g1217) & (g1218) & (g1222) & (!g1239)) + ((g202) & (!g759) & (!g1217) & (!g1218) & (!g1222) & (!g1239)) + ((g202) & (!g759) & (!g1217) & (!g1218) & (g1222) & (!g1239)) + ((g202) & (!g759) & (!g1217) & (g1218) & (g1222) & (!g1239)) + ((g202) & (!g759) & (g1217) & (!g1218) & (!g1222) & (!g1239)) + ((g202) & (!g759) & (g1217) & (!g1218) & (g1222) & (!g1239)) + ((g202) & (!g759) & (g1217) & (g1218) & (g1222) & (!g1239)) + ((g202) & (g759) & (!g1217) & (!g1218) & (!g1222) & (!g1239)) + ((g202) & (g759) & (!g1217) & (!g1218) & (g1222) & (!g1239)) + ((g202) & (g759) & (!g1217) & (g1218) & (!g1222) & (!g1239)) + ((g202) & (g759) & (!g1217) & (g1218) & (g1222) & (!g1239)) + ((g202) & (g759) & (g1217) & (!g1218) & (!g1222) & (!g1239)) + ((g202) & (g759) & (g1217) & (!g1218) & (g1222) & (!g1239)) + ((g202) & (g759) & (g1217) & (g1218) & (g1222) & (!g1239)));
	assign g1241 = (((!g764) & (!g762) & (!g765) & (!g962) & (!g963) & (!g971)) + ((!g764) & (!g762) & (!g765) & (!g962) & (!g963) & (g971)) + ((!g764) & (!g762) & (!g765) & (!g962) & (g963) & (!g971)) + ((!g764) & (!g762) & (!g765) & (!g962) & (g963) & (g971)) + ((!g764) & (!g762) & (!g765) & (g962) & (!g963) & (!g971)) + ((!g764) & (!g762) & (!g765) & (g962) & (!g963) & (g971)) + ((!g764) & (!g762) & (!g765) & (g962) & (g963) & (!g971)) + ((!g764) & (!g762) & (!g765) & (g962) & (g963) & (g971)) + ((!g764) & (!g762) & (g765) & (!g962) & (!g963) & (!g971)) + ((!g764) & (!g762) & (g765) & (!g962) & (!g963) & (g971)) + ((!g764) & (!g762) & (g765) & (g962) & (!g963) & (!g971)) + ((!g764) & (!g762) & (g765) & (g962) & (!g963) & (g971)) + ((!g764) & (g762) & (!g765) & (g962) & (!g963) & (!g971)) + ((!g764) & (g762) & (!g765) & (g962) & (!g963) & (g971)) + ((!g764) & (g762) & (!g765) & (g962) & (g963) & (!g971)) + ((!g764) & (g762) & (!g765) & (g962) & (g963) & (g971)) + ((!g764) & (g762) & (g765) & (g962) & (!g963) & (!g971)) + ((!g764) & (g762) & (g765) & (g962) & (!g963) & (g971)) + ((g764) & (!g762) & (!g765) & (!g962) & (!g963) & (!g971)) + ((g764) & (!g762) & (!g765) & (!g962) & (g963) & (!g971)) + ((g764) & (!g762) & (!g765) & (g962) & (!g963) & (!g971)) + ((g764) & (!g762) & (!g765) & (g962) & (g963) & (!g971)) + ((g764) & (!g762) & (g765) & (!g962) & (!g963) & (!g971)) + ((g764) & (!g762) & (g765) & (g962) & (!g963) & (!g971)) + ((g764) & (g762) & (!g765) & (g962) & (!g963) & (!g971)) + ((g764) & (g762) & (!g765) & (g962) & (g963) & (!g971)) + ((g764) & (g762) & (g765) & (g962) & (!g963) & (!g971)));
	assign g1242 = (((!g252) & (g683) & (!g681) & (!g719) & (!g729) & (!g1168)) + ((!g252) & (g683) & (!g681) & (!g719) & (g729) & (!g1168)) + ((!g252) & (g683) & (!g681) & (g719) & (!g729) & (!g1168)) + ((!g252) & (g683) & (!g681) & (g719) & (g729) & (!g1168)) + ((!g252) & (g683) & (g681) & (!g719) & (!g729) & (!g1168)) + ((!g252) & (g683) & (g681) & (!g719) & (g729) & (!g1168)) + ((!g252) & (g683) & (g681) & (g719) & (!g729) & (!g1168)) + ((!g252) & (g683) & (g681) & (g719) & (g729) & (!g1168)) + ((g252) & (!g683) & (!g681) & (!g719) & (!g729) & (g1168)) + ((g252) & (g683) & (!g681) & (!g719) & (!g729) & (!g1168)) + ((g252) & (g683) & (!g681) & (!g719) & (!g729) & (g1168)) + ((g252) & (g683) & (!g681) & (!g719) & (g729) & (!g1168)) + ((g252) & (g683) & (!g681) & (!g719) & (g729) & (g1168)) + ((g252) & (g683) & (!g681) & (g719) & (!g729) & (!g1168)) + ((g252) & (g683) & (!g681) & (g719) & (!g729) & (g1168)) + ((g252) & (g683) & (!g681) & (g719) & (g729) & (!g1168)) + ((g252) & (g683) & (!g681) & (g719) & (g729) & (g1168)) + ((g252) & (g683) & (g681) & (!g719) & (!g729) & (!g1168)) + ((g252) & (g683) & (g681) & (!g719) & (!g729) & (g1168)) + ((g252) & (g683) & (g681) & (!g719) & (g729) & (!g1168)) + ((g252) & (g683) & (g681) & (!g719) & (g729) & (g1168)) + ((g252) & (g683) & (g681) & (g719) & (!g729) & (!g1168)) + ((g252) & (g683) & (g681) & (g719) & (!g729) & (g1168)) + ((g252) & (g683) & (g681) & (g719) & (g729) & (g1168)));
	assign g1243 = (((!sk[101]) & (!g2) & (!g252) & (!g683) & (g718)) + ((!sk[101]) & (!g2) & (!g252) & (g683) & (g718)) + ((!sk[101]) & (!g2) & (g252) & (!g683) & (g718)) + ((!sk[101]) & (!g2) & (g252) & (g683) & (g718)) + ((!sk[101]) & (g2) & (!g252) & (!g683) & (!g718)) + ((!sk[101]) & (g2) & (!g252) & (!g683) & (g718)) + ((!sk[101]) & (g2) & (!g252) & (g683) & (!g718)) + ((!sk[101]) & (g2) & (!g252) & (g683) & (g718)) + ((!sk[101]) & (g2) & (g252) & (!g683) & (!g718)) + ((!sk[101]) & (g2) & (g252) & (!g683) & (g718)) + ((!sk[101]) & (g2) & (g252) & (g683) & (!g718)) + ((!sk[101]) & (g2) & (g252) & (g683) & (g718)) + ((sk[101]) & (!g2) & (!g252) & (g683) & (!g718)) + ((sk[101]) & (!g2) & (!g252) & (g683) & (g718)) + ((sk[101]) & (!g2) & (g252) & (!g683) & (g718)) + ((sk[101]) & (!g2) & (g252) & (g683) & (!g718)) + ((sk[101]) & (g2) & (!g252) & (!g683) & (!g718)) + ((sk[101]) & (g2) & (!g252) & (!g683) & (g718)) + ((sk[101]) & (g2) & (g252) & (!g683) & (!g718)) + ((sk[101]) & (g2) & (g252) & (g683) & (g718)));
	assign g1244 = (((!g869) & (!g847) & (!g845) & (!g870) & (!g848) & (!g863)) + ((!g869) & (!g847) & (!g845) & (!g870) & (!g848) & (g863)) + ((!g869) & (!g847) & (!g845) & (!g870) & (g848) & (!g863)) + ((!g869) & (!g847) & (!g845) & (!g870) & (g848) & (g863)) + ((!g869) & (!g847) & (!g845) & (g870) & (!g848) & (!g863)) + ((!g869) & (!g847) & (!g845) & (g870) & (!g848) & (g863)) + ((!g869) & (!g847) & (!g845) & (g870) & (g848) & (!g863)) + ((!g869) & (!g847) & (!g845) & (g870) & (g848) & (g863)) + ((!g869) & (!g847) & (g845) & (g870) & (!g848) & (!g863)) + ((!g869) & (!g847) & (g845) & (g870) & (!g848) & (g863)) + ((!g869) & (!g847) & (g845) & (g870) & (g848) & (!g863)) + ((!g869) & (!g847) & (g845) & (g870) & (g848) & (g863)) + ((!g869) & (g847) & (!g845) & (!g870) & (!g848) & (!g863)) + ((!g869) & (g847) & (!g845) & (!g870) & (g848) & (!g863)) + ((!g869) & (g847) & (!g845) & (g870) & (!g848) & (!g863)) + ((!g869) & (g847) & (!g845) & (g870) & (g848) & (!g863)) + ((!g869) & (g847) & (g845) & (g870) & (!g848) & (!g863)) + ((!g869) & (g847) & (g845) & (g870) & (g848) & (!g863)) + ((g869) & (!g847) & (!g845) & (!g870) & (!g848) & (!g863)) + ((g869) & (!g847) & (!g845) & (!g870) & (!g848) & (g863)) + ((g869) & (!g847) & (!g845) & (g870) & (!g848) & (!g863)) + ((g869) & (!g847) & (!g845) & (g870) & (!g848) & (g863)) + ((g869) & (!g847) & (g845) & (g870) & (!g848) & (!g863)) + ((g869) & (!g847) & (g845) & (g870) & (!g848) & (g863)) + ((g869) & (g847) & (!g845) & (!g870) & (!g848) & (!g863)) + ((g869) & (g847) & (!g845) & (g870) & (!g848) & (!g863)) + ((g869) & (g847) & (g845) & (g870) & (!g848) & (!g863)));
	assign g1245 = (((!g252) & (!g843) & (!g899) & (!g1242) & (!g1243) & (!g1244)) + ((!g252) & (!g843) & (!g899) & (!g1242) & (g1243) & (g1244)) + ((!g252) & (!g843) & (!g899) & (g1242) & (!g1243) & (g1244)) + ((!g252) & (!g843) & (!g899) & (g1242) & (g1243) & (!g1244)) + ((!g252) & (!g843) & (g899) & (!g1242) & (!g1243) & (!g1244)) + ((!g252) & (!g843) & (g899) & (!g1242) & (g1243) & (g1244)) + ((!g252) & (!g843) & (g899) & (g1242) & (!g1243) & (g1244)) + ((!g252) & (!g843) & (g899) & (g1242) & (g1243) & (!g1244)) + ((!g252) & (g843) & (!g899) & (!g1242) & (!g1243) & (!g1244)) + ((!g252) & (g843) & (!g899) & (!g1242) & (!g1243) & (g1244)) + ((!g252) & (g843) & (!g899) & (g1242) & (g1243) & (!g1244)) + ((!g252) & (g843) & (!g899) & (g1242) & (g1243) & (g1244)) + ((!g252) & (g843) & (g899) & (!g1242) & (!g1243) & (!g1244)) + ((!g252) & (g843) & (g899) & (!g1242) & (g1243) & (g1244)) + ((!g252) & (g843) & (g899) & (g1242) & (!g1243) & (g1244)) + ((!g252) & (g843) & (g899) & (g1242) & (g1243) & (!g1244)) + ((g252) & (!g843) & (!g899) & (!g1242) & (!g1243) & (g1244)) + ((g252) & (!g843) & (!g899) & (!g1242) & (g1243) & (!g1244)) + ((g252) & (!g843) & (!g899) & (g1242) & (!g1243) & (!g1244)) + ((g252) & (!g843) & (!g899) & (g1242) & (g1243) & (g1244)) + ((g252) & (!g843) & (g899) & (!g1242) & (!g1243) & (g1244)) + ((g252) & (!g843) & (g899) & (!g1242) & (g1243) & (!g1244)) + ((g252) & (!g843) & (g899) & (g1242) & (!g1243) & (!g1244)) + ((g252) & (!g843) & (g899) & (g1242) & (g1243) & (g1244)) + ((g252) & (g843) & (!g899) & (!g1242) & (g1243) & (!g1244)) + ((g252) & (g843) & (!g899) & (!g1242) & (g1243) & (g1244)) + ((g252) & (g843) & (!g899) & (g1242) & (!g1243) & (!g1244)) + ((g252) & (g843) & (!g899) & (g1242) & (!g1243) & (g1244)) + ((g252) & (g843) & (g899) & (!g1242) & (!g1243) & (g1244)) + ((g252) & (g843) & (g899) & (!g1242) & (g1243) & (!g1244)) + ((g252) & (g843) & (g899) & (g1242) & (!g1243) & (!g1244)) + ((g252) & (g843) & (g899) & (g1242) & (g1243) & (g1244)));
	assign g1246 = (((!g202) & (!g759) & (!g972) & (!g1241) & (sk[104]) & (g1245)) + ((!g202) & (!g759) & (!g972) & (g1241) & (!sk[104]) & (!g1245)) + ((!g202) & (!g759) & (!g972) & (g1241) & (!sk[104]) & (g1245)) + ((!g202) & (!g759) & (!g972) & (g1241) & (sk[104]) & (!g1245)) + ((!g202) & (!g759) & (g972) & (!g1241) & (!sk[104]) & (!g1245)) + ((!g202) & (!g759) & (g972) & (!g1241) & (!sk[104]) & (g1245)) + ((!g202) & (!g759) & (g972) & (!g1241) & (sk[104]) & (g1245)) + ((!g202) & (!g759) & (g972) & (g1241) & (!sk[104]) & (!g1245)) + ((!g202) & (!g759) & (g972) & (g1241) & (!sk[104]) & (g1245)) + ((!g202) & (!g759) & (g972) & (g1241) & (sk[104]) & (!g1245)) + ((!g202) & (g759) & (!g972) & (!g1241) & (!sk[104]) & (!g1245)) + ((!g202) & (g759) & (!g972) & (!g1241) & (!sk[104]) & (g1245)) + ((!g202) & (g759) & (!g972) & (!g1241) & (sk[104]) & (g1245)) + ((!g202) & (g759) & (!g972) & (g1241) & (!sk[104]) & (!g1245)) + ((!g202) & (g759) & (!g972) & (g1241) & (!sk[104]) & (g1245)) + ((!g202) & (g759) & (!g972) & (g1241) & (sk[104]) & (g1245)) + ((!g202) & (g759) & (g972) & (!g1241) & (!sk[104]) & (!g1245)) + ((!g202) & (g759) & (g972) & (!g1241) & (!sk[104]) & (g1245)) + ((!g202) & (g759) & (g972) & (!g1241) & (sk[104]) & (g1245)) + ((!g202) & (g759) & (g972) & (g1241) & (!sk[104]) & (!g1245)) + ((!g202) & (g759) & (g972) & (g1241) & (!sk[104]) & (g1245)) + ((!g202) & (g759) & (g972) & (g1241) & (sk[104]) & (!g1245)) + ((g202) & (!g759) & (!g972) & (!g1241) & (sk[104]) & (!g1245)) + ((g202) & (!g759) & (!g972) & (g1241) & (!sk[104]) & (!g1245)) + ((g202) & (!g759) & (!g972) & (g1241) & (!sk[104]) & (g1245)) + ((g202) & (!g759) & (!g972) & (g1241) & (sk[104]) & (g1245)) + ((g202) & (!g759) & (g972) & (!g1241) & (!sk[104]) & (!g1245)) + ((g202) & (!g759) & (g972) & (!g1241) & (!sk[104]) & (g1245)) + ((g202) & (!g759) & (g972) & (!g1241) & (sk[104]) & (!g1245)) + ((g202) & (!g759) & (g972) & (g1241) & (!sk[104]) & (!g1245)) + ((g202) & (!g759) & (g972) & (g1241) & (!sk[104]) & (g1245)) + ((g202) & (!g759) & (g972) & (g1241) & (sk[104]) & (g1245)) + ((g202) & (g759) & (!g972) & (!g1241) & (!sk[104]) & (!g1245)) + ((g202) & (g759) & (!g972) & (!g1241) & (!sk[104]) & (g1245)) + ((g202) & (g759) & (!g972) & (!g1241) & (sk[104]) & (!g1245)) + ((g202) & (g759) & (!g972) & (g1241) & (!sk[104]) & (!g1245)) + ((g202) & (g759) & (!g972) & (g1241) & (!sk[104]) & (g1245)) + ((g202) & (g759) & (!g972) & (g1241) & (sk[104]) & (!g1245)) + ((g202) & (g759) & (g972) & (!g1241) & (!sk[104]) & (!g1245)) + ((g202) & (g759) & (g972) & (!g1241) & (!sk[104]) & (g1245)) + ((g202) & (g759) & (g972) & (!g1241) & (sk[104]) & (!g1245)) + ((g202) & (g759) & (g972) & (g1241) & (!sk[104]) & (!g1245)) + ((g202) & (g759) & (g972) & (g1241) & (!sk[104]) & (g1245)) + ((g202) & (g759) & (g972) & (g1241) & (sk[104]) & (g1245)));
	assign g1247 = (((!g1215) & (!g1216) & (!g1223) & (!g1238) & (!g1240) & (!g1246)) + ((!g1215) & (!g1216) & (!g1223) & (!g1238) & (g1240) & (g1246)) + ((!g1215) & (!g1216) & (!g1223) & (g1238) & (!g1240) & (g1246)) + ((!g1215) & (!g1216) & (!g1223) & (g1238) & (g1240) & (!g1246)) + ((!g1215) & (!g1216) & (g1223) & (!g1238) & (!g1240) & (!g1246)) + ((!g1215) & (!g1216) & (g1223) & (!g1238) & (g1240) & (g1246)) + ((!g1215) & (!g1216) & (g1223) & (g1238) & (!g1240) & (g1246)) + ((!g1215) & (!g1216) & (g1223) & (g1238) & (g1240) & (!g1246)) + ((!g1215) & (g1216) & (!g1223) & (!g1238) & (!g1240) & (g1246)) + ((!g1215) & (g1216) & (!g1223) & (!g1238) & (g1240) & (!g1246)) + ((!g1215) & (g1216) & (!g1223) & (g1238) & (!g1240) & (!g1246)) + ((!g1215) & (g1216) & (!g1223) & (g1238) & (g1240) & (g1246)) + ((!g1215) & (g1216) & (g1223) & (!g1238) & (!g1240) & (!g1246)) + ((!g1215) & (g1216) & (g1223) & (!g1238) & (g1240) & (g1246)) + ((!g1215) & (g1216) & (g1223) & (g1238) & (!g1240) & (g1246)) + ((!g1215) & (g1216) & (g1223) & (g1238) & (g1240) & (!g1246)) + ((g1215) & (!g1216) & (!g1223) & (!g1238) & (!g1240) & (g1246)) + ((g1215) & (!g1216) & (!g1223) & (!g1238) & (g1240) & (!g1246)) + ((g1215) & (!g1216) & (!g1223) & (g1238) & (!g1240) & (!g1246)) + ((g1215) & (!g1216) & (!g1223) & (g1238) & (g1240) & (g1246)) + ((g1215) & (!g1216) & (g1223) & (!g1238) & (!g1240) & (!g1246)) + ((g1215) & (!g1216) & (g1223) & (!g1238) & (g1240) & (g1246)) + ((g1215) & (!g1216) & (g1223) & (g1238) & (!g1240) & (g1246)) + ((g1215) & (!g1216) & (g1223) & (g1238) & (g1240) & (!g1246)) + ((g1215) & (g1216) & (!g1223) & (!g1238) & (!g1240) & (g1246)) + ((g1215) & (g1216) & (!g1223) & (!g1238) & (g1240) & (!g1246)) + ((g1215) & (g1216) & (!g1223) & (g1238) & (!g1240) & (!g1246)) + ((g1215) & (g1216) & (!g1223) & (g1238) & (g1240) & (g1246)) + ((g1215) & (g1216) & (g1223) & (!g1238) & (!g1240) & (g1246)) + ((g1215) & (g1216) & (g1223) & (!g1238) & (g1240) & (!g1246)) + ((g1215) & (g1216) & (g1223) & (g1238) & (!g1240) & (!g1246)) + ((g1215) & (g1216) & (g1223) & (g1238) & (g1240) & (g1246)));
	assign g1248 = (((!sk[106]) & (g1236) & (g1247)) + ((sk[106]) & (!g1236) & (g1247)) + ((sk[106]) & (g1236) & (!g1247)));
	assign g1249 = (((!g601) & (!g231) & (!sk[107]) & (!g73) & (g162)) + ((!g601) & (!g231) & (!sk[107]) & (g73) & (g162)) + ((!g601) & (g231) & (!sk[107]) & (!g73) & (g162)) + ((!g601) & (g231) & (!sk[107]) & (g73) & (g162)) + ((!g601) & (g231) & (sk[107]) & (!g73) & (!g162)) + ((g601) & (!g231) & (!sk[107]) & (!g73) & (!g162)) + ((g601) & (!g231) & (!sk[107]) & (!g73) & (g162)) + ((g601) & (!g231) & (!sk[107]) & (g73) & (!g162)) + ((g601) & (!g231) & (!sk[107]) & (g73) & (g162)) + ((g601) & (g231) & (!sk[107]) & (!g73) & (!g162)) + ((g601) & (g231) & (!sk[107]) & (!g73) & (g162)) + ((g601) & (g231) & (!sk[107]) & (g73) & (!g162)) + ((g601) & (g231) & (!sk[107]) & (g73) & (g162)));
	assign g1250 = (((!g9) & (!g70) & (!g58) & (!sk[108]) & (g18) & (!g1202)) + ((!g9) & (!g70) & (!g58) & (!sk[108]) & (g18) & (g1202)) + ((!g9) & (!g70) & (!g58) & (sk[108]) & (!g18) & (g1202)) + ((!g9) & (!g70) & (!g58) & (sk[108]) & (g18) & (g1202)) + ((!g9) & (!g70) & (g58) & (!sk[108]) & (!g18) & (!g1202)) + ((!g9) & (!g70) & (g58) & (!sk[108]) & (!g18) & (g1202)) + ((!g9) & (!g70) & (g58) & (!sk[108]) & (g18) & (!g1202)) + ((!g9) & (!g70) & (g58) & (!sk[108]) & (g18) & (g1202)) + ((!g9) & (!g70) & (g58) & (sk[108]) & (!g18) & (g1202)) + ((!g9) & (!g70) & (g58) & (sk[108]) & (g18) & (g1202)) + ((!g9) & (g70) & (!g58) & (!sk[108]) & (!g18) & (!g1202)) + ((!g9) & (g70) & (!g58) & (!sk[108]) & (!g18) & (g1202)) + ((!g9) & (g70) & (!g58) & (!sk[108]) & (g18) & (!g1202)) + ((!g9) & (g70) & (!g58) & (!sk[108]) & (g18) & (g1202)) + ((!g9) & (g70) & (!g58) & (sk[108]) & (!g18) & (g1202)) + ((!g9) & (g70) & (g58) & (!sk[108]) & (!g18) & (!g1202)) + ((!g9) & (g70) & (g58) & (!sk[108]) & (!g18) & (g1202)) + ((!g9) & (g70) & (g58) & (!sk[108]) & (g18) & (!g1202)) + ((!g9) & (g70) & (g58) & (!sk[108]) & (g18) & (g1202)) + ((!g9) & (g70) & (g58) & (sk[108]) & (!g18) & (g1202)) + ((g9) & (!g70) & (!g58) & (!sk[108]) & (g18) & (!g1202)) + ((g9) & (!g70) & (!g58) & (!sk[108]) & (g18) & (g1202)) + ((g9) & (!g70) & (!g58) & (sk[108]) & (!g18) & (g1202)) + ((g9) & (!g70) & (!g58) & (sk[108]) & (g18) & (g1202)) + ((g9) & (!g70) & (g58) & (!sk[108]) & (!g18) & (!g1202)) + ((g9) & (!g70) & (g58) & (!sk[108]) & (!g18) & (g1202)) + ((g9) & (!g70) & (g58) & (!sk[108]) & (g18) & (!g1202)) + ((g9) & (!g70) & (g58) & (!sk[108]) & (g18) & (g1202)) + ((g9) & (g70) & (!g58) & (!sk[108]) & (!g18) & (!g1202)) + ((g9) & (g70) & (!g58) & (!sk[108]) & (!g18) & (g1202)) + ((g9) & (g70) & (!g58) & (!sk[108]) & (g18) & (!g1202)) + ((g9) & (g70) & (!g58) & (!sk[108]) & (g18) & (g1202)) + ((g9) & (g70) & (!g58) & (sk[108]) & (!g18) & (g1202)) + ((g9) & (g70) & (g58) & (!sk[108]) & (!g18) & (!g1202)) + ((g9) & (g70) & (g58) & (!sk[108]) & (!g18) & (g1202)) + ((g9) & (g70) & (g58) & (!sk[108]) & (g18) & (!g1202)) + ((g9) & (g70) & (g58) & (!sk[108]) & (g18) & (g1202)));
	assign g1251 = (((!g58) & (!g104) & (!g593) & (!g35) & (!g268) & (g334)) + ((!g58) & (g104) & (!g593) & (!g35) & (!g268) & (g334)) + ((g58) & (!g104) & (!g593) & (!g35) & (!g268) & (g334)));
	assign g1252 = (((!g557) & (!g1227) & (!g1249) & (!sk[110]) & (g1250) & (!g1251)) + ((!g557) & (!g1227) & (!g1249) & (!sk[110]) & (g1250) & (g1251)) + ((!g557) & (!g1227) & (g1249) & (!sk[110]) & (!g1250) & (!g1251)) + ((!g557) & (!g1227) & (g1249) & (!sk[110]) & (!g1250) & (g1251)) + ((!g557) & (!g1227) & (g1249) & (!sk[110]) & (g1250) & (!g1251)) + ((!g557) & (!g1227) & (g1249) & (!sk[110]) & (g1250) & (g1251)) + ((!g557) & (g1227) & (!g1249) & (!sk[110]) & (!g1250) & (!g1251)) + ((!g557) & (g1227) & (!g1249) & (!sk[110]) & (!g1250) & (g1251)) + ((!g557) & (g1227) & (!g1249) & (!sk[110]) & (g1250) & (!g1251)) + ((!g557) & (g1227) & (!g1249) & (!sk[110]) & (g1250) & (g1251)) + ((!g557) & (g1227) & (g1249) & (!sk[110]) & (!g1250) & (!g1251)) + ((!g557) & (g1227) & (g1249) & (!sk[110]) & (!g1250) & (g1251)) + ((!g557) & (g1227) & (g1249) & (!sk[110]) & (g1250) & (!g1251)) + ((!g557) & (g1227) & (g1249) & (!sk[110]) & (g1250) & (g1251)) + ((g557) & (!g1227) & (!g1249) & (!sk[110]) & (g1250) & (!g1251)) + ((g557) & (!g1227) & (!g1249) & (!sk[110]) & (g1250) & (g1251)) + ((g557) & (!g1227) & (g1249) & (!sk[110]) & (!g1250) & (!g1251)) + ((g557) & (!g1227) & (g1249) & (!sk[110]) & (!g1250) & (g1251)) + ((g557) & (!g1227) & (g1249) & (!sk[110]) & (g1250) & (!g1251)) + ((g557) & (!g1227) & (g1249) & (!sk[110]) & (g1250) & (g1251)) + ((g557) & (g1227) & (!g1249) & (!sk[110]) & (!g1250) & (!g1251)) + ((g557) & (g1227) & (!g1249) & (!sk[110]) & (!g1250) & (g1251)) + ((g557) & (g1227) & (!g1249) & (!sk[110]) & (g1250) & (!g1251)) + ((g557) & (g1227) & (!g1249) & (!sk[110]) & (g1250) & (g1251)) + ((g557) & (g1227) & (g1249) & (!sk[110]) & (!g1250) & (!g1251)) + ((g557) & (g1227) & (g1249) & (!sk[110]) & (!g1250) & (g1251)) + ((g557) & (g1227) & (g1249) & (!sk[110]) & (g1250) & (!g1251)) + ((g557) & (g1227) & (g1249) & (!sk[110]) & (g1250) & (g1251)) + ((g557) & (g1227) & (g1249) & (sk[110]) & (g1250) & (g1251)));
	assign g1253 = (((!sk[111]) & (!g1234) & (!g1235) & (!g1248) & (g1252)) + ((!sk[111]) & (!g1234) & (!g1235) & (g1248) & (g1252)) + ((!sk[111]) & (!g1234) & (g1235) & (!g1248) & (g1252)) + ((!sk[111]) & (!g1234) & (g1235) & (g1248) & (g1252)) + ((!sk[111]) & (g1234) & (!g1235) & (!g1248) & (!g1252)) + ((!sk[111]) & (g1234) & (!g1235) & (!g1248) & (g1252)) + ((!sk[111]) & (g1234) & (!g1235) & (g1248) & (!g1252)) + ((!sk[111]) & (g1234) & (!g1235) & (g1248) & (g1252)) + ((!sk[111]) & (g1234) & (g1235) & (!g1248) & (!g1252)) + ((!sk[111]) & (g1234) & (g1235) & (!g1248) & (g1252)) + ((!sk[111]) & (g1234) & (g1235) & (g1248) & (!g1252)) + ((!sk[111]) & (g1234) & (g1235) & (g1248) & (g1252)) + ((sk[111]) & (!g1234) & (!g1235) & (!g1248) & (!g1252)) + ((sk[111]) & (!g1234) & (!g1235) & (g1248) & (g1252)) + ((sk[111]) & (!g1234) & (g1235) & (!g1248) & (g1252)) + ((sk[111]) & (!g1234) & (g1235) & (g1248) & (!g1252)) + ((sk[111]) & (g1234) & (!g1235) & (!g1248) & (g1252)) + ((sk[111]) & (g1234) & (!g1235) & (g1248) & (!g1252)) + ((sk[111]) & (g1234) & (g1235) & (!g1248) & (g1252)) + ((sk[111]) & (g1234) & (g1235) & (g1248) & (!g1252)));
	assign g1254 = (((!sk[112]) & (!g1209) & (!g1230) & (!g1233) & (g1253)) + ((!sk[112]) & (!g1209) & (!g1230) & (g1233) & (g1253)) + ((!sk[112]) & (!g1209) & (g1230) & (!g1233) & (g1253)) + ((!sk[112]) & (!g1209) & (g1230) & (g1233) & (g1253)) + ((!sk[112]) & (g1209) & (!g1230) & (!g1233) & (!g1253)) + ((!sk[112]) & (g1209) & (!g1230) & (!g1233) & (g1253)) + ((!sk[112]) & (g1209) & (!g1230) & (g1233) & (!g1253)) + ((!sk[112]) & (g1209) & (!g1230) & (g1233) & (g1253)) + ((!sk[112]) & (g1209) & (g1230) & (!g1233) & (!g1253)) + ((!sk[112]) & (g1209) & (g1230) & (!g1233) & (g1253)) + ((!sk[112]) & (g1209) & (g1230) & (g1233) & (!g1253)) + ((!sk[112]) & (g1209) & (g1230) & (g1233) & (g1253)) + ((sk[112]) & (!g1209) & (!g1230) & (!g1233) & (g1253)) + ((sk[112]) & (!g1209) & (!g1230) & (g1233) & (!g1253)) + ((sk[112]) & (!g1209) & (g1230) & (!g1233) & (g1253)) + ((sk[112]) & (!g1209) & (g1230) & (g1233) & (!g1253)) + ((sk[112]) & (g1209) & (!g1230) & (!g1233) & (!g1253)) + ((sk[112]) & (g1209) & (!g1230) & (g1233) & (!g1253)) + ((sk[112]) & (g1209) & (g1230) & (!g1233) & (g1253)) + ((sk[112]) & (g1209) & (g1230) & (g1233) & (!g1253)));
	assign g1255 = (((!g1185) & (!g1186) & (!g1207) & (!sk[113]) & (g1209) & (!g1230)) + ((!g1185) & (!g1186) & (!g1207) & (!sk[113]) & (g1209) & (g1230)) + ((!g1185) & (!g1186) & (g1207) & (!sk[113]) & (!g1209) & (!g1230)) + ((!g1185) & (!g1186) & (g1207) & (!sk[113]) & (!g1209) & (g1230)) + ((!g1185) & (!g1186) & (g1207) & (!sk[113]) & (g1209) & (!g1230)) + ((!g1185) & (!g1186) & (g1207) & (!sk[113]) & (g1209) & (g1230)) + ((!g1185) & (g1186) & (!g1207) & (!sk[113]) & (!g1209) & (!g1230)) + ((!g1185) & (g1186) & (!g1207) & (!sk[113]) & (!g1209) & (g1230)) + ((!g1185) & (g1186) & (!g1207) & (!sk[113]) & (g1209) & (!g1230)) + ((!g1185) & (g1186) & (!g1207) & (!sk[113]) & (g1209) & (g1230)) + ((!g1185) & (g1186) & (g1207) & (!sk[113]) & (!g1209) & (!g1230)) + ((!g1185) & (g1186) & (g1207) & (!sk[113]) & (!g1209) & (g1230)) + ((!g1185) & (g1186) & (g1207) & (!sk[113]) & (g1209) & (!g1230)) + ((!g1185) & (g1186) & (g1207) & (!sk[113]) & (g1209) & (g1230)) + ((g1185) & (!g1186) & (!g1207) & (!sk[113]) & (g1209) & (!g1230)) + ((g1185) & (!g1186) & (!g1207) & (!sk[113]) & (g1209) & (g1230)) + ((g1185) & (!g1186) & (g1207) & (!sk[113]) & (!g1209) & (!g1230)) + ((g1185) & (!g1186) & (g1207) & (!sk[113]) & (!g1209) & (g1230)) + ((g1185) & (!g1186) & (g1207) & (!sk[113]) & (g1209) & (!g1230)) + ((g1185) & (!g1186) & (g1207) & (!sk[113]) & (g1209) & (g1230)) + ((g1185) & (!g1186) & (g1207) & (sk[113]) & (!g1209) & (g1230)) + ((g1185) & (!g1186) & (g1207) & (sk[113]) & (g1209) & (!g1230)) + ((g1185) & (g1186) & (!g1207) & (!sk[113]) & (!g1209) & (!g1230)) + ((g1185) & (g1186) & (!g1207) & (!sk[113]) & (!g1209) & (g1230)) + ((g1185) & (g1186) & (!g1207) & (!sk[113]) & (g1209) & (!g1230)) + ((g1185) & (g1186) & (!g1207) & (!sk[113]) & (g1209) & (g1230)) + ((g1185) & (g1186) & (!g1207) & (sk[113]) & (!g1209) & (!g1230)) + ((g1185) & (g1186) & (!g1207) & (sk[113]) & (g1209) & (g1230)) + ((g1185) & (g1186) & (g1207) & (!sk[113]) & (!g1209) & (!g1230)) + ((g1185) & (g1186) & (g1207) & (!sk[113]) & (!g1209) & (g1230)) + ((g1185) & (g1186) & (g1207) & (!sk[113]) & (g1209) & (!g1230)) + ((g1185) & (g1186) & (g1207) & (!sk[113]) & (g1209) & (g1230)));
	assign sinx7x = (((!g1068) & (!g1232) & (!g1254) & (!sk[114]) & (g1255)) + ((!g1068) & (!g1232) & (g1254) & (!sk[114]) & (g1255)) + ((!g1068) & (!g1232) & (g1254) & (sk[114]) & (!g1255)) + ((!g1068) & (!g1232) & (g1254) & (sk[114]) & (g1255)) + ((!g1068) & (g1232) & (!g1254) & (!sk[114]) & (g1255)) + ((!g1068) & (g1232) & (!g1254) & (sk[114]) & (!g1255)) + ((!g1068) & (g1232) & (!g1254) & (sk[114]) & (g1255)) + ((!g1068) & (g1232) & (g1254) & (!sk[114]) & (g1255)) + ((g1068) & (!g1232) & (!g1254) & (!sk[114]) & (!g1255)) + ((g1068) & (!g1232) & (!g1254) & (!sk[114]) & (g1255)) + ((g1068) & (!g1232) & (!g1254) & (sk[114]) & (!g1255)) + ((g1068) & (!g1232) & (g1254) & (!sk[114]) & (!g1255)) + ((g1068) & (!g1232) & (g1254) & (!sk[114]) & (g1255)) + ((g1068) & (!g1232) & (g1254) & (sk[114]) & (g1255)) + ((g1068) & (g1232) & (!g1254) & (!sk[114]) & (!g1255)) + ((g1068) & (g1232) & (!g1254) & (!sk[114]) & (g1255)) + ((g1068) & (g1232) & (!g1254) & (sk[114]) & (g1255)) + ((g1068) & (g1232) & (g1254) & (!sk[114]) & (!g1255)) + ((g1068) & (g1232) & (g1254) & (!sk[114]) & (g1255)) + ((g1068) & (g1232) & (g1254) & (sk[114]) & (!g1255)));
	assign g1257 = (((!sk[115]) & (!g1234) & (g1235) & (!g1248)) + ((!sk[115]) & (!g1234) & (g1235) & (g1248)) + ((!sk[115]) & (g1234) & (g1235) & (!g1248)) + ((!sk[115]) & (g1234) & (g1235) & (g1248)) + ((sk[115]) & (!g1234) & (!g1235) & (g1248)) + ((sk[115]) & (!g1234) & (g1235) & (!g1248)) + ((sk[115]) & (g1234) & (!g1235) & (!g1248)) + ((sk[115]) & (g1234) & (g1235) & (!g1248)));
	assign g1258 = (((!g1209) & (!g1230) & (!g1233) & (!g1257) & (sk[116]) & (!g1252)) + ((!g1209) & (!g1230) & (!g1233) & (!g1257) & (sk[116]) & (g1252)) + ((!g1209) & (!g1230) & (!g1233) & (g1257) & (!sk[116]) & (!g1252)) + ((!g1209) & (!g1230) & (!g1233) & (g1257) & (!sk[116]) & (g1252)) + ((!g1209) & (!g1230) & (!g1233) & (g1257) & (sk[116]) & (g1252)) + ((!g1209) & (!g1230) & (g1233) & (!g1257) & (!sk[116]) & (!g1252)) + ((!g1209) & (!g1230) & (g1233) & (!g1257) & (!sk[116]) & (g1252)) + ((!g1209) & (!g1230) & (g1233) & (!g1257) & (sk[116]) & (g1252)) + ((!g1209) & (!g1230) & (g1233) & (g1257) & (!sk[116]) & (!g1252)) + ((!g1209) & (!g1230) & (g1233) & (g1257) & (!sk[116]) & (g1252)) + ((!g1209) & (g1230) & (!g1233) & (!g1257) & (!sk[116]) & (!g1252)) + ((!g1209) & (g1230) & (!g1233) & (!g1257) & (!sk[116]) & (g1252)) + ((!g1209) & (g1230) & (!g1233) & (!g1257) & (sk[116]) & (!g1252)) + ((!g1209) & (g1230) & (!g1233) & (!g1257) & (sk[116]) & (g1252)) + ((!g1209) & (g1230) & (!g1233) & (g1257) & (!sk[116]) & (!g1252)) + ((!g1209) & (g1230) & (!g1233) & (g1257) & (!sk[116]) & (g1252)) + ((!g1209) & (g1230) & (!g1233) & (g1257) & (sk[116]) & (g1252)) + ((!g1209) & (g1230) & (g1233) & (!g1257) & (!sk[116]) & (!g1252)) + ((!g1209) & (g1230) & (g1233) & (!g1257) & (!sk[116]) & (g1252)) + ((!g1209) & (g1230) & (g1233) & (!g1257) & (sk[116]) & (g1252)) + ((!g1209) & (g1230) & (g1233) & (g1257) & (!sk[116]) & (!g1252)) + ((!g1209) & (g1230) & (g1233) & (g1257) & (!sk[116]) & (g1252)) + ((g1209) & (!g1230) & (!g1233) & (!g1257) & (sk[116]) & (g1252)) + ((g1209) & (!g1230) & (!g1233) & (g1257) & (!sk[116]) & (!g1252)) + ((g1209) & (!g1230) & (!g1233) & (g1257) & (!sk[116]) & (g1252)) + ((g1209) & (!g1230) & (g1233) & (!g1257) & (!sk[116]) & (!g1252)) + ((g1209) & (!g1230) & (g1233) & (!g1257) & (!sk[116]) & (g1252)) + ((g1209) & (!g1230) & (g1233) & (!g1257) & (sk[116]) & (g1252)) + ((g1209) & (!g1230) & (g1233) & (g1257) & (!sk[116]) & (!g1252)) + ((g1209) & (!g1230) & (g1233) & (g1257) & (!sk[116]) & (g1252)) + ((g1209) & (g1230) & (!g1233) & (!g1257) & (!sk[116]) & (!g1252)) + ((g1209) & (g1230) & (!g1233) & (!g1257) & (!sk[116]) & (g1252)) + ((g1209) & (g1230) & (!g1233) & (!g1257) & (sk[116]) & (!g1252)) + ((g1209) & (g1230) & (!g1233) & (!g1257) & (sk[116]) & (g1252)) + ((g1209) & (g1230) & (!g1233) & (g1257) & (!sk[116]) & (!g1252)) + ((g1209) & (g1230) & (!g1233) & (g1257) & (!sk[116]) & (g1252)) + ((g1209) & (g1230) & (!g1233) & (g1257) & (sk[116]) & (g1252)) + ((g1209) & (g1230) & (g1233) & (!g1257) & (!sk[116]) & (!g1252)) + ((g1209) & (g1230) & (g1233) & (!g1257) & (!sk[116]) & (g1252)) + ((g1209) & (g1230) & (g1233) & (!g1257) & (sk[116]) & (g1252)) + ((g1209) & (g1230) & (g1233) & (g1257) & (!sk[116]) & (!g1252)) + ((g1209) & (g1230) & (g1233) & (g1257) & (!sk[116]) & (g1252)));
	assign g1259 = (((!g1215) & (!g1216) & (!g1223) & (!g1238) & (!g1240) & (g1246)) + ((!g1215) & (!g1216) & (!g1223) & (!g1238) & (g1240) & (!g1246)) + ((!g1215) & (!g1216) & (g1223) & (!g1238) & (!g1240) & (g1246)) + ((!g1215) & (!g1216) & (g1223) & (!g1238) & (g1240) & (!g1246)) + ((!g1215) & (g1216) & (!g1223) & (!g1238) & (!g1240) & (!g1246)) + ((!g1215) & (g1216) & (!g1223) & (!g1238) & (!g1240) & (g1246)) + ((!g1215) & (g1216) & (!g1223) & (!g1238) & (g1240) & (!g1246)) + ((!g1215) & (g1216) & (!g1223) & (!g1238) & (g1240) & (g1246)) + ((!g1215) & (g1216) & (!g1223) & (g1238) & (!g1240) & (g1246)) + ((!g1215) & (g1216) & (!g1223) & (g1238) & (g1240) & (!g1246)) + ((!g1215) & (g1216) & (g1223) & (!g1238) & (!g1240) & (g1246)) + ((!g1215) & (g1216) & (g1223) & (!g1238) & (g1240) & (!g1246)) + ((g1215) & (!g1216) & (!g1223) & (!g1238) & (!g1240) & (!g1246)) + ((g1215) & (!g1216) & (!g1223) & (!g1238) & (!g1240) & (g1246)) + ((g1215) & (!g1216) & (!g1223) & (!g1238) & (g1240) & (!g1246)) + ((g1215) & (!g1216) & (!g1223) & (!g1238) & (g1240) & (g1246)) + ((g1215) & (!g1216) & (!g1223) & (g1238) & (!g1240) & (g1246)) + ((g1215) & (!g1216) & (!g1223) & (g1238) & (g1240) & (!g1246)) + ((g1215) & (!g1216) & (g1223) & (!g1238) & (!g1240) & (g1246)) + ((g1215) & (!g1216) & (g1223) & (!g1238) & (g1240) & (!g1246)) + ((g1215) & (g1216) & (!g1223) & (!g1238) & (!g1240) & (!g1246)) + ((g1215) & (g1216) & (!g1223) & (!g1238) & (!g1240) & (g1246)) + ((g1215) & (g1216) & (!g1223) & (!g1238) & (g1240) & (!g1246)) + ((g1215) & (g1216) & (!g1223) & (!g1238) & (g1240) & (g1246)) + ((g1215) & (g1216) & (!g1223) & (g1238) & (!g1240) & (g1246)) + ((g1215) & (g1216) & (!g1223) & (g1238) & (g1240) & (!g1246)) + ((g1215) & (g1216) & (g1223) & (!g1238) & (!g1240) & (!g1246)) + ((g1215) & (g1216) & (g1223) & (!g1238) & (!g1240) & (g1246)) + ((g1215) & (g1216) & (g1223) & (!g1238) & (g1240) & (!g1246)) + ((g1215) & (g1216) & (g1223) & (!g1238) & (g1240) & (g1246)) + ((g1215) & (g1216) & (g1223) & (g1238) & (!g1240) & (g1246)) + ((g1215) & (g1216) & (g1223) & (g1238) & (g1240) & (!g1246)));
	assign g1260 = (((!g202) & (!g759) & (!sk[118]) & (!g972) & (g1241)) + ((!g202) & (!g759) & (!sk[118]) & (g972) & (g1241)) + ((!g202) & (!g759) & (sk[118]) & (!g972) & (g1241)) + ((!g202) & (!g759) & (sk[118]) & (g972) & (g1241)) + ((!g202) & (g759) & (!sk[118]) & (!g972) & (g1241)) + ((!g202) & (g759) & (!sk[118]) & (g972) & (g1241)) + ((!g202) & (g759) & (sk[118]) & (g972) & (g1241)) + ((g202) & (!g759) & (!sk[118]) & (!g972) & (!g1241)) + ((g202) & (!g759) & (!sk[118]) & (!g972) & (g1241)) + ((g202) & (!g759) & (!sk[118]) & (g972) & (!g1241)) + ((g202) & (!g759) & (!sk[118]) & (g972) & (g1241)) + ((g202) & (!g759) & (sk[118]) & (!g972) & (!g1241)) + ((g202) & (!g759) & (sk[118]) & (g972) & (!g1241)) + ((g202) & (g759) & (!sk[118]) & (!g972) & (!g1241)) + ((g202) & (g759) & (!sk[118]) & (!g972) & (g1241)) + ((g202) & (g759) & (!sk[118]) & (g972) & (!g1241)) + ((g202) & (g759) & (!sk[118]) & (g972) & (g1241)) + ((g202) & (g759) & (sk[118]) & (!g972) & (!g1241)) + ((g202) & (g759) & (sk[118]) & (!g972) & (g1241)) + ((g202) & (g759) & (sk[118]) & (g972) & (!g1241)));
	assign g1261 = (((!g764) & (!g762) & (!g765) & (!g962) & (!g971) & (!g994)) + ((!g764) & (!g762) & (!g765) & (!g962) & (!g971) & (g994)) + ((!g764) & (!g762) & (!g765) & (!g962) & (g971) & (!g994)) + ((!g764) & (!g762) & (!g765) & (!g962) & (g971) & (g994)) + ((!g764) & (!g762) & (!g765) & (g962) & (!g971) & (!g994)) + ((!g764) & (!g762) & (!g765) & (g962) & (!g971) & (g994)) + ((!g764) & (!g762) & (!g765) & (g962) & (g971) & (!g994)) + ((!g764) & (!g762) & (!g765) & (g962) & (g971) & (g994)) + ((!g764) & (!g762) & (g765) & (g962) & (!g971) & (!g994)) + ((!g764) & (!g762) & (g765) & (g962) & (!g971) & (g994)) + ((!g764) & (!g762) & (g765) & (g962) & (g971) & (!g994)) + ((!g764) & (!g762) & (g765) & (g962) & (g971) & (g994)) + ((!g764) & (g762) & (!g765) & (!g962) & (!g971) & (!g994)) + ((!g764) & (g762) & (!g765) & (!g962) & (!g971) & (g994)) + ((!g764) & (g762) & (!g765) & (g962) & (!g971) & (!g994)) + ((!g764) & (g762) & (!g765) & (g962) & (!g971) & (g994)) + ((!g764) & (g762) & (g765) & (g962) & (!g971) & (!g994)) + ((!g764) & (g762) & (g765) & (g962) & (!g971) & (g994)) + ((g764) & (!g762) & (!g765) & (!g962) & (!g971) & (!g994)) + ((g764) & (!g762) & (!g765) & (!g962) & (g971) & (!g994)) + ((g764) & (!g762) & (!g765) & (g962) & (!g971) & (!g994)) + ((g764) & (!g762) & (!g765) & (g962) & (g971) & (!g994)) + ((g764) & (!g762) & (g765) & (g962) & (!g971) & (!g994)) + ((g764) & (!g762) & (g765) & (g962) & (g971) & (!g994)) + ((g764) & (g762) & (!g765) & (!g962) & (!g971) & (!g994)) + ((g764) & (g762) & (!g765) & (g962) & (!g971) & (!g994)) + ((g764) & (g762) & (g765) & (g962) & (!g971) & (!g994)));
	assign g1262 = (((!g252) & (!g843) & (!g899) & (!g1242) & (g1243) & (!g1244)) + ((!g252) & (!g843) & (!g899) & (g1242) & (!g1243) & (!g1244)) + ((!g252) & (!g843) & (!g899) & (g1242) & (g1243) & (!g1244)) + ((!g252) & (!g843) & (!g899) & (g1242) & (g1243) & (g1244)) + ((!g252) & (!g843) & (g899) & (!g1242) & (g1243) & (!g1244)) + ((!g252) & (!g843) & (g899) & (g1242) & (!g1243) & (!g1244)) + ((!g252) & (!g843) & (g899) & (g1242) & (g1243) & (!g1244)) + ((!g252) & (!g843) & (g899) & (g1242) & (g1243) & (g1244)) + ((!g252) & (g843) & (!g899) & (!g1242) & (g1243) & (!g1244)) + ((!g252) & (g843) & (!g899) & (!g1242) & (g1243) & (g1244)) + ((!g252) & (g843) & (!g899) & (g1242) & (!g1243) & (!g1244)) + ((!g252) & (g843) & (!g899) & (g1242) & (!g1243) & (g1244)) + ((!g252) & (g843) & (!g899) & (g1242) & (g1243) & (!g1244)) + ((!g252) & (g843) & (!g899) & (g1242) & (g1243) & (g1244)) + ((!g252) & (g843) & (g899) & (!g1242) & (g1243) & (!g1244)) + ((!g252) & (g843) & (g899) & (g1242) & (!g1243) & (!g1244)) + ((!g252) & (g843) & (g899) & (g1242) & (g1243) & (!g1244)) + ((!g252) & (g843) & (g899) & (g1242) & (g1243) & (g1244)) + ((g252) & (!g843) & (!g899) & (!g1242) & (g1243) & (g1244)) + ((g252) & (!g843) & (!g899) & (g1242) & (!g1243) & (g1244)) + ((g252) & (!g843) & (!g899) & (g1242) & (g1243) & (!g1244)) + ((g252) & (!g843) & (!g899) & (g1242) & (g1243) & (g1244)) + ((g252) & (!g843) & (g899) & (!g1242) & (g1243) & (g1244)) + ((g252) & (!g843) & (g899) & (g1242) & (!g1243) & (g1244)) + ((g252) & (!g843) & (g899) & (g1242) & (g1243) & (!g1244)) + ((g252) & (!g843) & (g899) & (g1242) & (g1243) & (g1244)) + ((g252) & (g843) & (!g899) & (g1242) & (g1243) & (!g1244)) + ((g252) & (g843) & (!g899) & (g1242) & (g1243) & (g1244)) + ((g252) & (g843) & (g899) & (!g1242) & (g1243) & (g1244)) + ((g252) & (g843) & (g899) & (g1242) & (!g1243) & (g1244)) + ((g252) & (g843) & (g899) & (g1242) & (g1243) & (!g1244)) + ((g252) & (g843) & (g899) & (g1242) & (g1243) & (g1244)));
	assign g1263 = (((!sk[121]) & (!g2) & (!g252) & (!g683) & (g718)) + ((!sk[121]) & (!g2) & (!g252) & (g683) & (g718)) + ((!sk[121]) & (!g2) & (g252) & (!g683) & (g718)) + ((!sk[121]) & (!g2) & (g252) & (g683) & (g718)) + ((!sk[121]) & (g2) & (!g252) & (!g683) & (!g718)) + ((!sk[121]) & (g2) & (!g252) & (!g683) & (g718)) + ((!sk[121]) & (g2) & (!g252) & (g683) & (!g718)) + ((!sk[121]) & (g2) & (!g252) & (g683) & (g718)) + ((!sk[121]) & (g2) & (g252) & (!g683) & (!g718)) + ((!sk[121]) & (g2) & (g252) & (!g683) & (g718)) + ((!sk[121]) & (g2) & (g252) & (g683) & (!g718)) + ((!sk[121]) & (g2) & (g252) & (g683) & (g718)) + ((sk[121]) & (!g2) & (!g252) & (!g683) & (!g718)) + ((sk[121]) & (!g2) & (!g252) & (!g683) & (g718)) + ((sk[121]) & (!g2) & (g252) & (!g683) & (!g718)) + ((sk[121]) & (!g2) & (g252) & (!g683) & (g718)) + ((sk[121]) & (!g2) & (g252) & (g683) & (g718)) + ((sk[121]) & (g2) & (g252) & (!g683) & (g718)));
	assign g1264 = (((!g698) & (!g706) & (!g717) & (!g825) & (!g832) & (g848)) + ((!g698) & (!g706) & (!g717) & (g825) & (g832) & (g848)) + ((!g698) & (!g706) & (g717) & (!g825) & (!g832) & (g848)) + ((!g698) & (!g706) & (g717) & (g825) & (g832) & (g848)) + ((!g698) & (g706) & (!g717) & (!g825) & (!g832) & (g848)) + ((!g698) & (g706) & (!g717) & (g825) & (g832) & (g848)) + ((!g698) & (g706) & (g717) & (!g825) & (g832) & (g848)) + ((!g698) & (g706) & (g717) & (g825) & (!g832) & (g848)) + ((g698) & (!g706) & (!g717) & (!g825) & (!g832) & (g848)) + ((g698) & (!g706) & (!g717) & (g825) & (g832) & (g848)) + ((g698) & (!g706) & (g717) & (!g825) & (g832) & (g848)) + ((g698) & (!g706) & (g717) & (g825) & (!g832) & (g848)) + ((g698) & (g706) & (!g717) & (!g825) & (g832) & (g848)) + ((g698) & (g706) & (!g717) & (g825) & (!g832) & (g848)) + ((g698) & (g706) & (g717) & (!g825) & (g832) & (g848)) + ((g698) & (g706) & (g717) & (g825) & (!g832) & (g848)));
	assign g1265 = (((!g847) & (!g845) & (!g871) & (!g883) & (!g863) & (!g1264)) + ((!g847) & (!g845) & (!g871) & (!g883) & (g863) & (!g1264)) + ((!g847) & (!g845) & (!g871) & (g883) & (!g863) & (!g1264)) + ((!g847) & (!g845) & (!g871) & (g883) & (g863) & (!g1264)) + ((!g847) & (!g845) & (g871) & (!g883) & (!g863) & (!g1264)) + ((!g847) & (!g845) & (g871) & (!g883) & (g863) & (!g1264)) + ((!g847) & (!g845) & (g871) & (g883) & (!g863) & (!g1264)) + ((!g847) & (!g845) & (g871) & (g883) & (g863) & (!g1264)) + ((!g847) & (g845) & (!g871) & (!g883) & (!g863) & (!g1264)) + ((!g847) & (g845) & (!g871) & (g883) & (!g863) & (!g1264)) + ((!g847) & (g845) & (g871) & (!g883) & (!g863) & (!g1264)) + ((!g847) & (g845) & (g871) & (g883) & (!g863) & (!g1264)) + ((g847) & (!g845) & (!g871) & (g883) & (!g863) & (!g1264)) + ((g847) & (!g845) & (!g871) & (g883) & (g863) & (!g1264)) + ((g847) & (!g845) & (g871) & (!g883) & (!g863) & (!g1264)) + ((g847) & (!g845) & (g871) & (!g883) & (g863) & (!g1264)) + ((g847) & (g845) & (!g871) & (g883) & (!g863) & (!g1264)) + ((g847) & (g845) & (g871) & (!g883) & (!g863) & (!g1264)));
	assign g1266 = (((!g252) & (!g869) & (!g843) & (!g895) & (!g1263) & (!g1265)) + ((!g252) & (!g869) & (!g843) & (!g895) & (g1263) & (g1265)) + ((!g252) & (!g869) & (!g843) & (g895) & (!g1263) & (!g1265)) + ((!g252) & (!g869) & (!g843) & (g895) & (g1263) & (g1265)) + ((!g252) & (!g869) & (g843) & (!g895) & (!g1263) & (!g1265)) + ((!g252) & (!g869) & (g843) & (!g895) & (g1263) & (g1265)) + ((!g252) & (!g869) & (g843) & (g895) & (!g1263) & (!g1265)) + ((!g252) & (!g869) & (g843) & (g895) & (!g1263) & (g1265)) + ((!g252) & (g869) & (!g843) & (!g895) & (!g1263) & (!g1265)) + ((!g252) & (g869) & (!g843) & (!g895) & (g1263) & (g1265)) + ((!g252) & (g869) & (!g843) & (g895) & (!g1263) & (!g1265)) + ((!g252) & (g869) & (!g843) & (g895) & (g1263) & (g1265)) + ((!g252) & (g869) & (g843) & (!g895) & (!g1263) & (!g1265)) + ((!g252) & (g869) & (g843) & (!g895) & (g1263) & (g1265)) + ((!g252) & (g869) & (g843) & (g895) & (!g1263) & (!g1265)) + ((!g252) & (g869) & (g843) & (g895) & (!g1263) & (g1265)) + ((g252) & (!g869) & (!g843) & (!g895) & (!g1263) & (g1265)) + ((g252) & (!g869) & (!g843) & (!g895) & (g1263) & (!g1265)) + ((g252) & (!g869) & (!g843) & (g895) & (!g1263) & (g1265)) + ((g252) & (!g869) & (!g843) & (g895) & (g1263) & (!g1265)) + ((g252) & (!g869) & (g843) & (!g895) & (!g1263) & (g1265)) + ((g252) & (!g869) & (g843) & (!g895) & (g1263) & (!g1265)) + ((g252) & (!g869) & (g843) & (g895) & (g1263) & (!g1265)) + ((g252) & (!g869) & (g843) & (g895) & (g1263) & (g1265)) + ((g252) & (g869) & (!g843) & (!g895) & (!g1263) & (!g1265)) + ((g252) & (g869) & (!g843) & (!g895) & (g1263) & (g1265)) + ((g252) & (g869) & (!g843) & (g895) & (!g1263) & (!g1265)) + ((g252) & (g869) & (!g843) & (g895) & (g1263) & (g1265)) + ((g252) & (g869) & (g843) & (!g895) & (!g1263) & (!g1265)) + ((g252) & (g869) & (g843) & (!g895) & (g1263) & (g1265)) + ((g252) & (g869) & (g843) & (g895) & (!g1263) & (!g1265)) + ((g252) & (g869) & (g843) & (g895) & (!g1263) & (g1265)));
	assign g1267 = (((!g202) & (!g759) & (!g995) & (!g1261) & (!g1262) & (!g1266)) + ((!g202) & (!g759) & (!g995) & (!g1261) & (g1262) & (g1266)) + ((!g202) & (!g759) & (!g995) & (g1261) & (!g1262) & (g1266)) + ((!g202) & (!g759) & (!g995) & (g1261) & (g1262) & (!g1266)) + ((!g202) & (!g759) & (g995) & (!g1261) & (!g1262) & (!g1266)) + ((!g202) & (!g759) & (g995) & (!g1261) & (g1262) & (g1266)) + ((!g202) & (!g759) & (g995) & (g1261) & (!g1262) & (g1266)) + ((!g202) & (!g759) & (g995) & (g1261) & (g1262) & (!g1266)) + ((!g202) & (g759) & (!g995) & (!g1261) & (!g1262) & (!g1266)) + ((!g202) & (g759) & (!g995) & (!g1261) & (g1262) & (g1266)) + ((!g202) & (g759) & (!g995) & (g1261) & (!g1262) & (g1266)) + ((!g202) & (g759) & (!g995) & (g1261) & (g1262) & (!g1266)) + ((!g202) & (g759) & (g995) & (!g1261) & (!g1262) & (!g1266)) + ((!g202) & (g759) & (g995) & (!g1261) & (g1262) & (g1266)) + ((!g202) & (g759) & (g995) & (g1261) & (!g1262) & (!g1266)) + ((!g202) & (g759) & (g995) & (g1261) & (g1262) & (g1266)) + ((g202) & (!g759) & (!g995) & (!g1261) & (!g1262) & (g1266)) + ((g202) & (!g759) & (!g995) & (!g1261) & (g1262) & (!g1266)) + ((g202) & (!g759) & (!g995) & (g1261) & (!g1262) & (!g1266)) + ((g202) & (!g759) & (!g995) & (g1261) & (g1262) & (g1266)) + ((g202) & (!g759) & (g995) & (!g1261) & (!g1262) & (g1266)) + ((g202) & (!g759) & (g995) & (!g1261) & (g1262) & (!g1266)) + ((g202) & (!g759) & (g995) & (g1261) & (!g1262) & (!g1266)) + ((g202) & (!g759) & (g995) & (g1261) & (g1262) & (g1266)) + ((g202) & (g759) & (!g995) & (!g1261) & (!g1262) & (g1266)) + ((g202) & (g759) & (!g995) & (!g1261) & (g1262) & (!g1266)) + ((g202) & (g759) & (!g995) & (g1261) & (!g1262) & (!g1266)) + ((g202) & (g759) & (!g995) & (g1261) & (g1262) & (g1266)) + ((g202) & (g759) & (g995) & (!g1261) & (!g1262) & (g1266)) + ((g202) & (g759) & (g995) & (!g1261) & (g1262) & (!g1266)) + ((g202) & (g759) & (g995) & (g1261) & (!g1262) & (g1266)) + ((g202) & (g759) & (g995) & (g1261) & (g1262) & (!g1266)));
	assign g1268 = (((!sk[126]) & (!g744) & (!g748) & (!g1040) & (g1079)) + ((!sk[126]) & (!g744) & (!g748) & (g1040) & (g1079)) + ((!sk[126]) & (!g744) & (g748) & (!g1040) & (g1079)) + ((!sk[126]) & (!g744) & (g748) & (g1040) & (g1079)) + ((!sk[126]) & (g744) & (!g748) & (!g1040) & (!g1079)) + ((!sk[126]) & (g744) & (!g748) & (!g1040) & (g1079)) + ((!sk[126]) & (g744) & (!g748) & (g1040) & (!g1079)) + ((!sk[126]) & (g744) & (!g748) & (g1040) & (g1079)) + ((!sk[126]) & (g744) & (g748) & (!g1040) & (!g1079)) + ((!sk[126]) & (g744) & (g748) & (!g1040) & (g1079)) + ((!sk[126]) & (g744) & (g748) & (g1040) & (!g1079)) + ((!sk[126]) & (g744) & (g748) & (g1040) & (g1079)) + ((sk[126]) & (!g744) & (g748) & (!g1040) & (!g1079)) + ((sk[126]) & (!g744) & (g748) & (!g1040) & (g1079)) + ((sk[126]) & (g744) & (!g748) & (!g1040) & (!g1079)) + ((sk[126]) & (g744) & (!g748) & (g1040) & (!g1079)) + ((sk[126]) & (g744) & (g748) & (!g1040) & (!g1079)) + ((sk[126]) & (g744) & (g748) & (!g1040) & (g1079)) + ((sk[126]) & (g744) & (g748) & (g1040) & (!g1079)));
	assign g1269 = (((!g200) & (!g742) & (!g1040) & (!g1079) & (!g1080) & (g1268)) + ((!g200) & (!g742) & (!g1040) & (!g1079) & (g1080) & (g1268)) + ((!g200) & (!g742) & (!g1040) & (g1079) & (!g1080) & (g1268)) + ((!g200) & (!g742) & (!g1040) & (g1079) & (g1080) & (g1268)) + ((!g200) & (!g742) & (g1040) & (!g1079) & (!g1080) & (g1268)) + ((!g200) & (!g742) & (g1040) & (!g1079) & (g1080) & (g1268)) + ((!g200) & (!g742) & (g1040) & (g1079) & (!g1080) & (g1268)) + ((!g200) & (!g742) & (g1040) & (g1079) & (g1080) & (g1268)) + ((!g200) & (g742) & (!g1040) & (!g1079) & (!g1080) & (g1268)) + ((!g200) & (g742) & (!g1040) & (!g1079) & (g1080) & (g1268)) + ((!g200) & (g742) & (!g1040) & (g1079) & (!g1080) & (g1268)) + ((!g200) & (g742) & (!g1040) & (g1079) & (g1080) & (!g1268)) + ((!g200) & (g742) & (!g1040) & (g1079) & (g1080) & (g1268)) + ((!g200) & (g742) & (g1040) & (!g1079) & (!g1080) & (!g1268)) + ((!g200) & (g742) & (g1040) & (!g1079) & (!g1080) & (g1268)) + ((!g200) & (g742) & (g1040) & (!g1079) & (g1080) & (g1268)) + ((!g200) & (g742) & (g1040) & (g1079) & (!g1080) & (g1268)) + ((!g200) & (g742) & (g1040) & (g1079) & (g1080) & (g1268)) + ((g200) & (!g742) & (!g1040) & (!g1079) & (!g1080) & (!g1268)) + ((g200) & (!g742) & (!g1040) & (!g1079) & (g1080) & (!g1268)) + ((g200) & (!g742) & (!g1040) & (g1079) & (!g1080) & (!g1268)) + ((g200) & (!g742) & (!g1040) & (g1079) & (g1080) & (!g1268)) + ((g200) & (!g742) & (g1040) & (!g1079) & (!g1080) & (!g1268)) + ((g200) & (!g742) & (g1040) & (!g1079) & (g1080) & (!g1268)) + ((g200) & (!g742) & (g1040) & (g1079) & (!g1080) & (!g1268)) + ((g200) & (!g742) & (g1040) & (g1079) & (g1080) & (!g1268)) + ((g200) & (g742) & (!g1040) & (!g1079) & (!g1080) & (!g1268)) + ((g200) & (g742) & (!g1040) & (!g1079) & (g1080) & (!g1268)) + ((g200) & (g742) & (!g1040) & (g1079) & (!g1080) & (!g1268)) + ((g200) & (g742) & (g1040) & (!g1079) & (g1080) & (!g1268)) + ((g200) & (g742) & (g1040) & (g1079) & (!g1080) & (!g1268)) + ((g200) & (g742) & (g1040) & (g1079) & (g1080) & (!g1268)));
	assign g1270 = (((!g1240) & (!sk[0]) & (!g1260) & (!g1245) & (g1267) & (!g1269)) + ((!g1240) & (!sk[0]) & (!g1260) & (!g1245) & (g1267) & (g1269)) + ((!g1240) & (!sk[0]) & (!g1260) & (g1245) & (!g1267) & (!g1269)) + ((!g1240) & (!sk[0]) & (!g1260) & (g1245) & (!g1267) & (g1269)) + ((!g1240) & (!sk[0]) & (!g1260) & (g1245) & (g1267) & (!g1269)) + ((!g1240) & (!sk[0]) & (!g1260) & (g1245) & (g1267) & (g1269)) + ((!g1240) & (!sk[0]) & (g1260) & (!g1245) & (!g1267) & (!g1269)) + ((!g1240) & (!sk[0]) & (g1260) & (!g1245) & (!g1267) & (g1269)) + ((!g1240) & (!sk[0]) & (g1260) & (!g1245) & (g1267) & (!g1269)) + ((!g1240) & (!sk[0]) & (g1260) & (!g1245) & (g1267) & (g1269)) + ((!g1240) & (!sk[0]) & (g1260) & (g1245) & (!g1267) & (!g1269)) + ((!g1240) & (!sk[0]) & (g1260) & (g1245) & (!g1267) & (g1269)) + ((!g1240) & (!sk[0]) & (g1260) & (g1245) & (g1267) & (!g1269)) + ((!g1240) & (!sk[0]) & (g1260) & (g1245) & (g1267) & (g1269)) + ((!g1240) & (sk[0]) & (!g1260) & (!g1245) & (!g1267) & (!g1269)) + ((!g1240) & (sk[0]) & (!g1260) & (!g1245) & (g1267) & (g1269)) + ((!g1240) & (sk[0]) & (!g1260) & (g1245) & (!g1267) & (!g1269)) + ((!g1240) & (sk[0]) & (!g1260) & (g1245) & (g1267) & (g1269)) + ((!g1240) & (sk[0]) & (g1260) & (!g1245) & (!g1267) & (g1269)) + ((!g1240) & (sk[0]) & (g1260) & (!g1245) & (g1267) & (!g1269)) + ((!g1240) & (sk[0]) & (g1260) & (g1245) & (!g1267) & (!g1269)) + ((!g1240) & (sk[0]) & (g1260) & (g1245) & (g1267) & (g1269)) + ((g1240) & (!sk[0]) & (!g1260) & (!g1245) & (g1267) & (!g1269)) + ((g1240) & (!sk[0]) & (!g1260) & (!g1245) & (g1267) & (g1269)) + ((g1240) & (!sk[0]) & (!g1260) & (g1245) & (!g1267) & (!g1269)) + ((g1240) & (!sk[0]) & (!g1260) & (g1245) & (!g1267) & (g1269)) + ((g1240) & (!sk[0]) & (!g1260) & (g1245) & (g1267) & (!g1269)) + ((g1240) & (!sk[0]) & (!g1260) & (g1245) & (g1267) & (g1269)) + ((g1240) & (!sk[0]) & (g1260) & (!g1245) & (!g1267) & (!g1269)) + ((g1240) & (!sk[0]) & (g1260) & (!g1245) & (!g1267) & (g1269)) + ((g1240) & (!sk[0]) & (g1260) & (!g1245) & (g1267) & (!g1269)) + ((g1240) & (!sk[0]) & (g1260) & (!g1245) & (g1267) & (g1269)) + ((g1240) & (!sk[0]) & (g1260) & (g1245) & (!g1267) & (!g1269)) + ((g1240) & (!sk[0]) & (g1260) & (g1245) & (!g1267) & (g1269)) + ((g1240) & (!sk[0]) & (g1260) & (g1245) & (g1267) & (!g1269)) + ((g1240) & (!sk[0]) & (g1260) & (g1245) & (g1267) & (g1269)) + ((g1240) & (sk[0]) & (!g1260) & (!g1245) & (!g1267) & (g1269)) + ((g1240) & (sk[0]) & (!g1260) & (!g1245) & (g1267) & (!g1269)) + ((g1240) & (sk[0]) & (!g1260) & (g1245) & (!g1267) & (!g1269)) + ((g1240) & (sk[0]) & (!g1260) & (g1245) & (g1267) & (g1269)) + ((g1240) & (sk[0]) & (g1260) & (!g1245) & (!g1267) & (g1269)) + ((g1240) & (sk[0]) & (g1260) & (!g1245) & (g1267) & (!g1269)) + ((g1240) & (sk[0]) & (g1260) & (g1245) & (!g1267) & (g1269)) + ((g1240) & (sk[0]) & (g1260) & (g1245) & (g1267) & (!g1269)));
	assign g1271 = (((!g1259) & (sk[1]) & (g1270)) + ((g1259) & (!sk[1]) & (g1270)) + ((g1259) & (sk[1]) & (!g1270)));
	assign g1272 = (((!g114) & (g115) & (!g8) & (!g40) & (g25) & (!g149)) + ((!g114) & (g115) & (!g8) & (!g40) & (g25) & (g149)) + ((!g114) & (g115) & (!g8) & (g40) & (g25) & (!g149)) + ((!g114) & (g115) & (!g8) & (g40) & (g25) & (g149)) + ((!g114) & (g115) & (g8) & (!g40) & (g25) & (!g149)) + ((!g114) & (g115) & (g8) & (!g40) & (g25) & (g149)) + ((!g114) & (g115) & (g8) & (g40) & (g25) & (!g149)) + ((!g114) & (g115) & (g8) & (g40) & (g25) & (g149)) + ((g114) & (g115) & (!g8) & (g40) & (!g25) & (!g149)) + ((g114) & (g115) & (!g8) & (g40) & (!g25) & (g149)) + ((g114) & (g115) & (!g8) & (g40) & (g25) & (!g149)) + ((g114) & (g115) & (!g8) & (g40) & (g25) & (g149)) + ((g114) & (g115) & (g8) & (!g40) & (!g25) & (g149)) + ((g114) & (g115) & (g8) & (!g40) & (g25) & (g149)) + ((g114) & (g115) & (g8) & (g40) & (!g25) & (!g149)) + ((g114) & (g115) & (g8) & (g40) & (!g25) & (g149)) + ((g114) & (g115) & (g8) & (g40) & (g25) & (!g149)) + ((g114) & (g115) & (g8) & (g40) & (g25) & (g149)));
	assign g1273 = (((!g550) & (!g291) & (!g228) & (!sk[3]) & (g229) & (!g1272)) + ((!g550) & (!g291) & (!g228) & (!sk[3]) & (g229) & (g1272)) + ((!g550) & (!g291) & (g228) & (!sk[3]) & (!g229) & (!g1272)) + ((!g550) & (!g291) & (g228) & (!sk[3]) & (!g229) & (g1272)) + ((!g550) & (!g291) & (g228) & (!sk[3]) & (g229) & (!g1272)) + ((!g550) & (!g291) & (g228) & (!sk[3]) & (g229) & (g1272)) + ((!g550) & (g291) & (!g228) & (!sk[3]) & (!g229) & (!g1272)) + ((!g550) & (g291) & (!g228) & (!sk[3]) & (!g229) & (g1272)) + ((!g550) & (g291) & (!g228) & (!sk[3]) & (g229) & (!g1272)) + ((!g550) & (g291) & (!g228) & (!sk[3]) & (g229) & (g1272)) + ((!g550) & (g291) & (g228) & (!sk[3]) & (!g229) & (!g1272)) + ((!g550) & (g291) & (g228) & (!sk[3]) & (!g229) & (g1272)) + ((!g550) & (g291) & (g228) & (!sk[3]) & (g229) & (!g1272)) + ((!g550) & (g291) & (g228) & (!sk[3]) & (g229) & (g1272)) + ((g550) & (!g291) & (!g228) & (!sk[3]) & (g229) & (!g1272)) + ((g550) & (!g291) & (!g228) & (!sk[3]) & (g229) & (g1272)) + ((g550) & (!g291) & (g228) & (!sk[3]) & (!g229) & (!g1272)) + ((g550) & (!g291) & (g228) & (!sk[3]) & (!g229) & (g1272)) + ((g550) & (!g291) & (g228) & (!sk[3]) & (g229) & (!g1272)) + ((g550) & (!g291) & (g228) & (!sk[3]) & (g229) & (g1272)) + ((g550) & (g291) & (!g228) & (!sk[3]) & (!g229) & (!g1272)) + ((g550) & (g291) & (!g228) & (!sk[3]) & (!g229) & (g1272)) + ((g550) & (g291) & (!g228) & (!sk[3]) & (g229) & (!g1272)) + ((g550) & (g291) & (!g228) & (!sk[3]) & (g229) & (g1272)) + ((g550) & (g291) & (g228) & (!sk[3]) & (!g229) & (!g1272)) + ((g550) & (g291) & (g228) & (!sk[3]) & (!g229) & (g1272)) + ((g550) & (g291) & (g228) & (!sk[3]) & (g229) & (!g1272)) + ((g550) & (g291) & (g228) & (!sk[3]) & (g229) & (g1272)) + ((g550) & (g291) & (g228) & (sk[3]) & (g229) & (!g1272)));
	assign g1274 = (((!g153) & (!g146) & (!g74) & (!sk[4]) & (g152)) + ((!g153) & (!g146) & (!g74) & (sk[4]) & (!g152)) + ((!g153) & (!g146) & (g74) & (!sk[4]) & (g152)) + ((!g153) & (g146) & (!g74) & (!sk[4]) & (g152)) + ((!g153) & (g146) & (g74) & (!sk[4]) & (g152)) + ((g153) & (!g146) & (!g74) & (!sk[4]) & (!g152)) + ((g153) & (!g146) & (!g74) & (!sk[4]) & (g152)) + ((g153) & (!g146) & (g74) & (!sk[4]) & (!g152)) + ((g153) & (!g146) & (g74) & (!sk[4]) & (g152)) + ((g153) & (g146) & (!g74) & (!sk[4]) & (!g152)) + ((g153) & (g146) & (!g74) & (!sk[4]) & (g152)) + ((g153) & (g146) & (g74) & (!sk[4]) & (!g152)) + ((g153) & (g146) & (g74) & (!sk[4]) & (g152)));
	assign g1275 = (((!sk[5]) & (!g38) & (!g71) & (!g58) & (g104) & (!g32)) + ((!sk[5]) & (!g38) & (!g71) & (!g58) & (g104) & (g32)) + ((!sk[5]) & (!g38) & (!g71) & (g58) & (!g104) & (!g32)) + ((!sk[5]) & (!g38) & (!g71) & (g58) & (!g104) & (g32)) + ((!sk[5]) & (!g38) & (!g71) & (g58) & (g104) & (!g32)) + ((!sk[5]) & (!g38) & (!g71) & (g58) & (g104) & (g32)) + ((!sk[5]) & (!g38) & (g71) & (!g58) & (!g104) & (!g32)) + ((!sk[5]) & (!g38) & (g71) & (!g58) & (!g104) & (g32)) + ((!sk[5]) & (!g38) & (g71) & (!g58) & (g104) & (!g32)) + ((!sk[5]) & (!g38) & (g71) & (!g58) & (g104) & (g32)) + ((!sk[5]) & (!g38) & (g71) & (g58) & (!g104) & (!g32)) + ((!sk[5]) & (!g38) & (g71) & (g58) & (!g104) & (g32)) + ((!sk[5]) & (!g38) & (g71) & (g58) & (g104) & (!g32)) + ((!sk[5]) & (!g38) & (g71) & (g58) & (g104) & (g32)) + ((!sk[5]) & (g38) & (!g71) & (!g58) & (g104) & (!g32)) + ((!sk[5]) & (g38) & (!g71) & (!g58) & (g104) & (g32)) + ((!sk[5]) & (g38) & (!g71) & (g58) & (!g104) & (!g32)) + ((!sk[5]) & (g38) & (!g71) & (g58) & (!g104) & (g32)) + ((!sk[5]) & (g38) & (!g71) & (g58) & (g104) & (!g32)) + ((!sk[5]) & (g38) & (!g71) & (g58) & (g104) & (g32)) + ((!sk[5]) & (g38) & (g71) & (!g58) & (!g104) & (!g32)) + ((!sk[5]) & (g38) & (g71) & (!g58) & (!g104) & (g32)) + ((!sk[5]) & (g38) & (g71) & (!g58) & (g104) & (!g32)) + ((!sk[5]) & (g38) & (g71) & (!g58) & (g104) & (g32)) + ((!sk[5]) & (g38) & (g71) & (g58) & (!g104) & (!g32)) + ((!sk[5]) & (g38) & (g71) & (g58) & (!g104) & (g32)) + ((!sk[5]) & (g38) & (g71) & (g58) & (g104) & (!g32)) + ((!sk[5]) & (g38) & (g71) & (g58) & (g104) & (g32)) + ((sk[5]) & (!g38) & (!g71) & (!g58) & (!g104) & (!g32)) + ((sk[5]) & (!g38) & (!g71) & (!g58) & (!g104) & (g32)) + ((sk[5]) & (!g38) & (!g71) & (!g58) & (g104) & (!g32)) + ((sk[5]) & (!g38) & (!g71) & (!g58) & (g104) & (g32)) + ((sk[5]) & (!g38) & (!g71) & (g58) & (!g104) & (!g32)) + ((sk[5]) & (!g38) & (!g71) & (g58) & (!g104) & (g32)) + ((sk[5]) & (!g38) & (g71) & (!g58) & (!g104) & (!g32)) + ((sk[5]) & (!g38) & (g71) & (!g58) & (g104) & (!g32)) + ((sk[5]) & (g38) & (!g71) & (!g58) & (!g104) & (!g32)) + ((sk[5]) & (g38) & (!g71) & (!g58) & (!g104) & (g32)) + ((sk[5]) & (g38) & (!g71) & (g58) & (!g104) & (!g32)) + ((sk[5]) & (g38) & (!g71) & (g58) & (!g104) & (g32)) + ((sk[5]) & (g38) & (g71) & (!g58) & (!g104) & (!g32)));
	assign g1276 = (((!sk[6]) & (!g9) & (!g62) & (!g18) & (g1275)) + ((!sk[6]) & (!g9) & (!g62) & (g18) & (g1275)) + ((!sk[6]) & (!g9) & (g62) & (!g18) & (g1275)) + ((!sk[6]) & (!g9) & (g62) & (g18) & (g1275)) + ((!sk[6]) & (g9) & (!g62) & (!g18) & (!g1275)) + ((!sk[6]) & (g9) & (!g62) & (!g18) & (g1275)) + ((!sk[6]) & (g9) & (!g62) & (g18) & (!g1275)) + ((!sk[6]) & (g9) & (!g62) & (g18) & (g1275)) + ((!sk[6]) & (g9) & (g62) & (!g18) & (!g1275)) + ((!sk[6]) & (g9) & (g62) & (!g18) & (g1275)) + ((!sk[6]) & (g9) & (g62) & (g18) & (!g1275)) + ((!sk[6]) & (g9) & (g62) & (g18) & (g1275)) + ((sk[6]) & (!g9) & (!g62) & (!g18) & (g1275)) + ((sk[6]) & (!g9) & (!g62) & (g18) & (g1275)) + ((sk[6]) & (!g9) & (g62) & (!g18) & (g1275)) + ((sk[6]) & (g9) & (!g62) & (!g18) & (g1275)) + ((sk[6]) & (g9) & (g62) & (!g18) & (g1275)));
	assign g1277 = (((!g47) & (!g93) & (!g80) & (g1274) & (!sk[7]) & (!g1276)) + ((!g47) & (!g93) & (!g80) & (g1274) & (!sk[7]) & (g1276)) + ((!g47) & (!g93) & (!g80) & (g1274) & (sk[7]) & (g1276)) + ((!g47) & (!g93) & (g80) & (!g1274) & (!sk[7]) & (!g1276)) + ((!g47) & (!g93) & (g80) & (!g1274) & (!sk[7]) & (g1276)) + ((!g47) & (!g93) & (g80) & (g1274) & (!sk[7]) & (!g1276)) + ((!g47) & (!g93) & (g80) & (g1274) & (!sk[7]) & (g1276)) + ((!g47) & (g93) & (!g80) & (!g1274) & (!sk[7]) & (!g1276)) + ((!g47) & (g93) & (!g80) & (!g1274) & (!sk[7]) & (g1276)) + ((!g47) & (g93) & (!g80) & (g1274) & (!sk[7]) & (!g1276)) + ((!g47) & (g93) & (!g80) & (g1274) & (!sk[7]) & (g1276)) + ((!g47) & (g93) & (g80) & (!g1274) & (!sk[7]) & (!g1276)) + ((!g47) & (g93) & (g80) & (!g1274) & (!sk[7]) & (g1276)) + ((!g47) & (g93) & (g80) & (g1274) & (!sk[7]) & (!g1276)) + ((!g47) & (g93) & (g80) & (g1274) & (!sk[7]) & (g1276)) + ((g47) & (!g93) & (!g80) & (g1274) & (!sk[7]) & (!g1276)) + ((g47) & (!g93) & (!g80) & (g1274) & (!sk[7]) & (g1276)) + ((g47) & (!g93) & (g80) & (!g1274) & (!sk[7]) & (!g1276)) + ((g47) & (!g93) & (g80) & (!g1274) & (!sk[7]) & (g1276)) + ((g47) & (!g93) & (g80) & (g1274) & (!sk[7]) & (!g1276)) + ((g47) & (!g93) & (g80) & (g1274) & (!sk[7]) & (g1276)) + ((g47) & (g93) & (!g80) & (!g1274) & (!sk[7]) & (!g1276)) + ((g47) & (g93) & (!g80) & (!g1274) & (!sk[7]) & (g1276)) + ((g47) & (g93) & (!g80) & (g1274) & (!sk[7]) & (!g1276)) + ((g47) & (g93) & (!g80) & (g1274) & (!sk[7]) & (g1276)) + ((g47) & (g93) & (g80) & (!g1274) & (!sk[7]) & (!g1276)) + ((g47) & (g93) & (g80) & (!g1274) & (!sk[7]) & (g1276)) + ((g47) & (g93) & (g80) & (g1274) & (!sk[7]) & (!g1276)) + ((g47) & (g93) & (g80) & (g1274) & (!sk[7]) & (g1276)));
	assign g1278 = (((!g297) & (!g602) & (!g1015) & (g1273) & (!sk[8]) & (!g1277)) + ((!g297) & (!g602) & (!g1015) & (g1273) & (!sk[8]) & (g1277)) + ((!g297) & (!g602) & (g1015) & (!g1273) & (!sk[8]) & (!g1277)) + ((!g297) & (!g602) & (g1015) & (!g1273) & (!sk[8]) & (g1277)) + ((!g297) & (!g602) & (g1015) & (g1273) & (!sk[8]) & (!g1277)) + ((!g297) & (!g602) & (g1015) & (g1273) & (!sk[8]) & (g1277)) + ((!g297) & (g602) & (!g1015) & (!g1273) & (!sk[8]) & (!g1277)) + ((!g297) & (g602) & (!g1015) & (!g1273) & (!sk[8]) & (g1277)) + ((!g297) & (g602) & (!g1015) & (g1273) & (!sk[8]) & (!g1277)) + ((!g297) & (g602) & (!g1015) & (g1273) & (!sk[8]) & (g1277)) + ((!g297) & (g602) & (g1015) & (!g1273) & (!sk[8]) & (!g1277)) + ((!g297) & (g602) & (g1015) & (!g1273) & (!sk[8]) & (g1277)) + ((!g297) & (g602) & (g1015) & (g1273) & (!sk[8]) & (!g1277)) + ((!g297) & (g602) & (g1015) & (g1273) & (!sk[8]) & (g1277)) + ((!g297) & (g602) & (g1015) & (g1273) & (sk[8]) & (g1277)) + ((g297) & (!g602) & (!g1015) & (g1273) & (!sk[8]) & (!g1277)) + ((g297) & (!g602) & (!g1015) & (g1273) & (!sk[8]) & (g1277)) + ((g297) & (!g602) & (g1015) & (!g1273) & (!sk[8]) & (!g1277)) + ((g297) & (!g602) & (g1015) & (!g1273) & (!sk[8]) & (g1277)) + ((g297) & (!g602) & (g1015) & (g1273) & (!sk[8]) & (!g1277)) + ((g297) & (!g602) & (g1015) & (g1273) & (!sk[8]) & (g1277)) + ((g297) & (g602) & (!g1015) & (!g1273) & (!sk[8]) & (!g1277)) + ((g297) & (g602) & (!g1015) & (!g1273) & (!sk[8]) & (g1277)) + ((g297) & (g602) & (!g1015) & (g1273) & (!sk[8]) & (!g1277)) + ((g297) & (g602) & (!g1015) & (g1273) & (!sk[8]) & (g1277)) + ((g297) & (g602) & (g1015) & (!g1273) & (!sk[8]) & (!g1277)) + ((g297) & (g602) & (g1015) & (!g1273) & (!sk[8]) & (g1277)) + ((g297) & (g602) & (g1015) & (g1273) & (!sk[8]) & (!g1277)) + ((g297) & (g602) & (g1015) & (g1273) & (!sk[8]) & (g1277)));
	assign g1279 = (((!g1234) & (!g1235) & (!g1236) & (!g1247) & (!g1271) & (!g1278)) + ((!g1234) & (!g1235) & (!g1236) & (!g1247) & (g1271) & (g1278)) + ((!g1234) & (!g1235) & (!g1236) & (g1247) & (!g1271) & (!g1278)) + ((!g1234) & (!g1235) & (!g1236) & (g1247) & (g1271) & (g1278)) + ((!g1234) & (!g1235) & (g1236) & (!g1247) & (!g1271) & (!g1278)) + ((!g1234) & (!g1235) & (g1236) & (!g1247) & (g1271) & (g1278)) + ((!g1234) & (!g1235) & (g1236) & (g1247) & (!g1271) & (g1278)) + ((!g1234) & (!g1235) & (g1236) & (g1247) & (g1271) & (!g1278)) + ((!g1234) & (g1235) & (!g1236) & (!g1247) & (!g1271) & (!g1278)) + ((!g1234) & (g1235) & (!g1236) & (!g1247) & (g1271) & (g1278)) + ((!g1234) & (g1235) & (!g1236) & (g1247) & (!g1271) & (g1278)) + ((!g1234) & (g1235) & (!g1236) & (g1247) & (g1271) & (!g1278)) + ((!g1234) & (g1235) & (g1236) & (!g1247) & (!g1271) & (g1278)) + ((!g1234) & (g1235) & (g1236) & (!g1247) & (g1271) & (!g1278)) + ((!g1234) & (g1235) & (g1236) & (g1247) & (!g1271) & (g1278)) + ((!g1234) & (g1235) & (g1236) & (g1247) & (g1271) & (!g1278)) + ((g1234) & (!g1235) & (!g1236) & (!g1247) & (!g1271) & (!g1278)) + ((g1234) & (!g1235) & (!g1236) & (!g1247) & (g1271) & (g1278)) + ((g1234) & (!g1235) & (!g1236) & (g1247) & (!g1271) & (g1278)) + ((g1234) & (!g1235) & (!g1236) & (g1247) & (g1271) & (!g1278)) + ((g1234) & (!g1235) & (g1236) & (!g1247) & (!g1271) & (g1278)) + ((g1234) & (!g1235) & (g1236) & (!g1247) & (g1271) & (!g1278)) + ((g1234) & (!g1235) & (g1236) & (g1247) & (!g1271) & (g1278)) + ((g1234) & (!g1235) & (g1236) & (g1247) & (g1271) & (!g1278)) + ((g1234) & (g1235) & (!g1236) & (!g1247) & (!g1271) & (!g1278)) + ((g1234) & (g1235) & (!g1236) & (!g1247) & (g1271) & (g1278)) + ((g1234) & (g1235) & (!g1236) & (g1247) & (!g1271) & (g1278)) + ((g1234) & (g1235) & (!g1236) & (g1247) & (g1271) & (!g1278)) + ((g1234) & (g1235) & (g1236) & (!g1247) & (!g1271) & (g1278)) + ((g1234) & (g1235) & (g1236) & (!g1247) & (g1271) & (!g1278)) + ((g1234) & (g1235) & (g1236) & (g1247) & (!g1271) & (g1278)) + ((g1234) & (g1235) & (g1236) & (g1247) & (g1271) & (!g1278)));
	assign g1280 = (((!g1068) & (!g1232) & (!g1254) & (!g1255) & (!g1258) & (!g1279)) + ((!g1068) & (!g1232) & (!g1254) & (!g1255) & (g1258) & (g1279)) + ((!g1068) & (!g1232) & (!g1254) & (g1255) & (!g1258) & (!g1279)) + ((!g1068) & (!g1232) & (!g1254) & (g1255) & (g1258) & (g1279)) + ((!g1068) & (!g1232) & (g1254) & (!g1255) & (!g1258) & (!g1279)) + ((!g1068) & (!g1232) & (g1254) & (!g1255) & (g1258) & (g1279)) + ((!g1068) & (!g1232) & (g1254) & (g1255) & (!g1258) & (!g1279)) + ((!g1068) & (!g1232) & (g1254) & (g1255) & (g1258) & (g1279)) + ((!g1068) & (g1232) & (!g1254) & (!g1255) & (!g1258) & (!g1279)) + ((!g1068) & (g1232) & (!g1254) & (!g1255) & (g1258) & (g1279)) + ((!g1068) & (g1232) & (!g1254) & (g1255) & (!g1258) & (!g1279)) + ((!g1068) & (g1232) & (!g1254) & (g1255) & (g1258) & (g1279)) + ((!g1068) & (g1232) & (g1254) & (!g1255) & (!g1258) & (g1279)) + ((!g1068) & (g1232) & (g1254) & (!g1255) & (g1258) & (!g1279)) + ((!g1068) & (g1232) & (g1254) & (g1255) & (!g1258) & (g1279)) + ((!g1068) & (g1232) & (g1254) & (g1255) & (g1258) & (!g1279)) + ((g1068) & (!g1232) & (!g1254) & (!g1255) & (!g1258) & (g1279)) + ((g1068) & (!g1232) & (!g1254) & (!g1255) & (g1258) & (!g1279)) + ((g1068) & (!g1232) & (!g1254) & (g1255) & (!g1258) & (!g1279)) + ((g1068) & (!g1232) & (!g1254) & (g1255) & (g1258) & (g1279)) + ((g1068) & (!g1232) & (g1254) & (!g1255) & (!g1258) & (g1279)) + ((g1068) & (!g1232) & (g1254) & (!g1255) & (g1258) & (!g1279)) + ((g1068) & (!g1232) & (g1254) & (g1255) & (!g1258) & (g1279)) + ((g1068) & (!g1232) & (g1254) & (g1255) & (g1258) & (!g1279)) + ((g1068) & (g1232) & (!g1254) & (!g1255) & (!g1258) & (g1279)) + ((g1068) & (g1232) & (!g1254) & (!g1255) & (g1258) & (!g1279)) + ((g1068) & (g1232) & (!g1254) & (g1255) & (!g1258) & (g1279)) + ((g1068) & (g1232) & (!g1254) & (g1255) & (g1258) & (!g1279)) + ((g1068) & (g1232) & (g1254) & (!g1255) & (!g1258) & (!g1279)) + ((g1068) & (g1232) & (g1254) & (!g1255) & (g1258) & (g1279)) + ((g1068) & (g1232) & (g1254) & (g1255) & (!g1258) & (g1279)) + ((g1068) & (g1232) & (g1254) & (g1255) & (g1258) & (!g1279)));
	assign g1281 = (((!g1232) & (!sk[11]) & (!g1254) & (!g1255) & (g1258) & (!g1279)) + ((!g1232) & (!sk[11]) & (!g1254) & (!g1255) & (g1258) & (g1279)) + ((!g1232) & (!sk[11]) & (!g1254) & (g1255) & (!g1258) & (!g1279)) + ((!g1232) & (!sk[11]) & (!g1254) & (g1255) & (!g1258) & (g1279)) + ((!g1232) & (!sk[11]) & (!g1254) & (g1255) & (g1258) & (!g1279)) + ((!g1232) & (!sk[11]) & (!g1254) & (g1255) & (g1258) & (g1279)) + ((!g1232) & (!sk[11]) & (g1254) & (!g1255) & (!g1258) & (!g1279)) + ((!g1232) & (!sk[11]) & (g1254) & (!g1255) & (!g1258) & (g1279)) + ((!g1232) & (!sk[11]) & (g1254) & (!g1255) & (g1258) & (!g1279)) + ((!g1232) & (!sk[11]) & (g1254) & (!g1255) & (g1258) & (g1279)) + ((!g1232) & (!sk[11]) & (g1254) & (g1255) & (!g1258) & (!g1279)) + ((!g1232) & (!sk[11]) & (g1254) & (g1255) & (!g1258) & (g1279)) + ((!g1232) & (!sk[11]) & (g1254) & (g1255) & (g1258) & (!g1279)) + ((!g1232) & (!sk[11]) & (g1254) & (g1255) & (g1258) & (g1279)) + ((!g1232) & (sk[11]) & (!g1254) & (g1255) & (!g1258) & (!g1279)) + ((!g1232) & (sk[11]) & (!g1254) & (g1255) & (g1258) & (g1279)) + ((g1232) & (!sk[11]) & (!g1254) & (!g1255) & (g1258) & (!g1279)) + ((g1232) & (!sk[11]) & (!g1254) & (!g1255) & (g1258) & (g1279)) + ((g1232) & (!sk[11]) & (!g1254) & (g1255) & (!g1258) & (!g1279)) + ((g1232) & (!sk[11]) & (!g1254) & (g1255) & (!g1258) & (g1279)) + ((g1232) & (!sk[11]) & (!g1254) & (g1255) & (g1258) & (!g1279)) + ((g1232) & (!sk[11]) & (!g1254) & (g1255) & (g1258) & (g1279)) + ((g1232) & (!sk[11]) & (g1254) & (!g1255) & (!g1258) & (!g1279)) + ((g1232) & (!sk[11]) & (g1254) & (!g1255) & (!g1258) & (g1279)) + ((g1232) & (!sk[11]) & (g1254) & (!g1255) & (g1258) & (!g1279)) + ((g1232) & (!sk[11]) & (g1254) & (!g1255) & (g1258) & (g1279)) + ((g1232) & (!sk[11]) & (g1254) & (g1255) & (!g1258) & (!g1279)) + ((g1232) & (!sk[11]) & (g1254) & (g1255) & (!g1258) & (g1279)) + ((g1232) & (!sk[11]) & (g1254) & (g1255) & (g1258) & (!g1279)) + ((g1232) & (!sk[11]) & (g1254) & (g1255) & (g1258) & (g1279)) + ((g1232) & (sk[11]) & (g1254) & (g1255) & (!g1258) & (g1279)) + ((g1232) & (sk[11]) & (g1254) & (g1255) & (g1258) & (!g1279)));
	assign g1282 = (((g1186) & (!g1207) & (!g1209) & (!g1230) & (!g1233) & (g1253)) + ((g1186) & (!g1207) & (!g1209) & (!g1230) & (g1233) & (!g1253)) + ((g1186) & (!g1207) & (g1209) & (g1230) & (!g1233) & (g1253)) + ((g1186) & (!g1207) & (g1209) & (g1230) & (g1233) & (!g1253)));
	assign g1283 = (((!g1282) & (!sk[13]) & (g1258) & (!g1279)) + ((!g1282) & (!sk[13]) & (g1258) & (g1279)) + ((g1282) & (!sk[13]) & (g1258) & (!g1279)) + ((g1282) & (!sk[13]) & (g1258) & (g1279)) + ((g1282) & (sk[13]) & (!g1258) & (g1279)) + ((g1282) & (sk[13]) & (g1258) & (!g1279)));
	assign g1284 = (((!g1234) & (!g1235) & (!g1236) & (!g1247) & (!g1271) & (!g1278)) + ((!g1234) & (!g1235) & (!g1236) & (g1247) & (!g1271) & (!g1278)) + ((!g1234) & (!g1235) & (g1236) & (!g1247) & (!g1271) & (!g1278)) + ((!g1234) & (!g1235) & (g1236) & (g1247) & (g1271) & (!g1278)) + ((!g1234) & (g1235) & (!g1236) & (!g1247) & (!g1271) & (!g1278)) + ((!g1234) & (g1235) & (!g1236) & (g1247) & (g1271) & (!g1278)) + ((!g1234) & (g1235) & (g1236) & (!g1247) & (g1271) & (!g1278)) + ((!g1234) & (g1235) & (g1236) & (g1247) & (g1271) & (!g1278)) + ((g1234) & (!g1235) & (!g1236) & (!g1247) & (!g1271) & (!g1278)) + ((g1234) & (!g1235) & (!g1236) & (g1247) & (g1271) & (!g1278)) + ((g1234) & (!g1235) & (g1236) & (!g1247) & (g1271) & (!g1278)) + ((g1234) & (!g1235) & (g1236) & (g1247) & (g1271) & (!g1278)) + ((g1234) & (g1235) & (!g1236) & (!g1247) & (!g1271) & (!g1278)) + ((g1234) & (g1235) & (!g1236) & (g1247) & (g1271) & (!g1278)) + ((g1234) & (g1235) & (g1236) & (!g1247) & (g1271) & (!g1278)) + ((g1234) & (g1235) & (g1236) & (g1247) & (g1271) & (!g1278)));
	assign g1285 = (((!g1209) & (!g1230) & (!g1233) & (g1257) & (!g1252) & (!g1279)) + ((!g1209) & (!g1230) & (g1233) & (!g1257) & (!g1252) & (!g1279)) + ((!g1209) & (!g1230) & (g1233) & (g1257) & (!g1252) & (!g1279)) + ((!g1209) & (!g1230) & (g1233) & (g1257) & (g1252) & (!g1279)) + ((!g1209) & (g1230) & (!g1233) & (g1257) & (!g1252) & (!g1279)) + ((!g1209) & (g1230) & (g1233) & (!g1257) & (!g1252) & (!g1279)) + ((!g1209) & (g1230) & (g1233) & (g1257) & (!g1252) & (!g1279)) + ((!g1209) & (g1230) & (g1233) & (g1257) & (g1252) & (!g1279)) + ((g1209) & (!g1230) & (!g1233) & (!g1257) & (!g1252) & (!g1279)) + ((g1209) & (!g1230) & (!g1233) & (g1257) & (!g1252) & (!g1279)) + ((g1209) & (!g1230) & (!g1233) & (g1257) & (g1252) & (!g1279)) + ((g1209) & (!g1230) & (g1233) & (!g1257) & (!g1252) & (!g1279)) + ((g1209) & (!g1230) & (g1233) & (g1257) & (!g1252) & (!g1279)) + ((g1209) & (!g1230) & (g1233) & (g1257) & (g1252) & (!g1279)) + ((g1209) & (g1230) & (!g1233) & (g1257) & (!g1252) & (!g1279)) + ((g1209) & (g1230) & (g1233) & (!g1257) & (!g1252) & (!g1279)) + ((g1209) & (g1230) & (g1233) & (g1257) & (!g1252) & (!g1279)) + ((g1209) & (g1230) & (g1233) & (g1257) & (g1252) & (!g1279)));
	assign g1286 = (((!g1234) & (!g1235) & (!g1236) & (!g1247) & (!g1259) & (!g1270)) + ((!g1234) & (!g1235) & (!g1236) & (!g1247) & (!g1259) & (g1270)) + ((!g1234) & (!g1235) & (!g1236) & (!g1247) & (g1259) & (g1270)) + ((!g1234) & (!g1235) & (!g1236) & (g1247) & (!g1259) & (!g1270)) + ((!g1234) & (!g1235) & (!g1236) & (g1247) & (!g1259) & (g1270)) + ((!g1234) & (!g1235) & (!g1236) & (g1247) & (g1259) & (g1270)) + ((!g1234) & (!g1235) & (g1236) & (!g1247) & (!g1259) & (!g1270)) + ((!g1234) & (!g1235) & (g1236) & (!g1247) & (!g1259) & (g1270)) + ((!g1234) & (!g1235) & (g1236) & (!g1247) & (g1259) & (g1270)) + ((!g1234) & (!g1235) & (g1236) & (g1247) & (!g1259) & (g1270)) + ((!g1234) & (g1235) & (!g1236) & (!g1247) & (!g1259) & (!g1270)) + ((!g1234) & (g1235) & (!g1236) & (!g1247) & (!g1259) & (g1270)) + ((!g1234) & (g1235) & (!g1236) & (!g1247) & (g1259) & (g1270)) + ((!g1234) & (g1235) & (!g1236) & (g1247) & (!g1259) & (g1270)) + ((!g1234) & (g1235) & (g1236) & (!g1247) & (!g1259) & (g1270)) + ((!g1234) & (g1235) & (g1236) & (g1247) & (!g1259) & (g1270)) + ((g1234) & (!g1235) & (!g1236) & (!g1247) & (!g1259) & (!g1270)) + ((g1234) & (!g1235) & (!g1236) & (!g1247) & (!g1259) & (g1270)) + ((g1234) & (!g1235) & (!g1236) & (!g1247) & (g1259) & (g1270)) + ((g1234) & (!g1235) & (!g1236) & (g1247) & (!g1259) & (g1270)) + ((g1234) & (!g1235) & (g1236) & (!g1247) & (!g1259) & (g1270)) + ((g1234) & (!g1235) & (g1236) & (g1247) & (!g1259) & (g1270)) + ((g1234) & (g1235) & (!g1236) & (!g1247) & (!g1259) & (!g1270)) + ((g1234) & (g1235) & (!g1236) & (!g1247) & (!g1259) & (g1270)) + ((g1234) & (g1235) & (!g1236) & (!g1247) & (g1259) & (g1270)) + ((g1234) & (g1235) & (!g1236) & (g1247) & (!g1259) & (g1270)) + ((g1234) & (g1235) & (g1236) & (!g1247) & (!g1259) & (g1270)) + ((g1234) & (g1235) & (g1236) & (g1247) & (!g1259) & (g1270)));
	assign g1287 = (((!g1240) & (!g1260) & (!g1245) & (!g1267) & (sk[17]) & (!g1269)) + ((!g1240) & (!g1260) & (!g1245) & (!g1267) & (sk[17]) & (g1269)) + ((!g1240) & (!g1260) & (!g1245) & (g1267) & (!sk[17]) & (!g1269)) + ((!g1240) & (!g1260) & (!g1245) & (g1267) & (!sk[17]) & (g1269)) + ((!g1240) & (!g1260) & (!g1245) & (g1267) & (sk[17]) & (g1269)) + ((!g1240) & (!g1260) & (g1245) & (!g1267) & (!sk[17]) & (!g1269)) + ((!g1240) & (!g1260) & (g1245) & (!g1267) & (!sk[17]) & (g1269)) + ((!g1240) & (!g1260) & (g1245) & (!g1267) & (sk[17]) & (!g1269)) + ((!g1240) & (!g1260) & (g1245) & (!g1267) & (sk[17]) & (g1269)) + ((!g1240) & (!g1260) & (g1245) & (g1267) & (!sk[17]) & (!g1269)) + ((!g1240) & (!g1260) & (g1245) & (g1267) & (!sk[17]) & (g1269)) + ((!g1240) & (!g1260) & (g1245) & (g1267) & (sk[17]) & (g1269)) + ((!g1240) & (g1260) & (!g1245) & (!g1267) & (!sk[17]) & (!g1269)) + ((!g1240) & (g1260) & (!g1245) & (!g1267) & (!sk[17]) & (g1269)) + ((!g1240) & (g1260) & (!g1245) & (!g1267) & (sk[17]) & (g1269)) + ((!g1240) & (g1260) & (!g1245) & (g1267) & (!sk[17]) & (!g1269)) + ((!g1240) & (g1260) & (!g1245) & (g1267) & (!sk[17]) & (g1269)) + ((!g1240) & (g1260) & (g1245) & (!g1267) & (!sk[17]) & (!g1269)) + ((!g1240) & (g1260) & (g1245) & (!g1267) & (!sk[17]) & (g1269)) + ((!g1240) & (g1260) & (g1245) & (!g1267) & (sk[17]) & (!g1269)) + ((!g1240) & (g1260) & (g1245) & (!g1267) & (sk[17]) & (g1269)) + ((!g1240) & (g1260) & (g1245) & (g1267) & (!sk[17]) & (!g1269)) + ((!g1240) & (g1260) & (g1245) & (g1267) & (!sk[17]) & (g1269)) + ((!g1240) & (g1260) & (g1245) & (g1267) & (sk[17]) & (g1269)) + ((g1240) & (!g1260) & (!g1245) & (!g1267) & (sk[17]) & (g1269)) + ((g1240) & (!g1260) & (!g1245) & (g1267) & (!sk[17]) & (!g1269)) + ((g1240) & (!g1260) & (!g1245) & (g1267) & (!sk[17]) & (g1269)) + ((g1240) & (!g1260) & (g1245) & (!g1267) & (!sk[17]) & (!g1269)) + ((g1240) & (!g1260) & (g1245) & (!g1267) & (!sk[17]) & (g1269)) + ((g1240) & (!g1260) & (g1245) & (!g1267) & (sk[17]) & (!g1269)) + ((g1240) & (!g1260) & (g1245) & (!g1267) & (sk[17]) & (g1269)) + ((g1240) & (!g1260) & (g1245) & (g1267) & (!sk[17]) & (!g1269)) + ((g1240) & (!g1260) & (g1245) & (g1267) & (!sk[17]) & (g1269)) + ((g1240) & (!g1260) & (g1245) & (g1267) & (sk[17]) & (g1269)) + ((g1240) & (g1260) & (!g1245) & (!g1267) & (!sk[17]) & (!g1269)) + ((g1240) & (g1260) & (!g1245) & (!g1267) & (!sk[17]) & (g1269)) + ((g1240) & (g1260) & (!g1245) & (!g1267) & (sk[17]) & (g1269)) + ((g1240) & (g1260) & (!g1245) & (g1267) & (!sk[17]) & (!g1269)) + ((g1240) & (g1260) & (!g1245) & (g1267) & (!sk[17]) & (g1269)) + ((g1240) & (g1260) & (g1245) & (!g1267) & (!sk[17]) & (!g1269)) + ((g1240) & (g1260) & (g1245) & (!g1267) & (!sk[17]) & (g1269)) + ((g1240) & (g1260) & (g1245) & (!g1267) & (sk[17]) & (g1269)) + ((g1240) & (g1260) & (g1245) & (g1267) & (!sk[17]) & (!g1269)) + ((g1240) & (g1260) & (g1245) & (g1267) & (!sk[17]) & (g1269)));
	assign g1288 = (((!g202) & (!g759) & (!g995) & (!g1261) & (!g1262) & (!g1266)) + ((!g202) & (!g759) & (!g995) & (!g1261) & (g1262) & (!g1266)) + ((!g202) & (!g759) & (!g995) & (!g1261) & (g1262) & (g1266)) + ((!g202) & (!g759) & (!g995) & (g1261) & (g1262) & (!g1266)) + ((!g202) & (!g759) & (g995) & (!g1261) & (!g1262) & (!g1266)) + ((!g202) & (!g759) & (g995) & (!g1261) & (g1262) & (!g1266)) + ((!g202) & (!g759) & (g995) & (!g1261) & (g1262) & (g1266)) + ((!g202) & (!g759) & (g995) & (g1261) & (g1262) & (!g1266)) + ((!g202) & (g759) & (!g995) & (!g1261) & (!g1262) & (!g1266)) + ((!g202) & (g759) & (!g995) & (!g1261) & (g1262) & (!g1266)) + ((!g202) & (g759) & (!g995) & (!g1261) & (g1262) & (g1266)) + ((!g202) & (g759) & (!g995) & (g1261) & (g1262) & (!g1266)) + ((!g202) & (g759) & (g995) & (!g1261) & (!g1262) & (!g1266)) + ((!g202) & (g759) & (g995) & (!g1261) & (g1262) & (!g1266)) + ((!g202) & (g759) & (g995) & (!g1261) & (g1262) & (g1266)) + ((!g202) & (g759) & (g995) & (g1261) & (!g1262) & (!g1266)) + ((!g202) & (g759) & (g995) & (g1261) & (g1262) & (!g1266)) + ((!g202) & (g759) & (g995) & (g1261) & (g1262) & (g1266)) + ((g202) & (!g759) & (!g995) & (!g1261) & (g1262) & (!g1266)) + ((g202) & (!g759) & (!g995) & (g1261) & (!g1262) & (!g1266)) + ((g202) & (!g759) & (!g995) & (g1261) & (g1262) & (!g1266)) + ((g202) & (!g759) & (!g995) & (g1261) & (g1262) & (g1266)) + ((g202) & (!g759) & (g995) & (!g1261) & (g1262) & (!g1266)) + ((g202) & (!g759) & (g995) & (g1261) & (!g1262) & (!g1266)) + ((g202) & (!g759) & (g995) & (g1261) & (g1262) & (!g1266)) + ((g202) & (!g759) & (g995) & (g1261) & (g1262) & (g1266)) + ((g202) & (g759) & (!g995) & (!g1261) & (g1262) & (!g1266)) + ((g202) & (g759) & (!g995) & (g1261) & (!g1262) & (!g1266)) + ((g202) & (g759) & (!g995) & (g1261) & (g1262) & (!g1266)) + ((g202) & (g759) & (!g995) & (g1261) & (g1262) & (g1266)) + ((g202) & (g759) & (g995) & (!g1261) & (g1262) & (!g1266)) + ((g202) & (g759) & (g995) & (g1261) & (g1262) & (!g1266)));
	assign g1289 = (((!g200) & (!g742) & (g748) & (!g1040) & (!g1079) & (!g1080)) + ((!g200) & (!g742) & (g748) & (!g1040) & (!g1079) & (g1080)) + ((!g200) & (!g742) & (g748) & (g1040) & (!g1079) & (!g1080)) + ((!g200) & (!g742) & (g748) & (g1040) & (!g1079) & (g1080)) + ((!g200) & (g742) & (!g748) & (!g1040) & (!g1079) & (!g1080)) + ((!g200) & (g742) & (!g748) & (!g1040) & (!g1079) & (g1080)) + ((!g200) & (g742) & (!g748) & (g1040) & (!g1079) & (g1080)) + ((!g200) & (g742) & (g748) & (!g1040) & (!g1079) & (!g1080)) + ((!g200) & (g742) & (g748) & (!g1040) & (!g1079) & (g1080)) + ((!g200) & (g742) & (g748) & (g1040) & (!g1079) & (!g1080)) + ((!g200) & (g742) & (g748) & (g1040) & (!g1079) & (g1080)) + ((g200) & (!g742) & (!g748) & (!g1040) & (!g1079) & (!g1080)) + ((g200) & (!g742) & (!g748) & (!g1040) & (!g1079) & (g1080)) + ((g200) & (!g742) & (!g748) & (!g1040) & (g1079) & (!g1080)) + ((g200) & (!g742) & (!g748) & (!g1040) & (g1079) & (g1080)) + ((g200) & (!g742) & (!g748) & (g1040) & (!g1079) & (!g1080)) + ((g200) & (!g742) & (!g748) & (g1040) & (!g1079) & (g1080)) + ((g200) & (!g742) & (!g748) & (g1040) & (g1079) & (!g1080)) + ((g200) & (!g742) & (!g748) & (g1040) & (g1079) & (g1080)) + ((g200) & (!g742) & (g748) & (!g1040) & (g1079) & (!g1080)) + ((g200) & (!g742) & (g748) & (!g1040) & (g1079) & (g1080)) + ((g200) & (!g742) & (g748) & (g1040) & (g1079) & (!g1080)) + ((g200) & (!g742) & (g748) & (g1040) & (g1079) & (g1080)) + ((g200) & (g742) & (!g748) & (!g1040) & (g1079) & (!g1080)) + ((g200) & (g742) & (!g748) & (!g1040) & (g1079) & (g1080)) + ((g200) & (g742) & (!g748) & (g1040) & (!g1079) & (!g1080)) + ((g200) & (g742) & (!g748) & (g1040) & (g1079) & (!g1080)) + ((g200) & (g742) & (!g748) & (g1040) & (g1079) & (g1080)) + ((g200) & (g742) & (g748) & (!g1040) & (g1079) & (!g1080)) + ((g200) & (g742) & (g748) & (!g1040) & (g1079) & (g1080)) + ((g200) & (g742) & (g748) & (g1040) & (g1079) & (!g1080)) + ((g200) & (g742) & (g748) & (g1040) & (g1079) & (g1080)));
	assign g1290 = (((!sk[20]) & (!g843) & (g884) & (!g890)) + ((!sk[20]) & (!g843) & (g884) & (g890)) + ((!sk[20]) & (g843) & (g884) & (!g890)) + ((!sk[20]) & (g843) & (g884) & (g890)) + ((sk[20]) & (g843) & (!g884) & (!g890)) + ((sk[20]) & (g843) & (g884) & (g890)));
	assign g1291 = (((!g847) & (!g845) & (!g848) & (!g962) & (!g863) & (!g963)) + ((!g847) & (!g845) & (!g848) & (!g962) & (!g863) & (g963)) + ((!g847) & (!g845) & (!g848) & (!g962) & (g863) & (!g963)) + ((!g847) & (!g845) & (!g848) & (!g962) & (g863) & (g963)) + ((!g847) & (!g845) & (!g848) & (g962) & (!g863) & (!g963)) + ((!g847) & (!g845) & (!g848) & (g962) & (!g863) & (g963)) + ((!g847) & (!g845) & (!g848) & (g962) & (g863) & (!g963)) + ((!g847) & (!g845) & (!g848) & (g962) & (g863) & (g963)) + ((!g847) & (!g845) & (g848) & (!g962) & (!g863) & (!g963)) + ((!g847) & (!g845) & (g848) & (!g962) & (!g863) & (g963)) + ((!g847) & (!g845) & (g848) & (g962) & (!g863) & (!g963)) + ((!g847) & (!g845) & (g848) & (g962) & (!g863) & (g963)) + ((!g847) & (g845) & (!g848) & (!g962) & (!g863) & (!g963)) + ((!g847) & (g845) & (!g848) & (!g962) & (g863) & (!g963)) + ((!g847) & (g845) & (!g848) & (g962) & (!g863) & (!g963)) + ((!g847) & (g845) & (!g848) & (g962) & (g863) & (!g963)) + ((!g847) & (g845) & (g848) & (!g962) & (!g863) & (!g963)) + ((!g847) & (g845) & (g848) & (g962) & (!g863) & (!g963)) + ((g847) & (!g845) & (!g848) & (g962) & (!g863) & (!g963)) + ((g847) & (!g845) & (!g848) & (g962) & (!g863) & (g963)) + ((g847) & (!g845) & (!g848) & (g962) & (g863) & (!g963)) + ((g847) & (!g845) & (!g848) & (g962) & (g863) & (g963)) + ((g847) & (!g845) & (g848) & (g962) & (!g863) & (!g963)) + ((g847) & (!g845) & (g848) & (g962) & (!g863) & (g963)) + ((g847) & (g845) & (!g848) & (g962) & (!g863) & (!g963)) + ((g847) & (g845) & (!g848) & (g962) & (g863) & (!g963)) + ((g847) & (g845) & (g848) & (g962) & (!g863) & (!g963)));
	assign g1292 = (((!g252) & (!g835) & (!g1290) & (!sk[22]) & (g1291)) + ((!g252) & (!g835) & (!g1290) & (sk[22]) & (g1291)) + ((!g252) & (!g835) & (g1290) & (!sk[22]) & (g1291)) + ((!g252) & (g835) & (!g1290) & (!sk[22]) & (g1291)) + ((!g252) & (g835) & (!g1290) & (sk[22]) & (g1291)) + ((!g252) & (g835) & (g1290) & (!sk[22]) & (g1291)) + ((g252) & (!g835) & (!g1290) & (!sk[22]) & (!g1291)) + ((g252) & (!g835) & (!g1290) & (!sk[22]) & (g1291)) + ((g252) & (!g835) & (!g1290) & (sk[22]) & (g1291)) + ((g252) & (!g835) & (g1290) & (!sk[22]) & (!g1291)) + ((g252) & (!g835) & (g1290) & (!sk[22]) & (g1291)) + ((g252) & (g835) & (!g1290) & (!sk[22]) & (!g1291)) + ((g252) & (g835) & (!g1290) & (!sk[22]) & (g1291)) + ((g252) & (g835) & (!g1290) & (sk[22]) & (!g1291)) + ((g252) & (g835) & (g1290) & (!sk[22]) & (!g1291)) + ((g252) & (g835) & (g1290) & (!sk[22]) & (g1291)) + ((g252) & (g835) & (g1290) & (sk[22]) & (!g1291)) + ((g252) & (g835) & (g1290) & (sk[22]) & (g1291)));
	assign g1293 = (((!g252) & (!g869) & (!g843) & (!g895) & (!g1263) & (g1265)) + ((!g252) & (!g869) & (!g843) & (g895) & (!g1263) & (g1265)) + ((!g252) & (!g869) & (g843) & (!g895) & (!g1263) & (g1265)) + ((!g252) & (g869) & (!g843) & (!g895) & (!g1263) & (g1265)) + ((!g252) & (g869) & (!g843) & (g895) & (!g1263) & (g1265)) + ((!g252) & (g869) & (g843) & (!g895) & (!g1263) & (g1265)) + ((g252) & (!g869) & (!g843) & (!g895) & (!g1263) & (!g1265)) + ((g252) & (!g869) & (!g843) & (g895) & (!g1263) & (!g1265)) + ((g252) & (!g869) & (g843) & (!g895) & (!g1263) & (!g1265)) + ((g252) & (!g869) & (g843) & (g895) & (!g1263) & (!g1265)) + ((g252) & (!g869) & (g843) & (g895) & (!g1263) & (g1265)) + ((g252) & (g869) & (!g843) & (!g895) & (!g1263) & (!g1265)) + ((g252) & (g869) & (!g843) & (!g895) & (!g1263) & (g1265)) + ((g252) & (g869) & (!g843) & (!g895) & (g1263) & (!g1265)) + ((g252) & (g869) & (!g843) & (g895) & (!g1263) & (!g1265)) + ((g252) & (g869) & (!g843) & (g895) & (!g1263) & (g1265)) + ((g252) & (g869) & (!g843) & (g895) & (g1263) & (!g1265)) + ((g252) & (g869) & (g843) & (!g895) & (!g1263) & (!g1265)) + ((g252) & (g869) & (g843) & (!g895) & (!g1263) & (g1265)) + ((g252) & (g869) & (g843) & (!g895) & (g1263) & (!g1265)) + ((g252) & (g869) & (g843) & (g895) & (!g1263) & (!g1265)) + ((g252) & (g869) & (g843) & (g895) & (!g1263) & (g1265)) + ((g252) & (g869) & (g843) & (g895) & (g1263) & (!g1265)) + ((g252) & (g869) & (g843) & (g895) & (g1263) & (g1265)));
	assign g1294 = (((!g764) & (!g762) & (!g994) & (!sk[24]) & (g1040)) + ((!g764) & (!g762) & (g994) & (!sk[24]) & (g1040)) + ((!g764) & (g762) & (!g994) & (!sk[24]) & (g1040)) + ((!g764) & (g762) & (g994) & (!sk[24]) & (g1040)) + ((!g764) & (g762) & (g994) & (sk[24]) & (!g1040)) + ((!g764) & (g762) & (g994) & (sk[24]) & (g1040)) + ((g764) & (!g762) & (!g994) & (!sk[24]) & (!g1040)) + ((g764) & (!g762) & (!g994) & (!sk[24]) & (g1040)) + ((g764) & (!g762) & (!g994) & (sk[24]) & (!g1040)) + ((g764) & (!g762) & (g994) & (!sk[24]) & (!g1040)) + ((g764) & (!g762) & (g994) & (!sk[24]) & (g1040)) + ((g764) & (!g762) & (g994) & (sk[24]) & (!g1040)) + ((g764) & (g762) & (!g994) & (!sk[24]) & (!g1040)) + ((g764) & (g762) & (!g994) & (!sk[24]) & (g1040)) + ((g764) & (g762) & (!g994) & (sk[24]) & (!g1040)) + ((g764) & (g762) & (g994) & (!sk[24]) & (!g1040)) + ((g764) & (g762) & (g994) & (!sk[24]) & (g1040)) + ((g764) & (g762) & (g994) & (sk[24]) & (!g1040)) + ((g764) & (g762) & (g994) & (sk[24]) & (g1040)));
	assign g1295 = (((!g202) & (!g759) & (!g765) & (!g971) & (!g1041) & (g1294)) + ((!g202) & (!g759) & (!g765) & (!g971) & (g1041) & (g1294)) + ((!g202) & (!g759) & (!g765) & (g971) & (!g1041) & (g1294)) + ((!g202) & (!g759) & (!g765) & (g971) & (g1041) & (g1294)) + ((!g202) & (!g759) & (g765) & (!g971) & (!g1041) & (g1294)) + ((!g202) & (!g759) & (g765) & (!g971) & (g1041) & (g1294)) + ((!g202) & (!g759) & (g765) & (g971) & (!g1041) & (!g1294)) + ((!g202) & (!g759) & (g765) & (g971) & (!g1041) & (g1294)) + ((!g202) & (!g759) & (g765) & (g971) & (g1041) & (!g1294)) + ((!g202) & (!g759) & (g765) & (g971) & (g1041) & (g1294)) + ((!g202) & (g759) & (!g765) & (!g971) & (!g1041) & (!g1294)) + ((!g202) & (g759) & (!g765) & (!g971) & (!g1041) & (g1294)) + ((!g202) & (g759) & (!g765) & (!g971) & (g1041) & (g1294)) + ((!g202) & (g759) & (!g765) & (g971) & (!g1041) & (!g1294)) + ((!g202) & (g759) & (!g765) & (g971) & (!g1041) & (g1294)) + ((!g202) & (g759) & (!g765) & (g971) & (g1041) & (g1294)) + ((!g202) & (g759) & (g765) & (!g971) & (!g1041) & (!g1294)) + ((!g202) & (g759) & (g765) & (!g971) & (!g1041) & (g1294)) + ((!g202) & (g759) & (g765) & (!g971) & (g1041) & (g1294)) + ((!g202) & (g759) & (g765) & (g971) & (!g1041) & (!g1294)) + ((!g202) & (g759) & (g765) & (g971) & (!g1041) & (g1294)) + ((!g202) & (g759) & (g765) & (g971) & (g1041) & (!g1294)) + ((!g202) & (g759) & (g765) & (g971) & (g1041) & (g1294)) + ((g202) & (!g759) & (!g765) & (!g971) & (!g1041) & (!g1294)) + ((g202) & (!g759) & (!g765) & (!g971) & (g1041) & (!g1294)) + ((g202) & (!g759) & (!g765) & (g971) & (!g1041) & (!g1294)) + ((g202) & (!g759) & (!g765) & (g971) & (g1041) & (!g1294)) + ((g202) & (!g759) & (g765) & (!g971) & (!g1041) & (!g1294)) + ((g202) & (!g759) & (g765) & (!g971) & (g1041) & (!g1294)) + ((g202) & (g759) & (!g765) & (!g971) & (g1041) & (!g1294)) + ((g202) & (g759) & (!g765) & (g971) & (g1041) & (!g1294)) + ((g202) & (g759) & (g765) & (!g971) & (g1041) & (!g1294)));
	assign g1296 = (((!g1288) & (!g1289) & (!g1292) & (!sk[26]) & (g1293) & (!g1295)) + ((!g1288) & (!g1289) & (!g1292) & (!sk[26]) & (g1293) & (g1295)) + ((!g1288) & (!g1289) & (!g1292) & (sk[26]) & (!g1293) & (g1295)) + ((!g1288) & (!g1289) & (!g1292) & (sk[26]) & (g1293) & (!g1295)) + ((!g1288) & (!g1289) & (g1292) & (!sk[26]) & (!g1293) & (!g1295)) + ((!g1288) & (!g1289) & (g1292) & (!sk[26]) & (!g1293) & (g1295)) + ((!g1288) & (!g1289) & (g1292) & (!sk[26]) & (g1293) & (!g1295)) + ((!g1288) & (!g1289) & (g1292) & (!sk[26]) & (g1293) & (g1295)) + ((!g1288) & (!g1289) & (g1292) & (sk[26]) & (!g1293) & (!g1295)) + ((!g1288) & (!g1289) & (g1292) & (sk[26]) & (g1293) & (g1295)) + ((!g1288) & (g1289) & (!g1292) & (!sk[26]) & (!g1293) & (!g1295)) + ((!g1288) & (g1289) & (!g1292) & (!sk[26]) & (!g1293) & (g1295)) + ((!g1288) & (g1289) & (!g1292) & (!sk[26]) & (g1293) & (!g1295)) + ((!g1288) & (g1289) & (!g1292) & (!sk[26]) & (g1293) & (g1295)) + ((!g1288) & (g1289) & (!g1292) & (sk[26]) & (!g1293) & (!g1295)) + ((!g1288) & (g1289) & (!g1292) & (sk[26]) & (g1293) & (g1295)) + ((!g1288) & (g1289) & (g1292) & (!sk[26]) & (!g1293) & (!g1295)) + ((!g1288) & (g1289) & (g1292) & (!sk[26]) & (!g1293) & (g1295)) + ((!g1288) & (g1289) & (g1292) & (!sk[26]) & (g1293) & (!g1295)) + ((!g1288) & (g1289) & (g1292) & (!sk[26]) & (g1293) & (g1295)) + ((!g1288) & (g1289) & (g1292) & (sk[26]) & (!g1293) & (g1295)) + ((!g1288) & (g1289) & (g1292) & (sk[26]) & (g1293) & (!g1295)) + ((g1288) & (!g1289) & (!g1292) & (!sk[26]) & (g1293) & (!g1295)) + ((g1288) & (!g1289) & (!g1292) & (!sk[26]) & (g1293) & (g1295)) + ((g1288) & (!g1289) & (!g1292) & (sk[26]) & (!g1293) & (!g1295)) + ((g1288) & (!g1289) & (!g1292) & (sk[26]) & (g1293) & (g1295)) + ((g1288) & (!g1289) & (g1292) & (!sk[26]) & (!g1293) & (!g1295)) + ((g1288) & (!g1289) & (g1292) & (!sk[26]) & (!g1293) & (g1295)) + ((g1288) & (!g1289) & (g1292) & (!sk[26]) & (g1293) & (!g1295)) + ((g1288) & (!g1289) & (g1292) & (!sk[26]) & (g1293) & (g1295)) + ((g1288) & (!g1289) & (g1292) & (sk[26]) & (!g1293) & (g1295)) + ((g1288) & (!g1289) & (g1292) & (sk[26]) & (g1293) & (!g1295)) + ((g1288) & (g1289) & (!g1292) & (!sk[26]) & (!g1293) & (!g1295)) + ((g1288) & (g1289) & (!g1292) & (!sk[26]) & (!g1293) & (g1295)) + ((g1288) & (g1289) & (!g1292) & (!sk[26]) & (g1293) & (!g1295)) + ((g1288) & (g1289) & (!g1292) & (!sk[26]) & (g1293) & (g1295)) + ((g1288) & (g1289) & (!g1292) & (sk[26]) & (!g1293) & (g1295)) + ((g1288) & (g1289) & (!g1292) & (sk[26]) & (g1293) & (!g1295)) + ((g1288) & (g1289) & (g1292) & (!sk[26]) & (!g1293) & (!g1295)) + ((g1288) & (g1289) & (g1292) & (!sk[26]) & (!g1293) & (g1295)) + ((g1288) & (g1289) & (g1292) & (!sk[26]) & (g1293) & (!g1295)) + ((g1288) & (g1289) & (g1292) & (!sk[26]) & (g1293) & (g1295)) + ((g1288) & (g1289) & (g1292) & (sk[26]) & (!g1293) & (!g1295)) + ((g1288) & (g1289) & (g1292) & (sk[26]) & (g1293) & (g1295)));
	assign g1297 = (((!g1286) & (!g1287) & (sk[27]) & (!g1296)) + ((!g1286) & (g1287) & (!sk[27]) & (!g1296)) + ((!g1286) & (g1287) & (!sk[27]) & (g1296)) + ((!g1286) & (g1287) & (sk[27]) & (g1296)) + ((g1286) & (!g1287) & (sk[27]) & (g1296)) + ((g1286) & (g1287) & (!sk[27]) & (!g1296)) + ((g1286) & (g1287) & (!sk[27]) & (g1296)) + ((g1286) & (g1287) & (sk[27]) & (!g1296)));
	assign g1298 = (((!g38) & (!g17) & (!sk[28]) & (!g30) & (g62) & (!g46)) + ((!g38) & (!g17) & (!sk[28]) & (!g30) & (g62) & (g46)) + ((!g38) & (!g17) & (!sk[28]) & (g30) & (!g62) & (!g46)) + ((!g38) & (!g17) & (!sk[28]) & (g30) & (!g62) & (g46)) + ((!g38) & (!g17) & (!sk[28]) & (g30) & (g62) & (!g46)) + ((!g38) & (!g17) & (!sk[28]) & (g30) & (g62) & (g46)) + ((!g38) & (!g17) & (sk[28]) & (!g30) & (!g62) & (!g46)) + ((!g38) & (!g17) & (sk[28]) & (!g30) & (!g62) & (g46)) + ((!g38) & (!g17) & (sk[28]) & (!g30) & (g62) & (!g46)) + ((!g38) & (!g17) & (sk[28]) & (!g30) & (g62) & (g46)) + ((!g38) & (!g17) & (sk[28]) & (g30) & (!g62) & (!g46)) + ((!g38) & (!g17) & (sk[28]) & (g30) & (!g62) & (g46)) + ((!g38) & (g17) & (!sk[28]) & (!g30) & (!g62) & (!g46)) + ((!g38) & (g17) & (!sk[28]) & (!g30) & (!g62) & (g46)) + ((!g38) & (g17) & (!sk[28]) & (!g30) & (g62) & (!g46)) + ((!g38) & (g17) & (!sk[28]) & (!g30) & (g62) & (g46)) + ((!g38) & (g17) & (!sk[28]) & (g30) & (!g62) & (!g46)) + ((!g38) & (g17) & (!sk[28]) & (g30) & (!g62) & (g46)) + ((!g38) & (g17) & (!sk[28]) & (g30) & (g62) & (!g46)) + ((!g38) & (g17) & (!sk[28]) & (g30) & (g62) & (g46)) + ((!g38) & (g17) & (sk[28]) & (!g30) & (!g62) & (!g46)) + ((!g38) & (g17) & (sk[28]) & (!g30) & (g62) & (!g46)) + ((!g38) & (g17) & (sk[28]) & (g30) & (!g62) & (!g46)) + ((g38) & (!g17) & (!sk[28]) & (!g30) & (g62) & (!g46)) + ((g38) & (!g17) & (!sk[28]) & (!g30) & (g62) & (g46)) + ((g38) & (!g17) & (!sk[28]) & (g30) & (!g62) & (!g46)) + ((g38) & (!g17) & (!sk[28]) & (g30) & (!g62) & (g46)) + ((g38) & (!g17) & (!sk[28]) & (g30) & (g62) & (!g46)) + ((g38) & (!g17) & (!sk[28]) & (g30) & (g62) & (g46)) + ((g38) & (!g17) & (sk[28]) & (!g30) & (!g62) & (!g46)) + ((g38) & (!g17) & (sk[28]) & (!g30) & (!g62) & (g46)) + ((g38) & (!g17) & (sk[28]) & (g30) & (!g62) & (!g46)) + ((g38) & (!g17) & (sk[28]) & (g30) & (!g62) & (g46)) + ((g38) & (g17) & (!sk[28]) & (!g30) & (!g62) & (!g46)) + ((g38) & (g17) & (!sk[28]) & (!g30) & (!g62) & (g46)) + ((g38) & (g17) & (!sk[28]) & (!g30) & (g62) & (!g46)) + ((g38) & (g17) & (!sk[28]) & (!g30) & (g62) & (g46)) + ((g38) & (g17) & (!sk[28]) & (g30) & (!g62) & (!g46)) + ((g38) & (g17) & (!sk[28]) & (g30) & (!g62) & (g46)) + ((g38) & (g17) & (!sk[28]) & (g30) & (g62) & (!g46)) + ((g38) & (g17) & (!sk[28]) & (g30) & (g62) & (g46)) + ((g38) & (g17) & (sk[28]) & (!g30) & (!g62) & (!g46)) + ((g38) & (g17) & (sk[28]) & (g30) & (!g62) & (!g46)));
	assign g1299 = (((!sk[29]) & (!g99) & (!g40) & (!g590) & (g1298)) + ((!sk[29]) & (!g99) & (!g40) & (g590) & (g1298)) + ((!sk[29]) & (!g99) & (g40) & (!g590) & (g1298)) + ((!sk[29]) & (!g99) & (g40) & (g590) & (g1298)) + ((!sk[29]) & (g99) & (!g40) & (!g590) & (!g1298)) + ((!sk[29]) & (g99) & (!g40) & (!g590) & (g1298)) + ((!sk[29]) & (g99) & (!g40) & (g590) & (!g1298)) + ((!sk[29]) & (g99) & (!g40) & (g590) & (g1298)) + ((!sk[29]) & (g99) & (g40) & (!g590) & (!g1298)) + ((!sk[29]) & (g99) & (g40) & (!g590) & (g1298)) + ((!sk[29]) & (g99) & (g40) & (g590) & (!g1298)) + ((!sk[29]) & (g99) & (g40) & (g590) & (g1298)) + ((sk[29]) & (!g99) & (!g40) & (g590) & (g1298)) + ((sk[29]) & (!g99) & (g40) & (g590) & (g1298)) + ((sk[29]) & (g99) & (!g40) & (g590) & (g1298)));
	assign g1300 = (((!g268) & (!g82) & (!sk[30]) & (!g876) & (g1299)) + ((!g268) & (!g82) & (!sk[30]) & (g876) & (g1299)) + ((!g268) & (g82) & (!sk[30]) & (!g876) & (g1299)) + ((!g268) & (g82) & (!sk[30]) & (g876) & (g1299)) + ((!g268) & (g82) & (sk[30]) & (g876) & (g1299)) + ((g268) & (!g82) & (!sk[30]) & (!g876) & (!g1299)) + ((g268) & (!g82) & (!sk[30]) & (!g876) & (g1299)) + ((g268) & (!g82) & (!sk[30]) & (g876) & (!g1299)) + ((g268) & (!g82) & (!sk[30]) & (g876) & (g1299)) + ((g268) & (g82) & (!sk[30]) & (!g876) & (!g1299)) + ((g268) & (g82) & (!sk[30]) & (!g876) & (g1299)) + ((g268) & (g82) & (!sk[30]) & (g876) & (!g1299)) + ((g268) & (g82) & (!sk[30]) & (g876) & (g1299)));
	assign g1301 = (((!g55) & (!g647) & (!g967) & (g1007) & (!sk[31]) & (!g1300)) + ((!g55) & (!g647) & (!g967) & (g1007) & (!sk[31]) & (g1300)) + ((!g55) & (!g647) & (g967) & (!g1007) & (!sk[31]) & (!g1300)) + ((!g55) & (!g647) & (g967) & (!g1007) & (!sk[31]) & (g1300)) + ((!g55) & (!g647) & (g967) & (g1007) & (!sk[31]) & (!g1300)) + ((!g55) & (!g647) & (g967) & (g1007) & (!sk[31]) & (g1300)) + ((!g55) & (g647) & (!g967) & (!g1007) & (!sk[31]) & (!g1300)) + ((!g55) & (g647) & (!g967) & (!g1007) & (!sk[31]) & (g1300)) + ((!g55) & (g647) & (!g967) & (g1007) & (!sk[31]) & (!g1300)) + ((!g55) & (g647) & (!g967) & (g1007) & (!sk[31]) & (g1300)) + ((!g55) & (g647) & (!g967) & (g1007) & (sk[31]) & (g1300)) + ((!g55) & (g647) & (g967) & (!g1007) & (!sk[31]) & (!g1300)) + ((!g55) & (g647) & (g967) & (!g1007) & (!sk[31]) & (g1300)) + ((!g55) & (g647) & (g967) & (g1007) & (!sk[31]) & (!g1300)) + ((!g55) & (g647) & (g967) & (g1007) & (!sk[31]) & (g1300)) + ((g55) & (!g647) & (!g967) & (g1007) & (!sk[31]) & (!g1300)) + ((g55) & (!g647) & (!g967) & (g1007) & (!sk[31]) & (g1300)) + ((g55) & (!g647) & (g967) & (!g1007) & (!sk[31]) & (!g1300)) + ((g55) & (!g647) & (g967) & (!g1007) & (!sk[31]) & (g1300)) + ((g55) & (!g647) & (g967) & (g1007) & (!sk[31]) & (!g1300)) + ((g55) & (!g647) & (g967) & (g1007) & (!sk[31]) & (g1300)) + ((g55) & (g647) & (!g967) & (!g1007) & (!sk[31]) & (!g1300)) + ((g55) & (g647) & (!g967) & (!g1007) & (!sk[31]) & (g1300)) + ((g55) & (g647) & (!g967) & (g1007) & (!sk[31]) & (!g1300)) + ((g55) & (g647) & (!g967) & (g1007) & (!sk[31]) & (g1300)) + ((g55) & (g647) & (g967) & (!g1007) & (!sk[31]) & (!g1300)) + ((g55) & (g647) & (g967) & (!g1007) & (!sk[31]) & (g1300)) + ((g55) & (g647) & (g967) & (g1007) & (!sk[31]) & (!g1300)) + ((g55) & (g647) & (g967) & (g1007) & (!sk[31]) & (g1300)));
	assign g1302 = (((!sk[32]) & (!g1284) & (!g1285) & (!g1297) & (g1301)) + ((!sk[32]) & (!g1284) & (!g1285) & (g1297) & (g1301)) + ((!sk[32]) & (!g1284) & (g1285) & (!g1297) & (g1301)) + ((!sk[32]) & (!g1284) & (g1285) & (g1297) & (g1301)) + ((!sk[32]) & (g1284) & (!g1285) & (!g1297) & (!g1301)) + ((!sk[32]) & (g1284) & (!g1285) & (!g1297) & (g1301)) + ((!sk[32]) & (g1284) & (!g1285) & (g1297) & (!g1301)) + ((!sk[32]) & (g1284) & (!g1285) & (g1297) & (g1301)) + ((!sk[32]) & (g1284) & (g1285) & (!g1297) & (!g1301)) + ((!sk[32]) & (g1284) & (g1285) & (!g1297) & (g1301)) + ((!sk[32]) & (g1284) & (g1285) & (g1297) & (!g1301)) + ((!sk[32]) & (g1284) & (g1285) & (g1297) & (g1301)) + ((sk[32]) & (!g1284) & (!g1285) & (!g1297) & (!g1301)) + ((sk[32]) & (!g1284) & (!g1285) & (g1297) & (g1301)) + ((sk[32]) & (!g1284) & (g1285) & (!g1297) & (g1301)) + ((sk[32]) & (!g1284) & (g1285) & (g1297) & (!g1301)) + ((sk[32]) & (g1284) & (!g1285) & (!g1297) & (g1301)) + ((sk[32]) & (g1284) & (!g1285) & (g1297) & (!g1301)) + ((sk[32]) & (g1284) & (g1285) & (!g1297) & (g1301)) + ((sk[32]) & (g1284) & (g1285) & (g1297) & (!g1301)));
	assign g1303 = (((!sk[33]) & (!g1068) & (!g1281) & (!g1283) & (g1302)) + ((!sk[33]) & (!g1068) & (!g1281) & (g1283) & (g1302)) + ((!sk[33]) & (!g1068) & (g1281) & (!g1283) & (g1302)) + ((!sk[33]) & (!g1068) & (g1281) & (g1283) & (g1302)) + ((!sk[33]) & (g1068) & (!g1281) & (!g1283) & (!g1302)) + ((!sk[33]) & (g1068) & (!g1281) & (!g1283) & (g1302)) + ((!sk[33]) & (g1068) & (!g1281) & (g1283) & (!g1302)) + ((!sk[33]) & (g1068) & (!g1281) & (g1283) & (g1302)) + ((!sk[33]) & (g1068) & (g1281) & (!g1283) & (!g1302)) + ((!sk[33]) & (g1068) & (g1281) & (!g1283) & (g1302)) + ((!sk[33]) & (g1068) & (g1281) & (g1283) & (!g1302)) + ((!sk[33]) & (g1068) & (g1281) & (g1283) & (g1302)) + ((sk[33]) & (!g1068) & (!g1281) & (!g1283) & (g1302)) + ((sk[33]) & (!g1068) & (!g1281) & (g1283) & (!g1302)) + ((sk[33]) & (!g1068) & (g1281) & (!g1283) & (g1302)) + ((sk[33]) & (!g1068) & (g1281) & (g1283) & (!g1302)) + ((sk[33]) & (g1068) & (!g1281) & (!g1283) & (!g1302)) + ((sk[33]) & (g1068) & (!g1281) & (g1283) & (g1302)) + ((sk[33]) & (g1068) & (g1281) & (!g1283) & (g1302)) + ((sk[33]) & (g1068) & (g1281) & (g1283) & (!g1302)));
	assign g1304 = (((!sk[34]) & (!g1284) & (!g1285) & (!g1297) & (g1301)) + ((!sk[34]) & (!g1284) & (!g1285) & (g1297) & (g1301)) + ((!sk[34]) & (!g1284) & (g1285) & (!g1297) & (g1301)) + ((!sk[34]) & (!g1284) & (g1285) & (g1297) & (g1301)) + ((!sk[34]) & (g1284) & (!g1285) & (!g1297) & (!g1301)) + ((!sk[34]) & (g1284) & (!g1285) & (!g1297) & (g1301)) + ((!sk[34]) & (g1284) & (!g1285) & (g1297) & (!g1301)) + ((!sk[34]) & (g1284) & (!g1285) & (g1297) & (g1301)) + ((!sk[34]) & (g1284) & (g1285) & (!g1297) & (!g1301)) + ((!sk[34]) & (g1284) & (g1285) & (!g1297) & (g1301)) + ((!sk[34]) & (g1284) & (g1285) & (g1297) & (!g1301)) + ((!sk[34]) & (g1284) & (g1285) & (g1297) & (g1301)) + ((sk[34]) & (!g1284) & (!g1285) & (!g1297) & (g1301)) + ((sk[34]) & (!g1284) & (!g1285) & (g1297) & (!g1301)) + ((sk[34]) & (!g1284) & (!g1285) & (g1297) & (g1301)) + ((sk[34]) & (!g1284) & (g1285) & (g1297) & (g1301)) + ((sk[34]) & (g1284) & (!g1285) & (g1297) & (g1301)) + ((sk[34]) & (g1284) & (g1285) & (g1297) & (g1301)));
	assign g1305 = (((!g1288) & (!g1289) & (!g1292) & (!sk[35]) & (g1293) & (!g1295)) + ((!g1288) & (!g1289) & (!g1292) & (!sk[35]) & (g1293) & (g1295)) + ((!g1288) & (!g1289) & (g1292) & (!sk[35]) & (!g1293) & (!g1295)) + ((!g1288) & (!g1289) & (g1292) & (!sk[35]) & (!g1293) & (g1295)) + ((!g1288) & (!g1289) & (g1292) & (!sk[35]) & (g1293) & (!g1295)) + ((!g1288) & (!g1289) & (g1292) & (!sk[35]) & (g1293) & (g1295)) + ((!g1288) & (g1289) & (!g1292) & (!sk[35]) & (!g1293) & (!g1295)) + ((!g1288) & (g1289) & (!g1292) & (!sk[35]) & (!g1293) & (g1295)) + ((!g1288) & (g1289) & (!g1292) & (!sk[35]) & (g1293) & (!g1295)) + ((!g1288) & (g1289) & (!g1292) & (!sk[35]) & (g1293) & (g1295)) + ((!g1288) & (g1289) & (!g1292) & (sk[35]) & (!g1293) & (!g1295)) + ((!g1288) & (g1289) & (!g1292) & (sk[35]) & (g1293) & (g1295)) + ((!g1288) & (g1289) & (g1292) & (!sk[35]) & (!g1293) & (!g1295)) + ((!g1288) & (g1289) & (g1292) & (!sk[35]) & (!g1293) & (g1295)) + ((!g1288) & (g1289) & (g1292) & (!sk[35]) & (g1293) & (!g1295)) + ((!g1288) & (g1289) & (g1292) & (!sk[35]) & (g1293) & (g1295)) + ((!g1288) & (g1289) & (g1292) & (sk[35]) & (!g1293) & (g1295)) + ((!g1288) & (g1289) & (g1292) & (sk[35]) & (g1293) & (!g1295)) + ((g1288) & (!g1289) & (!g1292) & (!sk[35]) & (g1293) & (!g1295)) + ((g1288) & (!g1289) & (!g1292) & (!sk[35]) & (g1293) & (g1295)) + ((g1288) & (!g1289) & (!g1292) & (sk[35]) & (!g1293) & (!g1295)) + ((g1288) & (!g1289) & (!g1292) & (sk[35]) & (g1293) & (g1295)) + ((g1288) & (!g1289) & (g1292) & (!sk[35]) & (!g1293) & (!g1295)) + ((g1288) & (!g1289) & (g1292) & (!sk[35]) & (!g1293) & (g1295)) + ((g1288) & (!g1289) & (g1292) & (!sk[35]) & (g1293) & (!g1295)) + ((g1288) & (!g1289) & (g1292) & (!sk[35]) & (g1293) & (g1295)) + ((g1288) & (!g1289) & (g1292) & (sk[35]) & (!g1293) & (g1295)) + ((g1288) & (!g1289) & (g1292) & (sk[35]) & (g1293) & (!g1295)) + ((g1288) & (g1289) & (!g1292) & (!sk[35]) & (!g1293) & (!g1295)) + ((g1288) & (g1289) & (!g1292) & (!sk[35]) & (!g1293) & (g1295)) + ((g1288) & (g1289) & (!g1292) & (!sk[35]) & (g1293) & (!g1295)) + ((g1288) & (g1289) & (!g1292) & (!sk[35]) & (g1293) & (g1295)) + ((g1288) & (g1289) & (!g1292) & (sk[35]) & (!g1293) & (!g1295)) + ((g1288) & (g1289) & (!g1292) & (sk[35]) & (!g1293) & (g1295)) + ((g1288) & (g1289) & (!g1292) & (sk[35]) & (g1293) & (!g1295)) + ((g1288) & (g1289) & (!g1292) & (sk[35]) & (g1293) & (g1295)) + ((g1288) & (g1289) & (g1292) & (!sk[35]) & (!g1293) & (!g1295)) + ((g1288) & (g1289) & (g1292) & (!sk[35]) & (!g1293) & (g1295)) + ((g1288) & (g1289) & (g1292) & (!sk[35]) & (g1293) & (!g1295)) + ((g1288) & (g1289) & (g1292) & (!sk[35]) & (g1293) & (g1295)) + ((g1288) & (g1289) & (g1292) & (sk[35]) & (!g1293) & (!g1295)) + ((g1288) & (g1289) & (g1292) & (sk[35]) & (!g1293) & (g1295)) + ((g1288) & (g1289) & (g1292) & (sk[35]) & (g1293) & (!g1295)) + ((g1288) & (g1289) & (g1292) & (sk[35]) & (g1293) & (g1295)));
	assign g1306 = (((!g847) & (!g845) & (!g848) & (!g962) & (!g963) & (!g971)) + ((!g847) & (!g845) & (!g848) & (!g962) & (!g963) & (g971)) + ((!g847) & (!g845) & (!g848) & (!g962) & (g963) & (!g971)) + ((!g847) & (!g845) & (!g848) & (!g962) & (g963) & (g971)) + ((!g847) & (!g845) & (!g848) & (g962) & (!g963) & (!g971)) + ((!g847) & (!g845) & (!g848) & (g962) & (!g963) & (g971)) + ((!g847) & (!g845) & (!g848) & (g962) & (g963) & (!g971)) + ((!g847) & (!g845) & (!g848) & (g962) & (g963) & (g971)) + ((!g847) & (!g845) & (g848) & (!g962) & (!g963) & (!g971)) + ((!g847) & (!g845) & (g848) & (!g962) & (!g963) & (g971)) + ((!g847) & (!g845) & (g848) & (g962) & (!g963) & (!g971)) + ((!g847) & (!g845) & (g848) & (g962) & (!g963) & (g971)) + ((!g847) & (g845) & (!g848) & (g962) & (!g963) & (!g971)) + ((!g847) & (g845) & (!g848) & (g962) & (!g963) & (g971)) + ((!g847) & (g845) & (!g848) & (g962) & (g963) & (!g971)) + ((!g847) & (g845) & (!g848) & (g962) & (g963) & (g971)) + ((!g847) & (g845) & (g848) & (g962) & (!g963) & (!g971)) + ((!g847) & (g845) & (g848) & (g962) & (!g963) & (g971)) + ((g847) & (!g845) & (!g848) & (!g962) & (!g963) & (!g971)) + ((g847) & (!g845) & (!g848) & (!g962) & (g963) & (!g971)) + ((g847) & (!g845) & (!g848) & (g962) & (!g963) & (!g971)) + ((g847) & (!g845) & (!g848) & (g962) & (g963) & (!g971)) + ((g847) & (!g845) & (g848) & (!g962) & (!g963) & (!g971)) + ((g847) & (!g845) & (g848) & (g962) & (!g963) & (!g971)) + ((g847) & (g845) & (!g848) & (g962) & (!g963) & (!g971)) + ((g847) & (g845) & (!g848) & (g962) & (g963) & (!g971)) + ((g847) & (g845) & (g848) & (g962) & (!g963) & (!g971)));
	assign g1307 = (((!g252) & (!g843) & (!sk[37]) & (!g972) & (g1306)) + ((!g252) & (!g843) & (!sk[37]) & (g972) & (g1306)) + ((!g252) & (!g843) & (sk[37]) & (!g972) & (!g1306)) + ((!g252) & (!g843) & (sk[37]) & (g972) & (!g1306)) + ((!g252) & (g843) & (!sk[37]) & (!g972) & (g1306)) + ((!g252) & (g843) & (!sk[37]) & (g972) & (g1306)) + ((!g252) & (g843) & (sk[37]) & (!g972) & (!g1306)) + ((!g252) & (g843) & (sk[37]) & (!g972) & (g1306)) + ((!g252) & (g843) & (sk[37]) & (g972) & (!g1306)) + ((g252) & (!g843) & (!sk[37]) & (!g972) & (!g1306)) + ((g252) & (!g843) & (!sk[37]) & (!g972) & (g1306)) + ((g252) & (!g843) & (!sk[37]) & (g972) & (!g1306)) + ((g252) & (!g843) & (!sk[37]) & (g972) & (g1306)) + ((g252) & (!g843) & (sk[37]) & (!g972) & (g1306)) + ((g252) & (!g843) & (sk[37]) & (g972) & (g1306)) + ((g252) & (g843) & (!sk[37]) & (!g972) & (!g1306)) + ((g252) & (g843) & (!sk[37]) & (!g972) & (g1306)) + ((g252) & (g843) & (!sk[37]) & (g972) & (!g1306)) + ((g252) & (g843) & (!sk[37]) & (g972) & (g1306)) + ((g252) & (g843) & (sk[37]) & (g972) & (g1306)));
	assign g1308 = (((!g252) & (!sk[38]) & (!g200) & (!g869) & (g863)) + ((!g252) & (!sk[38]) & (!g200) & (g869) & (g863)) + ((!g252) & (!sk[38]) & (g200) & (!g869) & (g863)) + ((!g252) & (!sk[38]) & (g200) & (g869) & (g863)) + ((!g252) & (sk[38]) & (!g200) & (!g869) & (!g863)) + ((!g252) & (sk[38]) & (!g200) & (!g869) & (g863)) + ((!g252) & (sk[38]) & (!g200) & (g869) & (!g863)) + ((!g252) & (sk[38]) & (!g200) & (g869) & (g863)) + ((g252) & (!sk[38]) & (!g200) & (!g869) & (!g863)) + ((g252) & (!sk[38]) & (!g200) & (!g869) & (g863)) + ((g252) & (!sk[38]) & (!g200) & (g869) & (!g863)) + ((g252) & (!sk[38]) & (!g200) & (g869) & (g863)) + ((g252) & (!sk[38]) & (g200) & (!g869) & (!g863)) + ((g252) & (!sk[38]) & (g200) & (!g869) & (g863)) + ((g252) & (!sk[38]) & (g200) & (g869) & (!g863)) + ((g252) & (!sk[38]) & (g200) & (g869) & (g863)) + ((g252) & (sk[38]) & (!g200) & (!g869) & (!g863)) + ((g252) & (sk[38]) & (!g200) & (g869) & (g863)) + ((g252) & (sk[38]) & (g200) & (!g869) & (g863)) + ((g252) & (sk[38]) & (g200) & (g869) & (!g863)));
	assign g1309 = (((!g252) & (!g869) & (!g870) & (!g1290) & (!g1291) & (!g1308)) + ((!g252) & (!g869) & (!g870) & (!g1290) & (g1291) & (g1308)) + ((!g252) & (!g869) & (!g870) & (g1290) & (!g1291) & (!g1308)) + ((!g252) & (!g869) & (!g870) & (g1290) & (g1291) & (!g1308)) + ((!g252) & (!g869) & (g870) & (!g1290) & (!g1291) & (!g1308)) + ((!g252) & (!g869) & (g870) & (!g1290) & (g1291) & (g1308)) + ((!g252) & (!g869) & (g870) & (g1290) & (!g1291) & (!g1308)) + ((!g252) & (!g869) & (g870) & (g1290) & (g1291) & (!g1308)) + ((!g252) & (g869) & (!g870) & (!g1290) & (!g1291) & (!g1308)) + ((!g252) & (g869) & (!g870) & (!g1290) & (g1291) & (g1308)) + ((!g252) & (g869) & (!g870) & (g1290) & (!g1291) & (!g1308)) + ((!g252) & (g869) & (!g870) & (g1290) & (g1291) & (!g1308)) + ((!g252) & (g869) & (g870) & (!g1290) & (!g1291) & (!g1308)) + ((!g252) & (g869) & (g870) & (!g1290) & (g1291) & (g1308)) + ((!g252) & (g869) & (g870) & (g1290) & (!g1291) & (!g1308)) + ((!g252) & (g869) & (g870) & (g1290) & (g1291) & (!g1308)) + ((g252) & (!g869) & (!g870) & (!g1290) & (!g1291) & (!g1308)) + ((g252) & (!g869) & (!g870) & (!g1290) & (g1291) & (!g1308)) + ((g252) & (!g869) & (!g870) & (g1290) & (!g1291) & (!g1308)) + ((g252) & (!g869) & (!g870) & (g1290) & (g1291) & (!g1308)) + ((g252) & (!g869) & (g870) & (!g1290) & (!g1291) & (g1308)) + ((g252) & (!g869) & (g870) & (!g1290) & (g1291) & (!g1308)) + ((g252) & (!g869) & (g870) & (g1290) & (!g1291) & (g1308)) + ((g252) & (!g869) & (g870) & (g1290) & (g1291) & (g1308)) + ((g252) & (g869) & (!g870) & (!g1290) & (!g1291) & (g1308)) + ((g252) & (g869) & (!g870) & (!g1290) & (g1291) & (!g1308)) + ((g252) & (g869) & (!g870) & (g1290) & (!g1291) & (g1308)) + ((g252) & (g869) & (!g870) & (g1290) & (g1291) & (g1308)) + ((g252) & (g869) & (g870) & (!g1290) & (!g1291) & (g1308)) + ((g252) & (g869) & (g870) & (!g1290) & (g1291) & (g1308)) + ((g252) & (g869) & (g870) & (g1290) & (!g1291) & (g1308)) + ((g252) & (g869) & (g870) & (g1290) & (g1291) & (g1308)));
	assign g1310 = (((!g764) & (!g762) & (!g765) & (!g994) & (!g1040) & (!g1079)) + ((!g764) & (!g762) & (!g765) & (!g994) & (!g1040) & (g1079)) + ((!g764) & (!g762) & (!g765) & (!g994) & (g1040) & (!g1079)) + ((!g764) & (!g762) & (!g765) & (!g994) & (g1040) & (g1079)) + ((!g764) & (!g762) & (!g765) & (g994) & (!g1040) & (!g1079)) + ((!g764) & (!g762) & (!g765) & (g994) & (!g1040) & (g1079)) + ((!g764) & (!g762) & (!g765) & (g994) & (g1040) & (!g1079)) + ((!g764) & (!g762) & (!g765) & (g994) & (g1040) & (g1079)) + ((!g764) & (!g762) & (g765) & (!g994) & (!g1040) & (!g1079)) + ((!g764) & (!g762) & (g765) & (!g994) & (!g1040) & (g1079)) + ((!g764) & (!g762) & (g765) & (!g994) & (g1040) & (!g1079)) + ((!g764) & (!g762) & (g765) & (!g994) & (g1040) & (g1079)) + ((!g764) & (g762) & (!g765) & (!g994) & (g1040) & (!g1079)) + ((!g764) & (g762) & (!g765) & (!g994) & (g1040) & (g1079)) + ((!g764) & (g762) & (!g765) & (g994) & (g1040) & (!g1079)) + ((!g764) & (g762) & (!g765) & (g994) & (g1040) & (g1079)) + ((!g764) & (g762) & (g765) & (!g994) & (g1040) & (!g1079)) + ((!g764) & (g762) & (g765) & (!g994) & (g1040) & (g1079)) + ((g764) & (!g762) & (!g765) & (!g994) & (!g1040) & (g1079)) + ((g764) & (!g762) & (!g765) & (!g994) & (g1040) & (g1079)) + ((g764) & (!g762) & (!g765) & (g994) & (!g1040) & (g1079)) + ((g764) & (!g762) & (!g765) & (g994) & (g1040) & (g1079)) + ((g764) & (!g762) & (g765) & (!g994) & (!g1040) & (g1079)) + ((g764) & (!g762) & (g765) & (!g994) & (g1040) & (g1079)) + ((g764) & (g762) & (!g765) & (!g994) & (g1040) & (g1079)) + ((g764) & (g762) & (!g765) & (g994) & (g1040) & (g1079)) + ((g764) & (g762) & (g765) & (!g994) & (g1040) & (g1079)));
	assign g1311 = (((!g202) & (!g759) & (!g1040) & (!g1079) & (!g1080) & (g1310)) + ((!g202) & (!g759) & (!g1040) & (!g1079) & (g1080) & (g1310)) + ((!g202) & (!g759) & (!g1040) & (g1079) & (!g1080) & (g1310)) + ((!g202) & (!g759) & (!g1040) & (g1079) & (g1080) & (g1310)) + ((!g202) & (!g759) & (g1040) & (!g1079) & (!g1080) & (g1310)) + ((!g202) & (!g759) & (g1040) & (!g1079) & (g1080) & (g1310)) + ((!g202) & (!g759) & (g1040) & (g1079) & (!g1080) & (g1310)) + ((!g202) & (!g759) & (g1040) & (g1079) & (g1080) & (g1310)) + ((!g202) & (g759) & (!g1040) & (!g1079) & (!g1080) & (g1310)) + ((!g202) & (g759) & (!g1040) & (g1079) & (g1080) & (g1310)) + ((!g202) & (g759) & (g1040) & (!g1079) & (g1080) & (g1310)) + ((!g202) & (g759) & (g1040) & (g1079) & (!g1080) & (g1310)) + ((g202) & (!g759) & (!g1040) & (!g1079) & (!g1080) & (!g1310)) + ((g202) & (!g759) & (!g1040) & (!g1079) & (g1080) & (!g1310)) + ((g202) & (!g759) & (!g1040) & (g1079) & (!g1080) & (!g1310)) + ((g202) & (!g759) & (!g1040) & (g1079) & (g1080) & (!g1310)) + ((g202) & (!g759) & (g1040) & (!g1079) & (!g1080) & (!g1310)) + ((g202) & (!g759) & (g1040) & (!g1079) & (g1080) & (!g1310)) + ((g202) & (!g759) & (g1040) & (g1079) & (!g1080) & (!g1310)) + ((g202) & (!g759) & (g1040) & (g1079) & (g1080) & (!g1310)) + ((g202) & (g759) & (!g1040) & (!g1079) & (!g1080) & (!g1310)) + ((g202) & (g759) & (!g1040) & (!g1079) & (g1080) & (!g1310)) + ((g202) & (g759) & (!g1040) & (!g1079) & (g1080) & (g1310)) + ((g202) & (g759) & (!g1040) & (g1079) & (!g1080) & (!g1310)) + ((g202) & (g759) & (!g1040) & (g1079) & (!g1080) & (g1310)) + ((g202) & (g759) & (!g1040) & (g1079) & (g1080) & (!g1310)) + ((g202) & (g759) & (g1040) & (!g1079) & (!g1080) & (!g1310)) + ((g202) & (g759) & (g1040) & (!g1079) & (!g1080) & (g1310)) + ((g202) & (g759) & (g1040) & (!g1079) & (g1080) & (!g1310)) + ((g202) & (g759) & (g1040) & (g1079) & (!g1080) & (!g1310)) + ((g202) & (g759) & (g1040) & (g1079) & (g1080) & (!g1310)) + ((g202) & (g759) & (g1040) & (g1079) & (g1080) & (g1310)));
	assign g1312 = (((!g1292) & (!g1293) & (!g1295) & (!g1307) & (!g1309) & (!g1311)) + ((!g1292) & (!g1293) & (!g1295) & (!g1307) & (g1309) & (g1311)) + ((!g1292) & (!g1293) & (!g1295) & (g1307) & (!g1309) & (g1311)) + ((!g1292) & (!g1293) & (!g1295) & (g1307) & (g1309) & (!g1311)) + ((!g1292) & (!g1293) & (g1295) & (!g1307) & (!g1309) & (g1311)) + ((!g1292) & (!g1293) & (g1295) & (!g1307) & (g1309) & (!g1311)) + ((!g1292) & (!g1293) & (g1295) & (g1307) & (!g1309) & (!g1311)) + ((!g1292) & (!g1293) & (g1295) & (g1307) & (g1309) & (g1311)) + ((!g1292) & (g1293) & (!g1295) & (!g1307) & (!g1309) & (!g1311)) + ((!g1292) & (g1293) & (!g1295) & (!g1307) & (g1309) & (g1311)) + ((!g1292) & (g1293) & (!g1295) & (g1307) & (!g1309) & (g1311)) + ((!g1292) & (g1293) & (!g1295) & (g1307) & (g1309) & (!g1311)) + ((!g1292) & (g1293) & (g1295) & (!g1307) & (!g1309) & (!g1311)) + ((!g1292) & (g1293) & (g1295) & (!g1307) & (g1309) & (g1311)) + ((!g1292) & (g1293) & (g1295) & (g1307) & (!g1309) & (g1311)) + ((!g1292) & (g1293) & (g1295) & (g1307) & (g1309) & (!g1311)) + ((g1292) & (!g1293) & (!g1295) & (!g1307) & (!g1309) & (g1311)) + ((g1292) & (!g1293) & (!g1295) & (!g1307) & (g1309) & (!g1311)) + ((g1292) & (!g1293) & (!g1295) & (g1307) & (!g1309) & (!g1311)) + ((g1292) & (!g1293) & (!g1295) & (g1307) & (g1309) & (g1311)) + ((g1292) & (!g1293) & (g1295) & (!g1307) & (!g1309) & (g1311)) + ((g1292) & (!g1293) & (g1295) & (!g1307) & (g1309) & (!g1311)) + ((g1292) & (!g1293) & (g1295) & (g1307) & (!g1309) & (!g1311)) + ((g1292) & (!g1293) & (g1295) & (g1307) & (g1309) & (g1311)) + ((g1292) & (g1293) & (!g1295) & (!g1307) & (!g1309) & (!g1311)) + ((g1292) & (g1293) & (!g1295) & (!g1307) & (g1309) & (g1311)) + ((g1292) & (g1293) & (!g1295) & (g1307) & (!g1309) & (g1311)) + ((g1292) & (g1293) & (!g1295) & (g1307) & (g1309) & (!g1311)) + ((g1292) & (g1293) & (g1295) & (!g1307) & (!g1309) & (g1311)) + ((g1292) & (g1293) & (g1295) & (!g1307) & (g1309) & (!g1311)) + ((g1292) & (g1293) & (g1295) & (g1307) & (!g1309) & (!g1311)) + ((g1292) & (g1293) & (g1295) & (g1307) & (g1309) & (g1311)));
	assign g1313 = (((!g9) & (!g30) & (!g131) & (!sk[43]) & (g282)) + ((!g9) & (!g30) & (!g131) & (sk[43]) & (g282)) + ((!g9) & (!g30) & (g131) & (!sk[43]) & (g282)) + ((!g9) & (g30) & (!g131) & (!sk[43]) & (g282)) + ((!g9) & (g30) & (!g131) & (sk[43]) & (g282)) + ((!g9) & (g30) & (g131) & (!sk[43]) & (g282)) + ((g9) & (!g30) & (!g131) & (!sk[43]) & (!g282)) + ((g9) & (!g30) & (!g131) & (!sk[43]) & (g282)) + ((g9) & (!g30) & (!g131) & (sk[43]) & (g282)) + ((g9) & (!g30) & (g131) & (!sk[43]) & (!g282)) + ((g9) & (!g30) & (g131) & (!sk[43]) & (g282)) + ((g9) & (g30) & (!g131) & (!sk[43]) & (!g282)) + ((g9) & (g30) & (!g131) & (!sk[43]) & (g282)) + ((g9) & (g30) & (g131) & (!sk[43]) & (!g282)) + ((g9) & (g30) & (g131) & (!sk[43]) & (g282)));
	assign g1314 = (((!g62) & (!g32) & (!sk[44]) & (!g185) & (g147)) + ((!g62) & (!g32) & (!sk[44]) & (g185) & (g147)) + ((!g62) & (!g32) & (sk[44]) & (!g185) & (!g147)) + ((!g62) & (g32) & (!sk[44]) & (!g185) & (g147)) + ((!g62) & (g32) & (!sk[44]) & (g185) & (g147)) + ((!g62) & (g32) & (sk[44]) & (!g185) & (!g147)) + ((g62) & (!g32) & (!sk[44]) & (!g185) & (!g147)) + ((g62) & (!g32) & (!sk[44]) & (!g185) & (g147)) + ((g62) & (!g32) & (!sk[44]) & (g185) & (!g147)) + ((g62) & (!g32) & (!sk[44]) & (g185) & (g147)) + ((g62) & (!g32) & (sk[44]) & (!g185) & (!g147)) + ((g62) & (g32) & (!sk[44]) & (!g185) & (!g147)) + ((g62) & (g32) & (!sk[44]) & (!g185) & (g147)) + ((g62) & (g32) & (!sk[44]) & (g185) & (!g147)) + ((g62) & (g32) & (!sk[44]) & (g185) & (g147)));
	assign g1315 = (((!g92) & (!g967) & (!sk[45]) & (!g1274) & (g1314)) + ((!g92) & (!g967) & (!sk[45]) & (g1274) & (g1314)) + ((!g92) & (g967) & (!sk[45]) & (!g1274) & (g1314)) + ((!g92) & (g967) & (!sk[45]) & (g1274) & (g1314)) + ((g92) & (!g967) & (!sk[45]) & (!g1274) & (!g1314)) + ((g92) & (!g967) & (!sk[45]) & (!g1274) & (g1314)) + ((g92) & (!g967) & (!sk[45]) & (g1274) & (!g1314)) + ((g92) & (!g967) & (!sk[45]) & (g1274) & (g1314)) + ((g92) & (!g967) & (sk[45]) & (g1274) & (g1314)) + ((g92) & (g967) & (!sk[45]) & (!g1274) & (!g1314)) + ((g92) & (g967) & (!sk[45]) & (!g1274) & (g1314)) + ((g92) & (g967) & (!sk[45]) & (g1274) & (!g1314)) + ((g92) & (g967) & (!sk[45]) & (g1274) & (g1314)));
	assign g1316 = (((!g879) & (!g29) & (!sk[46]) & (!g254) & (g1315)) + ((!g879) & (!g29) & (!sk[46]) & (g254) & (g1315)) + ((!g879) & (g29) & (!sk[46]) & (!g254) & (g1315)) + ((!g879) & (g29) & (!sk[46]) & (g254) & (g1315)) + ((g879) & (!g29) & (!sk[46]) & (!g254) & (!g1315)) + ((g879) & (!g29) & (!sk[46]) & (!g254) & (g1315)) + ((g879) & (!g29) & (!sk[46]) & (g254) & (!g1315)) + ((g879) & (!g29) & (!sk[46]) & (g254) & (g1315)) + ((g879) & (!g29) & (sk[46]) & (!g254) & (g1315)) + ((g879) & (g29) & (!sk[46]) & (!g254) & (!g1315)) + ((g879) & (g29) & (!sk[46]) & (!g254) & (g1315)) + ((g879) & (g29) & (!sk[46]) & (g254) & (!g1315)) + ((g879) & (g29) & (!sk[46]) & (g254) & (g1315)));
	assign g1317 = (((!g123) & (!g1313) & (!g709) & (g1019) & (!sk[47]) & (!g1316)) + ((!g123) & (!g1313) & (!g709) & (g1019) & (!sk[47]) & (g1316)) + ((!g123) & (!g1313) & (g709) & (!g1019) & (!sk[47]) & (!g1316)) + ((!g123) & (!g1313) & (g709) & (!g1019) & (!sk[47]) & (g1316)) + ((!g123) & (!g1313) & (g709) & (g1019) & (!sk[47]) & (!g1316)) + ((!g123) & (!g1313) & (g709) & (g1019) & (!sk[47]) & (g1316)) + ((!g123) & (g1313) & (!g709) & (!g1019) & (!sk[47]) & (!g1316)) + ((!g123) & (g1313) & (!g709) & (!g1019) & (!sk[47]) & (g1316)) + ((!g123) & (g1313) & (!g709) & (g1019) & (!sk[47]) & (!g1316)) + ((!g123) & (g1313) & (!g709) & (g1019) & (!sk[47]) & (g1316)) + ((!g123) & (g1313) & (g709) & (!g1019) & (!sk[47]) & (!g1316)) + ((!g123) & (g1313) & (g709) & (!g1019) & (!sk[47]) & (g1316)) + ((!g123) & (g1313) & (g709) & (g1019) & (!sk[47]) & (!g1316)) + ((!g123) & (g1313) & (g709) & (g1019) & (!sk[47]) & (g1316)) + ((g123) & (!g1313) & (!g709) & (g1019) & (!sk[47]) & (!g1316)) + ((g123) & (!g1313) & (!g709) & (g1019) & (!sk[47]) & (g1316)) + ((g123) & (!g1313) & (g709) & (!g1019) & (!sk[47]) & (!g1316)) + ((g123) & (!g1313) & (g709) & (!g1019) & (!sk[47]) & (g1316)) + ((g123) & (!g1313) & (g709) & (g1019) & (!sk[47]) & (!g1316)) + ((g123) & (!g1313) & (g709) & (g1019) & (!sk[47]) & (g1316)) + ((g123) & (g1313) & (!g709) & (!g1019) & (!sk[47]) & (!g1316)) + ((g123) & (g1313) & (!g709) & (!g1019) & (!sk[47]) & (g1316)) + ((g123) & (g1313) & (!g709) & (g1019) & (!sk[47]) & (!g1316)) + ((g123) & (g1313) & (!g709) & (g1019) & (!sk[47]) & (g1316)) + ((g123) & (g1313) & (g709) & (!g1019) & (!sk[47]) & (!g1316)) + ((g123) & (g1313) & (g709) & (!g1019) & (!sk[47]) & (g1316)) + ((g123) & (g1313) & (g709) & (g1019) & (!sk[47]) & (!g1316)) + ((g123) & (g1313) & (g709) & (g1019) & (!sk[47]) & (g1316)) + ((g123) & (g1313) & (g709) & (g1019) & (sk[47]) & (g1316)));
	assign g1318 = (((!g1286) & (!g1287) & (!g1296) & (!g1305) & (!g1312) & (g1317)) + ((!g1286) & (!g1287) & (!g1296) & (!g1305) & (g1312) & (!g1317)) + ((!g1286) & (!g1287) & (!g1296) & (g1305) & (!g1312) & (!g1317)) + ((!g1286) & (!g1287) & (!g1296) & (g1305) & (g1312) & (g1317)) + ((!g1286) & (!g1287) & (g1296) & (!g1305) & (!g1312) & (!g1317)) + ((!g1286) & (!g1287) & (g1296) & (!g1305) & (g1312) & (g1317)) + ((!g1286) & (!g1287) & (g1296) & (g1305) & (!g1312) & (g1317)) + ((!g1286) & (!g1287) & (g1296) & (g1305) & (g1312) & (!g1317)) + ((!g1286) & (g1287) & (!g1296) & (!g1305) & (!g1312) & (g1317)) + ((!g1286) & (g1287) & (!g1296) & (!g1305) & (g1312) & (!g1317)) + ((!g1286) & (g1287) & (!g1296) & (g1305) & (!g1312) & (!g1317)) + ((!g1286) & (g1287) & (!g1296) & (g1305) & (g1312) & (g1317)) + ((!g1286) & (g1287) & (g1296) & (!g1305) & (!g1312) & (g1317)) + ((!g1286) & (g1287) & (g1296) & (!g1305) & (g1312) & (!g1317)) + ((!g1286) & (g1287) & (g1296) & (g1305) & (!g1312) & (!g1317)) + ((!g1286) & (g1287) & (g1296) & (g1305) & (g1312) & (g1317)) + ((g1286) & (!g1287) & (!g1296) & (!g1305) & (!g1312) & (!g1317)) + ((g1286) & (!g1287) & (!g1296) & (!g1305) & (g1312) & (g1317)) + ((g1286) & (!g1287) & (!g1296) & (g1305) & (!g1312) & (g1317)) + ((g1286) & (!g1287) & (!g1296) & (g1305) & (g1312) & (!g1317)) + ((g1286) & (!g1287) & (g1296) & (!g1305) & (!g1312) & (!g1317)) + ((g1286) & (!g1287) & (g1296) & (!g1305) & (g1312) & (g1317)) + ((g1286) & (!g1287) & (g1296) & (g1305) & (!g1312) & (g1317)) + ((g1286) & (!g1287) & (g1296) & (g1305) & (g1312) & (!g1317)) + ((g1286) & (g1287) & (!g1296) & (!g1305) & (!g1312) & (g1317)) + ((g1286) & (g1287) & (!g1296) & (!g1305) & (g1312) & (!g1317)) + ((g1286) & (g1287) & (!g1296) & (g1305) & (!g1312) & (!g1317)) + ((g1286) & (g1287) & (!g1296) & (g1305) & (g1312) & (g1317)) + ((g1286) & (g1287) & (g1296) & (!g1305) & (!g1312) & (!g1317)) + ((g1286) & (g1287) & (g1296) & (!g1305) & (g1312) & (g1317)) + ((g1286) & (g1287) & (g1296) & (g1305) & (!g1312) & (g1317)) + ((g1286) & (g1287) & (g1296) & (g1305) & (g1312) & (!g1317)));
	assign sinx10x = (((!g1068) & (!g1281) & (!g1283) & (!g1302) & (!g1304) & (!g1318)) + ((!g1068) & (!g1281) & (!g1283) & (!g1302) & (g1304) & (g1318)) + ((!g1068) & (!g1281) & (!g1283) & (g1302) & (!g1304) & (!g1318)) + ((!g1068) & (!g1281) & (!g1283) & (g1302) & (g1304) & (g1318)) + ((!g1068) & (!g1281) & (g1283) & (!g1302) & (!g1304) & (g1318)) + ((!g1068) & (!g1281) & (g1283) & (!g1302) & (g1304) & (!g1318)) + ((!g1068) & (!g1281) & (g1283) & (g1302) & (!g1304) & (!g1318)) + ((!g1068) & (!g1281) & (g1283) & (g1302) & (g1304) & (g1318)) + ((!g1068) & (g1281) & (!g1283) & (!g1302) & (!g1304) & (!g1318)) + ((!g1068) & (g1281) & (!g1283) & (!g1302) & (g1304) & (g1318)) + ((!g1068) & (g1281) & (!g1283) & (g1302) & (!g1304) & (!g1318)) + ((!g1068) & (g1281) & (!g1283) & (g1302) & (g1304) & (g1318)) + ((!g1068) & (g1281) & (g1283) & (!g1302) & (!g1304) & (g1318)) + ((!g1068) & (g1281) & (g1283) & (!g1302) & (g1304) & (!g1318)) + ((!g1068) & (g1281) & (g1283) & (g1302) & (!g1304) & (!g1318)) + ((!g1068) & (g1281) & (g1283) & (g1302) & (g1304) & (g1318)) + ((g1068) & (!g1281) & (!g1283) & (!g1302) & (!g1304) & (g1318)) + ((g1068) & (!g1281) & (!g1283) & (!g1302) & (g1304) & (!g1318)) + ((g1068) & (!g1281) & (!g1283) & (g1302) & (!g1304) & (g1318)) + ((g1068) & (!g1281) & (!g1283) & (g1302) & (g1304) & (!g1318)) + ((g1068) & (!g1281) & (g1283) & (!g1302) & (!g1304) & (!g1318)) + ((g1068) & (!g1281) & (g1283) & (!g1302) & (g1304) & (g1318)) + ((g1068) & (!g1281) & (g1283) & (g1302) & (!g1304) & (g1318)) + ((g1068) & (!g1281) & (g1283) & (g1302) & (g1304) & (!g1318)) + ((g1068) & (g1281) & (!g1283) & (!g1302) & (!g1304) & (g1318)) + ((g1068) & (g1281) & (!g1283) & (!g1302) & (g1304) & (!g1318)) + ((g1068) & (g1281) & (!g1283) & (g1302) & (!g1304) & (!g1318)) + ((g1068) & (g1281) & (!g1283) & (g1302) & (g1304) & (g1318)) + ((g1068) & (g1281) & (g1283) & (!g1302) & (!g1304) & (g1318)) + ((g1068) & (g1281) & (g1283) & (!g1302) & (g1304) & (!g1318)) + ((g1068) & (g1281) & (g1283) & (g1302) & (!g1304) & (g1318)) + ((g1068) & (g1281) & (g1283) & (g1302) & (g1304) & (!g1318)));
	assign g1320 = (((g1282) & (!g1258) & (g1279) & (!g1284) & (!g1297) & (g1301)) + ((g1282) & (!g1258) & (g1279) & (!g1284) & (g1297) & (!g1301)) + ((g1282) & (!g1258) & (g1279) & (g1284) & (!g1297) & (!g1301)) + ((g1282) & (!g1258) & (g1279) & (g1284) & (g1297) & (g1301)) + ((g1282) & (g1258) & (!g1279) & (!g1284) & (!g1297) & (g1301)) + ((g1282) & (g1258) & (!g1279) & (!g1284) & (g1297) & (!g1301)) + ((g1282) & (g1258) & (!g1279) & (g1284) & (!g1297) & (!g1301)) + ((g1282) & (g1258) & (!g1279) & (g1284) & (g1297) & (g1301)));
	assign g1321 = (((!g1320) & (!sk[51]) & (g1304) & (!g1318)) + ((!g1320) & (!sk[51]) & (g1304) & (g1318)) + ((g1320) & (!sk[51]) & (g1304) & (!g1318)) + ((g1320) & (!sk[51]) & (g1304) & (g1318)) + ((g1320) & (sk[51]) & (!g1304) & (!g1318)) + ((g1320) & (sk[51]) & (g1304) & (g1318)));
	assign g1322 = (((!g1286) & (!g1287) & (!sk[52]) & (!g1296) & (g1305) & (!g1312)) + ((!g1286) & (!g1287) & (!sk[52]) & (!g1296) & (g1305) & (g1312)) + ((!g1286) & (!g1287) & (!sk[52]) & (g1296) & (!g1305) & (!g1312)) + ((!g1286) & (!g1287) & (!sk[52]) & (g1296) & (!g1305) & (g1312)) + ((!g1286) & (!g1287) & (!sk[52]) & (g1296) & (g1305) & (!g1312)) + ((!g1286) & (!g1287) & (!sk[52]) & (g1296) & (g1305) & (g1312)) + ((!g1286) & (!g1287) & (sk[52]) & (!g1296) & (!g1305) & (!g1312)) + ((!g1286) & (!g1287) & (sk[52]) & (!g1296) & (g1305) & (g1312)) + ((!g1286) & (!g1287) & (sk[52]) & (g1296) & (!g1305) & (g1312)) + ((!g1286) & (!g1287) & (sk[52]) & (g1296) & (g1305) & (!g1312)) + ((!g1286) & (g1287) & (!sk[52]) & (!g1296) & (!g1305) & (!g1312)) + ((!g1286) & (g1287) & (!sk[52]) & (!g1296) & (!g1305) & (g1312)) + ((!g1286) & (g1287) & (!sk[52]) & (!g1296) & (g1305) & (!g1312)) + ((!g1286) & (g1287) & (!sk[52]) & (!g1296) & (g1305) & (g1312)) + ((!g1286) & (g1287) & (!sk[52]) & (g1296) & (!g1305) & (!g1312)) + ((!g1286) & (g1287) & (!sk[52]) & (g1296) & (!g1305) & (g1312)) + ((!g1286) & (g1287) & (!sk[52]) & (g1296) & (g1305) & (!g1312)) + ((!g1286) & (g1287) & (!sk[52]) & (g1296) & (g1305) & (g1312)) + ((!g1286) & (g1287) & (sk[52]) & (!g1296) & (!g1305) & (!g1312)) + ((!g1286) & (g1287) & (sk[52]) & (!g1296) & (g1305) & (g1312)) + ((!g1286) & (g1287) & (sk[52]) & (g1296) & (!g1305) & (!g1312)) + ((!g1286) & (g1287) & (sk[52]) & (g1296) & (g1305) & (g1312)) + ((g1286) & (!g1287) & (!sk[52]) & (!g1296) & (g1305) & (!g1312)) + ((g1286) & (!g1287) & (!sk[52]) & (!g1296) & (g1305) & (g1312)) + ((g1286) & (!g1287) & (!sk[52]) & (g1296) & (!g1305) & (!g1312)) + ((g1286) & (!g1287) & (!sk[52]) & (g1296) & (!g1305) & (g1312)) + ((g1286) & (!g1287) & (!sk[52]) & (g1296) & (g1305) & (!g1312)) + ((g1286) & (!g1287) & (!sk[52]) & (g1296) & (g1305) & (g1312)) + ((g1286) & (!g1287) & (sk[52]) & (!g1296) & (!g1305) & (g1312)) + ((g1286) & (!g1287) & (sk[52]) & (!g1296) & (g1305) & (!g1312)) + ((g1286) & (!g1287) & (sk[52]) & (g1296) & (!g1305) & (g1312)) + ((g1286) & (!g1287) & (sk[52]) & (g1296) & (g1305) & (!g1312)) + ((g1286) & (g1287) & (!sk[52]) & (!g1296) & (!g1305) & (!g1312)) + ((g1286) & (g1287) & (!sk[52]) & (!g1296) & (!g1305) & (g1312)) + ((g1286) & (g1287) & (!sk[52]) & (!g1296) & (g1305) & (!g1312)) + ((g1286) & (g1287) & (!sk[52]) & (!g1296) & (g1305) & (g1312)) + ((g1286) & (g1287) & (!sk[52]) & (g1296) & (!g1305) & (!g1312)) + ((g1286) & (g1287) & (!sk[52]) & (g1296) & (!g1305) & (g1312)) + ((g1286) & (g1287) & (!sk[52]) & (g1296) & (g1305) & (!g1312)) + ((g1286) & (g1287) & (!sk[52]) & (g1296) & (g1305) & (g1312)) + ((g1286) & (g1287) & (sk[52]) & (!g1296) & (!g1305) & (!g1312)) + ((g1286) & (g1287) & (sk[52]) & (!g1296) & (g1305) & (g1312)) + ((g1286) & (g1287) & (sk[52]) & (g1296) & (!g1305) & (g1312)) + ((g1286) & (g1287) & (sk[52]) & (g1296) & (g1305) & (!g1312)));
	assign g1323 = (((!g1284) & (!g1285) & (!g1297) & (!g1301) & (!g1322) & (g1317)) + ((!g1284) & (!g1285) & (!g1297) & (g1301) & (!g1322) & (!g1317)) + ((!g1284) & (!g1285) & (!g1297) & (g1301) & (!g1322) & (g1317)) + ((!g1284) & (!g1285) & (!g1297) & (g1301) & (g1322) & (g1317)) + ((!g1284) & (!g1285) & (g1297) & (!g1301) & (!g1322) & (!g1317)) + ((!g1284) & (!g1285) & (g1297) & (!g1301) & (!g1322) & (g1317)) + ((!g1284) & (!g1285) & (g1297) & (!g1301) & (g1322) & (g1317)) + ((!g1284) & (!g1285) & (g1297) & (g1301) & (!g1322) & (!g1317)) + ((!g1284) & (!g1285) & (g1297) & (g1301) & (!g1322) & (g1317)) + ((!g1284) & (!g1285) & (g1297) & (g1301) & (g1322) & (g1317)) + ((!g1284) & (g1285) & (!g1297) & (!g1301) & (!g1322) & (g1317)) + ((!g1284) & (g1285) & (!g1297) & (g1301) & (!g1322) & (g1317)) + ((!g1284) & (g1285) & (g1297) & (!g1301) & (!g1322) & (g1317)) + ((!g1284) & (g1285) & (g1297) & (g1301) & (!g1322) & (!g1317)) + ((!g1284) & (g1285) & (g1297) & (g1301) & (!g1322) & (g1317)) + ((!g1284) & (g1285) & (g1297) & (g1301) & (g1322) & (g1317)) + ((g1284) & (!g1285) & (!g1297) & (!g1301) & (!g1322) & (g1317)) + ((g1284) & (!g1285) & (!g1297) & (g1301) & (!g1322) & (g1317)) + ((g1284) & (!g1285) & (g1297) & (!g1301) & (!g1322) & (g1317)) + ((g1284) & (!g1285) & (g1297) & (g1301) & (!g1322) & (!g1317)) + ((g1284) & (!g1285) & (g1297) & (g1301) & (!g1322) & (g1317)) + ((g1284) & (!g1285) & (g1297) & (g1301) & (g1322) & (g1317)) + ((g1284) & (g1285) & (!g1297) & (!g1301) & (!g1322) & (g1317)) + ((g1284) & (g1285) & (!g1297) & (g1301) & (!g1322) & (g1317)) + ((g1284) & (g1285) & (g1297) & (!g1301) & (!g1322) & (g1317)) + ((g1284) & (g1285) & (g1297) & (g1301) & (!g1322) & (!g1317)) + ((g1284) & (g1285) & (g1297) & (g1301) & (!g1322) & (g1317)) + ((g1284) & (g1285) & (g1297) & (g1301) & (g1322) & (g1317)));
	assign g1324 = (((!g252) & (!g869) & (!sk[54]) & (!g870) & (g1290) & (!g1291)) + ((!g252) & (!g869) & (!sk[54]) & (!g870) & (g1290) & (g1291)) + ((!g252) & (!g869) & (!sk[54]) & (g870) & (!g1290) & (!g1291)) + ((!g252) & (!g869) & (!sk[54]) & (g870) & (!g1290) & (g1291)) + ((!g252) & (!g869) & (!sk[54]) & (g870) & (g1290) & (!g1291)) + ((!g252) & (!g869) & (!sk[54]) & (g870) & (g1290) & (g1291)) + ((!g252) & (!g869) & (sk[54]) & (!g870) & (!g1290) & (g1291)) + ((!g252) & (!g869) & (sk[54]) & (g870) & (!g1290) & (g1291)) + ((!g252) & (g869) & (!sk[54]) & (!g870) & (!g1290) & (!g1291)) + ((!g252) & (g869) & (!sk[54]) & (!g870) & (!g1290) & (g1291)) + ((!g252) & (g869) & (!sk[54]) & (!g870) & (g1290) & (!g1291)) + ((!g252) & (g869) & (!sk[54]) & (!g870) & (g1290) & (g1291)) + ((!g252) & (g869) & (!sk[54]) & (g870) & (!g1290) & (!g1291)) + ((!g252) & (g869) & (!sk[54]) & (g870) & (!g1290) & (g1291)) + ((!g252) & (g869) & (!sk[54]) & (g870) & (g1290) & (!g1291)) + ((!g252) & (g869) & (!sk[54]) & (g870) & (g1290) & (g1291)) + ((!g252) & (g869) & (sk[54]) & (!g870) & (!g1290) & (g1291)) + ((!g252) & (g869) & (sk[54]) & (g870) & (!g1290) & (g1291)) + ((g252) & (!g869) & (!sk[54]) & (!g870) & (g1290) & (!g1291)) + ((g252) & (!g869) & (!sk[54]) & (!g870) & (g1290) & (g1291)) + ((g252) & (!g869) & (!sk[54]) & (g870) & (!g1290) & (!g1291)) + ((g252) & (!g869) & (!sk[54]) & (g870) & (!g1290) & (g1291)) + ((g252) & (!g869) & (!sk[54]) & (g870) & (g1290) & (!g1291)) + ((g252) & (!g869) & (!sk[54]) & (g870) & (g1290) & (g1291)) + ((g252) & (!g869) & (sk[54]) & (g870) & (!g1290) & (!g1291)) + ((g252) & (!g869) & (sk[54]) & (g870) & (g1290) & (!g1291)) + ((g252) & (!g869) & (sk[54]) & (g870) & (g1290) & (g1291)) + ((g252) & (g869) & (!sk[54]) & (!g870) & (!g1290) & (!g1291)) + ((g252) & (g869) & (!sk[54]) & (!g870) & (!g1290) & (g1291)) + ((g252) & (g869) & (!sk[54]) & (!g870) & (g1290) & (!g1291)) + ((g252) & (g869) & (!sk[54]) & (!g870) & (g1290) & (g1291)) + ((g252) & (g869) & (!sk[54]) & (g870) & (!g1290) & (!g1291)) + ((g252) & (g869) & (!sk[54]) & (g870) & (!g1290) & (g1291)) + ((g252) & (g869) & (!sk[54]) & (g870) & (g1290) & (!g1291)) + ((g252) & (g869) & (!sk[54]) & (g870) & (g1290) & (g1291)) + ((g252) & (g869) & (sk[54]) & (!g870) & (!g1290) & (!g1291)) + ((g252) & (g869) & (sk[54]) & (!g870) & (g1290) & (!g1291)) + ((g252) & (g869) & (sk[54]) & (!g870) & (g1290) & (g1291)) + ((g252) & (g869) & (sk[54]) & (g870) & (!g1290) & (!g1291)) + ((g252) & (g869) & (sk[54]) & (g870) & (!g1290) & (g1291)) + ((g252) & (g869) & (sk[54]) & (g870) & (g1290) & (!g1291)) + ((g252) & (g869) & (sk[54]) & (g870) & (g1290) & (g1291)));
	assign g1325 = (((!g762) & (!sk[55]) & (!g765) & (!g1040) & (g1079)) + ((!g762) & (!sk[55]) & (!g765) & (g1040) & (g1079)) + ((!g762) & (!sk[55]) & (g765) & (!g1040) & (g1079)) + ((!g762) & (!sk[55]) & (g765) & (g1040) & (g1079)) + ((!g762) & (sk[55]) & (g765) & (!g1040) & (!g1079)) + ((!g762) & (sk[55]) & (g765) & (!g1040) & (g1079)) + ((g762) & (!sk[55]) & (!g765) & (!g1040) & (!g1079)) + ((g762) & (!sk[55]) & (!g765) & (!g1040) & (g1079)) + ((g762) & (!sk[55]) & (!g765) & (g1040) & (!g1079)) + ((g762) & (!sk[55]) & (!g765) & (g1040) & (g1079)) + ((g762) & (!sk[55]) & (g765) & (!g1040) & (!g1079)) + ((g762) & (!sk[55]) & (g765) & (!g1040) & (g1079)) + ((g762) & (!sk[55]) & (g765) & (g1040) & (!g1079)) + ((g762) & (!sk[55]) & (g765) & (g1040) & (g1079)) + ((g762) & (sk[55]) & (!g765) & (!g1040) & (!g1079)) + ((g762) & (sk[55]) & (!g765) & (g1040) & (!g1079)) + ((g762) & (sk[55]) & (g765) & (!g1040) & (!g1079)) + ((g762) & (sk[55]) & (g765) & (!g1040) & (g1079)) + ((g762) & (sk[55]) & (g765) & (g1040) & (!g1079)));
	assign g1326 = (((!g202) & (!g759) & (!g1040) & (!g1079) & (!g1080) & (g1325)) + ((!g202) & (!g759) & (!g1040) & (!g1079) & (g1080) & (g1325)) + ((!g202) & (!g759) & (!g1040) & (g1079) & (!g1080) & (g1325)) + ((!g202) & (!g759) & (!g1040) & (g1079) & (g1080) & (g1325)) + ((!g202) & (!g759) & (g1040) & (!g1079) & (!g1080) & (g1325)) + ((!g202) & (!g759) & (g1040) & (!g1079) & (g1080) & (g1325)) + ((!g202) & (!g759) & (g1040) & (g1079) & (!g1080) & (g1325)) + ((!g202) & (!g759) & (g1040) & (g1079) & (g1080) & (g1325)) + ((!g202) & (g759) & (!g1040) & (!g1079) & (!g1080) & (g1325)) + ((!g202) & (g759) & (!g1040) & (!g1079) & (g1080) & (g1325)) + ((!g202) & (g759) & (!g1040) & (g1079) & (!g1080) & (g1325)) + ((!g202) & (g759) & (!g1040) & (g1079) & (g1080) & (!g1325)) + ((!g202) & (g759) & (!g1040) & (g1079) & (g1080) & (g1325)) + ((!g202) & (g759) & (g1040) & (!g1079) & (!g1080) & (!g1325)) + ((!g202) & (g759) & (g1040) & (!g1079) & (!g1080) & (g1325)) + ((!g202) & (g759) & (g1040) & (!g1079) & (g1080) & (g1325)) + ((!g202) & (g759) & (g1040) & (g1079) & (!g1080) & (g1325)) + ((!g202) & (g759) & (g1040) & (g1079) & (g1080) & (g1325)) + ((g202) & (!g759) & (!g1040) & (!g1079) & (!g1080) & (!g1325)) + ((g202) & (!g759) & (!g1040) & (!g1079) & (g1080) & (!g1325)) + ((g202) & (!g759) & (!g1040) & (g1079) & (!g1080) & (!g1325)) + ((g202) & (!g759) & (!g1040) & (g1079) & (g1080) & (!g1325)) + ((g202) & (!g759) & (g1040) & (!g1079) & (!g1080) & (!g1325)) + ((g202) & (!g759) & (g1040) & (!g1079) & (g1080) & (!g1325)) + ((g202) & (!g759) & (g1040) & (g1079) & (!g1080) & (!g1325)) + ((g202) & (!g759) & (g1040) & (g1079) & (g1080) & (!g1325)) + ((g202) & (g759) & (!g1040) & (!g1079) & (!g1080) & (!g1325)) + ((g202) & (g759) & (!g1040) & (!g1079) & (g1080) & (!g1325)) + ((g202) & (g759) & (!g1040) & (g1079) & (!g1080) & (!g1325)) + ((g202) & (g759) & (g1040) & (!g1079) & (g1080) & (!g1325)) + ((g202) & (g759) & (g1040) & (g1079) & (!g1080) & (!g1325)) + ((g202) & (g759) & (g1040) & (g1079) & (g1080) & (!g1325)));
	assign g1327 = (((!g252) & (!g200) & (!sk[57]) & (!g869) & (g863)) + ((!g252) & (!g200) & (!sk[57]) & (g869) & (g863)) + ((!g252) & (g200) & (!sk[57]) & (!g869) & (g863)) + ((!g252) & (g200) & (!sk[57]) & (g869) & (g863)) + ((g252) & (!g200) & (!sk[57]) & (!g869) & (!g863)) + ((g252) & (!g200) & (!sk[57]) & (!g869) & (g863)) + ((g252) & (!g200) & (!sk[57]) & (g869) & (!g863)) + ((g252) & (!g200) & (!sk[57]) & (g869) & (g863)) + ((g252) & (!g200) & (sk[57]) & (!g869) & (g863)) + ((g252) & (!g200) & (sk[57]) & (g869) & (!g863)) + ((g252) & (!g200) & (sk[57]) & (g869) & (g863)) + ((g252) & (g200) & (!sk[57]) & (!g869) & (!g863)) + ((g252) & (g200) & (!sk[57]) & (!g869) & (g863)) + ((g252) & (g200) & (!sk[57]) & (g869) & (!g863)) + ((g252) & (g200) & (!sk[57]) & (g869) & (g863)) + ((g252) & (g200) & (sk[57]) & (g869) & (g863)));
	assign g1328 = (((!g847) & (!g845) & (!g848) & (!g962) & (!g971) & (!g994)) + ((!g847) & (!g845) & (!g848) & (!g962) & (!g971) & (g994)) + ((!g847) & (!g845) & (!g848) & (!g962) & (g971) & (!g994)) + ((!g847) & (!g845) & (!g848) & (!g962) & (g971) & (g994)) + ((!g847) & (!g845) & (!g848) & (g962) & (!g971) & (!g994)) + ((!g847) & (!g845) & (!g848) & (g962) & (!g971) & (g994)) + ((!g847) & (!g845) & (!g848) & (g962) & (g971) & (!g994)) + ((!g847) & (!g845) & (!g848) & (g962) & (g971) & (g994)) + ((!g847) & (!g845) & (g848) & (g962) & (!g971) & (!g994)) + ((!g847) & (!g845) & (g848) & (g962) & (!g971) & (g994)) + ((!g847) & (!g845) & (g848) & (g962) & (g971) & (!g994)) + ((!g847) & (!g845) & (g848) & (g962) & (g971) & (g994)) + ((!g847) & (g845) & (!g848) & (!g962) & (!g971) & (!g994)) + ((!g847) & (g845) & (!g848) & (!g962) & (!g971) & (g994)) + ((!g847) & (g845) & (!g848) & (g962) & (!g971) & (!g994)) + ((!g847) & (g845) & (!g848) & (g962) & (!g971) & (g994)) + ((!g847) & (g845) & (g848) & (g962) & (!g971) & (!g994)) + ((!g847) & (g845) & (g848) & (g962) & (!g971) & (g994)) + ((g847) & (!g845) & (!g848) & (!g962) & (!g971) & (!g994)) + ((g847) & (!g845) & (!g848) & (!g962) & (g971) & (!g994)) + ((g847) & (!g845) & (!g848) & (g962) & (!g971) & (!g994)) + ((g847) & (!g845) & (!g848) & (g962) & (g971) & (!g994)) + ((g847) & (!g845) & (g848) & (g962) & (!g971) & (!g994)) + ((g847) & (!g845) & (g848) & (g962) & (g971) & (!g994)) + ((g847) & (g845) & (!g848) & (!g962) & (!g971) & (!g994)) + ((g847) & (g845) & (!g848) & (g962) & (!g971) & (!g994)) + ((g847) & (g845) & (g848) & (g962) & (!g971) & (!g994)));
	assign g1329 = (((!g252) & (!g843) & (!g963) & (!g995) & (!g1327) & (g1328)) + ((!g252) & (!g843) & (!g963) & (!g995) & (g1327) & (!g1328)) + ((!g252) & (!g843) & (!g963) & (g995) & (!g1327) & (g1328)) + ((!g252) & (!g843) & (!g963) & (g995) & (g1327) & (!g1328)) + ((!g252) & (!g843) & (g963) & (!g995) & (!g1327) & (g1328)) + ((!g252) & (!g843) & (g963) & (!g995) & (g1327) & (!g1328)) + ((!g252) & (!g843) & (g963) & (g995) & (!g1327) & (g1328)) + ((!g252) & (!g843) & (g963) & (g995) & (g1327) & (!g1328)) + ((!g252) & (g843) & (!g963) & (!g995) & (!g1327) & (g1328)) + ((!g252) & (g843) & (!g963) & (!g995) & (g1327) & (!g1328)) + ((!g252) & (g843) & (!g963) & (g995) & (g1327) & (!g1328)) + ((!g252) & (g843) & (!g963) & (g995) & (g1327) & (g1328)) + ((!g252) & (g843) & (g963) & (!g995) & (!g1327) & (g1328)) + ((!g252) & (g843) & (g963) & (!g995) & (g1327) & (!g1328)) + ((!g252) & (g843) & (g963) & (g995) & (g1327) & (!g1328)) + ((!g252) & (g843) & (g963) & (g995) & (g1327) & (g1328)) + ((g252) & (!g843) & (!g963) & (!g995) & (!g1327) & (!g1328)) + ((g252) & (!g843) & (!g963) & (!g995) & (g1327) & (g1328)) + ((g252) & (!g843) & (!g963) & (g995) & (!g1327) & (!g1328)) + ((g252) & (!g843) & (!g963) & (g995) & (g1327) & (g1328)) + ((g252) & (!g843) & (g963) & (!g995) & (!g1327) & (g1328)) + ((g252) & (!g843) & (g963) & (!g995) & (g1327) & (!g1328)) + ((g252) & (!g843) & (g963) & (g995) & (!g1327) & (g1328)) + ((g252) & (!g843) & (g963) & (g995) & (g1327) & (!g1328)) + ((g252) & (g843) & (!g963) & (!g995) & (!g1327) & (!g1328)) + ((g252) & (g843) & (!g963) & (!g995) & (g1327) & (g1328)) + ((g252) & (g843) & (!g963) & (g995) & (!g1327) & (!g1328)) + ((g252) & (g843) & (!g963) & (g995) & (!g1327) & (g1328)) + ((g252) & (g843) & (g963) & (!g995) & (!g1327) & (g1328)) + ((g252) & (g843) & (g963) & (!g995) & (g1327) & (!g1328)) + ((g252) & (g843) & (g963) & (g995) & (g1327) & (!g1328)) + ((g252) & (g843) & (g963) & (g995) & (g1327) & (g1328)));
	assign g1330 = (((!sk[60]) & (!g1307) & (!g1308) & (!g1324) & (g1326) & (!g1329)) + ((!sk[60]) & (!g1307) & (!g1308) & (!g1324) & (g1326) & (g1329)) + ((!sk[60]) & (!g1307) & (!g1308) & (g1324) & (!g1326) & (!g1329)) + ((!sk[60]) & (!g1307) & (!g1308) & (g1324) & (!g1326) & (g1329)) + ((!sk[60]) & (!g1307) & (!g1308) & (g1324) & (g1326) & (!g1329)) + ((!sk[60]) & (!g1307) & (!g1308) & (g1324) & (g1326) & (g1329)) + ((!sk[60]) & (!g1307) & (g1308) & (!g1324) & (!g1326) & (!g1329)) + ((!sk[60]) & (!g1307) & (g1308) & (!g1324) & (!g1326) & (g1329)) + ((!sk[60]) & (!g1307) & (g1308) & (!g1324) & (g1326) & (!g1329)) + ((!sk[60]) & (!g1307) & (g1308) & (!g1324) & (g1326) & (g1329)) + ((!sk[60]) & (!g1307) & (g1308) & (g1324) & (!g1326) & (!g1329)) + ((!sk[60]) & (!g1307) & (g1308) & (g1324) & (!g1326) & (g1329)) + ((!sk[60]) & (!g1307) & (g1308) & (g1324) & (g1326) & (!g1329)) + ((!sk[60]) & (!g1307) & (g1308) & (g1324) & (g1326) & (g1329)) + ((!sk[60]) & (g1307) & (!g1308) & (!g1324) & (g1326) & (!g1329)) + ((!sk[60]) & (g1307) & (!g1308) & (!g1324) & (g1326) & (g1329)) + ((!sk[60]) & (g1307) & (!g1308) & (g1324) & (!g1326) & (!g1329)) + ((!sk[60]) & (g1307) & (!g1308) & (g1324) & (!g1326) & (g1329)) + ((!sk[60]) & (g1307) & (!g1308) & (g1324) & (g1326) & (!g1329)) + ((!sk[60]) & (g1307) & (!g1308) & (g1324) & (g1326) & (g1329)) + ((!sk[60]) & (g1307) & (g1308) & (!g1324) & (!g1326) & (!g1329)) + ((!sk[60]) & (g1307) & (g1308) & (!g1324) & (!g1326) & (g1329)) + ((!sk[60]) & (g1307) & (g1308) & (!g1324) & (g1326) & (!g1329)) + ((!sk[60]) & (g1307) & (g1308) & (!g1324) & (g1326) & (g1329)) + ((!sk[60]) & (g1307) & (g1308) & (g1324) & (!g1326) & (!g1329)) + ((!sk[60]) & (g1307) & (g1308) & (g1324) & (!g1326) & (g1329)) + ((!sk[60]) & (g1307) & (g1308) & (g1324) & (g1326) & (!g1329)) + ((!sk[60]) & (g1307) & (g1308) & (g1324) & (g1326) & (g1329)) + ((sk[60]) & (!g1307) & (!g1308) & (!g1324) & (!g1326) & (g1329)) + ((sk[60]) & (!g1307) & (!g1308) & (!g1324) & (g1326) & (!g1329)) + ((sk[60]) & (!g1307) & (!g1308) & (g1324) & (!g1326) & (g1329)) + ((sk[60]) & (!g1307) & (!g1308) & (g1324) & (g1326) & (!g1329)) + ((sk[60]) & (!g1307) & (g1308) & (!g1324) & (!g1326) & (!g1329)) + ((sk[60]) & (!g1307) & (g1308) & (!g1324) & (g1326) & (g1329)) + ((sk[60]) & (!g1307) & (g1308) & (g1324) & (!g1326) & (g1329)) + ((sk[60]) & (!g1307) & (g1308) & (g1324) & (g1326) & (!g1329)) + ((sk[60]) & (g1307) & (!g1308) & (!g1324) & (!g1326) & (!g1329)) + ((sk[60]) & (g1307) & (!g1308) & (!g1324) & (g1326) & (g1329)) + ((sk[60]) & (g1307) & (!g1308) & (g1324) & (!g1326) & (g1329)) + ((sk[60]) & (g1307) & (!g1308) & (g1324) & (g1326) & (!g1329)) + ((sk[60]) & (g1307) & (g1308) & (!g1324) & (!g1326) & (!g1329)) + ((sk[60]) & (g1307) & (g1308) & (!g1324) & (g1326) & (g1329)) + ((sk[60]) & (g1307) & (g1308) & (g1324) & (!g1326) & (!g1329)) + ((sk[60]) & (g1307) & (g1308) & (g1324) & (g1326) & (g1329)));
	assign g1331 = (((!g1292) & (!g1293) & (!g1295) & (!g1307) & (!g1309) & (!g1311)) + ((!g1292) & (!g1293) & (!g1295) & (!g1307) & (!g1309) & (g1311)) + ((!g1292) & (!g1293) & (!g1295) & (!g1307) & (g1309) & (g1311)) + ((!g1292) & (!g1293) & (!g1295) & (g1307) & (!g1309) & (g1311)) + ((!g1292) & (!g1293) & (!g1295) & (g1307) & (g1309) & (!g1311)) + ((!g1292) & (!g1293) & (!g1295) & (g1307) & (g1309) & (g1311)) + ((!g1292) & (!g1293) & (g1295) & (!g1307) & (!g1309) & (g1311)) + ((!g1292) & (!g1293) & (g1295) & (g1307) & (g1309) & (g1311)) + ((!g1292) & (g1293) & (!g1295) & (!g1307) & (!g1309) & (!g1311)) + ((!g1292) & (g1293) & (!g1295) & (!g1307) & (!g1309) & (g1311)) + ((!g1292) & (g1293) & (!g1295) & (!g1307) & (g1309) & (g1311)) + ((!g1292) & (g1293) & (!g1295) & (g1307) & (!g1309) & (g1311)) + ((!g1292) & (g1293) & (!g1295) & (g1307) & (g1309) & (!g1311)) + ((!g1292) & (g1293) & (!g1295) & (g1307) & (g1309) & (g1311)) + ((!g1292) & (g1293) & (g1295) & (!g1307) & (!g1309) & (!g1311)) + ((!g1292) & (g1293) & (g1295) & (!g1307) & (!g1309) & (g1311)) + ((!g1292) & (g1293) & (g1295) & (!g1307) & (g1309) & (g1311)) + ((!g1292) & (g1293) & (g1295) & (g1307) & (!g1309) & (g1311)) + ((!g1292) & (g1293) & (g1295) & (g1307) & (g1309) & (!g1311)) + ((!g1292) & (g1293) & (g1295) & (g1307) & (g1309) & (g1311)) + ((g1292) & (!g1293) & (!g1295) & (!g1307) & (!g1309) & (g1311)) + ((g1292) & (!g1293) & (!g1295) & (g1307) & (g1309) & (g1311)) + ((g1292) & (!g1293) & (g1295) & (!g1307) & (!g1309) & (g1311)) + ((g1292) & (!g1293) & (g1295) & (g1307) & (g1309) & (g1311)) + ((g1292) & (g1293) & (!g1295) & (!g1307) & (!g1309) & (!g1311)) + ((g1292) & (g1293) & (!g1295) & (!g1307) & (!g1309) & (g1311)) + ((g1292) & (g1293) & (!g1295) & (!g1307) & (g1309) & (g1311)) + ((g1292) & (g1293) & (!g1295) & (g1307) & (!g1309) & (g1311)) + ((g1292) & (g1293) & (!g1295) & (g1307) & (g1309) & (!g1311)) + ((g1292) & (g1293) & (!g1295) & (g1307) & (g1309) & (g1311)) + ((g1292) & (g1293) & (g1295) & (!g1307) & (!g1309) & (g1311)) + ((g1292) & (g1293) & (g1295) & (g1307) & (g1309) & (g1311)));
	assign g1332 = (((!g1330) & (sk[62]) & (g1331)) + ((g1330) & (!sk[62]) & (g1331)) + ((g1330) & (sk[62]) & (!g1331)));
	assign g1333 = (((!g1286) & (!g1287) & (!g1296) & (!g1305) & (!g1312) & (g1332)) + ((!g1286) & (!g1287) & (!g1296) & (!g1305) & (g1312) & (!g1332)) + ((!g1286) & (!g1287) & (!g1296) & (g1305) & (!g1312) & (!g1332)) + ((!g1286) & (!g1287) & (!g1296) & (g1305) & (g1312) & (!g1332)) + ((!g1286) & (!g1287) & (g1296) & (!g1305) & (!g1312) & (g1332)) + ((!g1286) & (!g1287) & (g1296) & (!g1305) & (g1312) & (g1332)) + ((!g1286) & (!g1287) & (g1296) & (g1305) & (!g1312) & (g1332)) + ((!g1286) & (!g1287) & (g1296) & (g1305) & (g1312) & (!g1332)) + ((!g1286) & (g1287) & (!g1296) & (!g1305) & (!g1312) & (g1332)) + ((!g1286) & (g1287) & (!g1296) & (!g1305) & (g1312) & (!g1332)) + ((!g1286) & (g1287) & (!g1296) & (g1305) & (!g1312) & (!g1332)) + ((!g1286) & (g1287) & (!g1296) & (g1305) & (g1312) & (!g1332)) + ((!g1286) & (g1287) & (g1296) & (!g1305) & (!g1312) & (g1332)) + ((!g1286) & (g1287) & (g1296) & (!g1305) & (g1312) & (!g1332)) + ((!g1286) & (g1287) & (g1296) & (g1305) & (!g1312) & (!g1332)) + ((!g1286) & (g1287) & (g1296) & (g1305) & (g1312) & (!g1332)) + ((g1286) & (!g1287) & (!g1296) & (!g1305) & (!g1312) & (g1332)) + ((g1286) & (!g1287) & (!g1296) & (!g1305) & (g1312) & (g1332)) + ((g1286) & (!g1287) & (!g1296) & (g1305) & (!g1312) & (g1332)) + ((g1286) & (!g1287) & (!g1296) & (g1305) & (g1312) & (!g1332)) + ((g1286) & (!g1287) & (g1296) & (!g1305) & (!g1312) & (g1332)) + ((g1286) & (!g1287) & (g1296) & (!g1305) & (g1312) & (g1332)) + ((g1286) & (!g1287) & (g1296) & (g1305) & (!g1312) & (g1332)) + ((g1286) & (!g1287) & (g1296) & (g1305) & (g1312) & (!g1332)) + ((g1286) & (g1287) & (!g1296) & (!g1305) & (!g1312) & (g1332)) + ((g1286) & (g1287) & (!g1296) & (!g1305) & (g1312) & (!g1332)) + ((g1286) & (g1287) & (!g1296) & (g1305) & (!g1312) & (!g1332)) + ((g1286) & (g1287) & (!g1296) & (g1305) & (g1312) & (!g1332)) + ((g1286) & (g1287) & (g1296) & (!g1305) & (!g1312) & (g1332)) + ((g1286) & (g1287) & (g1296) & (!g1305) & (g1312) & (g1332)) + ((g1286) & (g1287) & (g1296) & (g1305) & (!g1312) & (g1332)) + ((g1286) & (g1287) & (g1296) & (g1305) & (g1312) & (!g1332)));
	assign g1334 = (((!g275) & (!g208) & (!sk[64]) & (!g964) & (g349) & (!g157)) + ((!g275) & (!g208) & (!sk[64]) & (!g964) & (g349) & (g157)) + ((!g275) & (!g208) & (!sk[64]) & (g964) & (!g349) & (!g157)) + ((!g275) & (!g208) & (!sk[64]) & (g964) & (!g349) & (g157)) + ((!g275) & (!g208) & (!sk[64]) & (g964) & (g349) & (!g157)) + ((!g275) & (!g208) & (!sk[64]) & (g964) & (g349) & (g157)) + ((!g275) & (g208) & (!sk[64]) & (!g964) & (!g349) & (!g157)) + ((!g275) & (g208) & (!sk[64]) & (!g964) & (!g349) & (g157)) + ((!g275) & (g208) & (!sk[64]) & (!g964) & (g349) & (!g157)) + ((!g275) & (g208) & (!sk[64]) & (!g964) & (g349) & (g157)) + ((!g275) & (g208) & (!sk[64]) & (g964) & (!g349) & (!g157)) + ((!g275) & (g208) & (!sk[64]) & (g964) & (!g349) & (g157)) + ((!g275) & (g208) & (!sk[64]) & (g964) & (g349) & (!g157)) + ((!g275) & (g208) & (!sk[64]) & (g964) & (g349) & (g157)) + ((!g275) & (g208) & (sk[64]) & (g964) & (g349) & (g157)) + ((g275) & (!g208) & (!sk[64]) & (!g964) & (g349) & (!g157)) + ((g275) & (!g208) & (!sk[64]) & (!g964) & (g349) & (g157)) + ((g275) & (!g208) & (!sk[64]) & (g964) & (!g349) & (!g157)) + ((g275) & (!g208) & (!sk[64]) & (g964) & (!g349) & (g157)) + ((g275) & (!g208) & (!sk[64]) & (g964) & (g349) & (!g157)) + ((g275) & (!g208) & (!sk[64]) & (g964) & (g349) & (g157)) + ((g275) & (g208) & (!sk[64]) & (!g964) & (!g349) & (!g157)) + ((g275) & (g208) & (!sk[64]) & (!g964) & (!g349) & (g157)) + ((g275) & (g208) & (!sk[64]) & (!g964) & (g349) & (!g157)) + ((g275) & (g208) & (!sk[64]) & (!g964) & (g349) & (g157)) + ((g275) & (g208) & (!sk[64]) & (g964) & (!g349) & (!g157)) + ((g275) & (g208) & (!sk[64]) & (g964) & (!g349) & (g157)) + ((g275) & (g208) & (!sk[64]) & (g964) & (g349) & (!g157)) + ((g275) & (g208) & (!sk[64]) & (g964) & (g349) & (g157)));
	assign g1335 = (((!g259) & (!g286) & (!sk[65]) & (!g293) & (g1035) & (!g1334)) + ((!g259) & (!g286) & (!sk[65]) & (!g293) & (g1035) & (g1334)) + ((!g259) & (!g286) & (!sk[65]) & (g293) & (!g1035) & (!g1334)) + ((!g259) & (!g286) & (!sk[65]) & (g293) & (!g1035) & (g1334)) + ((!g259) & (!g286) & (!sk[65]) & (g293) & (g1035) & (!g1334)) + ((!g259) & (!g286) & (!sk[65]) & (g293) & (g1035) & (g1334)) + ((!g259) & (g286) & (!sk[65]) & (!g293) & (!g1035) & (!g1334)) + ((!g259) & (g286) & (!sk[65]) & (!g293) & (!g1035) & (g1334)) + ((!g259) & (g286) & (!sk[65]) & (!g293) & (g1035) & (!g1334)) + ((!g259) & (g286) & (!sk[65]) & (!g293) & (g1035) & (g1334)) + ((!g259) & (g286) & (!sk[65]) & (g293) & (!g1035) & (!g1334)) + ((!g259) & (g286) & (!sk[65]) & (g293) & (!g1035) & (g1334)) + ((!g259) & (g286) & (!sk[65]) & (g293) & (g1035) & (!g1334)) + ((!g259) & (g286) & (!sk[65]) & (g293) & (g1035) & (g1334)) + ((g259) & (!g286) & (!sk[65]) & (!g293) & (g1035) & (!g1334)) + ((g259) & (!g286) & (!sk[65]) & (!g293) & (g1035) & (g1334)) + ((g259) & (!g286) & (!sk[65]) & (g293) & (!g1035) & (!g1334)) + ((g259) & (!g286) & (!sk[65]) & (g293) & (!g1035) & (g1334)) + ((g259) & (!g286) & (!sk[65]) & (g293) & (g1035) & (!g1334)) + ((g259) & (!g286) & (!sk[65]) & (g293) & (g1035) & (g1334)) + ((g259) & (g286) & (!sk[65]) & (!g293) & (!g1035) & (!g1334)) + ((g259) & (g286) & (!sk[65]) & (!g293) & (!g1035) & (g1334)) + ((g259) & (g286) & (!sk[65]) & (!g293) & (g1035) & (!g1334)) + ((g259) & (g286) & (!sk[65]) & (!g293) & (g1035) & (g1334)) + ((g259) & (g286) & (!sk[65]) & (g293) & (!g1035) & (!g1334)) + ((g259) & (g286) & (!sk[65]) & (g293) & (!g1035) & (g1334)) + ((g259) & (g286) & (!sk[65]) & (g293) & (g1035) & (!g1334)) + ((g259) & (g286) & (!sk[65]) & (g293) & (g1035) & (g1334)) + ((g259) & (g286) & (sk[65]) & (g293) & (g1035) & (g1334)));
	assign g1336 = (((!sk[66]) & (g1333) & (g1335)) + ((sk[66]) & (!g1333) & (!g1335)) + ((sk[66]) & (g1333) & (g1335)));
	assign g1337 = (((!g1323) & (sk[67]) & (!g1336)) + ((g1323) & (!sk[67]) & (g1336)) + ((g1323) & (sk[67]) & (g1336)));
	assign g1338 = (((!g1281) & (!sk[68]) & (!g1283) & (!g1302) & (g1304) & (!g1318)) + ((!g1281) & (!sk[68]) & (!g1283) & (!g1302) & (g1304) & (g1318)) + ((!g1281) & (!sk[68]) & (!g1283) & (g1302) & (!g1304) & (!g1318)) + ((!g1281) & (!sk[68]) & (!g1283) & (g1302) & (!g1304) & (g1318)) + ((!g1281) & (!sk[68]) & (!g1283) & (g1302) & (g1304) & (!g1318)) + ((!g1281) & (!sk[68]) & (!g1283) & (g1302) & (g1304) & (g1318)) + ((!g1281) & (!sk[68]) & (g1283) & (!g1302) & (!g1304) & (!g1318)) + ((!g1281) & (!sk[68]) & (g1283) & (!g1302) & (!g1304) & (g1318)) + ((!g1281) & (!sk[68]) & (g1283) & (!g1302) & (g1304) & (!g1318)) + ((!g1281) & (!sk[68]) & (g1283) & (!g1302) & (g1304) & (g1318)) + ((!g1281) & (!sk[68]) & (g1283) & (g1302) & (!g1304) & (!g1318)) + ((!g1281) & (!sk[68]) & (g1283) & (g1302) & (!g1304) & (g1318)) + ((!g1281) & (!sk[68]) & (g1283) & (g1302) & (g1304) & (!g1318)) + ((!g1281) & (!sk[68]) & (g1283) & (g1302) & (g1304) & (g1318)) + ((g1281) & (!sk[68]) & (!g1283) & (!g1302) & (g1304) & (!g1318)) + ((g1281) & (!sk[68]) & (!g1283) & (!g1302) & (g1304) & (g1318)) + ((g1281) & (!sk[68]) & (!g1283) & (g1302) & (!g1304) & (!g1318)) + ((g1281) & (!sk[68]) & (!g1283) & (g1302) & (!g1304) & (g1318)) + ((g1281) & (!sk[68]) & (!g1283) & (g1302) & (g1304) & (!g1318)) + ((g1281) & (!sk[68]) & (!g1283) & (g1302) & (g1304) & (g1318)) + ((g1281) & (!sk[68]) & (g1283) & (!g1302) & (!g1304) & (!g1318)) + ((g1281) & (!sk[68]) & (g1283) & (!g1302) & (!g1304) & (g1318)) + ((g1281) & (!sk[68]) & (g1283) & (!g1302) & (g1304) & (!g1318)) + ((g1281) & (!sk[68]) & (g1283) & (!g1302) & (g1304) & (g1318)) + ((g1281) & (!sk[68]) & (g1283) & (g1302) & (!g1304) & (!g1318)) + ((g1281) & (!sk[68]) & (g1283) & (g1302) & (!g1304) & (g1318)) + ((g1281) & (!sk[68]) & (g1283) & (g1302) & (g1304) & (!g1318)) + ((g1281) & (!sk[68]) & (g1283) & (g1302) & (g1304) & (g1318)) + ((g1281) & (sk[68]) & (!g1283) & (g1302) & (!g1304) & (g1318)) + ((g1281) & (sk[68]) & (!g1283) & (g1302) & (g1304) & (!g1318)) + ((g1281) & (sk[68]) & (g1283) & (!g1302) & (!g1304) & (!g1318)) + ((g1281) & (sk[68]) & (g1283) & (!g1302) & (g1304) & (g1318)));
	assign g1339 = (((!sk[69]) & (!g1068) & (!g1321) & (!g1337) & (g1338)) + ((!sk[69]) & (!g1068) & (!g1321) & (g1337) & (g1338)) + ((!sk[69]) & (!g1068) & (g1321) & (!g1337) & (g1338)) + ((!sk[69]) & (!g1068) & (g1321) & (g1337) & (g1338)) + ((!sk[69]) & (g1068) & (!g1321) & (!g1337) & (!g1338)) + ((!sk[69]) & (g1068) & (!g1321) & (!g1337) & (g1338)) + ((!sk[69]) & (g1068) & (!g1321) & (g1337) & (!g1338)) + ((!sk[69]) & (g1068) & (!g1321) & (g1337) & (g1338)) + ((!sk[69]) & (g1068) & (g1321) & (!g1337) & (!g1338)) + ((!sk[69]) & (g1068) & (g1321) & (!g1337) & (g1338)) + ((!sk[69]) & (g1068) & (g1321) & (g1337) & (!g1338)) + ((!sk[69]) & (g1068) & (g1321) & (g1337) & (g1338)) + ((sk[69]) & (!g1068) & (!g1321) & (g1337) & (!g1338)) + ((sk[69]) & (!g1068) & (!g1321) & (g1337) & (g1338)) + ((sk[69]) & (!g1068) & (g1321) & (!g1337) & (!g1338)) + ((sk[69]) & (!g1068) & (g1321) & (!g1337) & (g1338)) + ((sk[69]) & (g1068) & (!g1321) & (!g1337) & (!g1338)) + ((sk[69]) & (g1068) & (!g1321) & (g1337) & (g1338)) + ((sk[69]) & (g1068) & (g1321) & (!g1337) & (g1338)) + ((sk[69]) & (g1068) & (g1321) & (g1337) & (!g1338)));
	assign g1340 = (((!g1307) & (!g1308) & (!g1324) & (!sk[70]) & (g1326) & (!g1329)) + ((!g1307) & (!g1308) & (!g1324) & (!sk[70]) & (g1326) & (g1329)) + ((!g1307) & (!g1308) & (!g1324) & (sk[70]) & (g1326) & (g1329)) + ((!g1307) & (!g1308) & (g1324) & (!sk[70]) & (!g1326) & (!g1329)) + ((!g1307) & (!g1308) & (g1324) & (!sk[70]) & (!g1326) & (g1329)) + ((!g1307) & (!g1308) & (g1324) & (!sk[70]) & (g1326) & (!g1329)) + ((!g1307) & (!g1308) & (g1324) & (!sk[70]) & (g1326) & (g1329)) + ((!g1307) & (!g1308) & (g1324) & (sk[70]) & (g1326) & (g1329)) + ((!g1307) & (g1308) & (!g1324) & (!sk[70]) & (!g1326) & (!g1329)) + ((!g1307) & (g1308) & (!g1324) & (!sk[70]) & (!g1326) & (g1329)) + ((!g1307) & (g1308) & (!g1324) & (!sk[70]) & (g1326) & (!g1329)) + ((!g1307) & (g1308) & (!g1324) & (!sk[70]) & (g1326) & (g1329)) + ((!g1307) & (g1308) & (!g1324) & (sk[70]) & (!g1326) & (g1329)) + ((!g1307) & (g1308) & (!g1324) & (sk[70]) & (g1326) & (!g1329)) + ((!g1307) & (g1308) & (!g1324) & (sk[70]) & (g1326) & (g1329)) + ((!g1307) & (g1308) & (g1324) & (!sk[70]) & (!g1326) & (!g1329)) + ((!g1307) & (g1308) & (g1324) & (!sk[70]) & (!g1326) & (g1329)) + ((!g1307) & (g1308) & (g1324) & (!sk[70]) & (g1326) & (!g1329)) + ((!g1307) & (g1308) & (g1324) & (!sk[70]) & (g1326) & (g1329)) + ((!g1307) & (g1308) & (g1324) & (sk[70]) & (g1326) & (g1329)) + ((g1307) & (!g1308) & (!g1324) & (!sk[70]) & (g1326) & (!g1329)) + ((g1307) & (!g1308) & (!g1324) & (!sk[70]) & (g1326) & (g1329)) + ((g1307) & (!g1308) & (!g1324) & (sk[70]) & (!g1326) & (g1329)) + ((g1307) & (!g1308) & (!g1324) & (sk[70]) & (g1326) & (!g1329)) + ((g1307) & (!g1308) & (!g1324) & (sk[70]) & (g1326) & (g1329)) + ((g1307) & (!g1308) & (g1324) & (!sk[70]) & (!g1326) & (!g1329)) + ((g1307) & (!g1308) & (g1324) & (!sk[70]) & (!g1326) & (g1329)) + ((g1307) & (!g1308) & (g1324) & (!sk[70]) & (g1326) & (!g1329)) + ((g1307) & (!g1308) & (g1324) & (!sk[70]) & (g1326) & (g1329)) + ((g1307) & (!g1308) & (g1324) & (sk[70]) & (g1326) & (g1329)) + ((g1307) & (g1308) & (!g1324) & (!sk[70]) & (!g1326) & (!g1329)) + ((g1307) & (g1308) & (!g1324) & (!sk[70]) & (!g1326) & (g1329)) + ((g1307) & (g1308) & (!g1324) & (!sk[70]) & (g1326) & (!g1329)) + ((g1307) & (g1308) & (!g1324) & (!sk[70]) & (g1326) & (g1329)) + ((g1307) & (g1308) & (!g1324) & (sk[70]) & (!g1326) & (g1329)) + ((g1307) & (g1308) & (!g1324) & (sk[70]) & (g1326) & (!g1329)) + ((g1307) & (g1308) & (!g1324) & (sk[70]) & (g1326) & (g1329)) + ((g1307) & (g1308) & (g1324) & (!sk[70]) & (!g1326) & (!g1329)) + ((g1307) & (g1308) & (g1324) & (!sk[70]) & (!g1326) & (g1329)) + ((g1307) & (g1308) & (g1324) & (!sk[70]) & (g1326) & (!g1329)) + ((g1307) & (g1308) & (g1324) & (!sk[70]) & (g1326) & (g1329)) + ((g1307) & (g1308) & (g1324) & (sk[70]) & (!g1326) & (g1329)) + ((g1307) & (g1308) & (g1324) & (sk[70]) & (g1326) & (!g1329)) + ((g1307) & (g1308) & (g1324) & (sk[70]) & (g1326) & (g1329)));
	assign g1341 = (((!g202) & (!g759) & (g765) & (!g1040) & (!g1079) & (!g1080)) + ((!g202) & (!g759) & (g765) & (!g1040) & (!g1079) & (g1080)) + ((!g202) & (!g759) & (g765) & (g1040) & (!g1079) & (!g1080)) + ((!g202) & (!g759) & (g765) & (g1040) & (!g1079) & (g1080)) + ((!g202) & (g759) & (!g765) & (!g1040) & (!g1079) & (!g1080)) + ((!g202) & (g759) & (!g765) & (!g1040) & (!g1079) & (g1080)) + ((!g202) & (g759) & (!g765) & (g1040) & (!g1079) & (g1080)) + ((!g202) & (g759) & (g765) & (!g1040) & (!g1079) & (!g1080)) + ((!g202) & (g759) & (g765) & (!g1040) & (!g1079) & (g1080)) + ((!g202) & (g759) & (g765) & (g1040) & (!g1079) & (!g1080)) + ((!g202) & (g759) & (g765) & (g1040) & (!g1079) & (g1080)) + ((g202) & (!g759) & (!g765) & (!g1040) & (!g1079) & (!g1080)) + ((g202) & (!g759) & (!g765) & (!g1040) & (!g1079) & (g1080)) + ((g202) & (!g759) & (!g765) & (!g1040) & (g1079) & (!g1080)) + ((g202) & (!g759) & (!g765) & (!g1040) & (g1079) & (g1080)) + ((g202) & (!g759) & (!g765) & (g1040) & (!g1079) & (!g1080)) + ((g202) & (!g759) & (!g765) & (g1040) & (!g1079) & (g1080)) + ((g202) & (!g759) & (!g765) & (g1040) & (g1079) & (!g1080)) + ((g202) & (!g759) & (!g765) & (g1040) & (g1079) & (g1080)) + ((g202) & (!g759) & (g765) & (!g1040) & (g1079) & (!g1080)) + ((g202) & (!g759) & (g765) & (!g1040) & (g1079) & (g1080)) + ((g202) & (!g759) & (g765) & (g1040) & (g1079) & (!g1080)) + ((g202) & (!g759) & (g765) & (g1040) & (g1079) & (g1080)) + ((g202) & (g759) & (!g765) & (!g1040) & (g1079) & (!g1080)) + ((g202) & (g759) & (!g765) & (!g1040) & (g1079) & (g1080)) + ((g202) & (g759) & (!g765) & (g1040) & (!g1079) & (!g1080)) + ((g202) & (g759) & (!g765) & (g1040) & (g1079) & (!g1080)) + ((g202) & (g759) & (!g765) & (g1040) & (g1079) & (g1080)) + ((g202) & (g759) & (g765) & (!g1040) & (g1079) & (!g1080)) + ((g202) & (g759) & (g765) & (!g1040) & (g1079) & (g1080)) + ((g202) & (g759) & (g765) & (g1040) & (g1079) & (!g1080)) + ((g202) & (g759) & (g765) & (g1040) & (g1079) & (g1080)));
	assign g1342 = (((!g847) & (!sk[72]) & (!g845) & (!g994) & (g1040)) + ((!g847) & (!sk[72]) & (!g845) & (g994) & (g1040)) + ((!g847) & (!sk[72]) & (g845) & (!g994) & (g1040)) + ((!g847) & (!sk[72]) & (g845) & (g994) & (g1040)) + ((!g847) & (sk[72]) & (g845) & (g994) & (!g1040)) + ((!g847) & (sk[72]) & (g845) & (g994) & (g1040)) + ((g847) & (!sk[72]) & (!g845) & (!g994) & (!g1040)) + ((g847) & (!sk[72]) & (!g845) & (!g994) & (g1040)) + ((g847) & (!sk[72]) & (!g845) & (g994) & (!g1040)) + ((g847) & (!sk[72]) & (!g845) & (g994) & (g1040)) + ((g847) & (!sk[72]) & (g845) & (!g994) & (!g1040)) + ((g847) & (!sk[72]) & (g845) & (!g994) & (g1040)) + ((g847) & (!sk[72]) & (g845) & (g994) & (!g1040)) + ((g847) & (!sk[72]) & (g845) & (g994) & (g1040)) + ((g847) & (sk[72]) & (!g845) & (!g994) & (!g1040)) + ((g847) & (sk[72]) & (!g845) & (g994) & (!g1040)) + ((g847) & (sk[72]) & (g845) & (!g994) & (!g1040)) + ((g847) & (sk[72]) & (g845) & (g994) & (!g1040)) + ((g847) & (sk[72]) & (g845) & (g994) & (g1040)));
	assign g1343 = (((!g252) & (!g843) & (!g848) & (!g971) & (!g1041) & (g1342)) + ((!g252) & (!g843) & (!g848) & (!g971) & (g1041) & (g1342)) + ((!g252) & (!g843) & (!g848) & (g971) & (!g1041) & (g1342)) + ((!g252) & (!g843) & (!g848) & (g971) & (g1041) & (g1342)) + ((!g252) & (!g843) & (g848) & (!g971) & (!g1041) & (g1342)) + ((!g252) & (!g843) & (g848) & (!g971) & (g1041) & (g1342)) + ((!g252) & (!g843) & (g848) & (g971) & (!g1041) & (!g1342)) + ((!g252) & (!g843) & (g848) & (g971) & (!g1041) & (g1342)) + ((!g252) & (!g843) & (g848) & (g971) & (g1041) & (!g1342)) + ((!g252) & (!g843) & (g848) & (g971) & (g1041) & (g1342)) + ((!g252) & (g843) & (!g848) & (!g971) & (!g1041) & (!g1342)) + ((!g252) & (g843) & (!g848) & (!g971) & (!g1041) & (g1342)) + ((!g252) & (g843) & (!g848) & (!g971) & (g1041) & (g1342)) + ((!g252) & (g843) & (!g848) & (g971) & (!g1041) & (!g1342)) + ((!g252) & (g843) & (!g848) & (g971) & (!g1041) & (g1342)) + ((!g252) & (g843) & (!g848) & (g971) & (g1041) & (g1342)) + ((!g252) & (g843) & (g848) & (!g971) & (!g1041) & (!g1342)) + ((!g252) & (g843) & (g848) & (!g971) & (!g1041) & (g1342)) + ((!g252) & (g843) & (g848) & (!g971) & (g1041) & (g1342)) + ((!g252) & (g843) & (g848) & (g971) & (!g1041) & (!g1342)) + ((!g252) & (g843) & (g848) & (g971) & (!g1041) & (g1342)) + ((!g252) & (g843) & (g848) & (g971) & (g1041) & (!g1342)) + ((!g252) & (g843) & (g848) & (g971) & (g1041) & (g1342)) + ((g252) & (!g843) & (!g848) & (!g971) & (!g1041) & (!g1342)) + ((g252) & (!g843) & (!g848) & (!g971) & (g1041) & (!g1342)) + ((g252) & (!g843) & (!g848) & (g971) & (!g1041) & (!g1342)) + ((g252) & (!g843) & (!g848) & (g971) & (g1041) & (!g1342)) + ((g252) & (!g843) & (g848) & (!g971) & (!g1041) & (!g1342)) + ((g252) & (!g843) & (g848) & (!g971) & (g1041) & (!g1342)) + ((g252) & (g843) & (!g848) & (!g971) & (g1041) & (!g1342)) + ((g252) & (g843) & (!g848) & (g971) & (g1041) & (!g1342)) + ((g252) & (g843) & (g848) & (!g971) & (g1041) & (!g1342)));
	assign g1344 = (((!g252) & (!g843) & (!g963) & (!g995) & (!g1327) & (g1328)) + ((!g252) & (!g843) & (!g963) & (g995) & (!g1327) & (g1328)) + ((!g252) & (!g843) & (g963) & (!g995) & (!g1327) & (g1328)) + ((!g252) & (!g843) & (g963) & (g995) & (!g1327) & (g1328)) + ((!g252) & (g843) & (!g963) & (!g995) & (!g1327) & (g1328)) + ((!g252) & (g843) & (g963) & (!g995) & (!g1327) & (g1328)) + ((g252) & (!g843) & (!g963) & (!g995) & (!g1327) & (!g1328)) + ((g252) & (!g843) & (!g963) & (g995) & (!g1327) & (!g1328)) + ((g252) & (!g843) & (g963) & (!g995) & (!g1327) & (!g1328)) + ((g252) & (!g843) & (g963) & (!g995) & (!g1327) & (g1328)) + ((g252) & (!g843) & (g963) & (!g995) & (g1327) & (!g1328)) + ((g252) & (!g843) & (g963) & (g995) & (!g1327) & (!g1328)) + ((g252) & (!g843) & (g963) & (g995) & (!g1327) & (g1328)) + ((g252) & (!g843) & (g963) & (g995) & (g1327) & (!g1328)) + ((g252) & (g843) & (!g963) & (!g995) & (!g1327) & (!g1328)) + ((g252) & (g843) & (!g963) & (g995) & (!g1327) & (!g1328)) + ((g252) & (g843) & (!g963) & (g995) & (!g1327) & (g1328)) + ((g252) & (g843) & (g963) & (!g995) & (!g1327) & (!g1328)) + ((g252) & (g843) & (g963) & (!g995) & (!g1327) & (g1328)) + ((g252) & (g843) & (g963) & (!g995) & (g1327) & (!g1328)) + ((g252) & (g843) & (g963) & (g995) & (!g1327) & (!g1328)) + ((g252) & (g843) & (g963) & (g995) & (!g1327) & (g1328)) + ((g252) & (g843) & (g963) & (g995) & (g1327) & (!g1328)) + ((g252) & (g843) & (g963) & (g995) & (g1327) & (g1328)));
	assign g1345 = (((!g252) & (!g962) & (!g963) & (!g1341) & (!g1343) & (!g1344)) + ((!g252) & (!g962) & (!g963) & (!g1341) & (g1343) & (g1344)) + ((!g252) & (!g962) & (!g963) & (g1341) & (!g1343) & (g1344)) + ((!g252) & (!g962) & (!g963) & (g1341) & (g1343) & (!g1344)) + ((!g252) & (!g962) & (g963) & (!g1341) & (!g1343) & (!g1344)) + ((!g252) & (!g962) & (g963) & (!g1341) & (g1343) & (g1344)) + ((!g252) & (!g962) & (g963) & (g1341) & (!g1343) & (g1344)) + ((!g252) & (!g962) & (g963) & (g1341) & (g1343) & (!g1344)) + ((!g252) & (g962) & (!g963) & (!g1341) & (!g1343) & (!g1344)) + ((!g252) & (g962) & (!g963) & (!g1341) & (g1343) & (g1344)) + ((!g252) & (g962) & (!g963) & (g1341) & (!g1343) & (g1344)) + ((!g252) & (g962) & (!g963) & (g1341) & (g1343) & (!g1344)) + ((!g252) & (g962) & (g963) & (!g1341) & (!g1343) & (!g1344)) + ((!g252) & (g962) & (g963) & (!g1341) & (g1343) & (g1344)) + ((!g252) & (g962) & (g963) & (g1341) & (!g1343) & (g1344)) + ((!g252) & (g962) & (g963) & (g1341) & (g1343) & (!g1344)) + ((g252) & (!g962) & (!g963) & (!g1341) & (!g1343) & (g1344)) + ((g252) & (!g962) & (!g963) & (!g1341) & (g1343) & (!g1344)) + ((g252) & (!g962) & (!g963) & (g1341) & (!g1343) & (!g1344)) + ((g252) & (!g962) & (!g963) & (g1341) & (g1343) & (g1344)) + ((g252) & (!g962) & (g963) & (!g1341) & (!g1343) & (!g1344)) + ((g252) & (!g962) & (g963) & (!g1341) & (g1343) & (g1344)) + ((g252) & (!g962) & (g963) & (g1341) & (!g1343) & (g1344)) + ((g252) & (!g962) & (g963) & (g1341) & (g1343) & (!g1344)) + ((g252) & (g962) & (!g963) & (!g1341) & (!g1343) & (!g1344)) + ((g252) & (g962) & (!g963) & (!g1341) & (g1343) & (g1344)) + ((g252) & (g962) & (!g963) & (g1341) & (!g1343) & (g1344)) + ((g252) & (g962) & (!g963) & (g1341) & (g1343) & (!g1344)) + ((g252) & (g962) & (g963) & (!g1341) & (!g1343) & (g1344)) + ((g252) & (g962) & (g963) & (!g1341) & (g1343) & (!g1344)) + ((g252) & (g962) & (g963) & (g1341) & (!g1343) & (!g1344)) + ((g252) & (g962) & (g963) & (g1341) & (g1343) & (g1344)));
	assign g1346 = (((!sk[76]) & (g1330) & (g1331)) + ((sk[76]) & (g1330) & (!g1331)));
	assign g1347 = (((!g1286) & (!g1287) & (!g1296) & (!g1305) & (g1312) & (!g1332)) + ((!g1286) & (!g1287) & (!g1296) & (g1305) & (!g1312) & (!g1332)) + ((!g1286) & (!g1287) & (!g1296) & (g1305) & (g1312) & (!g1332)) + ((!g1286) & (!g1287) & (g1296) & (g1305) & (g1312) & (!g1332)) + ((!g1286) & (g1287) & (!g1296) & (!g1305) & (g1312) & (!g1332)) + ((!g1286) & (g1287) & (!g1296) & (g1305) & (!g1312) & (!g1332)) + ((!g1286) & (g1287) & (!g1296) & (g1305) & (g1312) & (!g1332)) + ((!g1286) & (g1287) & (g1296) & (!g1305) & (g1312) & (!g1332)) + ((!g1286) & (g1287) & (g1296) & (g1305) & (!g1312) & (!g1332)) + ((!g1286) & (g1287) & (g1296) & (g1305) & (g1312) & (!g1332)) + ((g1286) & (!g1287) & (!g1296) & (g1305) & (g1312) & (!g1332)) + ((g1286) & (!g1287) & (g1296) & (g1305) & (g1312) & (!g1332)) + ((g1286) & (g1287) & (!g1296) & (!g1305) & (g1312) & (!g1332)) + ((g1286) & (g1287) & (!g1296) & (g1305) & (!g1312) & (!g1332)) + ((g1286) & (g1287) & (!g1296) & (g1305) & (g1312) & (!g1332)) + ((g1286) & (g1287) & (g1296) & (g1305) & (g1312) & (!g1332)));
	assign g1348 = (((!sk[78]) & (!g1340) & (!g1345) & (!g1346) & (g1347)) + ((!sk[78]) & (!g1340) & (!g1345) & (g1346) & (g1347)) + ((!sk[78]) & (!g1340) & (g1345) & (!g1346) & (g1347)) + ((!sk[78]) & (!g1340) & (g1345) & (g1346) & (g1347)) + ((!sk[78]) & (g1340) & (!g1345) & (!g1346) & (!g1347)) + ((!sk[78]) & (g1340) & (!g1345) & (!g1346) & (g1347)) + ((!sk[78]) & (g1340) & (!g1345) & (g1346) & (!g1347)) + ((!sk[78]) & (g1340) & (!g1345) & (g1346) & (g1347)) + ((!sk[78]) & (g1340) & (g1345) & (!g1346) & (!g1347)) + ((!sk[78]) & (g1340) & (g1345) & (!g1346) & (g1347)) + ((!sk[78]) & (g1340) & (g1345) & (g1346) & (!g1347)) + ((!sk[78]) & (g1340) & (g1345) & (g1346) & (g1347)) + ((sk[78]) & (!g1340) & (!g1345) & (!g1346) & (!g1347)) + ((sk[78]) & (!g1340) & (g1345) & (!g1346) & (g1347)) + ((sk[78]) & (!g1340) & (g1345) & (g1346) & (!g1347)) + ((sk[78]) & (!g1340) & (g1345) & (g1346) & (g1347)) + ((sk[78]) & (g1340) & (!g1345) & (!g1346) & (g1347)) + ((sk[78]) & (g1340) & (!g1345) & (g1346) & (!g1347)) + ((sk[78]) & (g1340) & (!g1345) & (g1346) & (g1347)) + ((sk[78]) & (g1340) & (g1345) & (!g1346) & (!g1347)));
	assign g1349 = (((!g83) & (!g47) & (!g194) & (!sk[79]) & (g630)) + ((!g83) & (!g47) & (!g194) & (sk[79]) & (g630)) + ((!g83) & (!g47) & (g194) & (!sk[79]) & (g630)) + ((!g83) & (g47) & (!g194) & (!sk[79]) & (g630)) + ((!g83) & (g47) & (g194) & (!sk[79]) & (g630)) + ((g83) & (!g47) & (!g194) & (!sk[79]) & (!g630)) + ((g83) & (!g47) & (!g194) & (!sk[79]) & (g630)) + ((g83) & (!g47) & (g194) & (!sk[79]) & (!g630)) + ((g83) & (!g47) & (g194) & (!sk[79]) & (g630)) + ((g83) & (g47) & (!g194) & (!sk[79]) & (!g630)) + ((g83) & (g47) & (!g194) & (!sk[79]) & (g630)) + ((g83) & (g47) & (g194) & (!sk[79]) & (!g630)) + ((g83) & (g47) & (g194) & (!sk[79]) & (g630)));
	assign g1350 = (((!g9) & (!g12) & (!g146) & (!sk[80]) & (g554) & (!g618)) + ((!g9) & (!g12) & (!g146) & (!sk[80]) & (g554) & (g618)) + ((!g9) & (!g12) & (!g146) & (sk[80]) & (g554) & (g618)) + ((!g9) & (!g12) & (g146) & (!sk[80]) & (!g554) & (!g618)) + ((!g9) & (!g12) & (g146) & (!sk[80]) & (!g554) & (g618)) + ((!g9) & (!g12) & (g146) & (!sk[80]) & (g554) & (!g618)) + ((!g9) & (!g12) & (g146) & (!sk[80]) & (g554) & (g618)) + ((!g9) & (g12) & (!g146) & (!sk[80]) & (!g554) & (!g618)) + ((!g9) & (g12) & (!g146) & (!sk[80]) & (!g554) & (g618)) + ((!g9) & (g12) & (!g146) & (!sk[80]) & (g554) & (!g618)) + ((!g9) & (g12) & (!g146) & (!sk[80]) & (g554) & (g618)) + ((!g9) & (g12) & (!g146) & (sk[80]) & (g554) & (g618)) + ((!g9) & (g12) & (g146) & (!sk[80]) & (!g554) & (!g618)) + ((!g9) & (g12) & (g146) & (!sk[80]) & (!g554) & (g618)) + ((!g9) & (g12) & (g146) & (!sk[80]) & (g554) & (!g618)) + ((!g9) & (g12) & (g146) & (!sk[80]) & (g554) & (g618)) + ((g9) & (!g12) & (!g146) & (!sk[80]) & (g554) & (!g618)) + ((g9) & (!g12) & (!g146) & (!sk[80]) & (g554) & (g618)) + ((g9) & (!g12) & (!g146) & (sk[80]) & (g554) & (g618)) + ((g9) & (!g12) & (g146) & (!sk[80]) & (!g554) & (!g618)) + ((g9) & (!g12) & (g146) & (!sk[80]) & (!g554) & (g618)) + ((g9) & (!g12) & (g146) & (!sk[80]) & (g554) & (!g618)) + ((g9) & (!g12) & (g146) & (!sk[80]) & (g554) & (g618)) + ((g9) & (g12) & (!g146) & (!sk[80]) & (!g554) & (!g618)) + ((g9) & (g12) & (!g146) & (!sk[80]) & (!g554) & (g618)) + ((g9) & (g12) & (!g146) & (!sk[80]) & (g554) & (!g618)) + ((g9) & (g12) & (!g146) & (!sk[80]) & (g554) & (g618)) + ((g9) & (g12) & (g146) & (!sk[80]) & (!g554) & (!g618)) + ((g9) & (g12) & (g146) & (!sk[80]) & (!g554) & (g618)) + ((g9) & (g12) & (g146) & (!sk[80]) & (g554) & (!g618)) + ((g9) & (g12) & (g146) & (!sk[80]) & (g554) & (g618)));
	assign g1351 = (((!g562) & (!g615) & (!sk[81]) & (!g1128) & (g1349) & (!g1350)) + ((!g562) & (!g615) & (!sk[81]) & (!g1128) & (g1349) & (g1350)) + ((!g562) & (!g615) & (!sk[81]) & (g1128) & (!g1349) & (!g1350)) + ((!g562) & (!g615) & (!sk[81]) & (g1128) & (!g1349) & (g1350)) + ((!g562) & (!g615) & (!sk[81]) & (g1128) & (g1349) & (!g1350)) + ((!g562) & (!g615) & (!sk[81]) & (g1128) & (g1349) & (g1350)) + ((!g562) & (g615) & (!sk[81]) & (!g1128) & (!g1349) & (!g1350)) + ((!g562) & (g615) & (!sk[81]) & (!g1128) & (!g1349) & (g1350)) + ((!g562) & (g615) & (!sk[81]) & (!g1128) & (g1349) & (!g1350)) + ((!g562) & (g615) & (!sk[81]) & (!g1128) & (g1349) & (g1350)) + ((!g562) & (g615) & (!sk[81]) & (g1128) & (!g1349) & (!g1350)) + ((!g562) & (g615) & (!sk[81]) & (g1128) & (!g1349) & (g1350)) + ((!g562) & (g615) & (!sk[81]) & (g1128) & (g1349) & (!g1350)) + ((!g562) & (g615) & (!sk[81]) & (g1128) & (g1349) & (g1350)) + ((g562) & (!g615) & (!sk[81]) & (!g1128) & (g1349) & (!g1350)) + ((g562) & (!g615) & (!sk[81]) & (!g1128) & (g1349) & (g1350)) + ((g562) & (!g615) & (!sk[81]) & (g1128) & (!g1349) & (!g1350)) + ((g562) & (!g615) & (!sk[81]) & (g1128) & (!g1349) & (g1350)) + ((g562) & (!g615) & (!sk[81]) & (g1128) & (g1349) & (!g1350)) + ((g562) & (!g615) & (!sk[81]) & (g1128) & (g1349) & (g1350)) + ((g562) & (g615) & (!sk[81]) & (!g1128) & (!g1349) & (!g1350)) + ((g562) & (g615) & (!sk[81]) & (!g1128) & (!g1349) & (g1350)) + ((g562) & (g615) & (!sk[81]) & (!g1128) & (g1349) & (!g1350)) + ((g562) & (g615) & (!sk[81]) & (!g1128) & (g1349) & (g1350)) + ((g562) & (g615) & (!sk[81]) & (g1128) & (!g1349) & (!g1350)) + ((g562) & (g615) & (!sk[81]) & (g1128) & (!g1349) & (g1350)) + ((g562) & (g615) & (!sk[81]) & (g1128) & (g1349) & (!g1350)) + ((g562) & (g615) & (!sk[81]) & (g1128) & (g1349) & (g1350)) + ((g562) & (g615) & (sk[81]) & (g1128) & (g1349) & (g1350)));
	assign g1352 = (((!g1323) & (!g1333) & (!g1335) & (!g1348) & (sk[82]) & (g1351)) + ((!g1323) & (!g1333) & (!g1335) & (g1348) & (!sk[82]) & (!g1351)) + ((!g1323) & (!g1333) & (!g1335) & (g1348) & (!sk[82]) & (g1351)) + ((!g1323) & (!g1333) & (!g1335) & (g1348) & (sk[82]) & (!g1351)) + ((!g1323) & (!g1333) & (g1335) & (!g1348) & (!sk[82]) & (!g1351)) + ((!g1323) & (!g1333) & (g1335) & (!g1348) & (!sk[82]) & (g1351)) + ((!g1323) & (!g1333) & (g1335) & (!g1348) & (sk[82]) & (g1351)) + ((!g1323) & (!g1333) & (g1335) & (g1348) & (!sk[82]) & (!g1351)) + ((!g1323) & (!g1333) & (g1335) & (g1348) & (!sk[82]) & (g1351)) + ((!g1323) & (!g1333) & (g1335) & (g1348) & (sk[82]) & (!g1351)) + ((!g1323) & (g1333) & (!g1335) & (!g1348) & (!sk[82]) & (!g1351)) + ((!g1323) & (g1333) & (!g1335) & (!g1348) & (!sk[82]) & (g1351)) + ((!g1323) & (g1333) & (!g1335) & (!g1348) & (sk[82]) & (g1351)) + ((!g1323) & (g1333) & (!g1335) & (g1348) & (!sk[82]) & (!g1351)) + ((!g1323) & (g1333) & (!g1335) & (g1348) & (!sk[82]) & (g1351)) + ((!g1323) & (g1333) & (!g1335) & (g1348) & (sk[82]) & (!g1351)) + ((!g1323) & (g1333) & (g1335) & (!g1348) & (!sk[82]) & (!g1351)) + ((!g1323) & (g1333) & (g1335) & (!g1348) & (!sk[82]) & (g1351)) + ((!g1323) & (g1333) & (g1335) & (!g1348) & (sk[82]) & (!g1351)) + ((!g1323) & (g1333) & (g1335) & (g1348) & (!sk[82]) & (!g1351)) + ((!g1323) & (g1333) & (g1335) & (g1348) & (!sk[82]) & (g1351)) + ((!g1323) & (g1333) & (g1335) & (g1348) & (sk[82]) & (g1351)) + ((g1323) & (!g1333) & (!g1335) & (!g1348) & (sk[82]) & (g1351)) + ((g1323) & (!g1333) & (!g1335) & (g1348) & (!sk[82]) & (!g1351)) + ((g1323) & (!g1333) & (!g1335) & (g1348) & (!sk[82]) & (g1351)) + ((g1323) & (!g1333) & (!g1335) & (g1348) & (sk[82]) & (!g1351)) + ((g1323) & (!g1333) & (g1335) & (!g1348) & (!sk[82]) & (!g1351)) + ((g1323) & (!g1333) & (g1335) & (!g1348) & (!sk[82]) & (g1351)) + ((g1323) & (!g1333) & (g1335) & (!g1348) & (sk[82]) & (!g1351)) + ((g1323) & (!g1333) & (g1335) & (g1348) & (!sk[82]) & (!g1351)) + ((g1323) & (!g1333) & (g1335) & (g1348) & (!sk[82]) & (g1351)) + ((g1323) & (!g1333) & (g1335) & (g1348) & (sk[82]) & (g1351)) + ((g1323) & (g1333) & (!g1335) & (!g1348) & (!sk[82]) & (!g1351)) + ((g1323) & (g1333) & (!g1335) & (!g1348) & (!sk[82]) & (g1351)) + ((g1323) & (g1333) & (!g1335) & (!g1348) & (sk[82]) & (!g1351)) + ((g1323) & (g1333) & (!g1335) & (g1348) & (!sk[82]) & (!g1351)) + ((g1323) & (g1333) & (!g1335) & (g1348) & (!sk[82]) & (g1351)) + ((g1323) & (g1333) & (!g1335) & (g1348) & (sk[82]) & (g1351)) + ((g1323) & (g1333) & (g1335) & (!g1348) & (!sk[82]) & (!g1351)) + ((g1323) & (g1333) & (g1335) & (!g1348) & (!sk[82]) & (g1351)) + ((g1323) & (g1333) & (g1335) & (!g1348) & (sk[82]) & (!g1351)) + ((g1323) & (g1333) & (g1335) & (g1348) & (!sk[82]) & (!g1351)) + ((g1323) & (g1333) & (g1335) & (g1348) & (!sk[82]) & (g1351)) + ((g1323) & (g1333) & (g1335) & (g1348) & (sk[82]) & (g1351)));
	assign sinx12x = (((!sk[83]) & (!g1068) & (!g1321) & (!g1337) & (g1338) & (!g1352)) + ((!sk[83]) & (!g1068) & (!g1321) & (!g1337) & (g1338) & (g1352)) + ((!sk[83]) & (!g1068) & (!g1321) & (g1337) & (!g1338) & (!g1352)) + ((!sk[83]) & (!g1068) & (!g1321) & (g1337) & (!g1338) & (g1352)) + ((!sk[83]) & (!g1068) & (!g1321) & (g1337) & (g1338) & (!g1352)) + ((!sk[83]) & (!g1068) & (!g1321) & (g1337) & (g1338) & (g1352)) + ((!sk[83]) & (!g1068) & (g1321) & (!g1337) & (!g1338) & (!g1352)) + ((!sk[83]) & (!g1068) & (g1321) & (!g1337) & (!g1338) & (g1352)) + ((!sk[83]) & (!g1068) & (g1321) & (!g1337) & (g1338) & (!g1352)) + ((!sk[83]) & (!g1068) & (g1321) & (!g1337) & (g1338) & (g1352)) + ((!sk[83]) & (!g1068) & (g1321) & (g1337) & (!g1338) & (!g1352)) + ((!sk[83]) & (!g1068) & (g1321) & (g1337) & (!g1338) & (g1352)) + ((!sk[83]) & (!g1068) & (g1321) & (g1337) & (g1338) & (!g1352)) + ((!sk[83]) & (!g1068) & (g1321) & (g1337) & (g1338) & (g1352)) + ((!sk[83]) & (g1068) & (!g1321) & (!g1337) & (g1338) & (!g1352)) + ((!sk[83]) & (g1068) & (!g1321) & (!g1337) & (g1338) & (g1352)) + ((!sk[83]) & (g1068) & (!g1321) & (g1337) & (!g1338) & (!g1352)) + ((!sk[83]) & (g1068) & (!g1321) & (g1337) & (!g1338) & (g1352)) + ((!sk[83]) & (g1068) & (!g1321) & (g1337) & (g1338) & (!g1352)) + ((!sk[83]) & (g1068) & (!g1321) & (g1337) & (g1338) & (g1352)) + ((!sk[83]) & (g1068) & (g1321) & (!g1337) & (!g1338) & (!g1352)) + ((!sk[83]) & (g1068) & (g1321) & (!g1337) & (!g1338) & (g1352)) + ((!sk[83]) & (g1068) & (g1321) & (!g1337) & (g1338) & (!g1352)) + ((!sk[83]) & (g1068) & (g1321) & (!g1337) & (g1338) & (g1352)) + ((!sk[83]) & (g1068) & (g1321) & (g1337) & (!g1338) & (!g1352)) + ((!sk[83]) & (g1068) & (g1321) & (g1337) & (!g1338) & (g1352)) + ((!sk[83]) & (g1068) & (g1321) & (g1337) & (g1338) & (!g1352)) + ((!sk[83]) & (g1068) & (g1321) & (g1337) & (g1338) & (g1352)) + ((sk[83]) & (!g1068) & (!g1321) & (!g1337) & (!g1338) & (g1352)) + ((sk[83]) & (!g1068) & (!g1321) & (!g1337) & (g1338) & (g1352)) + ((sk[83]) & (!g1068) & (!g1321) & (g1337) & (!g1338) & (g1352)) + ((sk[83]) & (!g1068) & (!g1321) & (g1337) & (g1338) & (g1352)) + ((sk[83]) & (!g1068) & (g1321) & (!g1337) & (!g1338) & (!g1352)) + ((sk[83]) & (!g1068) & (g1321) & (!g1337) & (g1338) & (!g1352)) + ((sk[83]) & (!g1068) & (g1321) & (g1337) & (!g1338) & (g1352)) + ((sk[83]) & (!g1068) & (g1321) & (g1337) & (g1338) & (g1352)) + ((sk[83]) & (g1068) & (!g1321) & (!g1337) & (!g1338) & (!g1352)) + ((sk[83]) & (g1068) & (!g1321) & (!g1337) & (g1338) & (!g1352)) + ((sk[83]) & (g1068) & (!g1321) & (g1337) & (!g1338) & (!g1352)) + ((sk[83]) & (g1068) & (!g1321) & (g1337) & (g1338) & (g1352)) + ((sk[83]) & (g1068) & (g1321) & (!g1337) & (!g1338) & (g1352)) + ((sk[83]) & (g1068) & (g1321) & (!g1337) & (g1338) & (!g1352)) + ((sk[83]) & (g1068) & (g1321) & (g1337) & (!g1338) & (!g1352)) + ((sk[83]) & (g1068) & (g1321) & (g1337) & (g1338) & (!g1352)));
	assign g1354 = (((!sk[84]) & (!g1321) & (!g1337) & (!g1338) & (g1352)) + ((!sk[84]) & (!g1321) & (!g1337) & (g1338) & (g1352)) + ((!sk[84]) & (!g1321) & (g1337) & (!g1338) & (g1352)) + ((!sk[84]) & (!g1321) & (g1337) & (g1338) & (g1352)) + ((!sk[84]) & (g1321) & (!g1337) & (!g1338) & (!g1352)) + ((!sk[84]) & (g1321) & (!g1337) & (!g1338) & (g1352)) + ((!sk[84]) & (g1321) & (!g1337) & (g1338) & (!g1352)) + ((!sk[84]) & (g1321) & (!g1337) & (g1338) & (g1352)) + ((!sk[84]) & (g1321) & (g1337) & (!g1338) & (!g1352)) + ((!sk[84]) & (g1321) & (g1337) & (!g1338) & (g1352)) + ((!sk[84]) & (g1321) & (g1337) & (g1338) & (!g1352)) + ((!sk[84]) & (g1321) & (g1337) & (g1338) & (g1352)) + ((sk[84]) & (!g1321) & (g1337) & (g1338) & (!g1352)) + ((sk[84]) & (g1321) & (!g1337) & (g1338) & (g1352)));
	assign g1355 = (((!g1320) & (!g1304) & (!g1322) & (g1317) & (!sk[85]) & (!g1336)) + ((!g1320) & (!g1304) & (!g1322) & (g1317) & (!sk[85]) & (g1336)) + ((!g1320) & (!g1304) & (g1322) & (!g1317) & (!sk[85]) & (!g1336)) + ((!g1320) & (!g1304) & (g1322) & (!g1317) & (!sk[85]) & (g1336)) + ((!g1320) & (!g1304) & (g1322) & (g1317) & (!sk[85]) & (!g1336)) + ((!g1320) & (!g1304) & (g1322) & (g1317) & (!sk[85]) & (g1336)) + ((!g1320) & (g1304) & (!g1322) & (!g1317) & (!sk[85]) & (!g1336)) + ((!g1320) & (g1304) & (!g1322) & (!g1317) & (!sk[85]) & (g1336)) + ((!g1320) & (g1304) & (!g1322) & (g1317) & (!sk[85]) & (!g1336)) + ((!g1320) & (g1304) & (!g1322) & (g1317) & (!sk[85]) & (g1336)) + ((!g1320) & (g1304) & (g1322) & (!g1317) & (!sk[85]) & (!g1336)) + ((!g1320) & (g1304) & (g1322) & (!g1317) & (!sk[85]) & (g1336)) + ((!g1320) & (g1304) & (g1322) & (g1317) & (!sk[85]) & (!g1336)) + ((!g1320) & (g1304) & (g1322) & (g1317) & (!sk[85]) & (g1336)) + ((g1320) & (!g1304) & (!g1322) & (g1317) & (!sk[85]) & (!g1336)) + ((g1320) & (!g1304) & (!g1322) & (g1317) & (!sk[85]) & (g1336)) + ((g1320) & (!g1304) & (!g1322) & (g1317) & (sk[85]) & (!g1336)) + ((g1320) & (!g1304) & (g1322) & (!g1317) & (!sk[85]) & (!g1336)) + ((g1320) & (!g1304) & (g1322) & (!g1317) & (!sk[85]) & (g1336)) + ((g1320) & (!g1304) & (g1322) & (!g1317) & (sk[85]) & (g1336)) + ((g1320) & (!g1304) & (g1322) & (g1317) & (!sk[85]) & (!g1336)) + ((g1320) & (!g1304) & (g1322) & (g1317) & (!sk[85]) & (g1336)) + ((g1320) & (g1304) & (!g1322) & (!g1317) & (!sk[85]) & (!g1336)) + ((g1320) & (g1304) & (!g1322) & (!g1317) & (!sk[85]) & (g1336)) + ((g1320) & (g1304) & (!g1322) & (!g1317) & (sk[85]) & (!g1336)) + ((g1320) & (g1304) & (!g1322) & (g1317) & (!sk[85]) & (!g1336)) + ((g1320) & (g1304) & (!g1322) & (g1317) & (!sk[85]) & (g1336)) + ((g1320) & (g1304) & (g1322) & (!g1317) & (!sk[85]) & (!g1336)) + ((g1320) & (g1304) & (g1322) & (!g1317) & (!sk[85]) & (g1336)) + ((g1320) & (g1304) & (g1322) & (g1317) & (!sk[85]) & (!g1336)) + ((g1320) & (g1304) & (g1322) & (g1317) & (!sk[85]) & (g1336)) + ((g1320) & (g1304) & (g1322) & (g1317) & (sk[85]) & (!g1336)));
	assign g1356 = (((!g252) & (!g962) & (!g963) & (!g1341) & (g1343) & (g1344)) + ((!g252) & (!g962) & (!g963) & (g1341) & (!g1343) & (g1344)) + ((!g252) & (!g962) & (!g963) & (g1341) & (g1343) & (!g1344)) + ((!g252) & (!g962) & (!g963) & (g1341) & (g1343) & (g1344)) + ((!g252) & (!g962) & (g963) & (!g1341) & (g1343) & (g1344)) + ((!g252) & (!g962) & (g963) & (g1341) & (!g1343) & (g1344)) + ((!g252) & (!g962) & (g963) & (g1341) & (g1343) & (!g1344)) + ((!g252) & (!g962) & (g963) & (g1341) & (g1343) & (g1344)) + ((!g252) & (g962) & (!g963) & (!g1341) & (g1343) & (g1344)) + ((!g252) & (g962) & (!g963) & (g1341) & (!g1343) & (g1344)) + ((!g252) & (g962) & (!g963) & (g1341) & (g1343) & (!g1344)) + ((!g252) & (g962) & (!g963) & (g1341) & (g1343) & (g1344)) + ((!g252) & (g962) & (g963) & (!g1341) & (g1343) & (g1344)) + ((!g252) & (g962) & (g963) & (g1341) & (!g1343) & (g1344)) + ((!g252) & (g962) & (g963) & (g1341) & (g1343) & (!g1344)) + ((!g252) & (g962) & (g963) & (g1341) & (g1343) & (g1344)) + ((g252) & (!g962) & (!g963) & (!g1341) & (g1343) & (!g1344)) + ((g252) & (!g962) & (!g963) & (g1341) & (!g1343) & (!g1344)) + ((g252) & (!g962) & (!g963) & (g1341) & (g1343) & (!g1344)) + ((g252) & (!g962) & (!g963) & (g1341) & (g1343) & (g1344)) + ((g252) & (!g962) & (g963) & (!g1341) & (g1343) & (g1344)) + ((g252) & (!g962) & (g963) & (g1341) & (!g1343) & (g1344)) + ((g252) & (!g962) & (g963) & (g1341) & (g1343) & (!g1344)) + ((g252) & (!g962) & (g963) & (g1341) & (g1343) & (g1344)) + ((g252) & (g962) & (!g963) & (!g1341) & (g1343) & (g1344)) + ((g252) & (g962) & (!g963) & (g1341) & (!g1343) & (g1344)) + ((g252) & (g962) & (!g963) & (g1341) & (g1343) & (!g1344)) + ((g252) & (g962) & (!g963) & (g1341) & (g1343) & (g1344)) + ((g252) & (g962) & (g963) & (!g1341) & (g1343) & (!g1344)) + ((g252) & (g962) & (g963) & (g1341) & (!g1343) & (!g1344)) + ((g252) & (g962) & (g963) & (g1341) & (g1343) & (!g1344)) + ((g252) & (g962) & (g963) & (g1341) & (g1343) & (g1344)));
	assign g1357 = (((!g847) & (!g845) & (!g848) & (!g994) & (!g1040) & (!g1079)) + ((!g847) & (!g845) & (!g848) & (!g994) & (!g1040) & (g1079)) + ((!g847) & (!g845) & (!g848) & (!g994) & (g1040) & (!g1079)) + ((!g847) & (!g845) & (!g848) & (!g994) & (g1040) & (g1079)) + ((!g847) & (!g845) & (!g848) & (g994) & (!g1040) & (!g1079)) + ((!g847) & (!g845) & (!g848) & (g994) & (!g1040) & (g1079)) + ((!g847) & (!g845) & (!g848) & (g994) & (g1040) & (!g1079)) + ((!g847) & (!g845) & (!g848) & (g994) & (g1040) & (g1079)) + ((!g847) & (!g845) & (g848) & (!g994) & (!g1040) & (!g1079)) + ((!g847) & (!g845) & (g848) & (!g994) & (!g1040) & (g1079)) + ((!g847) & (!g845) & (g848) & (!g994) & (g1040) & (!g1079)) + ((!g847) & (!g845) & (g848) & (!g994) & (g1040) & (g1079)) + ((!g847) & (g845) & (!g848) & (!g994) & (g1040) & (!g1079)) + ((!g847) & (g845) & (!g848) & (!g994) & (g1040) & (g1079)) + ((!g847) & (g845) & (!g848) & (g994) & (g1040) & (!g1079)) + ((!g847) & (g845) & (!g848) & (g994) & (g1040) & (g1079)) + ((!g847) & (g845) & (g848) & (!g994) & (g1040) & (!g1079)) + ((!g847) & (g845) & (g848) & (!g994) & (g1040) & (g1079)) + ((g847) & (!g845) & (!g848) & (!g994) & (!g1040) & (g1079)) + ((g847) & (!g845) & (!g848) & (!g994) & (g1040) & (g1079)) + ((g847) & (!g845) & (!g848) & (g994) & (!g1040) & (g1079)) + ((g847) & (!g845) & (!g848) & (g994) & (g1040) & (g1079)) + ((g847) & (!g845) & (g848) & (!g994) & (!g1040) & (g1079)) + ((g847) & (!g845) & (g848) & (!g994) & (g1040) & (g1079)) + ((g847) & (g845) & (!g848) & (!g994) & (g1040) & (g1079)) + ((g847) & (g845) & (!g848) & (g994) & (g1040) & (g1079)) + ((g847) & (g845) & (g848) & (!g994) & (g1040) & (g1079)));
	assign g1358 = (((!g252) & (!g843) & (!g1040) & (!g1079) & (!g1080) & (!g1357)) + ((!g252) & (!g843) & (!g1040) & (!g1079) & (g1080) & (!g1357)) + ((!g252) & (!g843) & (!g1040) & (g1079) & (!g1080) & (!g1357)) + ((!g252) & (!g843) & (!g1040) & (g1079) & (g1080) & (!g1357)) + ((!g252) & (!g843) & (g1040) & (!g1079) & (!g1080) & (!g1357)) + ((!g252) & (!g843) & (g1040) & (!g1079) & (g1080) & (!g1357)) + ((!g252) & (!g843) & (g1040) & (g1079) & (!g1080) & (!g1357)) + ((!g252) & (!g843) & (g1040) & (g1079) & (g1080) & (!g1357)) + ((!g252) & (g843) & (!g1040) & (!g1079) & (!g1080) & (!g1357)) + ((!g252) & (g843) & (!g1040) & (!g1079) & (g1080) & (!g1357)) + ((!g252) & (g843) & (!g1040) & (!g1079) & (g1080) & (g1357)) + ((!g252) & (g843) & (!g1040) & (g1079) & (!g1080) & (!g1357)) + ((!g252) & (g843) & (!g1040) & (g1079) & (!g1080) & (g1357)) + ((!g252) & (g843) & (!g1040) & (g1079) & (g1080) & (!g1357)) + ((!g252) & (g843) & (g1040) & (!g1079) & (!g1080) & (!g1357)) + ((!g252) & (g843) & (g1040) & (!g1079) & (!g1080) & (g1357)) + ((!g252) & (g843) & (g1040) & (!g1079) & (g1080) & (!g1357)) + ((!g252) & (g843) & (g1040) & (g1079) & (!g1080) & (!g1357)) + ((!g252) & (g843) & (g1040) & (g1079) & (g1080) & (!g1357)) + ((!g252) & (g843) & (g1040) & (g1079) & (g1080) & (g1357)) + ((g252) & (!g843) & (!g1040) & (!g1079) & (!g1080) & (g1357)) + ((g252) & (!g843) & (!g1040) & (!g1079) & (g1080) & (g1357)) + ((g252) & (!g843) & (!g1040) & (g1079) & (!g1080) & (g1357)) + ((g252) & (!g843) & (!g1040) & (g1079) & (g1080) & (g1357)) + ((g252) & (!g843) & (g1040) & (!g1079) & (!g1080) & (g1357)) + ((g252) & (!g843) & (g1040) & (!g1079) & (g1080) & (g1357)) + ((g252) & (!g843) & (g1040) & (g1079) & (!g1080) & (g1357)) + ((g252) & (!g843) & (g1040) & (g1079) & (g1080) & (g1357)) + ((g252) & (g843) & (!g1040) & (!g1079) & (!g1080) & (g1357)) + ((g252) & (g843) & (!g1040) & (g1079) & (g1080) & (g1357)) + ((g252) & (g843) & (g1040) & (!g1079) & (g1080) & (g1357)) + ((g252) & (g843) & (g1040) & (g1079) & (!g1080) & (g1357)));
	assign g1359 = (((!sk[89]) & (!g202) & (!g252) & (!g962) & (g971)) + ((!sk[89]) & (!g202) & (!g252) & (g962) & (g971)) + ((!sk[89]) & (!g202) & (g252) & (!g962) & (g971)) + ((!sk[89]) & (!g202) & (g252) & (g962) & (g971)) + ((!sk[89]) & (g202) & (!g252) & (!g962) & (!g971)) + ((!sk[89]) & (g202) & (!g252) & (!g962) & (g971)) + ((!sk[89]) & (g202) & (!g252) & (g962) & (!g971)) + ((!sk[89]) & (g202) & (!g252) & (g962) & (g971)) + ((!sk[89]) & (g202) & (g252) & (!g962) & (!g971)) + ((!sk[89]) & (g202) & (g252) & (!g962) & (g971)) + ((!sk[89]) & (g202) & (g252) & (g962) & (!g971)) + ((!sk[89]) & (g202) & (g252) & (g962) & (g971)) + ((sk[89]) & (!g202) & (g252) & (!g962) & (!g971)) + ((sk[89]) & (!g202) & (g252) & (g962) & (g971)) + ((sk[89]) & (g202) & (!g252) & (!g962) & (!g971)) + ((sk[89]) & (g202) & (!g252) & (!g962) & (g971)) + ((sk[89]) & (g202) & (!g252) & (g962) & (!g971)) + ((sk[89]) & (g202) & (!g252) & (g962) & (g971)) + ((sk[89]) & (g202) & (g252) & (!g962) & (g971)) + ((sk[89]) & (g202) & (g252) & (g962) & (!g971)));
	assign g1360 = (((!g252) & (!g962) & (!g963) & (!g1344) & (!g1358) & (g1359)) + ((!g252) & (!g962) & (!g963) & (!g1344) & (g1358) & (!g1359)) + ((!g252) & (!g962) & (!g963) & (g1344) & (!g1358) & (!g1359)) + ((!g252) & (!g962) & (!g963) & (g1344) & (g1358) & (g1359)) + ((!g252) & (!g962) & (g963) & (!g1344) & (!g1358) & (g1359)) + ((!g252) & (!g962) & (g963) & (!g1344) & (g1358) & (!g1359)) + ((!g252) & (!g962) & (g963) & (g1344) & (!g1358) & (!g1359)) + ((!g252) & (!g962) & (g963) & (g1344) & (g1358) & (g1359)) + ((!g252) & (g962) & (!g963) & (!g1344) & (!g1358) & (g1359)) + ((!g252) & (g962) & (!g963) & (!g1344) & (g1358) & (!g1359)) + ((!g252) & (g962) & (!g963) & (g1344) & (!g1358) & (!g1359)) + ((!g252) & (g962) & (!g963) & (g1344) & (g1358) & (g1359)) + ((!g252) & (g962) & (g963) & (!g1344) & (!g1358) & (g1359)) + ((!g252) & (g962) & (g963) & (!g1344) & (g1358) & (!g1359)) + ((!g252) & (g962) & (g963) & (g1344) & (!g1358) & (!g1359)) + ((!g252) & (g962) & (g963) & (g1344) & (g1358) & (g1359)) + ((g252) & (!g962) & (!g963) & (!g1344) & (!g1358) & (!g1359)) + ((g252) & (!g962) & (!g963) & (!g1344) & (g1358) & (g1359)) + ((g252) & (!g962) & (!g963) & (g1344) & (!g1358) & (!g1359)) + ((g252) & (!g962) & (!g963) & (g1344) & (g1358) & (g1359)) + ((g252) & (!g962) & (g963) & (!g1344) & (!g1358) & (g1359)) + ((g252) & (!g962) & (g963) & (!g1344) & (g1358) & (!g1359)) + ((g252) & (!g962) & (g963) & (g1344) & (!g1358) & (!g1359)) + ((g252) & (!g962) & (g963) & (g1344) & (g1358) & (g1359)) + ((g252) & (g962) & (!g963) & (!g1344) & (!g1358) & (g1359)) + ((g252) & (g962) & (!g963) & (!g1344) & (g1358) & (!g1359)) + ((g252) & (g962) & (!g963) & (g1344) & (!g1358) & (!g1359)) + ((g252) & (g962) & (!g963) & (g1344) & (g1358) & (g1359)) + ((g252) & (g962) & (g963) & (!g1344) & (!g1358) & (g1359)) + ((g252) & (g962) & (g963) & (!g1344) & (g1358) & (!g1359)) + ((g252) & (g962) & (g963) & (g1344) & (!g1358) & (g1359)) + ((g252) & (g962) & (g963) & (g1344) & (g1358) & (!g1359)));
	assign g1361 = (((!g1356) & (sk[91]) & (g1360)) + ((g1356) & (!sk[91]) & (g1360)) + ((g1356) & (sk[91]) & (!g1360)));
	assign g1362 = (((!sk[92]) & (!g1340) & (!g1345) & (!g1346) & (g1347) & (!g1361)) + ((!sk[92]) & (!g1340) & (!g1345) & (!g1346) & (g1347) & (g1361)) + ((!sk[92]) & (!g1340) & (!g1345) & (g1346) & (!g1347) & (!g1361)) + ((!sk[92]) & (!g1340) & (!g1345) & (g1346) & (!g1347) & (g1361)) + ((!sk[92]) & (!g1340) & (!g1345) & (g1346) & (g1347) & (!g1361)) + ((!sk[92]) & (!g1340) & (!g1345) & (g1346) & (g1347) & (g1361)) + ((!sk[92]) & (!g1340) & (g1345) & (!g1346) & (!g1347) & (!g1361)) + ((!sk[92]) & (!g1340) & (g1345) & (!g1346) & (!g1347) & (g1361)) + ((!sk[92]) & (!g1340) & (g1345) & (!g1346) & (g1347) & (!g1361)) + ((!sk[92]) & (!g1340) & (g1345) & (!g1346) & (g1347) & (g1361)) + ((!sk[92]) & (!g1340) & (g1345) & (g1346) & (!g1347) & (!g1361)) + ((!sk[92]) & (!g1340) & (g1345) & (g1346) & (!g1347) & (g1361)) + ((!sk[92]) & (!g1340) & (g1345) & (g1346) & (g1347) & (!g1361)) + ((!sk[92]) & (!g1340) & (g1345) & (g1346) & (g1347) & (g1361)) + ((!sk[92]) & (g1340) & (!g1345) & (!g1346) & (g1347) & (!g1361)) + ((!sk[92]) & (g1340) & (!g1345) & (!g1346) & (g1347) & (g1361)) + ((!sk[92]) & (g1340) & (!g1345) & (g1346) & (!g1347) & (!g1361)) + ((!sk[92]) & (g1340) & (!g1345) & (g1346) & (!g1347) & (g1361)) + ((!sk[92]) & (g1340) & (!g1345) & (g1346) & (g1347) & (!g1361)) + ((!sk[92]) & (g1340) & (!g1345) & (g1346) & (g1347) & (g1361)) + ((!sk[92]) & (g1340) & (g1345) & (!g1346) & (!g1347) & (!g1361)) + ((!sk[92]) & (g1340) & (g1345) & (!g1346) & (!g1347) & (g1361)) + ((!sk[92]) & (g1340) & (g1345) & (!g1346) & (g1347) & (!g1361)) + ((!sk[92]) & (g1340) & (g1345) & (!g1346) & (g1347) & (g1361)) + ((!sk[92]) & (g1340) & (g1345) & (g1346) & (!g1347) & (!g1361)) + ((!sk[92]) & (g1340) & (g1345) & (g1346) & (!g1347) & (g1361)) + ((!sk[92]) & (g1340) & (g1345) & (g1346) & (g1347) & (!g1361)) + ((!sk[92]) & (g1340) & (g1345) & (g1346) & (g1347) & (g1361)) + ((sk[92]) & (!g1340) & (!g1345) & (!g1346) & (!g1347) & (!g1361)) + ((sk[92]) & (!g1340) & (!g1345) & (!g1346) & (g1347) & (g1361)) + ((sk[92]) & (!g1340) & (!g1345) & (g1346) & (!g1347) & (g1361)) + ((sk[92]) & (!g1340) & (!g1345) & (g1346) & (g1347) & (g1361)) + ((sk[92]) & (!g1340) & (g1345) & (!g1346) & (!g1347) & (!g1361)) + ((sk[92]) & (!g1340) & (g1345) & (!g1346) & (g1347) & (!g1361)) + ((sk[92]) & (!g1340) & (g1345) & (g1346) & (!g1347) & (!g1361)) + ((sk[92]) & (!g1340) & (g1345) & (g1346) & (g1347) & (!g1361)) + ((sk[92]) & (g1340) & (!g1345) & (!g1346) & (!g1347) & (g1361)) + ((sk[92]) & (g1340) & (!g1345) & (!g1346) & (g1347) & (g1361)) + ((sk[92]) & (g1340) & (!g1345) & (g1346) & (!g1347) & (g1361)) + ((sk[92]) & (g1340) & (!g1345) & (g1346) & (g1347) & (g1361)) + ((sk[92]) & (g1340) & (g1345) & (!g1346) & (!g1347) & (!g1361)) + ((sk[92]) & (g1340) & (g1345) & (!g1346) & (g1347) & (g1361)) + ((sk[92]) & (g1340) & (g1345) & (g1346) & (!g1347) & (g1361)) + ((sk[92]) & (g1340) & (g1345) & (g1346) & (g1347) & (g1361)));
	assign g1363 = (((!g9) & (!g10) & (!g16) & (!g62) & (!g42) & (!g133)) + ((!g9) & (!g10) & (!g16) & (!g62) & (!g42) & (g133)) + ((!g9) & (!g10) & (!g16) & (!g62) & (g42) & (!g133)) + ((!g9) & (!g10) & (!g16) & (!g62) & (g42) & (g133)) + ((!g9) & (!g10) & (!g16) & (g62) & (!g42) & (!g133)) + ((!g9) & (!g10) & (!g16) & (g62) & (!g42) & (g133)) + ((!g9) & (!g10) & (g16) & (!g62) & (!g42) & (!g133)) + ((!g9) & (!g10) & (g16) & (g62) & (!g42) & (!g133)) + ((!g9) & (g10) & (!g16) & (!g62) & (!g42) & (!g133)) + ((!g9) & (g10) & (!g16) & (!g62) & (!g42) & (g133)) + ((!g9) & (g10) & (!g16) & (!g62) & (g42) & (!g133)) + ((!g9) & (g10) & (!g16) & (!g62) & (g42) & (g133)) + ((!g9) & (g10) & (!g16) & (g62) & (!g42) & (!g133)) + ((!g9) & (g10) & (!g16) & (g62) & (!g42) & (g133)) + ((!g9) & (g10) & (g16) & (!g62) & (!g42) & (!g133)) + ((!g9) & (g10) & (g16) & (g62) & (!g42) & (!g133)) + ((g9) & (!g10) & (!g16) & (!g62) & (!g42) & (!g133)) + ((g9) & (!g10) & (!g16) & (g62) & (!g42) & (!g133)) + ((g9) & (!g10) & (g16) & (!g62) & (!g42) & (!g133)) + ((g9) & (!g10) & (g16) & (g62) & (!g42) & (!g133)));
	assign g1364 = (((!g297) & (!sk[94]) & (!g177) & (!g1073) & (g1363)) + ((!g297) & (!sk[94]) & (!g177) & (g1073) & (g1363)) + ((!g297) & (!sk[94]) & (g177) & (!g1073) & (g1363)) + ((!g297) & (!sk[94]) & (g177) & (g1073) & (g1363)) + ((!g297) & (sk[94]) & (!g177) & (g1073) & (g1363)) + ((g297) & (!sk[94]) & (!g177) & (!g1073) & (!g1363)) + ((g297) & (!sk[94]) & (!g177) & (!g1073) & (g1363)) + ((g297) & (!sk[94]) & (!g177) & (g1073) & (!g1363)) + ((g297) & (!sk[94]) & (!g177) & (g1073) & (g1363)) + ((g297) & (!sk[94]) & (g177) & (!g1073) & (!g1363)) + ((g297) & (!sk[94]) & (g177) & (!g1073) & (g1363)) + ((g297) & (!sk[94]) & (g177) & (g1073) & (!g1363)) + ((g297) & (!sk[94]) & (g177) & (g1073) & (g1363)));
	assign g1365 = (((!g703) & (!g829) & (!sk[95]) & (!g1028) & (g1364)) + ((!g703) & (!g829) & (!sk[95]) & (g1028) & (g1364)) + ((!g703) & (g829) & (!sk[95]) & (!g1028) & (g1364)) + ((!g703) & (g829) & (!sk[95]) & (g1028) & (g1364)) + ((g703) & (!g829) & (!sk[95]) & (!g1028) & (!g1364)) + ((g703) & (!g829) & (!sk[95]) & (!g1028) & (g1364)) + ((g703) & (!g829) & (!sk[95]) & (g1028) & (!g1364)) + ((g703) & (!g829) & (!sk[95]) & (g1028) & (g1364)) + ((g703) & (g829) & (!sk[95]) & (!g1028) & (!g1364)) + ((g703) & (g829) & (!sk[95]) & (!g1028) & (g1364)) + ((g703) & (g829) & (!sk[95]) & (g1028) & (!g1364)) + ((g703) & (g829) & (!sk[95]) & (g1028) & (g1364)) + ((g703) & (g829) & (sk[95]) & (g1028) & (g1364)));
	assign g1366 = (((!g1323) & (!sk[96]) & (!g1333) & (!g1335) & (g1348) & (!g1351)) + ((!g1323) & (!sk[96]) & (!g1333) & (!g1335) & (g1348) & (g1351)) + ((!g1323) & (!sk[96]) & (!g1333) & (g1335) & (!g1348) & (!g1351)) + ((!g1323) & (!sk[96]) & (!g1333) & (g1335) & (!g1348) & (g1351)) + ((!g1323) & (!sk[96]) & (!g1333) & (g1335) & (g1348) & (!g1351)) + ((!g1323) & (!sk[96]) & (!g1333) & (g1335) & (g1348) & (g1351)) + ((!g1323) & (!sk[96]) & (g1333) & (!g1335) & (!g1348) & (!g1351)) + ((!g1323) & (!sk[96]) & (g1333) & (!g1335) & (!g1348) & (g1351)) + ((!g1323) & (!sk[96]) & (g1333) & (!g1335) & (g1348) & (!g1351)) + ((!g1323) & (!sk[96]) & (g1333) & (!g1335) & (g1348) & (g1351)) + ((!g1323) & (!sk[96]) & (g1333) & (g1335) & (!g1348) & (!g1351)) + ((!g1323) & (!sk[96]) & (g1333) & (g1335) & (!g1348) & (g1351)) + ((!g1323) & (!sk[96]) & (g1333) & (g1335) & (g1348) & (!g1351)) + ((!g1323) & (!sk[96]) & (g1333) & (g1335) & (g1348) & (g1351)) + ((!g1323) & (sk[96]) & (!g1333) & (!g1335) & (!g1348) & (!g1351)) + ((!g1323) & (sk[96]) & (!g1333) & (!g1335) & (g1348) & (!g1351)) + ((!g1323) & (sk[96]) & (!g1333) & (!g1335) & (g1348) & (g1351)) + ((!g1323) & (sk[96]) & (!g1333) & (g1335) & (!g1348) & (!g1351)) + ((!g1323) & (sk[96]) & (!g1333) & (g1335) & (g1348) & (!g1351)) + ((!g1323) & (sk[96]) & (!g1333) & (g1335) & (g1348) & (g1351)) + ((!g1323) & (sk[96]) & (g1333) & (!g1335) & (!g1348) & (!g1351)) + ((!g1323) & (sk[96]) & (g1333) & (!g1335) & (g1348) & (!g1351)) + ((!g1323) & (sk[96]) & (g1333) & (!g1335) & (g1348) & (g1351)) + ((!g1323) & (sk[96]) & (g1333) & (g1335) & (g1348) & (!g1351)) + ((g1323) & (!sk[96]) & (!g1333) & (!g1335) & (g1348) & (!g1351)) + ((g1323) & (!sk[96]) & (!g1333) & (!g1335) & (g1348) & (g1351)) + ((g1323) & (!sk[96]) & (!g1333) & (g1335) & (!g1348) & (!g1351)) + ((g1323) & (!sk[96]) & (!g1333) & (g1335) & (!g1348) & (g1351)) + ((g1323) & (!sk[96]) & (!g1333) & (g1335) & (g1348) & (!g1351)) + ((g1323) & (!sk[96]) & (!g1333) & (g1335) & (g1348) & (g1351)) + ((g1323) & (!sk[96]) & (g1333) & (!g1335) & (!g1348) & (!g1351)) + ((g1323) & (!sk[96]) & (g1333) & (!g1335) & (!g1348) & (g1351)) + ((g1323) & (!sk[96]) & (g1333) & (!g1335) & (g1348) & (!g1351)) + ((g1323) & (!sk[96]) & (g1333) & (!g1335) & (g1348) & (g1351)) + ((g1323) & (!sk[96]) & (g1333) & (g1335) & (!g1348) & (!g1351)) + ((g1323) & (!sk[96]) & (g1333) & (g1335) & (!g1348) & (g1351)) + ((g1323) & (!sk[96]) & (g1333) & (g1335) & (g1348) & (!g1351)) + ((g1323) & (!sk[96]) & (g1333) & (g1335) & (g1348) & (g1351)) + ((g1323) & (sk[96]) & (!g1333) & (!g1335) & (!g1348) & (!g1351)) + ((g1323) & (sk[96]) & (!g1333) & (!g1335) & (g1348) & (!g1351)) + ((g1323) & (sk[96]) & (!g1333) & (!g1335) & (g1348) & (g1351)) + ((g1323) & (sk[96]) & (!g1333) & (g1335) & (g1348) & (!g1351)) + ((g1323) & (sk[96]) & (g1333) & (!g1335) & (g1348) & (!g1351)) + ((g1323) & (sk[96]) & (g1333) & (g1335) & (g1348) & (!g1351)));
	assign g1367 = (((!sk[97]) & (!g1355) & (!g1352) & (!g1362) & (g1365) & (!g1366)) + ((!sk[97]) & (!g1355) & (!g1352) & (!g1362) & (g1365) & (g1366)) + ((!sk[97]) & (!g1355) & (!g1352) & (g1362) & (!g1365) & (!g1366)) + ((!sk[97]) & (!g1355) & (!g1352) & (g1362) & (!g1365) & (g1366)) + ((!sk[97]) & (!g1355) & (!g1352) & (g1362) & (g1365) & (!g1366)) + ((!sk[97]) & (!g1355) & (!g1352) & (g1362) & (g1365) & (g1366)) + ((!sk[97]) & (!g1355) & (g1352) & (!g1362) & (!g1365) & (!g1366)) + ((!sk[97]) & (!g1355) & (g1352) & (!g1362) & (!g1365) & (g1366)) + ((!sk[97]) & (!g1355) & (g1352) & (!g1362) & (g1365) & (!g1366)) + ((!sk[97]) & (!g1355) & (g1352) & (!g1362) & (g1365) & (g1366)) + ((!sk[97]) & (!g1355) & (g1352) & (g1362) & (!g1365) & (!g1366)) + ((!sk[97]) & (!g1355) & (g1352) & (g1362) & (!g1365) & (g1366)) + ((!sk[97]) & (!g1355) & (g1352) & (g1362) & (g1365) & (!g1366)) + ((!sk[97]) & (!g1355) & (g1352) & (g1362) & (g1365) & (g1366)) + ((!sk[97]) & (g1355) & (!g1352) & (!g1362) & (g1365) & (!g1366)) + ((!sk[97]) & (g1355) & (!g1352) & (!g1362) & (g1365) & (g1366)) + ((!sk[97]) & (g1355) & (!g1352) & (g1362) & (!g1365) & (!g1366)) + ((!sk[97]) & (g1355) & (!g1352) & (g1362) & (!g1365) & (g1366)) + ((!sk[97]) & (g1355) & (!g1352) & (g1362) & (g1365) & (!g1366)) + ((!sk[97]) & (g1355) & (!g1352) & (g1362) & (g1365) & (g1366)) + ((!sk[97]) & (g1355) & (g1352) & (!g1362) & (!g1365) & (!g1366)) + ((!sk[97]) & (g1355) & (g1352) & (!g1362) & (!g1365) & (g1366)) + ((!sk[97]) & (g1355) & (g1352) & (!g1362) & (g1365) & (!g1366)) + ((!sk[97]) & (g1355) & (g1352) & (!g1362) & (g1365) & (g1366)) + ((!sk[97]) & (g1355) & (g1352) & (g1362) & (!g1365) & (!g1366)) + ((!sk[97]) & (g1355) & (g1352) & (g1362) & (!g1365) & (g1366)) + ((!sk[97]) & (g1355) & (g1352) & (g1362) & (g1365) & (!g1366)) + ((!sk[97]) & (g1355) & (g1352) & (g1362) & (g1365) & (g1366)) + ((sk[97]) & (!g1355) & (!g1352) & (!g1362) & (!g1365) & (g1366)) + ((sk[97]) & (!g1355) & (!g1352) & (!g1362) & (g1365) & (!g1366)) + ((sk[97]) & (!g1355) & (!g1352) & (g1362) & (!g1365) & (!g1366)) + ((sk[97]) & (!g1355) & (!g1352) & (g1362) & (g1365) & (g1366)) + ((sk[97]) & (!g1355) & (g1352) & (!g1362) & (!g1365) & (g1366)) + ((sk[97]) & (!g1355) & (g1352) & (!g1362) & (g1365) & (!g1366)) + ((sk[97]) & (!g1355) & (g1352) & (g1362) & (!g1365) & (!g1366)) + ((sk[97]) & (!g1355) & (g1352) & (g1362) & (g1365) & (g1366)) + ((sk[97]) & (g1355) & (!g1352) & (!g1362) & (!g1365) & (g1366)) + ((sk[97]) & (g1355) & (!g1352) & (!g1362) & (g1365) & (!g1366)) + ((sk[97]) & (g1355) & (!g1352) & (g1362) & (!g1365) & (!g1366)) + ((sk[97]) & (g1355) & (!g1352) & (g1362) & (g1365) & (g1366)) + ((sk[97]) & (g1355) & (g1352) & (!g1362) & (!g1365) & (!g1366)) + ((sk[97]) & (g1355) & (g1352) & (!g1362) & (g1365) & (g1366)) + ((sk[97]) & (g1355) & (g1352) & (g1362) & (!g1365) & (g1366)) + ((sk[97]) & (g1355) & (g1352) & (g1362) & (g1365) & (!g1366)));
	assign sinx13x = (((!sk[98]) & (!g1068) & (g1354) & (!g1367)) + ((!sk[98]) & (!g1068) & (g1354) & (g1367)) + ((!sk[98]) & (g1068) & (g1354) & (!g1367)) + ((!sk[98]) & (g1068) & (g1354) & (g1367)) + ((sk[98]) & (!g1068) & (!g1354) & (g1367)) + ((sk[98]) & (!g1068) & (g1354) & (g1367)) + ((sk[98]) & (g1068) & (!g1354) & (!g1367)) + ((sk[98]) & (g1068) & (g1354) & (g1367)));
	assign g1369 = (((!g1355) & (!g1352) & (!g1362) & (!sk[99]) & (g1365) & (!g1366)) + ((!g1355) & (!g1352) & (!g1362) & (!sk[99]) & (g1365) & (g1366)) + ((!g1355) & (!g1352) & (g1362) & (!sk[99]) & (!g1365) & (!g1366)) + ((!g1355) & (!g1352) & (g1362) & (!sk[99]) & (!g1365) & (g1366)) + ((!g1355) & (!g1352) & (g1362) & (!sk[99]) & (g1365) & (!g1366)) + ((!g1355) & (!g1352) & (g1362) & (!sk[99]) & (g1365) & (g1366)) + ((!g1355) & (g1352) & (!g1362) & (!sk[99]) & (!g1365) & (!g1366)) + ((!g1355) & (g1352) & (!g1362) & (!sk[99]) & (!g1365) & (g1366)) + ((!g1355) & (g1352) & (!g1362) & (!sk[99]) & (g1365) & (!g1366)) + ((!g1355) & (g1352) & (!g1362) & (!sk[99]) & (g1365) & (g1366)) + ((!g1355) & (g1352) & (g1362) & (!sk[99]) & (!g1365) & (!g1366)) + ((!g1355) & (g1352) & (g1362) & (!sk[99]) & (!g1365) & (g1366)) + ((!g1355) & (g1352) & (g1362) & (!sk[99]) & (g1365) & (!g1366)) + ((!g1355) & (g1352) & (g1362) & (!sk[99]) & (g1365) & (g1366)) + ((g1355) & (!g1352) & (!g1362) & (!sk[99]) & (g1365) & (!g1366)) + ((g1355) & (!g1352) & (!g1362) & (!sk[99]) & (g1365) & (g1366)) + ((g1355) & (!g1352) & (g1362) & (!sk[99]) & (!g1365) & (!g1366)) + ((g1355) & (!g1352) & (g1362) & (!sk[99]) & (!g1365) & (g1366)) + ((g1355) & (!g1352) & (g1362) & (!sk[99]) & (g1365) & (!g1366)) + ((g1355) & (!g1352) & (g1362) & (!sk[99]) & (g1365) & (g1366)) + ((g1355) & (g1352) & (!g1362) & (!sk[99]) & (!g1365) & (!g1366)) + ((g1355) & (g1352) & (!g1362) & (!sk[99]) & (!g1365) & (g1366)) + ((g1355) & (g1352) & (!g1362) & (!sk[99]) & (g1365) & (!g1366)) + ((g1355) & (g1352) & (!g1362) & (!sk[99]) & (g1365) & (g1366)) + ((g1355) & (g1352) & (!g1362) & (sk[99]) & (!g1365) & (g1366)) + ((g1355) & (g1352) & (!g1362) & (sk[99]) & (g1365) & (!g1366)) + ((g1355) & (g1352) & (g1362) & (!sk[99]) & (!g1365) & (!g1366)) + ((g1355) & (g1352) & (g1362) & (!sk[99]) & (!g1365) & (g1366)) + ((g1355) & (g1352) & (g1362) & (!sk[99]) & (g1365) & (!g1366)) + ((g1355) & (g1352) & (g1362) & (!sk[99]) & (g1365) & (g1366)) + ((g1355) & (g1352) & (g1362) & (sk[99]) & (!g1365) & (!g1366)) + ((g1355) & (g1352) & (g1362) & (sk[99]) & (g1365) & (g1366)));
	assign g1370 = (((!g1340) & (!g1345) & (!g1346) & (!g1347) & (g1361) & (!g1365)) + ((!g1340) & (!g1345) & (!g1346) & (g1347) & (!g1361) & (!g1365)) + ((!g1340) & (!g1345) & (g1346) & (!g1347) & (!g1361) & (!g1365)) + ((!g1340) & (!g1345) & (g1346) & (g1347) & (!g1361) & (!g1365)) + ((!g1340) & (g1345) & (!g1346) & (!g1347) & (g1361) & (!g1365)) + ((!g1340) & (g1345) & (!g1346) & (g1347) & (g1361) & (!g1365)) + ((!g1340) & (g1345) & (g1346) & (!g1347) & (g1361) & (!g1365)) + ((!g1340) & (g1345) & (g1346) & (g1347) & (g1361) & (!g1365)) + ((g1340) & (!g1345) & (!g1346) & (!g1347) & (!g1361) & (!g1365)) + ((g1340) & (!g1345) & (!g1346) & (g1347) & (!g1361) & (!g1365)) + ((g1340) & (!g1345) & (g1346) & (!g1347) & (!g1361) & (!g1365)) + ((g1340) & (!g1345) & (g1346) & (g1347) & (!g1361) & (!g1365)) + ((g1340) & (g1345) & (!g1346) & (!g1347) & (g1361) & (!g1365)) + ((g1340) & (g1345) & (!g1346) & (g1347) & (!g1361) & (!g1365)) + ((g1340) & (g1345) & (g1346) & (!g1347) & (!g1361) & (!g1365)) + ((g1340) & (g1345) & (g1346) & (g1347) & (!g1361) & (!g1365)));
	assign g1371 = (((!g1340) & (!g1345) & (!g1346) & (!g1347) & (!g1361) & (g1365)) + ((!g1340) & (!g1345) & (!g1346) & (g1347) & (g1361) & (g1365)) + ((!g1340) & (!g1345) & (g1346) & (!g1347) & (g1361) & (g1365)) + ((!g1340) & (!g1345) & (g1346) & (g1347) & (g1361) & (g1365)) + ((!g1340) & (g1345) & (!g1346) & (!g1347) & (!g1361) & (g1365)) + ((!g1340) & (g1345) & (!g1346) & (g1347) & (!g1361) & (g1365)) + ((!g1340) & (g1345) & (g1346) & (!g1347) & (!g1361) & (g1365)) + ((!g1340) & (g1345) & (g1346) & (g1347) & (!g1361) & (g1365)) + ((g1340) & (!g1345) & (!g1346) & (!g1347) & (g1361) & (g1365)) + ((g1340) & (!g1345) & (!g1346) & (g1347) & (g1361) & (g1365)) + ((g1340) & (!g1345) & (g1346) & (!g1347) & (g1361) & (g1365)) + ((g1340) & (!g1345) & (g1346) & (g1347) & (g1361) & (g1365)) + ((g1340) & (g1345) & (!g1346) & (!g1347) & (!g1361) & (g1365)) + ((g1340) & (g1345) & (!g1346) & (g1347) & (g1361) & (g1365)) + ((g1340) & (g1345) & (g1346) & (!g1347) & (g1361) & (g1365)) + ((g1340) & (g1345) & (g1346) & (g1347) & (g1361) & (g1365)));
	assign g1372 = (((!g1323) & (!g1333) & (!g1335) & (!g1348) & (!g1351) & (!g1371)) + ((!g1323) & (!g1333) & (!g1335) & (g1348) & (!g1351) & (!g1371)) + ((!g1323) & (!g1333) & (!g1335) & (g1348) & (g1351) & (!g1371)) + ((!g1323) & (!g1333) & (g1335) & (!g1348) & (!g1351) & (!g1371)) + ((!g1323) & (!g1333) & (g1335) & (g1348) & (!g1351) & (!g1371)) + ((!g1323) & (!g1333) & (g1335) & (g1348) & (g1351) & (!g1371)) + ((!g1323) & (g1333) & (!g1335) & (!g1348) & (!g1351) & (!g1371)) + ((!g1323) & (g1333) & (!g1335) & (g1348) & (!g1351) & (!g1371)) + ((!g1323) & (g1333) & (!g1335) & (g1348) & (g1351) & (!g1371)) + ((!g1323) & (g1333) & (g1335) & (g1348) & (!g1351) & (!g1371)) + ((g1323) & (!g1333) & (!g1335) & (!g1348) & (!g1351) & (!g1371)) + ((g1323) & (!g1333) & (!g1335) & (g1348) & (!g1351) & (!g1371)) + ((g1323) & (!g1333) & (!g1335) & (g1348) & (g1351) & (!g1371)) + ((g1323) & (!g1333) & (g1335) & (g1348) & (!g1351) & (!g1371)) + ((g1323) & (g1333) & (!g1335) & (g1348) & (!g1351) & (!g1371)) + ((g1323) & (g1333) & (g1335) & (g1348) & (!g1351) & (!g1371)));
	assign g1373 = (((!g252) & (!g962) & (!g963) & (!g1344) & (!g1358) & (!g1359)) + ((!g252) & (!g962) & (!g963) & (!g1344) & (g1358) & (!g1359)) + ((!g252) & (!g962) & (!g963) & (!g1344) & (g1358) & (g1359)) + ((!g252) & (!g962) & (!g963) & (g1344) & (g1358) & (!g1359)) + ((!g252) & (!g962) & (g963) & (!g1344) & (!g1358) & (!g1359)) + ((!g252) & (!g962) & (g963) & (!g1344) & (g1358) & (!g1359)) + ((!g252) & (!g962) & (g963) & (!g1344) & (g1358) & (g1359)) + ((!g252) & (!g962) & (g963) & (g1344) & (g1358) & (!g1359)) + ((!g252) & (g962) & (!g963) & (!g1344) & (!g1358) & (!g1359)) + ((!g252) & (g962) & (!g963) & (!g1344) & (g1358) & (!g1359)) + ((!g252) & (g962) & (!g963) & (!g1344) & (g1358) & (g1359)) + ((!g252) & (g962) & (!g963) & (g1344) & (g1358) & (!g1359)) + ((!g252) & (g962) & (g963) & (!g1344) & (!g1358) & (!g1359)) + ((!g252) & (g962) & (g963) & (!g1344) & (g1358) & (!g1359)) + ((!g252) & (g962) & (g963) & (!g1344) & (g1358) & (g1359)) + ((!g252) & (g962) & (g963) & (g1344) & (g1358) & (!g1359)) + ((g252) & (!g962) & (!g963) & (!g1344) & (g1358) & (!g1359)) + ((g252) & (!g962) & (!g963) & (g1344) & (g1358) & (!g1359)) + ((g252) & (!g962) & (g963) & (!g1344) & (!g1358) & (!g1359)) + ((g252) & (!g962) & (g963) & (!g1344) & (g1358) & (!g1359)) + ((g252) & (!g962) & (g963) & (!g1344) & (g1358) & (g1359)) + ((g252) & (!g962) & (g963) & (g1344) & (g1358) & (!g1359)) + ((g252) & (g962) & (!g963) & (!g1344) & (!g1358) & (!g1359)) + ((g252) & (g962) & (!g963) & (!g1344) & (g1358) & (!g1359)) + ((g252) & (g962) & (!g963) & (!g1344) & (g1358) & (g1359)) + ((g252) & (g962) & (!g963) & (g1344) & (g1358) & (!g1359)) + ((g252) & (g962) & (g963) & (!g1344) & (!g1358) & (!g1359)) + ((g252) & (g962) & (g963) & (!g1344) & (g1358) & (!g1359)) + ((g252) & (g962) & (g963) & (!g1344) & (g1358) & (g1359)) + ((g252) & (g962) & (g963) & (g1344) & (!g1358) & (!g1359)) + ((g252) & (g962) & (g963) & (g1344) & (g1358) & (!g1359)) + ((g252) & (g962) & (g963) & (g1344) & (g1358) & (g1359)));
	assign g1374 = (((!g845) & (!g848) & (!sk[104]) & (!g1040) & (g1079)) + ((!g845) & (!g848) & (!sk[104]) & (g1040) & (g1079)) + ((!g845) & (g848) & (!sk[104]) & (!g1040) & (g1079)) + ((!g845) & (g848) & (!sk[104]) & (g1040) & (g1079)) + ((!g845) & (g848) & (sk[104]) & (!g1040) & (!g1079)) + ((!g845) & (g848) & (sk[104]) & (!g1040) & (g1079)) + ((g845) & (!g848) & (!sk[104]) & (!g1040) & (!g1079)) + ((g845) & (!g848) & (!sk[104]) & (!g1040) & (g1079)) + ((g845) & (!g848) & (!sk[104]) & (g1040) & (!g1079)) + ((g845) & (!g848) & (!sk[104]) & (g1040) & (g1079)) + ((g845) & (!g848) & (sk[104]) & (!g1040) & (!g1079)) + ((g845) & (!g848) & (sk[104]) & (g1040) & (!g1079)) + ((g845) & (g848) & (!sk[104]) & (!g1040) & (!g1079)) + ((g845) & (g848) & (!sk[104]) & (!g1040) & (g1079)) + ((g845) & (g848) & (!sk[104]) & (g1040) & (!g1079)) + ((g845) & (g848) & (!sk[104]) & (g1040) & (g1079)) + ((g845) & (g848) & (sk[104]) & (!g1040) & (!g1079)) + ((g845) & (g848) & (sk[104]) & (!g1040) & (g1079)) + ((g845) & (g848) & (sk[104]) & (g1040) & (!g1079)));
	assign g1375 = (((!g252) & (!sk[105]) & (!g843) & (!g1188) & (g1374)) + ((!g252) & (!sk[105]) & (!g843) & (g1188) & (g1374)) + ((!g252) & (!sk[105]) & (g843) & (!g1188) & (g1374)) + ((!g252) & (!sk[105]) & (g843) & (g1188) & (g1374)) + ((!g252) & (sk[105]) & (!g843) & (!g1188) & (!g1374)) + ((!g252) & (sk[105]) & (!g843) & (g1188) & (!g1374)) + ((!g252) & (sk[105]) & (g843) & (!g1188) & (!g1374)) + ((g252) & (!sk[105]) & (!g843) & (!g1188) & (!g1374)) + ((g252) & (!sk[105]) & (!g843) & (!g1188) & (g1374)) + ((g252) & (!sk[105]) & (!g843) & (g1188) & (!g1374)) + ((g252) & (!sk[105]) & (!g843) & (g1188) & (g1374)) + ((g252) & (!sk[105]) & (g843) & (!g1188) & (!g1374)) + ((g252) & (!sk[105]) & (g843) & (!g1188) & (g1374)) + ((g252) & (!sk[105]) & (g843) & (g1188) & (!g1374)) + ((g252) & (!sk[105]) & (g843) & (g1188) & (g1374)) + ((g252) & (sk[105]) & (!g843) & (!g1188) & (g1374)) + ((g252) & (sk[105]) & (!g843) & (g1188) & (g1374)) + ((g252) & (sk[105]) & (g843) & (!g1188) & (g1374)) + ((g252) & (sk[105]) & (g843) & (g1188) & (!g1374)) + ((g252) & (sk[105]) & (g843) & (g1188) & (g1374)));
	assign g1376 = (((!g202) & (!g252) & (!sk[106]) & (!g962) & (g971)) + ((!g202) & (!g252) & (!sk[106]) & (g962) & (g971)) + ((!g202) & (g252) & (!sk[106]) & (!g962) & (g971)) + ((!g202) & (g252) & (!sk[106]) & (g962) & (g971)) + ((!g202) & (g252) & (sk[106]) & (!g962) & (!g971)) + ((!g202) & (g252) & (sk[106]) & (!g962) & (g971)) + ((!g202) & (g252) & (sk[106]) & (g962) & (g971)) + ((g202) & (!g252) & (!sk[106]) & (!g962) & (!g971)) + ((g202) & (!g252) & (!sk[106]) & (!g962) & (g971)) + ((g202) & (!g252) & (!sk[106]) & (g962) & (!g971)) + ((g202) & (!g252) & (!sk[106]) & (g962) & (g971)) + ((g202) & (g252) & (!sk[106]) & (!g962) & (!g971)) + ((g202) & (g252) & (!sk[106]) & (!g962) & (g971)) + ((g202) & (g252) & (!sk[106]) & (g962) & (!g971)) + ((g202) & (g252) & (!sk[106]) & (g962) & (g971)) + ((g202) & (g252) & (sk[106]) & (!g962) & (g971)));
	assign g1377 = (((!g252) & (!sk[107]) & (!g994) & (!g1375) & (g1376)) + ((!g252) & (!sk[107]) & (!g994) & (g1375) & (g1376)) + ((!g252) & (!sk[107]) & (g994) & (!g1375) & (g1376)) + ((!g252) & (!sk[107]) & (g994) & (g1375) & (g1376)) + ((!g252) & (sk[107]) & (!g994) & (!g1375) & (!g1376)) + ((!g252) & (sk[107]) & (!g994) & (g1375) & (g1376)) + ((!g252) & (sk[107]) & (g994) & (!g1375) & (!g1376)) + ((!g252) & (sk[107]) & (g994) & (g1375) & (g1376)) + ((g252) & (!sk[107]) & (!g994) & (!g1375) & (!g1376)) + ((g252) & (!sk[107]) & (!g994) & (!g1375) & (g1376)) + ((g252) & (!sk[107]) & (!g994) & (g1375) & (!g1376)) + ((g252) & (!sk[107]) & (!g994) & (g1375) & (g1376)) + ((g252) & (!sk[107]) & (g994) & (!g1375) & (!g1376)) + ((g252) & (!sk[107]) & (g994) & (!g1375) & (g1376)) + ((g252) & (!sk[107]) & (g994) & (g1375) & (!g1376)) + ((g252) & (!sk[107]) & (g994) & (g1375) & (g1376)) + ((g252) & (sk[107]) & (!g994) & (!g1375) & (!g1376)) + ((g252) & (sk[107]) & (!g994) & (g1375) & (g1376)) + ((g252) & (sk[107]) & (g994) & (!g1375) & (g1376)) + ((g252) & (sk[107]) & (g994) & (g1375) & (!g1376)));
	assign g1378 = (((!g1340) & (!g1345) & (!g1346) & (!g1347) & (!g1356) & (!g1360)) + ((!g1340) & (!g1345) & (!g1346) & (!g1347) & (!g1356) & (g1360)) + ((!g1340) & (!g1345) & (!g1346) & (!g1347) & (g1356) & (!g1360)) + ((!g1340) & (!g1345) & (!g1346) & (g1347) & (!g1356) & (!g1360)) + ((!g1340) & (!g1345) & (g1346) & (!g1347) & (!g1356) & (!g1360)) + ((!g1340) & (!g1345) & (g1346) & (g1347) & (!g1356) & (!g1360)) + ((!g1340) & (g1345) & (!g1346) & (!g1347) & (!g1356) & (!g1360)) + ((!g1340) & (g1345) & (!g1346) & (!g1347) & (!g1356) & (g1360)) + ((!g1340) & (g1345) & (!g1346) & (!g1347) & (g1356) & (!g1360)) + ((!g1340) & (g1345) & (!g1346) & (g1347) & (!g1356) & (!g1360)) + ((!g1340) & (g1345) & (!g1346) & (g1347) & (!g1356) & (g1360)) + ((!g1340) & (g1345) & (!g1346) & (g1347) & (g1356) & (!g1360)) + ((!g1340) & (g1345) & (g1346) & (!g1347) & (!g1356) & (!g1360)) + ((!g1340) & (g1345) & (g1346) & (!g1347) & (!g1356) & (g1360)) + ((!g1340) & (g1345) & (g1346) & (!g1347) & (g1356) & (!g1360)) + ((!g1340) & (g1345) & (g1346) & (g1347) & (!g1356) & (!g1360)) + ((!g1340) & (g1345) & (g1346) & (g1347) & (!g1356) & (g1360)) + ((!g1340) & (g1345) & (g1346) & (g1347) & (g1356) & (!g1360)) + ((g1340) & (!g1345) & (!g1346) & (!g1347) & (!g1356) & (!g1360)) + ((g1340) & (!g1345) & (!g1346) & (g1347) & (!g1356) & (!g1360)) + ((g1340) & (!g1345) & (g1346) & (!g1347) & (!g1356) & (!g1360)) + ((g1340) & (!g1345) & (g1346) & (g1347) & (!g1356) & (!g1360)) + ((g1340) & (g1345) & (!g1346) & (!g1347) & (!g1356) & (!g1360)) + ((g1340) & (g1345) & (!g1346) & (!g1347) & (!g1356) & (g1360)) + ((g1340) & (g1345) & (!g1346) & (!g1347) & (g1356) & (!g1360)) + ((g1340) & (g1345) & (!g1346) & (g1347) & (!g1356) & (!g1360)) + ((g1340) & (g1345) & (g1346) & (!g1347) & (!g1356) & (!g1360)) + ((g1340) & (g1345) & (g1346) & (g1347) & (!g1356) & (!g1360)));
	assign g1379 = (((!g10) & (!g99) & (!sk[109]) & (!g33) & (g288)) + ((!g10) & (!g99) & (!sk[109]) & (g33) & (g288)) + ((!g10) & (!g99) & (sk[109]) & (!g33) & (!g288)) + ((!g10) & (g99) & (!sk[109]) & (!g33) & (g288)) + ((!g10) & (g99) & (!sk[109]) & (g33) & (g288)) + ((!g10) & (g99) & (sk[109]) & (!g33) & (!g288)) + ((g10) & (!g99) & (!sk[109]) & (!g33) & (!g288)) + ((g10) & (!g99) & (!sk[109]) & (!g33) & (g288)) + ((g10) & (!g99) & (!sk[109]) & (g33) & (!g288)) + ((g10) & (!g99) & (!sk[109]) & (g33) & (g288)) + ((g10) & (!g99) & (sk[109]) & (!g33) & (!g288)) + ((g10) & (g99) & (!sk[109]) & (!g33) & (!g288)) + ((g10) & (g99) & (!sk[109]) & (!g33) & (g288)) + ((g10) & (g99) & (!sk[109]) & (g33) & (!g288)) + ((g10) & (g99) & (!sk[109]) & (g33) & (g288)));
	assign g1380 = (((!sk[110]) & (!g79) & (!g260) & (!g618) & (g967) & (!g1379)) + ((!sk[110]) & (!g79) & (!g260) & (!g618) & (g967) & (g1379)) + ((!sk[110]) & (!g79) & (!g260) & (g618) & (!g967) & (!g1379)) + ((!sk[110]) & (!g79) & (!g260) & (g618) & (!g967) & (g1379)) + ((!sk[110]) & (!g79) & (!g260) & (g618) & (g967) & (!g1379)) + ((!sk[110]) & (!g79) & (!g260) & (g618) & (g967) & (g1379)) + ((!sk[110]) & (!g79) & (g260) & (!g618) & (!g967) & (!g1379)) + ((!sk[110]) & (!g79) & (g260) & (!g618) & (!g967) & (g1379)) + ((!sk[110]) & (!g79) & (g260) & (!g618) & (g967) & (!g1379)) + ((!sk[110]) & (!g79) & (g260) & (!g618) & (g967) & (g1379)) + ((!sk[110]) & (!g79) & (g260) & (g618) & (!g967) & (!g1379)) + ((!sk[110]) & (!g79) & (g260) & (g618) & (!g967) & (g1379)) + ((!sk[110]) & (!g79) & (g260) & (g618) & (g967) & (!g1379)) + ((!sk[110]) & (!g79) & (g260) & (g618) & (g967) & (g1379)) + ((!sk[110]) & (g79) & (!g260) & (!g618) & (g967) & (!g1379)) + ((!sk[110]) & (g79) & (!g260) & (!g618) & (g967) & (g1379)) + ((!sk[110]) & (g79) & (!g260) & (g618) & (!g967) & (!g1379)) + ((!sk[110]) & (g79) & (!g260) & (g618) & (!g967) & (g1379)) + ((!sk[110]) & (g79) & (!g260) & (g618) & (g967) & (!g1379)) + ((!sk[110]) & (g79) & (!g260) & (g618) & (g967) & (g1379)) + ((!sk[110]) & (g79) & (g260) & (!g618) & (!g967) & (!g1379)) + ((!sk[110]) & (g79) & (g260) & (!g618) & (!g967) & (g1379)) + ((!sk[110]) & (g79) & (g260) & (!g618) & (g967) & (!g1379)) + ((!sk[110]) & (g79) & (g260) & (!g618) & (g967) & (g1379)) + ((!sk[110]) & (g79) & (g260) & (g618) & (!g967) & (!g1379)) + ((!sk[110]) & (g79) & (g260) & (g618) & (!g967) & (g1379)) + ((!sk[110]) & (g79) & (g260) & (g618) & (g967) & (!g1379)) + ((!sk[110]) & (g79) & (g260) & (g618) & (g967) & (g1379)) + ((sk[110]) & (!g79) & (g260) & (g618) & (!g967) & (g1379)));
	assign g1381 = (((!g699) & (!g145) & (!g421) & (g654) & (!sk[111]) & (!g1380)) + ((!g699) & (!g145) & (!g421) & (g654) & (!sk[111]) & (g1380)) + ((!g699) & (!g145) & (g421) & (!g654) & (!sk[111]) & (!g1380)) + ((!g699) & (!g145) & (g421) & (!g654) & (!sk[111]) & (g1380)) + ((!g699) & (!g145) & (g421) & (g654) & (!sk[111]) & (!g1380)) + ((!g699) & (!g145) & (g421) & (g654) & (!sk[111]) & (g1380)) + ((!g699) & (g145) & (!g421) & (!g654) & (!sk[111]) & (!g1380)) + ((!g699) & (g145) & (!g421) & (!g654) & (!sk[111]) & (g1380)) + ((!g699) & (g145) & (!g421) & (g654) & (!sk[111]) & (!g1380)) + ((!g699) & (g145) & (!g421) & (g654) & (!sk[111]) & (g1380)) + ((!g699) & (g145) & (g421) & (!g654) & (!sk[111]) & (!g1380)) + ((!g699) & (g145) & (g421) & (!g654) & (!sk[111]) & (g1380)) + ((!g699) & (g145) & (g421) & (g654) & (!sk[111]) & (!g1380)) + ((!g699) & (g145) & (g421) & (g654) & (!sk[111]) & (g1380)) + ((g699) & (!g145) & (!g421) & (g654) & (!sk[111]) & (!g1380)) + ((g699) & (!g145) & (!g421) & (g654) & (!sk[111]) & (g1380)) + ((g699) & (!g145) & (g421) & (!g654) & (!sk[111]) & (!g1380)) + ((g699) & (!g145) & (g421) & (!g654) & (!sk[111]) & (g1380)) + ((g699) & (!g145) & (g421) & (g654) & (!sk[111]) & (!g1380)) + ((g699) & (!g145) & (g421) & (g654) & (!sk[111]) & (g1380)) + ((g699) & (g145) & (!g421) & (!g654) & (!sk[111]) & (!g1380)) + ((g699) & (g145) & (!g421) & (!g654) & (!sk[111]) & (g1380)) + ((g699) & (g145) & (!g421) & (g654) & (!sk[111]) & (!g1380)) + ((g699) & (g145) & (!g421) & (g654) & (!sk[111]) & (g1380)) + ((g699) & (g145) & (g421) & (!g654) & (!sk[111]) & (!g1380)) + ((g699) & (g145) & (g421) & (!g654) & (!sk[111]) & (g1380)) + ((g699) & (g145) & (g421) & (g654) & (!sk[111]) & (!g1380)) + ((g699) & (g145) & (g421) & (g654) & (!sk[111]) & (g1380)) + ((g699) & (g145) & (g421) & (g654) & (sk[111]) & (g1380)));
	assign g1382 = (((!g1373) & (!g1377) & (!sk[112]) & (!g1378) & (g1381)) + ((!g1373) & (!g1377) & (!sk[112]) & (g1378) & (g1381)) + ((!g1373) & (!g1377) & (sk[112]) & (!g1378) & (!g1381)) + ((!g1373) & (!g1377) & (sk[112]) & (g1378) & (g1381)) + ((!g1373) & (g1377) & (!sk[112]) & (!g1378) & (g1381)) + ((!g1373) & (g1377) & (!sk[112]) & (g1378) & (g1381)) + ((!g1373) & (g1377) & (sk[112]) & (!g1378) & (g1381)) + ((!g1373) & (g1377) & (sk[112]) & (g1378) & (!g1381)) + ((g1373) & (!g1377) & (!sk[112]) & (!g1378) & (!g1381)) + ((g1373) & (!g1377) & (!sk[112]) & (!g1378) & (g1381)) + ((g1373) & (!g1377) & (!sk[112]) & (g1378) & (!g1381)) + ((g1373) & (!g1377) & (!sk[112]) & (g1378) & (g1381)) + ((g1373) & (!g1377) & (sk[112]) & (!g1378) & (g1381)) + ((g1373) & (!g1377) & (sk[112]) & (g1378) & (!g1381)) + ((g1373) & (g1377) & (!sk[112]) & (!g1378) & (!g1381)) + ((g1373) & (g1377) & (!sk[112]) & (!g1378) & (g1381)) + ((g1373) & (g1377) & (!sk[112]) & (g1378) & (!g1381)) + ((g1373) & (g1377) & (!sk[112]) & (g1378) & (g1381)) + ((g1373) & (g1377) & (sk[112]) & (!g1378) & (!g1381)) + ((g1373) & (g1377) & (sk[112]) & (g1378) & (g1381)));
	assign g1383 = (((!g1370) & (!sk[113]) & (g1372) & (!g1382)) + ((!g1370) & (!sk[113]) & (g1372) & (g1382)) + ((!g1370) & (sk[113]) & (!g1372) & (g1382)) + ((!g1370) & (sk[113]) & (g1372) & (!g1382)) + ((g1370) & (!sk[113]) & (g1372) & (!g1382)) + ((g1370) & (!sk[113]) & (g1372) & (g1382)) + ((g1370) & (sk[113]) & (!g1372) & (!g1382)) + ((g1370) & (sk[113]) & (g1372) & (!g1382)));
	assign sinx14x = (((!sk[114]) & (!g1068) & (!g1354) & (!g1367) & (g1369) & (!g1383)) + ((!sk[114]) & (!g1068) & (!g1354) & (!g1367) & (g1369) & (g1383)) + ((!sk[114]) & (!g1068) & (!g1354) & (g1367) & (!g1369) & (!g1383)) + ((!sk[114]) & (!g1068) & (!g1354) & (g1367) & (!g1369) & (g1383)) + ((!sk[114]) & (!g1068) & (!g1354) & (g1367) & (g1369) & (!g1383)) + ((!sk[114]) & (!g1068) & (!g1354) & (g1367) & (g1369) & (g1383)) + ((!sk[114]) & (!g1068) & (g1354) & (!g1367) & (!g1369) & (!g1383)) + ((!sk[114]) & (!g1068) & (g1354) & (!g1367) & (!g1369) & (g1383)) + ((!sk[114]) & (!g1068) & (g1354) & (!g1367) & (g1369) & (!g1383)) + ((!sk[114]) & (!g1068) & (g1354) & (!g1367) & (g1369) & (g1383)) + ((!sk[114]) & (!g1068) & (g1354) & (g1367) & (!g1369) & (!g1383)) + ((!sk[114]) & (!g1068) & (g1354) & (g1367) & (!g1369) & (g1383)) + ((!sk[114]) & (!g1068) & (g1354) & (g1367) & (g1369) & (!g1383)) + ((!sk[114]) & (!g1068) & (g1354) & (g1367) & (g1369) & (g1383)) + ((!sk[114]) & (g1068) & (!g1354) & (!g1367) & (g1369) & (!g1383)) + ((!sk[114]) & (g1068) & (!g1354) & (!g1367) & (g1369) & (g1383)) + ((!sk[114]) & (g1068) & (!g1354) & (g1367) & (!g1369) & (!g1383)) + ((!sk[114]) & (g1068) & (!g1354) & (g1367) & (!g1369) & (g1383)) + ((!sk[114]) & (g1068) & (!g1354) & (g1367) & (g1369) & (!g1383)) + ((!sk[114]) & (g1068) & (!g1354) & (g1367) & (g1369) & (g1383)) + ((!sk[114]) & (g1068) & (g1354) & (!g1367) & (!g1369) & (!g1383)) + ((!sk[114]) & (g1068) & (g1354) & (!g1367) & (!g1369) & (g1383)) + ((!sk[114]) & (g1068) & (g1354) & (!g1367) & (g1369) & (!g1383)) + ((!sk[114]) & (g1068) & (g1354) & (!g1367) & (g1369) & (g1383)) + ((!sk[114]) & (g1068) & (g1354) & (g1367) & (!g1369) & (!g1383)) + ((!sk[114]) & (g1068) & (g1354) & (g1367) & (!g1369) & (g1383)) + ((!sk[114]) & (g1068) & (g1354) & (g1367) & (g1369) & (!g1383)) + ((!sk[114]) & (g1068) & (g1354) & (g1367) & (g1369) & (g1383)) + ((sk[114]) & (!g1068) & (!g1354) & (!g1367) & (!g1369) & (g1383)) + ((sk[114]) & (!g1068) & (!g1354) & (!g1367) & (g1369) & (!g1383)) + ((sk[114]) & (!g1068) & (!g1354) & (g1367) & (!g1369) & (g1383)) + ((sk[114]) & (!g1068) & (!g1354) & (g1367) & (g1369) & (!g1383)) + ((sk[114]) & (!g1068) & (g1354) & (!g1367) & (!g1369) & (g1383)) + ((sk[114]) & (!g1068) & (g1354) & (!g1367) & (g1369) & (!g1383)) + ((sk[114]) & (!g1068) & (g1354) & (g1367) & (!g1369) & (g1383)) + ((sk[114]) & (!g1068) & (g1354) & (g1367) & (g1369) & (!g1383)) + ((sk[114]) & (g1068) & (!g1354) & (!g1367) & (!g1369) & (!g1383)) + ((sk[114]) & (g1068) & (!g1354) & (!g1367) & (g1369) & (g1383)) + ((sk[114]) & (g1068) & (!g1354) & (g1367) & (!g1369) & (!g1383)) + ((sk[114]) & (g1068) & (!g1354) & (g1367) & (g1369) & (g1383)) + ((sk[114]) & (g1068) & (g1354) & (!g1367) & (!g1369) & (g1383)) + ((sk[114]) & (g1068) & (g1354) & (!g1367) & (g1369) & (!g1383)) + ((sk[114]) & (g1068) & (g1354) & (g1367) & (!g1369) & (!g1383)) + ((sk[114]) & (g1068) & (g1354) & (g1367) & (g1369) & (g1383)));
	assign g1385 = (((!g1373) & (!sk[115]) & (g1377) & (!g1378)) + ((!g1373) & (!sk[115]) & (g1377) & (g1378)) + ((!g1373) & (sk[115]) & (!g1377) & (g1378)) + ((!g1373) & (sk[115]) & (g1377) & (!g1378)) + ((g1373) & (!sk[115]) & (g1377) & (!g1378)) + ((g1373) & (!sk[115]) & (g1377) & (g1378)) + ((g1373) & (sk[115]) & (!g1377) & (!g1378)) + ((g1373) & (sk[115]) & (g1377) & (g1378)));
	assign g1386 = (((!sk[116]) & (!g252) & (!g994) & (!g1375) & (g1376)) + ((!sk[116]) & (!g252) & (!g994) & (g1375) & (g1376)) + ((!sk[116]) & (!g252) & (g994) & (!g1375) & (g1376)) + ((!sk[116]) & (!g252) & (g994) & (g1375) & (g1376)) + ((!sk[116]) & (g252) & (!g994) & (!g1375) & (!g1376)) + ((!sk[116]) & (g252) & (!g994) & (!g1375) & (g1376)) + ((!sk[116]) & (g252) & (!g994) & (g1375) & (!g1376)) + ((!sk[116]) & (g252) & (!g994) & (g1375) & (g1376)) + ((!sk[116]) & (g252) & (g994) & (!g1375) & (!g1376)) + ((!sk[116]) & (g252) & (g994) & (!g1375) & (g1376)) + ((!sk[116]) & (g252) & (g994) & (g1375) & (!g1376)) + ((!sk[116]) & (g252) & (g994) & (g1375) & (g1376)) + ((sk[116]) & (!g252) & (!g994) & (g1375) & (!g1376)) + ((sk[116]) & (!g252) & (g994) & (g1375) & (!g1376)) + ((sk[116]) & (g252) & (!g994) & (g1375) & (!g1376)) + ((sk[116]) & (g252) & (g994) & (!g1375) & (!g1376)) + ((sk[116]) & (g252) & (g994) & (g1375) & (!g1376)) + ((sk[116]) & (g252) & (g994) & (g1375) & (g1376)));
	assign g1387 = (((!g252) & (!g843) & (g848) & (!g1040) & (!g1079) & (!g1080)) + ((!g252) & (!g843) & (g848) & (!g1040) & (!g1079) & (g1080)) + ((!g252) & (!g843) & (g848) & (g1040) & (!g1079) & (!g1080)) + ((!g252) & (!g843) & (g848) & (g1040) & (!g1079) & (g1080)) + ((!g252) & (g843) & (!g848) & (!g1040) & (!g1079) & (!g1080)) + ((!g252) & (g843) & (!g848) & (!g1040) & (!g1079) & (g1080)) + ((!g252) & (g843) & (!g848) & (g1040) & (!g1079) & (g1080)) + ((!g252) & (g843) & (g848) & (!g1040) & (!g1079) & (!g1080)) + ((!g252) & (g843) & (g848) & (!g1040) & (!g1079) & (g1080)) + ((!g252) & (g843) & (g848) & (g1040) & (!g1079) & (!g1080)) + ((!g252) & (g843) & (g848) & (g1040) & (!g1079) & (g1080)) + ((g252) & (!g843) & (!g848) & (!g1040) & (!g1079) & (!g1080)) + ((g252) & (!g843) & (!g848) & (!g1040) & (!g1079) & (g1080)) + ((g252) & (!g843) & (!g848) & (!g1040) & (g1079) & (!g1080)) + ((g252) & (!g843) & (!g848) & (!g1040) & (g1079) & (g1080)) + ((g252) & (!g843) & (!g848) & (g1040) & (!g1079) & (!g1080)) + ((g252) & (!g843) & (!g848) & (g1040) & (!g1079) & (g1080)) + ((g252) & (!g843) & (!g848) & (g1040) & (g1079) & (!g1080)) + ((g252) & (!g843) & (!g848) & (g1040) & (g1079) & (g1080)) + ((g252) & (!g843) & (g848) & (!g1040) & (g1079) & (!g1080)) + ((g252) & (!g843) & (g848) & (!g1040) & (g1079) & (g1080)) + ((g252) & (!g843) & (g848) & (g1040) & (g1079) & (!g1080)) + ((g252) & (!g843) & (g848) & (g1040) & (g1079) & (g1080)) + ((g252) & (g843) & (!g848) & (!g1040) & (g1079) & (!g1080)) + ((g252) & (g843) & (!g848) & (!g1040) & (g1079) & (g1080)) + ((g252) & (g843) & (!g848) & (g1040) & (!g1079) & (!g1080)) + ((g252) & (g843) & (!g848) & (g1040) & (g1079) & (!g1080)) + ((g252) & (g843) & (!g848) & (g1040) & (g1079) & (g1080)) + ((g252) & (g843) & (g848) & (!g1040) & (g1079) & (!g1080)) + ((g252) & (g843) & (g848) & (!g1040) & (g1079) & (g1080)) + ((g252) & (g843) & (g848) & (g1040) & (g1079) & (!g1080)) + ((g252) & (g843) & (g848) & (g1040) & (g1079) & (g1080)));
	assign g1388 = (((!g252) & (!g994) & (!g1040) & (!sk[118]) & (g1387)) + ((!g252) & (!g994) & (!g1040) & (sk[118]) & (!g1387)) + ((!g252) & (!g994) & (g1040) & (!sk[118]) & (g1387)) + ((!g252) & (!g994) & (g1040) & (sk[118]) & (!g1387)) + ((!g252) & (g994) & (!g1040) & (!sk[118]) & (g1387)) + ((!g252) & (g994) & (!g1040) & (sk[118]) & (!g1387)) + ((!g252) & (g994) & (g1040) & (!sk[118]) & (g1387)) + ((!g252) & (g994) & (g1040) & (sk[118]) & (!g1387)) + ((g252) & (!g994) & (!g1040) & (!sk[118]) & (!g1387)) + ((g252) & (!g994) & (!g1040) & (!sk[118]) & (g1387)) + ((g252) & (!g994) & (!g1040) & (sk[118]) & (g1387)) + ((g252) & (!g994) & (g1040) & (!sk[118]) & (!g1387)) + ((g252) & (!g994) & (g1040) & (!sk[118]) & (g1387)) + ((g252) & (!g994) & (g1040) & (sk[118]) & (!g1387)) + ((g252) & (g994) & (!g1040) & (!sk[118]) & (!g1387)) + ((g252) & (g994) & (!g1040) & (!sk[118]) & (g1387)) + ((g252) & (g994) & (!g1040) & (sk[118]) & (!g1387)) + ((g252) & (g994) & (g1040) & (!sk[118]) & (!g1387)) + ((g252) & (g994) & (g1040) & (!sk[118]) & (g1387)) + ((g252) & (g994) & (g1040) & (sk[118]) & (g1387)));
	assign g1389 = (((!g1373) & (!g1377) & (!g1378) & (!g1386) & (sk[119]) & (!g1388)) + ((!g1373) & (!g1377) & (!g1378) & (g1386) & (!sk[119]) & (!g1388)) + ((!g1373) & (!g1377) & (!g1378) & (g1386) & (!sk[119]) & (g1388)) + ((!g1373) & (!g1377) & (!g1378) & (g1386) & (sk[119]) & (g1388)) + ((!g1373) & (!g1377) & (g1378) & (!g1386) & (!sk[119]) & (!g1388)) + ((!g1373) & (!g1377) & (g1378) & (!g1386) & (!sk[119]) & (g1388)) + ((!g1373) & (!g1377) & (g1378) & (!g1386) & (sk[119]) & (g1388)) + ((!g1373) & (!g1377) & (g1378) & (g1386) & (!sk[119]) & (!g1388)) + ((!g1373) & (!g1377) & (g1378) & (g1386) & (!sk[119]) & (g1388)) + ((!g1373) & (!g1377) & (g1378) & (g1386) & (sk[119]) & (!g1388)) + ((!g1373) & (g1377) & (!g1378) & (!g1386) & (!sk[119]) & (!g1388)) + ((!g1373) & (g1377) & (!g1378) & (!g1386) & (!sk[119]) & (g1388)) + ((!g1373) & (g1377) & (!g1378) & (!g1386) & (sk[119]) & (g1388)) + ((!g1373) & (g1377) & (!g1378) & (g1386) & (!sk[119]) & (!g1388)) + ((!g1373) & (g1377) & (!g1378) & (g1386) & (!sk[119]) & (g1388)) + ((!g1373) & (g1377) & (!g1378) & (g1386) & (sk[119]) & (!g1388)) + ((!g1373) & (g1377) & (g1378) & (!g1386) & (!sk[119]) & (!g1388)) + ((!g1373) & (g1377) & (g1378) & (!g1386) & (!sk[119]) & (g1388)) + ((!g1373) & (g1377) & (g1378) & (!g1386) & (sk[119]) & (g1388)) + ((!g1373) & (g1377) & (g1378) & (g1386) & (!sk[119]) & (!g1388)) + ((!g1373) & (g1377) & (g1378) & (g1386) & (!sk[119]) & (g1388)) + ((!g1373) & (g1377) & (g1378) & (g1386) & (sk[119]) & (!g1388)) + ((g1373) & (!g1377) & (!g1378) & (!g1386) & (sk[119]) & (!g1388)) + ((g1373) & (!g1377) & (!g1378) & (g1386) & (!sk[119]) & (!g1388)) + ((g1373) & (!g1377) & (!g1378) & (g1386) & (!sk[119]) & (g1388)) + ((g1373) & (!g1377) & (!g1378) & (g1386) & (sk[119]) & (g1388)) + ((g1373) & (!g1377) & (g1378) & (!g1386) & (!sk[119]) & (!g1388)) + ((g1373) & (!g1377) & (g1378) & (!g1386) & (!sk[119]) & (g1388)) + ((g1373) & (!g1377) & (g1378) & (!g1386) & (sk[119]) & (!g1388)) + ((g1373) & (!g1377) & (g1378) & (g1386) & (!sk[119]) & (!g1388)) + ((g1373) & (!g1377) & (g1378) & (g1386) & (!sk[119]) & (g1388)) + ((g1373) & (!g1377) & (g1378) & (g1386) & (sk[119]) & (g1388)) + ((g1373) & (g1377) & (!g1378) & (!g1386) & (!sk[119]) & (!g1388)) + ((g1373) & (g1377) & (!g1378) & (!g1386) & (!sk[119]) & (g1388)) + ((g1373) & (g1377) & (!g1378) & (!g1386) & (sk[119]) & (!g1388)) + ((g1373) & (g1377) & (!g1378) & (g1386) & (!sk[119]) & (!g1388)) + ((g1373) & (g1377) & (!g1378) & (g1386) & (!sk[119]) & (g1388)) + ((g1373) & (g1377) & (!g1378) & (g1386) & (sk[119]) & (g1388)) + ((g1373) & (g1377) & (g1378) & (!g1386) & (!sk[119]) & (!g1388)) + ((g1373) & (g1377) & (g1378) & (!g1386) & (!sk[119]) & (g1388)) + ((g1373) & (g1377) & (g1378) & (!g1386) & (sk[119]) & (g1388)) + ((g1373) & (g1377) & (g1378) & (g1386) & (!sk[119]) & (!g1388)) + ((g1373) & (g1377) & (g1378) & (g1386) & (!sk[119]) & (g1388)) + ((g1373) & (g1377) & (g1378) & (g1386) & (sk[119]) & (!g1388)));
	assign g1390 = (((!g9) & (!g46) & (!g41) & (!g66) & (!g20) & (g357)) + ((!g9) & (!g46) & (!g41) & (!g66) & (g20) & (g357)) + ((!g9) & (!g46) & (!g41) & (g66) & (!g20) & (g357)) + ((!g9) & (!g46) & (!g41) & (g66) & (g20) & (g357)) + ((!g9) & (!g46) & (g41) & (!g66) & (!g20) & (g357)) + ((!g9) & (!g46) & (g41) & (!g66) & (g20) & (g357)) + ((!g9) & (!g46) & (g41) & (g66) & (!g20) & (g357)) + ((!g9) & (!g46) & (g41) & (g66) & (g20) & (g357)) + ((!g9) & (g46) & (!g41) & (!g66) & (!g20) & (g357)) + ((!g9) & (g46) & (!g41) & (!g66) & (g20) & (g357)) + ((!g9) & (g46) & (!g41) & (g66) & (!g20) & (g357)) + ((!g9) & (g46) & (!g41) & (g66) & (g20) & (g357)) + ((g9) & (!g46) & (!g41) & (!g66) & (!g20) & (g357)) + ((g9) & (!g46) & (g41) & (!g66) & (!g20) & (g357)) + ((g9) & (g46) & (!g41) & (!g66) & (!g20) & (g357)));
	assign g1391 = (((!g49) & (!g62) & (!g101) & (!sk[121]) & (g1177)) + ((!g49) & (!g62) & (!g101) & (sk[121]) & (!g1177)) + ((!g49) & (!g62) & (g101) & (!sk[121]) & (g1177)) + ((!g49) & (g62) & (!g101) & (!sk[121]) & (g1177)) + ((!g49) & (g62) & (!g101) & (sk[121]) & (!g1177)) + ((!g49) & (g62) & (g101) & (!sk[121]) & (g1177)) + ((g49) & (!g62) & (!g101) & (!sk[121]) & (!g1177)) + ((g49) & (!g62) & (!g101) & (!sk[121]) & (g1177)) + ((g49) & (!g62) & (!g101) & (sk[121]) & (!g1177)) + ((g49) & (!g62) & (g101) & (!sk[121]) & (!g1177)) + ((g49) & (!g62) & (g101) & (!sk[121]) & (g1177)) + ((g49) & (g62) & (!g101) & (!sk[121]) & (!g1177)) + ((g49) & (g62) & (!g101) & (!sk[121]) & (g1177)) + ((g49) & (g62) & (g101) & (!sk[121]) & (!g1177)) + ((g49) & (g62) & (g101) & (!sk[121]) & (g1177)));
	assign g1392 = (((!sk[122]) & (!g99) & (!g40) & (!g636) & (g1379) & (!g1391)) + ((!sk[122]) & (!g99) & (!g40) & (!g636) & (g1379) & (g1391)) + ((!sk[122]) & (!g99) & (!g40) & (g636) & (!g1379) & (!g1391)) + ((!sk[122]) & (!g99) & (!g40) & (g636) & (!g1379) & (g1391)) + ((!sk[122]) & (!g99) & (!g40) & (g636) & (g1379) & (!g1391)) + ((!sk[122]) & (!g99) & (!g40) & (g636) & (g1379) & (g1391)) + ((!sk[122]) & (!g99) & (g40) & (!g636) & (!g1379) & (!g1391)) + ((!sk[122]) & (!g99) & (g40) & (!g636) & (!g1379) & (g1391)) + ((!sk[122]) & (!g99) & (g40) & (!g636) & (g1379) & (!g1391)) + ((!sk[122]) & (!g99) & (g40) & (!g636) & (g1379) & (g1391)) + ((!sk[122]) & (!g99) & (g40) & (g636) & (!g1379) & (!g1391)) + ((!sk[122]) & (!g99) & (g40) & (g636) & (!g1379) & (g1391)) + ((!sk[122]) & (!g99) & (g40) & (g636) & (g1379) & (!g1391)) + ((!sk[122]) & (!g99) & (g40) & (g636) & (g1379) & (g1391)) + ((!sk[122]) & (g99) & (!g40) & (!g636) & (g1379) & (!g1391)) + ((!sk[122]) & (g99) & (!g40) & (!g636) & (g1379) & (g1391)) + ((!sk[122]) & (g99) & (!g40) & (g636) & (!g1379) & (!g1391)) + ((!sk[122]) & (g99) & (!g40) & (g636) & (!g1379) & (g1391)) + ((!sk[122]) & (g99) & (!g40) & (g636) & (g1379) & (!g1391)) + ((!sk[122]) & (g99) & (!g40) & (g636) & (g1379) & (g1391)) + ((!sk[122]) & (g99) & (g40) & (!g636) & (!g1379) & (!g1391)) + ((!sk[122]) & (g99) & (g40) & (!g636) & (!g1379) & (g1391)) + ((!sk[122]) & (g99) & (g40) & (!g636) & (g1379) & (!g1391)) + ((!sk[122]) & (g99) & (g40) & (!g636) & (g1379) & (g1391)) + ((!sk[122]) & (g99) & (g40) & (g636) & (!g1379) & (!g1391)) + ((!sk[122]) & (g99) & (g40) & (g636) & (!g1379) & (g1391)) + ((!sk[122]) & (g99) & (g40) & (g636) & (g1379) & (!g1391)) + ((!sk[122]) & (g99) & (g40) & (g636) & (g1379) & (g1391)) + ((sk[122]) & (!g99) & (!g40) & (g636) & (g1379) & (g1391)) + ((sk[122]) & (!g99) & (g40) & (g636) & (g1379) & (g1391)) + ((sk[122]) & (g99) & (!g40) & (g636) & (g1379) & (g1391)));
	assign g1393 = (((!sk[123]) & (!g333) & (!g620) & (!g1349) & (g1390) & (!g1392)) + ((!sk[123]) & (!g333) & (!g620) & (!g1349) & (g1390) & (g1392)) + ((!sk[123]) & (!g333) & (!g620) & (g1349) & (!g1390) & (!g1392)) + ((!sk[123]) & (!g333) & (!g620) & (g1349) & (!g1390) & (g1392)) + ((!sk[123]) & (!g333) & (!g620) & (g1349) & (g1390) & (!g1392)) + ((!sk[123]) & (!g333) & (!g620) & (g1349) & (g1390) & (g1392)) + ((!sk[123]) & (!g333) & (g620) & (!g1349) & (!g1390) & (!g1392)) + ((!sk[123]) & (!g333) & (g620) & (!g1349) & (!g1390) & (g1392)) + ((!sk[123]) & (!g333) & (g620) & (!g1349) & (g1390) & (!g1392)) + ((!sk[123]) & (!g333) & (g620) & (!g1349) & (g1390) & (g1392)) + ((!sk[123]) & (!g333) & (g620) & (g1349) & (!g1390) & (!g1392)) + ((!sk[123]) & (!g333) & (g620) & (g1349) & (!g1390) & (g1392)) + ((!sk[123]) & (!g333) & (g620) & (g1349) & (g1390) & (!g1392)) + ((!sk[123]) & (!g333) & (g620) & (g1349) & (g1390) & (g1392)) + ((!sk[123]) & (g333) & (!g620) & (!g1349) & (g1390) & (!g1392)) + ((!sk[123]) & (g333) & (!g620) & (!g1349) & (g1390) & (g1392)) + ((!sk[123]) & (g333) & (!g620) & (g1349) & (!g1390) & (!g1392)) + ((!sk[123]) & (g333) & (!g620) & (g1349) & (!g1390) & (g1392)) + ((!sk[123]) & (g333) & (!g620) & (g1349) & (g1390) & (!g1392)) + ((!sk[123]) & (g333) & (!g620) & (g1349) & (g1390) & (g1392)) + ((!sk[123]) & (g333) & (g620) & (!g1349) & (!g1390) & (!g1392)) + ((!sk[123]) & (g333) & (g620) & (!g1349) & (!g1390) & (g1392)) + ((!sk[123]) & (g333) & (g620) & (!g1349) & (g1390) & (!g1392)) + ((!sk[123]) & (g333) & (g620) & (!g1349) & (g1390) & (g1392)) + ((!sk[123]) & (g333) & (g620) & (g1349) & (!g1390) & (!g1392)) + ((!sk[123]) & (g333) & (g620) & (g1349) & (!g1390) & (g1392)) + ((!sk[123]) & (g333) & (g620) & (g1349) & (g1390) & (!g1392)) + ((!sk[123]) & (g333) & (g620) & (g1349) & (g1390) & (g1392)) + ((sk[123]) & (g333) & (g620) & (g1349) & (g1390) & (g1392)));
	assign g1394 = (((!g1370) & (!g1372) & (!g1385) & (!g1381) & (!g1389) & (g1393)) + ((!g1370) & (!g1372) & (!g1385) & (!g1381) & (g1389) & (!g1393)) + ((!g1370) & (!g1372) & (!g1385) & (g1381) & (!g1389) & (g1393)) + ((!g1370) & (!g1372) & (!g1385) & (g1381) & (g1389) & (!g1393)) + ((!g1370) & (!g1372) & (g1385) & (!g1381) & (!g1389) & (!g1393)) + ((!g1370) & (!g1372) & (g1385) & (!g1381) & (g1389) & (g1393)) + ((!g1370) & (!g1372) & (g1385) & (g1381) & (!g1389) & (g1393)) + ((!g1370) & (!g1372) & (g1385) & (g1381) & (g1389) & (!g1393)) + ((!g1370) & (g1372) & (!g1385) & (!g1381) & (!g1389) & (!g1393)) + ((!g1370) & (g1372) & (!g1385) & (!g1381) & (g1389) & (g1393)) + ((!g1370) & (g1372) & (!g1385) & (g1381) & (!g1389) & (g1393)) + ((!g1370) & (g1372) & (!g1385) & (g1381) & (g1389) & (!g1393)) + ((!g1370) & (g1372) & (g1385) & (!g1381) & (!g1389) & (!g1393)) + ((!g1370) & (g1372) & (g1385) & (!g1381) & (g1389) & (g1393)) + ((!g1370) & (g1372) & (g1385) & (g1381) & (!g1389) & (!g1393)) + ((!g1370) & (g1372) & (g1385) & (g1381) & (g1389) & (g1393)) + ((g1370) & (!g1372) & (!g1385) & (!g1381) & (!g1389) & (!g1393)) + ((g1370) & (!g1372) & (!g1385) & (!g1381) & (g1389) & (g1393)) + ((g1370) & (!g1372) & (!g1385) & (g1381) & (!g1389) & (g1393)) + ((g1370) & (!g1372) & (!g1385) & (g1381) & (g1389) & (!g1393)) + ((g1370) & (!g1372) & (g1385) & (!g1381) & (!g1389) & (!g1393)) + ((g1370) & (!g1372) & (g1385) & (!g1381) & (g1389) & (g1393)) + ((g1370) & (!g1372) & (g1385) & (g1381) & (!g1389) & (!g1393)) + ((g1370) & (!g1372) & (g1385) & (g1381) & (g1389) & (g1393)) + ((g1370) & (g1372) & (!g1385) & (!g1381) & (!g1389) & (!g1393)) + ((g1370) & (g1372) & (!g1385) & (!g1381) & (g1389) & (g1393)) + ((g1370) & (g1372) & (!g1385) & (g1381) & (!g1389) & (g1393)) + ((g1370) & (g1372) & (!g1385) & (g1381) & (g1389) & (!g1393)) + ((g1370) & (g1372) & (g1385) & (!g1381) & (!g1389) & (!g1393)) + ((g1370) & (g1372) & (g1385) & (!g1381) & (g1389) & (g1393)) + ((g1370) & (g1372) & (g1385) & (g1381) & (!g1389) & (!g1393)) + ((g1370) & (g1372) & (g1385) & (g1381) & (g1389) & (g1393)));
	assign sinx15x = (((!g1068) & (!g1354) & (!g1367) & (!g1369) & (!g1383) & (g1394)) + ((!g1068) & (!g1354) & (!g1367) & (!g1369) & (g1383) & (g1394)) + ((!g1068) & (!g1354) & (!g1367) & (g1369) & (!g1383) & (g1394)) + ((!g1068) & (!g1354) & (!g1367) & (g1369) & (g1383) & (!g1394)) + ((!g1068) & (!g1354) & (g1367) & (!g1369) & (!g1383) & (g1394)) + ((!g1068) & (!g1354) & (g1367) & (!g1369) & (g1383) & (g1394)) + ((!g1068) & (!g1354) & (g1367) & (g1369) & (!g1383) & (g1394)) + ((!g1068) & (!g1354) & (g1367) & (g1369) & (g1383) & (!g1394)) + ((!g1068) & (g1354) & (!g1367) & (!g1369) & (!g1383) & (g1394)) + ((!g1068) & (g1354) & (!g1367) & (!g1369) & (g1383) & (g1394)) + ((!g1068) & (g1354) & (!g1367) & (g1369) & (!g1383) & (g1394)) + ((!g1068) & (g1354) & (!g1367) & (g1369) & (g1383) & (!g1394)) + ((!g1068) & (g1354) & (g1367) & (!g1369) & (!g1383) & (g1394)) + ((!g1068) & (g1354) & (g1367) & (!g1369) & (g1383) & (g1394)) + ((!g1068) & (g1354) & (g1367) & (g1369) & (!g1383) & (g1394)) + ((!g1068) & (g1354) & (g1367) & (g1369) & (g1383) & (!g1394)) + ((g1068) & (!g1354) & (!g1367) & (!g1369) & (!g1383) & (!g1394)) + ((g1068) & (!g1354) & (!g1367) & (!g1369) & (g1383) & (!g1394)) + ((g1068) & (!g1354) & (!g1367) & (g1369) & (!g1383) & (!g1394)) + ((g1068) & (!g1354) & (!g1367) & (g1369) & (g1383) & (g1394)) + ((g1068) & (!g1354) & (g1367) & (!g1369) & (!g1383) & (!g1394)) + ((g1068) & (!g1354) & (g1367) & (!g1369) & (g1383) & (!g1394)) + ((g1068) & (!g1354) & (g1367) & (g1369) & (!g1383) & (!g1394)) + ((g1068) & (!g1354) & (g1367) & (g1369) & (g1383) & (g1394)) + ((g1068) & (g1354) & (!g1367) & (!g1369) & (!g1383) & (g1394)) + ((g1068) & (g1354) & (!g1367) & (!g1369) & (g1383) & (!g1394)) + ((g1068) & (g1354) & (!g1367) & (g1369) & (!g1383) & (!g1394)) + ((g1068) & (g1354) & (!g1367) & (g1369) & (g1383) & (!g1394)) + ((g1068) & (g1354) & (g1367) & (!g1369) & (!g1383) & (!g1394)) + ((g1068) & (g1354) & (g1367) & (!g1369) & (g1383) & (!g1394)) + ((g1068) & (g1354) & (g1367) & (g1369) & (!g1383) & (!g1394)) + ((g1068) & (g1354) & (g1367) & (g1369) & (g1383) & (g1394)));
	assign g1396 = (((g1355) & (g1352) & (!g1362) & (!g1365) & (g1366) & (!g1382)) + ((g1355) & (g1352) & (!g1362) & (g1365) & (!g1366) & (g1382)) + ((g1355) & (g1352) & (g1362) & (!g1365) & (!g1366) & (g1382)) + ((g1355) & (g1352) & (g1362) & (g1365) & (g1366) & (g1382)));
	assign g1397 = (((g1396) & (!sk[127]) & (g1394)) + ((g1396) & (sk[127]) & (g1394)));
	assign g1398 = (((!g1370) & (!g1372) & (!g1385) & (!sk[0]) & (g1381)) + ((!g1370) & (!g1372) & (!g1385) & (sk[0]) & (!g1381)) + ((!g1370) & (!g1372) & (!g1385) & (sk[0]) & (g1381)) + ((!g1370) & (!g1372) & (g1385) & (!sk[0]) & (g1381)) + ((!g1370) & (!g1372) & (g1385) & (sk[0]) & (g1381)) + ((!g1370) & (g1372) & (!g1385) & (!sk[0]) & (g1381)) + ((!g1370) & (g1372) & (!g1385) & (sk[0]) & (g1381)) + ((!g1370) & (g1372) & (g1385) & (!sk[0]) & (g1381)) + ((g1370) & (!g1372) & (!g1385) & (!sk[0]) & (!g1381)) + ((g1370) & (!g1372) & (!g1385) & (!sk[0]) & (g1381)) + ((g1370) & (!g1372) & (!g1385) & (sk[0]) & (g1381)) + ((g1370) & (!g1372) & (g1385) & (!sk[0]) & (!g1381)) + ((g1370) & (!g1372) & (g1385) & (!sk[0]) & (g1381)) + ((g1370) & (g1372) & (!g1385) & (!sk[0]) & (!g1381)) + ((g1370) & (g1372) & (!g1385) & (!sk[0]) & (g1381)) + ((g1370) & (g1372) & (!g1385) & (sk[0]) & (g1381)) + ((g1370) & (g1372) & (g1385) & (!sk[0]) & (!g1381)) + ((g1370) & (g1372) & (g1385) & (!sk[0]) & (g1381)));
	assign g1399 = (((!g252) & (!g994) & (!g1040) & (!g1079) & (sk[1]) & (g1387)) + ((!g252) & (!g994) & (!g1040) & (g1079) & (!sk[1]) & (!g1387)) + ((!g252) & (!g994) & (!g1040) & (g1079) & (!sk[1]) & (g1387)) + ((!g252) & (!g994) & (!g1040) & (g1079) & (sk[1]) & (g1387)) + ((!g252) & (!g994) & (g1040) & (!g1079) & (!sk[1]) & (!g1387)) + ((!g252) & (!g994) & (g1040) & (!g1079) & (!sk[1]) & (g1387)) + ((!g252) & (!g994) & (g1040) & (!g1079) & (sk[1]) & (g1387)) + ((!g252) & (!g994) & (g1040) & (g1079) & (!sk[1]) & (!g1387)) + ((!g252) & (!g994) & (g1040) & (g1079) & (!sk[1]) & (g1387)) + ((!g252) & (!g994) & (g1040) & (g1079) & (sk[1]) & (g1387)) + ((!g252) & (g994) & (!g1040) & (!g1079) & (!sk[1]) & (!g1387)) + ((!g252) & (g994) & (!g1040) & (!g1079) & (!sk[1]) & (g1387)) + ((!g252) & (g994) & (!g1040) & (!g1079) & (sk[1]) & (g1387)) + ((!g252) & (g994) & (!g1040) & (g1079) & (!sk[1]) & (!g1387)) + ((!g252) & (g994) & (!g1040) & (g1079) & (!sk[1]) & (g1387)) + ((!g252) & (g994) & (!g1040) & (g1079) & (sk[1]) & (g1387)) + ((!g252) & (g994) & (g1040) & (!g1079) & (!sk[1]) & (!g1387)) + ((!g252) & (g994) & (g1040) & (!g1079) & (!sk[1]) & (g1387)) + ((!g252) & (g994) & (g1040) & (!g1079) & (sk[1]) & (g1387)) + ((!g252) & (g994) & (g1040) & (g1079) & (!sk[1]) & (!g1387)) + ((!g252) & (g994) & (g1040) & (g1079) & (!sk[1]) & (g1387)) + ((!g252) & (g994) & (g1040) & (g1079) & (sk[1]) & (g1387)) + ((g252) & (!g994) & (!g1040) & (!g1079) & (sk[1]) & (!g1387)) + ((g252) & (!g994) & (!g1040) & (!g1079) & (sk[1]) & (g1387)) + ((g252) & (!g994) & (!g1040) & (g1079) & (!sk[1]) & (!g1387)) + ((g252) & (!g994) & (!g1040) & (g1079) & (!sk[1]) & (g1387)) + ((g252) & (!g994) & (g1040) & (!g1079) & (!sk[1]) & (!g1387)) + ((g252) & (!g994) & (g1040) & (!g1079) & (!sk[1]) & (g1387)) + ((g252) & (!g994) & (g1040) & (!g1079) & (sk[1]) & (g1387)) + ((g252) & (!g994) & (g1040) & (g1079) & (!sk[1]) & (!g1387)) + ((g252) & (!g994) & (g1040) & (g1079) & (!sk[1]) & (g1387)) + ((g252) & (!g994) & (g1040) & (g1079) & (sk[1]) & (!g1387)) + ((g252) & (g994) & (!g1040) & (!g1079) & (!sk[1]) & (!g1387)) + ((g252) & (g994) & (!g1040) & (!g1079) & (!sk[1]) & (g1387)) + ((g252) & (g994) & (!g1040) & (!g1079) & (sk[1]) & (!g1387)) + ((g252) & (g994) & (!g1040) & (g1079) & (!sk[1]) & (!g1387)) + ((g252) & (g994) & (!g1040) & (g1079) & (!sk[1]) & (g1387)) + ((g252) & (g994) & (!g1040) & (g1079) & (sk[1]) & (g1387)) + ((g252) & (g994) & (g1040) & (!g1079) & (!sk[1]) & (!g1387)) + ((g252) & (g994) & (g1040) & (!g1079) & (!sk[1]) & (g1387)) + ((g252) & (g994) & (g1040) & (!g1079) & (sk[1]) & (!g1387)) + ((g252) & (g994) & (g1040) & (!g1079) & (sk[1]) & (g1387)) + ((g252) & (g994) & (g1040) & (g1079) & (!sk[1]) & (!g1387)) + ((g252) & (g994) & (g1040) & (g1079) & (!sk[1]) & (g1387)));
	assign g1400 = (((!g1373) & (!g1377) & (!g1378) & (!g1386) & (!g1388) & (g1399)) + ((!g1373) & (!g1377) & (!g1378) & (!g1386) & (g1388) & (g1399)) + ((!g1373) & (!g1377) & (!g1378) & (g1386) & (!g1388) & (!g1399)) + ((!g1373) & (!g1377) & (!g1378) & (g1386) & (g1388) & (g1399)) + ((!g1373) & (!g1377) & (g1378) & (!g1386) & (!g1388) & (!g1399)) + ((!g1373) & (!g1377) & (g1378) & (!g1386) & (g1388) & (g1399)) + ((!g1373) & (!g1377) & (g1378) & (g1386) & (!g1388) & (!g1399)) + ((!g1373) & (!g1377) & (g1378) & (g1386) & (g1388) & (!g1399)) + ((!g1373) & (g1377) & (!g1378) & (!g1386) & (!g1388) & (!g1399)) + ((!g1373) & (g1377) & (!g1378) & (!g1386) & (g1388) & (g1399)) + ((!g1373) & (g1377) & (!g1378) & (g1386) & (!g1388) & (!g1399)) + ((!g1373) & (g1377) & (!g1378) & (g1386) & (g1388) & (!g1399)) + ((!g1373) & (g1377) & (g1378) & (!g1386) & (!g1388) & (!g1399)) + ((!g1373) & (g1377) & (g1378) & (!g1386) & (g1388) & (g1399)) + ((!g1373) & (g1377) & (g1378) & (g1386) & (!g1388) & (!g1399)) + ((!g1373) & (g1377) & (g1378) & (g1386) & (g1388) & (!g1399)) + ((g1373) & (!g1377) & (!g1378) & (!g1386) & (!g1388) & (g1399)) + ((g1373) & (!g1377) & (!g1378) & (!g1386) & (g1388) & (g1399)) + ((g1373) & (!g1377) & (!g1378) & (g1386) & (!g1388) & (!g1399)) + ((g1373) & (!g1377) & (!g1378) & (g1386) & (g1388) & (g1399)) + ((g1373) & (!g1377) & (g1378) & (!g1386) & (!g1388) & (g1399)) + ((g1373) & (!g1377) & (g1378) & (!g1386) & (g1388) & (g1399)) + ((g1373) & (!g1377) & (g1378) & (g1386) & (!g1388) & (!g1399)) + ((g1373) & (!g1377) & (g1378) & (g1386) & (g1388) & (g1399)) + ((g1373) & (g1377) & (!g1378) & (!g1386) & (!g1388) & (g1399)) + ((g1373) & (g1377) & (!g1378) & (!g1386) & (g1388) & (g1399)) + ((g1373) & (g1377) & (!g1378) & (g1386) & (!g1388) & (!g1399)) + ((g1373) & (g1377) & (!g1378) & (g1386) & (g1388) & (g1399)) + ((g1373) & (g1377) & (g1378) & (!g1386) & (!g1388) & (!g1399)) + ((g1373) & (g1377) & (g1378) & (!g1386) & (g1388) & (g1399)) + ((g1373) & (g1377) & (g1378) & (g1386) & (!g1388) & (!g1399)) + ((g1373) & (g1377) & (g1378) & (g1386) & (g1388) & (!g1399)));
	assign g1401 = (((!sk[3]) & (!g9) & (!g49) & (!g25) & (g826)) + ((!sk[3]) & (!g9) & (!g49) & (g25) & (g826)) + ((!sk[3]) & (!g9) & (g49) & (!g25) & (g826)) + ((!sk[3]) & (!g9) & (g49) & (g25) & (g826)) + ((!sk[3]) & (g9) & (!g49) & (!g25) & (!g826)) + ((!sk[3]) & (g9) & (!g49) & (!g25) & (g826)) + ((!sk[3]) & (g9) & (!g49) & (g25) & (!g826)) + ((!sk[3]) & (g9) & (!g49) & (g25) & (g826)) + ((!sk[3]) & (g9) & (g49) & (!g25) & (!g826)) + ((!sk[3]) & (g9) & (g49) & (!g25) & (g826)) + ((!sk[3]) & (g9) & (g49) & (g25) & (!g826)) + ((!sk[3]) & (g9) & (g49) & (g25) & (g826)) + ((sk[3]) & (!g9) & (!g49) & (!g25) & (g826)) + ((sk[3]) & (!g9) & (!g49) & (g25) & (g826)) + ((sk[3]) & (!g9) & (g49) & (!g25) & (g826)) + ((sk[3]) & (!g9) & (g49) & (g25) & (g826)) + ((sk[3]) & (g9) & (!g49) & (!g25) & (g826)));
	assign g1402 = (((!sk[4]) & (!g112) & (!g113) & (!g97) & (g98) & (!g16)) + ((!sk[4]) & (!g112) & (!g113) & (!g97) & (g98) & (g16)) + ((!sk[4]) & (!g112) & (!g113) & (g97) & (!g98) & (!g16)) + ((!sk[4]) & (!g112) & (!g113) & (g97) & (!g98) & (g16)) + ((!sk[4]) & (!g112) & (!g113) & (g97) & (g98) & (!g16)) + ((!sk[4]) & (!g112) & (!g113) & (g97) & (g98) & (g16)) + ((!sk[4]) & (!g112) & (g113) & (!g97) & (!g98) & (!g16)) + ((!sk[4]) & (!g112) & (g113) & (!g97) & (!g98) & (g16)) + ((!sk[4]) & (!g112) & (g113) & (!g97) & (g98) & (!g16)) + ((!sk[4]) & (!g112) & (g113) & (!g97) & (g98) & (g16)) + ((!sk[4]) & (!g112) & (g113) & (g97) & (!g98) & (!g16)) + ((!sk[4]) & (!g112) & (g113) & (g97) & (!g98) & (g16)) + ((!sk[4]) & (!g112) & (g113) & (g97) & (g98) & (!g16)) + ((!sk[4]) & (!g112) & (g113) & (g97) & (g98) & (g16)) + ((!sk[4]) & (g112) & (!g113) & (!g97) & (g98) & (!g16)) + ((!sk[4]) & (g112) & (!g113) & (!g97) & (g98) & (g16)) + ((!sk[4]) & (g112) & (!g113) & (g97) & (!g98) & (!g16)) + ((!sk[4]) & (g112) & (!g113) & (g97) & (!g98) & (g16)) + ((!sk[4]) & (g112) & (!g113) & (g97) & (g98) & (!g16)) + ((!sk[4]) & (g112) & (!g113) & (g97) & (g98) & (g16)) + ((!sk[4]) & (g112) & (g113) & (!g97) & (!g98) & (!g16)) + ((!sk[4]) & (g112) & (g113) & (!g97) & (!g98) & (g16)) + ((!sk[4]) & (g112) & (g113) & (!g97) & (g98) & (!g16)) + ((!sk[4]) & (g112) & (g113) & (!g97) & (g98) & (g16)) + ((!sk[4]) & (g112) & (g113) & (g97) & (!g98) & (!g16)) + ((!sk[4]) & (g112) & (g113) & (g97) & (!g98) & (g16)) + ((!sk[4]) & (g112) & (g113) & (g97) & (g98) & (!g16)) + ((!sk[4]) & (g112) & (g113) & (g97) & (g98) & (g16)) + ((sk[4]) & (!g112) & (!g113) & (!g97) & (g98) & (g16)) + ((sk[4]) & (!g112) & (g113) & (g97) & (g98) & (g16)) + ((sk[4]) & (g112) & (!g113) & (!g97) & (!g98) & (g16)) + ((sk[4]) & (g112) & (!g113) & (g97) & (g98) & (g16)) + ((sk[4]) & (g112) & (g113) & (g97) & (!g98) & (g16)) + ((sk[4]) & (g112) & (g113) & (g97) & (g98) & (g16)));
	assign g1403 = (((!g70) & (!g10) & (!sk[5]) & (!g99) & (g42) & (!g1402)) + ((!g70) & (!g10) & (!sk[5]) & (!g99) & (g42) & (g1402)) + ((!g70) & (!g10) & (!sk[5]) & (g99) & (!g42) & (!g1402)) + ((!g70) & (!g10) & (!sk[5]) & (g99) & (!g42) & (g1402)) + ((!g70) & (!g10) & (!sk[5]) & (g99) & (g42) & (!g1402)) + ((!g70) & (!g10) & (!sk[5]) & (g99) & (g42) & (g1402)) + ((!g70) & (!g10) & (sk[5]) & (!g99) & (!g42) & (!g1402)) + ((!g70) & (!g10) & (sk[5]) & (!g99) & (g42) & (!g1402)) + ((!g70) & (!g10) & (sk[5]) & (g99) & (!g42) & (!g1402)) + ((!g70) & (!g10) & (sk[5]) & (g99) & (g42) & (!g1402)) + ((!g70) & (g10) & (!sk[5]) & (!g99) & (!g42) & (!g1402)) + ((!g70) & (g10) & (!sk[5]) & (!g99) & (!g42) & (g1402)) + ((!g70) & (g10) & (!sk[5]) & (!g99) & (g42) & (!g1402)) + ((!g70) & (g10) & (!sk[5]) & (!g99) & (g42) & (g1402)) + ((!g70) & (g10) & (!sk[5]) & (g99) & (!g42) & (!g1402)) + ((!g70) & (g10) & (!sk[5]) & (g99) & (!g42) & (g1402)) + ((!g70) & (g10) & (!sk[5]) & (g99) & (g42) & (!g1402)) + ((!g70) & (g10) & (!sk[5]) & (g99) & (g42) & (g1402)) + ((!g70) & (g10) & (sk[5]) & (!g99) & (!g42) & (!g1402)) + ((!g70) & (g10) & (sk[5]) & (!g99) & (g42) & (!g1402)) + ((g70) & (!g10) & (!sk[5]) & (!g99) & (g42) & (!g1402)) + ((g70) & (!g10) & (!sk[5]) & (!g99) & (g42) & (g1402)) + ((g70) & (!g10) & (!sk[5]) & (g99) & (!g42) & (!g1402)) + ((g70) & (!g10) & (!sk[5]) & (g99) & (!g42) & (g1402)) + ((g70) & (!g10) & (!sk[5]) & (g99) & (g42) & (!g1402)) + ((g70) & (!g10) & (!sk[5]) & (g99) & (g42) & (g1402)) + ((g70) & (!g10) & (sk[5]) & (!g99) & (!g42) & (!g1402)) + ((g70) & (!g10) & (sk[5]) & (g99) & (!g42) & (!g1402)) + ((g70) & (g10) & (!sk[5]) & (!g99) & (!g42) & (!g1402)) + ((g70) & (g10) & (!sk[5]) & (!g99) & (!g42) & (g1402)) + ((g70) & (g10) & (!sk[5]) & (!g99) & (g42) & (!g1402)) + ((g70) & (g10) & (!sk[5]) & (!g99) & (g42) & (g1402)) + ((g70) & (g10) & (!sk[5]) & (g99) & (!g42) & (!g1402)) + ((g70) & (g10) & (!sk[5]) & (g99) & (!g42) & (g1402)) + ((g70) & (g10) & (!sk[5]) & (g99) & (g42) & (!g1402)) + ((g70) & (g10) & (!sk[5]) & (g99) & (g42) & (g1402)) + ((g70) & (g10) & (sk[5]) & (!g99) & (!g42) & (!g1402)));
	assign g1404 = (((!sk[6]) & (!g62) & (!g91) & (!g651) & (g1401) & (!g1403)) + ((!sk[6]) & (!g62) & (!g91) & (!g651) & (g1401) & (g1403)) + ((!sk[6]) & (!g62) & (!g91) & (g651) & (!g1401) & (!g1403)) + ((!sk[6]) & (!g62) & (!g91) & (g651) & (!g1401) & (g1403)) + ((!sk[6]) & (!g62) & (!g91) & (g651) & (g1401) & (!g1403)) + ((!sk[6]) & (!g62) & (!g91) & (g651) & (g1401) & (g1403)) + ((!sk[6]) & (!g62) & (g91) & (!g651) & (!g1401) & (!g1403)) + ((!sk[6]) & (!g62) & (g91) & (!g651) & (!g1401) & (g1403)) + ((!sk[6]) & (!g62) & (g91) & (!g651) & (g1401) & (!g1403)) + ((!sk[6]) & (!g62) & (g91) & (!g651) & (g1401) & (g1403)) + ((!sk[6]) & (!g62) & (g91) & (g651) & (!g1401) & (!g1403)) + ((!sk[6]) & (!g62) & (g91) & (g651) & (!g1401) & (g1403)) + ((!sk[6]) & (!g62) & (g91) & (g651) & (g1401) & (!g1403)) + ((!sk[6]) & (!g62) & (g91) & (g651) & (g1401) & (g1403)) + ((!sk[6]) & (g62) & (!g91) & (!g651) & (g1401) & (!g1403)) + ((!sk[6]) & (g62) & (!g91) & (!g651) & (g1401) & (g1403)) + ((!sk[6]) & (g62) & (!g91) & (g651) & (!g1401) & (!g1403)) + ((!sk[6]) & (g62) & (!g91) & (g651) & (!g1401) & (g1403)) + ((!sk[6]) & (g62) & (!g91) & (g651) & (g1401) & (!g1403)) + ((!sk[6]) & (g62) & (!g91) & (g651) & (g1401) & (g1403)) + ((!sk[6]) & (g62) & (g91) & (!g651) & (!g1401) & (!g1403)) + ((!sk[6]) & (g62) & (g91) & (!g651) & (!g1401) & (g1403)) + ((!sk[6]) & (g62) & (g91) & (!g651) & (g1401) & (!g1403)) + ((!sk[6]) & (g62) & (g91) & (!g651) & (g1401) & (g1403)) + ((!sk[6]) & (g62) & (g91) & (g651) & (!g1401) & (!g1403)) + ((!sk[6]) & (g62) & (g91) & (g651) & (!g1401) & (g1403)) + ((!sk[6]) & (g62) & (g91) & (g651) & (g1401) & (!g1403)) + ((!sk[6]) & (g62) & (g91) & (g651) & (g1401) & (g1403)) + ((sk[6]) & (!g62) & (!g91) & (!g651) & (g1401) & (g1403)) + ((sk[6]) & (!g62) & (g91) & (!g651) & (g1401) & (g1403)) + ((sk[6]) & (g62) & (!g91) & (!g651) & (g1401) & (g1403)));
	assign g1405 = (((!g270) & (!g125) & (!sk[7]) & (!g586) & (g1026) & (!g1404)) + ((!g270) & (!g125) & (!sk[7]) & (!g586) & (g1026) & (g1404)) + ((!g270) & (!g125) & (!sk[7]) & (g586) & (!g1026) & (!g1404)) + ((!g270) & (!g125) & (!sk[7]) & (g586) & (!g1026) & (g1404)) + ((!g270) & (!g125) & (!sk[7]) & (g586) & (g1026) & (!g1404)) + ((!g270) & (!g125) & (!sk[7]) & (g586) & (g1026) & (g1404)) + ((!g270) & (g125) & (!sk[7]) & (!g586) & (!g1026) & (!g1404)) + ((!g270) & (g125) & (!sk[7]) & (!g586) & (!g1026) & (g1404)) + ((!g270) & (g125) & (!sk[7]) & (!g586) & (g1026) & (!g1404)) + ((!g270) & (g125) & (!sk[7]) & (!g586) & (g1026) & (g1404)) + ((!g270) & (g125) & (!sk[7]) & (g586) & (!g1026) & (!g1404)) + ((!g270) & (g125) & (!sk[7]) & (g586) & (!g1026) & (g1404)) + ((!g270) & (g125) & (!sk[7]) & (g586) & (g1026) & (!g1404)) + ((!g270) & (g125) & (!sk[7]) & (g586) & (g1026) & (g1404)) + ((g270) & (!g125) & (!sk[7]) & (!g586) & (g1026) & (!g1404)) + ((g270) & (!g125) & (!sk[7]) & (!g586) & (g1026) & (g1404)) + ((g270) & (!g125) & (!sk[7]) & (g586) & (!g1026) & (!g1404)) + ((g270) & (!g125) & (!sk[7]) & (g586) & (!g1026) & (g1404)) + ((g270) & (!g125) & (!sk[7]) & (g586) & (g1026) & (!g1404)) + ((g270) & (!g125) & (!sk[7]) & (g586) & (g1026) & (g1404)) + ((g270) & (g125) & (!sk[7]) & (!g586) & (!g1026) & (!g1404)) + ((g270) & (g125) & (!sk[7]) & (!g586) & (!g1026) & (g1404)) + ((g270) & (g125) & (!sk[7]) & (!g586) & (g1026) & (!g1404)) + ((g270) & (g125) & (!sk[7]) & (!g586) & (g1026) & (g1404)) + ((g270) & (g125) & (!sk[7]) & (g586) & (!g1026) & (!g1404)) + ((g270) & (g125) & (!sk[7]) & (g586) & (!g1026) & (g1404)) + ((g270) & (g125) & (!sk[7]) & (g586) & (g1026) & (!g1404)) + ((g270) & (g125) & (!sk[7]) & (g586) & (g1026) & (g1404)) + ((g270) & (g125) & (sk[7]) & (g586) & (g1026) & (g1404)));
	assign g1406 = (((!sk[8]) & (!g1389) & (!g1393) & (!g1398) & (g1400) & (!g1405)) + ((!sk[8]) & (!g1389) & (!g1393) & (!g1398) & (g1400) & (g1405)) + ((!sk[8]) & (!g1389) & (!g1393) & (g1398) & (!g1400) & (!g1405)) + ((!sk[8]) & (!g1389) & (!g1393) & (g1398) & (!g1400) & (g1405)) + ((!sk[8]) & (!g1389) & (!g1393) & (g1398) & (g1400) & (!g1405)) + ((!sk[8]) & (!g1389) & (!g1393) & (g1398) & (g1400) & (g1405)) + ((!sk[8]) & (!g1389) & (g1393) & (!g1398) & (!g1400) & (!g1405)) + ((!sk[8]) & (!g1389) & (g1393) & (!g1398) & (!g1400) & (g1405)) + ((!sk[8]) & (!g1389) & (g1393) & (!g1398) & (g1400) & (!g1405)) + ((!sk[8]) & (!g1389) & (g1393) & (!g1398) & (g1400) & (g1405)) + ((!sk[8]) & (!g1389) & (g1393) & (g1398) & (!g1400) & (!g1405)) + ((!sk[8]) & (!g1389) & (g1393) & (g1398) & (!g1400) & (g1405)) + ((!sk[8]) & (!g1389) & (g1393) & (g1398) & (g1400) & (!g1405)) + ((!sk[8]) & (!g1389) & (g1393) & (g1398) & (g1400) & (g1405)) + ((!sk[8]) & (g1389) & (!g1393) & (!g1398) & (g1400) & (!g1405)) + ((!sk[8]) & (g1389) & (!g1393) & (!g1398) & (g1400) & (g1405)) + ((!sk[8]) & (g1389) & (!g1393) & (g1398) & (!g1400) & (!g1405)) + ((!sk[8]) & (g1389) & (!g1393) & (g1398) & (!g1400) & (g1405)) + ((!sk[8]) & (g1389) & (!g1393) & (g1398) & (g1400) & (!g1405)) + ((!sk[8]) & (g1389) & (!g1393) & (g1398) & (g1400) & (g1405)) + ((!sk[8]) & (g1389) & (g1393) & (!g1398) & (!g1400) & (!g1405)) + ((!sk[8]) & (g1389) & (g1393) & (!g1398) & (!g1400) & (g1405)) + ((!sk[8]) & (g1389) & (g1393) & (!g1398) & (g1400) & (!g1405)) + ((!sk[8]) & (g1389) & (g1393) & (!g1398) & (g1400) & (g1405)) + ((!sk[8]) & (g1389) & (g1393) & (g1398) & (!g1400) & (!g1405)) + ((!sk[8]) & (g1389) & (g1393) & (g1398) & (!g1400) & (g1405)) + ((!sk[8]) & (g1389) & (g1393) & (g1398) & (g1400) & (!g1405)) + ((!sk[8]) & (g1389) & (g1393) & (g1398) & (g1400) & (g1405)) + ((sk[8]) & (!g1389) & (!g1393) & (!g1398) & (!g1400) & (g1405)) + ((sk[8]) & (!g1389) & (!g1393) & (!g1398) & (g1400) & (!g1405)) + ((sk[8]) & (!g1389) & (!g1393) & (g1398) & (!g1400) & (g1405)) + ((sk[8]) & (!g1389) & (!g1393) & (g1398) & (g1400) & (!g1405)) + ((sk[8]) & (!g1389) & (g1393) & (!g1398) & (!g1400) & (g1405)) + ((sk[8]) & (!g1389) & (g1393) & (!g1398) & (g1400) & (!g1405)) + ((sk[8]) & (!g1389) & (g1393) & (g1398) & (!g1400) & (!g1405)) + ((sk[8]) & (!g1389) & (g1393) & (g1398) & (g1400) & (g1405)) + ((sk[8]) & (g1389) & (!g1393) & (!g1398) & (!g1400) & (g1405)) + ((sk[8]) & (g1389) & (!g1393) & (!g1398) & (g1400) & (!g1405)) + ((sk[8]) & (g1389) & (!g1393) & (g1398) & (!g1400) & (!g1405)) + ((sk[8]) & (g1389) & (!g1393) & (g1398) & (g1400) & (g1405)) + ((sk[8]) & (g1389) & (g1393) & (!g1398) & (!g1400) & (!g1405)) + ((sk[8]) & (g1389) & (g1393) & (!g1398) & (g1400) & (g1405)) + ((sk[8]) & (g1389) & (g1393) & (g1398) & (!g1400) & (!g1405)) + ((sk[8]) & (g1389) & (g1393) & (g1398) & (g1400) & (g1405)));
	assign g1407 = (((!sk[9]) & (!g1354) & (!g1367) & (!g1369) & (g1383) & (!g1394)) + ((!sk[9]) & (!g1354) & (!g1367) & (!g1369) & (g1383) & (g1394)) + ((!sk[9]) & (!g1354) & (!g1367) & (g1369) & (!g1383) & (!g1394)) + ((!sk[9]) & (!g1354) & (!g1367) & (g1369) & (!g1383) & (g1394)) + ((!sk[9]) & (!g1354) & (!g1367) & (g1369) & (g1383) & (!g1394)) + ((!sk[9]) & (!g1354) & (!g1367) & (g1369) & (g1383) & (g1394)) + ((!sk[9]) & (!g1354) & (g1367) & (!g1369) & (!g1383) & (!g1394)) + ((!sk[9]) & (!g1354) & (g1367) & (!g1369) & (!g1383) & (g1394)) + ((!sk[9]) & (!g1354) & (g1367) & (!g1369) & (g1383) & (!g1394)) + ((!sk[9]) & (!g1354) & (g1367) & (!g1369) & (g1383) & (g1394)) + ((!sk[9]) & (!g1354) & (g1367) & (g1369) & (!g1383) & (!g1394)) + ((!sk[9]) & (!g1354) & (g1367) & (g1369) & (!g1383) & (g1394)) + ((!sk[9]) & (!g1354) & (g1367) & (g1369) & (g1383) & (!g1394)) + ((!sk[9]) & (!g1354) & (g1367) & (g1369) & (g1383) & (g1394)) + ((!sk[9]) & (g1354) & (!g1367) & (!g1369) & (g1383) & (!g1394)) + ((!sk[9]) & (g1354) & (!g1367) & (!g1369) & (g1383) & (g1394)) + ((!sk[9]) & (g1354) & (!g1367) & (g1369) & (!g1383) & (!g1394)) + ((!sk[9]) & (g1354) & (!g1367) & (g1369) & (!g1383) & (g1394)) + ((!sk[9]) & (g1354) & (!g1367) & (g1369) & (g1383) & (!g1394)) + ((!sk[9]) & (g1354) & (!g1367) & (g1369) & (g1383) & (g1394)) + ((!sk[9]) & (g1354) & (g1367) & (!g1369) & (!g1383) & (!g1394)) + ((!sk[9]) & (g1354) & (g1367) & (!g1369) & (!g1383) & (g1394)) + ((!sk[9]) & (g1354) & (g1367) & (!g1369) & (g1383) & (!g1394)) + ((!sk[9]) & (g1354) & (g1367) & (!g1369) & (g1383) & (g1394)) + ((!sk[9]) & (g1354) & (g1367) & (g1369) & (!g1383) & (!g1394)) + ((!sk[9]) & (g1354) & (g1367) & (g1369) & (!g1383) & (g1394)) + ((!sk[9]) & (g1354) & (g1367) & (g1369) & (g1383) & (!g1394)) + ((!sk[9]) & (g1354) & (g1367) & (g1369) & (g1383) & (g1394)) + ((sk[9]) & (g1354) & (!g1367) & (!g1369) & (!g1383) & (!g1394)) + ((sk[9]) & (g1354) & (!g1367) & (g1369) & (g1383) & (g1394)));
	assign sinx16x = (((!g1068) & (!g1397) & (!g1406) & (!sk[10]) & (g1407)) + ((!g1068) & (!g1397) & (g1406) & (!sk[10]) & (g1407)) + ((!g1068) & (!g1397) & (g1406) & (sk[10]) & (!g1407)) + ((!g1068) & (!g1397) & (g1406) & (sk[10]) & (g1407)) + ((!g1068) & (g1397) & (!g1406) & (!sk[10]) & (g1407)) + ((!g1068) & (g1397) & (!g1406) & (sk[10]) & (!g1407)) + ((!g1068) & (g1397) & (!g1406) & (sk[10]) & (g1407)) + ((!g1068) & (g1397) & (g1406) & (!sk[10]) & (g1407)) + ((g1068) & (!g1397) & (!g1406) & (!sk[10]) & (!g1407)) + ((g1068) & (!g1397) & (!g1406) & (!sk[10]) & (g1407)) + ((g1068) & (!g1397) & (!g1406) & (sk[10]) & (!g1407)) + ((g1068) & (!g1397) & (g1406) & (!sk[10]) & (!g1407)) + ((g1068) & (!g1397) & (g1406) & (!sk[10]) & (g1407)) + ((g1068) & (!g1397) & (g1406) & (sk[10]) & (g1407)) + ((g1068) & (g1397) & (!g1406) & (!sk[10]) & (!g1407)) + ((g1068) & (g1397) & (!g1406) & (!sk[10]) & (g1407)) + ((g1068) & (g1397) & (!g1406) & (sk[10]) & (g1407)) + ((g1068) & (g1397) & (g1406) & (!sk[10]) & (!g1407)) + ((g1068) & (g1397) & (g1406) & (!sk[10]) & (g1407)) + ((g1068) & (g1397) & (g1406) & (sk[10]) & (!g1407)));
	assign g1409 = (((!g1389) & (!g1393) & (!sk[11]) & (!g1398) & (g1400) & (!g1405)) + ((!g1389) & (!g1393) & (!sk[11]) & (!g1398) & (g1400) & (g1405)) + ((!g1389) & (!g1393) & (!sk[11]) & (g1398) & (!g1400) & (!g1405)) + ((!g1389) & (!g1393) & (!sk[11]) & (g1398) & (!g1400) & (g1405)) + ((!g1389) & (!g1393) & (!sk[11]) & (g1398) & (g1400) & (!g1405)) + ((!g1389) & (!g1393) & (!sk[11]) & (g1398) & (g1400) & (g1405)) + ((!g1389) & (!g1393) & (sk[11]) & (!g1398) & (!g1400) & (!g1405)) + ((!g1389) & (!g1393) & (sk[11]) & (!g1398) & (g1400) & (!g1405)) + ((!g1389) & (!g1393) & (sk[11]) & (!g1398) & (g1400) & (g1405)) + ((!g1389) & (!g1393) & (sk[11]) & (g1398) & (!g1400) & (!g1405)) + ((!g1389) & (!g1393) & (sk[11]) & (g1398) & (g1400) & (!g1405)) + ((!g1389) & (!g1393) & (sk[11]) & (g1398) & (g1400) & (g1405)) + ((!g1389) & (g1393) & (!sk[11]) & (!g1398) & (!g1400) & (!g1405)) + ((!g1389) & (g1393) & (!sk[11]) & (!g1398) & (!g1400) & (g1405)) + ((!g1389) & (g1393) & (!sk[11]) & (!g1398) & (g1400) & (!g1405)) + ((!g1389) & (g1393) & (!sk[11]) & (!g1398) & (g1400) & (g1405)) + ((!g1389) & (g1393) & (!sk[11]) & (g1398) & (!g1400) & (!g1405)) + ((!g1389) & (g1393) & (!sk[11]) & (g1398) & (!g1400) & (g1405)) + ((!g1389) & (g1393) & (!sk[11]) & (g1398) & (g1400) & (!g1405)) + ((!g1389) & (g1393) & (!sk[11]) & (g1398) & (g1400) & (g1405)) + ((!g1389) & (g1393) & (sk[11]) & (!g1398) & (!g1400) & (!g1405)) + ((!g1389) & (g1393) & (sk[11]) & (!g1398) & (g1400) & (!g1405)) + ((!g1389) & (g1393) & (sk[11]) & (!g1398) & (g1400) & (g1405)) + ((!g1389) & (g1393) & (sk[11]) & (g1398) & (g1400) & (!g1405)) + ((g1389) & (!g1393) & (!sk[11]) & (!g1398) & (g1400) & (!g1405)) + ((g1389) & (!g1393) & (!sk[11]) & (!g1398) & (g1400) & (g1405)) + ((g1389) & (!g1393) & (!sk[11]) & (g1398) & (!g1400) & (!g1405)) + ((g1389) & (!g1393) & (!sk[11]) & (g1398) & (!g1400) & (g1405)) + ((g1389) & (!g1393) & (!sk[11]) & (g1398) & (g1400) & (!g1405)) + ((g1389) & (!g1393) & (!sk[11]) & (g1398) & (g1400) & (g1405)) + ((g1389) & (!g1393) & (sk[11]) & (!g1398) & (!g1400) & (!g1405)) + ((g1389) & (!g1393) & (sk[11]) & (!g1398) & (g1400) & (!g1405)) + ((g1389) & (!g1393) & (sk[11]) & (!g1398) & (g1400) & (g1405)) + ((g1389) & (!g1393) & (sk[11]) & (g1398) & (g1400) & (!g1405)) + ((g1389) & (g1393) & (!sk[11]) & (!g1398) & (!g1400) & (!g1405)) + ((g1389) & (g1393) & (!sk[11]) & (!g1398) & (!g1400) & (g1405)) + ((g1389) & (g1393) & (!sk[11]) & (!g1398) & (g1400) & (!g1405)) + ((g1389) & (g1393) & (!sk[11]) & (!g1398) & (g1400) & (g1405)) + ((g1389) & (g1393) & (!sk[11]) & (g1398) & (!g1400) & (!g1405)) + ((g1389) & (g1393) & (!sk[11]) & (g1398) & (!g1400) & (g1405)) + ((g1389) & (g1393) & (!sk[11]) & (g1398) & (g1400) & (!g1405)) + ((g1389) & (g1393) & (!sk[11]) & (g1398) & (g1400) & (g1405)) + ((g1389) & (g1393) & (sk[11]) & (!g1398) & (g1400) & (!g1405)) + ((g1389) & (g1393) & (sk[11]) & (g1398) & (g1400) & (!g1405)));
	assign g1410 = (((!g9) & (!g12) & (!sk[12]) & (!g23) & (g47)) + ((!g9) & (!g12) & (!sk[12]) & (g23) & (g47)) + ((!g9) & (!g12) & (sk[12]) & (!g23) & (!g47)) + ((!g9) & (!g12) & (sk[12]) & (g23) & (!g47)) + ((!g9) & (g12) & (!sk[12]) & (!g23) & (g47)) + ((!g9) & (g12) & (!sk[12]) & (g23) & (g47)) + ((!g9) & (g12) & (sk[12]) & (!g23) & (!g47)) + ((!g9) & (g12) & (sk[12]) & (g23) & (!g47)) + ((g9) & (!g12) & (!sk[12]) & (!g23) & (!g47)) + ((g9) & (!g12) & (!sk[12]) & (!g23) & (g47)) + ((g9) & (!g12) & (!sk[12]) & (g23) & (!g47)) + ((g9) & (!g12) & (!sk[12]) & (g23) & (g47)) + ((g9) & (!g12) & (sk[12]) & (!g23) & (!g47)) + ((g9) & (g12) & (!sk[12]) & (!g23) & (!g47)) + ((g9) & (g12) & (!sk[12]) & (!g23) & (g47)) + ((g9) & (g12) & (!sk[12]) & (g23) & (!g47)) + ((g9) & (g12) & (!sk[12]) & (g23) & (g47)));
	assign g1411 = (((!sk[13]) & (!g16) & (!g127) & (!g152) & (g119) & (!g1410)) + ((!sk[13]) & (!g16) & (!g127) & (!g152) & (g119) & (g1410)) + ((!sk[13]) & (!g16) & (!g127) & (g152) & (!g119) & (!g1410)) + ((!sk[13]) & (!g16) & (!g127) & (g152) & (!g119) & (g1410)) + ((!sk[13]) & (!g16) & (!g127) & (g152) & (g119) & (!g1410)) + ((!sk[13]) & (!g16) & (!g127) & (g152) & (g119) & (g1410)) + ((!sk[13]) & (!g16) & (g127) & (!g152) & (!g119) & (!g1410)) + ((!sk[13]) & (!g16) & (g127) & (!g152) & (!g119) & (g1410)) + ((!sk[13]) & (!g16) & (g127) & (!g152) & (g119) & (!g1410)) + ((!sk[13]) & (!g16) & (g127) & (!g152) & (g119) & (g1410)) + ((!sk[13]) & (!g16) & (g127) & (g152) & (!g119) & (!g1410)) + ((!sk[13]) & (!g16) & (g127) & (g152) & (!g119) & (g1410)) + ((!sk[13]) & (!g16) & (g127) & (g152) & (g119) & (!g1410)) + ((!sk[13]) & (!g16) & (g127) & (g152) & (g119) & (g1410)) + ((!sk[13]) & (g16) & (!g127) & (!g152) & (g119) & (!g1410)) + ((!sk[13]) & (g16) & (!g127) & (!g152) & (g119) & (g1410)) + ((!sk[13]) & (g16) & (!g127) & (g152) & (!g119) & (!g1410)) + ((!sk[13]) & (g16) & (!g127) & (g152) & (!g119) & (g1410)) + ((!sk[13]) & (g16) & (!g127) & (g152) & (g119) & (!g1410)) + ((!sk[13]) & (g16) & (!g127) & (g152) & (g119) & (g1410)) + ((!sk[13]) & (g16) & (g127) & (!g152) & (!g119) & (!g1410)) + ((!sk[13]) & (g16) & (g127) & (!g152) & (!g119) & (g1410)) + ((!sk[13]) & (g16) & (g127) & (!g152) & (g119) & (!g1410)) + ((!sk[13]) & (g16) & (g127) & (!g152) & (g119) & (g1410)) + ((!sk[13]) & (g16) & (g127) & (g152) & (!g119) & (!g1410)) + ((!sk[13]) & (g16) & (g127) & (g152) & (!g119) & (g1410)) + ((!sk[13]) & (g16) & (g127) & (g152) & (g119) & (!g1410)) + ((!sk[13]) & (g16) & (g127) & (g152) & (g119) & (g1410)) + ((sk[13]) & (!g16) & (!g127) & (!g152) & (!g119) & (g1410)) + ((sk[13]) & (!g16) & (!g127) & (!g152) & (g119) & (g1410)) + ((sk[13]) & (g16) & (!g127) & (!g152) & (!g119) & (g1410)));
	assign g1412 = (((g240) & (g75) & (g269) & (g878) & (g1020) & (g1411)));
	assign sinx17x = (((!g1068) & (!g1397) & (!g1409) & (!g1406) & (!g1407) & (!g1412)) + ((!g1068) & (!g1397) & (!g1409) & (!g1406) & (g1407) & (!g1412)) + ((!g1068) & (!g1397) & (!g1409) & (g1406) & (!g1407) & (!g1412)) + ((!g1068) & (!g1397) & (!g1409) & (g1406) & (g1407) & (!g1412)) + ((!g1068) & (!g1397) & (g1409) & (!g1406) & (!g1407) & (g1412)) + ((!g1068) & (!g1397) & (g1409) & (!g1406) & (g1407) & (g1412)) + ((!g1068) & (!g1397) & (g1409) & (g1406) & (!g1407) & (g1412)) + ((!g1068) & (!g1397) & (g1409) & (g1406) & (g1407) & (g1412)) + ((!g1068) & (g1397) & (!g1409) & (!g1406) & (!g1407) & (!g1412)) + ((!g1068) & (g1397) & (!g1409) & (!g1406) & (g1407) & (!g1412)) + ((!g1068) & (g1397) & (!g1409) & (g1406) & (!g1407) & (g1412)) + ((!g1068) & (g1397) & (!g1409) & (g1406) & (g1407) & (g1412)) + ((!g1068) & (g1397) & (g1409) & (!g1406) & (!g1407) & (g1412)) + ((!g1068) & (g1397) & (g1409) & (!g1406) & (g1407) & (g1412)) + ((!g1068) & (g1397) & (g1409) & (g1406) & (!g1407) & (!g1412)) + ((!g1068) & (g1397) & (g1409) & (g1406) & (g1407) & (!g1412)) + ((g1068) & (!g1397) & (!g1409) & (!g1406) & (!g1407) & (g1412)) + ((g1068) & (!g1397) & (!g1409) & (!g1406) & (g1407) & (!g1412)) + ((g1068) & (!g1397) & (!g1409) & (g1406) & (!g1407) & (g1412)) + ((g1068) & (!g1397) & (!g1409) & (g1406) & (g1407) & (g1412)) + ((g1068) & (!g1397) & (g1409) & (!g1406) & (!g1407) & (!g1412)) + ((g1068) & (!g1397) & (g1409) & (!g1406) & (g1407) & (g1412)) + ((g1068) & (!g1397) & (g1409) & (g1406) & (!g1407) & (!g1412)) + ((g1068) & (!g1397) & (g1409) & (g1406) & (g1407) & (!g1412)) + ((g1068) & (g1397) & (!g1409) & (!g1406) & (!g1407) & (g1412)) + ((g1068) & (g1397) & (!g1409) & (!g1406) & (g1407) & (g1412)) + ((g1068) & (g1397) & (!g1409) & (g1406) & (!g1407) & (!g1412)) + ((g1068) & (g1397) & (!g1409) & (g1406) & (g1407) & (g1412)) + ((g1068) & (g1397) & (g1409) & (!g1406) & (!g1407) & (!g1412)) + ((g1068) & (g1397) & (g1409) & (!g1406) & (g1407) & (!g1412)) + ((g1068) & (g1397) & (g1409) & (g1406) & (!g1407) & (g1412)) + ((g1068) & (g1397) & (g1409) & (g1406) & (g1407) & (!g1412)));
	assign g1414 = (((!sk[16]) & (!g1397) & (g1406) & (!g1407)) + ((!sk[16]) & (!g1397) & (g1406) & (g1407)) + ((!sk[16]) & (g1397) & (g1406) & (!g1407)) + ((!sk[16]) & (g1397) & (g1406) & (g1407)) + ((sk[16]) & (!g1397) & (!g1406) & (g1407)) + ((sk[16]) & (g1397) & (g1406) & (g1407)));
	assign g1415 = (((g1396) & (!g1389) & (!g1393) & (!g1398) & (!g1400) & (g1405)) + ((g1396) & (!g1389) & (!g1393) & (!g1398) & (g1400) & (!g1405)) + ((g1396) & (!g1389) & (g1393) & (g1398) & (!g1400) & (!g1405)) + ((g1396) & (!g1389) & (g1393) & (g1398) & (g1400) & (g1405)) + ((g1396) & (g1389) & (!g1393) & (g1398) & (!g1400) & (!g1405)) + ((g1396) & (g1389) & (!g1393) & (g1398) & (g1400) & (g1405)) + ((g1396) & (g1389) & (g1393) & (!g1398) & (!g1400) & (!g1405)) + ((g1396) & (g1389) & (g1393) & (!g1398) & (g1400) & (g1405)));
	assign g1416 = (((!g16) & (!g30) & (!g129) & (!sk[18]) & (g287) & (!g228)) + ((!g16) & (!g30) & (!g129) & (!sk[18]) & (g287) & (g228)) + ((!g16) & (!g30) & (!g129) & (sk[18]) & (!g287) & (g228)) + ((!g16) & (!g30) & (g129) & (!sk[18]) & (!g287) & (!g228)) + ((!g16) & (!g30) & (g129) & (!sk[18]) & (!g287) & (g228)) + ((!g16) & (!g30) & (g129) & (!sk[18]) & (g287) & (!g228)) + ((!g16) & (!g30) & (g129) & (!sk[18]) & (g287) & (g228)) + ((!g16) & (g30) & (!g129) & (!sk[18]) & (!g287) & (!g228)) + ((!g16) & (g30) & (!g129) & (!sk[18]) & (!g287) & (g228)) + ((!g16) & (g30) & (!g129) & (!sk[18]) & (g287) & (!g228)) + ((!g16) & (g30) & (!g129) & (!sk[18]) & (g287) & (g228)) + ((!g16) & (g30) & (!g129) & (sk[18]) & (!g287) & (g228)) + ((!g16) & (g30) & (g129) & (!sk[18]) & (!g287) & (!g228)) + ((!g16) & (g30) & (g129) & (!sk[18]) & (!g287) & (g228)) + ((!g16) & (g30) & (g129) & (!sk[18]) & (g287) & (!g228)) + ((!g16) & (g30) & (g129) & (!sk[18]) & (g287) & (g228)) + ((g16) & (!g30) & (!g129) & (!sk[18]) & (g287) & (!g228)) + ((g16) & (!g30) & (!g129) & (!sk[18]) & (g287) & (g228)) + ((g16) & (!g30) & (!g129) & (sk[18]) & (!g287) & (g228)) + ((g16) & (!g30) & (g129) & (!sk[18]) & (!g287) & (!g228)) + ((g16) & (!g30) & (g129) & (!sk[18]) & (!g287) & (g228)) + ((g16) & (!g30) & (g129) & (!sk[18]) & (g287) & (!g228)) + ((g16) & (!g30) & (g129) & (!sk[18]) & (g287) & (g228)) + ((g16) & (g30) & (!g129) & (!sk[18]) & (!g287) & (!g228)) + ((g16) & (g30) & (!g129) & (!sk[18]) & (!g287) & (g228)) + ((g16) & (g30) & (!g129) & (!sk[18]) & (g287) & (!g228)) + ((g16) & (g30) & (!g129) & (!sk[18]) & (g287) & (g228)) + ((g16) & (g30) & (g129) & (!sk[18]) & (!g287) & (!g228)) + ((g16) & (g30) & (g129) & (!sk[18]) & (!g287) & (g228)) + ((g16) & (g30) & (g129) & (!sk[18]) & (g287) & (!g228)) + ((g16) & (g30) & (g129) & (!sk[18]) & (g287) & (g228)));
	assign g1417 = (((!g47) & (!g93) & (g348) & (g349) & (g350) & (g701)));
	assign g1418 = (((g591) & (g224) & (g341) & (g1014) & (g1416) & (g1417)));
	assign g1419 = (((!g1068) & (!g1409) & (!g1414) & (!g1415) & (!g1412) & (g1418)) + ((!g1068) & (!g1409) & (!g1414) & (!g1415) & (g1412) & (g1418)) + ((!g1068) & (!g1409) & (!g1414) & (g1415) & (!g1412) & (!g1418)) + ((!g1068) & (!g1409) & (!g1414) & (g1415) & (g1412) & (g1418)) + ((!g1068) & (!g1409) & (g1414) & (!g1415) & (!g1412) & (g1418)) + ((!g1068) & (!g1409) & (g1414) & (!g1415) & (g1412) & (g1418)) + ((!g1068) & (!g1409) & (g1414) & (g1415) & (!g1412) & (!g1418)) + ((!g1068) & (!g1409) & (g1414) & (g1415) & (g1412) & (g1418)) + ((!g1068) & (g1409) & (!g1414) & (!g1415) & (!g1412) & (!g1418)) + ((!g1068) & (g1409) & (!g1414) & (!g1415) & (g1412) & (g1418)) + ((!g1068) & (g1409) & (!g1414) & (g1415) & (!g1412) & (!g1418)) + ((!g1068) & (g1409) & (!g1414) & (g1415) & (g1412) & (!g1418)) + ((!g1068) & (g1409) & (g1414) & (!g1415) & (!g1412) & (!g1418)) + ((!g1068) & (g1409) & (g1414) & (!g1415) & (g1412) & (g1418)) + ((!g1068) & (g1409) & (g1414) & (g1415) & (!g1412) & (!g1418)) + ((!g1068) & (g1409) & (g1414) & (g1415) & (g1412) & (!g1418)) + ((g1068) & (!g1409) & (!g1414) & (!g1415) & (!g1412) & (!g1418)) + ((g1068) & (!g1409) & (!g1414) & (!g1415) & (g1412) & (!g1418)) + ((g1068) & (!g1409) & (!g1414) & (g1415) & (!g1412) & (g1418)) + ((g1068) & (!g1409) & (!g1414) & (g1415) & (g1412) & (!g1418)) + ((g1068) & (!g1409) & (g1414) & (!g1415) & (!g1412) & (!g1418)) + ((g1068) & (!g1409) & (g1414) & (!g1415) & (g1412) & (g1418)) + ((g1068) & (!g1409) & (g1414) & (g1415) & (!g1412) & (!g1418)) + ((g1068) & (!g1409) & (g1414) & (g1415) & (g1412) & (!g1418)) + ((g1068) & (g1409) & (!g1414) & (!g1415) & (!g1412) & (g1418)) + ((g1068) & (g1409) & (!g1414) & (!g1415) & (g1412) & (!g1418)) + ((g1068) & (g1409) & (!g1414) & (g1415) & (!g1412) & (g1418)) + ((g1068) & (g1409) & (!g1414) & (g1415) & (g1412) & (g1418)) + ((g1068) & (g1409) & (g1414) & (!g1415) & (!g1412) & (!g1418)) + ((g1068) & (g1409) & (g1414) & (!g1415) & (g1412) & (!g1418)) + ((g1068) & (g1409) & (g1414) & (g1415) & (!g1412) & (g1418)) + ((g1068) & (g1409) & (g1414) & (g1415) & (g1412) & (!g1418)));
	assign g1420 = (((!g38) & (!g9) & (!sk[22]) & (!g10) & (g30) & (!g104)) + ((!g38) & (!g9) & (!sk[22]) & (!g10) & (g30) & (g104)) + ((!g38) & (!g9) & (!sk[22]) & (g10) & (!g30) & (!g104)) + ((!g38) & (!g9) & (!sk[22]) & (g10) & (!g30) & (g104)) + ((!g38) & (!g9) & (!sk[22]) & (g10) & (g30) & (!g104)) + ((!g38) & (!g9) & (!sk[22]) & (g10) & (g30) & (g104)) + ((!g38) & (!g9) & (sk[22]) & (!g10) & (!g30) & (!g104)) + ((!g38) & (!g9) & (sk[22]) & (!g10) & (!g30) & (g104)) + ((!g38) & (!g9) & (sk[22]) & (!g10) & (g30) & (!g104)) + ((!g38) & (!g9) & (sk[22]) & (!g10) & (g30) & (g104)) + ((!g38) & (!g9) & (sk[22]) & (g10) & (!g30) & (!g104)) + ((!g38) & (!g9) & (sk[22]) & (g10) & (!g30) & (g104)) + ((!g38) & (!g9) & (sk[22]) & (g10) & (g30) & (!g104)) + ((!g38) & (!g9) & (sk[22]) & (g10) & (g30) & (g104)) + ((!g38) & (g9) & (!sk[22]) & (!g10) & (!g30) & (!g104)) + ((!g38) & (g9) & (!sk[22]) & (!g10) & (!g30) & (g104)) + ((!g38) & (g9) & (!sk[22]) & (!g10) & (g30) & (!g104)) + ((!g38) & (g9) & (!sk[22]) & (!g10) & (g30) & (g104)) + ((!g38) & (g9) & (!sk[22]) & (g10) & (!g30) & (!g104)) + ((!g38) & (g9) & (!sk[22]) & (g10) & (!g30) & (g104)) + ((!g38) & (g9) & (!sk[22]) & (g10) & (g30) & (!g104)) + ((!g38) & (g9) & (!sk[22]) & (g10) & (g30) & (g104)) + ((!g38) & (g9) & (sk[22]) & (!g10) & (!g30) & (!g104)) + ((!g38) & (g9) & (sk[22]) & (!g10) & (!g30) & (g104)) + ((g38) & (!g9) & (!sk[22]) & (!g10) & (g30) & (!g104)) + ((g38) & (!g9) & (!sk[22]) & (!g10) & (g30) & (g104)) + ((g38) & (!g9) & (!sk[22]) & (g10) & (!g30) & (!g104)) + ((g38) & (!g9) & (!sk[22]) & (g10) & (!g30) & (g104)) + ((g38) & (!g9) & (!sk[22]) & (g10) & (g30) & (!g104)) + ((g38) & (!g9) & (!sk[22]) & (g10) & (g30) & (g104)) + ((g38) & (!g9) & (sk[22]) & (!g10) & (!g30) & (!g104)) + ((g38) & (!g9) & (sk[22]) & (!g10) & (g30) & (!g104)) + ((g38) & (!g9) & (sk[22]) & (g10) & (!g30) & (!g104)) + ((g38) & (!g9) & (sk[22]) & (g10) & (g30) & (!g104)) + ((g38) & (g9) & (!sk[22]) & (!g10) & (!g30) & (!g104)) + ((g38) & (g9) & (!sk[22]) & (!g10) & (!g30) & (g104)) + ((g38) & (g9) & (!sk[22]) & (!g10) & (g30) & (!g104)) + ((g38) & (g9) & (!sk[22]) & (!g10) & (g30) & (g104)) + ((g38) & (g9) & (!sk[22]) & (g10) & (!g30) & (!g104)) + ((g38) & (g9) & (!sk[22]) & (g10) & (!g30) & (g104)) + ((g38) & (g9) & (!sk[22]) & (g10) & (g30) & (!g104)) + ((g38) & (g9) & (!sk[22]) & (g10) & (g30) & (g104)) + ((g38) & (g9) & (sk[22]) & (!g10) & (!g30) & (!g104)));
	assign g1421 = (((!g71) & (!g66) & (!g59) & (!g20) & (!g137) & (g1420)) + ((!g71) & (!g66) & (!g59) & (g20) & (!g137) & (g1420)) + ((!g71) & (g66) & (!g59) & (!g20) & (!g137) & (g1420)) + ((!g71) & (g66) & (!g59) & (g20) & (!g137) & (g1420)) + ((g71) & (!g66) & (!g59) & (!g20) & (!g137) & (g1420)));
	assign g1422 = (((!g168) & (!g859) & (!g1250) & (!sk[24]) & (g1390) & (!g1421)) + ((!g168) & (!g859) & (!g1250) & (!sk[24]) & (g1390) & (g1421)) + ((!g168) & (!g859) & (g1250) & (!sk[24]) & (!g1390) & (!g1421)) + ((!g168) & (!g859) & (g1250) & (!sk[24]) & (!g1390) & (g1421)) + ((!g168) & (!g859) & (g1250) & (!sk[24]) & (g1390) & (!g1421)) + ((!g168) & (!g859) & (g1250) & (!sk[24]) & (g1390) & (g1421)) + ((!g168) & (g859) & (!g1250) & (!sk[24]) & (!g1390) & (!g1421)) + ((!g168) & (g859) & (!g1250) & (!sk[24]) & (!g1390) & (g1421)) + ((!g168) & (g859) & (!g1250) & (!sk[24]) & (g1390) & (!g1421)) + ((!g168) & (g859) & (!g1250) & (!sk[24]) & (g1390) & (g1421)) + ((!g168) & (g859) & (g1250) & (!sk[24]) & (!g1390) & (!g1421)) + ((!g168) & (g859) & (g1250) & (!sk[24]) & (!g1390) & (g1421)) + ((!g168) & (g859) & (g1250) & (!sk[24]) & (g1390) & (!g1421)) + ((!g168) & (g859) & (g1250) & (!sk[24]) & (g1390) & (g1421)) + ((g168) & (!g859) & (!g1250) & (!sk[24]) & (g1390) & (!g1421)) + ((g168) & (!g859) & (!g1250) & (!sk[24]) & (g1390) & (g1421)) + ((g168) & (!g859) & (g1250) & (!sk[24]) & (!g1390) & (!g1421)) + ((g168) & (!g859) & (g1250) & (!sk[24]) & (!g1390) & (g1421)) + ((g168) & (!g859) & (g1250) & (!sk[24]) & (g1390) & (!g1421)) + ((g168) & (!g859) & (g1250) & (!sk[24]) & (g1390) & (g1421)) + ((g168) & (g859) & (!g1250) & (!sk[24]) & (!g1390) & (!g1421)) + ((g168) & (g859) & (!g1250) & (!sk[24]) & (!g1390) & (g1421)) + ((g168) & (g859) & (!g1250) & (!sk[24]) & (g1390) & (!g1421)) + ((g168) & (g859) & (!g1250) & (!sk[24]) & (g1390) & (g1421)) + ((g168) & (g859) & (g1250) & (!sk[24]) & (!g1390) & (!g1421)) + ((g168) & (g859) & (g1250) & (!sk[24]) & (!g1390) & (g1421)) + ((g168) & (g859) & (g1250) & (!sk[24]) & (g1390) & (!g1421)) + ((g168) & (g859) & (g1250) & (!sk[24]) & (g1390) & (g1421)) + ((g168) & (g859) & (g1250) & (sk[24]) & (g1390) & (g1421)));
	assign g1423 = (((!g1409) & (!sk[25]) & (!g1415) & (!g1412) & (g1418) & (!g1422)) + ((!g1409) & (!sk[25]) & (!g1415) & (!g1412) & (g1418) & (g1422)) + ((!g1409) & (!sk[25]) & (!g1415) & (g1412) & (!g1418) & (!g1422)) + ((!g1409) & (!sk[25]) & (!g1415) & (g1412) & (!g1418) & (g1422)) + ((!g1409) & (!sk[25]) & (!g1415) & (g1412) & (g1418) & (!g1422)) + ((!g1409) & (!sk[25]) & (!g1415) & (g1412) & (g1418) & (g1422)) + ((!g1409) & (!sk[25]) & (g1415) & (!g1412) & (!g1418) & (!g1422)) + ((!g1409) & (!sk[25]) & (g1415) & (!g1412) & (!g1418) & (g1422)) + ((!g1409) & (!sk[25]) & (g1415) & (!g1412) & (g1418) & (!g1422)) + ((!g1409) & (!sk[25]) & (g1415) & (!g1412) & (g1418) & (g1422)) + ((!g1409) & (!sk[25]) & (g1415) & (g1412) & (!g1418) & (!g1422)) + ((!g1409) & (!sk[25]) & (g1415) & (g1412) & (!g1418) & (g1422)) + ((!g1409) & (!sk[25]) & (g1415) & (g1412) & (g1418) & (!g1422)) + ((!g1409) & (!sk[25]) & (g1415) & (g1412) & (g1418) & (g1422)) + ((!g1409) & (sk[25]) & (!g1415) & (!g1412) & (!g1418) & (!g1422)) + ((!g1409) & (sk[25]) & (!g1415) & (!g1412) & (g1418) & (!g1422)) + ((!g1409) & (sk[25]) & (!g1415) & (g1412) & (!g1418) & (!g1422)) + ((!g1409) & (sk[25]) & (!g1415) & (g1412) & (g1418) & (!g1422)) + ((!g1409) & (sk[25]) & (g1415) & (!g1412) & (!g1418) & (g1422)) + ((!g1409) & (sk[25]) & (g1415) & (!g1412) & (g1418) & (!g1422)) + ((!g1409) & (sk[25]) & (g1415) & (g1412) & (!g1418) & (!g1422)) + ((!g1409) & (sk[25]) & (g1415) & (g1412) & (g1418) & (!g1422)) + ((g1409) & (!sk[25]) & (!g1415) & (!g1412) & (g1418) & (!g1422)) + ((g1409) & (!sk[25]) & (!g1415) & (!g1412) & (g1418) & (g1422)) + ((g1409) & (!sk[25]) & (!g1415) & (g1412) & (!g1418) & (!g1422)) + ((g1409) & (!sk[25]) & (!g1415) & (g1412) & (!g1418) & (g1422)) + ((g1409) & (!sk[25]) & (!g1415) & (g1412) & (g1418) & (!g1422)) + ((g1409) & (!sk[25]) & (!g1415) & (g1412) & (g1418) & (g1422)) + ((g1409) & (!sk[25]) & (g1415) & (!g1412) & (!g1418) & (!g1422)) + ((g1409) & (!sk[25]) & (g1415) & (!g1412) & (!g1418) & (g1422)) + ((g1409) & (!sk[25]) & (g1415) & (!g1412) & (g1418) & (!g1422)) + ((g1409) & (!sk[25]) & (g1415) & (!g1412) & (g1418) & (g1422)) + ((g1409) & (!sk[25]) & (g1415) & (g1412) & (!g1418) & (!g1422)) + ((g1409) & (!sk[25]) & (g1415) & (g1412) & (!g1418) & (g1422)) + ((g1409) & (!sk[25]) & (g1415) & (g1412) & (g1418) & (!g1422)) + ((g1409) & (!sk[25]) & (g1415) & (g1412) & (g1418) & (g1422)) + ((g1409) & (sk[25]) & (!g1415) & (!g1412) & (!g1418) & (g1422)) + ((g1409) & (sk[25]) & (!g1415) & (!g1412) & (g1418) & (!g1422)) + ((g1409) & (sk[25]) & (!g1415) & (g1412) & (!g1418) & (!g1422)) + ((g1409) & (sk[25]) & (!g1415) & (g1412) & (g1418) & (!g1422)) + ((g1409) & (sk[25]) & (g1415) & (!g1412) & (!g1418) & (g1422)) + ((g1409) & (sk[25]) & (g1415) & (!g1412) & (g1418) & (!g1422)) + ((g1409) & (sk[25]) & (g1415) & (g1412) & (!g1418) & (g1422)) + ((g1409) & (sk[25]) & (g1415) & (g1412) & (g1418) & (!g1422)));
	assign g1424 = (((!g1397) & (!g1409) & (!g1406) & (g1407) & (g1412) & (g1418)) + ((!g1397) & (g1409) & (!g1406) & (g1407) & (!g1412) & (!g1418)) + ((g1397) & (!g1409) & (g1406) & (g1407) & (!g1412) & (!g1418)) + ((g1397) & (g1409) & (g1406) & (g1407) & (g1412) & (!g1418)));
	assign sinx19x = (((!g1068) & (g1423) & (!sk[27]) & (!g1424)) + ((!g1068) & (g1423) & (!sk[27]) & (g1424)) + ((!g1068) & (g1423) & (sk[27]) & (!g1424)) + ((!g1068) & (g1423) & (sk[27]) & (g1424)) + ((g1068) & (!g1423) & (sk[27]) & (!g1424)) + ((g1068) & (g1423) & (!sk[27]) & (!g1424)) + ((g1068) & (g1423) & (!sk[27]) & (g1424)) + ((g1068) & (g1423) & (sk[27]) & (g1424)));
	assign g1426 = (((!g593) & (!g1006) & (!g35) & (!sk[28]) & (g587)) + ((!g593) & (!g1006) & (g35) & (!sk[28]) & (g587)) + ((!g593) & (g1006) & (!g35) & (!sk[28]) & (g587)) + ((!g593) & (g1006) & (!g35) & (sk[28]) & (!g587)) + ((!g593) & (g1006) & (g35) & (!sk[28]) & (g587)) + ((g593) & (!g1006) & (!g35) & (!sk[28]) & (!g587)) + ((g593) & (!g1006) & (!g35) & (!sk[28]) & (g587)) + ((g593) & (!g1006) & (g35) & (!sk[28]) & (!g587)) + ((g593) & (!g1006) & (g35) & (!sk[28]) & (g587)) + ((g593) & (g1006) & (!g35) & (!sk[28]) & (!g587)) + ((g593) & (g1006) & (!g35) & (!sk[28]) & (g587)) + ((g593) & (g1006) & (g35) & (!sk[28]) & (!g587)) + ((g593) & (g1006) & (g35) & (!sk[28]) & (g587)));
	assign g1427 = (((!g112) & (!g113) & (!g97) & (!g98) & (!g62) & (g46)) + ((!g112) & (!g113) & (!g97) & (!g98) & (g62) & (g46)) + ((!g112) & (!g113) & (!g97) & (g98) & (g62) & (!g46)) + ((!g112) & (!g113) & (!g97) & (g98) & (g62) & (g46)) + ((!g112) & (!g113) & (g97) & (!g98) & (g62) & (!g46)) + ((!g112) & (!g113) & (g97) & (!g98) & (g62) & (g46)) + ((g112) & (g113) & (g97) & (g98) & (!g62) & (g46)) + ((g112) & (g113) & (g97) & (g98) & (g62) & (g46)));
	assign g1428 = (((!g85) & (!g236) & (!sk[30]) & (!g87) & (g965) & (!g1427)) + ((!g85) & (!g236) & (!sk[30]) & (!g87) & (g965) & (g1427)) + ((!g85) & (!g236) & (!sk[30]) & (g87) & (!g965) & (!g1427)) + ((!g85) & (!g236) & (!sk[30]) & (g87) & (!g965) & (g1427)) + ((!g85) & (!g236) & (!sk[30]) & (g87) & (g965) & (!g1427)) + ((!g85) & (!g236) & (!sk[30]) & (g87) & (g965) & (g1427)) + ((!g85) & (!g236) & (sk[30]) & (!g87) & (g965) & (!g1427)) + ((!g85) & (g236) & (!sk[30]) & (!g87) & (!g965) & (!g1427)) + ((!g85) & (g236) & (!sk[30]) & (!g87) & (!g965) & (g1427)) + ((!g85) & (g236) & (!sk[30]) & (!g87) & (g965) & (!g1427)) + ((!g85) & (g236) & (!sk[30]) & (!g87) & (g965) & (g1427)) + ((!g85) & (g236) & (!sk[30]) & (g87) & (!g965) & (!g1427)) + ((!g85) & (g236) & (!sk[30]) & (g87) & (!g965) & (g1427)) + ((!g85) & (g236) & (!sk[30]) & (g87) & (g965) & (!g1427)) + ((!g85) & (g236) & (!sk[30]) & (g87) & (g965) & (g1427)) + ((g85) & (!g236) & (!sk[30]) & (!g87) & (g965) & (!g1427)) + ((g85) & (!g236) & (!sk[30]) & (!g87) & (g965) & (g1427)) + ((g85) & (!g236) & (!sk[30]) & (g87) & (!g965) & (!g1427)) + ((g85) & (!g236) & (!sk[30]) & (g87) & (!g965) & (g1427)) + ((g85) & (!g236) & (!sk[30]) & (g87) & (g965) & (!g1427)) + ((g85) & (!g236) & (!sk[30]) & (g87) & (g965) & (g1427)) + ((g85) & (g236) & (!sk[30]) & (!g87) & (!g965) & (!g1427)) + ((g85) & (g236) & (!sk[30]) & (!g87) & (!g965) & (g1427)) + ((g85) & (g236) & (!sk[30]) & (!g87) & (g965) & (!g1427)) + ((g85) & (g236) & (!sk[30]) & (!g87) & (g965) & (g1427)) + ((g85) & (g236) & (!sk[30]) & (g87) & (!g965) & (!g1427)) + ((g85) & (g236) & (!sk[30]) & (g87) & (!g965) & (g1427)) + ((g85) & (g236) & (!sk[30]) & (g87) & (g965) & (!g1427)) + ((g85) & (g236) & (!sk[30]) & (g87) & (g965) & (g1427)));
	assign g1429 = (((!g599) & (!g136) & (!g1273) & (!sk[31]) & (g1426) & (!g1428)) + ((!g599) & (!g136) & (!g1273) & (!sk[31]) & (g1426) & (g1428)) + ((!g599) & (!g136) & (g1273) & (!sk[31]) & (!g1426) & (!g1428)) + ((!g599) & (!g136) & (g1273) & (!sk[31]) & (!g1426) & (g1428)) + ((!g599) & (!g136) & (g1273) & (!sk[31]) & (g1426) & (!g1428)) + ((!g599) & (!g136) & (g1273) & (!sk[31]) & (g1426) & (g1428)) + ((!g599) & (g136) & (!g1273) & (!sk[31]) & (!g1426) & (!g1428)) + ((!g599) & (g136) & (!g1273) & (!sk[31]) & (!g1426) & (g1428)) + ((!g599) & (g136) & (!g1273) & (!sk[31]) & (g1426) & (!g1428)) + ((!g599) & (g136) & (!g1273) & (!sk[31]) & (g1426) & (g1428)) + ((!g599) & (g136) & (g1273) & (!sk[31]) & (!g1426) & (!g1428)) + ((!g599) & (g136) & (g1273) & (!sk[31]) & (!g1426) & (g1428)) + ((!g599) & (g136) & (g1273) & (!sk[31]) & (g1426) & (!g1428)) + ((!g599) & (g136) & (g1273) & (!sk[31]) & (g1426) & (g1428)) + ((g599) & (!g136) & (!g1273) & (!sk[31]) & (g1426) & (!g1428)) + ((g599) & (!g136) & (!g1273) & (!sk[31]) & (g1426) & (g1428)) + ((g599) & (!g136) & (g1273) & (!sk[31]) & (!g1426) & (!g1428)) + ((g599) & (!g136) & (g1273) & (!sk[31]) & (!g1426) & (g1428)) + ((g599) & (!g136) & (g1273) & (!sk[31]) & (g1426) & (!g1428)) + ((g599) & (!g136) & (g1273) & (!sk[31]) & (g1426) & (g1428)) + ((g599) & (g136) & (!g1273) & (!sk[31]) & (!g1426) & (!g1428)) + ((g599) & (g136) & (!g1273) & (!sk[31]) & (!g1426) & (g1428)) + ((g599) & (g136) & (!g1273) & (!sk[31]) & (g1426) & (!g1428)) + ((g599) & (g136) & (!g1273) & (!sk[31]) & (g1426) & (g1428)) + ((g599) & (g136) & (g1273) & (!sk[31]) & (!g1426) & (!g1428)) + ((g599) & (g136) & (g1273) & (!sk[31]) & (!g1426) & (g1428)) + ((g599) & (g136) & (g1273) & (!sk[31]) & (g1426) & (!g1428)) + ((g599) & (g136) & (g1273) & (!sk[31]) & (g1426) & (g1428)) + ((g599) & (g136) & (g1273) & (sk[31]) & (g1426) & (g1428)));
	assign g1430 = (((!g1409) & (!g1415) & (!g1412) & (!g1418) & (!g1422) & (g1429)) + ((!g1409) & (!g1415) & (!g1412) & (!g1418) & (g1422) & (g1429)) + ((!g1409) & (!g1415) & (!g1412) & (g1418) & (!g1422) & (g1429)) + ((!g1409) & (!g1415) & (!g1412) & (g1418) & (g1422) & (g1429)) + ((!g1409) & (!g1415) & (g1412) & (!g1418) & (!g1422) & (g1429)) + ((!g1409) & (!g1415) & (g1412) & (!g1418) & (g1422) & (g1429)) + ((!g1409) & (!g1415) & (g1412) & (g1418) & (!g1422) & (g1429)) + ((!g1409) & (!g1415) & (g1412) & (g1418) & (g1422) & (g1429)) + ((!g1409) & (g1415) & (!g1412) & (!g1418) & (!g1422) & (!g1429)) + ((!g1409) & (g1415) & (!g1412) & (!g1418) & (g1422) & (g1429)) + ((!g1409) & (g1415) & (!g1412) & (g1418) & (!g1422) & (g1429)) + ((!g1409) & (g1415) & (!g1412) & (g1418) & (g1422) & (g1429)) + ((!g1409) & (g1415) & (g1412) & (!g1418) & (!g1422) & (g1429)) + ((!g1409) & (g1415) & (g1412) & (!g1418) & (g1422) & (g1429)) + ((!g1409) & (g1415) & (g1412) & (g1418) & (!g1422) & (g1429)) + ((!g1409) & (g1415) & (g1412) & (g1418) & (g1422) & (g1429)) + ((g1409) & (!g1415) & (!g1412) & (!g1418) & (!g1422) & (!g1429)) + ((g1409) & (!g1415) & (!g1412) & (!g1418) & (g1422) & (g1429)) + ((g1409) & (!g1415) & (!g1412) & (g1418) & (!g1422) & (g1429)) + ((g1409) & (!g1415) & (!g1412) & (g1418) & (g1422) & (g1429)) + ((g1409) & (!g1415) & (g1412) & (!g1418) & (!g1422) & (g1429)) + ((g1409) & (!g1415) & (g1412) & (!g1418) & (g1422) & (g1429)) + ((g1409) & (!g1415) & (g1412) & (g1418) & (!g1422) & (g1429)) + ((g1409) & (!g1415) & (g1412) & (g1418) & (g1422) & (g1429)) + ((g1409) & (g1415) & (!g1412) & (!g1418) & (!g1422) & (!g1429)) + ((g1409) & (g1415) & (!g1412) & (!g1418) & (g1422) & (g1429)) + ((g1409) & (g1415) & (!g1412) & (g1418) & (!g1422) & (g1429)) + ((g1409) & (g1415) & (!g1412) & (g1418) & (g1422) & (g1429)) + ((g1409) & (g1415) & (g1412) & (!g1418) & (!g1422) & (!g1429)) + ((g1409) & (g1415) & (g1412) & (!g1418) & (g1422) & (g1429)) + ((g1409) & (g1415) & (g1412) & (g1418) & (!g1422) & (g1429)) + ((g1409) & (g1415) & (g1412) & (g1418) & (g1422) & (g1429)));
	assign g1431 = (((!g1068) & (!g1423) & (!g1424) & (!sk[33]) & (g1430)) + ((!g1068) & (!g1423) & (!g1424) & (sk[33]) & (g1430)) + ((!g1068) & (!g1423) & (g1424) & (!sk[33]) & (g1430)) + ((!g1068) & (!g1423) & (g1424) & (sk[33]) & (g1430)) + ((!g1068) & (g1423) & (!g1424) & (!sk[33]) & (g1430)) + ((!g1068) & (g1423) & (!g1424) & (sk[33]) & (g1430)) + ((!g1068) & (g1423) & (g1424) & (!sk[33]) & (g1430)) + ((!g1068) & (g1423) & (g1424) & (sk[33]) & (g1430)) + ((g1068) & (!g1423) & (!g1424) & (!sk[33]) & (!g1430)) + ((g1068) & (!g1423) & (!g1424) & (!sk[33]) & (g1430)) + ((g1068) & (!g1423) & (!g1424) & (sk[33]) & (!g1430)) + ((g1068) & (!g1423) & (g1424) & (!sk[33]) & (!g1430)) + ((g1068) & (!g1423) & (g1424) & (!sk[33]) & (g1430)) + ((g1068) & (!g1423) & (g1424) & (sk[33]) & (g1430)) + ((g1068) & (g1423) & (!g1424) & (!sk[33]) & (!g1430)) + ((g1068) & (g1423) & (!g1424) & (!sk[33]) & (g1430)) + ((g1068) & (g1423) & (!g1424) & (sk[33]) & (!g1430)) + ((g1068) & (g1423) & (g1424) & (!sk[33]) & (!g1430)) + ((g1068) & (g1423) & (g1424) & (!sk[33]) & (g1430)) + ((g1068) & (g1423) & (g1424) & (sk[33]) & (!g1430)));
	assign g1432 = (((!g1409) & (g1415) & (!g1412) & (!g1418) & (!g1422) & (!g1429)) + ((g1409) & (g1415) & (g1412) & (!g1418) & (!g1422) & (!g1429)));
	assign g1433 = (((!g10) & (!g62) & (!g46) & (!sk[35]) & (g27)) + ((!g10) & (!g62) & (g46) & (!sk[35]) & (g27)) + ((!g10) & (!g62) & (g46) & (sk[35]) & (g27)) + ((!g10) & (g62) & (!g46) & (!sk[35]) & (g27)) + ((!g10) & (g62) & (!g46) & (sk[35]) & (g27)) + ((!g10) & (g62) & (g46) & (!sk[35]) & (g27)) + ((!g10) & (g62) & (g46) & (sk[35]) & (g27)) + ((g10) & (!g62) & (!g46) & (!sk[35]) & (!g27)) + ((g10) & (!g62) & (!g46) & (!sk[35]) & (g27)) + ((g10) & (!g62) & (g46) & (!sk[35]) & (!g27)) + ((g10) & (!g62) & (g46) & (!sk[35]) & (g27)) + ((g10) & (!g62) & (g46) & (sk[35]) & (!g27)) + ((g10) & (!g62) & (g46) & (sk[35]) & (g27)) + ((g10) & (g62) & (!g46) & (!sk[35]) & (!g27)) + ((g10) & (g62) & (!g46) & (!sk[35]) & (g27)) + ((g10) & (g62) & (!g46) & (sk[35]) & (g27)) + ((g10) & (g62) & (g46) & (!sk[35]) & (!g27)) + ((g10) & (g62) & (g46) & (!sk[35]) & (g27)) + ((g10) & (g62) & (g46) & (sk[35]) & (!g27)) + ((g10) & (g62) & (g46) & (sk[35]) & (g27)));
	assign g1434 = (((!sk[36]) & (!g69) & (!g885) & (!g213) & (g216) & (!g1433)) + ((!sk[36]) & (!g69) & (!g885) & (!g213) & (g216) & (g1433)) + ((!sk[36]) & (!g69) & (!g885) & (g213) & (!g216) & (!g1433)) + ((!sk[36]) & (!g69) & (!g885) & (g213) & (!g216) & (g1433)) + ((!sk[36]) & (!g69) & (!g885) & (g213) & (g216) & (!g1433)) + ((!sk[36]) & (!g69) & (!g885) & (g213) & (g216) & (g1433)) + ((!sk[36]) & (!g69) & (g885) & (!g213) & (!g216) & (!g1433)) + ((!sk[36]) & (!g69) & (g885) & (!g213) & (!g216) & (g1433)) + ((!sk[36]) & (!g69) & (g885) & (!g213) & (g216) & (!g1433)) + ((!sk[36]) & (!g69) & (g885) & (!g213) & (g216) & (g1433)) + ((!sk[36]) & (!g69) & (g885) & (g213) & (!g216) & (!g1433)) + ((!sk[36]) & (!g69) & (g885) & (g213) & (!g216) & (g1433)) + ((!sk[36]) & (!g69) & (g885) & (g213) & (g216) & (!g1433)) + ((!sk[36]) & (!g69) & (g885) & (g213) & (g216) & (g1433)) + ((!sk[36]) & (g69) & (!g885) & (!g213) & (g216) & (!g1433)) + ((!sk[36]) & (g69) & (!g885) & (!g213) & (g216) & (g1433)) + ((!sk[36]) & (g69) & (!g885) & (g213) & (!g216) & (!g1433)) + ((!sk[36]) & (g69) & (!g885) & (g213) & (!g216) & (g1433)) + ((!sk[36]) & (g69) & (!g885) & (g213) & (g216) & (!g1433)) + ((!sk[36]) & (g69) & (!g885) & (g213) & (g216) & (g1433)) + ((!sk[36]) & (g69) & (g885) & (!g213) & (!g216) & (!g1433)) + ((!sk[36]) & (g69) & (g885) & (!g213) & (!g216) & (g1433)) + ((!sk[36]) & (g69) & (g885) & (!g213) & (g216) & (!g1433)) + ((!sk[36]) & (g69) & (g885) & (!g213) & (g216) & (g1433)) + ((!sk[36]) & (g69) & (g885) & (g213) & (!g216) & (!g1433)) + ((!sk[36]) & (g69) & (g885) & (g213) & (!g216) & (g1433)) + ((!sk[36]) & (g69) & (g885) & (g213) & (g216) & (!g1433)) + ((!sk[36]) & (g69) & (g885) & (g213) & (g216) & (g1433)) + ((sk[36]) & (g69) & (g885) & (g213) & (!g216) & (!g1433)));
	assign g1435 = (((!g1409) & (!g1412) & (!g1418) & (!g1422) & (!g1429) & (!g1434)) + ((!g1409) & (!g1412) & (!g1418) & (!g1422) & (g1429) & (!g1434)) + ((!g1409) & (!g1412) & (!g1418) & (g1422) & (!g1429) & (!g1434)) + ((!g1409) & (!g1412) & (!g1418) & (g1422) & (g1429) & (!g1434)) + ((!g1409) & (!g1412) & (g1418) & (!g1422) & (!g1429) & (!g1434)) + ((!g1409) & (!g1412) & (g1418) & (!g1422) & (g1429) & (!g1434)) + ((!g1409) & (!g1412) & (g1418) & (g1422) & (!g1429) & (!g1434)) + ((!g1409) & (!g1412) & (g1418) & (g1422) & (g1429) & (!g1434)) + ((!g1409) & (g1412) & (!g1418) & (!g1422) & (!g1429) & (!g1434)) + ((!g1409) & (g1412) & (!g1418) & (!g1422) & (g1429) & (!g1434)) + ((!g1409) & (g1412) & (!g1418) & (g1422) & (!g1429) & (!g1434)) + ((!g1409) & (g1412) & (!g1418) & (g1422) & (g1429) & (!g1434)) + ((!g1409) & (g1412) & (g1418) & (!g1422) & (!g1429) & (!g1434)) + ((!g1409) & (g1412) & (g1418) & (!g1422) & (g1429) & (!g1434)) + ((!g1409) & (g1412) & (g1418) & (g1422) & (!g1429) & (!g1434)) + ((!g1409) & (g1412) & (g1418) & (g1422) & (g1429) & (!g1434)) + ((g1409) & (!g1412) & (!g1418) & (!g1422) & (!g1429) & (g1434)) + ((g1409) & (!g1412) & (!g1418) & (!g1422) & (g1429) & (!g1434)) + ((g1409) & (!g1412) & (!g1418) & (g1422) & (!g1429) & (!g1434)) + ((g1409) & (!g1412) & (!g1418) & (g1422) & (g1429) & (!g1434)) + ((g1409) & (!g1412) & (g1418) & (!g1422) & (!g1429) & (!g1434)) + ((g1409) & (!g1412) & (g1418) & (!g1422) & (g1429) & (!g1434)) + ((g1409) & (!g1412) & (g1418) & (g1422) & (!g1429) & (!g1434)) + ((g1409) & (!g1412) & (g1418) & (g1422) & (g1429) & (!g1434)) + ((g1409) & (g1412) & (!g1418) & (!g1422) & (!g1429) & (!g1434)) + ((g1409) & (g1412) & (!g1418) & (!g1422) & (g1429) & (!g1434)) + ((g1409) & (g1412) & (!g1418) & (g1422) & (!g1429) & (!g1434)) + ((g1409) & (g1412) & (!g1418) & (g1422) & (g1429) & (!g1434)) + ((g1409) & (g1412) & (g1418) & (!g1422) & (!g1429) & (!g1434)) + ((g1409) & (g1412) & (g1418) & (!g1422) & (g1429) & (!g1434)) + ((g1409) & (g1412) & (g1418) & (g1422) & (!g1429) & (!g1434)) + ((g1409) & (g1412) & (g1418) & (g1422) & (g1429) & (!g1434)));
	assign sinx21x = (((!g1068) & (!g1423) & (!g1424) & (!g1432) & (!g1430) & (g1435)) + ((!g1068) & (!g1423) & (!g1424) & (!g1432) & (g1430) & (g1435)) + ((!g1068) & (!g1423) & (!g1424) & (g1432) & (!g1430) & (!g1435)) + ((!g1068) & (!g1423) & (!g1424) & (g1432) & (g1430) & (!g1435)) + ((!g1068) & (!g1423) & (g1424) & (!g1432) & (!g1430) & (g1435)) + ((!g1068) & (!g1423) & (g1424) & (!g1432) & (g1430) & (g1435)) + ((!g1068) & (!g1423) & (g1424) & (g1432) & (!g1430) & (!g1435)) + ((!g1068) & (!g1423) & (g1424) & (g1432) & (g1430) & (!g1435)) + ((!g1068) & (g1423) & (!g1424) & (!g1432) & (!g1430) & (g1435)) + ((!g1068) & (g1423) & (!g1424) & (!g1432) & (g1430) & (g1435)) + ((!g1068) & (g1423) & (!g1424) & (g1432) & (!g1430) & (!g1435)) + ((!g1068) & (g1423) & (!g1424) & (g1432) & (g1430) & (!g1435)) + ((!g1068) & (g1423) & (g1424) & (!g1432) & (!g1430) & (g1435)) + ((!g1068) & (g1423) & (g1424) & (!g1432) & (g1430) & (g1435)) + ((!g1068) & (g1423) & (g1424) & (g1432) & (!g1430) & (!g1435)) + ((!g1068) & (g1423) & (g1424) & (g1432) & (g1430) & (!g1435)) + ((g1068) & (!g1423) & (!g1424) & (!g1432) & (!g1430) & (!g1435)) + ((g1068) & (!g1423) & (!g1424) & (!g1432) & (g1430) & (!g1435)) + ((g1068) & (!g1423) & (!g1424) & (g1432) & (!g1430) & (g1435)) + ((g1068) & (!g1423) & (!g1424) & (g1432) & (g1430) & (g1435)) + ((g1068) & (!g1423) & (g1424) & (!g1432) & (!g1430) & (!g1435)) + ((g1068) & (!g1423) & (g1424) & (!g1432) & (g1430) & (g1435)) + ((g1068) & (!g1423) & (g1424) & (g1432) & (!g1430) & (g1435)) + ((g1068) & (!g1423) & (g1424) & (g1432) & (g1430) & (!g1435)) + ((g1068) & (g1423) & (!g1424) & (!g1432) & (!g1430) & (!g1435)) + ((g1068) & (g1423) & (!g1424) & (!g1432) & (g1430) & (!g1435)) + ((g1068) & (g1423) & (!g1424) & (g1432) & (!g1430) & (g1435)) + ((g1068) & (g1423) & (!g1424) & (g1432) & (g1430) & (g1435)) + ((g1068) & (g1423) & (g1424) & (!g1432) & (!g1430) & (!g1435)) + ((g1068) & (g1423) & (g1424) & (!g1432) & (g1430) & (!g1435)) + ((g1068) & (g1423) & (g1424) & (g1432) & (!g1430) & (g1435)) + ((g1068) & (g1423) & (g1424) & (g1432) & (g1430) & (g1435)));
	assign g1437 = (((!g1409) & (!g1412) & (!g1418) & (g1422) & (!sk[39]) & (!g1429)) + ((!g1409) & (!g1412) & (!g1418) & (g1422) & (!sk[39]) & (g1429)) + ((!g1409) & (!g1412) & (g1418) & (!g1422) & (!sk[39]) & (!g1429)) + ((!g1409) & (!g1412) & (g1418) & (!g1422) & (!sk[39]) & (g1429)) + ((!g1409) & (!g1412) & (g1418) & (g1422) & (!sk[39]) & (!g1429)) + ((!g1409) & (!g1412) & (g1418) & (g1422) & (!sk[39]) & (g1429)) + ((!g1409) & (g1412) & (!g1418) & (!g1422) & (!sk[39]) & (!g1429)) + ((!g1409) & (g1412) & (!g1418) & (!g1422) & (!sk[39]) & (g1429)) + ((!g1409) & (g1412) & (!g1418) & (g1422) & (!sk[39]) & (!g1429)) + ((!g1409) & (g1412) & (!g1418) & (g1422) & (!sk[39]) & (g1429)) + ((!g1409) & (g1412) & (g1418) & (!g1422) & (!sk[39]) & (!g1429)) + ((!g1409) & (g1412) & (g1418) & (!g1422) & (!sk[39]) & (g1429)) + ((!g1409) & (g1412) & (g1418) & (g1422) & (!sk[39]) & (!g1429)) + ((!g1409) & (g1412) & (g1418) & (g1422) & (!sk[39]) & (g1429)) + ((g1409) & (!g1412) & (!g1418) & (!g1422) & (sk[39]) & (!g1429)) + ((g1409) & (!g1412) & (!g1418) & (g1422) & (!sk[39]) & (!g1429)) + ((g1409) & (!g1412) & (!g1418) & (g1422) & (!sk[39]) & (g1429)) + ((g1409) & (!g1412) & (g1418) & (!g1422) & (!sk[39]) & (!g1429)) + ((g1409) & (!g1412) & (g1418) & (!g1422) & (!sk[39]) & (g1429)) + ((g1409) & (!g1412) & (g1418) & (g1422) & (!sk[39]) & (!g1429)) + ((g1409) & (!g1412) & (g1418) & (g1422) & (!sk[39]) & (g1429)) + ((g1409) & (g1412) & (!g1418) & (!g1422) & (!sk[39]) & (!g1429)) + ((g1409) & (g1412) & (!g1418) & (!g1422) & (!sk[39]) & (g1429)) + ((g1409) & (g1412) & (!g1418) & (g1422) & (!sk[39]) & (!g1429)) + ((g1409) & (g1412) & (!g1418) & (g1422) & (!sk[39]) & (g1429)) + ((g1409) & (g1412) & (g1418) & (!g1422) & (!sk[39]) & (!g1429)) + ((g1409) & (g1412) & (g1418) & (!g1422) & (!sk[39]) & (g1429)) + ((g1409) & (g1412) & (g1418) & (g1422) & (!sk[39]) & (!g1429)) + ((g1409) & (g1412) & (g1418) & (g1422) & (!sk[39]) & (g1429)));
	assign g1438 = (((!g69) & (g209) & (!sk[40]) & (!g219)) + ((!g69) & (g209) & (!sk[40]) & (g219)) + ((g69) & (g209) & (!sk[40]) & (!g219)) + ((g69) & (g209) & (!sk[40]) & (g219)) + ((g69) & (g209) & (sk[40]) & (g219)));
	assign g1439 = (((!g1432) & (!g1437) & (!g1434) & (!sk[41]) & (g1438)) + ((!g1432) & (!g1437) & (!g1434) & (sk[41]) & (g1438)) + ((!g1432) & (!g1437) & (g1434) & (!sk[41]) & (g1438)) + ((!g1432) & (!g1437) & (g1434) & (sk[41]) & (g1438)) + ((!g1432) & (g1437) & (!g1434) & (!sk[41]) & (g1438)) + ((!g1432) & (g1437) & (!g1434) & (sk[41]) & (!g1438)) + ((!g1432) & (g1437) & (g1434) & (!sk[41]) & (g1438)) + ((!g1432) & (g1437) & (g1434) & (sk[41]) & (g1438)) + ((g1432) & (!g1437) & (!g1434) & (!sk[41]) & (!g1438)) + ((g1432) & (!g1437) & (!g1434) & (!sk[41]) & (g1438)) + ((g1432) & (!g1437) & (!g1434) & (sk[41]) & (!g1438)) + ((g1432) & (!g1437) & (g1434) & (!sk[41]) & (!g1438)) + ((g1432) & (!g1437) & (g1434) & (!sk[41]) & (g1438)) + ((g1432) & (!g1437) & (g1434) & (sk[41]) & (g1438)) + ((g1432) & (g1437) & (!g1434) & (!sk[41]) & (!g1438)) + ((g1432) & (g1437) & (!g1434) & (!sk[41]) & (g1438)) + ((g1432) & (g1437) & (!g1434) & (sk[41]) & (!g1438)) + ((g1432) & (g1437) & (g1434) & (!sk[41]) & (!g1438)) + ((g1432) & (g1437) & (g1434) & (!sk[41]) & (g1438)) + ((g1432) & (g1437) & (g1434) & (sk[41]) & (!g1438)));
	assign g1440 = (((!g1423) & (!sk[42]) & (!g1424) & (!g1432) & (g1430) & (!g1435)) + ((!g1423) & (!sk[42]) & (!g1424) & (!g1432) & (g1430) & (g1435)) + ((!g1423) & (!sk[42]) & (!g1424) & (g1432) & (!g1430) & (!g1435)) + ((!g1423) & (!sk[42]) & (!g1424) & (g1432) & (!g1430) & (g1435)) + ((!g1423) & (!sk[42]) & (!g1424) & (g1432) & (g1430) & (!g1435)) + ((!g1423) & (!sk[42]) & (!g1424) & (g1432) & (g1430) & (g1435)) + ((!g1423) & (!sk[42]) & (g1424) & (!g1432) & (!g1430) & (!g1435)) + ((!g1423) & (!sk[42]) & (g1424) & (!g1432) & (!g1430) & (g1435)) + ((!g1423) & (!sk[42]) & (g1424) & (!g1432) & (g1430) & (!g1435)) + ((!g1423) & (!sk[42]) & (g1424) & (!g1432) & (g1430) & (g1435)) + ((!g1423) & (!sk[42]) & (g1424) & (g1432) & (!g1430) & (!g1435)) + ((!g1423) & (!sk[42]) & (g1424) & (g1432) & (!g1430) & (g1435)) + ((!g1423) & (!sk[42]) & (g1424) & (g1432) & (g1430) & (!g1435)) + ((!g1423) & (!sk[42]) & (g1424) & (g1432) & (g1430) & (g1435)) + ((!g1423) & (sk[42]) & (g1424) & (!g1432) & (g1430) & (!g1435)) + ((!g1423) & (sk[42]) & (g1424) & (g1432) & (g1430) & (g1435)) + ((g1423) & (!sk[42]) & (!g1424) & (!g1432) & (g1430) & (!g1435)) + ((g1423) & (!sk[42]) & (!g1424) & (!g1432) & (g1430) & (g1435)) + ((g1423) & (!sk[42]) & (!g1424) & (g1432) & (!g1430) & (!g1435)) + ((g1423) & (!sk[42]) & (!g1424) & (g1432) & (!g1430) & (g1435)) + ((g1423) & (!sk[42]) & (!g1424) & (g1432) & (g1430) & (!g1435)) + ((g1423) & (!sk[42]) & (!g1424) & (g1432) & (g1430) & (g1435)) + ((g1423) & (!sk[42]) & (g1424) & (!g1432) & (!g1430) & (!g1435)) + ((g1423) & (!sk[42]) & (g1424) & (!g1432) & (!g1430) & (g1435)) + ((g1423) & (!sk[42]) & (g1424) & (!g1432) & (g1430) & (!g1435)) + ((g1423) & (!sk[42]) & (g1424) & (!g1432) & (g1430) & (g1435)) + ((g1423) & (!sk[42]) & (g1424) & (g1432) & (!g1430) & (!g1435)) + ((g1423) & (!sk[42]) & (g1424) & (g1432) & (!g1430) & (g1435)) + ((g1423) & (!sk[42]) & (g1424) & (g1432) & (g1430) & (!g1435)) + ((g1423) & (!sk[42]) & (g1424) & (g1432) & (g1430) & (g1435)));
	assign g1441 = (((!g1068) & (!sk[43]) & (g1439) & (!g1440)) + ((!g1068) & (!sk[43]) & (g1439) & (g1440)) + ((!g1068) & (sk[43]) & (g1439) & (!g1440)) + ((!g1068) & (sk[43]) & (g1439) & (g1440)) + ((g1068) & (!sk[43]) & (g1439) & (!g1440)) + ((g1068) & (!sk[43]) & (g1439) & (g1440)) + ((g1068) & (sk[43]) & (!g1439) & (!g1440)) + ((g1068) & (sk[43]) & (g1439) & (g1440)));
	assign g1442 = (((!sk[44]) & (!ax22x) & (!ax21x) & (!g6) & (ax20x)) + ((!sk[44]) & (!ax22x) & (!ax21x) & (g6) & (ax20x)) + ((!sk[44]) & (!ax22x) & (ax21x) & (!g6) & (ax20x)) + ((!sk[44]) & (!ax22x) & (ax21x) & (g6) & (ax20x)) + ((!sk[44]) & (ax22x) & (!ax21x) & (!g6) & (!ax20x)) + ((!sk[44]) & (ax22x) & (!ax21x) & (!g6) & (ax20x)) + ((!sk[44]) & (ax22x) & (!ax21x) & (g6) & (!ax20x)) + ((!sk[44]) & (ax22x) & (!ax21x) & (g6) & (ax20x)) + ((!sk[44]) & (ax22x) & (ax21x) & (!g6) & (!ax20x)) + ((!sk[44]) & (ax22x) & (ax21x) & (!g6) & (ax20x)) + ((!sk[44]) & (ax22x) & (ax21x) & (g6) & (!ax20x)) + ((!sk[44]) & (ax22x) & (ax21x) & (g6) & (ax20x)) + ((sk[44]) & (!ax22x) & (!ax21x) & (g6) & (!ax20x)));
	assign g1443 = (((!g1432) & (!sk[45]) & (!g1437) & (!g1434) & (g1438)) + ((!g1432) & (!sk[45]) & (!g1437) & (g1434) & (g1438)) + ((!g1432) & (!sk[45]) & (g1437) & (!g1434) & (g1438)) + ((!g1432) & (!sk[45]) & (g1437) & (g1434) & (g1438)) + ((!g1432) & (sk[45]) & (g1437) & (!g1434) & (!g1438)) + ((g1432) & (!sk[45]) & (!g1437) & (!g1434) & (!g1438)) + ((g1432) & (!sk[45]) & (!g1437) & (!g1434) & (g1438)) + ((g1432) & (!sk[45]) & (!g1437) & (g1434) & (!g1438)) + ((g1432) & (!sk[45]) & (!g1437) & (g1434) & (g1438)) + ((g1432) & (!sk[45]) & (g1437) & (!g1434) & (!g1438)) + ((g1432) & (!sk[45]) & (g1437) & (!g1434) & (g1438)) + ((g1432) & (!sk[45]) & (g1437) & (g1434) & (!g1438)) + ((g1432) & (!sk[45]) & (g1437) & (g1434) & (g1438)) + ((g1432) & (sk[45]) & (!g1437) & (!g1434) & (!g1438)) + ((g1432) & (sk[45]) & (g1437) & (!g1434) & (!g1438)) + ((g1432) & (sk[45]) & (g1437) & (g1434) & (!g1438)));
	assign sinx23x = (((!g1068) & (!g1439) & (!g1440) & (!sk[46]) & (g1442) & (!g1443)) + ((!g1068) & (!g1439) & (!g1440) & (!sk[46]) & (g1442) & (g1443)) + ((!g1068) & (!g1439) & (!g1440) & (sk[46]) & (!g1442) & (g1443)) + ((!g1068) & (!g1439) & (!g1440) & (sk[46]) & (g1442) & (!g1443)) + ((!g1068) & (!g1439) & (!g1440) & (sk[46]) & (g1442) & (g1443)) + ((!g1068) & (!g1439) & (g1440) & (!sk[46]) & (!g1442) & (!g1443)) + ((!g1068) & (!g1439) & (g1440) & (!sk[46]) & (!g1442) & (g1443)) + ((!g1068) & (!g1439) & (g1440) & (!sk[46]) & (g1442) & (!g1443)) + ((!g1068) & (!g1439) & (g1440) & (!sk[46]) & (g1442) & (g1443)) + ((!g1068) & (!g1439) & (g1440) & (sk[46]) & (!g1442) & (g1443)) + ((!g1068) & (!g1439) & (g1440) & (sk[46]) & (g1442) & (!g1443)) + ((!g1068) & (!g1439) & (g1440) & (sk[46]) & (g1442) & (g1443)) + ((!g1068) & (g1439) & (!g1440) & (!sk[46]) & (!g1442) & (!g1443)) + ((!g1068) & (g1439) & (!g1440) & (!sk[46]) & (!g1442) & (g1443)) + ((!g1068) & (g1439) & (!g1440) & (!sk[46]) & (g1442) & (!g1443)) + ((!g1068) & (g1439) & (!g1440) & (!sk[46]) & (g1442) & (g1443)) + ((!g1068) & (g1439) & (!g1440) & (sk[46]) & (!g1442) & (g1443)) + ((!g1068) & (g1439) & (!g1440) & (sk[46]) & (g1442) & (!g1443)) + ((!g1068) & (g1439) & (!g1440) & (sk[46]) & (g1442) & (g1443)) + ((!g1068) & (g1439) & (g1440) & (!sk[46]) & (!g1442) & (!g1443)) + ((!g1068) & (g1439) & (g1440) & (!sk[46]) & (!g1442) & (g1443)) + ((!g1068) & (g1439) & (g1440) & (!sk[46]) & (g1442) & (!g1443)) + ((!g1068) & (g1439) & (g1440) & (!sk[46]) & (g1442) & (g1443)) + ((!g1068) & (g1439) & (g1440) & (sk[46]) & (!g1442) & (g1443)) + ((!g1068) & (g1439) & (g1440) & (sk[46]) & (g1442) & (!g1443)) + ((!g1068) & (g1439) & (g1440) & (sk[46]) & (g1442) & (g1443)) + ((g1068) & (!g1439) & (!g1440) & (!sk[46]) & (g1442) & (!g1443)) + ((g1068) & (!g1439) & (!g1440) & (!sk[46]) & (g1442) & (g1443)) + ((g1068) & (!g1439) & (!g1440) & (sk[46]) & (!g1442) & (!g1443)) + ((g1068) & (!g1439) & (!g1440) & (sk[46]) & (g1442) & (!g1443)) + ((g1068) & (!g1439) & (!g1440) & (sk[46]) & (g1442) & (g1443)) + ((g1068) & (!g1439) & (g1440) & (!sk[46]) & (!g1442) & (!g1443)) + ((g1068) & (!g1439) & (g1440) & (!sk[46]) & (!g1442) & (g1443)) + ((g1068) & (!g1439) & (g1440) & (!sk[46]) & (g1442) & (!g1443)) + ((g1068) & (!g1439) & (g1440) & (!sk[46]) & (g1442) & (g1443)) + ((g1068) & (!g1439) & (g1440) & (sk[46]) & (!g1442) & (!g1443)) + ((g1068) & (!g1439) & (g1440) & (sk[46]) & (g1442) & (!g1443)) + ((g1068) & (!g1439) & (g1440) & (sk[46]) & (g1442) & (g1443)) + ((g1068) & (g1439) & (!g1440) & (!sk[46]) & (!g1442) & (!g1443)) + ((g1068) & (g1439) & (!g1440) & (!sk[46]) & (!g1442) & (g1443)) + ((g1068) & (g1439) & (!g1440) & (!sk[46]) & (g1442) & (!g1443)) + ((g1068) & (g1439) & (!g1440) & (!sk[46]) & (g1442) & (g1443)) + ((g1068) & (g1439) & (!g1440) & (sk[46]) & (!g1442) & (!g1443)) + ((g1068) & (g1439) & (!g1440) & (sk[46]) & (g1442) & (!g1443)) + ((g1068) & (g1439) & (!g1440) & (sk[46]) & (g1442) & (g1443)) + ((g1068) & (g1439) & (g1440) & (!sk[46]) & (!g1442) & (!g1443)) + ((g1068) & (g1439) & (g1440) & (!sk[46]) & (!g1442) & (g1443)) + ((g1068) & (g1439) & (g1440) & (!sk[46]) & (g1442) & (!g1443)) + ((g1068) & (g1439) & (g1440) & (!sk[46]) & (g1442) & (g1443)) + ((g1068) & (g1439) & (g1440) & (sk[46]) & (!g1442) & (g1443)) + ((g1068) & (g1439) & (g1440) & (sk[46]) & (g1442) & (!g1443)) + ((g1068) & (g1439) & (g1440) & (sk[46]) & (g1442) & (g1443)));
	assign g1445 = (((!g1432) & (!g1437) & (!g1434) & (!sk[47]) & (g1438) & (!g1442)) + ((!g1432) & (!g1437) & (!g1434) & (!sk[47]) & (g1438) & (g1442)) + ((!g1432) & (!g1437) & (!g1434) & (sk[47]) & (!g1438) & (!g1442)) + ((!g1432) & (!g1437) & (!g1434) & (sk[47]) & (g1438) & (!g1442)) + ((!g1432) & (!g1437) & (g1434) & (!sk[47]) & (!g1438) & (!g1442)) + ((!g1432) & (!g1437) & (g1434) & (!sk[47]) & (!g1438) & (g1442)) + ((!g1432) & (!g1437) & (g1434) & (!sk[47]) & (g1438) & (!g1442)) + ((!g1432) & (!g1437) & (g1434) & (!sk[47]) & (g1438) & (g1442)) + ((!g1432) & (!g1437) & (g1434) & (sk[47]) & (!g1438) & (!g1442)) + ((!g1432) & (!g1437) & (g1434) & (sk[47]) & (g1438) & (!g1442)) + ((!g1432) & (g1437) & (!g1434) & (!sk[47]) & (!g1438) & (!g1442)) + ((!g1432) & (g1437) & (!g1434) & (!sk[47]) & (!g1438) & (g1442)) + ((!g1432) & (g1437) & (!g1434) & (!sk[47]) & (g1438) & (!g1442)) + ((!g1432) & (g1437) & (!g1434) & (!sk[47]) & (g1438) & (g1442)) + ((!g1432) & (g1437) & (!g1434) & (sk[47]) & (g1438) & (!g1442)) + ((!g1432) & (g1437) & (g1434) & (!sk[47]) & (!g1438) & (!g1442)) + ((!g1432) & (g1437) & (g1434) & (!sk[47]) & (!g1438) & (g1442)) + ((!g1432) & (g1437) & (g1434) & (!sk[47]) & (g1438) & (!g1442)) + ((!g1432) & (g1437) & (g1434) & (!sk[47]) & (g1438) & (g1442)) + ((!g1432) & (g1437) & (g1434) & (sk[47]) & (!g1438) & (!g1442)) + ((!g1432) & (g1437) & (g1434) & (sk[47]) & (g1438) & (!g1442)) + ((g1432) & (!g1437) & (!g1434) & (!sk[47]) & (g1438) & (!g1442)) + ((g1432) & (!g1437) & (!g1434) & (!sk[47]) & (g1438) & (g1442)) + ((g1432) & (!g1437) & (!g1434) & (sk[47]) & (g1438) & (!g1442)) + ((g1432) & (!g1437) & (g1434) & (!sk[47]) & (!g1438) & (!g1442)) + ((g1432) & (!g1437) & (g1434) & (!sk[47]) & (!g1438) & (g1442)) + ((g1432) & (!g1437) & (g1434) & (!sk[47]) & (g1438) & (!g1442)) + ((g1432) & (!g1437) & (g1434) & (!sk[47]) & (g1438) & (g1442)) + ((g1432) & (!g1437) & (g1434) & (sk[47]) & (!g1438) & (!g1442)) + ((g1432) & (!g1437) & (g1434) & (sk[47]) & (g1438) & (!g1442)) + ((g1432) & (g1437) & (!g1434) & (!sk[47]) & (!g1438) & (!g1442)) + ((g1432) & (g1437) & (!g1434) & (!sk[47]) & (!g1438) & (g1442)) + ((g1432) & (g1437) & (!g1434) & (!sk[47]) & (g1438) & (!g1442)) + ((g1432) & (g1437) & (!g1434) & (!sk[47]) & (g1438) & (g1442)) + ((g1432) & (g1437) & (!g1434) & (sk[47]) & (g1438) & (!g1442)) + ((g1432) & (g1437) & (g1434) & (!sk[47]) & (!g1438) & (!g1442)) + ((g1432) & (g1437) & (g1434) & (!sk[47]) & (!g1438) & (g1442)) + ((g1432) & (g1437) & (g1434) & (!sk[47]) & (g1438) & (!g1442)) + ((g1432) & (g1437) & (g1434) & (!sk[47]) & (g1438) & (g1442)) + ((g1432) & (g1437) & (g1434) & (sk[47]) & (g1438) & (!g1442)));
	assign sinx24x = (((!g1068) & (!sk[48]) & (!g1439) & (!g1440) & (g1445)) + ((!g1068) & (!sk[48]) & (!g1439) & (g1440) & (g1445)) + ((!g1068) & (!sk[48]) & (g1439) & (!g1440) & (g1445)) + ((!g1068) & (!sk[48]) & (g1439) & (g1440) & (g1445)) + ((g1068) & (!sk[48]) & (!g1439) & (!g1440) & (!g1445)) + ((g1068) & (!sk[48]) & (!g1439) & (!g1440) & (g1445)) + ((g1068) & (!sk[48]) & (!g1439) & (g1440) & (!g1445)) + ((g1068) & (!sk[48]) & (!g1439) & (g1440) & (g1445)) + ((g1068) & (!sk[48]) & (g1439) & (!g1440) & (!g1445)) + ((g1068) & (!sk[48]) & (g1439) & (!g1440) & (g1445)) + ((g1068) & (!sk[48]) & (g1439) & (g1440) & (!g1445)) + ((g1068) & (!sk[48]) & (g1439) & (g1440) & (g1445)) + ((g1068) & (sk[48]) & (!g1439) & (!g1440) & (!g1445)) + ((g1068) & (sk[48]) & (!g1439) & (!g1440) & (g1445)) + ((g1068) & (sk[48]) & (!g1439) & (g1440) & (!g1445)) + ((g1068) & (sk[48]) & (!g1439) & (g1440) & (g1445)) + ((g1068) & (sk[48]) & (g1439) & (!g1440) & (!g1445)) + ((g1068) & (sk[48]) & (g1439) & (!g1440) & (g1445)) + ((g1068) & (sk[48]) & (g1439) & (g1440) & (!g1445)));
	assign g1447 = (((!sk[49]) & (g1448) & (g1449)) + ((sk[49]) & (!g1448) & (!g1449)));
	assign g1448 = (((!g722) & (sk[50]) & (g1450)) + ((g722) & (!sk[50]) & (g1450)));
	assign g1449 = (((!sk[51]) & (g722) & (g1453)) + ((sk[51]) & (g722) & (g1453)));
	assign g1450 = (((!g1451) & (sk[52]) & (!g1452)) + ((g1451) & (!sk[52]) & (g1452)));
	assign g1451 = (((!g844) & (sk[53]) & (g1456)) + ((g844) & (!sk[53]) & (g1456)));
	assign g1452 = (((g844) & (!sk[54]) & (g1457)) + ((g844) & (sk[54]) & (g1457)));
	assign g1453 = (((!g1454) & (sk[55]) & (!g1455)) + ((g1454) & (!sk[55]) & (g1455)));
	assign g1454 = (((!sk[56]) & (g844) & (g1458)) + ((sk[56]) & (!g844) & (g1458)));
	assign g1455 = (((!sk[57]) & (g844) & (g1459)) + ((sk[57]) & (g844) & (g1459)));
	assign g1456 = (((!sk[58]) & (!g842) & (!g777) & (!g724) & (g754)) + ((!sk[58]) & (!g842) & (!g777) & (g724) & (g754)) + ((!sk[58]) & (!g842) & (g777) & (!g724) & (g754)) + ((!sk[58]) & (!g842) & (g777) & (g724) & (g754)) + ((!sk[58]) & (g842) & (!g777) & (!g724) & (!g754)) + ((!sk[58]) & (g842) & (!g777) & (!g724) & (g754)) + ((!sk[58]) & (g842) & (!g777) & (g724) & (!g754)) + ((!sk[58]) & (g842) & (!g777) & (g724) & (g754)) + ((!sk[58]) & (g842) & (g777) & (!g724) & (!g754)) + ((!sk[58]) & (g842) & (g777) & (!g724) & (g754)) + ((!sk[58]) & (g842) & (g777) & (g724) & (!g754)) + ((!sk[58]) & (g842) & (g777) & (g724) & (g754)) + ((sk[58]) & (!g842) & (g777) & (!g724) & (!g754)) + ((sk[58]) & (!g842) & (g777) & (!g724) & (g754)) + ((sk[58]) & (!g842) & (g777) & (g724) & (!g754)) + ((sk[58]) & (!g842) & (g777) & (g724) & (g754)) + ((sk[58]) & (g842) & (!g777) & (!g724) & (!g754)) + ((sk[58]) & (g842) & (!g777) & (!g724) & (g754)) + ((sk[58]) & (g842) & (g777) & (!g724) & (g754)) + ((sk[58]) & (g842) & (g777) & (g724) & (g754)));
	assign g1457 = (((!g842) & (!g777) & (!g723) & (!sk[59]) & (g754)) + ((!g842) & (!g777) & (!g723) & (sk[59]) & (!g754)) + ((!g842) & (!g777) & (!g723) & (sk[59]) & (g754)) + ((!g842) & (!g777) & (g723) & (!sk[59]) & (g754)) + ((!g842) & (g777) & (!g723) & (!sk[59]) & (g754)) + ((!g842) & (g777) & (!g723) & (sk[59]) & (!g754)) + ((!g842) & (g777) & (!g723) & (sk[59]) & (g754)) + ((!g842) & (g777) & (g723) & (!sk[59]) & (g754)) + ((!g842) & (g777) & (g723) & (sk[59]) & (!g754)) + ((!g842) & (g777) & (g723) & (sk[59]) & (g754)) + ((g842) & (!g777) & (!g723) & (!sk[59]) & (!g754)) + ((g842) & (!g777) & (!g723) & (!sk[59]) & (g754)) + ((g842) & (!g777) & (!g723) & (sk[59]) & (!g754)) + ((g842) & (!g777) & (!g723) & (sk[59]) & (g754)) + ((g842) & (!g777) & (g723) & (!sk[59]) & (!g754)) + ((g842) & (!g777) & (g723) & (!sk[59]) & (g754)) + ((g842) & (g777) & (!g723) & (!sk[59]) & (!g754)) + ((g842) & (g777) & (!g723) & (!sk[59]) & (g754)) + ((g842) & (g777) & (!g723) & (sk[59]) & (g754)) + ((g842) & (g777) & (g723) & (!sk[59]) & (!g754)) + ((g842) & (g777) & (g723) & (!sk[59]) & (g754)) + ((g842) & (g777) & (g723) & (sk[59]) & (g754)));
	assign g1458 = (((!sk[60]) & (!g842) & (!g777) & (!g724) & (g754)) + ((!sk[60]) & (!g842) & (!g777) & (g724) & (g754)) + ((!sk[60]) & (!g842) & (g777) & (!g724) & (g754)) + ((!sk[60]) & (!g842) & (g777) & (g724) & (g754)) + ((!sk[60]) & (g842) & (!g777) & (!g724) & (!g754)) + ((!sk[60]) & (g842) & (!g777) & (!g724) & (g754)) + ((!sk[60]) & (g842) & (!g777) & (g724) & (!g754)) + ((!sk[60]) & (g842) & (!g777) & (g724) & (g754)) + ((!sk[60]) & (g842) & (g777) & (!g724) & (!g754)) + ((!sk[60]) & (g842) & (g777) & (!g724) & (g754)) + ((!sk[60]) & (g842) & (g777) & (g724) & (!g754)) + ((!sk[60]) & (g842) & (g777) & (g724) & (g754)) + ((sk[60]) & (g842) & (!g777) & (!g724) & (!g754)) + ((sk[60]) & (g842) & (!g777) & (!g724) & (g754)) + ((sk[60]) & (g842) & (g777) & (!g724) & (g754)) + ((sk[60]) & (g842) & (g777) & (g724) & (g754)));
	assign g1459 = (((!g842) & (!sk[61]) & (!g777) & (!g723) & (g754)) + ((!g842) & (!sk[61]) & (!g777) & (g723) & (g754)) + ((!g842) & (!sk[61]) & (g777) & (!g723) & (g754)) + ((!g842) & (!sk[61]) & (g777) & (g723) & (g754)) + ((!g842) & (sk[61]) & (!g777) & (!g723) & (!g754)) + ((!g842) & (sk[61]) & (!g777) & (!g723) & (g754)) + ((g842) & (!sk[61]) & (!g777) & (!g723) & (!g754)) + ((g842) & (!sk[61]) & (!g777) & (!g723) & (g754)) + ((g842) & (!sk[61]) & (!g777) & (g723) & (!g754)) + ((g842) & (!sk[61]) & (!g777) & (g723) & (g754)) + ((g842) & (!sk[61]) & (g777) & (!g723) & (!g754)) + ((g842) & (!sk[61]) & (g777) & (!g723) & (g754)) + ((g842) & (!sk[61]) & (g777) & (g723) & (!g754)) + ((g842) & (!sk[61]) & (g777) & (g723) & (g754)) + ((g842) & (sk[61]) & (!g777) & (!g723) & (!g754)) + ((g842) & (sk[61]) & (!g777) & (!g723) & (g754)) + ((g842) & (sk[61]) & (g777) & (!g723) & (g754)) + ((g842) & (sk[61]) & (g777) & (g723) & (g754)));

endmodule